
module round ( in, round_num, keyin, keyout, out );
  input [127:0] in;
  input [3:0] round_num;
  input [127:0] keyin;
  output [127:0] keyout;
  output [127:0] out;
  wire   n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, \_0_net_[127] ,
         \_0_net_[126] , \_0_net_[125] , \_0_net_[124] , \_0_net_[123] ,
         \_0_net_[122] , \_0_net_[121] , \_0_net_[120] , \_0_net_[119] ,
         \_0_net_[118] , \_0_net_[117] , \_0_net_[116] , \_0_net_[115] ,
         \_0_net_[114] , \_0_net_[113] , \_0_net_[112] , \_0_net_[111] ,
         \_0_net_[110] , \_0_net_[109] , \_0_net_[108] , \_0_net_[107] ,
         \_0_net_[106] , \_0_net_[105] , \_0_net_[104] , \_0_net_[103] ,
         \_0_net_[102] , \_0_net_[101] , \_0_net_[100] , \_0_net_[99] ,
         \_0_net_[98] , \_0_net_[97] , \_0_net_[96] , \_0_net_[95] ,
         \_0_net_[94] , \_0_net_[93] , \_0_net_[92] , \_0_net_[91] ,
         \_0_net_[90] , \_0_net_[89] , \_0_net_[88] , \_0_net_[87] ,
         \_0_net_[86] , \_0_net_[85] , \_0_net_[84] , \_0_net_[83] ,
         \_0_net_[82] , \_0_net_[81] , \_0_net_[80] , \_0_net_[79] ,
         \_0_net_[78] , \_0_net_[77] , \_0_net_[76] , \_0_net_[75] ,
         \_0_net_[74] , \_0_net_[73] , \_0_net_[72] , \_0_net_[71] ,
         \_0_net_[70] , \_0_net_[69] , \_0_net_[68] , \_0_net_[67] ,
         \_0_net_[66] , \_0_net_[65] , \_0_net_[64] , \_0_net_[63] ,
         \_0_net_[62] , \_0_net_[61] , \_0_net_[60] , \_0_net_[59] ,
         \_0_net_[58] , \_0_net_[57] , \_0_net_[56] , \_0_net_[55] ,
         \_0_net_[54] , \_0_net_[53] , \_0_net_[52] , \_0_net_[51] ,
         \_0_net_[50] , \_0_net_[49] , \_0_net_[48] , \_0_net_[47] ,
         \_0_net_[46] , \_0_net_[45] , \_0_net_[44] , \_0_net_[43] ,
         \_0_net_[42] , \_0_net_[41] , \_0_net_[40] , \_0_net_[39] ,
         \_0_net_[38] , \_0_net_[37] , \_0_net_[36] , \_0_net_[35] ,
         \_0_net_[34] , \_0_net_[33] , \_0_net_[32] , \_0_net_[31] ,
         \_0_net_[30] , \_0_net_[29] , \_0_net_[28] , \_0_net_[27] ,
         \_0_net_[26] , \_0_net_[25] , \_0_net_[24] , \_0_net_[23] ,
         \_0_net_[22] , \_0_net_[21] , \_0_net_[20] , \_0_net_[19] ,
         \_0_net_[18] , \_0_net_[17] , \_0_net_[16] , \_0_net_[15] ,
         \_0_net_[14] , \_0_net_[13] , \_0_net_[12] , \_0_net_[11] ,
         \_0_net_[10] , \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] ,
         \_0_net_[5] , \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] ,
         \_0_net_[0] , n3, n2, n4, n13, n14, n15, n16, n17, n19, n21, n23, n24,
         n25, n27, n29, n31, n32, n34, n35, n36, n38, n40, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n157, n158, n159,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n190, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n206, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n221, n222, n223, n224, n225, n226, n227, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n348, n349, n350, n351, n352, n354, n356, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n380, n381, n382, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n394, n396, n397,
         n399, n400, n402, n404, n405, n407, n408, n410, n412, n413, n414,
         n416, n417, n419, n421, n422, n423, n424, n426, n427, n428, n429,
         n430, n431, n432, n433;
  wire   [127:0] sb_out;
  wire   [127:0] sr_out;
  wire   [127:0] mc_out;

  keygen x ( .round_num({round_num[3:2], n74, n72}), .keyin(keyin), .keyout({
        keyout[127:126], n434, n435, keyout[123:96], n436, n437, n438, n439, 
        n440, keyout[90:88], n441, n442, n443, keyout[84:82], n444, n445, 
        keyout[79], n446, n447, keyout[76:75], n448, keyout[73:72], n449, n450, 
        keyout[69], n451, n452, keyout[66], n453, keyout[64:60], n454, 
        keyout[58:56], n455, n456, n457, keyout[52], n458, n459, keyout[49], 
        n460, keyout[47], n461, n462, keyout[44], n463, keyout[42], n464, n465, 
        keyout[39], n466, n467, n468, n469, n470, n471, n472, keyout[31], n473, 
        n474, keyout[28], n475, keyout[26], n476, n477, keyout[23:17], n478, 
        keyout[15], n479, n480, keyout[12:8], n481, n482, keyout[5], n483, 
        keyout[3:2], n484, keyout[0]}) );
  subbytes sb ( .in(in), .out(sb_out) );
  shift_rows sr ( .in(sb_out), .out(sr_out) );
  Mix_Column mc ( .in(sr_out), .out(mc_out) );
  add_round_keys_1 adk ( .state({\_0_net_[127] , \_0_net_[126] , 
        \_0_net_[125] , \_0_net_[124] , \_0_net_[123] , \_0_net_[122] , 
        \_0_net_[121] , \_0_net_[120] , \_0_net_[119] , \_0_net_[118] , 
        \_0_net_[117] , \_0_net_[116] , \_0_net_[115] , \_0_net_[114] , 
        \_0_net_[113] , \_0_net_[112] , \_0_net_[111] , \_0_net_[110] , 
        \_0_net_[109] , \_0_net_[108] , \_0_net_[107] , \_0_net_[106] , 
        \_0_net_[105] , \_0_net_[104] , \_0_net_[103] , \_0_net_[102] , 
        \_0_net_[101] , \_0_net_[100] , \_0_net_[99] , \_0_net_[98] , 
        \_0_net_[97] , \_0_net_[96] , \_0_net_[95] , \_0_net_[94] , 
        \_0_net_[93] , \_0_net_[92] , \_0_net_[91] , \_0_net_[90] , 
        \_0_net_[89] , \_0_net_[88] , \_0_net_[87] , \_0_net_[86] , 
        \_0_net_[85] , \_0_net_[84] , \_0_net_[83] , \_0_net_[82] , 
        \_0_net_[81] , \_0_net_[80] , \_0_net_[79] , \_0_net_[78] , 
        \_0_net_[77] , \_0_net_[76] , \_0_net_[75] , \_0_net_[74] , 
        \_0_net_[73] , \_0_net_[72] , \_0_net_[71] , \_0_net_[70] , 
        \_0_net_[69] , \_0_net_[68] , \_0_net_[67] , \_0_net_[66] , 
        \_0_net_[65] , \_0_net_[64] , \_0_net_[63] , \_0_net_[62] , 
        \_0_net_[61] , \_0_net_[60] , \_0_net_[59] , \_0_net_[58] , 
        \_0_net_[57] , \_0_net_[56] , \_0_net_[55] , \_0_net_[54] , 
        \_0_net_[53] , \_0_net_[52] , \_0_net_[51] , \_0_net_[50] , 
        \_0_net_[49] , \_0_net_[48] , \_0_net_[47] , \_0_net_[46] , 
        \_0_net_[45] , \_0_net_[44] , \_0_net_[43] , \_0_net_[42] , 
        \_0_net_[41] , \_0_net_[40] , \_0_net_[39] , \_0_net_[38] , 
        \_0_net_[37] , \_0_net_[36] , \_0_net_[35] , \_0_net_[34] , 
        \_0_net_[33] , \_0_net_[32] , \_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_0_net_[0] }), 
        .subkey({keyout[127:126], n434, n435, keyout[123:96], n436, n437, n438, 
        n439, n440, keyout[90:88], n441, n442, n443, keyout[84:82], n444, n445, 
        keyout[79], n446, n447, keyout[76:75], n448, keyout[73:72], n449, n450, 
        keyout[69], n451, n452, keyout[66], n453, keyout[64:60], n454, 
        keyout[58:56], n455, n456, n457, keyout[52], n458, n459, keyout[49], 
        n460, keyout[47], n461, n462, keyout[44], n463, keyout[42], n464, n465, 
        keyout[39], n466, n467, n468, n469, n470, n471, n472, keyout[31], n473, 
        n474, keyout[28], n475, keyout[26], n476, n477, keyout[23:17], n478, 
        keyout[15], n479, n480, keyout[12:8], n481, n482, keyout[5], n483, 
        keyout[3:2], n484, keyout[0]}), .out(out) );
  AO22X1_HVT U126 ( .A1(mc_out[102]), .A2(n113), .A3(sr_out[102]), .A4(n87), 
        .Y(\_0_net_[102] ) );
  NAND2X0_HVT U131 ( .A1(round_num[3]), .A2(round_num[1]), .Y(n3) );
  DELLN1X2_HVT U1 ( .A(sr_out[25]), .Y(n31) );
  DELLN1X2_HVT U2 ( .A(sr_out[72]), .Y(n289) );
  DELLN1X2_HVT U3 ( .A(sr_out[73]), .Y(n286) );
  DELLN1X2_HVT U4 ( .A(sr_out[127]), .Y(n336) );
  DELLN1X2_HVT U5 ( .A(sr_out[1]), .Y(n259) );
  DELLN1X2_HVT U6 ( .A(sr_out[5]), .Y(n272) );
  DELLN1X2_HVT U7 ( .A(sr_out[15]), .Y(n421) );
  NBUFFX2_HVT U8 ( .A(sr_out[16]), .Y(n416) );
  DELLN1X2_HVT U9 ( .A(sr_out[19]), .Y(n404) );
  DELLN1X2_HVT U10 ( .A(sr_out[28]), .Y(n130) );
  DELLN1X2_HVT U11 ( .A(sr_out[34]), .Y(n345) );
  DELLN1X2_HVT U12 ( .A(sr_out[39]), .Y(n384) );
  DELLN1X2_HVT U13 ( .A(sr_out[41]), .Y(n407) );
  NBUFFX2_HVT U14 ( .A(sr_out[55]), .Y(n319) );
  DELLN1X2_HVT U15 ( .A(sr_out[57]), .Y(n13) );
  DELLN1X2_HVT U16 ( .A(sr_out[71]), .Y(n331) );
  DELLN1X2_HVT U17 ( .A(sr_out[79]), .Y(n279) );
  NBUFFX2_HVT U18 ( .A(sr_out[81]), .Y(n396) );
  DELLN1X2_HVT U19 ( .A(sr_out[86]), .Y(n24) );
  DELLN1X2_HVT U20 ( .A(sr_out[97]), .Y(n179) );
  NBUFFX2_HVT U21 ( .A(sr_out[100]), .Y(n71) );
  DELLN1X2_HVT U22 ( .A(sr_out[108]), .Y(n42) );
  DELLN1X2_HVT U23 ( .A(sr_out[114]), .Y(n216) );
  INVX1_HVT U24 ( .A(n447), .Y(n410) );
  INVX1_HVT U25 ( .A(n459), .Y(n334) );
  INVX1_HVT U26 ( .A(n469), .Y(n159) );
  INVX1_HVT U27 ( .A(n470), .Y(n227) );
  INVX1_HVT U28 ( .A(n443), .Y(n38) );
  INVX1_HVT U29 ( .A(n434), .Y(n36) );
  INVX1_HVT U30 ( .A(n458), .Y(n69) );
  INVX1_HVT U31 ( .A(n438), .Y(n51) );
  INVX1_HVT U32 ( .A(n451), .Y(n29) );
  INVX1_HVT U33 ( .A(n449), .Y(n402) );
  INVX1_HVT U34 ( .A(n463), .Y(n354) );
  INVX1_HVT U35 ( .A(n474), .Y(n419) );
  INVX1_HVT U36 ( .A(n475), .Y(n17) );
  NBUFFX2_HVT U37 ( .A(n483), .Y(keyout[4]) );
  NAND2X0_HVT U38 ( .A1(mc_out[111]), .A2(n104), .Y(n2) );
  NAND2X0_HVT U39 ( .A1(sr_out[111]), .A2(n431), .Y(n4) );
  NAND2X0_HVT U40 ( .A1(n2), .A2(n4), .Y(\_0_net_[111] ) );
  DELLN1X2_HVT U41 ( .A(sr_out[119]), .Y(n306) );
  INVX1_HVT U42 ( .A(n436), .Y(n414) );
  NBUFFX2_HVT U43 ( .A(n460), .Y(keyout[48]) );
  DELLN1X2_HVT U44 ( .A(sr_out[4]), .Y(n399) );
  NBUFFX2_HVT U45 ( .A(n481), .Y(keyout[7]) );
  NBUFFX2_HVT U46 ( .A(n440), .Y(keyout[91]) );
  NBUFFX2_HVT U47 ( .A(n435), .Y(keyout[124]) );
  NBUFFX2_HVT U48 ( .A(n473), .Y(keyout[30]) );
  NBUFFX2_HVT U49 ( .A(n439), .Y(keyout[92]) );
  NBUFFX2_HVT U50 ( .A(n476), .Y(keyout[25]) );
  NBUFFX2_HVT U51 ( .A(n466), .Y(keyout[38]) );
  INVX1_HVT U52 ( .A(round_num[1]), .Y(n73) );
  INVX0_HVT U53 ( .A(n446), .Y(n366) );
  INVX1_HVT U54 ( .A(n456), .Y(n394) );
  INVX1_HVT U55 ( .A(n461), .Y(n155) );
  INVX1_HVT U56 ( .A(n465), .Y(n204) );
  INVX1_HVT U57 ( .A(n478), .Y(n346) );
  INVX1_HVT U58 ( .A(n479), .Y(n356) );
  INVX1_HVT U59 ( .A(n484), .Y(n253) );
  INVX1_HVT U60 ( .A(n14), .Y(n427) );
  NBUFFX2_HVT U61 ( .A(sr_out[20]), .Y(n79) );
  NBUFFX2_HVT U62 ( .A(sr_out[60]), .Y(n387) );
  INVX1_HVT U63 ( .A(n14), .Y(n112) );
  INVX1_HVT U64 ( .A(n427), .Y(n116) );
  DELLN1X2_HVT U65 ( .A(sr_out[103]), .Y(n23) );
  INVX1_HVT U66 ( .A(n111), .Y(n76) );
  INVX1_HVT U67 ( .A(n432), .Y(n120) );
  INVX1_HVT U68 ( .A(n427), .Y(n121) );
  INVX1_HVT U69 ( .A(n111), .Y(n122) );
  INVX1_HVT U70 ( .A(n112), .Y(n115) );
  INVX1_HVT U71 ( .A(n112), .Y(n119) );
  INVX1_HVT U72 ( .A(n427), .Y(n75) );
  INVX1_HVT U73 ( .A(n427), .Y(n114) );
  NAND2X0_HVT U74 ( .A1(sr_out[26]), .A2(n107), .Y(n201) );
  DELLN1X2_HVT U75 ( .A(sr_out[46]), .Y(n322) );
  NAND2X0_HVT U76 ( .A1(sr_out[67]), .A2(n107), .Y(n363) );
  NAND2X0_HVT U77 ( .A1(sr_out[74]), .A2(n83), .Y(n258) );
  NAND2X0_HVT U78 ( .A1(sr_out[104]), .A2(n106), .Y(n64) );
  INVX1_HVT U79 ( .A(n445), .Y(n32) );
  INVX1_HVT U80 ( .A(n452), .Y(n19) );
  INVX1_HVT U81 ( .A(n462), .Y(n27) );
  INVX1_HVT U82 ( .A(n454), .Y(n382) );
  INVX1_HVT U83 ( .A(n437), .Y(n417) );
  INVX1_HVT U84 ( .A(n441), .Y(n392) );
  INVX1_HVT U85 ( .A(n442), .Y(n188) );
  INVX1_HVT U86 ( .A(n444), .Y(n219) );
  INVX1_HVT U87 ( .A(n448), .Y(n190) );
  INVX1_HVT U88 ( .A(n450), .Y(n25) );
  INVX1_HVT U89 ( .A(n453), .Y(n405) );
  INVX1_HVT U90 ( .A(n455), .Y(n400) );
  INVX1_HVT U91 ( .A(n457), .Y(n397) );
  INVX1_HVT U92 ( .A(n464), .Y(n378) );
  INVX1_HVT U93 ( .A(n467), .Y(n408) );
  INVX1_HVT U94 ( .A(n468), .Y(n424) );
  INVX1_HVT U95 ( .A(n471), .Y(n21) );
  INVX1_HVT U96 ( .A(n472), .Y(n40) );
  INVX1_HVT U97 ( .A(n137), .Y(keyout[24]) );
  INVX1_HVT U98 ( .A(n477), .Y(n137) );
  INVX1_HVT U99 ( .A(n480), .Y(n206) );
  INVX1_HVT U100 ( .A(n352), .Y(keyout[6]) );
  INVX1_HVT U101 ( .A(n482), .Y(n352) );
  OR3X1_HVT U102 ( .A1(round_num[2]), .A2(round_num[0]), .A3(n3), .Y(n14) );
  INVX0_HVT U103 ( .A(n426), .Y(n433) );
  INVX0_HVT U104 ( .A(n82), .Y(n83) );
  INVX0_HVT U105 ( .A(n155), .Y(keyout[46]) );
  INVX1_HVT U106 ( .A(n206), .Y(keyout[13]) );
  INVX1_HVT U107 ( .A(n400), .Y(keyout[55]) );
  NAND2X0_HVT U108 ( .A1(mc_out[42]), .A2(n116), .Y(n15) );
  NAND2X0_HVT U109 ( .A1(sr_out[42]), .A2(n430), .Y(n16) );
  NAND2X0_HVT U110 ( .A1(n15), .A2(n16), .Y(\_0_net_[42] ) );
  INVX1_HVT U111 ( .A(n402), .Y(keyout[71]) );
  INVX0_HVT U112 ( .A(n17), .Y(keyout[27]) );
  INVX0_HVT U113 ( .A(n19), .Y(keyout[67]) );
  INVX0_HVT U114 ( .A(n21), .Y(keyout[33]) );
  INVX0_HVT U115 ( .A(n14), .Y(n111) );
  INVX0_HVT U116 ( .A(n25), .Y(keyout[70]) );
  NAND2X0_HVT U117 ( .A1(sr_out[36]), .A2(n106), .Y(n54) );
  INVX0_HVT U118 ( .A(n417), .Y(keyout[94]) );
  INVX0_HVT U119 ( .A(n27), .Y(keyout[45]) );
  INVX0_HVT U120 ( .A(n29), .Y(keyout[68]) );
  INVX0_HVT U121 ( .A(n32), .Y(keyout[80]) );
  NAND2X0_HVT U122 ( .A1(mc_out[86]), .A2(n115), .Y(n34) );
  NAND2X0_HVT U123 ( .A1(n24), .A2(n106), .Y(n35) );
  NAND2X0_HVT U124 ( .A1(n34), .A2(n35), .Y(\_0_net_[86] ) );
  INVX0_HVT U125 ( .A(n36), .Y(keyout[125]) );
  NAND2X0_HVT U127 ( .A1(sr_out[68]), .A2(n103), .Y(n56) );
  INVX0_HVT U128 ( .A(n38), .Y(keyout[85]) );
  NAND2X0_HVT U129 ( .A1(n13), .A2(n84), .Y(n321) );
  INVX0_HVT U130 ( .A(n40), .Y(keyout[32]) );
  INVX0_HVT U132 ( .A(n408), .Y(keyout[37]) );
  NAND2X0_HVT U133 ( .A1(mc_out[47]), .A2(n85), .Y(n43) );
  NAND2X0_HVT U134 ( .A1(sr_out[47]), .A2(n88), .Y(n44) );
  NAND2X0_HVT U135 ( .A1(n43), .A2(n44), .Y(\_0_net_[47] ) );
  NAND2X0_HVT U136 ( .A1(mc_out[82]), .A2(n119), .Y(n45) );
  NAND2X0_HVT U137 ( .A1(n429), .A2(sr_out[82]), .Y(n46) );
  NAND2X0_HVT U138 ( .A1(n45), .A2(n46), .Y(\_0_net_[82] ) );
  NAND2X0_HVT U139 ( .A1(mc_out[76]), .A2(n121), .Y(n47) );
  NAND2X0_HVT U140 ( .A1(sr_out[76]), .A2(n87), .Y(n48) );
  NAND2X0_HVT U141 ( .A1(n47), .A2(n48), .Y(\_0_net_[76] ) );
  NAND2X0_HVT U142 ( .A1(mc_out[38]), .A2(n116), .Y(n49) );
  NAND2X0_HVT U143 ( .A1(sr_out[38]), .A2(n97), .Y(n50) );
  NAND2X0_HVT U144 ( .A1(n49), .A2(n50), .Y(\_0_net_[38] ) );
  INVX0_HVT U145 ( .A(n51), .Y(keyout[93]) );
  NAND2X0_HVT U146 ( .A1(mc_out[36]), .A2(n89), .Y(n53) );
  NAND2X0_HVT U147 ( .A1(n53), .A2(n54), .Y(\_0_net_[36] ) );
  NAND2X0_HVT U148 ( .A1(mc_out[68]), .A2(n118), .Y(n55) );
  NAND2X0_HVT U149 ( .A1(n55), .A2(n56), .Y(\_0_net_[68] ) );
  NAND2X0_HVT U150 ( .A1(mc_out[122]), .A2(n115), .Y(n57) );
  NAND2X0_HVT U151 ( .A1(sr_out[122]), .A2(n83), .Y(n58) );
  NAND2X0_HVT U152 ( .A1(n57), .A2(n58), .Y(\_0_net_[122] ) );
  NAND2X0_HVT U153 ( .A1(mc_out[29]), .A2(n114), .Y(n59) );
  NAND2X0_HVT U154 ( .A1(sr_out[29]), .A2(n87), .Y(n60) );
  NAND2X0_HVT U155 ( .A1(n59), .A2(n60), .Y(\_0_net_[29] ) );
  INVX0_HVT U156 ( .A(n219), .Y(keyout[81]) );
  NAND2X0_HVT U157 ( .A1(mc_out[11]), .A2(n116), .Y(n61) );
  NAND2X0_HVT U158 ( .A1(sr_out[11]), .A2(n84), .Y(n62) );
  NAND2X0_HVT U159 ( .A1(n61), .A2(n62), .Y(\_0_net_[11] ) );
  NAND2X0_HVT U160 ( .A1(mc_out[104]), .A2(n89), .Y(n63) );
  NAND2X0_HVT U161 ( .A1(n63), .A2(n64), .Y(\_0_net_[104] ) );
  NAND2X0_HVT U162 ( .A1(mc_out[5]), .A2(n116), .Y(n65) );
  NAND2X0_HVT U163 ( .A1(n272), .A2(n91), .Y(n66) );
  NAND2X0_HVT U164 ( .A1(n65), .A2(n66), .Y(\_0_net_[5] ) );
  NAND2X0_HVT U165 ( .A1(mc_out[84]), .A2(n75), .Y(n67) );
  NAND2X0_HVT U166 ( .A1(sr_out[84]), .A2(n95), .Y(n68) );
  NAND2X0_HVT U167 ( .A1(n67), .A2(n68), .Y(\_0_net_[84] ) );
  NAND2X0_HVT U168 ( .A1(n431), .A2(sr_out[48]), .Y(n303) );
  INVX0_HVT U169 ( .A(n427), .Y(n82) );
  INVX0_HVT U170 ( .A(n69), .Y(keyout[51]) );
  INVX0_HVT U171 ( .A(n346), .Y(keyout[16]) );
  NBUFFX2_HVT U172 ( .A(round_num[0]), .Y(n72) );
  INVX0_HVT U173 ( .A(n111), .Y(n117) );
  INVX0_HVT U174 ( .A(n73), .Y(n74) );
  NAND2X0_HVT U175 ( .A1(mc_out[32]), .A2(n114), .Y(n77) );
  NAND2X0_HVT U176 ( .A1(n83), .A2(sr_out[32]), .Y(n78) );
  NAND2X0_HVT U177 ( .A1(n77), .A2(n78), .Y(\_0_net_[32] ) );
  INVX0_HVT U178 ( .A(n112), .Y(n113) );
  NAND2X0_HVT U179 ( .A1(mc_out[70]), .A2(n114), .Y(n80) );
  NAND2X0_HVT U180 ( .A1(sr_out[70]), .A2(n91), .Y(n81) );
  NAND2X0_HVT U181 ( .A1(n80), .A2(n81), .Y(\_0_net_[70] ) );
  INVX1_HVT U182 ( .A(n108), .Y(n84) );
  INVX0_HVT U183 ( .A(n111), .Y(n85) );
  INVX0_HVT U184 ( .A(n112), .Y(n86) );
  INVX1_HVT U185 ( .A(n85), .Y(n87) );
  INVX1_HVT U186 ( .A(n86), .Y(n88) );
  INVX0_HVT U187 ( .A(n431), .Y(n89) );
  INVX0_HVT U188 ( .A(n430), .Y(n90) );
  INVX1_HVT U189 ( .A(n90), .Y(n91) );
  INVX0_HVT U190 ( .A(n428), .Y(n92) );
  INVX0_HVT U191 ( .A(n428), .Y(n93) );
  INVX1_HVT U192 ( .A(n92), .Y(n94) );
  INVX1_HVT U193 ( .A(n93), .Y(n95) );
  INVX0_HVT U194 ( .A(n429), .Y(n96) );
  INVX1_HVT U195 ( .A(n96), .Y(n97) );
  INVX1_HVT U196 ( .A(n96), .Y(n98) );
  INVX0_HVT U197 ( .A(n433), .Y(n99) );
  INVX1_HVT U198 ( .A(n99), .Y(n100) );
  INVX0_HVT U199 ( .A(n111), .Y(n101) );
  INVX0_HVT U200 ( .A(n433), .Y(n102) );
  INVX1_HVT U201 ( .A(n101), .Y(n103) );
  INVX0_HVT U202 ( .A(n432), .Y(n104) );
  INVX0_HVT U203 ( .A(n432), .Y(n105) );
  INVX1_HVT U204 ( .A(n104), .Y(n106) );
  INVX1_HVT U205 ( .A(n105), .Y(n107) );
  INVX0_HVT U206 ( .A(n427), .Y(n108) );
  INVX0_HVT U207 ( .A(n432), .Y(n109) );
  INVX1_HVT U208 ( .A(n109), .Y(n110) );
  INVX0_HVT U209 ( .A(n111), .Y(n118) );
  INVX0_HVT U210 ( .A(n111), .Y(n426) );
  INVX0_HVT U211 ( .A(n82), .Y(n432) );
  INVX0_HVT U212 ( .A(n101), .Y(n429) );
  INVX0_HVT U213 ( .A(n426), .Y(n430) );
  INVX0_HVT U214 ( .A(n102), .Y(n431) );
  INVX0_HVT U215 ( .A(n104), .Y(n428) );
  NAND2X0_HVT U216 ( .A1(sr_out[2]), .A2(n431), .Y(n285) );
  NAND2X0_HVT U217 ( .A1(sr_out[75]), .A2(n110), .Y(n269) );
  NAND2X0_HVT U218 ( .A1(mc_out[14]), .A2(n115), .Y(n123) );
  NAND2X0_HVT U219 ( .A1(sr_out[14]), .A2(n433), .Y(n124) );
  NAND2X0_HVT U220 ( .A1(n123), .A2(n124), .Y(\_0_net_[14] ) );
  NAND2X0_HVT U221 ( .A1(mc_out[110]), .A2(n121), .Y(n125) );
  NAND2X0_HVT U222 ( .A1(sr_out[110]), .A2(n97), .Y(n126) );
  NAND2X0_HVT U223 ( .A1(n125), .A2(n126), .Y(\_0_net_[110] ) );
  DELLN2X2_HVT U224 ( .A(sr_out[7]), .Y(n127) );
  NAND2X0_HVT U225 ( .A1(mc_out[94]), .A2(n122), .Y(n128) );
  NAND2X0_HVT U226 ( .A1(sr_out[94]), .A2(n84), .Y(n129) );
  NAND2X0_HVT U227 ( .A1(n128), .A2(n129), .Y(\_0_net_[94] ) );
  NAND2X0_HVT U228 ( .A1(mc_out[18]), .A2(n116), .Y(n131) );
  NAND2X0_HVT U229 ( .A1(sr_out[18]), .A2(n100), .Y(n132) );
  NAND2X0_HVT U230 ( .A1(n131), .A2(n132), .Y(\_0_net_[18] ) );
  NAND2X0_HVT U231 ( .A1(n42), .A2(n95), .Y(n281) );
  NAND2X0_HVT U232 ( .A1(mc_out[16]), .A2(n102), .Y(n133) );
  NAND2X0_HVT U233 ( .A1(n416), .A2(n88), .Y(n134) );
  NAND2X0_HVT U234 ( .A1(n133), .A2(n134), .Y(\_0_net_[16] ) );
  NAND2X0_HVT U235 ( .A1(mc_out[95]), .A2(n117), .Y(n135) );
  NAND2X0_HVT U236 ( .A1(sr_out[95]), .A2(n83), .Y(n136) );
  NAND2X0_HVT U237 ( .A1(n135), .A2(n136), .Y(\_0_net_[95] ) );
  NAND2X0_HVT U238 ( .A1(mc_out[71]), .A2(n122), .Y(n139) );
  NAND2X0_HVT U239 ( .A1(n331), .A2(n433), .Y(n140) );
  NAND2X0_HVT U240 ( .A1(n139), .A2(n140), .Y(\_0_net_[71] ) );
  NAND2X0_HVT U241 ( .A1(mc_out[85]), .A2(n122), .Y(n141) );
  NAND2X0_HVT U242 ( .A1(sr_out[85]), .A2(n112), .Y(n142) );
  NAND2X0_HVT U243 ( .A1(n141), .A2(n142), .Y(\_0_net_[85] ) );
  NAND2X0_HVT U244 ( .A1(mc_out[10]), .A2(n115), .Y(n143) );
  NAND2X0_HVT U245 ( .A1(sr_out[10]), .A2(n83), .Y(n144) );
  NAND2X0_HVT U246 ( .A1(n143), .A2(n144), .Y(\_0_net_[10] ) );
  NAND2X0_HVT U247 ( .A1(mc_out[72]), .A2(n118), .Y(n145) );
  NAND2X0_HVT U248 ( .A1(n289), .A2(n112), .Y(n146) );
  NAND2X0_HVT U249 ( .A1(n145), .A2(n146), .Y(\_0_net_[72] ) );
  NAND2X0_HVT U250 ( .A1(mc_out[23]), .A2(n122), .Y(n147) );
  NAND2X0_HVT U251 ( .A1(sr_out[23]), .A2(n106), .Y(n148) );
  NAND2X0_HVT U252 ( .A1(n147), .A2(n148), .Y(\_0_net_[23] ) );
  NAND2X0_HVT U253 ( .A1(mc_out[77]), .A2(n75), .Y(n149) );
  NAND2X0_HVT U254 ( .A1(sr_out[77]), .A2(n87), .Y(n150) );
  NAND2X0_HVT U255 ( .A1(n149), .A2(n150), .Y(\_0_net_[77] ) );
  NAND2X0_HVT U256 ( .A1(mc_out[103]), .A2(n105), .Y(n151) );
  NAND2X0_HVT U257 ( .A1(n23), .A2(n106), .Y(n152) );
  NAND2X0_HVT U258 ( .A1(n151), .A2(n152), .Y(\_0_net_[103] ) );
  NAND2X0_HVT U259 ( .A1(mc_out[66]), .A2(n119), .Y(n153) );
  NAND2X0_HVT U260 ( .A1(sr_out[66]), .A2(n98), .Y(n154) );
  NAND2X0_HVT U261 ( .A1(n153), .A2(n154), .Y(\_0_net_[66] ) );
  NAND2X0_HVT U262 ( .A1(mc_out[93]), .A2(n117), .Y(n157) );
  NAND2X0_HVT U263 ( .A1(sr_out[93]), .A2(n87), .Y(n158) );
  NAND2X0_HVT U264 ( .A1(n157), .A2(n158), .Y(\_0_net_[93] ) );
  INVX1_HVT U265 ( .A(n159), .Y(keyout[35]) );
  NAND2X0_HVT U266 ( .A1(mc_out[83]), .A2(n114), .Y(n161) );
  NAND2X0_HVT U267 ( .A1(sr_out[83]), .A2(n103), .Y(n162) );
  NAND2X0_HVT U268 ( .A1(n161), .A2(n162), .Y(\_0_net_[83] ) );
  NAND2X0_HVT U269 ( .A1(mc_out[127]), .A2(n114), .Y(n163) );
  NAND2X0_HVT U270 ( .A1(n336), .A2(n100), .Y(n164) );
  NAND2X0_HVT U271 ( .A1(n163), .A2(n164), .Y(\_0_net_[127] ) );
  NAND2X0_HVT U272 ( .A1(n84), .A2(sr_out[62]), .Y(n252) );
  NAND2X0_HVT U273 ( .A1(mc_out[40]), .A2(n118), .Y(n165) );
  NAND2X0_HVT U274 ( .A1(sr_out[40]), .A2(n94), .Y(n166) );
  NAND2X0_HVT U275 ( .A1(n165), .A2(n166), .Y(\_0_net_[40] ) );
  NAND2X0_HVT U276 ( .A1(mc_out[8]), .A2(n114), .Y(n167) );
  NAND2X0_HVT U277 ( .A1(sr_out[8]), .A2(n98), .Y(n168) );
  NAND2X0_HVT U278 ( .A1(n167), .A2(n168), .Y(\_0_net_[8] ) );
  NAND2X0_HVT U279 ( .A1(mc_out[34]), .A2(n121), .Y(n169) );
  NAND2X0_HVT U280 ( .A1(n345), .A2(n103), .Y(n170) );
  NAND2X0_HVT U281 ( .A1(n169), .A2(n170), .Y(\_0_net_[34] ) );
  NAND2X0_HVT U282 ( .A1(mc_out[61]), .A2(n101), .Y(n171) );
  NAND2X0_HVT U283 ( .A1(sr_out[61]), .A2(n103), .Y(n172) );
  NAND2X0_HVT U284 ( .A1(n171), .A2(n172), .Y(\_0_net_[61] ) );
  NAND2X0_HVT U285 ( .A1(mc_out[0]), .A2(n76), .Y(n173) );
  NAND2X0_HVT U286 ( .A1(sr_out[0]), .A2(n83), .Y(n174) );
  NAND2X0_HVT U287 ( .A1(n173), .A2(n174), .Y(\_0_net_[0] ) );
  NAND2X0_HVT U288 ( .A1(n127), .A2(n94), .Y(n263) );
  NAND2X0_HVT U289 ( .A1(mc_out[21]), .A2(n117), .Y(n175) );
  NAND2X0_HVT U290 ( .A1(sr_out[21]), .A2(n110), .Y(n176) );
  NAND2X0_HVT U291 ( .A1(n175), .A2(n176), .Y(\_0_net_[21] ) );
  NAND2X0_HVT U292 ( .A1(mc_out[58]), .A2(n120), .Y(n177) );
  NAND2X0_HVT U293 ( .A1(n98), .A2(sr_out[58]), .Y(n178) );
  NAND2X0_HVT U294 ( .A1(n177), .A2(n178), .Y(\_0_net_[58] ) );
  NAND2X0_HVT U295 ( .A1(mc_out[45]), .A2(n116), .Y(n180) );
  NAND2X0_HVT U296 ( .A1(sr_out[45]), .A2(n97), .Y(n181) );
  NAND2X0_HVT U297 ( .A1(n180), .A2(n181), .Y(\_0_net_[45] ) );
  NAND2X0_HVT U298 ( .A1(mc_out[17]), .A2(n76), .Y(n182) );
  NAND2X0_HVT U299 ( .A1(n100), .A2(sr_out[17]), .Y(n183) );
  NAND2X0_HVT U300 ( .A1(n182), .A2(n183), .Y(\_0_net_[17] ) );
  NAND2X0_HVT U301 ( .A1(mc_out[37]), .A2(n114), .Y(n184) );
  NAND2X0_HVT U302 ( .A1(sr_out[37]), .A2(n429), .Y(n185) );
  NAND2X0_HVT U303 ( .A1(n184), .A2(n185), .Y(\_0_net_[37] ) );
  NAND2X0_HVT U304 ( .A1(mc_out[50]), .A2(n119), .Y(n186) );
  NAND2X0_HVT U305 ( .A1(n94), .A2(sr_out[50]), .Y(n187) );
  NAND2X0_HVT U306 ( .A1(n186), .A2(n187), .Y(\_0_net_[50] ) );
  INVX1_HVT U307 ( .A(n188), .Y(keyout[86]) );
  INVX1_HVT U308 ( .A(n190), .Y(keyout[74]) );
  NAND2X0_HVT U309 ( .A1(mc_out[52]), .A2(n105), .Y(n192) );
  NAND2X0_HVT U310 ( .A1(sr_out[52]), .A2(n83), .Y(n193) );
  NAND2X0_HVT U311 ( .A1(n192), .A2(n193), .Y(\_0_net_[52] ) );
  NAND2X0_HVT U312 ( .A1(sr_out[121]), .A2(n110), .Y(n301) );
  NAND2X0_HVT U313 ( .A1(mc_out[30]), .A2(n113), .Y(n194) );
  NAND2X0_HVT U314 ( .A1(sr_out[30]), .A2(n94), .Y(n195) );
  NAND2X0_HVT U315 ( .A1(n194), .A2(n195), .Y(\_0_net_[30] ) );
  NAND2X0_HVT U316 ( .A1(mc_out[25]), .A2(n117), .Y(n196) );
  NAND2X0_HVT U317 ( .A1(n31), .A2(n87), .Y(n197) );
  NAND2X0_HVT U318 ( .A1(n196), .A2(n197), .Y(\_0_net_[25] ) );
  NAND2X0_HVT U319 ( .A1(mc_out[15]), .A2(n113), .Y(n198) );
  NAND2X0_HVT U320 ( .A1(n421), .A2(n431), .Y(n199) );
  NAND2X0_HVT U321 ( .A1(n198), .A2(n199), .Y(\_0_net_[15] ) );
  NAND2X0_HVT U322 ( .A1(mc_out[26]), .A2(n120), .Y(n200) );
  NAND2X0_HVT U323 ( .A1(n200), .A2(n201), .Y(\_0_net_[26] ) );
  NAND2X0_HVT U324 ( .A1(mc_out[87]), .A2(n117), .Y(n202) );
  NAND2X0_HVT U325 ( .A1(sr_out[87]), .A2(n429), .Y(n203) );
  NAND2X0_HVT U326 ( .A1(n202), .A2(n203), .Y(\_0_net_[87] ) );
  INVX1_HVT U327 ( .A(n204), .Y(keyout[40]) );
  NAND2X0_HVT U328 ( .A1(sr_out[117]), .A2(n83), .Y(n297) );
  NAND2X0_HVT U329 ( .A1(n306), .A2(n84), .Y(n267) );
  NAND2X0_HVT U330 ( .A1(sr_out[27]), .A2(n430), .Y(n250) );
  NAND2X0_HVT U331 ( .A1(mc_out[65]), .A2(n76), .Y(n208) );
  NAND2X0_HVT U332 ( .A1(n112), .A2(sr_out[65]), .Y(n209) );
  NAND2X0_HVT U333 ( .A1(n208), .A2(n209), .Y(\_0_net_[65] ) );
  NAND2X0_HVT U334 ( .A1(mc_out[64]), .A2(n121), .Y(n210) );
  NAND2X0_HVT U335 ( .A1(n100), .A2(sr_out[64]), .Y(n211) );
  NAND2X0_HVT U336 ( .A1(n210), .A2(n211), .Y(\_0_net_[64] ) );
  NAND2X0_HVT U337 ( .A1(n216), .A2(n100), .Y(n215) );
  NAND2X0_HVT U338 ( .A1(n407), .A2(n110), .Y(n333) );
  NAND2X0_HVT U339 ( .A1(mc_out[80]), .A2(n120), .Y(n212) );
  NAND2X0_HVT U340 ( .A1(sr_out[80]), .A2(n84), .Y(n213) );
  NAND2X0_HVT U341 ( .A1(n212), .A2(n213), .Y(\_0_net_[80] ) );
  NAND2X0_HVT U342 ( .A1(mc_out[114]), .A2(n75), .Y(n214) );
  NAND2X0_HVT U343 ( .A1(n214), .A2(n215), .Y(\_0_net_[114] ) );
  NAND2X0_HVT U344 ( .A1(mc_out[92]), .A2(n117), .Y(n217) );
  NAND2X0_HVT U345 ( .A1(sr_out[92]), .A2(n103), .Y(n218) );
  NAND2X0_HVT U346 ( .A1(n217), .A2(n218), .Y(\_0_net_[92] ) );
  NAND2X0_HVT U347 ( .A1(n179), .A2(n103), .Y(n365) );
  NAND2X0_HVT U348 ( .A1(mc_out[59]), .A2(n85), .Y(n221) );
  NAND2X0_HVT U349 ( .A1(sr_out[59]), .A2(n107), .Y(n222) );
  NAND2X0_HVT U350 ( .A1(n221), .A2(n222), .Y(\_0_net_[59] ) );
  NAND2X0_HVT U351 ( .A1(mc_out[39]), .A2(n120), .Y(n223) );
  NAND2X0_HVT U352 ( .A1(n384), .A2(n97), .Y(n224) );
  NAND2X0_HVT U353 ( .A1(n223), .A2(n224), .Y(\_0_net_[39] ) );
  NAND2X0_HVT U354 ( .A1(mc_out[100]), .A2(n120), .Y(n225) );
  NAND2X0_HVT U355 ( .A1(n71), .A2(n110), .Y(n226) );
  NAND2X0_HVT U356 ( .A1(n225), .A2(n226), .Y(\_0_net_[100] ) );
  INVX1_HVT U357 ( .A(n227), .Y(keyout[34]) );
  NAND2X0_HVT U358 ( .A1(mc_out[54]), .A2(n76), .Y(n229) );
  NAND2X0_HVT U359 ( .A1(sr_out[54]), .A2(n87), .Y(n230) );
  NAND2X0_HVT U360 ( .A1(n229), .A2(n230), .Y(\_0_net_[54] ) );
  NAND2X0_HVT U361 ( .A1(mc_out[33]), .A2(n116), .Y(n231) );
  NAND2X0_HVT U362 ( .A1(sr_out[33]), .A2(n106), .Y(n232) );
  NAND2X0_HVT U363 ( .A1(n231), .A2(n232), .Y(\_0_net_[33] ) );
  NAND2X0_HVT U364 ( .A1(n107), .A2(sr_out[118]), .Y(n276) );
  NAND2X0_HVT U365 ( .A1(mc_out[56]), .A2(n118), .Y(n233) );
  NAND2X0_HVT U366 ( .A1(sr_out[56]), .A2(n100), .Y(n234) );
  NAND2X0_HVT U367 ( .A1(n233), .A2(n234), .Y(\_0_net_[56] ) );
  NAND2X0_HVT U368 ( .A1(sr_out[44]), .A2(n95), .Y(n291) );
  NAND2X0_HVT U369 ( .A1(mc_out[22]), .A2(n119), .Y(n235) );
  NAND2X0_HVT U370 ( .A1(sr_out[22]), .A2(n91), .Y(n236) );
  NAND2X0_HVT U371 ( .A1(n235), .A2(n236), .Y(\_0_net_[22] ) );
  NAND2X0_HVT U372 ( .A1(mc_out[35]), .A2(n75), .Y(n237) );
  NAND2X0_HVT U373 ( .A1(sr_out[35]), .A2(n106), .Y(n238) );
  NAND2X0_HVT U374 ( .A1(n237), .A2(n238), .Y(\_0_net_[35] ) );
  NAND2X0_HVT U375 ( .A1(mc_out[49]), .A2(n99), .Y(n239) );
  NAND2X0_HVT U376 ( .A1(sr_out[49]), .A2(n88), .Y(n240) );
  NAND2X0_HVT U377 ( .A1(n239), .A2(n240), .Y(\_0_net_[49] ) );
  NAND2X0_HVT U378 ( .A1(mc_out[55]), .A2(n115), .Y(n241) );
  NAND2X0_HVT U379 ( .A1(n319), .A2(n431), .Y(n242) );
  NAND2X0_HVT U380 ( .A1(n241), .A2(n242), .Y(\_0_net_[55] ) );
  NAND2X0_HVT U381 ( .A1(mc_out[24]), .A2(n118), .Y(n243) );
  NAND2X0_HVT U382 ( .A1(sr_out[24]), .A2(n91), .Y(n244) );
  NAND2X0_HVT U383 ( .A1(n243), .A2(n244), .Y(\_0_net_[24] ) );
  NAND2X0_HVT U384 ( .A1(mc_out[88]), .A2(n116), .Y(n245) );
  NAND2X0_HVT U385 ( .A1(n87), .A2(sr_out[88]), .Y(n246) );
  NAND2X0_HVT U386 ( .A1(n245), .A2(n246), .Y(\_0_net_[88] ) );
  NAND2X0_HVT U387 ( .A1(n387), .A2(n107), .Y(n283) );
  NAND2X0_HVT U388 ( .A1(mc_out[109]), .A2(n121), .Y(n247) );
  NAND2X0_HVT U389 ( .A1(sr_out[109]), .A2(n431), .Y(n248) );
  NAND2X0_HVT U390 ( .A1(n247), .A2(n248), .Y(\_0_net_[109] ) );
  NAND2X0_HVT U391 ( .A1(mc_out[27]), .A2(n105), .Y(n249) );
  NAND2X0_HVT U392 ( .A1(n249), .A2(n250), .Y(\_0_net_[27] ) );
  NAND2X0_HVT U393 ( .A1(mc_out[62]), .A2(n76), .Y(n251) );
  NAND2X0_HVT U394 ( .A1(n251), .A2(n252), .Y(\_0_net_[62] ) );
  INVX1_HVT U395 ( .A(n253), .Y(keyout[1]) );
  NAND2X0_HVT U396 ( .A1(mc_out[90]), .A2(n109), .Y(n255) );
  NAND2X0_HVT U397 ( .A1(sr_out[90]), .A2(n112), .Y(n256) );
  NAND2X0_HVT U398 ( .A1(n255), .A2(n256), .Y(\_0_net_[90] ) );
  NAND2X0_HVT U399 ( .A1(mc_out[74]), .A2(n114), .Y(n257) );
  NAND2X0_HVT U400 ( .A1(n257), .A2(n258), .Y(\_0_net_[74] ) );
  NAND2X0_HVT U401 ( .A1(mc_out[46]), .A2(n115), .Y(n260) );
  NAND2X0_HVT U402 ( .A1(n322), .A2(n95), .Y(n261) );
  NAND2X0_HVT U403 ( .A1(n260), .A2(n261), .Y(\_0_net_[46] ) );
  NAND2X0_HVT U404 ( .A1(mc_out[7]), .A2(n76), .Y(n262) );
  NAND2X0_HVT U405 ( .A1(n262), .A2(n263), .Y(\_0_net_[7] ) );
  NAND2X0_HVT U406 ( .A1(mc_out[126]), .A2(n75), .Y(n264) );
  NAND2X0_HVT U407 ( .A1(sr_out[126]), .A2(n98), .Y(n265) );
  NAND2X0_HVT U408 ( .A1(n264), .A2(n265), .Y(\_0_net_[126] ) );
  NAND2X0_HVT U409 ( .A1(mc_out[119]), .A2(n119), .Y(n266) );
  NAND2X0_HVT U410 ( .A1(n266), .A2(n267), .Y(\_0_net_[119] ) );
  NAND2X0_HVT U411 ( .A1(mc_out[75]), .A2(n109), .Y(n268) );
  NAND2X0_HVT U412 ( .A1(n268), .A2(n269), .Y(\_0_net_[75] ) );
  NAND2X0_HVT U413 ( .A1(n84), .A2(sr_out[51]), .Y(n299) );
  NAND2X0_HVT U414 ( .A1(mc_out[101]), .A2(n119), .Y(n270) );
  NAND2X0_HVT U415 ( .A1(n98), .A2(sr_out[101]), .Y(n271) );
  NAND2X0_HVT U416 ( .A1(n270), .A2(n271), .Y(\_0_net_[101] ) );
  NAND2X0_HVT U417 ( .A1(mc_out[6]), .A2(n122), .Y(n273) );
  NAND2X0_HVT U418 ( .A1(sr_out[6]), .A2(n106), .Y(n274) );
  NAND2X0_HVT U419 ( .A1(n273), .A2(n274), .Y(\_0_net_[6] ) );
  NAND2X0_HVT U420 ( .A1(mc_out[118]), .A2(n121), .Y(n275) );
  NAND2X0_HVT U421 ( .A1(n275), .A2(n276), .Y(\_0_net_[118] ) );
  NAND2X0_HVT U422 ( .A1(mc_out[9]), .A2(n99), .Y(n277) );
  NAND2X0_HVT U423 ( .A1(sr_out[9]), .A2(n107), .Y(n278) );
  NAND2X0_HVT U424 ( .A1(n277), .A2(n278), .Y(\_0_net_[9] ) );
  NAND2X0_HVT U425 ( .A1(mc_out[108]), .A2(n121), .Y(n280) );
  NAND2X0_HVT U426 ( .A1(n280), .A2(n281), .Y(\_0_net_[108] ) );
  NAND2X0_HVT U427 ( .A1(mc_out[60]), .A2(n75), .Y(n282) );
  NAND2X0_HVT U428 ( .A1(n282), .A2(n283), .Y(\_0_net_[60] ) );
  NAND2X0_HVT U429 ( .A1(mc_out[2]), .A2(n113), .Y(n284) );
  NAND2X0_HVT U430 ( .A1(n284), .A2(n285), .Y(\_0_net_[2] ) );
  NAND2X0_HVT U431 ( .A1(mc_out[123]), .A2(n119), .Y(n287) );
  NAND2X0_HVT U432 ( .A1(sr_out[123]), .A2(n100), .Y(n288) );
  NAND2X0_HVT U433 ( .A1(n287), .A2(n288), .Y(\_0_net_[123] ) );
  NAND2X0_HVT U434 ( .A1(mc_out[44]), .A2(n118), .Y(n290) );
  NAND2X0_HVT U435 ( .A1(n290), .A2(n291), .Y(\_0_net_[44] ) );
  NAND2X0_HVT U436 ( .A1(mc_out[98]), .A2(n122), .Y(n292) );
  NAND2X0_HVT U437 ( .A1(sr_out[98]), .A2(n88), .Y(n293) );
  NAND2X0_HVT U438 ( .A1(n292), .A2(n293), .Y(\_0_net_[98] ) );
  NAND2X0_HVT U439 ( .A1(mc_out[13]), .A2(n75), .Y(n294) );
  NAND2X0_HVT U440 ( .A1(n103), .A2(sr_out[13]), .Y(n295) );
  NAND2X0_HVT U441 ( .A1(n295), .A2(n294), .Y(\_0_net_[13] ) );
  NAND2X0_HVT U442 ( .A1(mc_out[117]), .A2(n105), .Y(n296) );
  NAND2X0_HVT U443 ( .A1(n296), .A2(n297), .Y(\_0_net_[117] ) );
  NAND2X0_HVT U444 ( .A1(mc_out[51]), .A2(n118), .Y(n298) );
  NAND2X0_HVT U445 ( .A1(n298), .A2(n299), .Y(\_0_net_[51] ) );
  NAND2X0_HVT U446 ( .A1(mc_out[121]), .A2(n122), .Y(n300) );
  NAND2X0_HVT U447 ( .A1(n300), .A2(n301), .Y(\_0_net_[121] ) );
  NAND2X0_HVT U448 ( .A1(mc_out[48]), .A2(n75), .Y(n302) );
  NAND2X0_HVT U449 ( .A1(n302), .A2(n303), .Y(\_0_net_[48] ) );
  NAND2X0_HVT U450 ( .A1(mc_out[69]), .A2(n121), .Y(n304) );
  NAND2X0_HVT U451 ( .A1(n91), .A2(sr_out[69]), .Y(n305) );
  NAND2X0_HVT U452 ( .A1(n304), .A2(n305), .Y(\_0_net_[69] ) );
  NAND2X0_HVT U453 ( .A1(n110), .A2(sr_out[107]), .Y(n324) );
  NAND2X0_HVT U454 ( .A1(mc_out[53]), .A2(n90), .Y(n307) );
  NAND2X0_HVT U455 ( .A1(n107), .A2(sr_out[53]), .Y(n308) );
  NAND2X0_HVT U456 ( .A1(n307), .A2(n308), .Y(\_0_net_[53] ) );
  NAND2X0_HVT U457 ( .A1(mc_out[96]), .A2(n115), .Y(n309) );
  NAND2X0_HVT U458 ( .A1(n98), .A2(sr_out[96]), .Y(n310) );
  NAND2X0_HVT U459 ( .A1(n309), .A2(n310), .Y(\_0_net_[96] ) );
  NAND2X0_HVT U460 ( .A1(mc_out[89]), .A2(n86), .Y(n311) );
  NAND2X0_HVT U461 ( .A1(n430), .A2(sr_out[89]), .Y(n312) );
  NAND2X0_HVT U462 ( .A1(n311), .A2(n312), .Y(\_0_net_[89] ) );
  NAND2X0_HVT U463 ( .A1(mc_out[19]), .A2(n118), .Y(n313) );
  NAND2X0_HVT U464 ( .A1(n404), .A2(n97), .Y(n314) );
  NAND2X0_HVT U465 ( .A1(n313), .A2(n314), .Y(\_0_net_[19] ) );
  NAND2X0_HVT U466 ( .A1(mc_out[79]), .A2(n93), .Y(n315) );
  NAND2X0_HVT U467 ( .A1(n279), .A2(n88), .Y(n316) );
  NAND2X0_HVT U468 ( .A1(n315), .A2(n316), .Y(\_0_net_[79] ) );
  NAND2X0_HVT U469 ( .A1(mc_out[113]), .A2(n115), .Y(n317) );
  NAND2X0_HVT U470 ( .A1(sr_out[113]), .A2(n429), .Y(n318) );
  NAND2X0_HVT U471 ( .A1(n317), .A2(n318), .Y(\_0_net_[113] ) );
  NAND2X0_HVT U472 ( .A1(mc_out[57]), .A2(n113), .Y(n320) );
  NAND2X0_HVT U473 ( .A1(n320), .A2(n321), .Y(\_0_net_[57] ) );
  NAND2X0_HVT U474 ( .A1(mc_out[107]), .A2(n122), .Y(n323) );
  NAND2X0_HVT U475 ( .A1(n323), .A2(n324), .Y(\_0_net_[107] ) );
  NAND2X0_HVT U476 ( .A1(mc_out[106]), .A2(n121), .Y(n325) );
  NAND2X0_HVT U477 ( .A1(n103), .A2(sr_out[106]), .Y(n326) );
  NAND2X0_HVT U478 ( .A1(n325), .A2(n326), .Y(\_0_net_[106] ) );
  NAND2X0_HVT U479 ( .A1(mc_out[91]), .A2(n99), .Y(n327) );
  NAND2X0_HVT U480 ( .A1(n88), .A2(sr_out[91]), .Y(n328) );
  NAND2X0_HVT U481 ( .A1(n327), .A2(n328), .Y(\_0_net_[91] ) );
  NAND2X0_HVT U482 ( .A1(mc_out[124]), .A2(n90), .Y(n329) );
  NAND2X0_HVT U483 ( .A1(n112), .A2(sr_out[124]), .Y(n330) );
  NAND2X0_HVT U484 ( .A1(n329), .A2(n330), .Y(\_0_net_[124] ) );
  NAND2X0_HVT U485 ( .A1(mc_out[41]), .A2(n122), .Y(n332) );
  NAND2X0_HVT U486 ( .A1(n332), .A2(n333), .Y(\_0_net_[41] ) );
  INVX1_HVT U487 ( .A(n334), .Y(keyout[50]) );
  NAND2X0_HVT U488 ( .A1(mc_out[31]), .A2(n92), .Y(n337) );
  NAND2X0_HVT U489 ( .A1(sr_out[31]), .A2(n84), .Y(n338) );
  NAND2X0_HVT U490 ( .A1(n337), .A2(n338), .Y(\_0_net_[31] ) );
  NAND2X0_HVT U491 ( .A1(mc_out[112]), .A2(n117), .Y(n339) );
  NAND2X0_HVT U492 ( .A1(sr_out[112]), .A2(n430), .Y(n340) );
  NAND2X0_HVT U493 ( .A1(n339), .A2(n340), .Y(\_0_net_[112] ) );
  NAND2X0_HVT U494 ( .A1(mc_out[116]), .A2(n120), .Y(n341) );
  NAND2X0_HVT U495 ( .A1(sr_out[116]), .A2(n83), .Y(n342) );
  NAND2X0_HVT U496 ( .A1(n341), .A2(n342), .Y(\_0_net_[116] ) );
  NAND2X0_HVT U497 ( .A1(mc_out[28]), .A2(n120), .Y(n343) );
  NAND2X0_HVT U498 ( .A1(n87), .A2(n130), .Y(n344) );
  NAND2X0_HVT U499 ( .A1(n343), .A2(n344), .Y(\_0_net_[28] ) );
  NAND2X0_HVT U500 ( .A1(mc_out[115]), .A2(n82), .Y(n348) );
  NAND2X0_HVT U501 ( .A1(n94), .A2(sr_out[115]), .Y(n349) );
  NAND2X0_HVT U502 ( .A1(n348), .A2(n349), .Y(\_0_net_[115] ) );
  NAND2X0_HVT U503 ( .A1(mc_out[120]), .A2(n113), .Y(n350) );
  NAND2X0_HVT U504 ( .A1(n103), .A2(sr_out[120]), .Y(n351) );
  NAND2X0_HVT U505 ( .A1(n350), .A2(n351), .Y(\_0_net_[120] ) );
  INVX1_HVT U506 ( .A(n354), .Y(keyout[43]) );
  INVX1_HVT U507 ( .A(n356), .Y(keyout[14]) );
  NAND2X0_HVT U508 ( .A1(mc_out[78]), .A2(n104), .Y(n358) );
  NAND2X0_HVT U509 ( .A1(sr_out[78]), .A2(n110), .Y(n359) );
  NAND2X0_HVT U510 ( .A1(n358), .A2(n359), .Y(\_0_net_[78] ) );
  NAND2X0_HVT U511 ( .A1(mc_out[73]), .A2(n120), .Y(n360) );
  NAND2X0_HVT U512 ( .A1(n286), .A2(n84), .Y(n361) );
  NAND2X0_HVT U513 ( .A1(n360), .A2(n361), .Y(\_0_net_[73] ) );
  NAND2X0_HVT U514 ( .A1(mc_out[67]), .A2(n108), .Y(n362) );
  NAND2X0_HVT U515 ( .A1(n362), .A2(n363), .Y(\_0_net_[67] ) );
  NAND2X0_HVT U516 ( .A1(mc_out[97]), .A2(n109), .Y(n364) );
  NAND2X0_HVT U517 ( .A1(n364), .A2(n365), .Y(\_0_net_[97] ) );
  INVX1_HVT U518 ( .A(n366), .Y(keyout[78]) );
  NAND2X0_HVT U519 ( .A1(sr_out[12]), .A2(n88), .Y(n375) );
  NAND2X0_HVT U520 ( .A1(sr_out[3]), .A2(n110), .Y(n371) );
  NAND2X0_HVT U521 ( .A1(mc_out[105]), .A2(n76), .Y(n368) );
  NAND2X0_HVT U522 ( .A1(sr_out[105]), .A2(n97), .Y(n369) );
  NAND2X0_HVT U523 ( .A1(n368), .A2(n369), .Y(\_0_net_[105] ) );
  NAND2X0_HVT U524 ( .A1(mc_out[3]), .A2(n76), .Y(n370) );
  NAND2X0_HVT U525 ( .A1(n370), .A2(n371), .Y(\_0_net_[3] ) );
  NAND2X0_HVT U526 ( .A1(mc_out[81]), .A2(n109), .Y(n372) );
  NAND2X0_HVT U527 ( .A1(n396), .A2(n428), .Y(n373) );
  NAND2X0_HVT U528 ( .A1(n372), .A2(n373), .Y(\_0_net_[81] ) );
  NAND2X0_HVT U529 ( .A1(mc_out[12]), .A2(n118), .Y(n374) );
  NAND2X0_HVT U530 ( .A1(n374), .A2(n375), .Y(\_0_net_[12] ) );
  NAND2X0_HVT U531 ( .A1(mc_out[99]), .A2(n114), .Y(n376) );
  NAND2X0_HVT U532 ( .A1(n83), .A2(sr_out[99]), .Y(n377) );
  NAND2X0_HVT U533 ( .A1(n376), .A2(n377), .Y(\_0_net_[99] ) );
  INVX1_HVT U534 ( .A(n378), .Y(keyout[41]) );
  NAND2X0_HVT U535 ( .A1(mc_out[4]), .A2(n120), .Y(n380) );
  NAND2X0_HVT U536 ( .A1(n399), .A2(n84), .Y(n381) );
  NAND2X0_HVT U537 ( .A1(n380), .A2(n381), .Y(\_0_net_[4] ) );
  INVX1_HVT U538 ( .A(n382), .Y(keyout[59]) );
  NAND2X0_HVT U539 ( .A1(mc_out[1]), .A2(n117), .Y(n385) );
  NAND2X0_HVT U540 ( .A1(n259), .A2(n91), .Y(n386) );
  NAND2X0_HVT U541 ( .A1(n385), .A2(n386), .Y(\_0_net_[1] ) );
  NAND2X0_HVT U542 ( .A1(mc_out[63]), .A2(n76), .Y(n388) );
  NAND2X0_HVT U543 ( .A1(sr_out[63]), .A2(n88), .Y(n389) );
  NAND2X0_HVT U544 ( .A1(n388), .A2(n389), .Y(\_0_net_[63] ) );
  NAND2X0_HVT U545 ( .A1(mc_out[43]), .A2(n117), .Y(n390) );
  NAND2X0_HVT U546 ( .A1(sr_out[43]), .A2(n429), .Y(n391) );
  NAND2X0_HVT U547 ( .A1(n390), .A2(n391), .Y(\_0_net_[43] ) );
  INVX1_HVT U548 ( .A(n392), .Y(keyout[87]) );
  INVX1_HVT U549 ( .A(n394), .Y(keyout[54]) );
  INVX1_HVT U550 ( .A(n397), .Y(keyout[53]) );
  INVX1_HVT U551 ( .A(n405), .Y(keyout[65]) );
  INVX1_HVT U552 ( .A(n410), .Y(keyout[77]) );
  NAND2X0_HVT U553 ( .A1(mc_out[125]), .A2(n75), .Y(n412) );
  NAND2X0_HVT U554 ( .A1(sr_out[125]), .A2(n430), .Y(n413) );
  NAND2X0_HVT U555 ( .A1(n412), .A2(n413), .Y(\_0_net_[125] ) );
  INVX1_HVT U556 ( .A(n414), .Y(keyout[95]) );
  INVX1_HVT U557 ( .A(n419), .Y(keyout[29]) );
  NAND2X0_HVT U558 ( .A1(mc_out[20]), .A2(n113), .Y(n422) );
  NAND2X0_HVT U559 ( .A1(n95), .A2(n79), .Y(n423) );
  NAND2X0_HVT U560 ( .A1(n422), .A2(n423), .Y(\_0_net_[20] ) );
  INVX1_HVT U561 ( .A(n424), .Y(keyout[36]) );
endmodule

