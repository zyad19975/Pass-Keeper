
module inv_sbox_6 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n196, n197, n198, n199, n200, n201, n202, n208, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623;

  NAND2X0_HVT U1 ( .A1(n303), .A2(n327), .Y(n623) );
  NAND2X0_HVT U3 ( .A1(n303), .A2(in[6]), .Y(n621) );
  NAND2X0_HVT U4 ( .A1(n286), .A2(n340), .Y(n620) );
  NAND2X0_HVT U6 ( .A1(n345), .A2(n305), .Y(n617) );
  NAND2X0_HVT U8 ( .A1(n347), .A2(n336), .Y(n615) );
  NAND2X0_HVT U9 ( .A1(n342), .A2(n615), .Y(n614) );
  NAND2X0_HVT U10 ( .A1(n304), .A2(n612), .Y(n613) );
  NAND2X0_HVT U11 ( .A1(n349), .A2(n341), .Y(n611) );
  NAND2X0_HVT U12 ( .A1(n345), .A2(n324), .Y(n610) );
  NAND2X0_HVT U13 ( .A1(n339), .A2(n615), .Y(n609) );
  NAND2X0_HVT U15 ( .A1(n333), .A2(n263), .Y(n607) );
  NAND2X0_HVT U19 ( .A1(n287), .A2(n412), .Y(n602) );
  NAND2X0_HVT U25 ( .A1(in[6]), .A2(n325), .Y(n618) );
  NAND2X0_HVT U32 ( .A1(n327), .A2(n349), .Y(n590) );
  NAND2X0_HVT U35 ( .A1(n615), .A2(n413), .Y(n587) );
  NAND2X0_HVT U38 ( .A1(n324), .A2(n349), .Y(n584) );
  NAND2X0_HVT U42 ( .A1(n617), .A2(n413), .Y(n580) );
  OA21X1_HVT U53 ( .A1(n302), .A2(n572), .A3(n248), .Y(n570) );
  NAND2X0_HVT U55 ( .A1(n339), .A2(n199), .Y(n568) );
  MUX41X1_HVT U56 ( .A1(n393), .A3(n334), .A2(n377), .A4(n198), .S0(n314), 
        .S1(n352), .Y(n567) );
  AO21X1_HVT U60 ( .A1(n562), .A2(n321), .A3(n601), .Y(n563) );
  NAND2X0_HVT U66 ( .A1(n263), .A2(n295), .Y(n556) );
  MUX41X1_HVT U67 ( .A1(n367), .A3(n394), .A2(n369), .A4(n556), .S0(n323), 
        .S1(n315), .Y(n555) );
  MUX41X1_HVT U68 ( .A1(n367), .A3(n239), .A2(n368), .A4(n304), .S0(n317), 
        .S1(n267), .Y(n554) );
  MUX41X1_HVT U69 ( .A1(n554), .A3(n557), .A2(n555), .A4(n558), .S0(n266), 
        .S1(n330), .Y(n553) );
  NAND2X0_HVT U72 ( .A1(n334), .A2(n247), .Y(n551) );
  MUX41X1_HVT U73 ( .A1(n595), .A3(n551), .A2(n395), .A4(n324), .S0(n322), 
        .S1(n314), .Y(n550) );
  MUX41X1_HVT U74 ( .A1(n613), .A3(n383), .A2(n382), .A4(n245), .S0(n314), 
        .S1(n268), .Y(n549) );
  MUX41X1_HVT U78 ( .A1(n546), .A3(n550), .A2(n549), .A4(n552), .S0(n266), 
        .S1(n330), .Y(n545) );
  MUX41X1_HVT U80 ( .A1(n397), .A3(n393), .A2(n614), .A4(n619), .S0(n317), 
        .S1(n352), .Y(n543) );
  NAND2X0_HVT U81 ( .A1(n341), .A2(n616), .Y(n542) );
  AND2X1_HVT U82 ( .A1(n617), .A2(n337), .Y(n541) );
  MUX41X1_HVT U83 ( .A1(n541), .A3(n380), .A2(n297), .A4(n542), .S0(n317), 
        .S1(n352), .Y(n540) );
  MUX41X1_HVT U84 ( .A1(n312), .A3(n379), .A2(n398), .A4(n253), .S0(n318), 
        .S1(n267), .Y(n539) );
  MUX41X1_HVT U85 ( .A1(n539), .A3(n543), .A2(n540), .A4(n544), .S0(n266), 
        .S1(n330), .Y(n538) );
  MUX41X1_HVT U87 ( .A1(n360), .A3(n312), .A2(n399), .A4(n377), .S0(n316), 
        .S1(n323), .Y(n537) );
  NAND2X0_HVT U89 ( .A1(n349), .A2(n409), .Y(n535) );
  MUX41X1_HVT U90 ( .A1(n411), .A3(n247), .A2(n575), .A4(n535), .S0(n317), 
        .S1(n267), .Y(n534) );
  MUX41X1_HVT U98 ( .A1(n527), .A3(n401), .A2(n385), .A4(n594), .S0(n315), 
        .S1(n353), .Y(n526) );
  MUX41X1_HVT U99 ( .A1(n590), .A3(n371), .A2(n574), .A4(n333), .S0(n268), 
        .S1(n315), .Y(n525) );
  NAND2X0_HVT U100 ( .A1(n349), .A2(n408), .Y(n524) );
  MUX41X1_HVT U101 ( .A1(n402), .A3(n610), .A2(n384), .A4(n524), .S0(n267), 
        .S1(n318), .Y(n523) );
  AND2X1_HVT U104 ( .A1(n616), .A2(n335), .Y(n521) );
  MUX41X1_HVT U105 ( .A1(n608), .A3(n403), .A2(n542), .A4(n521), .S0(n314), 
        .S1(n352), .Y(n520) );
  MUX41X1_HVT U107 ( .A1(n402), .A3(n337), .A2(n519), .A4(n361), .S0(n317), 
        .S1(n268), .Y(n518) );
  MUX41X1_HVT U108 ( .A1(n245), .A3(n333), .A2(n377), .A4(n341), .S0(n320), 
        .S1(n267), .Y(n517) );
  MUX41X1_HVT U109 ( .A1(n401), .A3(n357), .A2(n398), .A4(n391), .S0(n317), 
        .S1(n268), .Y(n516) );
  MUX41X1_HVT U110 ( .A1(n516), .A3(n518), .A2(n517), .A4(n520), .S0(n266), 
        .S1(n288), .Y(n515) );
  AO21X1_HVT U112 ( .A1(n387), .A2(n322), .A3(n598), .Y(n513) );
  NAND2X0_HVT U114 ( .A1(n342), .A2(n247), .Y(n511) );
  MUX41X1_HVT U115 ( .A1(n511), .A3(n611), .A2(n387), .A4(n337), .S0(n267), 
        .S1(n315), .Y(n510) );
  MUX41X1_HVT U116 ( .A1(n386), .A3(n379), .A2(n357), .A4(n607), .S0(n316), 
        .S1(n267), .Y(n509) );
  NAND2X0_HVT U118 ( .A1(n349), .A2(n239), .Y(n507) );
  MUX41X1_HVT U119 ( .A1(n404), .A3(n508), .A2(n585), .A4(n507), .S0(n316), 
        .S1(n353), .Y(n506) );
  MUX41X1_HVT U122 ( .A1(n392), .A3(n308), .A2(n576), .A4(n396), .S0(n316), 
        .S1(n353), .Y(n504) );
  MUX41X1_HVT U124 ( .A1(n310), .A3(n503), .A2(n599), .A4(n374), .S0(n321), 
        .S1(n316), .Y(n502) );
  AOI21X1_HVT U127 ( .A1(n320), .A2(n498), .A3(n362), .Y(n499) );
  NAND2X0_HVT U129 ( .A1(n319), .A2(n342), .Y(n496) );
  MUX41X1_HVT U130 ( .A1(n496), .A3(n497), .A2(n500), .A4(n499), .S0(n323), 
        .S1(n288), .Y(n495) );
  AND2X1_HVT U131 ( .A1(n295), .A2(n269), .Y(n494) );
  MUX41X1_HVT U132 ( .A1(n237), .A3(n494), .A2(n406), .A4(n367), .S0(n322), 
        .S1(n314), .Y(n493) );
  MUX41X1_HVT U133 ( .A1(n407), .A3(n361), .A2(n198), .A4(n292), .S0(n321), 
        .S1(n315), .Y(n492) );
  MUX41X1_HVT U136 ( .A1(n573), .A3(n524), .A2(n490), .A4(n365), .S0(n319), 
        .S1(n352), .Y(n489) );
  MUX41X1_HVT U137 ( .A1(n615), .A3(n593), .A2(n253), .A4(n400), .S0(n323), 
        .S1(n318), .Y(n488) );
  MUX41X1_HVT U139 ( .A1(n487), .A3(n491), .A2(n495), .A4(n501), .S0(n266), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n382), .A3(n309), .A2(n376), .A4(n611), .S0(n322), 
        .S1(n315), .Y(n486) );
  NAND2X0_HVT U141 ( .A1(n333), .A2(n349), .Y(n485) );
  MUX41X1_HVT U142 ( .A1(n485), .A3(n583), .A2(n405), .A4(n376), .S0(n320), 
        .S1(n353), .Y(n484) );
  MUX41X1_HVT U151 ( .A1(n297), .A3(n385), .A2(n296), .A4(n476), .S0(n321), 
        .S1(n315), .Y(n475) );
  MUX41X1_HVT U155 ( .A1(n376), .A3(n611), .A2(n603), .A4(n378), .S0(n318), 
        .S1(n353), .Y(n471) );
  NAND2X0_HVT U159 ( .A1(n467), .A2(n466), .Y(n468) );
  MUX41X1_HVT U162 ( .A1(n389), .A3(n372), .A2(n587), .A4(n464), .S0(n318), 
        .S1(n352), .Y(n463) );
  NAND2X0_HVT U163 ( .A1(n344), .A2(n409), .Y(n462) );
  MUX41X1_HVT U164 ( .A1(n614), .A3(n462), .A2(n585), .A4(n245), .S0(n316), 
        .S1(n352), .Y(n461) );
  NAND2X0_HVT U166 ( .A1(n612), .A2(n458), .Y(n459) );
  MUX41X1_HVT U172 ( .A1(n535), .A3(n453), .A2(n307), .A4(n600), .S0(n318), 
        .S1(n268), .Y(n452) );
  MUX41X1_HVT U174 ( .A1(n399), .A3(n198), .A2(n407), .A4(n413), .S0(n318), 
        .S1(n353), .Y(n450) );
  NAND2X0_HVT U177 ( .A1(n343), .A2(n239), .Y(n448) );
  AND2X1_HVT U179 ( .A1(n617), .A2(n335), .Y(n446) );
  MUX41X1_HVT U182 ( .A1(n361), .A3(n199), .A2(n360), .A4(n297), .S0(n316), 
        .S1(n353), .Y(n443) );
  MUX41X1_HVT U183 ( .A1(n388), .A3(n393), .A2(n373), .A4(n580), .S0(n321), 
        .S1(n314), .Y(n442) );
  AND2X1_HVT U185 ( .A1(n413), .A2(n269), .Y(n440) );
  NAND2X0_HVT U191 ( .A1(n270), .A2(n366), .Y(n434) );
  AND2X1_HVT U192 ( .A1(n383), .A2(n432), .Y(n433) );
  NAND2X0_HVT U194 ( .A1(n580), .A2(n432), .Y(n430) );
  MUX41X1_HVT U195 ( .A1(n431), .A3(n430), .A2(n433), .A4(n434), .S0(n317), 
        .S1(n331), .Y(n429) );
  NAND2X0_HVT U198 ( .A1(n345), .A2(n413), .Y(n612) );
  NAND2X0_HVT U200 ( .A1(n336), .A2(n349), .Y(n498) );
  NAND2X0_HVT U207 ( .A1(n349), .A2(n411), .Y(n562) );
  MUX41X1_HVT U2 ( .A1(n536), .A3(n530), .A2(n537), .A4(n534), .S0(n332), .S1(
        n330), .Y(n529) );
  INVX1_HVT U5 ( .A(n332), .Y(n266) );
  MUX41X1_HVT U7 ( .A1(n411), .A3(n342), .A2(n586), .A4(n341), .S0(n196), .S1(
        n268), .Y(n451) );
  IBUFFX16_HVT U14 ( .A(n318), .Y(n196) );
  IBUFFX2_HVT U16 ( .A(n576), .Y(n391) );
  MUX21X2_HVT U17 ( .A1(n395), .A2(n581), .S0(n322), .Y(n437) );
  INVX1_HVT U18 ( .A(n596), .Y(n377) );
  INVX0_HVT U20 ( .A(n296), .Y(n600) );
  MUX21X2_HVT U21 ( .A1(n340), .A2(n222), .S0(n269), .Y(n296) );
  INVX0_HVT U22 ( .A(n568), .Y(n197) );
  INVX1_HVT U23 ( .A(n197), .Y(n198) );
  INVX1_HVT U24 ( .A(n360), .Y(n199) );
  INVX0_HVT U26 ( .A(n620), .Y(n360) );
  MUX41X1_HVT U27 ( .A1(n457), .A3(n463), .A2(n461), .A4(n465), .S0(n200), 
        .S1(n201), .Y(n456) );
  IBUFFX16_HVT U28 ( .A(n332), .Y(n200) );
  IBUFFX16_HVT U29 ( .A(n272), .Y(n201) );
  IBUFFX2_HVT U30 ( .A(n410), .Y(n303) );
  IBUFFX2_HVT U31 ( .A(n324), .Y(n298) );
  MUX41X1_HVT U33 ( .A1(n565), .A3(n569), .A2(n561), .A4(n567), .S0(n266), 
        .S1(n202), .Y(n560) );
  IBUFFX16_HVT U34 ( .A(n330), .Y(n202) );
  INVX1_HVT U36 ( .A(n237), .Y(n619) );
  XNOR2X2_HVT U37 ( .A1(n302), .A2(n316), .Y(n313) );
  INVX0_HVT U39 ( .A(n599), .Y(n374) );
  MUX21X2_HVT U40 ( .A1(n619), .A2(n376), .S0(n261), .Y(n566) );
  INVX1_HVT U41 ( .A(n597), .Y(n376) );
  NAND2X0_HVT U43 ( .A1(n342), .A2(n208), .Y(n218) );
  NAND2X0_HVT U44 ( .A1(n341), .A2(n344), .Y(n219) );
  NAND2X0_HVT U45 ( .A1(n218), .A2(n219), .Y(n608) );
  IBUFFX2_HVT U46 ( .A(n344), .Y(n208) );
  MUX21X2_HVT U47 ( .A1(n568), .A2(n374), .S0(n220), .Y(n564) );
  IBUFFX16_HVT U48 ( .A(n322), .Y(n220) );
  INVX0_HVT U49 ( .A(n606), .Y(n221) );
  INVX0_HVT U50 ( .A(n221), .Y(n222) );
  NBUFFX4_HVT U51 ( .A(n414), .Y(n326) );
  MUX41X1_HVT U52 ( .A1(n576), .A3(n592), .A2(n357), .A4(n369), .S0(n244), 
        .S1(n354), .Y(n536) );
  IBUFFX2_HVT U54 ( .A(n354), .Y(n267) );
  INVX1_HVT U57 ( .A(n622), .Y(n408) );
  NAND2X0_HVT U58 ( .A1(n553), .A2(n249), .Y(n250) );
  MUX21X1_HVT U59 ( .A1(n296), .A2(n199), .S0(n319), .Y(n559) );
  MUX21X1_HVT U61 ( .A1(n328), .A2(n337), .S0(n262), .Y(n223) );
  IBUFFX16_HVT U62 ( .A(n223), .Y(n581) );
  MUX21X1_HVT U63 ( .A1(n223), .A2(n225), .S0(n226), .Y(n224) );
  IBUFFX16_HVT U64 ( .A(n224), .Y(n514) );
  IBUFFX16_HVT U65 ( .A(n362), .Y(n225) );
  IBUFFX16_HVT U70 ( .A(n323), .Y(n226) );
  INVX1_HVT U71 ( .A(n328), .Y(n295) );
  XNOR2X2_HVT U75 ( .A1(n326), .A2(n325), .Y(n606) );
  INVX0_HVT U76 ( .A(n606), .Y(n413) );
  MUX21X1_HVT U77 ( .A1(n312), .A2(n597), .S0(n270), .Y(n474) );
  NAND2X0_HVT U79 ( .A1(n480), .A2(n227), .Y(n228) );
  NAND2X0_HVT U86 ( .A1(n470), .A2(n235), .Y(n229) );
  NAND2X0_HVT U88 ( .A1(n228), .A2(n229), .Y(out[5]) );
  INVX1_HVT U91 ( .A(n235), .Y(n227) );
  IBUFFX2_HVT U92 ( .A(in[7]), .Y(n235) );
  MUX21X2_HVT U93 ( .A1(n245), .A2(n559), .S0(n313), .Y(n558) );
  MUX21X2_HVT U94 ( .A1(n563), .A2(n564), .S0(n230), .Y(n561) );
  IBUFFX16_HVT U95 ( .A(n319), .Y(n230) );
  MUX21X2_HVT U96 ( .A1(n411), .A2(n333), .S0(n231), .Y(n591) );
  IBUFFX16_HVT U97 ( .A(n240), .Y(n231) );
  NAND2X0_HVT U102 ( .A1(n443), .A2(n232), .Y(n233) );
  NAND2X0_HVT U103 ( .A1(n442), .A2(n259), .Y(n234) );
  NAND2X0_HVT U106 ( .A1(n233), .A2(n234), .Y(n441) );
  INVX0_HVT U111 ( .A(n259), .Y(n232) );
  IBUFFX2_HVT U113 ( .A(n331), .Y(n259) );
  NBUFFX4_HVT U117 ( .A(n410), .Y(n324) );
  AO21X1_HVT U120 ( .A1(n240), .A2(n408), .A3(n302), .Y(n432) );
  MUX21X1_HVT U121 ( .A1(n239), .A2(n408), .S0(n236), .Y(n599) );
  IBUFFX16_HVT U123 ( .A(n241), .Y(n236) );
  INVX1_HVT U125 ( .A(n416), .Y(n406) );
  INVX1_HVT U126 ( .A(in[5]), .Y(n258) );
  AND2X1_HVT U128 ( .A1(n620), .A2(n336), .Y(n237) );
  INVX1_HVT U134 ( .A(n303), .Y(n238) );
  INVX2_HVT U135 ( .A(n238), .Y(n239) );
  IBUFFX2_HVT U138 ( .A(n348), .Y(n240) );
  IBUFFX2_HVT U143 ( .A(n348), .Y(n241) );
  INVX2_HVT U144 ( .A(in[0]), .Y(n348) );
  MUX21X2_HVT U145 ( .A1(n459), .A2(n460), .S0(n319), .Y(n457) );
  MUX21X2_HVT U146 ( .A1(n396), .A2(n579), .S0(n270), .Y(n469) );
  MUX21X2_HVT U147 ( .A1(n515), .A2(n505), .S0(n242), .Y(out[3]) );
  IBUFFX16_HVT U148 ( .A(in[7]), .Y(n242) );
  INVX0_HVT U149 ( .A(n580), .Y(n361) );
  INVX1_HVT U150 ( .A(n248), .Y(n594) );
  INVX0_HVT U152 ( .A(n586), .Y(n384) );
  INVX0_HVT U153 ( .A(n597), .Y(n252) );
  MUX21X2_HVT U154 ( .A1(n479), .A2(n478), .S0(n319), .Y(n477) );
  INVX0_HVT U156 ( .A(n601), .Y(n373) );
  INVX1_HVT U157 ( .A(n348), .Y(n343) );
  INVX0_HVT U158 ( .A(n601), .Y(n245) );
  OA21X1_HVT U160 ( .A1(n359), .A2(n302), .A3(n601), .Y(n547) );
  MUX41X1_HVT U161 ( .A1(n436), .A3(n439), .A2(n437), .A4(n438), .S0(n243), 
        .S1(n280), .Y(n435) );
  IBUFFX16_HVT U165 ( .A(n279), .Y(n243) );
  IBUFFX16_HVT U167 ( .A(n317), .Y(n244) );
  INVX0_HVT U168 ( .A(n346), .Y(n269) );
  INVX0_HVT U169 ( .A(n346), .Y(n349) );
  MUX21X1_HVT U170 ( .A1(n333), .A2(n328), .S0(n322), .Y(n533) );
  INVX1_HVT U171 ( .A(n337), .Y(n412) );
  INVX2_HVT U173 ( .A(n348), .Y(n346) );
  INVX1_HVT U175 ( .A(n348), .Y(n345) );
  MUX21X2_HVT U176 ( .A1(n522), .A2(n529), .S0(n246), .Y(out[2]) );
  IBUFFX16_HVT U178 ( .A(n306), .Y(n246) );
  INVX0_HVT U180 ( .A(n362), .Y(n247) );
  MUX21X1_HVT U181 ( .A1(n305), .A2(n335), .S0(n287), .Y(n248) );
  NAND2X0_HVT U184 ( .A1(n560), .A2(in[7]), .Y(n251) );
  NAND2X0_HVT U186 ( .A1(n251), .A2(n250), .Y(out[0]) );
  IBUFFX2_HVT U187 ( .A(in[7]), .Y(n249) );
  INVX1_HVT U188 ( .A(n252), .Y(n253) );
  IBUFFX2_HVT U189 ( .A(n617), .Y(n292) );
  NAND2X0_HVT U190 ( .A1(n531), .A2(n254), .Y(n255) );
  NAND2X0_HVT U193 ( .A1(n532), .A2(n319), .Y(n256) );
  NAND2X0_HVT U196 ( .A1(n255), .A2(n256), .Y(n530) );
  IBUFFX2_HVT U197 ( .A(n319), .Y(n254) );
  MUX21X1_HVT U199 ( .A1(n533), .A2(n338), .S0(n286), .Y(n532) );
  MUX41X1_HVT U201 ( .A1(n452), .A3(n454), .A2(n450), .A4(n451), .S0(n257), 
        .S1(n258), .Y(n449) );
  IBUFFX16_HVT U202 ( .A(n279), .Y(n257) );
  MUX41X1_HVT U203 ( .A1(n481), .A3(n484), .A2(n483), .A4(n486), .S0(n266), 
        .S1(n260), .Y(n480) );
  IBUFFX16_HVT U204 ( .A(n329), .Y(n260) );
  IBUFFX16_HVT U205 ( .A(n320), .Y(n261) );
  MUX21X1_HVT U206 ( .A1(n411), .A2(n328), .S0(n262), .Y(n453) );
  NBUFFX2_HVT U208 ( .A(n343), .Y(n262) );
  NBUFFX2_HVT U209 ( .A(n346), .Y(n263) );
  IBUFFX2_HVT U210 ( .A(n348), .Y(n347) );
  INVX0_HVT U211 ( .A(n333), .Y(n277) );
  INVX2_HVT U212 ( .A(n305), .Y(n411) );
  NAND2X0_HVT U213 ( .A1(n343), .A2(n338), .Y(n616) );
  INVX0_HVT U214 ( .A(n585), .Y(n385) );
  INVX0_HVT U215 ( .A(n335), .Y(n278) );
  MUX21X1_HVT U216 ( .A1(n396), .A2(n356), .S0(n323), .Y(n548) );
  NAND2X0_HVT U217 ( .A1(n473), .A2(n284), .Y(n264) );
  INVX0_HVT U218 ( .A(in[5]), .Y(n332) );
  INVX1_HVT U219 ( .A(n322), .Y(n270) );
  INVX1_HVT U220 ( .A(n323), .Y(n273) );
  INVX0_HVT U221 ( .A(n331), .Y(n279) );
  INVX1_HVT U222 ( .A(n329), .Y(n331) );
  INVX1_HVT U223 ( .A(n288), .Y(n272) );
  INVX1_HVT U224 ( .A(in[1]), .Y(n329) );
  INVX1_HVT U225 ( .A(n354), .Y(n351) );
  INVX0_HVT U226 ( .A(n314), .Y(n284) );
  INVX1_HVT U227 ( .A(n314), .Y(n280) );
  MUX21X1_HVT U228 ( .A1(n328), .A2(n334), .S0(n269), .Y(n597) );
  NAND2X0_HVT U229 ( .A1(n474), .A2(n320), .Y(n265) );
  NAND2X0_HVT U230 ( .A1(n264), .A2(n265), .Y(n472) );
  MUX41X1_HVT U231 ( .A1(n472), .A3(n477), .A2(n471), .A4(n475), .S0(n266), 
        .S1(n272), .Y(n470) );
  IBUFFX2_HVT U232 ( .A(n591), .Y(n381) );
  MUX21X2_HVT U233 ( .A1(n375), .A2(n566), .S0(n313), .Y(n565) );
  INVX1_HVT U234 ( .A(n351), .Y(n271) );
  IBUFFX2_HVT U235 ( .A(n354), .Y(n268) );
  AO21X1_HVT U236 ( .A1(n269), .A2(n304), .A3(n271), .Y(n466) );
  INVX0_HVT U237 ( .A(n595), .Y(n378) );
  INVX1_HVT U238 ( .A(n348), .Y(n344) );
  MUX41X1_HVT U239 ( .A1(n542), .A3(n482), .A2(n403), .A4(n591), .S0(n280), 
        .S1(n271), .Y(n481) );
  MUX41X1_HVT U240 ( .A1(n512), .A3(n509), .A2(n510), .A4(n506), .S0(n332), 
        .S1(n272), .Y(n505) );
  NAND2X0_HVT U241 ( .A1(n596), .A2(n273), .Y(n274) );
  NAND2X0_HVT U242 ( .A1(n599), .A2(n268), .Y(n275) );
  NAND2X0_HVT U243 ( .A1(n274), .A2(n275), .Y(n460) );
  INVX0_HVT U244 ( .A(n276), .Y(n531) );
  INVX1_HVT U245 ( .A(n426), .Y(n395) );
  MUX21X1_HVT U246 ( .A1(n277), .A2(n587), .S0(n271), .Y(n276) );
  XNOR2X1_HVT U247 ( .A1(n278), .A2(n262), .Y(n574) );
  NAND2X0_HVT U248 ( .A1(n545), .A2(n281), .Y(n282) );
  NAND2X0_HVT U249 ( .A1(n538), .A2(n306), .Y(n283) );
  NAND2X0_HVT U250 ( .A1(n282), .A2(n283), .Y(out[1]) );
  INVX1_HVT U251 ( .A(n306), .Y(n281) );
  MUX21X2_HVT U252 ( .A1(n312), .A2(n574), .S0(n323), .Y(n438) );
  MUX21X2_HVT U253 ( .A1(n513), .A2(n514), .S0(n320), .Y(n512) );
  INVX0_HVT U254 ( .A(n615), .Y(n363) );
  MUX41X1_HVT U255 ( .A1(n584), .A3(n371), .A2(n372), .A4(n370), .S0(n284), 
        .S1(n271), .Y(n557) );
  IBUFFX2_HVT U256 ( .A(n354), .Y(n352) );
  INVX1_HVT U257 ( .A(n285), .Y(n571) );
  MUX21X1_HVT U258 ( .A1(n571), .A2(n570), .S0(n319), .Y(n569) );
  MUX21X1_HVT U259 ( .A1(n607), .A2(n595), .S0(n271), .Y(n285) );
  IBUFFX2_HVT U260 ( .A(n607), .Y(n368) );
  NBUFFX2_HVT U261 ( .A(n346), .Y(n286) );
  NBUFFX2_HVT U262 ( .A(n346), .Y(n287) );
  NBUFFX2_HVT U263 ( .A(n414), .Y(n327) );
  INVX1_HVT U264 ( .A(in[4]), .Y(n354) );
  INVX0_HVT U265 ( .A(n448), .Y(n301) );
  OA21X1_HVT U266 ( .A1(n379), .A2(n270), .A3(n562), .Y(n436) );
  INVX0_HVT U267 ( .A(n311), .Y(n300) );
  AO21X1_HVT U268 ( .A1(n334), .A2(n199), .A3(n302), .Y(n458) );
  OA21X1_HVT U269 ( .A1(n358), .A2(n271), .A3(n364), .Y(n473) );
  MUX41X1_HVT U270 ( .A1(n409), .A3(n388), .A2(n602), .A4(n599), .S0(n318), 
        .S1(n268), .Y(n483) );
  INVX1_HVT U271 ( .A(n279), .Y(n288) );
  INVX1_HVT U272 ( .A(in[3]), .Y(n410) );
  INVX1_HVT U273 ( .A(n321), .Y(n302) );
  INVX0_HVT U274 ( .A(in[7]), .Y(n306) );
  MUX41X1_HVT U275 ( .A1(n435), .A3(n429), .A2(n444), .A4(n441), .S0(n332), 
        .S1(n281), .Y(out[7]) );
  NAND2X0_HVT U276 ( .A1(n447), .A2(n288), .Y(n289) );
  NAND2X0_HVT U277 ( .A1(n445), .A2(n279), .Y(n290) );
  NAND2X0_HVT U278 ( .A1(n289), .A2(n290), .Y(n444) );
  MUX41X1_HVT U279 ( .A1(n528), .A3(n525), .A2(n526), .A4(n523), .S0(n332), 
        .S1(n279), .Y(n522) );
  MUX21X2_HVT U280 ( .A1(n548), .A2(n547), .S0(n320), .Y(n546) );
  MUX41X1_HVT U281 ( .A1(n400), .A3(n378), .A2(n609), .A4(n394), .S0(n284), 
        .S1(n271), .Y(n528) );
  INVX1_HVT U282 ( .A(n428), .Y(n393) );
  IBUFFX2_HVT U283 ( .A(n354), .Y(n353) );
  INVX1_HVT U284 ( .A(n291), .Y(n552) );
  MUX21X1_HVT U285 ( .A1(n409), .A2(n411), .S0(n345), .Y(n578) );
  MUX41X1_HVT U286 ( .A1(n587), .A3(n355), .A2(n304), .A4(n292), .S0(n284), 
        .S1(n273), .Y(n291) );
  MUX41X1_HVT U287 ( .A1(n577), .A3(n446), .A2(n355), .A4(n590), .S0(n284), 
        .S1(n270), .Y(n445) );
  MUX21X2_HVT U288 ( .A1(n502), .A2(n504), .S0(n331), .Y(n501) );
  MUX41X1_HVT U289 ( .A1(n605), .A3(n381), .A2(n604), .A4(n379), .S0(n280), 
        .S1(n270), .Y(n544) );
  NAND2X0_HVT U290 ( .A1(n456), .A2(n281), .Y(n293) );
  NAND2X0_HVT U291 ( .A1(n449), .A2(n306), .Y(n294) );
  NAND2X0_HVT U292 ( .A1(n293), .A2(n294), .Y(out[6]) );
  NBUFFX2_HVT U293 ( .A(n414), .Y(n328) );
  INVX0_HVT U294 ( .A(n299), .Y(n447) );
  MUX21X1_HVT U295 ( .A1(n333), .A2(n324), .S0(n344), .Y(n601) );
  XOR2X1_HVT U296 ( .A1(n304), .A2(n343), .Y(n585) );
  NBUFFX2_HVT U297 ( .A(n623), .Y(n304) );
  MUX21X1_HVT U298 ( .A1(n222), .A2(n298), .S0(n269), .Y(n297) );
  INVX1_HVT U299 ( .A(n578), .Y(n389) );
  MUX41X1_HVT U300 ( .A1(n389), .A3(n342), .A2(n301), .A4(n300), .S0(n280), 
        .S1(n302), .Y(n299) );
  MUX21X1_HVT U301 ( .A1(n411), .A2(n412), .S0(n344), .Y(n455) );
  NBUFFX2_HVT U302 ( .A(n622), .Y(n341) );
  MUX41X1_HVT U303 ( .A1(n455), .A3(n310), .A2(n307), .A4(n311), .S0(n280), 
        .S1(n271), .Y(n454) );
  AO21X2_HVT U304 ( .A1(n323), .A2(n363), .A3(n408), .Y(n478) );
  NBUFFX2_HVT U305 ( .A(n623), .Y(n305) );
  MUX21X2_HVT U306 ( .A1(n390), .A2(n310), .S0(n321), .Y(n431) );
  MUX21X2_HVT U307 ( .A1(n406), .A2(n237), .S0(n321), .Y(n479) );
  MUX21X2_HVT U308 ( .A1(n468), .A2(n469), .S0(n320), .Y(n465) );
  NBUFFX2_HVT U309 ( .A(n622), .Y(n340) );
  AND2X1_HVT U310 ( .A1(n617), .A2(n340), .Y(n307) );
  AND2X1_HVT U311 ( .A1(n340), .A2(n607), .Y(n308) );
  MUX21X1_HVT U312 ( .A1(n408), .A2(n327), .S0(n345), .Y(n426) );
  MUX21X1_HVT U313 ( .A1(n335), .A2(n338), .S0(n343), .Y(n464) );
  NAND2X0_HVT U314 ( .A1(n324), .A2(n326), .Y(n622) );
  MUX21X1_HVT U315 ( .A1(n411), .A2(n334), .S0(n240), .Y(n422) );
  MUX21X1_HVT U316 ( .A1(n326), .A2(n413), .S0(n263), .Y(n586) );
  MUX21X1_HVT U317 ( .A1(n327), .A2(n408), .S0(n262), .Y(n596) );
  MUX21X1_HVT U318 ( .A1(n408), .A2(n413), .S0(n345), .Y(n589) );
  MUX21X1_HVT U319 ( .A1(n325), .A2(n408), .S0(n240), .Y(n592) );
  MUX21X1_HVT U320 ( .A1(n326), .A2(n409), .S0(n240), .Y(n476) );
  MUX21X1_HVT U321 ( .A1(n413), .A2(n325), .S0(n263), .Y(n583) );
  MUX21X1_HVT U322 ( .A1(n405), .A2(n309), .S0(n319), .Y(n500) );
  MUX21X1_HVT U323 ( .A1(n413), .A2(n328), .S0(n344), .Y(n417) );
  MUX21X1_HVT U324 ( .A1(n589), .A2(n308), .S0(n320), .Y(n497) );
  MUX21X1_HVT U325 ( .A1(n326), .A2(n341), .S0(n241), .Y(n519) );
  XOR2X1_HVT U326 ( .A1(n337), .A2(n286), .Y(n575) );
  XOR2X1_HVT U327 ( .A1(n334), .A2(n344), .Y(n576) );
  MUX21X1_HVT U328 ( .A1(n334), .A2(n409), .S0(n343), .Y(n588) );
  MUX21X1_HVT U329 ( .A1(n324), .A2(n340), .S0(n241), .Y(n424) );
  INVX1_HVT U330 ( .A(n335), .Y(n409) );
  MUX21X1_HVT U331 ( .A1(n339), .A2(n340), .S0(n287), .Y(n604) );
  MUX21X1_HVT U332 ( .A1(n324), .A2(n412), .S0(n347), .Y(n579) );
  MUX21X1_HVT U333 ( .A1(n412), .A2(n324), .S0(n286), .Y(n425) );
  XNOR2X1_HVT U334 ( .A1(n341), .A2(n287), .Y(n309) );
  MUX21X1_HVT U335 ( .A1(n325), .A2(n327), .S0(n345), .Y(n577) );
  MUX21X1_HVT U336 ( .A1(n335), .A2(n341), .S0(n286), .Y(n416) );
  MUX21X1_HVT U337 ( .A1(n326), .A2(n334), .S0(n343), .Y(n582) );
  AND2X1_HVT U338 ( .A1(n263), .A2(n328), .Y(n310) );
  MUX21X1_HVT U339 ( .A1(n338), .A2(n325), .S0(n263), .Y(n603) );
  MUX21X1_HVT U340 ( .A1(n339), .A2(n327), .S0(n343), .Y(n503) );
  MUX21X1_HVT U341 ( .A1(n325), .A2(n338), .S0(n347), .Y(n419) );
  NBUFFX2_HVT U342 ( .A(n351), .Y(n321) );
  NBUFFX2_HVT U343 ( .A(n351), .Y(n323) );
  NBUFFX2_HVT U344 ( .A(n351), .Y(n322) );
  MUX21X1_HVT U345 ( .A1(n440), .A2(n397), .S0(n321), .Y(n439) );
  MUX21X1_HVT U346 ( .A1(n408), .A2(n412), .S0(n347), .Y(n572) );
  NBUFFX2_HVT U347 ( .A(n606), .Y(n333) );
  MUX21X1_HVT U348 ( .A1(n341), .A2(n336), .S0(n287), .Y(n482) );
  NBUFFX2_HVT U349 ( .A(n618), .Y(n335) );
  AND2X1_HVT U350 ( .A1(n412), .A2(n349), .Y(n311) );
  AND2X1_HVT U351 ( .A1(n339), .A2(n349), .Y(n312) );
  NBUFFX2_HVT U352 ( .A(n618), .Y(n336) );
  NBUFFX2_HVT U353 ( .A(n410), .Y(n325) );
  NBUFFX2_HVT U354 ( .A(n350), .Y(n318) );
  NBUFFX2_HVT U355 ( .A(n350), .Y(n320) );
  NBUFFX2_HVT U356 ( .A(n350), .Y(n319) );
  NBUFFX2_HVT U357 ( .A(in[2]), .Y(n316) );
  NBUFFX2_HVT U358 ( .A(n350), .Y(n314) );
  NBUFFX2_HVT U359 ( .A(n350), .Y(n317) );
  NBUFFX2_HVT U360 ( .A(n350), .Y(n315) );
  INVX1_HVT U361 ( .A(n329), .Y(n330) );
  MUX21X1_HVT U362 ( .A1(n492), .A2(n493), .S0(n288), .Y(n491) );
  MUX21X1_HVT U363 ( .A1(n488), .A2(n489), .S0(n331), .Y(n487) );
  MUX21X1_HVT U364 ( .A1(n412), .A2(n409), .S0(n262), .Y(n508) );
  NBUFFX2_HVT U365 ( .A(in[2]), .Y(n350) );
  MUX21X1_HVT U366 ( .A1(n408), .A2(n295), .S0(n240), .Y(n490) );
  XOR2X1_HVT U367 ( .A1(n241), .A2(n295), .Y(n573) );
  MUX21X1_HVT U368 ( .A1(n324), .A2(n295), .S0(n344), .Y(n418) );
  MUX21X1_HVT U369 ( .A1(n295), .A2(n411), .S0(n345), .Y(n598) );
  MUX21X1_HVT U370 ( .A1(n338), .A2(n295), .S0(n287), .Y(n423) );
  MUX21X1_HVT U371 ( .A1(n295), .A2(n339), .S0(n240), .Y(n427) );
  MUX21X1_HVT U372 ( .A1(n295), .A2(n342), .S0(n287), .Y(n605) );
  MUX21X1_HVT U373 ( .A1(n336), .A2(n295), .S0(n241), .Y(n593) );
  MUX21X1_HVT U374 ( .A1(n295), .A2(n409), .S0(n347), .Y(n428) );
  INVX0_HVT U375 ( .A(in[6]), .Y(n414) );
  NBUFFX2_HVT U376 ( .A(n623), .Y(n342) );
  MUX21X1_HVT U377 ( .A1(n411), .A2(n239), .S0(n241), .Y(n415) );
  MUX21X1_HVT U378 ( .A1(n304), .A2(n239), .S0(n263), .Y(n467) );
  MUX21X1_HVT U379 ( .A1(n239), .A2(n336), .S0(n287), .Y(n420) );
  MUX21X1_HVT U380 ( .A1(n239), .A2(n304), .S0(n286), .Y(n421) );
  MUX21X1_HVT U381 ( .A1(n336), .A2(n239), .S0(n347), .Y(n527) );
  MUX21X1_HVT U382 ( .A1(n328), .A2(n239), .S0(n241), .Y(n595) );
  NBUFFX2_HVT U383 ( .A(n606), .Y(n334) );
  NBUFFX2_HVT U384 ( .A(n621), .Y(n337) );
  NBUFFX2_HVT U385 ( .A(n621), .Y(n338) );
  NBUFFX2_HVT U386 ( .A(n621), .Y(n339) );
  INVX0_HVT U387 ( .A(n611), .Y(n355) );
  INVX0_HVT U388 ( .A(n590), .Y(n356) );
  INVX0_HVT U389 ( .A(n584), .Y(n357) );
  INVX0_HVT U390 ( .A(n524), .Y(n358) );
  INVX0_HVT U391 ( .A(n485), .Y(n359) );
  INVX0_HVT U392 ( .A(n616), .Y(n362) );
  INVX0_HVT U393 ( .A(n609), .Y(n364) );
  INVX0_HVT U394 ( .A(n614), .Y(n365) );
  INVX0_HVT U395 ( .A(n610), .Y(n366) );
  INVX0_HVT U396 ( .A(n608), .Y(n367) );
  INVX0_HVT U397 ( .A(n605), .Y(n369) );
  INVX0_HVT U398 ( .A(n604), .Y(n370) );
  INVX0_HVT U399 ( .A(n603), .Y(n371) );
  INVX0_HVT U400 ( .A(n602), .Y(n372) );
  INVX0_HVT U401 ( .A(n598), .Y(n375) );
  INVX0_HVT U402 ( .A(n593), .Y(n379) );
  INVX0_HVT U403 ( .A(n592), .Y(n380) );
  INVX0_HVT U404 ( .A(n589), .Y(n382) );
  INVX0_HVT U405 ( .A(n588), .Y(n383) );
  INVX0_HVT U406 ( .A(n583), .Y(n386) );
  INVX0_HVT U407 ( .A(n582), .Y(n387) );
  INVX0_HVT U408 ( .A(n579), .Y(n388) );
  INVX0_HVT U409 ( .A(n577), .Y(n390) );
  INVX0_HVT U410 ( .A(n613), .Y(n392) );
  INVX0_HVT U411 ( .A(n427), .Y(n394) );
  INVX0_HVT U412 ( .A(n425), .Y(n396) );
  INVX0_HVT U413 ( .A(n424), .Y(n397) );
  INVX0_HVT U414 ( .A(n423), .Y(n398) );
  INVX0_HVT U415 ( .A(n422), .Y(n399) );
  INVX0_HVT U416 ( .A(n421), .Y(n400) );
  INVX0_HVT U417 ( .A(n420), .Y(n401) );
  INVX0_HVT U418 ( .A(n419), .Y(n402) );
  INVX0_HVT U419 ( .A(n418), .Y(n403) );
  INVX0_HVT U420 ( .A(n467), .Y(n404) );
  INVX0_HVT U421 ( .A(n417), .Y(n405) );
  INVX0_HVT U422 ( .A(n415), .Y(n407) );
endmodule

