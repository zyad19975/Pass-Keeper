
module ram_dp_DATA_WIDTH4_ADDR_WIDTH4_25 ( clk, rst, write, a_addr, a_din, 
        b_din, b_dout );
  input [3:0] a_addr;
  input [3:0] a_din;
  input [3:0] b_din;
  output [15:0] b_dout;
  input clk, rst, write;
  wire   N17, N18, N19, N20, \mem[15][15] , \mem[15][14] , \mem[15][13] ,
         \mem[15][12] , \mem[15][11] , \mem[15][10] , \mem[15][9] ,
         \mem[15][8] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][15] ,
         \mem[14][14] , \mem[14][13] , \mem[14][12] , \mem[14][11] ,
         \mem[14][10] , \mem[14][9] , \mem[14][8] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][15] , \mem[13][14] , \mem[13][13] ,
         \mem[13][12] , \mem[13][11] , \mem[13][10] , \mem[13][9] ,
         \mem[13][8] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][15] ,
         \mem[12][14] , \mem[12][13] , \mem[12][12] , \mem[12][11] ,
         \mem[12][10] , \mem[12][9] , \mem[12][8] , \mem[12][7] , \mem[12][6] ,
         \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] , \mem[12][1] ,
         \mem[12][0] , \mem[11][15] , \mem[11][14] , \mem[11][13] ,
         \mem[11][12] , \mem[11][11] , \mem[11][10] , \mem[11][9] ,
         \mem[11][8] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][15] , \mem[9][14] , \mem[9][13] , \mem[9][12] ,
         \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] , \mem[9][7] ,
         \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] ,
         \mem[9][1] , \mem[9][0] , \mem[8][15] , \mem[8][14] , \mem[8][13] ,
         \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] , \mem[8][8] ,
         \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] , \mem[8][3] ,
         \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][15] , \mem[7][14] ,
         \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] ,
         \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][15] ,
         \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] ,
         \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][15] , \mem[3][14] , \mem[3][13] ,
         \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] ,
         \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] ,
         \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][15] ,
         \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N539, N540, N541, N542, N543, N544, N545, N546, N547,
         N548, N549, N550, N551, N552, N553, N554, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379;
  assign N17 = b_din[0];
  assign N18 = b_din[1];
  assign N19 = b_din[2];
  assign N20 = b_din[3];

  DFFNX1_HVT \b_dout_reg[15]  ( .D(N539), .CLK(clk), .Q(b_dout[15]) );
  DFFNX1_HVT \b_dout_reg[14]  ( .D(N540), .CLK(clk), .Q(b_dout[14]) );
  DFFNX1_HVT \b_dout_reg[13]  ( .D(N541), .CLK(clk), .Q(b_dout[13]) );
  DFFNX1_HVT \b_dout_reg[12]  ( .D(N542), .CLK(clk), .Q(b_dout[12]) );
  DFFNX1_HVT \b_dout_reg[11]  ( .D(N543), .CLK(clk), .Q(b_dout[11]) );
  DFFNX1_HVT \b_dout_reg[10]  ( .D(N544), .CLK(clk), .Q(b_dout[10]) );
  DFFNX1_HVT \b_dout_reg[9]  ( .D(N545), .CLK(clk), .Q(b_dout[9]) );
  DFFNX1_HVT \b_dout_reg[8]  ( .D(N546), .CLK(clk), .Q(b_dout[8]) );
  DFFNX1_HVT \b_dout_reg[7]  ( .D(N547), .CLK(clk), .Q(b_dout[7]) );
  DFFNX1_HVT \b_dout_reg[6]  ( .D(N548), .CLK(clk), .Q(b_dout[6]) );
  DFFNX1_HVT \b_dout_reg[5]  ( .D(N549), .CLK(clk), .Q(b_dout[5]) );
  DFFNX1_HVT \b_dout_reg[4]  ( .D(N550), .CLK(clk), .Q(b_dout[4]) );
  DFFNX1_HVT \b_dout_reg[3]  ( .D(N551), .CLK(clk), .Q(b_dout[3]) );
  DFFNX1_HVT \b_dout_reg[2]  ( .D(N552), .CLK(clk), .Q(b_dout[2]) );
  DFFNX1_HVT \b_dout_reg[1]  ( .D(N553), .CLK(clk), .Q(b_dout[1]) );
  DFFNX1_HVT \b_dout_reg[0]  ( .D(N554), .CLK(clk), .Q(b_dout[0]) );
  DFFNX1_HVT \mem_reg[15][15]  ( .D(n124), .CLK(clk), .Q(\mem[15][15] ) );
  DFFNX1_HVT \mem_reg[15][14]  ( .D(n125), .CLK(clk), .Q(\mem[15][14] ) );
  DFFNX1_HVT \mem_reg[15][13]  ( .D(n126), .CLK(clk), .Q(\mem[15][13] ) );
  DFFNX1_HVT \mem_reg[15][12]  ( .D(n127), .CLK(clk), .Q(\mem[15][12] ) );
  DFFNX1_HVT \mem_reg[15][11]  ( .D(n128), .CLK(clk), .Q(\mem[15][11] ) );
  DFFNX1_HVT \mem_reg[15][10]  ( .D(n129), .CLK(clk), .Q(\mem[15][10] ) );
  DFFNX1_HVT \mem_reg[15][9]  ( .D(n130), .CLK(clk), .Q(\mem[15][9] ) );
  DFFNX1_HVT \mem_reg[15][8]  ( .D(n131), .CLK(clk), .Q(\mem[15][8] ) );
  DFFNX1_HVT \mem_reg[15][7]  ( .D(n132), .CLK(clk), .Q(\mem[15][7] ) );
  DFFNX1_HVT \mem_reg[15][6]  ( .D(n133), .CLK(clk), .Q(\mem[15][6] ) );
  DFFNX1_HVT \mem_reg[15][5]  ( .D(n134), .CLK(clk), .Q(\mem[15][5] ) );
  DFFNX1_HVT \mem_reg[15][4]  ( .D(n135), .CLK(clk), .Q(\mem[15][4] ) );
  DFFNX1_HVT \mem_reg[15][3]  ( .D(n136), .CLK(clk), .Q(\mem[15][3] ) );
  DFFNX1_HVT \mem_reg[15][2]  ( .D(n137), .CLK(clk), .Q(\mem[15][2] ) );
  DFFNX1_HVT \mem_reg[15][1]  ( .D(n138), .CLK(clk), .Q(\mem[15][1] ) );
  DFFNX1_HVT \mem_reg[15][0]  ( .D(n139), .CLK(clk), .Q(\mem[15][0] ) );
  DFFNX1_HVT \mem_reg[14][15]  ( .D(n140), .CLK(clk), .Q(\mem[14][15] ) );
  DFFNX1_HVT \mem_reg[14][14]  ( .D(n141), .CLK(clk), .Q(\mem[14][14] ) );
  DFFNX1_HVT \mem_reg[14][13]  ( .D(n142), .CLK(clk), .Q(\mem[14][13] ) );
  DFFNX1_HVT \mem_reg[14][12]  ( .D(n143), .CLK(clk), .Q(\mem[14][12] ) );
  DFFNX1_HVT \mem_reg[14][11]  ( .D(n144), .CLK(clk), .Q(\mem[14][11] ) );
  DFFNX1_HVT \mem_reg[14][10]  ( .D(n145), .CLK(clk), .Q(\mem[14][10] ) );
  DFFNX1_HVT \mem_reg[14][9]  ( .D(n146), .CLK(clk), .Q(\mem[14][9] ) );
  DFFNX1_HVT \mem_reg[14][8]  ( .D(n147), .CLK(clk), .Q(\mem[14][8] ) );
  DFFNX1_HVT \mem_reg[14][7]  ( .D(n148), .CLK(clk), .Q(\mem[14][7] ) );
  DFFNX1_HVT \mem_reg[14][6]  ( .D(n149), .CLK(clk), .Q(\mem[14][6] ) );
  DFFNX1_HVT \mem_reg[14][5]  ( .D(n150), .CLK(clk), .Q(\mem[14][5] ) );
  DFFNX1_HVT \mem_reg[14][4]  ( .D(n151), .CLK(clk), .Q(\mem[14][4] ) );
  DFFNX1_HVT \mem_reg[14][3]  ( .D(n152), .CLK(clk), .Q(\mem[14][3] ) );
  DFFNX1_HVT \mem_reg[14][2]  ( .D(n153), .CLK(clk), .Q(\mem[14][2] ) );
  DFFNX1_HVT \mem_reg[14][1]  ( .D(n154), .CLK(clk), .Q(\mem[14][1] ) );
  DFFNX1_HVT \mem_reg[14][0]  ( .D(n155), .CLK(clk), .Q(\mem[14][0] ) );
  DFFNX1_HVT \mem_reg[13][15]  ( .D(n156), .CLK(clk), .Q(\mem[13][15] ) );
  DFFNX1_HVT \mem_reg[13][14]  ( .D(n157), .CLK(clk), .Q(\mem[13][14] ) );
  DFFNX1_HVT \mem_reg[13][13]  ( .D(n158), .CLK(clk), .Q(\mem[13][13] ) );
  DFFNX1_HVT \mem_reg[13][12]  ( .D(n159), .CLK(clk), .Q(\mem[13][12] ) );
  DFFNX1_HVT \mem_reg[13][11]  ( .D(n160), .CLK(clk), .Q(\mem[13][11] ) );
  DFFNX1_HVT \mem_reg[13][10]  ( .D(n161), .CLK(clk), .Q(\mem[13][10] ) );
  DFFNX1_HVT \mem_reg[13][9]  ( .D(n162), .CLK(clk), .Q(\mem[13][9] ) );
  DFFNX1_HVT \mem_reg[13][8]  ( .D(n163), .CLK(clk), .Q(\mem[13][8] ) );
  DFFNX1_HVT \mem_reg[13][7]  ( .D(n164), .CLK(clk), .Q(\mem[13][7] ) );
  DFFNX1_HVT \mem_reg[13][6]  ( .D(n165), .CLK(clk), .Q(\mem[13][6] ) );
  DFFNX1_HVT \mem_reg[13][5]  ( .D(n166), .CLK(clk), .Q(\mem[13][5] ) );
  DFFNX1_HVT \mem_reg[13][4]  ( .D(n167), .CLK(clk), .Q(\mem[13][4] ) );
  DFFNX1_HVT \mem_reg[13][3]  ( .D(n168), .CLK(clk), .Q(\mem[13][3] ) );
  DFFNX1_HVT \mem_reg[13][2]  ( .D(n169), .CLK(clk), .Q(\mem[13][2] ) );
  DFFNX1_HVT \mem_reg[13][1]  ( .D(n170), .CLK(clk), .Q(\mem[13][1] ) );
  DFFNX1_HVT \mem_reg[13][0]  ( .D(n171), .CLK(clk), .Q(\mem[13][0] ) );
  DFFNX1_HVT \mem_reg[12][15]  ( .D(n172), .CLK(clk), .Q(\mem[12][15] ) );
  DFFNX1_HVT \mem_reg[12][14]  ( .D(n173), .CLK(clk), .Q(\mem[12][14] ) );
  DFFNX1_HVT \mem_reg[12][13]  ( .D(n174), .CLK(clk), .Q(\mem[12][13] ) );
  DFFNX1_HVT \mem_reg[12][12]  ( .D(n175), .CLK(clk), .Q(\mem[12][12] ) );
  DFFNX1_HVT \mem_reg[12][11]  ( .D(n176), .CLK(clk), .Q(\mem[12][11] ) );
  DFFNX1_HVT \mem_reg[12][10]  ( .D(n177), .CLK(clk), .Q(\mem[12][10] ) );
  DFFNX1_HVT \mem_reg[12][9]  ( .D(n178), .CLK(clk), .Q(\mem[12][9] ) );
  DFFNX1_HVT \mem_reg[12][8]  ( .D(n179), .CLK(clk), .Q(\mem[12][8] ) );
  DFFNX1_HVT \mem_reg[12][7]  ( .D(n180), .CLK(clk), .Q(\mem[12][7] ) );
  DFFNX1_HVT \mem_reg[12][6]  ( .D(n181), .CLK(clk), .Q(\mem[12][6] ) );
  DFFNX1_HVT \mem_reg[12][5]  ( .D(n182), .CLK(clk), .Q(\mem[12][5] ) );
  DFFNX1_HVT \mem_reg[12][4]  ( .D(n183), .CLK(clk), .Q(\mem[12][4] ) );
  DFFNX1_HVT \mem_reg[12][3]  ( .D(n184), .CLK(clk), .Q(\mem[12][3] ) );
  DFFNX1_HVT \mem_reg[12][2]  ( .D(n185), .CLK(clk), .Q(\mem[12][2] ) );
  DFFNX1_HVT \mem_reg[12][1]  ( .D(n186), .CLK(clk), .Q(\mem[12][1] ) );
  DFFNX1_HVT \mem_reg[12][0]  ( .D(n187), .CLK(clk), .Q(\mem[12][0] ) );
  DFFNX1_HVT \mem_reg[11][15]  ( .D(n188), .CLK(clk), .Q(\mem[11][15] ) );
  DFFNX1_HVT \mem_reg[11][14]  ( .D(n189), .CLK(clk), .Q(\mem[11][14] ) );
  DFFNX1_HVT \mem_reg[11][13]  ( .D(n190), .CLK(clk), .Q(\mem[11][13] ) );
  DFFNX1_HVT \mem_reg[11][12]  ( .D(n191), .CLK(clk), .Q(\mem[11][12] ) );
  DFFNX1_HVT \mem_reg[11][11]  ( .D(n192), .CLK(clk), .Q(\mem[11][11] ) );
  DFFNX1_HVT \mem_reg[11][10]  ( .D(n193), .CLK(clk), .Q(\mem[11][10] ) );
  DFFNX1_HVT \mem_reg[11][9]  ( .D(n194), .CLK(clk), .Q(\mem[11][9] ) );
  DFFNX1_HVT \mem_reg[11][8]  ( .D(n195), .CLK(clk), .Q(\mem[11][8] ) );
  DFFNX1_HVT \mem_reg[11][7]  ( .D(n196), .CLK(clk), .Q(\mem[11][7] ) );
  DFFNX1_HVT \mem_reg[11][6]  ( .D(n197), .CLK(clk), .Q(\mem[11][6] ) );
  DFFNX1_HVT \mem_reg[11][5]  ( .D(n198), .CLK(clk), .Q(\mem[11][5] ) );
  DFFNX1_HVT \mem_reg[11][4]  ( .D(n199), .CLK(clk), .Q(\mem[11][4] ) );
  DFFNX1_HVT \mem_reg[11][3]  ( .D(n200), .CLK(clk), .Q(\mem[11][3] ) );
  DFFNX1_HVT \mem_reg[11][2]  ( .D(n201), .CLK(clk), .Q(\mem[11][2] ) );
  DFFNX1_HVT \mem_reg[11][1]  ( .D(n202), .CLK(clk), .Q(\mem[11][1] ) );
  DFFNX1_HVT \mem_reg[11][0]  ( .D(n203), .CLK(clk), .Q(\mem[11][0] ) );
  DFFNX1_HVT \mem_reg[10][15]  ( .D(n204), .CLK(clk), .Q(\mem[10][15] ) );
  DFFNX1_HVT \mem_reg[10][14]  ( .D(n205), .CLK(clk), .Q(\mem[10][14] ) );
  DFFNX1_HVT \mem_reg[10][13]  ( .D(n206), .CLK(clk), .Q(\mem[10][13] ) );
  DFFNX1_HVT \mem_reg[10][12]  ( .D(n207), .CLK(clk), .Q(\mem[10][12] ) );
  DFFNX1_HVT \mem_reg[10][11]  ( .D(n208), .CLK(clk), .Q(\mem[10][11] ) );
  DFFNX1_HVT \mem_reg[10][10]  ( .D(n209), .CLK(clk), .Q(\mem[10][10] ) );
  DFFNX1_HVT \mem_reg[10][9]  ( .D(n210), .CLK(clk), .Q(\mem[10][9] ) );
  DFFNX1_HVT \mem_reg[10][8]  ( .D(n211), .CLK(clk), .Q(\mem[10][8] ) );
  DFFNX1_HVT \mem_reg[10][7]  ( .D(n212), .CLK(clk), .Q(\mem[10][7] ) );
  DFFNX1_HVT \mem_reg[10][6]  ( .D(n213), .CLK(clk), .Q(\mem[10][6] ) );
  DFFNX1_HVT \mem_reg[10][5]  ( .D(n214), .CLK(clk), .Q(\mem[10][5] ) );
  DFFNX1_HVT \mem_reg[10][4]  ( .D(n215), .CLK(clk), .Q(\mem[10][4] ) );
  DFFNX1_HVT \mem_reg[10][3]  ( .D(n216), .CLK(clk), .Q(\mem[10][3] ) );
  DFFNX1_HVT \mem_reg[10][2]  ( .D(n217), .CLK(clk), .Q(\mem[10][2] ) );
  DFFNX1_HVT \mem_reg[10][1]  ( .D(n218), .CLK(clk), .Q(\mem[10][1] ) );
  DFFNX1_HVT \mem_reg[10][0]  ( .D(n219), .CLK(clk), .Q(\mem[10][0] ) );
  DFFNX1_HVT \mem_reg[9][15]  ( .D(n220), .CLK(clk), .Q(\mem[9][15] ) );
  DFFNX1_HVT \mem_reg[9][14]  ( .D(n221), .CLK(clk), .Q(\mem[9][14] ) );
  DFFNX1_HVT \mem_reg[9][13]  ( .D(n222), .CLK(clk), .Q(\mem[9][13] ) );
  DFFNX1_HVT \mem_reg[9][12]  ( .D(n223), .CLK(clk), .Q(\mem[9][12] ) );
  DFFNX1_HVT \mem_reg[9][11]  ( .D(n224), .CLK(clk), .Q(\mem[9][11] ) );
  DFFNX1_HVT \mem_reg[9][10]  ( .D(n225), .CLK(clk), .Q(\mem[9][10] ) );
  DFFNX1_HVT \mem_reg[9][9]  ( .D(n226), .CLK(clk), .Q(\mem[9][9] ) );
  DFFNX1_HVT \mem_reg[9][8]  ( .D(n227), .CLK(clk), .Q(\mem[9][8] ) );
  DFFNX1_HVT \mem_reg[9][7]  ( .D(n228), .CLK(clk), .Q(\mem[9][7] ) );
  DFFNX1_HVT \mem_reg[9][6]  ( .D(n229), .CLK(clk), .Q(\mem[9][6] ) );
  DFFNX1_HVT \mem_reg[9][5]  ( .D(n230), .CLK(clk), .Q(\mem[9][5] ) );
  DFFNX1_HVT \mem_reg[9][4]  ( .D(n231), .CLK(clk), .Q(\mem[9][4] ) );
  DFFNX1_HVT \mem_reg[9][3]  ( .D(n232), .CLK(clk), .Q(\mem[9][3] ) );
  DFFNX1_HVT \mem_reg[9][2]  ( .D(n233), .CLK(clk), .Q(\mem[9][2] ) );
  DFFNX1_HVT \mem_reg[9][1]  ( .D(n234), .CLK(clk), .Q(\mem[9][1] ) );
  DFFNX1_HVT \mem_reg[9][0]  ( .D(n235), .CLK(clk), .Q(\mem[9][0] ) );
  DFFNX1_HVT \mem_reg[8][15]  ( .D(n236), .CLK(clk), .Q(\mem[8][15] ) );
  DFFNX1_HVT \mem_reg[8][14]  ( .D(n237), .CLK(clk), .Q(\mem[8][14] ) );
  DFFNX1_HVT \mem_reg[8][13]  ( .D(n238), .CLK(clk), .Q(\mem[8][13] ) );
  DFFNX1_HVT \mem_reg[8][12]  ( .D(n239), .CLK(clk), .Q(\mem[8][12] ) );
  DFFNX1_HVT \mem_reg[8][11]  ( .D(n240), .CLK(clk), .Q(\mem[8][11] ) );
  DFFNX1_HVT \mem_reg[8][10]  ( .D(n241), .CLK(clk), .Q(\mem[8][10] ) );
  DFFNX1_HVT \mem_reg[8][9]  ( .D(n242), .CLK(clk), .Q(\mem[8][9] ) );
  DFFNX1_HVT \mem_reg[8][8]  ( .D(n243), .CLK(clk), .Q(\mem[8][8] ) );
  DFFNX1_HVT \mem_reg[8][7]  ( .D(n244), .CLK(clk), .Q(\mem[8][7] ) );
  DFFNX1_HVT \mem_reg[8][6]  ( .D(n245), .CLK(clk), .Q(\mem[8][6] ) );
  DFFNX1_HVT \mem_reg[8][5]  ( .D(n246), .CLK(clk), .Q(\mem[8][5] ) );
  DFFNX1_HVT \mem_reg[8][4]  ( .D(n247), .CLK(clk), .Q(\mem[8][4] ) );
  DFFNX1_HVT \mem_reg[8][3]  ( .D(n248), .CLK(clk), .Q(\mem[8][3] ) );
  DFFNX1_HVT \mem_reg[8][2]  ( .D(n249), .CLK(clk), .Q(\mem[8][2] ) );
  DFFNX1_HVT \mem_reg[8][1]  ( .D(n250), .CLK(clk), .Q(\mem[8][1] ) );
  DFFNX1_HVT \mem_reg[8][0]  ( .D(n251), .CLK(clk), .Q(\mem[8][0] ) );
  DFFNX1_HVT \mem_reg[7][15]  ( .D(n252), .CLK(clk), .Q(\mem[7][15] ) );
  DFFNX1_HVT \mem_reg[7][14]  ( .D(n253), .CLK(clk), .Q(\mem[7][14] ) );
  DFFNX1_HVT \mem_reg[7][13]  ( .D(n254), .CLK(clk), .Q(\mem[7][13] ) );
  DFFNX1_HVT \mem_reg[7][12]  ( .D(n255), .CLK(clk), .Q(\mem[7][12] ) );
  DFFNX1_HVT \mem_reg[7][11]  ( .D(n256), .CLK(clk), .Q(\mem[7][11] ) );
  DFFNX1_HVT \mem_reg[7][10]  ( .D(n257), .CLK(clk), .Q(\mem[7][10] ) );
  DFFNX1_HVT \mem_reg[7][9]  ( .D(n258), .CLK(clk), .Q(\mem[7][9] ) );
  DFFNX1_HVT \mem_reg[7][8]  ( .D(n259), .CLK(clk), .Q(\mem[7][8] ) );
  DFFNX1_HVT \mem_reg[7][7]  ( .D(n260), .CLK(clk), .Q(\mem[7][7] ) );
  DFFNX1_HVT \mem_reg[7][6]  ( .D(n261), .CLK(clk), .Q(\mem[7][6] ) );
  DFFNX1_HVT \mem_reg[7][5]  ( .D(n262), .CLK(clk), .Q(\mem[7][5] ) );
  DFFNX1_HVT \mem_reg[7][4]  ( .D(n263), .CLK(clk), .Q(\mem[7][4] ) );
  DFFNX1_HVT \mem_reg[7][3]  ( .D(n264), .CLK(clk), .Q(\mem[7][3] ) );
  DFFNX1_HVT \mem_reg[7][2]  ( .D(n265), .CLK(clk), .Q(\mem[7][2] ) );
  DFFNX1_HVT \mem_reg[7][1]  ( .D(n266), .CLK(clk), .Q(\mem[7][1] ) );
  DFFNX1_HVT \mem_reg[7][0]  ( .D(n267), .CLK(clk), .Q(\mem[7][0] ) );
  DFFNX1_HVT \mem_reg[6][15]  ( .D(n268), .CLK(clk), .Q(\mem[6][15] ) );
  DFFNX1_HVT \mem_reg[6][14]  ( .D(n269), .CLK(clk), .Q(\mem[6][14] ) );
  DFFNX1_HVT \mem_reg[6][13]  ( .D(n270), .CLK(clk), .Q(\mem[6][13] ) );
  DFFNX1_HVT \mem_reg[6][12]  ( .D(n271), .CLK(clk), .Q(\mem[6][12] ) );
  DFFNX1_HVT \mem_reg[6][11]  ( .D(n272), .CLK(clk), .Q(\mem[6][11] ) );
  DFFNX1_HVT \mem_reg[6][10]  ( .D(n273), .CLK(clk), .Q(\mem[6][10] ) );
  DFFNX1_HVT \mem_reg[6][9]  ( .D(n274), .CLK(clk), .Q(\mem[6][9] ) );
  DFFNX1_HVT \mem_reg[6][8]  ( .D(n275), .CLK(clk), .Q(\mem[6][8] ) );
  DFFNX1_HVT \mem_reg[6][7]  ( .D(n276), .CLK(clk), .Q(\mem[6][7] ) );
  DFFNX1_HVT \mem_reg[6][6]  ( .D(n277), .CLK(clk), .Q(\mem[6][6] ) );
  DFFNX1_HVT \mem_reg[6][5]  ( .D(n278), .CLK(clk), .Q(\mem[6][5] ) );
  DFFNX1_HVT \mem_reg[6][4]  ( .D(n279), .CLK(clk), .Q(\mem[6][4] ) );
  DFFNX1_HVT \mem_reg[6][3]  ( .D(n280), .CLK(clk), .Q(\mem[6][3] ) );
  DFFNX1_HVT \mem_reg[6][2]  ( .D(n281), .CLK(clk), .Q(\mem[6][2] ) );
  DFFNX1_HVT \mem_reg[6][1]  ( .D(n282), .CLK(clk), .Q(\mem[6][1] ) );
  DFFNX1_HVT \mem_reg[6][0]  ( .D(n283), .CLK(clk), .Q(\mem[6][0] ) );
  DFFNX1_HVT \mem_reg[5][15]  ( .D(n284), .CLK(clk), .Q(\mem[5][15] ) );
  DFFNX1_HVT \mem_reg[5][14]  ( .D(n285), .CLK(clk), .Q(\mem[5][14] ) );
  DFFNX1_HVT \mem_reg[5][13]  ( .D(n286), .CLK(clk), .Q(\mem[5][13] ) );
  DFFNX1_HVT \mem_reg[5][12]  ( .D(n287), .CLK(clk), .Q(\mem[5][12] ) );
  DFFNX1_HVT \mem_reg[5][11]  ( .D(n288), .CLK(clk), .Q(\mem[5][11] ) );
  DFFNX1_HVT \mem_reg[5][10]  ( .D(n289), .CLK(clk), .Q(\mem[5][10] ) );
  DFFNX1_HVT \mem_reg[5][9]  ( .D(n290), .CLK(clk), .Q(\mem[5][9] ) );
  DFFNX1_HVT \mem_reg[5][8]  ( .D(n291), .CLK(clk), .Q(\mem[5][8] ) );
  DFFNX1_HVT \mem_reg[5][7]  ( .D(n292), .CLK(clk), .Q(\mem[5][7] ) );
  DFFNX1_HVT \mem_reg[5][6]  ( .D(n293), .CLK(clk), .Q(\mem[5][6] ) );
  DFFNX1_HVT \mem_reg[5][5]  ( .D(n294), .CLK(clk), .Q(\mem[5][5] ) );
  DFFNX1_HVT \mem_reg[5][4]  ( .D(n295), .CLK(clk), .Q(\mem[5][4] ) );
  DFFNX1_HVT \mem_reg[5][3]  ( .D(n296), .CLK(clk), .Q(\mem[5][3] ) );
  DFFNX1_HVT \mem_reg[5][2]  ( .D(n297), .CLK(clk), .Q(\mem[5][2] ) );
  DFFNX1_HVT \mem_reg[5][1]  ( .D(n298), .CLK(clk), .Q(\mem[5][1] ) );
  DFFNX1_HVT \mem_reg[5][0]  ( .D(n299), .CLK(clk), .Q(\mem[5][0] ) );
  DFFNX1_HVT \mem_reg[4][15]  ( .D(n300), .CLK(clk), .Q(\mem[4][15] ) );
  DFFNX1_HVT \mem_reg[4][14]  ( .D(n301), .CLK(clk), .Q(\mem[4][14] ) );
  DFFNX1_HVT \mem_reg[4][13]  ( .D(n302), .CLK(clk), .Q(\mem[4][13] ) );
  DFFNX1_HVT \mem_reg[4][12]  ( .D(n303), .CLK(clk), .Q(\mem[4][12] ) );
  DFFNX1_HVT \mem_reg[4][11]  ( .D(n304), .CLK(clk), .Q(\mem[4][11] ) );
  DFFNX1_HVT \mem_reg[4][10]  ( .D(n305), .CLK(clk), .Q(\mem[4][10] ) );
  DFFNX1_HVT \mem_reg[4][9]  ( .D(n306), .CLK(clk), .Q(\mem[4][9] ) );
  DFFNX1_HVT \mem_reg[4][8]  ( .D(n307), .CLK(clk), .Q(\mem[4][8] ) );
  DFFNX1_HVT \mem_reg[4][7]  ( .D(n308), .CLK(clk), .Q(\mem[4][7] ) );
  DFFNX1_HVT \mem_reg[4][6]  ( .D(n309), .CLK(clk), .Q(\mem[4][6] ) );
  DFFNX1_HVT \mem_reg[4][5]  ( .D(n310), .CLK(clk), .Q(\mem[4][5] ) );
  DFFNX1_HVT \mem_reg[4][4]  ( .D(n311), .CLK(clk), .Q(\mem[4][4] ) );
  DFFNX1_HVT \mem_reg[4][3]  ( .D(n312), .CLK(clk), .Q(\mem[4][3] ) );
  DFFNX1_HVT \mem_reg[4][2]  ( .D(n313), .CLK(clk), .Q(\mem[4][2] ) );
  DFFNX1_HVT \mem_reg[4][1]  ( .D(n314), .CLK(clk), .Q(\mem[4][1] ) );
  DFFNX1_HVT \mem_reg[4][0]  ( .D(n315), .CLK(clk), .Q(\mem[4][0] ) );
  DFFNX1_HVT \mem_reg[3][15]  ( .D(n316), .CLK(clk), .Q(\mem[3][15] ) );
  DFFNX1_HVT \mem_reg[3][14]  ( .D(n317), .CLK(clk), .Q(\mem[3][14] ) );
  DFFNX1_HVT \mem_reg[3][13]  ( .D(n318), .CLK(clk), .Q(\mem[3][13] ) );
  DFFNX1_HVT \mem_reg[3][12]  ( .D(n319), .CLK(clk), .Q(\mem[3][12] ) );
  DFFNX1_HVT \mem_reg[3][11]  ( .D(n320), .CLK(clk), .Q(\mem[3][11] ) );
  DFFNX1_HVT \mem_reg[3][10]  ( .D(n321), .CLK(clk), .Q(\mem[3][10] ) );
  DFFNX1_HVT \mem_reg[3][9]  ( .D(n322), .CLK(clk), .Q(\mem[3][9] ) );
  DFFNX1_HVT \mem_reg[3][8]  ( .D(n323), .CLK(clk), .Q(\mem[3][8] ) );
  DFFNX1_HVT \mem_reg[3][7]  ( .D(n324), .CLK(clk), .Q(\mem[3][7] ) );
  DFFNX1_HVT \mem_reg[3][6]  ( .D(n325), .CLK(clk), .Q(\mem[3][6] ) );
  DFFNX1_HVT \mem_reg[3][5]  ( .D(n326), .CLK(clk), .Q(\mem[3][5] ) );
  DFFNX1_HVT \mem_reg[3][4]  ( .D(n327), .CLK(clk), .Q(\mem[3][4] ) );
  DFFNX1_HVT \mem_reg[3][3]  ( .D(n328), .CLK(clk), .Q(\mem[3][3] ) );
  DFFNX1_HVT \mem_reg[3][2]  ( .D(n329), .CLK(clk), .Q(\mem[3][2] ) );
  DFFNX1_HVT \mem_reg[3][1]  ( .D(n330), .CLK(clk), .Q(\mem[3][1] ) );
  DFFNX1_HVT \mem_reg[3][0]  ( .D(n331), .CLK(clk), .Q(\mem[3][0] ) );
  DFFNX1_HVT \mem_reg[2][15]  ( .D(n332), .CLK(clk), .Q(\mem[2][15] ) );
  DFFNX1_HVT \mem_reg[2][14]  ( .D(n333), .CLK(clk), .Q(\mem[2][14] ) );
  DFFNX1_HVT \mem_reg[2][13]  ( .D(n334), .CLK(clk), .Q(\mem[2][13] ) );
  DFFNX1_HVT \mem_reg[2][12]  ( .D(n335), .CLK(clk), .Q(\mem[2][12] ) );
  DFFNX1_HVT \mem_reg[2][11]  ( .D(n336), .CLK(clk), .Q(\mem[2][11] ) );
  DFFNX1_HVT \mem_reg[2][10]  ( .D(n337), .CLK(clk), .Q(\mem[2][10] ) );
  DFFNX1_HVT \mem_reg[2][9]  ( .D(n338), .CLK(clk), .Q(\mem[2][9] ) );
  DFFNX1_HVT \mem_reg[2][8]  ( .D(n339), .CLK(clk), .Q(\mem[2][8] ) );
  DFFNX1_HVT \mem_reg[2][7]  ( .D(n340), .CLK(clk), .Q(\mem[2][7] ) );
  DFFNX1_HVT \mem_reg[2][6]  ( .D(n341), .CLK(clk), .Q(\mem[2][6] ) );
  DFFNX1_HVT \mem_reg[2][5]  ( .D(n342), .CLK(clk), .Q(\mem[2][5] ) );
  DFFNX1_HVT \mem_reg[2][4]  ( .D(n343), .CLK(clk), .Q(\mem[2][4] ) );
  DFFNX1_HVT \mem_reg[2][3]  ( .D(n344), .CLK(clk), .Q(\mem[2][3] ) );
  DFFNX1_HVT \mem_reg[2][2]  ( .D(n345), .CLK(clk), .Q(\mem[2][2] ) );
  DFFNX1_HVT \mem_reg[2][1]  ( .D(n346), .CLK(clk), .Q(\mem[2][1] ) );
  DFFNX1_HVT \mem_reg[2][0]  ( .D(n347), .CLK(clk), .Q(\mem[2][0] ) );
  DFFNX1_HVT \mem_reg[1][15]  ( .D(n348), .CLK(clk), .Q(\mem[1][15] ) );
  DFFNX1_HVT \mem_reg[1][14]  ( .D(n349), .CLK(clk), .Q(\mem[1][14] ) );
  DFFNX1_HVT \mem_reg[1][13]  ( .D(n350), .CLK(clk), .Q(\mem[1][13] ) );
  DFFNX1_HVT \mem_reg[1][12]  ( .D(n351), .CLK(clk), .Q(\mem[1][12] ) );
  DFFNX1_HVT \mem_reg[1][11]  ( .D(n352), .CLK(clk), .Q(\mem[1][11] ) );
  DFFNX1_HVT \mem_reg[1][10]  ( .D(n353), .CLK(clk), .Q(\mem[1][10] ) );
  DFFNX1_HVT \mem_reg[1][9]  ( .D(n354), .CLK(clk), .Q(\mem[1][9] ) );
  DFFNX1_HVT \mem_reg[1][8]  ( .D(n355), .CLK(clk), .Q(\mem[1][8] ) );
  DFFNX1_HVT \mem_reg[1][7]  ( .D(n356), .CLK(clk), .Q(\mem[1][7] ) );
  DFFNX1_HVT \mem_reg[1][6]  ( .D(n357), .CLK(clk), .Q(\mem[1][6] ) );
  DFFNX1_HVT \mem_reg[1][5]  ( .D(n358), .CLK(clk), .Q(\mem[1][5] ) );
  DFFNX1_HVT \mem_reg[1][4]  ( .D(n359), .CLK(clk), .Q(\mem[1][4] ) );
  DFFNX1_HVT \mem_reg[1][3]  ( .D(n360), .CLK(clk), .Q(\mem[1][3] ) );
  DFFNX1_HVT \mem_reg[1][2]  ( .D(n361), .CLK(clk), .Q(\mem[1][2] ) );
  DFFNX1_HVT \mem_reg[1][1]  ( .D(n362), .CLK(clk), .Q(\mem[1][1] ) );
  DFFNX1_HVT \mem_reg[1][0]  ( .D(n363), .CLK(clk), .Q(\mem[1][0] ) );
  DFFNX1_HVT \mem_reg[0][15]  ( .D(n364), .CLK(clk), .Q(\mem[0][15] ) );
  DFFNX1_HVT \mem_reg[0][14]  ( .D(n365), .CLK(clk), .Q(\mem[0][14] ) );
  DFFNX1_HVT \mem_reg[0][13]  ( .D(n366), .CLK(clk), .Q(\mem[0][13] ) );
  DFFNX1_HVT \mem_reg[0][12]  ( .D(n367), .CLK(clk), .Q(\mem[0][12] ) );
  DFFNX1_HVT \mem_reg[0][11]  ( .D(n368), .CLK(clk), .Q(\mem[0][11] ) );
  DFFNX1_HVT \mem_reg[0][10]  ( .D(n369), .CLK(clk), .Q(\mem[0][10] ) );
  DFFNX1_HVT \mem_reg[0][9]  ( .D(n370), .CLK(clk), .Q(\mem[0][9] ) );
  DFFNX1_HVT \mem_reg[0][8]  ( .D(n371), .CLK(clk), .Q(\mem[0][8] ) );
  DFFNX1_HVT \mem_reg[0][7]  ( .D(n372), .CLK(clk), .Q(\mem[0][7] ) );
  DFFNX1_HVT \mem_reg[0][6]  ( .D(n373), .CLK(clk), .Q(\mem[0][6] ) );
  DFFNX1_HVT \mem_reg[0][5]  ( .D(n374), .CLK(clk), .Q(\mem[0][5] ) );
  DFFNX1_HVT \mem_reg[0][4]  ( .D(n375), .CLK(clk), .Q(\mem[0][4] ) );
  DFFNX1_HVT \mem_reg[0][3]  ( .D(n376), .CLK(clk), .Q(\mem[0][3] ) );
  DFFNX1_HVT \mem_reg[0][2]  ( .D(n377), .CLK(clk), .Q(\mem[0][2] ) );
  DFFNX1_HVT \mem_reg[0][1]  ( .D(n378), .CLK(clk), .Q(\mem[0][1] ) );
  DFFNX1_HVT \mem_reg[0][0]  ( .D(n379), .CLK(clk), .Q(\mem[0][0] ) );
  MUX41X1_HVT U3 ( .A1(\mem[12][0] ), .A3(\mem[14][0] ), .A2(\mem[13][0] ), 
        .A4(\mem[15][0] ), .S0(N18), .S1(N17), .Y(n1) );
  MUX41X1_HVT U4 ( .A1(\mem[8][0] ), .A3(\mem[10][0] ), .A2(\mem[9][0] ), .A4(
        \mem[11][0] ), .S0(N18), .S1(N17), .Y(n2) );
  MUX41X1_HVT U5 ( .A1(\mem[4][0] ), .A3(\mem[6][0] ), .A2(\mem[5][0] ), .A4(
        \mem[7][0] ), .S0(N18), .S1(N17), .Y(n3) );
  MUX41X1_HVT U6 ( .A1(\mem[0][0] ), .A3(\mem[2][0] ), .A2(\mem[1][0] ), .A4(
        \mem[3][0] ), .S0(N18), .S1(N17), .Y(n4) );
  MUX41X1_HVT U7 ( .A1(n4), .A3(n2), .A2(n3), .A4(n1), .S0(N20), .S1(N19), .Y(
        N554) );
  MUX41X1_HVT U8 ( .A1(\mem[12][1] ), .A3(\mem[14][1] ), .A2(\mem[13][1] ), 
        .A4(\mem[15][1] ), .S0(N18), .S1(N17), .Y(n5) );
  MUX41X1_HVT U9 ( .A1(\mem[8][1] ), .A3(\mem[10][1] ), .A2(\mem[9][1] ), .A4(
        \mem[11][1] ), .S0(N18), .S1(N17), .Y(n6) );
  MUX41X1_HVT U10 ( .A1(\mem[4][1] ), .A3(\mem[6][1] ), .A2(\mem[5][1] ), .A4(
        \mem[7][1] ), .S0(N18), .S1(N17), .Y(n7) );
  MUX41X1_HVT U11 ( .A1(\mem[0][1] ), .A3(\mem[2][1] ), .A2(\mem[1][1] ), .A4(
        \mem[3][1] ), .S0(N18), .S1(N17), .Y(n8) );
  MUX41X1_HVT U12 ( .A1(n8), .A3(n6), .A2(n7), .A4(n5), .S0(N20), .S1(N19), 
        .Y(N553) );
  MUX41X1_HVT U13 ( .A1(\mem[12][2] ), .A3(\mem[14][2] ), .A2(\mem[13][2] ), 
        .A4(\mem[15][2] ), .S0(N18), .S1(N17), .Y(n9) );
  MUX41X1_HVT U14 ( .A1(\mem[8][2] ), .A3(\mem[10][2] ), .A2(\mem[9][2] ), 
        .A4(\mem[11][2] ), .S0(N18), .S1(N17), .Y(n10) );
  MUX41X1_HVT U15 ( .A1(\mem[4][2] ), .A3(\mem[6][2] ), .A2(\mem[5][2] ), .A4(
        \mem[7][2] ), .S0(N18), .S1(N17), .Y(n11) );
  MUX41X1_HVT U16 ( .A1(\mem[0][2] ), .A3(\mem[2][2] ), .A2(\mem[1][2] ), .A4(
        \mem[3][2] ), .S0(N18), .S1(N17), .Y(n12) );
  MUX41X1_HVT U17 ( .A1(n12), .A3(n10), .A2(n11), .A4(n9), .S0(N20), .S1(N19), 
        .Y(N552) );
  MUX41X1_HVT U18 ( .A1(\mem[12][3] ), .A3(\mem[14][3] ), .A2(\mem[13][3] ), 
        .A4(\mem[15][3] ), .S0(N18), .S1(N17), .Y(n13) );
  MUX41X1_HVT U19 ( .A1(\mem[8][3] ), .A3(\mem[10][3] ), .A2(\mem[9][3] ), 
        .A4(\mem[11][3] ), .S0(N18), .S1(N17), .Y(n14) );
  MUX41X1_HVT U20 ( .A1(\mem[4][3] ), .A3(\mem[6][3] ), .A2(\mem[5][3] ), .A4(
        \mem[7][3] ), .S0(N18), .S1(N17), .Y(n15) );
  MUX41X1_HVT U21 ( .A1(\mem[0][3] ), .A3(\mem[2][3] ), .A2(\mem[1][3] ), .A4(
        \mem[3][3] ), .S0(N18), .S1(N17), .Y(n16) );
  MUX41X1_HVT U22 ( .A1(n16), .A3(n14), .A2(n15), .A4(n13), .S0(N20), .S1(N19), 
        .Y(N551) );
  MUX41X1_HVT U23 ( .A1(\mem[12][4] ), .A3(\mem[14][4] ), .A2(\mem[13][4] ), 
        .A4(\mem[15][4] ), .S0(N18), .S1(N17), .Y(n17) );
  MUX41X1_HVT U24 ( .A1(\mem[8][4] ), .A3(\mem[10][4] ), .A2(\mem[9][4] ), 
        .A4(\mem[11][4] ), .S0(N18), .S1(N17), .Y(n18) );
  MUX41X1_HVT U25 ( .A1(\mem[4][4] ), .A3(\mem[6][4] ), .A2(\mem[5][4] ), .A4(
        \mem[7][4] ), .S0(N18), .S1(N17), .Y(n19) );
  MUX41X1_HVT U26 ( .A1(\mem[0][4] ), .A3(\mem[2][4] ), .A2(\mem[1][4] ), .A4(
        \mem[3][4] ), .S0(N18), .S1(N17), .Y(n20) );
  MUX41X1_HVT U27 ( .A1(n20), .A3(n18), .A2(n19), .A4(n17), .S0(N20), .S1(N19), 
        .Y(N550) );
  MUX41X1_HVT U28 ( .A1(\mem[12][5] ), .A3(\mem[14][5] ), .A2(\mem[13][5] ), 
        .A4(\mem[15][5] ), .S0(N18), .S1(N17), .Y(n21) );
  MUX41X1_HVT U29 ( .A1(\mem[8][5] ), .A3(\mem[10][5] ), .A2(\mem[9][5] ), 
        .A4(\mem[11][5] ), .S0(N18), .S1(N17), .Y(n22) );
  MUX41X1_HVT U30 ( .A1(\mem[4][5] ), .A3(\mem[6][5] ), .A2(\mem[5][5] ), .A4(
        \mem[7][5] ), .S0(N18), .S1(N17), .Y(n23) );
  MUX41X1_HVT U31 ( .A1(\mem[0][5] ), .A3(\mem[2][5] ), .A2(\mem[1][5] ), .A4(
        \mem[3][5] ), .S0(N18), .S1(N17), .Y(n24) );
  MUX41X1_HVT U32 ( .A1(n24), .A3(n22), .A2(n23), .A4(n21), .S0(N20), .S1(N19), 
        .Y(N549) );
  MUX41X1_HVT U33 ( .A1(\mem[12][6] ), .A3(\mem[14][6] ), .A2(\mem[13][6] ), 
        .A4(\mem[15][6] ), .S0(N18), .S1(N17), .Y(n25) );
  MUX41X1_HVT U34 ( .A1(\mem[8][6] ), .A3(\mem[10][6] ), .A2(\mem[9][6] ), 
        .A4(\mem[11][6] ), .S0(N18), .S1(N17), .Y(n26) );
  MUX41X1_HVT U35 ( .A1(\mem[4][6] ), .A3(\mem[6][6] ), .A2(\mem[5][6] ), .A4(
        \mem[7][6] ), .S0(N18), .S1(N17), .Y(n27) );
  MUX41X1_HVT U36 ( .A1(\mem[0][6] ), .A3(\mem[2][6] ), .A2(\mem[1][6] ), .A4(
        \mem[3][6] ), .S0(N18), .S1(N17), .Y(n28) );
  MUX41X1_HVT U37 ( .A1(n28), .A3(n26), .A2(n27), .A4(n25), .S0(N20), .S1(N19), 
        .Y(N548) );
  MUX41X1_HVT U38 ( .A1(\mem[12][7] ), .A3(\mem[14][7] ), .A2(\mem[13][7] ), 
        .A4(\mem[15][7] ), .S0(N18), .S1(N17), .Y(n29) );
  MUX41X1_HVT U39 ( .A1(\mem[8][7] ), .A3(\mem[10][7] ), .A2(\mem[9][7] ), 
        .A4(\mem[11][7] ), .S0(N18), .S1(N17), .Y(n30) );
  MUX41X1_HVT U40 ( .A1(\mem[4][7] ), .A3(\mem[6][7] ), .A2(\mem[5][7] ), .A4(
        \mem[7][7] ), .S0(N18), .S1(N17), .Y(n31) );
  MUX41X1_HVT U41 ( .A1(\mem[0][7] ), .A3(\mem[2][7] ), .A2(\mem[1][7] ), .A4(
        \mem[3][7] ), .S0(N18), .S1(N17), .Y(n32) );
  MUX41X1_HVT U42 ( .A1(n32), .A3(n30), .A2(n31), .A4(n29), .S0(N20), .S1(N19), 
        .Y(N547) );
  MUX41X1_HVT U43 ( .A1(\mem[12][8] ), .A3(\mem[14][8] ), .A2(\mem[13][8] ), 
        .A4(\mem[15][8] ), .S0(N18), .S1(N17), .Y(n33) );
  MUX41X1_HVT U44 ( .A1(\mem[8][8] ), .A3(\mem[10][8] ), .A2(\mem[9][8] ), 
        .A4(\mem[11][8] ), .S0(N18), .S1(N17), .Y(n34) );
  MUX41X1_HVT U45 ( .A1(\mem[4][8] ), .A3(\mem[6][8] ), .A2(\mem[5][8] ), .A4(
        \mem[7][8] ), .S0(N18), .S1(N17), .Y(n35) );
  MUX41X1_HVT U46 ( .A1(\mem[0][8] ), .A3(\mem[2][8] ), .A2(\mem[1][8] ), .A4(
        \mem[3][8] ), .S0(N18), .S1(N17), .Y(n36) );
  MUX41X1_HVT U47 ( .A1(n36), .A3(n34), .A2(n35), .A4(n33), .S0(N20), .S1(N19), 
        .Y(N546) );
  MUX41X1_HVT U48 ( .A1(\mem[12][9] ), .A3(\mem[14][9] ), .A2(\mem[13][9] ), 
        .A4(\mem[15][9] ), .S0(N18), .S1(N17), .Y(n37) );
  MUX41X1_HVT U49 ( .A1(\mem[8][9] ), .A3(\mem[10][9] ), .A2(\mem[9][9] ), 
        .A4(\mem[11][9] ), .S0(N18), .S1(N17), .Y(n38) );
  MUX41X1_HVT U50 ( .A1(\mem[4][9] ), .A3(\mem[6][9] ), .A2(\mem[5][9] ), .A4(
        \mem[7][9] ), .S0(N18), .S1(N17), .Y(n39) );
  MUX41X1_HVT U51 ( .A1(\mem[0][9] ), .A3(\mem[2][9] ), .A2(\mem[1][9] ), .A4(
        \mem[3][9] ), .S0(N18), .S1(N17), .Y(n40) );
  MUX41X1_HVT U52 ( .A1(n40), .A3(n38), .A2(n39), .A4(n37), .S0(N20), .S1(N19), 
        .Y(N545) );
  MUX41X1_HVT U53 ( .A1(\mem[12][10] ), .A3(\mem[14][10] ), .A2(\mem[13][10] ), 
        .A4(\mem[15][10] ), .S0(N18), .S1(N17), .Y(n41) );
  MUX41X1_HVT U54 ( .A1(\mem[8][10] ), .A3(\mem[10][10] ), .A2(\mem[9][10] ), 
        .A4(\mem[11][10] ), .S0(N18), .S1(N17), .Y(n42) );
  MUX41X1_HVT U55 ( .A1(\mem[4][10] ), .A3(\mem[6][10] ), .A2(\mem[5][10] ), 
        .A4(\mem[7][10] ), .S0(N18), .S1(N17), .Y(n43) );
  MUX41X1_HVT U56 ( .A1(\mem[0][10] ), .A3(\mem[2][10] ), .A2(\mem[1][10] ), 
        .A4(\mem[3][10] ), .S0(N18), .S1(N17), .Y(n44) );
  MUX41X1_HVT U57 ( .A1(n44), .A3(n42), .A2(n43), .A4(n41), .S0(N20), .S1(N19), 
        .Y(N544) );
  MUX41X1_HVT U58 ( .A1(\mem[12][11] ), .A3(\mem[14][11] ), .A2(\mem[13][11] ), 
        .A4(\mem[15][11] ), .S0(N18), .S1(N17), .Y(n45) );
  MUX41X1_HVT U59 ( .A1(\mem[8][11] ), .A3(\mem[10][11] ), .A2(\mem[9][11] ), 
        .A4(\mem[11][11] ), .S0(N18), .S1(N17), .Y(n46) );
  MUX41X1_HVT U60 ( .A1(\mem[4][11] ), .A3(\mem[6][11] ), .A2(\mem[5][11] ), 
        .A4(\mem[7][11] ), .S0(N18), .S1(N17), .Y(n47) );
  MUX41X1_HVT U61 ( .A1(\mem[0][11] ), .A3(\mem[2][11] ), .A2(\mem[1][11] ), 
        .A4(\mem[3][11] ), .S0(N18), .S1(N17), .Y(n48) );
  MUX41X1_HVT U62 ( .A1(n48), .A3(n46), .A2(n47), .A4(n45), .S0(N20), .S1(N19), 
        .Y(N543) );
  MUX41X1_HVT U63 ( .A1(\mem[12][12] ), .A3(\mem[14][12] ), .A2(\mem[13][12] ), 
        .A4(\mem[15][12] ), .S0(N18), .S1(N17), .Y(n49) );
  MUX41X1_HVT U64 ( .A1(\mem[8][12] ), .A3(\mem[10][12] ), .A2(\mem[9][12] ), 
        .A4(\mem[11][12] ), .S0(N18), .S1(N17), .Y(n50) );
  MUX41X1_HVT U65 ( .A1(\mem[4][12] ), .A3(\mem[6][12] ), .A2(\mem[5][12] ), 
        .A4(\mem[7][12] ), .S0(N18), .S1(N17), .Y(n51) );
  MUX41X1_HVT U66 ( .A1(\mem[0][12] ), .A3(\mem[2][12] ), .A2(\mem[1][12] ), 
        .A4(\mem[3][12] ), .S0(N18), .S1(N17), .Y(n52) );
  MUX41X1_HVT U67 ( .A1(n52), .A3(n50), .A2(n51), .A4(n49), .S0(N20), .S1(N19), 
        .Y(N542) );
  MUX41X1_HVT U68 ( .A1(\mem[12][13] ), .A3(\mem[14][13] ), .A2(\mem[13][13] ), 
        .A4(\mem[15][13] ), .S0(N18), .S1(N17), .Y(n53) );
  MUX41X1_HVT U69 ( .A1(\mem[8][13] ), .A3(\mem[10][13] ), .A2(\mem[9][13] ), 
        .A4(\mem[11][13] ), .S0(N18), .S1(N17), .Y(n54) );
  MUX41X1_HVT U70 ( .A1(\mem[4][13] ), .A3(\mem[6][13] ), .A2(\mem[5][13] ), 
        .A4(\mem[7][13] ), .S0(N18), .S1(N17), .Y(n55) );
  MUX41X1_HVT U71 ( .A1(\mem[0][13] ), .A3(\mem[2][13] ), .A2(\mem[1][13] ), 
        .A4(\mem[3][13] ), .S0(N18), .S1(N17), .Y(n56) );
  MUX41X1_HVT U72 ( .A1(n56), .A3(n54), .A2(n55), .A4(n53), .S0(N20), .S1(N19), 
        .Y(N541) );
  MUX41X1_HVT U73 ( .A1(\mem[12][14] ), .A3(\mem[14][14] ), .A2(\mem[13][14] ), 
        .A4(\mem[15][14] ), .S0(N18), .S1(N17), .Y(n57) );
  MUX41X1_HVT U74 ( .A1(\mem[8][14] ), .A3(\mem[10][14] ), .A2(\mem[9][14] ), 
        .A4(\mem[11][14] ), .S0(N18), .S1(N17), .Y(n58) );
  MUX41X1_HVT U75 ( .A1(\mem[4][14] ), .A3(\mem[6][14] ), .A2(\mem[5][14] ), 
        .A4(\mem[7][14] ), .S0(N18), .S1(N17), .Y(n59) );
  MUX41X1_HVT U76 ( .A1(\mem[0][14] ), .A3(\mem[2][14] ), .A2(\mem[1][14] ), 
        .A4(\mem[3][14] ), .S0(N18), .S1(N17), .Y(n60) );
  MUX41X1_HVT U77 ( .A1(n60), .A3(n58), .A2(n59), .A4(n57), .S0(N20), .S1(N19), 
        .Y(N540) );
  MUX41X1_HVT U78 ( .A1(\mem[12][15] ), .A3(\mem[14][15] ), .A2(\mem[13][15] ), 
        .A4(\mem[15][15] ), .S0(N18), .S1(N17), .Y(n61) );
  MUX41X1_HVT U79 ( .A1(\mem[8][15] ), .A3(\mem[10][15] ), .A2(\mem[9][15] ), 
        .A4(\mem[11][15] ), .S0(N18), .S1(N17), .Y(n62) );
  MUX41X1_HVT U80 ( .A1(\mem[4][15] ), .A3(\mem[6][15] ), .A2(\mem[5][15] ), 
        .A4(\mem[7][15] ), .S0(N18), .S1(N17), .Y(n63) );
  MUX41X1_HVT U81 ( .A1(\mem[0][15] ), .A3(\mem[2][15] ), .A2(\mem[1][15] ), 
        .A4(\mem[3][15] ), .S0(N18), .S1(N17), .Y(n64) );
  MUX41X1_HVT U82 ( .A1(n64), .A3(n62), .A2(n63), .A4(n61), .S0(N20), .S1(N19), 
        .Y(N539) );
  AO22X1_HVT U83 ( .A1(\mem[15][15] ), .A2(n65), .A3(n66), .A4(n67), .Y(n124)
         );
  AO22X1_HVT U84 ( .A1(\mem[15][14] ), .A2(n65), .A3(n68), .A4(n66), .Y(n125)
         );
  AO22X1_HVT U85 ( .A1(\mem[15][13] ), .A2(n65), .A3(n69), .A4(n66), .Y(n126)
         );
  AO22X1_HVT U86 ( .A1(\mem[15][12] ), .A2(n65), .A3(n70), .A4(n66), .Y(n127)
         );
  AO22X1_HVT U87 ( .A1(\mem[15][11] ), .A2(n65), .A3(n71), .A4(n66), .Y(n128)
         );
  AO22X1_HVT U88 ( .A1(\mem[15][10] ), .A2(n65), .A3(n72), .A4(n66), .Y(n129)
         );
  AO22X1_HVT U89 ( .A1(\mem[15][9] ), .A2(n65), .A3(n73), .A4(n66), .Y(n130)
         );
  AO22X1_HVT U90 ( .A1(\mem[15][8] ), .A2(n65), .A3(n74), .A4(n66), .Y(n131)
         );
  AO22X1_HVT U91 ( .A1(\mem[15][7] ), .A2(n65), .A3(n75), .A4(n66), .Y(n132)
         );
  AO22X1_HVT U92 ( .A1(\mem[15][6] ), .A2(n65), .A3(n76), .A4(n66), .Y(n133)
         );
  AO22X1_HVT U93 ( .A1(\mem[15][5] ), .A2(n65), .A3(n77), .A4(n66), .Y(n134)
         );
  AO22X1_HVT U94 ( .A1(\mem[15][4] ), .A2(n65), .A3(n78), .A4(n66), .Y(n135)
         );
  AO22X1_HVT U95 ( .A1(\mem[15][3] ), .A2(n65), .A3(n79), .A4(n66), .Y(n136)
         );
  AO22X1_HVT U96 ( .A1(\mem[15][2] ), .A2(n65), .A3(n80), .A4(n66), .Y(n137)
         );
  AO22X1_HVT U97 ( .A1(\mem[15][1] ), .A2(n65), .A3(n81), .A4(n66), .Y(n138)
         );
  AO22X1_HVT U98 ( .A1(\mem[15][0] ), .A2(n65), .A3(n82), .A4(n66), .Y(n139)
         );
  AND2X1_HVT U99 ( .A1(n83), .A2(n84), .Y(n66) );
  AO22X1_HVT U100 ( .A1(\mem[14][15] ), .A2(n65), .A3(n85), .A4(n67), .Y(n140)
         );
  AO22X1_HVT U101 ( .A1(\mem[14][14] ), .A2(n65), .A3(n85), .A4(n68), .Y(n141)
         );
  AO22X1_HVT U102 ( .A1(\mem[14][13] ), .A2(n65), .A3(n85), .A4(n69), .Y(n142)
         );
  AO22X1_HVT U103 ( .A1(\mem[14][12] ), .A2(n65), .A3(n85), .A4(n70), .Y(n143)
         );
  AO22X1_HVT U104 ( .A1(\mem[14][11] ), .A2(n65), .A3(n85), .A4(n71), .Y(n144)
         );
  AO22X1_HVT U105 ( .A1(\mem[14][10] ), .A2(n65), .A3(n85), .A4(n72), .Y(n145)
         );
  AO22X1_HVT U106 ( .A1(\mem[14][9] ), .A2(n65), .A3(n85), .A4(n73), .Y(n146)
         );
  AO22X1_HVT U107 ( .A1(\mem[14][8] ), .A2(n65), .A3(n85), .A4(n74), .Y(n147)
         );
  AO22X1_HVT U108 ( .A1(\mem[14][7] ), .A2(n65), .A3(n85), .A4(n75), .Y(n148)
         );
  AO22X1_HVT U109 ( .A1(\mem[14][6] ), .A2(n65), .A3(n85), .A4(n76), .Y(n149)
         );
  AO22X1_HVT U110 ( .A1(\mem[14][5] ), .A2(n65), .A3(n85), .A4(n77), .Y(n150)
         );
  AO22X1_HVT U111 ( .A1(\mem[14][4] ), .A2(n65), .A3(n85), .A4(n78), .Y(n151)
         );
  AO22X1_HVT U112 ( .A1(\mem[14][3] ), .A2(n65), .A3(n85), .A4(n79), .Y(n152)
         );
  AO22X1_HVT U113 ( .A1(\mem[14][2] ), .A2(n65), .A3(n85), .A4(n80), .Y(n153)
         );
  AO22X1_HVT U114 ( .A1(\mem[14][1] ), .A2(n65), .A3(n85), .A4(n81), .Y(n154)
         );
  AO22X1_HVT U115 ( .A1(\mem[14][0] ), .A2(n65), .A3(n85), .A4(n82), .Y(n155)
         );
  AND2X1_HVT U116 ( .A1(n86), .A2(n83), .Y(n85) );
  AO22X1_HVT U117 ( .A1(\mem[13][15] ), .A2(n65), .A3(n87), .A4(n67), .Y(n156)
         );
  AO22X1_HVT U118 ( .A1(\mem[13][14] ), .A2(n65), .A3(n87), .A4(n68), .Y(n157)
         );
  AO22X1_HVT U119 ( .A1(\mem[13][13] ), .A2(n65), .A3(n87), .A4(n69), .Y(n158)
         );
  AO22X1_HVT U120 ( .A1(\mem[13][12] ), .A2(n65), .A3(n87), .A4(n70), .Y(n159)
         );
  AO22X1_HVT U121 ( .A1(\mem[13][11] ), .A2(n65), .A3(n87), .A4(n71), .Y(n160)
         );
  AO22X1_HVT U122 ( .A1(\mem[13][10] ), .A2(n65), .A3(n87), .A4(n72), .Y(n161)
         );
  AO22X1_HVT U123 ( .A1(\mem[13][9] ), .A2(n65), .A3(n87), .A4(n73), .Y(n162)
         );
  AO22X1_HVT U124 ( .A1(\mem[13][8] ), .A2(n65), .A3(n87), .A4(n74), .Y(n163)
         );
  AO22X1_HVT U125 ( .A1(\mem[13][7] ), .A2(n65), .A3(n87), .A4(n75), .Y(n164)
         );
  AO22X1_HVT U126 ( .A1(\mem[13][6] ), .A2(n65), .A3(n87), .A4(n76), .Y(n165)
         );
  AO22X1_HVT U127 ( .A1(\mem[13][5] ), .A2(n65), .A3(n87), .A4(n77), .Y(n166)
         );
  AO22X1_HVT U128 ( .A1(\mem[13][4] ), .A2(n65), .A3(n87), .A4(n78), .Y(n167)
         );
  AO22X1_HVT U129 ( .A1(\mem[13][3] ), .A2(n65), .A3(n87), .A4(n79), .Y(n168)
         );
  AO22X1_HVT U130 ( .A1(\mem[13][2] ), .A2(n65), .A3(n87), .A4(n80), .Y(n169)
         );
  AO22X1_HVT U131 ( .A1(\mem[13][1] ), .A2(n65), .A3(n87), .A4(n81), .Y(n170)
         );
  AO22X1_HVT U132 ( .A1(\mem[13][0] ), .A2(n65), .A3(n87), .A4(n82), .Y(n171)
         );
  AND2X1_HVT U133 ( .A1(n88), .A2(n84), .Y(n87) );
  AO22X1_HVT U134 ( .A1(\mem[12][15] ), .A2(n65), .A3(n89), .A4(n67), .Y(n172)
         );
  AO22X1_HVT U135 ( .A1(\mem[12][14] ), .A2(n65), .A3(n89), .A4(n68), .Y(n173)
         );
  AO22X1_HVT U136 ( .A1(\mem[12][13] ), .A2(n65), .A3(n89), .A4(n69), .Y(n174)
         );
  AO22X1_HVT U137 ( .A1(\mem[12][12] ), .A2(n65), .A3(n89), .A4(n70), .Y(n175)
         );
  AO22X1_HVT U138 ( .A1(\mem[12][11] ), .A2(n65), .A3(n89), .A4(n71), .Y(n176)
         );
  AO22X1_HVT U139 ( .A1(\mem[12][10] ), .A2(n65), .A3(n89), .A4(n72), .Y(n177)
         );
  AO22X1_HVT U140 ( .A1(\mem[12][9] ), .A2(n65), .A3(n89), .A4(n73), .Y(n178)
         );
  AO22X1_HVT U141 ( .A1(\mem[12][8] ), .A2(n65), .A3(n89), .A4(n74), .Y(n179)
         );
  AO22X1_HVT U142 ( .A1(\mem[12][7] ), .A2(n65), .A3(n89), .A4(n75), .Y(n180)
         );
  AO22X1_HVT U143 ( .A1(\mem[12][6] ), .A2(n65), .A3(n89), .A4(n76), .Y(n181)
         );
  AO22X1_HVT U144 ( .A1(\mem[12][5] ), .A2(n65), .A3(n89), .A4(n77), .Y(n182)
         );
  AO22X1_HVT U145 ( .A1(\mem[12][4] ), .A2(n65), .A3(n89), .A4(n78), .Y(n183)
         );
  AO22X1_HVT U146 ( .A1(\mem[12][3] ), .A2(n65), .A3(n89), .A4(n79), .Y(n184)
         );
  AO22X1_HVT U147 ( .A1(\mem[12][2] ), .A2(n65), .A3(n89), .A4(n80), .Y(n185)
         );
  AO22X1_HVT U148 ( .A1(\mem[12][1] ), .A2(n65), .A3(n89), .A4(n81), .Y(n186)
         );
  AO22X1_HVT U149 ( .A1(\mem[12][0] ), .A2(n65), .A3(n89), .A4(n82), .Y(n187)
         );
  AND2X1_HVT U150 ( .A1(n88), .A2(n86), .Y(n89) );
  AO22X1_HVT U151 ( .A1(\mem[11][15] ), .A2(n65), .A3(n90), .A4(n67), .Y(n188)
         );
  AO22X1_HVT U152 ( .A1(\mem[11][14] ), .A2(n65), .A3(n90), .A4(n68), .Y(n189)
         );
  AO22X1_HVT U153 ( .A1(\mem[11][13] ), .A2(n65), .A3(n90), .A4(n69), .Y(n190)
         );
  AO22X1_HVT U154 ( .A1(\mem[11][12] ), .A2(n65), .A3(n90), .A4(n70), .Y(n191)
         );
  AO22X1_HVT U155 ( .A1(\mem[11][11] ), .A2(n65), .A3(n90), .A4(n71), .Y(n192)
         );
  AO22X1_HVT U156 ( .A1(\mem[11][10] ), .A2(n65), .A3(n90), .A4(n72), .Y(n193)
         );
  AO22X1_HVT U157 ( .A1(\mem[11][9] ), .A2(n65), .A3(n90), .A4(n73), .Y(n194)
         );
  AO22X1_HVT U158 ( .A1(\mem[11][8] ), .A2(n65), .A3(n90), .A4(n74), .Y(n195)
         );
  AO22X1_HVT U159 ( .A1(\mem[11][7] ), .A2(n65), .A3(n90), .A4(n75), .Y(n196)
         );
  AO22X1_HVT U160 ( .A1(\mem[11][6] ), .A2(n65), .A3(n90), .A4(n76), .Y(n197)
         );
  AO22X1_HVT U161 ( .A1(\mem[11][5] ), .A2(n65), .A3(n90), .A4(n77), .Y(n198)
         );
  AO22X1_HVT U162 ( .A1(\mem[11][4] ), .A2(n65), .A3(n90), .A4(n78), .Y(n199)
         );
  AO22X1_HVT U163 ( .A1(\mem[11][3] ), .A2(n65), .A3(n90), .A4(n79), .Y(n200)
         );
  AO22X1_HVT U164 ( .A1(\mem[11][2] ), .A2(n65), .A3(n90), .A4(n80), .Y(n201)
         );
  AO22X1_HVT U165 ( .A1(\mem[11][1] ), .A2(n65), .A3(n90), .A4(n81), .Y(n202)
         );
  AO22X1_HVT U166 ( .A1(\mem[11][0] ), .A2(n65), .A3(n90), .A4(n82), .Y(n203)
         );
  AND2X1_HVT U167 ( .A1(n91), .A2(n84), .Y(n90) );
  AO22X1_HVT U168 ( .A1(\mem[10][15] ), .A2(n65), .A3(n92), .A4(n67), .Y(n204)
         );
  AO22X1_HVT U169 ( .A1(\mem[10][14] ), .A2(n65), .A3(n92), .A4(n68), .Y(n205)
         );
  AO22X1_HVT U170 ( .A1(\mem[10][13] ), .A2(n65), .A3(n92), .A4(n69), .Y(n206)
         );
  AO22X1_HVT U171 ( .A1(\mem[10][12] ), .A2(n65), .A3(n92), .A4(n70), .Y(n207)
         );
  AO22X1_HVT U172 ( .A1(\mem[10][11] ), .A2(n65), .A3(n92), .A4(n71), .Y(n208)
         );
  AO22X1_HVT U173 ( .A1(\mem[10][10] ), .A2(n65), .A3(n92), .A4(n72), .Y(n209)
         );
  AO22X1_HVT U174 ( .A1(\mem[10][9] ), .A2(n65), .A3(n92), .A4(n73), .Y(n210)
         );
  AO22X1_HVT U175 ( .A1(\mem[10][8] ), .A2(n65), .A3(n92), .A4(n74), .Y(n211)
         );
  AO22X1_HVT U176 ( .A1(\mem[10][7] ), .A2(n65), .A3(n92), .A4(n75), .Y(n212)
         );
  AO22X1_HVT U177 ( .A1(\mem[10][6] ), .A2(n65), .A3(n92), .A4(n76), .Y(n213)
         );
  AO22X1_HVT U178 ( .A1(\mem[10][5] ), .A2(n65), .A3(n92), .A4(n77), .Y(n214)
         );
  AO22X1_HVT U179 ( .A1(\mem[10][4] ), .A2(n65), .A3(n92), .A4(n78), .Y(n215)
         );
  AO22X1_HVT U180 ( .A1(\mem[10][3] ), .A2(n65), .A3(n92), .A4(n79), .Y(n216)
         );
  AO22X1_HVT U181 ( .A1(\mem[10][2] ), .A2(n65), .A3(n92), .A4(n80), .Y(n217)
         );
  AO22X1_HVT U182 ( .A1(\mem[10][1] ), .A2(n65), .A3(n92), .A4(n81), .Y(n218)
         );
  AO22X1_HVT U183 ( .A1(\mem[10][0] ), .A2(n65), .A3(n92), .A4(n82), .Y(n219)
         );
  AND2X1_HVT U184 ( .A1(n91), .A2(n86), .Y(n92) );
  AO22X1_HVT U185 ( .A1(\mem[9][15] ), .A2(n65), .A3(n93), .A4(n67), .Y(n220)
         );
  AO22X1_HVT U186 ( .A1(\mem[9][14] ), .A2(n65), .A3(n93), .A4(n68), .Y(n221)
         );
  AO22X1_HVT U187 ( .A1(\mem[9][13] ), .A2(n65), .A3(n93), .A4(n69), .Y(n222)
         );
  AO22X1_HVT U188 ( .A1(\mem[9][12] ), .A2(n65), .A3(n93), .A4(n70), .Y(n223)
         );
  AO22X1_HVT U189 ( .A1(\mem[9][11] ), .A2(n65), .A3(n93), .A4(n71), .Y(n224)
         );
  AO22X1_HVT U190 ( .A1(\mem[9][10] ), .A2(n65), .A3(n93), .A4(n72), .Y(n225)
         );
  AO22X1_HVT U191 ( .A1(\mem[9][9] ), .A2(n65), .A3(n93), .A4(n73), .Y(n226)
         );
  AO22X1_HVT U192 ( .A1(\mem[9][8] ), .A2(n65), .A3(n93), .A4(n74), .Y(n227)
         );
  AO22X1_HVT U193 ( .A1(\mem[9][7] ), .A2(n65), .A3(n93), .A4(n75), .Y(n228)
         );
  AO22X1_HVT U194 ( .A1(\mem[9][6] ), .A2(n65), .A3(n93), .A4(n76), .Y(n229)
         );
  AO22X1_HVT U195 ( .A1(\mem[9][5] ), .A2(n65), .A3(n93), .A4(n77), .Y(n230)
         );
  AO22X1_HVT U196 ( .A1(\mem[9][4] ), .A2(n65), .A3(n93), .A4(n78), .Y(n231)
         );
  AO22X1_HVT U197 ( .A1(\mem[9][3] ), .A2(n65), .A3(n93), .A4(n79), .Y(n232)
         );
  AO22X1_HVT U198 ( .A1(\mem[9][2] ), .A2(n65), .A3(n93), .A4(n80), .Y(n233)
         );
  AO22X1_HVT U199 ( .A1(\mem[9][1] ), .A2(n65), .A3(n93), .A4(n81), .Y(n234)
         );
  AO22X1_HVT U200 ( .A1(\mem[9][0] ), .A2(n65), .A3(n93), .A4(n82), .Y(n235)
         );
  AND2X1_HVT U201 ( .A1(n94), .A2(n84), .Y(n93) );
  AND2X1_HVT U202 ( .A1(a_din[0]), .A2(n95), .Y(n84) );
  AO22X1_HVT U203 ( .A1(\mem[8][15] ), .A2(n65), .A3(n96), .A4(n67), .Y(n236)
         );
  AO22X1_HVT U204 ( .A1(\mem[8][14] ), .A2(n65), .A3(n96), .A4(n68), .Y(n237)
         );
  AO22X1_HVT U205 ( .A1(\mem[8][13] ), .A2(n65), .A3(n96), .A4(n69), .Y(n238)
         );
  AO22X1_HVT U206 ( .A1(\mem[8][12] ), .A2(n65), .A3(n96), .A4(n70), .Y(n239)
         );
  AO22X1_HVT U207 ( .A1(\mem[8][11] ), .A2(n65), .A3(n96), .A4(n71), .Y(n240)
         );
  AO22X1_HVT U208 ( .A1(\mem[8][10] ), .A2(n65), .A3(n96), .A4(n72), .Y(n241)
         );
  AO22X1_HVT U209 ( .A1(\mem[8][9] ), .A2(n65), .A3(n96), .A4(n73), .Y(n242)
         );
  AO22X1_HVT U210 ( .A1(\mem[8][8] ), .A2(n65), .A3(n96), .A4(n74), .Y(n243)
         );
  AO22X1_HVT U211 ( .A1(\mem[8][7] ), .A2(n65), .A3(n96), .A4(n75), .Y(n244)
         );
  AO22X1_HVT U212 ( .A1(\mem[8][6] ), .A2(n65), .A3(n96), .A4(n76), .Y(n245)
         );
  AO22X1_HVT U213 ( .A1(\mem[8][5] ), .A2(n65), .A3(n96), .A4(n77), .Y(n246)
         );
  AO22X1_HVT U214 ( .A1(\mem[8][4] ), .A2(n65), .A3(n96), .A4(n78), .Y(n247)
         );
  AO22X1_HVT U215 ( .A1(\mem[8][3] ), .A2(n65), .A3(n96), .A4(n79), .Y(n248)
         );
  AO22X1_HVT U216 ( .A1(\mem[8][2] ), .A2(n65), .A3(n96), .A4(n80), .Y(n249)
         );
  AO22X1_HVT U217 ( .A1(\mem[8][1] ), .A2(n65), .A3(n96), .A4(n81), .Y(n250)
         );
  AO22X1_HVT U218 ( .A1(\mem[8][0] ), .A2(n65), .A3(n96), .A4(n82), .Y(n251)
         );
  AND2X1_HVT U219 ( .A1(n94), .A2(n86), .Y(n96) );
  AND2X1_HVT U220 ( .A1(n95), .A2(n97), .Y(n86) );
  AND2X1_HVT U221 ( .A1(write), .A2(a_din[3]), .Y(n95) );
  AO22X1_HVT U222 ( .A1(\mem[7][15] ), .A2(n65), .A3(n98), .A4(n67), .Y(n252)
         );
  AO22X1_HVT U223 ( .A1(\mem[7][14] ), .A2(n65), .A3(n98), .A4(n68), .Y(n253)
         );
  AO22X1_HVT U224 ( .A1(\mem[7][13] ), .A2(n65), .A3(n98), .A4(n69), .Y(n254)
         );
  AO22X1_HVT U225 ( .A1(\mem[7][12] ), .A2(n65), .A3(n98), .A4(n70), .Y(n255)
         );
  AO22X1_HVT U226 ( .A1(\mem[7][11] ), .A2(n65), .A3(n98), .A4(n71), .Y(n256)
         );
  AO22X1_HVT U227 ( .A1(\mem[7][10] ), .A2(n65), .A3(n98), .A4(n72), .Y(n257)
         );
  AO22X1_HVT U228 ( .A1(\mem[7][9] ), .A2(n65), .A3(n98), .A4(n73), .Y(n258)
         );
  AO22X1_HVT U229 ( .A1(\mem[7][8] ), .A2(n65), .A3(n98), .A4(n74), .Y(n259)
         );
  AO22X1_HVT U230 ( .A1(\mem[7][7] ), .A2(n65), .A3(n98), .A4(n75), .Y(n260)
         );
  AO22X1_HVT U231 ( .A1(\mem[7][6] ), .A2(n65), .A3(n98), .A4(n76), .Y(n261)
         );
  AO22X1_HVT U232 ( .A1(\mem[7][5] ), .A2(n65), .A3(n98), .A4(n77), .Y(n262)
         );
  AO22X1_HVT U233 ( .A1(\mem[7][4] ), .A2(n65), .A3(n98), .A4(n78), .Y(n263)
         );
  AO22X1_HVT U234 ( .A1(\mem[7][3] ), .A2(n65), .A3(n98), .A4(n79), .Y(n264)
         );
  AO22X1_HVT U235 ( .A1(\mem[7][2] ), .A2(n65), .A3(n98), .A4(n80), .Y(n265)
         );
  AO22X1_HVT U236 ( .A1(\mem[7][1] ), .A2(n65), .A3(n98), .A4(n81), .Y(n266)
         );
  AO22X1_HVT U237 ( .A1(\mem[7][0] ), .A2(n65), .A3(n98), .A4(n82), .Y(n267)
         );
  AND2X1_HVT U238 ( .A1(n99), .A2(n83), .Y(n98) );
  AO22X1_HVT U239 ( .A1(\mem[6][15] ), .A2(n65), .A3(n100), .A4(n67), .Y(n268)
         );
  AO22X1_HVT U240 ( .A1(\mem[6][14] ), .A2(n65), .A3(n100), .A4(n68), .Y(n269)
         );
  AO22X1_HVT U241 ( .A1(\mem[6][13] ), .A2(n65), .A3(n100), .A4(n69), .Y(n270)
         );
  AO22X1_HVT U242 ( .A1(\mem[6][12] ), .A2(n65), .A3(n100), .A4(n70), .Y(n271)
         );
  AO22X1_HVT U243 ( .A1(\mem[6][11] ), .A2(n65), .A3(n100), .A4(n71), .Y(n272)
         );
  AO22X1_HVT U244 ( .A1(\mem[6][10] ), .A2(n65), .A3(n100), .A4(n72), .Y(n273)
         );
  AO22X1_HVT U245 ( .A1(\mem[6][9] ), .A2(n65), .A3(n100), .A4(n73), .Y(n274)
         );
  AO22X1_HVT U246 ( .A1(\mem[6][8] ), .A2(n65), .A3(n100), .A4(n74), .Y(n275)
         );
  AO22X1_HVT U247 ( .A1(\mem[6][7] ), .A2(n65), .A3(n100), .A4(n75), .Y(n276)
         );
  AO22X1_HVT U248 ( .A1(\mem[6][6] ), .A2(n65), .A3(n100), .A4(n76), .Y(n277)
         );
  AO22X1_HVT U249 ( .A1(\mem[6][5] ), .A2(n65), .A3(n100), .A4(n77), .Y(n278)
         );
  AO22X1_HVT U250 ( .A1(\mem[6][4] ), .A2(n65), .A3(n100), .A4(n78), .Y(n279)
         );
  AO22X1_HVT U251 ( .A1(\mem[6][3] ), .A2(n65), .A3(n100), .A4(n79), .Y(n280)
         );
  AO22X1_HVT U252 ( .A1(\mem[6][2] ), .A2(n65), .A3(n100), .A4(n80), .Y(n281)
         );
  AO22X1_HVT U253 ( .A1(\mem[6][1] ), .A2(n65), .A3(n100), .A4(n81), .Y(n282)
         );
  AO22X1_HVT U254 ( .A1(\mem[6][0] ), .A2(n65), .A3(n100), .A4(n82), .Y(n283)
         );
  AND2X1_HVT U255 ( .A1(n101), .A2(n83), .Y(n100) );
  AND2X1_HVT U256 ( .A1(a_din[2]), .A2(a_din[1]), .Y(n83) );
  AO22X1_HVT U257 ( .A1(\mem[5][15] ), .A2(n65), .A3(n102), .A4(n67), .Y(n284)
         );
  AO22X1_HVT U258 ( .A1(\mem[5][14] ), .A2(n65), .A3(n102), .A4(n68), .Y(n285)
         );
  AO22X1_HVT U259 ( .A1(\mem[5][13] ), .A2(n65), .A3(n102), .A4(n69), .Y(n286)
         );
  AO22X1_HVT U260 ( .A1(\mem[5][12] ), .A2(n65), .A3(n102), .A4(n70), .Y(n287)
         );
  AO22X1_HVT U261 ( .A1(\mem[5][11] ), .A2(n65), .A3(n102), .A4(n71), .Y(n288)
         );
  AO22X1_HVT U262 ( .A1(\mem[5][10] ), .A2(n65), .A3(n102), .A4(n72), .Y(n289)
         );
  AO22X1_HVT U263 ( .A1(\mem[5][9] ), .A2(n65), .A3(n102), .A4(n73), .Y(n290)
         );
  AO22X1_HVT U264 ( .A1(\mem[5][8] ), .A2(n65), .A3(n102), .A4(n74), .Y(n291)
         );
  AO22X1_HVT U265 ( .A1(\mem[5][7] ), .A2(n65), .A3(n102), .A4(n75), .Y(n292)
         );
  AO22X1_HVT U266 ( .A1(\mem[5][6] ), .A2(n65), .A3(n102), .A4(n76), .Y(n293)
         );
  AO22X1_HVT U267 ( .A1(\mem[5][5] ), .A2(n65), .A3(n102), .A4(n77), .Y(n294)
         );
  AO22X1_HVT U268 ( .A1(\mem[5][4] ), .A2(n65), .A3(n102), .A4(n78), .Y(n295)
         );
  AO22X1_HVT U269 ( .A1(\mem[5][3] ), .A2(n65), .A3(n102), .A4(n79), .Y(n296)
         );
  AO22X1_HVT U270 ( .A1(\mem[5][2] ), .A2(n65), .A3(n102), .A4(n80), .Y(n297)
         );
  AO22X1_HVT U271 ( .A1(\mem[5][1] ), .A2(n65), .A3(n102), .A4(n81), .Y(n298)
         );
  AO22X1_HVT U272 ( .A1(\mem[5][0] ), .A2(n65), .A3(n102), .A4(n82), .Y(n299)
         );
  AND2X1_HVT U273 ( .A1(n99), .A2(n88), .Y(n102) );
  AO22X1_HVT U274 ( .A1(\mem[4][15] ), .A2(n65), .A3(n103), .A4(n67), .Y(n300)
         );
  AO22X1_HVT U275 ( .A1(\mem[4][14] ), .A2(n65), .A3(n103), .A4(n68), .Y(n301)
         );
  AO22X1_HVT U276 ( .A1(\mem[4][13] ), .A2(n65), .A3(n103), .A4(n69), .Y(n302)
         );
  AO22X1_HVT U277 ( .A1(\mem[4][12] ), .A2(n65), .A3(n103), .A4(n70), .Y(n303)
         );
  AO22X1_HVT U278 ( .A1(\mem[4][11] ), .A2(n65), .A3(n103), .A4(n71), .Y(n304)
         );
  AO22X1_HVT U279 ( .A1(\mem[4][10] ), .A2(n65), .A3(n103), .A4(n72), .Y(n305)
         );
  AO22X1_HVT U280 ( .A1(\mem[4][9] ), .A2(n65), .A3(n103), .A4(n73), .Y(n306)
         );
  AO22X1_HVT U281 ( .A1(\mem[4][8] ), .A2(n65), .A3(n103), .A4(n74), .Y(n307)
         );
  AO22X1_HVT U282 ( .A1(\mem[4][7] ), .A2(n65), .A3(n103), .A4(n75), .Y(n308)
         );
  AO22X1_HVT U283 ( .A1(\mem[4][6] ), .A2(n65), .A3(n103), .A4(n76), .Y(n309)
         );
  AO22X1_HVT U284 ( .A1(\mem[4][5] ), .A2(n65), .A3(n103), .A4(n77), .Y(n310)
         );
  AO22X1_HVT U285 ( .A1(\mem[4][4] ), .A2(n65), .A3(n103), .A4(n78), .Y(n311)
         );
  AO22X1_HVT U286 ( .A1(\mem[4][3] ), .A2(n65), .A3(n103), .A4(n79), .Y(n312)
         );
  AO22X1_HVT U287 ( .A1(\mem[4][2] ), .A2(n65), .A3(n103), .A4(n80), .Y(n313)
         );
  AO22X1_HVT U288 ( .A1(\mem[4][1] ), .A2(n65), .A3(n103), .A4(n81), .Y(n314)
         );
  AO22X1_HVT U289 ( .A1(\mem[4][0] ), .A2(n65), .A3(n103), .A4(n82), .Y(n315)
         );
  AND2X1_HVT U290 ( .A1(n101), .A2(n88), .Y(n103) );
  AND2X1_HVT U291 ( .A1(a_din[2]), .A2(n104), .Y(n88) );
  AO22X1_HVT U292 ( .A1(\mem[3][15] ), .A2(n65), .A3(n105), .A4(n67), .Y(n316)
         );
  AO22X1_HVT U293 ( .A1(\mem[3][14] ), .A2(n65), .A3(n105), .A4(n68), .Y(n317)
         );
  AO22X1_HVT U294 ( .A1(\mem[3][13] ), .A2(n65), .A3(n105), .A4(n69), .Y(n318)
         );
  AO22X1_HVT U295 ( .A1(\mem[3][12] ), .A2(n65), .A3(n105), .A4(n70), .Y(n319)
         );
  AO22X1_HVT U296 ( .A1(\mem[3][11] ), .A2(n65), .A3(n105), .A4(n71), .Y(n320)
         );
  AO22X1_HVT U297 ( .A1(\mem[3][10] ), .A2(n65), .A3(n105), .A4(n72), .Y(n321)
         );
  AO22X1_HVT U298 ( .A1(\mem[3][9] ), .A2(n65), .A3(n105), .A4(n73), .Y(n322)
         );
  AO22X1_HVT U299 ( .A1(\mem[3][8] ), .A2(n65), .A3(n105), .A4(n74), .Y(n323)
         );
  AO22X1_HVT U300 ( .A1(\mem[3][7] ), .A2(n65), .A3(n105), .A4(n75), .Y(n324)
         );
  AO22X1_HVT U301 ( .A1(\mem[3][6] ), .A2(n65), .A3(n105), .A4(n76), .Y(n325)
         );
  AO22X1_HVT U302 ( .A1(\mem[3][5] ), .A2(n65), .A3(n105), .A4(n77), .Y(n326)
         );
  AO22X1_HVT U303 ( .A1(\mem[3][4] ), .A2(n65), .A3(n105), .A4(n78), .Y(n327)
         );
  AO22X1_HVT U304 ( .A1(\mem[3][3] ), .A2(n65), .A3(n105), .A4(n79), .Y(n328)
         );
  AO22X1_HVT U305 ( .A1(\mem[3][2] ), .A2(n65), .A3(n105), .A4(n80), .Y(n329)
         );
  AO22X1_HVT U306 ( .A1(\mem[3][1] ), .A2(n65), .A3(n105), .A4(n81), .Y(n330)
         );
  AO22X1_HVT U307 ( .A1(\mem[3][0] ), .A2(n65), .A3(n105), .A4(n82), .Y(n331)
         );
  AND2X1_HVT U308 ( .A1(n99), .A2(n91), .Y(n105) );
  AO22X1_HVT U309 ( .A1(\mem[2][15] ), .A2(n65), .A3(n106), .A4(n67), .Y(n332)
         );
  AO22X1_HVT U310 ( .A1(\mem[2][14] ), .A2(n65), .A3(n106), .A4(n68), .Y(n333)
         );
  AO22X1_HVT U311 ( .A1(\mem[2][13] ), .A2(n65), .A3(n106), .A4(n69), .Y(n334)
         );
  AO22X1_HVT U312 ( .A1(\mem[2][12] ), .A2(n65), .A3(n106), .A4(n70), .Y(n335)
         );
  AO22X1_HVT U313 ( .A1(\mem[2][11] ), .A2(n65), .A3(n106), .A4(n71), .Y(n336)
         );
  AO22X1_HVT U314 ( .A1(\mem[2][10] ), .A2(n65), .A3(n106), .A4(n72), .Y(n337)
         );
  AO22X1_HVT U315 ( .A1(\mem[2][9] ), .A2(n65), .A3(n106), .A4(n73), .Y(n338)
         );
  AO22X1_HVT U316 ( .A1(\mem[2][8] ), .A2(n65), .A3(n106), .A4(n74), .Y(n339)
         );
  AO22X1_HVT U317 ( .A1(\mem[2][7] ), .A2(n65), .A3(n106), .A4(n75), .Y(n340)
         );
  AO22X1_HVT U318 ( .A1(\mem[2][6] ), .A2(n65), .A3(n106), .A4(n76), .Y(n341)
         );
  AO22X1_HVT U319 ( .A1(\mem[2][5] ), .A2(n65), .A3(n106), .A4(n77), .Y(n342)
         );
  AO22X1_HVT U320 ( .A1(\mem[2][4] ), .A2(n65), .A3(n106), .A4(n78), .Y(n343)
         );
  AO22X1_HVT U321 ( .A1(\mem[2][3] ), .A2(n65), .A3(n106), .A4(n79), .Y(n344)
         );
  AO22X1_HVT U322 ( .A1(\mem[2][2] ), .A2(n65), .A3(n106), .A4(n80), .Y(n345)
         );
  AO22X1_HVT U323 ( .A1(\mem[2][1] ), .A2(n65), .A3(n106), .A4(n81), .Y(n346)
         );
  AO22X1_HVT U324 ( .A1(\mem[2][0] ), .A2(n65), .A3(n106), .A4(n82), .Y(n347)
         );
  AND2X1_HVT U325 ( .A1(n101), .A2(n91), .Y(n106) );
  AND2X1_HVT U326 ( .A1(a_din[1]), .A2(n107), .Y(n91) );
  AO22X1_HVT U327 ( .A1(\mem[1][15] ), .A2(n65), .A3(n108), .A4(n67), .Y(n348)
         );
  AO22X1_HVT U328 ( .A1(\mem[1][14] ), .A2(n65), .A3(n108), .A4(n68), .Y(n349)
         );
  AO22X1_HVT U329 ( .A1(\mem[1][13] ), .A2(n65), .A3(n108), .A4(n69), .Y(n350)
         );
  AO22X1_HVT U330 ( .A1(\mem[1][12] ), .A2(n65), .A3(n108), .A4(n70), .Y(n351)
         );
  AO22X1_HVT U331 ( .A1(\mem[1][11] ), .A2(n65), .A3(n108), .A4(n71), .Y(n352)
         );
  AO22X1_HVT U332 ( .A1(\mem[1][10] ), .A2(n65), .A3(n108), .A4(n72), .Y(n353)
         );
  AO22X1_HVT U333 ( .A1(\mem[1][9] ), .A2(n65), .A3(n108), .A4(n73), .Y(n354)
         );
  AO22X1_HVT U334 ( .A1(\mem[1][8] ), .A2(n65), .A3(n108), .A4(n74), .Y(n355)
         );
  AO22X1_HVT U335 ( .A1(\mem[1][7] ), .A2(n65), .A3(n108), .A4(n75), .Y(n356)
         );
  AO22X1_HVT U336 ( .A1(\mem[1][6] ), .A2(n65), .A3(n108), .A4(n76), .Y(n357)
         );
  AO22X1_HVT U337 ( .A1(\mem[1][5] ), .A2(n65), .A3(n108), .A4(n77), .Y(n358)
         );
  AO22X1_HVT U338 ( .A1(\mem[1][4] ), .A2(n65), .A3(n108), .A4(n78), .Y(n359)
         );
  AO22X1_HVT U339 ( .A1(\mem[1][3] ), .A2(n65), .A3(n108), .A4(n79), .Y(n360)
         );
  AO22X1_HVT U340 ( .A1(\mem[1][2] ), .A2(n65), .A3(n108), .A4(n80), .Y(n361)
         );
  AO22X1_HVT U341 ( .A1(\mem[1][1] ), .A2(n65), .A3(n108), .A4(n81), .Y(n362)
         );
  AO22X1_HVT U342 ( .A1(\mem[1][0] ), .A2(n65), .A3(n108), .A4(n82), .Y(n363)
         );
  AND2X1_HVT U343 ( .A1(n99), .A2(n94), .Y(n108) );
  AND2X1_HVT U344 ( .A1(n109), .A2(a_din[0]), .Y(n99) );
  AO22X1_HVT U345 ( .A1(\mem[0][15] ), .A2(n65), .A3(n110), .A4(n67), .Y(n364)
         );
  AND2X1_HVT U346 ( .A1(n111), .A2(n112), .Y(n67) );
  AO22X1_HVT U347 ( .A1(\mem[0][14] ), .A2(n65), .A3(n110), .A4(n68), .Y(n365)
         );
  AND2X1_HVT U348 ( .A1(n113), .A2(n111), .Y(n68) );
  AO22X1_HVT U349 ( .A1(\mem[0][13] ), .A2(n65), .A3(n110), .A4(n69), .Y(n366)
         );
  AND2X1_HVT U350 ( .A1(n114), .A2(n111), .Y(n69) );
  AO22X1_HVT U351 ( .A1(\mem[0][12] ), .A2(n65), .A3(n110), .A4(n70), .Y(n367)
         );
  AND2X1_HVT U352 ( .A1(n115), .A2(n111), .Y(n70) );
  AND2X1_HVT U353 ( .A1(a_addr[3]), .A2(a_addr[2]), .Y(n111) );
  AO22X1_HVT U354 ( .A1(\mem[0][11] ), .A2(n65), .A3(n110), .A4(n71), .Y(n368)
         );
  AND2X1_HVT U355 ( .A1(n116), .A2(n112), .Y(n71) );
  AO22X1_HVT U356 ( .A1(\mem[0][10] ), .A2(n65), .A3(n110), .A4(n72), .Y(n369)
         );
  AND2X1_HVT U357 ( .A1(n116), .A2(n113), .Y(n72) );
  AO22X1_HVT U358 ( .A1(\mem[0][9] ), .A2(n65), .A3(n110), .A4(n73), .Y(n370)
         );
  AND2X1_HVT U359 ( .A1(n116), .A2(n114), .Y(n73) );
  AO22X1_HVT U360 ( .A1(\mem[0][8] ), .A2(n65), .A3(n110), .A4(n74), .Y(n371)
         );
  AND2X1_HVT U361 ( .A1(n116), .A2(n115), .Y(n74) );
  AND2X1_HVT U362 ( .A1(a_addr[3]), .A2(n117), .Y(n116) );
  AO22X1_HVT U363 ( .A1(\mem[0][7] ), .A2(n65), .A3(n110), .A4(n75), .Y(n372)
         );
  AND2X1_HVT U364 ( .A1(n118), .A2(n112), .Y(n75) );
  AO22X1_HVT U365 ( .A1(\mem[0][6] ), .A2(n65), .A3(n110), .A4(n76), .Y(n373)
         );
  AND2X1_HVT U366 ( .A1(n118), .A2(n113), .Y(n76) );
  AO22X1_HVT U367 ( .A1(\mem[0][5] ), .A2(n65), .A3(n110), .A4(n77), .Y(n374)
         );
  AND2X1_HVT U368 ( .A1(n118), .A2(n114), .Y(n77) );
  AO22X1_HVT U369 ( .A1(\mem[0][4] ), .A2(n65), .A3(n110), .A4(n78), .Y(n375)
         );
  AND2X1_HVT U370 ( .A1(n118), .A2(n115), .Y(n78) );
  AND2X1_HVT U371 ( .A1(a_addr[2]), .A2(n119), .Y(n118) );
  AO22X1_HVT U372 ( .A1(\mem[0][3] ), .A2(n65), .A3(n110), .A4(n79), .Y(n376)
         );
  AND2X1_HVT U373 ( .A1(n120), .A2(n112), .Y(n79) );
  AND3X1_HVT U374 ( .A1(a_addr[0]), .A2(n65), .A3(a_addr[1]), .Y(n112) );
  AO22X1_HVT U375 ( .A1(\mem[0][2] ), .A2(n65), .A3(n110), .A4(n80), .Y(n377)
         );
  AND2X1_HVT U376 ( .A1(n120), .A2(n113), .Y(n80) );
  AND3X1_HVT U377 ( .A1(n121), .A2(n65), .A3(a_addr[1]), .Y(n113) );
  AO22X1_HVT U378 ( .A1(\mem[0][1] ), .A2(n65), .A3(n110), .A4(n81), .Y(n378)
         );
  AND2X1_HVT U379 ( .A1(n120), .A2(n114), .Y(n81) );
  AND3X1_HVT U380 ( .A1(n122), .A2(n65), .A3(a_addr[0]), .Y(n114) );
  AO22X1_HVT U381 ( .A1(\mem[0][0] ), .A2(n65), .A3(n110), .A4(n82), .Y(n379)
         );
  AND2X1_HVT U382 ( .A1(n120), .A2(n115), .Y(n82) );
  AND3X1_HVT U383 ( .A1(n122), .A2(n65), .A3(n121), .Y(n115) );
  INVX0_HVT U384 ( .A(a_addr[0]), .Y(n121) );
  INVX0_HVT U385 ( .A(a_addr[1]), .Y(n122) );
  AND2X1_HVT U386 ( .A1(n117), .A2(n119), .Y(n120) );
  INVX0_HVT U387 ( .A(a_addr[3]), .Y(n119) );
  INVX0_HVT U388 ( .A(a_addr[2]), .Y(n117) );
  AND2X1_HVT U389 ( .A1(n101), .A2(n94), .Y(n110) );
  AND2X1_HVT U390 ( .A1(n104), .A2(n107), .Y(n94) );
  INVX0_HVT U391 ( .A(a_din[2]), .Y(n107) );
  INVX0_HVT U392 ( .A(a_din[1]), .Y(n104) );
  AND2X1_HVT U393 ( .A1(n109), .A2(n97), .Y(n101) );
  INVX0_HVT U394 ( .A(a_din[0]), .Y(n97) );
  AND2X1_HVT U395 ( .A1(write), .A2(n123), .Y(n109) );
  INVX0_HVT U396 ( .A(a_din[3]), .Y(n123) );
  INVX0_HVT U397 ( .A(rst), .Y(n65) );
endmodule

