
module inv_sbox_1 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n196, n197, n198, n199, n200, n201, n202, n208, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663;

  NAND2X0_HVT U4 ( .A1(n296), .A2(n382), .Y(n660) );
  NAND2X0_HVT U5 ( .A1(n660), .A2(n380), .Y(n659) );
  NAND2X0_HVT U7 ( .A1(n385), .A2(n661), .Y(n656) );
  NAND2X0_HVT U8 ( .A1(n296), .A2(n380), .Y(n655) );
  NAND2X0_HVT U9 ( .A1(n236), .A2(n655), .Y(n654) );
  NAND2X0_HVT U10 ( .A1(n235), .A2(n652), .Y(n653) );
  NAND2X0_HVT U11 ( .A1(n389), .A2(n382), .Y(n651) );
  NAND2X0_HVT U12 ( .A1(n297), .A2(n368), .Y(n650) );
  NAND2X0_HVT U13 ( .A1(n661), .A2(n248), .Y(n649) );
  NAND2X0_HVT U15 ( .A1(n378), .A2(n384), .Y(n647) );
  NAND2X0_HVT U19 ( .A1(n387), .A2(n282), .Y(n642) );
  NAND2X0_HVT U32 ( .A1(n370), .A2(n389), .Y(n630) );
  NAND2X0_HVT U35 ( .A1(n655), .A2(n261), .Y(n627) );
  NAND2X0_HVT U38 ( .A1(n368), .A2(n389), .Y(n624) );
  NAND2X0_HVT U42 ( .A1(n657), .A2(n261), .Y(n620) );
  OA21X1_HVT U53 ( .A1(n395), .A2(n612), .A3(n421), .Y(n610) );
  NAND2X0_HVT U55 ( .A1(n290), .A2(n660), .Y(n608) );
  MUX41X1_HVT U56 ( .A1(n435), .A3(n378), .A2(n420), .A4(n608), .S0(n361), 
        .S1(n345), .Y(n607) );
  AO21X1_HVT U60 ( .A1(n602), .A2(n334), .A3(n641), .Y(n603) );
  MUX41X1_HVT U62 ( .A1(n601), .A3(n607), .A2(n605), .A4(n609), .S0(n376), 
        .S1(n373), .Y(n600) );
  MUX41X1_HVT U65 ( .A1(n414), .A3(n416), .A2(n415), .A4(n624), .S0(n361), 
        .S1(n345), .Y(n597) );
  NAND2X0_HVT U66 ( .A1(n298), .A2(n356), .Y(n596) );
  MUX41X1_HVT U67 ( .A1(n411), .A3(n436), .A2(n413), .A4(n596), .S0(n364), 
        .S1(n358), .Y(n595) );
  MUX41X1_HVT U68 ( .A1(n411), .A3(n272), .A2(n412), .A4(n235), .S0(n360), 
        .S1(n345), .Y(n594) );
  MUX41X1_HVT U69 ( .A1(n594), .A3(n597), .A2(n595), .A4(n598), .S0(n376), 
        .S1(n373), .Y(n593) );
  NAND2X0_HVT U72 ( .A1(n378), .A2(n656), .Y(n591) );
  MUX41X1_HVT U73 ( .A1(n635), .A3(n591), .A2(n437), .A4(n367), .S0(n365), 
        .S1(n358), .Y(n590) );
  MUX41X1_HVT U80 ( .A1(n439), .A3(n435), .A2(n654), .A4(n659), .S0(n360), 
        .S1(n392), .Y(n583) );
  NAND2X0_HVT U81 ( .A1(n382), .A2(n656), .Y(n582) );
  AND2X1_HVT U82 ( .A1(n299), .A2(n661), .Y(n581) );
  MUX41X1_HVT U88 ( .A1(n413), .A3(n398), .A2(n632), .A4(n616), .S0(n360), 
        .S1(n393), .Y(n576) );
  NAND2X0_HVT U89 ( .A1(n322), .A2(n281), .Y(n575) );
  MUX41X1_HVT U90 ( .A1(n241), .A3(n656), .A2(n615), .A4(n575), .S0(n360), 
        .S1(n345), .Y(n574) );
  MUX41X1_HVT U99 ( .A1(n630), .A3(n415), .A2(n614), .A4(n378), .S0(n345), 
        .S1(n358), .Y(n565) );
  NAND2X0_HVT U100 ( .A1(n389), .A2(n450), .Y(n564) );
  MUX41X1_HVT U101 ( .A1(n444), .A3(n650), .A2(n426), .A4(n564), .S0(n345), 
        .S1(n357), .Y(n563) );
  AND2X1_HVT U104 ( .A1(n656), .A2(n379), .Y(n561) );
  MUX41X1_HVT U105 ( .A1(n648), .A3(n445), .A2(n582), .A4(n561), .S0(n361), 
        .S1(n393), .Y(n560) );
  MUX41X1_HVT U107 ( .A1(n444), .A3(n661), .A2(n559), .A4(n404), .S0(n360), 
        .S1(n391), .Y(n558) );
  MUX41X1_HVT U108 ( .A1(n417), .A3(n378), .A2(n420), .A4(n381), .S0(n361), 
        .S1(n393), .Y(n557) );
  MUX41X1_HVT U109 ( .A1(n443), .A3(n398), .A2(n440), .A4(n433), .S0(n360), 
        .S1(n391), .Y(n556) );
  MUX41X1_HVT U110 ( .A1(n556), .A3(n558), .A2(n557), .A4(n560), .S0(in[5]), 
        .S1(n374), .Y(n555) );
  AO21X1_HVT U112 ( .A1(n429), .A2(n365), .A3(n638), .Y(n553) );
  NAND2X0_HVT U114 ( .A1(n237), .A2(n656), .Y(n551) );
  MUX41X1_HVT U115 ( .A1(n551), .A3(n651), .A2(n429), .A4(n661), .S0(n345), 
        .S1(n358), .Y(n550) );
  MUX41X1_HVT U116 ( .A1(n428), .A3(n422), .A2(n398), .A4(n647), .S0(n359), 
        .S1(n393), .Y(n549) );
  NAND2X0_HVT U118 ( .A1(n322), .A2(n272), .Y(n547) );
  MUX41X1_HVT U119 ( .A1(n446), .A3(n548), .A2(n625), .A4(n547), .S0(n359), 
        .S1(n391), .Y(n546) );
  MUX41X1_HVT U122 ( .A1(n434), .A3(n350), .A2(n616), .A4(n438), .S0(n359), 
        .S1(n334), .Y(n544) );
  MUX41X1_HVT U124 ( .A1(n352), .A3(n543), .A2(n639), .A4(n231), .S0(n334), 
        .S1(n359), .Y(n542) );
  AOI21X1_HVT U127 ( .A1(n363), .A2(n538), .A3(n405), .Y(n539) );
  NAND2X0_HVT U129 ( .A1(n313), .A2(n235), .Y(n536) );
  MUX41X1_HVT U130 ( .A1(n536), .A3(n537), .A2(n540), .A4(n539), .S0(n364), 
        .S1(n374), .Y(n535) );
  AND2X1_HVT U131 ( .A1(n356), .A2(n388), .Y(n534) );
  MUX41X1_HVT U132 ( .A1(n402), .A3(n534), .A2(n448), .A4(n411), .S0(n365), 
        .S1(n361), .Y(n533) );
  MUX41X1_HVT U133 ( .A1(n449), .A3(n404), .A2(n608), .A4(n403), .S0(n334), 
        .S1(n357), .Y(n532) );
  MUX41X1_HVT U136 ( .A1(n613), .A3(n564), .A2(n530), .A4(n409), .S0(n313), 
        .S1(n345), .Y(n529) );
  MUX41X1_HVT U137 ( .A1(n248), .A3(n633), .A2(n637), .A4(n442), .S0(n364), 
        .S1(n357), .Y(n528) );
  NAND2X0_HVT U141 ( .A1(n378), .A2(n322), .Y(n525) );
  MUX41X1_HVT U142 ( .A1(n525), .A3(n623), .A2(n447), .A4(n419), .S0(n363), 
        .S1(n391), .Y(n524) );
  MUX41X1_HVT U143 ( .A1(n281), .A3(n430), .A2(n642), .A4(n639), .S0(n362), 
        .S1(n392), .Y(n523) );
  MUX41X1_HVT U145 ( .A1(n631), .A3(n445), .A2(n522), .A4(n582), .S0(n363), 
        .S1(n391), .Y(n521) );
  MUX41X1_HVT U146 ( .A1(n521), .A3(n523), .A2(n524), .A4(n526), .S0(n374), 
        .S1(n376), .Y(n520) );
  MUX41X1_HVT U151 ( .A1(n249), .A3(n427), .A2(n278), .A4(n516), .S0(n334), 
        .S1(n357), .Y(n515) );
  MUX41X1_HVT U155 ( .A1(n419), .A3(n651), .A2(n643), .A4(n310), .S0(n362), 
        .S1(n364), .Y(n511) );
  NAND2X0_HVT U159 ( .A1(n507), .A2(n506), .Y(n508) );
  NAND2X0_HVT U163 ( .A1(n385), .A2(n281), .Y(n502) );
  NAND2X0_HVT U166 ( .A1(n652), .A2(n498), .Y(n499) );
  NAND2X0_HVT U177 ( .A1(n297), .A2(n272), .Y(n488) );
  AND2X1_HVT U179 ( .A1(n299), .A2(n379), .Y(n486) );
  MUX41X1_HVT U180 ( .A1(n630), .A3(n396), .A2(n486), .A4(n617), .S0(n362), 
        .S1(n393), .Y(n485) );
  MUX41X1_HVT U182 ( .A1(n404), .A3(n316), .A2(n401), .A4(n249), .S0(n359), 
        .S1(n391), .Y(n483) );
  AND2X1_HVT U185 ( .A1(n453), .A2(n388), .Y(n480) );
  NAND2X0_HVT U191 ( .A1(n268), .A2(n410), .Y(n474) );
  AND2X1_HVT U192 ( .A1(n425), .A2(n472), .Y(n473) );
  NAND2X0_HVT U194 ( .A1(n620), .A2(n472), .Y(n470) );
  MUX41X1_HVT U195 ( .A1(n471), .A3(n470), .A2(n473), .A4(n474), .S0(n360), 
        .S1(n374), .Y(n469) );
  NAND2X0_HVT U198 ( .A1(n284), .A2(n261), .Y(n652) );
  NAND2X0_HVT U200 ( .A1(n380), .A2(n322), .Y(n538) );
  NAND2X0_HVT U207 ( .A1(n322), .A2(n241), .Y(n602) );
  MUX21X1_HVT U1 ( .A1(n261), .A2(n197), .S0(n198), .Y(n196) );
  IBUFFX16_HVT U2 ( .A(n196), .Y(n573) );
  IBUFFX16_HVT U3 ( .A(n371), .Y(n197) );
  IBUFFX16_HVT U6 ( .A(n268), .Y(n198) );
  INVX2_HVT U14 ( .A(n377), .Y(n261) );
  XOR2X2_HVT U16 ( .A1(n377), .A2(n385), .Y(n616) );
  INVX0_HVT U17 ( .A(n385), .Y(n226) );
  MUX41X1_HVT U18 ( .A1(n240), .A3(n236), .A2(n626), .A4(n381), .S0(n199), 
        .S1(n391), .Y(n491) );
  IBUFFX16_HVT U20 ( .A(n362), .Y(n199) );
  MUX21X1_HVT U21 ( .A1(n250), .A2(n377), .S0(n296), .Y(n249) );
  MUX41X1_HVT U22 ( .A1(n497), .A3(n503), .A2(n501), .A4(n505), .S0(n200), 
        .S1(n374), .Y(n496) );
  IBUFFX16_HVT U23 ( .A(n266), .Y(n200) );
  AO21X2_HVT U24 ( .A1(n366), .A2(n406), .A3(n450), .Y(n518) );
  AO21X1_HVT U25 ( .A1(n298), .A2(n450), .A3(n268), .Y(n472) );
  MUX21X2_HVT U26 ( .A1(n542), .A2(n544), .S0(n201), .Y(n541) );
  IBUFFX16_HVT U27 ( .A(n372), .Y(n201) );
  INVX1_HVT U28 ( .A(n244), .Y(n495) );
  IBUFFX2_HVT U29 ( .A(in[6]), .Y(n283) );
  MUX21X2_HVT U30 ( .A1(n639), .A2(n636), .S0(n233), .Y(n500) );
  IBUFFX2_HVT U31 ( .A(n362), .Y(n243) );
  MUX21X1_HVT U33 ( .A1(n290), .A2(n379), .S0(n265), .Y(n504) );
  IBUFFX2_HVT U34 ( .A(n296), .Y(n265) );
  INVX0_HVT U36 ( .A(n647), .Y(n412) );
  INVX1_HVT U37 ( .A(n231), .Y(n639) );
  MUX21X2_HVT U39 ( .A1(n370), .A2(n450), .S0(n285), .Y(n636) );
  MUX41X1_HVT U40 ( .A1(n425), .A3(n417), .A2(n653), .A4(n424), .S0(n392), 
        .S1(n227), .Y(n589) );
  NAND2X0_HVT U41 ( .A1(n281), .A2(n202), .Y(n208) );
  NAND2X0_HVT U43 ( .A1(n378), .A2(n226), .Y(n218) );
  NAND2X0_HVT U44 ( .A1(n208), .A2(n218), .Y(n628) );
  INVX0_HVT U45 ( .A(n226), .Y(n202) );
  INVX1_HVT U46 ( .A(n641), .Y(n417) );
  INVX2_HVT U47 ( .A(n629), .Y(n424) );
  IBUFFX2_HVT U48 ( .A(n361), .Y(n227) );
  INVX1_HVT U49 ( .A(n335), .Y(n392) );
  INVX1_HVT U50 ( .A(n658), .Y(n281) );
  INVX0_HVT U51 ( .A(n628), .Y(n425) );
  INVX4_HVT U52 ( .A(n335), .Y(n345) );
  INVX1_HVT U54 ( .A(in[5]), .Y(n223) );
  INVX0_HVT U57 ( .A(n387), .Y(n224) );
  INVX0_HVT U58 ( .A(n271), .Y(n219) );
  INVX1_HVT U59 ( .A(n347), .Y(n271) );
  NAND2X0_HVT U61 ( .A1(n240), .A2(n220), .Y(n221) );
  NAND2X0_HVT U63 ( .A1(n378), .A2(n387), .Y(n222) );
  NAND2X0_HVT U64 ( .A1(n221), .A2(n222), .Y(n462) );
  IBUFFX2_HVT U70 ( .A(n387), .Y(n220) );
  INVX0_HVT U71 ( .A(n462), .Y(n441) );
  MUX41X1_HVT U74 ( .A1(n566), .A3(n563), .A2(n568), .A4(n565), .S0(n223), 
        .S1(n373), .Y(n562) );
  INVX1_HVT U75 ( .A(n388), .Y(n385) );
  AO21X2_HVT U76 ( .A1(n378), .A2(n316), .A3(n395), .Y(n498) );
  IBUFFX2_HVT U77 ( .A(n342), .Y(n269) );
  INVX1_HVT U78 ( .A(n274), .Y(n270) );
  IBUFFX8_HVT U79 ( .A(n376), .Y(n274) );
  NBUFFX4_HVT U83 ( .A(n454), .Y(n369) );
  MUX21X1_HVT U84 ( .A1(n347), .A2(n380), .S0(n224), .Y(n567) );
  MUX41X1_HVT U85 ( .A1(n427), .A3(n634), .A2(n567), .A4(n443), .S0(n225), 
        .S1(n395), .Y(n566) );
  IBUFFX16_HVT U86 ( .A(n259), .Y(n225) );
  INVX1_HVT U87 ( .A(n367), .Y(n250) );
  INVX1_HVT U91 ( .A(n282), .Y(n245) );
  INVX1_HVT U92 ( .A(n347), .Y(n232) );
  MUX21X1_HVT U93 ( .A1(n241), .A2(n451), .S0(n228), .Y(n618) );
  IBUFFX16_HVT U94 ( .A(n386), .Y(n228) );
  MUX41X1_HVT U95 ( .A1(n416), .A3(n504), .A2(n431), .A4(n627), .S0(n229), 
        .S1(n243), .Y(n503) );
  IBUFFX16_HVT U96 ( .A(n242), .Y(n229) );
  MUX41X1_HVT U97 ( .A1(n442), .A3(n310), .A2(n649), .A4(n436), .S0(n230), 
        .S1(n269), .Y(n568) );
  IBUFFX16_HVT U98 ( .A(n361), .Y(n230) );
  MUX21X1_HVT U102 ( .A1(n381), .A2(n232), .S0(n386), .Y(n231) );
  IBUFFX16_HVT U103 ( .A(n334), .Y(n233) );
  INVX0_HVT U106 ( .A(n392), .Y(n276) );
  INVX0_HVT U111 ( .A(n392), .Y(n280) );
  IBUFFX2_HVT U113 ( .A(n663), .Y(n234) );
  INVX1_HVT U117 ( .A(n234), .Y(n235) );
  INVX1_HVT U120 ( .A(n234), .Y(n236) );
  INVX0_HVT U121 ( .A(n234), .Y(n237) );
  INVX0_HVT U123 ( .A(n452), .Y(n238) );
  INVX0_HVT U125 ( .A(n452), .Y(n239) );
  INVX1_HVT U126 ( .A(n238), .Y(n240) );
  INVX1_HVT U128 ( .A(n239), .Y(n241) );
  IBUFFX16_HVT U134 ( .A(n393), .Y(n242) );
  INVX2_HVT U135 ( .A(n394), .Y(n393) );
  XNOR2X2_HVT U138 ( .A1(n369), .A2(n346), .Y(n646) );
  IBUFFX2_HVT U139 ( .A(n346), .Y(n347) );
  MUX41X1_HVT U140 ( .A1(n449), .A3(n261), .A2(n441), .A4(n608), .S0(n362), 
        .S1(n394), .Y(n490) );
  INVX1_HVT U144 ( .A(n251), .Y(n493) );
  IBUFFX2_HVT U147 ( .A(n387), .Y(n253) );
  INVX1_HVT U148 ( .A(n388), .Y(n387) );
  IBUFFX2_HVT U149 ( .A(n384), .Y(n277) );
  INVX1_HVT U150 ( .A(n388), .Y(n384) );
  MUX21X1_HVT U152 ( .A1(n236), .A2(n245), .S0(n387), .Y(n244) );
  MUX41X1_HVT U153 ( .A1(n353), .A3(n349), .A2(n352), .A4(n495), .S0(n246), 
        .S1(n247), .Y(n494) );
  IBUFFX16_HVT U154 ( .A(n319), .Y(n246) );
  IBUFFX16_HVT U156 ( .A(n394), .Y(n247) );
  INVX0_HVT U157 ( .A(n387), .Y(n262) );
  MUX41X1_HVT U158 ( .A1(n654), .A3(n625), .A2(n502), .A4(n417), .S0(n391), 
        .S1(n359), .Y(n501) );
  INVX1_HVT U160 ( .A(n406), .Y(n248) );
  INVX2_HVT U161 ( .A(n335), .Y(n391) );
  INVX1_HVT U162 ( .A(n377), .Y(n453) );
  INVX0_HVT U164 ( .A(n626), .Y(n426) );
  MUX21X2_HVT U165 ( .A1(n369), .A2(n453), .S0(n296), .Y(n626) );
  MUX21X1_HVT U167 ( .A1(n252), .A2(n237), .S0(n253), .Y(n251) );
  IBUFFX16_HVT U168 ( .A(n371), .Y(n252) );
  MUX41X1_HVT U169 ( .A1(n640), .A3(n349), .A2(n493), .A4(n575), .S0(n254), 
        .S1(n268), .Y(n492) );
  IBUFFX16_HVT U170 ( .A(n362), .Y(n254) );
  MUX41X1_HVT U171 ( .A1(n492), .A3(n494), .A2(n490), .A4(n491), .S0(n255), 
        .S1(n375), .Y(n489) );
  IBUFFX16_HVT U172 ( .A(n372), .Y(n255) );
  INVX1_HVT U173 ( .A(n455), .Y(n449) );
  INVX2_HVT U174 ( .A(n342), .Y(n335) );
  AO21X1_HVT U175 ( .A1(n388), .A2(n237), .A3(n395), .Y(n506) );
  MUX41X1_HVT U176 ( .A1(n407), .A3(n651), .A2(n240), .A4(n299), .S0(n275), 
        .S1(n276), .Y(n592) );
  MUX21X1_HVT U178 ( .A1(n240), .A2(n451), .S0(n285), .Y(n634) );
  MUX21X1_HVT U181 ( .A1(n407), .A2(n378), .S0(n366), .Y(n571) );
  MUX41X1_HVT U183 ( .A1(n586), .A3(n589), .A2(n590), .A4(n592), .S0(n295), 
        .S1(n294), .Y(n585) );
  IBUFFX2_HVT U184 ( .A(n375), .Y(n294) );
  IBUFFX2_HVT U186 ( .A(n372), .Y(n295) );
  NAND2X1_HVT U187 ( .A1(n610), .A2(n256), .Y(n257) );
  NAND2X0_HVT U188 ( .A1(n611), .A2(n264), .Y(n258) );
  NAND2X0_HVT U189 ( .A1(n257), .A2(n258), .Y(n609) );
  INVX1_HVT U190 ( .A(n264), .Y(n256) );
  IBUFFX2_HVT U193 ( .A(n313), .Y(n264) );
  OR2X1_HVT U196 ( .A1(n371), .A2(n219), .Y(n658) );
  INVX1_HVT U197 ( .A(n371), .Y(n356) );
  IBUFFX16_HVT U199 ( .A(n361), .Y(n259) );
  MUX21X1_HVT U201 ( .A1(n237), .A2(n453), .S0(n262), .Y(n260) );
  IBUFFX16_HVT U202 ( .A(n260), .Y(n631) );
  MUX41X1_HVT U203 ( .A1(n583), .A3(n579), .A2(n584), .A4(n580), .S0(n263), 
        .S1(n373), .Y(n578) );
  IBUFFX16_HVT U204 ( .A(n376), .Y(n263) );
  INVX1_HVT U205 ( .A(n383), .Y(n452) );
  IBUFFX16_HVT U206 ( .A(n376), .Y(n266) );
  NBUFFX4_HVT U208 ( .A(n454), .Y(n371) );
  MUX21X1_HVT U209 ( .A1(n377), .A2(n371), .S0(n387), .Y(n637) );
  IBUFFX2_HVT U210 ( .A(n634), .Y(n421) );
  MUX41X1_HVT U211 ( .A1(n618), .A3(n240), .A2(n488), .A4(n353), .S0(n267), 
        .S1(n269), .Y(n487) );
  IBUFFX16_HVT U212 ( .A(n362), .Y(n267) );
  INVX2_HVT U213 ( .A(n269), .Y(n334) );
  INVX1_HVT U214 ( .A(n379), .Y(n451) );
  INVX1_HVT U215 ( .A(in[4]), .Y(n394) );
  INVX1_HVT U216 ( .A(n342), .Y(n268) );
  MUX21X1_HVT U217 ( .A1(n310), .A2(n412), .S0(n364), .Y(n611) );
  MUX41X1_HVT U218 ( .A1(n574), .A3(n570), .A2(n577), .A4(n576), .S0(n273), 
        .S1(n270), .Y(n569) );
  INVX1_HVT U219 ( .A(n271), .Y(n272) );
  MUX21X1_HVT U220 ( .A1(n368), .A2(n377), .S0(n277), .Y(n641) );
  INVX1_HVT U221 ( .A(n282), .Y(n661) );
  INVX2_HVT U222 ( .A(n342), .Y(n395) );
  IBUFFX16_HVT U223 ( .A(n373), .Y(n273) );
  NOR2X4_HVT U224 ( .A1(n346), .A2(n283), .Y(n282) );
  INVX1_HVT U225 ( .A(in[3]), .Y(n346) );
  IBUFFX16_HVT U226 ( .A(n360), .Y(n275) );
  MUX21X1_HVT U227 ( .A1(n377), .A2(n381), .S0(n386), .Y(n278) );
  IBUFFX16_HVT U228 ( .A(n278), .Y(n640) );
  MUX41X1_HVT U229 ( .A1(n637), .A3(n440), .A2(n422), .A4(n354), .S0(n279), 
        .S1(n280), .Y(n579) );
  IBUFFX16_HVT U230 ( .A(n361), .Y(n279) );
  INVX0_HVT U231 ( .A(n282), .Y(n290) );
  MUX41X1_HVT U232 ( .A1(n651), .A3(n419), .A2(n351), .A4(n424), .S0(n323), 
        .S1(n319), .Y(n526) );
  MUX21X1_HVT U233 ( .A1(n518), .A2(n519), .S0(n319), .Y(n517) );
  INVX1_HVT U234 ( .A(n388), .Y(n284) );
  INVX0_HVT U235 ( .A(n388), .Y(n285) );
  INVX0_HVT U236 ( .A(n388), .Y(n386) );
  NAND2X0_HVT U237 ( .A1(n437), .A2(n286), .Y(n287) );
  NAND2X0_HVT U238 ( .A1(n621), .A2(n365), .Y(n288) );
  NAND2X0_HVT U239 ( .A1(n287), .A2(n288), .Y(n477) );
  IBUFFX2_HVT U240 ( .A(n365), .Y(n286) );
  MUX21X1_HVT U241 ( .A1(n371), .A2(n290), .S0(n285), .Y(n289) );
  IBUFFX16_HVT U242 ( .A(n289), .Y(n621) );
  INVX0_HVT U243 ( .A(n466), .Y(n437) );
  INVX0_HVT U244 ( .A(n285), .Y(n322) );
  NAND2X0_HVT U245 ( .A1(n438), .A2(n291), .Y(n292) );
  NAND2X0_HVT U246 ( .A1(n619), .A2(n323), .Y(n293) );
  NAND2X0_HVT U247 ( .A1(n292), .A2(n293), .Y(n509) );
  IBUFFX2_HVT U248 ( .A(n323), .Y(n291) );
  INVX0_HVT U249 ( .A(n365), .Y(n323) );
  INVX0_HVT U250 ( .A(n619), .Y(n430) );
  IBUFFX2_HVT U251 ( .A(n616), .Y(n433) );
  INVX0_HVT U252 ( .A(n284), .Y(n389) );
  INVX2_HVT U253 ( .A(in[0]), .Y(n388) );
  NBUFFX2_HVT U254 ( .A(n386), .Y(n296) );
  NBUFFX2_HVT U255 ( .A(n386), .Y(n297) );
  NBUFFX2_HVT U256 ( .A(n386), .Y(n298) );
  MUX41X1_HVT U257 ( .A1(n401), .A3(n354), .A2(n441), .A4(n420), .S0(n359), 
        .S1(n345), .Y(n577) );
  INVX0_HVT U258 ( .A(n319), .Y(n313) );
  NAND2X0_HVT U259 ( .A1(n553), .A2(n306), .Y(n340) );
  INVX0_HVT U260 ( .A(n360), .Y(n306) );
  INVX1_HVT U261 ( .A(in[1]), .Y(n372) );
  INVX0_HVT U262 ( .A(n372), .Y(n373) );
  INVX1_HVT U263 ( .A(n300), .Y(n305) );
  INVX1_HVT U264 ( .A(in[7]), .Y(n300) );
  INVX1_HVT U265 ( .A(n635), .Y(n310) );
  INVX1_HVT U266 ( .A(n357), .Y(n319) );
  INVX1_HVT U267 ( .A(n375), .Y(n376) );
  INVX1_HVT U268 ( .A(in[5]), .Y(n375) );
  INVX0_HVT U269 ( .A(n618), .Y(n431) );
  INVX1_HVT U270 ( .A(n403), .Y(n299) );
  INVX1_HVT U271 ( .A(n657), .Y(n403) );
  NAND2X0_HVT U272 ( .A1(n284), .A2(n235), .Y(n657) );
  NAND2X0_HVT U273 ( .A1(n562), .A2(n300), .Y(n343) );
  NAND2X0_HVT U274 ( .A1(n510), .A2(n300), .Y(n301) );
  NAND2X0_HVT U275 ( .A1(n520), .A2(n305), .Y(n302) );
  NAND2X0_HVT U276 ( .A1(n301), .A2(n302), .Y(out[5]) );
  NAND2X0_HVT U277 ( .A1(n593), .A2(n300), .Y(n303) );
  NAND2X0_HVT U278 ( .A1(n600), .A2(in[7]), .Y(n304) );
  NAND2X0_HVT U279 ( .A1(n303), .A2(n304), .Y(out[0]) );
  INVX1_HVT U280 ( .A(n633), .Y(n422) );
  NAND2X0_HVT U281 ( .A1(n578), .A2(n300), .Y(n328) );
  INVX1_HVT U282 ( .A(n465), .Y(n438) );
  MUX41X1_HVT U283 ( .A1(n475), .A3(n484), .A2(n469), .A4(n481), .S0(n305), 
        .S1(n375), .Y(out[7]) );
  MUX41X1_HVT U284 ( .A1(n582), .A3(n249), .A2(n423), .A4(n581), .S0(n306), 
        .S1(n269), .Y(n580) );
  NAND2X0_HVT U285 ( .A1(n290), .A2(n307), .Y(n308) );
  NAND2X0_HVT U286 ( .A1(n573), .A2(n322), .Y(n309) );
  NAND2X0_HVT U287 ( .A1(n308), .A2(n309), .Y(n572) );
  IBUFFX2_HVT U288 ( .A(n322), .Y(n307) );
  NAND2X0_HVT U289 ( .A1(n499), .A2(n306), .Y(n311) );
  NAND2X0_HVT U290 ( .A1(n500), .A2(n358), .Y(n312) );
  NAND2X0_HVT U291 ( .A1(n311), .A2(n312), .Y(n497) );
  MUX41X1_HVT U292 ( .A1(n535), .A3(n541), .A2(n527), .A4(n531), .S0(n376), 
        .S1(n300), .Y(out[4]) );
  MUX41X1_HVT U293 ( .A1(n477), .A3(n478), .A2(n476), .A4(n479), .S0(n373), 
        .S1(n313), .Y(n475) );
  MUX21X2_HVT U294 ( .A1(n513), .A2(n514), .S0(n363), .Y(n512) );
  NAND2X0_HVT U295 ( .A1(n482), .A2(n372), .Y(n314) );
  NAND2X0_HVT U296 ( .A1(n483), .A2(n373), .Y(n315) );
  NAND2X0_HVT U297 ( .A1(n314), .A2(n315), .Y(n481) );
  OA21X1_HVT U298 ( .A1(n422), .A2(n395), .A3(n602), .Y(n476) );
  MUX41X1_HVT U299 ( .A1(n620), .A3(n417), .A2(n435), .A4(n430), .S0(n323), 
        .S1(n306), .Y(n482) );
  INVX1_HVT U300 ( .A(n401), .Y(n316) );
  INVX0_HVT U301 ( .A(n660), .Y(n401) );
  NAND2X0_HVT U302 ( .A1(n571), .A2(n306), .Y(n317) );
  NAND2X0_HVT U303 ( .A1(n572), .A2(n358), .Y(n318) );
  NAND2X0_HVT U304 ( .A1(n317), .A2(n318), .Y(n570) );
  NAND2X0_HVT U305 ( .A1(n533), .A2(in[1]), .Y(n320) );
  NAND2X0_HVT U306 ( .A1(n532), .A2(n372), .Y(n321) );
  NAND2X0_HVT U307 ( .A1(n320), .A2(n321), .Y(n531) );
  INVX0_HVT U308 ( .A(n620), .Y(n404) );
  NAND2X0_HVT U309 ( .A1(n637), .A2(n323), .Y(n324) );
  NAND2X0_HVT U310 ( .A1(n354), .A2(n365), .Y(n325) );
  NAND2X0_HVT U311 ( .A1(n324), .A2(n325), .Y(n514) );
  MUX41X1_HVT U312 ( .A1(n512), .A3(n517), .A2(n511), .A4(n515), .S0(n376), 
        .S1(n372), .Y(n510) );
  NAND2X0_HVT U313 ( .A1(n587), .A2(n358), .Y(n326) );
  NAND2X0_HVT U314 ( .A1(n588), .A2(n306), .Y(n327) );
  NAND2X0_HVT U315 ( .A1(n327), .A2(n326), .Y(n586) );
  NAND2X0_HVT U316 ( .A1(n585), .A2(n305), .Y(n329) );
  NAND2X0_HVT U317 ( .A1(n328), .A2(n329), .Y(out[1]) );
  OA21X1_HVT U318 ( .A1(n400), .A2(n268), .A3(n641), .Y(n587) );
  MUX21X1_HVT U319 ( .A1(n438), .A2(n397), .S0(n366), .Y(n588) );
  NAND2X0_HVT U320 ( .A1(n614), .A2(n365), .Y(n330) );
  NAND2X0_HVT U321 ( .A1(n354), .A2(n323), .Y(n331) );
  NAND2X0_HVT U322 ( .A1(n330), .A2(n331), .Y(n478) );
  INVX0_HVT U323 ( .A(n651), .Y(n396) );
  MUX21X2_HVT U324 ( .A1(n448), .A2(n402), .S0(n366), .Y(n519) );
  MUX21X2_HVT U325 ( .A1(n545), .A2(n555), .S0(n305), .Y(out[3]) );
  OA21X1_HVT U326 ( .A1(n399), .A2(n395), .A3(n408), .Y(n513) );
  MUX41X1_HVT U327 ( .A1(n552), .A3(n549), .A2(n550), .A4(n546), .S0(n375), 
        .S1(n372), .Y(n545) );
  NAND2X0_HVT U328 ( .A1(n487), .A2(n374), .Y(n332) );
  NAND2X0_HVT U329 ( .A1(n485), .A2(n372), .Y(n333) );
  NAND2X0_HVT U330 ( .A1(n332), .A2(n333), .Y(n484) );
  NBUFFX2_HVT U331 ( .A(in[4]), .Y(n342) );
  NAND2X0_HVT U332 ( .A1(n508), .A2(n306), .Y(n336) );
  NAND2X0_HVT U333 ( .A1(n509), .A2(n363), .Y(n337) );
  NAND2X0_HVT U334 ( .A1(n336), .A2(n337), .Y(n505) );
  NAND2X0_HVT U335 ( .A1(n496), .A2(n305), .Y(n338) );
  NAND2X0_HVT U336 ( .A1(n489), .A2(n300), .Y(n339) );
  NAND2X0_HVT U337 ( .A1(n339), .A2(n338), .Y(out[6]) );
  NAND2X0_HVT U338 ( .A1(n554), .A2(n363), .Y(n341) );
  NAND2X0_HVT U339 ( .A1(n340), .A2(n341), .Y(n552) );
  NAND2X0_HVT U340 ( .A1(n569), .A2(n305), .Y(n344) );
  NAND2X0_HVT U341 ( .A1(n344), .A2(n343), .Y(out[2]) );
  INVX0_HVT U342 ( .A(n370), .Y(n348) );
  MUX41X1_HVT U343 ( .A1(n645), .A3(n260), .A2(n644), .A4(n422), .S0(n319), 
        .S1(n268), .Y(n584) );
  OR2X1_HVT U344 ( .A1(n346), .A2(n348), .Y(n663) );
  INVX1_HVT U345 ( .A(n381), .Y(n450) );
  NBUFFX2_HVT U346 ( .A(n662), .Y(n381) );
  NBUFFX2_HVT U347 ( .A(n658), .Y(n379) );
  NBUFFX2_HVT U348 ( .A(n662), .Y(n382) );
  NBUFFX2_HVT U349 ( .A(n658), .Y(n380) );
  AND2X1_HVT U350 ( .A1(n657), .A2(n382), .Y(n349) );
  MUX21X1_HVT U351 ( .A1(n432), .A2(n352), .S0(n334), .Y(n471) );
  AND2X1_HVT U352 ( .A1(n382), .A2(n647), .Y(n350) );
  NAND2X0_HVT U353 ( .A1(n367), .A2(n369), .Y(n662) );
  MUX21X1_HVT U354 ( .A1(n450), .A2(n453), .S0(n285), .Y(n629) );
  MUX21X1_HVT U355 ( .A1(n369), .A2(n451), .S0(n298), .Y(n516) );
  MUX21X1_HVT U356 ( .A1(n368), .A2(n450), .S0(n298), .Y(n632) );
  MUX21X1_HVT U357 ( .A1(n368), .A2(n282), .S0(n387), .Y(n619) );
  MUX21X1_HVT U358 ( .A1(n417), .A2(n599), .S0(n355), .Y(n598) );
  MUX21X1_HVT U359 ( .A1(n278), .A2(n316), .S0(n357), .Y(n599) );
  MUX21X1_HVT U360 ( .A1(n604), .A2(n603), .S0(n313), .Y(n601) );
  MUX21X1_HVT U361 ( .A1(n231), .A2(n608), .S0(n365), .Y(n604) );
  MUX21X1_HVT U362 ( .A1(n381), .A2(n380), .S0(n387), .Y(n522) );
  MUX21X1_HVT U363 ( .A1(n282), .A2(n368), .S0(n284), .Y(n465) );
  MUX21X1_HVT U364 ( .A1(n379), .A2(n382), .S0(n297), .Y(n456) );
  MUX21X1_HVT U365 ( .A1(n453), .A2(n368), .S0(n284), .Y(n623) );
  MUX21X1_HVT U366 ( .A1(n405), .A2(n621), .S0(n366), .Y(n554) );
  MUX21X1_HVT U367 ( .A1(n450), .A2(n282), .S0(n385), .Y(n612) );
  MUX21X1_HVT U368 ( .A1(n629), .A2(n350), .S0(n363), .Y(n537) );
  MUX21X1_HVT U369 ( .A1(n447), .A2(n351), .S0(n363), .Y(n540) );
  XOR2X1_HVT U370 ( .A1(n379), .A2(n284), .Y(n614) );
  MUX21X1_HVT U371 ( .A1(n261), .A2(n371), .S0(n385), .Y(n457) );
  XNOR2X1_HVT U372 ( .A1(n381), .A2(n285), .Y(n351) );
  XOR2X1_HVT U373 ( .A1(n661), .A2(n284), .Y(n615) );
  MUX21X1_HVT U374 ( .A1(n368), .A2(n382), .S0(n384), .Y(n464) );
  MUX21X1_HVT U375 ( .A1(n290), .A2(n382), .S0(n384), .Y(n644) );
  MUX21X1_HVT U376 ( .A1(n290), .A2(n368), .S0(n297), .Y(n643) );
  MUX21X1_HVT U377 ( .A1(n369), .A2(n382), .S0(n385), .Y(n559) );
  XOR2X1_HVT U378 ( .A1(n236), .A2(n384), .Y(n625) );
  MUX21X1_HVT U379 ( .A1(n235), .A2(n382), .S0(n387), .Y(n648) );
  MUX21X1_HVT U380 ( .A1(n418), .A2(n606), .S0(n355), .Y(n605) );
  MUX21X1_HVT U381 ( .A1(n419), .A2(n659), .S0(n363), .Y(n606) );
  MUX21X1_HVT U382 ( .A1(n290), .A2(n370), .S0(n285), .Y(n543) );
  MUX21X1_HVT U383 ( .A1(n369), .A2(n378), .S0(n297), .Y(n622) );
  MUX21X1_HVT U384 ( .A1(n367), .A2(n290), .S0(n298), .Y(n459) );
  AND2X1_HVT U385 ( .A1(n298), .A2(n371), .Y(n352) );
  NBUFFX2_HVT U386 ( .A(n392), .Y(n365) );
  NBUFFX2_HVT U387 ( .A(n393), .Y(n364) );
  NBUFFX2_HVT U388 ( .A(n393), .Y(n366) );
  NBUFFX2_HVT U389 ( .A(n346), .Y(n367) );
  MUX21X1_HVT U390 ( .A1(n480), .A2(n439), .S0(n334), .Y(n479) );
  NBUFFX2_HVT U391 ( .A(n663), .Y(n383) );
  NBUFFX2_HVT U392 ( .A(n346), .Y(n368) );
  AND2X1_HVT U393 ( .A1(n282), .A2(n389), .Y(n353) );
  AND2X1_HVT U394 ( .A1(n661), .A2(n389), .Y(n354) );
  NBUFFX2_HVT U395 ( .A(n390), .Y(n362) );
  NBUFFX2_HVT U396 ( .A(n390), .Y(n363) );
  NBUFFX2_HVT U397 ( .A(n454), .Y(n370) );
  XNOR2X1_HVT U398 ( .A1(n395), .A2(n359), .Y(n355) );
  NBUFFX2_HVT U399 ( .A(n390), .Y(n359) );
  NBUFFX2_HVT U400 ( .A(n390), .Y(n361) );
  NBUFFX2_HVT U401 ( .A(n390), .Y(n358) );
  NBUFFX2_HVT U402 ( .A(n390), .Y(n357) );
  NBUFFX2_HVT U403 ( .A(n390), .Y(n360) );
  INVX1_HVT U404 ( .A(n372), .Y(n374) );
  MUX21X1_HVT U405 ( .A1(n528), .A2(n529), .S0(n374), .Y(n527) );
  MUX21X1_HVT U406 ( .A1(n282), .A2(n451), .S0(n296), .Y(n548) );
  MUX21X1_HVT U407 ( .A1(n236), .A2(n272), .S0(n285), .Y(n507) );
  MUX21X1_HVT U408 ( .A1(n347), .A2(n380), .S0(n384), .Y(n460) );
  MUX21X1_HVT U409 ( .A1(n347), .A2(n237), .S0(n284), .Y(n461) );
  MUX21X1_HVT U410 ( .A1(n371), .A2(n347), .S0(n297), .Y(n635) );
  INVX0_HVT U411 ( .A(in[6]), .Y(n454) );
  NBUFFX2_HVT U412 ( .A(in[2]), .Y(n390) );
  MUX21X1_HVT U413 ( .A1(n241), .A2(n347), .S0(n284), .Y(n455) );
  NBUFFX2_HVT U414 ( .A(n646), .Y(n377) );
  NBUFFX2_HVT U415 ( .A(n646), .Y(n378) );
  MUX21X1_HVT U416 ( .A1(n368), .A2(n370), .S0(n384), .Y(n617) );
  MUX21X1_HVT U417 ( .A1(n450), .A2(n370), .S0(n385), .Y(n466) );
  MUX21X1_HVT U418 ( .A1(n450), .A2(n356), .S0(n285), .Y(n530) );
  XOR2X1_HVT U419 ( .A1(n298), .A2(n356), .Y(n613) );
  MUX21X1_HVT U420 ( .A1(n356), .A2(n661), .S0(n284), .Y(n467) );
  MUX21X1_HVT U421 ( .A1(n290), .A2(n356), .S0(n385), .Y(n463) );
  MUX21X1_HVT U422 ( .A1(n367), .A2(n356), .S0(n384), .Y(n458) );
  MUX21X1_HVT U423 ( .A1(n356), .A2(n235), .S0(n384), .Y(n645) );
  MUX21X1_HVT U424 ( .A1(n356), .A2(n241), .S0(n385), .Y(n638) );
  MUX21X1_HVT U425 ( .A1(n380), .A2(n356), .S0(n386), .Y(n633) );
  MUX21X1_HVT U426 ( .A1(n356), .A2(n281), .S0(n297), .Y(n468) );
  INVX0_HVT U427 ( .A(n630), .Y(n397) );
  INVX0_HVT U428 ( .A(n624), .Y(n398) );
  INVX0_HVT U429 ( .A(n564), .Y(n399) );
  INVX0_HVT U430 ( .A(n525), .Y(n400) );
  INVX0_HVT U431 ( .A(n659), .Y(n402) );
  INVX0_HVT U432 ( .A(n656), .Y(n405) );
  INVX0_HVT U433 ( .A(n655), .Y(n406) );
  INVX0_HVT U434 ( .A(n627), .Y(n407) );
  INVX0_HVT U435 ( .A(n649), .Y(n408) );
  INVX0_HVT U436 ( .A(n654), .Y(n409) );
  INVX0_HVT U437 ( .A(n650), .Y(n410) );
  INVX0_HVT U438 ( .A(n648), .Y(n411) );
  INVX0_HVT U439 ( .A(n645), .Y(n413) );
  INVX0_HVT U440 ( .A(n644), .Y(n414) );
  INVX0_HVT U441 ( .A(n643), .Y(n415) );
  INVX0_HVT U442 ( .A(n642), .Y(n416) );
  INVX0_HVT U443 ( .A(n638), .Y(n418) );
  INVX0_HVT U444 ( .A(n637), .Y(n419) );
  INVX0_HVT U445 ( .A(n636), .Y(n420) );
  INVX0_HVT U446 ( .A(n632), .Y(n423) );
  INVX0_HVT U447 ( .A(n625), .Y(n427) );
  INVX0_HVT U448 ( .A(n623), .Y(n428) );
  INVX0_HVT U449 ( .A(n622), .Y(n429) );
  INVX0_HVT U450 ( .A(n617), .Y(n432) );
  INVX0_HVT U451 ( .A(n653), .Y(n434) );
  INVX0_HVT U452 ( .A(n468), .Y(n435) );
  INVX0_HVT U453 ( .A(n467), .Y(n436) );
  INVX0_HVT U454 ( .A(n464), .Y(n439) );
  INVX0_HVT U455 ( .A(n463), .Y(n440) );
  INVX0_HVT U456 ( .A(n461), .Y(n442) );
  INVX0_HVT U457 ( .A(n460), .Y(n443) );
  INVX0_HVT U458 ( .A(n459), .Y(n444) );
  INVX0_HVT U459 ( .A(n458), .Y(n445) );
  INVX0_HVT U460 ( .A(n507), .Y(n446) );
  INVX0_HVT U461 ( .A(n457), .Y(n447) );
  INVX0_HVT U462 ( .A(n456), .Y(n448) );
endmodule

