
module sbox_3 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n142, n210, n211, n212, n213, n216, n217, n218, n219, n227,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600;

  NAND2X0_HVT U4 ( .A1(n309), .A2(n598), .Y(n597) );
  NAND2X0_HVT U5 ( .A1(n317), .A2(n298), .Y(n595) );
  NAND2X0_HVT U13 ( .A1(n587), .A2(n313), .Y(n588) );
  NAND2X0_HVT U15 ( .A1(n598), .A2(n299), .Y(n585) );
  NAND2X0_HVT U21 ( .A1(n309), .A2(n319), .Y(n579) );
  NAND2X0_HVT U24 ( .A1(n305), .A2(n319), .Y(n577) );
  NAND2X0_HVT U33 ( .A1(n377), .A2(n319), .Y(n568) );
  NAND2X0_HVT U35 ( .A1(n303), .A2(n319), .Y(n566) );
  NAND2X0_HVT U42 ( .A1(n317), .A2(n305), .Y(n559) );
  MUX41X1_HVT U51 ( .A1(n366), .A3(n325), .A2(n343), .A4(n344), .S0(n247), 
        .S1(n292), .Y(n551) );
  NAND2X0_HVT U53 ( .A1(n548), .A2(n558), .Y(n549) );
  NAND2X0_HVT U56 ( .A1(n309), .A2(n544), .Y(n545) );
  MUX41X1_HVT U57 ( .A1(n367), .A3(n581), .A2(n545), .A4(n590), .S0(n321), 
        .S1(n292), .Y(n543) );
  NAND2X0_HVT U58 ( .A1(n313), .A2(n598), .Y(n542) );
  MUX41X1_HVT U59 ( .A1(n285), .A3(n542), .A2(n283), .A4(n342), .S0(n247), 
        .S1(n292), .Y(n541) );
  MUX41X1_HVT U61 ( .A1(n282), .A3(n341), .A2(n340), .A4(n299), .S0(n321), 
        .S1(n292), .Y(n539) );
  NAND2X0_HVT U62 ( .A1(n319), .A2(n311), .Y(n538) );
  MUX41X1_HVT U63 ( .A1(n538), .A3(n332), .A2(n361), .A4(n339), .S0(n267), 
        .S1(n292), .Y(n537) );
  AO21X1_HVT U66 ( .A1(n337), .A2(n294), .A3(n360), .Y(n534) );
  MUX41X1_HVT U68 ( .A1(n335), .A3(n534), .A2(n533), .A4(n535), .S0(n286), 
        .S1(n320), .Y(n532) );
  MUX41X1_HVT U69 ( .A1(n532), .A3(n540), .A2(n536), .A4(n546), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n306), .A2(n527), .Y(n528) );
  MUX41X1_HVT U74 ( .A1(n529), .A3(n575), .A2(n528), .A4(n577), .S0(n288), 
        .S1(n267), .Y(n526) );
  MUX41X1_HVT U75 ( .A1(n364), .A3(n369), .A2(n381), .A4(n346), .S0(n286), 
        .S1(n266), .Y(n525) );
  MUX41X1_HVT U77 ( .A1(n592), .A3(n371), .A2(n524), .A4(n370), .S0(n295), 
        .S1(n246), .Y(n523) );
  MUX41X1_HVT U78 ( .A1(n523), .A3(n526), .A2(n525), .A4(n530), .S0(in[0]), 
        .S1(n292), .Y(n522) );
  AND3X1_HVT U80 ( .A1(n310), .A2(n544), .A3(n519), .Y(n520) );
  MUX41X1_HVT U82 ( .A1(n556), .A3(n344), .A2(n326), .A4(n586), .S0(n286), 
        .S1(n321), .Y(n517) );
  AND2X1_HVT U83 ( .A1(n317), .A2(n261), .Y(n516) );
  MUX41X1_HVT U84 ( .A1(n345), .A3(n594), .A2(n584), .A4(n516), .S0(n286), 
        .S1(n267), .Y(n515) );
  NAND2X0_HVT U85 ( .A1(n319), .A2(n380), .Y(n514) );
  MUX41X1_HVT U86 ( .A1(n369), .A3(n514), .A2(n280), .A4(n278), .S0(n286), 
        .S1(n266), .Y(n513) );
  MUX41X1_HVT U87 ( .A1(n513), .A3(n517), .A2(n515), .A4(n518), .S0(n304), 
        .S1(in[5]), .Y(n512) );
  MUX41X1_HVT U90 ( .A1(n555), .A3(n559), .A2(n366), .A4(n511), .S0(n287), 
        .S1(n321), .Y(n510) );
  AO21X1_HVT U93 ( .A1(n297), .A2(n506), .A3(n365), .Y(n507) );
  MUX41X1_HVT U97 ( .A1(n364), .A3(n281), .A2(n317), .A4(n585), .S0(n286), 
        .S1(n321), .Y(n502) );
  NAND2X0_HVT U101 ( .A1(n497), .A2(n496), .Y(n498) );
  MUX41X1_HVT U103 ( .A1(n598), .A3(n336), .A2(n260), .A4(n566), .S0(n286), 
        .S1(n320), .Y(n494) );
  MUX41X1_HVT U105 ( .A1(n348), .A3(n554), .A2(n493), .A4(n363), .S0(n286), 
        .S1(n321), .Y(n492) );
  OA21X1_HVT U109 ( .A1(n354), .A2(n268), .A3(n342), .Y(n489) );
  NAND2X0_HVT U110 ( .A1(n310), .A2(n487), .Y(n488) );
  AND2X1_HVT U115 ( .A1(n317), .A2(n299), .Y(n482) );
  MUX41X1_HVT U116 ( .A1(n588), .A3(n482), .A2(n346), .A4(n570), .S0(n287), 
        .S1(n247), .Y(n481) );
  NAND2X0_HVT U123 ( .A1(n473), .A2(n472), .Y(n474) );
  MUX41X1_HVT U125 ( .A1(n579), .A3(n285), .A2(n335), .A4(n373), .S0(n287), 
        .S1(n247), .Y(n470) );
  MUX41X1_HVT U131 ( .A1(n465), .A3(n467), .A2(n466), .A4(n468), .S0(n294), 
        .S1(n321), .Y(n464) );
  MUX41X1_HVT U136 ( .A1(n278), .A3(n568), .A2(n374), .A4(n565), .S0(n287), 
        .S1(n320), .Y(n461) );
  MUX41X1_HVT U139 ( .A1(n459), .A3(n235), .A2(n461), .A4(n462), .S0(n304), 
        .S1(in[5]), .Y(n458) );
  AND2X1_HVT U140 ( .A1(n307), .A2(n249), .Y(n457) );
  NAND2X0_HVT U146 ( .A1(n317), .A2(n313), .Y(n527) );
  MUX41X1_HVT U153 ( .A1(n488), .A3(n282), .A2(n599), .A4(n328), .S0(n287), 
        .S1(n321), .Y(n445) );
  AND2X1_HVT U154 ( .A1(n297), .A2(n305), .Y(n444) );
  NAND2X0_HVT U158 ( .A1(n317), .A2(n380), .Y(n440) );
  MUX41X1_HVT U159 ( .A1(n588), .A3(n300), .A2(n440), .A4(n334), .S0(n246), 
        .S1(n267), .Y(n439) );
  MUX41X1_HVT U160 ( .A1(n439), .A3(n445), .A2(n441), .A4(n446), .S0(n304), 
        .S1(n293), .Y(n438) );
  AND2X1_HVT U162 ( .A1(n594), .A2(n527), .Y(n436) );
  MUX41X1_HVT U163 ( .A1(n341), .A3(n436), .A2(n279), .A4(n437), .S0(n289), 
        .S1(n320), .Y(n435) );
  MUX41X1_HVT U165 ( .A1(n579), .A3(n349), .A2(n555), .A4(n434), .S0(n267), 
        .S1(n289), .Y(n433) );
  NAND2X0_HVT U166 ( .A1(n313), .A2(n544), .Y(n432) );
  NAND2X0_HVT U167 ( .A1(n381), .A2(n319), .Y(n431) );
  MUX41X1_HVT U168 ( .A1(n367), .A3(n591), .A2(n431), .A4(n432), .S0(n290), 
        .S1(n266), .Y(n430) );
  MUX41X1_HVT U172 ( .A1(n427), .A3(n433), .A2(n430), .A4(n435), .S0(in[0]), 
        .S1(n293), .Y(n426) );
  NAND2X0_HVT U174 ( .A1(n317), .A2(n594), .Y(n587) );
  MUX41X1_HVT U176 ( .A1(n301), .A3(n425), .A2(n372), .A4(n587), .S0(n267), 
        .S1(n289), .Y(n424) );
  NAND2X0_HVT U177 ( .A1(n317), .A2(n302), .Y(n423) );
  MUX41X1_HVT U178 ( .A1(n583), .A3(n423), .A2(n375), .A4(n563), .S0(n288), 
        .S1(n267), .Y(n422) );
  MUX41X1_HVT U179 ( .A1(n573), .A3(n376), .A2(n330), .A4(n375), .S0(n246), 
        .S1(n266), .Y(n421) );
  MUX41X1_HVT U180 ( .A1(n333), .A3(n592), .A2(n588), .A4(n277), .S0(n295), 
        .S1(n246), .Y(n420) );
  MUX41X1_HVT U181 ( .A1(n420), .A3(n422), .A2(n421), .A4(n424), .S0(n304), 
        .S1(n293), .Y(n419) );
  MUX41X1_HVT U182 ( .A1(n356), .A3(n308), .A2(n358), .A4(n347), .S0(n266), 
        .S1(n291), .Y(n418) );
  MUX41X1_HVT U189 ( .A1(n412), .A3(n587), .A2(n413), .A4(n363), .S0(n295), 
        .S1(n288), .Y(n411) );
  MUX41X1_HVT U190 ( .A1(n411), .A3(n414), .A2(n415), .A4(n418), .S0(n293), 
        .S1(in[0]), .Y(n410) );
  MUX41X1_HVT U194 ( .A1(n560), .A3(n574), .A2(n233), .A4(n307), .S0(n295), 
        .S1(n290), .Y(n407) );
  MUX41X1_HVT U195 ( .A1(n594), .A3(n368), .A2(n312), .A4(n564), .S0(n288), 
        .S1(n267), .Y(n406) );
  AO21X1_HVT U197 ( .A1(n280), .A2(n296), .A3(n365), .Y(n404) );
  MUX41X1_HVT U199 ( .A1(n403), .A3(n407), .A2(n406), .A4(n408), .S0(in[0]), 
        .S1(n293), .Y(n402) );
  MUX41X1_HVT U203 ( .A1(n565), .A3(n357), .A2(n589), .A4(n569), .S0(n246), 
        .S1(n320), .Y(n398) );
  MUX41X1_HVT U204 ( .A1(n545), .A3(n588), .A2(n353), .A4(n578), .S0(n288), 
        .S1(n266), .Y(n397) );
  MUX41X1_HVT U205 ( .A1(n261), .A3(n598), .A2(n376), .A4(n351), .S0(n291), 
        .S1(n267), .Y(n396) );
  NAND2X0_HVT U208 ( .A1(n317), .A2(n309), .Y(n487) );
  NAND2X0_HVT U212 ( .A1(n317), .A2(n306), .Y(n544) );
  NAND2X0_HVT U214 ( .A1(n594), .A2(n319), .Y(n394) );
  NAND2X0_HVT U215 ( .A1(n487), .A2(n307), .Y(n393) );
  NAND2X0_HVT U218 ( .A1(n378), .A2(n317), .Y(n447) );
  NAND2X0_HVT U220 ( .A1(n296), .A2(n394), .Y(n519) );
  INVX2_HVT U1 ( .A(n318), .Y(n250) );
  MUX21X2_HVT U2 ( .A1(n350), .A2(n463), .S0(n290), .Y(n462) );
  NAND2X2_HVT U3 ( .A1(n258), .A2(n259), .Y(out[4]) );
  NAND2X1_HVT U6 ( .A1(n453), .A2(n23), .Y(n48) );
  NAND2X0_HVT U7 ( .A1(n454), .A2(n210), .Y(n142) );
  NAND2X0_HVT U8 ( .A1(n48), .A2(n142), .Y(n452) );
  IBUFFX2_HVT U9 ( .A(n210), .Y(n23) );
  IBUFFX2_HVT U10 ( .A(n290), .Y(n210) );
  MUX21X2_HVT U11 ( .A1(n331), .A2(n572), .S0(n257), .Y(n454) );
  NAND2X1_HVT U12 ( .A1(n317), .A2(n310), .Y(n598) );
  MUX21X1_HVT U14 ( .A1(n547), .A2(n551), .S0(n290), .Y(n546) );
  INVX2_HVT U16 ( .A(n248), .Y(n317) );
  MUX21X1_HVT U17 ( .A1(n400), .A2(n401), .S0(n289), .Y(n399) );
  MUX21X1_HVT U18 ( .A1(n597), .A2(n460), .S0(n268), .Y(n459) );
  MUX21X2_HVT U19 ( .A1(n410), .A2(n419), .S0(in[6]), .Y(out[6]) );
  MUX21X1_HVT U20 ( .A1(n474), .A2(n475), .S0(n257), .Y(n471) );
  XNOR2X1_HVT U22 ( .A1(n271), .A2(n249), .Y(n211) );
  IBUFFX16_HVT U23 ( .A(n211), .Y(n555) );
  MUX41X1_HVT U25 ( .A1(n562), .A3(n281), .A2(n555), .A4(n527), .S0(n212), 
        .S1(n266), .Y(n414) );
  IBUFFX16_HVT U26 ( .A(n291), .Y(n212) );
  INVX1_HVT U27 ( .A(n271), .Y(n594) );
  MUX41X1_HVT U28 ( .A1(n484), .A3(n490), .A2(n486), .A4(n489), .S0(n213), 
        .S1(n216), .Y(n483) );
  IBUFFX16_HVT U29 ( .A(n269), .Y(n213) );
  IBUFFX16_HVT U30 ( .A(n257), .Y(n216) );
  MUX21X2_HVT U31 ( .A1(n508), .A2(n507), .S0(n217), .Y(n505) );
  IBUFFX16_HVT U32 ( .A(n291), .Y(n217) );
  MUX41X1_HVT U34 ( .A1(n505), .A3(n502), .A2(n510), .A4(n503), .S0(n218), 
        .S1(n219), .Y(n501) );
  IBUFFX16_HVT U36 ( .A(n304), .Y(n218) );
  IBUFFX16_HVT U37 ( .A(n269), .Y(n219) );
  MUX21X1_HVT U38 ( .A1(n537), .A2(n539), .S0(n289), .Y(n536) );
  MUX41X1_HVT U39 ( .A1(n483), .A3(n469), .A2(n477), .A4(n464), .S0(n227), 
        .S1(n231), .Y(out[3]) );
  IBUFFX16_HVT U40 ( .A(in[6]), .Y(n227) );
  IBUFFX16_HVT U41 ( .A(in[0]), .Y(n231) );
  MUX21X1_HVT U43 ( .A1(n470), .A2(n471), .S0(n294), .Y(n469) );
  INVX1_HVT U44 ( .A(in[1]), .Y(n232) );
  INVX0_HVT U45 ( .A(in[1]), .Y(n248) );
  INVX1_HVT U46 ( .A(n250), .Y(n319) );
  MUX21X1_HVT U47 ( .A1(n234), .A2(n271), .S0(n232), .Y(n233) );
  IBUFFX16_HVT U48 ( .A(n378), .Y(n234) );
  MUX41X1_HVT U49 ( .A1(n574), .A3(n595), .A2(n236), .A4(n233), .S0(n237), 
        .S1(n238), .Y(n235) );
  IBUFFX16_HVT U50 ( .A(n307), .Y(n236) );
  IBUFFX16_HVT U52 ( .A(n246), .Y(n237) );
  IBUFFX16_HVT U54 ( .A(n247), .Y(n238) );
  INVX1_HVT U55 ( .A(n248), .Y(n245) );
  MUX21X2_HVT U60 ( .A1(n491), .A2(n501), .S0(n239), .Y(out[2]) );
  IBUFFX16_HVT U64 ( .A(n263), .Y(n239) );
  MUX21X2_HVT U65 ( .A1(n557), .A2(n531), .S0(n289), .Y(n530) );
  MUX21X2_HVT U67 ( .A1(n380), .A2(n368), .S0(n297), .Y(n531) );
  INVX2_HVT U70 ( .A(n232), .Y(n315) );
  NBUFFX2_HVT U71 ( .A(n316), .Y(n240) );
  NBUFFX2_HVT U72 ( .A(n316), .Y(n241) );
  IBUFFX2_HVT U76 ( .A(n318), .Y(n316) );
  INVX0_HVT U79 ( .A(n304), .Y(n262) );
  INVX0_HVT U81 ( .A(n260), .Y(n572) );
  INVX0_HVT U88 ( .A(n242), .Y(n565) );
  INVX0_HVT U89 ( .A(n323), .Y(n267) );
  INVX1_HVT U91 ( .A(in[5]), .Y(n269) );
  INVX1_HVT U92 ( .A(n297), .Y(n257) );
  INVX1_HVT U94 ( .A(n295), .Y(n243) );
  INVX1_HVT U95 ( .A(in[7]), .Y(n324) );
  INVX1_HVT U96 ( .A(n324), .Y(n247) );
  INVX1_HVT U98 ( .A(n303), .Y(n261) );
  INVX0_HVT U99 ( .A(in[6]), .Y(n263) );
  INVX0_HVT U100 ( .A(n288), .Y(n268) );
  INVX1_HVT U102 ( .A(n272), .Y(n246) );
  INVX0_HVT U104 ( .A(n287), .Y(n272) );
  MUX21X1_HVT U106 ( .A1(n303), .A2(n298), .S0(n232), .Y(n409) );
  MUX41X1_HVT U107 ( .A1(n409), .A3(n552), .A2(n566), .A4(n559), .S0(n268), 
        .S1(n323), .Y(n408) );
  IBUFFX2_HVT U108 ( .A(n323), .Y(n321) );
  INVX2_HVT U111 ( .A(n249), .Y(n314) );
  INVX1_HVT U112 ( .A(n245), .Y(n249) );
  MUX21X1_HVT U113 ( .A1(n312), .A2(n302), .S0(n318), .Y(n242) );
  INVX1_HVT U114 ( .A(n500), .Y(n275) );
  INVX0_HVT U117 ( .A(n273), .Y(n499) );
  MUX21X2_HVT U118 ( .A1(n371), .A2(n563), .S0(n243), .Y(n442) );
  MUX21X2_HVT U119 ( .A1(n442), .A2(n443), .S0(n291), .Y(n441) );
  MUX21X1_HVT U120 ( .A1(n274), .A2(n275), .S0(n244), .Y(n273) );
  IBUFFX16_HVT U121 ( .A(n276), .Y(n244) );
  OA21X1_HVT U122 ( .A1(n561), .A2(n257), .A3(n447), .Y(n448) );
  INVX1_HVT U124 ( .A(n561), .Y(n357) );
  INVX1_HVT U126 ( .A(in[1]), .Y(n318) );
  OA21X1_HVT U127 ( .A1(n567), .A2(n257), .A3(n345), .Y(n416) );
  OA21X1_HVT U128 ( .A1(n329), .A2(n324), .A3(n570), .Y(n453) );
  INVX1_HVT U129 ( .A(n570), .Y(n351) );
  IBUFFX2_HVT U130 ( .A(n578), .Y(n345) );
  NAND2X0_HVT U132 ( .A1(n488), .A2(n246), .Y(n251) );
  NAND2X0_HVT U133 ( .A1(n570), .A2(n268), .Y(n252) );
  NAND2X0_HVT U134 ( .A1(n251), .A2(n252), .Y(n486) );
  MUX21X1_HVT U135 ( .A1(n312), .A2(n306), .S0(n240), .Y(n570) );
  MUX21X2_HVT U137 ( .A1(n578), .A2(n356), .S0(n296), .Y(n460) );
  IBUFFX2_HVT U138 ( .A(n590), .Y(n337) );
  NAND2X0_HVT U141 ( .A1(n395), .A2(n263), .Y(n253) );
  NAND2X0_HVT U142 ( .A1(n402), .A2(n270), .Y(n254) );
  NAND2X0_HVT U143 ( .A1(n253), .A2(n254), .Y(out[7]) );
  INVX0_HVT U144 ( .A(n263), .Y(n270) );
  NAND2X0_HVT U145 ( .A1(n478), .A2(n269), .Y(n255) );
  NAND2X0_HVT U147 ( .A1(n481), .A2(n294), .Y(n256) );
  NAND2X0_HVT U148 ( .A1(n255), .A2(n256), .Y(n477) );
  NAND2X0_HVT U149 ( .A1(n450), .A2(n263), .Y(n258) );
  NAND2X0_HVT U150 ( .A1(n458), .A2(in[6]), .Y(n259) );
  OA21X2_HVT U151 ( .A1(n283), .A2(n243), .A3(n570), .Y(n428) );
  MUX21X1_HVT U152 ( .A1(n261), .A2(n308), .S0(n250), .Y(n260) );
  MUX21X2_HVT U155 ( .A1(n541), .A2(n543), .S0(n289), .Y(n540) );
  MUX41X1_HVT U156 ( .A1(n399), .A3(n397), .A2(n398), .A4(n396), .S0(n262), 
        .S1(n269), .Y(n395) );
  MUX21X1_HVT U157 ( .A1(n351), .A2(n586), .S0(n291), .Y(n500) );
  MUX21X2_HVT U161 ( .A1(n584), .A2(n277), .S0(n295), .Y(n401) );
  OA21X1_HVT U164 ( .A1(n593), .A2(n324), .A3(n355), .Y(n400) );
  NAND2X0_HVT U169 ( .A1(n512), .A2(n263), .Y(n264) );
  NAND2X0_HVT U170 ( .A1(n522), .A2(in[6]), .Y(n265) );
  NAND2X0_HVT U171 ( .A1(n264), .A2(n265), .Y(out[1]) );
  INVX0_HVT U173 ( .A(n323), .Y(n266) );
  INVX1_HVT U175 ( .A(in[7]), .Y(n323) );
  INVX0_HVT U183 ( .A(n323), .Y(n320) );
  MUX41X1_HVT U184 ( .A1(n452), .A3(n456), .A2(n451), .A4(n455), .S0(n304), 
        .S1(n269), .Y(n450) );
  MUX21X2_HVT U185 ( .A1(n327), .A2(n476), .S0(n288), .Y(n475) );
  MUX41X1_HVT U186 ( .A1(n555), .A3(n364), .A2(n527), .A4(n374), .S0(n268), 
        .S1(n243), .Y(n451) );
  MUX41X1_HVT U187 ( .A1(n281), .A3(n326), .A2(n504), .A4(n368), .S0(n268), 
        .S1(n266), .Y(n503) );
  INVX0_HVT U188 ( .A(n324), .Y(n322) );
  MUX41X1_HVT U191 ( .A1(n494), .A3(n499), .A2(n492), .A4(n495), .S0(in[0]), 
        .S1(n269), .Y(n491) );
  AO21X2_HVT U192 ( .A1(n318), .A2(n378), .A3(n324), .Y(n497) );
  MUX21X1_HVT U193 ( .A1(n299), .A2(n298), .S0(n250), .Y(n584) );
  NBUFFX2_HVT U196 ( .A(n271), .Y(n299) );
  MUX21X2_HVT U198 ( .A1(n426), .A2(n438), .S0(in[6]), .Y(out[5]) );
  NBUFFX2_HVT U200 ( .A(n382), .Y(n302) );
  NBUFFX2_HVT U201 ( .A(n382), .Y(n303) );
  XOR2X1_HVT U202 ( .A1(n257), .A2(n574), .Y(n557) );
  XNOR2X2_HVT U206 ( .A1(n301), .A2(in[3]), .Y(n271) );
  AND3X2_HVT U207 ( .A1(n290), .A2(n319), .A3(n261), .Y(n467) );
  AO21X2_HVT U209 ( .A1(n291), .A2(n306), .A3(n594), .Y(n479) );
  MUX41X1_HVT U210 ( .A1(n306), .A3(n362), .A2(n299), .A4(n345), .S0(n272), 
        .S1(n324), .Y(n455) );
  IBUFFX16_HVT U211 ( .A(n282), .Y(n274) );
  XNOR2X1_HVT U213 ( .A1(n290), .A2(n320), .Y(n276) );
  MUX41X1_HVT U216 ( .A1(n352), .A3(n457), .A2(n355), .A4(n576), .S0(n272), 
        .S1(n243), .Y(n456) );
  XOR2X1_HVT U217 ( .A1(n319), .A2(n272), .Y(n553) );
  MUX21X2_HVT U219 ( .A1(n485), .A2(n311), .S0(n553), .Y(n484) );
  INVX0_HVT U221 ( .A(in[3]), .Y(n379) );
  INVX1_HVT U222 ( .A(n308), .Y(n377) );
  NBUFFX2_HVT U223 ( .A(n271), .Y(n300) );
  AND2X1_HVT U224 ( .A1(n300), .A2(n544), .Y(n277) );
  MUX21X1_HVT U225 ( .A1(n279), .A2(n340), .S0(n287), .Y(n466) );
  NBUFFX2_HVT U226 ( .A(n596), .Y(n308) );
  INVX1_HVT U227 ( .A(n599), .Y(n381) );
  MUX21X1_HVT U228 ( .A1(n377), .A2(n380), .S0(n294), .Y(n548) );
  NBUFFX2_HVT U229 ( .A(n596), .Y(n309) );
  MUX21X1_HVT U230 ( .A1(n336), .A2(n378), .S0(n294), .Y(n533) );
  AND2X1_HVT U231 ( .A1(n310), .A2(n527), .Y(n278) );
  MUX21X1_HVT U232 ( .A1(n300), .A2(n380), .S0(n317), .Y(n593) );
  MUX21X1_HVT U233 ( .A1(n310), .A2(n299), .S0(n241), .Y(n560) );
  MUX21X1_HVT U234 ( .A1(n309), .A2(n594), .S0(n240), .Y(n564) );
  MUX21X1_HVT U235 ( .A1(n299), .A2(n303), .S0(n315), .Y(n496) );
  MUX21X1_HVT U236 ( .A1(n377), .A2(n381), .S0(n240), .Y(n425) );
  MUX21X1_HVT U237 ( .A1(n299), .A2(n377), .S0(n315), .Y(n504) );
  MUX21X1_HVT U238 ( .A1(n381), .A2(n380), .S0(n250), .Y(n574) );
  MUX21X1_HVT U239 ( .A1(n380), .A2(n377), .S0(n240), .Y(n563) );
  MUX21X1_HVT U240 ( .A1(n594), .A2(n381), .S0(n245), .Y(n576) );
  MUX21X1_HVT U241 ( .A1(n298), .A2(n381), .S0(n240), .Y(n561) );
  NAND2X0_HVT U242 ( .A1(n301), .A2(n379), .Y(n596) );
  MUX21X1_HVT U243 ( .A1(n380), .A2(n299), .S0(n315), .Y(n437) );
  MUX21X1_HVT U244 ( .A1(n309), .A2(n307), .S0(n241), .Y(n511) );
  MUX21X1_HVT U245 ( .A1(n594), .A2(n303), .S0(n241), .Y(n524) );
  INVX1_HVT U246 ( .A(n591), .Y(n378) );
  INVX1_HVT U247 ( .A(n312), .Y(n380) );
  MUX21X1_HVT U248 ( .A1(n380), .A2(n298), .S0(n240), .Y(n567) );
  MUX21X1_HVT U249 ( .A1(n373), .A2(n307), .S0(n296), .Y(n463) );
  MUX21X1_HVT U250 ( .A1(n479), .A2(n480), .S0(n296), .Y(n478) );
  MUX21X1_HVT U251 ( .A1(n328), .A2(n353), .S0(n287), .Y(n480) );
  NBUFFX2_HVT U252 ( .A(n599), .Y(n310) );
  XOR2X1_HVT U253 ( .A1(n311), .A2(n314), .Y(n552) );
  MUX21X1_HVT U254 ( .A1(n377), .A2(n302), .S0(n314), .Y(n386) );
  MUX21X1_HVT U255 ( .A1(n298), .A2(n594), .S0(n315), .Y(n388) );
  MUX21X1_HVT U256 ( .A1(n309), .A2(n298), .S0(n250), .Y(n589) );
  MUX21X1_HVT U257 ( .A1(n302), .A2(n298), .S0(n315), .Y(n476) );
  XOR2X1_HVT U258 ( .A1(n314), .A2(n378), .Y(n556) );
  MUX21X1_HVT U259 ( .A1(n298), .A2(n313), .S0(n315), .Y(n412) );
  MUX21X1_HVT U260 ( .A1(n312), .A2(n310), .S0(n315), .Y(n413) );
  MUX21X1_HVT U261 ( .A1(n378), .A2(n377), .S0(n245), .Y(n582) );
  MUX21X1_HVT U262 ( .A1(n311), .A2(n306), .S0(n250), .Y(n586) );
  MUX21X1_HVT U263 ( .A1(n308), .A2(n313), .S0(n314), .Y(n506) );
  MUX21X1_HVT U264 ( .A1(n298), .A2(n380), .S0(n250), .Y(n590) );
  NBUFFX2_HVT U265 ( .A(n599), .Y(n311) );
  MUX21X1_HVT U266 ( .A1(n306), .A2(n298), .S0(n315), .Y(n390) );
  MUX21X1_HVT U267 ( .A1(n311), .A2(n302), .S0(n315), .Y(n392) );
  XNOR2X1_HVT U268 ( .A1(n308), .A2(n314), .Y(n279) );
  XNOR2X1_HVT U269 ( .A1(n312), .A2(n314), .Y(n280) );
  AND2X1_HVT U270 ( .A1(n317), .A2(n381), .Y(n281) );
  MUX21X1_HVT U271 ( .A1(n310), .A2(n309), .S0(n314), .Y(n385) );
  AND2X1_HVT U272 ( .A1(n313), .A2(n487), .Y(n282) );
  MUX21X1_HVT U273 ( .A1(n307), .A2(n302), .S0(n241), .Y(n529) );
  MUX21X1_HVT U274 ( .A1(n307), .A2(n313), .S0(n290), .Y(n473) );
  XOR2X1_HVT U275 ( .A1(n301), .A2(n314), .Y(n575) );
  NBUFFX2_HVT U276 ( .A(n322), .Y(n295) );
  NBUFFX2_HVT U277 ( .A(n322), .Y(n296) );
  NBUFFX2_HVT U278 ( .A(n379), .Y(n298) );
  NBUFFX2_HVT U279 ( .A(n322), .Y(n297) );
  NBUFFX2_HVT U280 ( .A(in[2]), .Y(n287) );
  NBUFFX2_HVT U281 ( .A(in[5]), .Y(n294) );
  NBUFFX2_HVT U282 ( .A(in[2]), .Y(n289) );
  NBUFFX2_HVT U283 ( .A(in[2]), .Y(n288) );
  NBUFFX2_HVT U284 ( .A(in[5]), .Y(n293) );
  NBUFFX2_HVT U285 ( .A(in[2]), .Y(n290) );
  NBUFFX2_HVT U286 ( .A(in[2]), .Y(n291) );
  NBUFFX2_HVT U287 ( .A(in[5]), .Y(n292) );
  NBUFFX2_HVT U288 ( .A(n291), .Y(n286) );
  NBUFFX2_HVT U289 ( .A(n382), .Y(n301) );
  MUX21X1_HVT U290 ( .A1(n300), .A2(n305), .S0(n250), .Y(n578) );
  MUX21X1_HVT U291 ( .A1(n498), .A2(n350), .S0(n290), .Y(n495) );
  MUX21X1_HVT U292 ( .A1(n416), .A2(n417), .S0(n289), .Y(n415) );
  MUX21X1_HVT U293 ( .A1(n514), .A2(n305), .S0(n296), .Y(n417) );
  XOR2X1_HVT U294 ( .A1(n314), .A2(n305), .Y(n554) );
  MUX21X1_HVT U295 ( .A1(n306), .A2(n300), .S0(n241), .Y(n493) );
  NAND2X0_HVT U296 ( .A1(in[3]), .A2(n303), .Y(n599) );
  MUX21X1_HVT U297 ( .A1(n521), .A2(n520), .S0(n291), .Y(n518) );
  MUX21X1_HVT U298 ( .A1(n580), .A2(n307), .S0(n297), .Y(n521) );
  AND2X1_HVT U299 ( .A1(n300), .A2(n319), .Y(n283) );
  NBUFFX2_HVT U300 ( .A(n600), .Y(n312) );
  MUX21X1_HVT U301 ( .A1(n305), .A2(n377), .S0(n240), .Y(n562) );
  MUX21X1_HVT U302 ( .A1(n448), .A2(n449), .S0(n291), .Y(n446) );
  MUX21X1_HVT U303 ( .A1(n370), .A2(n378), .S0(n296), .Y(n449) );
  MUX21X1_HVT U304 ( .A1(n429), .A2(n428), .S0(n290), .Y(n427) );
  MUX21X1_HVT U305 ( .A1(n307), .A2(n368), .S0(n297), .Y(n429) );
  MUX21X1_HVT U306 ( .A1(n583), .A2(n352), .S0(n288), .Y(n465) );
  MUX21X1_HVT U307 ( .A1(n378), .A2(n381), .S0(n315), .Y(n434) );
  MUX21X1_HVT U308 ( .A1(n381), .A2(n305), .S0(n250), .Y(n581) );
  MUX21X1_HVT U309 ( .A1(n242), .A2(n598), .S0(n288), .Y(n490) );
  MUX21X1_HVT U310 ( .A1(n549), .A2(n550), .S0(n295), .Y(n547) );
  MUX21X1_HVT U311 ( .A1(n305), .A2(n566), .S0(n294), .Y(n550) );
  XOR2X1_HVT U312 ( .A1(n314), .A2(n293), .Y(n558) );
  MUX21X1_HVT U313 ( .A1(n598), .A2(n249), .S0(n289), .Y(n472) );
  NBUFFX2_HVT U314 ( .A(n591), .Y(n306) );
  MUX21X1_HVT U315 ( .A1(n444), .A2(n311), .S0(n284), .Y(n443) );
  MUX21X1_HVT U316 ( .A1(n359), .A2(n375), .S0(n296), .Y(n405) );
  MUX21X1_HVT U317 ( .A1(n305), .A2(n378), .S0(n315), .Y(n389) );
  MUX21X1_HVT U318 ( .A1(n571), .A2(n393), .S0(n295), .Y(n387) );
  MUX21X1_HVT U319 ( .A1(n309), .A2(n305), .S0(n245), .Y(n592) );
  MUX21X1_HVT U320 ( .A1(n338), .A2(n319), .S0(n294), .Y(n535) );
  NBUFFX2_HVT U321 ( .A(n600), .Y(n313) );
  MUX21X1_HVT U322 ( .A1(n348), .A2(n571), .S0(n288), .Y(n468) );
  MUX21X1_HVT U323 ( .A1(n311), .A2(n509), .S0(n284), .Y(n508) );
  MUX21X1_HVT U324 ( .A1(n305), .A2(n302), .S0(n297), .Y(n509) );
  NBUFFX2_HVT U325 ( .A(n591), .Y(n307) );
  XNOR2X1_HVT U326 ( .A1(n324), .A2(n314), .Y(n284) );
  AND2X1_HVT U327 ( .A1(n298), .A2(n319), .Y(n285) );
  MUX21X1_HVT U328 ( .A1(n405), .A2(n404), .S0(n289), .Y(n403) );
  INVX0_HVT U329 ( .A(in[4]), .Y(n382) );
  MUX21X1_HVT U330 ( .A1(n377), .A2(n261), .S0(n241), .Y(n569) );
  NAND2X0_HVT U331 ( .A1(in[4]), .A2(n379), .Y(n591) );
  NAND2X0_HVT U332 ( .A1(in[3]), .A2(in[4]), .Y(n600) );
  MUX21X1_HVT U333 ( .A1(n261), .A2(n594), .S0(n315), .Y(n391) );
  MUX21X1_HVT U334 ( .A1(n261), .A2(n378), .S0(n317), .Y(n583) );
  MUX21X1_HVT U335 ( .A1(n261), .A2(n311), .S0(n245), .Y(n580) );
  MUX21X1_HVT U336 ( .A1(n261), .A2(n306), .S0(n315), .Y(n384) );
  MUX21X1_HVT U337 ( .A1(n261), .A2(n313), .S0(n241), .Y(n383) );
  MUX21X1_HVT U338 ( .A1(n313), .A2(n261), .S0(n245), .Y(n573) );
  MUX21X1_HVT U339 ( .A1(n305), .A2(n261), .S0(n287), .Y(n485) );
  MUX21X1_HVT U340 ( .A1(n298), .A2(n261), .S0(n250), .Y(n571) );
  NBUFFX2_HVT U341 ( .A(in[3]), .Y(n305) );
  NBUFFX2_HVT U342 ( .A(in[0]), .Y(n304) );
  INVX0_HVT U343 ( .A(n579), .Y(n325) );
  INVX0_HVT U344 ( .A(n577), .Y(n326) );
  INVX0_HVT U345 ( .A(n568), .Y(n327) );
  INVX0_HVT U346 ( .A(n566), .Y(n328) );
  INVX0_HVT U347 ( .A(n431), .Y(n329) );
  INVX0_HVT U348 ( .A(n394), .Y(n330) );
  INVX0_HVT U349 ( .A(n598), .Y(n331) );
  INVX0_HVT U350 ( .A(n585), .Y(n332) );
  INVX0_HVT U351 ( .A(n597), .Y(n333) );
  INVX0_HVT U352 ( .A(n595), .Y(n334) );
  INVX0_HVT U353 ( .A(n593), .Y(n335) );
  INVX0_HVT U354 ( .A(n592), .Y(n336) );
  INVX0_HVT U355 ( .A(n589), .Y(n338) );
  INVX0_HVT U356 ( .A(n586), .Y(n339) );
  INVX0_HVT U357 ( .A(n584), .Y(n340) );
  INVX0_HVT U358 ( .A(n583), .Y(n341) );
  INVX0_HVT U359 ( .A(n582), .Y(n342) );
  INVX0_HVT U360 ( .A(n581), .Y(n343) );
  INVX0_HVT U361 ( .A(n580), .Y(n344) );
  INVX0_HVT U362 ( .A(n576), .Y(n346) );
  INVX0_HVT U363 ( .A(n575), .Y(n347) );
  INVX0_HVT U364 ( .A(n573), .Y(n348) );
  INVX0_HVT U365 ( .A(n571), .Y(n349) );
  INVX0_HVT U366 ( .A(n387), .Y(n350) );
  INVX0_HVT U367 ( .A(n569), .Y(n352) );
  INVX0_HVT U368 ( .A(n567), .Y(n353) );
  INVX0_HVT U369 ( .A(n564), .Y(n354) );
  INVX0_HVT U370 ( .A(n563), .Y(n355) );
  INVX0_HVT U371 ( .A(n562), .Y(n356) );
  INVX0_HVT U372 ( .A(n560), .Y(n358) );
  INVX0_HVT U373 ( .A(n559), .Y(n359) );
  INVX0_HVT U374 ( .A(n527), .Y(n360) );
  INVX0_HVT U375 ( .A(n588), .Y(n361) );
  INVX0_HVT U376 ( .A(n487), .Y(n362) );
  INVX0_HVT U377 ( .A(n393), .Y(n363) );
  INVX0_HVT U378 ( .A(n544), .Y(n364) );
  INVX0_HVT U379 ( .A(n447), .Y(n365) );
  INVX0_HVT U380 ( .A(n392), .Y(n366) );
  INVX0_HVT U381 ( .A(n391), .Y(n367) );
  INVX0_HVT U382 ( .A(n390), .Y(n368) );
  INVX0_HVT U383 ( .A(n389), .Y(n369) );
  INVX0_HVT U384 ( .A(n388), .Y(n370) );
  INVX0_HVT U385 ( .A(n506), .Y(n371) );
  INVX0_HVT U386 ( .A(n496), .Y(n372) );
  INVX0_HVT U387 ( .A(n386), .Y(n373) );
  INVX0_HVT U388 ( .A(n385), .Y(n374) );
  INVX0_HVT U389 ( .A(n384), .Y(n375) );
  INVX0_HVT U390 ( .A(n383), .Y(n376) );
endmodule

