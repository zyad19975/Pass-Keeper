
module sbox_15 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n50, n168, n210, n211, n212, n213, n216, n217, n218, n219,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582;

  NAND2X0_HVT U3 ( .A1(n294), .A2(n288), .Y(n580) );
  NAND2X0_HVT U4 ( .A1(n287), .A2(n241), .Y(n579) );
  NAND2X0_HVT U5 ( .A1(n218), .A2(n276), .Y(n577) );
  NAND2X0_HVT U13 ( .A1(n569), .A2(n289), .Y(n570) );
  NAND2X0_HVT U15 ( .A1(n239), .A2(n278), .Y(n567) );
  NAND2X0_HVT U21 ( .A1(n287), .A2(n296), .Y(n561) );
  NAND2X0_HVT U24 ( .A1(n284), .A2(n296), .Y(n559) );
  NAND2X0_HVT U33 ( .A1(n359), .A2(n296), .Y(n550) );
  NAND2X0_HVT U35 ( .A1(n282), .A2(n296), .Y(n548) );
  NAND2X0_HVT U42 ( .A1(n294), .A2(n284), .Y(n541) );
  MUX41X1_HVT U51 ( .A1(n347), .A3(n305), .A2(n322), .A4(n323), .S0(n302), 
        .S1(n298), .Y(n534) );
  NAND2X0_HVT U53 ( .A1(n531), .A2(n540), .Y(n532) );
  NAND2X0_HVT U56 ( .A1(n287), .A2(n527), .Y(n528) );
  MUX41X1_HVT U57 ( .A1(n348), .A3(n563), .A2(n528), .A4(n572), .S0(n302), 
        .S1(n298), .Y(n526) );
  NAND2X0_HVT U58 ( .A1(n289), .A2(n240), .Y(n525) );
  MUX41X1_HVT U59 ( .A1(n265), .A3(n525), .A2(n263), .A4(n321), .S0(n302), 
        .S1(n298), .Y(n524) );
  MUX41X1_HVT U61 ( .A1(n261), .A3(n320), .A2(n319), .A4(n277), .S0(n302), 
        .S1(n298), .Y(n522) );
  NAND2X0_HVT U62 ( .A1(n296), .A2(n581), .Y(n521) );
  MUX41X1_HVT U63 ( .A1(n521), .A3(n312), .A2(n342), .A4(n318), .S0(n302), 
        .S1(n298), .Y(n520) );
  AO21X1_HVT U66 ( .A1(n316), .A2(in[5]), .A3(n341), .Y(n517) );
  MUX41X1_HVT U68 ( .A1(n314), .A3(n517), .A2(n516), .A4(n518), .S0(n266), 
        .S1(n301), .Y(n515) );
  MUX41X1_HVT U69 ( .A1(n515), .A3(n523), .A2(n519), .A4(n529), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n286), .A2(n510), .Y(n511) );
  MUX41X1_HVT U74 ( .A1(n512), .A3(n557), .A2(n511), .A4(n559), .S0(n268), 
        .S1(n274), .Y(n509) );
  MUX41X1_HVT U75 ( .A1(n345), .A3(n350), .A2(n363), .A4(n325), .S0(n266), 
        .S1(n301), .Y(n508) );
  MUX41X1_HVT U77 ( .A1(n574), .A3(n352), .A2(n507), .A4(n351), .S0(n273), 
        .S1(n271), .Y(n506) );
  MUX41X1_HVT U78 ( .A1(n506), .A3(n509), .A2(n508), .A4(n513), .S0(in[0]), 
        .S1(n299), .Y(n505) );
  AND3X1_HVT U80 ( .A1(n288), .A2(n527), .A3(n502), .Y(n503) );
  MUX41X1_HVT U82 ( .A1(n538), .A3(n323), .A2(n306), .A4(n568), .S0(n266), 
        .S1(n273), .Y(n500) );
  AND2X1_HVT U83 ( .A1(n219), .A2(n248), .Y(n499) );
  MUX41X1_HVT U84 ( .A1(n324), .A3(n576), .A2(n566), .A4(n499), .S0(n266), 
        .S1(n301), .Y(n498) );
  NAND2X0_HVT U85 ( .A1(n296), .A2(n362), .Y(n497) );
  MUX41X1_HVT U86 ( .A1(n350), .A3(n497), .A2(n262), .A4(n258), .S0(n266), 
        .S1(n300), .Y(n496) );
  MUX41X1_HVT U87 ( .A1(n496), .A3(n500), .A2(n498), .A4(n501), .S0(in[0]), 
        .S1(n272), .Y(n495) );
  MUX41X1_HVT U90 ( .A1(n537), .A3(n541), .A2(n347), .A4(n494), .S0(n267), 
        .S1(n275), .Y(n493) );
  AO21X1_HVT U93 ( .A1(n275), .A2(n489), .A3(n346), .Y(n490) );
  MUX41X1_HVT U96 ( .A1(n306), .A3(n260), .A2(n349), .A4(n487), .S0(n266), 
        .S1(n301), .Y(n486) );
  MUX41X1_HVT U97 ( .A1(n345), .A3(n260), .A2(n218), .A4(n567), .S0(n266), 
        .S1(n275), .Y(n485) );
  NAND2X0_HVT U101 ( .A1(n480), .A2(n479), .Y(n481) );
  MUX41X1_HVT U103 ( .A1(n240), .A3(n315), .A2(n328), .A4(n548), .S0(n266), 
        .S1(n300), .Y(n477) );
  OA21X1_HVT U109 ( .A1(n335), .A2(n297), .A3(n321), .Y(n472) );
  NAND2X0_HVT U110 ( .A1(n288), .A2(n470), .Y(n471) );
  MUX41X1_HVT U114 ( .A1(n467), .A3(n473), .A2(n469), .A4(n472), .S0(n299), 
        .S1(n274), .Y(n466) );
  AND2X1_HVT U115 ( .A1(n219), .A2(n277), .Y(n465) );
  MUX41X1_HVT U116 ( .A1(n570), .A3(n465), .A2(n325), .A4(n552), .S0(n267), 
        .S1(n302), .Y(n464) );
  NAND2X0_HVT U123 ( .A1(n456), .A2(n455), .Y(n457) );
  MUX41X1_HVT U125 ( .A1(n561), .A3(n265), .A2(n314), .A4(n354), .S0(n267), 
        .S1(n302), .Y(n453) );
  AND3X1_HVT U128 ( .A1(n270), .A2(n296), .A3(n248), .Y(n450) );
  MUX41X1_HVT U131 ( .A1(n448), .A3(n450), .A2(n449), .A4(n451), .S0(in[5]), 
        .S1(n302), .Y(n447) );
  MUX41X1_HVT U132 ( .A1(n447), .A3(n460), .A2(n452), .A4(n466), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  AND2X1_HVT U140 ( .A1(n285), .A2(n296), .Y(n439) );
  MUX41X1_HVT U141 ( .A1(n558), .A3(n336), .A2(n439), .A4(n332), .S0(n268), 
        .S1(n302), .Y(n438) );
  MUX41X1_HVT U142 ( .A1(n324), .A3(n277), .A2(n343), .A4(n285), .S0(n267), 
        .S1(n302), .Y(n437) );
  NAND2X0_HVT U146 ( .A1(n294), .A2(n289), .Y(n510) );
  OA21X1_HVT U151 ( .A1(n543), .A2(n303), .A3(n429), .Y(n430) );
  MUX41X1_HVT U153 ( .A1(n471), .A3(n261), .A2(n581), .A4(n308), .S0(n267), 
        .S1(n274), .Y(n427) );
  AND2X1_HVT U154 ( .A1(n275), .A2(n284), .Y(n426) );
  NAND2X0_HVT U158 ( .A1(n291), .A2(n362), .Y(n422) );
  MUX41X1_HVT U159 ( .A1(n570), .A3(n277), .A2(n422), .A4(n251), .S0(n266), 
        .S1(n301), .Y(n421) );
  MUX41X1_HVT U160 ( .A1(n421), .A3(n427), .A2(n423), .A4(n428), .S0(in[0]), 
        .S1(n272), .Y(n420) );
  NAND2X0_HVT U166 ( .A1(n289), .A2(n527), .Y(n415) );
  NAND2X0_HVT U167 ( .A1(n363), .A2(n296), .Y(n414) );
  OA21X1_HVT U170 ( .A1(n263), .A2(n303), .A3(n552), .Y(n411) );
  NAND2X0_HVT U174 ( .A1(n292), .A2(n576), .Y(n569) );
  NAND2X0_HVT U177 ( .A1(n292), .A2(n281), .Y(n406) );
  MUX41X1_HVT U178 ( .A1(n565), .A3(n406), .A2(n357), .A4(n545), .S0(n268), 
        .S1(n300), .Y(n405) );
  MUX41X1_HVT U179 ( .A1(n555), .A3(n358), .A2(n310), .A4(n357), .S0(n271), 
        .S1(n273), .Y(n404) );
  MUX41X1_HVT U180 ( .A1(n313), .A3(n574), .A2(n570), .A4(n257), .S0(n273), 
        .S1(n269), .Y(n403) );
  MUX41X1_HVT U181 ( .A1(n403), .A3(n405), .A2(n404), .A4(n407), .S0(in[0]), 
        .S1(n272), .Y(n402) );
  OA21X1_HVT U184 ( .A1(n549), .A2(n303), .A3(n324), .Y(n399) );
  MUX41X1_HVT U186 ( .A1(n260), .A3(n544), .A2(n510), .A4(n537), .S0(n270), 
        .S1(n300), .Y(n397) );
  MUX41X1_HVT U189 ( .A1(n395), .A3(n569), .A2(n396), .A4(n344), .S0(n273), 
        .S1(n270), .Y(n394) );
  MUX41X1_HVT U190 ( .A1(n394), .A3(n397), .A2(n398), .A4(n401), .S0(n272), 
        .S1(in[0]), .Y(n393) );
  MUX41X1_HVT U193 ( .A1(n541), .A3(n548), .A2(n535), .A4(n392), .S0(n271), 
        .S1(n301), .Y(n391) );
  MUX41X1_HVT U195 ( .A1(n576), .A3(n349), .A2(n582), .A4(n546), .S0(n268), 
        .S1(n301), .Y(n389) );
  AO21X1_HVT U197 ( .A1(n262), .A2(n274), .A3(n346), .Y(n387) );
  MUX41X1_HVT U199 ( .A1(n386), .A3(n390), .A2(n389), .A4(n391), .S0(in[0]), 
        .S1(n272), .Y(n385) );
  MUX41X1_HVT U203 ( .A1(n547), .A3(n338), .A2(n571), .A4(n551), .S0(n269), 
        .S1(n300), .Y(n381) );
  MUX41X1_HVT U204 ( .A1(n528), .A3(n570), .A2(n333), .A4(n560), .S0(n270), 
        .S1(n273), .Y(n380) );
  MUX41X1_HVT U205 ( .A1(n248), .A3(n239), .A2(n358), .A4(n331), .S0(n266), 
        .S1(n300), .Y(n379) );
  NAND2X0_HVT U208 ( .A1(n218), .A2(n287), .Y(n470) );
  NAND2X0_HVT U212 ( .A1(n293), .A2(n286), .Y(n527) );
  NAND2X0_HVT U214 ( .A1(n576), .A2(n296), .Y(n377) );
  NAND2X0_HVT U215 ( .A1(n470), .A2(n286), .Y(n376) );
  AO21X1_HVT U216 ( .A1(n296), .A2(n360), .A3(n303), .Y(n480) );
  NAND2X0_HVT U218 ( .A1(n360), .A2(n211), .Y(n429) );
  NAND2X0_HVT U220 ( .A1(n274), .A2(n377), .Y(n502) );
  XOR2X2_HVT U1 ( .A1(n303), .A2(n556), .Y(n539) );
  INVX2_HVT U2 ( .A(n50), .Y(n576) );
  MUX41X1_HVT U6 ( .A1(n537), .A3(n345), .A2(n510), .A4(n356), .S0(n23), .S1(
        n304), .Y(n433) );
  IBUFFX16_HVT U7 ( .A(n268), .Y(n23) );
  INVX1_HVT U8 ( .A(n274), .Y(n237) );
  MUX21X1_HVT U9 ( .A1(n545), .A2(n352), .S0(n273), .Y(n424) );
  INVX1_HVT U10 ( .A(n273), .Y(n231) );
  INVX1_HVT U11 ( .A(n275), .Y(n216) );
  MUX21X1_HVT U12 ( .A1(n383), .A2(n384), .S0(n269), .Y(n382) );
  MUX21X1_HVT U14 ( .A1(n337), .A2(n560), .S0(n237), .Y(n442) );
  MUX21X1_HVT U16 ( .A1(n530), .A2(n534), .S0(n270), .Y(n529) );
  MUX21X1_HVT U17 ( .A1(n424), .A2(n425), .S0(n271), .Y(n423) );
  MUX21X1_HVT U18 ( .A1(n257), .A2(n566), .S0(n231), .Y(n384) );
  MUX21X1_HVT U19 ( .A1(n311), .A2(n554), .S0(n216), .Y(n436) );
  MUX21X2_HVT U20 ( .A1(n461), .A2(n464), .S0(n48), .Y(n460) );
  IBUFFX16_HVT U22 ( .A(n247), .Y(n48) );
  INVX4_HVT U23 ( .A(n304), .Y(n302) );
  XNOR2X2_HVT U25 ( .A1(n280), .A2(n283), .Y(n50) );
  MUX21X2_HVT U26 ( .A1(n278), .A2(n276), .S0(n293), .Y(n566) );
  NBUFFX2_HVT U27 ( .A(n50), .Y(n278) );
  INVX0_HVT U28 ( .A(n566), .Y(n319) );
  MUX21X2_HVT U29 ( .A1(n579), .A2(n442), .S0(n168), .Y(n441) );
  IBUFFX16_HVT U30 ( .A(n271), .Y(n168) );
  MUX21X2_HVT U31 ( .A1(n520), .A2(n522), .S0(n269), .Y(n519) );
  AO21X2_HVT U32 ( .A1(n271), .A2(n285), .A3(n576), .Y(n462) );
  MUX21X2_HVT U34 ( .A1(n279), .A2(n284), .S0(n293), .Y(n560) );
  INVX0_HVT U36 ( .A(n560), .Y(n324) );
  OA21X1_HVT U37 ( .A1(n575), .A2(n303), .A3(n336), .Y(n383) );
  INVX2_HVT U38 ( .A(n235), .Y(n210) );
  INVX2_HVT U39 ( .A(n235), .Y(n211) );
  MUX41X1_HVT U40 ( .A1(n493), .A3(n486), .A2(n488), .A4(n485), .S0(n212), 
        .S1(n213), .Y(n484) );
  IBUFFX16_HVT U41 ( .A(in[0]), .Y(n212) );
  IBUFFX16_HVT U43 ( .A(n298), .Y(n213) );
  IBUFFX2_HVT U44 ( .A(n554), .Y(n328) );
  MUX21X2_HVT U45 ( .A1(n435), .A2(n436), .S0(n217), .Y(n434) );
  IBUFFX16_HVT U46 ( .A(n270), .Y(n217) );
  NBUFFX2_HVT U47 ( .A(in[1]), .Y(n236) );
  INVX1_HVT U48 ( .A(n295), .Y(n218) );
  INVX1_HVT U49 ( .A(n295), .Y(n219) );
  IBUFFX2_HVT U50 ( .A(in[1]), .Y(n295) );
  INVX1_HVT U52 ( .A(n295), .Y(n293) );
  INVX2_HVT U54 ( .A(in[1]), .Y(n235) );
  INVX1_HVT U55 ( .A(in[7]), .Y(n304) );
  MUX41X1_HVT U60 ( .A1(n437), .A3(n433), .A2(n438), .A4(n434), .S0(n232), 
        .S1(n298), .Y(n432) );
  IBUFFX16_HVT U64 ( .A(in[0]), .Y(n232) );
  IBUFFX2_HVT U65 ( .A(n304), .Y(n300) );
  OA21X1_HVT U67 ( .A1(n309), .A2(n303), .A3(n552), .Y(n435) );
  INVX2_HVT U70 ( .A(n235), .Y(n291) );
  IBUFFX16_HVT U71 ( .A(n295), .Y(n294) );
  MUX41X1_HVT U72 ( .A1(n441), .A3(n444), .A2(n443), .A4(n445), .S0(n233), 
        .S1(n234), .Y(n440) );
  IBUFFX16_HVT U76 ( .A(n249), .Y(n233) );
  IBUFFX16_HVT U79 ( .A(n247), .Y(n234) );
  INVX4_HVT U81 ( .A(n236), .Y(n296) );
  INVX2_HVT U88 ( .A(n235), .Y(n292) );
  IBUFFX2_HVT U89 ( .A(in[7]), .Y(n303) );
  MUX21X2_HVT U91 ( .A1(n378), .A2(n385), .S0(in[6]), .Y(out[7]) );
  MUX21X2_HVT U92 ( .A1(n402), .A2(n393), .S0(n253), .Y(out[6]) );
  INVX1_HVT U94 ( .A(in[6]), .Y(n253) );
  INVX1_HVT U95 ( .A(n580), .Y(n238) );
  INVX0_HVT U98 ( .A(n238), .Y(n239) );
  INVX0_HVT U99 ( .A(n238), .Y(n240) );
  INVX0_HVT U100 ( .A(n238), .Y(n241) );
  MUX21X1_HVT U102 ( .A1(n539), .A2(n514), .S0(n269), .Y(n513) );
  INVX1_HVT U104 ( .A(in[2]), .Y(n297) );
  MUX41X1_HVT U105 ( .A1(n569), .A3(n353), .A2(n408), .A4(n280), .S0(n303), 
        .S1(n242), .Y(n407) );
  IBUFFX2_HVT U106 ( .A(n267), .Y(n242) );
  MUX21X2_HVT U107 ( .A1(n495), .A2(n505), .S0(in[6]), .Y(out[1]) );
  IBUFFX2_HVT U108 ( .A(n545), .Y(n336) );
  MUX41X1_HVT U111 ( .A1(n326), .A3(n339), .A2(n578), .A4(n337), .S0(n303), 
        .S1(n297), .Y(n401) );
  NBUFFX2_HVT U112 ( .A(in[2]), .Y(n267) );
  INVX1_HVT U113 ( .A(n259), .Y(n244) );
  INVX1_HVT U117 ( .A(n304), .Y(n301) );
  INVX1_HVT U118 ( .A(n419), .Y(n245) );
  INVX0_HVT U119 ( .A(n250), .Y(n444) );
  INVX0_HVT U120 ( .A(n556), .Y(n252) );
  INVX1_HVT U121 ( .A(n254), .Y(n255) );
  INVX1_HVT U122 ( .A(n298), .Y(n247) );
  INVX1_HVT U124 ( .A(in[0]), .Y(n249) );
  INVX0_HVT U126 ( .A(n577), .Y(n251) );
  MUX41X1_HVT U127 ( .A1(n547), .A3(n356), .A2(n550), .A4(n258), .S0(n242), 
        .S1(n303), .Y(n443) );
  MUX41X1_HVT U129 ( .A1(n285), .A3(n348), .A2(n415), .A4(n414), .S0(n297), 
        .S1(n301), .Y(n413) );
  INVX1_HVT U130 ( .A(n243), .Y(n418) );
  MUX41X1_HVT U133 ( .A1(n246), .A3(n565), .A2(n245), .A4(n244), .S0(n297), 
        .S1(n300), .Y(n243) );
  NAND2X0_HVT U134 ( .A1(n576), .A2(n510), .Y(n246) );
  MUX41X1_HVT U135 ( .A1(n418), .A3(n413), .A2(n416), .A4(n410), .S0(n249), 
        .S1(n247), .Y(n409) );
  MUX21X2_HVT U136 ( .A1(n420), .A2(n409), .S0(n253), .Y(out[5]) );
  IBUFFX2_HVT U137 ( .A(n280), .Y(n248) );
  MUX41X1_HVT U138 ( .A1(n382), .A3(n380), .A2(n381), .A4(n379), .S0(n249), 
        .S1(n247), .Y(n378) );
  NBUFFX4_HVT U139 ( .A(n364), .Y(n280) );
  MUX41X1_HVT U143 ( .A1(n252), .A3(n251), .A2(n285), .A4(n368), .S0(n242), 
        .S1(n303), .Y(n250) );
  MUX21X2_HVT U144 ( .A1(n440), .A2(n432), .S0(n253), .Y(out[4]) );
  MUX41X1_HVT U145 ( .A1(n327), .A3(n536), .A2(n476), .A4(n344), .S0(n266), 
        .S1(n300), .Y(n475) );
  XOR2X1_HVT U147 ( .A1(n297), .A2(n304), .Y(n254) );
  MUX41X1_HVT U148 ( .A1(n482), .A3(n478), .A2(n477), .A4(n475), .S0(n247), 
        .S1(n249), .Y(n474) );
  MUX21X2_HVT U149 ( .A1(n484), .A2(n474), .S0(n253), .Y(out[2]) );
  MUX41X1_HVT U150 ( .A1(n285), .A3(n355), .A2(n556), .A4(n542), .S0(n303), 
        .S1(n297), .Y(n390) );
  MUX41X1_HVT U152 ( .A1(n417), .A3(n537), .A2(n329), .A4(n561), .S0(n303), 
        .S1(n297), .Y(n416) );
  MUX21X1_HVT U155 ( .A1(n288), .A2(n468), .S0(n256), .Y(n467) );
  MUX21X2_HVT U156 ( .A1(n483), .A2(n261), .S0(n255), .Y(n482) );
  XNOR2X1_HVT U157 ( .A1(n296), .A2(n297), .Y(n256) );
  IBUFFX2_HVT U161 ( .A(n235), .Y(n290) );
  INVX0_HVT U162 ( .A(n283), .Y(n361) );
  INVX1_HVT U163 ( .A(n578), .Y(n359) );
  MUX21X1_HVT U164 ( .A1(n259), .A2(n319), .S0(n267), .Y(n449) );
  NBUFFX2_HVT U165 ( .A(n50), .Y(n279) );
  NBUFFX2_HVT U168 ( .A(n50), .Y(n277) );
  AND2X1_HVT U169 ( .A1(n279), .A2(n527), .Y(n257) );
  INVX1_HVT U171 ( .A(n581), .Y(n363) );
  MUX21X1_HVT U172 ( .A1(n359), .A2(n362), .S0(n299), .Y(n531) );
  NBUFFX2_HVT U173 ( .A(n578), .Y(n287) );
  MUX21X1_HVT U175 ( .A1(n552), .A2(n471), .S0(n267), .Y(n469) );
  MUX21X1_HVT U176 ( .A1(n315), .A2(n360), .S0(in[5]), .Y(n516) );
  AND2X1_HVT U182 ( .A1(n288), .A2(n510), .Y(n258) );
  MUX21X1_HVT U183 ( .A1(n279), .A2(n362), .S0(n293), .Y(n575) );
  MUX21X1_HVT U185 ( .A1(n453), .A2(n454), .S0(in[5]), .Y(n452) );
  MUX21X1_HVT U187 ( .A1(n458), .A2(n457), .S0(n275), .Y(n454) );
  MUX21X1_HVT U188 ( .A1(n288), .A2(n278), .S0(n290), .Y(n542) );
  MUX21X1_HVT U191 ( .A1(n277), .A2(n282), .S0(n292), .Y(n479) );
  MUX21X1_HVT U192 ( .A1(n278), .A2(n359), .S0(n290), .Y(n487) );
  MUX21X1_HVT U194 ( .A1(n287), .A2(n576), .S0(n219), .Y(n546) );
  MUX21X1_HVT U196 ( .A1(n359), .A2(n363), .S0(n218), .Y(n408) );
  MUX21X1_HVT U198 ( .A1(n362), .A2(n278), .S0(n218), .Y(n419) );
  MUX21X1_HVT U200 ( .A1(n576), .A2(n360), .S0(n211), .Y(n368) );
  MUX21X1_HVT U201 ( .A1(n576), .A2(n363), .S0(n218), .Y(n558) );
  MUX21X1_HVT U202 ( .A1(n287), .A2(n286), .S0(n210), .Y(n494) );
  MUX21X1_HVT U206 ( .A1(n576), .A2(n282), .S0(n218), .Y(n507) );
  XOR2X1_HVT U207 ( .A1(n576), .A2(n210), .Y(n537) );
  MUX21X1_HVT U209 ( .A1(n276), .A2(n576), .S0(n210), .Y(n371) );
  MUX21X1_HVT U210 ( .A1(n363), .A2(n362), .S0(n293), .Y(n556) );
  MUX21X1_HVT U211 ( .A1(n362), .A2(n359), .S0(n292), .Y(n545) );
  MUX21X1_HVT U213 ( .A1(n362), .A2(n276), .S0(n211), .Y(n549) );
  MUX21X1_HVT U217 ( .A1(n276), .A2(n363), .S0(n290), .Y(n543) );
  MUX21X1_HVT U219 ( .A1(n282), .A2(n359), .S0(n291), .Y(n554) );
  MUX21X1_HVT U221 ( .A1(n462), .A2(n463), .S0(n274), .Y(n461) );
  MUX21X1_HVT U222 ( .A1(n308), .A2(n333), .S0(n267), .Y(n463) );
  MUX21X1_HVT U223 ( .A1(n330), .A2(n446), .S0(n270), .Y(n445) );
  MUX21X1_HVT U224 ( .A1(n354), .A2(n573), .S0(n274), .Y(n446) );
  NAND2X0_HVT U225 ( .A1(n280), .A2(n361), .Y(n578) );
  MUX21X1_HVT U226 ( .A1(n359), .A2(n281), .S0(n291), .Y(n369) );
  INVX1_HVT U227 ( .A(n582), .Y(n362) );
  MUX21X1_HVT U228 ( .A1(n288), .A2(n286), .S0(n293), .Y(n568) );
  MUX21X1_HVT U229 ( .A1(n360), .A2(n359), .S0(n290), .Y(n564) );
  MUX21X1_HVT U230 ( .A1(n331), .A2(n568), .S0(n271), .Y(n483) );
  MUX21X1_HVT U231 ( .A1(n307), .A2(n459), .S0(n268), .Y(n458) );
  MUX21X1_HVT U232 ( .A1(n281), .A2(n276), .S0(n293), .Y(n459) );
  NBUFFX2_HVT U233 ( .A(n581), .Y(n288) );
  INVX1_HVT U234 ( .A(n285), .Y(n360) );
  MUX21X1_HVT U235 ( .A1(n287), .A2(n289), .S0(n292), .Y(n489) );
  MUX21X1_HVT U236 ( .A1(n276), .A2(n362), .S0(n292), .Y(n572) );
  MUX21X1_HVT U237 ( .A1(n276), .A2(n282), .S0(n210), .Y(n392) );
  XOR2X1_HVT U238 ( .A1(n581), .A2(n211), .Y(n535) );
  MUX21X1_HVT U239 ( .A1(n276), .A2(n289), .S0(n290), .Y(n395) );
  MUX21X1_HVT U240 ( .A1(n582), .A2(n288), .S0(n218), .Y(n396) );
  XOR2X1_HVT U241 ( .A1(n219), .A2(n360), .Y(n538) );
  MUX21X1_HVT U242 ( .A1(n581), .A2(n281), .S0(n210), .Y(n375) );
  XNOR2X1_HVT U243 ( .A1(n578), .A2(n219), .Y(n259) );
  AND2X1_HVT U244 ( .A1(n290), .A2(n363), .Y(n260) );
  MUX21X1_HVT U245 ( .A1(n289), .A2(n286), .S0(n290), .Y(n552) );
  MUX21X1_HVT U246 ( .A1(n287), .A2(n276), .S0(n210), .Y(n571) );
  MUX21X1_HVT U247 ( .A1(n581), .A2(n287), .S0(n219), .Y(n367) );
  AND2X1_HVT U248 ( .A1(n289), .A2(n470), .Y(n261) );
  XNOR2X1_HVT U249 ( .A1(n582), .A2(n219), .Y(n262) );
  MUX21X1_HVT U250 ( .A1(n286), .A2(n276), .S0(n293), .Y(n373) );
  MUX21X1_HVT U251 ( .A1(n286), .A2(n281), .S0(n291), .Y(n512) );
  MUX21X1_HVT U252 ( .A1(n573), .A2(n289), .S0(n270), .Y(n456) );
  XOR2X1_HVT U253 ( .A1(n280), .A2(n211), .Y(n557) );
  NBUFFX2_HVT U254 ( .A(in[7]), .Y(n275) );
  NBUFFX2_HVT U255 ( .A(in[7]), .Y(n273) );
  NBUFFX2_HVT U256 ( .A(in[7]), .Y(n274) );
  NBUFFX2_HVT U257 ( .A(n361), .Y(n276) );
  NBUFFX2_HVT U258 ( .A(in[2]), .Y(n268) );
  NBUFFX2_HVT U259 ( .A(n299), .Y(n272) );
  NBUFFX2_HVT U260 ( .A(in[2]), .Y(n270) );
  NBUFFX2_HVT U261 ( .A(in[2]), .Y(n271) );
  NBUFFX2_HVT U262 ( .A(in[2]), .Y(n269) );
  NBUFFX2_HVT U263 ( .A(in[2]), .Y(n266) );
  MUX21X1_HVT U264 ( .A1(n481), .A2(n330), .S0(n270), .Y(n478) );
  MUX21X1_HVT U265 ( .A1(n399), .A2(n400), .S0(n269), .Y(n398) );
  MUX21X1_HVT U266 ( .A1(n497), .A2(n284), .S0(n274), .Y(n400) );
  XOR2X1_HVT U267 ( .A1(n291), .A2(n283), .Y(n536) );
  MUX21X1_HVT U268 ( .A1(n286), .A2(n279), .S0(n291), .Y(n476) );
  MUX21X1_HVT U269 ( .A1(n430), .A2(n431), .S0(n271), .Y(n428) );
  MUX21X1_HVT U270 ( .A1(n351), .A2(n360), .S0(n274), .Y(n431) );
  MUX21X1_HVT U271 ( .A1(n504), .A2(n503), .S0(n271), .Y(n501) );
  MUX21X1_HVT U272 ( .A1(n562), .A2(n286), .S0(n275), .Y(n504) );
  MUX21X1_HVT U273 ( .A1(n412), .A2(n411), .S0(n270), .Y(n410) );
  MUX21X1_HVT U274 ( .A1(n286), .A2(n349), .S0(n275), .Y(n412) );
  AND2X1_HVT U275 ( .A1(n279), .A2(n296), .Y(n263) );
  MUX21X1_HVT U276 ( .A1(n284), .A2(n359), .S0(n218), .Y(n544) );
  MUX21X1_HVT U277 ( .A1(n362), .A2(n349), .S0(n275), .Y(n514) );
  MUX21X1_HVT U278 ( .A1(n360), .A2(n363), .S0(n294), .Y(n417) );
  NAND2X0_HVT U279 ( .A1(n283), .A2(n282), .Y(n581) );
  NBUFFX2_HVT U280 ( .A(n364), .Y(n282) );
  MUX21X1_HVT U281 ( .A1(n363), .A2(n284), .S0(n291), .Y(n563) );
  MUX21X1_HVT U282 ( .A1(n334), .A2(n241), .S0(n268), .Y(n473) );
  MUX21X1_HVT U283 ( .A1(n426), .A2(n288), .S0(n264), .Y(n425) );
  MUX21X1_HVT U284 ( .A1(n565), .A2(n332), .S0(n268), .Y(n448) );
  MUX21X1_HVT U285 ( .A1(n532), .A2(n533), .S0(n273), .Y(n530) );
  MUX21X1_HVT U286 ( .A1(n284), .A2(n548), .S0(n299), .Y(n533) );
  XOR2X1_HVT U287 ( .A1(n292), .A2(n272), .Y(n540) );
  MUX21X1_HVT U288 ( .A1(n240), .A2(n296), .S0(n269), .Y(n455) );
  NBUFFX2_HVT U289 ( .A(n573), .Y(n285) );
  MUX21X1_HVT U290 ( .A1(n284), .A2(n360), .S0(n210), .Y(n372) );
  MUX21X1_HVT U291 ( .A1(n553), .A2(n376), .S0(n273), .Y(n370) );
  MUX21X1_HVT U292 ( .A1(n287), .A2(n284), .S0(n219), .Y(n574) );
  MUX21X1_HVT U293 ( .A1(n317), .A2(n296), .S0(in[5]), .Y(n518) );
  NBUFFX2_HVT U294 ( .A(n573), .Y(n286) );
  MUX21X1_HVT U295 ( .A1(n327), .A2(n553), .S0(n268), .Y(n451) );
  MUX21X1_HVT U296 ( .A1(n340), .A2(n357), .S0(n274), .Y(n388) );
  MUX21X1_HVT U297 ( .A1(n288), .A2(n492), .S0(n264), .Y(n491) );
  MUX21X1_HVT U298 ( .A1(n284), .A2(n281), .S0(n275), .Y(n492) );
  NBUFFX2_HVT U299 ( .A(n582), .Y(n289) );
  NBUFFX2_HVT U300 ( .A(n364), .Y(n281) );
  XNOR2X1_HVT U301 ( .A1(n304), .A2(n211), .Y(n264) );
  AND2X1_HVT U302 ( .A1(n276), .A2(n296), .Y(n265) );
  NBUFFX2_HVT U303 ( .A(in[5]), .Y(n299) );
  NBUFFX2_HVT U304 ( .A(in[5]), .Y(n298) );
  MUX21X1_HVT U305 ( .A1(n388), .A2(n387), .S0(n269), .Y(n386) );
  INVX0_HVT U306 ( .A(in[4]), .Y(n364) );
  MUX21X1_HVT U307 ( .A1(n490), .A2(n491), .S0(n271), .Y(n488) );
  MUX21X1_HVT U308 ( .A1(n524), .A2(n526), .S0(n269), .Y(n523) );
  MUX21X1_HVT U309 ( .A1(n359), .A2(n248), .S0(n211), .Y(n551) );
  NAND2X0_HVT U310 ( .A1(n283), .A2(in[4]), .Y(n582) );
  MUX21X1_HVT U311 ( .A1(n248), .A2(n576), .S0(n211), .Y(n374) );
  MUX21X1_HVT U312 ( .A1(n248), .A2(n362), .S0(n291), .Y(n547) );
  MUX21X1_HVT U313 ( .A1(n248), .A2(n360), .S0(n291), .Y(n565) );
  NAND2X0_HVT U314 ( .A1(in[4]), .A2(n361), .Y(n573) );
  MUX21X1_HVT U315 ( .A1(n248), .A2(n288), .S0(n292), .Y(n562) );
  MUX21X1_HVT U316 ( .A1(n289), .A2(n248), .S0(n292), .Y(n555) );
  MUX21X1_HVT U317 ( .A1(n284), .A2(n248), .S0(n267), .Y(n468) );
  MUX21X1_HVT U318 ( .A1(n248), .A2(n286), .S0(n290), .Y(n366) );
  MUX21X1_HVT U319 ( .A1(n248), .A2(n289), .S0(n219), .Y(n365) );
  MUX21X1_HVT U320 ( .A1(n276), .A2(n248), .S0(n210), .Y(n553) );
  NBUFFX2_HVT U321 ( .A(in[3]), .Y(n283) );
  NBUFFX2_HVT U322 ( .A(in[3]), .Y(n284) );
  INVX0_HVT U323 ( .A(n561), .Y(n305) );
  INVX0_HVT U324 ( .A(n559), .Y(n306) );
  INVX0_HVT U325 ( .A(n550), .Y(n307) );
  INVX0_HVT U326 ( .A(n548), .Y(n308) );
  INVX0_HVT U327 ( .A(n414), .Y(n309) );
  INVX0_HVT U328 ( .A(n377), .Y(n310) );
  INVX0_HVT U329 ( .A(n241), .Y(n311) );
  INVX0_HVT U330 ( .A(n567), .Y(n312) );
  INVX0_HVT U331 ( .A(n579), .Y(n313) );
  INVX0_HVT U332 ( .A(n575), .Y(n314) );
  INVX0_HVT U333 ( .A(n574), .Y(n315) );
  INVX0_HVT U334 ( .A(n572), .Y(n316) );
  INVX0_HVT U335 ( .A(n571), .Y(n317) );
  INVX0_HVT U336 ( .A(n568), .Y(n318) );
  INVX0_HVT U337 ( .A(n565), .Y(n320) );
  INVX0_HVT U338 ( .A(n564), .Y(n321) );
  INVX0_HVT U339 ( .A(n563), .Y(n322) );
  INVX0_HVT U340 ( .A(n562), .Y(n323) );
  INVX0_HVT U341 ( .A(n558), .Y(n325) );
  INVX0_HVT U342 ( .A(n557), .Y(n326) );
  INVX0_HVT U343 ( .A(n555), .Y(n327) );
  INVX0_HVT U344 ( .A(n553), .Y(n329) );
  INVX0_HVT U345 ( .A(n370), .Y(n330) );
  INVX0_HVT U346 ( .A(n552), .Y(n331) );
  INVX0_HVT U347 ( .A(n551), .Y(n332) );
  INVX0_HVT U348 ( .A(n549), .Y(n333) );
  INVX0_HVT U349 ( .A(n547), .Y(n334) );
  INVX0_HVT U350 ( .A(n546), .Y(n335) );
  INVX0_HVT U351 ( .A(n544), .Y(n337) );
  INVX0_HVT U352 ( .A(n543), .Y(n338) );
  INVX0_HVT U353 ( .A(n542), .Y(n339) );
  INVX0_HVT U354 ( .A(n541), .Y(n340) );
  INVX0_HVT U355 ( .A(n510), .Y(n341) );
  INVX0_HVT U356 ( .A(n570), .Y(n342) );
  INVX0_HVT U357 ( .A(n470), .Y(n343) );
  INVX0_HVT U358 ( .A(n376), .Y(n344) );
  INVX0_HVT U359 ( .A(n527), .Y(n345) );
  INVX0_HVT U360 ( .A(n429), .Y(n346) );
  INVX0_HVT U361 ( .A(n375), .Y(n347) );
  INVX0_HVT U362 ( .A(n374), .Y(n348) );
  INVX0_HVT U363 ( .A(n373), .Y(n349) );
  INVX0_HVT U364 ( .A(n372), .Y(n350) );
  INVX0_HVT U365 ( .A(n371), .Y(n351) );
  INVX0_HVT U366 ( .A(n489), .Y(n352) );
  INVX0_HVT U367 ( .A(n479), .Y(n353) );
  INVX0_HVT U368 ( .A(n369), .Y(n354) );
  INVX0_HVT U369 ( .A(n368), .Y(n355) );
  INVX0_HVT U370 ( .A(n367), .Y(n356) );
  INVX0_HVT U371 ( .A(n366), .Y(n357) );
  INVX0_HVT U372 ( .A(n365), .Y(n358) );
endmodule

