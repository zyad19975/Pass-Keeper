
module sbox_10 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n50, n210, n211, n212, n213, n216, n217, n218, n219, n229, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605;

  NAND2X0_HVT U3 ( .A1(n321), .A2(n314), .Y(n603) );
  NAND2X0_HVT U4 ( .A1(n312), .A2(n603), .Y(n602) );
  NAND2X0_HVT U5 ( .A1(n321), .A2(n301), .Y(n600) );
  NAND2X0_HVT U13 ( .A1(n592), .A2(n316), .Y(n593) );
  NAND2X0_HVT U15 ( .A1(n603), .A2(n303), .Y(n590) );
  NAND2X0_HVT U21 ( .A1(n312), .A2(n255), .Y(n584) );
  NAND2X0_HVT U24 ( .A1(n309), .A2(n255), .Y(n582) );
  NAND2X0_HVT U33 ( .A1(n381), .A2(n255), .Y(n573) );
  NAND2X0_HVT U35 ( .A1(n307), .A2(n255), .Y(n571) );
  NAND2X0_HVT U42 ( .A1(n321), .A2(n309), .Y(n564) );
  MUX41X1_HVT U51 ( .A1(n370), .A3(n331), .A2(n346), .A4(n347), .S0(n327), 
        .S1(n297), .Y(n556) );
  NAND2X0_HVT U53 ( .A1(n553), .A2(n563), .Y(n554) );
  NAND2X0_HVT U56 ( .A1(n312), .A2(n549), .Y(n550) );
  MUX41X1_HVT U57 ( .A1(n371), .A3(n586), .A2(n550), .A4(n595), .S0(n327), 
        .S1(n297), .Y(n548) );
  NAND2X0_HVT U58 ( .A1(n316), .A2(n603), .Y(n547) );
  MUX41X1_HVT U61 ( .A1(n286), .A3(n344), .A2(n343), .A4(n302), .S0(n327), 
        .S1(n297), .Y(n544) );
  NAND2X0_HVT U62 ( .A1(n255), .A2(n604), .Y(n543) );
  AO21X1_HVT U66 ( .A1(n256), .A2(in[5]), .A3(n364), .Y(n539) );
  MUX41X1_HVT U68 ( .A1(n340), .A3(n539), .A2(n538), .A4(n540), .S0(n291), 
        .S1(n272), .Y(n537) );
  NAND2X0_HVT U73 ( .A1(n311), .A2(n532), .Y(n533) );
  MUX41X1_HVT U74 ( .A1(n534), .A3(n580), .A2(n533), .A4(n582), .S0(n293), 
        .S1(n326), .Y(n531) );
  MUX41X1_HVT U75 ( .A1(n368), .A3(n373), .A2(n385), .A4(n349), .S0(n291), 
        .S1(n272), .Y(n530) );
  MUX41X1_HVT U77 ( .A1(n597), .A3(n375), .A2(n529), .A4(n374), .S0(n299), 
        .S1(n324), .Y(n528) );
  MUX41X1_HVT U78 ( .A1(n528), .A3(n531), .A2(n530), .A4(n535), .S0(n308), 
        .S1(n297), .Y(n527) );
  AND3X1_HVT U80 ( .A1(n314), .A2(n549), .A3(n524), .Y(n525) );
  MUX41X1_HVT U82 ( .A1(n561), .A3(n347), .A2(n332), .A4(n591), .S0(n291), 
        .S1(n326), .Y(n522) );
  AND2X1_HVT U83 ( .A1(n321), .A2(n273), .Y(n521) );
  MUX41X1_HVT U84 ( .A1(n348), .A3(n599), .A2(n589), .A4(n521), .S0(n291), 
        .S1(n325), .Y(n520) );
  NAND2X0_HVT U85 ( .A1(n255), .A2(n384), .Y(n519) );
  MUX41X1_HVT U86 ( .A1(n373), .A3(n519), .A2(n287), .A4(n283), .S0(n291), 
        .S1(n326), .Y(n518) );
  MUX41X1_HVT U90 ( .A1(n560), .A3(n564), .A2(n370), .A4(n516), .S0(n292), 
        .S1(n325), .Y(n515) );
  AO21X1_HVT U93 ( .A1(n328), .A2(n511), .A3(n369), .Y(n512) );
  MUX41X1_HVT U96 ( .A1(n332), .A3(n285), .A2(n372), .A4(n509), .S0(n291), 
        .S1(n325), .Y(n508) );
  MUX41X1_HVT U97 ( .A1(n368), .A3(n285), .A2(n321), .A4(n590), .S0(n291), 
        .S1(n272), .Y(n507) );
  MUX41X1_HVT U98 ( .A1(n507), .A3(n510), .A2(n508), .A4(n515), .S0(n308), 
        .S1(n296), .Y(n506) );
  NAND2X0_HVT U101 ( .A1(n502), .A2(n501), .Y(n503) );
  MUX41X1_HVT U103 ( .A1(n603), .A3(n341), .A2(n352), .A4(n571), .S0(n291), 
        .S1(n326), .Y(n499) );
  MUX41X1_HVT U105 ( .A1(n351), .A3(n558), .A2(n498), .A4(n367), .S0(n291), 
        .S1(n325), .Y(n497) );
  MUX41X1_HVT U106 ( .A1(n497), .A3(n500), .A2(n499), .A4(n504), .S0(in[0]), 
        .S1(n296), .Y(n496) );
  OA21X1_HVT U109 ( .A1(n358), .A2(n268), .A3(n345), .Y(n494) );
  NAND2X0_HVT U110 ( .A1(n314), .A2(n492), .Y(n493) );
  MUX41X1_HVT U114 ( .A1(n489), .A3(n495), .A2(n491), .A4(n494), .S0(in[5]), 
        .S1(n325), .Y(n488) );
  AND2X1_HVT U115 ( .A1(n321), .A2(n302), .Y(n487) );
  NAND2X0_HVT U123 ( .A1(n478), .A2(n477), .Y(n479) );
  MUX41X1_HVT U125 ( .A1(n584), .A3(n290), .A2(n340), .A4(n377), .S0(n292), 
        .S1(n327), .Y(n475) );
  MUX41X1_HVT U131 ( .A1(n470), .A3(n472), .A2(n471), .A4(n473), .S0(in[5]), 
        .S1(n327), .Y(n469) );
  MUX41X1_HVT U132 ( .A1(n469), .A3(n482), .A2(n474), .A4(n488), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  MUX41X1_HVT U136 ( .A1(n283), .A3(n573), .A2(n379), .A4(n570), .S0(n292), 
        .S1(n327), .Y(n465) );
  MUX41X1_HVT U139 ( .A1(n463), .A3(n466), .A2(n465), .A4(n467), .S0(n308), 
        .S1(n296), .Y(n462) );
  AND2X1_HVT U140 ( .A1(n310), .A2(n265), .Y(n461) );
  OA21X1_HVT U144 ( .A1(n335), .A2(n329), .A3(n575), .Y(n457) );
  NAND2X0_HVT U146 ( .A1(n321), .A2(n316), .Y(n532) );
  MUX41X1_HVT U147 ( .A1(n379), .A3(n532), .A2(n368), .A4(n560), .S0(n293), 
        .S1(n327), .Y(n455) );
  MUX41X1_HVT U148 ( .A1(n455), .A3(n459), .A2(n456), .A4(n460), .S0(in[0]), 
        .S1(n296), .Y(n454) );
  OA21X1_HVT U151 ( .A1(n566), .A2(n329), .A3(n451), .Y(n452) );
  MUX41X1_HVT U153 ( .A1(n493), .A3(n286), .A2(n313), .A4(n334), .S0(n292), 
        .S1(n325), .Y(n449) );
  AND2X1_HVT U154 ( .A1(n328), .A2(n309), .Y(n448) );
  NAND2X0_HVT U158 ( .A1(n321), .A2(n384), .Y(n444) );
  MUX41X1_HVT U159 ( .A1(n593), .A3(n302), .A2(n444), .A4(n275), .S0(n324), 
        .S1(n326), .Y(n443) );
  MUX41X1_HVT U160 ( .A1(n443), .A3(n449), .A2(n445), .A4(n450), .S0(n308), 
        .S1(n298), .Y(n442) );
  AND2X1_HVT U162 ( .A1(n599), .A2(n532), .Y(n440) );
  MUX41X1_HVT U163 ( .A1(n344), .A3(n440), .A2(n284), .A4(n441), .S0(n324), 
        .S1(n272), .Y(n439) );
  MUX41X1_HVT U165 ( .A1(n584), .A3(n353), .A2(n560), .A4(n438), .S0(n327), 
        .S1(n323), .Y(n437) );
  NAND2X0_HVT U166 ( .A1(n316), .A2(n549), .Y(n436) );
  NAND2X0_HVT U167 ( .A1(n385), .A2(n255), .Y(n435) );
  MUX41X1_HVT U168 ( .A1(n371), .A3(n310), .A2(n435), .A4(n436), .S0(n323), 
        .S1(n272), .Y(n434) );
  OA21X1_HVT U170 ( .A1(n288), .A2(n329), .A3(n575), .Y(n432) );
  MUX41X1_HVT U172 ( .A1(n431), .A3(n437), .A2(n434), .A4(n439), .S0(n308), 
        .S1(n296), .Y(n430) );
  NAND2X0_HVT U174 ( .A1(n321), .A2(n599), .Y(n592) );
  MUX41X1_HVT U176 ( .A1(n305), .A3(n429), .A2(n376), .A4(n592), .S0(n327), 
        .S1(n324), .Y(n428) );
  NAND2X0_HVT U177 ( .A1(n321), .A2(n306), .Y(n427) );
  MUX41X1_HVT U178 ( .A1(n588), .A3(n427), .A2(n50), .A4(n568), .S0(n293), 
        .S1(n326), .Y(n426) );
  MUX41X1_HVT U179 ( .A1(n578), .A3(n380), .A2(n336), .A4(n50), .S0(n323), 
        .S1(n326), .Y(n425) );
  MUX41X1_HVT U180 ( .A1(n339), .A3(n597), .A2(n593), .A4(n282), .S0(n299), 
        .S1(n323), .Y(n424) );
  MUX41X1_HVT U186 ( .A1(n285), .A3(n567), .A2(n532), .A4(n560), .S0(n324), 
        .S1(n272), .Y(n418) );
  MUX41X1_HVT U189 ( .A1(n416), .A3(n592), .A2(n417), .A4(n367), .S0(n299), 
        .S1(n323), .Y(n415) );
  MUX41X1_HVT U193 ( .A1(n564), .A3(n571), .A2(n557), .A4(n413), .S0(n323), 
        .S1(n272), .Y(n412) );
  MUX41X1_HVT U194 ( .A1(n565), .A3(n263), .A2(n378), .A4(n310), .S0(n299), 
        .S1(n323), .Y(n411) );
  MUX41X1_HVT U195 ( .A1(n599), .A3(n372), .A2(n315), .A4(n569), .S0(n323), 
        .S1(n326), .Y(n410) );
  AO21X1_HVT U197 ( .A1(n287), .A2(n300), .A3(n369), .Y(n408) );
  MUX41X1_HVT U199 ( .A1(n407), .A3(n411), .A2(n410), .A4(n412), .S0(n308), 
        .S1(n298), .Y(n406) );
  OA21X1_HVT U201 ( .A1(n598), .A2(n329), .A3(n359), .Y(n404) );
  MUX41X1_HVT U203 ( .A1(n570), .A3(n361), .A2(n594), .A4(n574), .S0(n324), 
        .S1(n325), .Y(n402) );
  MUX41X1_HVT U204 ( .A1(n550), .A3(n593), .A2(n262), .A4(n583), .S0(n323), 
        .S1(n272), .Y(n401) );
  MUX41X1_HVT U205 ( .A1(n273), .A3(n603), .A2(n380), .A4(n355), .S0(n324), 
        .S1(n325), .Y(n400) );
  MUX41X1_HVT U206 ( .A1(n400), .A3(n402), .A2(n401), .A4(n403), .S0(n308), 
        .S1(n298), .Y(n399) );
  MUX21X2_HVT U207 ( .A1(n399), .A2(n406), .S0(in[6]), .Y(out[7]) );
  NAND2X0_HVT U208 ( .A1(n321), .A2(n312), .Y(n492) );
  NAND2X0_HVT U212 ( .A1(n321), .A2(n311), .Y(n549) );
  NAND2X0_HVT U214 ( .A1(n599), .A2(n255), .Y(n398) );
  NAND2X0_HVT U215 ( .A1(n492), .A2(n311), .Y(n397) );
  NAND2X0_HVT U218 ( .A1(n382), .A2(n321), .Y(n451) );
  NAND2X0_HVT U220 ( .A1(n300), .A2(n398), .Y(n524) );
  XNOR2X2_HVT U1 ( .A1(n241), .A2(in[3]), .Y(n23) );
  INVX8_HVT U2 ( .A(n23), .Y(n599) );
  NBUFFX2_HVT U6 ( .A(n23), .Y(n304) );
  MUX21X2_HVT U7 ( .A1(n604), .A2(n514), .S0(n289), .Y(n513) );
  XNOR2X2_HVT U8 ( .A1(n329), .A2(n317), .Y(n289) );
  MUX21X1_HVT U9 ( .A1(n583), .A2(n360), .S0(n300), .Y(n464) );
  INVX1_HVT U10 ( .A(n583), .Y(n348) );
  MUX21X2_HVT U11 ( .A1(n301), .A2(n303), .S0(n216), .Y(n589) );
  MUX21X2_HVT U12 ( .A1(n309), .A2(n304), .S0(n217), .Y(n583) );
  IBUFFX2_HVT U14 ( .A(n329), .Y(n326) );
  MUX21X1_HVT U16 ( .A1(n210), .A2(n386), .S0(n266), .Y(n50) );
  IBUFFX16_HVT U17 ( .A(n311), .Y(n210) );
  INVX1_HVT U18 ( .A(n266), .Y(n318) );
  NAND2X0_HVT U19 ( .A1(n546), .A2(n211), .Y(n212) );
  NAND2X0_HVT U20 ( .A1(n548), .A2(n257), .Y(n213) );
  NAND2X0_HVT U22 ( .A1(n212), .A2(n213), .Y(n545) );
  IBUFFX2_HVT U23 ( .A(n257), .Y(n211) );
  IBUFFX16_HVT U25 ( .A(n319), .Y(n216) );
  IBUFFX16_HVT U26 ( .A(n319), .Y(n217) );
  INVX1_HVT U27 ( .A(n562), .Y(n246) );
  MUX21X2_HVT U28 ( .A1(n408), .A2(n409), .S0(n218), .Y(n407) );
  IBUFFX16_HVT U29 ( .A(n294), .Y(n218) );
  NAND2X0_HVT U30 ( .A1(n475), .A2(n219), .Y(n229) );
  NAND2X0_HVT U31 ( .A1(n476), .A2(n233), .Y(n231) );
  NAND2X0_HVT U32 ( .A1(n229), .A2(n231), .Y(n474) );
  INVX0_HVT U34 ( .A(n233), .Y(n219) );
  MUX21X1_HVT U36 ( .A1(n479), .A2(n480), .S0(n271), .Y(n476) );
  INVX1_HVT U37 ( .A(n239), .Y(n233) );
  XOR2X1_HVT U38 ( .A1(n599), .A2(n265), .Y(n232) );
  IBUFFX16_HVT U39 ( .A(n232), .Y(n560) );
  IBUFFX2_HVT U40 ( .A(n265), .Y(n317) );
  MUX41X1_HVT U41 ( .A1(n310), .A3(n366), .A2(n302), .A4(n348), .S0(n234), 
        .S1(n330), .Y(n459) );
  IBUFFX16_HVT U43 ( .A(n292), .Y(n234) );
  INVX0_HVT U44 ( .A(in[1]), .Y(n322) );
  INVX0_HVT U45 ( .A(in[1]), .Y(n266) );
  NBUFFX4_HVT U46 ( .A(n23), .Y(n303) );
  INVX4_HVT U47 ( .A(n330), .Y(n327) );
  INVX4_HVT U48 ( .A(in[7]), .Y(n330) );
  MUX21X2_HVT U49 ( .A1(n512), .A2(n513), .S0(n295), .Y(n510) );
  MUX21X2_HVT U50 ( .A1(n602), .A2(n464), .S0(n235), .Y(n463) );
  IBUFFX16_HVT U52 ( .A(n295), .Y(n235) );
  MUX21X2_HVT U54 ( .A1(n282), .A2(n589), .S0(n271), .Y(n405) );
  AO21X2_HVT U55 ( .A1(n295), .A2(n310), .A3(n599), .Y(n484) );
  NAND2X0_HVT U59 ( .A1(n542), .A2(n236), .Y(n237) );
  NAND2X0_HVT U60 ( .A1(n544), .A2(n291), .Y(n238) );
  NAND2X0_HVT U63 ( .A1(n237), .A2(n238), .Y(n541) );
  IBUFFX2_HVT U64 ( .A(n291), .Y(n236) );
  MUX21X2_HVT U65 ( .A1(n363), .A2(n50), .S0(n300), .Y(n409) );
  IBUFFX16_HVT U67 ( .A(in[5]), .Y(n239) );
  INVX0_HVT U69 ( .A(in[1]), .Y(n265) );
  MUX21X2_HVT U70 ( .A1(n496), .A2(n506), .S0(in[6]), .Y(out[2]) );
  INVX1_HVT U71 ( .A(n329), .Y(n272) );
  AO21X1_HVT U72 ( .A1(n266), .A2(n382), .A3(n329), .Y(n502) );
  INVX2_HVT U76 ( .A(in[7]), .Y(n329) );
  INVX1_HVT U79 ( .A(n245), .Y(n535) );
  INVX0_HVT U81 ( .A(n306), .Y(n240) );
  INVX0_HVT U87 ( .A(in[4]), .Y(n241) );
  NBUFFX2_HVT U88 ( .A(n386), .Y(n306) );
  INVX0_HVT U89 ( .A(n322), .Y(n242) );
  INVX1_HVT U91 ( .A(n322), .Y(n243) );
  INVX1_HVT U92 ( .A(n322), .Y(n319) );
  MUX21X2_HVT U94 ( .A1(n423), .A2(n414), .S0(n244), .Y(out[6]) );
  IBUFFX16_HVT U95 ( .A(in[6]), .Y(n244) );
  INVX0_HVT U99 ( .A(n589), .Y(n343) );
  MUX21X1_HVT U100 ( .A1(n301), .A2(n311), .S0(n266), .Y(n394) );
  MUX21X1_HVT U102 ( .A1(n247), .A2(n246), .S0(n248), .Y(n245) );
  IBUFFX16_HVT U104 ( .A(n536), .Y(n247) );
  IBUFFX16_HVT U107 ( .A(n257), .Y(n248) );
  MUX41X1_HVT U108 ( .A1(n342), .A3(n365), .A2(n338), .A4(n543), .S0(n330), 
        .S1(n249), .Y(n542) );
  IBUFFX16_HVT U111 ( .A(n297), .Y(n249) );
  MUX21X1_HVT U112 ( .A1(n301), .A2(n312), .S0(n255), .Y(n594) );
  MUX21X1_HVT U113 ( .A1(n243), .A2(n594), .S0(n251), .Y(n250) );
  IBUFFX16_HVT U116 ( .A(n250), .Y(n540) );
  IBUFFX16_HVT U117 ( .A(n298), .Y(n251) );
  INVX2_HVT U118 ( .A(n322), .Y(n320) );
  MUX41X1_HVT U119 ( .A1(n551), .A3(n541), .A2(n545), .A4(n537), .S0(n252), 
        .S1(n253), .Y(out[0]) );
  IBUFFX16_HVT U120 ( .A(in[6]), .Y(n252) );
  IBUFFX16_HVT U121 ( .A(n308), .Y(n253) );
  INVX0_HVT U122 ( .A(n597), .Y(n341) );
  MUX21X1_HVT U124 ( .A1(n309), .A2(n519), .S0(n271), .Y(n421) );
  OA21X1_HVT U126 ( .A1(n572), .A2(n329), .A3(n348), .Y(n420) );
  INVX0_HVT U127 ( .A(n262), .Y(n572) );
  XOR2X1_HVT U128 ( .A1(n329), .A2(n579), .Y(n562) );
  INVX1_HVT U129 ( .A(in[0]), .Y(n254) );
  INVX1_HVT U130 ( .A(n295), .Y(n268) );
  INVX1_HVT U133 ( .A(n296), .Y(n267) );
  INVX1_HVT U134 ( .A(n328), .Y(n271) );
  INVX0_HVT U135 ( .A(n264), .Y(n324) );
  INVX0_HVT U137 ( .A(n293), .Y(n264) );
  MUX21X1_HVT U138 ( .A1(n312), .A2(n309), .S0(n319), .Y(n597) );
  IBUFFX2_HVT U141 ( .A(n567), .Y(n360) );
  MUX41X1_HVT U142 ( .A1(n419), .A3(n422), .A2(n415), .A4(n418), .S0(n298), 
        .S1(n254), .Y(n414) );
  MUX21X2_HVT U143 ( .A1(n486), .A2(n483), .S0(n267), .Y(n482) );
  INVX0_HVT U145 ( .A(n256), .Y(n595) );
  IBUFFX2_HVT U149 ( .A(n586), .Y(n346) );
  MUX21X2_HVT U150 ( .A1(n420), .A2(n421), .S0(n294), .Y(n419) );
  NBUFFX2_HVT U152 ( .A(n322), .Y(n255) );
  MUX41X1_HVT U155 ( .A1(n290), .A3(n547), .A2(n288), .A4(n345), .S0(n327), 
        .S1(n297), .Y(n546) );
  MUX21X1_HVT U156 ( .A1(n309), .A2(n315), .S0(n319), .Y(n256) );
  NAND2X0_HVT U157 ( .A1(n556), .A2(n257), .Y(n258) );
  NAND2X0_HVT U161 ( .A1(n552), .A2(n268), .Y(n259) );
  NAND2X0_HVT U164 ( .A1(n258), .A2(n259), .Y(n551) );
  INVX0_HVT U169 ( .A(n268), .Y(n257) );
  INVX0_HVT U171 ( .A(n571), .Y(n334) );
  NAND2X0_HVT U173 ( .A1(n554), .A2(n271), .Y(n260) );
  NAND2X0_HVT U175 ( .A1(n555), .A2(n299), .Y(n261) );
  NAND2X0_HVT U181 ( .A1(n260), .A2(n261), .Y(n552) );
  MUX21X1_HVT U182 ( .A1(n309), .A2(n571), .S0(n296), .Y(n555) );
  MUX21X1_HVT U183 ( .A1(n307), .A2(n301), .S0(n266), .Y(n413) );
  MUX21X2_HVT U184 ( .A1(n384), .A2(n372), .S0(n328), .Y(n536) );
  MUX21X1_HVT U185 ( .A1(n309), .A2(n315), .S0(n255), .Y(n262) );
  INVX2_HVT U187 ( .A(n265), .Y(n321) );
  MUX21X1_HVT U188 ( .A1(n384), .A2(n385), .S0(n255), .Y(n579) );
  INVX0_HVT U190 ( .A(n389), .Y(n378) );
  MUX41X1_HVT U191 ( .A1(n428), .A3(n425), .A2(n426), .A4(n424), .S0(n254), 
        .S1(n267), .Y(n423) );
  INVX0_HVT U192 ( .A(n276), .Y(n263) );
  INVX1_HVT U196 ( .A(n579), .Y(n276) );
  MUX41X1_HVT U198 ( .A1(n356), .A3(n461), .A2(n359), .A4(n581), .S0(n264), 
        .S1(n330), .Y(n460) );
  INVX1_HVT U200 ( .A(n585), .Y(n347) );
  MUX21X1_HVT U202 ( .A1(n311), .A2(n585), .S0(n271), .Y(n526) );
  MUX41X1_HVT U209 ( .A1(n523), .A3(n520), .A2(n522), .A4(n518), .S0(n254), 
        .S1(n267), .Y(n517) );
  INVX1_HVT U210 ( .A(n394), .Y(n372) );
  MUX21X2_HVT U211 ( .A1(n525), .A2(n526), .S0(n268), .Y(n523) );
  IBUFFX2_HVT U213 ( .A(n574), .Y(n356) );
  NAND2X0_HVT U216 ( .A1(n404), .A2(n268), .Y(n269) );
  NAND2X0_HVT U217 ( .A1(n405), .A2(n257), .Y(n270) );
  NAND2X0_HVT U219 ( .A1(n269), .A2(n270), .Y(n403) );
  MUX21X2_HVT U221 ( .A1(n517), .A2(n527), .S0(in[6]), .Y(out[1]) );
  MUX41X1_HVT U222 ( .A1(n575), .A3(n349), .A2(n487), .A4(n593), .S0(n268), 
        .S1(n271), .Y(n486) );
  INVX1_HVT U223 ( .A(n329), .Y(n325) );
  INVX0_HVT U224 ( .A(n274), .Y(n466) );
  MUX21X1_HVT U225 ( .A1(n355), .A2(n591), .S0(n295), .Y(n505) );
  INVX0_HVT U226 ( .A(in[6]), .Y(n277) );
  INVX0_HVT U227 ( .A(n600), .Y(n275) );
  IBUFFX2_HVT U228 ( .A(n386), .Y(n273) );
  INVX1_HVT U229 ( .A(in[4]), .Y(n386) );
  MUX41X1_HVT U230 ( .A1(n276), .A3(n275), .A2(n310), .A4(n389), .S0(n264), 
        .S1(n330), .Y(n274) );
  AND3X2_HVT U231 ( .A1(n294), .A2(n255), .A3(n273), .Y(n472) );
  MUX41X1_HVT U232 ( .A1(n350), .A3(n362), .A2(n601), .A4(n360), .S0(n330), 
        .S1(n264), .Y(n422) );
  MUX21X2_HVT U233 ( .A1(n430), .A2(n442), .S0(in[6]), .Y(out[5]) );
  MUX21X2_HVT U234 ( .A1(n462), .A2(n454), .S0(n277), .Y(out[4]) );
  IBUFFX2_HVT U235 ( .A(n330), .Y(n328) );
  XOR2X1_HVT U236 ( .A1(n264), .A2(n330), .Y(n559) );
  NAND2X0_HVT U237 ( .A1(n604), .A2(n278), .Y(n279) );
  NAND2X0_HVT U238 ( .A1(n490), .A2(n281), .Y(n280) );
  NAND2X0_HVT U239 ( .A1(n280), .A2(n279), .Y(n489) );
  INVX0_HVT U240 ( .A(n281), .Y(n278) );
  XNOR2X1_HVT U241 ( .A1(n317), .A2(n324), .Y(n281) );
  INVX0_HVT U242 ( .A(in[3]), .Y(n383) );
  MUX21X2_HVT U243 ( .A1(n286), .A2(n505), .S0(n559), .Y(n504) );
  INVX1_HVT U244 ( .A(n601), .Y(n381) );
  MUX21X1_HVT U245 ( .A1(n284), .A2(n343), .S0(n292), .Y(n471) );
  NBUFFX2_HVT U246 ( .A(n23), .Y(n302) );
  AND2X1_HVT U247 ( .A1(n304), .A2(n549), .Y(n282) );
  INVX1_HVT U248 ( .A(n313), .Y(n385) );
  MUX21X1_HVT U249 ( .A1(n381), .A2(n384), .S0(in[5]), .Y(n553) );
  NBUFFX2_HVT U250 ( .A(n601), .Y(n312) );
  MUX21X1_HVT U251 ( .A1(n341), .A2(n382), .S0(n298), .Y(n538) );
  MUX21X1_HVT U252 ( .A1(n575), .A2(n493), .S0(n292), .Y(n491) );
  AND2X1_HVT U253 ( .A1(n314), .A2(n532), .Y(n283) );
  MUX21X1_HVT U254 ( .A1(n304), .A2(n384), .S0(n321), .Y(n598) );
  MUX21X1_HVT U255 ( .A1(n314), .A2(n303), .S0(n320), .Y(n565) );
  MUX21X1_HVT U256 ( .A1(n302), .A2(n307), .S0(n318), .Y(n501) );
  MUX21X1_HVT U257 ( .A1(n381), .A2(n385), .S0(n243), .Y(n429) );
  MUX21X1_HVT U258 ( .A1(n312), .A2(n599), .S0(n242), .Y(n569) );
  MUX21X1_HVT U259 ( .A1(n384), .A2(n303), .S0(n318), .Y(n441) );
  MUX21X1_HVT U260 ( .A1(n303), .A2(n381), .S0(n318), .Y(n509) );
  MUX21X1_HVT U261 ( .A1(n599), .A2(n382), .S0(n318), .Y(n389) );
  MUX21X1_HVT U262 ( .A1(n599), .A2(n385), .S0(n242), .Y(n581) );
  MUX21X1_HVT U263 ( .A1(n599), .A2(n307), .S0(n242), .Y(n529) );
  MUX21X1_HVT U264 ( .A1(n301), .A2(n599), .S0(n318), .Y(n392) );
  MUX21X1_HVT U265 ( .A1(n384), .A2(n381), .S0(n243), .Y(n568) );
  MUX21X1_HVT U266 ( .A1(n301), .A2(n385), .S0(n320), .Y(n566) );
  MUX21X1_HVT U267 ( .A1(n307), .A2(n381), .S0(n243), .Y(n577) );
  MUX21X1_HVT U268 ( .A1(n382), .A2(n381), .S0(n242), .Y(n587) );
  MUX21X1_HVT U269 ( .A1(n354), .A2(n468), .S0(n294), .Y(n467) );
  MUX21X1_HVT U270 ( .A1(n377), .A2(n311), .S0(n300), .Y(n468) );
  MUX21X1_HVT U271 ( .A1(n484), .A2(n485), .S0(n300), .Y(n483) );
  MUX21X1_HVT U272 ( .A1(n334), .A2(n262), .S0(n292), .Y(n485) );
  MUX21X1_HVT U273 ( .A1(n312), .A2(n311), .S0(n242), .Y(n516) );
  NAND2X0_HVT U274 ( .A1(n305), .A2(n383), .Y(n601) );
  MUX21X1_HVT U275 ( .A1(n381), .A2(n306), .S0(n317), .Y(n390) );
  NBUFFX2_HVT U276 ( .A(n604), .Y(n313) );
  INVX1_HVT U277 ( .A(n315), .Y(n384) );
  MUX21X1_HVT U278 ( .A1(n333), .A2(n481), .S0(n293), .Y(n480) );
  MUX21X1_HVT U279 ( .A1(n306), .A2(n301), .S0(n318), .Y(n481) );
  NBUFFX2_HVT U280 ( .A(n604), .Y(n314) );
  XOR2X1_HVT U281 ( .A1(n317), .A2(n382), .Y(n561) );
  MUX21X1_HVT U282 ( .A1(n383), .A2(n316), .S0(n318), .Y(n416) );
  MUX21X1_HVT U283 ( .A1(n315), .A2(n314), .S0(n318), .Y(n417) );
  INVX1_HVT U284 ( .A(n310), .Y(n382) );
  MUX21X1_HVT U285 ( .A1(n314), .A2(n311), .S0(n319), .Y(n591) );
  MUX21X1_HVT U286 ( .A1(n601), .A2(n316), .S0(n317), .Y(n511) );
  XOR2X1_HVT U287 ( .A1(n313), .A2(n317), .Y(n557) );
  MUX21X1_HVT U288 ( .A1(n313), .A2(n306), .S0(n318), .Y(n396) );
  XNOR2X1_HVT U289 ( .A1(n601), .A2(n317), .Y(n284) );
  AND2X1_HVT U290 ( .A1(n321), .A2(n385), .Y(n285) );
  MUX21X1_HVT U291 ( .A1(n315), .A2(n311), .S0(n320), .Y(n575) );
  AND2X1_HVT U292 ( .A1(n316), .A2(n492), .Y(n286) );
  MUX21X1_HVT U293 ( .A1(n313), .A2(n312), .S0(n317), .Y(n388) );
  XNOR2X1_HVT U294 ( .A1(n315), .A2(n317), .Y(n287) );
  MUX21X1_HVT U295 ( .A1(n311), .A2(n306), .S0(n320), .Y(n534) );
  MUX21X1_HVT U296 ( .A1(n596), .A2(n316), .S0(n294), .Y(n478) );
  XOR2X1_HVT U297 ( .A1(n305), .A2(n317), .Y(n580) );
  NBUFFX2_HVT U298 ( .A(n328), .Y(n299) );
  NBUFFX2_HVT U299 ( .A(n328), .Y(n300) );
  NBUFFX2_HVT U300 ( .A(n383), .Y(n301) );
  NBUFFX2_HVT U301 ( .A(in[2]), .Y(n292) );
  NBUFFX2_HVT U302 ( .A(in[2]), .Y(n293) );
  NBUFFX2_HVT U303 ( .A(in[5]), .Y(n298) );
  NBUFFX2_HVT U304 ( .A(in[2]), .Y(n294) );
  NBUFFX2_HVT U305 ( .A(in[2]), .Y(n295) );
  NBUFFX2_HVT U306 ( .A(in[5]), .Y(n297) );
  NBUFFX2_HVT U307 ( .A(in[2]), .Y(n291) );
  NBUFFX2_HVT U308 ( .A(in[5]), .Y(n296) );
  NBUFFX2_HVT U309 ( .A(n386), .Y(n305) );
  MUX21X1_HVT U310 ( .A1(n503), .A2(n354), .S0(n294), .Y(n500) );
  XOR2X1_HVT U311 ( .A1(n317), .A2(n309), .Y(n558) );
  MUX21X1_HVT U312 ( .A1(n311), .A2(n304), .S0(n320), .Y(n498) );
  MUX21X1_HVT U313 ( .A1(n433), .A2(n432), .S0(n294), .Y(n431) );
  MUX21X1_HVT U314 ( .A1(n596), .A2(n372), .S0(n328), .Y(n433) );
  MUX21X1_HVT U315 ( .A1(n452), .A2(n453), .S0(n295), .Y(n450) );
  MUX21X1_HVT U316 ( .A1(n374), .A2(n382), .S0(n300), .Y(n453) );
  AND2X1_HVT U317 ( .A1(n304), .A2(n255), .Y(n288) );
  MUX21X1_HVT U318 ( .A1(n309), .A2(n381), .S0(n242), .Y(n567) );
  MUX21X1_HVT U319 ( .A1(n458), .A2(n457), .S0(n294), .Y(n456) );
  MUX21X1_HVT U320 ( .A1(n577), .A2(n337), .S0(n299), .Y(n458) );
  MUX21X1_HVT U321 ( .A1(n588), .A2(n356), .S0(n293), .Y(n470) );
  MUX21X1_HVT U322 ( .A1(n382), .A2(n385), .S0(n318), .Y(n438) );
  NAND2X0_HVT U323 ( .A1(in[3]), .A2(n307), .Y(n604) );
  NBUFFX2_HVT U324 ( .A(n386), .Y(n307) );
  NBUFFX2_HVT U325 ( .A(n605), .Y(n315) );
  MUX21X1_HVT U326 ( .A1(n385), .A2(n309), .S0(n319), .Y(n586) );
  MUX21X1_HVT U327 ( .A1(n357), .A2(n603), .S0(n293), .Y(n495) );
  MUX21X1_HVT U328 ( .A1(n446), .A2(n447), .S0(n295), .Y(n445) );
  MUX21X1_HVT U329 ( .A1(n448), .A2(n604), .S0(n289), .Y(n447) );
  MUX21X1_HVT U330 ( .A1(n568), .A2(n375), .S0(n299), .Y(n446) );
  XOR2X1_HVT U331 ( .A1(n317), .A2(n298), .Y(n563) );
  MUX21X1_HVT U332 ( .A1(n603), .A2(n266), .S0(n294), .Y(n477) );
  NBUFFX2_HVT U333 ( .A(n596), .Y(n310) );
  NBUFFX2_HVT U334 ( .A(n596), .Y(n311) );
  MUX21X1_HVT U335 ( .A1(n309), .A2(n382), .S0(n318), .Y(n393) );
  MUX21X1_HVT U336 ( .A1(n576), .A2(n397), .S0(n299), .Y(n391) );
  MUX21X1_HVT U337 ( .A1(n351), .A2(n576), .S0(n293), .Y(n473) );
  MUX21X1_HVT U338 ( .A1(n309), .A2(n306), .S0(n328), .Y(n514) );
  NBUFFX2_HVT U339 ( .A(n605), .Y(n316) );
  AND2X1_HVT U340 ( .A1(n301), .A2(n255), .Y(n290) );
  INVX1_HVT U341 ( .A(n268), .Y(n323) );
  MUX21X1_HVT U342 ( .A1(n381), .A2(n273), .S0(n242), .Y(n574) );
  NAND2X0_HVT U343 ( .A1(in[3]), .A2(n240), .Y(n605) );
  MUX21X1_HVT U344 ( .A1(n273), .A2(n599), .S0(n318), .Y(n395) );
  MUX21X1_HVT U345 ( .A1(n273), .A2(n384), .S0(n243), .Y(n570) );
  MUX21X1_HVT U346 ( .A1(n273), .A2(n382), .S0(n320), .Y(n588) );
  NAND2X0_HVT U347 ( .A1(in[4]), .A2(n383), .Y(n596) );
  MUX21X1_HVT U348 ( .A1(n273), .A2(n314), .S0(n319), .Y(n585) );
  MUX21X1_HVT U349 ( .A1(n316), .A2(n273), .S0(n320), .Y(n578) );
  MUX21X1_HVT U350 ( .A1(n309), .A2(n273), .S0(n292), .Y(n490) );
  MUX21X1_HVT U351 ( .A1(n273), .A2(n316), .S0(n243), .Y(n387) );
  MUX21X1_HVT U352 ( .A1(n301), .A2(n273), .S0(n243), .Y(n576) );
  NBUFFX2_HVT U353 ( .A(in[3]), .Y(n309) );
  NBUFFX2_HVT U354 ( .A(in[0]), .Y(n308) );
  INVX0_HVT U355 ( .A(n584), .Y(n331) );
  INVX0_HVT U356 ( .A(n582), .Y(n332) );
  INVX0_HVT U357 ( .A(n573), .Y(n333) );
  INVX0_HVT U358 ( .A(n435), .Y(n335) );
  INVX0_HVT U359 ( .A(n398), .Y(n336) );
  INVX0_HVT U360 ( .A(n603), .Y(n337) );
  INVX0_HVT U361 ( .A(n590), .Y(n338) );
  INVX0_HVT U362 ( .A(n602), .Y(n339) );
  INVX0_HVT U363 ( .A(n598), .Y(n340) );
  INVX0_HVT U364 ( .A(n591), .Y(n342) );
  INVX0_HVT U365 ( .A(n588), .Y(n344) );
  INVX0_HVT U366 ( .A(n587), .Y(n345) );
  INVX0_HVT U367 ( .A(n581), .Y(n349) );
  INVX0_HVT U368 ( .A(n580), .Y(n350) );
  INVX0_HVT U369 ( .A(n578), .Y(n351) );
  INVX0_HVT U370 ( .A(n577), .Y(n352) );
  INVX0_HVT U371 ( .A(n576), .Y(n353) );
  INVX0_HVT U372 ( .A(n391), .Y(n354) );
  INVX0_HVT U373 ( .A(n575), .Y(n355) );
  INVX0_HVT U374 ( .A(n570), .Y(n357) );
  INVX0_HVT U375 ( .A(n569), .Y(n358) );
  INVX0_HVT U376 ( .A(n568), .Y(n359) );
  INVX0_HVT U377 ( .A(n566), .Y(n361) );
  INVX0_HVT U378 ( .A(n565), .Y(n362) );
  INVX0_HVT U379 ( .A(n564), .Y(n363) );
  INVX0_HVT U380 ( .A(n532), .Y(n364) );
  INVX0_HVT U381 ( .A(n593), .Y(n365) );
  INVX0_HVT U382 ( .A(n492), .Y(n366) );
  INVX0_HVT U383 ( .A(n397), .Y(n367) );
  INVX0_HVT U384 ( .A(n549), .Y(n368) );
  INVX0_HVT U385 ( .A(n451), .Y(n369) );
  INVX0_HVT U386 ( .A(n396), .Y(n370) );
  INVX0_HVT U387 ( .A(n395), .Y(n371) );
  INVX0_HVT U388 ( .A(n393), .Y(n373) );
  INVX0_HVT U389 ( .A(n392), .Y(n374) );
  INVX0_HVT U390 ( .A(n511), .Y(n375) );
  INVX0_HVT U391 ( .A(n501), .Y(n376) );
  INVX0_HVT U392 ( .A(n390), .Y(n377) );
  INVX0_HVT U393 ( .A(n388), .Y(n379) );
  INVX0_HVT U394 ( .A(n387), .Y(n380) );
endmodule

