
module Get_key ( clk, rest, local_key, rount_no, key_round, done );
  input [127:0] local_key;
  input [3:0] rount_no;
  output [127:0] key_round;
  input clk, rest;
  output done;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192;
  wire   [3:0] round_number;
  wire   [127:0] prev_key;
  wire   [127:0] keyout;
  wire   [3:0] state;

  DFFX1_HVT \state_reg[0]  ( .D(n3797), .CLK(clk), .Q(state[0]), .QN(n1) );
  DFFX1_HVT \state_reg[3]  ( .D(n3796), .CLK(clk), .Q(state[3]), .QN(n4) );
  DFFX1_HVT \state_reg[2]  ( .D(n3794), .CLK(clk), .Q(state[2]), .QN(n2) );
  DFFX1_HVT \state_reg[1]  ( .D(n3795), .CLK(clk), .Q(state[1]), .QN(n3) );
  DFFX1_HVT done_reg ( .D(n3793), .CLK(clk), .Q(done) );
  DFFX1_HVT \round_number_reg[2]  ( .D(n3790), .CLK(clk), .Q(round_number[2])
         );
  DFFX1_HVT \round_number_reg[3]  ( .D(n3789), .CLK(clk), .Q(round_number[3])
         );
  DFFX1_HVT \round_number_reg[0]  ( .D(n3792), .CLK(clk), .Q(round_number[0])
         );
  DFFX1_HVT \round_number_reg[1]  ( .D(n3791), .CLK(clk), .Q(round_number[1])
         );
  DFFX1_HVT \prev_key_reg[0]  ( .D(n3788), .CLK(clk), .Q(prev_key[0]) );
  DFFX1_HVT \prev_key_reg[1]  ( .D(n3787), .CLK(clk), .Q(prev_key[1]) );
  DFFX1_HVT \prev_key_reg[2]  ( .D(n3786), .CLK(clk), .Q(prev_key[2]) );
  DFFX1_HVT \prev_key_reg[3]  ( .D(n3785), .CLK(clk), .Q(prev_key[3]) );
  DFFX1_HVT \prev_key_reg[4]  ( .D(n3784), .CLK(clk), .Q(prev_key[4]) );
  DFFX1_HVT \prev_key_reg[5]  ( .D(n3783), .CLK(clk), .Q(prev_key[5]) );
  DFFX1_HVT \prev_key_reg[6]  ( .D(n3782), .CLK(clk), .Q(prev_key[6]) );
  DFFX1_HVT \prev_key_reg[7]  ( .D(n3781), .CLK(clk), .Q(prev_key[7]) );
  DFFX1_HVT \prev_key_reg[8]  ( .D(n3780), .CLK(clk), .Q(prev_key[8]) );
  DFFX1_HVT \prev_key_reg[9]  ( .D(n3779), .CLK(clk), .Q(prev_key[9]) );
  DFFX1_HVT \prev_key_reg[10]  ( .D(n3778), .CLK(clk), .Q(prev_key[10]) );
  DFFX1_HVT \prev_key_reg[11]  ( .D(n3777), .CLK(clk), .Q(prev_key[11]) );
  DFFX1_HVT \prev_key_reg[12]  ( .D(n3776), .CLK(clk), .Q(prev_key[12]) );
  DFFX1_HVT \prev_key_reg[13]  ( .D(n3775), .CLK(clk), .Q(prev_key[13]) );
  DFFX1_HVT \prev_key_reg[14]  ( .D(n3774), .CLK(clk), .Q(prev_key[14]) );
  DFFX1_HVT \prev_key_reg[15]  ( .D(n3773), .CLK(clk), .Q(prev_key[15]) );
  DFFX1_HVT \prev_key_reg[16]  ( .D(n3772), .CLK(clk), .Q(prev_key[16]) );
  DFFX1_HVT \prev_key_reg[17]  ( .D(n3771), .CLK(clk), .Q(prev_key[17]) );
  DFFX1_HVT \prev_key_reg[18]  ( .D(n3770), .CLK(clk), .Q(prev_key[18]) );
  DFFX1_HVT \prev_key_reg[19]  ( .D(n3769), .CLK(clk), .Q(prev_key[19]) );
  DFFX1_HVT \prev_key_reg[20]  ( .D(n3768), .CLK(clk), .Q(prev_key[20]) );
  DFFX1_HVT \prev_key_reg[21]  ( .D(n3767), .CLK(clk), .Q(prev_key[21]) );
  DFFX1_HVT \prev_key_reg[22]  ( .D(n3766), .CLK(clk), .Q(prev_key[22]) );
  DFFX1_HVT \prev_key_reg[23]  ( .D(n3765), .CLK(clk), .Q(prev_key[23]) );
  DFFX1_HVT \prev_key_reg[24]  ( .D(n3764), .CLK(clk), .Q(prev_key[24]) );
  DFFX1_HVT \prev_key_reg[25]  ( .D(n3763), .CLK(clk), .Q(prev_key[25]) );
  DFFX1_HVT \prev_key_reg[26]  ( .D(n3762), .CLK(clk), .Q(prev_key[26]) );
  DFFX1_HVT \prev_key_reg[27]  ( .D(n3761), .CLK(clk), .Q(prev_key[27]) );
  DFFX1_HVT \prev_key_reg[28]  ( .D(n3760), .CLK(clk), .Q(prev_key[28]) );
  DFFX1_HVT \prev_key_reg[29]  ( .D(n3759), .CLK(clk), .Q(prev_key[29]) );
  DFFX1_HVT \prev_key_reg[30]  ( .D(n3758), .CLK(clk), .Q(prev_key[30]) );
  DFFX1_HVT \prev_key_reg[31]  ( .D(n3757), .CLK(clk), .Q(prev_key[31]) );
  DFFX1_HVT \prev_key_reg[32]  ( .D(n3756), .CLK(clk), .Q(prev_key[32]) );
  DFFX1_HVT \prev_key_reg[33]  ( .D(n3755), .CLK(clk), .Q(prev_key[33]) );
  DFFX1_HVT \prev_key_reg[34]  ( .D(n3754), .CLK(clk), .Q(prev_key[34]) );
  DFFX1_HVT \prev_key_reg[35]  ( .D(n3753), .CLK(clk), .Q(prev_key[35]) );
  DFFX1_HVT \prev_key_reg[36]  ( .D(n3752), .CLK(clk), .Q(prev_key[36]) );
  DFFX1_HVT \prev_key_reg[37]  ( .D(n3751), .CLK(clk), .Q(prev_key[37]) );
  DFFX1_HVT \prev_key_reg[38]  ( .D(n3750), .CLK(clk), .Q(prev_key[38]) );
  DFFX1_HVT \prev_key_reg[39]  ( .D(n3749), .CLK(clk), .Q(prev_key[39]) );
  DFFX1_HVT \prev_key_reg[40]  ( .D(n3748), .CLK(clk), .Q(prev_key[40]) );
  DFFX1_HVT \prev_key_reg[41]  ( .D(n3747), .CLK(clk), .Q(prev_key[41]) );
  DFFX1_HVT \prev_key_reg[42]  ( .D(n3746), .CLK(clk), .Q(prev_key[42]) );
  DFFX1_HVT \prev_key_reg[43]  ( .D(n3745), .CLK(clk), .Q(prev_key[43]) );
  DFFX1_HVT \prev_key_reg[44]  ( .D(n3744), .CLK(clk), .Q(prev_key[44]) );
  DFFX1_HVT \prev_key_reg[45]  ( .D(n3743), .CLK(clk), .Q(prev_key[45]) );
  DFFX1_HVT \prev_key_reg[46]  ( .D(n3742), .CLK(clk), .Q(prev_key[46]) );
  DFFX1_HVT \prev_key_reg[47]  ( .D(n3741), .CLK(clk), .Q(prev_key[47]) );
  DFFX1_HVT \prev_key_reg[48]  ( .D(n3740), .CLK(clk), .Q(prev_key[48]) );
  DFFX1_HVT \prev_key_reg[49]  ( .D(n3739), .CLK(clk), .Q(prev_key[49]) );
  DFFX1_HVT \prev_key_reg[50]  ( .D(n3738), .CLK(clk), .Q(prev_key[50]) );
  DFFX1_HVT \prev_key_reg[51]  ( .D(n3737), .CLK(clk), .Q(prev_key[51]) );
  DFFX1_HVT \prev_key_reg[52]  ( .D(n3736), .CLK(clk), .Q(prev_key[52]) );
  DFFX1_HVT \prev_key_reg[53]  ( .D(n3735), .CLK(clk), .Q(prev_key[53]) );
  DFFX1_HVT \prev_key_reg[54]  ( .D(n3734), .CLK(clk), .Q(prev_key[54]) );
  DFFX1_HVT \prev_key_reg[55]  ( .D(n3733), .CLK(clk), .Q(prev_key[55]) );
  DFFX1_HVT \prev_key_reg[56]  ( .D(n3732), .CLK(clk), .Q(prev_key[56]) );
  DFFX1_HVT \prev_key_reg[57]  ( .D(n3731), .CLK(clk), .Q(prev_key[57]) );
  DFFX1_HVT \prev_key_reg[58]  ( .D(n3730), .CLK(clk), .Q(prev_key[58]) );
  DFFX1_HVT \prev_key_reg[59]  ( .D(n3729), .CLK(clk), .Q(prev_key[59]) );
  DFFX1_HVT \prev_key_reg[60]  ( .D(n3728), .CLK(clk), .Q(prev_key[60]) );
  DFFX1_HVT \prev_key_reg[61]  ( .D(n3727), .CLK(clk), .Q(prev_key[61]) );
  DFFX1_HVT \prev_key_reg[62]  ( .D(n3726), .CLK(clk), .Q(prev_key[62]) );
  DFFX1_HVT \prev_key_reg[63]  ( .D(n3725), .CLK(clk), .Q(prev_key[63]) );
  DFFX1_HVT \prev_key_reg[64]  ( .D(n3724), .CLK(clk), .Q(prev_key[64]) );
  DFFX1_HVT \prev_key_reg[65]  ( .D(n3723), .CLK(clk), .Q(prev_key[65]) );
  DFFX1_HVT \prev_key_reg[66]  ( .D(n3722), .CLK(clk), .Q(prev_key[66]) );
  DFFX1_HVT \prev_key_reg[67]  ( .D(n3721), .CLK(clk), .Q(prev_key[67]) );
  DFFX1_HVT \prev_key_reg[68]  ( .D(n3720), .CLK(clk), .Q(prev_key[68]) );
  DFFX1_HVT \prev_key_reg[69]  ( .D(n3719), .CLK(clk), .Q(prev_key[69]) );
  DFFX1_HVT \prev_key_reg[70]  ( .D(n3718), .CLK(clk), .Q(prev_key[70]) );
  DFFX1_HVT \prev_key_reg[71]  ( .D(n3717), .CLK(clk), .Q(prev_key[71]) );
  DFFX1_HVT \prev_key_reg[72]  ( .D(n3716), .CLK(clk), .Q(prev_key[72]) );
  DFFX1_HVT \prev_key_reg[73]  ( .D(n3715), .CLK(clk), .Q(prev_key[73]) );
  DFFX1_HVT \prev_key_reg[74]  ( .D(n3714), .CLK(clk), .Q(prev_key[74]) );
  DFFX1_HVT \prev_key_reg[75]  ( .D(n3713), .CLK(clk), .Q(prev_key[75]) );
  DFFX1_HVT \prev_key_reg[76]  ( .D(n3712), .CLK(clk), .Q(prev_key[76]) );
  DFFX1_HVT \prev_key_reg[77]  ( .D(n3711), .CLK(clk), .Q(prev_key[77]) );
  DFFX1_HVT \prev_key_reg[78]  ( .D(n3710), .CLK(clk), .Q(prev_key[78]) );
  DFFX1_HVT \prev_key_reg[79]  ( .D(n3709), .CLK(clk), .Q(prev_key[79]) );
  DFFX1_HVT \prev_key_reg[80]  ( .D(n3708), .CLK(clk), .Q(prev_key[80]) );
  DFFX1_HVT \prev_key_reg[81]  ( .D(n3707), .CLK(clk), .Q(prev_key[81]) );
  DFFX1_HVT \prev_key_reg[82]  ( .D(n3706), .CLK(clk), .Q(prev_key[82]) );
  DFFX1_HVT \prev_key_reg[83]  ( .D(n3705), .CLK(clk), .Q(prev_key[83]) );
  DFFX1_HVT \prev_key_reg[84]  ( .D(n3704), .CLK(clk), .Q(prev_key[84]) );
  DFFX1_HVT \prev_key_reg[85]  ( .D(n3703), .CLK(clk), .Q(prev_key[85]) );
  DFFX1_HVT \prev_key_reg[86]  ( .D(n3702), .CLK(clk), .Q(prev_key[86]) );
  DFFX1_HVT \prev_key_reg[87]  ( .D(n3701), .CLK(clk), .Q(prev_key[87]) );
  DFFX1_HVT \prev_key_reg[88]  ( .D(n3700), .CLK(clk), .Q(prev_key[88]) );
  DFFX1_HVT \prev_key_reg[89]  ( .D(n3699), .CLK(clk), .Q(prev_key[89]) );
  DFFX1_HVT \prev_key_reg[90]  ( .D(n3698), .CLK(clk), .Q(prev_key[90]) );
  DFFX1_HVT \prev_key_reg[91]  ( .D(n3697), .CLK(clk), .Q(prev_key[91]) );
  DFFX1_HVT \prev_key_reg[92]  ( .D(n3696), .CLK(clk), .Q(prev_key[92]) );
  DFFX1_HVT \prev_key_reg[93]  ( .D(n3695), .CLK(clk), .Q(prev_key[93]) );
  DFFX1_HVT \prev_key_reg[94]  ( .D(n3694), .CLK(clk), .Q(prev_key[94]) );
  DFFX1_HVT \prev_key_reg[95]  ( .D(n3693), .CLK(clk), .Q(prev_key[95]) );
  DFFX1_HVT \prev_key_reg[96]  ( .D(n3692), .CLK(clk), .Q(prev_key[96]) );
  DFFX1_HVT \prev_key_reg[97]  ( .D(n3691), .CLK(clk), .Q(prev_key[97]) );
  DFFX1_HVT \prev_key_reg[98]  ( .D(n3690), .CLK(clk), .Q(prev_key[98]) );
  DFFX1_HVT \prev_key_reg[99]  ( .D(n3689), .CLK(clk), .Q(prev_key[99]) );
  DFFX1_HVT \prev_key_reg[100]  ( .D(n3688), .CLK(clk), .Q(prev_key[100]) );
  DFFX1_HVT \prev_key_reg[101]  ( .D(n3687), .CLK(clk), .Q(prev_key[101]) );
  DFFX1_HVT \prev_key_reg[102]  ( .D(n3686), .CLK(clk), .Q(prev_key[102]) );
  DFFX1_HVT \prev_key_reg[103]  ( .D(n3685), .CLK(clk), .Q(prev_key[103]) );
  DFFX1_HVT \prev_key_reg[104]  ( .D(n3684), .CLK(clk), .Q(prev_key[104]) );
  DFFX1_HVT \prev_key_reg[105]  ( .D(n3683), .CLK(clk), .Q(prev_key[105]) );
  DFFX1_HVT \prev_key_reg[106]  ( .D(n3682), .CLK(clk), .Q(prev_key[106]) );
  DFFX1_HVT \prev_key_reg[107]  ( .D(n3681), .CLK(clk), .Q(prev_key[107]) );
  DFFX1_HVT \prev_key_reg[108]  ( .D(n3680), .CLK(clk), .Q(prev_key[108]) );
  DFFX1_HVT \prev_key_reg[109]  ( .D(n3679), .CLK(clk), .Q(prev_key[109]) );
  DFFX1_HVT \prev_key_reg[110]  ( .D(n3678), .CLK(clk), .Q(prev_key[110]) );
  DFFX1_HVT \prev_key_reg[111]  ( .D(n3677), .CLK(clk), .Q(prev_key[111]) );
  DFFX1_HVT \prev_key_reg[112]  ( .D(n3676), .CLK(clk), .Q(prev_key[112]) );
  DFFX1_HVT \prev_key_reg[113]  ( .D(n3675), .CLK(clk), .Q(prev_key[113]) );
  DFFX1_HVT \prev_key_reg[114]  ( .D(n3674), .CLK(clk), .Q(prev_key[114]) );
  DFFX1_HVT \prev_key_reg[115]  ( .D(n3673), .CLK(clk), .Q(prev_key[115]) );
  DFFX1_HVT \prev_key_reg[116]  ( .D(n3672), .CLK(clk), .Q(prev_key[116]) );
  DFFX1_HVT \prev_key_reg[117]  ( .D(n3671), .CLK(clk), .Q(prev_key[117]) );
  DFFX1_HVT \prev_key_reg[118]  ( .D(n3670), .CLK(clk), .Q(prev_key[118]) );
  DFFX1_HVT \prev_key_reg[119]  ( .D(n3669), .CLK(clk), .Q(prev_key[119]) );
  DFFX1_HVT \prev_key_reg[120]  ( .D(n3668), .CLK(clk), .Q(prev_key[120]) );
  DFFX1_HVT \prev_key_reg[121]  ( .D(n3667), .CLK(clk), .Q(prev_key[121]) );
  DFFX1_HVT \prev_key_reg[122]  ( .D(n3666), .CLK(clk), .Q(prev_key[122]) );
  DFFX1_HVT \prev_key_reg[123]  ( .D(n3665), .CLK(clk), .Q(prev_key[123]) );
  DFFX1_HVT \prev_key_reg[124]  ( .D(n3664), .CLK(clk), .Q(prev_key[124]) );
  DFFX1_HVT \prev_key_reg[125]  ( .D(n3663), .CLK(clk), .Q(prev_key[125]) );
  DFFX1_HVT \prev_key_reg[126]  ( .D(n3662), .CLK(clk), .Q(prev_key[126]) );
  DFFX1_HVT \prev_key_reg[127]  ( .D(n3661), .CLK(clk), .Q(prev_key[127]) );
  DFFX1_HVT \keys_reg[0][127]  ( .D(n3660), .CLK(clk), .Q(n4366), .QN(n19) );
  DFFX1_HVT \keys_reg[0][126]  ( .D(n3659), .CLK(clk), .Q(n4367), .QN(n20) );
  DFFX1_HVT \keys_reg[0][125]  ( .D(n3658), .CLK(clk), .Q(n4368), .QN(n21) );
  DFFX1_HVT \keys_reg[0][124]  ( .D(n3657), .CLK(clk), .Q(n4369), .QN(n22) );
  DFFX1_HVT \keys_reg[0][123]  ( .D(n3656), .CLK(clk), .Q(n4370), .QN(n23) );
  DFFX1_HVT \keys_reg[0][122]  ( .D(n3655), .CLK(clk), .Q(n4371), .QN(n24) );
  DFFX1_HVT \keys_reg[0][121]  ( .D(n3654), .CLK(clk), .Q(n4372), .QN(n25) );
  DFFX1_HVT \keys_reg[0][120]  ( .D(n3653), .CLK(clk), .Q(n4373), .QN(n26) );
  DFFX1_HVT \keys_reg[0][119]  ( .D(n3652), .CLK(clk), .Q(n4374), .QN(n27) );
  DFFX1_HVT \keys_reg[0][118]  ( .D(n3651), .CLK(clk), .Q(n4375), .QN(n28) );
  DFFX1_HVT \keys_reg[0][117]  ( .D(n3650), .CLK(clk), .Q(n4376), .QN(n29) );
  DFFX1_HVT \keys_reg[0][116]  ( .D(n3649), .CLK(clk), .Q(n4377), .QN(n30) );
  DFFX1_HVT \keys_reg[0][115]  ( .D(n3648), .CLK(clk), .Q(n4378), .QN(n31) );
  DFFX1_HVT \keys_reg[0][114]  ( .D(n3647), .CLK(clk), .Q(n4379), .QN(n32) );
  DFFX1_HVT \keys_reg[0][113]  ( .D(n3646), .CLK(clk), .Q(n4380), .QN(n33) );
  DFFX1_HVT \keys_reg[0][112]  ( .D(n3645), .CLK(clk), .Q(n4381), .QN(n34) );
  DFFX1_HVT \keys_reg[0][111]  ( .D(n3644), .CLK(clk), .Q(n4382), .QN(n35) );
  DFFX1_HVT \keys_reg[0][110]  ( .D(n3643), .CLK(clk), .Q(n4383), .QN(n36) );
  DFFX1_HVT \keys_reg[0][109]  ( .D(n3642), .CLK(clk), .Q(n4384), .QN(n37) );
  DFFX1_HVT \keys_reg[0][108]  ( .D(n3641), .CLK(clk), .Q(n4385), .QN(n38) );
  DFFX1_HVT \keys_reg[0][107]  ( .D(n3640), .CLK(clk), .Q(n4386), .QN(n39) );
  DFFX1_HVT \keys_reg[0][106]  ( .D(n3639), .CLK(clk), .Q(n4387), .QN(n40) );
  DFFX1_HVT \keys_reg[0][105]  ( .D(n3638), .CLK(clk), .Q(n4388), .QN(n41) );
  DFFX1_HVT \keys_reg[0][104]  ( .D(n3637), .CLK(clk), .Q(n4389), .QN(n42) );
  DFFX1_HVT \keys_reg[0][103]  ( .D(n3636), .CLK(clk), .Q(n4390), .QN(n43) );
  DFFX1_HVT \keys_reg[0][102]  ( .D(n3635), .CLK(clk), .Q(n4391), .QN(n44) );
  DFFX1_HVT \keys_reg[0][101]  ( .D(n3634), .CLK(clk), .Q(n4392), .QN(n45) );
  DFFX1_HVT \keys_reg[0][100]  ( .D(n3633), .CLK(clk), .Q(n4393), .QN(n46) );
  DFFX1_HVT \keys_reg[0][99]  ( .D(n3632), .CLK(clk), .Q(n4394), .QN(n47) );
  DFFX1_HVT \keys_reg[0][98]  ( .D(n3631), .CLK(clk), .Q(n4395), .QN(n48) );
  DFFX1_HVT \keys_reg[0][97]  ( .D(n3630), .CLK(clk), .Q(n4396), .QN(n49) );
  DFFX1_HVT \keys_reg[0][96]  ( .D(n3629), .CLK(clk), .Q(n4397), .QN(n50) );
  DFFX1_HVT \keys_reg[0][95]  ( .D(n3628), .CLK(clk), .Q(n4398), .QN(n51) );
  DFFX1_HVT \keys_reg[0][94]  ( .D(n3627), .CLK(clk), .Q(n4399), .QN(n52) );
  DFFX1_HVT \keys_reg[0][93]  ( .D(n3626), .CLK(clk), .Q(n4400), .QN(n53) );
  DFFX1_HVT \keys_reg[0][92]  ( .D(n3625), .CLK(clk), .Q(n4401), .QN(n54) );
  DFFX1_HVT \keys_reg[0][91]  ( .D(n3624), .CLK(clk), .Q(n4402), .QN(n55) );
  DFFX1_HVT \keys_reg[0][90]  ( .D(n3623), .CLK(clk), .Q(n4403), .QN(n56) );
  DFFX1_HVT \keys_reg[0][89]  ( .D(n3622), .CLK(clk), .Q(n4404), .QN(n57) );
  DFFX1_HVT \keys_reg[0][88]  ( .D(n3621), .CLK(clk), .Q(n4405), .QN(n58) );
  DFFX1_HVT \keys_reg[0][87]  ( .D(n3620), .CLK(clk), .Q(n4406), .QN(n59) );
  DFFX1_HVT \keys_reg[0][86]  ( .D(n3619), .CLK(clk), .Q(n4407), .QN(n60) );
  DFFX1_HVT \keys_reg[0][85]  ( .D(n3618), .CLK(clk), .Q(n4408), .QN(n61) );
  DFFX1_HVT \keys_reg[0][84]  ( .D(n3617), .CLK(clk), .Q(n4409), .QN(n62) );
  DFFX1_HVT \keys_reg[0][83]  ( .D(n3616), .CLK(clk), .Q(n4410), .QN(n63) );
  DFFX1_HVT \keys_reg[0][82]  ( .D(n3615), .CLK(clk), .Q(n4411), .QN(n64) );
  DFFX1_HVT \keys_reg[0][81]  ( .D(n3614), .CLK(clk), .Q(n4412), .QN(n65) );
  DFFX1_HVT \keys_reg[0][80]  ( .D(n3613), .CLK(clk), .Q(n4413), .QN(n66) );
  DFFX1_HVT \keys_reg[0][79]  ( .D(n3612), .CLK(clk), .Q(n4414), .QN(n67) );
  DFFX1_HVT \keys_reg[0][78]  ( .D(n3611), .CLK(clk), .Q(n4415), .QN(n68) );
  DFFX1_HVT \keys_reg[0][77]  ( .D(n3610), .CLK(clk), .Q(n4416), .QN(n69) );
  DFFX1_HVT \keys_reg[0][76]  ( .D(n3609), .CLK(clk), .Q(n4417), .QN(n70) );
  DFFX1_HVT \keys_reg[0][75]  ( .D(n3608), .CLK(clk), .Q(n4418), .QN(n71) );
  DFFX1_HVT \keys_reg[0][74]  ( .D(n3607), .CLK(clk), .Q(n4419), .QN(n72) );
  DFFX1_HVT \keys_reg[0][73]  ( .D(n3606), .CLK(clk), .Q(n4420), .QN(n73) );
  DFFX1_HVT \keys_reg[0][72]  ( .D(n3605), .CLK(clk), .Q(n4421), .QN(n74) );
  DFFX1_HVT \keys_reg[0][71]  ( .D(n3604), .CLK(clk), .Q(n4422), .QN(n75) );
  DFFX1_HVT \keys_reg[0][70]  ( .D(n3603), .CLK(clk), .Q(n4423), .QN(n76) );
  DFFX1_HVT \keys_reg[0][69]  ( .D(n3602), .CLK(clk), .Q(n4424), .QN(n77) );
  DFFX1_HVT \keys_reg[0][68]  ( .D(n3601), .CLK(clk), .Q(n4425), .QN(n78) );
  DFFX1_HVT \keys_reg[0][67]  ( .D(n3600), .CLK(clk), .Q(n4426), .QN(n79) );
  DFFX1_HVT \keys_reg[0][66]  ( .D(n3599), .CLK(clk), .Q(n4427), .QN(n80) );
  DFFX1_HVT \keys_reg[0][65]  ( .D(n3598), .CLK(clk), .Q(n4428), .QN(n81) );
  DFFX1_HVT \keys_reg[0][64]  ( .D(n3597), .CLK(clk), .Q(n4429), .QN(n82) );
  DFFX1_HVT \keys_reg[0][63]  ( .D(n3596), .CLK(clk), .Q(n4430), .QN(n83) );
  DFFX1_HVT \keys_reg[0][62]  ( .D(n3595), .CLK(clk), .Q(n4431), .QN(n84) );
  DFFX1_HVT \keys_reg[0][61]  ( .D(n3594), .CLK(clk), .Q(n4432), .QN(n85) );
  DFFX1_HVT \keys_reg[0][60]  ( .D(n3593), .CLK(clk), .Q(n4433), .QN(n86) );
  DFFX1_HVT \keys_reg[0][59]  ( .D(n3592), .CLK(clk), .Q(n4434), .QN(n87) );
  DFFX1_HVT \keys_reg[0][58]  ( .D(n3591), .CLK(clk), .Q(n4435), .QN(n88) );
  DFFX1_HVT \keys_reg[0][57]  ( .D(n3590), .CLK(clk), .Q(n4436), .QN(n89) );
  DFFX1_HVT \keys_reg[0][56]  ( .D(n3589), .CLK(clk), .Q(n4437), .QN(n90) );
  DFFX1_HVT \keys_reg[0][55]  ( .D(n3588), .CLK(clk), .Q(n4438), .QN(n91) );
  DFFX1_HVT \keys_reg[0][54]  ( .D(n3587), .CLK(clk), .Q(n4439), .QN(n92) );
  DFFX1_HVT \keys_reg[0][53]  ( .D(n3586), .CLK(clk), .Q(n4440), .QN(n93) );
  DFFX1_HVT \keys_reg[0][52]  ( .D(n3585), .CLK(clk), .Q(n4441), .QN(n94) );
  DFFX1_HVT \keys_reg[0][51]  ( .D(n3584), .CLK(clk), .Q(n4442), .QN(n95) );
  DFFX1_HVT \keys_reg[0][50]  ( .D(n3583), .CLK(clk), .Q(n4443), .QN(n96) );
  DFFX1_HVT \keys_reg[0][49]  ( .D(n3582), .CLK(clk), .Q(n4444), .QN(n97) );
  DFFX1_HVT \keys_reg[0][48]  ( .D(n3581), .CLK(clk), .Q(n4445), .QN(n98) );
  DFFX1_HVT \keys_reg[0][47]  ( .D(n3580), .CLK(clk), .Q(n4446), .QN(n99) );
  DFFX1_HVT \keys_reg[0][46]  ( .D(n3579), .CLK(clk), .Q(n4447), .QN(n100) );
  DFFX1_HVT \keys_reg[0][45]  ( .D(n3578), .CLK(clk), .Q(n4448), .QN(n101) );
  DFFX1_HVT \keys_reg[0][44]  ( .D(n3577), .CLK(clk), .Q(n4449), .QN(n102) );
  DFFX1_HVT \keys_reg[0][43]  ( .D(n3576), .CLK(clk), .Q(n4450), .QN(n103) );
  DFFX1_HVT \keys_reg[0][42]  ( .D(n3575), .CLK(clk), .Q(n4451), .QN(n104) );
  DFFX1_HVT \keys_reg[0][41]  ( .D(n3574), .CLK(clk), .Q(n4452), .QN(n105) );
  DFFX1_HVT \keys_reg[0][40]  ( .D(n3573), .CLK(clk), .Q(n4453), .QN(n106) );
  DFFX1_HVT \keys_reg[0][39]  ( .D(n3572), .CLK(clk), .Q(n4454), .QN(n107) );
  DFFX1_HVT \keys_reg[0][38]  ( .D(n3571), .CLK(clk), .Q(n4455), .QN(n108) );
  DFFX1_HVT \keys_reg[0][37]  ( .D(n3570), .CLK(clk), .Q(n4456), .QN(n109) );
  DFFX1_HVT \keys_reg[0][36]  ( .D(n3569), .CLK(clk), .Q(n4457), .QN(n110) );
  DFFX1_HVT \keys_reg[0][35]  ( .D(n3568), .CLK(clk), .Q(n4458), .QN(n111) );
  DFFX1_HVT \keys_reg[0][34]  ( .D(n3567), .CLK(clk), .Q(n4459), .QN(n112) );
  DFFX1_HVT \keys_reg[0][33]  ( .D(n3566), .CLK(clk), .Q(n4460), .QN(n113) );
  DFFX1_HVT \keys_reg[0][32]  ( .D(n3565), .CLK(clk), .Q(n4461), .QN(n114) );
  DFFX1_HVT \keys_reg[0][31]  ( .D(n3564), .CLK(clk), .Q(n4462), .QN(n115) );
  DFFX1_HVT \keys_reg[0][30]  ( .D(n3563), .CLK(clk), .Q(n4463), .QN(n116) );
  DFFX1_HVT \keys_reg[0][29]  ( .D(n3562), .CLK(clk), .Q(n4464), .QN(n117) );
  DFFX1_HVT \keys_reg[0][28]  ( .D(n3561), .CLK(clk), .Q(n4465), .QN(n118) );
  DFFX1_HVT \keys_reg[0][27]  ( .D(n3560), .CLK(clk), .Q(n4466), .QN(n119) );
  DFFX1_HVT \keys_reg[0][26]  ( .D(n3559), .CLK(clk), .Q(n4467), .QN(n120) );
  DFFX1_HVT \keys_reg[0][25]  ( .D(n3558), .CLK(clk), .Q(n4468), .QN(n121) );
  DFFX1_HVT \keys_reg[0][24]  ( .D(n3557), .CLK(clk), .Q(n4469), .QN(n122) );
  DFFX1_HVT \keys_reg[0][23]  ( .D(n3556), .CLK(clk), .Q(n4470), .QN(n123) );
  DFFX1_HVT \keys_reg[0][22]  ( .D(n3555), .CLK(clk), .Q(n4471), .QN(n124) );
  DFFX1_HVT \keys_reg[0][21]  ( .D(n3554), .CLK(clk), .Q(n4472), .QN(n125) );
  DFFX1_HVT \keys_reg[0][20]  ( .D(n3553), .CLK(clk), .Q(n4473), .QN(n126) );
  DFFX1_HVT \keys_reg[0][19]  ( .D(n3552), .CLK(clk), .Q(n4474), .QN(n127) );
  DFFX1_HVT \keys_reg[0][18]  ( .D(n3551), .CLK(clk), .Q(n4475), .QN(n128) );
  DFFX1_HVT \keys_reg[0][17]  ( .D(n3550), .CLK(clk), .Q(n4476), .QN(n129) );
  DFFX1_HVT \keys_reg[0][16]  ( .D(n3549), .CLK(clk), .Q(n4477), .QN(n130) );
  DFFX1_HVT \keys_reg[0][15]  ( .D(n3548), .CLK(clk), .Q(n4478), .QN(n131) );
  DFFX1_HVT \keys_reg[0][14]  ( .D(n3547), .CLK(clk), .Q(n4479), .QN(n132) );
  DFFX1_HVT \keys_reg[0][13]  ( .D(n3546), .CLK(clk), .Q(n4480), .QN(n133) );
  DFFX1_HVT \keys_reg[0][12]  ( .D(n3545), .CLK(clk), .Q(n4481), .QN(n134) );
  DFFX1_HVT \keys_reg[0][11]  ( .D(n3544), .CLK(clk), .Q(n4482), .QN(n135) );
  DFFX1_HVT \keys_reg[0][10]  ( .D(n3543), .CLK(clk), .Q(n4483), .QN(n136) );
  DFFX1_HVT \keys_reg[0][9]  ( .D(n3542), .CLK(clk), .Q(n4484), .QN(n137) );
  DFFX1_HVT \keys_reg[0][8]  ( .D(n3541), .CLK(clk), .Q(n4485), .QN(n138) );
  DFFX1_HVT \keys_reg[0][7]  ( .D(n3540), .CLK(clk), .Q(n4486), .QN(n139) );
  DFFX1_HVT \keys_reg[0][6]  ( .D(n3539), .CLK(clk), .Q(n4487), .QN(n140) );
  DFFX1_HVT \keys_reg[0][5]  ( .D(n3538), .CLK(clk), .Q(n4488), .QN(n141) );
  DFFX1_HVT \keys_reg[0][4]  ( .D(n3537), .CLK(clk), .Q(n4489), .QN(n142) );
  DFFX1_HVT \keys_reg[0][3]  ( .D(n3536), .CLK(clk), .Q(n4490), .QN(n143) );
  DFFX1_HVT \keys_reg[0][2]  ( .D(n3535), .CLK(clk), .Q(n4491), .QN(n144) );
  DFFX1_HVT \keys_reg[0][1]  ( .D(n3534), .CLK(clk), .Q(n4492), .QN(n145) );
  DFFX1_HVT \keys_reg[0][0]  ( .D(n3533), .CLK(clk), .Q(n4493), .QN(n146) );
  DFFX1_HVT \keys_reg[1][127]  ( .D(n3532), .CLK(clk), .Q(n5), .QN(n147) );
  DFFX1_HVT \keys_reg[1][126]  ( .D(n3531), .CLK(clk), .Q(n6), .QN(n148) );
  DFFX1_HVT \keys_reg[1][125]  ( .D(n3530), .CLK(clk), .Q(n7), .QN(n149) );
  DFFX1_HVT \keys_reg[1][124]  ( .D(n3529), .CLK(clk), .Q(n8), .QN(n150) );
  DFFX1_HVT \keys_reg[1][123]  ( .D(n3528), .CLK(clk), .Q(n9), .QN(n151) );
  DFFX1_HVT \keys_reg[1][122]  ( .D(n3527), .CLK(clk), .Q(n10), .QN(n152) );
  DFFX1_HVT \keys_reg[1][121]  ( .D(n3526), .CLK(clk), .Q(n11), .QN(n153) );
  DFFX1_HVT \keys_reg[1][120]  ( .D(n3525), .CLK(clk), .Q(n12), .QN(n154) );
  DFFX1_HVT \keys_reg[1][119]  ( .D(n3524), .CLK(clk), .Q(n13), .QN(n155) );
  DFFX1_HVT \keys_reg[1][118]  ( .D(n3523), .CLK(clk), .Q(n14), .QN(n156) );
  DFFX1_HVT \keys_reg[1][117]  ( .D(n3522), .CLK(clk), .Q(n15), .QN(n157) );
  DFFX1_HVT \keys_reg[1][116]  ( .D(n3521), .CLK(clk), .Q(n16), .QN(n158) );
  DFFX1_HVT \keys_reg[1][115]  ( .D(n3520), .CLK(clk), .Q(n17), .QN(n159) );
  DFFX1_HVT \keys_reg[1][114]  ( .D(n3519), .CLK(clk), .Q(n18), .QN(n160) );
  DFFX1_HVT \keys_reg[1][113]  ( .D(n3518), .CLK(clk), .Q(n1427), .QN(n161) );
  DFFX1_HVT \keys_reg[1][112]  ( .D(n3517), .CLK(clk), .Q(n1428), .QN(n162) );
  DFFX1_HVT \keys_reg[1][111]  ( .D(n3516), .CLK(clk), .Q(n1429), .QN(n163) );
  DFFX1_HVT \keys_reg[1][110]  ( .D(n3515), .CLK(clk), .Q(n1430), .QN(n164) );
  DFFX1_HVT \keys_reg[1][109]  ( .D(n3514), .CLK(clk), .Q(n1431), .QN(n165) );
  DFFX1_HVT \keys_reg[1][108]  ( .D(n3513), .CLK(clk), .Q(n1432), .QN(n166) );
  DFFX1_HVT \keys_reg[1][107]  ( .D(n3512), .CLK(clk), .Q(n1433), .QN(n167) );
  DFFX1_HVT \keys_reg[1][106]  ( .D(n3511), .CLK(clk), .Q(n1434), .QN(n168) );
  DFFX1_HVT \keys_reg[1][105]  ( .D(n3510), .CLK(clk), .Q(n1435), .QN(n169) );
  DFFX1_HVT \keys_reg[1][104]  ( .D(n3509), .CLK(clk), .Q(n1436), .QN(n170) );
  DFFX1_HVT \keys_reg[1][103]  ( .D(n3508), .CLK(clk), .Q(n1437), .QN(n171) );
  DFFX1_HVT \keys_reg[1][102]  ( .D(n3507), .CLK(clk), .Q(n1438), .QN(n172) );
  DFFX1_HVT \keys_reg[1][101]  ( .D(n3506), .CLK(clk), .Q(n1439), .QN(n173) );
  DFFX1_HVT \keys_reg[1][100]  ( .D(n3505), .CLK(clk), .Q(n1440), .QN(n174) );
  DFFX1_HVT \keys_reg[1][99]  ( .D(n3504), .CLK(clk), .Q(n1441), .QN(n175) );
  DFFX1_HVT \keys_reg[1][98]  ( .D(n3503), .CLK(clk), .Q(n1442), .QN(n176) );
  DFFX1_HVT \keys_reg[1][97]  ( .D(n3502), .CLK(clk), .Q(n1443), .QN(n177) );
  DFFX1_HVT \keys_reg[1][96]  ( .D(n3501), .CLK(clk), .Q(n1444), .QN(n178) );
  DFFX1_HVT \keys_reg[1][95]  ( .D(n3500), .CLK(clk), .Q(n1445), .QN(n179) );
  DFFX1_HVT \keys_reg[1][94]  ( .D(n3499), .CLK(clk), .Q(n1446), .QN(n180) );
  DFFX1_HVT \keys_reg[1][93]  ( .D(n3498), .CLK(clk), .Q(n1447), .QN(n181) );
  DFFX1_HVT \keys_reg[1][92]  ( .D(n3497), .CLK(clk), .Q(n1448), .QN(n182) );
  DFFX1_HVT \keys_reg[1][91]  ( .D(n3496), .CLK(clk), .Q(n1449), .QN(n183) );
  DFFX1_HVT \keys_reg[1][90]  ( .D(n3495), .CLK(clk), .Q(n1450), .QN(n184) );
  DFFX1_HVT \keys_reg[1][89]  ( .D(n3494), .CLK(clk), .Q(n1451), .QN(n185) );
  DFFX1_HVT \keys_reg[1][88]  ( .D(n3493), .CLK(clk), .Q(n1452), .QN(n186) );
  DFFX1_HVT \keys_reg[1][87]  ( .D(n3492), .CLK(clk), .Q(n1453), .QN(n187) );
  DFFX1_HVT \keys_reg[1][86]  ( .D(n3491), .CLK(clk), .Q(n1454), .QN(n188) );
  DFFX1_HVT \keys_reg[1][85]  ( .D(n3490), .CLK(clk), .Q(n1455), .QN(n189) );
  DFFX1_HVT \keys_reg[1][84]  ( .D(n3489), .CLK(clk), .Q(n1456), .QN(n190) );
  DFFX1_HVT \keys_reg[1][83]  ( .D(n3488), .CLK(clk), .Q(n1457), .QN(n191) );
  DFFX1_HVT \keys_reg[1][82]  ( .D(n3487), .CLK(clk), .Q(n1458), .QN(n192) );
  DFFX1_HVT \keys_reg[1][81]  ( .D(n3486), .CLK(clk), .Q(n1459), .QN(n193) );
  DFFX1_HVT \keys_reg[1][80]  ( .D(n3485), .CLK(clk), .Q(n1460), .QN(n194) );
  DFFX1_HVT \keys_reg[1][79]  ( .D(n3484), .CLK(clk), .Q(n1461), .QN(n195) );
  DFFX1_HVT \keys_reg[1][78]  ( .D(n3483), .CLK(clk), .Q(n1462), .QN(n196) );
  DFFX1_HVT \keys_reg[1][77]  ( .D(n3482), .CLK(clk), .Q(n1463), .QN(n197) );
  DFFX1_HVT \keys_reg[1][76]  ( .D(n3481), .CLK(clk), .Q(n1464), .QN(n198) );
  DFFX1_HVT \keys_reg[1][75]  ( .D(n3480), .CLK(clk), .Q(n1465), .QN(n199) );
  DFFX1_HVT \keys_reg[1][74]  ( .D(n3479), .CLK(clk), .Q(n1466), .QN(n200) );
  DFFX1_HVT \keys_reg[1][73]  ( .D(n3478), .CLK(clk), .Q(n1467), .QN(n201) );
  DFFX1_HVT \keys_reg[1][72]  ( .D(n3477), .CLK(clk), .Q(n1468), .QN(n202) );
  DFFX1_HVT \keys_reg[1][71]  ( .D(n3476), .CLK(clk), .Q(n1469), .QN(n203) );
  DFFX1_HVT \keys_reg[1][70]  ( .D(n3475), .CLK(clk), .Q(n1470), .QN(n204) );
  DFFX1_HVT \keys_reg[1][69]  ( .D(n3474), .CLK(clk), .Q(n1471), .QN(n205) );
  DFFX1_HVT \keys_reg[1][68]  ( .D(n3473), .CLK(clk), .Q(n1472), .QN(n206) );
  DFFX1_HVT \keys_reg[1][67]  ( .D(n3472), .CLK(clk), .Q(n1473), .QN(n207) );
  DFFX1_HVT \keys_reg[1][66]  ( .D(n3471), .CLK(clk), .Q(n1474), .QN(n208) );
  DFFX1_HVT \keys_reg[1][65]  ( .D(n3470), .CLK(clk), .Q(n1475), .QN(n209) );
  DFFX1_HVT \keys_reg[1][64]  ( .D(n3469), .CLK(clk), .Q(n1476), .QN(n210) );
  DFFX1_HVT \keys_reg[1][63]  ( .D(n3468), .CLK(clk), .Q(n1477), .QN(n211) );
  DFFX1_HVT \keys_reg[1][62]  ( .D(n3467), .CLK(clk), .Q(n1478), .QN(n212) );
  DFFX1_HVT \keys_reg[1][61]  ( .D(n3466), .CLK(clk), .Q(n1479), .QN(n213) );
  DFFX1_HVT \keys_reg[1][60]  ( .D(n3465), .CLK(clk), .Q(n1480), .QN(n214) );
  DFFX1_HVT \keys_reg[1][59]  ( .D(n3464), .CLK(clk), .Q(n1481), .QN(n215) );
  DFFX1_HVT \keys_reg[1][58]  ( .D(n3463), .CLK(clk), .Q(n1482), .QN(n216) );
  DFFX1_HVT \keys_reg[1][57]  ( .D(n3462), .CLK(clk), .Q(n1483), .QN(n217) );
  DFFX1_HVT \keys_reg[1][56]  ( .D(n3461), .CLK(clk), .Q(n1484), .QN(n218) );
  DFFX1_HVT \keys_reg[1][55]  ( .D(n3460), .CLK(clk), .Q(n1485), .QN(n219) );
  DFFX1_HVT \keys_reg[1][54]  ( .D(n3459), .CLK(clk), .Q(n1486), .QN(n220) );
  DFFX1_HVT \keys_reg[1][53]  ( .D(n3458), .CLK(clk), .Q(n1487), .QN(n221) );
  DFFX1_HVT \keys_reg[1][52]  ( .D(n3457), .CLK(clk), .Q(n1488), .QN(n222) );
  DFFX1_HVT \keys_reg[1][51]  ( .D(n3456), .CLK(clk), .Q(n1489), .QN(n223) );
  DFFX1_HVT \keys_reg[1][50]  ( .D(n3455), .CLK(clk), .Q(n1490), .QN(n224) );
  DFFX1_HVT \keys_reg[1][49]  ( .D(n3454), .CLK(clk), .Q(n1491), .QN(n225) );
  DFFX1_HVT \keys_reg[1][48]  ( .D(n3453), .CLK(clk), .Q(n1492), .QN(n226) );
  DFFX1_HVT \keys_reg[1][47]  ( .D(n3452), .CLK(clk), .Q(n1493), .QN(n227) );
  DFFX1_HVT \keys_reg[1][46]  ( .D(n3451), .CLK(clk), .Q(n1494), .QN(n228) );
  DFFX1_HVT \keys_reg[1][45]  ( .D(n3450), .CLK(clk), .Q(n1495), .QN(n229) );
  DFFX1_HVT \keys_reg[1][44]  ( .D(n3449), .CLK(clk), .Q(n1496), .QN(n230) );
  DFFX1_HVT \keys_reg[1][43]  ( .D(n3448), .CLK(clk), .Q(n1497), .QN(n231) );
  DFFX1_HVT \keys_reg[1][42]  ( .D(n3447), .CLK(clk), .Q(n1498), .QN(n232) );
  DFFX1_HVT \keys_reg[1][41]  ( .D(n3446), .CLK(clk), .Q(n1499), .QN(n233) );
  DFFX1_HVT \keys_reg[1][40]  ( .D(n3445), .CLK(clk), .Q(n1500), .QN(n234) );
  DFFX1_HVT \keys_reg[1][39]  ( .D(n3444), .CLK(clk), .Q(n1501), .QN(n235) );
  DFFX1_HVT \keys_reg[1][38]  ( .D(n3443), .CLK(clk), .Q(n1502), .QN(n236) );
  DFFX1_HVT \keys_reg[1][37]  ( .D(n3442), .CLK(clk), .Q(n1503), .QN(n237) );
  DFFX1_HVT \keys_reg[1][36]  ( .D(n3441), .CLK(clk), .Q(n1504), .QN(n238) );
  DFFX1_HVT \keys_reg[1][35]  ( .D(n3440), .CLK(clk), .Q(n1505), .QN(n239) );
  DFFX1_HVT \keys_reg[1][34]  ( .D(n3439), .CLK(clk), .Q(n1506), .QN(n240) );
  DFFX1_HVT \keys_reg[1][33]  ( .D(n3438), .CLK(clk), .Q(n1507), .QN(n241) );
  DFFX1_HVT \keys_reg[1][32]  ( .D(n3437), .CLK(clk), .Q(n1508), .QN(n242) );
  DFFX1_HVT \keys_reg[1][31]  ( .D(n3436), .CLK(clk), .Q(n1509), .QN(n243) );
  DFFX1_HVT \keys_reg[1][30]  ( .D(n3435), .CLK(clk), .Q(n1510), .QN(n244) );
  DFFX1_HVT \keys_reg[1][29]  ( .D(n3434), .CLK(clk), .Q(n1511), .QN(n245) );
  DFFX1_HVT \keys_reg[1][28]  ( .D(n3433), .CLK(clk), .Q(n1512), .QN(n246) );
  DFFX1_HVT \keys_reg[1][27]  ( .D(n3432), .CLK(clk), .Q(n1513), .QN(n247) );
  DFFX1_HVT \keys_reg[1][26]  ( .D(n3431), .CLK(clk), .Q(n1514), .QN(n248) );
  DFFX1_HVT \keys_reg[1][25]  ( .D(n3430), .CLK(clk), .Q(n1515), .QN(n249) );
  DFFX1_HVT \keys_reg[1][24]  ( .D(n3429), .CLK(clk), .Q(n1516), .QN(n250) );
  DFFX1_HVT \keys_reg[1][23]  ( .D(n3428), .CLK(clk), .Q(n1517), .QN(n251) );
  DFFX1_HVT \keys_reg[1][22]  ( .D(n3427), .CLK(clk), .Q(n1518), .QN(n252) );
  DFFX1_HVT \keys_reg[1][21]  ( .D(n3426), .CLK(clk), .Q(n1519), .QN(n253) );
  DFFX1_HVT \keys_reg[1][20]  ( .D(n3425), .CLK(clk), .Q(n1520), .QN(n254) );
  DFFX1_HVT \keys_reg[1][19]  ( .D(n3424), .CLK(clk), .Q(n1521), .QN(n255) );
  DFFX1_HVT \keys_reg[1][18]  ( .D(n3423), .CLK(clk), .Q(n1522), .QN(n256) );
  DFFX1_HVT \keys_reg[1][17]  ( .D(n3422), .CLK(clk), .Q(n1523), .QN(n257) );
  DFFX1_HVT \keys_reg[1][16]  ( .D(n3421), .CLK(clk), .Q(n1524), .QN(n258) );
  DFFX1_HVT \keys_reg[1][15]  ( .D(n3420), .CLK(clk), .Q(n1525), .QN(n259) );
  DFFX1_HVT \keys_reg[1][14]  ( .D(n3419), .CLK(clk), .Q(n1526), .QN(n260) );
  DFFX1_HVT \keys_reg[1][13]  ( .D(n3418), .CLK(clk), .Q(n1527), .QN(n261) );
  DFFX1_HVT \keys_reg[1][12]  ( .D(n3417), .CLK(clk), .Q(n1528), .QN(n262) );
  DFFX1_HVT \keys_reg[1][11]  ( .D(n3416), .CLK(clk), .Q(n1529), .QN(n263) );
  DFFX1_HVT \keys_reg[1][10]  ( .D(n3415), .CLK(clk), .Q(n1530), .QN(n264) );
  DFFX1_HVT \keys_reg[1][9]  ( .D(n3414), .CLK(clk), .Q(n1531), .QN(n265) );
  DFFX1_HVT \keys_reg[1][8]  ( .D(n3413), .CLK(clk), .Q(n1532), .QN(n266) );
  DFFX1_HVT \keys_reg[1][7]  ( .D(n3412), .CLK(clk), .Q(n1533), .QN(n267) );
  DFFX1_HVT \keys_reg[1][6]  ( .D(n3411), .CLK(clk), .Q(n1534), .QN(n268) );
  DFFX1_HVT \keys_reg[1][5]  ( .D(n3410), .CLK(clk), .Q(n1535), .QN(n269) );
  DFFX1_HVT \keys_reg[1][4]  ( .D(n3409), .CLK(clk), .Q(n1536), .QN(n270) );
  DFFX1_HVT \keys_reg[1][3]  ( .D(n3408), .CLK(clk), .Q(n1537), .QN(n271) );
  DFFX1_HVT \keys_reg[1][2]  ( .D(n3407), .CLK(clk), .Q(n1538), .QN(n272) );
  DFFX1_HVT \keys_reg[1][1]  ( .D(n3406), .CLK(clk), .Q(n1539), .QN(n273) );
  DFFX1_HVT \keys_reg[1][0]  ( .D(n3405), .CLK(clk), .Q(n1540), .QN(n274) );
  DFFX1_HVT \keys_reg[2][127]  ( .D(n3404), .CLK(clk), .Q(n3982), .QN(n275) );
  DFFX1_HVT \keys_reg[2][126]  ( .D(n3403), .CLK(clk), .Q(n3983), .QN(n276) );
  DFFX1_HVT \keys_reg[2][125]  ( .D(n3402), .CLK(clk), .Q(n3984), .QN(n277) );
  DFFX1_HVT \keys_reg[2][124]  ( .D(n3401), .CLK(clk), .Q(n3985), .QN(n278) );
  DFFX1_HVT \keys_reg[2][123]  ( .D(n3400), .CLK(clk), .Q(n3986), .QN(n279) );
  DFFX1_HVT \keys_reg[2][122]  ( .D(n3399), .CLK(clk), .Q(n3987), .QN(n280) );
  DFFX1_HVT \keys_reg[2][121]  ( .D(n3398), .CLK(clk), .Q(n3988), .QN(n281) );
  DFFX1_HVT \keys_reg[2][120]  ( .D(n3397), .CLK(clk), .Q(n3989), .QN(n282) );
  DFFX1_HVT \keys_reg[2][119]  ( .D(n3396), .CLK(clk), .Q(n3990), .QN(n283) );
  DFFX1_HVT \keys_reg[2][118]  ( .D(n3395), .CLK(clk), .Q(n3991), .QN(n284) );
  DFFX1_HVT \keys_reg[2][117]  ( .D(n3394), .CLK(clk), .Q(n3992), .QN(n285) );
  DFFX1_HVT \keys_reg[2][116]  ( .D(n3393), .CLK(clk), .Q(n3993), .QN(n286) );
  DFFX1_HVT \keys_reg[2][115]  ( .D(n3392), .CLK(clk), .Q(n3994), .QN(n287) );
  DFFX1_HVT \keys_reg[2][114]  ( .D(n3391), .CLK(clk), .Q(n3995), .QN(n288) );
  DFFX1_HVT \keys_reg[2][113]  ( .D(n3390), .CLK(clk), .Q(n3996), .QN(n289) );
  DFFX1_HVT \keys_reg[2][112]  ( .D(n3389), .CLK(clk), .Q(n3997), .QN(n290) );
  DFFX1_HVT \keys_reg[2][111]  ( .D(n3388), .CLK(clk), .Q(n3998), .QN(n291) );
  DFFX1_HVT \keys_reg[2][110]  ( .D(n3387), .CLK(clk), .Q(n3999), .QN(n292) );
  DFFX1_HVT \keys_reg[2][109]  ( .D(n3386), .CLK(clk), .Q(n4000), .QN(n293) );
  DFFX1_HVT \keys_reg[2][108]  ( .D(n3385), .CLK(clk), .Q(n4001), .QN(n294) );
  DFFX1_HVT \keys_reg[2][107]  ( .D(n3384), .CLK(clk), .Q(n4002), .QN(n295) );
  DFFX1_HVT \keys_reg[2][106]  ( .D(n3383), .CLK(clk), .Q(n4003), .QN(n296) );
  DFFX1_HVT \keys_reg[2][105]  ( .D(n3382), .CLK(clk), .Q(n4004), .QN(n297) );
  DFFX1_HVT \keys_reg[2][104]  ( .D(n3381), .CLK(clk), .Q(n4005), .QN(n298) );
  DFFX1_HVT \keys_reg[2][103]  ( .D(n3380), .CLK(clk), .Q(n4006), .QN(n299) );
  DFFX1_HVT \keys_reg[2][102]  ( .D(n3379), .CLK(clk), .Q(n4007), .QN(n300) );
  DFFX1_HVT \keys_reg[2][101]  ( .D(n3378), .CLK(clk), .Q(n4008), .QN(n301) );
  DFFX1_HVT \keys_reg[2][100]  ( .D(n3377), .CLK(clk), .Q(n4009), .QN(n302) );
  DFFX1_HVT \keys_reg[2][99]  ( .D(n3376), .CLK(clk), .Q(n4010), .QN(n303) );
  DFFX1_HVT \keys_reg[2][98]  ( .D(n3375), .CLK(clk), .Q(n4011), .QN(n304) );
  DFFX1_HVT \keys_reg[2][97]  ( .D(n3374), .CLK(clk), .Q(n4012), .QN(n305) );
  DFFX1_HVT \keys_reg[2][96]  ( .D(n3373), .CLK(clk), .Q(n4013), .QN(n306) );
  DFFX1_HVT \keys_reg[2][95]  ( .D(n3372), .CLK(clk), .Q(n4014), .QN(n307) );
  DFFX1_HVT \keys_reg[2][94]  ( .D(n3371), .CLK(clk), .Q(n4015), .QN(n308) );
  DFFX1_HVT \keys_reg[2][93]  ( .D(n3370), .CLK(clk), .Q(n4016), .QN(n309) );
  DFFX1_HVT \keys_reg[2][92]  ( .D(n3369), .CLK(clk), .Q(n4017), .QN(n310) );
  DFFX1_HVT \keys_reg[2][91]  ( .D(n3368), .CLK(clk), .Q(n4018), .QN(n311) );
  DFFX1_HVT \keys_reg[2][90]  ( .D(n3367), .CLK(clk), .Q(n4019), .QN(n312) );
  DFFX1_HVT \keys_reg[2][89]  ( .D(n3366), .CLK(clk), .Q(n4020), .QN(n313) );
  DFFX1_HVT \keys_reg[2][88]  ( .D(n3365), .CLK(clk), .Q(n4021), .QN(n314) );
  DFFX1_HVT \keys_reg[2][87]  ( .D(n3364), .CLK(clk), .Q(n4022), .QN(n315) );
  DFFX1_HVT \keys_reg[2][86]  ( .D(n3363), .CLK(clk), .Q(n4023), .QN(n316) );
  DFFX1_HVT \keys_reg[2][85]  ( .D(n3362), .CLK(clk), .Q(n4024), .QN(n317) );
  DFFX1_HVT \keys_reg[2][84]  ( .D(n3361), .CLK(clk), .Q(n4025), .QN(n318) );
  DFFX1_HVT \keys_reg[2][83]  ( .D(n3360), .CLK(clk), .Q(n4026), .QN(n319) );
  DFFX1_HVT \keys_reg[2][82]  ( .D(n3359), .CLK(clk), .Q(n4027), .QN(n320) );
  DFFX1_HVT \keys_reg[2][81]  ( .D(n3358), .CLK(clk), .Q(n4028), .QN(n321) );
  DFFX1_HVT \keys_reg[2][80]  ( .D(n3357), .CLK(clk), .Q(n4029), .QN(n322) );
  DFFX1_HVT \keys_reg[2][79]  ( .D(n3356), .CLK(clk), .Q(n4030), .QN(n323) );
  DFFX1_HVT \keys_reg[2][78]  ( .D(n3355), .CLK(clk), .Q(n4031), .QN(n324) );
  DFFX1_HVT \keys_reg[2][77]  ( .D(n3354), .CLK(clk), .Q(n4032), .QN(n325) );
  DFFX1_HVT \keys_reg[2][76]  ( .D(n3353), .CLK(clk), .Q(n4033), .QN(n326) );
  DFFX1_HVT \keys_reg[2][75]  ( .D(n3352), .CLK(clk), .Q(n4034), .QN(n327) );
  DFFX1_HVT \keys_reg[2][74]  ( .D(n3351), .CLK(clk), .Q(n4035), .QN(n328) );
  DFFX1_HVT \keys_reg[2][73]  ( .D(n3350), .CLK(clk), .Q(n4036), .QN(n329) );
  DFFX1_HVT \keys_reg[2][72]  ( .D(n3349), .CLK(clk), .Q(n4037), .QN(n330) );
  DFFX1_HVT \keys_reg[2][71]  ( .D(n3348), .CLK(clk), .Q(n4038), .QN(n331) );
  DFFX1_HVT \keys_reg[2][70]  ( .D(n3347), .CLK(clk), .Q(n4039), .QN(n332) );
  DFFX1_HVT \keys_reg[2][69]  ( .D(n3346), .CLK(clk), .Q(n4040), .QN(n333) );
  DFFX1_HVT \keys_reg[2][68]  ( .D(n3345), .CLK(clk), .Q(n4041), .QN(n334) );
  DFFX1_HVT \keys_reg[2][67]  ( .D(n3344), .CLK(clk), .Q(n4042), .QN(n335) );
  DFFX1_HVT \keys_reg[2][66]  ( .D(n3343), .CLK(clk), .Q(n4043), .QN(n336) );
  DFFX1_HVT \keys_reg[2][65]  ( .D(n3342), .CLK(clk), .Q(n4044), .QN(n337) );
  DFFX1_HVT \keys_reg[2][64]  ( .D(n3341), .CLK(clk), .Q(n4045), .QN(n338) );
  DFFX1_HVT \keys_reg[2][63]  ( .D(n3340), .CLK(clk), .Q(n4046), .QN(n339) );
  DFFX1_HVT \keys_reg[2][62]  ( .D(n3339), .CLK(clk), .Q(n4047), .QN(n340) );
  DFFX1_HVT \keys_reg[2][61]  ( .D(n3338), .CLK(clk), .Q(n4048), .QN(n341) );
  DFFX1_HVT \keys_reg[2][60]  ( .D(n3337), .CLK(clk), .Q(n4049), .QN(n342) );
  DFFX1_HVT \keys_reg[2][59]  ( .D(n3336), .CLK(clk), .Q(n4050), .QN(n343) );
  DFFX1_HVT \keys_reg[2][58]  ( .D(n3335), .CLK(clk), .Q(n4051), .QN(n344) );
  DFFX1_HVT \keys_reg[2][57]  ( .D(n3334), .CLK(clk), .Q(n4052), .QN(n345) );
  DFFX1_HVT \keys_reg[2][56]  ( .D(n3333), .CLK(clk), .Q(n4053), .QN(n346) );
  DFFX1_HVT \keys_reg[2][55]  ( .D(n3332), .CLK(clk), .Q(n4054), .QN(n347) );
  DFFX1_HVT \keys_reg[2][54]  ( .D(n3331), .CLK(clk), .Q(n4055), .QN(n348) );
  DFFX1_HVT \keys_reg[2][53]  ( .D(n3330), .CLK(clk), .Q(n4056), .QN(n349) );
  DFFX1_HVT \keys_reg[2][52]  ( .D(n3329), .CLK(clk), .Q(n4057), .QN(n350) );
  DFFX1_HVT \keys_reg[2][51]  ( .D(n3328), .CLK(clk), .Q(n4058), .QN(n351) );
  DFFX1_HVT \keys_reg[2][50]  ( .D(n3327), .CLK(clk), .Q(n4059), .QN(n352) );
  DFFX1_HVT \keys_reg[2][49]  ( .D(n3326), .CLK(clk), .Q(n4060), .QN(n353) );
  DFFX1_HVT \keys_reg[2][48]  ( .D(n3325), .CLK(clk), .Q(n4061), .QN(n354) );
  DFFX1_HVT \keys_reg[2][47]  ( .D(n3324), .CLK(clk), .Q(n4062), .QN(n355) );
  DFFX1_HVT \keys_reg[2][46]  ( .D(n3323), .CLK(clk), .Q(n4063), .QN(n356) );
  DFFX1_HVT \keys_reg[2][45]  ( .D(n3322), .CLK(clk), .Q(n4064), .QN(n357) );
  DFFX1_HVT \keys_reg[2][44]  ( .D(n3321), .CLK(clk), .Q(n4065), .QN(n358) );
  DFFX1_HVT \keys_reg[2][43]  ( .D(n3320), .CLK(clk), .Q(n4066), .QN(n359) );
  DFFX1_HVT \keys_reg[2][42]  ( .D(n3319), .CLK(clk), .Q(n4067), .QN(n360) );
  DFFX1_HVT \keys_reg[2][41]  ( .D(n3318), .CLK(clk), .Q(n4068), .QN(n361) );
  DFFX1_HVT \keys_reg[2][40]  ( .D(n3317), .CLK(clk), .Q(n4069), .QN(n362) );
  DFFX1_HVT \keys_reg[2][39]  ( .D(n3316), .CLK(clk), .Q(n4070), .QN(n363) );
  DFFX1_HVT \keys_reg[2][38]  ( .D(n3315), .CLK(clk), .Q(n4071), .QN(n364) );
  DFFX1_HVT \keys_reg[2][37]  ( .D(n3314), .CLK(clk), .Q(n4072), .QN(n365) );
  DFFX1_HVT \keys_reg[2][36]  ( .D(n3313), .CLK(clk), .Q(n4073), .QN(n366) );
  DFFX1_HVT \keys_reg[2][35]  ( .D(n3312), .CLK(clk), .Q(n4074), .QN(n367) );
  DFFX1_HVT \keys_reg[2][34]  ( .D(n3311), .CLK(clk), .Q(n4075), .QN(n368) );
  DFFX1_HVT \keys_reg[2][33]  ( .D(n3310), .CLK(clk), .Q(n4076), .QN(n369) );
  DFFX1_HVT \keys_reg[2][32]  ( .D(n3309), .CLK(clk), .Q(n4077), .QN(n370) );
  DFFX1_HVT \keys_reg[2][31]  ( .D(n3308), .CLK(clk), .Q(n4078), .QN(n371) );
  DFFX1_HVT \keys_reg[2][30]  ( .D(n3307), .CLK(clk), .Q(n4079), .QN(n372) );
  DFFX1_HVT \keys_reg[2][29]  ( .D(n3306), .CLK(clk), .Q(n4080), .QN(n373) );
  DFFX1_HVT \keys_reg[2][28]  ( .D(n3305), .CLK(clk), .Q(n4081), .QN(n374) );
  DFFX1_HVT \keys_reg[2][27]  ( .D(n3304), .CLK(clk), .Q(n4082), .QN(n375) );
  DFFX1_HVT \keys_reg[2][26]  ( .D(n3303), .CLK(clk), .Q(n4083), .QN(n376) );
  DFFX1_HVT \keys_reg[2][25]  ( .D(n3302), .CLK(clk), .Q(n4084), .QN(n377) );
  DFFX1_HVT \keys_reg[2][24]  ( .D(n3301), .CLK(clk), .Q(n4085), .QN(n378) );
  DFFX1_HVT \keys_reg[2][23]  ( .D(n3300), .CLK(clk), .Q(n4086), .QN(n379) );
  DFFX1_HVT \keys_reg[2][22]  ( .D(n3299), .CLK(clk), .Q(n4087), .QN(n380) );
  DFFX1_HVT \keys_reg[2][21]  ( .D(n3298), .CLK(clk), .Q(n4088), .QN(n381) );
  DFFX1_HVT \keys_reg[2][20]  ( .D(n3297), .CLK(clk), .Q(n4089), .QN(n382) );
  DFFX1_HVT \keys_reg[2][19]  ( .D(n3296), .CLK(clk), .Q(n4090), .QN(n383) );
  DFFX1_HVT \keys_reg[2][18]  ( .D(n3295), .CLK(clk), .Q(n4091), .QN(n384) );
  DFFX1_HVT \keys_reg[2][17]  ( .D(n3294), .CLK(clk), .Q(n4092), .QN(n385) );
  DFFX1_HVT \keys_reg[2][16]  ( .D(n3293), .CLK(clk), .Q(n4093), .QN(n386) );
  DFFX1_HVT \keys_reg[2][15]  ( .D(n3292), .CLK(clk), .Q(n4094), .QN(n387) );
  DFFX1_HVT \keys_reg[2][14]  ( .D(n3291), .CLK(clk), .Q(n4095), .QN(n388) );
  DFFX1_HVT \keys_reg[2][13]  ( .D(n3290), .CLK(clk), .Q(n4096), .QN(n389) );
  DFFX1_HVT \keys_reg[2][12]  ( .D(n3289), .CLK(clk), .Q(n4097), .QN(n390) );
  DFFX1_HVT \keys_reg[2][11]  ( .D(n3288), .CLK(clk), .Q(n4098), .QN(n391) );
  DFFX1_HVT \keys_reg[2][10]  ( .D(n3287), .CLK(clk), .Q(n4099), .QN(n392) );
  DFFX1_HVT \keys_reg[2][9]  ( .D(n3286), .CLK(clk), .Q(n4100), .QN(n393) );
  DFFX1_HVT \keys_reg[2][8]  ( .D(n3285), .CLK(clk), .Q(n4101), .QN(n394) );
  DFFX1_HVT \keys_reg[2][7]  ( .D(n3284), .CLK(clk), .Q(n4102), .QN(n395) );
  DFFX1_HVT \keys_reg[2][6]  ( .D(n3283), .CLK(clk), .Q(n4103), .QN(n396) );
  DFFX1_HVT \keys_reg[2][5]  ( .D(n3282), .CLK(clk), .Q(n4104), .QN(n397) );
  DFFX1_HVT \keys_reg[2][4]  ( .D(n3281), .CLK(clk), .Q(n4105), .QN(n398) );
  DFFX1_HVT \keys_reg[2][3]  ( .D(n3280), .CLK(clk), .Q(n4106), .QN(n399) );
  DFFX1_HVT \keys_reg[2][2]  ( .D(n3279), .CLK(clk), .Q(n4107), .QN(n400) );
  DFFX1_HVT \keys_reg[2][1]  ( .D(n3278), .CLK(clk), .Q(n4108), .QN(n401) );
  DFFX1_HVT \keys_reg[2][0]  ( .D(n3277), .CLK(clk), .Q(n4109), .QN(n402) );
  DFFX1_HVT \keys_reg[3][127]  ( .D(n3276), .CLK(clk), .Q(n1669), .QN(n403) );
  DFFX1_HVT \keys_reg[3][126]  ( .D(n3275), .CLK(clk), .Q(n1670), .QN(n404) );
  DFFX1_HVT \keys_reg[3][125]  ( .D(n3274), .CLK(clk), .Q(n1671), .QN(n405) );
  DFFX1_HVT \keys_reg[3][124]  ( .D(n3273), .CLK(clk), .Q(n1672), .QN(n406) );
  DFFX1_HVT \keys_reg[3][123]  ( .D(n3272), .CLK(clk), .Q(n1673), .QN(n407) );
  DFFX1_HVT \keys_reg[3][122]  ( .D(n3271), .CLK(clk), .Q(n1674), .QN(n408) );
  DFFX1_HVT \keys_reg[3][121]  ( .D(n3270), .CLK(clk), .Q(n1675), .QN(n409) );
  DFFX1_HVT \keys_reg[3][120]  ( .D(n3269), .CLK(clk), .Q(n1676), .QN(n410) );
  DFFX1_HVT \keys_reg[3][119]  ( .D(n3268), .CLK(clk), .Q(n1677), .QN(n411) );
  DFFX1_HVT \keys_reg[3][118]  ( .D(n3267), .CLK(clk), .Q(n1678), .QN(n412) );
  DFFX1_HVT \keys_reg[3][117]  ( .D(n3266), .CLK(clk), .Q(n1679), .QN(n413) );
  DFFX1_HVT \keys_reg[3][116]  ( .D(n3265), .CLK(clk), .Q(n1680), .QN(n414) );
  DFFX1_HVT \keys_reg[3][115]  ( .D(n3264), .CLK(clk), .Q(n1681), .QN(n415) );
  DFFX1_HVT \keys_reg[3][114]  ( .D(n3263), .CLK(clk), .Q(n1682), .QN(n416) );
  DFFX1_HVT \keys_reg[3][113]  ( .D(n3262), .CLK(clk), .Q(n1683), .QN(n417) );
  DFFX1_HVT \keys_reg[3][112]  ( .D(n3261), .CLK(clk), .Q(n1684), .QN(n418) );
  DFFX1_HVT \keys_reg[3][111]  ( .D(n3260), .CLK(clk), .Q(n1685), .QN(n419) );
  DFFX1_HVT \keys_reg[3][110]  ( .D(n3259), .CLK(clk), .Q(n1686), .QN(n420) );
  DFFX1_HVT \keys_reg[3][109]  ( .D(n3258), .CLK(clk), .Q(n1687), .QN(n421) );
  DFFX1_HVT \keys_reg[3][108]  ( .D(n3257), .CLK(clk), .Q(n1688), .QN(n422) );
  DFFX1_HVT \keys_reg[3][107]  ( .D(n3256), .CLK(clk), .Q(n1689), .QN(n423) );
  DFFX1_HVT \keys_reg[3][106]  ( .D(n3255), .CLK(clk), .Q(n1690), .QN(n424) );
  DFFX1_HVT \keys_reg[3][105]  ( .D(n3254), .CLK(clk), .Q(n1691), .QN(n425) );
  DFFX1_HVT \keys_reg[3][104]  ( .D(n3253), .CLK(clk), .Q(n1692), .QN(n426) );
  DFFX1_HVT \keys_reg[3][103]  ( .D(n3252), .CLK(clk), .Q(n1693), .QN(n427) );
  DFFX1_HVT \keys_reg[3][102]  ( .D(n3251), .CLK(clk), .Q(n1694), .QN(n428) );
  DFFX1_HVT \keys_reg[3][101]  ( .D(n3250), .CLK(clk), .Q(n1695), .QN(n429) );
  DFFX1_HVT \keys_reg[3][100]  ( .D(n3249), .CLK(clk), .Q(n1696), .QN(n430) );
  DFFX1_HVT \keys_reg[3][99]  ( .D(n3248), .CLK(clk), .Q(n1697), .QN(n431) );
  DFFX1_HVT \keys_reg[3][98]  ( .D(n3247), .CLK(clk), .Q(n1698), .QN(n432) );
  DFFX1_HVT \keys_reg[3][97]  ( .D(n3246), .CLK(clk), .Q(n1699), .QN(n433) );
  DFFX1_HVT \keys_reg[3][96]  ( .D(n3245), .CLK(clk), .Q(n1700), .QN(n434) );
  DFFX1_HVT \keys_reg[3][95]  ( .D(n3244), .CLK(clk), .Q(n1701), .QN(n435) );
  DFFX1_HVT \keys_reg[3][94]  ( .D(n3243), .CLK(clk), .Q(n1702), .QN(n436) );
  DFFX1_HVT \keys_reg[3][93]  ( .D(n3242), .CLK(clk), .Q(n1703), .QN(n437) );
  DFFX1_HVT \keys_reg[3][92]  ( .D(n3241), .CLK(clk), .Q(n1704), .QN(n438) );
  DFFX1_HVT \keys_reg[3][91]  ( .D(n3240), .CLK(clk), .Q(n1705), .QN(n439) );
  DFFX1_HVT \keys_reg[3][90]  ( .D(n3239), .CLK(clk), .Q(n1706), .QN(n440) );
  DFFX1_HVT \keys_reg[3][89]  ( .D(n3238), .CLK(clk), .Q(n1707), .QN(n441) );
  DFFX1_HVT \keys_reg[3][88]  ( .D(n3237), .CLK(clk), .Q(n1708), .QN(n442) );
  DFFX1_HVT \keys_reg[3][87]  ( .D(n3236), .CLK(clk), .Q(n1709), .QN(n443) );
  DFFX1_HVT \keys_reg[3][86]  ( .D(n3235), .CLK(clk), .Q(n1710), .QN(n444) );
  DFFX1_HVT \keys_reg[3][85]  ( .D(n3234), .CLK(clk), .Q(n1711), .QN(n445) );
  DFFX1_HVT \keys_reg[3][84]  ( .D(n3233), .CLK(clk), .Q(n1712), .QN(n446) );
  DFFX1_HVT \keys_reg[3][83]  ( .D(n3232), .CLK(clk), .Q(n1713), .QN(n447) );
  DFFX1_HVT \keys_reg[3][82]  ( .D(n3231), .CLK(clk), .Q(n1714), .QN(n448) );
  DFFX1_HVT \keys_reg[3][81]  ( .D(n3230), .CLK(clk), .Q(n1715), .QN(n449) );
  DFFX1_HVT \keys_reg[3][80]  ( .D(n3229), .CLK(clk), .Q(n1716), .QN(n450) );
  DFFX1_HVT \keys_reg[3][79]  ( .D(n3228), .CLK(clk), .Q(n1717), .QN(n451) );
  DFFX1_HVT \keys_reg[3][78]  ( .D(n3227), .CLK(clk), .Q(n1718), .QN(n452) );
  DFFX1_HVT \keys_reg[3][77]  ( .D(n3226), .CLK(clk), .Q(n1719), .QN(n453) );
  DFFX1_HVT \keys_reg[3][76]  ( .D(n3225), .CLK(clk), .Q(n1720), .QN(n454) );
  DFFX1_HVT \keys_reg[3][75]  ( .D(n3224), .CLK(clk), .Q(n1721), .QN(n455) );
  DFFX1_HVT \keys_reg[3][74]  ( .D(n3223), .CLK(clk), .Q(n1722), .QN(n456) );
  DFFX1_HVT \keys_reg[3][73]  ( .D(n3222), .CLK(clk), .Q(n1723), .QN(n457) );
  DFFX1_HVT \keys_reg[3][72]  ( .D(n3221), .CLK(clk), .Q(n1724), .QN(n458) );
  DFFX1_HVT \keys_reg[3][71]  ( .D(n3220), .CLK(clk), .Q(n1725), .QN(n459) );
  DFFX1_HVT \keys_reg[3][70]  ( .D(n3219), .CLK(clk), .Q(n1726), .QN(n460) );
  DFFX1_HVT \keys_reg[3][69]  ( .D(n3218), .CLK(clk), .Q(n1727), .QN(n461) );
  DFFX1_HVT \keys_reg[3][68]  ( .D(n3217), .CLK(clk), .Q(n1728), .QN(n462) );
  DFFX1_HVT \keys_reg[3][67]  ( .D(n3216), .CLK(clk), .Q(n1729), .QN(n463) );
  DFFX1_HVT \keys_reg[3][66]  ( .D(n3215), .CLK(clk), .Q(n1730), .QN(n464) );
  DFFX1_HVT \keys_reg[3][65]  ( .D(n3214), .CLK(clk), .Q(n1731), .QN(n465) );
  DFFX1_HVT \keys_reg[3][64]  ( .D(n3213), .CLK(clk), .Q(n1732), .QN(n466) );
  DFFX1_HVT \keys_reg[3][63]  ( .D(n3212), .CLK(clk), .Q(n1733), .QN(n467) );
  DFFX1_HVT \keys_reg[3][62]  ( .D(n3211), .CLK(clk), .Q(n1734), .QN(n468) );
  DFFX1_HVT \keys_reg[3][61]  ( .D(n3210), .CLK(clk), .Q(n1735), .QN(n469) );
  DFFX1_HVT \keys_reg[3][60]  ( .D(n3209), .CLK(clk), .Q(n1736), .QN(n470) );
  DFFX1_HVT \keys_reg[3][59]  ( .D(n3208), .CLK(clk), .Q(n1737), .QN(n471) );
  DFFX1_HVT \keys_reg[3][58]  ( .D(n3207), .CLK(clk), .Q(n1738), .QN(n472) );
  DFFX1_HVT \keys_reg[3][57]  ( .D(n3206), .CLK(clk), .Q(n1739), .QN(n473) );
  DFFX1_HVT \keys_reg[3][56]  ( .D(n3205), .CLK(clk), .Q(n1740), .QN(n474) );
  DFFX1_HVT \keys_reg[3][55]  ( .D(n3204), .CLK(clk), .Q(n1741), .QN(n475) );
  DFFX1_HVT \keys_reg[3][54]  ( .D(n3203), .CLK(clk), .Q(n1742), .QN(n476) );
  DFFX1_HVT \keys_reg[3][53]  ( .D(n3202), .CLK(clk), .Q(n1743), .QN(n477) );
  DFFX1_HVT \keys_reg[3][52]  ( .D(n3201), .CLK(clk), .Q(n1744), .QN(n478) );
  DFFX1_HVT \keys_reg[3][51]  ( .D(n3200), .CLK(clk), .Q(n1745), .QN(n479) );
  DFFX1_HVT \keys_reg[3][50]  ( .D(n3199), .CLK(clk), .Q(n1746), .QN(n480) );
  DFFX1_HVT \keys_reg[3][49]  ( .D(n3198), .CLK(clk), .Q(n1747), .QN(n481) );
  DFFX1_HVT \keys_reg[3][48]  ( .D(n3197), .CLK(clk), .Q(n1748), .QN(n482) );
  DFFX1_HVT \keys_reg[3][47]  ( .D(n3196), .CLK(clk), .Q(n1749), .QN(n483) );
  DFFX1_HVT \keys_reg[3][46]  ( .D(n3195), .CLK(clk), .Q(n1750), .QN(n484) );
  DFFX1_HVT \keys_reg[3][45]  ( .D(n3194), .CLK(clk), .Q(n1751), .QN(n485) );
  DFFX1_HVT \keys_reg[3][44]  ( .D(n3193), .CLK(clk), .Q(n1752), .QN(n486) );
  DFFX1_HVT \keys_reg[3][43]  ( .D(n3192), .CLK(clk), .Q(n1753), .QN(n487) );
  DFFX1_HVT \keys_reg[3][42]  ( .D(n3191), .CLK(clk), .Q(n1754), .QN(n488) );
  DFFX1_HVT \keys_reg[3][41]  ( .D(n3190), .CLK(clk), .Q(n1755), .QN(n489) );
  DFFX1_HVT \keys_reg[3][40]  ( .D(n3189), .CLK(clk), .Q(n1756), .QN(n490) );
  DFFX1_HVT \keys_reg[3][39]  ( .D(n3188), .CLK(clk), .Q(n1757), .QN(n491) );
  DFFX1_HVT \keys_reg[3][38]  ( .D(n3187), .CLK(clk), .Q(n1758), .QN(n492) );
  DFFX1_HVT \keys_reg[3][37]  ( .D(n3186), .CLK(clk), .Q(n1759), .QN(n493) );
  DFFX1_HVT \keys_reg[3][36]  ( .D(n3185), .CLK(clk), .Q(n1760), .QN(n494) );
  DFFX1_HVT \keys_reg[3][35]  ( .D(n3184), .CLK(clk), .Q(n1761), .QN(n495) );
  DFFX1_HVT \keys_reg[3][34]  ( .D(n3183), .CLK(clk), .Q(n1762), .QN(n496) );
  DFFX1_HVT \keys_reg[3][33]  ( .D(n3182), .CLK(clk), .Q(n1763), .QN(n497) );
  DFFX1_HVT \keys_reg[3][32]  ( .D(n3181), .CLK(clk), .Q(n1764), .QN(n498) );
  DFFX1_HVT \keys_reg[3][31]  ( .D(n3180), .CLK(clk), .Q(n1765), .QN(n499) );
  DFFX1_HVT \keys_reg[3][30]  ( .D(n3179), .CLK(clk), .Q(n1766), .QN(n500) );
  DFFX1_HVT \keys_reg[3][29]  ( .D(n3178), .CLK(clk), .Q(n1767), .QN(n501) );
  DFFX1_HVT \keys_reg[3][28]  ( .D(n3177), .CLK(clk), .Q(n1768), .QN(n502) );
  DFFX1_HVT \keys_reg[3][27]  ( .D(n3176), .CLK(clk), .Q(n1769), .QN(n503) );
  DFFX1_HVT \keys_reg[3][26]  ( .D(n3175), .CLK(clk), .Q(n1770), .QN(n504) );
  DFFX1_HVT \keys_reg[3][25]  ( .D(n3174), .CLK(clk), .Q(n1771), .QN(n505) );
  DFFX1_HVT \keys_reg[3][24]  ( .D(n3173), .CLK(clk), .Q(n1772), .QN(n506) );
  DFFX1_HVT \keys_reg[3][23]  ( .D(n3172), .CLK(clk), .Q(n1773), .QN(n507) );
  DFFX1_HVT \keys_reg[3][22]  ( .D(n3171), .CLK(clk), .Q(n1774), .QN(n508) );
  DFFX1_HVT \keys_reg[3][21]  ( .D(n3170), .CLK(clk), .Q(n1775), .QN(n509) );
  DFFX1_HVT \keys_reg[3][20]  ( .D(n3169), .CLK(clk), .Q(n1776), .QN(n510) );
  DFFX1_HVT \keys_reg[3][19]  ( .D(n3168), .CLK(clk), .Q(n1777), .QN(n511) );
  DFFX1_HVT \keys_reg[3][18]  ( .D(n3167), .CLK(clk), .Q(n1778), .QN(n512) );
  DFFX1_HVT \keys_reg[3][17]  ( .D(n3166), .CLK(clk), .Q(n1779), .QN(n513) );
  DFFX1_HVT \keys_reg[3][16]  ( .D(n3165), .CLK(clk), .Q(n1780), .QN(n514) );
  DFFX1_HVT \keys_reg[3][15]  ( .D(n3164), .CLK(clk), .Q(n1781), .QN(n515) );
  DFFX1_HVT \keys_reg[3][14]  ( .D(n3163), .CLK(clk), .Q(n1782), .QN(n516) );
  DFFX1_HVT \keys_reg[3][13]  ( .D(n3162), .CLK(clk), .Q(n1783), .QN(n517) );
  DFFX1_HVT \keys_reg[3][12]  ( .D(n3161), .CLK(clk), .Q(n1784), .QN(n518) );
  DFFX1_HVT \keys_reg[3][11]  ( .D(n3160), .CLK(clk), .Q(n1785), .QN(n519) );
  DFFX1_HVT \keys_reg[3][10]  ( .D(n3159), .CLK(clk), .Q(n1786), .QN(n520) );
  DFFX1_HVT \keys_reg[3][9]  ( .D(n3158), .CLK(clk), .Q(n1787), .QN(n521) );
  DFFX1_HVT \keys_reg[3][8]  ( .D(n3157), .CLK(clk), .Q(n1788), .QN(n522) );
  DFFX1_HVT \keys_reg[3][7]  ( .D(n3156), .CLK(clk), .Q(n1789), .QN(n523) );
  DFFX1_HVT \keys_reg[3][6]  ( .D(n3155), .CLK(clk), .Q(n1790), .QN(n524) );
  DFFX1_HVT \keys_reg[3][5]  ( .D(n3154), .CLK(clk), .Q(n1791), .QN(n525) );
  DFFX1_HVT \keys_reg[3][4]  ( .D(n3153), .CLK(clk), .Q(n1792), .QN(n526) );
  DFFX1_HVT \keys_reg[3][3]  ( .D(n3152), .CLK(clk), .Q(n1793), .QN(n527) );
  DFFX1_HVT \keys_reg[3][2]  ( .D(n3151), .CLK(clk), .Q(n1794), .QN(n528) );
  DFFX1_HVT \keys_reg[3][1]  ( .D(n3150), .CLK(clk), .Q(n1795), .QN(n529) );
  DFFX1_HVT \keys_reg[3][0]  ( .D(n3149), .CLK(clk), .Q(n1796), .QN(n530) );
  DFFX1_HVT \keys_reg[4][127]  ( .D(n3148), .CLK(clk), .Q(n2053), .QN(n531) );
  DFFX1_HVT \keys_reg[4][126]  ( .D(n3147), .CLK(clk), .Q(n2054), .QN(n532) );
  DFFX1_HVT \keys_reg[4][125]  ( .D(n3146), .CLK(clk), .Q(n2055), .QN(n533) );
  DFFX1_HVT \keys_reg[4][124]  ( .D(n3145), .CLK(clk), .Q(n2056), .QN(n534) );
  DFFX1_HVT \keys_reg[4][123]  ( .D(n3144), .CLK(clk), .Q(n2057), .QN(n535) );
  DFFX1_HVT \keys_reg[4][122]  ( .D(n3143), .CLK(clk), .Q(n2058), .QN(n536) );
  DFFX1_HVT \keys_reg[4][121]  ( .D(n3142), .CLK(clk), .Q(n2059), .QN(n537) );
  DFFX1_HVT \keys_reg[4][120]  ( .D(n3141), .CLK(clk), .Q(n2060), .QN(n538) );
  DFFX1_HVT \keys_reg[4][119]  ( .D(n3140), .CLK(clk), .Q(n2061), .QN(n539) );
  DFFX1_HVT \keys_reg[4][118]  ( .D(n3139), .CLK(clk), .Q(n2062), .QN(n540) );
  DFFX1_HVT \keys_reg[4][117]  ( .D(n3138), .CLK(clk), .Q(n2063), .QN(n541) );
  DFFX1_HVT \keys_reg[4][116]  ( .D(n3137), .CLK(clk), .Q(n2064), .QN(n542) );
  DFFX1_HVT \keys_reg[4][115]  ( .D(n3136), .CLK(clk), .Q(n2065), .QN(n543) );
  DFFX1_HVT \keys_reg[4][114]  ( .D(n3135), .CLK(clk), .Q(n2066), .QN(n544) );
  DFFX1_HVT \keys_reg[4][113]  ( .D(n3134), .CLK(clk), .Q(n2067), .QN(n545) );
  DFFX1_HVT \keys_reg[4][112]  ( .D(n3133), .CLK(clk), .Q(n2068), .QN(n546) );
  DFFX1_HVT \keys_reg[4][111]  ( .D(n3132), .CLK(clk), .Q(n2069), .QN(n547) );
  DFFX1_HVT \keys_reg[4][110]  ( .D(n3131), .CLK(clk), .Q(n2070), .QN(n548) );
  DFFX1_HVT \keys_reg[4][109]  ( .D(n3130), .CLK(clk), .Q(n2071), .QN(n549) );
  DFFX1_HVT \keys_reg[4][108]  ( .D(n3129), .CLK(clk), .Q(n2072), .QN(n550) );
  DFFX1_HVT \keys_reg[4][107]  ( .D(n3128), .CLK(clk), .Q(n2073), .QN(n551) );
  DFFX1_HVT \keys_reg[4][106]  ( .D(n3127), .CLK(clk), .Q(n2074), .QN(n552) );
  DFFX1_HVT \keys_reg[4][105]  ( .D(n3126), .CLK(clk), .Q(n2075), .QN(n553) );
  DFFX1_HVT \keys_reg[4][104]  ( .D(n3125), .CLK(clk), .Q(n2076), .QN(n554) );
  DFFX1_HVT \keys_reg[4][103]  ( .D(n3124), .CLK(clk), .Q(n2077), .QN(n555) );
  DFFX1_HVT \keys_reg[4][102]  ( .D(n3123), .CLK(clk), .Q(n2078), .QN(n556) );
  DFFX1_HVT \keys_reg[4][101]  ( .D(n3122), .CLK(clk), .Q(n2079), .QN(n557) );
  DFFX1_HVT \keys_reg[4][100]  ( .D(n3121), .CLK(clk), .Q(n2080), .QN(n558) );
  DFFX1_HVT \keys_reg[4][99]  ( .D(n3120), .CLK(clk), .Q(n2081), .QN(n559) );
  DFFX1_HVT \keys_reg[4][98]  ( .D(n3119), .CLK(clk), .Q(n2082), .QN(n560) );
  DFFX1_HVT \keys_reg[4][97]  ( .D(n3118), .CLK(clk), .Q(n2083), .QN(n561) );
  DFFX1_HVT \keys_reg[4][96]  ( .D(n3117), .CLK(clk), .Q(n2084), .QN(n562) );
  DFFX1_HVT \keys_reg[4][95]  ( .D(n3116), .CLK(clk), .Q(n2085), .QN(n563) );
  DFFX1_HVT \keys_reg[4][94]  ( .D(n3115), .CLK(clk), .Q(n2086), .QN(n564) );
  DFFX1_HVT \keys_reg[4][93]  ( .D(n3114), .CLK(clk), .Q(n2087), .QN(n565) );
  DFFX1_HVT \keys_reg[4][92]  ( .D(n3113), .CLK(clk), .Q(n2088), .QN(n566) );
  DFFX1_HVT \keys_reg[4][91]  ( .D(n3112), .CLK(clk), .Q(n2089), .QN(n567) );
  DFFX1_HVT \keys_reg[4][90]  ( .D(n3111), .CLK(clk), .Q(n2090), .QN(n568) );
  DFFX1_HVT \keys_reg[4][89]  ( .D(n3110), .CLK(clk), .Q(n2091), .QN(n569) );
  DFFX1_HVT \keys_reg[4][88]  ( .D(n3109), .CLK(clk), .Q(n2092), .QN(n570) );
  DFFX1_HVT \keys_reg[4][87]  ( .D(n3108), .CLK(clk), .Q(n2093), .QN(n571) );
  DFFX1_HVT \keys_reg[4][86]  ( .D(n3107), .CLK(clk), .Q(n2094), .QN(n572) );
  DFFX1_HVT \keys_reg[4][85]  ( .D(n3106), .CLK(clk), .Q(n2095), .QN(n573) );
  DFFX1_HVT \keys_reg[4][84]  ( .D(n3105), .CLK(clk), .Q(n2096), .QN(n574) );
  DFFX1_HVT \keys_reg[4][83]  ( .D(n3104), .CLK(clk), .Q(n2097), .QN(n575) );
  DFFX1_HVT \keys_reg[4][82]  ( .D(n3103), .CLK(clk), .Q(n2098), .QN(n576) );
  DFFX1_HVT \keys_reg[4][81]  ( .D(n3102), .CLK(clk), .Q(n2099), .QN(n577) );
  DFFX1_HVT \keys_reg[4][80]  ( .D(n3101), .CLK(clk), .Q(n2100), .QN(n578) );
  DFFX1_HVT \keys_reg[4][79]  ( .D(n3100), .CLK(clk), .Q(n2101), .QN(n579) );
  DFFX1_HVT \keys_reg[4][78]  ( .D(n3099), .CLK(clk), .Q(n2102), .QN(n580) );
  DFFX1_HVT \keys_reg[4][77]  ( .D(n3098), .CLK(clk), .Q(n2103), .QN(n581) );
  DFFX1_HVT \keys_reg[4][76]  ( .D(n3097), .CLK(clk), .Q(n2104), .QN(n582) );
  DFFX1_HVT \keys_reg[4][75]  ( .D(n3096), .CLK(clk), .Q(n2105), .QN(n583) );
  DFFX1_HVT \keys_reg[4][74]  ( .D(n3095), .CLK(clk), .Q(n2106), .QN(n584) );
  DFFX1_HVT \keys_reg[4][73]  ( .D(n3094), .CLK(clk), .Q(n2107), .QN(n585) );
  DFFX1_HVT \keys_reg[4][72]  ( .D(n3093), .CLK(clk), .Q(n2108), .QN(n586) );
  DFFX1_HVT \keys_reg[4][71]  ( .D(n3092), .CLK(clk), .Q(n2109), .QN(n587) );
  DFFX1_HVT \keys_reg[4][70]  ( .D(n3091), .CLK(clk), .Q(n2110), .QN(n588) );
  DFFX1_HVT \keys_reg[4][69]  ( .D(n3090), .CLK(clk), .Q(n2111), .QN(n589) );
  DFFX1_HVT \keys_reg[4][68]  ( .D(n3089), .CLK(clk), .Q(n2112), .QN(n590) );
  DFFX1_HVT \keys_reg[4][67]  ( .D(n3088), .CLK(clk), .Q(n2113), .QN(n591) );
  DFFX1_HVT \keys_reg[4][66]  ( .D(n3087), .CLK(clk), .Q(n2114), .QN(n592) );
  DFFX1_HVT \keys_reg[4][65]  ( .D(n3086), .CLK(clk), .Q(n2115), .QN(n593) );
  DFFX1_HVT \keys_reg[4][64]  ( .D(n3085), .CLK(clk), .Q(n2116), .QN(n594) );
  DFFX1_HVT \keys_reg[4][63]  ( .D(n3084), .CLK(clk), .Q(n2117), .QN(n595) );
  DFFX1_HVT \keys_reg[4][62]  ( .D(n3083), .CLK(clk), .Q(n2118), .QN(n596) );
  DFFX1_HVT \keys_reg[4][61]  ( .D(n3082), .CLK(clk), .Q(n2119), .QN(n597) );
  DFFX1_HVT \keys_reg[4][60]  ( .D(n3081), .CLK(clk), .Q(n2120), .QN(n598) );
  DFFX1_HVT \keys_reg[4][59]  ( .D(n3080), .CLK(clk), .Q(n2121), .QN(n599) );
  DFFX1_HVT \keys_reg[4][58]  ( .D(n3079), .CLK(clk), .Q(n2122), .QN(n600) );
  DFFX1_HVT \keys_reg[4][57]  ( .D(n3078), .CLK(clk), .Q(n2123), .QN(n601) );
  DFFX1_HVT \keys_reg[4][56]  ( .D(n3077), .CLK(clk), .Q(n2124), .QN(n602) );
  DFFX1_HVT \keys_reg[4][55]  ( .D(n3076), .CLK(clk), .Q(n3798), .QN(n603) );
  DFFX1_HVT \keys_reg[4][54]  ( .D(n3075), .CLK(clk), .Q(n3799), .QN(n604) );
  DFFX1_HVT \keys_reg[4][53]  ( .D(n3074), .CLK(clk), .Q(n3800), .QN(n605) );
  DFFX1_HVT \keys_reg[4][52]  ( .D(n3073), .CLK(clk), .Q(n3801), .QN(n606) );
  DFFX1_HVT \keys_reg[4][51]  ( .D(n3072), .CLK(clk), .Q(n3802), .QN(n607) );
  DFFX1_HVT \keys_reg[4][50]  ( .D(n3071), .CLK(clk), .Q(n3803), .QN(n608) );
  DFFX1_HVT \keys_reg[4][49]  ( .D(n3070), .CLK(clk), .Q(n3804), .QN(n609) );
  DFFX1_HVT \keys_reg[4][48]  ( .D(n3069), .CLK(clk), .Q(n3805), .QN(n610) );
  DFFX1_HVT \keys_reg[4][47]  ( .D(n3068), .CLK(clk), .Q(n3806), .QN(n611) );
  DFFX1_HVT \keys_reg[4][46]  ( .D(n3067), .CLK(clk), .Q(n3807), .QN(n612) );
  DFFX1_HVT \keys_reg[4][45]  ( .D(n3066), .CLK(clk), .Q(n3808), .QN(n613) );
  DFFX1_HVT \keys_reg[4][44]  ( .D(n3065), .CLK(clk), .Q(n3809), .QN(n614) );
  DFFX1_HVT \keys_reg[4][43]  ( .D(n3064), .CLK(clk), .Q(n3810), .QN(n615) );
  DFFX1_HVT \keys_reg[4][42]  ( .D(n3063), .CLK(clk), .Q(n3811), .QN(n616) );
  DFFX1_HVT \keys_reg[4][41]  ( .D(n3062), .CLK(clk), .Q(n3812), .QN(n617) );
  DFFX1_HVT \keys_reg[4][40]  ( .D(n3061), .CLK(clk), .Q(n3813), .QN(n618) );
  DFFX1_HVT \keys_reg[4][39]  ( .D(n3060), .CLK(clk), .Q(n3814), .QN(n619) );
  DFFX1_HVT \keys_reg[4][38]  ( .D(n3059), .CLK(clk), .Q(n3815), .QN(n620) );
  DFFX1_HVT \keys_reg[4][37]  ( .D(n3058), .CLK(clk), .Q(n3816), .QN(n621) );
  DFFX1_HVT \keys_reg[4][36]  ( .D(n3057), .CLK(clk), .Q(n3817), .QN(n622) );
  DFFX1_HVT \keys_reg[4][35]  ( .D(n3056), .CLK(clk), .Q(n3818), .QN(n623) );
  DFFX1_HVT \keys_reg[4][34]  ( .D(n3055), .CLK(clk), .Q(n3819), .QN(n624) );
  DFFX1_HVT \keys_reg[4][33]  ( .D(n3054), .CLK(clk), .Q(n3820), .QN(n625) );
  DFFX1_HVT \keys_reg[4][32]  ( .D(n3053), .CLK(clk), .Q(n3821), .QN(n626) );
  DFFX1_HVT \keys_reg[4][31]  ( .D(n3052), .CLK(clk), .Q(n3822), .QN(n627) );
  DFFX1_HVT \keys_reg[4][30]  ( .D(n3051), .CLK(clk), .Q(n3823), .QN(n628) );
  DFFX1_HVT \keys_reg[4][29]  ( .D(n3050), .CLK(clk), .Q(n3824), .QN(n629) );
  DFFX1_HVT \keys_reg[4][28]  ( .D(n3049), .CLK(clk), .Q(n3825), .QN(n630) );
  DFFX1_HVT \keys_reg[4][27]  ( .D(n3048), .CLK(clk), .Q(n3826), .QN(n631) );
  DFFX1_HVT \keys_reg[4][26]  ( .D(n3047), .CLK(clk), .Q(n3827), .QN(n632) );
  DFFX1_HVT \keys_reg[4][25]  ( .D(n3046), .CLK(clk), .Q(n3828), .QN(n633) );
  DFFX1_HVT \keys_reg[4][24]  ( .D(n3045), .CLK(clk), .Q(n3829), .QN(n634) );
  DFFX1_HVT \keys_reg[4][23]  ( .D(n3044), .CLK(clk), .Q(n3830), .QN(n635) );
  DFFX1_HVT \keys_reg[4][22]  ( .D(n3043), .CLK(clk), .Q(n3831), .QN(n636) );
  DFFX1_HVT \keys_reg[4][21]  ( .D(n3042), .CLK(clk), .Q(n3832), .QN(n637) );
  DFFX1_HVT \keys_reg[4][20]  ( .D(n3041), .CLK(clk), .Q(n3833), .QN(n638) );
  DFFX1_HVT \keys_reg[4][19]  ( .D(n3040), .CLK(clk), .Q(n3834), .QN(n639) );
  DFFX1_HVT \keys_reg[4][18]  ( .D(n3039), .CLK(clk), .Q(n3835), .QN(n640) );
  DFFX1_HVT \keys_reg[4][17]  ( .D(n3038), .CLK(clk), .Q(n3836), .QN(n641) );
  DFFX1_HVT \keys_reg[4][16]  ( .D(n3037), .CLK(clk), .Q(n3837), .QN(n642) );
  DFFX1_HVT \keys_reg[4][15]  ( .D(n3036), .CLK(clk), .Q(n3838), .QN(n643) );
  DFFX1_HVT \keys_reg[4][14]  ( .D(n3035), .CLK(clk), .Q(n3839), .QN(n644) );
  DFFX1_HVT \keys_reg[4][13]  ( .D(n3034), .CLK(clk), .Q(n3840), .QN(n645) );
  DFFX1_HVT \keys_reg[4][12]  ( .D(n3033), .CLK(clk), .Q(n3841), .QN(n646) );
  DFFX1_HVT \keys_reg[4][11]  ( .D(n3032), .CLK(clk), .Q(n3842), .QN(n647) );
  DFFX1_HVT \keys_reg[4][10]  ( .D(n3031), .CLK(clk), .Q(n3843), .QN(n648) );
  DFFX1_HVT \keys_reg[4][9]  ( .D(n3030), .CLK(clk), .Q(n3844), .QN(n649) );
  DFFX1_HVT \keys_reg[4][8]  ( .D(n3029), .CLK(clk), .Q(n3845), .QN(n650) );
  DFFX1_HVT \keys_reg[4][7]  ( .D(n3028), .CLK(clk), .Q(n3846), .QN(n651) );
  DFFX1_HVT \keys_reg[4][6]  ( .D(n3027), .CLK(clk), .Q(n3847), .QN(n652) );
  DFFX1_HVT \keys_reg[4][5]  ( .D(n3026), .CLK(clk), .Q(n3848), .QN(n653) );
  DFFX1_HVT \keys_reg[4][4]  ( .D(n3025), .CLK(clk), .Q(n3849), .QN(n654) );
  DFFX1_HVT \keys_reg[4][3]  ( .D(n3024), .CLK(clk), .Q(n3850), .QN(n655) );
  DFFX1_HVT \keys_reg[4][2]  ( .D(n3023), .CLK(clk), .Q(n3851), .QN(n656) );
  DFFX1_HVT \keys_reg[4][1]  ( .D(n3022), .CLK(clk), .Q(n3852), .QN(n657) );
  DFFX1_HVT \keys_reg[4][0]  ( .D(n3021), .CLK(clk), .Q(n3853), .QN(n658) );
  DFFX1_HVT \keys_reg[5][127]  ( .D(n3020), .CLK(clk), .Q(n4110), .QN(n659) );
  DFFX1_HVT \keys_reg[5][126]  ( .D(n3019), .CLK(clk), .Q(n4111), .QN(n660) );
  DFFX1_HVT \keys_reg[5][125]  ( .D(n3018), .CLK(clk), .Q(n4112), .QN(n661) );
  DFFX1_HVT \keys_reg[5][124]  ( .D(n3017), .CLK(clk), .Q(n4113), .QN(n662) );
  DFFX1_HVT \keys_reg[5][123]  ( .D(n3016), .CLK(clk), .Q(n4114), .QN(n663) );
  DFFX1_HVT \keys_reg[5][122]  ( .D(n3015), .CLK(clk), .Q(n4115), .QN(n664) );
  DFFX1_HVT \keys_reg[5][121]  ( .D(n3014), .CLK(clk), .Q(n4116), .QN(n665) );
  DFFX1_HVT \keys_reg[5][120]  ( .D(n3013), .CLK(clk), .Q(n4117), .QN(n666) );
  DFFX1_HVT \keys_reg[5][119]  ( .D(n3012), .CLK(clk), .Q(n4118), .QN(n667) );
  DFFX1_HVT \keys_reg[5][118]  ( .D(n3011), .CLK(clk), .Q(n4119), .QN(n668) );
  DFFX1_HVT \keys_reg[5][117]  ( .D(n3010), .CLK(clk), .Q(n4120), .QN(n669) );
  DFFX1_HVT \keys_reg[5][116]  ( .D(n3009), .CLK(clk), .Q(n4121), .QN(n670) );
  DFFX1_HVT \keys_reg[5][115]  ( .D(n3008), .CLK(clk), .Q(n4122), .QN(n671) );
  DFFX1_HVT \keys_reg[5][114]  ( .D(n3007), .CLK(clk), .Q(n4123), .QN(n672) );
  DFFX1_HVT \keys_reg[5][113]  ( .D(n3006), .CLK(clk), .Q(n4124), .QN(n673) );
  DFFX1_HVT \keys_reg[5][112]  ( .D(n3005), .CLK(clk), .Q(n4125), .QN(n674) );
  DFFX1_HVT \keys_reg[5][111]  ( .D(n3004), .CLK(clk), .Q(n4126), .QN(n675) );
  DFFX1_HVT \keys_reg[5][110]  ( .D(n3003), .CLK(clk), .Q(n4127), .QN(n676) );
  DFFX1_HVT \keys_reg[5][109]  ( .D(n3002), .CLK(clk), .Q(n4128), .QN(n677) );
  DFFX1_HVT \keys_reg[5][108]  ( .D(n3001), .CLK(clk), .Q(n4129), .QN(n678) );
  DFFX1_HVT \keys_reg[5][107]  ( .D(n3000), .CLK(clk), .Q(n4130), .QN(n679) );
  DFFX1_HVT \keys_reg[5][106]  ( .D(n2999), .CLK(clk), .Q(n4131), .QN(n680) );
  DFFX1_HVT \keys_reg[5][105]  ( .D(n2998), .CLK(clk), .Q(n4132), .QN(n681) );
  DFFX1_HVT \keys_reg[5][104]  ( .D(n2997), .CLK(clk), .Q(n4133), .QN(n682) );
  DFFX1_HVT \keys_reg[5][103]  ( .D(n2996), .CLK(clk), .Q(n4134), .QN(n683) );
  DFFX1_HVT \keys_reg[5][102]  ( .D(n2995), .CLK(clk), .Q(n4135), .QN(n684) );
  DFFX1_HVT \keys_reg[5][101]  ( .D(n2994), .CLK(clk), .Q(n4136), .QN(n685) );
  DFFX1_HVT \keys_reg[5][100]  ( .D(n2993), .CLK(clk), .Q(n4137), .QN(n686) );
  DFFX1_HVT \keys_reg[5][99]  ( .D(n2992), .CLK(clk), .Q(n4138), .QN(n687) );
  DFFX1_HVT \keys_reg[5][98]  ( .D(n2991), .CLK(clk), .Q(n4139), .QN(n688) );
  DFFX1_HVT \keys_reg[5][97]  ( .D(n2990), .CLK(clk), .Q(n4140), .QN(n689) );
  DFFX1_HVT \keys_reg[5][96]  ( .D(n2989), .CLK(clk), .Q(n4141), .QN(n690) );
  DFFX1_HVT \keys_reg[5][95]  ( .D(n2988), .CLK(clk), .Q(n4142), .QN(n691) );
  DFFX1_HVT \keys_reg[5][94]  ( .D(n2987), .CLK(clk), .Q(n4143), .QN(n692) );
  DFFX1_HVT \keys_reg[5][93]  ( .D(n2986), .CLK(clk), .Q(n4144), .QN(n693) );
  DFFX1_HVT \keys_reg[5][92]  ( .D(n2985), .CLK(clk), .Q(n4145), .QN(n694) );
  DFFX1_HVT \keys_reg[5][91]  ( .D(n2984), .CLK(clk), .Q(n4146), .QN(n695) );
  DFFX1_HVT \keys_reg[5][90]  ( .D(n2983), .CLK(clk), .Q(n4147), .QN(n696) );
  DFFX1_HVT \keys_reg[5][89]  ( .D(n2982), .CLK(clk), .Q(n4148), .QN(n697) );
  DFFX1_HVT \keys_reg[5][88]  ( .D(n2981), .CLK(clk), .Q(n4149), .QN(n698) );
  DFFX1_HVT \keys_reg[5][87]  ( .D(n2980), .CLK(clk), .Q(n4150), .QN(n699) );
  DFFX1_HVT \keys_reg[5][86]  ( .D(n2979), .CLK(clk), .Q(n4151), .QN(n700) );
  DFFX1_HVT \keys_reg[5][85]  ( .D(n2978), .CLK(clk), .Q(n4152), .QN(n701) );
  DFFX1_HVT \keys_reg[5][84]  ( .D(n2977), .CLK(clk), .Q(n4153), .QN(n702) );
  DFFX1_HVT \keys_reg[5][83]  ( .D(n2976), .CLK(clk), .Q(n4154), .QN(n703) );
  DFFX1_HVT \keys_reg[5][82]  ( .D(n2975), .CLK(clk), .Q(n4155), .QN(n704) );
  DFFX1_HVT \keys_reg[5][81]  ( .D(n2974), .CLK(clk), .Q(n4156), .QN(n705) );
  DFFX1_HVT \keys_reg[5][80]  ( .D(n2973), .CLK(clk), .Q(n4157), .QN(n706) );
  DFFX1_HVT \keys_reg[5][79]  ( .D(n2972), .CLK(clk), .Q(n4158), .QN(n707) );
  DFFX1_HVT \keys_reg[5][78]  ( .D(n2971), .CLK(clk), .Q(n4159), .QN(n708) );
  DFFX1_HVT \keys_reg[5][77]  ( .D(n2970), .CLK(clk), .Q(n4160), .QN(n709) );
  DFFX1_HVT \keys_reg[5][76]  ( .D(n2969), .CLK(clk), .Q(n4161), .QN(n710) );
  DFFX1_HVT \keys_reg[5][75]  ( .D(n2968), .CLK(clk), .Q(n4162), .QN(n711) );
  DFFX1_HVT \keys_reg[5][74]  ( .D(n2967), .CLK(clk), .Q(n4163), .QN(n712) );
  DFFX1_HVT \keys_reg[5][73]  ( .D(n2966), .CLK(clk), .Q(n4164), .QN(n713) );
  DFFX1_HVT \keys_reg[5][72]  ( .D(n2965), .CLK(clk), .Q(n4165), .QN(n714) );
  DFFX1_HVT \keys_reg[5][71]  ( .D(n2964), .CLK(clk), .Q(n4166), .QN(n715) );
  DFFX1_HVT \keys_reg[5][70]  ( .D(n2963), .CLK(clk), .Q(n4167), .QN(n716) );
  DFFX1_HVT \keys_reg[5][69]  ( .D(n2962), .CLK(clk), .Q(n4168), .QN(n717) );
  DFFX1_HVT \keys_reg[5][68]  ( .D(n2961), .CLK(clk), .Q(n4169), .QN(n718) );
  DFFX1_HVT \keys_reg[5][67]  ( .D(n2960), .CLK(clk), .Q(n4170), .QN(n719) );
  DFFX1_HVT \keys_reg[5][66]  ( .D(n2959), .CLK(clk), .Q(n4171), .QN(n720) );
  DFFX1_HVT \keys_reg[5][65]  ( .D(n2958), .CLK(clk), .Q(n4172), .QN(n721) );
  DFFX1_HVT \keys_reg[5][64]  ( .D(n2957), .CLK(clk), .Q(n4173), .QN(n722) );
  DFFX1_HVT \keys_reg[5][63]  ( .D(n2956), .CLK(clk), .Q(n4174), .QN(n723) );
  DFFX1_HVT \keys_reg[5][62]  ( .D(n2955), .CLK(clk), .Q(n4175), .QN(n724) );
  DFFX1_HVT \keys_reg[5][61]  ( .D(n2954), .CLK(clk), .Q(n4176), .QN(n725) );
  DFFX1_HVT \keys_reg[5][60]  ( .D(n2953), .CLK(clk), .Q(n4177), .QN(n726) );
  DFFX1_HVT \keys_reg[5][59]  ( .D(n2952), .CLK(clk), .Q(n4178), .QN(n727) );
  DFFX1_HVT \keys_reg[5][58]  ( .D(n2951), .CLK(clk), .Q(n4179), .QN(n728) );
  DFFX1_HVT \keys_reg[5][57]  ( .D(n2950), .CLK(clk), .Q(n4180), .QN(n729) );
  DFFX1_HVT \keys_reg[5][56]  ( .D(n2949), .CLK(clk), .Q(n4181), .QN(n730) );
  DFFX1_HVT \keys_reg[5][55]  ( .D(n2948), .CLK(clk), .Q(n4182), .QN(n731) );
  DFFX1_HVT \keys_reg[5][54]  ( .D(n2947), .CLK(clk), .Q(n4183), .QN(n732) );
  DFFX1_HVT \keys_reg[5][53]  ( .D(n2946), .CLK(clk), .Q(n4184), .QN(n733) );
  DFFX1_HVT \keys_reg[5][52]  ( .D(n2945), .CLK(clk), .Q(n4185), .QN(n734) );
  DFFX1_HVT \keys_reg[5][51]  ( .D(n2944), .CLK(clk), .Q(n4186), .QN(n735) );
  DFFX1_HVT \keys_reg[5][50]  ( .D(n2943), .CLK(clk), .Q(n4187), .QN(n736) );
  DFFX1_HVT \keys_reg[5][49]  ( .D(n2942), .CLK(clk), .Q(n4188), .QN(n737) );
  DFFX1_HVT \keys_reg[5][48]  ( .D(n2941), .CLK(clk), .Q(n4189), .QN(n738) );
  DFFX1_HVT \keys_reg[5][47]  ( .D(n2940), .CLK(clk), .Q(n4190), .QN(n739) );
  DFFX1_HVT \keys_reg[5][46]  ( .D(n2939), .CLK(clk), .Q(n4191), .QN(n740) );
  DFFX1_HVT \keys_reg[5][45]  ( .D(n2938), .CLK(clk), .Q(n4192), .QN(n741) );
  DFFX1_HVT \keys_reg[5][44]  ( .D(n2937), .CLK(clk), .Q(n4193), .QN(n742) );
  DFFX1_HVT \keys_reg[5][43]  ( .D(n2936), .CLK(clk), .Q(n4194), .QN(n743) );
  DFFX1_HVT \keys_reg[5][42]  ( .D(n2935), .CLK(clk), .Q(n4195), .QN(n744) );
  DFFX1_HVT \keys_reg[5][41]  ( .D(n2934), .CLK(clk), .Q(n4196), .QN(n745) );
  DFFX1_HVT \keys_reg[5][40]  ( .D(n2933), .CLK(clk), .Q(n4197), .QN(n746) );
  DFFX1_HVT \keys_reg[5][39]  ( .D(n2932), .CLK(clk), .Q(n4198), .QN(n747) );
  DFFX1_HVT \keys_reg[5][38]  ( .D(n2931), .CLK(clk), .Q(n4199), .QN(n748) );
  DFFX1_HVT \keys_reg[5][37]  ( .D(n2930), .CLK(clk), .Q(n4200), .QN(n749) );
  DFFX1_HVT \keys_reg[5][36]  ( .D(n2929), .CLK(clk), .Q(n4201), .QN(n750) );
  DFFX1_HVT \keys_reg[5][35]  ( .D(n2928), .CLK(clk), .Q(n4202), .QN(n751) );
  DFFX1_HVT \keys_reg[5][34]  ( .D(n2927), .CLK(clk), .Q(n4203), .QN(n752) );
  DFFX1_HVT \keys_reg[5][33]  ( .D(n2926), .CLK(clk), .Q(n4204), .QN(n753) );
  DFFX1_HVT \keys_reg[5][32]  ( .D(n2925), .CLK(clk), .Q(n4205), .QN(n754) );
  DFFX1_HVT \keys_reg[5][31]  ( .D(n2924), .CLK(clk), .Q(n4206), .QN(n755) );
  DFFX1_HVT \keys_reg[5][30]  ( .D(n2923), .CLK(clk), .Q(n4207), .QN(n756) );
  DFFX1_HVT \keys_reg[5][29]  ( .D(n2922), .CLK(clk), .Q(n4208), .QN(n757) );
  DFFX1_HVT \keys_reg[5][28]  ( .D(n2921), .CLK(clk), .Q(n4209), .QN(n758) );
  DFFX1_HVT \keys_reg[5][27]  ( .D(n2920), .CLK(clk), .Q(n4210), .QN(n759) );
  DFFX1_HVT \keys_reg[5][26]  ( .D(n2919), .CLK(clk), .Q(n4211), .QN(n760) );
  DFFX1_HVT \keys_reg[5][25]  ( .D(n2918), .CLK(clk), .Q(n4212), .QN(n761) );
  DFFX1_HVT \keys_reg[5][24]  ( .D(n2917), .CLK(clk), .Q(n4213), .QN(n762) );
  DFFX1_HVT \keys_reg[5][23]  ( .D(n2916), .CLK(clk), .Q(n4214), .QN(n763) );
  DFFX1_HVT \keys_reg[5][22]  ( .D(n2915), .CLK(clk), .Q(n4215), .QN(n764) );
  DFFX1_HVT \keys_reg[5][21]  ( .D(n2914), .CLK(clk), .Q(n4216), .QN(n765) );
  DFFX1_HVT \keys_reg[5][20]  ( .D(n2913), .CLK(clk), .Q(n4217), .QN(n766) );
  DFFX1_HVT \keys_reg[5][19]  ( .D(n2912), .CLK(clk), .Q(n4218), .QN(n767) );
  DFFX1_HVT \keys_reg[5][18]  ( .D(n2911), .CLK(clk), .Q(n4219), .QN(n768) );
  DFFX1_HVT \keys_reg[5][17]  ( .D(n2910), .CLK(clk), .Q(n4220), .QN(n769) );
  DFFX1_HVT \keys_reg[5][16]  ( .D(n2909), .CLK(clk), .Q(n4221), .QN(n770) );
  DFFX1_HVT \keys_reg[5][15]  ( .D(n2908), .CLK(clk), .Q(n4222), .QN(n771) );
  DFFX1_HVT \keys_reg[5][14]  ( .D(n2907), .CLK(clk), .Q(n4223), .QN(n772) );
  DFFX1_HVT \keys_reg[5][13]  ( .D(n2906), .CLK(clk), .Q(n4224), .QN(n773) );
  DFFX1_HVT \keys_reg[5][12]  ( .D(n2905), .CLK(clk), .Q(n4225), .QN(n774) );
  DFFX1_HVT \keys_reg[5][11]  ( .D(n2904), .CLK(clk), .Q(n4226), .QN(n775) );
  DFFX1_HVT \keys_reg[5][10]  ( .D(n2903), .CLK(clk), .Q(n4227), .QN(n776) );
  DFFX1_HVT \keys_reg[5][9]  ( .D(n2902), .CLK(clk), .Q(n4228), .QN(n777) );
  DFFX1_HVT \keys_reg[5][8]  ( .D(n2901), .CLK(clk), .Q(n4229), .QN(n778) );
  DFFX1_HVT \keys_reg[5][7]  ( .D(n2900), .CLK(clk), .Q(n4230), .QN(n779) );
  DFFX1_HVT \keys_reg[5][6]  ( .D(n2899), .CLK(clk), .Q(n4231), .QN(n780) );
  DFFX1_HVT \keys_reg[5][5]  ( .D(n2898), .CLK(clk), .Q(n4232), .QN(n781) );
  DFFX1_HVT \keys_reg[5][4]  ( .D(n2897), .CLK(clk), .Q(n4233), .QN(n782) );
  DFFX1_HVT \keys_reg[5][3]  ( .D(n2896), .CLK(clk), .Q(n4234), .QN(n783) );
  DFFX1_HVT \keys_reg[5][2]  ( .D(n2895), .CLK(clk), .Q(n4235), .QN(n784) );
  DFFX1_HVT \keys_reg[5][1]  ( .D(n2894), .CLK(clk), .Q(n4236), .QN(n785) );
  DFFX1_HVT \keys_reg[5][0]  ( .D(n2893), .CLK(clk), .Q(n4237), .QN(n786) );
  DFFX1_HVT \keys_reg[6][127]  ( .D(n2892), .CLK(clk), .Q(n1797), .QN(n787) );
  DFFX1_HVT \keys_reg[6][126]  ( .D(n2891), .CLK(clk), .Q(n1798), .QN(n788) );
  DFFX1_HVT \keys_reg[6][125]  ( .D(n2890), .CLK(clk), .Q(n1799), .QN(n789) );
  DFFX1_HVT \keys_reg[6][124]  ( .D(n2889), .CLK(clk), .Q(n1800), .QN(n790) );
  DFFX1_HVT \keys_reg[6][123]  ( .D(n2888), .CLK(clk), .Q(n1801), .QN(n791) );
  DFFX1_HVT \keys_reg[6][122]  ( .D(n2887), .CLK(clk), .Q(n1802), .QN(n792) );
  DFFX1_HVT \keys_reg[6][121]  ( .D(n2886), .CLK(clk), .Q(n1803), .QN(n793) );
  DFFX1_HVT \keys_reg[6][120]  ( .D(n2885), .CLK(clk), .Q(n1804), .QN(n794) );
  DFFX1_HVT \keys_reg[6][119]  ( .D(n2884), .CLK(clk), .Q(n1805), .QN(n795) );
  DFFX1_HVT \keys_reg[6][118]  ( .D(n2883), .CLK(clk), .Q(n1806), .QN(n796) );
  DFFX1_HVT \keys_reg[6][117]  ( .D(n2882), .CLK(clk), .Q(n1807), .QN(n797) );
  DFFX1_HVT \keys_reg[6][116]  ( .D(n2881), .CLK(clk), .Q(n1808), .QN(n798) );
  DFFX1_HVT \keys_reg[6][115]  ( .D(n2880), .CLK(clk), .Q(n1809), .QN(n799) );
  DFFX1_HVT \keys_reg[6][114]  ( .D(n2879), .CLK(clk), .Q(n1810), .QN(n800) );
  DFFX1_HVT \keys_reg[6][113]  ( .D(n2878), .CLK(clk), .Q(n1811), .QN(n801) );
  DFFX1_HVT \keys_reg[6][112]  ( .D(n2877), .CLK(clk), .Q(n1812), .QN(n802) );
  DFFX1_HVT \keys_reg[6][111]  ( .D(n2876), .CLK(clk), .Q(n1813), .QN(n803) );
  DFFX1_HVT \keys_reg[6][110]  ( .D(n2875), .CLK(clk), .Q(n1814), .QN(n804) );
  DFFX1_HVT \keys_reg[6][109]  ( .D(n2874), .CLK(clk), .Q(n1815), .QN(n805) );
  DFFX1_HVT \keys_reg[6][108]  ( .D(n2873), .CLK(clk), .Q(n1816), .QN(n806) );
  DFFX1_HVT \keys_reg[6][107]  ( .D(n2872), .CLK(clk), .Q(n1817), .QN(n807) );
  DFFX1_HVT \keys_reg[6][106]  ( .D(n2871), .CLK(clk), .Q(n1818), .QN(n808) );
  DFFX1_HVT \keys_reg[6][105]  ( .D(n2870), .CLK(clk), .Q(n1819), .QN(n809) );
  DFFX1_HVT \keys_reg[6][104]  ( .D(n2869), .CLK(clk), .Q(n1820), .QN(n810) );
  DFFX1_HVT \keys_reg[6][103]  ( .D(n2868), .CLK(clk), .Q(n1821), .QN(n811) );
  DFFX1_HVT \keys_reg[6][102]  ( .D(n2867), .CLK(clk), .Q(n1822), .QN(n812) );
  DFFX1_HVT \keys_reg[6][101]  ( .D(n2866), .CLK(clk), .Q(n1823), .QN(n813) );
  DFFX1_HVT \keys_reg[6][100]  ( .D(n2865), .CLK(clk), .Q(n1824), .QN(n814) );
  DFFX1_HVT \keys_reg[6][99]  ( .D(n2864), .CLK(clk), .Q(n1825), .QN(n815) );
  DFFX1_HVT \keys_reg[6][98]  ( .D(n2863), .CLK(clk), .Q(n1826), .QN(n816) );
  DFFX1_HVT \keys_reg[6][97]  ( .D(n2862), .CLK(clk), .Q(n1827), .QN(n817) );
  DFFX1_HVT \keys_reg[6][96]  ( .D(n2861), .CLK(clk), .Q(n1828), .QN(n818) );
  DFFX1_HVT \keys_reg[6][95]  ( .D(n2860), .CLK(clk), .Q(n1829), .QN(n819) );
  DFFX1_HVT \keys_reg[6][94]  ( .D(n2859), .CLK(clk), .Q(n1830), .QN(n820) );
  DFFX1_HVT \keys_reg[6][93]  ( .D(n2858), .CLK(clk), .Q(n1831), .QN(n821) );
  DFFX1_HVT \keys_reg[6][92]  ( .D(n2857), .CLK(clk), .Q(n1832), .QN(n822) );
  DFFX1_HVT \keys_reg[6][91]  ( .D(n2856), .CLK(clk), .Q(n1833), .QN(n823) );
  DFFX1_HVT \keys_reg[6][90]  ( .D(n2855), .CLK(clk), .Q(n1834), .QN(n824) );
  DFFX1_HVT \keys_reg[6][89]  ( .D(n2854), .CLK(clk), .Q(n1835), .QN(n825) );
  DFFX1_HVT \keys_reg[6][88]  ( .D(n2853), .CLK(clk), .Q(n1836), .QN(n826) );
  DFFX1_HVT \keys_reg[6][87]  ( .D(n2852), .CLK(clk), .Q(n1837), .QN(n827) );
  DFFX1_HVT \keys_reg[6][86]  ( .D(n2851), .CLK(clk), .Q(n1838), .QN(n828) );
  DFFX1_HVT \keys_reg[6][85]  ( .D(n2850), .CLK(clk), .Q(n1839), .QN(n829) );
  DFFX1_HVT \keys_reg[6][84]  ( .D(n2849), .CLK(clk), .Q(n1840), .QN(n830) );
  DFFX1_HVT \keys_reg[6][83]  ( .D(n2848), .CLK(clk), .Q(n1841), .QN(n831) );
  DFFX1_HVT \keys_reg[6][82]  ( .D(n2847), .CLK(clk), .Q(n1842), .QN(n832) );
  DFFX1_HVT \keys_reg[6][81]  ( .D(n2846), .CLK(clk), .Q(n1843), .QN(n833) );
  DFFX1_HVT \keys_reg[6][80]  ( .D(n2845), .CLK(clk), .Q(n1844), .QN(n834) );
  DFFX1_HVT \keys_reg[6][79]  ( .D(n2844), .CLK(clk), .Q(n1845), .QN(n835) );
  DFFX1_HVT \keys_reg[6][78]  ( .D(n2843), .CLK(clk), .Q(n1846), .QN(n836) );
  DFFX1_HVT \keys_reg[6][77]  ( .D(n2842), .CLK(clk), .Q(n1847), .QN(n837) );
  DFFX1_HVT \keys_reg[6][76]  ( .D(n2841), .CLK(clk), .Q(n1848), .QN(n838) );
  DFFX1_HVT \keys_reg[6][75]  ( .D(n2840), .CLK(clk), .Q(n1849), .QN(n839) );
  DFFX1_HVT \keys_reg[6][74]  ( .D(n2839), .CLK(clk), .Q(n1850), .QN(n840) );
  DFFX1_HVT \keys_reg[6][73]  ( .D(n2838), .CLK(clk), .Q(n1851), .QN(n841) );
  DFFX1_HVT \keys_reg[6][72]  ( .D(n2837), .CLK(clk), .Q(n1852), .QN(n842) );
  DFFX1_HVT \keys_reg[6][71]  ( .D(n2836), .CLK(clk), .Q(n1853), .QN(n843) );
  DFFX1_HVT \keys_reg[6][70]  ( .D(n2835), .CLK(clk), .Q(n1854), .QN(n844) );
  DFFX1_HVT \keys_reg[6][69]  ( .D(n2834), .CLK(clk), .Q(n1855), .QN(n845) );
  DFFX1_HVT \keys_reg[6][68]  ( .D(n2833), .CLK(clk), .Q(n1856), .QN(n846) );
  DFFX1_HVT \keys_reg[6][67]  ( .D(n2832), .CLK(clk), .Q(n1857), .QN(n847) );
  DFFX1_HVT \keys_reg[6][66]  ( .D(n2831), .CLK(clk), .Q(n1858), .QN(n848) );
  DFFX1_HVT \keys_reg[6][65]  ( .D(n2830), .CLK(clk), .Q(n1859), .QN(n849) );
  DFFX1_HVT \keys_reg[6][64]  ( .D(n2829), .CLK(clk), .Q(n1860), .QN(n850) );
  DFFX1_HVT \keys_reg[6][63]  ( .D(n2828), .CLK(clk), .Q(n1861), .QN(n851) );
  DFFX1_HVT \keys_reg[6][62]  ( .D(n2827), .CLK(clk), .Q(n1862), .QN(n852) );
  DFFX1_HVT \keys_reg[6][61]  ( .D(n2826), .CLK(clk), .Q(n1863), .QN(n853) );
  DFFX1_HVT \keys_reg[6][60]  ( .D(n2825), .CLK(clk), .Q(n1864), .QN(n854) );
  DFFX1_HVT \keys_reg[6][59]  ( .D(n2824), .CLK(clk), .Q(n1865), .QN(n855) );
  DFFX1_HVT \keys_reg[6][58]  ( .D(n2823), .CLK(clk), .Q(n1866), .QN(n856) );
  DFFX1_HVT \keys_reg[6][57]  ( .D(n2822), .CLK(clk), .Q(n1867), .QN(n857) );
  DFFX1_HVT \keys_reg[6][56]  ( .D(n2821), .CLK(clk), .Q(n1868), .QN(n858) );
  DFFX1_HVT \keys_reg[6][55]  ( .D(n2820), .CLK(clk), .Q(n1869), .QN(n859) );
  DFFX1_HVT \keys_reg[6][54]  ( .D(n2819), .CLK(clk), .Q(n1870), .QN(n860) );
  DFFX1_HVT \keys_reg[6][53]  ( .D(n2818), .CLK(clk), .Q(n1871), .QN(n861) );
  DFFX1_HVT \keys_reg[6][52]  ( .D(n2817), .CLK(clk), .Q(n1872), .QN(n862) );
  DFFX1_HVT \keys_reg[6][51]  ( .D(n2816), .CLK(clk), .Q(n1873), .QN(n863) );
  DFFX1_HVT \keys_reg[6][50]  ( .D(n2815), .CLK(clk), .Q(n1874), .QN(n864) );
  DFFX1_HVT \keys_reg[6][49]  ( .D(n2814), .CLK(clk), .Q(n1875), .QN(n865) );
  DFFX1_HVT \keys_reg[6][48]  ( .D(n2813), .CLK(clk), .Q(n1876), .QN(n866) );
  DFFX1_HVT \keys_reg[6][47]  ( .D(n2812), .CLK(clk), .Q(n1877), .QN(n867) );
  DFFX1_HVT \keys_reg[6][46]  ( .D(n2811), .CLK(clk), .Q(n1878), .QN(n868) );
  DFFX1_HVT \keys_reg[6][45]  ( .D(n2810), .CLK(clk), .Q(n1879), .QN(n869) );
  DFFX1_HVT \keys_reg[6][44]  ( .D(n2809), .CLK(clk), .Q(n1880), .QN(n870) );
  DFFX1_HVT \keys_reg[6][43]  ( .D(n2808), .CLK(clk), .Q(n1881), .QN(n871) );
  DFFX1_HVT \keys_reg[6][42]  ( .D(n2807), .CLK(clk), .Q(n1882), .QN(n872) );
  DFFX1_HVT \keys_reg[6][41]  ( .D(n2806), .CLK(clk), .Q(n1883), .QN(n873) );
  DFFX1_HVT \keys_reg[6][40]  ( .D(n2805), .CLK(clk), .Q(n1884), .QN(n874) );
  DFFX1_HVT \keys_reg[6][39]  ( .D(n2804), .CLK(clk), .Q(n1885), .QN(n875) );
  DFFX1_HVT \keys_reg[6][38]  ( .D(n2803), .CLK(clk), .Q(n1886), .QN(n876) );
  DFFX1_HVT \keys_reg[6][37]  ( .D(n2802), .CLK(clk), .Q(n1887), .QN(n877) );
  DFFX1_HVT \keys_reg[6][36]  ( .D(n2801), .CLK(clk), .Q(n1888), .QN(n878) );
  DFFX1_HVT \keys_reg[6][35]  ( .D(n2800), .CLK(clk), .Q(n1889), .QN(n879) );
  DFFX1_HVT \keys_reg[6][34]  ( .D(n2799), .CLK(clk), .Q(n1890), .QN(n880) );
  DFFX1_HVT \keys_reg[6][33]  ( .D(n2798), .CLK(clk), .Q(n1891), .QN(n881) );
  DFFX1_HVT \keys_reg[6][32]  ( .D(n2797), .CLK(clk), .Q(n1892), .QN(n882) );
  DFFX1_HVT \keys_reg[6][31]  ( .D(n2796), .CLK(clk), .Q(n1893), .QN(n883) );
  DFFX1_HVT \keys_reg[6][30]  ( .D(n2795), .CLK(clk), .Q(n1894), .QN(n884) );
  DFFX1_HVT \keys_reg[6][29]  ( .D(n2794), .CLK(clk), .Q(n1895), .QN(n885) );
  DFFX1_HVT \keys_reg[6][28]  ( .D(n2793), .CLK(clk), .Q(n1896), .QN(n886) );
  DFFX1_HVT \keys_reg[6][27]  ( .D(n2792), .CLK(clk), .Q(n1897), .QN(n887) );
  DFFX1_HVT \keys_reg[6][26]  ( .D(n2791), .CLK(clk), .Q(n1898), .QN(n888) );
  DFFX1_HVT \keys_reg[6][25]  ( .D(n2790), .CLK(clk), .Q(n1899), .QN(n889) );
  DFFX1_HVT \keys_reg[6][24]  ( .D(n2789), .CLK(clk), .Q(n1900), .QN(n890) );
  DFFX1_HVT \keys_reg[6][23]  ( .D(n2788), .CLK(clk), .Q(n1901), .QN(n891) );
  DFFX1_HVT \keys_reg[6][22]  ( .D(n2787), .CLK(clk), .Q(n1902), .QN(n892) );
  DFFX1_HVT \keys_reg[6][21]  ( .D(n2786), .CLK(clk), .Q(n1903), .QN(n893) );
  DFFX1_HVT \keys_reg[6][20]  ( .D(n2785), .CLK(clk), .Q(n1904), .QN(n894) );
  DFFX1_HVT \keys_reg[6][19]  ( .D(n2784), .CLK(clk), .Q(n1905), .QN(n895) );
  DFFX1_HVT \keys_reg[6][18]  ( .D(n2783), .CLK(clk), .Q(n1906), .QN(n896) );
  DFFX1_HVT \keys_reg[6][17]  ( .D(n2782), .CLK(clk), .Q(n1907), .QN(n897) );
  DFFX1_HVT \keys_reg[6][16]  ( .D(n2781), .CLK(clk), .Q(n1908), .QN(n898) );
  DFFX1_HVT \keys_reg[6][15]  ( .D(n2780), .CLK(clk), .Q(n1909), .QN(n899) );
  DFFX1_HVT \keys_reg[6][14]  ( .D(n2779), .CLK(clk), .Q(n1910), .QN(n900) );
  DFFX1_HVT \keys_reg[6][13]  ( .D(n2778), .CLK(clk), .Q(n1911), .QN(n901) );
  DFFX1_HVT \keys_reg[6][12]  ( .D(n2777), .CLK(clk), .Q(n1912), .QN(n902) );
  DFFX1_HVT \keys_reg[6][11]  ( .D(n2776), .CLK(clk), .Q(n1913), .QN(n903) );
  DFFX1_HVT \keys_reg[6][10]  ( .D(n2775), .CLK(clk), .Q(n1914), .QN(n904) );
  DFFX1_HVT \keys_reg[6][9]  ( .D(n2774), .CLK(clk), .Q(n1915), .QN(n905) );
  DFFX1_HVT \keys_reg[6][8]  ( .D(n2773), .CLK(clk), .Q(n1916), .QN(n906) );
  DFFX1_HVT \keys_reg[6][7]  ( .D(n2772), .CLK(clk), .Q(n1917), .QN(n907) );
  DFFX1_HVT \keys_reg[6][6]  ( .D(n2771), .CLK(clk), .Q(n1918), .QN(n908) );
  DFFX1_HVT \keys_reg[6][5]  ( .D(n2770), .CLK(clk), .Q(n1919), .QN(n909) );
  DFFX1_HVT \keys_reg[6][4]  ( .D(n2769), .CLK(clk), .Q(n1920), .QN(n910) );
  DFFX1_HVT \keys_reg[6][3]  ( .D(n2768), .CLK(clk), .Q(n1921), .QN(n911) );
  DFFX1_HVT \keys_reg[6][2]  ( .D(n2767), .CLK(clk), .Q(n1922), .QN(n912) );
  DFFX1_HVT \keys_reg[6][1]  ( .D(n2766), .CLK(clk), .Q(n1923), .QN(n913) );
  DFFX1_HVT \keys_reg[6][0]  ( .D(n2765), .CLK(clk), .Q(n1924), .QN(n914) );
  DFFX1_HVT \keys_reg[7][127]  ( .D(n2764), .CLK(clk), .Q(n3854), .QN(n915) );
  DFFX1_HVT \keys_reg[7][126]  ( .D(n2763), .CLK(clk), .Q(n3855), .QN(n916) );
  DFFX1_HVT \keys_reg[7][125]  ( .D(n2762), .CLK(clk), .Q(n3856), .QN(n917) );
  DFFX1_HVT \keys_reg[7][124]  ( .D(n2761), .CLK(clk), .Q(n3857), .QN(n918) );
  DFFX1_HVT \keys_reg[7][123]  ( .D(n2760), .CLK(clk), .Q(n3858), .QN(n919) );
  DFFX1_HVT \keys_reg[7][122]  ( .D(n2759), .CLK(clk), .Q(n3859), .QN(n920) );
  DFFX1_HVT \keys_reg[7][121]  ( .D(n2758), .CLK(clk), .Q(n3860), .QN(n921) );
  DFFX1_HVT \keys_reg[7][120]  ( .D(n2757), .CLK(clk), .Q(n3861), .QN(n922) );
  DFFX1_HVT \keys_reg[7][119]  ( .D(n2756), .CLK(clk), .Q(n3862), .QN(n923) );
  DFFX1_HVT \keys_reg[7][118]  ( .D(n2755), .CLK(clk), .Q(n3863), .QN(n924) );
  DFFX1_HVT \keys_reg[7][117]  ( .D(n2754), .CLK(clk), .Q(n3864), .QN(n925) );
  DFFX1_HVT \keys_reg[7][116]  ( .D(n2753), .CLK(clk), .Q(n3865), .QN(n926) );
  DFFX1_HVT \keys_reg[7][115]  ( .D(n2752), .CLK(clk), .Q(n3866), .QN(n927) );
  DFFX1_HVT \keys_reg[7][114]  ( .D(n2751), .CLK(clk), .Q(n3867), .QN(n928) );
  DFFX1_HVT \keys_reg[7][113]  ( .D(n2750), .CLK(clk), .Q(n3868), .QN(n929) );
  DFFX1_HVT \keys_reg[7][112]  ( .D(n2749), .CLK(clk), .Q(n3869), .QN(n930) );
  DFFX1_HVT \keys_reg[7][111]  ( .D(n2748), .CLK(clk), .Q(n3870), .QN(n931) );
  DFFX1_HVT \keys_reg[7][110]  ( .D(n2747), .CLK(clk), .Q(n3871), .QN(n932) );
  DFFX1_HVT \keys_reg[7][109]  ( .D(n2746), .CLK(clk), .Q(n3872), .QN(n933) );
  DFFX1_HVT \keys_reg[7][108]  ( .D(n2745), .CLK(clk), .Q(n3873), .QN(n934) );
  DFFX1_HVT \keys_reg[7][107]  ( .D(n2744), .CLK(clk), .Q(n3874), .QN(n935) );
  DFFX1_HVT \keys_reg[7][106]  ( .D(n2743), .CLK(clk), .Q(n3875), .QN(n936) );
  DFFX1_HVT \keys_reg[7][105]  ( .D(n2742), .CLK(clk), .Q(n3876), .QN(n937) );
  DFFX1_HVT \keys_reg[7][104]  ( .D(n2741), .CLK(clk), .Q(n3877), .QN(n938) );
  DFFX1_HVT \keys_reg[7][103]  ( .D(n2740), .CLK(clk), .Q(n3878), .QN(n939) );
  DFFX1_HVT \keys_reg[7][102]  ( .D(n2739), .CLK(clk), .Q(n3879), .QN(n940) );
  DFFX1_HVT \keys_reg[7][101]  ( .D(n2738), .CLK(clk), .Q(n3880), .QN(n941) );
  DFFX1_HVT \keys_reg[7][100]  ( .D(n2737), .CLK(clk), .Q(n3881), .QN(n942) );
  DFFX1_HVT \keys_reg[7][99]  ( .D(n2736), .CLK(clk), .Q(n3882), .QN(n943) );
  DFFX1_HVT \keys_reg[7][98]  ( .D(n2735), .CLK(clk), .Q(n3883), .QN(n944) );
  DFFX1_HVT \keys_reg[7][97]  ( .D(n2734), .CLK(clk), .Q(n3884), .QN(n945) );
  DFFX1_HVT \keys_reg[7][96]  ( .D(n2733), .CLK(clk), .Q(n3885), .QN(n946) );
  DFFX1_HVT \keys_reg[7][95]  ( .D(n2732), .CLK(clk), .Q(n3886), .QN(n947) );
  DFFX1_HVT \keys_reg[7][94]  ( .D(n2731), .CLK(clk), .Q(n3887), .QN(n948) );
  DFFX1_HVT \keys_reg[7][93]  ( .D(n2730), .CLK(clk), .Q(n3888), .QN(n949) );
  DFFX1_HVT \keys_reg[7][92]  ( .D(n2729), .CLK(clk), .Q(n3889), .QN(n950) );
  DFFX1_HVT \keys_reg[7][91]  ( .D(n2728), .CLK(clk), .Q(n3890), .QN(n951) );
  DFFX1_HVT \keys_reg[7][90]  ( .D(n2727), .CLK(clk), .Q(n3891), .QN(n952) );
  DFFX1_HVT \keys_reg[7][89]  ( .D(n2726), .CLK(clk), .Q(n3892), .QN(n953) );
  DFFX1_HVT \keys_reg[7][88]  ( .D(n2725), .CLK(clk), .Q(n3893), .QN(n954) );
  DFFX1_HVT \keys_reg[7][87]  ( .D(n2724), .CLK(clk), .Q(n3894), .QN(n955) );
  DFFX1_HVT \keys_reg[7][86]  ( .D(n2723), .CLK(clk), .Q(n3895), .QN(n956) );
  DFFX1_HVT \keys_reg[7][85]  ( .D(n2722), .CLK(clk), .Q(n3896), .QN(n957) );
  DFFX1_HVT \keys_reg[7][84]  ( .D(n2721), .CLK(clk), .Q(n3897), .QN(n958) );
  DFFX1_HVT \keys_reg[7][83]  ( .D(n2720), .CLK(clk), .Q(n3898), .QN(n959) );
  DFFX1_HVT \keys_reg[7][82]  ( .D(n2719), .CLK(clk), .Q(n3899), .QN(n960) );
  DFFX1_HVT \keys_reg[7][81]  ( .D(n2718), .CLK(clk), .Q(n3900), .QN(n961) );
  DFFX1_HVT \keys_reg[7][80]  ( .D(n2717), .CLK(clk), .Q(n3901), .QN(n962) );
  DFFX1_HVT \keys_reg[7][79]  ( .D(n2716), .CLK(clk), .Q(n3902), .QN(n963) );
  DFFX1_HVT \keys_reg[7][78]  ( .D(n2715), .CLK(clk), .Q(n3903), .QN(n964) );
  DFFX1_HVT \keys_reg[7][77]  ( .D(n2714), .CLK(clk), .Q(n3904), .QN(n965) );
  DFFX1_HVT \keys_reg[7][76]  ( .D(n2713), .CLK(clk), .Q(n3905), .QN(n966) );
  DFFX1_HVT \keys_reg[7][75]  ( .D(n2712), .CLK(clk), .Q(n3906), .QN(n967) );
  DFFX1_HVT \keys_reg[7][74]  ( .D(n2711), .CLK(clk), .Q(n3907), .QN(n968) );
  DFFX1_HVT \keys_reg[7][73]  ( .D(n2710), .CLK(clk), .Q(n3908), .QN(n969) );
  DFFX1_HVT \keys_reg[7][72]  ( .D(n2709), .CLK(clk), .Q(n3909), .QN(n970) );
  DFFX1_HVT \keys_reg[7][71]  ( .D(n2708), .CLK(clk), .Q(n3910), .QN(n971) );
  DFFX1_HVT \keys_reg[7][70]  ( .D(n2707), .CLK(clk), .Q(n3911), .QN(n972) );
  DFFX1_HVT \keys_reg[7][69]  ( .D(n2706), .CLK(clk), .Q(n3912), .QN(n973) );
  DFFX1_HVT \keys_reg[7][68]  ( .D(n2705), .CLK(clk), .Q(n3913), .QN(n974) );
  DFFX1_HVT \keys_reg[7][67]  ( .D(n2704), .CLK(clk), .Q(n3914), .QN(n975) );
  DFFX1_HVT \keys_reg[7][66]  ( .D(n2703), .CLK(clk), .Q(n3915), .QN(n976) );
  DFFX1_HVT \keys_reg[7][65]  ( .D(n2702), .CLK(clk), .Q(n3916), .QN(n977) );
  DFFX1_HVT \keys_reg[7][64]  ( .D(n2701), .CLK(clk), .Q(n3917), .QN(n978) );
  DFFX1_HVT \keys_reg[7][63]  ( .D(n2700), .CLK(clk), .Q(n3918), .QN(n979) );
  DFFX1_HVT \keys_reg[7][62]  ( .D(n2699), .CLK(clk), .Q(n3919), .QN(n980) );
  DFFX1_HVT \keys_reg[7][61]  ( .D(n2698), .CLK(clk), .Q(n3920), .QN(n981) );
  DFFX1_HVT \keys_reg[7][60]  ( .D(n2697), .CLK(clk), .Q(n3921), .QN(n982) );
  DFFX1_HVT \keys_reg[7][59]  ( .D(n2696), .CLK(clk), .Q(n3922), .QN(n983) );
  DFFX1_HVT \keys_reg[7][58]  ( .D(n2695), .CLK(clk), .Q(n3923), .QN(n984) );
  DFFX1_HVT \keys_reg[7][57]  ( .D(n2694), .CLK(clk), .Q(n3924), .QN(n985) );
  DFFX1_HVT \keys_reg[7][56]  ( .D(n2693), .CLK(clk), .Q(n3925), .QN(n986) );
  DFFX1_HVT \keys_reg[7][55]  ( .D(n2692), .CLK(clk), .Q(n3926), .QN(n987) );
  DFFX1_HVT \keys_reg[7][54]  ( .D(n2691), .CLK(clk), .Q(n3927), .QN(n988) );
  DFFX1_HVT \keys_reg[7][53]  ( .D(n2690), .CLK(clk), .Q(n3928), .QN(n989) );
  DFFX1_HVT \keys_reg[7][52]  ( .D(n2689), .CLK(clk), .Q(n3929), .QN(n990) );
  DFFX1_HVT \keys_reg[7][51]  ( .D(n2688), .CLK(clk), .Q(n3930), .QN(n991) );
  DFFX1_HVT \keys_reg[7][50]  ( .D(n2687), .CLK(clk), .Q(n3931), .QN(n992) );
  DFFX1_HVT \keys_reg[7][49]  ( .D(n2686), .CLK(clk), .Q(n3932), .QN(n993) );
  DFFX1_HVT \keys_reg[7][48]  ( .D(n2685), .CLK(clk), .Q(n3933), .QN(n994) );
  DFFX1_HVT \keys_reg[7][47]  ( .D(n2684), .CLK(clk), .Q(n3934), .QN(n995) );
  DFFX1_HVT \keys_reg[7][46]  ( .D(n2683), .CLK(clk), .Q(n3935), .QN(n996) );
  DFFX1_HVT \keys_reg[7][45]  ( .D(n2682), .CLK(clk), .Q(n3936), .QN(n997) );
  DFFX1_HVT \keys_reg[7][44]  ( .D(n2681), .CLK(clk), .Q(n3937), .QN(n998) );
  DFFX1_HVT \keys_reg[7][43]  ( .D(n2680), .CLK(clk), .Q(n3938), .QN(n999) );
  DFFX1_HVT \keys_reg[7][42]  ( .D(n2679), .CLK(clk), .Q(n3939), .QN(n1000) );
  DFFX1_HVT \keys_reg[7][41]  ( .D(n2678), .CLK(clk), .Q(n3940), .QN(n1001) );
  DFFX1_HVT \keys_reg[7][40]  ( .D(n2677), .CLK(clk), .Q(n3941), .QN(n1002) );
  DFFX1_HVT \keys_reg[7][39]  ( .D(n2676), .CLK(clk), .Q(n3942), .QN(n1003) );
  DFFX1_HVT \keys_reg[7][38]  ( .D(n2675), .CLK(clk), .Q(n3943), .QN(n1004) );
  DFFX1_HVT \keys_reg[7][37]  ( .D(n2674), .CLK(clk), .Q(n3944), .QN(n1005) );
  DFFX1_HVT \keys_reg[7][36]  ( .D(n2673), .CLK(clk), .Q(n3945), .QN(n1006) );
  DFFX1_HVT \keys_reg[7][35]  ( .D(n2672), .CLK(clk), .Q(n3946), .QN(n1007) );
  DFFX1_HVT \keys_reg[7][34]  ( .D(n2671), .CLK(clk), .Q(n3947), .QN(n1008) );
  DFFX1_HVT \keys_reg[7][33]  ( .D(n2670), .CLK(clk), .Q(n3948), .QN(n1009) );
  DFFX1_HVT \keys_reg[7][32]  ( .D(n2669), .CLK(clk), .Q(n3949), .QN(n1010) );
  DFFX1_HVT \keys_reg[7][31]  ( .D(n2668), .CLK(clk), .Q(n3950), .QN(n1011) );
  DFFX1_HVT \keys_reg[7][30]  ( .D(n2667), .CLK(clk), .Q(n3951), .QN(n1012) );
  DFFX1_HVT \keys_reg[7][29]  ( .D(n2666), .CLK(clk), .Q(n3952), .QN(n1013) );
  DFFX1_HVT \keys_reg[7][28]  ( .D(n2665), .CLK(clk), .Q(n3953), .QN(n1014) );
  DFFX1_HVT \keys_reg[7][27]  ( .D(n2664), .CLK(clk), .Q(n3954), .QN(n1015) );
  DFFX1_HVT \keys_reg[7][26]  ( .D(n2663), .CLK(clk), .Q(n3955), .QN(n1016) );
  DFFX1_HVT \keys_reg[7][25]  ( .D(n2662), .CLK(clk), .Q(n3956), .QN(n1017) );
  DFFX1_HVT \keys_reg[7][24]  ( .D(n2661), .CLK(clk), .Q(n3957), .QN(n1018) );
  DFFX1_HVT \keys_reg[7][23]  ( .D(n2660), .CLK(clk), .Q(n3958), .QN(n1019) );
  DFFX1_HVT \keys_reg[7][22]  ( .D(n2659), .CLK(clk), .Q(n3959), .QN(n1020) );
  DFFX1_HVT \keys_reg[7][21]  ( .D(n2658), .CLK(clk), .Q(n3960), .QN(n1021) );
  DFFX1_HVT \keys_reg[7][20]  ( .D(n2657), .CLK(clk), .Q(n3961), .QN(n1022) );
  DFFX1_HVT \keys_reg[7][19]  ( .D(n2656), .CLK(clk), .Q(n3962), .QN(n1023) );
  DFFX1_HVT \keys_reg[7][18]  ( .D(n2655), .CLK(clk), .Q(n3963), .QN(n1024) );
  DFFX1_HVT \keys_reg[7][17]  ( .D(n2654), .CLK(clk), .Q(n3964), .QN(n1025) );
  DFFX1_HVT \keys_reg[7][16]  ( .D(n2653), .CLK(clk), .Q(n3965), .QN(n1026) );
  DFFX1_HVT \keys_reg[7][15]  ( .D(n2652), .CLK(clk), .Q(n3966), .QN(n1027) );
  DFFX1_HVT \keys_reg[7][14]  ( .D(n2651), .CLK(clk), .Q(n3967), .QN(n1028) );
  DFFX1_HVT \keys_reg[7][13]  ( .D(n2650), .CLK(clk), .Q(n3968), .QN(n1029) );
  DFFX1_HVT \keys_reg[7][12]  ( .D(n2649), .CLK(clk), .Q(n3969), .QN(n1030) );
  DFFX1_HVT \keys_reg[7][11]  ( .D(n2648), .CLK(clk), .Q(n3970), .QN(n1031) );
  DFFX1_HVT \keys_reg[7][10]  ( .D(n2647), .CLK(clk), .Q(n3971), .QN(n1032) );
  DFFX1_HVT \keys_reg[7][9]  ( .D(n2646), .CLK(clk), .Q(n3972), .QN(n1033) );
  DFFX1_HVT \keys_reg[7][8]  ( .D(n2645), .CLK(clk), .Q(n3973), .QN(n1034) );
  DFFX1_HVT \keys_reg[7][7]  ( .D(n2644), .CLK(clk), .Q(n3974), .QN(n1035) );
  DFFX1_HVT \keys_reg[7][6]  ( .D(n2643), .CLK(clk), .Q(n3975), .QN(n1036) );
  DFFX1_HVT \keys_reg[7][5]  ( .D(n2642), .CLK(clk), .Q(n3976), .QN(n1037) );
  DFFX1_HVT \keys_reg[7][4]  ( .D(n2641), .CLK(clk), .Q(n3977), .QN(n1038) );
  DFFX1_HVT \keys_reg[7][3]  ( .D(n2640), .CLK(clk), .Q(n3978), .QN(n1039) );
  DFFX1_HVT \keys_reg[7][2]  ( .D(n2639), .CLK(clk), .Q(n3979), .QN(n1040) );
  DFFX1_HVT \keys_reg[7][1]  ( .D(n2638), .CLK(clk), .Q(n3980), .QN(n1041) );
  DFFX1_HVT \keys_reg[7][0]  ( .D(n2637), .CLK(clk), .Q(n3981), .QN(n1042) );
  DFFX1_HVT \keys_reg[8][127]  ( .D(n2636), .CLK(clk), .Q(n4238), .QN(n1043)
         );
  DFFX1_HVT \keys_reg[8][126]  ( .D(n2635), .CLK(clk), .Q(n4239), .QN(n1044)
         );
  DFFX1_HVT \keys_reg[8][125]  ( .D(n2634), .CLK(clk), .Q(n4240), .QN(n1045)
         );
  DFFX1_HVT \keys_reg[8][124]  ( .D(n2633), .CLK(clk), .Q(n4241), .QN(n1046)
         );
  DFFX1_HVT \keys_reg[8][123]  ( .D(n2632), .CLK(clk), .Q(n4242), .QN(n1047)
         );
  DFFX1_HVT \keys_reg[8][122]  ( .D(n2631), .CLK(clk), .Q(n4243), .QN(n1048)
         );
  DFFX1_HVT \keys_reg[8][121]  ( .D(n2630), .CLK(clk), .Q(n4244), .QN(n1049)
         );
  DFFX1_HVT \keys_reg[8][120]  ( .D(n2629), .CLK(clk), .Q(n4245), .QN(n1050)
         );
  DFFX1_HVT \keys_reg[8][119]  ( .D(n2628), .CLK(clk), .Q(n4246), .QN(n1051)
         );
  DFFX1_HVT \keys_reg[8][118]  ( .D(n2627), .CLK(clk), .Q(n4247), .QN(n1052)
         );
  DFFX1_HVT \keys_reg[8][117]  ( .D(n2626), .CLK(clk), .Q(n4248), .QN(n1053)
         );
  DFFX1_HVT \keys_reg[8][116]  ( .D(n2625), .CLK(clk), .Q(n4249), .QN(n1054)
         );
  DFFX1_HVT \keys_reg[8][115]  ( .D(n2624), .CLK(clk), .Q(n4250), .QN(n1055)
         );
  DFFX1_HVT \keys_reg[8][114]  ( .D(n2623), .CLK(clk), .Q(n4251), .QN(n1056)
         );
  DFFX1_HVT \keys_reg[8][113]  ( .D(n2622), .CLK(clk), .Q(n4252), .QN(n1057)
         );
  DFFX1_HVT \keys_reg[8][112]  ( .D(n2621), .CLK(clk), .Q(n4253), .QN(n1058)
         );
  DFFX1_HVT \keys_reg[8][111]  ( .D(n2620), .CLK(clk), .Q(n4254), .QN(n1059)
         );
  DFFX1_HVT \keys_reg[8][110]  ( .D(n2619), .CLK(clk), .Q(n4255), .QN(n1060)
         );
  DFFX1_HVT \keys_reg[8][109]  ( .D(n2618), .CLK(clk), .Q(n4256), .QN(n1061)
         );
  DFFX1_HVT \keys_reg[8][108]  ( .D(n2617), .CLK(clk), .Q(n4257), .QN(n1062)
         );
  DFFX1_HVT \keys_reg[8][107]  ( .D(n2616), .CLK(clk), .Q(n4258), .QN(n1063)
         );
  DFFX1_HVT \keys_reg[8][106]  ( .D(n2615), .CLK(clk), .Q(n4259), .QN(n1064)
         );
  DFFX1_HVT \keys_reg[8][105]  ( .D(n2614), .CLK(clk), .Q(n4260), .QN(n1065)
         );
  DFFX1_HVT \keys_reg[8][104]  ( .D(n2613), .CLK(clk), .Q(n4261), .QN(n1066)
         );
  DFFX1_HVT \keys_reg[8][103]  ( .D(n2612), .CLK(clk), .Q(n4262), .QN(n1067)
         );
  DFFX1_HVT \keys_reg[8][102]  ( .D(n2611), .CLK(clk), .Q(n4263), .QN(n1068)
         );
  DFFX1_HVT \keys_reg[8][101]  ( .D(n2610), .CLK(clk), .Q(n4264), .QN(n1069)
         );
  DFFX1_HVT \keys_reg[8][100]  ( .D(n2609), .CLK(clk), .Q(n4265), .QN(n1070)
         );
  DFFX1_HVT \keys_reg[8][99]  ( .D(n2608), .CLK(clk), .Q(n4266), .QN(n1071) );
  DFFX1_HVT \keys_reg[8][98]  ( .D(n2607), .CLK(clk), .Q(n4267), .QN(n1072) );
  DFFX1_HVT \keys_reg[8][97]  ( .D(n2606), .CLK(clk), .Q(n4268), .QN(n1073) );
  DFFX1_HVT \keys_reg[8][96]  ( .D(n2605), .CLK(clk), .Q(n4269), .QN(n1074) );
  DFFX1_HVT \keys_reg[8][95]  ( .D(n2604), .CLK(clk), .Q(n4270), .QN(n1075) );
  DFFX1_HVT \keys_reg[8][94]  ( .D(n2603), .CLK(clk), .Q(n4271), .QN(n1076) );
  DFFX1_HVT \keys_reg[8][93]  ( .D(n2602), .CLK(clk), .Q(n4272), .QN(n1077) );
  DFFX1_HVT \keys_reg[8][92]  ( .D(n2601), .CLK(clk), .Q(n4273), .QN(n1078) );
  DFFX1_HVT \keys_reg[8][91]  ( .D(n2600), .CLK(clk), .Q(n4274), .QN(n1079) );
  DFFX1_HVT \keys_reg[8][90]  ( .D(n2599), .CLK(clk), .Q(n4275), .QN(n1080) );
  DFFX1_HVT \keys_reg[8][89]  ( .D(n2598), .CLK(clk), .Q(n4276), .QN(n1081) );
  DFFX1_HVT \keys_reg[8][88]  ( .D(n2597), .CLK(clk), .Q(n4277), .QN(n1082) );
  DFFX1_HVT \keys_reg[8][87]  ( .D(n2596), .CLK(clk), .Q(n4278), .QN(n1083) );
  DFFX1_HVT \keys_reg[8][86]  ( .D(n2595), .CLK(clk), .Q(n4279), .QN(n1084) );
  DFFX1_HVT \keys_reg[8][85]  ( .D(n2594), .CLK(clk), .Q(n4280), .QN(n1085) );
  DFFX1_HVT \keys_reg[8][84]  ( .D(n2593), .CLK(clk), .Q(n4281), .QN(n1086) );
  DFFX1_HVT \keys_reg[8][83]  ( .D(n2592), .CLK(clk), .Q(n4282), .QN(n1087) );
  DFFX1_HVT \keys_reg[8][82]  ( .D(n2591), .CLK(clk), .Q(n4283), .QN(n1088) );
  DFFX1_HVT \keys_reg[8][81]  ( .D(n2590), .CLK(clk), .Q(n4284), .QN(n1089) );
  DFFX1_HVT \keys_reg[8][80]  ( .D(n2589), .CLK(clk), .Q(n4285), .QN(n1090) );
  DFFX1_HVT \keys_reg[8][79]  ( .D(n2588), .CLK(clk), .Q(n4286), .QN(n1091) );
  DFFX1_HVT \keys_reg[8][78]  ( .D(n2587), .CLK(clk), .Q(n4287), .QN(n1092) );
  DFFX1_HVT \keys_reg[8][77]  ( .D(n2586), .CLK(clk), .Q(n4288), .QN(n1093) );
  DFFX1_HVT \keys_reg[8][76]  ( .D(n2585), .CLK(clk), .Q(n4289), .QN(n1094) );
  DFFX1_HVT \keys_reg[8][75]  ( .D(n2584), .CLK(clk), .Q(n4290), .QN(n1095) );
  DFFX1_HVT \keys_reg[8][74]  ( .D(n2583), .CLK(clk), .Q(n4291), .QN(n1096) );
  DFFX1_HVT \keys_reg[8][73]  ( .D(n2582), .CLK(clk), .Q(n4292), .QN(n1097) );
  DFFX1_HVT \keys_reg[8][72]  ( .D(n2581), .CLK(clk), .Q(n4293), .QN(n1098) );
  DFFX1_HVT \keys_reg[8][71]  ( .D(n2580), .CLK(clk), .Q(n4294), .QN(n1099) );
  DFFX1_HVT \keys_reg[8][70]  ( .D(n2579), .CLK(clk), .Q(n4295), .QN(n1100) );
  DFFX1_HVT \keys_reg[8][69]  ( .D(n2578), .CLK(clk), .Q(n4296), .QN(n1101) );
  DFFX1_HVT \keys_reg[8][68]  ( .D(n2577), .CLK(clk), .Q(n4297), .QN(n1102) );
  DFFX1_HVT \keys_reg[8][67]  ( .D(n2576), .CLK(clk), .Q(n4298), .QN(n1103) );
  DFFX1_HVT \keys_reg[8][66]  ( .D(n2575), .CLK(clk), .Q(n4299), .QN(n1104) );
  DFFX1_HVT \keys_reg[8][65]  ( .D(n2574), .CLK(clk), .Q(n4300), .QN(n1105) );
  DFFX1_HVT \keys_reg[8][64]  ( .D(n2573), .CLK(clk), .Q(n4301), .QN(n1106) );
  DFFX1_HVT \keys_reg[8][63]  ( .D(n2572), .CLK(clk), .Q(n4302), .QN(n1107) );
  DFFX1_HVT \keys_reg[8][62]  ( .D(n2571), .CLK(clk), .Q(n4303), .QN(n1108) );
  DFFX1_HVT \keys_reg[8][61]  ( .D(n2570), .CLK(clk), .Q(n4304), .QN(n1109) );
  DFFX1_HVT \keys_reg[8][60]  ( .D(n2569), .CLK(clk), .Q(n4305), .QN(n1110) );
  DFFX1_HVT \keys_reg[8][59]  ( .D(n2568), .CLK(clk), .Q(n4306), .QN(n1111) );
  DFFX1_HVT \keys_reg[8][58]  ( .D(n2567), .CLK(clk), .Q(n4307), .QN(n1112) );
  DFFX1_HVT \keys_reg[8][57]  ( .D(n2566), .CLK(clk), .Q(n4308), .QN(n1113) );
  DFFX1_HVT \keys_reg[8][56]  ( .D(n2565), .CLK(clk), .Q(n4309), .QN(n1114) );
  DFFX1_HVT \keys_reg[8][55]  ( .D(n2564), .CLK(clk), .Q(n4310), .QN(n1115) );
  DFFX1_HVT \keys_reg[8][54]  ( .D(n2563), .CLK(clk), .Q(n4311), .QN(n1116) );
  DFFX1_HVT \keys_reg[8][53]  ( .D(n2562), .CLK(clk), .Q(n4312), .QN(n1117) );
  DFFX1_HVT \keys_reg[8][52]  ( .D(n2561), .CLK(clk), .Q(n4313), .QN(n1118) );
  DFFX1_HVT \keys_reg[8][51]  ( .D(n2560), .CLK(clk), .Q(n4314), .QN(n1119) );
  DFFX1_HVT \keys_reg[8][50]  ( .D(n2559), .CLK(clk), .Q(n4315), .QN(n1120) );
  DFFX1_HVT \keys_reg[8][49]  ( .D(n2558), .CLK(clk), .Q(n4316), .QN(n1121) );
  DFFX1_HVT \keys_reg[8][48]  ( .D(n2557), .CLK(clk), .Q(n4317), .QN(n1122) );
  DFFX1_HVT \keys_reg[8][47]  ( .D(n2556), .CLK(clk), .Q(n4318), .QN(n1123) );
  DFFX1_HVT \keys_reg[8][46]  ( .D(n2555), .CLK(clk), .Q(n4319), .QN(n1124) );
  DFFX1_HVT \keys_reg[8][45]  ( .D(n2554), .CLK(clk), .Q(n4320), .QN(n1125) );
  DFFX1_HVT \keys_reg[8][44]  ( .D(n2553), .CLK(clk), .Q(n4321), .QN(n1126) );
  DFFX1_HVT \keys_reg[8][43]  ( .D(n2552), .CLK(clk), .Q(n4322), .QN(n1127) );
  DFFX1_HVT \keys_reg[8][42]  ( .D(n2551), .CLK(clk), .Q(n4323), .QN(n1128) );
  DFFX1_HVT \keys_reg[8][41]  ( .D(n2550), .CLK(clk), .Q(n4324), .QN(n1129) );
  DFFX1_HVT \keys_reg[8][40]  ( .D(n2549), .CLK(clk), .Q(n4325), .QN(n1130) );
  DFFX1_HVT \keys_reg[8][39]  ( .D(n2548), .CLK(clk), .Q(n4326), .QN(n1131) );
  DFFX1_HVT \keys_reg[8][38]  ( .D(n2547), .CLK(clk), .Q(n4327), .QN(n1132) );
  DFFX1_HVT \keys_reg[8][37]  ( .D(n2546), .CLK(clk), .Q(n4328), .QN(n1133) );
  DFFX1_HVT \keys_reg[8][36]  ( .D(n2545), .CLK(clk), .Q(n4329), .QN(n1134) );
  DFFX1_HVT \keys_reg[8][35]  ( .D(n2544), .CLK(clk), .Q(n4330), .QN(n1135) );
  DFFX1_HVT \keys_reg[8][34]  ( .D(n2543), .CLK(clk), .Q(n4331), .QN(n1136) );
  DFFX1_HVT \keys_reg[8][33]  ( .D(n2542), .CLK(clk), .Q(n4332), .QN(n1137) );
  DFFX1_HVT \keys_reg[8][32]  ( .D(n2541), .CLK(clk), .Q(n4333), .QN(n1138) );
  DFFX1_HVT \keys_reg[8][31]  ( .D(n2540), .CLK(clk), .Q(n4334), .QN(n1139) );
  DFFX1_HVT \keys_reg[8][30]  ( .D(n2539), .CLK(clk), .Q(n4335), .QN(n1140) );
  DFFX1_HVT \keys_reg[8][29]  ( .D(n2538), .CLK(clk), .Q(n4336), .QN(n1141) );
  DFFX1_HVT \keys_reg[8][28]  ( .D(n2537), .CLK(clk), .Q(n4337), .QN(n1142) );
  DFFX1_HVT \keys_reg[8][27]  ( .D(n2536), .CLK(clk), .Q(n4338), .QN(n1143) );
  DFFX1_HVT \keys_reg[8][26]  ( .D(n2535), .CLK(clk), .Q(n4339), .QN(n1144) );
  DFFX1_HVT \keys_reg[8][25]  ( .D(n2534), .CLK(clk), .Q(n4340), .QN(n1145) );
  DFFX1_HVT \keys_reg[8][24]  ( .D(n2533), .CLK(clk), .Q(n4341), .QN(n1146) );
  DFFX1_HVT \keys_reg[8][23]  ( .D(n2532), .CLK(clk), .Q(n4342), .QN(n1147) );
  DFFX1_HVT \keys_reg[8][22]  ( .D(n2531), .CLK(clk), .Q(n4343), .QN(n1148) );
  DFFX1_HVT \keys_reg[8][21]  ( .D(n2530), .CLK(clk), .Q(n4344), .QN(n1149) );
  DFFX1_HVT \keys_reg[8][20]  ( .D(n2529), .CLK(clk), .Q(n4345), .QN(n1150) );
  DFFX1_HVT \keys_reg[8][19]  ( .D(n2528), .CLK(clk), .Q(n4346), .QN(n1151) );
  DFFX1_HVT \keys_reg[8][18]  ( .D(n2527), .CLK(clk), .Q(n4347), .QN(n1152) );
  DFFX1_HVT \keys_reg[8][17]  ( .D(n2526), .CLK(clk), .Q(n4348), .QN(n1153) );
  DFFX1_HVT \keys_reg[8][16]  ( .D(n2525), .CLK(clk), .Q(n4349), .QN(n1154) );
  DFFX1_HVT \keys_reg[8][15]  ( .D(n2524), .CLK(clk), .Q(n4350), .QN(n1155) );
  DFFX1_HVT \keys_reg[8][14]  ( .D(n2523), .CLK(clk), .Q(n4351), .QN(n1156) );
  DFFX1_HVT \keys_reg[8][13]  ( .D(n2522), .CLK(clk), .Q(n4352), .QN(n1157) );
  DFFX1_HVT \keys_reg[8][12]  ( .D(n2521), .CLK(clk), .Q(n4353), .QN(n1158) );
  DFFX1_HVT \keys_reg[8][11]  ( .D(n2520), .CLK(clk), .Q(n4354), .QN(n1159) );
  DFFX1_HVT \keys_reg[8][10]  ( .D(n2519), .CLK(clk), .Q(n4355), .QN(n1160) );
  DFFX1_HVT \keys_reg[8][9]  ( .D(n2518), .CLK(clk), .Q(n4356), .QN(n1161) );
  DFFX1_HVT \keys_reg[8][8]  ( .D(n2517), .CLK(clk), .Q(n4357), .QN(n1162) );
  DFFX1_HVT \keys_reg[8][7]  ( .D(n2516), .CLK(clk), .Q(n4358), .QN(n1163) );
  DFFX1_HVT \keys_reg[8][6]  ( .D(n2515), .CLK(clk), .Q(n4359), .QN(n1164) );
  DFFX1_HVT \keys_reg[8][5]  ( .D(n2514), .CLK(clk), .Q(n4360), .QN(n1165) );
  DFFX1_HVT \keys_reg[8][4]  ( .D(n2513), .CLK(clk), .Q(n4361), .QN(n1166) );
  DFFX1_HVT \keys_reg[8][3]  ( .D(n2512), .CLK(clk), .Q(n4362), .QN(n1167) );
  DFFX1_HVT \keys_reg[8][2]  ( .D(n2511), .CLK(clk), .Q(n4363), .QN(n1168) );
  DFFX1_HVT \keys_reg[8][1]  ( .D(n2510), .CLK(clk), .Q(n4364), .QN(n1169) );
  DFFX1_HVT \keys_reg[8][0]  ( .D(n2509), .CLK(clk), .Q(n4365), .QN(n1170) );
  DFFX1_HVT \keys_reg[9][127]  ( .D(n2508), .CLK(clk), .Q(n1925), .QN(n1171)
         );
  DFFX1_HVT \keys_reg[9][126]  ( .D(n2507), .CLK(clk), .Q(n1926), .QN(n1172)
         );
  DFFX1_HVT \keys_reg[9][125]  ( .D(n2506), .CLK(clk), .Q(n1927), .QN(n1173)
         );
  DFFX1_HVT \keys_reg[9][124]  ( .D(n2505), .CLK(clk), .Q(n1928), .QN(n1174)
         );
  DFFX1_HVT \keys_reg[9][123]  ( .D(n2504), .CLK(clk), .Q(n1929), .QN(n1175)
         );
  DFFX1_HVT \keys_reg[9][122]  ( .D(n2503), .CLK(clk), .Q(n1930), .QN(n1176)
         );
  DFFX1_HVT \keys_reg[9][121]  ( .D(n2502), .CLK(clk), .Q(n1931), .QN(n1177)
         );
  DFFX1_HVT \keys_reg[9][120]  ( .D(n2501), .CLK(clk), .Q(n1932), .QN(n1178)
         );
  DFFX1_HVT \keys_reg[9][119]  ( .D(n2500), .CLK(clk), .Q(n1933), .QN(n1179)
         );
  DFFX1_HVT \keys_reg[9][118]  ( .D(n2499), .CLK(clk), .Q(n1934), .QN(n1180)
         );
  DFFX1_HVT \keys_reg[9][117]  ( .D(n2498), .CLK(clk), .Q(n1935), .QN(n1181)
         );
  DFFX1_HVT \keys_reg[9][116]  ( .D(n2497), .CLK(clk), .Q(n1936), .QN(n1182)
         );
  DFFX1_HVT \keys_reg[9][115]  ( .D(n2496), .CLK(clk), .Q(n1937), .QN(n1183)
         );
  DFFX1_HVT \keys_reg[9][114]  ( .D(n2495), .CLK(clk), .Q(n1938), .QN(n1184)
         );
  DFFX1_HVT \keys_reg[9][113]  ( .D(n2494), .CLK(clk), .Q(n1939), .QN(n1185)
         );
  DFFX1_HVT \keys_reg[9][112]  ( .D(n2493), .CLK(clk), .Q(n1940), .QN(n1186)
         );
  DFFX1_HVT \keys_reg[9][111]  ( .D(n2492), .CLK(clk), .Q(n1941), .QN(n1187)
         );
  DFFX1_HVT \keys_reg[9][110]  ( .D(n2491), .CLK(clk), .Q(n1942), .QN(n1188)
         );
  DFFX1_HVT \keys_reg[9][109]  ( .D(n2490), .CLK(clk), .Q(n1943), .QN(n1189)
         );
  DFFX1_HVT \keys_reg[9][108]  ( .D(n2489), .CLK(clk), .Q(n1944), .QN(n1190)
         );
  DFFX1_HVT \keys_reg[9][107]  ( .D(n2488), .CLK(clk), .Q(n1945), .QN(n1191)
         );
  DFFX1_HVT \keys_reg[9][106]  ( .D(n2487), .CLK(clk), .Q(n1946), .QN(n1192)
         );
  DFFX1_HVT \keys_reg[9][105]  ( .D(n2486), .CLK(clk), .Q(n1947), .QN(n1193)
         );
  DFFX1_HVT \keys_reg[9][104]  ( .D(n2485), .CLK(clk), .Q(n1948), .QN(n1194)
         );
  DFFX1_HVT \keys_reg[9][103]  ( .D(n2484), .CLK(clk), .Q(n1949), .QN(n1195)
         );
  DFFX1_HVT \keys_reg[9][102]  ( .D(n2483), .CLK(clk), .Q(n1950), .QN(n1196)
         );
  DFFX1_HVT \keys_reg[9][101]  ( .D(n2482), .CLK(clk), .Q(n1951), .QN(n1197)
         );
  DFFX1_HVT \keys_reg[9][100]  ( .D(n2481), .CLK(clk), .Q(n1952), .QN(n1198)
         );
  DFFX1_HVT \keys_reg[9][99]  ( .D(n2480), .CLK(clk), .Q(n1953), .QN(n1199) );
  DFFX1_HVT \keys_reg[9][98]  ( .D(n2479), .CLK(clk), .Q(n1954), .QN(n1200) );
  DFFX1_HVT \keys_reg[9][97]  ( .D(n2478), .CLK(clk), .Q(n1955), .QN(n1201) );
  DFFX1_HVT \keys_reg[9][96]  ( .D(n2477), .CLK(clk), .Q(n1956), .QN(n1202) );
  DFFX1_HVT \keys_reg[9][95]  ( .D(n2476), .CLK(clk), .Q(n1957), .QN(n1203) );
  DFFX1_HVT \keys_reg[9][94]  ( .D(n2475), .CLK(clk), .Q(n1958), .QN(n1204) );
  DFFX1_HVT \keys_reg[9][93]  ( .D(n2474), .CLK(clk), .Q(n1959), .QN(n1205) );
  DFFX1_HVT \keys_reg[9][92]  ( .D(n2473), .CLK(clk), .Q(n1960), .QN(n1206) );
  DFFX1_HVT \keys_reg[9][91]  ( .D(n2472), .CLK(clk), .Q(n1961), .QN(n1207) );
  DFFX1_HVT \keys_reg[9][90]  ( .D(n2471), .CLK(clk), .Q(n1962), .QN(n1208) );
  DFFX1_HVT \keys_reg[9][89]  ( .D(n2470), .CLK(clk), .Q(n1963), .QN(n1209) );
  DFFX1_HVT \keys_reg[9][88]  ( .D(n2469), .CLK(clk), .Q(n1964), .QN(n1210) );
  DFFX1_HVT \keys_reg[9][87]  ( .D(n2468), .CLK(clk), .Q(n1965), .QN(n1211) );
  DFFX1_HVT \keys_reg[9][86]  ( .D(n2467), .CLK(clk), .Q(n1966), .QN(n1212) );
  DFFX1_HVT \keys_reg[9][85]  ( .D(n2466), .CLK(clk), .Q(n1967), .QN(n1213) );
  DFFX1_HVT \keys_reg[9][84]  ( .D(n2465), .CLK(clk), .Q(n1968), .QN(n1214) );
  DFFX1_HVT \keys_reg[9][83]  ( .D(n2464), .CLK(clk), .Q(n1969), .QN(n1215) );
  DFFX1_HVT \keys_reg[9][82]  ( .D(n2463), .CLK(clk), .Q(n1970), .QN(n1216) );
  DFFX1_HVT \keys_reg[9][81]  ( .D(n2462), .CLK(clk), .Q(n1971), .QN(n1217) );
  DFFX1_HVT \keys_reg[9][80]  ( .D(n2461), .CLK(clk), .Q(n1972), .QN(n1218) );
  DFFX1_HVT \keys_reg[9][79]  ( .D(n2460), .CLK(clk), .Q(n1973), .QN(n1219) );
  DFFX1_HVT \keys_reg[9][78]  ( .D(n2459), .CLK(clk), .Q(n1974), .QN(n1220) );
  DFFX1_HVT \keys_reg[9][77]  ( .D(n2458), .CLK(clk), .Q(n1975), .QN(n1221) );
  DFFX1_HVT \keys_reg[9][76]  ( .D(n2457), .CLK(clk), .Q(n1976), .QN(n1222) );
  DFFX1_HVT \keys_reg[9][75]  ( .D(n2456), .CLK(clk), .Q(n1977), .QN(n1223) );
  DFFX1_HVT \keys_reg[9][74]  ( .D(n2455), .CLK(clk), .Q(n1978), .QN(n1224) );
  DFFX1_HVT \keys_reg[9][73]  ( .D(n2454), .CLK(clk), .Q(n1979), .QN(n1225) );
  DFFX1_HVT \keys_reg[9][72]  ( .D(n2453), .CLK(clk), .Q(n1980), .QN(n1226) );
  DFFX1_HVT \keys_reg[9][71]  ( .D(n2452), .CLK(clk), .Q(n1981), .QN(n1227) );
  DFFX1_HVT \keys_reg[9][70]  ( .D(n2451), .CLK(clk), .Q(n1982), .QN(n1228) );
  DFFX1_HVT \keys_reg[9][69]  ( .D(n2450), .CLK(clk), .Q(n1983), .QN(n1229) );
  DFFX1_HVT \keys_reg[9][68]  ( .D(n2449), .CLK(clk), .Q(n1984), .QN(n1230) );
  DFFX1_HVT \keys_reg[9][67]  ( .D(n2448), .CLK(clk), .Q(n1985), .QN(n1231) );
  DFFX1_HVT \keys_reg[9][66]  ( .D(n2447), .CLK(clk), .Q(n1986), .QN(n1232) );
  DFFX1_HVT \keys_reg[9][65]  ( .D(n2446), .CLK(clk), .Q(n1987), .QN(n1233) );
  DFFX1_HVT \keys_reg[9][64]  ( .D(n2445), .CLK(clk), .Q(n1988), .QN(n1234) );
  DFFX1_HVT \keys_reg[9][63]  ( .D(n2444), .CLK(clk), .Q(n1989), .QN(n1235) );
  DFFX1_HVT \keys_reg[9][62]  ( .D(n2443), .CLK(clk), .Q(n1990), .QN(n1236) );
  DFFX1_HVT \keys_reg[9][61]  ( .D(n2442), .CLK(clk), .Q(n1991), .QN(n1237) );
  DFFX1_HVT \keys_reg[9][60]  ( .D(n2441), .CLK(clk), .Q(n1992), .QN(n1238) );
  DFFX1_HVT \keys_reg[9][59]  ( .D(n2440), .CLK(clk), .Q(n1993), .QN(n1239) );
  DFFX1_HVT \keys_reg[9][58]  ( .D(n2439), .CLK(clk), .Q(n1994), .QN(n1240) );
  DFFX1_HVT \keys_reg[9][57]  ( .D(n2438), .CLK(clk), .Q(n1995), .QN(n1241) );
  DFFX1_HVT \keys_reg[9][56]  ( .D(n2437), .CLK(clk), .Q(n1996), .QN(n1242) );
  DFFX1_HVT \keys_reg[9][55]  ( .D(n2436), .CLK(clk), .Q(n1997), .QN(n1243) );
  DFFX1_HVT \keys_reg[9][54]  ( .D(n2435), .CLK(clk), .Q(n1998), .QN(n1244) );
  DFFX1_HVT \keys_reg[9][53]  ( .D(n2434), .CLK(clk), .Q(n1999), .QN(n1245) );
  DFFX1_HVT \keys_reg[9][52]  ( .D(n2433), .CLK(clk), .Q(n2000), .QN(n1246) );
  DFFX1_HVT \keys_reg[9][51]  ( .D(n2432), .CLK(clk), .Q(n2001), .QN(n1247) );
  DFFX1_HVT \keys_reg[9][50]  ( .D(n2431), .CLK(clk), .Q(n2002), .QN(n1248) );
  DFFX1_HVT \keys_reg[9][49]  ( .D(n2430), .CLK(clk), .Q(n2003), .QN(n1249) );
  DFFX1_HVT \keys_reg[9][48]  ( .D(n2429), .CLK(clk), .Q(n2004), .QN(n1250) );
  DFFX1_HVT \keys_reg[9][47]  ( .D(n2428), .CLK(clk), .Q(n2005), .QN(n1251) );
  DFFX1_HVT \keys_reg[9][46]  ( .D(n2427), .CLK(clk), .Q(n2006), .QN(n1252) );
  DFFX1_HVT \keys_reg[9][45]  ( .D(n2426), .CLK(clk), .Q(n2007), .QN(n1253) );
  DFFX1_HVT \keys_reg[9][44]  ( .D(n2425), .CLK(clk), .Q(n2008), .QN(n1254) );
  DFFX1_HVT \keys_reg[9][43]  ( .D(n2424), .CLK(clk), .Q(n2009), .QN(n1255) );
  DFFX1_HVT \keys_reg[9][42]  ( .D(n2423), .CLK(clk), .Q(n2010), .QN(n1256) );
  DFFX1_HVT \keys_reg[9][41]  ( .D(n2422), .CLK(clk), .Q(n2011), .QN(n1257) );
  DFFX1_HVT \keys_reg[9][40]  ( .D(n2421), .CLK(clk), .Q(n2012), .QN(n1258) );
  DFFX1_HVT \keys_reg[9][39]  ( .D(n2420), .CLK(clk), .Q(n2013), .QN(n1259) );
  DFFX1_HVT \keys_reg[9][38]  ( .D(n2419), .CLK(clk), .Q(n2014), .QN(n1260) );
  DFFX1_HVT \keys_reg[9][37]  ( .D(n2418), .CLK(clk), .Q(n2015), .QN(n1261) );
  DFFX1_HVT \keys_reg[9][36]  ( .D(n2417), .CLK(clk), .Q(n2016), .QN(n1262) );
  DFFX1_HVT \keys_reg[9][35]  ( .D(n2416), .CLK(clk), .Q(n2017), .QN(n1263) );
  DFFX1_HVT \keys_reg[9][34]  ( .D(n2415), .CLK(clk), .Q(n2018), .QN(n1264) );
  DFFX1_HVT \keys_reg[9][33]  ( .D(n2414), .CLK(clk), .Q(n2019), .QN(n1265) );
  DFFX1_HVT \keys_reg[9][32]  ( .D(n2413), .CLK(clk), .Q(n2020), .QN(n1266) );
  DFFX1_HVT \keys_reg[9][31]  ( .D(n2412), .CLK(clk), .Q(n2021), .QN(n1267) );
  DFFX1_HVT \keys_reg[9][30]  ( .D(n2411), .CLK(clk), .Q(n2022), .QN(n1268) );
  DFFX1_HVT \keys_reg[9][29]  ( .D(n2410), .CLK(clk), .Q(n2023), .QN(n1269) );
  DFFX1_HVT \keys_reg[9][28]  ( .D(n2409), .CLK(clk), .Q(n2024), .QN(n1270) );
  DFFX1_HVT \keys_reg[9][27]  ( .D(n2408), .CLK(clk), .Q(n2025), .QN(n1271) );
  DFFX1_HVT \keys_reg[9][26]  ( .D(n2407), .CLK(clk), .Q(n2026), .QN(n1272) );
  DFFX1_HVT \keys_reg[9][25]  ( .D(n2406), .CLK(clk), .Q(n2027), .QN(n1273) );
  DFFX1_HVT \keys_reg[9][24]  ( .D(n2405), .CLK(clk), .Q(n2028), .QN(n1274) );
  DFFX1_HVT \keys_reg[9][23]  ( .D(n2404), .CLK(clk), .Q(n2029), .QN(n1275) );
  DFFX1_HVT \keys_reg[9][22]  ( .D(n2403), .CLK(clk), .Q(n2030), .QN(n1276) );
  DFFX1_HVT \keys_reg[9][21]  ( .D(n2402), .CLK(clk), .Q(n2031), .QN(n1277) );
  DFFX1_HVT \keys_reg[9][20]  ( .D(n2401), .CLK(clk), .Q(n2032), .QN(n1278) );
  DFFX1_HVT \keys_reg[9][19]  ( .D(n2400), .CLK(clk), .Q(n2033), .QN(n1279) );
  DFFX1_HVT \keys_reg[9][18]  ( .D(n2399), .CLK(clk), .Q(n2034), .QN(n1280) );
  DFFX1_HVT \keys_reg[9][17]  ( .D(n2398), .CLK(clk), .Q(n2035), .QN(n1281) );
  DFFX1_HVT \keys_reg[9][16]  ( .D(n2397), .CLK(clk), .Q(n2036), .QN(n1282) );
  DFFX1_HVT \keys_reg[9][15]  ( .D(n2396), .CLK(clk), .Q(n2037), .QN(n1283) );
  DFFX1_HVT \keys_reg[9][14]  ( .D(n2395), .CLK(clk), .Q(n2038), .QN(n1284) );
  DFFX1_HVT \keys_reg[9][13]  ( .D(n2394), .CLK(clk), .Q(n2039), .QN(n1285) );
  DFFX1_HVT \keys_reg[9][12]  ( .D(n2393), .CLK(clk), .Q(n2040), .QN(n1286) );
  DFFX1_HVT \keys_reg[9][11]  ( .D(n2392), .CLK(clk), .Q(n2041), .QN(n1287) );
  DFFX1_HVT \keys_reg[9][10]  ( .D(n2391), .CLK(clk), .Q(n2042), .QN(n1288) );
  DFFX1_HVT \keys_reg[9][9]  ( .D(n2390), .CLK(clk), .Q(n2043), .QN(n1289) );
  DFFX1_HVT \keys_reg[9][8]  ( .D(n2389), .CLK(clk), .Q(n2044), .QN(n1290) );
  DFFX1_HVT \keys_reg[9][7]  ( .D(n2388), .CLK(clk), .Q(n2045), .QN(n1291) );
  DFFX1_HVT \keys_reg[9][6]  ( .D(n2387), .CLK(clk), .Q(n2046), .QN(n1292) );
  DFFX1_HVT \keys_reg[9][5]  ( .D(n2386), .CLK(clk), .Q(n2047), .QN(n1293) );
  DFFX1_HVT \keys_reg[9][4]  ( .D(n2385), .CLK(clk), .Q(n2048), .QN(n1294) );
  DFFX1_HVT \keys_reg[9][3]  ( .D(n2384), .CLK(clk), .Q(n2049), .QN(n1295) );
  DFFX1_HVT \keys_reg[9][2]  ( .D(n2383), .CLK(clk), .Q(n2050), .QN(n1296) );
  DFFX1_HVT \keys_reg[9][1]  ( .D(n2382), .CLK(clk), .Q(n2051), .QN(n1297) );
  DFFX1_HVT \keys_reg[9][0]  ( .D(n2381), .CLK(clk), .Q(n2052), .QN(n1298) );
  DFFX1_HVT \keys_reg[10][127]  ( .D(n2380), .CLK(clk), .Q(n1541), .QN(n1299)
         );
  DFFX1_HVT \keys_reg[10][126]  ( .D(n2379), .CLK(clk), .Q(n1542), .QN(n1300)
         );
  DFFX1_HVT \keys_reg[10][125]  ( .D(n2378), .CLK(clk), .Q(n1543), .QN(n1301)
         );
  DFFX1_HVT \keys_reg[10][124]  ( .D(n2377), .CLK(clk), .Q(n1544), .QN(n1302)
         );
  DFFX1_HVT \keys_reg[10][123]  ( .D(n2376), .CLK(clk), .Q(n1545), .QN(n1303)
         );
  DFFX1_HVT \keys_reg[10][122]  ( .D(n2375), .CLK(clk), .Q(n1546), .QN(n1304)
         );
  DFFX1_HVT \keys_reg[10][121]  ( .D(n2374), .CLK(clk), .Q(n1547), .QN(n1305)
         );
  DFFX1_HVT \keys_reg[10][120]  ( .D(n2373), .CLK(clk), .Q(n1548), .QN(n1306)
         );
  DFFX1_HVT \keys_reg[10][119]  ( .D(n2372), .CLK(clk), .Q(n1549), .QN(n1307)
         );
  DFFX1_HVT \keys_reg[10][118]  ( .D(n2371), .CLK(clk), .Q(n1550), .QN(n1308)
         );
  DFFX1_HVT \keys_reg[10][117]  ( .D(n2370), .CLK(clk), .Q(n1551), .QN(n1309)
         );
  DFFX1_HVT \keys_reg[10][116]  ( .D(n2369), .CLK(clk), .Q(n1552), .QN(n1310)
         );
  DFFX1_HVT \keys_reg[10][115]  ( .D(n2368), .CLK(clk), .Q(n1553), .QN(n1311)
         );
  DFFX1_HVT \keys_reg[10][114]  ( .D(n2367), .CLK(clk), .Q(n1554), .QN(n1312)
         );
  DFFX1_HVT \keys_reg[10][113]  ( .D(n2366), .CLK(clk), .Q(n1555), .QN(n1313)
         );
  DFFX1_HVT \keys_reg[10][112]  ( .D(n2365), .CLK(clk), .Q(n1556), .QN(n1314)
         );
  DFFX1_HVT \keys_reg[10][111]  ( .D(n2364), .CLK(clk), .Q(n1557), .QN(n1315)
         );
  DFFX1_HVT \keys_reg[10][110]  ( .D(n2363), .CLK(clk), .Q(n1558), .QN(n1316)
         );
  DFFX1_HVT \keys_reg[10][109]  ( .D(n2362), .CLK(clk), .Q(n1559), .QN(n1317)
         );
  DFFX1_HVT \keys_reg[10][108]  ( .D(n2361), .CLK(clk), .Q(n1560), .QN(n1318)
         );
  DFFX1_HVT \keys_reg[10][107]  ( .D(n2360), .CLK(clk), .Q(n1561), .QN(n1319)
         );
  DFFX1_HVT \keys_reg[10][106]  ( .D(n2359), .CLK(clk), .Q(n1562), .QN(n1320)
         );
  DFFX1_HVT \keys_reg[10][105]  ( .D(n2358), .CLK(clk), .Q(n1563), .QN(n1321)
         );
  DFFX1_HVT \keys_reg[10][104]  ( .D(n2357), .CLK(clk), .Q(n1564), .QN(n1322)
         );
  DFFX1_HVT \keys_reg[10][103]  ( .D(n2356), .CLK(clk), .Q(n1565), .QN(n1323)
         );
  DFFX1_HVT \keys_reg[10][102]  ( .D(n2355), .CLK(clk), .Q(n1566), .QN(n1324)
         );
  DFFX1_HVT \keys_reg[10][101]  ( .D(n2354), .CLK(clk), .Q(n1567), .QN(n1325)
         );
  DFFX1_HVT \keys_reg[10][100]  ( .D(n2353), .CLK(clk), .Q(n1568), .QN(n1326)
         );
  DFFX1_HVT \keys_reg[10][99]  ( .D(n2352), .CLK(clk), .Q(n1569), .QN(n1327)
         );
  DFFX1_HVT \keys_reg[10][98]  ( .D(n2351), .CLK(clk), .Q(n1570), .QN(n1328)
         );
  DFFX1_HVT \keys_reg[10][97]  ( .D(n2350), .CLK(clk), .Q(n1571), .QN(n1329)
         );
  DFFX1_HVT \keys_reg[10][96]  ( .D(n2349), .CLK(clk), .Q(n1572), .QN(n1330)
         );
  DFFX1_HVT \keys_reg[10][95]  ( .D(n2348), .CLK(clk), .Q(n1573), .QN(n1331)
         );
  DFFX1_HVT \keys_reg[10][94]  ( .D(n2347), .CLK(clk), .Q(n1574), .QN(n1332)
         );
  DFFX1_HVT \keys_reg[10][93]  ( .D(n2346), .CLK(clk), .Q(n1575), .QN(n1333)
         );
  DFFX1_HVT \keys_reg[10][92]  ( .D(n2345), .CLK(clk), .Q(n1576), .QN(n1334)
         );
  DFFX1_HVT \keys_reg[10][91]  ( .D(n2344), .CLK(clk), .Q(n1577), .QN(n1335)
         );
  DFFX1_HVT \keys_reg[10][90]  ( .D(n2343), .CLK(clk), .Q(n1578), .QN(n1336)
         );
  DFFX1_HVT \keys_reg[10][89]  ( .D(n2342), .CLK(clk), .Q(n1579), .QN(n1337)
         );
  DFFX1_HVT \keys_reg[10][88]  ( .D(n2341), .CLK(clk), .Q(n1580), .QN(n1338)
         );
  DFFX1_HVT \keys_reg[10][87]  ( .D(n2340), .CLK(clk), .Q(n1581), .QN(n1339)
         );
  DFFX1_HVT \keys_reg[10][86]  ( .D(n2339), .CLK(clk), .Q(n1582), .QN(n1340)
         );
  DFFX1_HVT \keys_reg[10][85]  ( .D(n2338), .CLK(clk), .Q(n1583), .QN(n1341)
         );
  DFFX1_HVT \keys_reg[10][84]  ( .D(n2337), .CLK(clk), .Q(n1584), .QN(n1342)
         );
  DFFX1_HVT \keys_reg[10][83]  ( .D(n2336), .CLK(clk), .Q(n1585), .QN(n1343)
         );
  DFFX1_HVT \keys_reg[10][82]  ( .D(n2335), .CLK(clk), .Q(n1586), .QN(n1344)
         );
  DFFX1_HVT \keys_reg[10][81]  ( .D(n2334), .CLK(clk), .Q(n1587), .QN(n1345)
         );
  DFFX1_HVT \keys_reg[10][80]  ( .D(n2333), .CLK(clk), .Q(n1588), .QN(n1346)
         );
  DFFX1_HVT \keys_reg[10][79]  ( .D(n2332), .CLK(clk), .Q(n1589), .QN(n1347)
         );
  DFFX1_HVT \keys_reg[10][78]  ( .D(n2331), .CLK(clk), .Q(n1590), .QN(n1348)
         );
  DFFX1_HVT \keys_reg[10][77]  ( .D(n2330), .CLK(clk), .Q(n1591), .QN(n1349)
         );
  DFFX1_HVT \keys_reg[10][76]  ( .D(n2329), .CLK(clk), .Q(n1592), .QN(n1350)
         );
  DFFX1_HVT \keys_reg[10][75]  ( .D(n2328), .CLK(clk), .Q(n1593), .QN(n1351)
         );
  DFFX1_HVT \keys_reg[10][74]  ( .D(n2327), .CLK(clk), .Q(n1594), .QN(n1352)
         );
  DFFX1_HVT \keys_reg[10][73]  ( .D(n2326), .CLK(clk), .Q(n1595), .QN(n1353)
         );
  DFFX1_HVT \keys_reg[10][72]  ( .D(n2325), .CLK(clk), .Q(n1596), .QN(n1354)
         );
  DFFX1_HVT \keys_reg[10][71]  ( .D(n2324), .CLK(clk), .Q(n1597), .QN(n1355)
         );
  DFFX1_HVT \keys_reg[10][70]  ( .D(n2323), .CLK(clk), .Q(n1598), .QN(n1356)
         );
  DFFX1_HVT \keys_reg[10][69]  ( .D(n2322), .CLK(clk), .Q(n1599), .QN(n1357)
         );
  DFFX1_HVT \keys_reg[10][68]  ( .D(n2321), .CLK(clk), .Q(n1600), .QN(n1358)
         );
  DFFX1_HVT \keys_reg[10][67]  ( .D(n2320), .CLK(clk), .Q(n1601), .QN(n1359)
         );
  DFFX1_HVT \keys_reg[10][66]  ( .D(n2319), .CLK(clk), .Q(n1602), .QN(n1360)
         );
  DFFX1_HVT \keys_reg[10][65]  ( .D(n2318), .CLK(clk), .Q(n1603), .QN(n1361)
         );
  DFFX1_HVT \keys_reg[10][64]  ( .D(n2317), .CLK(clk), .Q(n1604), .QN(n1362)
         );
  DFFX1_HVT \keys_reg[10][63]  ( .D(n2316), .CLK(clk), .Q(n1605), .QN(n1363)
         );
  DFFX1_HVT \keys_reg[10][62]  ( .D(n2315), .CLK(clk), .Q(n1606), .QN(n1364)
         );
  DFFX1_HVT \keys_reg[10][61]  ( .D(n2314), .CLK(clk), .Q(n1607), .QN(n1365)
         );
  DFFX1_HVT \keys_reg[10][60]  ( .D(n2313), .CLK(clk), .Q(n1608), .QN(n1366)
         );
  DFFX1_HVT \keys_reg[10][59]  ( .D(n2312), .CLK(clk), .Q(n1609), .QN(n1367)
         );
  DFFX1_HVT \keys_reg[10][58]  ( .D(n2311), .CLK(clk), .Q(n1610), .QN(n1368)
         );
  DFFX1_HVT \keys_reg[10][57]  ( .D(n2310), .CLK(clk), .Q(n1611), .QN(n1369)
         );
  DFFX1_HVT \keys_reg[10][56]  ( .D(n2309), .CLK(clk), .Q(n1612), .QN(n1370)
         );
  DFFX1_HVT \keys_reg[10][55]  ( .D(n2308), .CLK(clk), .Q(n1613), .QN(n1371)
         );
  DFFX1_HVT \keys_reg[10][54]  ( .D(n2307), .CLK(clk), .Q(n1614), .QN(n1372)
         );
  DFFX1_HVT \keys_reg[10][53]  ( .D(n2306), .CLK(clk), .Q(n1615), .QN(n1373)
         );
  DFFX1_HVT \keys_reg[10][52]  ( .D(n2305), .CLK(clk), .Q(n1616), .QN(n1374)
         );
  DFFX1_HVT \keys_reg[10][51]  ( .D(n2304), .CLK(clk), .Q(n1617), .QN(n1375)
         );
  DFFX1_HVT \keys_reg[10][50]  ( .D(n2303), .CLK(clk), .Q(n1618), .QN(n1376)
         );
  DFFX1_HVT \keys_reg[10][49]  ( .D(n2302), .CLK(clk), .Q(n1619), .QN(n1377)
         );
  DFFX1_HVT \keys_reg[10][48]  ( .D(n2301), .CLK(clk), .Q(n1620), .QN(n1378)
         );
  DFFX1_HVT \keys_reg[10][47]  ( .D(n2300), .CLK(clk), .Q(n1621), .QN(n1379)
         );
  DFFX1_HVT \keys_reg[10][46]  ( .D(n2299), .CLK(clk), .Q(n1622), .QN(n1380)
         );
  DFFX1_HVT \keys_reg[10][45]  ( .D(n2298), .CLK(clk), .Q(n1623), .QN(n1381)
         );
  DFFX1_HVT \keys_reg[10][44]  ( .D(n2297), .CLK(clk), .Q(n1624), .QN(n1382)
         );
  DFFX1_HVT \keys_reg[10][43]  ( .D(n2296), .CLK(clk), .Q(n1625), .QN(n1383)
         );
  DFFX1_HVT \keys_reg[10][42]  ( .D(n2295), .CLK(clk), .Q(n1626), .QN(n1384)
         );
  DFFX1_HVT \keys_reg[10][41]  ( .D(n2294), .CLK(clk), .Q(n1627), .QN(n1385)
         );
  DFFX1_HVT \keys_reg[10][40]  ( .D(n2293), .CLK(clk), .Q(n1628), .QN(n1386)
         );
  DFFX1_HVT \keys_reg[10][39]  ( .D(n2292), .CLK(clk), .Q(n1629), .QN(n1387)
         );
  DFFX1_HVT \keys_reg[10][38]  ( .D(n2291), .CLK(clk), .Q(n1630), .QN(n1388)
         );
  DFFX1_HVT \keys_reg[10][37]  ( .D(n2290), .CLK(clk), .Q(n1631), .QN(n1389)
         );
  DFFX1_HVT \keys_reg[10][36]  ( .D(n2289), .CLK(clk), .Q(n1632), .QN(n1390)
         );
  DFFX1_HVT \keys_reg[10][35]  ( .D(n2288), .CLK(clk), .Q(n1633), .QN(n1391)
         );
  DFFX1_HVT \keys_reg[10][34]  ( .D(n2287), .CLK(clk), .Q(n1634), .QN(n1392)
         );
  DFFX1_HVT \keys_reg[10][33]  ( .D(n2286), .CLK(clk), .Q(n1635), .QN(n1393)
         );
  DFFX1_HVT \keys_reg[10][32]  ( .D(n2285), .CLK(clk), .Q(n1636), .QN(n1394)
         );
  DFFX1_HVT \keys_reg[10][31]  ( .D(n2284), .CLK(clk), .Q(n1637), .QN(n1395)
         );
  DFFX1_HVT \keys_reg[10][30]  ( .D(n2283), .CLK(clk), .Q(n1638), .QN(n1396)
         );
  DFFX1_HVT \keys_reg[10][29]  ( .D(n2282), .CLK(clk), .Q(n1639), .QN(n1397)
         );
  DFFX1_HVT \keys_reg[10][28]  ( .D(n2281), .CLK(clk), .Q(n1640), .QN(n1398)
         );
  DFFX1_HVT \keys_reg[10][27]  ( .D(n2280), .CLK(clk), .Q(n1641), .QN(n1399)
         );
  DFFX1_HVT \keys_reg[10][26]  ( .D(n2279), .CLK(clk), .Q(n1642), .QN(n1400)
         );
  DFFX1_HVT \keys_reg[10][25]  ( .D(n2278), .CLK(clk), .Q(n1643), .QN(n1401)
         );
  DFFX1_HVT \keys_reg[10][24]  ( .D(n2277), .CLK(clk), .Q(n1644), .QN(n1402)
         );
  DFFX1_HVT \keys_reg[10][23]  ( .D(n2276), .CLK(clk), .Q(n1645), .QN(n1403)
         );
  DFFX1_HVT \keys_reg[10][22]  ( .D(n2275), .CLK(clk), .Q(n1646), .QN(n1404)
         );
  DFFX1_HVT \keys_reg[10][21]  ( .D(n2274), .CLK(clk), .Q(n1647), .QN(n1405)
         );
  DFFX1_HVT \keys_reg[10][20]  ( .D(n2273), .CLK(clk), .Q(n1648), .QN(n1406)
         );
  DFFX1_HVT \keys_reg[10][19]  ( .D(n2272), .CLK(clk), .Q(n1649), .QN(n1407)
         );
  DFFX1_HVT \keys_reg[10][18]  ( .D(n2271), .CLK(clk), .Q(n1650), .QN(n1408)
         );
  DFFX1_HVT \keys_reg[10][17]  ( .D(n2270), .CLK(clk), .Q(n1651), .QN(n1409)
         );
  DFFX1_HVT \keys_reg[10][16]  ( .D(n2269), .CLK(clk), .Q(n1652), .QN(n1410)
         );
  DFFX1_HVT \keys_reg[10][15]  ( .D(n2268), .CLK(clk), .Q(n1653), .QN(n1411)
         );
  DFFX1_HVT \keys_reg[10][14]  ( .D(n2267), .CLK(clk), .Q(n1654), .QN(n1412)
         );
  DFFX1_HVT \keys_reg[10][13]  ( .D(n2266), .CLK(clk), .Q(n1655), .QN(n1413)
         );
  DFFX1_HVT \keys_reg[10][12]  ( .D(n2265), .CLK(clk), .Q(n1656), .QN(n1414)
         );
  DFFX1_HVT \keys_reg[10][11]  ( .D(n2264), .CLK(clk), .Q(n1657), .QN(n1415)
         );
  DFFX1_HVT \keys_reg[10][10]  ( .D(n2263), .CLK(clk), .Q(n1658), .QN(n1416)
         );
  DFFX1_HVT \keys_reg[10][9]  ( .D(n2262), .CLK(clk), .Q(n1659), .QN(n1417) );
  DFFX1_HVT \keys_reg[10][8]  ( .D(n2261), .CLK(clk), .Q(n1660), .QN(n1418) );
  DFFX1_HVT \keys_reg[10][7]  ( .D(n2260), .CLK(clk), .Q(n1661), .QN(n1419) );
  DFFX1_HVT \keys_reg[10][6]  ( .D(n2259), .CLK(clk), .Q(n1662), .QN(n1420) );
  DFFX1_HVT \keys_reg[10][5]  ( .D(n2258), .CLK(clk), .Q(n1663), .QN(n1421) );
  DFFX1_HVT \keys_reg[10][4]  ( .D(n2257), .CLK(clk), .Q(n1664), .QN(n1422) );
  DFFX1_HVT \keys_reg[10][3]  ( .D(n2256), .CLK(clk), .Q(n1665), .QN(n1423) );
  DFFX1_HVT \keys_reg[10][2]  ( .D(n2255), .CLK(clk), .Q(n1666), .QN(n1424) );
  DFFX1_HVT \keys_reg[10][1]  ( .D(n2254), .CLK(clk), .Q(n1667), .QN(n1425) );
  DFFX1_HVT \keys_reg[10][0]  ( .D(n2253), .CLK(clk), .Q(n1668), .QN(n1426) );
  DFFX1_HVT \key_round_reg[127]  ( .D(n2252), .CLK(clk), .Q(key_round[127]) );
  DFFX1_HVT \key_round_reg[126]  ( .D(n2251), .CLK(clk), .Q(key_round[126]) );
  DFFX1_HVT \key_round_reg[125]  ( .D(n2250), .CLK(clk), .Q(key_round[125]) );
  DFFX1_HVT \key_round_reg[124]  ( .D(n2249), .CLK(clk), .Q(key_round[124]) );
  DFFX1_HVT \key_round_reg[123]  ( .D(n2248), .CLK(clk), .Q(key_round[123]) );
  DFFX1_HVT \key_round_reg[122]  ( .D(n2247), .CLK(clk), .Q(key_round[122]) );
  DFFX1_HVT \key_round_reg[121]  ( .D(n2246), .CLK(clk), .Q(key_round[121]) );
  DFFX1_HVT \key_round_reg[120]  ( .D(n2245), .CLK(clk), .Q(key_round[120]) );
  DFFX1_HVT \key_round_reg[119]  ( .D(n2244), .CLK(clk), .Q(key_round[119]) );
  DFFX1_HVT \key_round_reg[118]  ( .D(n2243), .CLK(clk), .Q(key_round[118]) );
  DFFX1_HVT \key_round_reg[117]  ( .D(n2242), .CLK(clk), .Q(key_round[117]) );
  DFFX1_HVT \key_round_reg[116]  ( .D(n2241), .CLK(clk), .Q(key_round[116]) );
  DFFX1_HVT \key_round_reg[115]  ( .D(n2240), .CLK(clk), .Q(key_round[115]) );
  DFFX1_HVT \key_round_reg[114]  ( .D(n2239), .CLK(clk), .Q(key_round[114]) );
  DFFX1_HVT \key_round_reg[113]  ( .D(n2238), .CLK(clk), .Q(key_round[113]) );
  DFFX1_HVT \key_round_reg[112]  ( .D(n2237), .CLK(clk), .Q(key_round[112]) );
  DFFX1_HVT \key_round_reg[111]  ( .D(n2236), .CLK(clk), .Q(key_round[111]) );
  DFFX1_HVT \key_round_reg[110]  ( .D(n2235), .CLK(clk), .Q(key_round[110]) );
  DFFX1_HVT \key_round_reg[109]  ( .D(n2234), .CLK(clk), .Q(key_round[109]) );
  DFFX1_HVT \key_round_reg[108]  ( .D(n2233), .CLK(clk), .Q(key_round[108]) );
  DFFX1_HVT \key_round_reg[107]  ( .D(n2232), .CLK(clk), .Q(key_round[107]) );
  DFFX1_HVT \key_round_reg[106]  ( .D(n2231), .CLK(clk), .Q(key_round[106]) );
  DFFX1_HVT \key_round_reg[105]  ( .D(n2230), .CLK(clk), .Q(key_round[105]) );
  DFFX1_HVT \key_round_reg[104]  ( .D(n2229), .CLK(clk), .Q(key_round[104]) );
  DFFX1_HVT \key_round_reg[103]  ( .D(n2228), .CLK(clk), .Q(key_round[103]) );
  DFFX1_HVT \key_round_reg[102]  ( .D(n2227), .CLK(clk), .Q(key_round[102]) );
  DFFX1_HVT \key_round_reg[101]  ( .D(n2226), .CLK(clk), .Q(key_round[101]) );
  DFFX1_HVT \key_round_reg[100]  ( .D(n2225), .CLK(clk), .Q(key_round[100]) );
  DFFX1_HVT \key_round_reg[99]  ( .D(n2224), .CLK(clk), .Q(key_round[99]) );
  DFFX1_HVT \key_round_reg[98]  ( .D(n2223), .CLK(clk), .Q(key_round[98]) );
  DFFX1_HVT \key_round_reg[97]  ( .D(n2222), .CLK(clk), .Q(key_round[97]) );
  DFFX1_HVT \key_round_reg[96]  ( .D(n2221), .CLK(clk), .Q(key_round[96]) );
  DFFX1_HVT \key_round_reg[95]  ( .D(n2220), .CLK(clk), .Q(key_round[95]) );
  DFFX1_HVT \key_round_reg[94]  ( .D(n2219), .CLK(clk), .Q(key_round[94]) );
  DFFX1_HVT \key_round_reg[93]  ( .D(n2218), .CLK(clk), .Q(key_round[93]) );
  DFFX1_HVT \key_round_reg[92]  ( .D(n2217), .CLK(clk), .Q(key_round[92]) );
  DFFX1_HVT \key_round_reg[91]  ( .D(n2216), .CLK(clk), .Q(key_round[91]) );
  DFFX1_HVT \key_round_reg[90]  ( .D(n2215), .CLK(clk), .Q(key_round[90]) );
  DFFX1_HVT \key_round_reg[89]  ( .D(n2214), .CLK(clk), .Q(key_round[89]) );
  DFFX1_HVT \key_round_reg[88]  ( .D(n2213), .CLK(clk), .Q(key_round[88]) );
  DFFX1_HVT \key_round_reg[87]  ( .D(n2212), .CLK(clk), .Q(key_round[87]) );
  DFFX1_HVT \key_round_reg[86]  ( .D(n2211), .CLK(clk), .Q(key_round[86]) );
  DFFX1_HVT \key_round_reg[85]  ( .D(n2210), .CLK(clk), .Q(key_round[85]) );
  DFFX1_HVT \key_round_reg[84]  ( .D(n2209), .CLK(clk), .Q(key_round[84]) );
  DFFX1_HVT \key_round_reg[83]  ( .D(n2208), .CLK(clk), .Q(key_round[83]) );
  DFFX1_HVT \key_round_reg[82]  ( .D(n2207), .CLK(clk), .Q(key_round[82]) );
  DFFX1_HVT \key_round_reg[81]  ( .D(n2206), .CLK(clk), .Q(key_round[81]) );
  DFFX1_HVT \key_round_reg[80]  ( .D(n2205), .CLK(clk), .Q(key_round[80]) );
  DFFX1_HVT \key_round_reg[79]  ( .D(n2204), .CLK(clk), .Q(key_round[79]) );
  DFFX1_HVT \key_round_reg[78]  ( .D(n2203), .CLK(clk), .Q(key_round[78]) );
  DFFX1_HVT \key_round_reg[77]  ( .D(n2202), .CLK(clk), .Q(key_round[77]) );
  DFFX1_HVT \key_round_reg[76]  ( .D(n2201), .CLK(clk), .Q(key_round[76]) );
  DFFX1_HVT \key_round_reg[75]  ( .D(n2200), .CLK(clk), .Q(key_round[75]) );
  DFFX1_HVT \key_round_reg[74]  ( .D(n2199), .CLK(clk), .Q(key_round[74]) );
  DFFX1_HVT \key_round_reg[73]  ( .D(n2198), .CLK(clk), .Q(key_round[73]) );
  DFFX1_HVT \key_round_reg[72]  ( .D(n2197), .CLK(clk), .Q(key_round[72]) );
  DFFX1_HVT \key_round_reg[71]  ( .D(n2196), .CLK(clk), .Q(key_round[71]) );
  DFFX1_HVT \key_round_reg[70]  ( .D(n2195), .CLK(clk), .Q(key_round[70]) );
  DFFX1_HVT \key_round_reg[69]  ( .D(n2194), .CLK(clk), .Q(key_round[69]) );
  DFFX1_HVT \key_round_reg[68]  ( .D(n2193), .CLK(clk), .Q(key_round[68]) );
  DFFX1_HVT \key_round_reg[67]  ( .D(n2192), .CLK(clk), .Q(key_round[67]) );
  DFFX1_HVT \key_round_reg[66]  ( .D(n2191), .CLK(clk), .Q(key_round[66]) );
  DFFX1_HVT \key_round_reg[65]  ( .D(n2190), .CLK(clk), .Q(key_round[65]) );
  DFFX1_HVT \key_round_reg[64]  ( .D(n2189), .CLK(clk), .Q(key_round[64]) );
  DFFX1_HVT \key_round_reg[63]  ( .D(n2188), .CLK(clk), .Q(key_round[63]) );
  DFFX1_HVT \key_round_reg[62]  ( .D(n2187), .CLK(clk), .Q(key_round[62]) );
  DFFX1_HVT \key_round_reg[61]  ( .D(n2186), .CLK(clk), .Q(key_round[61]) );
  DFFX1_HVT \key_round_reg[60]  ( .D(n2185), .CLK(clk), .Q(key_round[60]) );
  DFFX1_HVT \key_round_reg[59]  ( .D(n2184), .CLK(clk), .Q(key_round[59]) );
  DFFX1_HVT \key_round_reg[58]  ( .D(n2183), .CLK(clk), .Q(key_round[58]) );
  DFFX1_HVT \key_round_reg[57]  ( .D(n2182), .CLK(clk), .Q(key_round[57]) );
  DFFX1_HVT \key_round_reg[56]  ( .D(n2181), .CLK(clk), .Q(key_round[56]) );
  DFFX1_HVT \key_round_reg[55]  ( .D(n2180), .CLK(clk), .Q(key_round[55]) );
  DFFX1_HVT \key_round_reg[54]  ( .D(n2179), .CLK(clk), .Q(key_round[54]) );
  DFFX1_HVT \key_round_reg[53]  ( .D(n2178), .CLK(clk), .Q(key_round[53]) );
  DFFX1_HVT \key_round_reg[52]  ( .D(n2177), .CLK(clk), .Q(key_round[52]) );
  DFFX1_HVT \key_round_reg[51]  ( .D(n2176), .CLK(clk), .Q(key_round[51]) );
  DFFX1_HVT \key_round_reg[50]  ( .D(n2175), .CLK(clk), .Q(key_round[50]) );
  DFFX1_HVT \key_round_reg[49]  ( .D(n2174), .CLK(clk), .Q(key_round[49]) );
  DFFX1_HVT \key_round_reg[48]  ( .D(n2173), .CLK(clk), .Q(key_round[48]) );
  DFFX1_HVT \key_round_reg[47]  ( .D(n2172), .CLK(clk), .Q(key_round[47]) );
  DFFX1_HVT \key_round_reg[46]  ( .D(n2171), .CLK(clk), .Q(key_round[46]) );
  DFFX1_HVT \key_round_reg[45]  ( .D(n2170), .CLK(clk), .Q(key_round[45]) );
  DFFX1_HVT \key_round_reg[44]  ( .D(n2169), .CLK(clk), .Q(key_round[44]) );
  DFFX1_HVT \key_round_reg[43]  ( .D(n2168), .CLK(clk), .Q(key_round[43]) );
  DFFX1_HVT \key_round_reg[42]  ( .D(n2167), .CLK(clk), .Q(key_round[42]) );
  DFFX1_HVT \key_round_reg[41]  ( .D(n2166), .CLK(clk), .Q(key_round[41]) );
  DFFX1_HVT \key_round_reg[40]  ( .D(n2165), .CLK(clk), .Q(key_round[40]) );
  DFFX1_HVT \key_round_reg[39]  ( .D(n2164), .CLK(clk), .Q(key_round[39]) );
  DFFX1_HVT \key_round_reg[38]  ( .D(n2163), .CLK(clk), .Q(key_round[38]) );
  DFFX1_HVT \key_round_reg[37]  ( .D(n2162), .CLK(clk), .Q(key_round[37]) );
  DFFX1_HVT \key_round_reg[36]  ( .D(n2161), .CLK(clk), .Q(key_round[36]) );
  DFFX1_HVT \key_round_reg[35]  ( .D(n2160), .CLK(clk), .Q(key_round[35]) );
  DFFX1_HVT \key_round_reg[34]  ( .D(n2159), .CLK(clk), .Q(key_round[34]) );
  DFFX1_HVT \key_round_reg[33]  ( .D(n2158), .CLK(clk), .Q(key_round[33]) );
  DFFX1_HVT \key_round_reg[32]  ( .D(n2157), .CLK(clk), .Q(key_round[32]) );
  DFFX1_HVT \key_round_reg[31]  ( .D(n2156), .CLK(clk), .Q(key_round[31]) );
  DFFX1_HVT \key_round_reg[30]  ( .D(n2155), .CLK(clk), .Q(key_round[30]) );
  DFFX1_HVT \key_round_reg[29]  ( .D(n2154), .CLK(clk), .Q(key_round[29]) );
  DFFX1_HVT \key_round_reg[28]  ( .D(n2153), .CLK(clk), .Q(key_round[28]) );
  DFFX1_HVT \key_round_reg[27]  ( .D(n2152), .CLK(clk), .Q(key_round[27]) );
  DFFX1_HVT \key_round_reg[26]  ( .D(n2151), .CLK(clk), .Q(key_round[26]) );
  DFFX1_HVT \key_round_reg[25]  ( .D(n2150), .CLK(clk), .Q(key_round[25]) );
  DFFX1_HVT \key_round_reg[24]  ( .D(n2149), .CLK(clk), .Q(key_round[24]) );
  DFFX1_HVT \key_round_reg[23]  ( .D(n2148), .CLK(clk), .Q(key_round[23]) );
  DFFX1_HVT \key_round_reg[22]  ( .D(n2147), .CLK(clk), .Q(key_round[22]) );
  DFFX1_HVT \key_round_reg[21]  ( .D(n2146), .CLK(clk), .Q(key_round[21]) );
  DFFX1_HVT \key_round_reg[20]  ( .D(n2145), .CLK(clk), .Q(key_round[20]) );
  DFFX1_HVT \key_round_reg[19]  ( .D(n2144), .CLK(clk), .Q(key_round[19]) );
  DFFX1_HVT \key_round_reg[18]  ( .D(n2143), .CLK(clk), .Q(key_round[18]) );
  DFFX1_HVT \key_round_reg[17]  ( .D(n2142), .CLK(clk), .Q(key_round[17]) );
  DFFX1_HVT \key_round_reg[16]  ( .D(n2141), .CLK(clk), .Q(key_round[16]) );
  DFFX1_HVT \key_round_reg[15]  ( .D(n2140), .CLK(clk), .Q(key_round[15]) );
  DFFX1_HVT \key_round_reg[14]  ( .D(n2139), .CLK(clk), .Q(key_round[14]) );
  DFFX1_HVT \key_round_reg[13]  ( .D(n2138), .CLK(clk), .Q(key_round[13]) );
  DFFX1_HVT \key_round_reg[12]  ( .D(n2137), .CLK(clk), .Q(key_round[12]) );
  DFFX1_HVT \key_round_reg[11]  ( .D(n2136), .CLK(clk), .Q(key_round[11]) );
  DFFX1_HVT \key_round_reg[10]  ( .D(n2135), .CLK(clk), .Q(key_round[10]) );
  DFFX1_HVT \key_round_reg[9]  ( .D(n2134), .CLK(clk), .Q(key_round[9]) );
  DFFX1_HVT \key_round_reg[8]  ( .D(n2133), .CLK(clk), .Q(key_round[8]) );
  DFFX1_HVT \key_round_reg[7]  ( .D(n2132), .CLK(clk), .Q(key_round[7]) );
  DFFX1_HVT \key_round_reg[6]  ( .D(n2131), .CLK(clk), .Q(key_round[6]) );
  DFFX1_HVT \key_round_reg[5]  ( .D(n2130), .CLK(clk), .Q(key_round[5]) );
  DFFX1_HVT \key_round_reg[4]  ( .D(n2129), .CLK(clk), .Q(key_round[4]) );
  DFFX1_HVT \key_round_reg[3]  ( .D(n2128), .CLK(clk), .Q(key_round[3]) );
  DFFX1_HVT \key_round_reg[2]  ( .D(n2127), .CLK(clk), .Q(key_round[2]) );
  DFFX1_HVT \key_round_reg[1]  ( .D(n2126), .CLK(clk), .Q(key_round[1]) );
  DFFX1_HVT \key_round_reg[0]  ( .D(n2125), .CLK(clk), .Q(key_round[0]) );
  keygen_1 key ( .round_num(round_number), .keyin(prev_key), .keyout(keyout)
         );
  NAND4X1_HVT U3 ( .A1(n4494), .A2(n4495), .A3(n4496), .A4(n4497), .Y(n3797)
         );
  AND3X2_HVT U4 ( .A1(n4506), .A2(n4499), .A3(n4507), .Y(n4494) );
  NAND4X1_HVT U5 ( .A1(n4499), .A2(n4497), .A3(n4500), .A4(n4501), .Y(n3796)
         );
  NAND4X1_HVT U6 ( .A1(n4506), .A2(n4496), .A3(n4503), .A4(n4508), .Y(n3794)
         );
  NAND4X1_HVT U7 ( .A1(n4503), .A2(n4500), .A3(n4504), .A4(n4505), .Y(n3795)
         );
  OR2X1_HVT U8 ( .A1(n4498), .A2(n1), .Y(n4495) );
  OA21X1_HVT U9 ( .A1(n4), .A2(n4498), .A3(n4502), .Y(n4501) );
  OA21X1_HVT U10 ( .A1(n3), .A2(n4498), .A3(n4494), .Y(n4505) );
  OA21X1_HVT U11 ( .A1(n2), .A2(n4498), .A3(n4509), .Y(n4508) );
  OR2X1_HVT U12 ( .A1(n4510), .A2(rest), .Y(n4498) );
  AO21X1_HVT U13 ( .A1(done), .A2(n4511), .A3(n4512), .Y(n3793) );
  OR2X1_HVT U14 ( .A1(n4513), .A2(n4514), .Y(n3792) );
  MUX21X1_HVT U15 ( .A1(round_number[0]), .A2(n4515), .S0(n4516), .Y(n4514) );
  NAND3X0_HVT U16 ( .A1(n4517), .A2(n4518), .A3(n4519), .Y(n4515) );
  MUX21X1_HVT U17 ( .A1(round_number[1]), .A2(n4520), .S0(n4516), .Y(n3791) );
  MUX21X1_HVT U18 ( .A1(round_number[2]), .A2(n4521), .S0(n4516), .Y(n3790) );
  NAND3X0_HVT U19 ( .A1(n4522), .A2(n4523), .A3(n4519), .Y(n4521) );
  AND2X1_HVT U20 ( .A1(n4524), .A2(n4525), .Y(n4519) );
  MUX21X1_HVT U21 ( .A1(round_number[3]), .A2(n4526), .S0(n4516), .Y(n3789) );
  NAND2X0_HVT U22 ( .A1(n4527), .A2(n4528), .Y(n4526) );
  AO222X1_HVT U23 ( .A1(local_key[0]), .A2(n4513), .A3(keyout[0]), .A4(n4529), 
        .A5(prev_key[0]), .A6(n4530), .Y(n3788) );
  AO222X1_HVT U24 ( .A1(local_key[1]), .A2(n4513), .A3(keyout[1]), .A4(n4529), 
        .A5(prev_key[1]), .A6(n4530), .Y(n3787) );
  AO222X1_HVT U25 ( .A1(local_key[2]), .A2(n4513), .A3(keyout[2]), .A4(n4529), 
        .A5(prev_key[2]), .A6(n4530), .Y(n3786) );
  AO222X1_HVT U26 ( .A1(local_key[3]), .A2(n4513), .A3(keyout[3]), .A4(n4529), 
        .A5(prev_key[3]), .A6(n4530), .Y(n3785) );
  AO222X1_HVT U27 ( .A1(local_key[4]), .A2(n4513), .A3(keyout[4]), .A4(n4529), 
        .A5(prev_key[4]), .A6(n4530), .Y(n3784) );
  AO222X1_HVT U28 ( .A1(local_key[5]), .A2(n4513), .A3(keyout[5]), .A4(n4529), 
        .A5(prev_key[5]), .A6(n4530), .Y(n3783) );
  AO222X1_HVT U29 ( .A1(local_key[6]), .A2(n4513), .A3(keyout[6]), .A4(n4529), 
        .A5(prev_key[6]), .A6(n4530), .Y(n3782) );
  AO222X1_HVT U30 ( .A1(local_key[7]), .A2(n4513), .A3(keyout[7]), .A4(n4529), 
        .A5(prev_key[7]), .A6(n4530), .Y(n3781) );
  AO222X1_HVT U31 ( .A1(local_key[8]), .A2(n4513), .A3(keyout[8]), .A4(n4529), 
        .A5(prev_key[8]), .A6(n4530), .Y(n3780) );
  AO222X1_HVT U32 ( .A1(local_key[9]), .A2(n4513), .A3(keyout[9]), .A4(n4529), 
        .A5(prev_key[9]), .A6(n4530), .Y(n3779) );
  AO222X1_HVT U33 ( .A1(local_key[10]), .A2(n4513), .A3(keyout[10]), .A4(n4529), .A5(prev_key[10]), .A6(n4530), .Y(n3778) );
  AO222X1_HVT U34 ( .A1(local_key[11]), .A2(n4513), .A3(keyout[11]), .A4(n4529), .A5(prev_key[11]), .A6(n4530), .Y(n3777) );
  AO222X1_HVT U35 ( .A1(local_key[12]), .A2(n4513), .A3(keyout[12]), .A4(n4529), .A5(prev_key[12]), .A6(n4530), .Y(n3776) );
  AO222X1_HVT U36 ( .A1(local_key[13]), .A2(n4513), .A3(keyout[13]), .A4(n4529), .A5(prev_key[13]), .A6(n4530), .Y(n3775) );
  AO222X1_HVT U37 ( .A1(local_key[14]), .A2(n4513), .A3(keyout[14]), .A4(n4529), .A5(prev_key[14]), .A6(n4530), .Y(n3774) );
  AO222X1_HVT U38 ( .A1(local_key[15]), .A2(n4513), .A3(keyout[15]), .A4(n4529), .A5(prev_key[15]), .A6(n4530), .Y(n3773) );
  AO222X1_HVT U39 ( .A1(local_key[16]), .A2(n4513), .A3(keyout[16]), .A4(n4529), .A5(prev_key[16]), .A6(n4530), .Y(n3772) );
  AO222X1_HVT U40 ( .A1(local_key[17]), .A2(n4513), .A3(keyout[17]), .A4(n4529), .A5(prev_key[17]), .A6(n4530), .Y(n3771) );
  AO222X1_HVT U41 ( .A1(local_key[18]), .A2(n4513), .A3(keyout[18]), .A4(n4529), .A5(prev_key[18]), .A6(n4530), .Y(n3770) );
  AO222X1_HVT U42 ( .A1(local_key[19]), .A2(n4513), .A3(keyout[19]), .A4(n4529), .A5(prev_key[19]), .A6(n4530), .Y(n3769) );
  AO222X1_HVT U43 ( .A1(local_key[20]), .A2(n4513), .A3(keyout[20]), .A4(n4529), .A5(prev_key[20]), .A6(n4530), .Y(n3768) );
  AO222X1_HVT U44 ( .A1(local_key[21]), .A2(n4513), .A3(keyout[21]), .A4(n4529), .A5(prev_key[21]), .A6(n4530), .Y(n3767) );
  AO222X1_HVT U45 ( .A1(local_key[22]), .A2(n4513), .A3(keyout[22]), .A4(n4529), .A5(prev_key[22]), .A6(n4530), .Y(n3766) );
  AO222X1_HVT U46 ( .A1(local_key[23]), .A2(n4513), .A3(keyout[23]), .A4(n4529), .A5(prev_key[23]), .A6(n4530), .Y(n3765) );
  AO222X1_HVT U47 ( .A1(local_key[24]), .A2(n4513), .A3(keyout[24]), .A4(n4529), .A5(prev_key[24]), .A6(n4530), .Y(n3764) );
  AO222X1_HVT U48 ( .A1(local_key[25]), .A2(n4513), .A3(keyout[25]), .A4(n4529), .A5(prev_key[25]), .A6(n4530), .Y(n3763) );
  AO222X1_HVT U49 ( .A1(local_key[26]), .A2(n4513), .A3(keyout[26]), .A4(n4529), .A5(prev_key[26]), .A6(n4530), .Y(n3762) );
  AO222X1_HVT U50 ( .A1(local_key[27]), .A2(n4513), .A3(keyout[27]), .A4(n4529), .A5(prev_key[27]), .A6(n4530), .Y(n3761) );
  AO222X1_HVT U51 ( .A1(local_key[28]), .A2(n4513), .A3(keyout[28]), .A4(n4529), .A5(prev_key[28]), .A6(n4530), .Y(n3760) );
  AO222X1_HVT U52 ( .A1(local_key[29]), .A2(n4513), .A3(keyout[29]), .A4(n4529), .A5(prev_key[29]), .A6(n4530), .Y(n3759) );
  AO222X1_HVT U53 ( .A1(local_key[30]), .A2(n4513), .A3(keyout[30]), .A4(n4529), .A5(prev_key[30]), .A6(n4530), .Y(n3758) );
  AO222X1_HVT U54 ( .A1(local_key[31]), .A2(n4513), .A3(keyout[31]), .A4(n4529), .A5(prev_key[31]), .A6(n4530), .Y(n3757) );
  AO222X1_HVT U55 ( .A1(local_key[32]), .A2(n4513), .A3(keyout[32]), .A4(n4529), .A5(prev_key[32]), .A6(n4530), .Y(n3756) );
  AO222X1_HVT U56 ( .A1(local_key[33]), .A2(n4513), .A3(keyout[33]), .A4(n4529), .A5(prev_key[33]), .A6(n4530), .Y(n3755) );
  AO222X1_HVT U57 ( .A1(local_key[34]), .A2(n4513), .A3(keyout[34]), .A4(n4529), .A5(prev_key[34]), .A6(n4530), .Y(n3754) );
  AO222X1_HVT U58 ( .A1(local_key[35]), .A2(n4513), .A3(keyout[35]), .A4(n4529), .A5(prev_key[35]), .A6(n4530), .Y(n3753) );
  AO222X1_HVT U59 ( .A1(local_key[36]), .A2(n4513), .A3(keyout[36]), .A4(n4529), .A5(prev_key[36]), .A6(n4530), .Y(n3752) );
  AO222X1_HVT U60 ( .A1(local_key[37]), .A2(n4513), .A3(keyout[37]), .A4(n4529), .A5(prev_key[37]), .A6(n4530), .Y(n3751) );
  AO222X1_HVT U61 ( .A1(local_key[38]), .A2(n4513), .A3(keyout[38]), .A4(n4529), .A5(prev_key[38]), .A6(n4530), .Y(n3750) );
  AO222X1_HVT U62 ( .A1(local_key[39]), .A2(n4513), .A3(keyout[39]), .A4(n4529), .A5(prev_key[39]), .A6(n4530), .Y(n3749) );
  AO222X1_HVT U63 ( .A1(local_key[40]), .A2(n4513), .A3(keyout[40]), .A4(n4529), .A5(prev_key[40]), .A6(n4530), .Y(n3748) );
  AO222X1_HVT U64 ( .A1(local_key[41]), .A2(n4513), .A3(keyout[41]), .A4(n4529), .A5(prev_key[41]), .A6(n4530), .Y(n3747) );
  AO222X1_HVT U65 ( .A1(local_key[42]), .A2(n4513), .A3(keyout[42]), .A4(n4529), .A5(prev_key[42]), .A6(n4530), .Y(n3746) );
  AO222X1_HVT U66 ( .A1(local_key[43]), .A2(n4513), .A3(keyout[43]), .A4(n4529), .A5(prev_key[43]), .A6(n4530), .Y(n3745) );
  AO222X1_HVT U67 ( .A1(local_key[44]), .A2(n4513), .A3(keyout[44]), .A4(n4529), .A5(prev_key[44]), .A6(n4530), .Y(n3744) );
  AO222X1_HVT U68 ( .A1(local_key[45]), .A2(n4513), .A3(keyout[45]), .A4(n4529), .A5(prev_key[45]), .A6(n4530), .Y(n3743) );
  AO222X1_HVT U69 ( .A1(local_key[46]), .A2(n4513), .A3(keyout[46]), .A4(n4529), .A5(prev_key[46]), .A6(n4530), .Y(n3742) );
  AO222X1_HVT U70 ( .A1(local_key[47]), .A2(n4513), .A3(keyout[47]), .A4(n4529), .A5(prev_key[47]), .A6(n4530), .Y(n3741) );
  AO222X1_HVT U71 ( .A1(local_key[48]), .A2(n4513), .A3(keyout[48]), .A4(n4529), .A5(prev_key[48]), .A6(n4530), .Y(n3740) );
  AO222X1_HVT U72 ( .A1(local_key[49]), .A2(n4513), .A3(keyout[49]), .A4(n4529), .A5(prev_key[49]), .A6(n4530), .Y(n3739) );
  AO222X1_HVT U73 ( .A1(local_key[50]), .A2(n4513), .A3(keyout[50]), .A4(n4529), .A5(prev_key[50]), .A6(n4530), .Y(n3738) );
  AO222X1_HVT U74 ( .A1(local_key[51]), .A2(n4513), .A3(keyout[51]), .A4(n4529), .A5(prev_key[51]), .A6(n4530), .Y(n3737) );
  AO222X1_HVT U75 ( .A1(local_key[52]), .A2(n4513), .A3(keyout[52]), .A4(n4529), .A5(prev_key[52]), .A6(n4530), .Y(n3736) );
  AO222X1_HVT U76 ( .A1(local_key[53]), .A2(n4513), .A3(keyout[53]), .A4(n4529), .A5(prev_key[53]), .A6(n4530), .Y(n3735) );
  AO222X1_HVT U77 ( .A1(local_key[54]), .A2(n4513), .A3(keyout[54]), .A4(n4529), .A5(prev_key[54]), .A6(n4530), .Y(n3734) );
  AO222X1_HVT U78 ( .A1(local_key[55]), .A2(n4513), .A3(keyout[55]), .A4(n4529), .A5(prev_key[55]), .A6(n4530), .Y(n3733) );
  AO222X1_HVT U79 ( .A1(local_key[56]), .A2(n4513), .A3(keyout[56]), .A4(n4529), .A5(prev_key[56]), .A6(n4530), .Y(n3732) );
  AO222X1_HVT U80 ( .A1(local_key[57]), .A2(n4513), .A3(keyout[57]), .A4(n4529), .A5(prev_key[57]), .A6(n4530), .Y(n3731) );
  AO222X1_HVT U81 ( .A1(local_key[58]), .A2(n4513), .A3(keyout[58]), .A4(n4529), .A5(prev_key[58]), .A6(n4530), .Y(n3730) );
  AO222X1_HVT U82 ( .A1(local_key[59]), .A2(n4513), .A3(keyout[59]), .A4(n4529), .A5(prev_key[59]), .A6(n4530), .Y(n3729) );
  AO222X1_HVT U83 ( .A1(local_key[60]), .A2(n4513), .A3(keyout[60]), .A4(n4529), .A5(prev_key[60]), .A6(n4530), .Y(n3728) );
  AO222X1_HVT U84 ( .A1(local_key[61]), .A2(n4513), .A3(keyout[61]), .A4(n4529), .A5(prev_key[61]), .A6(n4530), .Y(n3727) );
  AO222X1_HVT U85 ( .A1(local_key[62]), .A2(n4513), .A3(keyout[62]), .A4(n4529), .A5(prev_key[62]), .A6(n4530), .Y(n3726) );
  AO222X1_HVT U86 ( .A1(local_key[63]), .A2(n4513), .A3(keyout[63]), .A4(n4529), .A5(prev_key[63]), .A6(n4530), .Y(n3725) );
  AO222X1_HVT U87 ( .A1(local_key[64]), .A2(n4513), .A3(keyout[64]), .A4(n4529), .A5(prev_key[64]), .A6(n4530), .Y(n3724) );
  AO222X1_HVT U88 ( .A1(local_key[65]), .A2(n4513), .A3(keyout[65]), .A4(n4529), .A5(prev_key[65]), .A6(n4530), .Y(n3723) );
  AO222X1_HVT U89 ( .A1(local_key[66]), .A2(n4513), .A3(keyout[66]), .A4(n4529), .A5(prev_key[66]), .A6(n4530), .Y(n3722) );
  AO222X1_HVT U90 ( .A1(local_key[67]), .A2(n4513), .A3(keyout[67]), .A4(n4529), .A5(prev_key[67]), .A6(n4530), .Y(n3721) );
  AO222X1_HVT U91 ( .A1(local_key[68]), .A2(n4513), .A3(keyout[68]), .A4(n4529), .A5(prev_key[68]), .A6(n4530), .Y(n3720) );
  AO222X1_HVT U92 ( .A1(local_key[69]), .A2(n4513), .A3(keyout[69]), .A4(n4529), .A5(prev_key[69]), .A6(n4530), .Y(n3719) );
  AO222X1_HVT U93 ( .A1(local_key[70]), .A2(n4513), .A3(keyout[70]), .A4(n4529), .A5(prev_key[70]), .A6(n4530), .Y(n3718) );
  AO222X1_HVT U94 ( .A1(local_key[71]), .A2(n4513), .A3(keyout[71]), .A4(n4529), .A5(prev_key[71]), .A6(n4530), .Y(n3717) );
  AO222X1_HVT U95 ( .A1(local_key[72]), .A2(n4513), .A3(keyout[72]), .A4(n4529), .A5(prev_key[72]), .A6(n4530), .Y(n3716) );
  AO222X1_HVT U96 ( .A1(local_key[73]), .A2(n4513), .A3(keyout[73]), .A4(n4529), .A5(prev_key[73]), .A6(n4530), .Y(n3715) );
  AO222X1_HVT U97 ( .A1(local_key[74]), .A2(n4513), .A3(keyout[74]), .A4(n4529), .A5(prev_key[74]), .A6(n4530), .Y(n3714) );
  AO222X1_HVT U98 ( .A1(local_key[75]), .A2(n4513), .A3(keyout[75]), .A4(n4529), .A5(prev_key[75]), .A6(n4530), .Y(n3713) );
  AO222X1_HVT U99 ( .A1(local_key[76]), .A2(n4513), .A3(keyout[76]), .A4(n4529), .A5(prev_key[76]), .A6(n4530), .Y(n3712) );
  AO222X1_HVT U100 ( .A1(local_key[77]), .A2(n4513), .A3(keyout[77]), .A4(
        n4529), .A5(prev_key[77]), .A6(n4530), .Y(n3711) );
  AO222X1_HVT U101 ( .A1(local_key[78]), .A2(n4513), .A3(keyout[78]), .A4(
        n4529), .A5(prev_key[78]), .A6(n4530), .Y(n3710) );
  AO222X1_HVT U102 ( .A1(local_key[79]), .A2(n4513), .A3(keyout[79]), .A4(
        n4529), .A5(prev_key[79]), .A6(n4530), .Y(n3709) );
  AO222X1_HVT U103 ( .A1(local_key[80]), .A2(n4513), .A3(keyout[80]), .A4(
        n4529), .A5(prev_key[80]), .A6(n4530), .Y(n3708) );
  AO222X1_HVT U104 ( .A1(local_key[81]), .A2(n4513), .A3(keyout[81]), .A4(
        n4529), .A5(prev_key[81]), .A6(n4530), .Y(n3707) );
  AO222X1_HVT U105 ( .A1(local_key[82]), .A2(n4513), .A3(keyout[82]), .A4(
        n4529), .A5(prev_key[82]), .A6(n4530), .Y(n3706) );
  AO222X1_HVT U106 ( .A1(local_key[83]), .A2(n4513), .A3(keyout[83]), .A4(
        n4529), .A5(prev_key[83]), .A6(n4530), .Y(n3705) );
  AO222X1_HVT U107 ( .A1(local_key[84]), .A2(n4513), .A3(keyout[84]), .A4(
        n4529), .A5(prev_key[84]), .A6(n4530), .Y(n3704) );
  AO222X1_HVT U108 ( .A1(local_key[85]), .A2(n4513), .A3(keyout[85]), .A4(
        n4529), .A5(prev_key[85]), .A6(n4530), .Y(n3703) );
  AO222X1_HVT U109 ( .A1(local_key[86]), .A2(n4513), .A3(keyout[86]), .A4(
        n4529), .A5(prev_key[86]), .A6(n4530), .Y(n3702) );
  AO222X1_HVT U110 ( .A1(local_key[87]), .A2(n4513), .A3(keyout[87]), .A4(
        n4529), .A5(prev_key[87]), .A6(n4530), .Y(n3701) );
  AO222X1_HVT U111 ( .A1(local_key[88]), .A2(n4513), .A3(keyout[88]), .A4(
        n4529), .A5(prev_key[88]), .A6(n4530), .Y(n3700) );
  AO222X1_HVT U112 ( .A1(local_key[89]), .A2(n4513), .A3(keyout[89]), .A4(
        n4529), .A5(prev_key[89]), .A6(n4530), .Y(n3699) );
  AO222X1_HVT U113 ( .A1(local_key[90]), .A2(n4513), .A3(keyout[90]), .A4(
        n4529), .A5(prev_key[90]), .A6(n4530), .Y(n3698) );
  AO222X1_HVT U114 ( .A1(local_key[91]), .A2(n4513), .A3(keyout[91]), .A4(
        n4529), .A5(prev_key[91]), .A6(n4530), .Y(n3697) );
  AO222X1_HVT U115 ( .A1(local_key[92]), .A2(n4513), .A3(keyout[92]), .A4(
        n4529), .A5(prev_key[92]), .A6(n4530), .Y(n3696) );
  AO222X1_HVT U116 ( .A1(local_key[93]), .A2(n4513), .A3(keyout[93]), .A4(
        n4529), .A5(prev_key[93]), .A6(n4530), .Y(n3695) );
  AO222X1_HVT U117 ( .A1(local_key[94]), .A2(n4513), .A3(keyout[94]), .A4(
        n4529), .A5(prev_key[94]), .A6(n4530), .Y(n3694) );
  AO222X1_HVT U118 ( .A1(local_key[95]), .A2(n4513), .A3(keyout[95]), .A4(
        n4529), .A5(prev_key[95]), .A6(n4530), .Y(n3693) );
  AO222X1_HVT U119 ( .A1(local_key[96]), .A2(n4513), .A3(keyout[96]), .A4(
        n4529), .A5(prev_key[96]), .A6(n4530), .Y(n3692) );
  AO222X1_HVT U120 ( .A1(local_key[97]), .A2(n4513), .A3(keyout[97]), .A4(
        n4529), .A5(prev_key[97]), .A6(n4530), .Y(n3691) );
  AO222X1_HVT U121 ( .A1(local_key[98]), .A2(n4513), .A3(keyout[98]), .A4(
        n4529), .A5(prev_key[98]), .A6(n4530), .Y(n3690) );
  AO222X1_HVT U122 ( .A1(local_key[99]), .A2(n4513), .A3(keyout[99]), .A4(
        n4529), .A5(prev_key[99]), .A6(n4530), .Y(n3689) );
  AO222X1_HVT U123 ( .A1(local_key[100]), .A2(n4513), .A3(keyout[100]), .A4(
        n4529), .A5(prev_key[100]), .A6(n4530), .Y(n3688) );
  AO222X1_HVT U124 ( .A1(local_key[101]), .A2(n4513), .A3(keyout[101]), .A4(
        n4529), .A5(prev_key[101]), .A6(n4530), .Y(n3687) );
  AO222X1_HVT U125 ( .A1(local_key[102]), .A2(n4513), .A3(keyout[102]), .A4(
        n4529), .A5(prev_key[102]), .A6(n4530), .Y(n3686) );
  AO222X1_HVT U126 ( .A1(local_key[103]), .A2(n4513), .A3(keyout[103]), .A4(
        n4529), .A5(prev_key[103]), .A6(n4530), .Y(n3685) );
  AO222X1_HVT U127 ( .A1(local_key[104]), .A2(n4513), .A3(keyout[104]), .A4(
        n4529), .A5(prev_key[104]), .A6(n4530), .Y(n3684) );
  AO222X1_HVT U128 ( .A1(local_key[105]), .A2(n4513), .A3(keyout[105]), .A4(
        n4529), .A5(prev_key[105]), .A6(n4530), .Y(n3683) );
  AO222X1_HVT U129 ( .A1(local_key[106]), .A2(n4513), .A3(keyout[106]), .A4(
        n4529), .A5(prev_key[106]), .A6(n4530), .Y(n3682) );
  AO222X1_HVT U130 ( .A1(local_key[107]), .A2(n4513), .A3(keyout[107]), .A4(
        n4529), .A5(prev_key[107]), .A6(n4530), .Y(n3681) );
  AO222X1_HVT U131 ( .A1(local_key[108]), .A2(n4513), .A3(keyout[108]), .A4(
        n4529), .A5(prev_key[108]), .A6(n4530), .Y(n3680) );
  AO222X1_HVT U132 ( .A1(local_key[109]), .A2(n4513), .A3(keyout[109]), .A4(
        n4529), .A5(prev_key[109]), .A6(n4530), .Y(n3679) );
  AO222X1_HVT U133 ( .A1(local_key[110]), .A2(n4513), .A3(keyout[110]), .A4(
        n4529), .A5(prev_key[110]), .A6(n4530), .Y(n3678) );
  AO222X1_HVT U134 ( .A1(local_key[111]), .A2(n4513), .A3(keyout[111]), .A4(
        n4529), .A5(prev_key[111]), .A6(n4530), .Y(n3677) );
  AO222X1_HVT U135 ( .A1(local_key[112]), .A2(n4513), .A3(keyout[112]), .A4(
        n4529), .A5(prev_key[112]), .A6(n4530), .Y(n3676) );
  AO222X1_HVT U136 ( .A1(local_key[113]), .A2(n4513), .A3(keyout[113]), .A4(
        n4529), .A5(prev_key[113]), .A6(n4530), .Y(n3675) );
  AO222X1_HVT U137 ( .A1(local_key[114]), .A2(n4513), .A3(keyout[114]), .A4(
        n4529), .A5(prev_key[114]), .A6(n4530), .Y(n3674) );
  AO222X1_HVT U138 ( .A1(local_key[115]), .A2(n4513), .A3(keyout[115]), .A4(
        n4529), .A5(prev_key[115]), .A6(n4530), .Y(n3673) );
  AO222X1_HVT U139 ( .A1(local_key[116]), .A2(n4513), .A3(keyout[116]), .A4(
        n4529), .A5(prev_key[116]), .A6(n4530), .Y(n3672) );
  AO222X1_HVT U140 ( .A1(local_key[117]), .A2(n4513), .A3(keyout[117]), .A4(
        n4529), .A5(prev_key[117]), .A6(n4530), .Y(n3671) );
  AO222X1_HVT U141 ( .A1(local_key[118]), .A2(n4513), .A3(keyout[118]), .A4(
        n4529), .A5(prev_key[118]), .A6(n4530), .Y(n3670) );
  AO222X1_HVT U142 ( .A1(local_key[119]), .A2(n4513), .A3(keyout[119]), .A4(
        n4529), .A5(prev_key[119]), .A6(n4530), .Y(n3669) );
  AO222X1_HVT U143 ( .A1(local_key[120]), .A2(n4513), .A3(keyout[120]), .A4(
        n4529), .A5(prev_key[120]), .A6(n4530), .Y(n3668) );
  AO222X1_HVT U144 ( .A1(local_key[121]), .A2(n4513), .A3(keyout[121]), .A4(
        n4529), .A5(prev_key[121]), .A6(n4530), .Y(n3667) );
  AO222X1_HVT U145 ( .A1(local_key[122]), .A2(n4513), .A3(keyout[122]), .A4(
        n4529), .A5(prev_key[122]), .A6(n4530), .Y(n3666) );
  AO222X1_HVT U146 ( .A1(local_key[123]), .A2(n4513), .A3(keyout[123]), .A4(
        n4529), .A5(prev_key[123]), .A6(n4530), .Y(n3665) );
  AO222X1_HVT U147 ( .A1(local_key[124]), .A2(n4513), .A3(keyout[124]), .A4(
        n4529), .A5(prev_key[124]), .A6(n4530), .Y(n3664) );
  AO222X1_HVT U148 ( .A1(local_key[125]), .A2(n4513), .A3(keyout[125]), .A4(
        n4529), .A5(prev_key[125]), .A6(n4530), .Y(n3663) );
  AO222X1_HVT U149 ( .A1(local_key[126]), .A2(n4513), .A3(keyout[126]), .A4(
        n4529), .A5(prev_key[126]), .A6(n4530), .Y(n3662) );
  AO222X1_HVT U150 ( .A1(local_key[127]), .A2(n4513), .A3(keyout[127]), .A4(
        n4529), .A5(prev_key[127]), .A6(n4530), .Y(n3661) );
  INVX0_HVT U151 ( .A(n4516), .Y(n4530) );
  AND2X1_HVT U152 ( .A1(n4516), .A2(n4510), .Y(n4529) );
  AND2X1_HVT U153 ( .A1(n4516), .A2(n4531), .Y(n4513) );
  OA21X1_HVT U154 ( .A1(n4510), .A2(n4531), .A3(n4511), .Y(n4516) );
  NAND4X0_HVT U155 ( .A1(n4532), .A2(n4527), .A3(n4525), .A4(n4523), .Y(n4510)
         );
  AND2X1_HVT U156 ( .A1(n4517), .A2(n4533), .Y(n4527) );
  INVX0_HVT U157 ( .A(n4520), .Y(n4532) );
  NAND2X0_HVT U158 ( .A1(n4534), .A2(n4528), .Y(n4520) );
  MUX21X1_HVT U159 ( .A1(local_key[127]), .A2(n4366), .S0(n4504), .Y(n3660) );
  MUX21X1_HVT U160 ( .A1(local_key[126]), .A2(n4367), .S0(n4504), .Y(n3659) );
  MUX21X1_HVT U161 ( .A1(local_key[125]), .A2(n4368), .S0(n4504), .Y(n3658) );
  MUX21X1_HVT U162 ( .A1(local_key[124]), .A2(n4369), .S0(n4504), .Y(n3657) );
  MUX21X1_HVT U163 ( .A1(local_key[123]), .A2(n4370), .S0(n4504), .Y(n3656) );
  MUX21X1_HVT U164 ( .A1(local_key[122]), .A2(n4371), .S0(n4504), .Y(n3655) );
  MUX21X1_HVT U165 ( .A1(local_key[121]), .A2(n4372), .S0(n4504), .Y(n3654) );
  MUX21X1_HVT U166 ( .A1(local_key[120]), .A2(n4373), .S0(n4504), .Y(n3653) );
  MUX21X1_HVT U167 ( .A1(local_key[119]), .A2(n4374), .S0(n4504), .Y(n3652) );
  MUX21X1_HVT U168 ( .A1(local_key[118]), .A2(n4375), .S0(n4504), .Y(n3651) );
  MUX21X1_HVT U169 ( .A1(local_key[117]), .A2(n4376), .S0(n4504), .Y(n3650) );
  MUX21X1_HVT U170 ( .A1(local_key[116]), .A2(n4377), .S0(n4504), .Y(n3649) );
  MUX21X1_HVT U171 ( .A1(local_key[115]), .A2(n4378), .S0(n4504), .Y(n3648) );
  MUX21X1_HVT U172 ( .A1(local_key[114]), .A2(n4379), .S0(n4504), .Y(n3647) );
  MUX21X1_HVT U173 ( .A1(local_key[113]), .A2(n4380), .S0(n4504), .Y(n3646) );
  MUX21X1_HVT U174 ( .A1(local_key[112]), .A2(n4381), .S0(n4504), .Y(n3645) );
  MUX21X1_HVT U175 ( .A1(local_key[111]), .A2(n4382), .S0(n4504), .Y(n3644) );
  MUX21X1_HVT U176 ( .A1(local_key[110]), .A2(n4383), .S0(n4504), .Y(n3643) );
  MUX21X1_HVT U177 ( .A1(local_key[109]), .A2(n4384), .S0(n4504), .Y(n3642) );
  MUX21X1_HVT U178 ( .A1(local_key[108]), .A2(n4385), .S0(n4504), .Y(n3641) );
  MUX21X1_HVT U179 ( .A1(local_key[107]), .A2(n4386), .S0(n4504), .Y(n3640) );
  MUX21X1_HVT U180 ( .A1(local_key[106]), .A2(n4387), .S0(n4504), .Y(n3639) );
  MUX21X1_HVT U181 ( .A1(local_key[105]), .A2(n4388), .S0(n4504), .Y(n3638) );
  MUX21X1_HVT U182 ( .A1(local_key[104]), .A2(n4389), .S0(n4504), .Y(n3637) );
  MUX21X1_HVT U183 ( .A1(local_key[103]), .A2(n4390), .S0(n4504), .Y(n3636) );
  MUX21X1_HVT U184 ( .A1(local_key[102]), .A2(n4391), .S0(n4504), .Y(n3635) );
  MUX21X1_HVT U185 ( .A1(local_key[101]), .A2(n4392), .S0(n4504), .Y(n3634) );
  MUX21X1_HVT U186 ( .A1(local_key[100]), .A2(n4393), .S0(n4504), .Y(n3633) );
  MUX21X1_HVT U187 ( .A1(local_key[99]), .A2(n4394), .S0(n4504), .Y(n3632) );
  MUX21X1_HVT U188 ( .A1(local_key[98]), .A2(n4395), .S0(n4504), .Y(n3631) );
  MUX21X1_HVT U189 ( .A1(local_key[97]), .A2(n4396), .S0(n4504), .Y(n3630) );
  MUX21X1_HVT U190 ( .A1(local_key[96]), .A2(n4397), .S0(n4504), .Y(n3629) );
  MUX21X1_HVT U191 ( .A1(local_key[95]), .A2(n4398), .S0(n4504), .Y(n3628) );
  MUX21X1_HVT U192 ( .A1(local_key[94]), .A2(n4399), .S0(n4504), .Y(n3627) );
  MUX21X1_HVT U193 ( .A1(local_key[93]), .A2(n4400), .S0(n4504), .Y(n3626) );
  MUX21X1_HVT U194 ( .A1(local_key[92]), .A2(n4401), .S0(n4504), .Y(n3625) );
  MUX21X1_HVT U195 ( .A1(local_key[91]), .A2(n4402), .S0(n4504), .Y(n3624) );
  MUX21X1_HVT U196 ( .A1(local_key[90]), .A2(n4403), .S0(n4504), .Y(n3623) );
  MUX21X1_HVT U197 ( .A1(local_key[89]), .A2(n4404), .S0(n4504), .Y(n3622) );
  MUX21X1_HVT U198 ( .A1(local_key[88]), .A2(n4405), .S0(n4504), .Y(n3621) );
  MUX21X1_HVT U199 ( .A1(local_key[87]), .A2(n4406), .S0(n4504), .Y(n3620) );
  MUX21X1_HVT U200 ( .A1(local_key[86]), .A2(n4407), .S0(n4504), .Y(n3619) );
  MUX21X1_HVT U201 ( .A1(local_key[85]), .A2(n4408), .S0(n4504), .Y(n3618) );
  MUX21X1_HVT U202 ( .A1(local_key[84]), .A2(n4409), .S0(n4504), .Y(n3617) );
  MUX21X1_HVT U203 ( .A1(local_key[83]), .A2(n4410), .S0(n4504), .Y(n3616) );
  MUX21X1_HVT U204 ( .A1(local_key[82]), .A2(n4411), .S0(n4504), .Y(n3615) );
  MUX21X1_HVT U205 ( .A1(local_key[81]), .A2(n4412), .S0(n4504), .Y(n3614) );
  MUX21X1_HVT U206 ( .A1(local_key[80]), .A2(n4413), .S0(n4504), .Y(n3613) );
  MUX21X1_HVT U207 ( .A1(local_key[79]), .A2(n4414), .S0(n4504), .Y(n3612) );
  MUX21X1_HVT U208 ( .A1(local_key[78]), .A2(n4415), .S0(n4504), .Y(n3611) );
  MUX21X1_HVT U209 ( .A1(local_key[77]), .A2(n4416), .S0(n4504), .Y(n3610) );
  MUX21X1_HVT U210 ( .A1(local_key[76]), .A2(n4417), .S0(n4504), .Y(n3609) );
  MUX21X1_HVT U211 ( .A1(local_key[75]), .A2(n4418), .S0(n4504), .Y(n3608) );
  MUX21X1_HVT U212 ( .A1(local_key[74]), .A2(n4419), .S0(n4504), .Y(n3607) );
  MUX21X1_HVT U213 ( .A1(local_key[73]), .A2(n4420), .S0(n4504), .Y(n3606) );
  MUX21X1_HVT U214 ( .A1(local_key[72]), .A2(n4421), .S0(n4504), .Y(n3605) );
  MUX21X1_HVT U215 ( .A1(local_key[71]), .A2(n4422), .S0(n4504), .Y(n3604) );
  MUX21X1_HVT U216 ( .A1(local_key[70]), .A2(n4423), .S0(n4504), .Y(n3603) );
  MUX21X1_HVT U217 ( .A1(local_key[69]), .A2(n4424), .S0(n4504), .Y(n3602) );
  MUX21X1_HVT U218 ( .A1(local_key[68]), .A2(n4425), .S0(n4504), .Y(n3601) );
  MUX21X1_HVT U219 ( .A1(local_key[67]), .A2(n4426), .S0(n4504), .Y(n3600) );
  MUX21X1_HVT U220 ( .A1(local_key[66]), .A2(n4427), .S0(n4504), .Y(n3599) );
  MUX21X1_HVT U221 ( .A1(local_key[65]), .A2(n4428), .S0(n4504), .Y(n3598) );
  MUX21X1_HVT U222 ( .A1(local_key[64]), .A2(n4429), .S0(n4504), .Y(n3597) );
  MUX21X1_HVT U223 ( .A1(local_key[63]), .A2(n4430), .S0(n4504), .Y(n3596) );
  MUX21X1_HVT U224 ( .A1(local_key[62]), .A2(n4431), .S0(n4504), .Y(n3595) );
  MUX21X1_HVT U225 ( .A1(local_key[61]), .A2(n4432), .S0(n4504), .Y(n3594) );
  MUX21X1_HVT U226 ( .A1(local_key[60]), .A2(n4433), .S0(n4504), .Y(n3593) );
  MUX21X1_HVT U227 ( .A1(local_key[59]), .A2(n4434), .S0(n4504), .Y(n3592) );
  MUX21X1_HVT U228 ( .A1(local_key[58]), .A2(n4435), .S0(n4504), .Y(n3591) );
  MUX21X1_HVT U229 ( .A1(local_key[57]), .A2(n4436), .S0(n4504), .Y(n3590) );
  MUX21X1_HVT U230 ( .A1(local_key[56]), .A2(n4437), .S0(n4504), .Y(n3589) );
  MUX21X1_HVT U231 ( .A1(local_key[55]), .A2(n4438), .S0(n4504), .Y(n3588) );
  MUX21X1_HVT U232 ( .A1(local_key[54]), .A2(n4439), .S0(n4504), .Y(n3587) );
  MUX21X1_HVT U233 ( .A1(local_key[53]), .A2(n4440), .S0(n4504), .Y(n3586) );
  MUX21X1_HVT U234 ( .A1(local_key[52]), .A2(n4441), .S0(n4504), .Y(n3585) );
  MUX21X1_HVT U235 ( .A1(local_key[51]), .A2(n4442), .S0(n4504), .Y(n3584) );
  MUX21X1_HVT U236 ( .A1(local_key[50]), .A2(n4443), .S0(n4504), .Y(n3583) );
  MUX21X1_HVT U237 ( .A1(local_key[49]), .A2(n4444), .S0(n4504), .Y(n3582) );
  MUX21X1_HVT U238 ( .A1(local_key[48]), .A2(n4445), .S0(n4504), .Y(n3581) );
  MUX21X1_HVT U239 ( .A1(local_key[47]), .A2(n4446), .S0(n4504), .Y(n3580) );
  MUX21X1_HVT U240 ( .A1(local_key[46]), .A2(n4447), .S0(n4504), .Y(n3579) );
  MUX21X1_HVT U241 ( .A1(local_key[45]), .A2(n4448), .S0(n4504), .Y(n3578) );
  MUX21X1_HVT U242 ( .A1(local_key[44]), .A2(n4449), .S0(n4504), .Y(n3577) );
  MUX21X1_HVT U243 ( .A1(local_key[43]), .A2(n4450), .S0(n4504), .Y(n3576) );
  MUX21X1_HVT U244 ( .A1(local_key[42]), .A2(n4451), .S0(n4504), .Y(n3575) );
  MUX21X1_HVT U245 ( .A1(local_key[41]), .A2(n4452), .S0(n4504), .Y(n3574) );
  MUX21X1_HVT U246 ( .A1(local_key[40]), .A2(n4453), .S0(n4504), .Y(n3573) );
  MUX21X1_HVT U247 ( .A1(local_key[39]), .A2(n4454), .S0(n4504), .Y(n3572) );
  MUX21X1_HVT U248 ( .A1(local_key[38]), .A2(n4455), .S0(n4504), .Y(n3571) );
  MUX21X1_HVT U249 ( .A1(local_key[37]), .A2(n4456), .S0(n4504), .Y(n3570) );
  MUX21X1_HVT U250 ( .A1(local_key[36]), .A2(n4457), .S0(n4504), .Y(n3569) );
  MUX21X1_HVT U251 ( .A1(local_key[35]), .A2(n4458), .S0(n4504), .Y(n3568) );
  MUX21X1_HVT U252 ( .A1(local_key[34]), .A2(n4459), .S0(n4504), .Y(n3567) );
  MUX21X1_HVT U253 ( .A1(local_key[33]), .A2(n4460), .S0(n4504), .Y(n3566) );
  MUX21X1_HVT U254 ( .A1(local_key[32]), .A2(n4461), .S0(n4504), .Y(n3565) );
  MUX21X1_HVT U255 ( .A1(local_key[31]), .A2(n4462), .S0(n4504), .Y(n3564) );
  MUX21X1_HVT U256 ( .A1(local_key[30]), .A2(n4463), .S0(n4504), .Y(n3563) );
  MUX21X1_HVT U257 ( .A1(local_key[29]), .A2(n4464), .S0(n4504), .Y(n3562) );
  MUX21X1_HVT U258 ( .A1(local_key[28]), .A2(n4465), .S0(n4504), .Y(n3561) );
  MUX21X1_HVT U259 ( .A1(local_key[27]), .A2(n4466), .S0(n4504), .Y(n3560) );
  MUX21X1_HVT U260 ( .A1(local_key[26]), .A2(n4467), .S0(n4504), .Y(n3559) );
  MUX21X1_HVT U261 ( .A1(local_key[25]), .A2(n4468), .S0(n4504), .Y(n3558) );
  MUX21X1_HVT U262 ( .A1(local_key[24]), .A2(n4469), .S0(n4504), .Y(n3557) );
  MUX21X1_HVT U263 ( .A1(local_key[23]), .A2(n4470), .S0(n4504), .Y(n3556) );
  MUX21X1_HVT U264 ( .A1(local_key[22]), .A2(n4471), .S0(n4504), .Y(n3555) );
  MUX21X1_HVT U265 ( .A1(local_key[21]), .A2(n4472), .S0(n4504), .Y(n3554) );
  MUX21X1_HVT U266 ( .A1(local_key[20]), .A2(n4473), .S0(n4504), .Y(n3553) );
  MUX21X1_HVT U267 ( .A1(local_key[19]), .A2(n4474), .S0(n4504), .Y(n3552) );
  MUX21X1_HVT U268 ( .A1(local_key[18]), .A2(n4475), .S0(n4504), .Y(n3551) );
  MUX21X1_HVT U269 ( .A1(local_key[17]), .A2(n4476), .S0(n4504), .Y(n3550) );
  MUX21X1_HVT U270 ( .A1(local_key[16]), .A2(n4477), .S0(n4504), .Y(n3549) );
  MUX21X1_HVT U271 ( .A1(local_key[15]), .A2(n4478), .S0(n4504), .Y(n3548) );
  MUX21X1_HVT U272 ( .A1(local_key[14]), .A2(n4479), .S0(n4504), .Y(n3547) );
  MUX21X1_HVT U273 ( .A1(local_key[13]), .A2(n4480), .S0(n4504), .Y(n3546) );
  MUX21X1_HVT U274 ( .A1(local_key[12]), .A2(n4481), .S0(n4504), .Y(n3545) );
  MUX21X1_HVT U275 ( .A1(local_key[11]), .A2(n4482), .S0(n4504), .Y(n3544) );
  MUX21X1_HVT U276 ( .A1(local_key[10]), .A2(n4483), .S0(n4504), .Y(n3543) );
  MUX21X1_HVT U277 ( .A1(local_key[9]), .A2(n4484), .S0(n4504), .Y(n3542) );
  MUX21X1_HVT U278 ( .A1(local_key[8]), .A2(n4485), .S0(n4504), .Y(n3541) );
  MUX21X1_HVT U279 ( .A1(local_key[7]), .A2(n4486), .S0(n4504), .Y(n3540) );
  MUX21X1_HVT U280 ( .A1(local_key[6]), .A2(n4487), .S0(n4504), .Y(n3539) );
  MUX21X1_HVT U281 ( .A1(local_key[5]), .A2(n4488), .S0(n4504), .Y(n3538) );
  MUX21X1_HVT U282 ( .A1(local_key[4]), .A2(n4489), .S0(n4504), .Y(n3537) );
  MUX21X1_HVT U283 ( .A1(local_key[3]), .A2(n4490), .S0(n4504), .Y(n3536) );
  MUX21X1_HVT U284 ( .A1(local_key[2]), .A2(n4491), .S0(n4504), .Y(n3535) );
  MUX21X1_HVT U285 ( .A1(local_key[1]), .A2(n4492), .S0(n4504), .Y(n3534) );
  MUX21X1_HVT U286 ( .A1(local_key[0]), .A2(n4493), .S0(n4504), .Y(n3533) );
  NAND2X0_HVT U287 ( .A1(n4531), .A2(n4511), .Y(n4504) );
  AND4X1_HVT U288 ( .A1(n1), .A2(n3), .A3(n2), .A4(n4), .Y(n4531) );
  MUX21X1_HVT U289 ( .A1(keyout[127]), .A2(n5), .S0(n4507), .Y(n3532) );
  MUX21X1_HVT U290 ( .A1(keyout[126]), .A2(n6), .S0(n4507), .Y(n3531) );
  MUX21X1_HVT U291 ( .A1(keyout[125]), .A2(n7), .S0(n4507), .Y(n3530) );
  MUX21X1_HVT U292 ( .A1(keyout[124]), .A2(n8), .S0(n4507), .Y(n3529) );
  MUX21X1_HVT U293 ( .A1(keyout[123]), .A2(n9), .S0(n4507), .Y(n3528) );
  MUX21X1_HVT U294 ( .A1(keyout[122]), .A2(n10), .S0(n4507), .Y(n3527) );
  MUX21X1_HVT U295 ( .A1(keyout[121]), .A2(n11), .S0(n4507), .Y(n3526) );
  MUX21X1_HVT U296 ( .A1(keyout[120]), .A2(n12), .S0(n4507), .Y(n3525) );
  MUX21X1_HVT U297 ( .A1(keyout[119]), .A2(n13), .S0(n4507), .Y(n3524) );
  MUX21X1_HVT U298 ( .A1(keyout[118]), .A2(n14), .S0(n4507), .Y(n3523) );
  MUX21X1_HVT U299 ( .A1(keyout[117]), .A2(n15), .S0(n4507), .Y(n3522) );
  MUX21X1_HVT U300 ( .A1(keyout[116]), .A2(n16), .S0(n4507), .Y(n3521) );
  MUX21X1_HVT U301 ( .A1(keyout[115]), .A2(n17), .S0(n4507), .Y(n3520) );
  MUX21X1_HVT U302 ( .A1(keyout[114]), .A2(n18), .S0(n4507), .Y(n3519) );
  MUX21X1_HVT U303 ( .A1(keyout[113]), .A2(n1427), .S0(n4507), .Y(n3518) );
  MUX21X1_HVT U304 ( .A1(keyout[112]), .A2(n1428), .S0(n4507), .Y(n3517) );
  MUX21X1_HVT U305 ( .A1(keyout[111]), .A2(n1429), .S0(n4507), .Y(n3516) );
  MUX21X1_HVT U306 ( .A1(keyout[110]), .A2(n1430), .S0(n4507), .Y(n3515) );
  MUX21X1_HVT U307 ( .A1(keyout[109]), .A2(n1431), .S0(n4507), .Y(n3514) );
  MUX21X1_HVT U308 ( .A1(keyout[108]), .A2(n1432), .S0(n4507), .Y(n3513) );
  MUX21X1_HVT U309 ( .A1(keyout[107]), .A2(n1433), .S0(n4507), .Y(n3512) );
  MUX21X1_HVT U310 ( .A1(keyout[106]), .A2(n1434), .S0(n4507), .Y(n3511) );
  MUX21X1_HVT U311 ( .A1(keyout[105]), .A2(n1435), .S0(n4507), .Y(n3510) );
  MUX21X1_HVT U312 ( .A1(keyout[104]), .A2(n1436), .S0(n4507), .Y(n3509) );
  MUX21X1_HVT U313 ( .A1(keyout[103]), .A2(n1437), .S0(n4507), .Y(n3508) );
  MUX21X1_HVT U314 ( .A1(keyout[102]), .A2(n1438), .S0(n4507), .Y(n3507) );
  MUX21X1_HVT U315 ( .A1(keyout[101]), .A2(n1439), .S0(n4507), .Y(n3506) );
  MUX21X1_HVT U316 ( .A1(keyout[100]), .A2(n1440), .S0(n4507), .Y(n3505) );
  MUX21X1_HVT U317 ( .A1(keyout[99]), .A2(n1441), .S0(n4507), .Y(n3504) );
  MUX21X1_HVT U318 ( .A1(keyout[98]), .A2(n1442), .S0(n4507), .Y(n3503) );
  MUX21X1_HVT U319 ( .A1(keyout[97]), .A2(n1443), .S0(n4507), .Y(n3502) );
  MUX21X1_HVT U320 ( .A1(keyout[96]), .A2(n1444), .S0(n4507), .Y(n3501) );
  MUX21X1_HVT U321 ( .A1(keyout[95]), .A2(n1445), .S0(n4507), .Y(n3500) );
  MUX21X1_HVT U322 ( .A1(keyout[94]), .A2(n1446), .S0(n4507), .Y(n3499) );
  MUX21X1_HVT U323 ( .A1(keyout[93]), .A2(n1447), .S0(n4507), .Y(n3498) );
  MUX21X1_HVT U324 ( .A1(keyout[92]), .A2(n1448), .S0(n4507), .Y(n3497) );
  MUX21X1_HVT U325 ( .A1(keyout[91]), .A2(n1449), .S0(n4507), .Y(n3496) );
  MUX21X1_HVT U326 ( .A1(keyout[90]), .A2(n1450), .S0(n4507), .Y(n3495) );
  MUX21X1_HVT U327 ( .A1(keyout[89]), .A2(n1451), .S0(n4507), .Y(n3494) );
  MUX21X1_HVT U328 ( .A1(keyout[88]), .A2(n1452), .S0(n4507), .Y(n3493) );
  MUX21X1_HVT U329 ( .A1(keyout[87]), .A2(n1453), .S0(n4507), .Y(n3492) );
  MUX21X1_HVT U330 ( .A1(keyout[86]), .A2(n1454), .S0(n4507), .Y(n3491) );
  MUX21X1_HVT U331 ( .A1(keyout[85]), .A2(n1455), .S0(n4507), .Y(n3490) );
  MUX21X1_HVT U332 ( .A1(keyout[84]), .A2(n1456), .S0(n4507), .Y(n3489) );
  MUX21X1_HVT U333 ( .A1(keyout[83]), .A2(n1457), .S0(n4507), .Y(n3488) );
  MUX21X1_HVT U334 ( .A1(keyout[82]), .A2(n1458), .S0(n4507), .Y(n3487) );
  MUX21X1_HVT U335 ( .A1(keyout[81]), .A2(n1459), .S0(n4507), .Y(n3486) );
  MUX21X1_HVT U336 ( .A1(keyout[80]), .A2(n1460), .S0(n4507), .Y(n3485) );
  MUX21X1_HVT U337 ( .A1(keyout[79]), .A2(n1461), .S0(n4507), .Y(n3484) );
  MUX21X1_HVT U338 ( .A1(keyout[78]), .A2(n1462), .S0(n4507), .Y(n3483) );
  MUX21X1_HVT U339 ( .A1(keyout[77]), .A2(n1463), .S0(n4507), .Y(n3482) );
  MUX21X1_HVT U340 ( .A1(keyout[76]), .A2(n1464), .S0(n4507), .Y(n3481) );
  MUX21X1_HVT U341 ( .A1(keyout[75]), .A2(n1465), .S0(n4507), .Y(n3480) );
  MUX21X1_HVT U342 ( .A1(keyout[74]), .A2(n1466), .S0(n4507), .Y(n3479) );
  MUX21X1_HVT U343 ( .A1(keyout[73]), .A2(n1467), .S0(n4507), .Y(n3478) );
  MUX21X1_HVT U344 ( .A1(keyout[72]), .A2(n1468), .S0(n4507), .Y(n3477) );
  MUX21X1_HVT U345 ( .A1(keyout[71]), .A2(n1469), .S0(n4507), .Y(n3476) );
  MUX21X1_HVT U346 ( .A1(keyout[70]), .A2(n1470), .S0(n4507), .Y(n3475) );
  MUX21X1_HVT U347 ( .A1(keyout[69]), .A2(n1471), .S0(n4507), .Y(n3474) );
  MUX21X1_HVT U348 ( .A1(keyout[68]), .A2(n1472), .S0(n4507), .Y(n3473) );
  MUX21X1_HVT U349 ( .A1(keyout[67]), .A2(n1473), .S0(n4507), .Y(n3472) );
  MUX21X1_HVT U350 ( .A1(keyout[66]), .A2(n1474), .S0(n4507), .Y(n3471) );
  MUX21X1_HVT U351 ( .A1(keyout[65]), .A2(n1475), .S0(n4507), .Y(n3470) );
  MUX21X1_HVT U352 ( .A1(keyout[64]), .A2(n1476), .S0(n4507), .Y(n3469) );
  MUX21X1_HVT U353 ( .A1(keyout[63]), .A2(n1477), .S0(n4507), .Y(n3468) );
  MUX21X1_HVT U354 ( .A1(keyout[62]), .A2(n1478), .S0(n4507), .Y(n3467) );
  MUX21X1_HVT U355 ( .A1(keyout[61]), .A2(n1479), .S0(n4507), .Y(n3466) );
  MUX21X1_HVT U356 ( .A1(keyout[60]), .A2(n1480), .S0(n4507), .Y(n3465) );
  MUX21X1_HVT U357 ( .A1(keyout[59]), .A2(n1481), .S0(n4507), .Y(n3464) );
  MUX21X1_HVT U358 ( .A1(keyout[58]), .A2(n1482), .S0(n4507), .Y(n3463) );
  MUX21X1_HVT U359 ( .A1(keyout[57]), .A2(n1483), .S0(n4507), .Y(n3462) );
  MUX21X1_HVT U360 ( .A1(keyout[56]), .A2(n1484), .S0(n4507), .Y(n3461) );
  MUX21X1_HVT U361 ( .A1(keyout[55]), .A2(n1485), .S0(n4507), .Y(n3460) );
  MUX21X1_HVT U362 ( .A1(keyout[54]), .A2(n1486), .S0(n4507), .Y(n3459) );
  MUX21X1_HVT U363 ( .A1(keyout[53]), .A2(n1487), .S0(n4507), .Y(n3458) );
  MUX21X1_HVT U364 ( .A1(keyout[52]), .A2(n1488), .S0(n4507), .Y(n3457) );
  MUX21X1_HVT U365 ( .A1(keyout[51]), .A2(n1489), .S0(n4507), .Y(n3456) );
  MUX21X1_HVT U366 ( .A1(keyout[50]), .A2(n1490), .S0(n4507), .Y(n3455) );
  MUX21X1_HVT U367 ( .A1(keyout[49]), .A2(n1491), .S0(n4507), .Y(n3454) );
  MUX21X1_HVT U368 ( .A1(keyout[48]), .A2(n1492), .S0(n4507), .Y(n3453) );
  MUX21X1_HVT U369 ( .A1(keyout[47]), .A2(n1493), .S0(n4507), .Y(n3452) );
  MUX21X1_HVT U370 ( .A1(keyout[46]), .A2(n1494), .S0(n4507), .Y(n3451) );
  MUX21X1_HVT U371 ( .A1(keyout[45]), .A2(n1495), .S0(n4507), .Y(n3450) );
  MUX21X1_HVT U372 ( .A1(keyout[44]), .A2(n1496), .S0(n4507), .Y(n3449) );
  MUX21X1_HVT U373 ( .A1(keyout[43]), .A2(n1497), .S0(n4507), .Y(n3448) );
  MUX21X1_HVT U374 ( .A1(keyout[42]), .A2(n1498), .S0(n4507), .Y(n3447) );
  MUX21X1_HVT U375 ( .A1(keyout[41]), .A2(n1499), .S0(n4507), .Y(n3446) );
  MUX21X1_HVT U376 ( .A1(keyout[40]), .A2(n1500), .S0(n4507), .Y(n3445) );
  MUX21X1_HVT U377 ( .A1(keyout[39]), .A2(n1501), .S0(n4507), .Y(n3444) );
  MUX21X1_HVT U378 ( .A1(keyout[38]), .A2(n1502), .S0(n4507), .Y(n3443) );
  MUX21X1_HVT U379 ( .A1(keyout[37]), .A2(n1503), .S0(n4507), .Y(n3442) );
  MUX21X1_HVT U380 ( .A1(keyout[36]), .A2(n1504), .S0(n4507), .Y(n3441) );
  MUX21X1_HVT U381 ( .A1(keyout[35]), .A2(n1505), .S0(n4507), .Y(n3440) );
  MUX21X1_HVT U382 ( .A1(keyout[34]), .A2(n1506), .S0(n4507), .Y(n3439) );
  MUX21X1_HVT U383 ( .A1(keyout[33]), .A2(n1507), .S0(n4507), .Y(n3438) );
  MUX21X1_HVT U384 ( .A1(keyout[32]), .A2(n1508), .S0(n4507), .Y(n3437) );
  MUX21X1_HVT U385 ( .A1(keyout[31]), .A2(n1509), .S0(n4507), .Y(n3436) );
  MUX21X1_HVT U386 ( .A1(keyout[30]), .A2(n1510), .S0(n4507), .Y(n3435) );
  MUX21X1_HVT U387 ( .A1(keyout[29]), .A2(n1511), .S0(n4507), .Y(n3434) );
  MUX21X1_HVT U388 ( .A1(keyout[28]), .A2(n1512), .S0(n4507), .Y(n3433) );
  MUX21X1_HVT U389 ( .A1(keyout[27]), .A2(n1513), .S0(n4507), .Y(n3432) );
  MUX21X1_HVT U390 ( .A1(keyout[26]), .A2(n1514), .S0(n4507), .Y(n3431) );
  MUX21X1_HVT U391 ( .A1(keyout[25]), .A2(n1515), .S0(n4507), .Y(n3430) );
  MUX21X1_HVT U392 ( .A1(keyout[24]), .A2(n1516), .S0(n4507), .Y(n3429) );
  MUX21X1_HVT U393 ( .A1(keyout[23]), .A2(n1517), .S0(n4507), .Y(n3428) );
  MUX21X1_HVT U394 ( .A1(keyout[22]), .A2(n1518), .S0(n4507), .Y(n3427) );
  MUX21X1_HVT U395 ( .A1(keyout[21]), .A2(n1519), .S0(n4507), .Y(n3426) );
  MUX21X1_HVT U396 ( .A1(keyout[20]), .A2(n1520), .S0(n4507), .Y(n3425) );
  MUX21X1_HVT U397 ( .A1(keyout[19]), .A2(n1521), .S0(n4507), .Y(n3424) );
  MUX21X1_HVT U398 ( .A1(keyout[18]), .A2(n1522), .S0(n4507), .Y(n3423) );
  MUX21X1_HVT U399 ( .A1(keyout[17]), .A2(n1523), .S0(n4507), .Y(n3422) );
  MUX21X1_HVT U400 ( .A1(keyout[16]), .A2(n1524), .S0(n4507), .Y(n3421) );
  MUX21X1_HVT U401 ( .A1(keyout[15]), .A2(n1525), .S0(n4507), .Y(n3420) );
  MUX21X1_HVT U402 ( .A1(keyout[14]), .A2(n1526), .S0(n4507), .Y(n3419) );
  MUX21X1_HVT U403 ( .A1(keyout[13]), .A2(n1527), .S0(n4507), .Y(n3418) );
  MUX21X1_HVT U404 ( .A1(keyout[12]), .A2(n1528), .S0(n4507), .Y(n3417) );
  MUX21X1_HVT U405 ( .A1(keyout[11]), .A2(n1529), .S0(n4507), .Y(n3416) );
  MUX21X1_HVT U406 ( .A1(keyout[10]), .A2(n1530), .S0(n4507), .Y(n3415) );
  MUX21X1_HVT U407 ( .A1(keyout[9]), .A2(n1531), .S0(n4507), .Y(n3414) );
  MUX21X1_HVT U408 ( .A1(keyout[8]), .A2(n1532), .S0(n4507), .Y(n3413) );
  MUX21X1_HVT U409 ( .A1(keyout[7]), .A2(n1533), .S0(n4507), .Y(n3412) );
  MUX21X1_HVT U410 ( .A1(keyout[6]), .A2(n1534), .S0(n4507), .Y(n3411) );
  MUX21X1_HVT U411 ( .A1(keyout[5]), .A2(n1535), .S0(n4507), .Y(n3410) );
  MUX21X1_HVT U412 ( .A1(keyout[4]), .A2(n1536), .S0(n4507), .Y(n3409) );
  MUX21X1_HVT U413 ( .A1(keyout[3]), .A2(n1537), .S0(n4507), .Y(n3408) );
  MUX21X1_HVT U414 ( .A1(keyout[2]), .A2(n1538), .S0(n4507), .Y(n3407) );
  MUX21X1_HVT U415 ( .A1(keyout[1]), .A2(n1539), .S0(n4507), .Y(n3406) );
  MUX21X1_HVT U416 ( .A1(keyout[0]), .A2(n1540), .S0(n4507), .Y(n3405) );
  NAND4X0_HVT U417 ( .A1(n4535), .A2(n4511), .A3(n1), .A4(n2), .Y(n4507) );
  MUX21X1_HVT U418 ( .A1(keyout[127]), .A2(n3982), .S0(n4509), .Y(n3404) );
  MUX21X1_HVT U419 ( .A1(keyout[126]), .A2(n3983), .S0(n4509), .Y(n3403) );
  MUX21X1_HVT U420 ( .A1(keyout[125]), .A2(n3984), .S0(n4509), .Y(n3402) );
  MUX21X1_HVT U421 ( .A1(keyout[124]), .A2(n3985), .S0(n4509), .Y(n3401) );
  MUX21X1_HVT U422 ( .A1(keyout[123]), .A2(n3986), .S0(n4509), .Y(n3400) );
  MUX21X1_HVT U423 ( .A1(keyout[122]), .A2(n3987), .S0(n4509), .Y(n3399) );
  MUX21X1_HVT U424 ( .A1(keyout[121]), .A2(n3988), .S0(n4509), .Y(n3398) );
  MUX21X1_HVT U425 ( .A1(keyout[120]), .A2(n3989), .S0(n4509), .Y(n3397) );
  MUX21X1_HVT U426 ( .A1(keyout[119]), .A2(n3990), .S0(n4509), .Y(n3396) );
  MUX21X1_HVT U427 ( .A1(keyout[118]), .A2(n3991), .S0(n4509), .Y(n3395) );
  MUX21X1_HVT U428 ( .A1(keyout[117]), .A2(n3992), .S0(n4509), .Y(n3394) );
  MUX21X1_HVT U429 ( .A1(keyout[116]), .A2(n3993), .S0(n4509), .Y(n3393) );
  MUX21X1_HVT U430 ( .A1(keyout[115]), .A2(n3994), .S0(n4509), .Y(n3392) );
  MUX21X1_HVT U431 ( .A1(keyout[114]), .A2(n3995), .S0(n4509), .Y(n3391) );
  MUX21X1_HVT U432 ( .A1(keyout[113]), .A2(n3996), .S0(n4509), .Y(n3390) );
  MUX21X1_HVT U433 ( .A1(keyout[112]), .A2(n3997), .S0(n4509), .Y(n3389) );
  MUX21X1_HVT U434 ( .A1(keyout[111]), .A2(n3998), .S0(n4509), .Y(n3388) );
  MUX21X1_HVT U435 ( .A1(keyout[110]), .A2(n3999), .S0(n4509), .Y(n3387) );
  MUX21X1_HVT U436 ( .A1(keyout[109]), .A2(n4000), .S0(n4509), .Y(n3386) );
  MUX21X1_HVT U437 ( .A1(keyout[108]), .A2(n4001), .S0(n4509), .Y(n3385) );
  MUX21X1_HVT U438 ( .A1(keyout[107]), .A2(n4002), .S0(n4509), .Y(n3384) );
  MUX21X1_HVT U439 ( .A1(keyout[106]), .A2(n4003), .S0(n4509), .Y(n3383) );
  MUX21X1_HVT U440 ( .A1(keyout[105]), .A2(n4004), .S0(n4509), .Y(n3382) );
  MUX21X1_HVT U441 ( .A1(keyout[104]), .A2(n4005), .S0(n4509), .Y(n3381) );
  MUX21X1_HVT U442 ( .A1(keyout[103]), .A2(n4006), .S0(n4509), .Y(n3380) );
  MUX21X1_HVT U443 ( .A1(keyout[102]), .A2(n4007), .S0(n4509), .Y(n3379) );
  MUX21X1_HVT U444 ( .A1(keyout[101]), .A2(n4008), .S0(n4509), .Y(n3378) );
  MUX21X1_HVT U445 ( .A1(keyout[100]), .A2(n4009), .S0(n4509), .Y(n3377) );
  MUX21X1_HVT U446 ( .A1(keyout[99]), .A2(n4010), .S0(n4509), .Y(n3376) );
  MUX21X1_HVT U447 ( .A1(keyout[98]), .A2(n4011), .S0(n4509), .Y(n3375) );
  MUX21X1_HVT U448 ( .A1(keyout[97]), .A2(n4012), .S0(n4509), .Y(n3374) );
  MUX21X1_HVT U449 ( .A1(keyout[96]), .A2(n4013), .S0(n4509), .Y(n3373) );
  MUX21X1_HVT U450 ( .A1(keyout[95]), .A2(n4014), .S0(n4509), .Y(n3372) );
  MUX21X1_HVT U451 ( .A1(keyout[94]), .A2(n4015), .S0(n4509), .Y(n3371) );
  MUX21X1_HVT U452 ( .A1(keyout[93]), .A2(n4016), .S0(n4509), .Y(n3370) );
  MUX21X1_HVT U453 ( .A1(keyout[92]), .A2(n4017), .S0(n4509), .Y(n3369) );
  MUX21X1_HVT U454 ( .A1(keyout[91]), .A2(n4018), .S0(n4509), .Y(n3368) );
  MUX21X1_HVT U455 ( .A1(keyout[90]), .A2(n4019), .S0(n4509), .Y(n3367) );
  MUX21X1_HVT U456 ( .A1(keyout[89]), .A2(n4020), .S0(n4509), .Y(n3366) );
  MUX21X1_HVT U457 ( .A1(keyout[88]), .A2(n4021), .S0(n4509), .Y(n3365) );
  MUX21X1_HVT U458 ( .A1(keyout[87]), .A2(n4022), .S0(n4509), .Y(n3364) );
  MUX21X1_HVT U459 ( .A1(keyout[86]), .A2(n4023), .S0(n4509), .Y(n3363) );
  MUX21X1_HVT U460 ( .A1(keyout[85]), .A2(n4024), .S0(n4509), .Y(n3362) );
  MUX21X1_HVT U461 ( .A1(keyout[84]), .A2(n4025), .S0(n4509), .Y(n3361) );
  MUX21X1_HVT U462 ( .A1(keyout[83]), .A2(n4026), .S0(n4509), .Y(n3360) );
  MUX21X1_HVT U463 ( .A1(keyout[82]), .A2(n4027), .S0(n4509), .Y(n3359) );
  MUX21X1_HVT U464 ( .A1(keyout[81]), .A2(n4028), .S0(n4509), .Y(n3358) );
  MUX21X1_HVT U465 ( .A1(keyout[80]), .A2(n4029), .S0(n4509), .Y(n3357) );
  MUX21X1_HVT U466 ( .A1(keyout[79]), .A2(n4030), .S0(n4509), .Y(n3356) );
  MUX21X1_HVT U467 ( .A1(keyout[78]), .A2(n4031), .S0(n4509), .Y(n3355) );
  MUX21X1_HVT U468 ( .A1(keyout[77]), .A2(n4032), .S0(n4509), .Y(n3354) );
  MUX21X1_HVT U469 ( .A1(keyout[76]), .A2(n4033), .S0(n4509), .Y(n3353) );
  MUX21X1_HVT U470 ( .A1(keyout[75]), .A2(n4034), .S0(n4509), .Y(n3352) );
  MUX21X1_HVT U471 ( .A1(keyout[74]), .A2(n4035), .S0(n4509), .Y(n3351) );
  MUX21X1_HVT U472 ( .A1(keyout[73]), .A2(n4036), .S0(n4509), .Y(n3350) );
  MUX21X1_HVT U473 ( .A1(keyout[72]), .A2(n4037), .S0(n4509), .Y(n3349) );
  MUX21X1_HVT U474 ( .A1(keyout[71]), .A2(n4038), .S0(n4509), .Y(n3348) );
  MUX21X1_HVT U475 ( .A1(keyout[70]), .A2(n4039), .S0(n4509), .Y(n3347) );
  MUX21X1_HVT U476 ( .A1(keyout[69]), .A2(n4040), .S0(n4509), .Y(n3346) );
  MUX21X1_HVT U477 ( .A1(keyout[68]), .A2(n4041), .S0(n4509), .Y(n3345) );
  MUX21X1_HVT U478 ( .A1(keyout[67]), .A2(n4042), .S0(n4509), .Y(n3344) );
  MUX21X1_HVT U479 ( .A1(keyout[66]), .A2(n4043), .S0(n4509), .Y(n3343) );
  MUX21X1_HVT U480 ( .A1(keyout[65]), .A2(n4044), .S0(n4509), .Y(n3342) );
  MUX21X1_HVT U481 ( .A1(keyout[64]), .A2(n4045), .S0(n4509), .Y(n3341) );
  MUX21X1_HVT U482 ( .A1(keyout[63]), .A2(n4046), .S0(n4509), .Y(n3340) );
  MUX21X1_HVT U483 ( .A1(keyout[62]), .A2(n4047), .S0(n4509), .Y(n3339) );
  MUX21X1_HVT U484 ( .A1(keyout[61]), .A2(n4048), .S0(n4509), .Y(n3338) );
  MUX21X1_HVT U485 ( .A1(keyout[60]), .A2(n4049), .S0(n4509), .Y(n3337) );
  MUX21X1_HVT U486 ( .A1(keyout[59]), .A2(n4050), .S0(n4509), .Y(n3336) );
  MUX21X1_HVT U487 ( .A1(keyout[58]), .A2(n4051), .S0(n4509), .Y(n3335) );
  MUX21X1_HVT U488 ( .A1(keyout[57]), .A2(n4052), .S0(n4509), .Y(n3334) );
  MUX21X1_HVT U489 ( .A1(keyout[56]), .A2(n4053), .S0(n4509), .Y(n3333) );
  MUX21X1_HVT U490 ( .A1(keyout[55]), .A2(n4054), .S0(n4509), .Y(n3332) );
  MUX21X1_HVT U491 ( .A1(keyout[54]), .A2(n4055), .S0(n4509), .Y(n3331) );
  MUX21X1_HVT U492 ( .A1(keyout[53]), .A2(n4056), .S0(n4509), .Y(n3330) );
  MUX21X1_HVT U493 ( .A1(keyout[52]), .A2(n4057), .S0(n4509), .Y(n3329) );
  MUX21X1_HVT U494 ( .A1(keyout[51]), .A2(n4058), .S0(n4509), .Y(n3328) );
  MUX21X1_HVT U495 ( .A1(keyout[50]), .A2(n4059), .S0(n4509), .Y(n3327) );
  MUX21X1_HVT U496 ( .A1(keyout[49]), .A2(n4060), .S0(n4509), .Y(n3326) );
  MUX21X1_HVT U497 ( .A1(keyout[48]), .A2(n4061), .S0(n4509), .Y(n3325) );
  MUX21X1_HVT U498 ( .A1(keyout[47]), .A2(n4062), .S0(n4509), .Y(n3324) );
  MUX21X1_HVT U499 ( .A1(keyout[46]), .A2(n4063), .S0(n4509), .Y(n3323) );
  MUX21X1_HVT U500 ( .A1(keyout[45]), .A2(n4064), .S0(n4509), .Y(n3322) );
  MUX21X1_HVT U501 ( .A1(keyout[44]), .A2(n4065), .S0(n4509), .Y(n3321) );
  MUX21X1_HVT U502 ( .A1(keyout[43]), .A2(n4066), .S0(n4509), .Y(n3320) );
  MUX21X1_HVT U503 ( .A1(keyout[42]), .A2(n4067), .S0(n4509), .Y(n3319) );
  MUX21X1_HVT U504 ( .A1(keyout[41]), .A2(n4068), .S0(n4509), .Y(n3318) );
  MUX21X1_HVT U505 ( .A1(keyout[40]), .A2(n4069), .S0(n4509), .Y(n3317) );
  MUX21X1_HVT U506 ( .A1(keyout[39]), .A2(n4070), .S0(n4509), .Y(n3316) );
  MUX21X1_HVT U507 ( .A1(keyout[38]), .A2(n4071), .S0(n4509), .Y(n3315) );
  MUX21X1_HVT U508 ( .A1(keyout[37]), .A2(n4072), .S0(n4509), .Y(n3314) );
  MUX21X1_HVT U509 ( .A1(keyout[36]), .A2(n4073), .S0(n4509), .Y(n3313) );
  MUX21X1_HVT U510 ( .A1(keyout[35]), .A2(n4074), .S0(n4509), .Y(n3312) );
  MUX21X1_HVT U511 ( .A1(keyout[34]), .A2(n4075), .S0(n4509), .Y(n3311) );
  MUX21X1_HVT U512 ( .A1(keyout[33]), .A2(n4076), .S0(n4509), .Y(n3310) );
  MUX21X1_HVT U513 ( .A1(keyout[32]), .A2(n4077), .S0(n4509), .Y(n3309) );
  MUX21X1_HVT U514 ( .A1(keyout[31]), .A2(n4078), .S0(n4509), .Y(n3308) );
  MUX21X1_HVT U515 ( .A1(keyout[30]), .A2(n4079), .S0(n4509), .Y(n3307) );
  MUX21X1_HVT U516 ( .A1(keyout[29]), .A2(n4080), .S0(n4509), .Y(n3306) );
  MUX21X1_HVT U517 ( .A1(keyout[28]), .A2(n4081), .S0(n4509), .Y(n3305) );
  MUX21X1_HVT U518 ( .A1(keyout[27]), .A2(n4082), .S0(n4509), .Y(n3304) );
  MUX21X1_HVT U519 ( .A1(keyout[26]), .A2(n4083), .S0(n4509), .Y(n3303) );
  MUX21X1_HVT U520 ( .A1(keyout[25]), .A2(n4084), .S0(n4509), .Y(n3302) );
  MUX21X1_HVT U521 ( .A1(keyout[24]), .A2(n4085), .S0(n4509), .Y(n3301) );
  MUX21X1_HVT U522 ( .A1(keyout[23]), .A2(n4086), .S0(n4509), .Y(n3300) );
  MUX21X1_HVT U523 ( .A1(keyout[22]), .A2(n4087), .S0(n4509), .Y(n3299) );
  MUX21X1_HVT U524 ( .A1(keyout[21]), .A2(n4088), .S0(n4509), .Y(n3298) );
  MUX21X1_HVT U525 ( .A1(keyout[20]), .A2(n4089), .S0(n4509), .Y(n3297) );
  MUX21X1_HVT U526 ( .A1(keyout[19]), .A2(n4090), .S0(n4509), .Y(n3296) );
  MUX21X1_HVT U527 ( .A1(keyout[18]), .A2(n4091), .S0(n4509), .Y(n3295) );
  MUX21X1_HVT U528 ( .A1(keyout[17]), .A2(n4092), .S0(n4509), .Y(n3294) );
  MUX21X1_HVT U529 ( .A1(keyout[16]), .A2(n4093), .S0(n4509), .Y(n3293) );
  MUX21X1_HVT U530 ( .A1(keyout[15]), .A2(n4094), .S0(n4509), .Y(n3292) );
  MUX21X1_HVT U531 ( .A1(keyout[14]), .A2(n4095), .S0(n4509), .Y(n3291) );
  MUX21X1_HVT U532 ( .A1(keyout[13]), .A2(n4096), .S0(n4509), .Y(n3290) );
  MUX21X1_HVT U533 ( .A1(keyout[12]), .A2(n4097), .S0(n4509), .Y(n3289) );
  MUX21X1_HVT U534 ( .A1(keyout[11]), .A2(n4098), .S0(n4509), .Y(n3288) );
  MUX21X1_HVT U535 ( .A1(keyout[10]), .A2(n4099), .S0(n4509), .Y(n3287) );
  MUX21X1_HVT U536 ( .A1(keyout[9]), .A2(n4100), .S0(n4509), .Y(n3286) );
  MUX21X1_HVT U537 ( .A1(keyout[8]), .A2(n4101), .S0(n4509), .Y(n3285) );
  MUX21X1_HVT U538 ( .A1(keyout[7]), .A2(n4102), .S0(n4509), .Y(n3284) );
  MUX21X1_HVT U539 ( .A1(keyout[6]), .A2(n4103), .S0(n4509), .Y(n3283) );
  MUX21X1_HVT U540 ( .A1(keyout[5]), .A2(n4104), .S0(n4509), .Y(n3282) );
  MUX21X1_HVT U541 ( .A1(keyout[4]), .A2(n4105), .S0(n4509), .Y(n3281) );
  MUX21X1_HVT U542 ( .A1(keyout[3]), .A2(n4106), .S0(n4509), .Y(n3280) );
  MUX21X1_HVT U543 ( .A1(keyout[2]), .A2(n4107), .S0(n4509), .Y(n3279) );
  MUX21X1_HVT U544 ( .A1(keyout[1]), .A2(n4108), .S0(n4509), .Y(n3278) );
  MUX21X1_HVT U545 ( .A1(keyout[0]), .A2(n4109), .S0(n4509), .Y(n3277) );
  OR2X1_HVT U546 ( .A1(n4518), .A2(rest), .Y(n4509) );
  NAND3X0_HVT U547 ( .A1(n4535), .A2(n2), .A3(state[0]), .Y(n4518) );
  MUX21X1_HVT U548 ( .A1(keyout[127]), .A2(n1669), .S0(n4496), .Y(n3276) );
  MUX21X1_HVT U549 ( .A1(keyout[126]), .A2(n1670), .S0(n4496), .Y(n3275) );
  MUX21X1_HVT U550 ( .A1(keyout[125]), .A2(n1671), .S0(n4496), .Y(n3274) );
  MUX21X1_HVT U551 ( .A1(keyout[124]), .A2(n1672), .S0(n4496), .Y(n3273) );
  MUX21X1_HVT U552 ( .A1(keyout[123]), .A2(n1673), .S0(n4496), .Y(n3272) );
  MUX21X1_HVT U553 ( .A1(keyout[122]), .A2(n1674), .S0(n4496), .Y(n3271) );
  MUX21X1_HVT U554 ( .A1(keyout[121]), .A2(n1675), .S0(n4496), .Y(n3270) );
  MUX21X1_HVT U555 ( .A1(keyout[120]), .A2(n1676), .S0(n4496), .Y(n3269) );
  MUX21X1_HVT U556 ( .A1(keyout[119]), .A2(n1677), .S0(n4496), .Y(n3268) );
  MUX21X1_HVT U557 ( .A1(keyout[118]), .A2(n1678), .S0(n4496), .Y(n3267) );
  MUX21X1_HVT U558 ( .A1(keyout[117]), .A2(n1679), .S0(n4496), .Y(n3266) );
  MUX21X1_HVT U559 ( .A1(keyout[116]), .A2(n1680), .S0(n4496), .Y(n3265) );
  MUX21X1_HVT U560 ( .A1(keyout[115]), .A2(n1681), .S0(n4496), .Y(n3264) );
  MUX21X1_HVT U561 ( .A1(keyout[114]), .A2(n1682), .S0(n4496), .Y(n3263) );
  MUX21X1_HVT U562 ( .A1(keyout[113]), .A2(n1683), .S0(n4496), .Y(n3262) );
  MUX21X1_HVT U563 ( .A1(keyout[112]), .A2(n1684), .S0(n4496), .Y(n3261) );
  MUX21X1_HVT U564 ( .A1(keyout[111]), .A2(n1685), .S0(n4496), .Y(n3260) );
  MUX21X1_HVT U565 ( .A1(keyout[110]), .A2(n1686), .S0(n4496), .Y(n3259) );
  MUX21X1_HVT U566 ( .A1(keyout[109]), .A2(n1687), .S0(n4496), .Y(n3258) );
  MUX21X1_HVT U567 ( .A1(keyout[108]), .A2(n1688), .S0(n4496), .Y(n3257) );
  MUX21X1_HVT U568 ( .A1(keyout[107]), .A2(n1689), .S0(n4496), .Y(n3256) );
  MUX21X1_HVT U569 ( .A1(keyout[106]), .A2(n1690), .S0(n4496), .Y(n3255) );
  MUX21X1_HVT U570 ( .A1(keyout[105]), .A2(n1691), .S0(n4496), .Y(n3254) );
  MUX21X1_HVT U571 ( .A1(keyout[104]), .A2(n1692), .S0(n4496), .Y(n3253) );
  MUX21X1_HVT U572 ( .A1(keyout[103]), .A2(n1693), .S0(n4496), .Y(n3252) );
  MUX21X1_HVT U573 ( .A1(keyout[102]), .A2(n1694), .S0(n4496), .Y(n3251) );
  MUX21X1_HVT U574 ( .A1(keyout[101]), .A2(n1695), .S0(n4496), .Y(n3250) );
  MUX21X1_HVT U575 ( .A1(keyout[100]), .A2(n1696), .S0(n4496), .Y(n3249) );
  MUX21X1_HVT U576 ( .A1(keyout[99]), .A2(n1697), .S0(n4496), .Y(n3248) );
  MUX21X1_HVT U577 ( .A1(keyout[98]), .A2(n1698), .S0(n4496), .Y(n3247) );
  MUX21X1_HVT U578 ( .A1(keyout[97]), .A2(n1699), .S0(n4496), .Y(n3246) );
  MUX21X1_HVT U579 ( .A1(keyout[96]), .A2(n1700), .S0(n4496), .Y(n3245) );
  MUX21X1_HVT U580 ( .A1(keyout[95]), .A2(n1701), .S0(n4496), .Y(n3244) );
  MUX21X1_HVT U581 ( .A1(keyout[94]), .A2(n1702), .S0(n4496), .Y(n3243) );
  MUX21X1_HVT U582 ( .A1(keyout[93]), .A2(n1703), .S0(n4496), .Y(n3242) );
  MUX21X1_HVT U583 ( .A1(keyout[92]), .A2(n1704), .S0(n4496), .Y(n3241) );
  MUX21X1_HVT U584 ( .A1(keyout[91]), .A2(n1705), .S0(n4496), .Y(n3240) );
  MUX21X1_HVT U585 ( .A1(keyout[90]), .A2(n1706), .S0(n4496), .Y(n3239) );
  MUX21X1_HVT U586 ( .A1(keyout[89]), .A2(n1707), .S0(n4496), .Y(n3238) );
  MUX21X1_HVT U587 ( .A1(keyout[88]), .A2(n1708), .S0(n4496), .Y(n3237) );
  MUX21X1_HVT U588 ( .A1(keyout[87]), .A2(n1709), .S0(n4496), .Y(n3236) );
  MUX21X1_HVT U589 ( .A1(keyout[86]), .A2(n1710), .S0(n4496), .Y(n3235) );
  MUX21X1_HVT U590 ( .A1(keyout[85]), .A2(n1711), .S0(n4496), .Y(n3234) );
  MUX21X1_HVT U591 ( .A1(keyout[84]), .A2(n1712), .S0(n4496), .Y(n3233) );
  MUX21X1_HVT U592 ( .A1(keyout[83]), .A2(n1713), .S0(n4496), .Y(n3232) );
  MUX21X1_HVT U593 ( .A1(keyout[82]), .A2(n1714), .S0(n4496), .Y(n3231) );
  MUX21X1_HVT U594 ( .A1(keyout[81]), .A2(n1715), .S0(n4496), .Y(n3230) );
  MUX21X1_HVT U595 ( .A1(keyout[80]), .A2(n1716), .S0(n4496), .Y(n3229) );
  MUX21X1_HVT U596 ( .A1(keyout[79]), .A2(n1717), .S0(n4496), .Y(n3228) );
  MUX21X1_HVT U597 ( .A1(keyout[78]), .A2(n1718), .S0(n4496), .Y(n3227) );
  MUX21X1_HVT U598 ( .A1(keyout[77]), .A2(n1719), .S0(n4496), .Y(n3226) );
  MUX21X1_HVT U599 ( .A1(keyout[76]), .A2(n1720), .S0(n4496), .Y(n3225) );
  MUX21X1_HVT U600 ( .A1(keyout[75]), .A2(n1721), .S0(n4496), .Y(n3224) );
  MUX21X1_HVT U601 ( .A1(keyout[74]), .A2(n1722), .S0(n4496), .Y(n3223) );
  MUX21X1_HVT U602 ( .A1(keyout[73]), .A2(n1723), .S0(n4496), .Y(n3222) );
  MUX21X1_HVT U603 ( .A1(keyout[72]), .A2(n1724), .S0(n4496), .Y(n3221) );
  MUX21X1_HVT U604 ( .A1(keyout[71]), .A2(n1725), .S0(n4496), .Y(n3220) );
  MUX21X1_HVT U605 ( .A1(keyout[70]), .A2(n1726), .S0(n4496), .Y(n3219) );
  MUX21X1_HVT U606 ( .A1(keyout[69]), .A2(n1727), .S0(n4496), .Y(n3218) );
  MUX21X1_HVT U607 ( .A1(keyout[68]), .A2(n1728), .S0(n4496), .Y(n3217) );
  MUX21X1_HVT U608 ( .A1(keyout[67]), .A2(n1729), .S0(n4496), .Y(n3216) );
  MUX21X1_HVT U609 ( .A1(keyout[66]), .A2(n1730), .S0(n4496), .Y(n3215) );
  MUX21X1_HVT U610 ( .A1(keyout[65]), .A2(n1731), .S0(n4496), .Y(n3214) );
  MUX21X1_HVT U611 ( .A1(keyout[64]), .A2(n1732), .S0(n4496), .Y(n3213) );
  MUX21X1_HVT U612 ( .A1(keyout[63]), .A2(n1733), .S0(n4496), .Y(n3212) );
  MUX21X1_HVT U613 ( .A1(keyout[62]), .A2(n1734), .S0(n4496), .Y(n3211) );
  MUX21X1_HVT U614 ( .A1(keyout[61]), .A2(n1735), .S0(n4496), .Y(n3210) );
  MUX21X1_HVT U615 ( .A1(keyout[60]), .A2(n1736), .S0(n4496), .Y(n3209) );
  MUX21X1_HVT U616 ( .A1(keyout[59]), .A2(n1737), .S0(n4496), .Y(n3208) );
  MUX21X1_HVT U617 ( .A1(keyout[58]), .A2(n1738), .S0(n4496), .Y(n3207) );
  MUX21X1_HVT U618 ( .A1(keyout[57]), .A2(n1739), .S0(n4496), .Y(n3206) );
  MUX21X1_HVT U619 ( .A1(keyout[56]), .A2(n1740), .S0(n4496), .Y(n3205) );
  MUX21X1_HVT U620 ( .A1(keyout[55]), .A2(n1741), .S0(n4496), .Y(n3204) );
  MUX21X1_HVT U621 ( .A1(keyout[54]), .A2(n1742), .S0(n4496), .Y(n3203) );
  MUX21X1_HVT U622 ( .A1(keyout[53]), .A2(n1743), .S0(n4496), .Y(n3202) );
  MUX21X1_HVT U623 ( .A1(keyout[52]), .A2(n1744), .S0(n4496), .Y(n3201) );
  MUX21X1_HVT U624 ( .A1(keyout[51]), .A2(n1745), .S0(n4496), .Y(n3200) );
  MUX21X1_HVT U625 ( .A1(keyout[50]), .A2(n1746), .S0(n4496), .Y(n3199) );
  MUX21X1_HVT U626 ( .A1(keyout[49]), .A2(n1747), .S0(n4496), .Y(n3198) );
  MUX21X1_HVT U627 ( .A1(keyout[48]), .A2(n1748), .S0(n4496), .Y(n3197) );
  MUX21X1_HVT U628 ( .A1(keyout[47]), .A2(n1749), .S0(n4496), .Y(n3196) );
  MUX21X1_HVT U629 ( .A1(keyout[46]), .A2(n1750), .S0(n4496), .Y(n3195) );
  MUX21X1_HVT U630 ( .A1(keyout[45]), .A2(n1751), .S0(n4496), .Y(n3194) );
  MUX21X1_HVT U631 ( .A1(keyout[44]), .A2(n1752), .S0(n4496), .Y(n3193) );
  MUX21X1_HVT U632 ( .A1(keyout[43]), .A2(n1753), .S0(n4496), .Y(n3192) );
  MUX21X1_HVT U633 ( .A1(keyout[42]), .A2(n1754), .S0(n4496), .Y(n3191) );
  MUX21X1_HVT U634 ( .A1(keyout[41]), .A2(n1755), .S0(n4496), .Y(n3190) );
  MUX21X1_HVT U635 ( .A1(keyout[40]), .A2(n1756), .S0(n4496), .Y(n3189) );
  MUX21X1_HVT U636 ( .A1(keyout[39]), .A2(n1757), .S0(n4496), .Y(n3188) );
  MUX21X1_HVT U637 ( .A1(keyout[38]), .A2(n1758), .S0(n4496), .Y(n3187) );
  MUX21X1_HVT U638 ( .A1(keyout[37]), .A2(n1759), .S0(n4496), .Y(n3186) );
  MUX21X1_HVT U639 ( .A1(keyout[36]), .A2(n1760), .S0(n4496), .Y(n3185) );
  MUX21X1_HVT U640 ( .A1(keyout[35]), .A2(n1761), .S0(n4496), .Y(n3184) );
  MUX21X1_HVT U641 ( .A1(keyout[34]), .A2(n1762), .S0(n4496), .Y(n3183) );
  MUX21X1_HVT U642 ( .A1(keyout[33]), .A2(n1763), .S0(n4496), .Y(n3182) );
  MUX21X1_HVT U643 ( .A1(keyout[32]), .A2(n1764), .S0(n4496), .Y(n3181) );
  MUX21X1_HVT U644 ( .A1(keyout[31]), .A2(n1765), .S0(n4496), .Y(n3180) );
  MUX21X1_HVT U645 ( .A1(keyout[30]), .A2(n1766), .S0(n4496), .Y(n3179) );
  MUX21X1_HVT U646 ( .A1(keyout[29]), .A2(n1767), .S0(n4496), .Y(n3178) );
  MUX21X1_HVT U647 ( .A1(keyout[28]), .A2(n1768), .S0(n4496), .Y(n3177) );
  MUX21X1_HVT U648 ( .A1(keyout[27]), .A2(n1769), .S0(n4496), .Y(n3176) );
  MUX21X1_HVT U649 ( .A1(keyout[26]), .A2(n1770), .S0(n4496), .Y(n3175) );
  MUX21X1_HVT U650 ( .A1(keyout[25]), .A2(n1771), .S0(n4496), .Y(n3174) );
  MUX21X1_HVT U651 ( .A1(keyout[24]), .A2(n1772), .S0(n4496), .Y(n3173) );
  MUX21X1_HVT U652 ( .A1(keyout[23]), .A2(n1773), .S0(n4496), .Y(n3172) );
  MUX21X1_HVT U653 ( .A1(keyout[22]), .A2(n1774), .S0(n4496), .Y(n3171) );
  MUX21X1_HVT U654 ( .A1(keyout[21]), .A2(n1775), .S0(n4496), .Y(n3170) );
  MUX21X1_HVT U655 ( .A1(keyout[20]), .A2(n1776), .S0(n4496), .Y(n3169) );
  MUX21X1_HVT U656 ( .A1(keyout[19]), .A2(n1777), .S0(n4496), .Y(n3168) );
  MUX21X1_HVT U657 ( .A1(keyout[18]), .A2(n1778), .S0(n4496), .Y(n3167) );
  MUX21X1_HVT U658 ( .A1(keyout[17]), .A2(n1779), .S0(n4496), .Y(n3166) );
  MUX21X1_HVT U659 ( .A1(keyout[16]), .A2(n1780), .S0(n4496), .Y(n3165) );
  MUX21X1_HVT U660 ( .A1(keyout[15]), .A2(n1781), .S0(n4496), .Y(n3164) );
  MUX21X1_HVT U661 ( .A1(keyout[14]), .A2(n1782), .S0(n4496), .Y(n3163) );
  MUX21X1_HVT U662 ( .A1(keyout[13]), .A2(n1783), .S0(n4496), .Y(n3162) );
  MUX21X1_HVT U663 ( .A1(keyout[12]), .A2(n1784), .S0(n4496), .Y(n3161) );
  MUX21X1_HVT U664 ( .A1(keyout[11]), .A2(n1785), .S0(n4496), .Y(n3160) );
  MUX21X1_HVT U665 ( .A1(keyout[10]), .A2(n1786), .S0(n4496), .Y(n3159) );
  MUX21X1_HVT U666 ( .A1(keyout[9]), .A2(n1787), .S0(n4496), .Y(n3158) );
  MUX21X1_HVT U667 ( .A1(keyout[8]), .A2(n1788), .S0(n4496), .Y(n3157) );
  MUX21X1_HVT U668 ( .A1(keyout[7]), .A2(n1789), .S0(n4496), .Y(n3156) );
  MUX21X1_HVT U669 ( .A1(keyout[6]), .A2(n1790), .S0(n4496), .Y(n3155) );
  MUX21X1_HVT U670 ( .A1(keyout[5]), .A2(n1791), .S0(n4496), .Y(n3154) );
  MUX21X1_HVT U671 ( .A1(keyout[4]), .A2(n1792), .S0(n4496), .Y(n3153) );
  MUX21X1_HVT U672 ( .A1(keyout[3]), .A2(n1793), .S0(n4496), .Y(n3152) );
  MUX21X1_HVT U673 ( .A1(keyout[2]), .A2(n1794), .S0(n4496), .Y(n3151) );
  MUX21X1_HVT U674 ( .A1(keyout[1]), .A2(n1795), .S0(n4496), .Y(n3150) );
  MUX21X1_HVT U675 ( .A1(keyout[0]), .A2(n1796), .S0(n4496), .Y(n3149) );
  OR2X1_HVT U676 ( .A1(n4523), .A2(rest), .Y(n4496) );
  NAND2X0_HVT U677 ( .A1(n4536), .A2(n1), .Y(n4523) );
  MUX21X1_HVT U678 ( .A1(keyout[127]), .A2(n2053), .S0(n4503), .Y(n3148) );
  MUX21X1_HVT U679 ( .A1(keyout[126]), .A2(n2054), .S0(n4503), .Y(n3147) );
  MUX21X1_HVT U680 ( .A1(keyout[125]), .A2(n2055), .S0(n4503), .Y(n3146) );
  MUX21X1_HVT U681 ( .A1(keyout[124]), .A2(n2056), .S0(n4503), .Y(n3145) );
  MUX21X1_HVT U682 ( .A1(keyout[123]), .A2(n2057), .S0(n4503), .Y(n3144) );
  MUX21X1_HVT U683 ( .A1(keyout[122]), .A2(n2058), .S0(n4503), .Y(n3143) );
  MUX21X1_HVT U684 ( .A1(keyout[121]), .A2(n2059), .S0(n4503), .Y(n3142) );
  MUX21X1_HVT U685 ( .A1(keyout[120]), .A2(n2060), .S0(n4503), .Y(n3141) );
  MUX21X1_HVT U686 ( .A1(keyout[119]), .A2(n2061), .S0(n4503), .Y(n3140) );
  MUX21X1_HVT U687 ( .A1(keyout[118]), .A2(n2062), .S0(n4503), .Y(n3139) );
  MUX21X1_HVT U688 ( .A1(keyout[117]), .A2(n2063), .S0(n4503), .Y(n3138) );
  MUX21X1_HVT U689 ( .A1(keyout[116]), .A2(n2064), .S0(n4503), .Y(n3137) );
  MUX21X1_HVT U690 ( .A1(keyout[115]), .A2(n2065), .S0(n4503), .Y(n3136) );
  MUX21X1_HVT U691 ( .A1(keyout[114]), .A2(n2066), .S0(n4503), .Y(n3135) );
  MUX21X1_HVT U692 ( .A1(keyout[113]), .A2(n2067), .S0(n4503), .Y(n3134) );
  MUX21X1_HVT U693 ( .A1(keyout[112]), .A2(n2068), .S0(n4503), .Y(n3133) );
  MUX21X1_HVT U694 ( .A1(keyout[111]), .A2(n2069), .S0(n4503), .Y(n3132) );
  MUX21X1_HVT U695 ( .A1(keyout[110]), .A2(n2070), .S0(n4503), .Y(n3131) );
  MUX21X1_HVT U696 ( .A1(keyout[109]), .A2(n2071), .S0(n4503), .Y(n3130) );
  MUX21X1_HVT U697 ( .A1(keyout[108]), .A2(n2072), .S0(n4503), .Y(n3129) );
  MUX21X1_HVT U698 ( .A1(keyout[107]), .A2(n2073), .S0(n4503), .Y(n3128) );
  MUX21X1_HVT U699 ( .A1(keyout[106]), .A2(n2074), .S0(n4503), .Y(n3127) );
  MUX21X1_HVT U700 ( .A1(keyout[105]), .A2(n2075), .S0(n4503), .Y(n3126) );
  MUX21X1_HVT U701 ( .A1(keyout[104]), .A2(n2076), .S0(n4503), .Y(n3125) );
  MUX21X1_HVT U702 ( .A1(keyout[103]), .A2(n2077), .S0(n4503), .Y(n3124) );
  MUX21X1_HVT U703 ( .A1(keyout[102]), .A2(n2078), .S0(n4503), .Y(n3123) );
  MUX21X1_HVT U704 ( .A1(keyout[101]), .A2(n2079), .S0(n4503), .Y(n3122) );
  MUX21X1_HVT U705 ( .A1(keyout[100]), .A2(n2080), .S0(n4503), .Y(n3121) );
  MUX21X1_HVT U706 ( .A1(keyout[99]), .A2(n2081), .S0(n4503), .Y(n3120) );
  MUX21X1_HVT U707 ( .A1(keyout[98]), .A2(n2082), .S0(n4503), .Y(n3119) );
  MUX21X1_HVT U708 ( .A1(keyout[97]), .A2(n2083), .S0(n4503), .Y(n3118) );
  MUX21X1_HVT U709 ( .A1(keyout[96]), .A2(n2084), .S0(n4503), .Y(n3117) );
  MUX21X1_HVT U710 ( .A1(keyout[95]), .A2(n2085), .S0(n4503), .Y(n3116) );
  MUX21X1_HVT U711 ( .A1(keyout[94]), .A2(n2086), .S0(n4503), .Y(n3115) );
  MUX21X1_HVT U712 ( .A1(keyout[93]), .A2(n2087), .S0(n4503), .Y(n3114) );
  MUX21X1_HVT U713 ( .A1(keyout[92]), .A2(n2088), .S0(n4503), .Y(n3113) );
  MUX21X1_HVT U714 ( .A1(keyout[91]), .A2(n2089), .S0(n4503), .Y(n3112) );
  MUX21X1_HVT U715 ( .A1(keyout[90]), .A2(n2090), .S0(n4503), .Y(n3111) );
  MUX21X1_HVT U716 ( .A1(keyout[89]), .A2(n2091), .S0(n4503), .Y(n3110) );
  MUX21X1_HVT U717 ( .A1(keyout[88]), .A2(n2092), .S0(n4503), .Y(n3109) );
  MUX21X1_HVT U718 ( .A1(keyout[87]), .A2(n2093), .S0(n4503), .Y(n3108) );
  MUX21X1_HVT U719 ( .A1(keyout[86]), .A2(n2094), .S0(n4503), .Y(n3107) );
  MUX21X1_HVT U720 ( .A1(keyout[85]), .A2(n2095), .S0(n4503), .Y(n3106) );
  MUX21X1_HVT U721 ( .A1(keyout[84]), .A2(n2096), .S0(n4503), .Y(n3105) );
  MUX21X1_HVT U722 ( .A1(keyout[83]), .A2(n2097), .S0(n4503), .Y(n3104) );
  MUX21X1_HVT U723 ( .A1(keyout[82]), .A2(n2098), .S0(n4503), .Y(n3103) );
  MUX21X1_HVT U724 ( .A1(keyout[81]), .A2(n2099), .S0(n4503), .Y(n3102) );
  MUX21X1_HVT U725 ( .A1(keyout[80]), .A2(n2100), .S0(n4503), .Y(n3101) );
  MUX21X1_HVT U726 ( .A1(keyout[79]), .A2(n2101), .S0(n4503), .Y(n3100) );
  MUX21X1_HVT U727 ( .A1(keyout[78]), .A2(n2102), .S0(n4503), .Y(n3099) );
  MUX21X1_HVT U728 ( .A1(keyout[77]), .A2(n2103), .S0(n4503), .Y(n3098) );
  MUX21X1_HVT U729 ( .A1(keyout[76]), .A2(n2104), .S0(n4503), .Y(n3097) );
  MUX21X1_HVT U730 ( .A1(keyout[75]), .A2(n2105), .S0(n4503), .Y(n3096) );
  MUX21X1_HVT U731 ( .A1(keyout[74]), .A2(n2106), .S0(n4503), .Y(n3095) );
  MUX21X1_HVT U732 ( .A1(keyout[73]), .A2(n2107), .S0(n4503), .Y(n3094) );
  MUX21X1_HVT U733 ( .A1(keyout[72]), .A2(n2108), .S0(n4503), .Y(n3093) );
  MUX21X1_HVT U734 ( .A1(keyout[71]), .A2(n2109), .S0(n4503), .Y(n3092) );
  MUX21X1_HVT U735 ( .A1(keyout[70]), .A2(n2110), .S0(n4503), .Y(n3091) );
  MUX21X1_HVT U736 ( .A1(keyout[69]), .A2(n2111), .S0(n4503), .Y(n3090) );
  MUX21X1_HVT U737 ( .A1(keyout[68]), .A2(n2112), .S0(n4503), .Y(n3089) );
  MUX21X1_HVT U738 ( .A1(keyout[67]), .A2(n2113), .S0(n4503), .Y(n3088) );
  MUX21X1_HVT U739 ( .A1(keyout[66]), .A2(n2114), .S0(n4503), .Y(n3087) );
  MUX21X1_HVT U740 ( .A1(keyout[65]), .A2(n2115), .S0(n4503), .Y(n3086) );
  MUX21X1_HVT U741 ( .A1(keyout[64]), .A2(n2116), .S0(n4503), .Y(n3085) );
  MUX21X1_HVT U742 ( .A1(keyout[63]), .A2(n2117), .S0(n4503), .Y(n3084) );
  MUX21X1_HVT U743 ( .A1(keyout[62]), .A2(n2118), .S0(n4503), .Y(n3083) );
  MUX21X1_HVT U744 ( .A1(keyout[61]), .A2(n2119), .S0(n4503), .Y(n3082) );
  MUX21X1_HVT U745 ( .A1(keyout[60]), .A2(n2120), .S0(n4503), .Y(n3081) );
  MUX21X1_HVT U746 ( .A1(keyout[59]), .A2(n2121), .S0(n4503), .Y(n3080) );
  MUX21X1_HVT U747 ( .A1(keyout[58]), .A2(n2122), .S0(n4503), .Y(n3079) );
  MUX21X1_HVT U748 ( .A1(keyout[57]), .A2(n2123), .S0(n4503), .Y(n3078) );
  MUX21X1_HVT U749 ( .A1(keyout[56]), .A2(n2124), .S0(n4503), .Y(n3077) );
  MUX21X1_HVT U750 ( .A1(keyout[55]), .A2(n3798), .S0(n4503), .Y(n3076) );
  MUX21X1_HVT U751 ( .A1(keyout[54]), .A2(n3799), .S0(n4503), .Y(n3075) );
  MUX21X1_HVT U752 ( .A1(keyout[53]), .A2(n3800), .S0(n4503), .Y(n3074) );
  MUX21X1_HVT U753 ( .A1(keyout[52]), .A2(n3801), .S0(n4503), .Y(n3073) );
  MUX21X1_HVT U754 ( .A1(keyout[51]), .A2(n3802), .S0(n4503), .Y(n3072) );
  MUX21X1_HVT U755 ( .A1(keyout[50]), .A2(n3803), .S0(n4503), .Y(n3071) );
  MUX21X1_HVT U756 ( .A1(keyout[49]), .A2(n3804), .S0(n4503), .Y(n3070) );
  MUX21X1_HVT U757 ( .A1(keyout[48]), .A2(n3805), .S0(n4503), .Y(n3069) );
  MUX21X1_HVT U758 ( .A1(keyout[47]), .A2(n3806), .S0(n4503), .Y(n3068) );
  MUX21X1_HVT U759 ( .A1(keyout[46]), .A2(n3807), .S0(n4503), .Y(n3067) );
  MUX21X1_HVT U760 ( .A1(keyout[45]), .A2(n3808), .S0(n4503), .Y(n3066) );
  MUX21X1_HVT U761 ( .A1(keyout[44]), .A2(n3809), .S0(n4503), .Y(n3065) );
  MUX21X1_HVT U762 ( .A1(keyout[43]), .A2(n3810), .S0(n4503), .Y(n3064) );
  MUX21X1_HVT U763 ( .A1(keyout[42]), .A2(n3811), .S0(n4503), .Y(n3063) );
  MUX21X1_HVT U764 ( .A1(keyout[41]), .A2(n3812), .S0(n4503), .Y(n3062) );
  MUX21X1_HVT U765 ( .A1(keyout[40]), .A2(n3813), .S0(n4503), .Y(n3061) );
  MUX21X1_HVT U766 ( .A1(keyout[39]), .A2(n3814), .S0(n4503), .Y(n3060) );
  MUX21X1_HVT U767 ( .A1(keyout[38]), .A2(n3815), .S0(n4503), .Y(n3059) );
  MUX21X1_HVT U768 ( .A1(keyout[37]), .A2(n3816), .S0(n4503), .Y(n3058) );
  MUX21X1_HVT U769 ( .A1(keyout[36]), .A2(n3817), .S0(n4503), .Y(n3057) );
  MUX21X1_HVT U770 ( .A1(keyout[35]), .A2(n3818), .S0(n4503), .Y(n3056) );
  MUX21X1_HVT U771 ( .A1(keyout[34]), .A2(n3819), .S0(n4503), .Y(n3055) );
  MUX21X1_HVT U772 ( .A1(keyout[33]), .A2(n3820), .S0(n4503), .Y(n3054) );
  MUX21X1_HVT U773 ( .A1(keyout[32]), .A2(n3821), .S0(n4503), .Y(n3053) );
  MUX21X1_HVT U774 ( .A1(keyout[31]), .A2(n3822), .S0(n4503), .Y(n3052) );
  MUX21X1_HVT U775 ( .A1(keyout[30]), .A2(n3823), .S0(n4503), .Y(n3051) );
  MUX21X1_HVT U776 ( .A1(keyout[29]), .A2(n3824), .S0(n4503), .Y(n3050) );
  MUX21X1_HVT U777 ( .A1(keyout[28]), .A2(n3825), .S0(n4503), .Y(n3049) );
  MUX21X1_HVT U778 ( .A1(keyout[27]), .A2(n3826), .S0(n4503), .Y(n3048) );
  MUX21X1_HVT U779 ( .A1(keyout[26]), .A2(n3827), .S0(n4503), .Y(n3047) );
  MUX21X1_HVT U780 ( .A1(keyout[25]), .A2(n3828), .S0(n4503), .Y(n3046) );
  MUX21X1_HVT U781 ( .A1(keyout[24]), .A2(n3829), .S0(n4503), .Y(n3045) );
  MUX21X1_HVT U782 ( .A1(keyout[23]), .A2(n3830), .S0(n4503), .Y(n3044) );
  MUX21X1_HVT U783 ( .A1(keyout[22]), .A2(n3831), .S0(n4503), .Y(n3043) );
  MUX21X1_HVT U784 ( .A1(keyout[21]), .A2(n3832), .S0(n4503), .Y(n3042) );
  MUX21X1_HVT U785 ( .A1(keyout[20]), .A2(n3833), .S0(n4503), .Y(n3041) );
  MUX21X1_HVT U786 ( .A1(keyout[19]), .A2(n3834), .S0(n4503), .Y(n3040) );
  MUX21X1_HVT U787 ( .A1(keyout[18]), .A2(n3835), .S0(n4503), .Y(n3039) );
  MUX21X1_HVT U788 ( .A1(keyout[17]), .A2(n3836), .S0(n4503), .Y(n3038) );
  MUX21X1_HVT U789 ( .A1(keyout[16]), .A2(n3837), .S0(n4503), .Y(n3037) );
  MUX21X1_HVT U790 ( .A1(keyout[15]), .A2(n3838), .S0(n4503), .Y(n3036) );
  MUX21X1_HVT U791 ( .A1(keyout[14]), .A2(n3839), .S0(n4503), .Y(n3035) );
  MUX21X1_HVT U792 ( .A1(keyout[13]), .A2(n3840), .S0(n4503), .Y(n3034) );
  MUX21X1_HVT U793 ( .A1(keyout[12]), .A2(n3841), .S0(n4503), .Y(n3033) );
  MUX21X1_HVT U794 ( .A1(keyout[11]), .A2(n3842), .S0(n4503), .Y(n3032) );
  MUX21X1_HVT U795 ( .A1(keyout[10]), .A2(n3843), .S0(n4503), .Y(n3031) );
  MUX21X1_HVT U796 ( .A1(keyout[9]), .A2(n3844), .S0(n4503), .Y(n3030) );
  MUX21X1_HVT U797 ( .A1(keyout[8]), .A2(n3845), .S0(n4503), .Y(n3029) );
  MUX21X1_HVT U798 ( .A1(keyout[7]), .A2(n3846), .S0(n4503), .Y(n3028) );
  MUX21X1_HVT U799 ( .A1(keyout[6]), .A2(n3847), .S0(n4503), .Y(n3027) );
  MUX21X1_HVT U800 ( .A1(keyout[5]), .A2(n3848), .S0(n4503), .Y(n3026) );
  MUX21X1_HVT U801 ( .A1(keyout[4]), .A2(n3849), .S0(n4503), .Y(n3025) );
  MUX21X1_HVT U802 ( .A1(keyout[3]), .A2(n3850), .S0(n4503), .Y(n3024) );
  MUX21X1_HVT U803 ( .A1(keyout[2]), .A2(n3851), .S0(n4503), .Y(n3023) );
  MUX21X1_HVT U804 ( .A1(keyout[1]), .A2(n3852), .S0(n4503), .Y(n3022) );
  MUX21X1_HVT U805 ( .A1(keyout[0]), .A2(n3853), .S0(n4503), .Y(n3021) );
  OR2X1_HVT U806 ( .A1(n4525), .A2(rest), .Y(n4503) );
  NAND2X0_HVT U807 ( .A1(state[0]), .A2(n4536), .Y(n4525) );
  AND3X1_HVT U808 ( .A1(n3), .A2(n4), .A3(state[2]), .Y(n4536) );
  MUX21X1_HVT U809 ( .A1(keyout[127]), .A2(n4110), .S0(n4506), .Y(n3020) );
  MUX21X1_HVT U810 ( .A1(keyout[126]), .A2(n4111), .S0(n4506), .Y(n3019) );
  MUX21X1_HVT U811 ( .A1(keyout[125]), .A2(n4112), .S0(n4506), .Y(n3018) );
  MUX21X1_HVT U812 ( .A1(keyout[124]), .A2(n4113), .S0(n4506), .Y(n3017) );
  MUX21X1_HVT U813 ( .A1(keyout[123]), .A2(n4114), .S0(n4506), .Y(n3016) );
  MUX21X1_HVT U814 ( .A1(keyout[122]), .A2(n4115), .S0(n4506), .Y(n3015) );
  MUX21X1_HVT U815 ( .A1(keyout[121]), .A2(n4116), .S0(n4506), .Y(n3014) );
  MUX21X1_HVT U816 ( .A1(keyout[120]), .A2(n4117), .S0(n4506), .Y(n3013) );
  MUX21X1_HVT U817 ( .A1(keyout[119]), .A2(n4118), .S0(n4506), .Y(n3012) );
  MUX21X1_HVT U818 ( .A1(keyout[118]), .A2(n4119), .S0(n4506), .Y(n3011) );
  MUX21X1_HVT U819 ( .A1(keyout[117]), .A2(n4120), .S0(n4506), .Y(n3010) );
  MUX21X1_HVT U820 ( .A1(keyout[116]), .A2(n4121), .S0(n4506), .Y(n3009) );
  MUX21X1_HVT U821 ( .A1(keyout[115]), .A2(n4122), .S0(n4506), .Y(n3008) );
  MUX21X1_HVT U822 ( .A1(keyout[114]), .A2(n4123), .S0(n4506), .Y(n3007) );
  MUX21X1_HVT U823 ( .A1(keyout[113]), .A2(n4124), .S0(n4506), .Y(n3006) );
  MUX21X1_HVT U824 ( .A1(keyout[112]), .A2(n4125), .S0(n4506), .Y(n3005) );
  MUX21X1_HVT U825 ( .A1(keyout[111]), .A2(n4126), .S0(n4506), .Y(n3004) );
  MUX21X1_HVT U826 ( .A1(keyout[110]), .A2(n4127), .S0(n4506), .Y(n3003) );
  MUX21X1_HVT U827 ( .A1(keyout[109]), .A2(n4128), .S0(n4506), .Y(n3002) );
  MUX21X1_HVT U828 ( .A1(keyout[108]), .A2(n4129), .S0(n4506), .Y(n3001) );
  MUX21X1_HVT U829 ( .A1(keyout[107]), .A2(n4130), .S0(n4506), .Y(n3000) );
  MUX21X1_HVT U830 ( .A1(keyout[106]), .A2(n4131), .S0(n4506), .Y(n2999) );
  MUX21X1_HVT U831 ( .A1(keyout[105]), .A2(n4132), .S0(n4506), .Y(n2998) );
  MUX21X1_HVT U832 ( .A1(keyout[104]), .A2(n4133), .S0(n4506), .Y(n2997) );
  MUX21X1_HVT U833 ( .A1(keyout[103]), .A2(n4134), .S0(n4506), .Y(n2996) );
  MUX21X1_HVT U834 ( .A1(keyout[102]), .A2(n4135), .S0(n4506), .Y(n2995) );
  MUX21X1_HVT U835 ( .A1(keyout[101]), .A2(n4136), .S0(n4506), .Y(n2994) );
  MUX21X1_HVT U836 ( .A1(keyout[100]), .A2(n4137), .S0(n4506), .Y(n2993) );
  MUX21X1_HVT U837 ( .A1(keyout[99]), .A2(n4138), .S0(n4506), .Y(n2992) );
  MUX21X1_HVT U838 ( .A1(keyout[98]), .A2(n4139), .S0(n4506), .Y(n2991) );
  MUX21X1_HVT U839 ( .A1(keyout[97]), .A2(n4140), .S0(n4506), .Y(n2990) );
  MUX21X1_HVT U840 ( .A1(keyout[96]), .A2(n4141), .S0(n4506), .Y(n2989) );
  MUX21X1_HVT U841 ( .A1(keyout[95]), .A2(n4142), .S0(n4506), .Y(n2988) );
  MUX21X1_HVT U842 ( .A1(keyout[94]), .A2(n4143), .S0(n4506), .Y(n2987) );
  MUX21X1_HVT U843 ( .A1(keyout[93]), .A2(n4144), .S0(n4506), .Y(n2986) );
  MUX21X1_HVT U844 ( .A1(keyout[92]), .A2(n4145), .S0(n4506), .Y(n2985) );
  MUX21X1_HVT U845 ( .A1(keyout[91]), .A2(n4146), .S0(n4506), .Y(n2984) );
  MUX21X1_HVT U846 ( .A1(keyout[90]), .A2(n4147), .S0(n4506), .Y(n2983) );
  MUX21X1_HVT U847 ( .A1(keyout[89]), .A2(n4148), .S0(n4506), .Y(n2982) );
  MUX21X1_HVT U848 ( .A1(keyout[88]), .A2(n4149), .S0(n4506), .Y(n2981) );
  MUX21X1_HVT U849 ( .A1(keyout[87]), .A2(n4150), .S0(n4506), .Y(n2980) );
  MUX21X1_HVT U850 ( .A1(keyout[86]), .A2(n4151), .S0(n4506), .Y(n2979) );
  MUX21X1_HVT U851 ( .A1(keyout[85]), .A2(n4152), .S0(n4506), .Y(n2978) );
  MUX21X1_HVT U852 ( .A1(keyout[84]), .A2(n4153), .S0(n4506), .Y(n2977) );
  MUX21X1_HVT U853 ( .A1(keyout[83]), .A2(n4154), .S0(n4506), .Y(n2976) );
  MUX21X1_HVT U854 ( .A1(keyout[82]), .A2(n4155), .S0(n4506), .Y(n2975) );
  MUX21X1_HVT U855 ( .A1(keyout[81]), .A2(n4156), .S0(n4506), .Y(n2974) );
  MUX21X1_HVT U856 ( .A1(keyout[80]), .A2(n4157), .S0(n4506), .Y(n2973) );
  MUX21X1_HVT U857 ( .A1(keyout[79]), .A2(n4158), .S0(n4506), .Y(n2972) );
  MUX21X1_HVT U858 ( .A1(keyout[78]), .A2(n4159), .S0(n4506), .Y(n2971) );
  MUX21X1_HVT U859 ( .A1(keyout[77]), .A2(n4160), .S0(n4506), .Y(n2970) );
  MUX21X1_HVT U860 ( .A1(keyout[76]), .A2(n4161), .S0(n4506), .Y(n2969) );
  MUX21X1_HVT U861 ( .A1(keyout[75]), .A2(n4162), .S0(n4506), .Y(n2968) );
  MUX21X1_HVT U862 ( .A1(keyout[74]), .A2(n4163), .S0(n4506), .Y(n2967) );
  MUX21X1_HVT U863 ( .A1(keyout[73]), .A2(n4164), .S0(n4506), .Y(n2966) );
  MUX21X1_HVT U864 ( .A1(keyout[72]), .A2(n4165), .S0(n4506), .Y(n2965) );
  MUX21X1_HVT U865 ( .A1(keyout[71]), .A2(n4166), .S0(n4506), .Y(n2964) );
  MUX21X1_HVT U866 ( .A1(keyout[70]), .A2(n4167), .S0(n4506), .Y(n2963) );
  MUX21X1_HVT U867 ( .A1(keyout[69]), .A2(n4168), .S0(n4506), .Y(n2962) );
  MUX21X1_HVT U868 ( .A1(keyout[68]), .A2(n4169), .S0(n4506), .Y(n2961) );
  MUX21X1_HVT U869 ( .A1(keyout[67]), .A2(n4170), .S0(n4506), .Y(n2960) );
  MUX21X1_HVT U870 ( .A1(keyout[66]), .A2(n4171), .S0(n4506), .Y(n2959) );
  MUX21X1_HVT U871 ( .A1(keyout[65]), .A2(n4172), .S0(n4506), .Y(n2958) );
  MUX21X1_HVT U872 ( .A1(keyout[64]), .A2(n4173), .S0(n4506), .Y(n2957) );
  MUX21X1_HVT U873 ( .A1(keyout[63]), .A2(n4174), .S0(n4506), .Y(n2956) );
  MUX21X1_HVT U874 ( .A1(keyout[62]), .A2(n4175), .S0(n4506), .Y(n2955) );
  MUX21X1_HVT U875 ( .A1(keyout[61]), .A2(n4176), .S0(n4506), .Y(n2954) );
  MUX21X1_HVT U876 ( .A1(keyout[60]), .A2(n4177), .S0(n4506), .Y(n2953) );
  MUX21X1_HVT U877 ( .A1(keyout[59]), .A2(n4178), .S0(n4506), .Y(n2952) );
  MUX21X1_HVT U878 ( .A1(keyout[58]), .A2(n4179), .S0(n4506), .Y(n2951) );
  MUX21X1_HVT U879 ( .A1(keyout[57]), .A2(n4180), .S0(n4506), .Y(n2950) );
  MUX21X1_HVT U880 ( .A1(keyout[56]), .A2(n4181), .S0(n4506), .Y(n2949) );
  MUX21X1_HVT U881 ( .A1(keyout[55]), .A2(n4182), .S0(n4506), .Y(n2948) );
  MUX21X1_HVT U882 ( .A1(keyout[54]), .A2(n4183), .S0(n4506), .Y(n2947) );
  MUX21X1_HVT U883 ( .A1(keyout[53]), .A2(n4184), .S0(n4506), .Y(n2946) );
  MUX21X1_HVT U884 ( .A1(keyout[52]), .A2(n4185), .S0(n4506), .Y(n2945) );
  MUX21X1_HVT U885 ( .A1(keyout[51]), .A2(n4186), .S0(n4506), .Y(n2944) );
  MUX21X1_HVT U886 ( .A1(keyout[50]), .A2(n4187), .S0(n4506), .Y(n2943) );
  MUX21X1_HVT U887 ( .A1(keyout[49]), .A2(n4188), .S0(n4506), .Y(n2942) );
  MUX21X1_HVT U888 ( .A1(keyout[48]), .A2(n4189), .S0(n4506), .Y(n2941) );
  MUX21X1_HVT U889 ( .A1(keyout[47]), .A2(n4190), .S0(n4506), .Y(n2940) );
  MUX21X1_HVT U890 ( .A1(keyout[46]), .A2(n4191), .S0(n4506), .Y(n2939) );
  MUX21X1_HVT U891 ( .A1(keyout[45]), .A2(n4192), .S0(n4506), .Y(n2938) );
  MUX21X1_HVT U892 ( .A1(keyout[44]), .A2(n4193), .S0(n4506), .Y(n2937) );
  MUX21X1_HVT U893 ( .A1(keyout[43]), .A2(n4194), .S0(n4506), .Y(n2936) );
  MUX21X1_HVT U894 ( .A1(keyout[42]), .A2(n4195), .S0(n4506), .Y(n2935) );
  MUX21X1_HVT U895 ( .A1(keyout[41]), .A2(n4196), .S0(n4506), .Y(n2934) );
  MUX21X1_HVT U896 ( .A1(keyout[40]), .A2(n4197), .S0(n4506), .Y(n2933) );
  MUX21X1_HVT U897 ( .A1(keyout[39]), .A2(n4198), .S0(n4506), .Y(n2932) );
  MUX21X1_HVT U898 ( .A1(keyout[38]), .A2(n4199), .S0(n4506), .Y(n2931) );
  MUX21X1_HVT U899 ( .A1(keyout[37]), .A2(n4200), .S0(n4506), .Y(n2930) );
  MUX21X1_HVT U900 ( .A1(keyout[36]), .A2(n4201), .S0(n4506), .Y(n2929) );
  MUX21X1_HVT U901 ( .A1(keyout[35]), .A2(n4202), .S0(n4506), .Y(n2928) );
  MUX21X1_HVT U902 ( .A1(keyout[34]), .A2(n4203), .S0(n4506), .Y(n2927) );
  MUX21X1_HVT U903 ( .A1(keyout[33]), .A2(n4204), .S0(n4506), .Y(n2926) );
  MUX21X1_HVT U904 ( .A1(keyout[32]), .A2(n4205), .S0(n4506), .Y(n2925) );
  MUX21X1_HVT U905 ( .A1(keyout[31]), .A2(n4206), .S0(n4506), .Y(n2924) );
  MUX21X1_HVT U906 ( .A1(keyout[30]), .A2(n4207), .S0(n4506), .Y(n2923) );
  MUX21X1_HVT U907 ( .A1(keyout[29]), .A2(n4208), .S0(n4506), .Y(n2922) );
  MUX21X1_HVT U908 ( .A1(keyout[28]), .A2(n4209), .S0(n4506), .Y(n2921) );
  MUX21X1_HVT U909 ( .A1(keyout[27]), .A2(n4210), .S0(n4506), .Y(n2920) );
  MUX21X1_HVT U910 ( .A1(keyout[26]), .A2(n4211), .S0(n4506), .Y(n2919) );
  MUX21X1_HVT U911 ( .A1(keyout[25]), .A2(n4212), .S0(n4506), .Y(n2918) );
  MUX21X1_HVT U912 ( .A1(keyout[24]), .A2(n4213), .S0(n4506), .Y(n2917) );
  MUX21X1_HVT U913 ( .A1(keyout[23]), .A2(n4214), .S0(n4506), .Y(n2916) );
  MUX21X1_HVT U914 ( .A1(keyout[22]), .A2(n4215), .S0(n4506), .Y(n2915) );
  MUX21X1_HVT U915 ( .A1(keyout[21]), .A2(n4216), .S0(n4506), .Y(n2914) );
  MUX21X1_HVT U916 ( .A1(keyout[20]), .A2(n4217), .S0(n4506), .Y(n2913) );
  MUX21X1_HVT U917 ( .A1(keyout[19]), .A2(n4218), .S0(n4506), .Y(n2912) );
  MUX21X1_HVT U918 ( .A1(keyout[18]), .A2(n4219), .S0(n4506), .Y(n2911) );
  MUX21X1_HVT U919 ( .A1(keyout[17]), .A2(n4220), .S0(n4506), .Y(n2910) );
  MUX21X1_HVT U920 ( .A1(keyout[16]), .A2(n4221), .S0(n4506), .Y(n2909) );
  MUX21X1_HVT U921 ( .A1(keyout[15]), .A2(n4222), .S0(n4506), .Y(n2908) );
  MUX21X1_HVT U922 ( .A1(keyout[14]), .A2(n4223), .S0(n4506), .Y(n2907) );
  MUX21X1_HVT U923 ( .A1(keyout[13]), .A2(n4224), .S0(n4506), .Y(n2906) );
  MUX21X1_HVT U924 ( .A1(keyout[12]), .A2(n4225), .S0(n4506), .Y(n2905) );
  MUX21X1_HVT U925 ( .A1(keyout[11]), .A2(n4226), .S0(n4506), .Y(n2904) );
  MUX21X1_HVT U926 ( .A1(keyout[10]), .A2(n4227), .S0(n4506), .Y(n2903) );
  MUX21X1_HVT U927 ( .A1(keyout[9]), .A2(n4228), .S0(n4506), .Y(n2902) );
  MUX21X1_HVT U928 ( .A1(keyout[8]), .A2(n4229), .S0(n4506), .Y(n2901) );
  MUX21X1_HVT U929 ( .A1(keyout[7]), .A2(n4230), .S0(n4506), .Y(n2900) );
  MUX21X1_HVT U930 ( .A1(keyout[6]), .A2(n4231), .S0(n4506), .Y(n2899) );
  MUX21X1_HVT U931 ( .A1(keyout[5]), .A2(n4232), .S0(n4506), .Y(n2898) );
  MUX21X1_HVT U932 ( .A1(keyout[4]), .A2(n4233), .S0(n4506), .Y(n2897) );
  MUX21X1_HVT U933 ( .A1(keyout[3]), .A2(n4234), .S0(n4506), .Y(n2896) );
  MUX21X1_HVT U934 ( .A1(keyout[2]), .A2(n4235), .S0(n4506), .Y(n2895) );
  MUX21X1_HVT U935 ( .A1(keyout[1]), .A2(n4236), .S0(n4506), .Y(n2894) );
  MUX21X1_HVT U936 ( .A1(keyout[0]), .A2(n4237), .S0(n4506), .Y(n2893) );
  OR2X1_HVT U937 ( .A1(n4522), .A2(rest), .Y(n4506) );
  NAND3X0_HVT U938 ( .A1(state[2]), .A2(n1), .A3(n4535), .Y(n4522) );
  MUX21X1_HVT U939 ( .A1(keyout[127]), .A2(n1797), .S0(n4502), .Y(n2892) );
  MUX21X1_HVT U940 ( .A1(keyout[126]), .A2(n1798), .S0(n4502), .Y(n2891) );
  MUX21X1_HVT U941 ( .A1(keyout[125]), .A2(n1799), .S0(n4502), .Y(n2890) );
  MUX21X1_HVT U942 ( .A1(keyout[124]), .A2(n1800), .S0(n4502), .Y(n2889) );
  MUX21X1_HVT U943 ( .A1(keyout[123]), .A2(n1801), .S0(n4502), .Y(n2888) );
  MUX21X1_HVT U944 ( .A1(keyout[122]), .A2(n1802), .S0(n4502), .Y(n2887) );
  MUX21X1_HVT U945 ( .A1(keyout[121]), .A2(n1803), .S0(n4502), .Y(n2886) );
  MUX21X1_HVT U946 ( .A1(keyout[120]), .A2(n1804), .S0(n4502), .Y(n2885) );
  MUX21X1_HVT U947 ( .A1(keyout[119]), .A2(n1805), .S0(n4502), .Y(n2884) );
  MUX21X1_HVT U948 ( .A1(keyout[118]), .A2(n1806), .S0(n4502), .Y(n2883) );
  MUX21X1_HVT U949 ( .A1(keyout[117]), .A2(n1807), .S0(n4502), .Y(n2882) );
  MUX21X1_HVT U950 ( .A1(keyout[116]), .A2(n1808), .S0(n4502), .Y(n2881) );
  MUX21X1_HVT U951 ( .A1(keyout[115]), .A2(n1809), .S0(n4502), .Y(n2880) );
  MUX21X1_HVT U952 ( .A1(keyout[114]), .A2(n1810), .S0(n4502), .Y(n2879) );
  MUX21X1_HVT U953 ( .A1(keyout[113]), .A2(n1811), .S0(n4502), .Y(n2878) );
  MUX21X1_HVT U954 ( .A1(keyout[112]), .A2(n1812), .S0(n4502), .Y(n2877) );
  MUX21X1_HVT U955 ( .A1(keyout[111]), .A2(n1813), .S0(n4502), .Y(n2876) );
  MUX21X1_HVT U956 ( .A1(keyout[110]), .A2(n1814), .S0(n4502), .Y(n2875) );
  MUX21X1_HVT U957 ( .A1(keyout[109]), .A2(n1815), .S0(n4502), .Y(n2874) );
  MUX21X1_HVT U958 ( .A1(keyout[108]), .A2(n1816), .S0(n4502), .Y(n2873) );
  MUX21X1_HVT U959 ( .A1(keyout[107]), .A2(n1817), .S0(n4502), .Y(n2872) );
  MUX21X1_HVT U960 ( .A1(keyout[106]), .A2(n1818), .S0(n4502), .Y(n2871) );
  MUX21X1_HVT U961 ( .A1(keyout[105]), .A2(n1819), .S0(n4502), .Y(n2870) );
  MUX21X1_HVT U962 ( .A1(keyout[104]), .A2(n1820), .S0(n4502), .Y(n2869) );
  MUX21X1_HVT U963 ( .A1(keyout[103]), .A2(n1821), .S0(n4502), .Y(n2868) );
  MUX21X1_HVT U964 ( .A1(keyout[102]), .A2(n1822), .S0(n4502), .Y(n2867) );
  MUX21X1_HVT U965 ( .A1(keyout[101]), .A2(n1823), .S0(n4502), .Y(n2866) );
  MUX21X1_HVT U966 ( .A1(keyout[100]), .A2(n1824), .S0(n4502), .Y(n2865) );
  MUX21X1_HVT U967 ( .A1(keyout[99]), .A2(n1825), .S0(n4502), .Y(n2864) );
  MUX21X1_HVT U968 ( .A1(keyout[98]), .A2(n1826), .S0(n4502), .Y(n2863) );
  MUX21X1_HVT U969 ( .A1(keyout[97]), .A2(n1827), .S0(n4502), .Y(n2862) );
  MUX21X1_HVT U970 ( .A1(keyout[96]), .A2(n1828), .S0(n4502), .Y(n2861) );
  MUX21X1_HVT U971 ( .A1(keyout[95]), .A2(n1829), .S0(n4502), .Y(n2860) );
  MUX21X1_HVT U972 ( .A1(keyout[94]), .A2(n1830), .S0(n4502), .Y(n2859) );
  MUX21X1_HVT U973 ( .A1(keyout[93]), .A2(n1831), .S0(n4502), .Y(n2858) );
  MUX21X1_HVT U974 ( .A1(keyout[92]), .A2(n1832), .S0(n4502), .Y(n2857) );
  MUX21X1_HVT U975 ( .A1(keyout[91]), .A2(n1833), .S0(n4502), .Y(n2856) );
  MUX21X1_HVT U976 ( .A1(keyout[90]), .A2(n1834), .S0(n4502), .Y(n2855) );
  MUX21X1_HVT U977 ( .A1(keyout[89]), .A2(n1835), .S0(n4502), .Y(n2854) );
  MUX21X1_HVT U978 ( .A1(keyout[88]), .A2(n1836), .S0(n4502), .Y(n2853) );
  MUX21X1_HVT U979 ( .A1(keyout[87]), .A2(n1837), .S0(n4502), .Y(n2852) );
  MUX21X1_HVT U980 ( .A1(keyout[86]), .A2(n1838), .S0(n4502), .Y(n2851) );
  MUX21X1_HVT U981 ( .A1(keyout[85]), .A2(n1839), .S0(n4502), .Y(n2850) );
  MUX21X1_HVT U982 ( .A1(keyout[84]), .A2(n1840), .S0(n4502), .Y(n2849) );
  MUX21X1_HVT U983 ( .A1(keyout[83]), .A2(n1841), .S0(n4502), .Y(n2848) );
  MUX21X1_HVT U984 ( .A1(keyout[82]), .A2(n1842), .S0(n4502), .Y(n2847) );
  MUX21X1_HVT U985 ( .A1(keyout[81]), .A2(n1843), .S0(n4502), .Y(n2846) );
  MUX21X1_HVT U986 ( .A1(keyout[80]), .A2(n1844), .S0(n4502), .Y(n2845) );
  MUX21X1_HVT U987 ( .A1(keyout[79]), .A2(n1845), .S0(n4502), .Y(n2844) );
  MUX21X1_HVT U988 ( .A1(keyout[78]), .A2(n1846), .S0(n4502), .Y(n2843) );
  MUX21X1_HVT U989 ( .A1(keyout[77]), .A2(n1847), .S0(n4502), .Y(n2842) );
  MUX21X1_HVT U990 ( .A1(keyout[76]), .A2(n1848), .S0(n4502), .Y(n2841) );
  MUX21X1_HVT U991 ( .A1(keyout[75]), .A2(n1849), .S0(n4502), .Y(n2840) );
  MUX21X1_HVT U992 ( .A1(keyout[74]), .A2(n1850), .S0(n4502), .Y(n2839) );
  MUX21X1_HVT U993 ( .A1(keyout[73]), .A2(n1851), .S0(n4502), .Y(n2838) );
  MUX21X1_HVT U994 ( .A1(keyout[72]), .A2(n1852), .S0(n4502), .Y(n2837) );
  MUX21X1_HVT U995 ( .A1(keyout[71]), .A2(n1853), .S0(n4502), .Y(n2836) );
  MUX21X1_HVT U996 ( .A1(keyout[70]), .A2(n1854), .S0(n4502), .Y(n2835) );
  MUX21X1_HVT U997 ( .A1(keyout[69]), .A2(n1855), .S0(n4502), .Y(n2834) );
  MUX21X1_HVT U998 ( .A1(keyout[68]), .A2(n1856), .S0(n4502), .Y(n2833) );
  MUX21X1_HVT U999 ( .A1(keyout[67]), .A2(n1857), .S0(n4502), .Y(n2832) );
  MUX21X1_HVT U1000 ( .A1(keyout[66]), .A2(n1858), .S0(n4502), .Y(n2831) );
  MUX21X1_HVT U1001 ( .A1(keyout[65]), .A2(n1859), .S0(n4502), .Y(n2830) );
  MUX21X1_HVT U1002 ( .A1(keyout[64]), .A2(n1860), .S0(n4502), .Y(n2829) );
  MUX21X1_HVT U1003 ( .A1(keyout[63]), .A2(n1861), .S0(n4502), .Y(n2828) );
  MUX21X1_HVT U1004 ( .A1(keyout[62]), .A2(n1862), .S0(n4502), .Y(n2827) );
  MUX21X1_HVT U1005 ( .A1(keyout[61]), .A2(n1863), .S0(n4502), .Y(n2826) );
  MUX21X1_HVT U1006 ( .A1(keyout[60]), .A2(n1864), .S0(n4502), .Y(n2825) );
  MUX21X1_HVT U1007 ( .A1(keyout[59]), .A2(n1865), .S0(n4502), .Y(n2824) );
  MUX21X1_HVT U1008 ( .A1(keyout[58]), .A2(n1866), .S0(n4502), .Y(n2823) );
  MUX21X1_HVT U1009 ( .A1(keyout[57]), .A2(n1867), .S0(n4502), .Y(n2822) );
  MUX21X1_HVT U1010 ( .A1(keyout[56]), .A2(n1868), .S0(n4502), .Y(n2821) );
  MUX21X1_HVT U1011 ( .A1(keyout[55]), .A2(n1869), .S0(n4502), .Y(n2820) );
  MUX21X1_HVT U1012 ( .A1(keyout[54]), .A2(n1870), .S0(n4502), .Y(n2819) );
  MUX21X1_HVT U1013 ( .A1(keyout[53]), .A2(n1871), .S0(n4502), .Y(n2818) );
  MUX21X1_HVT U1014 ( .A1(keyout[52]), .A2(n1872), .S0(n4502), .Y(n2817) );
  MUX21X1_HVT U1015 ( .A1(keyout[51]), .A2(n1873), .S0(n4502), .Y(n2816) );
  MUX21X1_HVT U1016 ( .A1(keyout[50]), .A2(n1874), .S0(n4502), .Y(n2815) );
  MUX21X1_HVT U1017 ( .A1(keyout[49]), .A2(n1875), .S0(n4502), .Y(n2814) );
  MUX21X1_HVT U1018 ( .A1(keyout[48]), .A2(n1876), .S0(n4502), .Y(n2813) );
  MUX21X1_HVT U1019 ( .A1(keyout[47]), .A2(n1877), .S0(n4502), .Y(n2812) );
  MUX21X1_HVT U1020 ( .A1(keyout[46]), .A2(n1878), .S0(n4502), .Y(n2811) );
  MUX21X1_HVT U1021 ( .A1(keyout[45]), .A2(n1879), .S0(n4502), .Y(n2810) );
  MUX21X1_HVT U1022 ( .A1(keyout[44]), .A2(n1880), .S0(n4502), .Y(n2809) );
  MUX21X1_HVT U1023 ( .A1(keyout[43]), .A2(n1881), .S0(n4502), .Y(n2808) );
  MUX21X1_HVT U1024 ( .A1(keyout[42]), .A2(n1882), .S0(n4502), .Y(n2807) );
  MUX21X1_HVT U1025 ( .A1(keyout[41]), .A2(n1883), .S0(n4502), .Y(n2806) );
  MUX21X1_HVT U1026 ( .A1(keyout[40]), .A2(n1884), .S0(n4502), .Y(n2805) );
  MUX21X1_HVT U1027 ( .A1(keyout[39]), .A2(n1885), .S0(n4502), .Y(n2804) );
  MUX21X1_HVT U1028 ( .A1(keyout[38]), .A2(n1886), .S0(n4502), .Y(n2803) );
  MUX21X1_HVT U1029 ( .A1(keyout[37]), .A2(n1887), .S0(n4502), .Y(n2802) );
  MUX21X1_HVT U1030 ( .A1(keyout[36]), .A2(n1888), .S0(n4502), .Y(n2801) );
  MUX21X1_HVT U1031 ( .A1(keyout[35]), .A2(n1889), .S0(n4502), .Y(n2800) );
  MUX21X1_HVT U1032 ( .A1(keyout[34]), .A2(n1890), .S0(n4502), .Y(n2799) );
  MUX21X1_HVT U1033 ( .A1(keyout[33]), .A2(n1891), .S0(n4502), .Y(n2798) );
  MUX21X1_HVT U1034 ( .A1(keyout[32]), .A2(n1892), .S0(n4502), .Y(n2797) );
  MUX21X1_HVT U1035 ( .A1(keyout[31]), .A2(n1893), .S0(n4502), .Y(n2796) );
  MUX21X1_HVT U1036 ( .A1(keyout[30]), .A2(n1894), .S0(n4502), .Y(n2795) );
  MUX21X1_HVT U1037 ( .A1(keyout[29]), .A2(n1895), .S0(n4502), .Y(n2794) );
  MUX21X1_HVT U1038 ( .A1(keyout[28]), .A2(n1896), .S0(n4502), .Y(n2793) );
  MUX21X1_HVT U1039 ( .A1(keyout[27]), .A2(n1897), .S0(n4502), .Y(n2792) );
  MUX21X1_HVT U1040 ( .A1(keyout[26]), .A2(n1898), .S0(n4502), .Y(n2791) );
  MUX21X1_HVT U1041 ( .A1(keyout[25]), .A2(n1899), .S0(n4502), .Y(n2790) );
  MUX21X1_HVT U1042 ( .A1(keyout[24]), .A2(n1900), .S0(n4502), .Y(n2789) );
  MUX21X1_HVT U1043 ( .A1(keyout[23]), .A2(n1901), .S0(n4502), .Y(n2788) );
  MUX21X1_HVT U1044 ( .A1(keyout[22]), .A2(n1902), .S0(n4502), .Y(n2787) );
  MUX21X1_HVT U1045 ( .A1(keyout[21]), .A2(n1903), .S0(n4502), .Y(n2786) );
  MUX21X1_HVT U1046 ( .A1(keyout[20]), .A2(n1904), .S0(n4502), .Y(n2785) );
  MUX21X1_HVT U1047 ( .A1(keyout[19]), .A2(n1905), .S0(n4502), .Y(n2784) );
  MUX21X1_HVT U1048 ( .A1(keyout[18]), .A2(n1906), .S0(n4502), .Y(n2783) );
  MUX21X1_HVT U1049 ( .A1(keyout[17]), .A2(n1907), .S0(n4502), .Y(n2782) );
  MUX21X1_HVT U1050 ( .A1(keyout[16]), .A2(n1908), .S0(n4502), .Y(n2781) );
  MUX21X1_HVT U1051 ( .A1(keyout[15]), .A2(n1909), .S0(n4502), .Y(n2780) );
  MUX21X1_HVT U1052 ( .A1(keyout[14]), .A2(n1910), .S0(n4502), .Y(n2779) );
  MUX21X1_HVT U1053 ( .A1(keyout[13]), .A2(n1911), .S0(n4502), .Y(n2778) );
  MUX21X1_HVT U1054 ( .A1(keyout[12]), .A2(n1912), .S0(n4502), .Y(n2777) );
  MUX21X1_HVT U1055 ( .A1(keyout[11]), .A2(n1913), .S0(n4502), .Y(n2776) );
  MUX21X1_HVT U1056 ( .A1(keyout[10]), .A2(n1914), .S0(n4502), .Y(n2775) );
  MUX21X1_HVT U1057 ( .A1(keyout[9]), .A2(n1915), .S0(n4502), .Y(n2774) );
  MUX21X1_HVT U1058 ( .A1(keyout[8]), .A2(n1916), .S0(n4502), .Y(n2773) );
  MUX21X1_HVT U1059 ( .A1(keyout[7]), .A2(n1917), .S0(n4502), .Y(n2772) );
  MUX21X1_HVT U1060 ( .A1(keyout[6]), .A2(n1918), .S0(n4502), .Y(n2771) );
  MUX21X1_HVT U1061 ( .A1(keyout[5]), .A2(n1919), .S0(n4502), .Y(n2770) );
  MUX21X1_HVT U1062 ( .A1(keyout[4]), .A2(n1920), .S0(n4502), .Y(n2769) );
  MUX21X1_HVT U1063 ( .A1(keyout[3]), .A2(n1921), .S0(n4502), .Y(n2768) );
  MUX21X1_HVT U1064 ( .A1(keyout[2]), .A2(n1922), .S0(n4502), .Y(n2767) );
  MUX21X1_HVT U1065 ( .A1(keyout[1]), .A2(n1923), .S0(n4502), .Y(n2766) );
  MUX21X1_HVT U1066 ( .A1(keyout[0]), .A2(n1924), .S0(n4502), .Y(n2765) );
  OR2X1_HVT U1067 ( .A1(n4524), .A2(rest), .Y(n4502) );
  NAND3X0_HVT U1068 ( .A1(n4535), .A2(state[2]), .A3(state[0]), .Y(n4524) );
  INVX0_HVT U1069 ( .A(n4534), .Y(n4535) );
  NAND2X0_HVT U1070 ( .A1(state[1]), .A2(n4), .Y(n4534) );
  MUX21X1_HVT U1071 ( .A1(keyout[127]), .A2(n3854), .S0(n4497), .Y(n2764) );
  MUX21X1_HVT U1072 ( .A1(keyout[126]), .A2(n3855), .S0(n4497), .Y(n2763) );
  MUX21X1_HVT U1073 ( .A1(keyout[125]), .A2(n3856), .S0(n4497), .Y(n2762) );
  MUX21X1_HVT U1074 ( .A1(keyout[124]), .A2(n3857), .S0(n4497), .Y(n2761) );
  MUX21X1_HVT U1075 ( .A1(keyout[123]), .A2(n3858), .S0(n4497), .Y(n2760) );
  MUX21X1_HVT U1076 ( .A1(keyout[122]), .A2(n3859), .S0(n4497), .Y(n2759) );
  MUX21X1_HVT U1077 ( .A1(keyout[121]), .A2(n3860), .S0(n4497), .Y(n2758) );
  MUX21X1_HVT U1078 ( .A1(keyout[120]), .A2(n3861), .S0(n4497), .Y(n2757) );
  MUX21X1_HVT U1079 ( .A1(keyout[119]), .A2(n3862), .S0(n4497), .Y(n2756) );
  MUX21X1_HVT U1080 ( .A1(keyout[118]), .A2(n3863), .S0(n4497), .Y(n2755) );
  MUX21X1_HVT U1081 ( .A1(keyout[117]), .A2(n3864), .S0(n4497), .Y(n2754) );
  MUX21X1_HVT U1082 ( .A1(keyout[116]), .A2(n3865), .S0(n4497), .Y(n2753) );
  MUX21X1_HVT U1083 ( .A1(keyout[115]), .A2(n3866), .S0(n4497), .Y(n2752) );
  MUX21X1_HVT U1084 ( .A1(keyout[114]), .A2(n3867), .S0(n4497), .Y(n2751) );
  MUX21X1_HVT U1085 ( .A1(keyout[113]), .A2(n3868), .S0(n4497), .Y(n2750) );
  MUX21X1_HVT U1086 ( .A1(keyout[112]), .A2(n3869), .S0(n4497), .Y(n2749) );
  MUX21X1_HVT U1087 ( .A1(keyout[111]), .A2(n3870), .S0(n4497), .Y(n2748) );
  MUX21X1_HVT U1088 ( .A1(keyout[110]), .A2(n3871), .S0(n4497), .Y(n2747) );
  MUX21X1_HVT U1089 ( .A1(keyout[109]), .A2(n3872), .S0(n4497), .Y(n2746) );
  MUX21X1_HVT U1090 ( .A1(keyout[108]), .A2(n3873), .S0(n4497), .Y(n2745) );
  MUX21X1_HVT U1091 ( .A1(keyout[107]), .A2(n3874), .S0(n4497), .Y(n2744) );
  MUX21X1_HVT U1092 ( .A1(keyout[106]), .A2(n3875), .S0(n4497), .Y(n2743) );
  MUX21X1_HVT U1093 ( .A1(keyout[105]), .A2(n3876), .S0(n4497), .Y(n2742) );
  MUX21X1_HVT U1094 ( .A1(keyout[104]), .A2(n3877), .S0(n4497), .Y(n2741) );
  MUX21X1_HVT U1095 ( .A1(keyout[103]), .A2(n3878), .S0(n4497), .Y(n2740) );
  MUX21X1_HVT U1096 ( .A1(keyout[102]), .A2(n3879), .S0(n4497), .Y(n2739) );
  MUX21X1_HVT U1097 ( .A1(keyout[101]), .A2(n3880), .S0(n4497), .Y(n2738) );
  MUX21X1_HVT U1098 ( .A1(keyout[100]), .A2(n3881), .S0(n4497), .Y(n2737) );
  MUX21X1_HVT U1099 ( .A1(keyout[99]), .A2(n3882), .S0(n4497), .Y(n2736) );
  MUX21X1_HVT U1100 ( .A1(keyout[98]), .A2(n3883), .S0(n4497), .Y(n2735) );
  MUX21X1_HVT U1101 ( .A1(keyout[97]), .A2(n3884), .S0(n4497), .Y(n2734) );
  MUX21X1_HVT U1102 ( .A1(keyout[96]), .A2(n3885), .S0(n4497), .Y(n2733) );
  MUX21X1_HVT U1103 ( .A1(keyout[95]), .A2(n3886), .S0(n4497), .Y(n2732) );
  MUX21X1_HVT U1104 ( .A1(keyout[94]), .A2(n3887), .S0(n4497), .Y(n2731) );
  MUX21X1_HVT U1105 ( .A1(keyout[93]), .A2(n3888), .S0(n4497), .Y(n2730) );
  MUX21X1_HVT U1106 ( .A1(keyout[92]), .A2(n3889), .S0(n4497), .Y(n2729) );
  MUX21X1_HVT U1107 ( .A1(keyout[91]), .A2(n3890), .S0(n4497), .Y(n2728) );
  MUX21X1_HVT U1108 ( .A1(keyout[90]), .A2(n3891), .S0(n4497), .Y(n2727) );
  MUX21X1_HVT U1109 ( .A1(keyout[89]), .A2(n3892), .S0(n4497), .Y(n2726) );
  MUX21X1_HVT U1110 ( .A1(keyout[88]), .A2(n3893), .S0(n4497), .Y(n2725) );
  MUX21X1_HVT U1111 ( .A1(keyout[87]), .A2(n3894), .S0(n4497), .Y(n2724) );
  MUX21X1_HVT U1112 ( .A1(keyout[86]), .A2(n3895), .S0(n4497), .Y(n2723) );
  MUX21X1_HVT U1113 ( .A1(keyout[85]), .A2(n3896), .S0(n4497), .Y(n2722) );
  MUX21X1_HVT U1114 ( .A1(keyout[84]), .A2(n3897), .S0(n4497), .Y(n2721) );
  MUX21X1_HVT U1115 ( .A1(keyout[83]), .A2(n3898), .S0(n4497), .Y(n2720) );
  MUX21X1_HVT U1116 ( .A1(keyout[82]), .A2(n3899), .S0(n4497), .Y(n2719) );
  MUX21X1_HVT U1117 ( .A1(keyout[81]), .A2(n3900), .S0(n4497), .Y(n2718) );
  MUX21X1_HVT U1118 ( .A1(keyout[80]), .A2(n3901), .S0(n4497), .Y(n2717) );
  MUX21X1_HVT U1119 ( .A1(keyout[79]), .A2(n3902), .S0(n4497), .Y(n2716) );
  MUX21X1_HVT U1120 ( .A1(keyout[78]), .A2(n3903), .S0(n4497), .Y(n2715) );
  MUX21X1_HVT U1121 ( .A1(keyout[77]), .A2(n3904), .S0(n4497), .Y(n2714) );
  MUX21X1_HVT U1122 ( .A1(keyout[76]), .A2(n3905), .S0(n4497), .Y(n2713) );
  MUX21X1_HVT U1123 ( .A1(keyout[75]), .A2(n3906), .S0(n4497), .Y(n2712) );
  MUX21X1_HVT U1124 ( .A1(keyout[74]), .A2(n3907), .S0(n4497), .Y(n2711) );
  MUX21X1_HVT U1125 ( .A1(keyout[73]), .A2(n3908), .S0(n4497), .Y(n2710) );
  MUX21X1_HVT U1126 ( .A1(keyout[72]), .A2(n3909), .S0(n4497), .Y(n2709) );
  MUX21X1_HVT U1127 ( .A1(keyout[71]), .A2(n3910), .S0(n4497), .Y(n2708) );
  MUX21X1_HVT U1128 ( .A1(keyout[70]), .A2(n3911), .S0(n4497), .Y(n2707) );
  MUX21X1_HVT U1129 ( .A1(keyout[69]), .A2(n3912), .S0(n4497), .Y(n2706) );
  MUX21X1_HVT U1130 ( .A1(keyout[68]), .A2(n3913), .S0(n4497), .Y(n2705) );
  MUX21X1_HVT U1131 ( .A1(keyout[67]), .A2(n3914), .S0(n4497), .Y(n2704) );
  MUX21X1_HVT U1132 ( .A1(keyout[66]), .A2(n3915), .S0(n4497), .Y(n2703) );
  MUX21X1_HVT U1133 ( .A1(keyout[65]), .A2(n3916), .S0(n4497), .Y(n2702) );
  MUX21X1_HVT U1134 ( .A1(keyout[64]), .A2(n3917), .S0(n4497), .Y(n2701) );
  MUX21X1_HVT U1135 ( .A1(keyout[63]), .A2(n3918), .S0(n4497), .Y(n2700) );
  MUX21X1_HVT U1136 ( .A1(keyout[62]), .A2(n3919), .S0(n4497), .Y(n2699) );
  MUX21X1_HVT U1137 ( .A1(keyout[61]), .A2(n3920), .S0(n4497), .Y(n2698) );
  MUX21X1_HVT U1138 ( .A1(keyout[60]), .A2(n3921), .S0(n4497), .Y(n2697) );
  MUX21X1_HVT U1139 ( .A1(keyout[59]), .A2(n3922), .S0(n4497), .Y(n2696) );
  MUX21X1_HVT U1140 ( .A1(keyout[58]), .A2(n3923), .S0(n4497), .Y(n2695) );
  MUX21X1_HVT U1141 ( .A1(keyout[57]), .A2(n3924), .S0(n4497), .Y(n2694) );
  MUX21X1_HVT U1142 ( .A1(keyout[56]), .A2(n3925), .S0(n4497), .Y(n2693) );
  MUX21X1_HVT U1143 ( .A1(keyout[55]), .A2(n3926), .S0(n4497), .Y(n2692) );
  MUX21X1_HVT U1144 ( .A1(keyout[54]), .A2(n3927), .S0(n4497), .Y(n2691) );
  MUX21X1_HVT U1145 ( .A1(keyout[53]), .A2(n3928), .S0(n4497), .Y(n2690) );
  MUX21X1_HVT U1146 ( .A1(keyout[52]), .A2(n3929), .S0(n4497), .Y(n2689) );
  MUX21X1_HVT U1147 ( .A1(keyout[51]), .A2(n3930), .S0(n4497), .Y(n2688) );
  MUX21X1_HVT U1148 ( .A1(keyout[50]), .A2(n3931), .S0(n4497), .Y(n2687) );
  MUX21X1_HVT U1149 ( .A1(keyout[49]), .A2(n3932), .S0(n4497), .Y(n2686) );
  MUX21X1_HVT U1150 ( .A1(keyout[48]), .A2(n3933), .S0(n4497), .Y(n2685) );
  MUX21X1_HVT U1151 ( .A1(keyout[47]), .A2(n3934), .S0(n4497), .Y(n2684) );
  MUX21X1_HVT U1152 ( .A1(keyout[46]), .A2(n3935), .S0(n4497), .Y(n2683) );
  MUX21X1_HVT U1153 ( .A1(keyout[45]), .A2(n3936), .S0(n4497), .Y(n2682) );
  MUX21X1_HVT U1154 ( .A1(keyout[44]), .A2(n3937), .S0(n4497), .Y(n2681) );
  MUX21X1_HVT U1155 ( .A1(keyout[43]), .A2(n3938), .S0(n4497), .Y(n2680) );
  MUX21X1_HVT U1156 ( .A1(keyout[42]), .A2(n3939), .S0(n4497), .Y(n2679) );
  MUX21X1_HVT U1157 ( .A1(keyout[41]), .A2(n3940), .S0(n4497), .Y(n2678) );
  MUX21X1_HVT U1158 ( .A1(keyout[40]), .A2(n3941), .S0(n4497), .Y(n2677) );
  MUX21X1_HVT U1159 ( .A1(keyout[39]), .A2(n3942), .S0(n4497), .Y(n2676) );
  MUX21X1_HVT U1160 ( .A1(keyout[38]), .A2(n3943), .S0(n4497), .Y(n2675) );
  MUX21X1_HVT U1161 ( .A1(keyout[37]), .A2(n3944), .S0(n4497), .Y(n2674) );
  MUX21X1_HVT U1162 ( .A1(keyout[36]), .A2(n3945), .S0(n4497), .Y(n2673) );
  MUX21X1_HVT U1163 ( .A1(keyout[35]), .A2(n3946), .S0(n4497), .Y(n2672) );
  MUX21X1_HVT U1164 ( .A1(keyout[34]), .A2(n3947), .S0(n4497), .Y(n2671) );
  MUX21X1_HVT U1165 ( .A1(keyout[33]), .A2(n3948), .S0(n4497), .Y(n2670) );
  MUX21X1_HVT U1166 ( .A1(keyout[32]), .A2(n3949), .S0(n4497), .Y(n2669) );
  MUX21X1_HVT U1167 ( .A1(keyout[31]), .A2(n3950), .S0(n4497), .Y(n2668) );
  MUX21X1_HVT U1168 ( .A1(keyout[30]), .A2(n3951), .S0(n4497), .Y(n2667) );
  MUX21X1_HVT U1169 ( .A1(keyout[29]), .A2(n3952), .S0(n4497), .Y(n2666) );
  MUX21X1_HVT U1170 ( .A1(keyout[28]), .A2(n3953), .S0(n4497), .Y(n2665) );
  MUX21X1_HVT U1171 ( .A1(keyout[27]), .A2(n3954), .S0(n4497), .Y(n2664) );
  MUX21X1_HVT U1172 ( .A1(keyout[26]), .A2(n3955), .S0(n4497), .Y(n2663) );
  MUX21X1_HVT U1173 ( .A1(keyout[25]), .A2(n3956), .S0(n4497), .Y(n2662) );
  MUX21X1_HVT U1174 ( .A1(keyout[24]), .A2(n3957), .S0(n4497), .Y(n2661) );
  MUX21X1_HVT U1175 ( .A1(keyout[23]), .A2(n3958), .S0(n4497), .Y(n2660) );
  MUX21X1_HVT U1176 ( .A1(keyout[22]), .A2(n3959), .S0(n4497), .Y(n2659) );
  MUX21X1_HVT U1177 ( .A1(keyout[21]), .A2(n3960), .S0(n4497), .Y(n2658) );
  MUX21X1_HVT U1178 ( .A1(keyout[20]), .A2(n3961), .S0(n4497), .Y(n2657) );
  MUX21X1_HVT U1179 ( .A1(keyout[19]), .A2(n3962), .S0(n4497), .Y(n2656) );
  MUX21X1_HVT U1180 ( .A1(keyout[18]), .A2(n3963), .S0(n4497), .Y(n2655) );
  MUX21X1_HVT U1181 ( .A1(keyout[17]), .A2(n3964), .S0(n4497), .Y(n2654) );
  MUX21X1_HVT U1182 ( .A1(keyout[16]), .A2(n3965), .S0(n4497), .Y(n2653) );
  MUX21X1_HVT U1183 ( .A1(keyout[15]), .A2(n3966), .S0(n4497), .Y(n2652) );
  MUX21X1_HVT U1184 ( .A1(keyout[14]), .A2(n3967), .S0(n4497), .Y(n2651) );
  MUX21X1_HVT U1185 ( .A1(keyout[13]), .A2(n3968), .S0(n4497), .Y(n2650) );
  MUX21X1_HVT U1186 ( .A1(keyout[12]), .A2(n3969), .S0(n4497), .Y(n2649) );
  MUX21X1_HVT U1187 ( .A1(keyout[11]), .A2(n3970), .S0(n4497), .Y(n2648) );
  MUX21X1_HVT U1188 ( .A1(keyout[10]), .A2(n3971), .S0(n4497), .Y(n2647) );
  MUX21X1_HVT U1189 ( .A1(keyout[9]), .A2(n3972), .S0(n4497), .Y(n2646) );
  MUX21X1_HVT U1190 ( .A1(keyout[8]), .A2(n3973), .S0(n4497), .Y(n2645) );
  MUX21X1_HVT U1191 ( .A1(keyout[7]), .A2(n3974), .S0(n4497), .Y(n2644) );
  MUX21X1_HVT U1192 ( .A1(keyout[6]), .A2(n3975), .S0(n4497), .Y(n2643) );
  MUX21X1_HVT U1193 ( .A1(keyout[5]), .A2(n3976), .S0(n4497), .Y(n2642) );
  MUX21X1_HVT U1194 ( .A1(keyout[4]), .A2(n3977), .S0(n4497), .Y(n2641) );
  MUX21X1_HVT U1195 ( .A1(keyout[3]), .A2(n3978), .S0(n4497), .Y(n2640) );
  MUX21X1_HVT U1196 ( .A1(keyout[2]), .A2(n3979), .S0(n4497), .Y(n2639) );
  MUX21X1_HVT U1197 ( .A1(keyout[1]), .A2(n3980), .S0(n4497), .Y(n2638) );
  MUX21X1_HVT U1198 ( .A1(keyout[0]), .A2(n3981), .S0(n4497), .Y(n2637) );
  OR2X1_HVT U1199 ( .A1(n4533), .A2(rest), .Y(n4497) );
  NAND3X0_HVT U1200 ( .A1(n1), .A2(n3), .A3(n4537), .Y(n4533) );
  MUX21X1_HVT U1201 ( .A1(keyout[127]), .A2(n4238), .S0(n4500), .Y(n2636) );
  MUX21X1_HVT U1202 ( .A1(keyout[126]), .A2(n4239), .S0(n4500), .Y(n2635) );
  MUX21X1_HVT U1203 ( .A1(keyout[125]), .A2(n4240), .S0(n4500), .Y(n2634) );
  MUX21X1_HVT U1204 ( .A1(keyout[124]), .A2(n4241), .S0(n4500), .Y(n2633) );
  MUX21X1_HVT U1205 ( .A1(keyout[123]), .A2(n4242), .S0(n4500), .Y(n2632) );
  MUX21X1_HVT U1206 ( .A1(keyout[122]), .A2(n4243), .S0(n4500), .Y(n2631) );
  MUX21X1_HVT U1207 ( .A1(keyout[121]), .A2(n4244), .S0(n4500), .Y(n2630) );
  MUX21X1_HVT U1208 ( .A1(keyout[120]), .A2(n4245), .S0(n4500), .Y(n2629) );
  MUX21X1_HVT U1209 ( .A1(keyout[119]), .A2(n4246), .S0(n4500), .Y(n2628) );
  MUX21X1_HVT U1210 ( .A1(keyout[118]), .A2(n4247), .S0(n4500), .Y(n2627) );
  MUX21X1_HVT U1211 ( .A1(keyout[117]), .A2(n4248), .S0(n4500), .Y(n2626) );
  MUX21X1_HVT U1212 ( .A1(keyout[116]), .A2(n4249), .S0(n4500), .Y(n2625) );
  MUX21X1_HVT U1213 ( .A1(keyout[115]), .A2(n4250), .S0(n4500), .Y(n2624) );
  MUX21X1_HVT U1214 ( .A1(keyout[114]), .A2(n4251), .S0(n4500), .Y(n2623) );
  MUX21X1_HVT U1215 ( .A1(keyout[113]), .A2(n4252), .S0(n4500), .Y(n2622) );
  MUX21X1_HVT U1216 ( .A1(keyout[112]), .A2(n4253), .S0(n4500), .Y(n2621) );
  MUX21X1_HVT U1217 ( .A1(keyout[111]), .A2(n4254), .S0(n4500), .Y(n2620) );
  MUX21X1_HVT U1218 ( .A1(keyout[110]), .A2(n4255), .S0(n4500), .Y(n2619) );
  MUX21X1_HVT U1219 ( .A1(keyout[109]), .A2(n4256), .S0(n4500), .Y(n2618) );
  MUX21X1_HVT U1220 ( .A1(keyout[108]), .A2(n4257), .S0(n4500), .Y(n2617) );
  MUX21X1_HVT U1221 ( .A1(keyout[107]), .A2(n4258), .S0(n4500), .Y(n2616) );
  MUX21X1_HVT U1222 ( .A1(keyout[106]), .A2(n4259), .S0(n4500), .Y(n2615) );
  MUX21X1_HVT U1223 ( .A1(keyout[105]), .A2(n4260), .S0(n4500), .Y(n2614) );
  MUX21X1_HVT U1224 ( .A1(keyout[104]), .A2(n4261), .S0(n4500), .Y(n2613) );
  MUX21X1_HVT U1225 ( .A1(keyout[103]), .A2(n4262), .S0(n4500), .Y(n2612) );
  MUX21X1_HVT U1226 ( .A1(keyout[102]), .A2(n4263), .S0(n4500), .Y(n2611) );
  MUX21X1_HVT U1227 ( .A1(keyout[101]), .A2(n4264), .S0(n4500), .Y(n2610) );
  MUX21X1_HVT U1228 ( .A1(keyout[100]), .A2(n4265), .S0(n4500), .Y(n2609) );
  MUX21X1_HVT U1229 ( .A1(keyout[99]), .A2(n4266), .S0(n4500), .Y(n2608) );
  MUX21X1_HVT U1230 ( .A1(keyout[98]), .A2(n4267), .S0(n4500), .Y(n2607) );
  MUX21X1_HVT U1231 ( .A1(keyout[97]), .A2(n4268), .S0(n4500), .Y(n2606) );
  MUX21X1_HVT U1232 ( .A1(keyout[96]), .A2(n4269), .S0(n4500), .Y(n2605) );
  MUX21X1_HVT U1233 ( .A1(keyout[95]), .A2(n4270), .S0(n4500), .Y(n2604) );
  MUX21X1_HVT U1234 ( .A1(keyout[94]), .A2(n4271), .S0(n4500), .Y(n2603) );
  MUX21X1_HVT U1235 ( .A1(keyout[93]), .A2(n4272), .S0(n4500), .Y(n2602) );
  MUX21X1_HVT U1236 ( .A1(keyout[92]), .A2(n4273), .S0(n4500), .Y(n2601) );
  MUX21X1_HVT U1237 ( .A1(keyout[91]), .A2(n4274), .S0(n4500), .Y(n2600) );
  MUX21X1_HVT U1238 ( .A1(keyout[90]), .A2(n4275), .S0(n4500), .Y(n2599) );
  MUX21X1_HVT U1239 ( .A1(keyout[89]), .A2(n4276), .S0(n4500), .Y(n2598) );
  MUX21X1_HVT U1240 ( .A1(keyout[88]), .A2(n4277), .S0(n4500), .Y(n2597) );
  MUX21X1_HVT U1241 ( .A1(keyout[87]), .A2(n4278), .S0(n4500), .Y(n2596) );
  MUX21X1_HVT U1242 ( .A1(keyout[86]), .A2(n4279), .S0(n4500), .Y(n2595) );
  MUX21X1_HVT U1243 ( .A1(keyout[85]), .A2(n4280), .S0(n4500), .Y(n2594) );
  MUX21X1_HVT U1244 ( .A1(keyout[84]), .A2(n4281), .S0(n4500), .Y(n2593) );
  MUX21X1_HVT U1245 ( .A1(keyout[83]), .A2(n4282), .S0(n4500), .Y(n2592) );
  MUX21X1_HVT U1246 ( .A1(keyout[82]), .A2(n4283), .S0(n4500), .Y(n2591) );
  MUX21X1_HVT U1247 ( .A1(keyout[81]), .A2(n4284), .S0(n4500), .Y(n2590) );
  MUX21X1_HVT U1248 ( .A1(keyout[80]), .A2(n4285), .S0(n4500), .Y(n2589) );
  MUX21X1_HVT U1249 ( .A1(keyout[79]), .A2(n4286), .S0(n4500), .Y(n2588) );
  MUX21X1_HVT U1250 ( .A1(keyout[78]), .A2(n4287), .S0(n4500), .Y(n2587) );
  MUX21X1_HVT U1251 ( .A1(keyout[77]), .A2(n4288), .S0(n4500), .Y(n2586) );
  MUX21X1_HVT U1252 ( .A1(keyout[76]), .A2(n4289), .S0(n4500), .Y(n2585) );
  MUX21X1_HVT U1253 ( .A1(keyout[75]), .A2(n4290), .S0(n4500), .Y(n2584) );
  MUX21X1_HVT U1254 ( .A1(keyout[74]), .A2(n4291), .S0(n4500), .Y(n2583) );
  MUX21X1_HVT U1255 ( .A1(keyout[73]), .A2(n4292), .S0(n4500), .Y(n2582) );
  MUX21X1_HVT U1256 ( .A1(keyout[72]), .A2(n4293), .S0(n4500), .Y(n2581) );
  MUX21X1_HVT U1257 ( .A1(keyout[71]), .A2(n4294), .S0(n4500), .Y(n2580) );
  MUX21X1_HVT U1258 ( .A1(keyout[70]), .A2(n4295), .S0(n4500), .Y(n2579) );
  MUX21X1_HVT U1259 ( .A1(keyout[69]), .A2(n4296), .S0(n4500), .Y(n2578) );
  MUX21X1_HVT U1260 ( .A1(keyout[68]), .A2(n4297), .S0(n4500), .Y(n2577) );
  MUX21X1_HVT U1261 ( .A1(keyout[67]), .A2(n4298), .S0(n4500), .Y(n2576) );
  MUX21X1_HVT U1262 ( .A1(keyout[66]), .A2(n4299), .S0(n4500), .Y(n2575) );
  MUX21X1_HVT U1263 ( .A1(keyout[65]), .A2(n4300), .S0(n4500), .Y(n2574) );
  MUX21X1_HVT U1264 ( .A1(keyout[64]), .A2(n4301), .S0(n4500), .Y(n2573) );
  MUX21X1_HVT U1265 ( .A1(keyout[63]), .A2(n4302), .S0(n4500), .Y(n2572) );
  MUX21X1_HVT U1266 ( .A1(keyout[62]), .A2(n4303), .S0(n4500), .Y(n2571) );
  MUX21X1_HVT U1267 ( .A1(keyout[61]), .A2(n4304), .S0(n4500), .Y(n2570) );
  MUX21X1_HVT U1268 ( .A1(keyout[60]), .A2(n4305), .S0(n4500), .Y(n2569) );
  MUX21X1_HVT U1269 ( .A1(keyout[59]), .A2(n4306), .S0(n4500), .Y(n2568) );
  MUX21X1_HVT U1270 ( .A1(keyout[58]), .A2(n4307), .S0(n4500), .Y(n2567) );
  MUX21X1_HVT U1271 ( .A1(keyout[57]), .A2(n4308), .S0(n4500), .Y(n2566) );
  MUX21X1_HVT U1272 ( .A1(keyout[56]), .A2(n4309), .S0(n4500), .Y(n2565) );
  MUX21X1_HVT U1273 ( .A1(keyout[55]), .A2(n4310), .S0(n4500), .Y(n2564) );
  MUX21X1_HVT U1274 ( .A1(keyout[54]), .A2(n4311), .S0(n4500), .Y(n2563) );
  MUX21X1_HVT U1275 ( .A1(keyout[53]), .A2(n4312), .S0(n4500), .Y(n2562) );
  MUX21X1_HVT U1276 ( .A1(keyout[52]), .A2(n4313), .S0(n4500), .Y(n2561) );
  MUX21X1_HVT U1277 ( .A1(keyout[51]), .A2(n4314), .S0(n4500), .Y(n2560) );
  MUX21X1_HVT U1278 ( .A1(keyout[50]), .A2(n4315), .S0(n4500), .Y(n2559) );
  MUX21X1_HVT U1279 ( .A1(keyout[49]), .A2(n4316), .S0(n4500), .Y(n2558) );
  MUX21X1_HVT U1280 ( .A1(keyout[48]), .A2(n4317), .S0(n4500), .Y(n2557) );
  MUX21X1_HVT U1281 ( .A1(keyout[47]), .A2(n4318), .S0(n4500), .Y(n2556) );
  MUX21X1_HVT U1282 ( .A1(keyout[46]), .A2(n4319), .S0(n4500), .Y(n2555) );
  MUX21X1_HVT U1283 ( .A1(keyout[45]), .A2(n4320), .S0(n4500), .Y(n2554) );
  MUX21X1_HVT U1284 ( .A1(keyout[44]), .A2(n4321), .S0(n4500), .Y(n2553) );
  MUX21X1_HVT U1285 ( .A1(keyout[43]), .A2(n4322), .S0(n4500), .Y(n2552) );
  MUX21X1_HVT U1286 ( .A1(keyout[42]), .A2(n4323), .S0(n4500), .Y(n2551) );
  MUX21X1_HVT U1287 ( .A1(keyout[41]), .A2(n4324), .S0(n4500), .Y(n2550) );
  MUX21X1_HVT U1288 ( .A1(keyout[40]), .A2(n4325), .S0(n4500), .Y(n2549) );
  MUX21X1_HVT U1289 ( .A1(keyout[39]), .A2(n4326), .S0(n4500), .Y(n2548) );
  MUX21X1_HVT U1290 ( .A1(keyout[38]), .A2(n4327), .S0(n4500), .Y(n2547) );
  MUX21X1_HVT U1291 ( .A1(keyout[37]), .A2(n4328), .S0(n4500), .Y(n2546) );
  MUX21X1_HVT U1292 ( .A1(keyout[36]), .A2(n4329), .S0(n4500), .Y(n2545) );
  MUX21X1_HVT U1293 ( .A1(keyout[35]), .A2(n4330), .S0(n4500), .Y(n2544) );
  MUX21X1_HVT U1294 ( .A1(keyout[34]), .A2(n4331), .S0(n4500), .Y(n2543) );
  MUX21X1_HVT U1295 ( .A1(keyout[33]), .A2(n4332), .S0(n4500), .Y(n2542) );
  MUX21X1_HVT U1296 ( .A1(keyout[32]), .A2(n4333), .S0(n4500), .Y(n2541) );
  MUX21X1_HVT U1297 ( .A1(keyout[31]), .A2(n4334), .S0(n4500), .Y(n2540) );
  MUX21X1_HVT U1298 ( .A1(keyout[30]), .A2(n4335), .S0(n4500), .Y(n2539) );
  MUX21X1_HVT U1299 ( .A1(keyout[29]), .A2(n4336), .S0(n4500), .Y(n2538) );
  MUX21X1_HVT U1300 ( .A1(keyout[28]), .A2(n4337), .S0(n4500), .Y(n2537) );
  MUX21X1_HVT U1301 ( .A1(keyout[27]), .A2(n4338), .S0(n4500), .Y(n2536) );
  MUX21X1_HVT U1302 ( .A1(keyout[26]), .A2(n4339), .S0(n4500), .Y(n2535) );
  MUX21X1_HVT U1303 ( .A1(keyout[25]), .A2(n4340), .S0(n4500), .Y(n2534) );
  MUX21X1_HVT U1304 ( .A1(keyout[24]), .A2(n4341), .S0(n4500), .Y(n2533) );
  MUX21X1_HVT U1305 ( .A1(keyout[23]), .A2(n4342), .S0(n4500), .Y(n2532) );
  MUX21X1_HVT U1306 ( .A1(keyout[22]), .A2(n4343), .S0(n4500), .Y(n2531) );
  MUX21X1_HVT U1307 ( .A1(keyout[21]), .A2(n4344), .S0(n4500), .Y(n2530) );
  MUX21X1_HVT U1308 ( .A1(keyout[20]), .A2(n4345), .S0(n4500), .Y(n2529) );
  MUX21X1_HVT U1309 ( .A1(keyout[19]), .A2(n4346), .S0(n4500), .Y(n2528) );
  MUX21X1_HVT U1310 ( .A1(keyout[18]), .A2(n4347), .S0(n4500), .Y(n2527) );
  MUX21X1_HVT U1311 ( .A1(keyout[17]), .A2(n4348), .S0(n4500), .Y(n2526) );
  MUX21X1_HVT U1312 ( .A1(keyout[16]), .A2(n4349), .S0(n4500), .Y(n2525) );
  MUX21X1_HVT U1313 ( .A1(keyout[15]), .A2(n4350), .S0(n4500), .Y(n2524) );
  MUX21X1_HVT U1314 ( .A1(keyout[14]), .A2(n4351), .S0(n4500), .Y(n2523) );
  MUX21X1_HVT U1315 ( .A1(keyout[13]), .A2(n4352), .S0(n4500), .Y(n2522) );
  MUX21X1_HVT U1316 ( .A1(keyout[12]), .A2(n4353), .S0(n4500), .Y(n2521) );
  MUX21X1_HVT U1317 ( .A1(keyout[11]), .A2(n4354), .S0(n4500), .Y(n2520) );
  MUX21X1_HVT U1318 ( .A1(keyout[10]), .A2(n4355), .S0(n4500), .Y(n2519) );
  MUX21X1_HVT U1319 ( .A1(keyout[9]), .A2(n4356), .S0(n4500), .Y(n2518) );
  MUX21X1_HVT U1320 ( .A1(keyout[8]), .A2(n4357), .S0(n4500), .Y(n2517) );
  MUX21X1_HVT U1321 ( .A1(keyout[7]), .A2(n4358), .S0(n4500), .Y(n2516) );
  MUX21X1_HVT U1322 ( .A1(keyout[6]), .A2(n4359), .S0(n4500), .Y(n2515) );
  MUX21X1_HVT U1323 ( .A1(keyout[5]), .A2(n4360), .S0(n4500), .Y(n2514) );
  MUX21X1_HVT U1324 ( .A1(keyout[4]), .A2(n4361), .S0(n4500), .Y(n2513) );
  MUX21X1_HVT U1325 ( .A1(keyout[3]), .A2(n4362), .S0(n4500), .Y(n2512) );
  MUX21X1_HVT U1326 ( .A1(keyout[2]), .A2(n4363), .S0(n4500), .Y(n2511) );
  MUX21X1_HVT U1327 ( .A1(keyout[1]), .A2(n4364), .S0(n4500), .Y(n2510) );
  MUX21X1_HVT U1328 ( .A1(keyout[0]), .A2(n4365), .S0(n4500), .Y(n2509) );
  OR2X1_HVT U1329 ( .A1(n4517), .A2(rest), .Y(n4500) );
  NAND3X0_HVT U1330 ( .A1(n4537), .A2(n3), .A3(state[0]), .Y(n4517) );
  MUX21X1_HVT U1331 ( .A1(keyout[127]), .A2(n1925), .S0(n4499), .Y(n2508) );
  MUX21X1_HVT U1332 ( .A1(keyout[126]), .A2(n1926), .S0(n4499), .Y(n2507) );
  MUX21X1_HVT U1333 ( .A1(keyout[125]), .A2(n1927), .S0(n4499), .Y(n2506) );
  MUX21X1_HVT U1334 ( .A1(keyout[124]), .A2(n1928), .S0(n4499), .Y(n2505) );
  MUX21X1_HVT U1335 ( .A1(keyout[123]), .A2(n1929), .S0(n4499), .Y(n2504) );
  MUX21X1_HVT U1336 ( .A1(keyout[122]), .A2(n1930), .S0(n4499), .Y(n2503) );
  MUX21X1_HVT U1337 ( .A1(keyout[121]), .A2(n1931), .S0(n4499), .Y(n2502) );
  MUX21X1_HVT U1338 ( .A1(keyout[120]), .A2(n1932), .S0(n4499), .Y(n2501) );
  MUX21X1_HVT U1339 ( .A1(keyout[119]), .A2(n1933), .S0(n4499), .Y(n2500) );
  MUX21X1_HVT U1340 ( .A1(keyout[118]), .A2(n1934), .S0(n4499), .Y(n2499) );
  MUX21X1_HVT U1341 ( .A1(keyout[117]), .A2(n1935), .S0(n4499), .Y(n2498) );
  MUX21X1_HVT U1342 ( .A1(keyout[116]), .A2(n1936), .S0(n4499), .Y(n2497) );
  MUX21X1_HVT U1343 ( .A1(keyout[115]), .A2(n1937), .S0(n4499), .Y(n2496) );
  MUX21X1_HVT U1344 ( .A1(keyout[114]), .A2(n1938), .S0(n4499), .Y(n2495) );
  MUX21X1_HVT U1345 ( .A1(keyout[113]), .A2(n1939), .S0(n4499), .Y(n2494) );
  MUX21X1_HVT U1346 ( .A1(keyout[112]), .A2(n1940), .S0(n4499), .Y(n2493) );
  MUX21X1_HVT U1347 ( .A1(keyout[111]), .A2(n1941), .S0(n4499), .Y(n2492) );
  MUX21X1_HVT U1348 ( .A1(keyout[110]), .A2(n1942), .S0(n4499), .Y(n2491) );
  MUX21X1_HVT U1349 ( .A1(keyout[109]), .A2(n1943), .S0(n4499), .Y(n2490) );
  MUX21X1_HVT U1350 ( .A1(keyout[108]), .A2(n1944), .S0(n4499), .Y(n2489) );
  MUX21X1_HVT U1351 ( .A1(keyout[107]), .A2(n1945), .S0(n4499), .Y(n2488) );
  MUX21X1_HVT U1352 ( .A1(keyout[106]), .A2(n1946), .S0(n4499), .Y(n2487) );
  MUX21X1_HVT U1353 ( .A1(keyout[105]), .A2(n1947), .S0(n4499), .Y(n2486) );
  MUX21X1_HVT U1354 ( .A1(keyout[104]), .A2(n1948), .S0(n4499), .Y(n2485) );
  MUX21X1_HVT U1355 ( .A1(keyout[103]), .A2(n1949), .S0(n4499), .Y(n2484) );
  MUX21X1_HVT U1356 ( .A1(keyout[102]), .A2(n1950), .S0(n4499), .Y(n2483) );
  MUX21X1_HVT U1357 ( .A1(keyout[101]), .A2(n1951), .S0(n4499), .Y(n2482) );
  MUX21X1_HVT U1358 ( .A1(keyout[100]), .A2(n1952), .S0(n4499), .Y(n2481) );
  MUX21X1_HVT U1359 ( .A1(keyout[99]), .A2(n1953), .S0(n4499), .Y(n2480) );
  MUX21X1_HVT U1360 ( .A1(keyout[98]), .A2(n1954), .S0(n4499), .Y(n2479) );
  MUX21X1_HVT U1361 ( .A1(keyout[97]), .A2(n1955), .S0(n4499), .Y(n2478) );
  MUX21X1_HVT U1362 ( .A1(keyout[96]), .A2(n1956), .S0(n4499), .Y(n2477) );
  MUX21X1_HVT U1363 ( .A1(keyout[95]), .A2(n1957), .S0(n4499), .Y(n2476) );
  MUX21X1_HVT U1364 ( .A1(keyout[94]), .A2(n1958), .S0(n4499), .Y(n2475) );
  MUX21X1_HVT U1365 ( .A1(keyout[93]), .A2(n1959), .S0(n4499), .Y(n2474) );
  MUX21X1_HVT U1366 ( .A1(keyout[92]), .A2(n1960), .S0(n4499), .Y(n2473) );
  MUX21X1_HVT U1367 ( .A1(keyout[91]), .A2(n1961), .S0(n4499), .Y(n2472) );
  MUX21X1_HVT U1368 ( .A1(keyout[90]), .A2(n1962), .S0(n4499), .Y(n2471) );
  MUX21X1_HVT U1369 ( .A1(keyout[89]), .A2(n1963), .S0(n4499), .Y(n2470) );
  MUX21X1_HVT U1370 ( .A1(keyout[88]), .A2(n1964), .S0(n4499), .Y(n2469) );
  MUX21X1_HVT U1371 ( .A1(keyout[87]), .A2(n1965), .S0(n4499), .Y(n2468) );
  MUX21X1_HVT U1372 ( .A1(keyout[86]), .A2(n1966), .S0(n4499), .Y(n2467) );
  MUX21X1_HVT U1373 ( .A1(keyout[85]), .A2(n1967), .S0(n4499), .Y(n2466) );
  MUX21X1_HVT U1374 ( .A1(keyout[84]), .A2(n1968), .S0(n4499), .Y(n2465) );
  MUX21X1_HVT U1375 ( .A1(keyout[83]), .A2(n1969), .S0(n4499), .Y(n2464) );
  MUX21X1_HVT U1376 ( .A1(keyout[82]), .A2(n1970), .S0(n4499), .Y(n2463) );
  MUX21X1_HVT U1377 ( .A1(keyout[81]), .A2(n1971), .S0(n4499), .Y(n2462) );
  MUX21X1_HVT U1378 ( .A1(keyout[80]), .A2(n1972), .S0(n4499), .Y(n2461) );
  MUX21X1_HVT U1379 ( .A1(keyout[79]), .A2(n1973), .S0(n4499), .Y(n2460) );
  MUX21X1_HVT U1380 ( .A1(keyout[78]), .A2(n1974), .S0(n4499), .Y(n2459) );
  MUX21X1_HVT U1381 ( .A1(keyout[77]), .A2(n1975), .S0(n4499), .Y(n2458) );
  MUX21X1_HVT U1382 ( .A1(keyout[76]), .A2(n1976), .S0(n4499), .Y(n2457) );
  MUX21X1_HVT U1383 ( .A1(keyout[75]), .A2(n1977), .S0(n4499), .Y(n2456) );
  MUX21X1_HVT U1384 ( .A1(keyout[74]), .A2(n1978), .S0(n4499), .Y(n2455) );
  MUX21X1_HVT U1385 ( .A1(keyout[73]), .A2(n1979), .S0(n4499), .Y(n2454) );
  MUX21X1_HVT U1386 ( .A1(keyout[72]), .A2(n1980), .S0(n4499), .Y(n2453) );
  MUX21X1_HVT U1387 ( .A1(keyout[71]), .A2(n1981), .S0(n4499), .Y(n2452) );
  MUX21X1_HVT U1388 ( .A1(keyout[70]), .A2(n1982), .S0(n4499), .Y(n2451) );
  MUX21X1_HVT U1389 ( .A1(keyout[69]), .A2(n1983), .S0(n4499), .Y(n2450) );
  MUX21X1_HVT U1390 ( .A1(keyout[68]), .A2(n1984), .S0(n4499), .Y(n2449) );
  MUX21X1_HVT U1391 ( .A1(keyout[67]), .A2(n1985), .S0(n4499), .Y(n2448) );
  MUX21X1_HVT U1392 ( .A1(keyout[66]), .A2(n1986), .S0(n4499), .Y(n2447) );
  MUX21X1_HVT U1393 ( .A1(keyout[65]), .A2(n1987), .S0(n4499), .Y(n2446) );
  MUX21X1_HVT U1394 ( .A1(keyout[64]), .A2(n1988), .S0(n4499), .Y(n2445) );
  MUX21X1_HVT U1395 ( .A1(keyout[63]), .A2(n1989), .S0(n4499), .Y(n2444) );
  MUX21X1_HVT U1396 ( .A1(keyout[62]), .A2(n1990), .S0(n4499), .Y(n2443) );
  MUX21X1_HVT U1397 ( .A1(keyout[61]), .A2(n1991), .S0(n4499), .Y(n2442) );
  MUX21X1_HVT U1398 ( .A1(keyout[60]), .A2(n1992), .S0(n4499), .Y(n2441) );
  MUX21X1_HVT U1399 ( .A1(keyout[59]), .A2(n1993), .S0(n4499), .Y(n2440) );
  MUX21X1_HVT U1400 ( .A1(keyout[58]), .A2(n1994), .S0(n4499), .Y(n2439) );
  MUX21X1_HVT U1401 ( .A1(keyout[57]), .A2(n1995), .S0(n4499), .Y(n2438) );
  MUX21X1_HVT U1402 ( .A1(keyout[56]), .A2(n1996), .S0(n4499), .Y(n2437) );
  MUX21X1_HVT U1403 ( .A1(keyout[55]), .A2(n1997), .S0(n4499), .Y(n2436) );
  MUX21X1_HVT U1404 ( .A1(keyout[54]), .A2(n1998), .S0(n4499), .Y(n2435) );
  MUX21X1_HVT U1405 ( .A1(keyout[53]), .A2(n1999), .S0(n4499), .Y(n2434) );
  MUX21X1_HVT U1406 ( .A1(keyout[52]), .A2(n2000), .S0(n4499), .Y(n2433) );
  MUX21X1_HVT U1407 ( .A1(keyout[51]), .A2(n2001), .S0(n4499), .Y(n2432) );
  MUX21X1_HVT U1408 ( .A1(keyout[50]), .A2(n2002), .S0(n4499), .Y(n2431) );
  MUX21X1_HVT U1409 ( .A1(keyout[49]), .A2(n2003), .S0(n4499), .Y(n2430) );
  MUX21X1_HVT U1410 ( .A1(keyout[48]), .A2(n2004), .S0(n4499), .Y(n2429) );
  MUX21X1_HVT U1411 ( .A1(keyout[47]), .A2(n2005), .S0(n4499), .Y(n2428) );
  MUX21X1_HVT U1412 ( .A1(keyout[46]), .A2(n2006), .S0(n4499), .Y(n2427) );
  MUX21X1_HVT U1413 ( .A1(keyout[45]), .A2(n2007), .S0(n4499), .Y(n2426) );
  MUX21X1_HVT U1414 ( .A1(keyout[44]), .A2(n2008), .S0(n4499), .Y(n2425) );
  MUX21X1_HVT U1415 ( .A1(keyout[43]), .A2(n2009), .S0(n4499), .Y(n2424) );
  MUX21X1_HVT U1416 ( .A1(keyout[42]), .A2(n2010), .S0(n4499), .Y(n2423) );
  MUX21X1_HVT U1417 ( .A1(keyout[41]), .A2(n2011), .S0(n4499), .Y(n2422) );
  MUX21X1_HVT U1418 ( .A1(keyout[40]), .A2(n2012), .S0(n4499), .Y(n2421) );
  MUX21X1_HVT U1419 ( .A1(keyout[39]), .A2(n2013), .S0(n4499), .Y(n2420) );
  MUX21X1_HVT U1420 ( .A1(keyout[38]), .A2(n2014), .S0(n4499), .Y(n2419) );
  MUX21X1_HVT U1421 ( .A1(keyout[37]), .A2(n2015), .S0(n4499), .Y(n2418) );
  MUX21X1_HVT U1422 ( .A1(keyout[36]), .A2(n2016), .S0(n4499), .Y(n2417) );
  MUX21X1_HVT U1423 ( .A1(keyout[35]), .A2(n2017), .S0(n4499), .Y(n2416) );
  MUX21X1_HVT U1424 ( .A1(keyout[34]), .A2(n2018), .S0(n4499), .Y(n2415) );
  MUX21X1_HVT U1425 ( .A1(keyout[33]), .A2(n2019), .S0(n4499), .Y(n2414) );
  MUX21X1_HVT U1426 ( .A1(keyout[32]), .A2(n2020), .S0(n4499), .Y(n2413) );
  MUX21X1_HVT U1427 ( .A1(keyout[31]), .A2(n2021), .S0(n4499), .Y(n2412) );
  MUX21X1_HVT U1428 ( .A1(keyout[30]), .A2(n2022), .S0(n4499), .Y(n2411) );
  MUX21X1_HVT U1429 ( .A1(keyout[29]), .A2(n2023), .S0(n4499), .Y(n2410) );
  MUX21X1_HVT U1430 ( .A1(keyout[28]), .A2(n2024), .S0(n4499), .Y(n2409) );
  MUX21X1_HVT U1431 ( .A1(keyout[27]), .A2(n2025), .S0(n4499), .Y(n2408) );
  MUX21X1_HVT U1432 ( .A1(keyout[26]), .A2(n2026), .S0(n4499), .Y(n2407) );
  MUX21X1_HVT U1433 ( .A1(keyout[25]), .A2(n2027), .S0(n4499), .Y(n2406) );
  MUX21X1_HVT U1434 ( .A1(keyout[24]), .A2(n2028), .S0(n4499), .Y(n2405) );
  MUX21X1_HVT U1435 ( .A1(keyout[23]), .A2(n2029), .S0(n4499), .Y(n2404) );
  MUX21X1_HVT U1436 ( .A1(keyout[22]), .A2(n2030), .S0(n4499), .Y(n2403) );
  MUX21X1_HVT U1437 ( .A1(keyout[21]), .A2(n2031), .S0(n4499), .Y(n2402) );
  MUX21X1_HVT U1438 ( .A1(keyout[20]), .A2(n2032), .S0(n4499), .Y(n2401) );
  MUX21X1_HVT U1439 ( .A1(keyout[19]), .A2(n2033), .S0(n4499), .Y(n2400) );
  MUX21X1_HVT U1440 ( .A1(keyout[18]), .A2(n2034), .S0(n4499), .Y(n2399) );
  MUX21X1_HVT U1441 ( .A1(keyout[17]), .A2(n2035), .S0(n4499), .Y(n2398) );
  MUX21X1_HVT U1442 ( .A1(keyout[16]), .A2(n2036), .S0(n4499), .Y(n2397) );
  MUX21X1_HVT U1443 ( .A1(keyout[15]), .A2(n2037), .S0(n4499), .Y(n2396) );
  MUX21X1_HVT U1444 ( .A1(keyout[14]), .A2(n2038), .S0(n4499), .Y(n2395) );
  MUX21X1_HVT U1445 ( .A1(keyout[13]), .A2(n2039), .S0(n4499), .Y(n2394) );
  MUX21X1_HVT U1446 ( .A1(keyout[12]), .A2(n2040), .S0(n4499), .Y(n2393) );
  MUX21X1_HVT U1447 ( .A1(keyout[11]), .A2(n2041), .S0(n4499), .Y(n2392) );
  MUX21X1_HVT U1448 ( .A1(keyout[10]), .A2(n2042), .S0(n4499), .Y(n2391) );
  MUX21X1_HVT U1449 ( .A1(keyout[9]), .A2(n2043), .S0(n4499), .Y(n2390) );
  MUX21X1_HVT U1450 ( .A1(keyout[8]), .A2(n2044), .S0(n4499), .Y(n2389) );
  MUX21X1_HVT U1451 ( .A1(keyout[7]), .A2(n2045), .S0(n4499), .Y(n2388) );
  MUX21X1_HVT U1452 ( .A1(keyout[6]), .A2(n2046), .S0(n4499), .Y(n2387) );
  MUX21X1_HVT U1453 ( .A1(keyout[5]), .A2(n2047), .S0(n4499), .Y(n2386) );
  MUX21X1_HVT U1454 ( .A1(keyout[4]), .A2(n2048), .S0(n4499), .Y(n2385) );
  MUX21X1_HVT U1455 ( .A1(keyout[3]), .A2(n2049), .S0(n4499), .Y(n2384) );
  MUX21X1_HVT U1456 ( .A1(keyout[2]), .A2(n2050), .S0(n4499), .Y(n2383) );
  MUX21X1_HVT U1457 ( .A1(keyout[1]), .A2(n2051), .S0(n4499), .Y(n2382) );
  MUX21X1_HVT U1458 ( .A1(keyout[0]), .A2(n2052), .S0(n4499), .Y(n2381) );
  OR2X1_HVT U1459 ( .A1(n4528), .A2(rest), .Y(n4499) );
  NAND3X0_HVT U1460 ( .A1(n4537), .A2(n1), .A3(state[1]), .Y(n4528) );
  MUX21X1_HVT U1461 ( .A1(n1541), .A2(keyout[127]), .S0(n4512), .Y(n2380) );
  MUX21X1_HVT U1462 ( .A1(n1542), .A2(keyout[126]), .S0(n4512), .Y(n2379) );
  MUX21X1_HVT U1463 ( .A1(n1543), .A2(keyout[125]), .S0(n4512), .Y(n2378) );
  MUX21X1_HVT U1464 ( .A1(n1544), .A2(keyout[124]), .S0(n4512), .Y(n2377) );
  MUX21X1_HVT U1465 ( .A1(n1545), .A2(keyout[123]), .S0(n4512), .Y(n2376) );
  MUX21X1_HVT U1466 ( .A1(n1546), .A2(keyout[122]), .S0(n4512), .Y(n2375) );
  MUX21X1_HVT U1467 ( .A1(n1547), .A2(keyout[121]), .S0(n4512), .Y(n2374) );
  MUX21X1_HVT U1468 ( .A1(n1548), .A2(keyout[120]), .S0(n4512), .Y(n2373) );
  MUX21X1_HVT U1469 ( .A1(n1549), .A2(keyout[119]), .S0(n4512), .Y(n2372) );
  MUX21X1_HVT U1470 ( .A1(n1550), .A2(keyout[118]), .S0(n4512), .Y(n2371) );
  MUX21X1_HVT U1471 ( .A1(n1551), .A2(keyout[117]), .S0(n4512), .Y(n2370) );
  MUX21X1_HVT U1472 ( .A1(n1552), .A2(keyout[116]), .S0(n4512), .Y(n2369) );
  MUX21X1_HVT U1473 ( .A1(n1553), .A2(keyout[115]), .S0(n4512), .Y(n2368) );
  MUX21X1_HVT U1474 ( .A1(n1554), .A2(keyout[114]), .S0(n4512), .Y(n2367) );
  MUX21X1_HVT U1475 ( .A1(n1555), .A2(keyout[113]), .S0(n4512), .Y(n2366) );
  MUX21X1_HVT U1476 ( .A1(n1556), .A2(keyout[112]), .S0(n4512), .Y(n2365) );
  MUX21X1_HVT U1477 ( .A1(n1557), .A2(keyout[111]), .S0(n4512), .Y(n2364) );
  MUX21X1_HVT U1478 ( .A1(n1558), .A2(keyout[110]), .S0(n4512), .Y(n2363) );
  MUX21X1_HVT U1479 ( .A1(n1559), .A2(keyout[109]), .S0(n4512), .Y(n2362) );
  MUX21X1_HVT U1480 ( .A1(n1560), .A2(keyout[108]), .S0(n4512), .Y(n2361) );
  MUX21X1_HVT U1481 ( .A1(n1561), .A2(keyout[107]), .S0(n4512), .Y(n2360) );
  MUX21X1_HVT U1482 ( .A1(n1562), .A2(keyout[106]), .S0(n4512), .Y(n2359) );
  MUX21X1_HVT U1483 ( .A1(n1563), .A2(keyout[105]), .S0(n4512), .Y(n2358) );
  MUX21X1_HVT U1484 ( .A1(n1564), .A2(keyout[104]), .S0(n4512), .Y(n2357) );
  MUX21X1_HVT U1485 ( .A1(n1565), .A2(keyout[103]), .S0(n4512), .Y(n2356) );
  MUX21X1_HVT U1486 ( .A1(n1566), .A2(keyout[102]), .S0(n4512), .Y(n2355) );
  MUX21X1_HVT U1487 ( .A1(n1567), .A2(keyout[101]), .S0(n4512), .Y(n2354) );
  MUX21X1_HVT U1488 ( .A1(n1568), .A2(keyout[100]), .S0(n4512), .Y(n2353) );
  MUX21X1_HVT U1489 ( .A1(n1569), .A2(keyout[99]), .S0(n4512), .Y(n2352) );
  MUX21X1_HVT U1490 ( .A1(n1570), .A2(keyout[98]), .S0(n4512), .Y(n2351) );
  MUX21X1_HVT U1491 ( .A1(n1571), .A2(keyout[97]), .S0(n4512), .Y(n2350) );
  MUX21X1_HVT U1492 ( .A1(n1572), .A2(keyout[96]), .S0(n4512), .Y(n2349) );
  MUX21X1_HVT U1493 ( .A1(n1573), .A2(keyout[95]), .S0(n4512), .Y(n2348) );
  MUX21X1_HVT U1494 ( .A1(n1574), .A2(keyout[94]), .S0(n4512), .Y(n2347) );
  MUX21X1_HVT U1495 ( .A1(n1575), .A2(keyout[93]), .S0(n4512), .Y(n2346) );
  MUX21X1_HVT U1496 ( .A1(n1576), .A2(keyout[92]), .S0(n4512), .Y(n2345) );
  MUX21X1_HVT U1497 ( .A1(n1577), .A2(keyout[91]), .S0(n4512), .Y(n2344) );
  MUX21X1_HVT U1498 ( .A1(n1578), .A2(keyout[90]), .S0(n4512), .Y(n2343) );
  MUX21X1_HVT U1499 ( .A1(n1579), .A2(keyout[89]), .S0(n4512), .Y(n2342) );
  MUX21X1_HVT U1500 ( .A1(n1580), .A2(keyout[88]), .S0(n4512), .Y(n2341) );
  MUX21X1_HVT U1501 ( .A1(n1581), .A2(keyout[87]), .S0(n4512), .Y(n2340) );
  MUX21X1_HVT U1502 ( .A1(n1582), .A2(keyout[86]), .S0(n4512), .Y(n2339) );
  MUX21X1_HVT U1503 ( .A1(n1583), .A2(keyout[85]), .S0(n4512), .Y(n2338) );
  MUX21X1_HVT U1504 ( .A1(n1584), .A2(keyout[84]), .S0(n4512), .Y(n2337) );
  MUX21X1_HVT U1505 ( .A1(n1585), .A2(keyout[83]), .S0(n4512), .Y(n2336) );
  MUX21X1_HVT U1506 ( .A1(n1586), .A2(keyout[82]), .S0(n4512), .Y(n2335) );
  MUX21X1_HVT U1507 ( .A1(n1587), .A2(keyout[81]), .S0(n4512), .Y(n2334) );
  MUX21X1_HVT U1508 ( .A1(n1588), .A2(keyout[80]), .S0(n4512), .Y(n2333) );
  MUX21X1_HVT U1509 ( .A1(n1589), .A2(keyout[79]), .S0(n4512), .Y(n2332) );
  MUX21X1_HVT U1510 ( .A1(n1590), .A2(keyout[78]), .S0(n4512), .Y(n2331) );
  MUX21X1_HVT U1511 ( .A1(n1591), .A2(keyout[77]), .S0(n4512), .Y(n2330) );
  MUX21X1_HVT U1512 ( .A1(n1592), .A2(keyout[76]), .S0(n4512), .Y(n2329) );
  MUX21X1_HVT U1513 ( .A1(n1593), .A2(keyout[75]), .S0(n4512), .Y(n2328) );
  MUX21X1_HVT U1514 ( .A1(n1594), .A2(keyout[74]), .S0(n4512), .Y(n2327) );
  MUX21X1_HVT U1515 ( .A1(n1595), .A2(keyout[73]), .S0(n4512), .Y(n2326) );
  MUX21X1_HVT U1516 ( .A1(n1596), .A2(keyout[72]), .S0(n4512), .Y(n2325) );
  MUX21X1_HVT U1517 ( .A1(n1597), .A2(keyout[71]), .S0(n4512), .Y(n2324) );
  MUX21X1_HVT U1518 ( .A1(n1598), .A2(keyout[70]), .S0(n4512), .Y(n2323) );
  MUX21X1_HVT U1519 ( .A1(n1599), .A2(keyout[69]), .S0(n4512), .Y(n2322) );
  MUX21X1_HVT U1520 ( .A1(n1600), .A2(keyout[68]), .S0(n4512), .Y(n2321) );
  MUX21X1_HVT U1521 ( .A1(n1601), .A2(keyout[67]), .S0(n4512), .Y(n2320) );
  MUX21X1_HVT U1522 ( .A1(n1602), .A2(keyout[66]), .S0(n4512), .Y(n2319) );
  MUX21X1_HVT U1523 ( .A1(n1603), .A2(keyout[65]), .S0(n4512), .Y(n2318) );
  MUX21X1_HVT U1524 ( .A1(n1604), .A2(keyout[64]), .S0(n4512), .Y(n2317) );
  MUX21X1_HVT U1525 ( .A1(n1605), .A2(keyout[63]), .S0(n4512), .Y(n2316) );
  MUX21X1_HVT U1526 ( .A1(n1606), .A2(keyout[62]), .S0(n4512), .Y(n2315) );
  MUX21X1_HVT U1527 ( .A1(n1607), .A2(keyout[61]), .S0(n4512), .Y(n2314) );
  MUX21X1_HVT U1528 ( .A1(n1608), .A2(keyout[60]), .S0(n4512), .Y(n2313) );
  MUX21X1_HVT U1529 ( .A1(n1609), .A2(keyout[59]), .S0(n4512), .Y(n2312) );
  MUX21X1_HVT U1530 ( .A1(n1610), .A2(keyout[58]), .S0(n4512), .Y(n2311) );
  MUX21X1_HVT U1531 ( .A1(n1611), .A2(keyout[57]), .S0(n4512), .Y(n2310) );
  MUX21X1_HVT U1532 ( .A1(n1612), .A2(keyout[56]), .S0(n4512), .Y(n2309) );
  MUX21X1_HVT U1533 ( .A1(n1613), .A2(keyout[55]), .S0(n4512), .Y(n2308) );
  MUX21X1_HVT U1534 ( .A1(n1614), .A2(keyout[54]), .S0(n4512), .Y(n2307) );
  MUX21X1_HVT U1535 ( .A1(n1615), .A2(keyout[53]), .S0(n4512), .Y(n2306) );
  MUX21X1_HVT U1536 ( .A1(n1616), .A2(keyout[52]), .S0(n4512), .Y(n2305) );
  MUX21X1_HVT U1537 ( .A1(n1617), .A2(keyout[51]), .S0(n4512), .Y(n2304) );
  MUX21X1_HVT U1538 ( .A1(n1618), .A2(keyout[50]), .S0(n4512), .Y(n2303) );
  MUX21X1_HVT U1539 ( .A1(n1619), .A2(keyout[49]), .S0(n4512), .Y(n2302) );
  MUX21X1_HVT U1540 ( .A1(n1620), .A2(keyout[48]), .S0(n4512), .Y(n2301) );
  MUX21X1_HVT U1541 ( .A1(n1621), .A2(keyout[47]), .S0(n4512), .Y(n2300) );
  MUX21X1_HVT U1542 ( .A1(n1622), .A2(keyout[46]), .S0(n4512), .Y(n2299) );
  MUX21X1_HVT U1543 ( .A1(n1623), .A2(keyout[45]), .S0(n4512), .Y(n2298) );
  MUX21X1_HVT U1544 ( .A1(n1624), .A2(keyout[44]), .S0(n4512), .Y(n2297) );
  MUX21X1_HVT U1545 ( .A1(n1625), .A2(keyout[43]), .S0(n4512), .Y(n2296) );
  MUX21X1_HVT U1546 ( .A1(n1626), .A2(keyout[42]), .S0(n4512), .Y(n2295) );
  MUX21X1_HVT U1547 ( .A1(n1627), .A2(keyout[41]), .S0(n4512), .Y(n2294) );
  MUX21X1_HVT U1548 ( .A1(n1628), .A2(keyout[40]), .S0(n4512), .Y(n2293) );
  MUX21X1_HVT U1549 ( .A1(n1629), .A2(keyout[39]), .S0(n4512), .Y(n2292) );
  MUX21X1_HVT U1550 ( .A1(n1630), .A2(keyout[38]), .S0(n4512), .Y(n2291) );
  MUX21X1_HVT U1551 ( .A1(n1631), .A2(keyout[37]), .S0(n4512), .Y(n2290) );
  MUX21X1_HVT U1552 ( .A1(n1632), .A2(keyout[36]), .S0(n4512), .Y(n2289) );
  MUX21X1_HVT U1553 ( .A1(n1633), .A2(keyout[35]), .S0(n4512), .Y(n2288) );
  MUX21X1_HVT U1554 ( .A1(n1634), .A2(keyout[34]), .S0(n4512), .Y(n2287) );
  MUX21X1_HVT U1555 ( .A1(n1635), .A2(keyout[33]), .S0(n4512), .Y(n2286) );
  MUX21X1_HVT U1556 ( .A1(n1636), .A2(keyout[32]), .S0(n4512), .Y(n2285) );
  MUX21X1_HVT U1557 ( .A1(n1637), .A2(keyout[31]), .S0(n4512), .Y(n2284) );
  MUX21X1_HVT U1558 ( .A1(n1638), .A2(keyout[30]), .S0(n4512), .Y(n2283) );
  MUX21X1_HVT U1559 ( .A1(n1639), .A2(keyout[29]), .S0(n4512), .Y(n2282) );
  MUX21X1_HVT U1560 ( .A1(n1640), .A2(keyout[28]), .S0(n4512), .Y(n2281) );
  MUX21X1_HVT U1561 ( .A1(n1641), .A2(keyout[27]), .S0(n4512), .Y(n2280) );
  MUX21X1_HVT U1562 ( .A1(n1642), .A2(keyout[26]), .S0(n4512), .Y(n2279) );
  MUX21X1_HVT U1563 ( .A1(n1643), .A2(keyout[25]), .S0(n4512), .Y(n2278) );
  MUX21X1_HVT U1564 ( .A1(n1644), .A2(keyout[24]), .S0(n4512), .Y(n2277) );
  MUX21X1_HVT U1565 ( .A1(n1645), .A2(keyout[23]), .S0(n4512), .Y(n2276) );
  MUX21X1_HVT U1566 ( .A1(n1646), .A2(keyout[22]), .S0(n4512), .Y(n2275) );
  MUX21X1_HVT U1567 ( .A1(n1647), .A2(keyout[21]), .S0(n4512), .Y(n2274) );
  MUX21X1_HVT U1568 ( .A1(n1648), .A2(keyout[20]), .S0(n4512), .Y(n2273) );
  MUX21X1_HVT U1569 ( .A1(n1649), .A2(keyout[19]), .S0(n4512), .Y(n2272) );
  MUX21X1_HVT U1570 ( .A1(n1650), .A2(keyout[18]), .S0(n4512), .Y(n2271) );
  MUX21X1_HVT U1571 ( .A1(n1651), .A2(keyout[17]), .S0(n4512), .Y(n2270) );
  MUX21X1_HVT U1572 ( .A1(n1652), .A2(keyout[16]), .S0(n4512), .Y(n2269) );
  MUX21X1_HVT U1573 ( .A1(n1653), .A2(keyout[15]), .S0(n4512), .Y(n2268) );
  MUX21X1_HVT U1574 ( .A1(n1654), .A2(keyout[14]), .S0(n4512), .Y(n2267) );
  MUX21X1_HVT U1575 ( .A1(n1655), .A2(keyout[13]), .S0(n4512), .Y(n2266) );
  MUX21X1_HVT U1576 ( .A1(n1656), .A2(keyout[12]), .S0(n4512), .Y(n2265) );
  MUX21X1_HVT U1577 ( .A1(n1657), .A2(keyout[11]), .S0(n4512), .Y(n2264) );
  MUX21X1_HVT U1578 ( .A1(n1658), .A2(keyout[10]), .S0(n4512), .Y(n2263) );
  MUX21X1_HVT U1579 ( .A1(n1659), .A2(keyout[9]), .S0(n4512), .Y(n2262) );
  MUX21X1_HVT U1580 ( .A1(n1660), .A2(keyout[8]), .S0(n4512), .Y(n2261) );
  MUX21X1_HVT U1581 ( .A1(n1661), .A2(keyout[7]), .S0(n4512), .Y(n2260) );
  MUX21X1_HVT U1582 ( .A1(n1662), .A2(keyout[6]), .S0(n4512), .Y(n2259) );
  MUX21X1_HVT U1583 ( .A1(n1663), .A2(keyout[5]), .S0(n4512), .Y(n2258) );
  MUX21X1_HVT U1584 ( .A1(n1664), .A2(keyout[4]), .S0(n4512), .Y(n2257) );
  MUX21X1_HVT U1585 ( .A1(n1665), .A2(keyout[3]), .S0(n4512), .Y(n2256) );
  MUX21X1_HVT U1586 ( .A1(n1666), .A2(keyout[2]), .S0(n4512), .Y(n2255) );
  MUX21X1_HVT U1587 ( .A1(n1667), .A2(keyout[1]), .S0(n4512), .Y(n2254) );
  MUX21X1_HVT U1588 ( .A1(n1668), .A2(keyout[0]), .S0(n4512), .Y(n2253) );
  MUX21X1_HVT U1589 ( .A1(key_round[127]), .A2(n4538), .S0(n4512), .Y(n2252)
         );
  NAND4X0_HVT U1590 ( .A1(n4539), .A2(n4540), .A3(n4541), .A4(n4542), .Y(n4538) );
  OA222X1_HVT U1591 ( .A1(n1043), .A2(n4543), .A3(n1171), .A4(n4544), .A5(
        n1299), .A6(n4545), .Y(n4542) );
  OA222X1_HVT U1592 ( .A1(n659), .A2(n4546), .A3(n787), .A4(n4547), .A5(n915), 
        .A6(n4548), .Y(n4541) );
  OA222X1_HVT U1593 ( .A1(n275), .A2(n4549), .A3(n403), .A4(n4550), .A5(n531), 
        .A6(n4551), .Y(n4540) );
  OA22X1_HVT U1594 ( .A1(n19), .A2(n4552), .A3(n147), .A4(n4553), .Y(n4539) );
  MUX21X1_HVT U1595 ( .A1(key_round[126]), .A2(n4554), .S0(n4512), .Y(n2251)
         );
  NAND4X0_HVT U1596 ( .A1(n4555), .A2(n4556), .A3(n4557), .A4(n4558), .Y(n4554) );
  OA222X1_HVT U1597 ( .A1(n1044), .A2(n4543), .A3(n1172), .A4(n4544), .A5(
        n1300), .A6(n4545), .Y(n4558) );
  OA222X1_HVT U1598 ( .A1(n660), .A2(n4546), .A3(n788), .A4(n4547), .A5(n916), 
        .A6(n4548), .Y(n4557) );
  OA222X1_HVT U1599 ( .A1(n276), .A2(n4549), .A3(n404), .A4(n4550), .A5(n532), 
        .A6(n4551), .Y(n4556) );
  OA22X1_HVT U1600 ( .A1(n20), .A2(n4552), .A3(n148), .A4(n4553), .Y(n4555) );
  MUX21X1_HVT U1601 ( .A1(key_round[125]), .A2(n4559), .S0(n4512), .Y(n2250)
         );
  NAND4X0_HVT U1602 ( .A1(n4560), .A2(n4561), .A3(n4562), .A4(n4563), .Y(n4559) );
  OA222X1_HVT U1603 ( .A1(n1045), .A2(n4543), .A3(n1173), .A4(n4544), .A5(
        n1301), .A6(n4545), .Y(n4563) );
  OA222X1_HVT U1604 ( .A1(n661), .A2(n4546), .A3(n789), .A4(n4547), .A5(n917), 
        .A6(n4548), .Y(n4562) );
  OA222X1_HVT U1605 ( .A1(n277), .A2(n4549), .A3(n405), .A4(n4550), .A5(n533), 
        .A6(n4551), .Y(n4561) );
  OA22X1_HVT U1606 ( .A1(n21), .A2(n4552), .A3(n149), .A4(n4553), .Y(n4560) );
  MUX21X1_HVT U1607 ( .A1(key_round[124]), .A2(n4564), .S0(n4512), .Y(n2249)
         );
  NAND4X0_HVT U1608 ( .A1(n4565), .A2(n4566), .A3(n4567), .A4(n4568), .Y(n4564) );
  OA222X1_HVT U1609 ( .A1(n1046), .A2(n4543), .A3(n1174), .A4(n4544), .A5(
        n1302), .A6(n4545), .Y(n4568) );
  OA222X1_HVT U1610 ( .A1(n662), .A2(n4546), .A3(n790), .A4(n4547), .A5(n918), 
        .A6(n4548), .Y(n4567) );
  OA222X1_HVT U1611 ( .A1(n278), .A2(n4549), .A3(n406), .A4(n4550), .A5(n534), 
        .A6(n4551), .Y(n4566) );
  OA22X1_HVT U1612 ( .A1(n22), .A2(n4552), .A3(n150), .A4(n4553), .Y(n4565) );
  MUX21X1_HVT U1613 ( .A1(key_round[123]), .A2(n4569), .S0(n4512), .Y(n2248)
         );
  NAND4X0_HVT U1614 ( .A1(n4570), .A2(n4571), .A3(n4572), .A4(n4573), .Y(n4569) );
  OA222X1_HVT U1615 ( .A1(n1047), .A2(n4543), .A3(n1175), .A4(n4544), .A5(
        n1303), .A6(n4545), .Y(n4573) );
  OA222X1_HVT U1616 ( .A1(n663), .A2(n4546), .A3(n791), .A4(n4547), .A5(n919), 
        .A6(n4548), .Y(n4572) );
  OA222X1_HVT U1617 ( .A1(n279), .A2(n4549), .A3(n407), .A4(n4550), .A5(n535), 
        .A6(n4551), .Y(n4571) );
  OA22X1_HVT U1618 ( .A1(n23), .A2(n4552), .A3(n151), .A4(n4553), .Y(n4570) );
  MUX21X1_HVT U1619 ( .A1(key_round[122]), .A2(n4574), .S0(n4512), .Y(n2247)
         );
  NAND4X0_HVT U1620 ( .A1(n4575), .A2(n4576), .A3(n4577), .A4(n4578), .Y(n4574) );
  OA222X1_HVT U1621 ( .A1(n1048), .A2(n4543), .A3(n1176), .A4(n4544), .A5(
        n1304), .A6(n4545), .Y(n4578) );
  OA222X1_HVT U1622 ( .A1(n664), .A2(n4546), .A3(n792), .A4(n4547), .A5(n920), 
        .A6(n4548), .Y(n4577) );
  OA222X1_HVT U1623 ( .A1(n280), .A2(n4549), .A3(n408), .A4(n4550), .A5(n536), 
        .A6(n4551), .Y(n4576) );
  OA22X1_HVT U1624 ( .A1(n24), .A2(n4552), .A3(n152), .A4(n4553), .Y(n4575) );
  MUX21X1_HVT U1625 ( .A1(key_round[121]), .A2(n4579), .S0(n4512), .Y(n2246)
         );
  NAND4X0_HVT U1626 ( .A1(n4580), .A2(n4581), .A3(n4582), .A4(n4583), .Y(n4579) );
  OA222X1_HVT U1627 ( .A1(n1049), .A2(n4543), .A3(n1177), .A4(n4544), .A5(
        n1305), .A6(n4545), .Y(n4583) );
  OA222X1_HVT U1628 ( .A1(n665), .A2(n4546), .A3(n793), .A4(n4547), .A5(n921), 
        .A6(n4548), .Y(n4582) );
  OA222X1_HVT U1629 ( .A1(n281), .A2(n4549), .A3(n409), .A4(n4550), .A5(n537), 
        .A6(n4551), .Y(n4581) );
  OA22X1_HVT U1630 ( .A1(n25), .A2(n4552), .A3(n153), .A4(n4553), .Y(n4580) );
  MUX21X1_HVT U1631 ( .A1(key_round[120]), .A2(n4584), .S0(n4512), .Y(n2245)
         );
  NAND4X0_HVT U1632 ( .A1(n4585), .A2(n4586), .A3(n4587), .A4(n4588), .Y(n4584) );
  OA222X1_HVT U1633 ( .A1(n1050), .A2(n4543), .A3(n1178), .A4(n4544), .A5(
        n1306), .A6(n4545), .Y(n4588) );
  OA222X1_HVT U1634 ( .A1(n666), .A2(n4546), .A3(n794), .A4(n4547), .A5(n922), 
        .A6(n4548), .Y(n4587) );
  OA222X1_HVT U1635 ( .A1(n282), .A2(n4549), .A3(n410), .A4(n4550), .A5(n538), 
        .A6(n4551), .Y(n4586) );
  OA22X1_HVT U1636 ( .A1(n26), .A2(n4552), .A3(n154), .A4(n4553), .Y(n4585) );
  MUX21X1_HVT U1637 ( .A1(key_round[119]), .A2(n4589), .S0(n4512), .Y(n2244)
         );
  NAND4X0_HVT U1638 ( .A1(n4590), .A2(n4591), .A3(n4592), .A4(n4593), .Y(n4589) );
  OA222X1_HVT U1639 ( .A1(n1051), .A2(n4543), .A3(n1179), .A4(n4544), .A5(
        n1307), .A6(n4545), .Y(n4593) );
  OA222X1_HVT U1640 ( .A1(n667), .A2(n4546), .A3(n795), .A4(n4547), .A5(n923), 
        .A6(n4548), .Y(n4592) );
  OA222X1_HVT U1641 ( .A1(n283), .A2(n4549), .A3(n411), .A4(n4550), .A5(n539), 
        .A6(n4551), .Y(n4591) );
  OA22X1_HVT U1642 ( .A1(n27), .A2(n4552), .A3(n155), .A4(n4553), .Y(n4590) );
  MUX21X1_HVT U1643 ( .A1(key_round[118]), .A2(n4594), .S0(n4512), .Y(n2243)
         );
  NAND4X0_HVT U1644 ( .A1(n4595), .A2(n4596), .A3(n4597), .A4(n4598), .Y(n4594) );
  OA222X1_HVT U1645 ( .A1(n1052), .A2(n4543), .A3(n1180), .A4(n4544), .A5(
        n1308), .A6(n4545), .Y(n4598) );
  OA222X1_HVT U1646 ( .A1(n668), .A2(n4546), .A3(n796), .A4(n4547), .A5(n924), 
        .A6(n4548), .Y(n4597) );
  OA222X1_HVT U1647 ( .A1(n284), .A2(n4549), .A3(n412), .A4(n4550), .A5(n540), 
        .A6(n4551), .Y(n4596) );
  OA22X1_HVT U1648 ( .A1(n28), .A2(n4552), .A3(n156), .A4(n4553), .Y(n4595) );
  MUX21X1_HVT U1649 ( .A1(key_round[117]), .A2(n4599), .S0(n4512), .Y(n2242)
         );
  NAND4X0_HVT U1650 ( .A1(n4600), .A2(n4601), .A3(n4602), .A4(n4603), .Y(n4599) );
  OA222X1_HVT U1651 ( .A1(n1053), .A2(n4543), .A3(n1181), .A4(n4544), .A5(
        n1309), .A6(n4545), .Y(n4603) );
  OA222X1_HVT U1652 ( .A1(n669), .A2(n4546), .A3(n797), .A4(n4547), .A5(n925), 
        .A6(n4548), .Y(n4602) );
  OA222X1_HVT U1653 ( .A1(n285), .A2(n4549), .A3(n413), .A4(n4550), .A5(n541), 
        .A6(n4551), .Y(n4601) );
  OA22X1_HVT U1654 ( .A1(n29), .A2(n4552), .A3(n157), .A4(n4553), .Y(n4600) );
  MUX21X1_HVT U1655 ( .A1(key_round[116]), .A2(n4604), .S0(n4512), .Y(n2241)
         );
  NAND4X0_HVT U1656 ( .A1(n4605), .A2(n4606), .A3(n4607), .A4(n4608), .Y(n4604) );
  OA222X1_HVT U1657 ( .A1(n1054), .A2(n4543), .A3(n1182), .A4(n4544), .A5(
        n1310), .A6(n4545), .Y(n4608) );
  OA222X1_HVT U1658 ( .A1(n670), .A2(n4546), .A3(n798), .A4(n4547), .A5(n926), 
        .A6(n4548), .Y(n4607) );
  OA222X1_HVT U1659 ( .A1(n286), .A2(n4549), .A3(n414), .A4(n4550), .A5(n542), 
        .A6(n4551), .Y(n4606) );
  OA22X1_HVT U1660 ( .A1(n30), .A2(n4552), .A3(n158), .A4(n4553), .Y(n4605) );
  MUX21X1_HVT U1661 ( .A1(key_round[115]), .A2(n4609), .S0(n4512), .Y(n2240)
         );
  NAND4X0_HVT U1662 ( .A1(n4610), .A2(n4611), .A3(n4612), .A4(n4613), .Y(n4609) );
  OA222X1_HVT U1663 ( .A1(n1055), .A2(n4543), .A3(n1183), .A4(n4544), .A5(
        n1311), .A6(n4545), .Y(n4613) );
  OA222X1_HVT U1664 ( .A1(n671), .A2(n4546), .A3(n799), .A4(n4547), .A5(n927), 
        .A6(n4548), .Y(n4612) );
  OA222X1_HVT U1665 ( .A1(n287), .A2(n4549), .A3(n415), .A4(n4550), .A5(n543), 
        .A6(n4551), .Y(n4611) );
  OA22X1_HVT U1666 ( .A1(n31), .A2(n4552), .A3(n159), .A4(n4553), .Y(n4610) );
  MUX21X1_HVT U1667 ( .A1(key_round[114]), .A2(n4614), .S0(n4512), .Y(n2239)
         );
  NAND4X0_HVT U1668 ( .A1(n4615), .A2(n4616), .A3(n4617), .A4(n4618), .Y(n4614) );
  OA222X1_HVT U1669 ( .A1(n1056), .A2(n4543), .A3(n1184), .A4(n4544), .A5(
        n1312), .A6(n4545), .Y(n4618) );
  OA222X1_HVT U1670 ( .A1(n672), .A2(n4546), .A3(n800), .A4(n4547), .A5(n928), 
        .A6(n4548), .Y(n4617) );
  OA222X1_HVT U1671 ( .A1(n288), .A2(n4549), .A3(n416), .A4(n4550), .A5(n544), 
        .A6(n4551), .Y(n4616) );
  OA22X1_HVT U1672 ( .A1(n32), .A2(n4552), .A3(n160), .A4(n4553), .Y(n4615) );
  MUX21X1_HVT U1673 ( .A1(key_round[113]), .A2(n4619), .S0(n4512), .Y(n2238)
         );
  NAND4X0_HVT U1674 ( .A1(n4620), .A2(n4621), .A3(n4622), .A4(n4623), .Y(n4619) );
  OA222X1_HVT U1675 ( .A1(n1057), .A2(n4543), .A3(n1185), .A4(n4544), .A5(
        n1313), .A6(n4545), .Y(n4623) );
  OA222X1_HVT U1676 ( .A1(n673), .A2(n4546), .A3(n801), .A4(n4547), .A5(n929), 
        .A6(n4548), .Y(n4622) );
  OA222X1_HVT U1677 ( .A1(n289), .A2(n4549), .A3(n417), .A4(n4550), .A5(n545), 
        .A6(n4551), .Y(n4621) );
  OA22X1_HVT U1678 ( .A1(n33), .A2(n4552), .A3(n161), .A4(n4553), .Y(n4620) );
  MUX21X1_HVT U1679 ( .A1(key_round[112]), .A2(n4624), .S0(n4512), .Y(n2237)
         );
  NAND4X0_HVT U1680 ( .A1(n4625), .A2(n4626), .A3(n4627), .A4(n4628), .Y(n4624) );
  OA222X1_HVT U1681 ( .A1(n1058), .A2(n4543), .A3(n1186), .A4(n4544), .A5(
        n1314), .A6(n4545), .Y(n4628) );
  OA222X1_HVT U1682 ( .A1(n674), .A2(n4546), .A3(n802), .A4(n4547), .A5(n930), 
        .A6(n4548), .Y(n4627) );
  OA222X1_HVT U1683 ( .A1(n290), .A2(n4549), .A3(n418), .A4(n4550), .A5(n546), 
        .A6(n4551), .Y(n4626) );
  OA22X1_HVT U1684 ( .A1(n34), .A2(n4552), .A3(n162), .A4(n4553), .Y(n4625) );
  MUX21X1_HVT U1685 ( .A1(key_round[111]), .A2(n4629), .S0(n4512), .Y(n2236)
         );
  NAND4X0_HVT U1686 ( .A1(n4630), .A2(n4631), .A3(n4632), .A4(n4633), .Y(n4629) );
  OA222X1_HVT U1687 ( .A1(n1059), .A2(n4543), .A3(n1187), .A4(n4544), .A5(
        n1315), .A6(n4545), .Y(n4633) );
  OA222X1_HVT U1688 ( .A1(n675), .A2(n4546), .A3(n803), .A4(n4547), .A5(n931), 
        .A6(n4548), .Y(n4632) );
  OA222X1_HVT U1689 ( .A1(n291), .A2(n4549), .A3(n419), .A4(n4550), .A5(n547), 
        .A6(n4551), .Y(n4631) );
  OA22X1_HVT U1690 ( .A1(n35), .A2(n4552), .A3(n163), .A4(n4553), .Y(n4630) );
  MUX21X1_HVT U1691 ( .A1(key_round[110]), .A2(n4634), .S0(n4512), .Y(n2235)
         );
  NAND4X0_HVT U1692 ( .A1(n4635), .A2(n4636), .A3(n4637), .A4(n4638), .Y(n4634) );
  OA222X1_HVT U1693 ( .A1(n1060), .A2(n4543), .A3(n1188), .A4(n4544), .A5(
        n1316), .A6(n4545), .Y(n4638) );
  OA222X1_HVT U1694 ( .A1(n676), .A2(n4546), .A3(n804), .A4(n4547), .A5(n932), 
        .A6(n4548), .Y(n4637) );
  OA222X1_HVT U1695 ( .A1(n292), .A2(n4549), .A3(n420), .A4(n4550), .A5(n548), 
        .A6(n4551), .Y(n4636) );
  OA22X1_HVT U1696 ( .A1(n36), .A2(n4552), .A3(n164), .A4(n4553), .Y(n4635) );
  MUX21X1_HVT U1697 ( .A1(key_round[109]), .A2(n4639), .S0(n4512), .Y(n2234)
         );
  NAND4X0_HVT U1698 ( .A1(n4640), .A2(n4641), .A3(n4642), .A4(n4643), .Y(n4639) );
  OA222X1_HVT U1699 ( .A1(n1061), .A2(n4543), .A3(n1189), .A4(n4544), .A5(
        n1317), .A6(n4545), .Y(n4643) );
  OA222X1_HVT U1700 ( .A1(n677), .A2(n4546), .A3(n805), .A4(n4547), .A5(n933), 
        .A6(n4548), .Y(n4642) );
  OA222X1_HVT U1701 ( .A1(n293), .A2(n4549), .A3(n421), .A4(n4550), .A5(n549), 
        .A6(n4551), .Y(n4641) );
  OA22X1_HVT U1702 ( .A1(n37), .A2(n4552), .A3(n165), .A4(n4553), .Y(n4640) );
  MUX21X1_HVT U1703 ( .A1(key_round[108]), .A2(n4644), .S0(n4512), .Y(n2233)
         );
  NAND4X0_HVT U1704 ( .A1(n4645), .A2(n4646), .A3(n4647), .A4(n4648), .Y(n4644) );
  OA222X1_HVT U1705 ( .A1(n1062), .A2(n4543), .A3(n1190), .A4(n4544), .A5(
        n1318), .A6(n4545), .Y(n4648) );
  OA222X1_HVT U1706 ( .A1(n678), .A2(n4546), .A3(n806), .A4(n4547), .A5(n934), 
        .A6(n4548), .Y(n4647) );
  OA222X1_HVT U1707 ( .A1(n294), .A2(n4549), .A3(n422), .A4(n4550), .A5(n550), 
        .A6(n4551), .Y(n4646) );
  OA22X1_HVT U1708 ( .A1(n38), .A2(n4552), .A3(n166), .A4(n4553), .Y(n4645) );
  MUX21X1_HVT U1709 ( .A1(key_round[107]), .A2(n4649), .S0(n4512), .Y(n2232)
         );
  NAND4X0_HVT U1710 ( .A1(n4650), .A2(n4651), .A3(n4652), .A4(n4653), .Y(n4649) );
  OA222X1_HVT U1711 ( .A1(n1063), .A2(n4543), .A3(n1191), .A4(n4544), .A5(
        n1319), .A6(n4545), .Y(n4653) );
  OA222X1_HVT U1712 ( .A1(n679), .A2(n4546), .A3(n807), .A4(n4547), .A5(n935), 
        .A6(n4548), .Y(n4652) );
  OA222X1_HVT U1713 ( .A1(n295), .A2(n4549), .A3(n423), .A4(n4550), .A5(n551), 
        .A6(n4551), .Y(n4651) );
  OA22X1_HVT U1714 ( .A1(n39), .A2(n4552), .A3(n167), .A4(n4553), .Y(n4650) );
  MUX21X1_HVT U1715 ( .A1(key_round[106]), .A2(n4654), .S0(n4512), .Y(n2231)
         );
  NAND4X0_HVT U1716 ( .A1(n4655), .A2(n4656), .A3(n4657), .A4(n4658), .Y(n4654) );
  OA222X1_HVT U1717 ( .A1(n1064), .A2(n4543), .A3(n1192), .A4(n4544), .A5(
        n1320), .A6(n4545), .Y(n4658) );
  OA222X1_HVT U1718 ( .A1(n680), .A2(n4546), .A3(n808), .A4(n4547), .A5(n936), 
        .A6(n4548), .Y(n4657) );
  OA222X1_HVT U1719 ( .A1(n296), .A2(n4549), .A3(n424), .A4(n4550), .A5(n552), 
        .A6(n4551), .Y(n4656) );
  OA22X1_HVT U1720 ( .A1(n40), .A2(n4552), .A3(n168), .A4(n4553), .Y(n4655) );
  MUX21X1_HVT U1721 ( .A1(key_round[105]), .A2(n4659), .S0(n4512), .Y(n2230)
         );
  NAND4X0_HVT U1722 ( .A1(n4660), .A2(n4661), .A3(n4662), .A4(n4663), .Y(n4659) );
  OA222X1_HVT U1723 ( .A1(n1065), .A2(n4543), .A3(n1193), .A4(n4544), .A5(
        n1321), .A6(n4545), .Y(n4663) );
  OA222X1_HVT U1724 ( .A1(n681), .A2(n4546), .A3(n809), .A4(n4547), .A5(n937), 
        .A6(n4548), .Y(n4662) );
  OA222X1_HVT U1725 ( .A1(n297), .A2(n4549), .A3(n425), .A4(n4550), .A5(n553), 
        .A6(n4551), .Y(n4661) );
  OA22X1_HVT U1726 ( .A1(n41), .A2(n4552), .A3(n169), .A4(n4553), .Y(n4660) );
  MUX21X1_HVT U1727 ( .A1(key_round[104]), .A2(n4664), .S0(n4512), .Y(n2229)
         );
  NAND4X0_HVT U1728 ( .A1(n4665), .A2(n4666), .A3(n4667), .A4(n4668), .Y(n4664) );
  OA222X1_HVT U1729 ( .A1(n1066), .A2(n4543), .A3(n1194), .A4(n4544), .A5(
        n1322), .A6(n4545), .Y(n4668) );
  OA222X1_HVT U1730 ( .A1(n682), .A2(n4546), .A3(n810), .A4(n4547), .A5(n938), 
        .A6(n4548), .Y(n4667) );
  OA222X1_HVT U1731 ( .A1(n298), .A2(n4549), .A3(n426), .A4(n4550), .A5(n554), 
        .A6(n4551), .Y(n4666) );
  OA22X1_HVT U1732 ( .A1(n42), .A2(n4552), .A3(n170), .A4(n4553), .Y(n4665) );
  MUX21X1_HVT U1733 ( .A1(key_round[103]), .A2(n4669), .S0(n4512), .Y(n2228)
         );
  NAND4X0_HVT U1734 ( .A1(n4670), .A2(n4671), .A3(n4672), .A4(n4673), .Y(n4669) );
  OA222X1_HVT U1735 ( .A1(n1067), .A2(n4543), .A3(n1195), .A4(n4544), .A5(
        n1323), .A6(n4545), .Y(n4673) );
  OA222X1_HVT U1736 ( .A1(n683), .A2(n4546), .A3(n811), .A4(n4547), .A5(n939), 
        .A6(n4548), .Y(n4672) );
  OA222X1_HVT U1737 ( .A1(n299), .A2(n4549), .A3(n427), .A4(n4550), .A5(n555), 
        .A6(n4551), .Y(n4671) );
  OA22X1_HVT U1738 ( .A1(n43), .A2(n4552), .A3(n171), .A4(n4553), .Y(n4670) );
  MUX21X1_HVT U1739 ( .A1(key_round[102]), .A2(n4674), .S0(n4512), .Y(n2227)
         );
  NAND4X0_HVT U1740 ( .A1(n4675), .A2(n4676), .A3(n4677), .A4(n4678), .Y(n4674) );
  OA222X1_HVT U1741 ( .A1(n1068), .A2(n4543), .A3(n1196), .A4(n4544), .A5(
        n1324), .A6(n4545), .Y(n4678) );
  OA222X1_HVT U1742 ( .A1(n684), .A2(n4546), .A3(n812), .A4(n4547), .A5(n940), 
        .A6(n4548), .Y(n4677) );
  OA222X1_HVT U1743 ( .A1(n300), .A2(n4549), .A3(n428), .A4(n4550), .A5(n556), 
        .A6(n4551), .Y(n4676) );
  OA22X1_HVT U1744 ( .A1(n44), .A2(n4552), .A3(n172), .A4(n4553), .Y(n4675) );
  MUX21X1_HVT U1745 ( .A1(key_round[101]), .A2(n4679), .S0(n4512), .Y(n2226)
         );
  NAND4X0_HVT U1746 ( .A1(n4680), .A2(n4681), .A3(n4682), .A4(n4683), .Y(n4679) );
  OA222X1_HVT U1747 ( .A1(n1069), .A2(n4543), .A3(n1197), .A4(n4544), .A5(
        n1325), .A6(n4545), .Y(n4683) );
  OA222X1_HVT U1748 ( .A1(n685), .A2(n4546), .A3(n813), .A4(n4547), .A5(n941), 
        .A6(n4548), .Y(n4682) );
  OA222X1_HVT U1749 ( .A1(n301), .A2(n4549), .A3(n429), .A4(n4550), .A5(n557), 
        .A6(n4551), .Y(n4681) );
  OA22X1_HVT U1750 ( .A1(n45), .A2(n4552), .A3(n173), .A4(n4553), .Y(n4680) );
  MUX21X1_HVT U1751 ( .A1(key_round[100]), .A2(n4684), .S0(n4512), .Y(n2225)
         );
  NAND4X0_HVT U1752 ( .A1(n4685), .A2(n4686), .A3(n4687), .A4(n4688), .Y(n4684) );
  OA222X1_HVT U1753 ( .A1(n1070), .A2(n4543), .A3(n1198), .A4(n4544), .A5(
        n1326), .A6(n4545), .Y(n4688) );
  OA222X1_HVT U1754 ( .A1(n686), .A2(n4546), .A3(n814), .A4(n4547), .A5(n942), 
        .A6(n4548), .Y(n4687) );
  OA222X1_HVT U1755 ( .A1(n302), .A2(n4549), .A3(n430), .A4(n4550), .A5(n558), 
        .A6(n4551), .Y(n4686) );
  OA22X1_HVT U1756 ( .A1(n46), .A2(n4552), .A3(n174), .A4(n4553), .Y(n4685) );
  MUX21X1_HVT U1757 ( .A1(key_round[99]), .A2(n4689), .S0(n4512), .Y(n2224) );
  NAND4X0_HVT U1758 ( .A1(n4690), .A2(n4691), .A3(n4692), .A4(n4693), .Y(n4689) );
  OA222X1_HVT U1759 ( .A1(n1071), .A2(n4543), .A3(n1199), .A4(n4544), .A5(
        n1327), .A6(n4545), .Y(n4693) );
  OA222X1_HVT U1760 ( .A1(n687), .A2(n4546), .A3(n815), .A4(n4547), .A5(n943), 
        .A6(n4548), .Y(n4692) );
  OA222X1_HVT U1761 ( .A1(n303), .A2(n4549), .A3(n431), .A4(n4550), .A5(n559), 
        .A6(n4551), .Y(n4691) );
  OA22X1_HVT U1762 ( .A1(n47), .A2(n4552), .A3(n175), .A4(n4553), .Y(n4690) );
  MUX21X1_HVT U1763 ( .A1(key_round[98]), .A2(n4694), .S0(n4512), .Y(n2223) );
  NAND4X0_HVT U1764 ( .A1(n4695), .A2(n4696), .A3(n4697), .A4(n4698), .Y(n4694) );
  OA222X1_HVT U1765 ( .A1(n1072), .A2(n4543), .A3(n1200), .A4(n4544), .A5(
        n1328), .A6(n4545), .Y(n4698) );
  OA222X1_HVT U1766 ( .A1(n688), .A2(n4546), .A3(n816), .A4(n4547), .A5(n944), 
        .A6(n4548), .Y(n4697) );
  OA222X1_HVT U1767 ( .A1(n304), .A2(n4549), .A3(n432), .A4(n4550), .A5(n560), 
        .A6(n4551), .Y(n4696) );
  OA22X1_HVT U1768 ( .A1(n48), .A2(n4552), .A3(n176), .A4(n4553), .Y(n4695) );
  MUX21X1_HVT U1769 ( .A1(key_round[97]), .A2(n4699), .S0(n4512), .Y(n2222) );
  NAND4X0_HVT U1770 ( .A1(n4700), .A2(n4701), .A3(n4702), .A4(n4703), .Y(n4699) );
  OA222X1_HVT U1771 ( .A1(n1073), .A2(n4543), .A3(n1201), .A4(n4544), .A5(
        n1329), .A6(n4545), .Y(n4703) );
  OA222X1_HVT U1772 ( .A1(n689), .A2(n4546), .A3(n817), .A4(n4547), .A5(n945), 
        .A6(n4548), .Y(n4702) );
  OA222X1_HVT U1773 ( .A1(n305), .A2(n4549), .A3(n433), .A4(n4550), .A5(n561), 
        .A6(n4551), .Y(n4701) );
  OA22X1_HVT U1774 ( .A1(n49), .A2(n4552), .A3(n177), .A4(n4553), .Y(n4700) );
  MUX21X1_HVT U1775 ( .A1(key_round[96]), .A2(n4704), .S0(n4512), .Y(n2221) );
  NAND4X0_HVT U1776 ( .A1(n4705), .A2(n4706), .A3(n4707), .A4(n4708), .Y(n4704) );
  OA222X1_HVT U1777 ( .A1(n1074), .A2(n4543), .A3(n1202), .A4(n4544), .A5(
        n1330), .A6(n4545), .Y(n4708) );
  OA222X1_HVT U1778 ( .A1(n690), .A2(n4546), .A3(n818), .A4(n4547), .A5(n946), 
        .A6(n4548), .Y(n4707) );
  OA222X1_HVT U1779 ( .A1(n306), .A2(n4549), .A3(n434), .A4(n4550), .A5(n562), 
        .A6(n4551), .Y(n4706) );
  OA22X1_HVT U1780 ( .A1(n50), .A2(n4552), .A3(n178), .A4(n4553), .Y(n4705) );
  MUX21X1_HVT U1781 ( .A1(key_round[95]), .A2(n4709), .S0(n4512), .Y(n2220) );
  NAND4X0_HVT U1782 ( .A1(n4710), .A2(n4711), .A3(n4712), .A4(n4713), .Y(n4709) );
  OA222X1_HVT U1783 ( .A1(n1075), .A2(n4543), .A3(n1203), .A4(n4544), .A5(
        n1331), .A6(n4545), .Y(n4713) );
  OA222X1_HVT U1784 ( .A1(n691), .A2(n4546), .A3(n819), .A4(n4547), .A5(n947), 
        .A6(n4548), .Y(n4712) );
  OA222X1_HVT U1785 ( .A1(n307), .A2(n4549), .A3(n435), .A4(n4550), .A5(n563), 
        .A6(n4551), .Y(n4711) );
  OA22X1_HVT U1786 ( .A1(n51), .A2(n4552), .A3(n179), .A4(n4553), .Y(n4710) );
  MUX21X1_HVT U1787 ( .A1(key_round[94]), .A2(n4714), .S0(n4512), .Y(n2219) );
  NAND4X0_HVT U1788 ( .A1(n4715), .A2(n4716), .A3(n4717), .A4(n4718), .Y(n4714) );
  OA222X1_HVT U1789 ( .A1(n1076), .A2(n4543), .A3(n1204), .A4(n4544), .A5(
        n1332), .A6(n4545), .Y(n4718) );
  OA222X1_HVT U1790 ( .A1(n692), .A2(n4546), .A3(n820), .A4(n4547), .A5(n948), 
        .A6(n4548), .Y(n4717) );
  OA222X1_HVT U1791 ( .A1(n308), .A2(n4549), .A3(n436), .A4(n4550), .A5(n564), 
        .A6(n4551), .Y(n4716) );
  OA22X1_HVT U1792 ( .A1(n52), .A2(n4552), .A3(n180), .A4(n4553), .Y(n4715) );
  MUX21X1_HVT U1793 ( .A1(key_round[93]), .A2(n4719), .S0(n4512), .Y(n2218) );
  NAND4X0_HVT U1794 ( .A1(n4720), .A2(n4721), .A3(n4722), .A4(n4723), .Y(n4719) );
  OA222X1_HVT U1795 ( .A1(n1077), .A2(n4543), .A3(n1205), .A4(n4544), .A5(
        n1333), .A6(n4545), .Y(n4723) );
  OA222X1_HVT U1796 ( .A1(n693), .A2(n4546), .A3(n821), .A4(n4547), .A5(n949), 
        .A6(n4548), .Y(n4722) );
  OA222X1_HVT U1797 ( .A1(n309), .A2(n4549), .A3(n437), .A4(n4550), .A5(n565), 
        .A6(n4551), .Y(n4721) );
  OA22X1_HVT U1798 ( .A1(n53), .A2(n4552), .A3(n181), .A4(n4553), .Y(n4720) );
  MUX21X1_HVT U1799 ( .A1(key_round[92]), .A2(n4724), .S0(n4512), .Y(n2217) );
  NAND4X0_HVT U1800 ( .A1(n4725), .A2(n4726), .A3(n4727), .A4(n4728), .Y(n4724) );
  OA222X1_HVT U1801 ( .A1(n1078), .A2(n4543), .A3(n1206), .A4(n4544), .A5(
        n1334), .A6(n4545), .Y(n4728) );
  OA222X1_HVT U1802 ( .A1(n694), .A2(n4546), .A3(n822), .A4(n4547), .A5(n950), 
        .A6(n4548), .Y(n4727) );
  OA222X1_HVT U1803 ( .A1(n310), .A2(n4549), .A3(n438), .A4(n4550), .A5(n566), 
        .A6(n4551), .Y(n4726) );
  OA22X1_HVT U1804 ( .A1(n54), .A2(n4552), .A3(n182), .A4(n4553), .Y(n4725) );
  MUX21X1_HVT U1805 ( .A1(key_round[91]), .A2(n4729), .S0(n4512), .Y(n2216) );
  NAND4X0_HVT U1806 ( .A1(n4730), .A2(n4731), .A3(n4732), .A4(n4733), .Y(n4729) );
  OA222X1_HVT U1807 ( .A1(n1079), .A2(n4543), .A3(n1207), .A4(n4544), .A5(
        n1335), .A6(n4545), .Y(n4733) );
  OA222X1_HVT U1808 ( .A1(n695), .A2(n4546), .A3(n823), .A4(n4547), .A5(n951), 
        .A6(n4548), .Y(n4732) );
  OA222X1_HVT U1809 ( .A1(n311), .A2(n4549), .A3(n439), .A4(n4550), .A5(n567), 
        .A6(n4551), .Y(n4731) );
  OA22X1_HVT U1810 ( .A1(n55), .A2(n4552), .A3(n183), .A4(n4553), .Y(n4730) );
  MUX21X1_HVT U1811 ( .A1(key_round[90]), .A2(n4734), .S0(n4512), .Y(n2215) );
  NAND4X0_HVT U1812 ( .A1(n4735), .A2(n4736), .A3(n4737), .A4(n4738), .Y(n4734) );
  OA222X1_HVT U1813 ( .A1(n1080), .A2(n4543), .A3(n1208), .A4(n4544), .A5(
        n1336), .A6(n4545), .Y(n4738) );
  OA222X1_HVT U1814 ( .A1(n696), .A2(n4546), .A3(n824), .A4(n4547), .A5(n952), 
        .A6(n4548), .Y(n4737) );
  OA222X1_HVT U1815 ( .A1(n312), .A2(n4549), .A3(n440), .A4(n4550), .A5(n568), 
        .A6(n4551), .Y(n4736) );
  OA22X1_HVT U1816 ( .A1(n56), .A2(n4552), .A3(n184), .A4(n4553), .Y(n4735) );
  MUX21X1_HVT U1817 ( .A1(key_round[89]), .A2(n4739), .S0(n4512), .Y(n2214) );
  NAND4X0_HVT U1818 ( .A1(n4740), .A2(n4741), .A3(n4742), .A4(n4743), .Y(n4739) );
  OA222X1_HVT U1819 ( .A1(n1081), .A2(n4543), .A3(n1209), .A4(n4544), .A5(
        n1337), .A6(n4545), .Y(n4743) );
  OA222X1_HVT U1820 ( .A1(n697), .A2(n4546), .A3(n825), .A4(n4547), .A5(n953), 
        .A6(n4548), .Y(n4742) );
  OA222X1_HVT U1821 ( .A1(n313), .A2(n4549), .A3(n441), .A4(n4550), .A5(n569), 
        .A6(n4551), .Y(n4741) );
  OA22X1_HVT U1822 ( .A1(n57), .A2(n4552), .A3(n185), .A4(n4553), .Y(n4740) );
  MUX21X1_HVT U1823 ( .A1(key_round[88]), .A2(n4744), .S0(n4512), .Y(n2213) );
  NAND4X0_HVT U1824 ( .A1(n4745), .A2(n4746), .A3(n4747), .A4(n4748), .Y(n4744) );
  OA222X1_HVT U1825 ( .A1(n1082), .A2(n4543), .A3(n1210), .A4(n4544), .A5(
        n1338), .A6(n4545), .Y(n4748) );
  OA222X1_HVT U1826 ( .A1(n698), .A2(n4546), .A3(n826), .A4(n4547), .A5(n954), 
        .A6(n4548), .Y(n4747) );
  OA222X1_HVT U1827 ( .A1(n314), .A2(n4549), .A3(n442), .A4(n4550), .A5(n570), 
        .A6(n4551), .Y(n4746) );
  OA22X1_HVT U1828 ( .A1(n58), .A2(n4552), .A3(n186), .A4(n4553), .Y(n4745) );
  MUX21X1_HVT U1829 ( .A1(key_round[87]), .A2(n4749), .S0(n4512), .Y(n2212) );
  NAND4X0_HVT U1830 ( .A1(n4750), .A2(n4751), .A3(n4752), .A4(n4753), .Y(n4749) );
  OA222X1_HVT U1831 ( .A1(n1083), .A2(n4543), .A3(n1211), .A4(n4544), .A5(
        n1339), .A6(n4545), .Y(n4753) );
  OA222X1_HVT U1832 ( .A1(n699), .A2(n4546), .A3(n827), .A4(n4547), .A5(n955), 
        .A6(n4548), .Y(n4752) );
  OA222X1_HVT U1833 ( .A1(n315), .A2(n4549), .A3(n443), .A4(n4550), .A5(n571), 
        .A6(n4551), .Y(n4751) );
  OA22X1_HVT U1834 ( .A1(n59), .A2(n4552), .A3(n187), .A4(n4553), .Y(n4750) );
  MUX21X1_HVT U1835 ( .A1(key_round[86]), .A2(n4754), .S0(n4512), .Y(n2211) );
  NAND4X0_HVT U1836 ( .A1(n4755), .A2(n4756), .A3(n4757), .A4(n4758), .Y(n4754) );
  OA222X1_HVT U1837 ( .A1(n1084), .A2(n4543), .A3(n1212), .A4(n4544), .A5(
        n1340), .A6(n4545), .Y(n4758) );
  OA222X1_HVT U1838 ( .A1(n700), .A2(n4546), .A3(n828), .A4(n4547), .A5(n956), 
        .A6(n4548), .Y(n4757) );
  OA222X1_HVT U1839 ( .A1(n316), .A2(n4549), .A3(n444), .A4(n4550), .A5(n572), 
        .A6(n4551), .Y(n4756) );
  OA22X1_HVT U1840 ( .A1(n60), .A2(n4552), .A3(n188), .A4(n4553), .Y(n4755) );
  MUX21X1_HVT U1841 ( .A1(key_round[85]), .A2(n4759), .S0(n4512), .Y(n2210) );
  NAND4X0_HVT U1842 ( .A1(n4760), .A2(n4761), .A3(n4762), .A4(n4763), .Y(n4759) );
  OA222X1_HVT U1843 ( .A1(n1085), .A2(n4543), .A3(n1213), .A4(n4544), .A5(
        n1341), .A6(n4545), .Y(n4763) );
  OA222X1_HVT U1844 ( .A1(n701), .A2(n4546), .A3(n829), .A4(n4547), .A5(n957), 
        .A6(n4548), .Y(n4762) );
  OA222X1_HVT U1845 ( .A1(n317), .A2(n4549), .A3(n445), .A4(n4550), .A5(n573), 
        .A6(n4551), .Y(n4761) );
  OA22X1_HVT U1846 ( .A1(n61), .A2(n4552), .A3(n189), .A4(n4553), .Y(n4760) );
  MUX21X1_HVT U1847 ( .A1(key_round[84]), .A2(n4764), .S0(n4512), .Y(n2209) );
  NAND4X0_HVT U1848 ( .A1(n4765), .A2(n4766), .A3(n4767), .A4(n4768), .Y(n4764) );
  OA222X1_HVT U1849 ( .A1(n1086), .A2(n4543), .A3(n1214), .A4(n4544), .A5(
        n1342), .A6(n4545), .Y(n4768) );
  OA222X1_HVT U1850 ( .A1(n702), .A2(n4546), .A3(n830), .A4(n4547), .A5(n958), 
        .A6(n4548), .Y(n4767) );
  OA222X1_HVT U1851 ( .A1(n318), .A2(n4549), .A3(n446), .A4(n4550), .A5(n574), 
        .A6(n4551), .Y(n4766) );
  OA22X1_HVT U1852 ( .A1(n62), .A2(n4552), .A3(n190), .A4(n4553), .Y(n4765) );
  MUX21X1_HVT U1853 ( .A1(key_round[83]), .A2(n4769), .S0(n4512), .Y(n2208) );
  NAND4X0_HVT U1854 ( .A1(n4770), .A2(n4771), .A3(n4772), .A4(n4773), .Y(n4769) );
  OA222X1_HVT U1855 ( .A1(n1087), .A2(n4543), .A3(n1215), .A4(n4544), .A5(
        n1343), .A6(n4545), .Y(n4773) );
  OA222X1_HVT U1856 ( .A1(n703), .A2(n4546), .A3(n831), .A4(n4547), .A5(n959), 
        .A6(n4548), .Y(n4772) );
  OA222X1_HVT U1857 ( .A1(n319), .A2(n4549), .A3(n447), .A4(n4550), .A5(n575), 
        .A6(n4551), .Y(n4771) );
  OA22X1_HVT U1858 ( .A1(n63), .A2(n4552), .A3(n191), .A4(n4553), .Y(n4770) );
  MUX21X1_HVT U1859 ( .A1(key_round[82]), .A2(n4774), .S0(n4512), .Y(n2207) );
  NAND4X0_HVT U1860 ( .A1(n4775), .A2(n4776), .A3(n4777), .A4(n4778), .Y(n4774) );
  OA222X1_HVT U1861 ( .A1(n1088), .A2(n4543), .A3(n1216), .A4(n4544), .A5(
        n1344), .A6(n4545), .Y(n4778) );
  OA222X1_HVT U1862 ( .A1(n704), .A2(n4546), .A3(n832), .A4(n4547), .A5(n960), 
        .A6(n4548), .Y(n4777) );
  OA222X1_HVT U1863 ( .A1(n320), .A2(n4549), .A3(n448), .A4(n4550), .A5(n576), 
        .A6(n4551), .Y(n4776) );
  OA22X1_HVT U1864 ( .A1(n64), .A2(n4552), .A3(n192), .A4(n4553), .Y(n4775) );
  MUX21X1_HVT U1865 ( .A1(key_round[81]), .A2(n4779), .S0(n4512), .Y(n2206) );
  NAND4X0_HVT U1866 ( .A1(n4780), .A2(n4781), .A3(n4782), .A4(n4783), .Y(n4779) );
  OA222X1_HVT U1867 ( .A1(n1089), .A2(n4543), .A3(n1217), .A4(n4544), .A5(
        n1345), .A6(n4545), .Y(n4783) );
  OA222X1_HVT U1868 ( .A1(n705), .A2(n4546), .A3(n833), .A4(n4547), .A5(n961), 
        .A6(n4548), .Y(n4782) );
  OA222X1_HVT U1869 ( .A1(n321), .A2(n4549), .A3(n449), .A4(n4550), .A5(n577), 
        .A6(n4551), .Y(n4781) );
  OA22X1_HVT U1870 ( .A1(n65), .A2(n4552), .A3(n193), .A4(n4553), .Y(n4780) );
  MUX21X1_HVT U1871 ( .A1(key_round[80]), .A2(n4784), .S0(n4512), .Y(n2205) );
  NAND4X0_HVT U1872 ( .A1(n4785), .A2(n4786), .A3(n4787), .A4(n4788), .Y(n4784) );
  OA222X1_HVT U1873 ( .A1(n1090), .A2(n4543), .A3(n1218), .A4(n4544), .A5(
        n1346), .A6(n4545), .Y(n4788) );
  OA222X1_HVT U1874 ( .A1(n706), .A2(n4546), .A3(n834), .A4(n4547), .A5(n962), 
        .A6(n4548), .Y(n4787) );
  OA222X1_HVT U1875 ( .A1(n322), .A2(n4549), .A3(n450), .A4(n4550), .A5(n578), 
        .A6(n4551), .Y(n4786) );
  OA22X1_HVT U1876 ( .A1(n66), .A2(n4552), .A3(n194), .A4(n4553), .Y(n4785) );
  MUX21X1_HVT U1877 ( .A1(key_round[79]), .A2(n4789), .S0(n4512), .Y(n2204) );
  NAND4X0_HVT U1878 ( .A1(n4790), .A2(n4791), .A3(n4792), .A4(n4793), .Y(n4789) );
  OA222X1_HVT U1879 ( .A1(n1091), .A2(n4543), .A3(n1219), .A4(n4544), .A5(
        n1347), .A6(n4545), .Y(n4793) );
  OA222X1_HVT U1880 ( .A1(n707), .A2(n4546), .A3(n835), .A4(n4547), .A5(n963), 
        .A6(n4548), .Y(n4792) );
  OA222X1_HVT U1881 ( .A1(n323), .A2(n4549), .A3(n451), .A4(n4550), .A5(n579), 
        .A6(n4551), .Y(n4791) );
  OA22X1_HVT U1882 ( .A1(n67), .A2(n4552), .A3(n195), .A4(n4553), .Y(n4790) );
  MUX21X1_HVT U1883 ( .A1(key_round[78]), .A2(n4794), .S0(n4512), .Y(n2203) );
  NAND4X0_HVT U1884 ( .A1(n4795), .A2(n4796), .A3(n4797), .A4(n4798), .Y(n4794) );
  OA222X1_HVT U1885 ( .A1(n1092), .A2(n4543), .A3(n1220), .A4(n4544), .A5(
        n1348), .A6(n4545), .Y(n4798) );
  OA222X1_HVT U1886 ( .A1(n708), .A2(n4546), .A3(n836), .A4(n4547), .A5(n964), 
        .A6(n4548), .Y(n4797) );
  OA222X1_HVT U1887 ( .A1(n324), .A2(n4549), .A3(n452), .A4(n4550), .A5(n580), 
        .A6(n4551), .Y(n4796) );
  OA22X1_HVT U1888 ( .A1(n68), .A2(n4552), .A3(n196), .A4(n4553), .Y(n4795) );
  MUX21X1_HVT U1889 ( .A1(key_round[77]), .A2(n4799), .S0(n4512), .Y(n2202) );
  NAND4X0_HVT U1890 ( .A1(n4800), .A2(n4801), .A3(n4802), .A4(n4803), .Y(n4799) );
  OA222X1_HVT U1891 ( .A1(n1093), .A2(n4543), .A3(n1221), .A4(n4544), .A5(
        n1349), .A6(n4545), .Y(n4803) );
  OA222X1_HVT U1892 ( .A1(n709), .A2(n4546), .A3(n837), .A4(n4547), .A5(n965), 
        .A6(n4548), .Y(n4802) );
  OA222X1_HVT U1893 ( .A1(n325), .A2(n4549), .A3(n453), .A4(n4550), .A5(n581), 
        .A6(n4551), .Y(n4801) );
  OA22X1_HVT U1894 ( .A1(n69), .A2(n4552), .A3(n197), .A4(n4553), .Y(n4800) );
  MUX21X1_HVT U1895 ( .A1(key_round[76]), .A2(n4804), .S0(n4512), .Y(n2201) );
  NAND4X0_HVT U1896 ( .A1(n4805), .A2(n4806), .A3(n4807), .A4(n4808), .Y(n4804) );
  OA222X1_HVT U1897 ( .A1(n1094), .A2(n4543), .A3(n1222), .A4(n4544), .A5(
        n1350), .A6(n4545), .Y(n4808) );
  OA222X1_HVT U1898 ( .A1(n710), .A2(n4546), .A3(n838), .A4(n4547), .A5(n966), 
        .A6(n4548), .Y(n4807) );
  OA222X1_HVT U1899 ( .A1(n326), .A2(n4549), .A3(n454), .A4(n4550), .A5(n582), 
        .A6(n4551), .Y(n4806) );
  OA22X1_HVT U1900 ( .A1(n70), .A2(n4552), .A3(n198), .A4(n4553), .Y(n4805) );
  MUX21X1_HVT U1901 ( .A1(key_round[75]), .A2(n4809), .S0(n4512), .Y(n2200) );
  NAND4X0_HVT U1902 ( .A1(n4810), .A2(n4811), .A3(n4812), .A4(n4813), .Y(n4809) );
  OA222X1_HVT U1903 ( .A1(n1095), .A2(n4543), .A3(n1223), .A4(n4544), .A5(
        n1351), .A6(n4545), .Y(n4813) );
  OA222X1_HVT U1904 ( .A1(n711), .A2(n4546), .A3(n839), .A4(n4547), .A5(n967), 
        .A6(n4548), .Y(n4812) );
  OA222X1_HVT U1905 ( .A1(n327), .A2(n4549), .A3(n455), .A4(n4550), .A5(n583), 
        .A6(n4551), .Y(n4811) );
  OA22X1_HVT U1906 ( .A1(n71), .A2(n4552), .A3(n199), .A4(n4553), .Y(n4810) );
  MUX21X1_HVT U1907 ( .A1(key_round[74]), .A2(n4814), .S0(n4512), .Y(n2199) );
  NAND4X0_HVT U1908 ( .A1(n4815), .A2(n4816), .A3(n4817), .A4(n4818), .Y(n4814) );
  OA222X1_HVT U1909 ( .A1(n1096), .A2(n4543), .A3(n1224), .A4(n4544), .A5(
        n1352), .A6(n4545), .Y(n4818) );
  OA222X1_HVT U1910 ( .A1(n712), .A2(n4546), .A3(n840), .A4(n4547), .A5(n968), 
        .A6(n4548), .Y(n4817) );
  OA222X1_HVT U1911 ( .A1(n328), .A2(n4549), .A3(n456), .A4(n4550), .A5(n584), 
        .A6(n4551), .Y(n4816) );
  OA22X1_HVT U1912 ( .A1(n72), .A2(n4552), .A3(n200), .A4(n4553), .Y(n4815) );
  MUX21X1_HVT U1913 ( .A1(key_round[73]), .A2(n4819), .S0(n4512), .Y(n2198) );
  NAND4X0_HVT U1914 ( .A1(n4820), .A2(n4821), .A3(n4822), .A4(n4823), .Y(n4819) );
  OA222X1_HVT U1915 ( .A1(n1097), .A2(n4543), .A3(n1225), .A4(n4544), .A5(
        n1353), .A6(n4545), .Y(n4823) );
  OA222X1_HVT U1916 ( .A1(n713), .A2(n4546), .A3(n841), .A4(n4547), .A5(n969), 
        .A6(n4548), .Y(n4822) );
  OA222X1_HVT U1917 ( .A1(n329), .A2(n4549), .A3(n457), .A4(n4550), .A5(n585), 
        .A6(n4551), .Y(n4821) );
  OA22X1_HVT U1918 ( .A1(n73), .A2(n4552), .A3(n201), .A4(n4553), .Y(n4820) );
  MUX21X1_HVT U1919 ( .A1(key_round[72]), .A2(n4824), .S0(n4512), .Y(n2197) );
  NAND4X0_HVT U1920 ( .A1(n4825), .A2(n4826), .A3(n4827), .A4(n4828), .Y(n4824) );
  OA222X1_HVT U1921 ( .A1(n1098), .A2(n4543), .A3(n1226), .A4(n4544), .A5(
        n1354), .A6(n4545), .Y(n4828) );
  OA222X1_HVT U1922 ( .A1(n714), .A2(n4546), .A3(n842), .A4(n4547), .A5(n970), 
        .A6(n4548), .Y(n4827) );
  OA222X1_HVT U1923 ( .A1(n330), .A2(n4549), .A3(n458), .A4(n4550), .A5(n586), 
        .A6(n4551), .Y(n4826) );
  OA22X1_HVT U1924 ( .A1(n74), .A2(n4552), .A3(n202), .A4(n4553), .Y(n4825) );
  MUX21X1_HVT U1925 ( .A1(key_round[71]), .A2(n4829), .S0(n4512), .Y(n2196) );
  NAND4X0_HVT U1926 ( .A1(n4830), .A2(n4831), .A3(n4832), .A4(n4833), .Y(n4829) );
  OA222X1_HVT U1927 ( .A1(n1099), .A2(n4543), .A3(n1227), .A4(n4544), .A5(
        n1355), .A6(n4545), .Y(n4833) );
  OA222X1_HVT U1928 ( .A1(n715), .A2(n4546), .A3(n843), .A4(n4547), .A5(n971), 
        .A6(n4548), .Y(n4832) );
  OA222X1_HVT U1929 ( .A1(n331), .A2(n4549), .A3(n459), .A4(n4550), .A5(n587), 
        .A6(n4551), .Y(n4831) );
  OA22X1_HVT U1930 ( .A1(n75), .A2(n4552), .A3(n203), .A4(n4553), .Y(n4830) );
  MUX21X1_HVT U1931 ( .A1(key_round[70]), .A2(n4834), .S0(n4512), .Y(n2195) );
  NAND4X0_HVT U1932 ( .A1(n4835), .A2(n4836), .A3(n4837), .A4(n4838), .Y(n4834) );
  OA222X1_HVT U1933 ( .A1(n1100), .A2(n4543), .A3(n1228), .A4(n4544), .A5(
        n1356), .A6(n4545), .Y(n4838) );
  OA222X1_HVT U1934 ( .A1(n716), .A2(n4546), .A3(n844), .A4(n4547), .A5(n972), 
        .A6(n4548), .Y(n4837) );
  OA222X1_HVT U1935 ( .A1(n332), .A2(n4549), .A3(n460), .A4(n4550), .A5(n588), 
        .A6(n4551), .Y(n4836) );
  OA22X1_HVT U1936 ( .A1(n76), .A2(n4552), .A3(n204), .A4(n4553), .Y(n4835) );
  MUX21X1_HVT U1937 ( .A1(key_round[69]), .A2(n4839), .S0(n4512), .Y(n2194) );
  NAND4X0_HVT U1938 ( .A1(n4840), .A2(n4841), .A3(n4842), .A4(n4843), .Y(n4839) );
  OA222X1_HVT U1939 ( .A1(n1101), .A2(n4543), .A3(n1229), .A4(n4544), .A5(
        n1357), .A6(n4545), .Y(n4843) );
  OA222X1_HVT U1940 ( .A1(n717), .A2(n4546), .A3(n845), .A4(n4547), .A5(n973), 
        .A6(n4548), .Y(n4842) );
  OA222X1_HVT U1941 ( .A1(n333), .A2(n4549), .A3(n461), .A4(n4550), .A5(n589), 
        .A6(n4551), .Y(n4841) );
  OA22X1_HVT U1942 ( .A1(n77), .A2(n4552), .A3(n205), .A4(n4553), .Y(n4840) );
  MUX21X1_HVT U1943 ( .A1(key_round[68]), .A2(n4844), .S0(n4512), .Y(n2193) );
  NAND4X0_HVT U1944 ( .A1(n4845), .A2(n4846), .A3(n4847), .A4(n4848), .Y(n4844) );
  OA222X1_HVT U1945 ( .A1(n1102), .A2(n4543), .A3(n1230), .A4(n4544), .A5(
        n1358), .A6(n4545), .Y(n4848) );
  OA222X1_HVT U1946 ( .A1(n718), .A2(n4546), .A3(n846), .A4(n4547), .A5(n974), 
        .A6(n4548), .Y(n4847) );
  OA222X1_HVT U1947 ( .A1(n334), .A2(n4549), .A3(n462), .A4(n4550), .A5(n590), 
        .A6(n4551), .Y(n4846) );
  OA22X1_HVT U1948 ( .A1(n78), .A2(n4552), .A3(n206), .A4(n4553), .Y(n4845) );
  MUX21X1_HVT U1949 ( .A1(key_round[67]), .A2(n4849), .S0(n4512), .Y(n2192) );
  NAND4X0_HVT U1950 ( .A1(n4850), .A2(n4851), .A3(n4852), .A4(n4853), .Y(n4849) );
  OA222X1_HVT U1951 ( .A1(n1103), .A2(n4543), .A3(n1231), .A4(n4544), .A5(
        n1359), .A6(n4545), .Y(n4853) );
  OA222X1_HVT U1952 ( .A1(n719), .A2(n4546), .A3(n847), .A4(n4547), .A5(n975), 
        .A6(n4548), .Y(n4852) );
  OA222X1_HVT U1953 ( .A1(n335), .A2(n4549), .A3(n463), .A4(n4550), .A5(n591), 
        .A6(n4551), .Y(n4851) );
  OA22X1_HVT U1954 ( .A1(n79), .A2(n4552), .A3(n207), .A4(n4553), .Y(n4850) );
  MUX21X1_HVT U1955 ( .A1(key_round[66]), .A2(n4854), .S0(n4512), .Y(n2191) );
  NAND4X0_HVT U1956 ( .A1(n4855), .A2(n4856), .A3(n4857), .A4(n4858), .Y(n4854) );
  OA222X1_HVT U1957 ( .A1(n1104), .A2(n4543), .A3(n1232), .A4(n4544), .A5(
        n1360), .A6(n4545), .Y(n4858) );
  OA222X1_HVT U1958 ( .A1(n720), .A2(n4546), .A3(n848), .A4(n4547), .A5(n976), 
        .A6(n4548), .Y(n4857) );
  OA222X1_HVT U1959 ( .A1(n336), .A2(n4549), .A3(n464), .A4(n4550), .A5(n592), 
        .A6(n4551), .Y(n4856) );
  OA22X1_HVT U1960 ( .A1(n80), .A2(n4552), .A3(n208), .A4(n4553), .Y(n4855) );
  MUX21X1_HVT U1961 ( .A1(key_round[65]), .A2(n4859), .S0(n4512), .Y(n2190) );
  NAND4X0_HVT U1962 ( .A1(n4860), .A2(n4861), .A3(n4862), .A4(n4863), .Y(n4859) );
  OA222X1_HVT U1963 ( .A1(n1105), .A2(n4543), .A3(n1233), .A4(n4544), .A5(
        n1361), .A6(n4545), .Y(n4863) );
  OA222X1_HVT U1964 ( .A1(n721), .A2(n4546), .A3(n849), .A4(n4547), .A5(n977), 
        .A6(n4548), .Y(n4862) );
  OA222X1_HVT U1965 ( .A1(n337), .A2(n4549), .A3(n465), .A4(n4550), .A5(n593), 
        .A6(n4551), .Y(n4861) );
  OA22X1_HVT U1966 ( .A1(n81), .A2(n4552), .A3(n209), .A4(n4553), .Y(n4860) );
  MUX21X1_HVT U1967 ( .A1(key_round[64]), .A2(n4864), .S0(n4512), .Y(n2189) );
  NAND4X0_HVT U1968 ( .A1(n4865), .A2(n4866), .A3(n4867), .A4(n4868), .Y(n4864) );
  OA222X1_HVT U1969 ( .A1(n1106), .A2(n4543), .A3(n1234), .A4(n4544), .A5(
        n1362), .A6(n4545), .Y(n4868) );
  OA222X1_HVT U1970 ( .A1(n722), .A2(n4546), .A3(n850), .A4(n4547), .A5(n978), 
        .A6(n4548), .Y(n4867) );
  OA222X1_HVT U1971 ( .A1(n338), .A2(n4549), .A3(n466), .A4(n4550), .A5(n594), 
        .A6(n4551), .Y(n4866) );
  OA22X1_HVT U1972 ( .A1(n82), .A2(n4552), .A3(n210), .A4(n4553), .Y(n4865) );
  MUX21X1_HVT U1973 ( .A1(key_round[63]), .A2(n4869), .S0(n4512), .Y(n2188) );
  NAND4X0_HVT U1974 ( .A1(n4870), .A2(n4871), .A3(n4872), .A4(n4873), .Y(n4869) );
  OA222X1_HVT U1975 ( .A1(n1107), .A2(n4543), .A3(n1235), .A4(n4544), .A5(
        n1363), .A6(n4545), .Y(n4873) );
  OA222X1_HVT U1976 ( .A1(n723), .A2(n4546), .A3(n851), .A4(n4547), .A5(n979), 
        .A6(n4548), .Y(n4872) );
  OA222X1_HVT U1977 ( .A1(n339), .A2(n4549), .A3(n467), .A4(n4550), .A5(n595), 
        .A6(n4551), .Y(n4871) );
  OA22X1_HVT U1978 ( .A1(n83), .A2(n4552), .A3(n211), .A4(n4553), .Y(n4870) );
  MUX21X1_HVT U1979 ( .A1(key_round[62]), .A2(n4874), .S0(n4512), .Y(n2187) );
  NAND4X0_HVT U1980 ( .A1(n4875), .A2(n4876), .A3(n4877), .A4(n4878), .Y(n4874) );
  OA222X1_HVT U1981 ( .A1(n1108), .A2(n4543), .A3(n1236), .A4(n4544), .A5(
        n1364), .A6(n4545), .Y(n4878) );
  OA222X1_HVT U1982 ( .A1(n724), .A2(n4546), .A3(n852), .A4(n4547), .A5(n980), 
        .A6(n4548), .Y(n4877) );
  OA222X1_HVT U1983 ( .A1(n340), .A2(n4549), .A3(n468), .A4(n4550), .A5(n596), 
        .A6(n4551), .Y(n4876) );
  OA22X1_HVT U1984 ( .A1(n84), .A2(n4552), .A3(n212), .A4(n4553), .Y(n4875) );
  MUX21X1_HVT U1985 ( .A1(key_round[61]), .A2(n4879), .S0(n4512), .Y(n2186) );
  NAND4X0_HVT U1986 ( .A1(n4880), .A2(n4881), .A3(n4882), .A4(n4883), .Y(n4879) );
  OA222X1_HVT U1987 ( .A1(n1109), .A2(n4543), .A3(n1237), .A4(n4544), .A5(
        n1365), .A6(n4545), .Y(n4883) );
  OA222X1_HVT U1988 ( .A1(n725), .A2(n4546), .A3(n853), .A4(n4547), .A5(n981), 
        .A6(n4548), .Y(n4882) );
  OA222X1_HVT U1989 ( .A1(n341), .A2(n4549), .A3(n469), .A4(n4550), .A5(n597), 
        .A6(n4551), .Y(n4881) );
  OA22X1_HVT U1990 ( .A1(n85), .A2(n4552), .A3(n213), .A4(n4553), .Y(n4880) );
  MUX21X1_HVT U1991 ( .A1(key_round[60]), .A2(n4884), .S0(n4512), .Y(n2185) );
  NAND4X0_HVT U1992 ( .A1(n4885), .A2(n4886), .A3(n4887), .A4(n4888), .Y(n4884) );
  OA222X1_HVT U1993 ( .A1(n1110), .A2(n4543), .A3(n1238), .A4(n4544), .A5(
        n1366), .A6(n4545), .Y(n4888) );
  OA222X1_HVT U1994 ( .A1(n726), .A2(n4546), .A3(n854), .A4(n4547), .A5(n982), 
        .A6(n4548), .Y(n4887) );
  OA222X1_HVT U1995 ( .A1(n342), .A2(n4549), .A3(n470), .A4(n4550), .A5(n598), 
        .A6(n4551), .Y(n4886) );
  OA22X1_HVT U1996 ( .A1(n86), .A2(n4552), .A3(n214), .A4(n4553), .Y(n4885) );
  MUX21X1_HVT U1997 ( .A1(key_round[59]), .A2(n4889), .S0(n4512), .Y(n2184) );
  NAND4X0_HVT U1998 ( .A1(n4890), .A2(n4891), .A3(n4892), .A4(n4893), .Y(n4889) );
  OA222X1_HVT U1999 ( .A1(n1111), .A2(n4543), .A3(n1239), .A4(n4544), .A5(
        n1367), .A6(n4545), .Y(n4893) );
  OA222X1_HVT U2000 ( .A1(n727), .A2(n4546), .A3(n855), .A4(n4547), .A5(n983), 
        .A6(n4548), .Y(n4892) );
  OA222X1_HVT U2001 ( .A1(n343), .A2(n4549), .A3(n471), .A4(n4550), .A5(n599), 
        .A6(n4551), .Y(n4891) );
  OA22X1_HVT U2002 ( .A1(n87), .A2(n4552), .A3(n215), .A4(n4553), .Y(n4890) );
  MUX21X1_HVT U2003 ( .A1(key_round[58]), .A2(n4894), .S0(n4512), .Y(n2183) );
  NAND4X0_HVT U2004 ( .A1(n4895), .A2(n4896), .A3(n4897), .A4(n4898), .Y(n4894) );
  OA222X1_HVT U2005 ( .A1(n1112), .A2(n4543), .A3(n1240), .A4(n4544), .A5(
        n1368), .A6(n4545), .Y(n4898) );
  OA222X1_HVT U2006 ( .A1(n728), .A2(n4546), .A3(n856), .A4(n4547), .A5(n984), 
        .A6(n4548), .Y(n4897) );
  OA222X1_HVT U2007 ( .A1(n344), .A2(n4549), .A3(n472), .A4(n4550), .A5(n600), 
        .A6(n4551), .Y(n4896) );
  OA22X1_HVT U2008 ( .A1(n88), .A2(n4552), .A3(n216), .A4(n4553), .Y(n4895) );
  MUX21X1_HVT U2009 ( .A1(key_round[57]), .A2(n4899), .S0(n4512), .Y(n2182) );
  NAND4X0_HVT U2010 ( .A1(n4900), .A2(n4901), .A3(n4902), .A4(n4903), .Y(n4899) );
  OA222X1_HVT U2011 ( .A1(n1113), .A2(n4543), .A3(n1241), .A4(n4544), .A5(
        n1369), .A6(n4545), .Y(n4903) );
  OA222X1_HVT U2012 ( .A1(n729), .A2(n4546), .A3(n857), .A4(n4547), .A5(n985), 
        .A6(n4548), .Y(n4902) );
  OA222X1_HVT U2013 ( .A1(n345), .A2(n4549), .A3(n473), .A4(n4550), .A5(n601), 
        .A6(n4551), .Y(n4901) );
  OA22X1_HVT U2014 ( .A1(n89), .A2(n4552), .A3(n217), .A4(n4553), .Y(n4900) );
  MUX21X1_HVT U2015 ( .A1(key_round[56]), .A2(n4904), .S0(n4512), .Y(n2181) );
  NAND4X0_HVT U2016 ( .A1(n4905), .A2(n4906), .A3(n4907), .A4(n4908), .Y(n4904) );
  OA222X1_HVT U2017 ( .A1(n1114), .A2(n4543), .A3(n1242), .A4(n4544), .A5(
        n1370), .A6(n4545), .Y(n4908) );
  OA222X1_HVT U2018 ( .A1(n730), .A2(n4546), .A3(n858), .A4(n4547), .A5(n986), 
        .A6(n4548), .Y(n4907) );
  OA222X1_HVT U2019 ( .A1(n346), .A2(n4549), .A3(n474), .A4(n4550), .A5(n602), 
        .A6(n4551), .Y(n4906) );
  OA22X1_HVT U2020 ( .A1(n90), .A2(n4552), .A3(n218), .A4(n4553), .Y(n4905) );
  MUX21X1_HVT U2021 ( .A1(key_round[55]), .A2(n4909), .S0(n4512), .Y(n2180) );
  NAND4X0_HVT U2022 ( .A1(n4910), .A2(n4911), .A3(n4912), .A4(n4913), .Y(n4909) );
  OA222X1_HVT U2023 ( .A1(n1115), .A2(n4543), .A3(n1243), .A4(n4544), .A5(
        n1371), .A6(n4545), .Y(n4913) );
  OA222X1_HVT U2024 ( .A1(n731), .A2(n4546), .A3(n859), .A4(n4547), .A5(n987), 
        .A6(n4548), .Y(n4912) );
  OA222X1_HVT U2025 ( .A1(n347), .A2(n4549), .A3(n475), .A4(n4550), .A5(n603), 
        .A6(n4551), .Y(n4911) );
  OA22X1_HVT U2026 ( .A1(n91), .A2(n4552), .A3(n219), .A4(n4553), .Y(n4910) );
  MUX21X1_HVT U2027 ( .A1(key_round[54]), .A2(n4914), .S0(n4512), .Y(n2179) );
  NAND4X0_HVT U2028 ( .A1(n4915), .A2(n4916), .A3(n4917), .A4(n4918), .Y(n4914) );
  OA222X1_HVT U2029 ( .A1(n1116), .A2(n4543), .A3(n1244), .A4(n4544), .A5(
        n1372), .A6(n4545), .Y(n4918) );
  OA222X1_HVT U2030 ( .A1(n732), .A2(n4546), .A3(n860), .A4(n4547), .A5(n988), 
        .A6(n4548), .Y(n4917) );
  OA222X1_HVT U2031 ( .A1(n348), .A2(n4549), .A3(n476), .A4(n4550), .A5(n604), 
        .A6(n4551), .Y(n4916) );
  OA22X1_HVT U2032 ( .A1(n92), .A2(n4552), .A3(n220), .A4(n4553), .Y(n4915) );
  MUX21X1_HVT U2033 ( .A1(key_round[53]), .A2(n4919), .S0(n4512), .Y(n2178) );
  NAND4X0_HVT U2034 ( .A1(n4920), .A2(n4921), .A3(n4922), .A4(n4923), .Y(n4919) );
  OA222X1_HVT U2035 ( .A1(n1117), .A2(n4543), .A3(n1245), .A4(n4544), .A5(
        n1373), .A6(n4545), .Y(n4923) );
  OA222X1_HVT U2036 ( .A1(n733), .A2(n4546), .A3(n861), .A4(n4547), .A5(n989), 
        .A6(n4548), .Y(n4922) );
  OA222X1_HVT U2037 ( .A1(n349), .A2(n4549), .A3(n477), .A4(n4550), .A5(n605), 
        .A6(n4551), .Y(n4921) );
  OA22X1_HVT U2038 ( .A1(n93), .A2(n4552), .A3(n221), .A4(n4553), .Y(n4920) );
  MUX21X1_HVT U2039 ( .A1(key_round[52]), .A2(n4924), .S0(n4512), .Y(n2177) );
  NAND4X0_HVT U2040 ( .A1(n4925), .A2(n4926), .A3(n4927), .A4(n4928), .Y(n4924) );
  OA222X1_HVT U2041 ( .A1(n1118), .A2(n4543), .A3(n1246), .A4(n4544), .A5(
        n1374), .A6(n4545), .Y(n4928) );
  OA222X1_HVT U2042 ( .A1(n734), .A2(n4546), .A3(n862), .A4(n4547), .A5(n990), 
        .A6(n4548), .Y(n4927) );
  OA222X1_HVT U2043 ( .A1(n350), .A2(n4549), .A3(n478), .A4(n4550), .A5(n606), 
        .A6(n4551), .Y(n4926) );
  OA22X1_HVT U2044 ( .A1(n94), .A2(n4552), .A3(n222), .A4(n4553), .Y(n4925) );
  MUX21X1_HVT U2045 ( .A1(key_round[51]), .A2(n4929), .S0(n4512), .Y(n2176) );
  NAND4X0_HVT U2046 ( .A1(n4930), .A2(n4931), .A3(n4932), .A4(n4933), .Y(n4929) );
  OA222X1_HVT U2047 ( .A1(n1119), .A2(n4543), .A3(n1247), .A4(n4544), .A5(
        n1375), .A6(n4545), .Y(n4933) );
  OA222X1_HVT U2048 ( .A1(n735), .A2(n4546), .A3(n863), .A4(n4547), .A5(n991), 
        .A6(n4548), .Y(n4932) );
  OA222X1_HVT U2049 ( .A1(n351), .A2(n4549), .A3(n479), .A4(n4550), .A5(n607), 
        .A6(n4551), .Y(n4931) );
  OA22X1_HVT U2050 ( .A1(n95), .A2(n4552), .A3(n223), .A4(n4553), .Y(n4930) );
  MUX21X1_HVT U2051 ( .A1(key_round[50]), .A2(n4934), .S0(n4512), .Y(n2175) );
  NAND4X0_HVT U2052 ( .A1(n4935), .A2(n4936), .A3(n4937), .A4(n4938), .Y(n4934) );
  OA222X1_HVT U2053 ( .A1(n1120), .A2(n4543), .A3(n1248), .A4(n4544), .A5(
        n1376), .A6(n4545), .Y(n4938) );
  OA222X1_HVT U2054 ( .A1(n736), .A2(n4546), .A3(n864), .A4(n4547), .A5(n992), 
        .A6(n4548), .Y(n4937) );
  OA222X1_HVT U2055 ( .A1(n352), .A2(n4549), .A3(n480), .A4(n4550), .A5(n608), 
        .A6(n4551), .Y(n4936) );
  OA22X1_HVT U2056 ( .A1(n96), .A2(n4552), .A3(n224), .A4(n4553), .Y(n4935) );
  MUX21X1_HVT U2057 ( .A1(key_round[49]), .A2(n4939), .S0(n4512), .Y(n2174) );
  NAND4X0_HVT U2058 ( .A1(n4940), .A2(n4941), .A3(n4942), .A4(n4943), .Y(n4939) );
  OA222X1_HVT U2059 ( .A1(n1121), .A2(n4543), .A3(n1249), .A4(n4544), .A5(
        n1377), .A6(n4545), .Y(n4943) );
  OA222X1_HVT U2060 ( .A1(n737), .A2(n4546), .A3(n865), .A4(n4547), .A5(n993), 
        .A6(n4548), .Y(n4942) );
  OA222X1_HVT U2061 ( .A1(n353), .A2(n4549), .A3(n481), .A4(n4550), .A5(n609), 
        .A6(n4551), .Y(n4941) );
  OA22X1_HVT U2062 ( .A1(n97), .A2(n4552), .A3(n225), .A4(n4553), .Y(n4940) );
  MUX21X1_HVT U2063 ( .A1(key_round[48]), .A2(n4944), .S0(n4512), .Y(n2173) );
  NAND4X0_HVT U2064 ( .A1(n4945), .A2(n4946), .A3(n4947), .A4(n4948), .Y(n4944) );
  OA222X1_HVT U2065 ( .A1(n1122), .A2(n4543), .A3(n1250), .A4(n4544), .A5(
        n1378), .A6(n4545), .Y(n4948) );
  OA222X1_HVT U2066 ( .A1(n738), .A2(n4546), .A3(n866), .A4(n4547), .A5(n994), 
        .A6(n4548), .Y(n4947) );
  OA222X1_HVT U2067 ( .A1(n354), .A2(n4549), .A3(n482), .A4(n4550), .A5(n610), 
        .A6(n4551), .Y(n4946) );
  OA22X1_HVT U2068 ( .A1(n98), .A2(n4552), .A3(n226), .A4(n4553), .Y(n4945) );
  MUX21X1_HVT U2069 ( .A1(key_round[47]), .A2(n4949), .S0(n4512), .Y(n2172) );
  NAND4X0_HVT U2070 ( .A1(n4950), .A2(n4951), .A3(n4952), .A4(n4953), .Y(n4949) );
  OA222X1_HVT U2071 ( .A1(n1123), .A2(n4543), .A3(n1251), .A4(n4544), .A5(
        n1379), .A6(n4545), .Y(n4953) );
  OA222X1_HVT U2072 ( .A1(n739), .A2(n4546), .A3(n867), .A4(n4547), .A5(n995), 
        .A6(n4548), .Y(n4952) );
  OA222X1_HVT U2073 ( .A1(n355), .A2(n4549), .A3(n483), .A4(n4550), .A5(n611), 
        .A6(n4551), .Y(n4951) );
  OA22X1_HVT U2074 ( .A1(n99), .A2(n4552), .A3(n227), .A4(n4553), .Y(n4950) );
  MUX21X1_HVT U2075 ( .A1(key_round[46]), .A2(n4954), .S0(n4512), .Y(n2171) );
  NAND4X0_HVT U2076 ( .A1(n4955), .A2(n4956), .A3(n4957), .A4(n4958), .Y(n4954) );
  OA222X1_HVT U2077 ( .A1(n1124), .A2(n4543), .A3(n1252), .A4(n4544), .A5(
        n1380), .A6(n4545), .Y(n4958) );
  OA222X1_HVT U2078 ( .A1(n740), .A2(n4546), .A3(n868), .A4(n4547), .A5(n996), 
        .A6(n4548), .Y(n4957) );
  OA222X1_HVT U2079 ( .A1(n356), .A2(n4549), .A3(n484), .A4(n4550), .A5(n612), 
        .A6(n4551), .Y(n4956) );
  OA22X1_HVT U2080 ( .A1(n100), .A2(n4552), .A3(n228), .A4(n4553), .Y(n4955)
         );
  MUX21X1_HVT U2081 ( .A1(key_round[45]), .A2(n4959), .S0(n4512), .Y(n2170) );
  NAND4X0_HVT U2082 ( .A1(n4960), .A2(n4961), .A3(n4962), .A4(n4963), .Y(n4959) );
  OA222X1_HVT U2083 ( .A1(n1125), .A2(n4543), .A3(n1253), .A4(n4544), .A5(
        n1381), .A6(n4545), .Y(n4963) );
  OA222X1_HVT U2084 ( .A1(n741), .A2(n4546), .A3(n869), .A4(n4547), .A5(n997), 
        .A6(n4548), .Y(n4962) );
  OA222X1_HVT U2085 ( .A1(n357), .A2(n4549), .A3(n485), .A4(n4550), .A5(n613), 
        .A6(n4551), .Y(n4961) );
  OA22X1_HVT U2086 ( .A1(n101), .A2(n4552), .A3(n229), .A4(n4553), .Y(n4960)
         );
  MUX21X1_HVT U2087 ( .A1(key_round[44]), .A2(n4964), .S0(n4512), .Y(n2169) );
  NAND4X0_HVT U2088 ( .A1(n4965), .A2(n4966), .A3(n4967), .A4(n4968), .Y(n4964) );
  OA222X1_HVT U2089 ( .A1(n1126), .A2(n4543), .A3(n1254), .A4(n4544), .A5(
        n1382), .A6(n4545), .Y(n4968) );
  OA222X1_HVT U2090 ( .A1(n742), .A2(n4546), .A3(n870), .A4(n4547), .A5(n998), 
        .A6(n4548), .Y(n4967) );
  OA222X1_HVT U2091 ( .A1(n358), .A2(n4549), .A3(n486), .A4(n4550), .A5(n614), 
        .A6(n4551), .Y(n4966) );
  OA22X1_HVT U2092 ( .A1(n102), .A2(n4552), .A3(n230), .A4(n4553), .Y(n4965)
         );
  MUX21X1_HVT U2093 ( .A1(key_round[43]), .A2(n4969), .S0(n4512), .Y(n2168) );
  NAND4X0_HVT U2094 ( .A1(n4970), .A2(n4971), .A3(n4972), .A4(n4973), .Y(n4969) );
  OA222X1_HVT U2095 ( .A1(n1127), .A2(n4543), .A3(n1255), .A4(n4544), .A5(
        n1383), .A6(n4545), .Y(n4973) );
  OA222X1_HVT U2096 ( .A1(n743), .A2(n4546), .A3(n871), .A4(n4547), .A5(n999), 
        .A6(n4548), .Y(n4972) );
  OA222X1_HVT U2097 ( .A1(n359), .A2(n4549), .A3(n487), .A4(n4550), .A5(n615), 
        .A6(n4551), .Y(n4971) );
  OA22X1_HVT U2098 ( .A1(n103), .A2(n4552), .A3(n231), .A4(n4553), .Y(n4970)
         );
  MUX21X1_HVT U2099 ( .A1(key_round[42]), .A2(n4974), .S0(n4512), .Y(n2167) );
  NAND4X0_HVT U2100 ( .A1(n4975), .A2(n4976), .A3(n4977), .A4(n4978), .Y(n4974) );
  OA222X1_HVT U2101 ( .A1(n1128), .A2(n4543), .A3(n1256), .A4(n4544), .A5(
        n1384), .A6(n4545), .Y(n4978) );
  OA222X1_HVT U2102 ( .A1(n744), .A2(n4546), .A3(n872), .A4(n4547), .A5(n1000), 
        .A6(n4548), .Y(n4977) );
  OA222X1_HVT U2103 ( .A1(n360), .A2(n4549), .A3(n488), .A4(n4550), .A5(n616), 
        .A6(n4551), .Y(n4976) );
  OA22X1_HVT U2104 ( .A1(n104), .A2(n4552), .A3(n232), .A4(n4553), .Y(n4975)
         );
  MUX21X1_HVT U2105 ( .A1(key_round[41]), .A2(n4979), .S0(n4512), .Y(n2166) );
  NAND4X0_HVT U2106 ( .A1(n4980), .A2(n4981), .A3(n4982), .A4(n4983), .Y(n4979) );
  OA222X1_HVT U2107 ( .A1(n1129), .A2(n4543), .A3(n1257), .A4(n4544), .A5(
        n1385), .A6(n4545), .Y(n4983) );
  OA222X1_HVT U2108 ( .A1(n745), .A2(n4546), .A3(n873), .A4(n4547), .A5(n1001), 
        .A6(n4548), .Y(n4982) );
  OA222X1_HVT U2109 ( .A1(n361), .A2(n4549), .A3(n489), .A4(n4550), .A5(n617), 
        .A6(n4551), .Y(n4981) );
  OA22X1_HVT U2110 ( .A1(n105), .A2(n4552), .A3(n233), .A4(n4553), .Y(n4980)
         );
  MUX21X1_HVT U2111 ( .A1(key_round[40]), .A2(n4984), .S0(n4512), .Y(n2165) );
  NAND4X0_HVT U2112 ( .A1(n4985), .A2(n4986), .A3(n4987), .A4(n4988), .Y(n4984) );
  OA222X1_HVT U2113 ( .A1(n1130), .A2(n4543), .A3(n1258), .A4(n4544), .A5(
        n1386), .A6(n4545), .Y(n4988) );
  OA222X1_HVT U2114 ( .A1(n746), .A2(n4546), .A3(n874), .A4(n4547), .A5(n1002), 
        .A6(n4548), .Y(n4987) );
  OA222X1_HVT U2115 ( .A1(n362), .A2(n4549), .A3(n490), .A4(n4550), .A5(n618), 
        .A6(n4551), .Y(n4986) );
  OA22X1_HVT U2116 ( .A1(n106), .A2(n4552), .A3(n234), .A4(n4553), .Y(n4985)
         );
  MUX21X1_HVT U2117 ( .A1(key_round[39]), .A2(n4989), .S0(n4512), .Y(n2164) );
  NAND4X0_HVT U2118 ( .A1(n4990), .A2(n4991), .A3(n4992), .A4(n4993), .Y(n4989) );
  OA222X1_HVT U2119 ( .A1(n1131), .A2(n4543), .A3(n1259), .A4(n4544), .A5(
        n1387), .A6(n4545), .Y(n4993) );
  OA222X1_HVT U2120 ( .A1(n747), .A2(n4546), .A3(n875), .A4(n4547), .A5(n1003), 
        .A6(n4548), .Y(n4992) );
  OA222X1_HVT U2121 ( .A1(n363), .A2(n4549), .A3(n491), .A4(n4550), .A5(n619), 
        .A6(n4551), .Y(n4991) );
  OA22X1_HVT U2122 ( .A1(n107), .A2(n4552), .A3(n235), .A4(n4553), .Y(n4990)
         );
  MUX21X1_HVT U2123 ( .A1(key_round[38]), .A2(n4994), .S0(n4512), .Y(n2163) );
  NAND4X0_HVT U2124 ( .A1(n4995), .A2(n4996), .A3(n4997), .A4(n4998), .Y(n4994) );
  OA222X1_HVT U2125 ( .A1(n1132), .A2(n4543), .A3(n1260), .A4(n4544), .A5(
        n1388), .A6(n4545), .Y(n4998) );
  OA222X1_HVT U2126 ( .A1(n748), .A2(n4546), .A3(n876), .A4(n4547), .A5(n1004), 
        .A6(n4548), .Y(n4997) );
  OA222X1_HVT U2127 ( .A1(n364), .A2(n4549), .A3(n492), .A4(n4550), .A5(n620), 
        .A6(n4551), .Y(n4996) );
  OA22X1_HVT U2128 ( .A1(n108), .A2(n4552), .A3(n236), .A4(n4553), .Y(n4995)
         );
  MUX21X1_HVT U2129 ( .A1(key_round[37]), .A2(n4999), .S0(n4512), .Y(n2162) );
  NAND4X0_HVT U2130 ( .A1(n5000), .A2(n5001), .A3(n5002), .A4(n5003), .Y(n4999) );
  OA222X1_HVT U2131 ( .A1(n1133), .A2(n4543), .A3(n1261), .A4(n4544), .A5(
        n1389), .A6(n4545), .Y(n5003) );
  OA222X1_HVT U2132 ( .A1(n749), .A2(n4546), .A3(n877), .A4(n4547), .A5(n1005), 
        .A6(n4548), .Y(n5002) );
  OA222X1_HVT U2133 ( .A1(n365), .A2(n4549), .A3(n493), .A4(n4550), .A5(n621), 
        .A6(n4551), .Y(n5001) );
  OA22X1_HVT U2134 ( .A1(n109), .A2(n4552), .A3(n237), .A4(n4553), .Y(n5000)
         );
  MUX21X1_HVT U2135 ( .A1(key_round[36]), .A2(n5004), .S0(n4512), .Y(n2161) );
  NAND4X0_HVT U2136 ( .A1(n5005), .A2(n5006), .A3(n5007), .A4(n5008), .Y(n5004) );
  OA222X1_HVT U2137 ( .A1(n1134), .A2(n4543), .A3(n1262), .A4(n4544), .A5(
        n1390), .A6(n4545), .Y(n5008) );
  OA222X1_HVT U2138 ( .A1(n750), .A2(n4546), .A3(n878), .A4(n4547), .A5(n1006), 
        .A6(n4548), .Y(n5007) );
  OA222X1_HVT U2139 ( .A1(n366), .A2(n4549), .A3(n494), .A4(n4550), .A5(n622), 
        .A6(n4551), .Y(n5006) );
  OA22X1_HVT U2140 ( .A1(n110), .A2(n4552), .A3(n238), .A4(n4553), .Y(n5005)
         );
  MUX21X1_HVT U2141 ( .A1(key_round[35]), .A2(n5009), .S0(n4512), .Y(n2160) );
  NAND4X0_HVT U2142 ( .A1(n5010), .A2(n5011), .A3(n5012), .A4(n5013), .Y(n5009) );
  OA222X1_HVT U2143 ( .A1(n1135), .A2(n4543), .A3(n1263), .A4(n4544), .A5(
        n1391), .A6(n4545), .Y(n5013) );
  OA222X1_HVT U2144 ( .A1(n751), .A2(n4546), .A3(n879), .A4(n4547), .A5(n1007), 
        .A6(n4548), .Y(n5012) );
  OA222X1_HVT U2145 ( .A1(n367), .A2(n4549), .A3(n495), .A4(n4550), .A5(n623), 
        .A6(n4551), .Y(n5011) );
  OA22X1_HVT U2146 ( .A1(n111), .A2(n4552), .A3(n239), .A4(n4553), .Y(n5010)
         );
  MUX21X1_HVT U2147 ( .A1(key_round[34]), .A2(n5014), .S0(n4512), .Y(n2159) );
  NAND4X0_HVT U2148 ( .A1(n5015), .A2(n5016), .A3(n5017), .A4(n5018), .Y(n5014) );
  OA222X1_HVT U2149 ( .A1(n1136), .A2(n4543), .A3(n1264), .A4(n4544), .A5(
        n1392), .A6(n4545), .Y(n5018) );
  OA222X1_HVT U2150 ( .A1(n752), .A2(n4546), .A3(n880), .A4(n4547), .A5(n1008), 
        .A6(n4548), .Y(n5017) );
  OA222X1_HVT U2151 ( .A1(n368), .A2(n4549), .A3(n496), .A4(n4550), .A5(n624), 
        .A6(n4551), .Y(n5016) );
  OA22X1_HVT U2152 ( .A1(n112), .A2(n4552), .A3(n240), .A4(n4553), .Y(n5015)
         );
  MUX21X1_HVT U2153 ( .A1(key_round[33]), .A2(n5019), .S0(n4512), .Y(n2158) );
  NAND4X0_HVT U2154 ( .A1(n5020), .A2(n5021), .A3(n5022), .A4(n5023), .Y(n5019) );
  OA222X1_HVT U2155 ( .A1(n1137), .A2(n4543), .A3(n1265), .A4(n4544), .A5(
        n1393), .A6(n4545), .Y(n5023) );
  OA222X1_HVT U2156 ( .A1(n753), .A2(n4546), .A3(n881), .A4(n4547), .A5(n1009), 
        .A6(n4548), .Y(n5022) );
  OA222X1_HVT U2157 ( .A1(n369), .A2(n4549), .A3(n497), .A4(n4550), .A5(n625), 
        .A6(n4551), .Y(n5021) );
  OA22X1_HVT U2158 ( .A1(n113), .A2(n4552), .A3(n241), .A4(n4553), .Y(n5020)
         );
  MUX21X1_HVT U2159 ( .A1(key_round[32]), .A2(n5024), .S0(n4512), .Y(n2157) );
  NAND4X0_HVT U2160 ( .A1(n5025), .A2(n5026), .A3(n5027), .A4(n5028), .Y(n5024) );
  OA222X1_HVT U2161 ( .A1(n1138), .A2(n4543), .A3(n1266), .A4(n4544), .A5(
        n1394), .A6(n4545), .Y(n5028) );
  OA222X1_HVT U2162 ( .A1(n754), .A2(n4546), .A3(n882), .A4(n4547), .A5(n1010), 
        .A6(n4548), .Y(n5027) );
  OA222X1_HVT U2163 ( .A1(n370), .A2(n4549), .A3(n498), .A4(n4550), .A5(n626), 
        .A6(n4551), .Y(n5026) );
  OA22X1_HVT U2164 ( .A1(n114), .A2(n4552), .A3(n242), .A4(n4553), .Y(n5025)
         );
  MUX21X1_HVT U2165 ( .A1(key_round[31]), .A2(n5029), .S0(n4512), .Y(n2156) );
  NAND4X0_HVT U2166 ( .A1(n5030), .A2(n5031), .A3(n5032), .A4(n5033), .Y(n5029) );
  OA222X1_HVT U2167 ( .A1(n1139), .A2(n4543), .A3(n1267), .A4(n4544), .A5(
        n1395), .A6(n4545), .Y(n5033) );
  OA222X1_HVT U2168 ( .A1(n755), .A2(n4546), .A3(n883), .A4(n4547), .A5(n1011), 
        .A6(n4548), .Y(n5032) );
  OA222X1_HVT U2169 ( .A1(n371), .A2(n4549), .A3(n499), .A4(n4550), .A5(n627), 
        .A6(n4551), .Y(n5031) );
  OA22X1_HVT U2170 ( .A1(n115), .A2(n4552), .A3(n243), .A4(n4553), .Y(n5030)
         );
  MUX21X1_HVT U2171 ( .A1(key_round[30]), .A2(n5034), .S0(n4512), .Y(n2155) );
  NAND4X0_HVT U2172 ( .A1(n5035), .A2(n5036), .A3(n5037), .A4(n5038), .Y(n5034) );
  OA222X1_HVT U2173 ( .A1(n1140), .A2(n4543), .A3(n1268), .A4(n4544), .A5(
        n1396), .A6(n4545), .Y(n5038) );
  OA222X1_HVT U2174 ( .A1(n756), .A2(n4546), .A3(n884), .A4(n4547), .A5(n1012), 
        .A6(n4548), .Y(n5037) );
  OA222X1_HVT U2175 ( .A1(n372), .A2(n4549), .A3(n500), .A4(n4550), .A5(n628), 
        .A6(n4551), .Y(n5036) );
  OA22X1_HVT U2176 ( .A1(n116), .A2(n4552), .A3(n244), .A4(n4553), .Y(n5035)
         );
  MUX21X1_HVT U2177 ( .A1(key_round[29]), .A2(n5039), .S0(n4512), .Y(n2154) );
  NAND4X0_HVT U2178 ( .A1(n5040), .A2(n5041), .A3(n5042), .A4(n5043), .Y(n5039) );
  OA222X1_HVT U2179 ( .A1(n1141), .A2(n4543), .A3(n1269), .A4(n4544), .A5(
        n1397), .A6(n4545), .Y(n5043) );
  OA222X1_HVT U2180 ( .A1(n757), .A2(n4546), .A3(n885), .A4(n4547), .A5(n1013), 
        .A6(n4548), .Y(n5042) );
  OA222X1_HVT U2181 ( .A1(n373), .A2(n4549), .A3(n501), .A4(n4550), .A5(n629), 
        .A6(n4551), .Y(n5041) );
  OA22X1_HVT U2182 ( .A1(n117), .A2(n4552), .A3(n245), .A4(n4553), .Y(n5040)
         );
  MUX21X1_HVT U2183 ( .A1(key_round[28]), .A2(n5044), .S0(n4512), .Y(n2153) );
  NAND4X0_HVT U2184 ( .A1(n5045), .A2(n5046), .A3(n5047), .A4(n5048), .Y(n5044) );
  OA222X1_HVT U2185 ( .A1(n1142), .A2(n4543), .A3(n1270), .A4(n4544), .A5(
        n1398), .A6(n4545), .Y(n5048) );
  OA222X1_HVT U2186 ( .A1(n758), .A2(n4546), .A3(n886), .A4(n4547), .A5(n1014), 
        .A6(n4548), .Y(n5047) );
  OA222X1_HVT U2187 ( .A1(n374), .A2(n4549), .A3(n502), .A4(n4550), .A5(n630), 
        .A6(n4551), .Y(n5046) );
  OA22X1_HVT U2188 ( .A1(n118), .A2(n4552), .A3(n246), .A4(n4553), .Y(n5045)
         );
  MUX21X1_HVT U2189 ( .A1(key_round[27]), .A2(n5049), .S0(n4512), .Y(n2152) );
  NAND4X0_HVT U2190 ( .A1(n5050), .A2(n5051), .A3(n5052), .A4(n5053), .Y(n5049) );
  OA222X1_HVT U2191 ( .A1(n1143), .A2(n4543), .A3(n1271), .A4(n4544), .A5(
        n1399), .A6(n4545), .Y(n5053) );
  OA222X1_HVT U2192 ( .A1(n759), .A2(n4546), .A3(n887), .A4(n4547), .A5(n1015), 
        .A6(n4548), .Y(n5052) );
  OA222X1_HVT U2193 ( .A1(n375), .A2(n4549), .A3(n503), .A4(n4550), .A5(n631), 
        .A6(n4551), .Y(n5051) );
  OA22X1_HVT U2194 ( .A1(n119), .A2(n4552), .A3(n247), .A4(n4553), .Y(n5050)
         );
  MUX21X1_HVT U2195 ( .A1(key_round[26]), .A2(n5054), .S0(n4512), .Y(n2151) );
  NAND4X0_HVT U2196 ( .A1(n5055), .A2(n5056), .A3(n5057), .A4(n5058), .Y(n5054) );
  OA222X1_HVT U2197 ( .A1(n1144), .A2(n4543), .A3(n1272), .A4(n4544), .A5(
        n1400), .A6(n4545), .Y(n5058) );
  OA222X1_HVT U2198 ( .A1(n760), .A2(n4546), .A3(n888), .A4(n4547), .A5(n1016), 
        .A6(n4548), .Y(n5057) );
  OA222X1_HVT U2199 ( .A1(n376), .A2(n4549), .A3(n504), .A4(n4550), .A5(n632), 
        .A6(n4551), .Y(n5056) );
  OA22X1_HVT U2200 ( .A1(n120), .A2(n4552), .A3(n248), .A4(n4553), .Y(n5055)
         );
  MUX21X1_HVT U2201 ( .A1(key_round[25]), .A2(n5059), .S0(n4512), .Y(n2150) );
  NAND4X0_HVT U2202 ( .A1(n5060), .A2(n5061), .A3(n5062), .A4(n5063), .Y(n5059) );
  OA222X1_HVT U2203 ( .A1(n1145), .A2(n4543), .A3(n1273), .A4(n4544), .A5(
        n1401), .A6(n4545), .Y(n5063) );
  OA222X1_HVT U2204 ( .A1(n761), .A2(n4546), .A3(n889), .A4(n4547), .A5(n1017), 
        .A6(n4548), .Y(n5062) );
  OA222X1_HVT U2205 ( .A1(n377), .A2(n4549), .A3(n505), .A4(n4550), .A5(n633), 
        .A6(n4551), .Y(n5061) );
  OA22X1_HVT U2206 ( .A1(n121), .A2(n4552), .A3(n249), .A4(n4553), .Y(n5060)
         );
  MUX21X1_HVT U2207 ( .A1(key_round[24]), .A2(n5064), .S0(n4512), .Y(n2149) );
  NAND4X0_HVT U2208 ( .A1(n5065), .A2(n5066), .A3(n5067), .A4(n5068), .Y(n5064) );
  OA222X1_HVT U2209 ( .A1(n1146), .A2(n4543), .A3(n1274), .A4(n4544), .A5(
        n1402), .A6(n4545), .Y(n5068) );
  OA222X1_HVT U2210 ( .A1(n762), .A2(n4546), .A3(n890), .A4(n4547), .A5(n1018), 
        .A6(n4548), .Y(n5067) );
  OA222X1_HVT U2211 ( .A1(n378), .A2(n4549), .A3(n506), .A4(n4550), .A5(n634), 
        .A6(n4551), .Y(n5066) );
  OA22X1_HVT U2212 ( .A1(n122), .A2(n4552), .A3(n250), .A4(n4553), .Y(n5065)
         );
  MUX21X1_HVT U2213 ( .A1(key_round[23]), .A2(n5069), .S0(n4512), .Y(n2148) );
  NAND4X0_HVT U2214 ( .A1(n5070), .A2(n5071), .A3(n5072), .A4(n5073), .Y(n5069) );
  OA222X1_HVT U2215 ( .A1(n1147), .A2(n4543), .A3(n1275), .A4(n4544), .A5(
        n1403), .A6(n4545), .Y(n5073) );
  OA222X1_HVT U2216 ( .A1(n763), .A2(n4546), .A3(n891), .A4(n4547), .A5(n1019), 
        .A6(n4548), .Y(n5072) );
  OA222X1_HVT U2217 ( .A1(n379), .A2(n4549), .A3(n507), .A4(n4550), .A5(n635), 
        .A6(n4551), .Y(n5071) );
  OA22X1_HVT U2218 ( .A1(n123), .A2(n4552), .A3(n251), .A4(n4553), .Y(n5070)
         );
  MUX21X1_HVT U2219 ( .A1(key_round[22]), .A2(n5074), .S0(n4512), .Y(n2147) );
  NAND4X0_HVT U2220 ( .A1(n5075), .A2(n5076), .A3(n5077), .A4(n5078), .Y(n5074) );
  OA222X1_HVT U2221 ( .A1(n1148), .A2(n4543), .A3(n1276), .A4(n4544), .A5(
        n1404), .A6(n4545), .Y(n5078) );
  OA222X1_HVT U2222 ( .A1(n764), .A2(n4546), .A3(n892), .A4(n4547), .A5(n1020), 
        .A6(n4548), .Y(n5077) );
  OA222X1_HVT U2223 ( .A1(n380), .A2(n4549), .A3(n508), .A4(n4550), .A5(n636), 
        .A6(n4551), .Y(n5076) );
  OA22X1_HVT U2224 ( .A1(n124), .A2(n4552), .A3(n252), .A4(n4553), .Y(n5075)
         );
  MUX21X1_HVT U2225 ( .A1(key_round[21]), .A2(n5079), .S0(n4512), .Y(n2146) );
  NAND4X0_HVT U2226 ( .A1(n5080), .A2(n5081), .A3(n5082), .A4(n5083), .Y(n5079) );
  OA222X1_HVT U2227 ( .A1(n1149), .A2(n4543), .A3(n1277), .A4(n4544), .A5(
        n1405), .A6(n4545), .Y(n5083) );
  OA222X1_HVT U2228 ( .A1(n765), .A2(n4546), .A3(n893), .A4(n4547), .A5(n1021), 
        .A6(n4548), .Y(n5082) );
  OA222X1_HVT U2229 ( .A1(n381), .A2(n4549), .A3(n509), .A4(n4550), .A5(n637), 
        .A6(n4551), .Y(n5081) );
  OA22X1_HVT U2230 ( .A1(n125), .A2(n4552), .A3(n253), .A4(n4553), .Y(n5080)
         );
  MUX21X1_HVT U2231 ( .A1(key_round[20]), .A2(n5084), .S0(n4512), .Y(n2145) );
  NAND4X0_HVT U2232 ( .A1(n5085), .A2(n5086), .A3(n5087), .A4(n5088), .Y(n5084) );
  OA222X1_HVT U2233 ( .A1(n1150), .A2(n4543), .A3(n1278), .A4(n4544), .A5(
        n1406), .A6(n4545), .Y(n5088) );
  OA222X1_HVT U2234 ( .A1(n766), .A2(n4546), .A3(n894), .A4(n4547), .A5(n1022), 
        .A6(n4548), .Y(n5087) );
  OA222X1_HVT U2235 ( .A1(n382), .A2(n4549), .A3(n510), .A4(n4550), .A5(n638), 
        .A6(n4551), .Y(n5086) );
  OA22X1_HVT U2236 ( .A1(n126), .A2(n4552), .A3(n254), .A4(n4553), .Y(n5085)
         );
  MUX21X1_HVT U2237 ( .A1(key_round[19]), .A2(n5089), .S0(n4512), .Y(n2144) );
  NAND4X0_HVT U2238 ( .A1(n5090), .A2(n5091), .A3(n5092), .A4(n5093), .Y(n5089) );
  OA222X1_HVT U2239 ( .A1(n1151), .A2(n4543), .A3(n1279), .A4(n4544), .A5(
        n1407), .A6(n4545), .Y(n5093) );
  OA222X1_HVT U2240 ( .A1(n767), .A2(n4546), .A3(n895), .A4(n4547), .A5(n1023), 
        .A6(n4548), .Y(n5092) );
  OA222X1_HVT U2241 ( .A1(n383), .A2(n4549), .A3(n511), .A4(n4550), .A5(n639), 
        .A6(n4551), .Y(n5091) );
  OA22X1_HVT U2242 ( .A1(n127), .A2(n4552), .A3(n255), .A4(n4553), .Y(n5090)
         );
  MUX21X1_HVT U2243 ( .A1(key_round[18]), .A2(n5094), .S0(n4512), .Y(n2143) );
  NAND4X0_HVT U2244 ( .A1(n5095), .A2(n5096), .A3(n5097), .A4(n5098), .Y(n5094) );
  OA222X1_HVT U2245 ( .A1(n1152), .A2(n4543), .A3(n1280), .A4(n4544), .A5(
        n1408), .A6(n4545), .Y(n5098) );
  OA222X1_HVT U2246 ( .A1(n768), .A2(n4546), .A3(n896), .A4(n4547), .A5(n1024), 
        .A6(n4548), .Y(n5097) );
  OA222X1_HVT U2247 ( .A1(n384), .A2(n4549), .A3(n512), .A4(n4550), .A5(n640), 
        .A6(n4551), .Y(n5096) );
  OA22X1_HVT U2248 ( .A1(n128), .A2(n4552), .A3(n256), .A4(n4553), .Y(n5095)
         );
  MUX21X1_HVT U2249 ( .A1(key_round[17]), .A2(n5099), .S0(n4512), .Y(n2142) );
  NAND4X0_HVT U2250 ( .A1(n5100), .A2(n5101), .A3(n5102), .A4(n5103), .Y(n5099) );
  OA222X1_HVT U2251 ( .A1(n1153), .A2(n4543), .A3(n1281), .A4(n4544), .A5(
        n1409), .A6(n4545), .Y(n5103) );
  OA222X1_HVT U2252 ( .A1(n769), .A2(n4546), .A3(n897), .A4(n4547), .A5(n1025), 
        .A6(n4548), .Y(n5102) );
  OA222X1_HVT U2253 ( .A1(n385), .A2(n4549), .A3(n513), .A4(n4550), .A5(n641), 
        .A6(n4551), .Y(n5101) );
  OA22X1_HVT U2254 ( .A1(n129), .A2(n4552), .A3(n257), .A4(n4553), .Y(n5100)
         );
  MUX21X1_HVT U2255 ( .A1(key_round[16]), .A2(n5104), .S0(n4512), .Y(n2141) );
  NAND4X0_HVT U2256 ( .A1(n5105), .A2(n5106), .A3(n5107), .A4(n5108), .Y(n5104) );
  OA222X1_HVT U2257 ( .A1(n1154), .A2(n4543), .A3(n1282), .A4(n4544), .A5(
        n1410), .A6(n4545), .Y(n5108) );
  OA222X1_HVT U2258 ( .A1(n770), .A2(n4546), .A3(n898), .A4(n4547), .A5(n1026), 
        .A6(n4548), .Y(n5107) );
  OA222X1_HVT U2259 ( .A1(n386), .A2(n4549), .A3(n514), .A4(n4550), .A5(n642), 
        .A6(n4551), .Y(n5106) );
  OA22X1_HVT U2260 ( .A1(n130), .A2(n4552), .A3(n258), .A4(n4553), .Y(n5105)
         );
  MUX21X1_HVT U2261 ( .A1(key_round[15]), .A2(n5109), .S0(n4512), .Y(n2140) );
  NAND4X0_HVT U2262 ( .A1(n5110), .A2(n5111), .A3(n5112), .A4(n5113), .Y(n5109) );
  OA222X1_HVT U2263 ( .A1(n1155), .A2(n4543), .A3(n1283), .A4(n4544), .A5(
        n1411), .A6(n4545), .Y(n5113) );
  OA222X1_HVT U2264 ( .A1(n771), .A2(n4546), .A3(n899), .A4(n4547), .A5(n1027), 
        .A6(n4548), .Y(n5112) );
  OA222X1_HVT U2265 ( .A1(n387), .A2(n4549), .A3(n515), .A4(n4550), .A5(n643), 
        .A6(n4551), .Y(n5111) );
  OA22X1_HVT U2266 ( .A1(n131), .A2(n4552), .A3(n259), .A4(n4553), .Y(n5110)
         );
  MUX21X1_HVT U2267 ( .A1(key_round[14]), .A2(n5114), .S0(n4512), .Y(n2139) );
  NAND4X0_HVT U2268 ( .A1(n5115), .A2(n5116), .A3(n5117), .A4(n5118), .Y(n5114) );
  OA222X1_HVT U2269 ( .A1(n1156), .A2(n4543), .A3(n1284), .A4(n4544), .A5(
        n1412), .A6(n4545), .Y(n5118) );
  OA222X1_HVT U2270 ( .A1(n772), .A2(n4546), .A3(n900), .A4(n4547), .A5(n1028), 
        .A6(n4548), .Y(n5117) );
  OA222X1_HVT U2271 ( .A1(n388), .A2(n4549), .A3(n516), .A4(n4550), .A5(n644), 
        .A6(n4551), .Y(n5116) );
  OA22X1_HVT U2272 ( .A1(n132), .A2(n4552), .A3(n260), .A4(n4553), .Y(n5115)
         );
  MUX21X1_HVT U2273 ( .A1(key_round[13]), .A2(n5119), .S0(n4512), .Y(n2138) );
  NAND4X0_HVT U2274 ( .A1(n5120), .A2(n5121), .A3(n5122), .A4(n5123), .Y(n5119) );
  OA222X1_HVT U2275 ( .A1(n1157), .A2(n4543), .A3(n1285), .A4(n4544), .A5(
        n1413), .A6(n4545), .Y(n5123) );
  OA222X1_HVT U2276 ( .A1(n773), .A2(n4546), .A3(n901), .A4(n4547), .A5(n1029), 
        .A6(n4548), .Y(n5122) );
  OA222X1_HVT U2277 ( .A1(n389), .A2(n4549), .A3(n517), .A4(n4550), .A5(n645), 
        .A6(n4551), .Y(n5121) );
  OA22X1_HVT U2278 ( .A1(n133), .A2(n4552), .A3(n261), .A4(n4553), .Y(n5120)
         );
  MUX21X1_HVT U2279 ( .A1(key_round[12]), .A2(n5124), .S0(n4512), .Y(n2137) );
  NAND4X0_HVT U2280 ( .A1(n5125), .A2(n5126), .A3(n5127), .A4(n5128), .Y(n5124) );
  OA222X1_HVT U2281 ( .A1(n1158), .A2(n4543), .A3(n1286), .A4(n4544), .A5(
        n1414), .A6(n4545), .Y(n5128) );
  OA222X1_HVT U2282 ( .A1(n774), .A2(n4546), .A3(n902), .A4(n4547), .A5(n1030), 
        .A6(n4548), .Y(n5127) );
  OA222X1_HVT U2283 ( .A1(n390), .A2(n4549), .A3(n518), .A4(n4550), .A5(n646), 
        .A6(n4551), .Y(n5126) );
  OA22X1_HVT U2284 ( .A1(n134), .A2(n4552), .A3(n262), .A4(n4553), .Y(n5125)
         );
  MUX21X1_HVT U2285 ( .A1(key_round[11]), .A2(n5129), .S0(n4512), .Y(n2136) );
  NAND4X0_HVT U2286 ( .A1(n5130), .A2(n5131), .A3(n5132), .A4(n5133), .Y(n5129) );
  OA222X1_HVT U2287 ( .A1(n1159), .A2(n4543), .A3(n1287), .A4(n4544), .A5(
        n1415), .A6(n4545), .Y(n5133) );
  OA222X1_HVT U2288 ( .A1(n775), .A2(n4546), .A3(n903), .A4(n4547), .A5(n1031), 
        .A6(n4548), .Y(n5132) );
  OA222X1_HVT U2289 ( .A1(n391), .A2(n4549), .A3(n519), .A4(n4550), .A5(n647), 
        .A6(n4551), .Y(n5131) );
  OA22X1_HVT U2290 ( .A1(n135), .A2(n4552), .A3(n263), .A4(n4553), .Y(n5130)
         );
  MUX21X1_HVT U2291 ( .A1(key_round[10]), .A2(n5134), .S0(n4512), .Y(n2135) );
  NAND4X0_HVT U2292 ( .A1(n5135), .A2(n5136), .A3(n5137), .A4(n5138), .Y(n5134) );
  OA222X1_HVT U2293 ( .A1(n1160), .A2(n4543), .A3(n1288), .A4(n4544), .A5(
        n1416), .A6(n4545), .Y(n5138) );
  OA222X1_HVT U2294 ( .A1(n776), .A2(n4546), .A3(n904), .A4(n4547), .A5(n1032), 
        .A6(n4548), .Y(n5137) );
  OA222X1_HVT U2295 ( .A1(n392), .A2(n4549), .A3(n520), .A4(n4550), .A5(n648), 
        .A6(n4551), .Y(n5136) );
  OA22X1_HVT U2296 ( .A1(n136), .A2(n4552), .A3(n264), .A4(n4553), .Y(n5135)
         );
  MUX21X1_HVT U2297 ( .A1(key_round[9]), .A2(n5139), .S0(n4512), .Y(n2134) );
  NAND4X0_HVT U2298 ( .A1(n5140), .A2(n5141), .A3(n5142), .A4(n5143), .Y(n5139) );
  OA222X1_HVT U2299 ( .A1(n1161), .A2(n4543), .A3(n1289), .A4(n4544), .A5(
        n1417), .A6(n4545), .Y(n5143) );
  OA222X1_HVT U2300 ( .A1(n777), .A2(n4546), .A3(n905), .A4(n4547), .A5(n1033), 
        .A6(n4548), .Y(n5142) );
  OA222X1_HVT U2301 ( .A1(n393), .A2(n4549), .A3(n521), .A4(n4550), .A5(n649), 
        .A6(n4551), .Y(n5141) );
  OA22X1_HVT U2302 ( .A1(n137), .A2(n4552), .A3(n265), .A4(n4553), .Y(n5140)
         );
  MUX21X1_HVT U2303 ( .A1(key_round[8]), .A2(n5144), .S0(n4512), .Y(n2133) );
  NAND4X0_HVT U2304 ( .A1(n5145), .A2(n5146), .A3(n5147), .A4(n5148), .Y(n5144) );
  OA222X1_HVT U2305 ( .A1(n1162), .A2(n4543), .A3(n1290), .A4(n4544), .A5(
        n1418), .A6(n4545), .Y(n5148) );
  OA222X1_HVT U2306 ( .A1(n778), .A2(n4546), .A3(n906), .A4(n4547), .A5(n1034), 
        .A6(n4548), .Y(n5147) );
  OA222X1_HVT U2307 ( .A1(n394), .A2(n4549), .A3(n522), .A4(n4550), .A5(n650), 
        .A6(n4551), .Y(n5146) );
  OA22X1_HVT U2308 ( .A1(n138), .A2(n4552), .A3(n266), .A4(n4553), .Y(n5145)
         );
  MUX21X1_HVT U2309 ( .A1(key_round[7]), .A2(n5149), .S0(n4512), .Y(n2132) );
  NAND4X0_HVT U2310 ( .A1(n5150), .A2(n5151), .A3(n5152), .A4(n5153), .Y(n5149) );
  OA222X1_HVT U2311 ( .A1(n1163), .A2(n4543), .A3(n1291), .A4(n4544), .A5(
        n1419), .A6(n4545), .Y(n5153) );
  OA222X1_HVT U2312 ( .A1(n779), .A2(n4546), .A3(n907), .A4(n4547), .A5(n1035), 
        .A6(n4548), .Y(n5152) );
  OA222X1_HVT U2313 ( .A1(n395), .A2(n4549), .A3(n523), .A4(n4550), .A5(n651), 
        .A6(n4551), .Y(n5151) );
  OA22X1_HVT U2314 ( .A1(n139), .A2(n4552), .A3(n267), .A4(n4553), .Y(n5150)
         );
  MUX21X1_HVT U2315 ( .A1(key_round[6]), .A2(n5154), .S0(n4512), .Y(n2131) );
  NAND4X0_HVT U2316 ( .A1(n5155), .A2(n5156), .A3(n5157), .A4(n5158), .Y(n5154) );
  OA222X1_HVT U2317 ( .A1(n1164), .A2(n4543), .A3(n1292), .A4(n4544), .A5(
        n1420), .A6(n4545), .Y(n5158) );
  OA222X1_HVT U2318 ( .A1(n780), .A2(n4546), .A3(n908), .A4(n4547), .A5(n1036), 
        .A6(n4548), .Y(n5157) );
  OA222X1_HVT U2319 ( .A1(n396), .A2(n4549), .A3(n524), .A4(n4550), .A5(n652), 
        .A6(n4551), .Y(n5156) );
  OA22X1_HVT U2320 ( .A1(n140), .A2(n4552), .A3(n268), .A4(n4553), .Y(n5155)
         );
  MUX21X1_HVT U2321 ( .A1(key_round[5]), .A2(n5159), .S0(n4512), .Y(n2130) );
  NAND4X0_HVT U2322 ( .A1(n5160), .A2(n5161), .A3(n5162), .A4(n5163), .Y(n5159) );
  OA222X1_HVT U2323 ( .A1(n1165), .A2(n4543), .A3(n1293), .A4(n4544), .A5(
        n1421), .A6(n4545), .Y(n5163) );
  OA222X1_HVT U2324 ( .A1(n781), .A2(n4546), .A3(n909), .A4(n4547), .A5(n1037), 
        .A6(n4548), .Y(n5162) );
  OA222X1_HVT U2325 ( .A1(n397), .A2(n4549), .A3(n525), .A4(n4550), .A5(n653), 
        .A6(n4551), .Y(n5161) );
  OA22X1_HVT U2326 ( .A1(n141), .A2(n4552), .A3(n269), .A4(n4553), .Y(n5160)
         );
  MUX21X1_HVT U2327 ( .A1(key_round[4]), .A2(n5164), .S0(n4512), .Y(n2129) );
  NAND4X0_HVT U2328 ( .A1(n5165), .A2(n5166), .A3(n5167), .A4(n5168), .Y(n5164) );
  OA222X1_HVT U2329 ( .A1(n1166), .A2(n4543), .A3(n1294), .A4(n4544), .A5(
        n1422), .A6(n4545), .Y(n5168) );
  OA222X1_HVT U2330 ( .A1(n782), .A2(n4546), .A3(n910), .A4(n4547), .A5(n1038), 
        .A6(n4548), .Y(n5167) );
  OA222X1_HVT U2331 ( .A1(n398), .A2(n4549), .A3(n526), .A4(n4550), .A5(n654), 
        .A6(n4551), .Y(n5166) );
  OA22X1_HVT U2332 ( .A1(n142), .A2(n4552), .A3(n270), .A4(n4553), .Y(n5165)
         );
  MUX21X1_HVT U2333 ( .A1(key_round[3]), .A2(n5169), .S0(n4512), .Y(n2128) );
  NAND4X0_HVT U2334 ( .A1(n5170), .A2(n5171), .A3(n5172), .A4(n5173), .Y(n5169) );
  OA222X1_HVT U2335 ( .A1(n1167), .A2(n4543), .A3(n1295), .A4(n4544), .A5(
        n1423), .A6(n4545), .Y(n5173) );
  OA222X1_HVT U2336 ( .A1(n783), .A2(n4546), .A3(n911), .A4(n4547), .A5(n1039), 
        .A6(n4548), .Y(n5172) );
  OA222X1_HVT U2337 ( .A1(n399), .A2(n4549), .A3(n527), .A4(n4550), .A5(n655), 
        .A6(n4551), .Y(n5171) );
  OA22X1_HVT U2338 ( .A1(n143), .A2(n4552), .A3(n271), .A4(n4553), .Y(n5170)
         );
  MUX21X1_HVT U2339 ( .A1(key_round[2]), .A2(n5174), .S0(n4512), .Y(n2127) );
  NAND4X0_HVT U2340 ( .A1(n5175), .A2(n5176), .A3(n5177), .A4(n5178), .Y(n5174) );
  OA222X1_HVT U2341 ( .A1(n1168), .A2(n4543), .A3(n1296), .A4(n4544), .A5(
        n1424), .A6(n4545), .Y(n5178) );
  OA222X1_HVT U2342 ( .A1(n784), .A2(n4546), .A3(n912), .A4(n4547), .A5(n1040), 
        .A6(n4548), .Y(n5177) );
  OA222X1_HVT U2343 ( .A1(n400), .A2(n4549), .A3(n528), .A4(n4550), .A5(n656), 
        .A6(n4551), .Y(n5176) );
  OA22X1_HVT U2344 ( .A1(n144), .A2(n4552), .A3(n272), .A4(n4553), .Y(n5175)
         );
  MUX21X1_HVT U2345 ( .A1(key_round[1]), .A2(n5179), .S0(n4512), .Y(n2126) );
  NAND4X0_HVT U2346 ( .A1(n5180), .A2(n5181), .A3(n5182), .A4(n5183), .Y(n5179) );
  OA222X1_HVT U2347 ( .A1(n1169), .A2(n4543), .A3(n1297), .A4(n4544), .A5(
        n1425), .A6(n4545), .Y(n5183) );
  OA222X1_HVT U2348 ( .A1(n785), .A2(n4546), .A3(n913), .A4(n4547), .A5(n1041), 
        .A6(n4548), .Y(n5182) );
  OA222X1_HVT U2349 ( .A1(n401), .A2(n4549), .A3(n529), .A4(n4550), .A5(n657), 
        .A6(n4551), .Y(n5181) );
  OA22X1_HVT U2350 ( .A1(n145), .A2(n4552), .A3(n273), .A4(n4553), .Y(n5180)
         );
  MUX21X1_HVT U2351 ( .A1(key_round[0]), .A2(n5184), .S0(n4512), .Y(n2125) );
  AND4X1_HVT U2352 ( .A1(state[0]), .A2(state[1]), .A3(n4537), .A4(n4511), .Y(
        n4512) );
  INVX0_HVT U2353 ( .A(rest), .Y(n4511) );
  AND2X1_HVT U2354 ( .A1(state[3]), .A2(n2), .Y(n4537) );
  NAND4X0_HVT U2355 ( .A1(n5185), .A2(n5186), .A3(n5187), .A4(n5188), .Y(n5184) );
  OA222X1_HVT U2356 ( .A1(n1170), .A2(n4543), .A3(n1298), .A4(n4544), .A5(
        n1426), .A6(n4545), .Y(n5188) );
  NAND2X0_HVT U2357 ( .A1(rount_no[1]), .A2(rount_no[3]), .Y(n4545) );
  NAND2X0_HVT U2358 ( .A1(rount_no[3]), .A2(rount_no[0]), .Y(n4544) );
  NAND2X0_HVT U2359 ( .A1(n5189), .A2(rount_no[3]), .Y(n4543) );
  OA222X1_HVT U2360 ( .A1(n786), .A2(n4546), .A3(n914), .A4(n4547), .A5(n1042), 
        .A6(n4548), .Y(n5187) );
  NAND3X0_HVT U2361 ( .A1(rount_no[1]), .A2(rount_no[0]), .A3(rount_no[2]), 
        .Y(n4548) );
  NAND3X0_HVT U2362 ( .A1(rount_no[1]), .A2(n5190), .A3(rount_no[2]), .Y(n4547) );
  NAND3X0_HVT U2363 ( .A1(rount_no[0]), .A2(n5191), .A3(rount_no[2]), .Y(n4546) );
  OA222X1_HVT U2364 ( .A1(n402), .A2(n4549), .A3(n530), .A4(n4550), .A5(n658), 
        .A6(n4551), .Y(n5186) );
  NAND2X0_HVT U2365 ( .A1(rount_no[2]), .A2(n5189), .Y(n4551) );
  OR3X1_HVT U2366 ( .A1(n5190), .A2(rount_no[2]), .A3(n5191), .Y(n4550) );
  NAND3X0_HVT U2367 ( .A1(rount_no[1]), .A2(n5190), .A3(n5192), .Y(n4549) );
  OA22X1_HVT U2368 ( .A1(n146), .A2(n4552), .A3(n274), .A4(n4553), .Y(n5185)
         );
  NAND3X0_HVT U2369 ( .A1(rount_no[0]), .A2(n5191), .A3(n5192), .Y(n4553) );
  NAND2X0_HVT U2370 ( .A1(n5192), .A2(n5189), .Y(n4552) );
  AND2X1_HVT U2371 ( .A1(n5191), .A2(n5190), .Y(n5189) );
  INVX0_HVT U2372 ( .A(rount_no[0]), .Y(n5190) );
  INVX0_HVT U2373 ( .A(rount_no[1]), .Y(n5191) );
  NOR2X0_HVT U2374 ( .A1(rount_no[3]), .A2(rount_no[2]), .Y(n5192) );
endmodule

