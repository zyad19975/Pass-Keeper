
module cde ( clk, rst, cam_start, pass, start_dec, start_enc, master_key, 
        account, data_flash, flash_pass_reg, flash_acc_reg, flash_or_acc_reg, 
        flash_or_acc_sel, pass_enc_reg, new_old_pass_sel, plain_reg, 
        local_master_reg, local_master_sel, out_reg, write_en, write_add, 
        boot_lood, match, dec_done, ready_encryption, write_data_flash, 
        add_flash, final_output );
  input [127:0] pass;
  input [127:0] master_key;
  input [127:0] account;
  input [255:0] data_flash;
  input [3:0] write_add;
  output [255:0] write_data_flash;
  output [3:0] add_flash;
  output [127:0] final_output;
  input clk, rst, cam_start, start_dec, start_enc, flash_pass_reg,
         flash_acc_reg, flash_or_acc_reg, flash_or_acc_sel, pass_enc_reg,
         new_old_pass_sel, plain_reg, local_master_reg, local_master_sel,
         out_reg, write_en, boot_lood;
  output match, dec_done, ready_encryption;

  wire   [127:0] out_flash_or_acc_sel;
  wire   [3:0] match_add;
  wire   [127:0] out_new_old_pass_sel;
  wire   [127:0] out_decry;
  wire   [127:0] out_local_master_sel;
  wire   [127:0] out_reg_flash_or_acc;
  wire   [127:0] out_encryption;
  wire   [127:0] out_reg_pass_enc;
  wire   [127:0] out_reg_plain_reg;
  wire   [127:0] out_local_master_reg;

  reg_D_0 reg_flash_or_acc ( .clk(clk), .rst(rst), .enable(flash_or_acc_reg), 
        .in(out_flash_or_acc_sel), .out(out_reg_flash_or_acc) );
  reg_D_6 reg_flash_account ( .clk(clk), .rst(rst), .enable(flash_acc_reg), 
        .in(out_reg_flash_or_acc), .out(write_data_flash[255:128]) );
  reg_D_5 reg_flash_pass ( .clk(clk), .rst(rst), .enable(flash_pass_reg), .in(
        out_encryption), .out(write_data_flash[127:0]) );
  reg_D_4 reg_pass_enc ( .clk(clk), .rst(rst), .enable(pass_enc_reg), .in(
        data_flash[127:0]), .out(out_reg_pass_enc) );
  reg_D_3 reg_plain_reg ( .clk(clk), .rst(rst), .enable(plain_reg), .in(
        out_new_old_pass_sel), .out(out_reg_plain_reg) );
  reg_D_2 reg_local_master ( .clk(clk), .rst(rst), .enable(local_master_reg), 
        .in(out_local_master_sel), .out(out_local_master_reg) );
  reg_D_1 reg_out_reg ( .clk(clk), .rst(rst), .enable(out_reg), .in(
        out_encryption), .out(final_output) );
  cam_DATA_WIDTH128_ADDR_WIDTH4 cam_inst ( .clk(clk), .rst(rst), .start(
        cam_start), .write_enable(write_en), .din(out_reg_flash_or_acc), 
        .write_addr(write_add), .match(match), .match_addr(match_add) );
  aes ENC ( .plaintext(out_reg_plain_reg), .key(out_local_master_reg), .clk(
        clk), .reset(rst), .start(start_enc), .cipher_text(out_encryption), 
        .ready(ready_encryption) );
  inv_aes DEC ( .clk(clk), .rest(rst), .start(start_dec), .plaintext1(
        out_reg_pass_enc), .local_key({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cipher_text(out_decry), .done(dec_done) );
  MUX21X1_HVT U2 ( .A1(pass[9]), .A2(out_decry[9]), .S0(new_old_pass_sel), .Y(
        out_new_old_pass_sel[9]) );
  MUX21X1_HVT U3 ( .A1(pass[99]), .A2(out_decry[99]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[99]) );
  MUX21X1_HVT U4 ( .A1(pass[98]), .A2(out_decry[98]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[98]) );
  MUX21X1_HVT U5 ( .A1(pass[97]), .A2(out_decry[97]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[97]) );
  MUX21X1_HVT U6 ( .A1(pass[96]), .A2(out_decry[96]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[96]) );
  MUX21X1_HVT U7 ( .A1(pass[95]), .A2(out_decry[95]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[95]) );
  MUX21X1_HVT U8 ( .A1(pass[94]), .A2(out_decry[94]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[94]) );
  MUX21X1_HVT U9 ( .A1(pass[93]), .A2(out_decry[93]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[93]) );
  MUX21X1_HVT U10 ( .A1(pass[92]), .A2(out_decry[92]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[92]) );
  MUX21X1_HVT U11 ( .A1(pass[91]), .A2(out_decry[91]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[91]) );
  MUX21X1_HVT U12 ( .A1(pass[90]), .A2(out_decry[90]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[90]) );
  MUX21X1_HVT U13 ( .A1(pass[8]), .A2(out_decry[8]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[8]) );
  MUX21X1_HVT U14 ( .A1(pass[89]), .A2(out_decry[89]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[89]) );
  MUX21X1_HVT U15 ( .A1(pass[88]), .A2(out_decry[88]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[88]) );
  MUX21X1_HVT U16 ( .A1(pass[87]), .A2(out_decry[87]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[87]) );
  MUX21X1_HVT U17 ( .A1(pass[86]), .A2(out_decry[86]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[86]) );
  MUX21X1_HVT U18 ( .A1(pass[85]), .A2(out_decry[85]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[85]) );
  MUX21X1_HVT U19 ( .A1(pass[84]), .A2(out_decry[84]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[84]) );
  MUX21X1_HVT U20 ( .A1(pass[83]), .A2(out_decry[83]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[83]) );
  MUX21X1_HVT U21 ( .A1(pass[82]), .A2(out_decry[82]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[82]) );
  MUX21X1_HVT U22 ( .A1(pass[81]), .A2(out_decry[81]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[81]) );
  MUX21X1_HVT U23 ( .A1(pass[80]), .A2(out_decry[80]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[80]) );
  MUX21X1_HVT U24 ( .A1(pass[7]), .A2(out_decry[7]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[7]) );
  MUX21X1_HVT U25 ( .A1(pass[79]), .A2(out_decry[79]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[79]) );
  MUX21X1_HVT U26 ( .A1(pass[78]), .A2(out_decry[78]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[78]) );
  MUX21X1_HVT U27 ( .A1(pass[77]), .A2(out_decry[77]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[77]) );
  MUX21X1_HVT U28 ( .A1(pass[76]), .A2(out_decry[76]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[76]) );
  MUX21X1_HVT U29 ( .A1(pass[75]), .A2(out_decry[75]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[75]) );
  MUX21X1_HVT U30 ( .A1(pass[74]), .A2(out_decry[74]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[74]) );
  MUX21X1_HVT U31 ( .A1(pass[73]), .A2(out_decry[73]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[73]) );
  MUX21X1_HVT U32 ( .A1(pass[72]), .A2(out_decry[72]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[72]) );
  MUX21X1_HVT U33 ( .A1(pass[71]), .A2(out_decry[71]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[71]) );
  MUX21X1_HVT U34 ( .A1(pass[70]), .A2(out_decry[70]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[70]) );
  MUX21X1_HVT U35 ( .A1(pass[6]), .A2(out_decry[6]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[6]) );
  MUX21X1_HVT U36 ( .A1(pass[69]), .A2(out_decry[69]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[69]) );
  MUX21X1_HVT U37 ( .A1(pass[68]), .A2(out_decry[68]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[68]) );
  MUX21X1_HVT U38 ( .A1(pass[67]), .A2(out_decry[67]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[67]) );
  MUX21X1_HVT U39 ( .A1(pass[66]), .A2(out_decry[66]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[66]) );
  MUX21X1_HVT U40 ( .A1(pass[65]), .A2(out_decry[65]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[65]) );
  MUX21X1_HVT U41 ( .A1(pass[64]), .A2(out_decry[64]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[64]) );
  MUX21X1_HVT U42 ( .A1(pass[63]), .A2(out_decry[63]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[63]) );
  MUX21X1_HVT U43 ( .A1(pass[62]), .A2(out_decry[62]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[62]) );
  MUX21X1_HVT U44 ( .A1(pass[61]), .A2(out_decry[61]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[61]) );
  MUX21X1_HVT U45 ( .A1(pass[60]), .A2(out_decry[60]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[60]) );
  MUX21X1_HVT U46 ( .A1(pass[5]), .A2(out_decry[5]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[5]) );
  MUX21X1_HVT U47 ( .A1(pass[59]), .A2(out_decry[59]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[59]) );
  MUX21X1_HVT U48 ( .A1(pass[58]), .A2(out_decry[58]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[58]) );
  MUX21X1_HVT U49 ( .A1(pass[57]), .A2(out_decry[57]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[57]) );
  MUX21X1_HVT U50 ( .A1(pass[56]), .A2(out_decry[56]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[56]) );
  MUX21X1_HVT U51 ( .A1(pass[55]), .A2(out_decry[55]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[55]) );
  MUX21X1_HVT U52 ( .A1(pass[54]), .A2(out_decry[54]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[54]) );
  MUX21X1_HVT U53 ( .A1(pass[53]), .A2(out_decry[53]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[53]) );
  MUX21X1_HVT U54 ( .A1(pass[52]), .A2(out_decry[52]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[52]) );
  MUX21X1_HVT U55 ( .A1(pass[51]), .A2(out_decry[51]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[51]) );
  MUX21X1_HVT U56 ( .A1(pass[50]), .A2(out_decry[50]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[50]) );
  MUX21X1_HVT U57 ( .A1(pass[4]), .A2(out_decry[4]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[4]) );
  MUX21X1_HVT U58 ( .A1(pass[49]), .A2(out_decry[49]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[49]) );
  MUX21X1_HVT U59 ( .A1(pass[48]), .A2(out_decry[48]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[48]) );
  MUX21X1_HVT U60 ( .A1(pass[47]), .A2(out_decry[47]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[47]) );
  MUX21X1_HVT U61 ( .A1(pass[46]), .A2(out_decry[46]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[46]) );
  MUX21X1_HVT U62 ( .A1(pass[45]), .A2(out_decry[45]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[45]) );
  MUX21X1_HVT U63 ( .A1(pass[44]), .A2(out_decry[44]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[44]) );
  MUX21X1_HVT U64 ( .A1(pass[43]), .A2(out_decry[43]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[43]) );
  MUX21X1_HVT U65 ( .A1(pass[42]), .A2(out_decry[42]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[42]) );
  MUX21X1_HVT U66 ( .A1(pass[41]), .A2(out_decry[41]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[41]) );
  MUX21X1_HVT U67 ( .A1(pass[40]), .A2(out_decry[40]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[40]) );
  MUX21X1_HVT U68 ( .A1(pass[3]), .A2(out_decry[3]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[3]) );
  MUX21X1_HVT U69 ( .A1(pass[39]), .A2(out_decry[39]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[39]) );
  MUX21X1_HVT U70 ( .A1(pass[38]), .A2(out_decry[38]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[38]) );
  MUX21X1_HVT U71 ( .A1(pass[37]), .A2(out_decry[37]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[37]) );
  MUX21X1_HVT U72 ( .A1(pass[36]), .A2(out_decry[36]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[36]) );
  MUX21X1_HVT U73 ( .A1(pass[35]), .A2(out_decry[35]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[35]) );
  MUX21X1_HVT U74 ( .A1(pass[34]), .A2(out_decry[34]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[34]) );
  MUX21X1_HVT U75 ( .A1(pass[33]), .A2(out_decry[33]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[33]) );
  MUX21X1_HVT U76 ( .A1(pass[32]), .A2(out_decry[32]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[32]) );
  MUX21X1_HVT U77 ( .A1(pass[31]), .A2(out_decry[31]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[31]) );
  MUX21X1_HVT U78 ( .A1(pass[30]), .A2(out_decry[30]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[30]) );
  MUX21X1_HVT U79 ( .A1(pass[2]), .A2(out_decry[2]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[2]) );
  MUX21X1_HVT U80 ( .A1(pass[29]), .A2(out_decry[29]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[29]) );
  MUX21X1_HVT U81 ( .A1(pass[28]), .A2(out_decry[28]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[28]) );
  MUX21X1_HVT U82 ( .A1(pass[27]), .A2(out_decry[27]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[27]) );
  MUX21X1_HVT U83 ( .A1(pass[26]), .A2(out_decry[26]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[26]) );
  MUX21X1_HVT U84 ( .A1(pass[25]), .A2(out_decry[25]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[25]) );
  MUX21X1_HVT U85 ( .A1(pass[24]), .A2(out_decry[24]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[24]) );
  MUX21X1_HVT U86 ( .A1(pass[23]), .A2(out_decry[23]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[23]) );
  MUX21X1_HVT U87 ( .A1(pass[22]), .A2(out_decry[22]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[22]) );
  MUX21X1_HVT U88 ( .A1(pass[21]), .A2(out_decry[21]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[21]) );
  MUX21X1_HVT U89 ( .A1(pass[20]), .A2(out_decry[20]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[20]) );
  MUX21X1_HVT U90 ( .A1(pass[1]), .A2(out_decry[1]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[1]) );
  MUX21X1_HVT U91 ( .A1(pass[19]), .A2(out_decry[19]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[19]) );
  MUX21X1_HVT U92 ( .A1(pass[18]), .A2(out_decry[18]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[18]) );
  MUX21X1_HVT U93 ( .A1(pass[17]), .A2(out_decry[17]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[17]) );
  MUX21X1_HVT U94 ( .A1(pass[16]), .A2(out_decry[16]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[16]) );
  MUX21X1_HVT U95 ( .A1(pass[15]), .A2(out_decry[15]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[15]) );
  MUX21X1_HVT U96 ( .A1(pass[14]), .A2(out_decry[14]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[14]) );
  MUX21X1_HVT U97 ( .A1(pass[13]), .A2(out_decry[13]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[13]) );
  MUX21X1_HVT U98 ( .A1(pass[12]), .A2(out_decry[12]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[12]) );
  MUX21X1_HVT U99 ( .A1(pass[127]), .A2(out_decry[127]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[127]) );
  MUX21X1_HVT U100 ( .A1(pass[126]), .A2(out_decry[126]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[126]) );
  MUX21X1_HVT U101 ( .A1(pass[125]), .A2(out_decry[125]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[125]) );
  MUX21X1_HVT U102 ( .A1(pass[124]), .A2(out_decry[124]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[124]) );
  MUX21X1_HVT U103 ( .A1(pass[123]), .A2(out_decry[123]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[123]) );
  MUX21X1_HVT U104 ( .A1(pass[122]), .A2(out_decry[122]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[122]) );
  MUX21X1_HVT U105 ( .A1(pass[121]), .A2(out_decry[121]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[121]) );
  MUX21X1_HVT U106 ( .A1(pass[120]), .A2(out_decry[120]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[120]) );
  MUX21X1_HVT U107 ( .A1(pass[11]), .A2(out_decry[11]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[11]) );
  MUX21X1_HVT U108 ( .A1(pass[119]), .A2(out_decry[119]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[119]) );
  MUX21X1_HVT U109 ( .A1(pass[118]), .A2(out_decry[118]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[118]) );
  MUX21X1_HVT U110 ( .A1(pass[117]), .A2(out_decry[117]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[117]) );
  MUX21X1_HVT U111 ( .A1(pass[116]), .A2(out_decry[116]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[116]) );
  MUX21X1_HVT U112 ( .A1(pass[115]), .A2(out_decry[115]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[115]) );
  MUX21X1_HVT U113 ( .A1(pass[114]), .A2(out_decry[114]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[114]) );
  MUX21X1_HVT U114 ( .A1(pass[113]), .A2(out_decry[113]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[113]) );
  MUX21X1_HVT U115 ( .A1(pass[112]), .A2(out_decry[112]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[112]) );
  MUX21X1_HVT U116 ( .A1(pass[111]), .A2(out_decry[111]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[111]) );
  MUX21X1_HVT U117 ( .A1(pass[110]), .A2(out_decry[110]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[110]) );
  MUX21X1_HVT U118 ( .A1(pass[10]), .A2(out_decry[10]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[10]) );
  MUX21X1_HVT U119 ( .A1(pass[109]), .A2(out_decry[109]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[109]) );
  MUX21X1_HVT U120 ( .A1(pass[108]), .A2(out_decry[108]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[108]) );
  MUX21X1_HVT U121 ( .A1(pass[107]), .A2(out_decry[107]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[107]) );
  MUX21X1_HVT U122 ( .A1(pass[106]), .A2(out_decry[106]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[106]) );
  MUX21X1_HVT U123 ( .A1(pass[105]), .A2(out_decry[105]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[105]) );
  MUX21X1_HVT U124 ( .A1(pass[104]), .A2(out_decry[104]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[104]) );
  MUX21X1_HVT U125 ( .A1(pass[103]), .A2(out_decry[103]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[103]) );
  MUX21X1_HVT U126 ( .A1(pass[102]), .A2(out_decry[102]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[102]) );
  MUX21X1_HVT U127 ( .A1(pass[101]), .A2(out_decry[101]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[101]) );
  MUX21X1_HVT U128 ( .A1(pass[100]), .A2(out_decry[100]), .S0(new_old_pass_sel), .Y(out_new_old_pass_sel[100]) );
  MUX21X1_HVT U129 ( .A1(pass[0]), .A2(out_decry[0]), .S0(new_old_pass_sel), 
        .Y(out_new_old_pass_sel[0]) );
  AND2X1_HVT U130 ( .A1(master_key[9]), .A2(local_master_sel), .Y(
        out_local_master_sel[9]) );
  AND2X1_HVT U131 ( .A1(master_key[99]), .A2(local_master_sel), .Y(
        out_local_master_sel[99]) );
  AND2X1_HVT U132 ( .A1(master_key[98]), .A2(local_master_sel), .Y(
        out_local_master_sel[98]) );
  AND2X1_HVT U133 ( .A1(master_key[97]), .A2(local_master_sel), .Y(
        out_local_master_sel[97]) );
  AND2X1_HVT U134 ( .A1(master_key[96]), .A2(local_master_sel), .Y(
        out_local_master_sel[96]) );
  AND2X1_HVT U135 ( .A1(master_key[95]), .A2(local_master_sel), .Y(
        out_local_master_sel[95]) );
  AND2X1_HVT U136 ( .A1(master_key[94]), .A2(local_master_sel), .Y(
        out_local_master_sel[94]) );
  AND2X1_HVT U137 ( .A1(master_key[93]), .A2(local_master_sel), .Y(
        out_local_master_sel[93]) );
  AND2X1_HVT U138 ( .A1(master_key[92]), .A2(local_master_sel), .Y(
        out_local_master_sel[92]) );
  AND2X1_HVT U139 ( .A1(master_key[91]), .A2(local_master_sel), .Y(
        out_local_master_sel[91]) );
  AND2X1_HVT U140 ( .A1(master_key[90]), .A2(local_master_sel), .Y(
        out_local_master_sel[90]) );
  AND2X1_HVT U141 ( .A1(master_key[8]), .A2(local_master_sel), .Y(
        out_local_master_sel[8]) );
  AND2X1_HVT U142 ( .A1(master_key[89]), .A2(local_master_sel), .Y(
        out_local_master_sel[89]) );
  AND2X1_HVT U143 ( .A1(master_key[88]), .A2(local_master_sel), .Y(
        out_local_master_sel[88]) );
  AND2X1_HVT U144 ( .A1(master_key[87]), .A2(local_master_sel), .Y(
        out_local_master_sel[87]) );
  AND2X1_HVT U145 ( .A1(master_key[86]), .A2(local_master_sel), .Y(
        out_local_master_sel[86]) );
  AND2X1_HVT U146 ( .A1(master_key[85]), .A2(local_master_sel), .Y(
        out_local_master_sel[85]) );
  AND2X1_HVT U147 ( .A1(master_key[84]), .A2(local_master_sel), .Y(
        out_local_master_sel[84]) );
  AND2X1_HVT U148 ( .A1(master_key[83]), .A2(local_master_sel), .Y(
        out_local_master_sel[83]) );
  AND2X1_HVT U149 ( .A1(master_key[82]), .A2(local_master_sel), .Y(
        out_local_master_sel[82]) );
  AND2X1_HVT U150 ( .A1(master_key[81]), .A2(local_master_sel), .Y(
        out_local_master_sel[81]) );
  AND2X1_HVT U151 ( .A1(master_key[80]), .A2(local_master_sel), .Y(
        out_local_master_sel[80]) );
  AND2X1_HVT U152 ( .A1(master_key[7]), .A2(local_master_sel), .Y(
        out_local_master_sel[7]) );
  AND2X1_HVT U153 ( .A1(master_key[79]), .A2(local_master_sel), .Y(
        out_local_master_sel[79]) );
  AND2X1_HVT U154 ( .A1(master_key[78]), .A2(local_master_sel), .Y(
        out_local_master_sel[78]) );
  AND2X1_HVT U155 ( .A1(master_key[77]), .A2(local_master_sel), .Y(
        out_local_master_sel[77]) );
  AND2X1_HVT U156 ( .A1(master_key[76]), .A2(local_master_sel), .Y(
        out_local_master_sel[76]) );
  AND2X1_HVT U157 ( .A1(master_key[75]), .A2(local_master_sel), .Y(
        out_local_master_sel[75]) );
  AND2X1_HVT U158 ( .A1(master_key[74]), .A2(local_master_sel), .Y(
        out_local_master_sel[74]) );
  AND2X1_HVT U159 ( .A1(master_key[73]), .A2(local_master_sel), .Y(
        out_local_master_sel[73]) );
  AND2X1_HVT U160 ( .A1(master_key[72]), .A2(local_master_sel), .Y(
        out_local_master_sel[72]) );
  AND2X1_HVT U161 ( .A1(master_key[71]), .A2(local_master_sel), .Y(
        out_local_master_sel[71]) );
  AND2X1_HVT U162 ( .A1(master_key[70]), .A2(local_master_sel), .Y(
        out_local_master_sel[70]) );
  AND2X1_HVT U163 ( .A1(master_key[6]), .A2(local_master_sel), .Y(
        out_local_master_sel[6]) );
  AND2X1_HVT U164 ( .A1(master_key[69]), .A2(local_master_sel), .Y(
        out_local_master_sel[69]) );
  AND2X1_HVT U165 ( .A1(master_key[68]), .A2(local_master_sel), .Y(
        out_local_master_sel[68]) );
  AND2X1_HVT U166 ( .A1(master_key[67]), .A2(local_master_sel), .Y(
        out_local_master_sel[67]) );
  AND2X1_HVT U167 ( .A1(master_key[66]), .A2(local_master_sel), .Y(
        out_local_master_sel[66]) );
  AND2X1_HVT U168 ( .A1(master_key[65]), .A2(local_master_sel), .Y(
        out_local_master_sel[65]) );
  AND2X1_HVT U169 ( .A1(master_key[64]), .A2(local_master_sel), .Y(
        out_local_master_sel[64]) );
  AND2X1_HVT U170 ( .A1(master_key[63]), .A2(local_master_sel), .Y(
        out_local_master_sel[63]) );
  AND2X1_HVT U171 ( .A1(master_key[62]), .A2(local_master_sel), .Y(
        out_local_master_sel[62]) );
  AND2X1_HVT U172 ( .A1(master_key[61]), .A2(local_master_sel), .Y(
        out_local_master_sel[61]) );
  AND2X1_HVT U173 ( .A1(master_key[60]), .A2(local_master_sel), .Y(
        out_local_master_sel[60]) );
  AND2X1_HVT U174 ( .A1(master_key[5]), .A2(local_master_sel), .Y(
        out_local_master_sel[5]) );
  AND2X1_HVT U175 ( .A1(master_key[59]), .A2(local_master_sel), .Y(
        out_local_master_sel[59]) );
  AND2X1_HVT U176 ( .A1(master_key[58]), .A2(local_master_sel), .Y(
        out_local_master_sel[58]) );
  AND2X1_HVT U177 ( .A1(master_key[57]), .A2(local_master_sel), .Y(
        out_local_master_sel[57]) );
  AND2X1_HVT U178 ( .A1(master_key[56]), .A2(local_master_sel), .Y(
        out_local_master_sel[56]) );
  AND2X1_HVT U179 ( .A1(master_key[55]), .A2(local_master_sel), .Y(
        out_local_master_sel[55]) );
  AND2X1_HVT U180 ( .A1(master_key[54]), .A2(local_master_sel), .Y(
        out_local_master_sel[54]) );
  AND2X1_HVT U181 ( .A1(master_key[53]), .A2(local_master_sel), .Y(
        out_local_master_sel[53]) );
  AND2X1_HVT U182 ( .A1(master_key[52]), .A2(local_master_sel), .Y(
        out_local_master_sel[52]) );
  AND2X1_HVT U183 ( .A1(master_key[51]), .A2(local_master_sel), .Y(
        out_local_master_sel[51]) );
  AND2X1_HVT U184 ( .A1(master_key[50]), .A2(local_master_sel), .Y(
        out_local_master_sel[50]) );
  AND2X1_HVT U185 ( .A1(master_key[4]), .A2(local_master_sel), .Y(
        out_local_master_sel[4]) );
  AND2X1_HVT U186 ( .A1(master_key[49]), .A2(local_master_sel), .Y(
        out_local_master_sel[49]) );
  AND2X1_HVT U187 ( .A1(master_key[48]), .A2(local_master_sel), .Y(
        out_local_master_sel[48]) );
  AND2X1_HVT U188 ( .A1(master_key[47]), .A2(local_master_sel), .Y(
        out_local_master_sel[47]) );
  AND2X1_HVT U189 ( .A1(master_key[46]), .A2(local_master_sel), .Y(
        out_local_master_sel[46]) );
  AND2X1_HVT U190 ( .A1(master_key[45]), .A2(local_master_sel), .Y(
        out_local_master_sel[45]) );
  AND2X1_HVT U191 ( .A1(master_key[44]), .A2(local_master_sel), .Y(
        out_local_master_sel[44]) );
  AND2X1_HVT U192 ( .A1(master_key[43]), .A2(local_master_sel), .Y(
        out_local_master_sel[43]) );
  AND2X1_HVT U193 ( .A1(master_key[42]), .A2(local_master_sel), .Y(
        out_local_master_sel[42]) );
  AND2X1_HVT U194 ( .A1(master_key[41]), .A2(local_master_sel), .Y(
        out_local_master_sel[41]) );
  AND2X1_HVT U195 ( .A1(master_key[40]), .A2(local_master_sel), .Y(
        out_local_master_sel[40]) );
  AND2X1_HVT U196 ( .A1(master_key[3]), .A2(local_master_sel), .Y(
        out_local_master_sel[3]) );
  AND2X1_HVT U197 ( .A1(master_key[39]), .A2(local_master_sel), .Y(
        out_local_master_sel[39]) );
  AND2X1_HVT U198 ( .A1(master_key[38]), .A2(local_master_sel), .Y(
        out_local_master_sel[38]) );
  AND2X1_HVT U199 ( .A1(master_key[37]), .A2(local_master_sel), .Y(
        out_local_master_sel[37]) );
  AND2X1_HVT U200 ( .A1(master_key[36]), .A2(local_master_sel), .Y(
        out_local_master_sel[36]) );
  AND2X1_HVT U201 ( .A1(master_key[35]), .A2(local_master_sel), .Y(
        out_local_master_sel[35]) );
  AND2X1_HVT U202 ( .A1(master_key[34]), .A2(local_master_sel), .Y(
        out_local_master_sel[34]) );
  AND2X1_HVT U203 ( .A1(master_key[33]), .A2(local_master_sel), .Y(
        out_local_master_sel[33]) );
  AND2X1_HVT U204 ( .A1(master_key[32]), .A2(local_master_sel), .Y(
        out_local_master_sel[32]) );
  AND2X1_HVT U205 ( .A1(master_key[31]), .A2(local_master_sel), .Y(
        out_local_master_sel[31]) );
  AND2X1_HVT U206 ( .A1(master_key[30]), .A2(local_master_sel), .Y(
        out_local_master_sel[30]) );
  AND2X1_HVT U207 ( .A1(master_key[2]), .A2(local_master_sel), .Y(
        out_local_master_sel[2]) );
  AND2X1_HVT U208 ( .A1(master_key[29]), .A2(local_master_sel), .Y(
        out_local_master_sel[29]) );
  AND2X1_HVT U209 ( .A1(master_key[28]), .A2(local_master_sel), .Y(
        out_local_master_sel[28]) );
  AND2X1_HVT U210 ( .A1(master_key[27]), .A2(local_master_sel), .Y(
        out_local_master_sel[27]) );
  AND2X1_HVT U211 ( .A1(master_key[26]), .A2(local_master_sel), .Y(
        out_local_master_sel[26]) );
  AND2X1_HVT U212 ( .A1(master_key[25]), .A2(local_master_sel), .Y(
        out_local_master_sel[25]) );
  AND2X1_HVT U213 ( .A1(master_key[24]), .A2(local_master_sel), .Y(
        out_local_master_sel[24]) );
  AND2X1_HVT U214 ( .A1(master_key[23]), .A2(local_master_sel), .Y(
        out_local_master_sel[23]) );
  AND2X1_HVT U215 ( .A1(master_key[22]), .A2(local_master_sel), .Y(
        out_local_master_sel[22]) );
  AND2X1_HVT U216 ( .A1(master_key[21]), .A2(local_master_sel), .Y(
        out_local_master_sel[21]) );
  AND2X1_HVT U217 ( .A1(master_key[20]), .A2(local_master_sel), .Y(
        out_local_master_sel[20]) );
  AND2X1_HVT U218 ( .A1(master_key[1]), .A2(local_master_sel), .Y(
        out_local_master_sel[1]) );
  AND2X1_HVT U219 ( .A1(master_key[19]), .A2(local_master_sel), .Y(
        out_local_master_sel[19]) );
  AND2X1_HVT U220 ( .A1(master_key[18]), .A2(local_master_sel), .Y(
        out_local_master_sel[18]) );
  AND2X1_HVT U221 ( .A1(master_key[17]), .A2(local_master_sel), .Y(
        out_local_master_sel[17]) );
  AND2X1_HVT U222 ( .A1(master_key[16]), .A2(local_master_sel), .Y(
        out_local_master_sel[16]) );
  AND2X1_HVT U223 ( .A1(master_key[15]), .A2(local_master_sel), .Y(
        out_local_master_sel[15]) );
  AND2X1_HVT U224 ( .A1(master_key[14]), .A2(local_master_sel), .Y(
        out_local_master_sel[14]) );
  AND2X1_HVT U225 ( .A1(master_key[13]), .A2(local_master_sel), .Y(
        out_local_master_sel[13]) );
  AND2X1_HVT U226 ( .A1(master_key[12]), .A2(local_master_sel), .Y(
        out_local_master_sel[12]) );
  AND2X1_HVT U227 ( .A1(master_key[127]), .A2(local_master_sel), .Y(
        out_local_master_sel[127]) );
  AND2X1_HVT U228 ( .A1(master_key[126]), .A2(local_master_sel), .Y(
        out_local_master_sel[126]) );
  AND2X1_HVT U229 ( .A1(master_key[125]), .A2(local_master_sel), .Y(
        out_local_master_sel[125]) );
  AND2X1_HVT U230 ( .A1(master_key[124]), .A2(local_master_sel), .Y(
        out_local_master_sel[124]) );
  AND2X1_HVT U231 ( .A1(master_key[123]), .A2(local_master_sel), .Y(
        out_local_master_sel[123]) );
  AND2X1_HVT U232 ( .A1(master_key[122]), .A2(local_master_sel), .Y(
        out_local_master_sel[122]) );
  AND2X1_HVT U233 ( .A1(master_key[121]), .A2(local_master_sel), .Y(
        out_local_master_sel[121]) );
  AND2X1_HVT U234 ( .A1(master_key[120]), .A2(local_master_sel), .Y(
        out_local_master_sel[120]) );
  AND2X1_HVT U235 ( .A1(master_key[11]), .A2(local_master_sel), .Y(
        out_local_master_sel[11]) );
  AND2X1_HVT U236 ( .A1(master_key[119]), .A2(local_master_sel), .Y(
        out_local_master_sel[119]) );
  AND2X1_HVT U237 ( .A1(master_key[118]), .A2(local_master_sel), .Y(
        out_local_master_sel[118]) );
  AND2X1_HVT U238 ( .A1(master_key[117]), .A2(local_master_sel), .Y(
        out_local_master_sel[117]) );
  AND2X1_HVT U239 ( .A1(master_key[116]), .A2(local_master_sel), .Y(
        out_local_master_sel[116]) );
  AND2X1_HVT U240 ( .A1(master_key[115]), .A2(local_master_sel), .Y(
        out_local_master_sel[115]) );
  AND2X1_HVT U241 ( .A1(master_key[114]), .A2(local_master_sel), .Y(
        out_local_master_sel[114]) );
  AND2X1_HVT U242 ( .A1(master_key[113]), .A2(local_master_sel), .Y(
        out_local_master_sel[113]) );
  AND2X1_HVT U243 ( .A1(master_key[112]), .A2(local_master_sel), .Y(
        out_local_master_sel[112]) );
  AND2X1_HVT U244 ( .A1(master_key[111]), .A2(local_master_sel), .Y(
        out_local_master_sel[111]) );
  AND2X1_HVT U245 ( .A1(master_key[110]), .A2(local_master_sel), .Y(
        out_local_master_sel[110]) );
  AND2X1_HVT U246 ( .A1(master_key[10]), .A2(local_master_sel), .Y(
        out_local_master_sel[10]) );
  AND2X1_HVT U247 ( .A1(master_key[109]), .A2(local_master_sel), .Y(
        out_local_master_sel[109]) );
  AND2X1_HVT U248 ( .A1(master_key[108]), .A2(local_master_sel), .Y(
        out_local_master_sel[108]) );
  AND2X1_HVT U249 ( .A1(master_key[107]), .A2(local_master_sel), .Y(
        out_local_master_sel[107]) );
  AND2X1_HVT U250 ( .A1(master_key[106]), .A2(local_master_sel), .Y(
        out_local_master_sel[106]) );
  AND2X1_HVT U251 ( .A1(master_key[105]), .A2(local_master_sel), .Y(
        out_local_master_sel[105]) );
  AND2X1_HVT U252 ( .A1(master_key[104]), .A2(local_master_sel), .Y(
        out_local_master_sel[104]) );
  AND2X1_HVT U253 ( .A1(master_key[103]), .A2(local_master_sel), .Y(
        out_local_master_sel[103]) );
  AND2X1_HVT U254 ( .A1(master_key[102]), .A2(local_master_sel), .Y(
        out_local_master_sel[102]) );
  AND2X1_HVT U255 ( .A1(master_key[101]), .A2(local_master_sel), .Y(
        out_local_master_sel[101]) );
  AND2X1_HVT U256 ( .A1(master_key[100]), .A2(local_master_sel), .Y(
        out_local_master_sel[100]) );
  AND2X1_HVT U257 ( .A1(master_key[0]), .A2(local_master_sel), .Y(
        out_local_master_sel[0]) );
  MUX21X1_HVT U258 ( .A1(data_flash[137]), .A2(account[9]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[9]) );
  MUX21X1_HVT U259 ( .A1(data_flash[227]), .A2(account[99]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[99]) );
  MUX21X1_HVT U260 ( .A1(data_flash[226]), .A2(account[98]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[98]) );
  MUX21X1_HVT U261 ( .A1(data_flash[225]), .A2(account[97]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[97]) );
  MUX21X1_HVT U262 ( .A1(data_flash[224]), .A2(account[96]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[96]) );
  MUX21X1_HVT U263 ( .A1(data_flash[223]), .A2(account[95]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[95]) );
  MUX21X1_HVT U264 ( .A1(data_flash[222]), .A2(account[94]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[94]) );
  MUX21X1_HVT U265 ( .A1(data_flash[221]), .A2(account[93]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[93]) );
  MUX21X1_HVT U266 ( .A1(data_flash[220]), .A2(account[92]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[92]) );
  MUX21X1_HVT U267 ( .A1(data_flash[219]), .A2(account[91]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[91]) );
  MUX21X1_HVT U268 ( .A1(data_flash[218]), .A2(account[90]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[90]) );
  MUX21X1_HVT U269 ( .A1(data_flash[136]), .A2(account[8]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[8]) );
  MUX21X1_HVT U270 ( .A1(data_flash[217]), .A2(account[89]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[89]) );
  MUX21X1_HVT U271 ( .A1(data_flash[216]), .A2(account[88]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[88]) );
  MUX21X1_HVT U272 ( .A1(data_flash[215]), .A2(account[87]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[87]) );
  MUX21X1_HVT U273 ( .A1(data_flash[214]), .A2(account[86]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[86]) );
  MUX21X1_HVT U274 ( .A1(data_flash[213]), .A2(account[85]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[85]) );
  MUX21X1_HVT U275 ( .A1(data_flash[212]), .A2(account[84]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[84]) );
  MUX21X1_HVT U276 ( .A1(data_flash[211]), .A2(account[83]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[83]) );
  MUX21X1_HVT U277 ( .A1(data_flash[210]), .A2(account[82]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[82]) );
  MUX21X1_HVT U278 ( .A1(data_flash[209]), .A2(account[81]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[81]) );
  MUX21X1_HVT U279 ( .A1(data_flash[208]), .A2(account[80]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[80]) );
  MUX21X1_HVT U280 ( .A1(data_flash[135]), .A2(account[7]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[7]) );
  MUX21X1_HVT U281 ( .A1(data_flash[207]), .A2(account[79]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[79]) );
  MUX21X1_HVT U282 ( .A1(data_flash[206]), .A2(account[78]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[78]) );
  MUX21X1_HVT U283 ( .A1(data_flash[205]), .A2(account[77]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[77]) );
  MUX21X1_HVT U284 ( .A1(data_flash[204]), .A2(account[76]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[76]) );
  MUX21X1_HVT U285 ( .A1(data_flash[203]), .A2(account[75]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[75]) );
  MUX21X1_HVT U286 ( .A1(data_flash[202]), .A2(account[74]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[74]) );
  MUX21X1_HVT U287 ( .A1(data_flash[201]), .A2(account[73]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[73]) );
  MUX21X1_HVT U288 ( .A1(data_flash[200]), .A2(account[72]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[72]) );
  MUX21X1_HVT U289 ( .A1(data_flash[199]), .A2(account[71]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[71]) );
  MUX21X1_HVT U290 ( .A1(data_flash[198]), .A2(account[70]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[70]) );
  MUX21X1_HVT U291 ( .A1(data_flash[134]), .A2(account[6]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[6]) );
  MUX21X1_HVT U292 ( .A1(data_flash[197]), .A2(account[69]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[69]) );
  MUX21X1_HVT U293 ( .A1(data_flash[196]), .A2(account[68]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[68]) );
  MUX21X1_HVT U294 ( .A1(data_flash[195]), .A2(account[67]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[67]) );
  MUX21X1_HVT U295 ( .A1(data_flash[194]), .A2(account[66]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[66]) );
  MUX21X1_HVT U296 ( .A1(data_flash[193]), .A2(account[65]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[65]) );
  MUX21X1_HVT U297 ( .A1(data_flash[192]), .A2(account[64]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[64]) );
  MUX21X1_HVT U298 ( .A1(data_flash[191]), .A2(account[63]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[63]) );
  MUX21X1_HVT U299 ( .A1(data_flash[190]), .A2(account[62]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[62]) );
  MUX21X1_HVT U300 ( .A1(data_flash[189]), .A2(account[61]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[61]) );
  MUX21X1_HVT U301 ( .A1(data_flash[188]), .A2(account[60]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[60]) );
  MUX21X1_HVT U302 ( .A1(data_flash[133]), .A2(account[5]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[5]) );
  MUX21X1_HVT U303 ( .A1(data_flash[187]), .A2(account[59]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[59]) );
  MUX21X1_HVT U304 ( .A1(data_flash[186]), .A2(account[58]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[58]) );
  MUX21X1_HVT U305 ( .A1(data_flash[185]), .A2(account[57]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[57]) );
  MUX21X1_HVT U306 ( .A1(data_flash[184]), .A2(account[56]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[56]) );
  MUX21X1_HVT U307 ( .A1(data_flash[183]), .A2(account[55]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[55]) );
  MUX21X1_HVT U308 ( .A1(data_flash[182]), .A2(account[54]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[54]) );
  MUX21X1_HVT U309 ( .A1(data_flash[181]), .A2(account[53]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[53]) );
  MUX21X1_HVT U310 ( .A1(data_flash[180]), .A2(account[52]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[52]) );
  MUX21X1_HVT U311 ( .A1(data_flash[179]), .A2(account[51]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[51]) );
  MUX21X1_HVT U312 ( .A1(data_flash[178]), .A2(account[50]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[50]) );
  MUX21X1_HVT U313 ( .A1(data_flash[132]), .A2(account[4]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[4]) );
  MUX21X1_HVT U314 ( .A1(data_flash[177]), .A2(account[49]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[49]) );
  MUX21X1_HVT U315 ( .A1(data_flash[176]), .A2(account[48]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[48]) );
  MUX21X1_HVT U316 ( .A1(data_flash[175]), .A2(account[47]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[47]) );
  MUX21X1_HVT U317 ( .A1(data_flash[174]), .A2(account[46]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[46]) );
  MUX21X1_HVT U318 ( .A1(data_flash[173]), .A2(account[45]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[45]) );
  MUX21X1_HVT U319 ( .A1(data_flash[172]), .A2(account[44]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[44]) );
  MUX21X1_HVT U320 ( .A1(data_flash[171]), .A2(account[43]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[43]) );
  MUX21X1_HVT U321 ( .A1(data_flash[170]), .A2(account[42]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[42]) );
  MUX21X1_HVT U322 ( .A1(data_flash[169]), .A2(account[41]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[41]) );
  MUX21X1_HVT U323 ( .A1(data_flash[168]), .A2(account[40]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[40]) );
  MUX21X1_HVT U324 ( .A1(data_flash[131]), .A2(account[3]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[3]) );
  MUX21X1_HVT U325 ( .A1(data_flash[167]), .A2(account[39]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[39]) );
  MUX21X1_HVT U326 ( .A1(data_flash[166]), .A2(account[38]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[38]) );
  MUX21X1_HVT U327 ( .A1(data_flash[165]), .A2(account[37]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[37]) );
  MUX21X1_HVT U328 ( .A1(data_flash[164]), .A2(account[36]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[36]) );
  MUX21X1_HVT U329 ( .A1(data_flash[163]), .A2(account[35]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[35]) );
  MUX21X1_HVT U330 ( .A1(data_flash[162]), .A2(account[34]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[34]) );
  MUX21X1_HVT U331 ( .A1(data_flash[161]), .A2(account[33]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[33]) );
  MUX21X1_HVT U332 ( .A1(data_flash[160]), .A2(account[32]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[32]) );
  MUX21X1_HVT U333 ( .A1(data_flash[159]), .A2(account[31]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[31]) );
  MUX21X1_HVT U334 ( .A1(data_flash[158]), .A2(account[30]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[30]) );
  MUX21X1_HVT U335 ( .A1(data_flash[130]), .A2(account[2]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[2]) );
  MUX21X1_HVT U336 ( .A1(data_flash[157]), .A2(account[29]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[29]) );
  MUX21X1_HVT U337 ( .A1(data_flash[156]), .A2(account[28]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[28]) );
  MUX21X1_HVT U338 ( .A1(data_flash[155]), .A2(account[27]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[27]) );
  MUX21X1_HVT U339 ( .A1(data_flash[154]), .A2(account[26]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[26]) );
  MUX21X1_HVT U340 ( .A1(data_flash[153]), .A2(account[25]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[25]) );
  MUX21X1_HVT U341 ( .A1(data_flash[152]), .A2(account[24]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[24]) );
  MUX21X1_HVT U342 ( .A1(data_flash[151]), .A2(account[23]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[23]) );
  MUX21X1_HVT U343 ( .A1(data_flash[150]), .A2(account[22]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[22]) );
  MUX21X1_HVT U344 ( .A1(data_flash[149]), .A2(account[21]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[21]) );
  MUX21X1_HVT U345 ( .A1(data_flash[148]), .A2(account[20]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[20]) );
  MUX21X1_HVT U346 ( .A1(data_flash[129]), .A2(account[1]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[1]) );
  MUX21X1_HVT U347 ( .A1(data_flash[147]), .A2(account[19]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[19]) );
  MUX21X1_HVT U348 ( .A1(data_flash[146]), .A2(account[18]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[18]) );
  MUX21X1_HVT U349 ( .A1(data_flash[145]), .A2(account[17]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[17]) );
  MUX21X1_HVT U350 ( .A1(data_flash[144]), .A2(account[16]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[16]) );
  MUX21X1_HVT U351 ( .A1(data_flash[143]), .A2(account[15]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[15]) );
  MUX21X1_HVT U352 ( .A1(data_flash[142]), .A2(account[14]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[14]) );
  MUX21X1_HVT U353 ( .A1(data_flash[141]), .A2(account[13]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[13]) );
  MUX21X1_HVT U354 ( .A1(data_flash[140]), .A2(account[12]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[12]) );
  MUX21X1_HVT U355 ( .A1(data_flash[255]), .A2(account[127]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[127]) );
  MUX21X1_HVT U356 ( .A1(data_flash[254]), .A2(account[126]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[126]) );
  MUX21X1_HVT U357 ( .A1(data_flash[253]), .A2(account[125]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[125]) );
  MUX21X1_HVT U358 ( .A1(data_flash[252]), .A2(account[124]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[124]) );
  MUX21X1_HVT U359 ( .A1(data_flash[251]), .A2(account[123]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[123]) );
  MUX21X1_HVT U360 ( .A1(data_flash[250]), .A2(account[122]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[122]) );
  MUX21X1_HVT U361 ( .A1(data_flash[249]), .A2(account[121]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[121]) );
  MUX21X1_HVT U362 ( .A1(data_flash[248]), .A2(account[120]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[120]) );
  MUX21X1_HVT U363 ( .A1(data_flash[139]), .A2(account[11]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[11]) );
  MUX21X1_HVT U364 ( .A1(data_flash[247]), .A2(account[119]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[119]) );
  MUX21X1_HVT U365 ( .A1(data_flash[246]), .A2(account[118]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[118]) );
  MUX21X1_HVT U366 ( .A1(data_flash[245]), .A2(account[117]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[117]) );
  MUX21X1_HVT U367 ( .A1(data_flash[244]), .A2(account[116]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[116]) );
  MUX21X1_HVT U368 ( .A1(data_flash[243]), .A2(account[115]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[115]) );
  MUX21X1_HVT U369 ( .A1(data_flash[242]), .A2(account[114]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[114]) );
  MUX21X1_HVT U370 ( .A1(data_flash[241]), .A2(account[113]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[113]) );
  MUX21X1_HVT U371 ( .A1(data_flash[240]), .A2(account[112]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[112]) );
  MUX21X1_HVT U372 ( .A1(data_flash[239]), .A2(account[111]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[111]) );
  MUX21X1_HVT U373 ( .A1(data_flash[238]), .A2(account[110]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[110]) );
  MUX21X1_HVT U374 ( .A1(data_flash[138]), .A2(account[10]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[10]) );
  MUX21X1_HVT U375 ( .A1(data_flash[237]), .A2(account[109]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[109]) );
  MUX21X1_HVT U376 ( .A1(data_flash[236]), .A2(account[108]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[108]) );
  MUX21X1_HVT U377 ( .A1(data_flash[235]), .A2(account[107]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[107]) );
  MUX21X1_HVT U378 ( .A1(data_flash[234]), .A2(account[106]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[106]) );
  MUX21X1_HVT U379 ( .A1(data_flash[233]), .A2(account[105]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[105]) );
  MUX21X1_HVT U380 ( .A1(data_flash[232]), .A2(account[104]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[104]) );
  MUX21X1_HVT U381 ( .A1(data_flash[231]), .A2(account[103]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[103]) );
  MUX21X1_HVT U382 ( .A1(data_flash[230]), .A2(account[102]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[102]) );
  MUX21X1_HVT U383 ( .A1(data_flash[229]), .A2(account[101]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[101]) );
  MUX21X1_HVT U384 ( .A1(data_flash[228]), .A2(account[100]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[100]) );
  MUX21X1_HVT U385 ( .A1(data_flash[128]), .A2(account[0]), .S0(
        flash_or_acc_sel), .Y(out_flash_or_acc_sel[0]) );
  MUX21X1_HVT U386 ( .A1(write_add[3]), .A2(match_add[3]), .S0(boot_lood), .Y(
        add_flash[3]) );
  MUX21X1_HVT U387 ( .A1(write_add[2]), .A2(match_add[2]), .S0(boot_lood), .Y(
        add_flash[2]) );
  MUX21X1_HVT U388 ( .A1(write_add[1]), .A2(match_add[1]), .S0(boot_lood), .Y(
        add_flash[1]) );
  MUX21X1_HVT U389 ( .A1(write_add[0]), .A2(match_add[0]), .S0(boot_lood), .Y(
        add_flash[0]) );
endmodule

