
module inv_sbox_11 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n1, n2, n24, n77, n93, n196, n197, n198, n199, n200, n201, n202, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642;

  NAND2X0_HVT U3 ( .A1(in[3]), .A2(n330), .Y(n642) );
  NAND2X0_HVT U7 ( .A1(n371), .A2(n365), .Y(n637) );
  NAND2X0_HVT U8 ( .A1(n371), .A2(n364), .Y(n636) );
  NAND2X0_HVT U9 ( .A1(n319), .A2(n636), .Y(n635) );
  NAND2X0_HVT U10 ( .A1(n319), .A2(n633), .Y(n634) );
  NAND2X0_HVT U11 ( .A1(n373), .A2(n326), .Y(n632) );
  NAND2X0_HVT U12 ( .A1(n368), .A2(n310), .Y(n631) );
  NAND2X0_HVT U13 ( .A1(n366), .A2(n248), .Y(n630) );
  NAND2X0_HVT U15 ( .A1(n361), .A2(n371), .Y(n628) );
  NAND2X0_HVT U19 ( .A1(n368), .A2(n435), .Y(n623) );
  NAND2X0_HVT U32 ( .A1(n353), .A2(n373), .Y(n612) );
  NAND2X0_HVT U35 ( .A1(n636), .A2(n436), .Y(n609) );
  NAND2X0_HVT U38 ( .A1(n351), .A2(n373), .Y(n606) );
  NAND2X0_HVT U42 ( .A1(n638), .A2(n436), .Y(n602) );
  OA21X1_HVT U53 ( .A1(n294), .A2(n594), .A3(n403), .Y(n592) );
  NAND2X0_HVT U55 ( .A1(n366), .A2(n641), .Y(n590) );
  MUX41X1_HVT U56 ( .A1(n417), .A3(n360), .A2(n401), .A4(n241), .S0(n344), 
        .S1(n295), .Y(n589) );
  AO21X1_HVT U60 ( .A1(n584), .A2(n350), .A3(n622), .Y(n585) );
  MUX41X1_HVT U62 ( .A1(n583), .A3(n589), .A2(n587), .A4(n591), .S0(n358), 
        .S1(n355), .Y(n582) );
  MUX41X1_HVT U65 ( .A1(n394), .A3(n396), .A2(n395), .A4(n606), .S0(n344), 
        .S1(n295), .Y(n579) );
  NAND2X0_HVT U66 ( .A1(n227), .A2(n338), .Y(n578) );
  MUX41X1_HVT U67 ( .A1(n392), .A3(n418), .A2(n220), .A4(n578), .S0(n349), 
        .S1(n341), .Y(n577) );
  MUX41X1_HVT U68 ( .A1(n392), .A3(n307), .A2(n393), .A4(n319), .S0(n343), 
        .S1(n295), .Y(n576) );
  MUX41X1_HVT U69 ( .A1(n576), .A3(n579), .A2(n577), .A4(n580), .S0(n358), 
        .S1(n355), .Y(n575) );
  NAND2X0_HVT U72 ( .A1(n362), .A2(n637), .Y(n573) );
  MUX41X1_HVT U73 ( .A1(n617), .A3(n573), .A2(n419), .A4(n310), .S0(n350), 
        .S1(n340), .Y(n572) );
  MUX41X1_HVT U74 ( .A1(n634), .A3(n408), .A2(n407), .A4(n1), .S0(n344), .S1(
        n377), .Y(n571) );
  MUX41X1_HVT U78 ( .A1(n569), .A3(n572), .A2(n571), .A4(n574), .S0(n358), 
        .S1(n355), .Y(n568) );
  NAND2X0_HVT U81 ( .A1(n326), .A2(n637), .Y(n565) );
  AND2X1_HVT U82 ( .A1(n638), .A2(n365), .Y(n564) );
  MUX41X1_HVT U83 ( .A1(n564), .A3(n405), .A2(n422), .A4(n565), .S0(n343), 
        .S1(n377), .Y(n563) );
  MUX41X1_HVT U85 ( .A1(n562), .A3(n566), .A2(n563), .A4(n567), .S0(n358), 
        .S1(n355), .Y(n561) );
  MUX41X1_HVT U88 ( .A1(n220), .A3(n382), .A2(n614), .A4(n598), .S0(n343), 
        .S1(n378), .Y(n559) );
  NAND2X0_HVT U89 ( .A1(n373), .A2(n313), .Y(n558) );
  MUX41X1_HVT U90 ( .A1(n316), .A3(n637), .A2(n597), .A4(n558), .S0(n343), 
        .S1(n295), .Y(n557) );
  MUX41X1_HVT U96 ( .A1(n418), .A3(n630), .A2(n402), .A4(n425), .S0(n344), 
        .S1(n293), .Y(n552) );
  MUX41X1_HVT U98 ( .A1(n551), .A3(n426), .A2(n409), .A4(n616), .S0(n344), 
        .S1(n293), .Y(n550) );
  MUX41X1_HVT U99 ( .A1(n612), .A3(n395), .A2(n596), .A4(n360), .S0(n295), 
        .S1(n341), .Y(n549) );
  NAND2X0_HVT U100 ( .A1(n373), .A2(n322), .Y(n548) );
  MUX41X1_HVT U101 ( .A1(n427), .A3(n631), .A2(n320), .A4(n548), .S0(n295), 
        .S1(n339), .Y(n547) );
  MUX41X1_HVT U102 ( .A1(n547), .A3(n550), .A2(n549), .A4(n552), .S0(n359), 
        .S1(n355), .Y(n546) );
  AND2X1_HVT U104 ( .A1(n637), .A2(n363), .Y(n545) );
  MUX41X1_HVT U105 ( .A1(n629), .A3(n428), .A2(n565), .A4(n545), .S0(n344), 
        .S1(n377), .Y(n544) );
  MUX41X1_HVT U107 ( .A1(n427), .A3(n365), .A2(n543), .A4(n386), .S0(n343), 
        .S1(n349), .Y(n542) );
  MUX41X1_HVT U108 ( .A1(n1), .A3(n360), .A2(n401), .A4(n325), .S0(n344), .S1(
        n377), .Y(n541) );
  MUX41X1_HVT U109 ( .A1(n426), .A3(n382), .A2(n423), .A4(n415), .S0(n343), 
        .S1(n293), .Y(n540) );
  MUX41X1_HVT U110 ( .A1(n540), .A3(n542), .A2(n541), .A4(n544), .S0(n359), 
        .S1(in[1]), .Y(n539) );
  AO21X1_HVT U112 ( .A1(n411), .A2(n349), .A3(n620), .Y(n537) );
  NAND2X0_HVT U114 ( .A1(n319), .A2(n637), .Y(n535) );
  MUX41X1_HVT U115 ( .A1(n535), .A3(n632), .A2(n411), .A4(n366), .S0(n295), 
        .S1(n341), .Y(n534) );
  MUX41X1_HVT U116 ( .A1(n410), .A3(n404), .A2(n382), .A4(n628), .S0(n342), 
        .S1(n378), .Y(n533) );
  NAND2X0_HVT U118 ( .A1(n373), .A2(n307), .Y(n531) );
  MUX41X1_HVT U119 ( .A1(n429), .A3(n532), .A2(n607), .A4(n531), .S0(n342), 
        .S1(n350), .Y(n530) );
  MUX41X1_HVT U120 ( .A1(n530), .A3(n534), .A2(n533), .A4(n536), .S0(n359), 
        .S1(n355), .Y(n529) );
  MUX41X1_HVT U122 ( .A1(n416), .A3(n332), .A2(n598), .A4(n420), .S0(n342), 
        .S1(n293), .Y(n528) );
  MUX41X1_HVT U124 ( .A1(n334), .A3(n527), .A2(n621), .A4(n398), .S0(n350), 
        .S1(n342), .Y(n526) );
  AOI21X1_HVT U127 ( .A1(n347), .A2(n522), .A3(n387), .Y(n523) );
  NAND2X0_HVT U129 ( .A1(n346), .A2(n318), .Y(n520) );
  MUX41X1_HVT U130 ( .A1(n520), .A3(n521), .A2(n524), .A4(n523), .S0(n350), 
        .S1(n356), .Y(n519) );
  AND2X1_HVT U131 ( .A1(n338), .A2(n292), .Y(n518) );
  MUX41X1_HVT U132 ( .A1(n276), .A3(n518), .A2(n431), .A4(n392), .S0(n350), 
        .S1(n340), .Y(n517) );
  MUX41X1_HVT U133 ( .A1(n432), .A3(n386), .A2(n241), .A4(n300), .S0(n349), 
        .S1(n339), .Y(n516) );
  MUX41X1_HVT U136 ( .A1(n595), .A3(n548), .A2(n514), .A4(n390), .S0(n346), 
        .S1(n378), .Y(n513) );
  MUX41X1_HVT U137 ( .A1(n248), .A3(n615), .A2(n619), .A4(n425), .S0(n349), 
        .S1(n339), .Y(n512) );
  MUX41X1_HVT U139 ( .A1(n511), .A3(n515), .A2(n519), .A4(n525), .S0(n359), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n407), .A3(n333), .A2(n400), .A4(n632), .S0(n349), 
        .S1(n341), .Y(n510) );
  NAND2X0_HVT U141 ( .A1(n361), .A2(n373), .Y(n509) );
  MUX41X1_HVT U142 ( .A1(n509), .A3(n605), .A2(n430), .A4(n400), .S0(n347), 
        .S1(n378), .Y(n508) );
  MUX41X1_HVT U143 ( .A1(n433), .A3(n412), .A2(n623), .A4(n621), .S0(n345), 
        .S1(n378), .Y(n507) );
  MUX41X1_HVT U145 ( .A1(n613), .A3(n428), .A2(n506), .A4(n565), .S0(n347), 
        .S1(n378), .Y(n505) );
  MUX41X1_HVT U146 ( .A1(n505), .A3(n507), .A2(n508), .A4(n510), .S0(n356), 
        .S1(n358), .Y(n504) );
  AO21X1_HVT U148 ( .A1(n349), .A2(n388), .A3(n322), .Y(n502) );
  MUX41X1_HVT U155 ( .A1(n400), .A3(n632), .A2(n624), .A4(n402), .S0(n345), 
        .S1(n293), .Y(n495) );
  MUX41X1_HVT U156 ( .A1(n495), .A3(n499), .A2(n496), .A4(n501), .S0(n359), 
        .S1(n355), .Y(n494) );
  NAND2X0_HVT U159 ( .A1(n491), .A2(n490), .Y(n492) );
  NAND2X0_HVT U163 ( .A1(n290), .A2(n433), .Y(n486) );
  MUX41X1_HVT U164 ( .A1(n635), .A3(n486), .A2(n607), .A4(n397), .S0(n342), 
        .S1(n293), .Y(n485) );
  NAND2X0_HVT U166 ( .A1(n633), .A2(n482), .Y(n483) );
  MUX41X1_HVT U173 ( .A1(n318), .A3(n316), .A2(n326), .A4(n608), .S0(n345), 
        .S1(n378), .Y(n475) );
  NAND2X0_HVT U177 ( .A1(n368), .A2(n307), .Y(n472) );
  MUX41X1_HVT U178 ( .A1(n335), .A3(n472), .A2(n315), .A4(n600), .S0(n345), 
        .S1(n293), .Y(n471) );
  AND2X1_HVT U179 ( .A1(n638), .A2(n363), .Y(n470) );
  MUX41X1_HVT U180 ( .A1(n612), .A3(n301), .A2(n470), .A4(n599), .S0(n345), 
        .S1(n293), .Y(n469) );
  MUX41X1_HVT U182 ( .A1(n386), .A3(n242), .A2(n385), .A4(n422), .S0(n342), 
        .S1(n378), .Y(n467) );
  AND2X1_HVT U185 ( .A1(n436), .A2(n292), .Y(n464) );
  NAND2X0_HVT U191 ( .A1(n380), .A2(n391), .Y(n458) );
  AND2X1_HVT U192 ( .A1(n408), .A2(n456), .Y(n457) );
  NAND2X0_HVT U194 ( .A1(n602), .A2(n456), .Y(n454) );
  MUX41X1_HVT U195 ( .A1(n455), .A3(n454), .A2(n457), .A4(n458), .S0(n343), 
        .S1(n356), .Y(n453) );
  NAND2X0_HVT U198 ( .A1(n227), .A2(n436), .Y(n633) );
  NAND2X0_HVT U200 ( .A1(n364), .A2(n373), .Y(n522) );
  NAND2X0_HVT U207 ( .A1(n373), .A2(n316), .Y(n584) );
  IBUFFX2_HVT U1 ( .A(n616), .Y(n403) );
  INVX2_HVT U2 ( .A(n360), .Y(n436) );
  IBUFFX2_HVT U4 ( .A(n345), .Y(n244) );
  MUX41X1_HVT U5 ( .A1(n554), .A3(n557), .A2(n559), .A4(n560), .S0(n355), .S1(
        n358), .Y(n553) );
  MUX41X2_HVT U6 ( .A1(n401), .A3(n424), .A2(n336), .A4(n385), .S0(n223), .S1(
        n252), .Y(n560) );
  INVX2_HVT U14 ( .A(n354), .Y(n355) );
  NBUFFX4_HVT U16 ( .A(n376), .Y(n350) );
  MUX21X1_HVT U17 ( .A1(n398), .A2(n590), .S0(n350), .Y(n586) );
  INVX0_HVT U18 ( .A(n350), .Y(n221) );
  MUX21X1_HVT U20 ( .A1(n353), .A2(n310), .S0(n312), .Y(n599) );
  IBUFFX2_HVT U21 ( .A(n372), .Y(n290) );
  NBUFFX2_HVT U22 ( .A(n376), .Y(n348) );
  INVX1_HVT U23 ( .A(n622), .Y(n1) );
  IBUFFX2_HVT U24 ( .A(n348), .Y(n252) );
  INVX1_HVT U25 ( .A(n380), .Y(n218) );
  IBUFFX2_HVT U26 ( .A(n350), .Y(n274) );
  MUX21X1_HVT U27 ( .A1(n414), .A2(n334), .S0(n348), .Y(n455) );
  MUX41X1_HVT U28 ( .A1(n489), .A3(n487), .A2(n485), .A4(n481), .S0(n2), .S1(
        n289), .Y(n480) );
  IBUFFX16_HVT U29 ( .A(n219), .Y(n2) );
  MUX21X2_HVT U30 ( .A1(n419), .A2(n603), .S0(n222), .Y(n461) );
  INVX2_HVT U31 ( .A(n372), .Y(n291) );
  NAND2X0_HVT U33 ( .A1(n568), .A2(n24), .Y(n77) );
  NAND2X0_HVT U34 ( .A1(n561), .A2(n303), .Y(n93) );
  NAND2X0_HVT U36 ( .A1(n77), .A2(n93), .Y(out[1]) );
  IBUFFX2_HVT U37 ( .A(n303), .Y(n24) );
  MUX21X2_HVT U39 ( .A1(n402), .A2(n393), .S0(n348), .Y(n593) );
  NAND2X0_HVT U40 ( .A1(n504), .A2(n196), .Y(n197) );
  NAND2X0_HVT U41 ( .A1(n494), .A2(n273), .Y(n198) );
  NAND2X0_HVT U43 ( .A1(n197), .A2(n198), .Y(out[5]) );
  INVX1_HVT U44 ( .A(n273), .Y(n196) );
  IBUFFX2_HVT U45 ( .A(in[7]), .Y(n273) );
  MUX21X1_HVT U46 ( .A1(n1), .A2(n581), .S0(n337), .Y(n580) );
  MUX41X1_HVT U47 ( .A1(n404), .A3(n336), .A2(n619), .A4(n423), .S0(n199), 
        .S1(n377), .Y(n562) );
  IBUFFX16_HVT U48 ( .A(n344), .Y(n199) );
  NAND2X0_HVT U49 ( .A1(n336), .A2(n200), .Y(n201) );
  NAND2X0_HVT U50 ( .A1(n619), .A2(n221), .Y(n202) );
  NAND2X0_HVT U51 ( .A1(n201), .A2(n202), .Y(n498) );
  INVX0_HVT U52 ( .A(n221), .Y(n200) );
  MUX21X1_HVT U54 ( .A1(n497), .A2(n498), .S0(n347), .Y(n496) );
  INVX0_HVT U57 ( .A(n220), .Y(n626) );
  INVX0_HVT U58 ( .A(n619), .Y(n400) );
  MUX21X1_HVT U59 ( .A1(n310), .A2(n435), .S0(n370), .Y(n601) );
  MUX21X1_HVT U61 ( .A1(n601), .A2(n420), .S0(n218), .Y(n493) );
  IBUFFX16_HVT U63 ( .A(n354), .Y(n219) );
  IBUFFX2_HVT U64 ( .A(n349), .Y(n283) );
  MUX21X2_HVT U70 ( .A1(n387), .A2(n603), .S0(n348), .Y(n538) );
  INVX4_HVT U71 ( .A(n370), .Y(n373) );
  MUX21X1_HVT U75 ( .A1(n437), .A2(n317), .S0(n291), .Y(n220) );
  INVX0_HVT U76 ( .A(n317), .Y(n319) );
  IBUFFX16_HVT U77 ( .A(n252), .Y(n222) );
  MUX21X2_HVT U79 ( .A1(n537), .A2(n538), .S0(n347), .Y(n536) );
  MUX21X1_HVT U80 ( .A1(n313), .A2(n315), .S0(n367), .Y(n600) );
  XOR2X1_HVT U84 ( .A1(n363), .A2(n369), .Y(n596) );
  INVX0_HVT U86 ( .A(n348), .Y(n279) );
  INVX1_HVT U87 ( .A(n555), .Y(n281) );
  IBUFFX16_HVT U91 ( .A(n342), .Y(n223) );
  IBUFFX2_HVT U92 ( .A(n380), .Y(n295) );
  INVX1_HVT U93 ( .A(in[1]), .Y(n354) );
  NAND2X0_HVT U94 ( .A1(n575), .A2(n224), .Y(n225) );
  NAND2X0_HVT U95 ( .A1(n582), .A2(in[7]), .Y(n226) );
  NAND2X0_HVT U97 ( .A1(n225), .A2(n226), .Y(out[0]) );
  IBUFFX2_HVT U103 ( .A(in[7]), .Y(n224) );
  MUX21X2_HVT U106 ( .A1(n281), .A2(n277), .S0(n282), .Y(n280) );
  INVX1_HVT U111 ( .A(n292), .Y(n227) );
  INVX1_HVT U113 ( .A(n641), .Y(n385) );
  MUX41X1_HVT U117 ( .A1(n331), .A3(n558), .A2(n327), .A4(n477), .S0(n379), 
        .S1(n345), .Y(n476) );
  IBUFFX2_HVT U121 ( .A(n379), .Y(n378) );
  MUX21X2_HVT U123 ( .A1(n483), .A2(n484), .S0(n346), .Y(n481) );
  INVX1_HVT U125 ( .A(n292), .Y(n368) );
  MUX21X2_HVT U126 ( .A1(n399), .A2(n588), .S0(n337), .Y(n587) );
  NAND2X0_HVT U128 ( .A1(n471), .A2(n228), .Y(n229) );
  NAND2X0_HVT U134 ( .A1(n469), .A2(n243), .Y(n230) );
  NAND2X0_HVT U135 ( .A1(n229), .A2(n230), .Y(n468) );
  INVX0_HVT U138 ( .A(n243), .Y(n228) );
  MUX41X1_HVT U144 ( .A1(n421), .A3(n635), .A2(n417), .A4(n640), .S0(n377), 
        .S1(n343), .Y(n566) );
  IBUFFX2_HVT U147 ( .A(n380), .Y(n377) );
  NAND2X0_HVT U149 ( .A1(n328), .A2(n231), .Y(n232) );
  NAND2X0_HVT U150 ( .A1(n362), .A2(n312), .Y(n233) );
  NAND2X0_HVT U151 ( .A1(n232), .A2(n233), .Y(n311) );
  INVX0_HVT U152 ( .A(n312), .Y(n231) );
  NAND2X0_HVT U153 ( .A1(n528), .A2(n234), .Y(n235) );
  NAND2X0_HVT U154 ( .A1(n526), .A2(n238), .Y(n236) );
  NAND2X0_HVT U157 ( .A1(n235), .A2(n236), .Y(n525) );
  INVX0_HVT U158 ( .A(n238), .Y(n234) );
  IBUFFX2_HVT U160 ( .A(n356), .Y(n238) );
  MUX41X1_HVT U161 ( .A1(n625), .A3(n626), .A2(n404), .A4(n406), .S0(n377), 
        .S1(n237), .Y(n567) );
  IBUFFX2_HVT U162 ( .A(n344), .Y(n237) );
  INVX1_HVT U165 ( .A(n372), .Y(n370) );
  OR2X1_HVT U167 ( .A1(n437), .A2(n239), .Y(n639) );
  IBUFFX16_HVT U168 ( .A(n351), .Y(n239) );
  IBUFFX2_HVT U169 ( .A(n437), .Y(n338) );
  INVX0_HVT U170 ( .A(n590), .Y(n240) );
  INVX0_HVT U171 ( .A(n240), .Y(n241) );
  INVX1_HVT U172 ( .A(n385), .Y(n242) );
  IBUFFX2_HVT U174 ( .A(n356), .Y(n243) );
  INVX1_HVT U175 ( .A(n639), .Y(n313) );
  INVX0_HVT U176 ( .A(n600), .Y(n413) );
  MUX21X2_HVT U181 ( .A1(n336), .A2(n596), .S0(n348), .Y(n462) );
  INVX0_HVT U183 ( .A(n599), .Y(n414) );
  INVX0_HVT U184 ( .A(n311), .Y(n327) );
  NAND2X0_HVT U186 ( .A1(n371), .A2(n298), .Y(n641) );
  INVX0_HVT U187 ( .A(n371), .Y(n312) );
  MUX41X1_HVT U188 ( .A1(n590), .A3(n424), .A2(n436), .A4(n432), .S0(n244), 
        .S1(n376), .Y(n474) );
  MUX21X2_HVT U189 ( .A1(n362), .A2(n353), .S0(n291), .Y(n619) );
  NAND2X0_HVT U190 ( .A1(n546), .A2(n245), .Y(n246) );
  NAND2X0_HVT U193 ( .A1(n553), .A2(n253), .Y(n247) );
  NAND2X0_HVT U196 ( .A1(n246), .A2(n247), .Y(out[2]) );
  INVX1_HVT U197 ( .A(n253), .Y(n245) );
  INVX0_HVT U199 ( .A(n388), .Y(n248) );
  IBUFFX2_HVT U201 ( .A(n303), .Y(n253) );
  INVX0_HVT U202 ( .A(n636), .Y(n388) );
  NAND2X0_HVT U203 ( .A1(n467), .A2(n249), .Y(n250) );
  NAND2X0_HVT U204 ( .A1(n466), .A2(n254), .Y(n251) );
  NAND2X0_HVT U205 ( .A1(n250), .A2(n251), .Y(n465) );
  INVX0_HVT U206 ( .A(n254), .Y(n249) );
  IBUFFX2_HVT U208 ( .A(n356), .Y(n254) );
  IBUFFX2_HVT U209 ( .A(n638), .Y(n300) );
  MUX21X1_HVT U210 ( .A1(n353), .A2(n322), .S0(n292), .Y(n450) );
  INVX1_HVT U211 ( .A(n615), .Y(n404) );
  INVX1_HVT U212 ( .A(n450), .Y(n419) );
  INVX1_HVT U213 ( .A(n363), .Y(n433) );
  INVX2_HVT U214 ( .A(n376), .Y(n380) );
  NAND2X0_HVT U215 ( .A1(n502), .A2(n255), .Y(n256) );
  NAND2X0_HVT U216 ( .A1(n503), .A2(n267), .Y(n257) );
  NAND2X0_HVT U217 ( .A1(n256), .A2(n257), .Y(n501) );
  INVX0_HVT U218 ( .A(n267), .Y(n255) );
  NAND2X0_HVT U219 ( .A1(n325), .A2(n258), .Y(n259) );
  NAND2X0_HVT U220 ( .A1(n363), .A2(n272), .Y(n260) );
  NAND2X0_HVT U221 ( .A1(n259), .A2(n260), .Y(n439) );
  INVX0_HVT U222 ( .A(n272), .Y(n258) );
  MUX21X1_HVT U223 ( .A1(n431), .A2(n276), .S0(n349), .Y(n503) );
  IBUFFX2_HVT U224 ( .A(n346), .Y(n267) );
  INVX0_HVT U225 ( .A(n323), .Y(n325) );
  INVX0_HVT U226 ( .A(n439), .Y(n431) );
  INVX0_HVT U227 ( .A(n601), .Y(n412) );
  OA21X1_HVT U228 ( .A1(n383), .A2(n294), .A3(n389), .Y(n497) );
  NAND2X0_HVT U229 ( .A1(n464), .A2(n261), .Y(n262) );
  NAND2X0_HVT U230 ( .A1(n421), .A2(n350), .Y(n263) );
  NAND2X0_HVT U231 ( .A1(n262), .A2(n263), .Y(n463) );
  IBUFFX2_HVT U232 ( .A(n350), .Y(n261) );
  NAND2X0_HVT U233 ( .A1(n242), .A2(n264), .Y(n265) );
  NAND2X0_HVT U234 ( .A1(n311), .A2(n271), .Y(n266) );
  NAND2X0_HVT U235 ( .A1(n266), .A2(n265), .Y(n581) );
  INVX0_HVT U236 ( .A(n271), .Y(n264) );
  IBUFFX2_HVT U237 ( .A(n346), .Y(n271) );
  INVX1_HVT U238 ( .A(n280), .Y(n554) );
  IBUFFX2_HVT U239 ( .A(n367), .Y(n272) );
  MUX41X1_HVT U240 ( .A1(n461), .A3(n460), .A2(n462), .A4(n463), .S0(n340), 
        .S1(n356), .Y(n459) );
  OA21X1_HVT U241 ( .A1(n404), .A2(n294), .A3(n584), .Y(n460) );
  INVX1_HVT U242 ( .A(n354), .Y(n356) );
  NAND2X0_HVT U243 ( .A1(n492), .A2(n268), .Y(n269) );
  NAND2X0_HVT U244 ( .A1(n493), .A2(n347), .Y(n270) );
  NAND2X0_HVT U245 ( .A1(n269), .A2(n270), .Y(n489) );
  IBUFFX2_HVT U246 ( .A(n347), .Y(n268) );
  INVX0_HVT U247 ( .A(n276), .Y(n640) );
  MUX41X1_HVT U248 ( .A1(n500), .A3(n311), .A2(n409), .A4(n422), .S0(n274), 
        .S1(n275), .Y(n499) );
  IBUFFX16_HVT U249 ( .A(n339), .Y(n275) );
  INVX1_HVT U250 ( .A(n285), .Y(n569) );
  INVX1_HVT U251 ( .A(n570), .Y(n286) );
  MUX21X1_HVT U252 ( .A1(n420), .A2(n381), .S0(n349), .Y(n570) );
  AND2X1_HVT U253 ( .A1(n641), .A2(n364), .Y(n276) );
  AO21X1_HVT U254 ( .A1(n362), .A2(n242), .A3(n294), .Y(n482) );
  MUX21X1_HVT U255 ( .A1(n278), .A2(n609), .S0(n279), .Y(n277) );
  IBUFFX16_HVT U256 ( .A(n361), .Y(n278) );
  IBUFFX16_HVT U257 ( .A(n346), .Y(n282) );
  INVX1_HVT U258 ( .A(in[4]), .Y(n379) );
  INVX1_HVT U259 ( .A(n292), .Y(n371) );
  INVX2_HVT U260 ( .A(n370), .Y(n292) );
  INVX1_HVT U261 ( .A(n448), .Y(n421) );
  MUX21X1_HVT U262 ( .A1(n433), .A2(n338), .S0(n292), .Y(n452) );
  MUX41X1_HVT U263 ( .A1(n602), .A3(n397), .A2(n417), .A4(n412), .S0(n283), 
        .S1(n284), .Y(n466) );
  IBUFFX16_HVT U264 ( .A(n340), .Y(n284) );
  INVX1_HVT U265 ( .A(n452), .Y(n417) );
  MUX21X1_HVT U266 ( .A1(n310), .A2(n435), .S0(n292), .Y(n449) );
  MUX21X1_HVT U267 ( .A1(n288), .A2(n286), .S0(n287), .Y(n285) );
  IBUFFX16_HVT U268 ( .A(n347), .Y(n287) );
  OAI21X1_HVT U269 ( .A1(n384), .A2(n294), .A3(n622), .Y(n288) );
  IBUFFX16_HVT U270 ( .A(n359), .Y(n289) );
  INVX1_HVT U271 ( .A(in[0]), .Y(n372) );
  INVX1_HVT U272 ( .A(n449), .Y(n420) );
  NAND2X0_HVT U273 ( .A1(n529), .A2(n303), .Y(n296) );
  INVX0_HVT U274 ( .A(n317), .Y(n314) );
  INVX0_HVT U275 ( .A(n328), .Y(n324) );
  INVX1_HVT U276 ( .A(in[5]), .Y(n357) );
  INVX1_HVT U277 ( .A(n376), .Y(n294) );
  INVX0_HVT U278 ( .A(in[6]), .Y(n437) );
  INVX2_HVT U279 ( .A(n379), .Y(n376) );
  INVX1_HVT U280 ( .A(n617), .Y(n402) );
  IBUFFX2_HVT U281 ( .A(n372), .Y(n367) );
  IBUFFX2_HVT U282 ( .A(n372), .Y(n369) );
  INVX1_HVT U283 ( .A(n622), .Y(n397) );
  INVX0_HVT U284 ( .A(n621), .Y(n398) );
  XNOR2X1_HVT U285 ( .A1(n352), .A2(n434), .Y(n627) );
  IBUFFX2_HVT U286 ( .A(n379), .Y(n293) );
  AO21X2_HVT U287 ( .A1(n292), .A2(n318), .A3(n294), .Y(n490) );
  AO21X2_HVT U288 ( .A1(n369), .A2(n324), .A3(n294), .Y(n456) );
  MUX21X1_HVT U289 ( .A1(n593), .A2(n592), .S0(n346), .Y(n591) );
  NAND2X0_HVT U290 ( .A1(n539), .A2(in[7]), .Y(n297) );
  NAND2X0_HVT U291 ( .A1(n296), .A2(n297), .Y(out[3]) );
  INVX1_HVT U292 ( .A(n329), .Y(n477) );
  INVX0_HVT U293 ( .A(n320), .Y(n608) );
  INVX0_HVT U294 ( .A(n299), .Y(n574) );
  NAND2X0_HVT U295 ( .A1(n351), .A2(n352), .Y(n298) );
  INVX1_HVT U296 ( .A(n352), .Y(n330) );
  INVX0_HVT U297 ( .A(in[7]), .Y(n303) );
  OR2X1_HVT U298 ( .A1(n330), .A2(n434), .Y(n321) );
  INVX1_HVT U299 ( .A(n321), .Y(n317) );
  INVX0_HVT U300 ( .A(n632), .Y(n301) );
  NAND2X0_HVT U301 ( .A1(n371), .A2(n319), .Y(n638) );
  INVX0_HVT U302 ( .A(n343), .Y(n302) );
  MUX41X1_HVT U303 ( .A1(n468), .A3(n465), .A2(n459), .A4(n453), .S0(n357), 
        .S1(n303), .Y(out[7]) );
  INVX1_HVT U304 ( .A(n357), .Y(n359) );
  MUX41X1_HVT U305 ( .A1(n609), .A3(n301), .A2(n314), .A4(n300), .S0(n302), 
        .S1(n380), .Y(n299) );
  NAND2X0_HVT U306 ( .A1(n480), .A2(n304), .Y(n305) );
  NAND2X0_HVT U307 ( .A1(n473), .A2(n303), .Y(n306) );
  NAND2X0_HVT U308 ( .A1(n305), .A2(n306), .Y(out[6]) );
  INVX1_HVT U309 ( .A(n303), .Y(n304) );
  INVX1_HVT U310 ( .A(n351), .Y(n307) );
  NAND2X0_HVT U311 ( .A1(n618), .A2(n294), .Y(n308) );
  NAND2X0_HVT U312 ( .A1(n621), .A2(n348), .Y(n309) );
  NAND2X0_HVT U313 ( .A1(n308), .A2(n309), .Y(n484) );
  INVX1_HVT U314 ( .A(n447), .Y(n422) );
  MUX41X1_HVT U315 ( .A1(n609), .A3(n488), .A2(n413), .A4(n396), .S0(n345), 
        .S1(n380), .Y(n487) );
  NBUFFX2_HVT U316 ( .A(n434), .Y(n310) );
  INVX1_HVT U317 ( .A(n314), .Y(n315) );
  INVX1_HVT U318 ( .A(n314), .Y(n316) );
  INVX1_HVT U319 ( .A(n317), .Y(n318) );
  MUX21X1_HVT U320 ( .A1(n361), .A2(n330), .S0(n373), .Y(n320) );
  INVX1_HVT U321 ( .A(n298), .Y(n322) );
  INVX1_HVT U322 ( .A(n298), .Y(n323) );
  INVX1_HVT U323 ( .A(n322), .Y(n326) );
  NAND2X0_HVT U324 ( .A1(n351), .A2(n352), .Y(n328) );
  INVX1_HVT U325 ( .A(n438), .Y(n432) );
  MUX21X1_HVT U326 ( .A1(n435), .A2(n316), .S0(n373), .Y(n479) );
  MUX41X1_HVT U327 ( .A1(n479), .A3(n334), .A2(n331), .A4(n335), .S0(n302), 
        .S1(n294), .Y(n478) );
  NBUFFX2_HVT U328 ( .A(n434), .Y(n351) );
  MUX21X1_HVT U329 ( .A1(n330), .A2(n318), .S0(n312), .Y(n329) );
  INVX0_HVT U330 ( .A(in[3]), .Y(n434) );
  MUX41X1_HVT U331 ( .A1(n478), .A3(n476), .A2(n475), .A4(n474), .S0(n354), 
        .S1(n357), .Y(n473) );
  MUX21X2_HVT U332 ( .A1(n512), .A2(n513), .S0(n356), .Y(n511) );
  NBUFFX2_HVT U333 ( .A(n639), .Y(n363) );
  AND2X1_HVT U334 ( .A1(n638), .A2(n326), .Y(n331) );
  NBUFFX2_HVT U335 ( .A(n639), .Y(n364) );
  AND2X1_HVT U336 ( .A1(n326), .A2(n628), .Y(n332) );
  MUX21X1_HVT U337 ( .A1(n363), .A2(n365), .S0(n290), .Y(n488) );
  MUX21X1_HVT U338 ( .A1(n323), .A2(n436), .S0(n291), .Y(n611) );
  MUX21X1_HVT U339 ( .A1(n310), .A2(n323), .S0(n369), .Y(n614) );
  MUX21X1_HVT U340 ( .A1(n586), .A2(n585), .S0(n346), .Y(n583) );
  MUX21X1_HVT U341 ( .A1(n310), .A2(n436), .S0(n290), .Y(n447) );
  MUX21X1_HVT U342 ( .A1(n362), .A2(n313), .S0(n290), .Y(n610) );
  MUX21X1_HVT U343 ( .A1(n316), .A2(n362), .S0(n367), .Y(n445) );
  MUX21X1_HVT U344 ( .A1(n315), .A2(n313), .S0(n291), .Y(n616) );
  MUX21X1_HVT U345 ( .A1(n324), .A2(n435), .S0(n369), .Y(n594) );
  XOR2X1_HVT U346 ( .A1(n366), .A2(n290), .Y(n597) );
  MUX21X1_HVT U347 ( .A1(n310), .A2(n325), .S0(n368), .Y(n448) );
  MUX21X1_HVT U348 ( .A1(n361), .A2(n310), .S0(n290), .Y(n622) );
  MUX21X1_HVT U349 ( .A1(n361), .A2(n315), .S0(n369), .Y(n613) );
  MUX21X1_HVT U350 ( .A1(n436), .A2(n353), .S0(n291), .Y(n440) );
  MUX21X1_HVT U351 ( .A1(n556), .A2(n365), .S0(n291), .Y(n555) );
  MUX21X1_HVT U352 ( .A1(n361), .A2(n353), .S0(n348), .Y(n556) );
  MUX21X1_HVT U353 ( .A1(n328), .A2(n364), .S0(n368), .Y(n506) );
  XNOR2X1_HVT U354 ( .A1(n326), .A2(n291), .Y(n333) );
  MUX21X1_HVT U355 ( .A1(n366), .A2(n328), .S0(n367), .Y(n625) );
  MUX21X1_HVT U356 ( .A1(n436), .A2(n310), .S0(n369), .Y(n605) );
  MUX21X1_HVT U357 ( .A1(n611), .A2(n332), .S0(n347), .Y(n521) );
  MUX21X1_HVT U358 ( .A1(n400), .A2(n640), .S0(n347), .Y(n588) );
  MUX21X1_HVT U359 ( .A1(n353), .A2(n325), .S0(n227), .Y(n543) );
  XOR2X1_HVT U360 ( .A1(n318), .A2(n369), .Y(n607) );
  MUX21X1_HVT U361 ( .A1(n318), .A2(n328), .S0(n290), .Y(n629) );
  XOR2X1_HVT U362 ( .A1(n360), .A2(n369), .Y(n598) );
  MUX21X1_HVT U363 ( .A1(n365), .A2(n310), .S0(n369), .Y(n624) );
  MUX21X1_HVT U364 ( .A1(n430), .A2(n333), .S0(n346), .Y(n524) );
  MUX21X1_HVT U365 ( .A1(n310), .A2(n365), .S0(n368), .Y(n442) );
  MUX21X1_HVT U366 ( .A1(n353), .A2(n362), .S0(n367), .Y(n604) );
  NBUFFX2_HVT U367 ( .A(n376), .Y(n349) );
  AND2X1_HVT U368 ( .A1(n227), .A2(n353), .Y(n334) );
  AND2X1_HVT U369 ( .A1(n435), .A2(n373), .Y(n335) );
  AND2X1_HVT U370 ( .A1(n366), .A2(n373), .Y(n336) );
  NBUFFX2_HVT U371 ( .A(n341), .Y(n345) );
  NBUFFX2_HVT U372 ( .A(n374), .Y(n347) );
  NBUFFX2_HVT U373 ( .A(n374), .Y(n346) );
  XNOR2X1_HVT U374 ( .A1(n294), .A2(n342), .Y(n337) );
  NBUFFX2_HVT U375 ( .A(n437), .Y(n352) );
  NBUFFX2_HVT U376 ( .A(n375), .Y(n342) );
  NBUFFX2_HVT U377 ( .A(n375), .Y(n344) );
  NBUFFX2_HVT U378 ( .A(n374), .Y(n340) );
  NBUFFX2_HVT U379 ( .A(n375), .Y(n343) );
  NBUFFX2_HVT U380 ( .A(n437), .Y(n353) );
  NBUFFX2_HVT U381 ( .A(n374), .Y(n341) );
  NBUFFX2_HVT U382 ( .A(n374), .Y(n339) );
  INVX1_HVT U383 ( .A(n357), .Y(n358) );
  MUX21X1_HVT U384 ( .A1(n435), .A2(n313), .S0(n368), .Y(n532) );
  MUX21X1_HVT U385 ( .A1(n516), .A2(n517), .S0(in[1]), .Y(n515) );
  NBUFFX2_HVT U386 ( .A(in[2]), .Y(n375) );
  NBUFFX2_HVT U387 ( .A(in[2]), .Y(n374) );
  MUX21X1_HVT U388 ( .A1(n315), .A2(n307), .S0(n290), .Y(n438) );
  MUX21X1_HVT U389 ( .A1(n318), .A2(n307), .S0(n367), .Y(n491) );
  MUX21X1_HVT U390 ( .A1(n307), .A2(n364), .S0(n291), .Y(n443) );
  MUX21X1_HVT U391 ( .A1(n307), .A2(n319), .S0(n291), .Y(n444) );
  MUX21X1_HVT U392 ( .A1(n364), .A2(n307), .S0(n367), .Y(n551) );
  MUX21X1_HVT U393 ( .A1(n353), .A2(n307), .S0(n291), .Y(n617) );
  NBUFFX2_HVT U394 ( .A(n642), .Y(n365) );
  NBUFFX2_HVT U395 ( .A(n642), .Y(n366) );
  NBUFFX2_HVT U396 ( .A(n627), .Y(n360) );
  NBUFFX2_HVT U397 ( .A(n627), .Y(n361) );
  NBUFFX2_HVT U398 ( .A(n627), .Y(n362) );
  MUX21X1_HVT U399 ( .A1(n322), .A2(n307), .S0(n367), .Y(n621) );
  MUX21X1_HVT U400 ( .A1(n353), .A2(n433), .S0(n227), .Y(n500) );
  MUX21X1_HVT U401 ( .A1(n366), .A2(n353), .S0(n227), .Y(n527) );
  MUX21X1_HVT U402 ( .A1(n353), .A2(n323), .S0(n367), .Y(n618) );
  MUX21X1_HVT U403 ( .A1(n323), .A2(n338), .S0(n227), .Y(n514) );
  XOR2X1_HVT U404 ( .A1(n290), .A2(n338), .Y(n595) );
  MUX21X1_HVT U405 ( .A1(n365), .A2(n338), .S0(n227), .Y(n446) );
  MUX21X1_HVT U406 ( .A1(n338), .A2(n366), .S0(n368), .Y(n451) );
  MUX21X1_HVT U407 ( .A1(n351), .A2(n338), .S0(n290), .Y(n441) );
  MUX21X1_HVT U408 ( .A1(n338), .A2(n316), .S0(n367), .Y(n620) );
  MUX21X1_HVT U409 ( .A1(n364), .A2(n338), .S0(n369), .Y(n615) );
  MUX21X1_HVT U410 ( .A1(n338), .A2(n435), .S0(n291), .Y(n603) );
  INVX0_HVT U411 ( .A(n612), .Y(n381) );
  INVX0_HVT U412 ( .A(n606), .Y(n382) );
  INVX0_HVT U413 ( .A(n548), .Y(n383) );
  INVX0_HVT U414 ( .A(n509), .Y(n384) );
  INVX0_HVT U415 ( .A(n602), .Y(n386) );
  INVX0_HVT U416 ( .A(n637), .Y(n387) );
  INVX0_HVT U417 ( .A(n630), .Y(n389) );
  INVX0_HVT U418 ( .A(n635), .Y(n390) );
  INVX0_HVT U419 ( .A(n631), .Y(n391) );
  INVX0_HVT U420 ( .A(n629), .Y(n392) );
  INVX0_HVT U421 ( .A(n628), .Y(n393) );
  INVX0_HVT U422 ( .A(n625), .Y(n394) );
  INVX0_HVT U423 ( .A(n624), .Y(n395) );
  INVX0_HVT U424 ( .A(n623), .Y(n396) );
  INVX0_HVT U425 ( .A(n620), .Y(n399) );
  INVX0_HVT U426 ( .A(n618), .Y(n401) );
  INVX0_HVT U427 ( .A(n614), .Y(n405) );
  INVX0_HVT U428 ( .A(n613), .Y(n406) );
  INVX0_HVT U429 ( .A(n611), .Y(n407) );
  INVX0_HVT U430 ( .A(n610), .Y(n408) );
  INVX0_HVT U431 ( .A(n607), .Y(n409) );
  INVX0_HVT U432 ( .A(n605), .Y(n410) );
  INVX0_HVT U433 ( .A(n604), .Y(n411) );
  INVX0_HVT U434 ( .A(n598), .Y(n415) );
  INVX0_HVT U435 ( .A(n634), .Y(n416) );
  INVX0_HVT U436 ( .A(n451), .Y(n418) );
  INVX0_HVT U437 ( .A(n446), .Y(n423) );
  INVX0_HVT U438 ( .A(n445), .Y(n424) );
  INVX0_HVT U439 ( .A(n444), .Y(n425) );
  INVX0_HVT U440 ( .A(n443), .Y(n426) );
  INVX0_HVT U441 ( .A(n442), .Y(n427) );
  INVX0_HVT U442 ( .A(n441), .Y(n428) );
  INVX0_HVT U443 ( .A(n491), .Y(n429) );
  INVX0_HVT U444 ( .A(n440), .Y(n430) );
  INVX0_HVT U445 ( .A(n642), .Y(n435) );
endmodule

