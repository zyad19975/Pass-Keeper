
module inv_sbox_9 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346;

  MUX41X1_HVT U1 ( .A1(n1), .A3(n2), .A2(n3), .A4(n4), .S0(in[7]), .S1(n5), 
        .Y(out[7]) );
  MUX21X1_HVT U2 ( .A1(n6), .A2(n7), .S0(n8), .Y(n4) );
  AO221X1_HVT U3 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .A5(n13), .Y(n7) );
  AO22X1_HVT U4 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .Y(n13) );
  AO221X1_HVT U5 ( .A1(n18), .A2(n12), .A3(n19), .A4(n16), .A5(n20), .Y(n6) );
  AO21X1_HVT U6 ( .A1(n10), .A2(n21), .A3(n22), .Y(n20) );
  OR3X1_HVT U7 ( .A1(n23), .A2(n24), .A3(n25), .Y(n3) );
  MUX21X1_HVT U8 ( .A1(n26), .A2(n27), .S0(n8), .Y(n25) );
  AO221X1_HVT U9 ( .A1(n12), .A2(n28), .A3(n18), .A4(in[2]), .A5(n29), .Y(n27)
         );
  INVX0_HVT U10 ( .A(n30), .Y(n29) );
  NAND2X0_HVT U11 ( .A1(n31), .A2(n32), .Y(n28) );
  AO221X1_HVT U12 ( .A1(n33), .A2(n34), .A3(in[2]), .A4(n35), .A5(n16), .Y(n26) );
  OAI21X1_HVT U13 ( .A1(n36), .A2(in[2]), .A3(n37), .Y(n34) );
  MUX21X1_HVT U14 ( .A1(n38), .A2(n39), .S0(n8), .Y(n2) );
  NAND3X0_HVT U15 ( .A1(n40), .A2(n41), .A3(n42), .Y(n39) );
  OA22X1_HVT U16 ( .A1(n43), .A2(n44), .A3(n45), .A4(n37), .Y(n42) );
  NAND3X0_HVT U17 ( .A1(n46), .A2(n47), .A3(n15), .Y(n41) );
  AO21X1_HVT U18 ( .A1(n48), .A2(n49), .A3(n50), .Y(n40) );
  NAND4X0_HVT U19 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .Y(n38) );
  OA22X1_HVT U20 ( .A1(n55), .A2(n50), .A3(n56), .A4(n57), .Y(n54) );
  NAND2X0_HVT U21 ( .A1(n10), .A2(n58), .Y(n53) );
  MUX21X1_HVT U22 ( .A1(n59), .A2(n60), .S0(n8), .Y(n1) );
  AO221X1_HVT U23 ( .A1(n61), .A2(n15), .A3(n62), .A4(n12), .A5(n63), .Y(n60)
         );
  AO21X1_HVT U24 ( .A1(n64), .A2(n65), .A3(n66), .Y(n63) );
  AO21X1_HVT U25 ( .A1(n67), .A2(in[2]), .A3(n10), .Y(n64) );
  AO221X1_HVT U26 ( .A1(n68), .A2(n16), .A3(n15), .A4(n69), .A5(n70), .Y(n59)
         );
  AO22X1_HVT U27 ( .A1(n71), .A2(n12), .A3(n72), .A4(n73), .Y(n70) );
  MUX21X1_HVT U28 ( .A1(n74), .A2(n75), .S0(in[7]), .Y(out[6]) );
  AO221X1_HVT U29 ( .A1(n76), .A2(n77), .A3(n78), .A4(n79), .A5(n80), .Y(n75)
         );
  AO22X1_HVT U30 ( .A1(n81), .A2(n82), .A3(n83), .A4(n84), .Y(n80) );
  AO221X1_HVT U31 ( .A1(n15), .A2(n85), .A3(n55), .A4(n12), .A5(n86), .Y(n84)
         );
  AO21X1_HVT U32 ( .A1(n16), .A2(n87), .A3(n88), .Y(n86) );
  NAND2X0_HVT U33 ( .A1(n89), .A2(n90), .Y(n87) );
  AND2X1_HVT U34 ( .A1(n91), .A2(n92), .Y(n55) );
  NAND2X0_HVT U35 ( .A1(n73), .A2(n93), .Y(n85) );
  AO221X1_HVT U36 ( .A1(n94), .A2(n95), .A3(n10), .A4(n96), .A5(n97), .Y(n82)
         );
  AO22X1_HVT U37 ( .A1(n15), .A2(in[0]), .A3(n98), .A4(n16), .Y(n97) );
  AO221X1_HVT U38 ( .A1(n9), .A2(n16), .A3(n15), .A4(n99), .A5(n100), .Y(n79)
         );
  AO221X1_HVT U39 ( .A1(n10), .A2(n46), .A3(n12), .A4(n101), .A5(n72), .Y(n100) );
  AO221X1_HVT U40 ( .A1(n16), .A2(n102), .A3(n73), .A4(n15), .A5(n103), .Y(n77) );
  AO221X1_HVT U41 ( .A1(n104), .A2(n95), .A3(n10), .A4(n105), .A5(n22), .Y(
        n103) );
  INVX0_HVT U42 ( .A(n106), .Y(n104) );
  AO221X1_HVT U43 ( .A1(n76), .A2(n107), .A3(n78), .A4(n108), .A5(n109), .Y(
        n74) );
  AO22X1_HVT U44 ( .A1(n81), .A2(n110), .A3(n83), .A4(n111), .Y(n109) );
  NAND3X0_HVT U45 ( .A1(n112), .A2(n65), .A3(n113), .Y(n111) );
  OA221X1_HVT U46 ( .A1(n114), .A2(n37), .A3(in[4]), .A4(n49), .A5(n115), .Y(
        n113) );
  NAND3X0_HVT U47 ( .A1(n47), .A2(n116), .A3(n15), .Y(n115) );
  NAND2X0_HVT U48 ( .A1(n16), .A2(n117), .Y(n112) );
  NAND4X0_HVT U49 ( .A1(n118), .A2(n119), .A3(n51), .A4(n30), .Y(n110) );
  NAND2X0_HVT U50 ( .A1(n120), .A2(n15), .Y(n30) );
  NAND3X0_HVT U51 ( .A1(n12), .A2(n121), .A3(n122), .Y(n51) );
  NAND3X0_HVT U52 ( .A1(n47), .A2(n116), .A3(n10), .Y(n119) );
  AO21X1_HVT U53 ( .A1(n65), .A2(n123), .A3(n50), .Y(n118) );
  AO221X1_HVT U54 ( .A1(n16), .A2(n124), .A3(n15), .A4(n116), .A5(n125), .Y(
        n108) );
  MUX21X1_HVT U55 ( .A1(n10), .A2(n12), .S0(n57), .Y(n125) );
  AO221X1_HVT U56 ( .A1(n10), .A2(n126), .A3(n127), .A4(n12), .A5(n128), .Y(
        n107) );
  AO22X1_HVT U57 ( .A1(n129), .A2(n15), .A3(n73), .A4(n16), .Y(n128) );
  MUX21X1_HVT U58 ( .A1(n130), .A2(n131), .S0(in[7]), .Y(out[5]) );
  AO221X1_HVT U59 ( .A1(n81), .A2(n132), .A3(n83), .A4(n133), .A5(n134), .Y(
        n131) );
  AO22X1_HVT U60 ( .A1(n78), .A2(n135), .A3(n76), .A4(n136), .Y(n134) );
  AO221X1_HVT U61 ( .A1(n15), .A2(n137), .A3(n138), .A4(n10), .A5(n139), .Y(
        n136) );
  AO22X1_HVT U62 ( .A1(n16), .A2(n140), .A3(n12), .A4(n141), .Y(n139) );
  NAND2X0_HVT U63 ( .A1(n93), .A2(n43), .Y(n137) );
  AO221X1_HVT U64 ( .A1(n142), .A2(n12), .A3(n16), .A4(n102), .A5(n143), .Y(
        n135) );
  AO22X1_HVT U65 ( .A1(n11), .A2(n10), .A3(n15), .A4(n123), .Y(n143) );
  INVX0_HVT U66 ( .A(n96), .Y(n11) );
  NAND2X0_HVT U67 ( .A1(n48), .A2(n123), .Y(n96) );
  AO221X1_HVT U68 ( .A1(n144), .A2(n16), .A3(n145), .A4(n15), .A5(n146), .Y(
        n133) );
  AO22X1_HVT U69 ( .A1(n10), .A2(n147), .A3(n12), .A4(n148), .Y(n146) );
  AO221X1_HVT U70 ( .A1(n144), .A2(n10), .A3(n149), .A4(n12), .A5(n150), .Y(
        n132) );
  AO22X1_HVT U71 ( .A1(n151), .A2(n15), .A3(n16), .A4(n43), .Y(n150) );
  AO221X1_HVT U72 ( .A1(n76), .A2(n152), .A3(n83), .A4(n153), .A5(n154), .Y(
        n130) );
  AO22X1_HVT U73 ( .A1(n81), .A2(n155), .A3(n78), .A4(n156), .Y(n154) );
  AO22X1_HVT U74 ( .A1(n10), .A2(n157), .A3(n158), .A4(n159), .Y(n156) );
  NAND3X0_HVT U75 ( .A1(n160), .A2(n161), .A3(n162), .Y(n158) );
  AO221X1_HVT U76 ( .A1(n163), .A2(n15), .A3(n164), .A4(in[2]), .A5(n165), .Y(
        n155) );
  AO22X1_HVT U77 ( .A1(n166), .A2(n16), .A3(n167), .A4(n12), .Y(n165) );
  INVX0_HVT U78 ( .A(n93), .Y(n166) );
  AO221X1_HVT U79 ( .A1(n19), .A2(n12), .A3(n168), .A4(n15), .A5(n169), .Y(
        n153) );
  AO22X1_HVT U80 ( .A1(n170), .A2(n10), .A3(n16), .A4(n171), .Y(n169) );
  NAND2X0_HVT U81 ( .A1(n172), .A2(n173), .Y(n171) );
  AO221X1_HVT U82 ( .A1(n10), .A2(n43), .A3(n144), .A4(n12), .A5(n174), .Y(
        n152) );
  AO22X1_HVT U83 ( .A1(n15), .A2(n175), .A3(n176), .A4(n16), .Y(n174) );
  MUX41X1_HVT U84 ( .A1(n177), .A3(n178), .A2(n179), .A4(n180), .S0(n5), .S1(
        in[7]), .Y(out[4]) );
  AO21X1_HVT U85 ( .A1(n145), .A2(n12), .A3(n181), .Y(n180) );
  MUX21X1_HVT U86 ( .A1(n182), .A2(n183), .S0(n8), .Y(n181) );
  AO221X1_HVT U87 ( .A1(n184), .A2(n95), .A3(n185), .A4(n186), .A5(n187), .Y(
        n183) );
  AO21X1_HVT U88 ( .A1(n24), .A2(n188), .A3(n12), .Y(n187) );
  INVX0_HVT U89 ( .A(n189), .Y(n24) );
  AO22X1_HVT U90 ( .A1(n151), .A2(n10), .A3(n190), .A4(n89), .Y(n182) );
  OAI21X1_HVT U91 ( .A1(n90), .A2(n186), .A3(n56), .Y(n190) );
  AND2X1_HVT U92 ( .A1(n43), .A2(n36), .Y(n151) );
  AND2X1_HVT U93 ( .A1(n191), .A2(n49), .Y(n145) );
  MUX21X1_HVT U94 ( .A1(n192), .A2(n193), .S0(n8), .Y(n179) );
  NAND3X0_HVT U95 ( .A1(n194), .A2(n195), .A3(n196), .Y(n193) );
  MUX21X1_HVT U96 ( .A1(n50), .A2(n44), .S0(n102), .Y(n196) );
  NAND2X0_HVT U97 ( .A1(n120), .A2(n95), .Y(n194) );
  INVX0_HVT U98 ( .A(n49), .Y(n120) );
  AO221X1_HVT U99 ( .A1(n197), .A2(n10), .A3(n198), .A4(n12), .A5(n199), .Y(
        n192) );
  AO22X1_HVT U100 ( .A1(n15), .A2(n200), .A3(n98), .A4(n16), .Y(n199) );
  INVX0_HVT U101 ( .A(n201), .Y(n198) );
  AND2X1_HVT U102 ( .A1(n188), .A2(n116), .Y(n197) );
  MUX21X1_HVT U103 ( .A1(n202), .A2(n203), .S0(n8), .Y(n178) );
  AO221X1_HVT U104 ( .A1(n204), .A2(n16), .A3(n15), .A4(n205), .A5(n206), .Y(
        n203) );
  AO21X1_HVT U105 ( .A1(n10), .A2(n157), .A3(n207), .Y(n206) );
  AO221X1_HVT U106 ( .A1(n10), .A2(n162), .A3(n208), .A4(n16), .A5(n209), .Y(
        n202) );
  AO22X1_HVT U107 ( .A1(n15), .A2(n210), .A3(n12), .A4(n211), .Y(n209) );
  NAND2X0_HVT U108 ( .A1(n212), .A2(n49), .Y(n211) );
  NAND2X0_HVT U109 ( .A1(n162), .A2(n31), .Y(n210) );
  INVX0_HVT U110 ( .A(n101), .Y(n208) );
  MUX21X1_HVT U111 ( .A1(n213), .A2(n214), .S0(n8), .Y(n177) );
  AO221X1_HVT U112 ( .A1(n215), .A2(n16), .A3(n18), .A4(n15), .A5(n216), .Y(
        n214) );
  AO22X1_HVT U113 ( .A1(n129), .A2(n12), .A3(n10), .A4(n126), .Y(n216) );
  AND2X1_HVT U114 ( .A1(n65), .A2(n217), .Y(n129) );
  INVX0_HVT U115 ( .A(n47), .Y(n215) );
  AO221X1_HVT U116 ( .A1(n163), .A2(n12), .A3(n218), .A4(n16), .A5(n219), .Y(
        n213) );
  AO21X1_HVT U117 ( .A1(n167), .A2(n10), .A3(n66), .Y(n219) );
  AND2X1_HVT U118 ( .A1(n220), .A2(n15), .Y(n66) );
  AND2X1_HVT U119 ( .A1(n21), .A2(n90), .Y(n167) );
  INVX0_HVT U120 ( .A(n221), .Y(n163) );
  MUX21X1_HVT U121 ( .A1(n222), .A2(n223), .S0(in[7]), .Y(out[3]) );
  AO221X1_HVT U122 ( .A1(n76), .A2(n224), .A3(n83), .A4(n225), .A5(n226), .Y(
        n223) );
  AO22X1_HVT U123 ( .A1(n81), .A2(n227), .A3(n78), .A4(n228), .Y(n226) );
  NAND3X0_HVT U124 ( .A1(n229), .A2(n189), .A3(n230), .Y(n228) );
  NAND2X0_HVT U125 ( .A1(n16), .A2(n116), .Y(n189) );
  NAND2X0_HVT U126 ( .A1(n9), .A2(n12), .Y(n229) );
  AO221X1_HVT U127 ( .A1(n12), .A2(n231), .A3(n15), .A4(n140), .A5(n232), .Y(
        n227) );
  AO22X1_HVT U128 ( .A1(n138), .A2(n10), .A3(n233), .A4(n16), .Y(n232) );
  AND2X1_HVT U129 ( .A1(n89), .A2(n46), .Y(n233) );
  AND2X1_HVT U130 ( .A1(n48), .A2(n31), .Y(n138) );
  INVX0_HVT U131 ( .A(n218), .Y(n231) );
  AO221X1_HVT U132 ( .A1(n18), .A2(n16), .A3(n45), .A4(n15), .A5(n234), .Y(
        n225) );
  AO221X1_HVT U133 ( .A1(n10), .A2(n159), .A3(n235), .A4(n12), .A5(n22), .Y(
        n234) );
  AND2X1_HVT U134 ( .A1(n236), .A2(n15), .Y(n22) );
  INVX0_HVT U135 ( .A(n17), .Y(n18) );
  NAND2X0_HVT U136 ( .A1(n73), .A2(n47), .Y(n17) );
  AO221X1_HVT U137 ( .A1(n237), .A2(n16), .A3(n238), .A4(n15), .A5(n239), .Y(
        n224) );
  AO22X1_HVT U138 ( .A1(n240), .A2(n12), .A3(n241), .A4(n10), .Y(n239) );
  INVX0_HVT U139 ( .A(n200), .Y(n237) );
  AO221X1_HVT U140 ( .A1(n81), .A2(n242), .A3(n76), .A4(n243), .A5(n244), .Y(
        n222) );
  AO22X1_HVT U141 ( .A1(n83), .A2(n245), .A3(n78), .A4(n246), .Y(n244) );
  AO221X1_HVT U142 ( .A1(n67), .A2(n10), .A3(n247), .A4(n12), .A5(n248), .Y(
        n246) );
  AO22X1_HVT U143 ( .A1(n241), .A2(n15), .A3(n16), .A4(n188), .Y(n248) );
  INVX0_HVT U144 ( .A(n147), .Y(n247) );
  NAND2X0_HVT U145 ( .A1(n35), .A2(n191), .Y(n147) );
  AO221X1_HVT U146 ( .A1(n12), .A2(n249), .A3(n250), .A4(n10), .A5(n251), .Y(
        n245) );
  AO22X1_HVT U147 ( .A1(n15), .A2(n43), .A3(n16), .A4(n159), .Y(n251) );
  NAND2X0_HVT U148 ( .A1(n57), .A2(n89), .Y(n249) );
  AO221X1_HVT U149 ( .A1(n252), .A2(in[2]), .A3(n15), .A4(n99), .A5(n253), .Y(
        n243) );
  AO222X1_HVT U150 ( .A1(n12), .A2(n94), .A3(n72), .A4(n122), .A5(n16), .A6(
        n32), .Y(n253) );
  NAND2X0_HVT U151 ( .A1(n65), .A2(n35), .Y(n94) );
  INVX0_HVT U152 ( .A(n168), .Y(n99) );
  INVX0_HVT U153 ( .A(n173), .Y(n252) );
  AO221X1_HVT U154 ( .A1(n254), .A2(n95), .A3(n61), .A4(n16), .A5(n255), .Y(
        n242) );
  AO21X1_HVT U155 ( .A1(n250), .A2(n15), .A3(n256), .Y(n255) );
  MUX21X1_HVT U156 ( .A1(n257), .A2(n220), .S0(n44), .Y(n256) );
  INVX0_HVT U157 ( .A(n212), .Y(n220) );
  AND2X1_HVT U158 ( .A1(n188), .A2(n172), .Y(n250) );
  INVX0_HVT U159 ( .A(n92), .Y(n254) );
  MUX21X1_HVT U160 ( .A1(n258), .A2(n259), .S0(in[7]), .Y(out[2]) );
  AO221X1_HVT U161 ( .A1(n76), .A2(n260), .A3(n78), .A4(n261), .A5(n262), .Y(
        n259) );
  AO22X1_HVT U162 ( .A1(n81), .A2(n263), .A3(n83), .A4(n264), .Y(n262) );
  AO221X1_HVT U163 ( .A1(n241), .A2(n10), .A3(n265), .A4(n12), .A5(n266), .Y(
        n264) );
  AO22X1_HVT U164 ( .A1(n15), .A2(n267), .A3(n16), .A4(n200), .Y(n266) );
  NAND2X0_HVT U165 ( .A1(n148), .A2(n106), .Y(n200) );
  INVX0_HVT U166 ( .A(n48), .Y(n241) );
  AO221X1_HVT U167 ( .A1(n268), .A2(n16), .A3(n127), .A4(n15), .A5(n269), .Y(
        n263) );
  AO22X1_HVT U168 ( .A1(n236), .A2(n12), .A3(n72), .A4(n159), .Y(n269) );
  INVX0_HVT U169 ( .A(n52), .Y(n72) );
  INVX0_HVT U170 ( .A(n21), .Y(n236) );
  AND2X1_HVT U171 ( .A1(n188), .A2(n65), .Y(n127) );
  INVX0_HVT U172 ( .A(n105), .Y(n268) );
  AO221X1_HVT U173 ( .A1(n10), .A2(n89), .A3(n185), .A4(n12), .A5(n270), .Y(
        n261) );
  OAI221X1_HVT U174 ( .A1(n123), .A2(n186), .A3(n50), .A4(n114), .A5(n195), 
        .Y(n270) );
  NAND2X0_HVT U175 ( .A1(n71), .A2(n15), .Y(n195) );
  INVX0_HVT U176 ( .A(n91), .Y(n114) );
  NAND2X0_HVT U177 ( .A1(n142), .A2(n121), .Y(n91) );
  AO221X1_HVT U178 ( .A1(n45), .A2(n16), .A3(n257), .A4(in[2]), .A5(n271), .Y(
        n260) );
  MUX21X1_HVT U179 ( .A1(n207), .A2(n272), .S0(n273), .Y(n271) );
  NAND2X0_HVT U180 ( .A1(n56), .A2(n52), .Y(n272) );
  NAND2X0_HVT U181 ( .A1(n10), .A2(n121), .Y(n52) );
  INVX0_HVT U182 ( .A(n160), .Y(n207) );
  NAND2X0_HVT U183 ( .A1(n12), .A2(n93), .Y(n160) );
  INVX0_HVT U184 ( .A(n89), .Y(n257) );
  AO221X1_HVT U185 ( .A1(n81), .A2(n274), .A3(n76), .A4(n275), .A5(n276), .Y(
        n258) );
  AO22X1_HVT U186 ( .A1(n83), .A2(n277), .A3(n78), .A4(n278), .Y(n276) );
  AO221X1_HVT U187 ( .A1(n16), .A2(n273), .A3(n279), .A4(n15), .A5(n280), .Y(
        n278) );
  AO22X1_HVT U188 ( .A1(n12), .A2(n172), .A3(n10), .A4(n69), .Y(n280) );
  NAND2X0_HVT U189 ( .A1(n173), .A2(n90), .Y(n69) );
  AO221X1_HVT U190 ( .A1(n12), .A2(n281), .A3(n240), .A4(n10), .A5(n282), .Y(
        n277) );
  AO22X1_HVT U191 ( .A1(n168), .A2(n15), .A3(n16), .A4(n283), .Y(n282) );
  OA21X1_HVT U192 ( .A1(n185), .A2(in[0]), .A3(n92), .Y(n168) );
  AND2X1_HVT U193 ( .A1(n93), .A2(n32), .Y(n240) );
  NAND2X0_HVT U194 ( .A1(n90), .A2(n217), .Y(n281) );
  AO221X1_HVT U195 ( .A1(n15), .A2(n35), .A3(n284), .A4(n10), .A5(n285), .Y(
        n275) );
  AO22X1_HVT U196 ( .A1(n16), .A2(n162), .A3(n235), .A4(n12), .Y(n285) );
  AND2X1_HVT U197 ( .A1(n48), .A2(n89), .Y(n235) );
  INVX0_HVT U198 ( .A(n124), .Y(n284) );
  NAND2X0_HVT U199 ( .A1(n172), .A2(n106), .Y(n124) );
  AO221X1_HVT U200 ( .A1(n10), .A2(n286), .A3(n287), .A4(n12), .A5(n288), .Y(
        n274) );
  AO22X1_HVT U201 ( .A1(n176), .A2(n15), .A3(n204), .A4(n16), .Y(n288) );
  AND2X1_HVT U202 ( .A1(n47), .A2(n32), .Y(n204) );
  NAND2X0_HVT U203 ( .A1(in[3]), .A2(n121), .Y(n32) );
  NAND2X0_HVT U204 ( .A1(n159), .A2(n93), .Y(n286) );
  MUX21X1_HVT U205 ( .A1(n289), .A2(n290), .S0(in[7]), .Y(out[1]) );
  AO221X1_HVT U206 ( .A1(n81), .A2(n291), .A3(n76), .A4(n292), .A5(n293), .Y(
        n290) );
  AO22X1_HVT U207 ( .A1(n83), .A2(n294), .A3(n78), .A4(n295), .Y(n293) );
  AO221X1_HVT U208 ( .A1(n9), .A2(n16), .A3(n149), .A4(n15), .A5(n296), .Y(
        n295) );
  AO22X1_HVT U209 ( .A1(n12), .A2(n201), .A3(n33), .A4(n10), .Y(n296) );
  AND2X1_HVT U210 ( .A1(n148), .A2(n173), .Y(n33) );
  NAND2X0_HVT U211 ( .A1(n57), .A2(n106), .Y(n201) );
  INVX0_HVT U212 ( .A(n184), .Y(n149) );
  NAND2X0_HVT U213 ( .A1(n162), .A2(n106), .Y(n184) );
  AO221X1_HVT U214 ( .A1(n15), .A2(n297), .A3(n62), .A4(n10), .A5(n298), .Y(
        n294) );
  AO22X1_HVT U215 ( .A1(n16), .A2(n58), .A3(n12), .A4(n299), .Y(n298) );
  AND2X1_HVT U216 ( .A1(n162), .A2(n49), .Y(n62) );
  NAND2X0_HVT U217 ( .A1(n273), .A2(n89), .Y(n297) );
  AO222X1_HVT U218 ( .A1(n98), .A2(n12), .A3(n300), .A4(n301), .A5(n45), .A6(
        n15), .Y(n292) );
  INVX0_HVT U219 ( .A(n172), .Y(n45) );
  OAI21X1_HVT U220 ( .A1(n148), .A2(n95), .A3(n44), .Y(n300) );
  OA21X1_HVT U221 ( .A1(n159), .A2(in[0]), .A3(n35), .Y(n98) );
  AO221X1_HVT U222 ( .A1(n302), .A2(n73), .A3(n185), .A4(n10), .A5(n303), .Y(
        n291) );
  AO22X1_HVT U223 ( .A1(n15), .A2(n43), .A3(n12), .A4(n47), .Y(n303) );
  NAND2X0_HVT U224 ( .A1(n121), .A2(n116), .Y(n43) );
  AND2X1_HVT U225 ( .A1(n16), .A2(n93), .Y(n302) );
  AO221X1_HVT U226 ( .A1(n16), .A2(n304), .A3(n15), .A4(n305), .A5(n306), .Y(
        n289) );
  AO22X1_HVT U227 ( .A1(n12), .A2(n307), .A3(n10), .A4(n308), .Y(n306) );
  AO221X1_HVT U228 ( .A1(n83), .A2(n14), .A3(n81), .A4(n309), .A5(n310), .Y(
        n308) );
  AO22X1_HVT U229 ( .A1(n311), .A2(n78), .A3(n76), .A4(n67), .Y(n310) );
  INVX0_HVT U230 ( .A(n267), .Y(n311) );
  NAND2X0_HVT U231 ( .A1(n48), .A2(n36), .Y(n267) );
  AO221X1_HVT U232 ( .A1(n83), .A2(n68), .A3(n81), .A4(n67), .A5(n312), .Y(
        n307) );
  AO22X1_HVT U233 ( .A1(n76), .A2(n71), .A3(n313), .A4(n78), .Y(n312) );
  AND2X1_HVT U234 ( .A1(n47), .A2(n159), .Y(n313) );
  INVX0_HVT U235 ( .A(n314), .Y(n71) );
  INVX0_HVT U236 ( .A(n205), .Y(n67) );
  NAND2X0_HVT U237 ( .A1(n90), .A2(n31), .Y(n205) );
  NAND2X0_HVT U238 ( .A1(n46), .A2(n121), .Y(n90) );
  AND2X1_HVT U239 ( .A1(n48), .A2(n21), .Y(n68) );
  AO221X1_HVT U240 ( .A1(n83), .A2(n101), .A3(n315), .A4(n81), .A5(n316), .Y(
        n305) );
  AO22X1_HVT U241 ( .A1(n78), .A2(n19), .A3(n238), .A4(n76), .Y(n316) );
  AND2X1_HVT U242 ( .A1(n31), .A2(n314), .Y(n238) );
  NAND2X0_HVT U243 ( .A1(in[6]), .A2(in[0]), .Y(n31) );
  AND2X1_HVT U244 ( .A1(n48), .A2(n106), .Y(n19) );
  NAND2X0_HVT U245 ( .A1(n73), .A2(in[0]), .Y(n106) );
  INVX0_HVT U246 ( .A(n141), .Y(n315) );
  NAND2X0_HVT U247 ( .A1(n148), .A2(n92), .Y(n141) );
  NAND2X0_HVT U248 ( .A1(n185), .A2(in[0]), .Y(n92) );
  NAND2X0_HVT U249 ( .A1(n57), .A2(n93), .Y(n101) );
  NAND2X0_HVT U250 ( .A1(in[0]), .A2(n46), .Y(n93) );
  AO221X1_HVT U251 ( .A1(n83), .A2(n221), .A3(n81), .A4(n317), .A5(n318), .Y(
        n304) );
  AO22X1_HVT U252 ( .A1(n78), .A2(n140), .A3(n76), .A4(n157), .Y(n318) );
  NAND2X0_HVT U253 ( .A1(n116), .A2(n89), .Y(n140) );
  MUX21X1_HVT U254 ( .A1(n319), .A2(n320), .S0(in[7]), .Y(out[0]) );
  AO221X1_HVT U255 ( .A1(n83), .A2(n321), .A3(n76), .A4(n322), .A5(n323), .Y(
        n320) );
  AO22X1_HVT U256 ( .A1(n81), .A2(n324), .A3(n325), .A4(n78), .Y(n323) );
  MUX21X1_HVT U257 ( .A1(n326), .A2(n327), .S0(n328), .Y(n325) );
  MUX21X1_HVT U258 ( .A1(n221), .A2(n144), .S0(n95), .Y(n327) );
  INVX0_HVT U259 ( .A(n157), .Y(n144) );
  NAND2X0_HVT U260 ( .A1(n148), .A2(n49), .Y(n157) );
  NAND2X0_HVT U261 ( .A1(in[0]), .A2(n329), .Y(n49) );
  NAND2X0_HVT U262 ( .A1(n21), .A2(n46), .Y(n221) );
  NAND2X0_HVT U263 ( .A1(n172), .A2(n47), .Y(n326) );
  AO222X1_HVT U264 ( .A1(n176), .A2(n12), .A3(n330), .A4(n331), .A5(n332), 
        .A6(n15), .Y(n324) );
  AO21X1_HVT U265 ( .A1(in[2]), .A2(n333), .A3(n10), .Y(n331) );
  NAND2X0_HVT U266 ( .A1(n162), .A2(n123), .Y(n333) );
  INVX0_HVT U267 ( .A(n283), .Y(n330) );
  NAND2X0_HVT U268 ( .A1(n65), .A2(n173), .Y(n283) );
  INVX0_HVT U269 ( .A(n299), .Y(n176) );
  NAND2X0_HVT U270 ( .A1(n172), .A2(n217), .Y(n299) );
  AO221X1_HVT U271 ( .A1(n15), .A2(n126), .A3(in[2]), .A4(n301), .A5(n334), 
        .Y(n322) );
  AO22X1_HVT U272 ( .A1(n16), .A2(n65), .A3(n335), .A4(n12), .Y(n334) );
  INVX0_HVT U273 ( .A(n102), .Y(n335) );
  NAND2X0_HVT U274 ( .A1(n162), .A2(n217), .Y(n102) );
  NAND2X0_HVT U275 ( .A1(in[0]), .A2(in[3]), .Y(n217) );
  NAND2X0_HVT U276 ( .A1(n164), .A2(n121), .Y(n162) );
  NAND2X0_HVT U277 ( .A1(n185), .A2(n121), .Y(n65) );
  AO221X1_HVT U278 ( .A1(n14), .A2(n12), .A3(n16), .A4(n126), .A5(n336), .Y(
        n321) );
  INVX0_HVT U279 ( .A(n230), .Y(n336) );
  OA22X1_HVT U280 ( .A1(n105), .A2(n56), .A3(n44), .A4(n73), .Y(n230) );
  NAND2X0_HVT U281 ( .A1(n172), .A2(n36), .Y(n105) );
  NAND2X0_HVT U282 ( .A1(n329), .A2(n121), .Y(n172) );
  NAND2X0_HVT U283 ( .A1(n159), .A2(n21), .Y(n126) );
  AND2X1_HVT U284 ( .A1(n173), .A2(n212), .Y(n14) );
  NAND2X0_HVT U285 ( .A1(n142), .A2(in[0]), .Y(n173) );
  INVX0_HVT U286 ( .A(n46), .Y(n142) );
  NAND2X0_HVT U287 ( .A1(in[6]), .A2(n58), .Y(n46) );
  AO221X1_HVT U288 ( .A1(n76), .A2(n337), .A3(n78), .A4(n338), .A5(n339), .Y(
        n319) );
  AO22X1_HVT U289 ( .A1(n83), .A2(n340), .A3(n341), .A4(n81), .Y(n339) );
  AND2X1_HVT U290 ( .A1(in[5]), .A2(in[1]), .Y(n81) );
  MUX21X1_HVT U291 ( .A1(n9), .A2(n342), .S0(n328), .Y(n341) );
  AND2X1_HVT U292 ( .A1(n50), .A2(n37), .Y(n328) );
  MUX21X1_HVT U293 ( .A1(n21), .A2(n170), .S0(n95), .Y(n342) );
  INVX0_HVT U294 ( .A(n117), .Y(n170) );
  NAND2X0_HVT U295 ( .A1(n36), .A2(n191), .Y(n117) );
  NAND2X0_HVT U296 ( .A1(n73), .A2(n121), .Y(n191) );
  INVX0_HVT U297 ( .A(n273), .Y(n73) );
  NAND2X0_HVT U298 ( .A1(n164), .A2(in[0]), .Y(n36) );
  INVX0_HVT U299 ( .A(n116), .Y(n164) );
  INVX0_HVT U300 ( .A(n301), .Y(n9) );
  NAND2X0_HVT U301 ( .A1(n35), .A2(n148), .Y(n301) );
  NAND2X0_HVT U302 ( .A1(n273), .A2(n121), .Y(n148) );
  AO221X1_HVT U303 ( .A1(n16), .A2(n48), .A3(n279), .A4(n15), .A5(n343), .Y(
        n340) );
  AO21X1_HVT U304 ( .A1(n344), .A2(n12), .A3(n88), .Y(n343) );
  AND2X1_HVT U305 ( .A1(n61), .A2(n10), .Y(n88) );
  INVX0_HVT U306 ( .A(n123), .Y(n61) );
  NAND2X0_HVT U307 ( .A1(n122), .A2(in[0]), .Y(n123) );
  INVX0_HVT U308 ( .A(n159), .Y(n122) );
  INVX0_HVT U309 ( .A(n309), .Y(n344) );
  NAND2X0_HVT U310 ( .A1(n21), .A2(n314), .Y(n309) );
  INVX0_HVT U311 ( .A(n175), .Y(n279) );
  NAND2X0_HVT U312 ( .A1(n35), .A2(n314), .Y(n175) );
  NAND2X0_HVT U313 ( .A1(n159), .A2(n121), .Y(n314) );
  NAND2X0_HVT U314 ( .A1(in[0]), .A2(n58), .Y(n35) );
  NAND2X0_HVT U315 ( .A1(n58), .A2(n121), .Y(n48) );
  AND2X1_HVT U316 ( .A1(in[5]), .A2(n8), .Y(n83) );
  AO221X1_HVT U317 ( .A1(n16), .A2(n329), .A3(n287), .A4(n15), .A5(n345), .Y(
        n338) );
  AO221X1_HVT U318 ( .A1(n265), .A2(n10), .A3(n218), .A4(n12), .A5(n23), .Y(
        n345) );
  INVX0_HVT U319 ( .A(n161), .Y(n23) );
  NAND2X0_HVT U320 ( .A1(n16), .A2(n121), .Y(n161) );
  INVX0_HVT U321 ( .A(n317), .Y(n265) );
  NAND2X0_HVT U322 ( .A1(n47), .A2(n212), .Y(n317) );
  NAND2X0_HVT U323 ( .A1(in[0]), .A2(n57), .Y(n47) );
  AND2X1_HVT U324 ( .A1(n89), .A2(n212), .Y(n287) );
  NAND2X0_HVT U325 ( .A1(in[6]), .A2(n121), .Y(n212) );
  INVX0_HVT U326 ( .A(in[0]), .Y(n121) );
  NAND2X0_HVT U327 ( .A1(in[0]), .A2(n159), .Y(n89) );
  AND2X1_HVT U328 ( .A1(in[1]), .A2(n5), .Y(n78) );
  AO221X1_HVT U329 ( .A1(n16), .A2(n57), .A3(n332), .A4(n15), .A5(n346), .Y(
        n337) );
  AO22X1_HVT U330 ( .A1(n218), .A2(n12), .A3(n10), .A4(in[3]), .Y(n346) );
  INVX0_HVT U331 ( .A(n44), .Y(n10) );
  NAND2X0_HVT U332 ( .A1(in[2]), .A2(n186), .Y(n44) );
  INVX0_HVT U333 ( .A(n37), .Y(n12) );
  NAND2X0_HVT U334 ( .A1(n95), .A2(n186), .Y(n37) );
  INVX0_HVT U335 ( .A(in[4]), .Y(n186) );
  OA21X1_HVT U336 ( .A1(n185), .A2(in[0]), .A3(n21), .Y(n218) );
  NAND2X0_HVT U337 ( .A1(in[0]), .A2(n116), .Y(n21) );
  INVX0_HVT U338 ( .A(n57), .Y(n185) );
  INVX0_HVT U339 ( .A(n56), .Y(n15) );
  NAND2X0_HVT U340 ( .A1(in[4]), .A2(n95), .Y(n56) );
  INVX0_HVT U341 ( .A(in[2]), .Y(n95) );
  INVX0_HVT U342 ( .A(n188), .Y(n332) );
  NAND2X0_HVT U343 ( .A1(in[0]), .A2(n273), .Y(n188) );
  NAND2X0_HVT U344 ( .A1(n116), .A2(n159), .Y(n273) );
  NAND2X0_HVT U345 ( .A1(in[6]), .A2(in[3]), .Y(n159) );
  NAND2X0_HVT U346 ( .A1(n329), .A2(n58), .Y(n116) );
  INVX0_HVT U347 ( .A(in[3]), .Y(n58) );
  NAND2X0_HVT U348 ( .A1(in[3]), .A2(n329), .Y(n57) );
  INVX0_HVT U349 ( .A(in[6]), .Y(n329) );
  INVX0_HVT U350 ( .A(n50), .Y(n16) );
  NAND2X0_HVT U351 ( .A1(in[2]), .A2(in[4]), .Y(n50) );
  AND2X1_HVT U352 ( .A1(n8), .A2(n5), .Y(n76) );
  INVX0_HVT U353 ( .A(in[5]), .Y(n5) );
  INVX0_HVT U354 ( .A(in[1]), .Y(n8) );
endmodule

