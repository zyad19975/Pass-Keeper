
module sbox_11 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n210, n211, n212, n213, n216, n217, n218, n219, n224, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609;

  NAND2X0_HVT U4 ( .A1(n315), .A2(n237), .Y(n606) );
  NAND2X0_HVT U5 ( .A1(n321), .A2(n387), .Y(n604) );
  NAND2X0_HVT U13 ( .A1(n596), .A2(n318), .Y(n597) );
  NAND2X0_HVT U15 ( .A1(n236), .A2(n306), .Y(n594) );
  NAND2X0_HVT U21 ( .A1(n315), .A2(n325), .Y(n588) );
  NAND2X0_HVT U24 ( .A1(n270), .A2(n325), .Y(n586) );
  NAND2X0_HVT U33 ( .A1(n385), .A2(n325), .Y(n577) );
  NAND2X0_HVT U42 ( .A1(n323), .A2(n311), .Y(n568) );
  MUX41X1_HVT U51 ( .A1(n374), .A3(n335), .A2(n351), .A4(n352), .S0(n265), 
        .S1(n328), .Y(n560) );
  NAND2X0_HVT U53 ( .A1(n557), .A2(n567), .Y(n558) );
  NAND2X0_HVT U56 ( .A1(n315), .A2(n553), .Y(n554) );
  MUX41X1_HVT U57 ( .A1(n375), .A3(n590), .A2(n554), .A4(n599), .S0(n265), 
        .S1(n328), .Y(n552) );
  NAND2X0_HVT U58 ( .A1(n318), .A2(n236), .Y(n551) );
  MUX41X1_HVT U59 ( .A1(n298), .A3(n551), .A2(n296), .A4(n350), .S0(n266), 
        .S1(n328), .Y(n550) );
  MUX41X1_HVT U61 ( .A1(n295), .A3(n349), .A2(n348), .A4(n306), .S0(n266), 
        .S1(n329), .Y(n548) );
  NAND2X0_HVT U62 ( .A1(n325), .A2(n608), .Y(n547) );
  MUX41X1_HVT U63 ( .A1(n547), .A3(n341), .A2(n369), .A4(n347), .S0(n266), 
        .S1(n301), .Y(n546) );
  AO21X1_HVT U66 ( .A1(n253), .A2(in[5]), .A3(n232), .Y(n543) );
  MUX41X1_HVT U68 ( .A1(n344), .A3(n543), .A2(n542), .A4(n544), .S0(n299), 
        .S1(n265), .Y(n541) );
  MUX41X1_HVT U69 ( .A1(n541), .A3(n549), .A2(n545), .A4(n555), .S0(in[6]), 
        .S1(n271), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n313), .A2(n536), .Y(n537) );
  MUX41X1_HVT U74 ( .A1(n538), .A3(n584), .A2(n537), .A4(n586), .S0(n280), 
        .S1(n331), .Y(n535) );
  MUX41X1_HVT U77 ( .A1(n601), .A3(n378), .A2(n533), .A4(n269), .S0(n302), 
        .S1(n326), .Y(n532) );
  MUX41X1_HVT U78 ( .A1(n532), .A3(n535), .A2(n534), .A4(n539), .S0(n310), 
        .S1(n328), .Y(n531) );
  AND3X1_HVT U80 ( .A1(n317), .A2(n553), .A3(n528), .Y(n529) );
  MUX41X1_HVT U82 ( .A1(n565), .A3(n352), .A2(n336), .A4(n595), .S0(n299), 
        .S1(n332), .Y(n526) );
  AND2X1_HVT U83 ( .A1(n322), .A2(n256), .Y(n525) );
  MUX41X1_HVT U84 ( .A1(n353), .A3(n603), .A2(n593), .A4(n525), .S0(n299), 
        .S1(n265), .Y(n524) );
  NAND2X0_HVT U85 ( .A1(n325), .A2(n388), .Y(n523) );
  MUX41X1_HVT U90 ( .A1(n564), .A3(n568), .A2(n374), .A4(n520), .S0(n300), 
        .S1(n303), .Y(n519) );
  AO21X1_HVT U93 ( .A1(n304), .A2(n515), .A3(n373), .Y(n516) );
  MUX41X1_HVT U96 ( .A1(n336), .A3(n294), .A2(n376), .A4(n513), .S0(n299), 
        .S1(n265), .Y(n512) );
  MUX41X1_HVT U97 ( .A1(n372), .A3(n294), .A2(n216), .A4(n594), .S0(n299), 
        .S1(n330), .Y(n511) );
  MUX41X1_HVT U98 ( .A1(n511), .A3(n514), .A2(n512), .A4(n519), .S0(n310), 
        .S1(n328), .Y(n510) );
  NAND2X0_HVT U101 ( .A1(n506), .A2(n505), .Y(n507) );
  MUX41X1_HVT U103 ( .A1(n237), .A3(n345), .A2(n357), .A4(n575), .S0(n299), 
        .S1(n266), .Y(n503) );
  MUX41X1_HVT U105 ( .A1(n356), .A3(n563), .A2(n502), .A4(n371), .S0(n299), 
        .S1(n265), .Y(n501) );
  OA21X1_HVT U109 ( .A1(n276), .A2(n251), .A3(n350), .Y(n498) );
  NAND2X0_HVT U110 ( .A1(n317), .A2(n496), .Y(n497) );
  MUX41X1_HVT U114 ( .A1(n493), .A3(n499), .A2(n495), .A4(n498), .S0(in[5]), 
        .S1(n331), .Y(n492) );
  AND2X1_HVT U115 ( .A1(n320), .A2(n307), .Y(n491) );
  MUX41X1_HVT U116 ( .A1(n263), .A3(n491), .A2(n354), .A4(n579), .S0(n300), 
        .S1(n331), .Y(n490) );
  AO21X1_HVT U118 ( .A1(n242), .A2(n312), .A3(n603), .Y(n488) );
  NAND2X0_HVT U123 ( .A1(n482), .A2(n481), .Y(n483) );
  MUX41X1_HVT U125 ( .A1(n588), .A3(n298), .A2(n344), .A4(n380), .S0(n300), 
        .S1(n266), .Y(n479) );
  MUX41X1_HVT U131 ( .A1(n474), .A3(n476), .A2(n475), .A4(n477), .S0(in[5]), 
        .S1(n265), .Y(n473) );
  MUX41X1_HVT U135 ( .A1(n381), .A3(n386), .A2(n604), .A4(n583), .S0(n280), 
        .S1(n332), .Y(n470) );
  MUX41X1_HVT U136 ( .A1(n291), .A3(n577), .A2(n382), .A4(n574), .S0(n300), 
        .S1(n331), .Y(n469) );
  MUX41X1_HVT U139 ( .A1(n467), .A3(n470), .A2(n469), .A4(n471), .S0(n310), 
        .S1(n328), .Y(n466) );
  AND2X1_HVT U140 ( .A1(n312), .A2(n325), .Y(n465) );
  OA21X1_HVT U144 ( .A1(n338), .A2(n333), .A3(n579), .Y(n461) );
  MUX41X1_HVT U147 ( .A1(n382), .A3(n536), .A2(n372), .A4(n564), .S0(n280), 
        .S1(n331), .Y(n459) );
  OA21X1_HVT U151 ( .A1(n570), .A2(n333), .A3(n455), .Y(n456) );
  MUX41X1_HVT U153 ( .A1(n497), .A3(n295), .A2(n316), .A4(n23), .S0(n300), 
        .S1(n331), .Y(n453) );
  AND2X1_HVT U154 ( .A1(n304), .A2(n270), .Y(n452) );
  NAND2X0_HVT U158 ( .A1(n323), .A2(n388), .Y(n448) );
  MUX41X1_HVT U159 ( .A1(n263), .A3(n306), .A2(n448), .A4(n343), .S0(n327), 
        .S1(n266), .Y(n447) );
  MUX41X1_HVT U160 ( .A1(n447), .A3(n453), .A2(n449), .A4(n454), .S0(n310), 
        .S1(n301), .Y(n446) );
  AND2X1_HVT U162 ( .A1(n603), .A2(n536), .Y(n444) );
  MUX41X1_HVT U163 ( .A1(n349), .A3(n444), .A2(n292), .A4(n445), .S0(n212), 
        .S1(n304), .Y(n443) );
  MUX41X1_HVT U165 ( .A1(n588), .A3(n358), .A2(n564), .A4(n442), .S0(n331), 
        .S1(n326), .Y(n441) );
  NAND2X0_HVT U166 ( .A1(n318), .A2(n553), .Y(n440) );
  NAND2X0_HVT U167 ( .A1(n389), .A2(n325), .Y(n439) );
  MUX41X1_HVT U168 ( .A1(n375), .A3(n312), .A2(n439), .A4(n440), .S0(n212), 
        .S1(n330), .Y(n438) );
  OA21X1_HVT U170 ( .A1(n296), .A2(n333), .A3(n579), .Y(n436) );
  MUX41X1_HVT U172 ( .A1(n435), .A3(n441), .A2(n438), .A4(n443), .S0(in[0]), 
        .S1(n328), .Y(n434) );
  NAND2X0_HVT U174 ( .A1(n319), .A2(n603), .Y(n596) );
  NAND2X0_HVT U177 ( .A1(n320), .A2(n309), .Y(n431) );
  MUX41X1_HVT U178 ( .A1(n592), .A3(n431), .A2(n383), .A4(n572), .S0(n242), 
        .S1(n331), .Y(n430) );
  MUX41X1_HVT U179 ( .A1(n582), .A3(n384), .A2(n339), .A4(n383), .S0(n212), 
        .S1(n265), .Y(n429) );
  MUX41X1_HVT U181 ( .A1(n428), .A3(n430), .A2(n429), .A4(n432), .S0(n310), 
        .S1(n301), .Y(n427) );
  MUX41X1_HVT U182 ( .A1(n365), .A3(n314), .A2(n367), .A4(n355), .S0(n331), 
        .S1(n327), .Y(n426) );
  OA21X1_HVT U184 ( .A1(n576), .A2(n333), .A3(n353), .Y(n424) );
  MUX41X1_HVT U189 ( .A1(n420), .A3(n596), .A2(n421), .A4(n371), .S0(n302), 
        .S1(n327), .Y(n419) );
  MUX41X1_HVT U194 ( .A1(n569), .A3(n583), .A2(n381), .A4(n312), .S0(n302), 
        .S1(n327), .Y(n415) );
  MUX41X1_HVT U195 ( .A1(n603), .A3(n376), .A2(n609), .A4(n573), .S0(n212), 
        .S1(n265), .Y(n414) );
  AO21X1_HVT U197 ( .A1(n293), .A2(n303), .A3(n373), .Y(n412) );
  MUX41X1_HVT U203 ( .A1(n574), .A3(n366), .A2(n598), .A4(n578), .S0(n327), 
        .S1(n303), .Y(n406) );
  MUX41X1_HVT U204 ( .A1(n554), .A3(n597), .A2(n362), .A4(n587), .S0(n212), 
        .S1(n266), .Y(n405) );
  MUX41X1_HVT U205 ( .A1(n256), .A3(n237), .A2(n384), .A4(n360), .S0(n327), 
        .S1(n266), .Y(n404) );
  MUX41X1_HVT U206 ( .A1(n404), .A3(n406), .A2(n405), .A4(n407), .S0(n310), 
        .S1(n301), .Y(n403) );
  NAND2X0_HVT U208 ( .A1(n319), .A2(n315), .Y(n496) );
  NAND2X0_HVT U212 ( .A1(n319), .A2(n313), .Y(n553) );
  NAND2X0_HVT U214 ( .A1(n603), .A2(n325), .Y(n402) );
  NAND2X0_HVT U215 ( .A1(n496), .A2(n313), .Y(n401) );
  AO21X1_HVT U216 ( .A1(n325), .A2(n386), .A3(n333), .Y(n506) );
  NAND2X0_HVT U218 ( .A1(n386), .A2(n217), .Y(n455) );
  NAND2X0_HVT U220 ( .A1(n303), .A2(n402), .Y(n528) );
  NOR2X1_HVT U1 ( .A1(n48), .A2(in[1]), .Y(n23) );
  IBUFFX4_HVT U2 ( .A(n23), .Y(n575) );
  IBUFFX16_HVT U3 ( .A(n309), .Y(n48) );
  MUX21X2_HVT U6 ( .A1(n560), .A2(n556), .S0(n210), .Y(n555) );
  IBUFFX16_HVT U7 ( .A(n264), .Y(n210) );
  INVX1_HVT U8 ( .A(n326), .Y(n211) );
  INVX2_HVT U9 ( .A(n211), .Y(n212) );
  MUX41X1_HVT U10 ( .A1(n433), .A3(n308), .A2(n596), .A4(n379), .S0(n213), 
        .S1(n326), .Y(n432) );
  IBUFFX16_HVT U11 ( .A(n266), .Y(n213) );
  INVX2_HVT U12 ( .A(in[1]), .Y(n325) );
  INVX1_HVT U14 ( .A(n324), .Y(n216) );
  INVX1_HVT U16 ( .A(n324), .Y(n217) );
  INVX1_HVT U17 ( .A(n324), .Y(n319) );
  MUX21X1_HVT U18 ( .A1(n572), .A2(n378), .S0(n302), .Y(n450) );
  INVX2_HVT U19 ( .A(n324), .Y(n323) );
  MUX21X1_HVT U20 ( .A1(n385), .A2(n311), .S0(n324), .Y(n571) );
  IBUFFX2_HVT U22 ( .A(n324), .Y(n320) );
  MUX41X1_HVT U23 ( .A1(n526), .A3(n522), .A2(n527), .A4(n524), .S0(n285), 
        .S1(n218), .Y(n521) );
  IBUFFX16_HVT U25 ( .A(n275), .Y(n218) );
  MUX21X1_HVT U26 ( .A1(n589), .A2(n600), .S0(in[7]), .Y(n530) );
  NAND2X0_HVT U27 ( .A1(n521), .A2(n219), .Y(n224) );
  NAND2X0_HVT U28 ( .A1(n531), .A2(in[6]), .Y(n231) );
  NAND2X2_HVT U29 ( .A1(n224), .A2(n231), .Y(out[1]) );
  IBUFFX2_HVT U30 ( .A(in[6]), .Y(n219) );
  INVX2_HVT U31 ( .A(in[7]), .Y(n333) );
  NOR2X2_HVT U32 ( .A1(n325), .A2(n233), .Y(n232) );
  INVX8_HVT U34 ( .A(n232), .Y(n536) );
  IBUFFX16_HVT U35 ( .A(n318), .Y(n233) );
  INVX2_HVT U36 ( .A(in[1]), .Y(n324) );
  MUX21X2_HVT U37 ( .A1(n487), .A2(n490), .S0(n329), .Y(n486) );
  MUX21X2_HVT U38 ( .A1(n530), .A2(n529), .S0(n300), .Y(n527) );
  MUX41X1_HVT U39 ( .A1(n564), .A3(n536), .A2(n571), .A4(n294), .S0(n234), 
        .S1(n235), .Y(n422) );
  IBUFFX16_HVT U40 ( .A(n327), .Y(n234) );
  IBUFFX16_HVT U41 ( .A(n332), .Y(n235) );
  IBUFFX2_HVT U43 ( .A(n571), .Y(n365) );
  INVX1_HVT U44 ( .A(n324), .Y(n322) );
  NBUFFX2_HVT U45 ( .A(n607), .Y(n236) );
  NBUFFX2_HVT U46 ( .A(n607), .Y(n237) );
  NBUFFX2_HVT U47 ( .A(n605), .Y(n314) );
  INVX0_HVT U48 ( .A(n334), .Y(n332) );
  INVX1_HVT U49 ( .A(n316), .Y(n389) );
  MUX21X1_HVT U50 ( .A1(n359), .A2(n472), .S0(n280), .Y(n471) );
  INVX0_HVT U52 ( .A(n313), .Y(n260) );
  NAND2X0_HVT U54 ( .A1(n322), .A2(n317), .Y(n607) );
  INVX0_HVT U55 ( .A(n315), .Y(n277) );
  INVX0_HVT U60 ( .A(n585), .Y(n354) );
  NAND2X0_HVT U64 ( .A1(n248), .A2(n249), .Y(out[2]) );
  INVX0_HVT U65 ( .A(n587), .Y(n353) );
  INVX0_HVT U67 ( .A(n372), .Y(n262) );
  INVX1_HVT U70 ( .A(n283), .Y(n327) );
  INVX1_HVT U71 ( .A(n251), .Y(n326) );
  MUX21X1_HVT U72 ( .A1(n606), .A2(n468), .S0(n283), .Y(n467) );
  INVX1_HVT U75 ( .A(n299), .Y(n251) );
  INVX0_HVT U76 ( .A(n251), .Y(n264) );
  INVX1_HVT U79 ( .A(n324), .Y(n321) );
  NBUFFX2_HVT U81 ( .A(n284), .Y(n307) );
  INVX0_HVT U86 ( .A(n580), .Y(n358) );
  INVX1_HVT U87 ( .A(n305), .Y(n270) );
  INVX1_HVT U88 ( .A(in[3]), .Y(n387) );
  INVX1_HVT U89 ( .A(n266), .Y(n252) );
  INVX0_HVT U91 ( .A(in[6]), .Y(n286) );
  INVX1_HVT U92 ( .A(n285), .Y(n271) );
  INVX1_HVT U94 ( .A(in[2]), .Y(n283) );
  INVX0_HVT U95 ( .A(in[5]), .Y(n275) );
  MUX21X1_HVT U99 ( .A1(n389), .A2(n603), .S0(n325), .Y(n585) );
  INVX0_HVT U100 ( .A(n589), .Y(n352) );
  XOR2X2_HVT U102 ( .A1(n284), .A2(n279), .Y(n564) );
  MUX21X2_HVT U104 ( .A1(n593), .A2(n290), .S0(n302), .Y(n409) );
  NAND2X0_HVT U106 ( .A1(n246), .A2(n247), .Y(out[4]) );
  INVX1_HVT U107 ( .A(n261), .Y(n534) );
  NAND2X0_HVT U108 ( .A1(n479), .A2(n275), .Y(n238) );
  NAND2X0_HVT U111 ( .A1(n480), .A2(n328), .Y(n239) );
  NAND2X0_HVT U112 ( .A1(n238), .A2(n239), .Y(n478) );
  MUX21X1_HVT U113 ( .A1(n484), .A2(n483), .S0(n304), .Y(n480) );
  NAND2X0_HVT U117 ( .A1(n356), .A2(n251), .Y(n240) );
  NAND2X0_HVT U119 ( .A1(n580), .A2(n299), .Y(n241) );
  NAND2X0_HVT U120 ( .A1(n240), .A2(n241), .Y(n477) );
  NAND2X0_HVT U121 ( .A1(n552), .A2(n242), .Y(n243) );
  NAND2X0_HVT U122 ( .A1(n550), .A2(n283), .Y(n244) );
  NAND2X0_HVT U124 ( .A1(n243), .A2(n244), .Y(n549) );
  INVX0_HVT U126 ( .A(n283), .Y(n242) );
  NAND2X0_HVT U127 ( .A1(n466), .A2(n245), .Y(n246) );
  NAND2X0_HVT U128 ( .A1(n458), .A2(n286), .Y(n247) );
  INVX1_HVT U129 ( .A(n286), .Y(n245) );
  MUX21X2_HVT U130 ( .A1(n595), .A2(n360), .S0(n283), .Y(n509) );
  NAND2X0_HVT U132 ( .A1(n510), .A2(n245), .Y(n248) );
  NAND2X0_HVT U133 ( .A1(n500), .A2(n286), .Y(n249) );
  IBUFFX2_HVT U134 ( .A(n595), .Y(n347) );
  INVX1_HVT U137 ( .A(n253), .Y(n599) );
  INVX1_HVT U138 ( .A(n276), .Y(n573) );
  MUX21X2_HVT U141 ( .A1(n295), .A2(n509), .S0(n250), .Y(n508) );
  XOR2X1_HVT U142 ( .A1(n251), .A2(n333), .Y(n250) );
  MUX41X1_HVT U143 ( .A1(n291), .A3(n293), .A2(n523), .A4(n377), .S0(n251), 
        .S1(n252), .Y(n522) );
  MUX21X1_HVT U145 ( .A1(n270), .A2(n609), .S0(n216), .Y(n253) );
  NAND2X0_HVT U146 ( .A1(n456), .A2(n283), .Y(n254) );
  NAND2X0_HVT U148 ( .A1(n457), .A2(n264), .Y(n255) );
  NAND2X0_HVT U149 ( .A1(n254), .A2(n255), .Y(n454) );
  MUX21X1_HVT U150 ( .A1(n269), .A2(n386), .S0(n303), .Y(n457) );
  MUX21X2_HVT U152 ( .A1(n566), .A2(n540), .S0(n280), .Y(n539) );
  MUX21X1_HVT U155 ( .A1(n307), .A2(n270), .S0(n319), .Y(n587) );
  INVX0_HVT U156 ( .A(n321), .Y(n279) );
  MUX21X1_HVT U157 ( .A1(n389), .A2(n388), .S0(n216), .Y(n583) );
  MUX21X2_HVT U161 ( .A1(n337), .A2(n485), .S0(n242), .Y(n484) );
  IBUFFX2_HVT U164 ( .A(n390), .Y(n256) );
  INVX1_HVT U169 ( .A(in[4]), .Y(n390) );
  INVX1_HVT U171 ( .A(n399), .Y(n375) );
  MUX21X2_HVT U173 ( .A1(n450), .A2(n451), .S0(n264), .Y(n449) );
  MUX21X2_HVT U175 ( .A1(n581), .A2(n340), .S0(n304), .Y(n462) );
  MUX21X2_HVT U176 ( .A1(n365), .A2(n587), .S0(n333), .Y(n468) );
  MUX21X2_HVT U180 ( .A1(n462), .A2(n461), .S0(n264), .Y(n460) );
  NAND2X0_HVT U183 ( .A1(n408), .A2(n283), .Y(n257) );
  NAND2X0_HVT U185 ( .A1(n409), .A2(n264), .Y(n258) );
  NAND2X0_HVT U186 ( .A1(n257), .A2(n258), .Y(n407) );
  INVX0_HVT U187 ( .A(n593), .Y(n348) );
  MUX21X1_HVT U188 ( .A1(n306), .A2(n305), .S0(n322), .Y(n593) );
  MUX41X1_HVT U190 ( .A1(n263), .A3(n290), .A2(n342), .A4(n601), .S0(n302), 
        .S1(n283), .Y(n428) );
  INVX0_HVT U191 ( .A(n395), .Y(n380) );
  INVX1_HVT U192 ( .A(n259), .Y(n472) );
  MUX21X1_HVT U193 ( .A1(n260), .A2(n395), .S0(n333), .Y(n259) );
  MUX41X1_HVT U196 ( .A1(n460), .A3(n464), .A2(n459), .A4(n463), .S0(in[0]), 
        .S1(n275), .Y(n458) );
  MUX41X1_HVT U198 ( .A1(n585), .A3(n608), .A2(n397), .A4(n262), .S0(n251), 
        .S1(n252), .Y(n261) );
  MUX21X1_HVT U199 ( .A1(n284), .A2(n277), .S0(n278), .Y(n276) );
  INVX0_HVT U200 ( .A(n217), .Y(n278) );
  NAND2X0_HVT U201 ( .A1(n403), .A2(n286), .Y(n267) );
  OA21X1_HVT U202 ( .A1(n602), .A2(n333), .A3(n364), .Y(n408) );
  INVX1_HVT U207 ( .A(n369), .Y(n263) );
  MUX41X1_HVT U209 ( .A1(n585), .A3(n364), .A2(n465), .A4(n361), .S0(n264), 
        .S1(in[7]), .Y(n464) );
  XOR2X2_HVT U210 ( .A1(n583), .A2(n333), .Y(n566) );
  INVX2_HVT U211 ( .A(n334), .Y(n265) );
  INVX2_HVT U213 ( .A(n334), .Y(n266) );
  MUX41X1_HVT U217 ( .A1(n411), .A3(n414), .A2(n415), .A4(n416), .S0(n301), 
        .S1(n271), .Y(n410) );
  NAND2X0_HVT U219 ( .A1(n410), .A2(in[6]), .Y(n268) );
  NAND2X0_HVT U221 ( .A1(n267), .A2(n268), .Y(out[7]) );
  MUX41X1_HVT U222 ( .A1(n568), .A3(n575), .A2(n561), .A4(n417), .S0(n327), 
        .S1(n302), .Y(n416) );
  MUX21X1_HVT U223 ( .A1(n270), .A2(n284), .S0(n217), .Y(n269) );
  MUX21X2_HVT U224 ( .A1(n413), .A2(n412), .S0(n264), .Y(n411) );
  NAND2X0_HVT U225 ( .A1(n317), .A2(n272), .Y(n273) );
  NAND2X0_HVT U226 ( .A1(n518), .A2(n297), .Y(n274) );
  NAND2X0_HVT U227 ( .A1(n273), .A2(n274), .Y(n517) );
  INVX0_HVT U228 ( .A(n297), .Y(n272) );
  MUX21X2_HVT U229 ( .A1(n517), .A2(n516), .S0(n283), .Y(n514) );
  INVX2_HVT U230 ( .A(in[7]), .Y(n334) );
  INVX1_HVT U231 ( .A(n284), .Y(n603) );
  MUX21X2_HVT U232 ( .A1(n434), .A2(n446), .S0(in[6]), .Y(out[5]) );
  AND3X2_HVT U233 ( .A1(n242), .A2(n325), .A3(n256), .Y(n476) );
  NAND2X0_HVT U234 ( .A1(n548), .A2(n280), .Y(n281) );
  NAND2X0_HVT U235 ( .A1(n546), .A2(n283), .Y(n282) );
  NAND2X0_HVT U236 ( .A1(n281), .A2(n282), .Y(n545) );
  INVX0_HVT U237 ( .A(n283), .Y(n280) );
  IBUFFX4_HVT U238 ( .A(n334), .Y(n330) );
  INVX2_HVT U239 ( .A(n334), .Y(n331) );
  INVX1_HVT U240 ( .A(in[0]), .Y(n285) );
  XNOR2X2_HVT U241 ( .A1(n308), .A2(in[3]), .Y(n284) );
  MUX41X1_HVT U242 ( .A1(n312), .A3(n370), .A2(n284), .A4(n353), .S0(n251), 
        .S1(n333), .Y(n463) );
  MUX41X1_HVT U243 ( .A1(n508), .A3(n503), .A2(n504), .A4(n501), .S0(n285), 
        .S1(n275), .Y(n500) );
  MUX41X1_HVT U244 ( .A1(n423), .A3(n426), .A2(n419), .A4(n422), .S0(n301), 
        .S1(n285), .Y(n418) );
  MUX41X1_HVT U245 ( .A1(n492), .A3(n478), .A2(n486), .A4(n473), .S0(n286), 
        .S1(n285), .Y(out[3]) );
  MUX21X2_HVT U246 ( .A1(n418), .A2(n427), .S0(in[6]), .Y(out[6]) );
  NAND2X0_HVT U247 ( .A1(n494), .A2(n287), .Y(n288) );
  NAND2X0_HVT U248 ( .A1(n608), .A2(n562), .Y(n289) );
  NAND2X0_HVT U249 ( .A1(n288), .A2(n289), .Y(n493) );
  INVX0_HVT U250 ( .A(n562), .Y(n287) );
  XOR2X1_HVT U251 ( .A1(n319), .A2(in[2]), .Y(n562) );
  NBUFFX16_HVT U252 ( .A(n329), .Y(n301) );
  INVX1_HVT U253 ( .A(n314), .Y(n385) );
  NBUFFX2_HVT U254 ( .A(n284), .Y(n306) );
  MUX21X1_HVT U255 ( .A1(n292), .A2(n348), .S0(n300), .Y(n475) );
  AND2X1_HVT U256 ( .A1(n307), .A2(n553), .Y(n290) );
  MUX21X1_HVT U257 ( .A1(n385), .A2(n388), .S0(n329), .Y(n557) );
  NBUFFX2_HVT U258 ( .A(n605), .Y(n315) );
  MUX21X1_HVT U259 ( .A1(n345), .A2(n386), .S0(in[5]), .Y(n542) );
  MUX21X1_HVT U260 ( .A1(n579), .A2(n497), .S0(n300), .Y(n495) );
  AND2X1_HVT U261 ( .A1(n317), .A2(n536), .Y(n291) );
  MUX21X1_HVT U262 ( .A1(n307), .A2(n388), .S0(n216), .Y(n602) );
  MUX21X1_HVT U263 ( .A1(n317), .A2(n306), .S0(n321), .Y(n569) );
  MUX21X1_HVT U264 ( .A1(n306), .A2(n309), .S0(n323), .Y(n505) );
  MUX21X1_HVT U265 ( .A1(n385), .A2(n389), .S0(n323), .Y(n433) );
  MUX21X1_HVT U266 ( .A1(n306), .A2(n385), .S0(n217), .Y(n513) );
  MUX21X1_HVT U267 ( .A1(n388), .A2(n385), .S0(n321), .Y(n572) );
  MUX21X1_HVT U268 ( .A1(n305), .A2(n389), .S0(n320), .Y(n570) );
  MUX21X1_HVT U269 ( .A1(n388), .A2(n306), .S0(n321), .Y(n445) );
  NAND2X0_HVT U270 ( .A1(n308), .A2(n387), .Y(n605) );
  MUX21X1_HVT U271 ( .A1(n603), .A2(n386), .S0(n216), .Y(n394) );
  NBUFFX2_HVT U272 ( .A(n608), .Y(n316) );
  MUX21X1_HVT U273 ( .A1(n315), .A2(n313), .S0(n321), .Y(n520) );
  MUX21X1_HVT U274 ( .A1(n603), .A2(n309), .S0(n323), .Y(n533) );
  INVX1_HVT U275 ( .A(n312), .Y(n386) );
  INVX1_HVT U276 ( .A(n609), .Y(n388) );
  MUX21X1_HVT U277 ( .A1(n388), .A2(n305), .S0(n322), .Y(n576) );
  MUX21X1_HVT U278 ( .A1(n309), .A2(n385), .S0(n320), .Y(n581) );
  MUX21X1_HVT U279 ( .A1(n488), .A2(n489), .S0(n303), .Y(n487) );
  MUX21X1_HVT U280 ( .A1(n23), .A2(n362), .S0(n300), .Y(n489) );
  NBUFFX2_HVT U281 ( .A(n608), .Y(n317) );
  MUX21X1_HVT U282 ( .A1(n305), .A2(n309), .S0(n217), .Y(n417) );
  XOR2X1_HVT U283 ( .A1(n316), .A2(n322), .Y(n561) );
  MUX21X1_HVT U284 ( .A1(n385), .A2(n309), .S0(n322), .Y(n395) );
  MUX21X1_HVT U285 ( .A1(n317), .A2(n313), .S0(n323), .Y(n595) );
  MUX21X1_HVT U286 ( .A1(n314), .A2(n318), .S0(n319), .Y(n515) );
  MUX21X1_HVT U287 ( .A1(n315), .A2(n305), .S0(n323), .Y(n598) );
  MUX21X1_HVT U288 ( .A1(n386), .A2(n385), .S0(n322), .Y(n591) );
  MUX21X1_HVT U289 ( .A1(n309), .A2(n305), .S0(n323), .Y(n485) );
  MUX21X1_HVT U290 ( .A1(n305), .A2(n318), .S0(n216), .Y(n420) );
  MUX21X1_HVT U291 ( .A1(n609), .A2(n317), .S0(n216), .Y(n421) );
  XOR2X1_HVT U292 ( .A1(n217), .A2(n386), .Y(n565) );
  MUX21X1_HVT U293 ( .A1(n609), .A2(n313), .S0(n217), .Y(n579) );
  MUX21X1_HVT U294 ( .A1(n316), .A2(n309), .S0(n319), .Y(n400) );
  XNOR2X1_HVT U295 ( .A1(n314), .A2(n321), .Y(n292) );
  XNOR2X1_HVT U296 ( .A1(n609), .A2(n322), .Y(n293) );
  AND2X1_HVT U297 ( .A1(n217), .A2(n389), .Y(n294) );
  MUX21X1_HVT U298 ( .A1(n313), .A2(n305), .S0(n320), .Y(n398) );
  MUX21X1_HVT U299 ( .A1(n316), .A2(n315), .S0(n321), .Y(n393) );
  AND2X1_HVT U300 ( .A1(n318), .A2(n496), .Y(n295) );
  MUX21X1_HVT U301 ( .A1(n313), .A2(n309), .S0(n320), .Y(n538) );
  MUX21X1_HVT U302 ( .A1(n600), .A2(n318), .S0(n280), .Y(n482) );
  XOR2X1_HVT U303 ( .A1(n308), .A2(n323), .Y(n584) );
  NBUFFX2_HVT U304 ( .A(n332), .Y(n303) );
  NBUFFX2_HVT U305 ( .A(n332), .Y(n302) );
  NBUFFX2_HVT U306 ( .A(n332), .Y(n304) );
  NBUFFX2_HVT U307 ( .A(n387), .Y(n305) );
  NBUFFX2_HVT U308 ( .A(in[2]), .Y(n300) );
  NBUFFX2_HVT U309 ( .A(in[2]), .Y(n299) );
  NBUFFX2_HVT U310 ( .A(n390), .Y(n308) );
  MUX21X1_HVT U311 ( .A1(n507), .A2(n359), .S0(n242), .Y(n504) );
  MUX21X1_HVT U312 ( .A1(n424), .A2(n425), .S0(n299), .Y(n423) );
  MUX21X1_HVT U313 ( .A1(n523), .A2(n311), .S0(n303), .Y(n425) );
  XOR2X1_HVT U314 ( .A1(n320), .A2(n270), .Y(n563) );
  MUX21X1_HVT U315 ( .A1(n313), .A2(n307), .S0(n320), .Y(n502) );
  NAND2X0_HVT U316 ( .A1(n311), .A2(n390), .Y(n608) );
  MUX21X1_HVT U317 ( .A1(n437), .A2(n436), .S0(n242), .Y(n435) );
  MUX21X1_HVT U318 ( .A1(n313), .A2(n376), .S0(n304), .Y(n437) );
  AND2X1_HVT U319 ( .A1(n307), .A2(n325), .Y(n296) );
  NBUFFX2_HVT U320 ( .A(n600), .Y(n312) );
  MUX21X1_HVT U321 ( .A1(n388), .A2(n376), .S0(n304), .Y(n540) );
  MUX21X1_HVT U322 ( .A1(n592), .A2(n361), .S0(n242), .Y(n474) );
  MUX21X1_HVT U323 ( .A1(n386), .A2(n389), .S0(n319), .Y(n442) );
  MUX21X1_HVT U324 ( .A1(n389), .A2(n311), .S0(n323), .Y(n590) );
  MUX21X1_HVT U325 ( .A1(n363), .A2(n237), .S0(n300), .Y(n499) );
  MUX21X1_HVT U326 ( .A1(n452), .A2(n317), .S0(n297), .Y(n451) );
  MUX21X1_HVT U327 ( .A1(n558), .A2(n559), .S0(n302), .Y(n556) );
  MUX21X1_HVT U328 ( .A1(n270), .A2(n575), .S0(in[5]), .Y(n559) );
  XOR2X1_HVT U329 ( .A1(n320), .A2(n301), .Y(n567) );
  MUX21X1_HVT U330 ( .A1(n237), .A2(n325), .S0(n280), .Y(n481) );
  NBUFFX2_HVT U331 ( .A(n600), .Y(n313) );
  MUX21X1_HVT U332 ( .A1(n368), .A2(n383), .S0(n303), .Y(n413) );
  MUX21X1_HVT U333 ( .A1(n311), .A2(n386), .S0(n322), .Y(n397) );
  MUX21X1_HVT U334 ( .A1(n580), .A2(n401), .S0(n302), .Y(n396) );
  MUX21X1_HVT U335 ( .A1(n315), .A2(n270), .S0(n216), .Y(n601) );
  MUX21X1_HVT U336 ( .A1(n346), .A2(n325), .S0(in[5]), .Y(n544) );
  MUX21X1_HVT U337 ( .A1(n311), .A2(n309), .S0(n304), .Y(n518) );
  NBUFFX2_HVT U338 ( .A(n609), .Y(n318) );
  NBUFFX2_HVT U339 ( .A(n390), .Y(n309) );
  XNOR2X1_HVT U340 ( .A1(n333), .A2(n322), .Y(n297) );
  AND2X1_HVT U341 ( .A1(n305), .A2(n325), .Y(n298) );
  NBUFFX2_HVT U342 ( .A(in[5]), .Y(n329) );
  NBUFFX2_HVT U343 ( .A(in[5]), .Y(n328) );
  MUX21X1_HVT U344 ( .A1(n385), .A2(n256), .S0(n321), .Y(n578) );
  NAND2X0_HVT U345 ( .A1(in[4]), .A2(n387), .Y(n600) );
  NAND2X0_HVT U346 ( .A1(in[3]), .A2(in[4]), .Y(n609) );
  MUX21X1_HVT U347 ( .A1(n256), .A2(n388), .S0(n217), .Y(n574) );
  MUX21X1_HVT U348 ( .A1(n256), .A2(n603), .S0(n216), .Y(n399) );
  MUX21X1_HVT U349 ( .A1(n256), .A2(n386), .S0(n321), .Y(n592) );
  MUX21X1_HVT U350 ( .A1(n256), .A2(n317), .S0(n320), .Y(n589) );
  MUX21X1_HVT U351 ( .A1(n256), .A2(n313), .S0(n319), .Y(n392) );
  MUX21X1_HVT U352 ( .A1(n256), .A2(n318), .S0(n319), .Y(n391) );
  MUX21X1_HVT U353 ( .A1(n318), .A2(n256), .S0(n217), .Y(n582) );
  MUX21X1_HVT U354 ( .A1(n270), .A2(n256), .S0(n300), .Y(n494) );
  MUX21X1_HVT U355 ( .A1(n305), .A2(n256), .S0(n216), .Y(n580) );
  NBUFFX2_HVT U356 ( .A(in[3]), .Y(n311) );
  NBUFFX2_HVT U357 ( .A(in[0]), .Y(n310) );
  INVX0_HVT U358 ( .A(n588), .Y(n335) );
  INVX0_HVT U359 ( .A(n586), .Y(n336) );
  INVX0_HVT U360 ( .A(n577), .Y(n337) );
  INVX0_HVT U361 ( .A(n439), .Y(n338) );
  INVX0_HVT U362 ( .A(n402), .Y(n339) );
  INVX0_HVT U363 ( .A(n236), .Y(n340) );
  INVX0_HVT U364 ( .A(n594), .Y(n341) );
  INVX0_HVT U365 ( .A(n606), .Y(n342) );
  INVX0_HVT U366 ( .A(n604), .Y(n343) );
  INVX0_HVT U367 ( .A(n602), .Y(n344) );
  INVX0_HVT U368 ( .A(n601), .Y(n345) );
  INVX0_HVT U369 ( .A(n598), .Y(n346) );
  INVX0_HVT U370 ( .A(n592), .Y(n349) );
  INVX0_HVT U371 ( .A(n591), .Y(n350) );
  INVX0_HVT U372 ( .A(n590), .Y(n351) );
  INVX0_HVT U373 ( .A(n584), .Y(n355) );
  INVX0_HVT U374 ( .A(n582), .Y(n356) );
  INVX0_HVT U375 ( .A(n581), .Y(n357) );
  INVX0_HVT U376 ( .A(n396), .Y(n359) );
  INVX0_HVT U377 ( .A(n579), .Y(n360) );
  INVX0_HVT U378 ( .A(n578), .Y(n361) );
  INVX0_HVT U379 ( .A(n576), .Y(n362) );
  INVX0_HVT U380 ( .A(n574), .Y(n363) );
  INVX0_HVT U381 ( .A(n572), .Y(n364) );
  INVX0_HVT U382 ( .A(n570), .Y(n366) );
  INVX0_HVT U383 ( .A(n569), .Y(n367) );
  INVX0_HVT U384 ( .A(n568), .Y(n368) );
  INVX0_HVT U385 ( .A(n597), .Y(n369) );
  INVX0_HVT U386 ( .A(n496), .Y(n370) );
  INVX0_HVT U387 ( .A(n401), .Y(n371) );
  INVX0_HVT U388 ( .A(n553), .Y(n372) );
  INVX0_HVT U389 ( .A(n455), .Y(n373) );
  INVX0_HVT U390 ( .A(n400), .Y(n374) );
  INVX0_HVT U391 ( .A(n398), .Y(n376) );
  INVX0_HVT U392 ( .A(n397), .Y(n377) );
  INVX0_HVT U393 ( .A(n515), .Y(n378) );
  INVX0_HVT U394 ( .A(n505), .Y(n379) );
  INVX0_HVT U395 ( .A(n394), .Y(n381) );
  INVX0_HVT U396 ( .A(n393), .Y(n382) );
  INVX0_HVT U397 ( .A(n392), .Y(n383) );
  INVX0_HVT U398 ( .A(n391), .Y(n384) );
endmodule

