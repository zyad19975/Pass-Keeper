
module sbox_14 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n50, n87, n210, n211, n212, n213, n216, n217, n218, n219, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608;

  NAND2X0_HVT U4 ( .A1(n313), .A2(n606), .Y(n605) );
  NAND2X0_HVT U5 ( .A1(n322), .A2(n303), .Y(n603) );
  NAND2X0_HVT U13 ( .A1(n595), .A2(n318), .Y(n596) );
  NAND2X0_HVT U15 ( .A1(n606), .A2(n216), .Y(n593) );
  NAND2X0_HVT U21 ( .A1(n313), .A2(n325), .Y(n587) );
  NAND2X0_HVT U24 ( .A1(n309), .A2(n325), .Y(n585) );
  NAND2X0_HVT U33 ( .A1(n385), .A2(n325), .Y(n576) );
  NAND2X0_HVT U35 ( .A1(n217), .A2(n325), .Y(n574) );
  NAND2X0_HVT U42 ( .A1(n320), .A2(n309), .Y(n567) );
  MUX41X1_HVT U51 ( .A1(n373), .A3(n332), .A2(n350), .A4(n351), .S0(n330), 
        .S1(n300), .Y(n559) );
  NAND2X0_HVT U53 ( .A1(n556), .A2(n566), .Y(n557) );
  NAND2X0_HVT U56 ( .A1(n313), .A2(n552), .Y(n553) );
  MUX41X1_HVT U57 ( .A1(n374), .A3(n589), .A2(n553), .A4(n598), .S0(n330), 
        .S1(n300), .Y(n551) );
  NAND2X0_HVT U58 ( .A1(n318), .A2(n606), .Y(n550) );
  MUX41X1_HVT U59 ( .A1(n293), .A3(n550), .A2(n291), .A4(n349), .S0(n330), 
        .S1(n300), .Y(n549) );
  MUX41X1_HVT U61 ( .A1(n289), .A3(n348), .A2(n347), .A4(n216), .S0(n277), 
        .S1(n300), .Y(n547) );
  NAND2X0_HVT U62 ( .A1(n325), .A2(n316), .Y(n546) );
  AO21X1_HVT U66 ( .A1(n344), .A2(n328), .A3(n367), .Y(n542) );
  MUX41X1_HVT U68 ( .A1(n342), .A3(n542), .A2(n541), .A4(n543), .S0(n294), 
        .S1(n278), .Y(n540) );
  MUX41X1_HVT U69 ( .A1(n540), .A3(n548), .A2(n544), .A4(n554), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n311), .A2(n535), .Y(n536) );
  MUX41X1_HVT U74 ( .A1(n537), .A3(n583), .A2(n536), .A4(n585), .S0(n296), 
        .S1(n329), .Y(n534) );
  MUX41X1_HVT U75 ( .A1(n371), .A3(n376), .A2(n388), .A4(n353), .S0(n294), 
        .S1(n264), .Y(n533) );
  MUX41X1_HVT U77 ( .A1(n600), .A3(n378), .A2(n532), .A4(n377), .S0(n301), 
        .S1(in[2]), .Y(n531) );
  AND3X1_HVT U80 ( .A1(n315), .A2(n552), .A3(n527), .Y(n528) );
  MUX41X1_HVT U82 ( .A1(n564), .A3(n351), .A2(n333), .A4(n594), .S0(n294), 
        .S1(n264), .Y(n525) );
  NAND2X0_HVT U85 ( .A1(n325), .A2(n274), .Y(n523) );
  MUX41X1_HVT U90 ( .A1(n563), .A3(n567), .A2(n373), .A4(n520), .S0(n295), 
        .S1(n264), .Y(n519) );
  AO21X1_HVT U93 ( .A1(n302), .A2(n515), .A3(n372), .Y(n516) );
  MUX41X1_HVT U96 ( .A1(n333), .A3(n288), .A2(n375), .A4(n513), .S0(n294), 
        .S1(n264), .Y(n512) );
  MUX41X1_HVT U97 ( .A1(n371), .A3(n288), .A2(n235), .A4(n593), .S0(n294), 
        .S1(n329), .Y(n511) );
  NAND2X0_HVT U101 ( .A1(n506), .A2(n505), .Y(n507) );
  MUX41X1_HVT U103 ( .A1(n606), .A3(n343), .A2(n356), .A4(n574), .S0(n294), 
        .S1(n329), .Y(n503) );
  MUX41X1_HVT U105 ( .A1(n355), .A3(n561), .A2(n502), .A4(n370), .S0(n294), 
        .S1(n329), .Y(n501) );
  OA21X1_HVT U109 ( .A1(n361), .A2(n275), .A3(n349), .Y(n498) );
  NAND2X0_HVT U110 ( .A1(n315), .A2(n496), .Y(n497) );
  MUX41X1_HVT U114 ( .A1(n493), .A3(n499), .A2(n495), .A4(n498), .S0(n328), 
        .S1(n329), .Y(n492) );
  AND2X1_HVT U115 ( .A1(n323), .A2(n216), .Y(n491) );
  MUX41X1_HVT U116 ( .A1(n596), .A3(n491), .A2(n353), .A4(n578), .S0(n295), 
        .S1(n277), .Y(n490) );
  AO21X1_HVT U118 ( .A1(n298), .A2(n310), .A3(n602), .Y(n488) );
  NAND2X0_HVT U123 ( .A1(n482), .A2(n481), .Y(n483) );
  MUX41X1_HVT U125 ( .A1(n587), .A3(n293), .A2(n342), .A4(n380), .S0(n295), 
        .S1(n277), .Y(n479) );
  AND3X1_HVT U128 ( .A1(n297), .A2(n325), .A3(n280), .Y(n476) );
  MUX41X1_HVT U131 ( .A1(n474), .A3(n476), .A2(n475), .A4(n477), .S0(n300), 
        .S1(n277), .Y(n473) );
  MUX41X1_HVT U135 ( .A1(n381), .A3(n386), .A2(n603), .A4(n582), .S0(n296), 
        .S1(n330), .Y(n470) );
  MUX41X1_HVT U139 ( .A1(n467), .A3(n470), .A2(n469), .A4(n471), .S0(n307), 
        .S1(n299), .Y(n466) );
  AND2X1_HVT U140 ( .A1(n310), .A2(n236), .Y(n465) );
  OA21X1_HVT U144 ( .A1(n336), .A2(n265), .A3(n578), .Y(n461) );
  NAND2X0_HVT U146 ( .A1(n323), .A2(n318), .Y(n535) );
  MUX41X1_HVT U147 ( .A1(n382), .A3(n535), .A2(n371), .A4(n563), .S0(n296), 
        .S1(n330), .Y(n459) );
  MUX41X1_HVT U148 ( .A1(n459), .A3(n463), .A2(n460), .A4(n464), .S0(in[0]), 
        .S1(n299), .Y(n458) );
  OA21X1_HVT U151 ( .A1(n569), .A2(n246), .A3(n455), .Y(n456) );
  MUX41X1_HVT U153 ( .A1(n497), .A3(n289), .A2(n314), .A4(n335), .S0(n295), 
        .S1(n264), .Y(n453) );
  AND2X1_HVT U154 ( .A1(n302), .A2(n309), .Y(n452) );
  NAND2X0_HVT U158 ( .A1(n322), .A2(n274), .Y(n448) );
  MUX41X1_HVT U159 ( .A1(n596), .A3(n23), .A2(n448), .A4(n341), .S0(n297), 
        .S1(n329), .Y(n447) );
  AND2X1_HVT U162 ( .A1(n602), .A2(n535), .Y(n444) );
  MUX41X1_HVT U163 ( .A1(n348), .A3(n444), .A2(n287), .A4(n445), .S0(in[2]), 
        .S1(n264), .Y(n443) );
  MUX41X1_HVT U165 ( .A1(n587), .A3(n357), .A2(n563), .A4(n442), .S0(n277), 
        .S1(n327), .Y(n441) );
  NAND2X0_HVT U166 ( .A1(n318), .A2(n552), .Y(n440) );
  NAND2X0_HVT U167 ( .A1(n388), .A2(n325), .Y(n439) );
  MUX41X1_HVT U168 ( .A1(n374), .A3(n310), .A2(n439), .A4(n440), .S0(n326), 
        .S1(n264), .Y(n438) );
  OA21X1_HVT U170 ( .A1(n291), .A2(n265), .A3(n578), .Y(n436) );
  MUX41X1_HVT U172 ( .A1(n435), .A3(n441), .A2(n438), .A4(n443), .S0(n307), 
        .S1(n299), .Y(n434) );
  NAND2X0_HVT U174 ( .A1(n233), .A2(n602), .Y(n595) );
  MUX41X1_HVT U176 ( .A1(n305), .A3(n433), .A2(n379), .A4(n595), .S0(n277), 
        .S1(in[2]), .Y(n432) );
  NAND2X0_HVT U177 ( .A1(n322), .A2(n306), .Y(n431) );
  MUX41X1_HVT U178 ( .A1(n591), .A3(n431), .A2(n383), .A4(n571), .S0(n296), 
        .S1(n278), .Y(n430) );
  MUX41X1_HVT U179 ( .A1(n581), .A3(n384), .A2(n337), .A4(n383), .S0(n327), 
        .S1(n279), .Y(n429) );
  MUX41X1_HVT U180 ( .A1(n340), .A3(n600), .A2(n596), .A4(n285), .S0(n301), 
        .S1(n294), .Y(n428) );
  MUX41X1_HVT U182 ( .A1(n363), .A3(n312), .A2(n365), .A4(n354), .S0(n277), 
        .S1(n327), .Y(n426) );
  OA21X1_HVT U184 ( .A1(n575), .A2(n265), .A3(n352), .Y(n424) );
  MUX41X1_HVT U186 ( .A1(n288), .A3(n570), .A2(n535), .A4(n563), .S0(in[2]), 
        .S1(n279), .Y(n422) );
  MUX41X1_HVT U189 ( .A1(n420), .A3(n595), .A2(n421), .A4(n370), .S0(n301), 
        .S1(in[2]), .Y(n419) );
  MUX41X1_HVT U194 ( .A1(n568), .A3(n582), .A2(n381), .A4(n310), .S0(n301), 
        .S1(n261), .Y(n415) );
  MUX41X1_HVT U195 ( .A1(n602), .A3(n375), .A2(n317), .A4(n572), .S0(n296), 
        .S1(n264), .Y(n414) );
  AO21X1_HVT U197 ( .A1(n290), .A2(n278), .A3(n372), .Y(n412) );
  OA21X1_HVT U201 ( .A1(n601), .A2(n265), .A3(n362), .Y(n408) );
  MUX41X1_HVT U204 ( .A1(n553), .A3(n596), .A2(n360), .A4(n586), .S0(in[2]), 
        .S1(n329), .Y(n405) );
  NAND2X0_HVT U208 ( .A1(n321), .A2(n313), .Y(n496) );
  NAND2X0_HVT U214 ( .A1(n602), .A2(n325), .Y(n402) );
  NAND2X0_HVT U215 ( .A1(n496), .A2(n311), .Y(n401) );
  NAND2X0_HVT U218 ( .A1(n386), .A2(n322), .Y(n455) );
  NAND2X0_HVT U220 ( .A1(n279), .A2(n402), .Y(n527) );
  XOR2X2_HVT U1 ( .A1(n50), .A2(n308), .Y(n23) );
  IBUFFX16_HVT U2 ( .A(n23), .Y(n602) );
  INVX8_HVT U3 ( .A(n389), .Y(n50) );
  XOR2X2_HVT U6 ( .A1(n582), .A2(n246), .Y(n565) );
  MUX21X2_HVT U7 ( .A1(n500), .A2(n510), .S0(n87), .Y(out[2]) );
  IBUFFX16_HVT U8 ( .A(n250), .Y(n87) );
  INVX1_HVT U9 ( .A(in[1]), .Y(n324) );
  INVX1_HVT U10 ( .A(in[1]), .Y(n236) );
  MUX21X1_HVT U11 ( .A1(n580), .A2(n338), .S0(n302), .Y(n462) );
  MUX21X2_HVT U12 ( .A1(n446), .A2(n434), .S0(n210), .Y(out[5]) );
  IBUFFX16_HVT U14 ( .A(in[6]), .Y(n210) );
  MUX41X1_HVT U16 ( .A1(n426), .A3(n423), .A2(n422), .A4(n419), .S0(n211), 
        .S1(n212), .Y(n418) );
  IBUFFX16_HVT U17 ( .A(n328), .Y(n211) );
  IBUFFX16_HVT U18 ( .A(in[0]), .Y(n212) );
  INVX0_HVT U19 ( .A(n23), .Y(n213) );
  INVX1_HVT U20 ( .A(n213), .Y(n216) );
  MUX21X1_HVT U22 ( .A1(n304), .A2(n23), .S0(n236), .Y(n592) );
  INVX2_HVT U23 ( .A(n331), .Y(n330) );
  MUX21X1_HVT U25 ( .A1(n565), .A2(n539), .S0(n298), .Y(n538) );
  INVX1_HVT U26 ( .A(in[4]), .Y(n217) );
  INVX1_HVT U27 ( .A(in[4]), .Y(n389) );
  INVX1_HVT U28 ( .A(n324), .Y(n319) );
  INVX1_HVT U29 ( .A(n324), .Y(n320) );
  INVX1_HVT U30 ( .A(n324), .Y(n322) );
  INVX1_HVT U31 ( .A(n324), .Y(n321) );
  OR2X1_HVT U32 ( .A1(n324), .A2(n218), .Y(n552) );
  IBUFFX16_HVT U34 ( .A(n311), .Y(n218) );
  MUX41X1_HVT U36 ( .A1(n526), .A3(n524), .A2(n525), .A4(n522), .S0(n219), 
        .S1(n231), .Y(n521) );
  IBUFFX16_HVT U37 ( .A(in[0]), .Y(n219) );
  IBUFFX16_HVT U38 ( .A(n299), .Y(n231) );
  MUX21X2_HVT U39 ( .A1(n311), .A2(n588), .S0(n232), .Y(n529) );
  IBUFFX16_HVT U40 ( .A(n302), .Y(n232) );
  NAND2X2_HVT U41 ( .A1(n319), .A2(n315), .Y(n606) );
  INVX2_HVT U43 ( .A(n236), .Y(n323) );
  NBUFFX2_HVT U44 ( .A(n319), .Y(n233) );
  NBUFFX2_HVT U45 ( .A(n319), .Y(n234) );
  NBUFFX2_HVT U46 ( .A(n319), .Y(n235) );
  NAND2X0_HVT U47 ( .A1(n483), .A2(n254), .Y(n255) );
  INVX0_HVT U48 ( .A(n352), .Y(n248) );
  NAND2X0_HVT U49 ( .A1(n334), .A2(n275), .Y(n252) );
  MUX21X1_HVT U50 ( .A1(n605), .A2(n468), .S0(n271), .Y(n467) );
  INVX1_HVT U52 ( .A(n298), .Y(n271) );
  INVX1_HVT U54 ( .A(n297), .Y(n243) );
  INVX1_HVT U55 ( .A(in[6]), .Y(n250) );
  NBUFFX2_HVT U60 ( .A(in[7]), .Y(n302) );
  INVX1_HVT U63 ( .A(in[7]), .Y(n331) );
  INVX0_HVT U64 ( .A(n275), .Y(n261) );
  INVX1_HVT U65 ( .A(n317), .Y(n274) );
  INVX1_HVT U67 ( .A(n307), .Y(n251) );
  INVX1_HVT U70 ( .A(n299), .Y(n272) );
  INVX1_HVT U71 ( .A(n326), .Y(n275) );
  INVX1_HVT U72 ( .A(in[2]), .Y(n260) );
  INVX1_HVT U76 ( .A(n265), .Y(n254) );
  MUX21X2_HVT U78 ( .A1(n418), .A2(n427), .S0(in[6]), .Y(out[6]) );
  MUX41X1_HVT U79 ( .A1(n405), .A3(n407), .A2(n404), .A4(n406), .S0(n307), 
        .S1(n272), .Y(n403) );
  MUX41X1_HVT U81 ( .A1(n606), .A3(n273), .A2(n280), .A4(n384), .S0(n329), 
        .S1(n260), .Y(n404) );
  MUX41X1_HVT U83 ( .A1(n364), .A3(n573), .A2(n577), .A4(n597), .S0(n275), 
        .S1(n264), .Y(n406) );
  INVX1_HVT U84 ( .A(n217), .Y(n280) );
  INVX2_HVT U86 ( .A(n331), .Y(n329) );
  INVX1_HVT U87 ( .A(n330), .Y(n246) );
  DELLN1X2_HVT U88 ( .A(in[7]), .Y(n301) );
  MUX41X1_HVT U89 ( .A1(n376), .A3(n523), .A2(n290), .A4(n286), .S0(n261), 
        .S1(n329), .Y(n522) );
  IBUFFX2_HVT U91 ( .A(n265), .Y(n278) );
  INVX1_HVT U92 ( .A(n588), .Y(n351) );
  MUX21X1_HVT U94 ( .A1(n571), .A2(n378), .S0(n301), .Y(n450) );
  IBUFFX2_HVT U95 ( .A(n571), .Y(n362) );
  MUX21X2_HVT U98 ( .A1(n551), .A2(n549), .S0(n271), .Y(n548) );
  MUX21X1_HVT U99 ( .A1(n592), .A2(n285), .S0(n301), .Y(n409) );
  INVX1_HVT U100 ( .A(n592), .Y(n347) );
  INVX1_HVT U102 ( .A(n247), .Y(n524) );
  NAND2X0_HVT U104 ( .A1(n452), .A2(n237), .Y(n238) );
  NAND2X0_HVT U106 ( .A1(n316), .A2(n292), .Y(n239) );
  NAND2X0_HVT U107 ( .A1(n238), .A2(n239), .Y(n451) );
  INVX0_HVT U108 ( .A(n292), .Y(n237) );
  NAND2X0_HVT U111 ( .A1(n410), .A2(n240), .Y(n241) );
  NAND2X0_HVT U112 ( .A1(n403), .A2(n250), .Y(n242) );
  NAND2X0_HVT U113 ( .A1(n241), .A2(n242), .Y(out[7]) );
  INVX1_HVT U117 ( .A(n250), .Y(n240) );
  MUX21X1_HVT U119 ( .A1(n408), .A2(n409), .S0(n261), .Y(n407) );
  IBUFFX2_HVT U120 ( .A(n601), .Y(n342) );
  MUX21X2_HVT U121 ( .A1(n461), .A2(n462), .S0(n243), .Y(n460) );
  NAND2X0_HVT U122 ( .A1(n516), .A2(n243), .Y(n244) );
  NAND2X0_HVT U124 ( .A1(n517), .A2(n298), .Y(n245) );
  NAND2X0_HVT U126 ( .A1(n244), .A2(n245), .Y(n514) );
  MUX21X1_HVT U127 ( .A1(n316), .A2(n518), .S0(n292), .Y(n517) );
  XNOR2X1_HVT U129 ( .A1(n265), .A2(n234), .Y(n292) );
  MUX41X1_HVT U130 ( .A1(n346), .A3(n368), .A2(n339), .A4(n546), .S0(n246), 
        .S1(n272), .Y(n545) );
  MUX41X1_HVT U132 ( .A1(n449), .A3(n454), .A2(n447), .A4(n453), .S0(n307), 
        .S1(n272), .Y(n446) );
  MUX21X2_HVT U133 ( .A1(n545), .A2(n547), .S0(n326), .Y(n544) );
  MUX41X1_HVT U134 ( .A1(n249), .A3(n347), .A2(n216), .A4(n248), .S0(n271), 
        .S1(n246), .Y(n247) );
  NAND2X0_HVT U136 ( .A1(n234), .A2(n280), .Y(n249) );
  MUX41X1_HVT U137 ( .A1(n514), .A3(n511), .A2(n519), .A4(n512), .S0(n251), 
        .S1(n328), .Y(n510) );
  NBUFFX4_HVT U138 ( .A(in[7]), .Y(n264) );
  NAND2X0_HVT U141 ( .A1(n485), .A2(n296), .Y(n253) );
  NAND2X0_HVT U142 ( .A1(n252), .A2(n253), .Y(n484) );
  NAND2X0_HVT U143 ( .A1(n484), .A2(n265), .Y(n256) );
  NAND2X0_HVT U145 ( .A1(n255), .A2(n256), .Y(n480) );
  NAND2X0_HVT U149 ( .A1(n289), .A2(n257), .Y(n258) );
  NAND2X0_HVT U150 ( .A1(n509), .A2(n562), .Y(n259) );
  NAND2X0_HVT U152 ( .A1(n258), .A2(n259), .Y(n508) );
  INVX0_HVT U155 ( .A(n562), .Y(n257) );
  MUX21X1_HVT U156 ( .A1(n273), .A2(n594), .S0(n298), .Y(n509) );
  INVX1_HVT U157 ( .A(n273), .Y(n578) );
  NAND2X0_HVT U160 ( .A1(n425), .A2(n261), .Y(n262) );
  NAND2X0_HVT U161 ( .A1(n424), .A2(n275), .Y(n263) );
  NAND2X0_HVT U164 ( .A1(n262), .A2(n263), .Y(n423) );
  INVX1_HVT U169 ( .A(n270), .Y(n573) );
  NAND2X0_HVT U171 ( .A1(n586), .A2(n265), .Y(n266) );
  NAND2X0_HVT U173 ( .A1(n363), .A2(n254), .Y(n267) );
  NAND2X0_HVT U175 ( .A1(n266), .A2(n267), .Y(n468) );
  IBUFFX2_HVT U181 ( .A(n330), .Y(n265) );
  NAND2X0_HVT U183 ( .A1(n458), .A2(n250), .Y(n268) );
  NAND2X0_HVT U185 ( .A1(n466), .A2(in[6]), .Y(n269) );
  NAND2X0_HVT U187 ( .A1(n268), .A2(n269), .Y(out[4]) );
  INVX1_HVT U188 ( .A(n570), .Y(n363) );
  MUX21X1_HVT U190 ( .A1(n398), .A2(n317), .S0(n246), .Y(n276) );
  INVX1_HVT U191 ( .A(n398), .Y(n375) );
  INVX1_HVT U192 ( .A(n276), .Y(n539) );
  MUX21X2_HVT U193 ( .A1(n366), .A2(n383), .S0(n279), .Y(n413) );
  MUX21X2_HVT U196 ( .A1(n456), .A2(n457), .S0(n298), .Y(n454) );
  INVX1_HVT U198 ( .A(n396), .Y(n377) );
  MUX41X1_HVT U199 ( .A1(n432), .A3(n429), .A2(n430), .A4(n428), .S0(n251), 
        .S1(n272), .Y(n427) );
  MUX21X2_HVT U200 ( .A1(n521), .A2(n530), .S0(in[6]), .Y(out[1]) );
  MUX21X2_HVT U202 ( .A1(n479), .A2(n480), .S0(n300), .Y(n478) );
  MUX21X1_HVT U203 ( .A1(n305), .A2(n317), .S0(n320), .Y(n270) );
  MUX21X2_HVT U205 ( .A1(n451), .A2(n450), .S0(n271), .Y(n449) );
  INVX1_HVT U206 ( .A(n577), .Y(n359) );
  AO21X2_HVT U207 ( .A1(n236), .A2(n386), .A3(n246), .Y(n506) );
  MUX41X1_HVT U209 ( .A1(n573), .A3(n382), .A2(n576), .A4(n286), .S0(n275), 
        .S1(n331), .Y(n469) );
  MUX21X2_HVT U210 ( .A1(n555), .A2(n559), .S0(n297), .Y(n554) );
  MUX41X1_HVT U211 ( .A1(n508), .A3(n503), .A2(n504), .A4(n501), .S0(n251), 
        .S1(n272), .Y(n500) );
  MUX21X1_HVT U212 ( .A1(n274), .A2(n386), .S0(n235), .Y(n273) );
  MUX21X2_HVT U213 ( .A1(n412), .A2(n413), .S0(n271), .Y(n411) );
  MUX41X1_HVT U216 ( .A1(n574), .A3(n567), .A2(n417), .A4(n560), .S0(n275), 
        .S1(n264), .Y(n416) );
  INVX1_HVT U217 ( .A(n391), .Y(n383) );
  MUX41X1_HVT U219 ( .A1(n538), .A3(n533), .A2(n534), .A4(n531), .S0(n251), 
        .S1(n272), .Y(n530) );
  MUX41X1_HVT U221 ( .A1(n414), .A3(n416), .A2(n411), .A4(n415), .S0(in[0]), 
        .S1(n272), .Y(n410) );
  NBUFFX2_HVT U222 ( .A(n330), .Y(n277) );
  INVX0_HVT U223 ( .A(n265), .Y(n279) );
  MUX21X1_HVT U224 ( .A1(n309), .A2(n23), .S0(n236), .Y(n586) );
  MUX41X1_HVT U225 ( .A1(n310), .A3(n369), .A2(n216), .A4(n352), .S0(n271), 
        .S1(n246), .Y(n463) );
  MUX41X1_HVT U226 ( .A1(n359), .A3(n465), .A2(n362), .A4(n584), .S0(n271), 
        .S1(n246), .Y(n464) );
  INVX2_HVT U227 ( .A(n260), .Y(n327) );
  NAND2X0_HVT U228 ( .A1(n316), .A2(n281), .Y(n282) );
  NAND2X0_HVT U229 ( .A1(n494), .A2(n284), .Y(n283) );
  NAND2X0_HVT U230 ( .A1(n282), .A2(n283), .Y(n493) );
  INVX0_HVT U231 ( .A(n284), .Y(n281) );
  MUX41X1_HVT U232 ( .A1(n492), .A3(n486), .A2(n478), .A4(n473), .S0(n251), 
        .S1(n250), .Y(out[3]) );
  XNOR2X1_HVT U233 ( .A1(n322), .A2(n327), .Y(n284) );
  XOR2X1_HVT U234 ( .A1(n275), .A2(n246), .Y(n562) );
  INVX0_HVT U235 ( .A(n308), .Y(n387) );
  INVX1_HVT U236 ( .A(n312), .Y(n385) );
  MUX21X1_HVT U237 ( .A1(n287), .A2(n347), .S0(n295), .Y(n475) );
  AND2X1_HVT U238 ( .A1(n216), .A2(n552), .Y(n285) );
  NBUFFX2_HVT U239 ( .A(n604), .Y(n312) );
  INVX1_HVT U240 ( .A(n314), .Y(n388) );
  MUX21X1_HVT U241 ( .A1(n385), .A2(n274), .S0(n328), .Y(n556) );
  NBUFFX2_HVT U242 ( .A(n604), .Y(n313) );
  MUX21X1_HVT U243 ( .A1(n343), .A2(n386), .S0(n299), .Y(n541) );
  MUX21X1_HVT U244 ( .A1(n578), .A2(n497), .S0(n295), .Y(n495) );
  AND2X1_HVT U245 ( .A1(n315), .A2(n535), .Y(n286) );
  MUX21X1_HVT U246 ( .A1(n23), .A2(n274), .S0(n319), .Y(n601) );
  MUX21X1_HVT U247 ( .A1(n315), .A2(n216), .S0(n321), .Y(n568) );
  MUX21X1_HVT U248 ( .A1(n216), .A2(n217), .S0(n323), .Y(n505) );
  MUX21X1_HVT U249 ( .A1(n385), .A2(n388), .S0(n320), .Y(n433) );
  MUX21X1_HVT U250 ( .A1(n274), .A2(n216), .S0(n322), .Y(n445) );
  MUX21X1_HVT U251 ( .A1(n216), .A2(n385), .S0(n233), .Y(n513) );
  MUX21X1_HVT U252 ( .A1(n602), .A2(n388), .S0(n320), .Y(n584) );
  MUX21X1_HVT U253 ( .A1(n313), .A2(n602), .S0(n321), .Y(n572) );
  MUX21X1_HVT U254 ( .A1(n602), .A2(n386), .S0(n234), .Y(n393) );
  MUX21X1_HVT U255 ( .A1(n313), .A2(n311), .S0(n234), .Y(n520) );
  MUX21X1_HVT U256 ( .A1(n602), .A2(n217), .S0(n235), .Y(n532) );
  XOR2X1_HVT U257 ( .A1(n602), .A2(n319), .Y(n563) );
  MUX21X1_HVT U258 ( .A1(n303), .A2(n602), .S0(n320), .Y(n396) );
  MUX21X1_HVT U259 ( .A1(n388), .A2(n274), .S0(n319), .Y(n582) );
  MUX21X1_HVT U260 ( .A1(n274), .A2(n385), .S0(n233), .Y(n571) );
  MUX21X1_HVT U261 ( .A1(n274), .A2(n303), .S0(n322), .Y(n575) );
  MUX21X1_HVT U262 ( .A1(n304), .A2(n388), .S0(n233), .Y(n569) );
  MUX21X1_HVT U263 ( .A1(n305), .A2(n385), .S0(n323), .Y(n580) );
  MUX21X1_HVT U264 ( .A1(n358), .A2(n472), .S0(n297), .Y(n471) );
  MUX21X1_HVT U265 ( .A1(n380), .A2(n311), .S0(n330), .Y(n472) );
  MUX21X1_HVT U266 ( .A1(n488), .A2(n489), .S0(n254), .Y(n487) );
  MUX21X1_HVT U267 ( .A1(n335), .A2(n360), .S0(n295), .Y(n489) );
  NAND2X0_HVT U268 ( .A1(n306), .A2(n387), .Y(n604) );
  MUX21X1_HVT U269 ( .A1(n385), .A2(n306), .S0(n319), .Y(n394) );
  NBUFFX2_HVT U270 ( .A(n607), .Y(n314) );
  MUX21X1_HVT U271 ( .A1(n316), .A2(n311), .S0(n323), .Y(n594) );
  MUX21X1_HVT U272 ( .A1(n312), .A2(n318), .S0(n321), .Y(n515) );
  MUX21X1_HVT U273 ( .A1(n305), .A2(n304), .S0(n234), .Y(n485) );
  NBUFFX2_HVT U274 ( .A(n607), .Y(n315) );
  NBUFFX2_HVT U275 ( .A(n607), .Y(n316) );
  XOR2X1_HVT U276 ( .A1(n322), .A2(n386), .Y(n564) );
  MUX21X1_HVT U277 ( .A1(n304), .A2(n318), .S0(n235), .Y(n420) );
  MUX21X1_HVT U278 ( .A1(n317), .A2(n315), .S0(n321), .Y(n421) );
  MUX21X1_HVT U279 ( .A1(n386), .A2(n385), .S0(n320), .Y(n590) );
  INVX1_HVT U280 ( .A(n310), .Y(n386) );
  MUX21X1_HVT U281 ( .A1(n304), .A2(n274), .S0(n319), .Y(n598) );
  MUX21X1_HVT U282 ( .A1(n313), .A2(n303), .S0(n321), .Y(n597) );
  MUX21X1_HVT U283 ( .A1(n303), .A2(n306), .S0(n321), .Y(n417) );
  XOR2X1_HVT U284 ( .A1(n314), .A2(n320), .Y(n560) );
  MUX21X1_HVT U285 ( .A1(n314), .A2(n305), .S0(n323), .Y(n400) );
  XNOR2X1_HVT U286 ( .A1(n312), .A2(n322), .Y(n287) );
  AND2X1_HVT U287 ( .A1(n320), .A2(n388), .Y(n288) );
  MUX21X1_HVT U288 ( .A1(n314), .A2(n313), .S0(n321), .Y(n392) );
  AND2X1_HVT U289 ( .A1(n318), .A2(n496), .Y(n289) );
  XNOR2X1_HVT U290 ( .A1(n317), .A2(n320), .Y(n290) );
  MUX21X1_HVT U291 ( .A1(n311), .A2(n303), .S0(n323), .Y(n398) );
  MUX21X1_HVT U292 ( .A1(n311), .A2(n306), .S0(n320), .Y(n537) );
  MUX21X1_HVT U293 ( .A1(n311), .A2(n318), .S0(n297), .Y(n482) );
  XOR2X1_HVT U294 ( .A1(n306), .A2(n320), .Y(n583) );
  NBUFFX2_HVT U295 ( .A(n387), .Y(n303) );
  NBUFFX2_HVT U296 ( .A(n387), .Y(n304) );
  NBUFFX2_HVT U297 ( .A(n326), .Y(n295) );
  NBUFFX2_HVT U298 ( .A(n326), .Y(n296) );
  NBUFFX2_HVT U299 ( .A(n327), .Y(n297) );
  NBUFFX2_HVT U300 ( .A(n327), .Y(n298) );
  NBUFFX2_HVT U301 ( .A(in[5]), .Y(n300) );
  NBUFFX2_HVT U302 ( .A(n326), .Y(n294) );
  NBUFFX2_HVT U303 ( .A(in[5]), .Y(n299) );
  MUX21X1_HVT U304 ( .A1(n507), .A2(n358), .S0(n297), .Y(n504) );
  MUX21X1_HVT U305 ( .A1(n523), .A2(n309), .S0(n302), .Y(n425) );
  XOR2X1_HVT U306 ( .A1(n323), .A2(n308), .Y(n561) );
  MUX21X1_HVT U307 ( .A1(n311), .A2(n216), .S0(n323), .Y(n502) );
  MUX21X1_HVT U308 ( .A1(n377), .A2(n386), .S0(n278), .Y(n457) );
  MUX21X1_HVT U309 ( .A1(n529), .A2(n528), .S0(n298), .Y(n526) );
  MUX21X1_HVT U310 ( .A1(n437), .A2(n436), .S0(n297), .Y(n435) );
  MUX21X1_HVT U311 ( .A1(n311), .A2(n375), .S0(n302), .Y(n437) );
  MUX21X1_HVT U312 ( .A1(n386), .A2(n388), .S0(n322), .Y(n442) );
  AND2X1_HVT U313 ( .A1(n216), .A2(n325), .Y(n291) );
  MUX21X1_HVT U314 ( .A1(n309), .A2(n385), .S0(n321), .Y(n570) );
  MUX21X1_HVT U315 ( .A1(n591), .A2(n359), .S0(n296), .Y(n474) );
  NAND2X0_HVT U316 ( .A1(n308), .A2(n305), .Y(n607) );
  NBUFFX2_HVT U317 ( .A(n389), .Y(n306) );
  NBUFFX2_HVT U318 ( .A(n608), .Y(n317) );
  MUX21X1_HVT U319 ( .A1(n388), .A2(n309), .S0(n323), .Y(n589) );
  MUX21X1_HVT U320 ( .A1(n270), .A2(n606), .S0(n296), .Y(n499) );
  MUX21X1_HVT U321 ( .A1(n557), .A2(n558), .S0(n301), .Y(n555) );
  MUX21X1_HVT U322 ( .A1(n309), .A2(n574), .S0(n328), .Y(n558) );
  XOR2X1_HVT U323 ( .A1(n235), .A2(n328), .Y(n566) );
  MUX21X1_HVT U324 ( .A1(n606), .A2(n236), .S0(n261), .Y(n481) );
  NBUFFX2_HVT U325 ( .A(n599), .Y(n310) );
  MUX21X1_HVT U326 ( .A1(n309), .A2(n386), .S0(n322), .Y(n397) );
  MUX21X1_HVT U327 ( .A1(n579), .A2(n401), .S0(n301), .Y(n395) );
  MUX21X1_HVT U328 ( .A1(n313), .A2(n309), .S0(n323), .Y(n600) );
  MUX21X1_HVT U329 ( .A1(n345), .A2(n325), .S0(n328), .Y(n543) );
  MUX21X1_HVT U330 ( .A1(n309), .A2(n217), .S0(n302), .Y(n518) );
  NBUFFX2_HVT U331 ( .A(n599), .Y(n311) );
  MUX21X1_HVT U332 ( .A1(n355), .A2(n579), .S0(n296), .Y(n477) );
  NBUFFX2_HVT U333 ( .A(n608), .Y(n318) );
  NBUFFX2_HVT U334 ( .A(n389), .Y(n305) );
  AND2X1_HVT U335 ( .A1(n304), .A2(n325), .Y(n293) );
  INVX1_HVT U336 ( .A(n260), .Y(n326) );
  NBUFFX2_HVT U337 ( .A(in[5]), .Y(n328) );
  MUX21X1_HVT U338 ( .A1(n487), .A2(n490), .S0(n300), .Y(n486) );
  MUX21X1_HVT U339 ( .A1(n385), .A2(n280), .S0(n323), .Y(n577) );
  NAND2X0_HVT U340 ( .A1(n308), .A2(in[4]), .Y(n608) );
  MUX21X1_HVT U341 ( .A1(n280), .A2(n602), .S0(n321), .Y(n399) );
  MUX21X1_HVT U342 ( .A1(n280), .A2(n386), .S0(n233), .Y(n591) );
  NAND2X0_HVT U343 ( .A1(in[4]), .A2(n387), .Y(n599) );
  MUX21X1_HVT U344 ( .A1(n280), .A2(n316), .S0(n319), .Y(n588) );
  MUX21X1_HVT U345 ( .A1(n280), .A2(n311), .S0(n322), .Y(n391) );
  MUX21X1_HVT U346 ( .A1(n318), .A2(n280), .S0(n321), .Y(n581) );
  MUX21X1_HVT U347 ( .A1(n309), .A2(n280), .S0(n295), .Y(n494) );
  MUX21X1_HVT U348 ( .A1(n280), .A2(n318), .S0(n323), .Y(n390) );
  MUX21X1_HVT U349 ( .A1(n303), .A2(n280), .S0(n319), .Y(n579) );
  NBUFFX2_HVT U350 ( .A(in[3]), .Y(n308) );
  INVX0_HVT U351 ( .A(in[1]), .Y(n325) );
  NBUFFX2_HVT U352 ( .A(in[3]), .Y(n309) );
  NBUFFX2_HVT U353 ( .A(in[0]), .Y(n307) );
  INVX0_HVT U354 ( .A(n587), .Y(n332) );
  INVX0_HVT U355 ( .A(n585), .Y(n333) );
  INVX0_HVT U356 ( .A(n576), .Y(n334) );
  INVX0_HVT U357 ( .A(n574), .Y(n335) );
  INVX0_HVT U358 ( .A(n439), .Y(n336) );
  INVX0_HVT U359 ( .A(n402), .Y(n337) );
  INVX0_HVT U360 ( .A(n606), .Y(n338) );
  INVX0_HVT U361 ( .A(n593), .Y(n339) );
  INVX0_HVT U362 ( .A(n605), .Y(n340) );
  INVX0_HVT U363 ( .A(n603), .Y(n341) );
  INVX0_HVT U364 ( .A(n600), .Y(n343) );
  INVX0_HVT U365 ( .A(n598), .Y(n344) );
  INVX0_HVT U366 ( .A(n597), .Y(n345) );
  INVX0_HVT U367 ( .A(n594), .Y(n346) );
  INVX0_HVT U368 ( .A(n591), .Y(n348) );
  INVX0_HVT U369 ( .A(n590), .Y(n349) );
  INVX0_HVT U370 ( .A(n589), .Y(n350) );
  INVX0_HVT U371 ( .A(n586), .Y(n352) );
  INVX0_HVT U372 ( .A(n584), .Y(n353) );
  INVX0_HVT U373 ( .A(n583), .Y(n354) );
  INVX0_HVT U374 ( .A(n581), .Y(n355) );
  INVX0_HVT U375 ( .A(n580), .Y(n356) );
  INVX0_HVT U376 ( .A(n579), .Y(n357) );
  INVX0_HVT U377 ( .A(n395), .Y(n358) );
  INVX0_HVT U378 ( .A(n575), .Y(n360) );
  INVX0_HVT U379 ( .A(n572), .Y(n361) );
  INVX0_HVT U380 ( .A(n569), .Y(n364) );
  INVX0_HVT U381 ( .A(n568), .Y(n365) );
  INVX0_HVT U382 ( .A(n567), .Y(n366) );
  INVX0_HVT U383 ( .A(n535), .Y(n367) );
  INVX0_HVT U384 ( .A(n596), .Y(n368) );
  INVX0_HVT U385 ( .A(n496), .Y(n369) );
  INVX0_HVT U386 ( .A(n401), .Y(n370) );
  INVX0_HVT U387 ( .A(n552), .Y(n371) );
  INVX0_HVT U388 ( .A(n455), .Y(n372) );
  INVX0_HVT U389 ( .A(n400), .Y(n373) );
  INVX0_HVT U390 ( .A(n399), .Y(n374) );
  INVX0_HVT U391 ( .A(n397), .Y(n376) );
  INVX0_HVT U392 ( .A(n515), .Y(n378) );
  INVX0_HVT U393 ( .A(n505), .Y(n379) );
  INVX0_HVT U394 ( .A(n394), .Y(n380) );
  INVX0_HVT U395 ( .A(n393), .Y(n381) );
  INVX0_HVT U396 ( .A(n392), .Y(n382) );
  INVX0_HVT U397 ( .A(n390), .Y(n384) );
endmodule

