
module sbox_9 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n45, n48, n50, n72, n210, n211, n212, n213, n216, n217, n218,
         n219, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584;

  NAND2X0_HVT U3 ( .A1(n238), .A2(n285), .Y(n582) );
  NAND2X0_HVT U4 ( .A1(n283), .A2(n582), .Y(n581) );
  NAND2X0_HVT U5 ( .A1(n290), .A2(n272), .Y(n579) );
  NAND2X0_HVT U13 ( .A1(n571), .A2(n584), .Y(n572) );
  NAND2X0_HVT U15 ( .A1(n582), .A2(n274), .Y(n569) );
  NAND2X0_HVT U21 ( .A1(n282), .A2(n295), .Y(n563) );
  NAND2X0_HVT U24 ( .A1(n279), .A2(n295), .Y(n561) );
  NAND2X0_HVT U33 ( .A1(n361), .A2(n295), .Y(n552) );
  NAND2X0_HVT U35 ( .A1(n277), .A2(n295), .Y(n550) );
  NAND2X0_HVT U42 ( .A1(n239), .A2(n279), .Y(n543) );
  MUX41X1_HVT U51 ( .A1(n349), .A3(n306), .A2(n324), .A4(n325), .S0(n302), 
        .S1(n299), .Y(n537) );
  NAND2X0_HVT U53 ( .A1(n534), .A2(n542), .Y(n535) );
  NAND2X0_HVT U56 ( .A1(n283), .A2(n530), .Y(n531) );
  MUX41X1_HVT U57 ( .A1(n350), .A3(n565), .A2(n531), .A4(n574), .S0(n245), 
        .S1(n299), .Y(n529) );
  NAND2X0_HVT U58 ( .A1(n584), .A2(n582), .Y(n528) );
  MUX41X1_HVT U59 ( .A1(n260), .A3(n528), .A2(n258), .A4(n323), .S0(n304), 
        .S1(n299), .Y(n527) );
  MUX41X1_HVT U61 ( .A1(n257), .A3(n322), .A2(n321), .A4(n273), .S0(n245), 
        .S1(in[5]), .Y(n525) );
  NAND2X0_HVT U62 ( .A1(n295), .A2(n286), .Y(n524) );
  MUX41X1_HVT U63 ( .A1(n524), .A3(n313), .A2(n344), .A4(n320), .S0(n245), 
        .S1(n299), .Y(n523) );
  AO21X1_HVT U66 ( .A1(n318), .A2(n268), .A3(n343), .Y(n520) );
  MUX41X1_HVT U68 ( .A1(n316), .A3(n520), .A2(n519), .A4(n521), .S0(n261), 
        .S1(n302), .Y(n518) );
  MUX41X1_HVT U69 ( .A1(n518), .A3(n526), .A2(n522), .A4(n532), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n280), .A2(n514), .Y(n515) );
  MUX41X1_HVT U75 ( .A1(n347), .A3(n352), .A2(n365), .A4(n327), .S0(n261), 
        .S1(n303), .Y(n512) );
  MUX41X1_HVT U77 ( .A1(n576), .A3(n354), .A2(n511), .A4(n353), .S0(n269), 
        .S1(n297), .Y(n510) );
  MUX41X1_HVT U78 ( .A1(n510), .A3(n513), .A2(n512), .A4(n517), .S0(in[0]), 
        .S1(n300), .Y(n509) );
  AND3X1_HVT U80 ( .A1(n285), .A2(n530), .A3(n506), .Y(n507) );
  AND2X1_HVT U83 ( .A1(n238), .A2(n244), .Y(n503) );
  MUX41X1_HVT U84 ( .A1(n326), .A3(n578), .A2(n568), .A4(n503), .S0(n261), 
        .S1(n302), .Y(n502) );
  NAND2X0_HVT U85 ( .A1(n295), .A2(n364), .Y(n501) );
  MUX41X1_HVT U86 ( .A1(n352), .A3(n501), .A2(n255), .A4(n253), .S0(n261), 
        .S1(n304), .Y(n500) );
  MUX41X1_HVT U87 ( .A1(n500), .A3(n504), .A2(n502), .A4(n505), .S0(in[0]), 
        .S1(n299), .Y(n499) );
  MUX41X1_HVT U90 ( .A1(n540), .A3(n543), .A2(n349), .A4(n498), .S0(n262), 
        .S1(n303), .Y(n497) );
  AO21X1_HVT U93 ( .A1(n271), .A2(n493), .A3(n348), .Y(n494) );
  MUX41X1_HVT U96 ( .A1(n307), .A3(n256), .A2(n351), .A4(n491), .S0(n261), 
        .S1(n302), .Y(n490) );
  MUX41X1_HVT U97 ( .A1(n347), .A3(n256), .A2(n238), .A4(n569), .S0(n261), 
        .S1(n303), .Y(n489) );
  MUX41X1_HVT U98 ( .A1(n489), .A3(n492), .A2(n490), .A4(n497), .S0(n278), 
        .S1(n299), .Y(n488) );
  NAND2X0_HVT U101 ( .A1(n484), .A2(n483), .Y(n485) );
  MUX41X1_HVT U103 ( .A1(n582), .A3(n317), .A2(n330), .A4(n550), .S0(n261), 
        .S1(n304), .Y(n481) );
  MUX41X1_HVT U105 ( .A1(n329), .A3(n539), .A2(n480), .A4(n346), .S0(n261), 
        .S1(n303), .Y(n479) );
  NAND2X0_HVT U110 ( .A1(n285), .A2(n474), .Y(n475) );
  AND2X1_HVT U115 ( .A1(n291), .A2(n273), .Y(n469) );
  MUX41X1_HVT U116 ( .A1(n572), .A3(n469), .A2(n327), .A4(n554), .S0(n262), 
        .S1(n245), .Y(n468) );
  NAND2X0_HVT U123 ( .A1(n460), .A2(n459), .Y(n461) );
  MUX41X1_HVT U125 ( .A1(n563), .A3(n260), .A2(n316), .A4(n356), .S0(n262), 
        .S1(n245), .Y(n457) );
  AND3X1_HVT U128 ( .A1(n265), .A2(n295), .A3(n244), .Y(n454) );
  MUX41X1_HVT U131 ( .A1(n452), .A3(n454), .A2(n453), .A4(n455), .S0(n268), 
        .S1(n245), .Y(n451) );
  MUX41X1_HVT U132 ( .A1(n451), .A3(n464), .A2(n456), .A4(n470), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  MUX41X1_HVT U135 ( .A1(n357), .A3(n362), .A2(n579), .A4(n558), .S0(n263), 
        .S1(n302), .Y(n448) );
  MUX41X1_HVT U136 ( .A1(n253), .A3(n552), .A2(n358), .A4(n549), .S0(n262), 
        .S1(n303), .Y(n447) );
  MUX41X1_HVT U139 ( .A1(n445), .A3(n448), .A2(n447), .A4(n449), .S0(n278), 
        .S1(n299), .Y(n444) );
  AND2X1_HVT U140 ( .A1(n281), .A2(n294), .Y(n443) );
  MUX41X1_HVT U142 ( .A1(n326), .A3(n273), .A2(n345), .A4(n281), .S0(n262), 
        .S1(n302), .Y(n441) );
  NAND2X0_HVT U146 ( .A1(n290), .A2(n288), .Y(n514) );
  MUX41X1_HVT U147 ( .A1(n358), .A3(n514), .A2(n347), .A4(n540), .S0(n263), 
        .S1(n302), .Y(n437) );
  MUX41X1_HVT U148 ( .A1(n437), .A3(n441), .A2(n438), .A4(n442), .S0(in[0]), 
        .S1(n267), .Y(n436) );
  OA21X1_HVT U151 ( .A1(n545), .A2(n249), .A3(n433), .Y(n434) );
  MUX41X1_HVT U153 ( .A1(n475), .A3(n257), .A2(n284), .A4(n309), .S0(n262), 
        .S1(n304), .Y(n431) );
  AND2X1_HVT U154 ( .A1(n271), .A2(n279), .Y(n430) );
  NAND2X0_HVT U158 ( .A1(n239), .A2(n364), .Y(n426) );
  MUX41X1_HVT U159 ( .A1(n572), .A3(n273), .A2(n426), .A4(n315), .S0(in[2]), 
        .S1(n303), .Y(n425) );
  MUX41X1_HVT U160 ( .A1(n425), .A3(n431), .A2(n427), .A4(n432), .S0(n278), 
        .S1(n267), .Y(n424) );
  AND2X1_HVT U162 ( .A1(n578), .A2(n514), .Y(n422) );
  MUX41X1_HVT U163 ( .A1(n322), .A3(n422), .A2(n254), .A4(n423), .S0(in[2]), 
        .S1(n303), .Y(n421) );
  MUX41X1_HVT U165 ( .A1(n563), .A3(n331), .A2(n540), .A4(n420), .S0(n304), 
        .S1(n266), .Y(n419) );
  NAND2X0_HVT U166 ( .A1(n584), .A2(n530), .Y(n418) );
  NAND2X0_HVT U167 ( .A1(n365), .A2(n295), .Y(n417) );
  MUX41X1_HVT U168 ( .A1(n350), .A3(n280), .A2(n417), .A4(n418), .S0(in[2]), 
        .S1(n304), .Y(n416) );
  MUX41X1_HVT U172 ( .A1(n413), .A3(n419), .A2(n416), .A4(n421), .S0(in[0]), 
        .S1(n300), .Y(n412) );
  NAND2X0_HVT U174 ( .A1(n239), .A2(n578), .Y(n571) );
  MUX41X1_HVT U176 ( .A1(n276), .A3(n411), .A2(n355), .A4(n571), .S0(n245), 
        .S1(n297), .Y(n410) );
  NAND2X0_HVT U177 ( .A1(n292), .A2(n276), .Y(n409) );
  MUX41X1_HVT U178 ( .A1(n567), .A3(n409), .A2(n359), .A4(n547), .S0(n263), 
        .S1(n304), .Y(n408) );
  MUX41X1_HVT U179 ( .A1(n557), .A3(n360), .A2(n311), .A4(n359), .S0(in[2]), 
        .S1(n304), .Y(n407) );
  MUX41X1_HVT U180 ( .A1(n314), .A3(n576), .A2(n572), .A4(n252), .S0(n269), 
        .S1(n261), .Y(n406) );
  MUX41X1_HVT U181 ( .A1(n406), .A3(n408), .A2(n407), .A4(n410), .S0(n278), 
        .S1(n267), .Y(n405) );
  MUX41X1_HVT U182 ( .A1(n339), .A3(n283), .A2(n341), .A4(n328), .S0(n245), 
        .S1(n297), .Y(n404) );
  OA21X1_HVT U184 ( .A1(n551), .A2(n241), .A3(n326), .Y(n402) );
  MUX41X1_HVT U186 ( .A1(n256), .A3(n546), .A2(n514), .A4(n540), .S0(n296), 
        .S1(n302), .Y(n400) );
  MUX41X1_HVT U189 ( .A1(n398), .A3(n571), .A2(n399), .A4(n346), .S0(n269), 
        .S1(n263), .Y(n397) );
  MUX41X1_HVT U190 ( .A1(n397), .A3(n400), .A2(n401), .A4(n404), .S0(n267), 
        .S1(n278), .Y(n396) );
  MUX41X1_HVT U193 ( .A1(n543), .A3(n550), .A2(n538), .A4(n395), .S0(n296), 
        .S1(n303), .Y(n394) );
  MUX41X1_HVT U195 ( .A1(n578), .A3(n351), .A2(n287), .A4(n548), .S0(in[2]), 
        .S1(n304), .Y(n392) );
  AO21X1_HVT U197 ( .A1(n255), .A2(n270), .A3(n348), .Y(n390) );
  MUX41X1_HVT U199 ( .A1(n389), .A3(n393), .A2(n392), .A4(n394), .S0(in[0]), 
        .S1(n267), .Y(n388) );
  OA21X1_HVT U201 ( .A1(n577), .A2(n241), .A3(n338), .Y(n386) );
  MUX41X1_HVT U203 ( .A1(n549), .A3(n340), .A2(n573), .A4(n553), .S0(in[2]), 
        .S1(n302), .Y(n384) );
  MUX41X1_HVT U204 ( .A1(n531), .A3(n572), .A2(n335), .A4(n562), .S0(in[2]), 
        .S1(n301), .Y(n383) );
  MUX41X1_HVT U205 ( .A1(n244), .A3(n582), .A2(n360), .A4(n333), .S0(in[2]), 
        .S1(n301), .Y(n382) );
  NAND2X0_HVT U208 ( .A1(n239), .A2(n282), .Y(n474) );
  NAND2X0_HVT U212 ( .A1(n289), .A2(n280), .Y(n530) );
  NAND2X0_HVT U214 ( .A1(n578), .A2(n295), .Y(n380) );
  NAND2X0_HVT U215 ( .A1(n474), .A2(n281), .Y(n379) );
  AO21X1_HVT U216 ( .A1(n294), .A2(n362), .A3(n241), .Y(n484) );
  NAND2X0_HVT U218 ( .A1(n362), .A2(n293), .Y(n433) );
  NAND2X0_HVT U220 ( .A1(n270), .A2(n380), .Y(n506) );
  MUX21X1_HVT U1 ( .A1(n45), .A2(n240), .S0(n264), .Y(n23) );
  IBUFFX16_HVT U2 ( .A(n23), .Y(n517) );
  XNOR2X2_HVT U6 ( .A1(n249), .A2(n558), .Y(n45) );
  MUX21X2_HVT U7 ( .A1(n275), .A2(n364), .S0(n289), .Y(n577) );
  MUX21X2_HVT U8 ( .A1(n274), .A2(n361), .S0(n238), .Y(n491) );
  NBUFFX2_HVT U9 ( .A(n366), .Y(n275) );
  MUX21X2_HVT U10 ( .A1(n288), .A2(n284), .S0(n295), .Y(n242) );
  MUX41X1_HVT U11 ( .A1(n471), .A3(n473), .A2(n477), .A4(n476), .S0(n303), 
        .S1(n268), .Y(n470) );
  INVX0_HVT U12 ( .A(n568), .Y(n321) );
  NAND2X0_HVT U14 ( .A1(n279), .A2(n48), .Y(n50) );
  NAND2X0_HVT U16 ( .A1(n275), .A2(n216), .Y(n72) );
  NAND2X0_HVT U17 ( .A1(n50), .A2(n72), .Y(n562) );
  INVX8_HVT U18 ( .A(n216), .Y(n48) );
  MUX21X2_HVT U19 ( .A1(n444), .A2(n436), .S0(n210), .Y(out[4]) );
  IBUFFX16_HVT U20 ( .A(in[6]), .Y(n210) );
  IBUFFX2_HVT U22 ( .A(n293), .Y(n216) );
  MUX21X1_HVT U23 ( .A1(n562), .A2(n339), .S0(n270), .Y(n446) );
  NAND2X0_HVT U25 ( .A1(n487), .A2(n211), .Y(n212) );
  NAND2X0_HVT U26 ( .A1(n257), .A2(n250), .Y(n213) );
  NAND2X0_HVT U27 ( .A1(n212), .A2(n213), .Y(n486) );
  INVX0_HVT U28 ( .A(n250), .Y(n211) );
  XNOR2X1_HVT U29 ( .A1(n243), .A2(n305), .Y(n250) );
  MUX21X2_HVT U30 ( .A1(n424), .A2(n412), .S0(n247), .Y(out[5]) );
  INVX2_HVT U31 ( .A(n305), .Y(n301) );
  NBUFFX4_HVT U32 ( .A(n301), .Y(n269) );
  INVX2_HVT U34 ( .A(n242), .Y(n558) );
  MUX21X2_HVT U36 ( .A1(n465), .A2(n468), .S0(n268), .Y(n464) );
  NAND2X0_HVT U37 ( .A1(n388), .A2(n217), .Y(n218) );
  NAND2X0_HVT U38 ( .A1(n381), .A2(n247), .Y(n219) );
  NAND2X0_HVT U39 ( .A1(n218), .A2(n219), .Y(out[7]) );
  IBUFFX2_HVT U40 ( .A(n247), .Y(n217) );
  INVX2_HVT U41 ( .A(n305), .Y(n303) );
  INVX4_HVT U43 ( .A(in[7]), .Y(n305) );
  NAND2X0_HVT U44 ( .A1(n252), .A2(n231), .Y(n232) );
  NAND2X0_HVT U45 ( .A1(n568), .A2(n241), .Y(n233) );
  NAND2X0_HVT U46 ( .A1(n232), .A2(n233), .Y(n387) );
  IBUFFX2_HVT U47 ( .A(n241), .Y(n231) );
  MUX21X2_HVT U48 ( .A1(n387), .A2(n386), .S0(n234), .Y(n385) );
  IBUFFX16_HVT U49 ( .A(n264), .Y(n234) );
  MUX21X1_HVT U50 ( .A1(n274), .A2(n272), .S0(n293), .Y(n568) );
  AO21X2_HVT U52 ( .A1(n266), .A2(n281), .A3(n578), .Y(n466) );
  OA21X1_HVT U54 ( .A1(n310), .A2(n249), .A3(n554), .Y(n439) );
  INVX2_HVT U55 ( .A(n269), .Y(n249) );
  INVX2_HVT U60 ( .A(n298), .Y(n297) );
  INVX2_HVT U64 ( .A(in[2]), .Y(n298) );
  MUX21X1_HVT U65 ( .A1(n396), .A2(n405), .S0(in[6]), .Y(out[6]) );
  NBUFFX4_HVT U67 ( .A(n366), .Y(n274) );
  NAND2X0_HVT U70 ( .A1(n286), .A2(n235), .Y(n236) );
  NAND2X0_HVT U71 ( .A1(n472), .A2(n251), .Y(n237) );
  NAND2X0_HVT U72 ( .A1(n236), .A2(n237), .Y(n471) );
  INVX0_HVT U74 ( .A(n251), .Y(n235) );
  MUX21X1_HVT U76 ( .A1(n508), .A2(n507), .S0(n266), .Y(n505) );
  INVX1_HVT U79 ( .A(n298), .Y(n296) );
  INVX1_HVT U81 ( .A(in[6]), .Y(n247) );
  INVX1_HVT U82 ( .A(n294), .Y(n291) );
  INVX1_HVT U88 ( .A(in[1]), .Y(n294) );
  INVX0_HVT U89 ( .A(n294), .Y(n238) );
  INVX0_HVT U91 ( .A(n294), .Y(n239) );
  INVX0_HVT U92 ( .A(n294), .Y(n290) );
  INVX0_HVT U94 ( .A(n376), .Y(n351) );
  INVX1_HVT U95 ( .A(n271), .Y(n241) );
  INVX0_HVT U99 ( .A(n263), .Y(n243) );
  INVX1_HVT U100 ( .A(in[4]), .Y(n367) );
  OA21X2_HVT U102 ( .A1(n258), .A2(n241), .A3(n554), .Y(n414) );
  MUX21X1_HVT U104 ( .A1(n376), .A2(n287), .S0(n241), .Y(n240) );
  INVX0_HVT U106 ( .A(n284), .Y(n365) );
  INVX1_HVT U107 ( .A(n294), .Y(n292) );
  IBUFFX2_HVT U108 ( .A(in[1]), .Y(n295) );
  MUX41X1_HVT U109 ( .A1(n570), .A3(n307), .A2(n325), .A4(n541), .S0(n243), 
        .S1(n305), .Y(n504) );
  IBUFFX2_HVT U111 ( .A(n305), .Y(n302) );
  MUX41X1_HVT U112 ( .A1(n561), .A3(n515), .A2(n559), .A4(n516), .S0(n243), 
        .S1(n241), .Y(n513) );
  MUX21X2_HVT U113 ( .A1(n509), .A2(n499), .S0(n247), .Y(out[1]) );
  IBUFFX2_HVT U114 ( .A(n305), .Y(n304) );
  XNOR2X1_HVT U117 ( .A1(n292), .A2(n297), .Y(n251) );
  INVX1_HVT U118 ( .A(n299), .Y(n248) );
  INVX1_HVT U119 ( .A(n278), .Y(n246) );
  INVX1_HVT U120 ( .A(n277), .Y(n244) );
  XOR2X2_HVT U121 ( .A1(n367), .A2(in[3]), .Y(n578) );
  INVX2_HVT U122 ( .A(n249), .Y(n245) );
  MUX41X1_HVT U124 ( .A1(n385), .A3(n383), .A2(n384), .A4(n382), .S0(n246), 
        .S1(n248), .Y(n381) );
  MUX21X2_HVT U126 ( .A1(n488), .A2(n478), .S0(n247), .Y(out[2]) );
  MUX41X1_HVT U127 ( .A1(n486), .A3(n481), .A2(n482), .A4(n479), .S0(n246), 
        .S1(n248), .Y(n478) );
  MUX41X1_HVT U129 ( .A1(n334), .A3(n443), .A2(n338), .A4(n560), .S0(n243), 
        .S1(n305), .Y(n442) );
  OA21X2_HVT U130 ( .A1(n337), .A2(n298), .A3(n323), .Y(n476) );
  NBUFFX2_HVT U133 ( .A(n296), .Y(n262) );
  MUX41X1_HVT U134 ( .A1(n280), .A3(n357), .A2(n558), .A4(n544), .S0(n249), 
        .S1(n298), .Y(n393) );
  INVX0_HVT U137 ( .A(n578), .Y(n366) );
  INVX0_HVT U138 ( .A(n294), .Y(n293) );
  INVX0_HVT U141 ( .A(n294), .Y(n289) );
  INVX0_HVT U143 ( .A(in[3]), .Y(n363) );
  INVX1_HVT U144 ( .A(n580), .Y(n361) );
  MUX21X1_HVT U145 ( .A1(n254), .A2(n321), .S0(n262), .Y(n453) );
  NBUFFX2_HVT U149 ( .A(n366), .Y(n273) );
  AND2X1_HVT U150 ( .A1(n275), .A2(n530), .Y(n252) );
  MUX21X1_HVT U152 ( .A1(n361), .A2(n364), .S0(n268), .Y(n534) );
  NBUFFX2_HVT U155 ( .A(n580), .Y(n282) );
  MUX21X1_HVT U156 ( .A1(n554), .A2(n475), .S0(n262), .Y(n473) );
  NBUFFX2_HVT U157 ( .A(n580), .Y(n283) );
  MUX21X1_HVT U161 ( .A1(n317), .A2(n362), .S0(n268), .Y(n519) );
  AND2X1_HVT U164 ( .A1(n285), .A2(n514), .Y(n253) );
  MUX21X1_HVT U169 ( .A1(n457), .A2(n458), .S0(n268), .Y(n456) );
  MUX21X1_HVT U170 ( .A1(n462), .A2(n461), .S0(n271), .Y(n458) );
  MUX21X1_HVT U171 ( .A1(n285), .A2(n274), .S0(n290), .Y(n544) );
  MUX21X1_HVT U173 ( .A1(n273), .A2(n277), .S0(n291), .Y(n483) );
  MUX21X1_HVT U175 ( .A1(n446), .A2(n581), .S0(n266), .Y(n445) );
  MUX21X1_HVT U183 ( .A1(n361), .A2(n365), .S0(n238), .Y(n411) );
  MUX21X1_HVT U185 ( .A1(n283), .A2(n578), .S0(n239), .Y(n548) );
  MUX21X1_HVT U187 ( .A1(n364), .A2(n274), .S0(n291), .Y(n423) );
  MUX21X1_HVT U188 ( .A1(n578), .A2(n362), .S0(n291), .Y(n371) );
  MUX21X1_HVT U191 ( .A1(n578), .A2(n365), .S0(n289), .Y(n560) );
  MUX21X1_HVT U192 ( .A1(n578), .A2(n277), .S0(n291), .Y(n511) );
  XOR2X1_HVT U194 ( .A1(n578), .A2(n291), .Y(n540) );
  MUX21X1_HVT U196 ( .A1(n272), .A2(n578), .S0(n238), .Y(n374) );
  MUX21X1_HVT U198 ( .A1(n364), .A2(n361), .S0(n238), .Y(n547) );
  MUX21X1_HVT U200 ( .A1(n272), .A2(n365), .S0(n290), .Y(n545) );
  MUX21X1_HVT U202 ( .A1(n277), .A2(n361), .S0(n238), .Y(n556) );
  MUX21X1_HVT U206 ( .A1(n332), .A2(n450), .S0(n265), .Y(n449) );
  MUX21X1_HVT U207 ( .A1(n356), .A2(n281), .S0(n270), .Y(n450) );
  MUX21X1_HVT U209 ( .A1(n466), .A2(n467), .S0(n270), .Y(n465) );
  MUX21X1_HVT U210 ( .A1(n309), .A2(n335), .S0(n262), .Y(n467) );
  MUX21X1_HVT U211 ( .A1(n282), .A2(n281), .S0(n238), .Y(n498) );
  NAND2X0_HVT U213 ( .A1(n276), .A2(n363), .Y(n580) );
  MUX21X1_HVT U217 ( .A1(n361), .A2(n276), .S0(n289), .Y(n372) );
  NBUFFX2_HVT U219 ( .A(n583), .Y(n284) );
  INVX1_HVT U221 ( .A(n287), .Y(n364) );
  MUX21X1_HVT U222 ( .A1(n364), .A2(n272), .S0(n290), .Y(n551) );
  MUX21X1_HVT U223 ( .A1(n308), .A2(n463), .S0(n263), .Y(n462) );
  MUX21X1_HVT U224 ( .A1(n276), .A2(n272), .S0(n289), .Y(n463) );
  NBUFFX2_HVT U225 ( .A(n583), .Y(n285) );
  XOR2X1_HVT U226 ( .A1(n292), .A2(n362), .Y(n541) );
  MUX21X1_HVT U227 ( .A1(n272), .A2(n288), .S0(n293), .Y(n398) );
  MUX21X1_HVT U228 ( .A1(n287), .A2(n285), .S0(n292), .Y(n399) );
  MUX21X1_HVT U229 ( .A1(n362), .A2(n361), .S0(n239), .Y(n566) );
  INVX1_HVT U230 ( .A(n575), .Y(n362) );
  MUX21X1_HVT U231 ( .A1(n286), .A2(n280), .S0(n293), .Y(n570) );
  MUX21X1_HVT U232 ( .A1(n283), .A2(n288), .S0(n293), .Y(n493) );
  MUX21X1_HVT U233 ( .A1(n272), .A2(n364), .S0(n292), .Y(n574) );
  MUX21X1_HVT U234 ( .A1(n282), .A2(n272), .S0(n293), .Y(n573) );
  MUX21X1_HVT U235 ( .A1(n333), .A2(n570), .S0(n266), .Y(n487) );
  NBUFFX2_HVT U236 ( .A(n583), .Y(n286) );
  MUX21X1_HVT U237 ( .A1(n272), .A2(n277), .S0(n293), .Y(n395) );
  XOR2X1_HVT U238 ( .A1(n284), .A2(n290), .Y(n538) );
  XNOR2X1_HVT U239 ( .A1(n282), .A2(n292), .Y(n254) );
  MUX21X1_HVT U240 ( .A1(n287), .A2(n280), .S0(n289), .Y(n554) );
  MUX21X1_HVT U241 ( .A1(n284), .A2(n276), .S0(n290), .Y(n378) );
  MUX21X1_HVT U242 ( .A1(n284), .A2(n282), .S0(n292), .Y(n370) );
  XNOR2X1_HVT U243 ( .A1(n287), .A2(n239), .Y(n255) );
  AND2X1_HVT U244 ( .A1(n289), .A2(n365), .Y(n256) );
  MUX21X1_HVT U245 ( .A1(n280), .A2(n272), .S0(n239), .Y(n376) );
  AND2X1_HVT U246 ( .A1(n584), .A2(n474), .Y(n257) );
  MUX21X1_HVT U247 ( .A1(n281), .A2(n276), .S0(n239), .Y(n516) );
  MUX21X1_HVT U248 ( .A1(n281), .A2(n288), .S0(n265), .Y(n460) );
  XOR2X1_HVT U249 ( .A1(n276), .A2(n292), .Y(n559) );
  NBUFFX2_HVT U250 ( .A(n301), .Y(n271) );
  NBUFFX2_HVT U251 ( .A(n301), .Y(n270) );
  NBUFFX2_HVT U252 ( .A(n363), .Y(n272) );
  NBUFFX2_HVT U253 ( .A(n300), .Y(n268) );
  NBUFFX2_HVT U254 ( .A(n296), .Y(n263) );
  NBUFFX2_HVT U255 ( .A(n297), .Y(n265) );
  NBUFFX2_HVT U256 ( .A(n297), .Y(n264) );
  NBUFFX2_HVT U257 ( .A(n300), .Y(n267) );
  NBUFFX2_HVT U258 ( .A(n297), .Y(n266) );
  NBUFFX2_HVT U259 ( .A(n296), .Y(n261) );
  MUX21X1_HVT U260 ( .A1(n402), .A2(n403), .S0(n264), .Y(n401) );
  MUX21X1_HVT U261 ( .A1(n501), .A2(n279), .S0(n270), .Y(n403) );
  MUX21X1_HVT U262 ( .A1(n485), .A2(n332), .S0(n265), .Y(n482) );
  MUX21X1_HVT U263 ( .A1(n523), .A2(n525), .S0(n264), .Y(n522) );
  XOR2X1_HVT U264 ( .A1(n293), .A2(in[3]), .Y(n539) );
  MUX21X1_HVT U265 ( .A1(n280), .A2(n275), .S0(n291), .Y(n480) );
  MUX21X1_HVT U266 ( .A1(n434), .A2(n435), .S0(n266), .Y(n432) );
  MUX21X1_HVT U267 ( .A1(n353), .A2(n362), .S0(n270), .Y(n435) );
  MUX21X1_HVT U268 ( .A1(n564), .A2(n281), .S0(n271), .Y(n508) );
  MUX21X1_HVT U269 ( .A1(n415), .A2(n414), .S0(n265), .Y(n413) );
  MUX21X1_HVT U270 ( .A1(n281), .A2(n351), .S0(n271), .Y(n415) );
  AND2X1_HVT U271 ( .A1(n275), .A2(n295), .Y(n258) );
  MUX21X1_HVT U272 ( .A1(n440), .A2(n439), .S0(n265), .Y(n438) );
  MUX21X1_HVT U273 ( .A1(n556), .A2(n312), .S0(n271), .Y(n440) );
  MUX21X1_HVT U274 ( .A1(n362), .A2(n365), .S0(n291), .Y(n420) );
  NAND2X0_HVT U275 ( .A1(n279), .A2(n277), .Y(n583) );
  NBUFFX2_HVT U276 ( .A(n367), .Y(n277) );
  NBUFFX2_HVT U277 ( .A(n584), .Y(n287) );
  MUX21X1_HVT U278 ( .A1(n365), .A2(n279), .S0(n291), .Y(n565) );
  MUX21X1_HVT U279 ( .A1(n279), .A2(n361), .S0(n239), .Y(n546) );
  MUX21X1_HVT U280 ( .A1(n336), .A2(n582), .S0(n263), .Y(n477) );
  MUX21X1_HVT U281 ( .A1(n428), .A2(n429), .S0(n266), .Y(n427) );
  MUX21X1_HVT U282 ( .A1(n430), .A2(n286), .S0(n259), .Y(n429) );
  MUX21X1_HVT U283 ( .A1(n547), .A2(n354), .S0(n269), .Y(n428) );
  MUX21X1_HVT U284 ( .A1(n567), .A2(n334), .S0(n263), .Y(n452) );
  MUX21X1_HVT U285 ( .A1(n582), .A2(n294), .S0(n264), .Y(n459) );
  MUX21X1_HVT U286 ( .A1(n535), .A2(n536), .S0(n269), .Y(n533) );
  MUX21X1_HVT U287 ( .A1(n279), .A2(n550), .S0(n268), .Y(n536) );
  XOR2X1_HVT U288 ( .A1(n238), .A2(n267), .Y(n542) );
  MUX21X1_HVT U289 ( .A1(n279), .A2(n362), .S0(n289), .Y(n375) );
  MUX21X1_HVT U290 ( .A1(n342), .A2(n359), .S0(n270), .Y(n391) );
  NBUFFX2_HVT U291 ( .A(n575), .Y(n280) );
  MUX21X1_HVT U292 ( .A1(n555), .A2(n379), .S0(n269), .Y(n373) );
  MUX21X1_HVT U293 ( .A1(n283), .A2(n279), .S0(n293), .Y(n576) );
  MUX21X1_HVT U294 ( .A1(n329), .A2(n555), .S0(n263), .Y(n455) );
  MUX21X1_HVT U295 ( .A1(n319), .A2(n295), .S0(n268), .Y(n521) );
  MUX21X1_HVT U296 ( .A1(n286), .A2(n496), .S0(n259), .Y(n495) );
  MUX21X1_HVT U297 ( .A1(n279), .A2(n276), .S0(n271), .Y(n496) );
  NBUFFX2_HVT U298 ( .A(n584), .Y(n288) );
  NBUFFX2_HVT U299 ( .A(n367), .Y(n276) );
  NBUFFX2_HVT U300 ( .A(n575), .Y(n281) );
  XNOR2X1_HVT U301 ( .A1(n249), .A2(n292), .Y(n259) );
  AND2X1_HVT U302 ( .A1(n363), .A2(n295), .Y(n260) );
  NBUFFX2_HVT U303 ( .A(in[5]), .Y(n300) );
  NBUFFX2_HVT U304 ( .A(in[5]), .Y(n299) );
  MUX21X1_HVT U305 ( .A1(n391), .A2(n390), .S0(n264), .Y(n389) );
  MUX21X1_HVT U306 ( .A1(n494), .A2(n495), .S0(n266), .Y(n492) );
  MUX21X1_HVT U307 ( .A1(n533), .A2(n537), .S0(n265), .Y(n532) );
  MUX21X1_HVT U308 ( .A1(n527), .A2(n529), .S0(n264), .Y(n526) );
  MUX21X1_HVT U309 ( .A1(n361), .A2(n244), .S0(n290), .Y(n553) );
  NAND2X0_HVT U310 ( .A1(in[3]), .A2(in[4]), .Y(n584) );
  MUX21X1_HVT U311 ( .A1(n244), .A2(n578), .S0(n239), .Y(n377) );
  MUX21X1_HVT U312 ( .A1(n244), .A2(n364), .S0(n238), .Y(n549) );
  MUX21X1_HVT U313 ( .A1(n244), .A2(n362), .S0(n292), .Y(n567) );
  NAND2X0_HVT U314 ( .A1(in[4]), .A2(n363), .Y(n575) );
  MUX21X1_HVT U315 ( .A1(n244), .A2(n286), .S0(n289), .Y(n564) );
  MUX21X1_HVT U316 ( .A1(n244), .A2(n280), .S0(n290), .Y(n369) );
  MUX21X1_HVT U317 ( .A1(n288), .A2(n244), .S0(n290), .Y(n557) );
  MUX21X1_HVT U318 ( .A1(n279), .A2(n244), .S0(n262), .Y(n472) );
  MUX21X1_HVT U319 ( .A1(n244), .A2(n584), .S0(n291), .Y(n368) );
  MUX21X1_HVT U320 ( .A1(n272), .A2(n244), .S0(n289), .Y(n555) );
  NBUFFX2_HVT U321 ( .A(in[3]), .Y(n279) );
  NBUFFX2_HVT U322 ( .A(in[0]), .Y(n278) );
  INVX0_HVT U323 ( .A(n563), .Y(n306) );
  INVX0_HVT U324 ( .A(n561), .Y(n307) );
  INVX0_HVT U325 ( .A(n552), .Y(n308) );
  INVX0_HVT U326 ( .A(n550), .Y(n309) );
  INVX0_HVT U327 ( .A(n417), .Y(n310) );
  INVX0_HVT U328 ( .A(n380), .Y(n311) );
  INVX0_HVT U329 ( .A(n582), .Y(n312) );
  INVX0_HVT U330 ( .A(n569), .Y(n313) );
  INVX0_HVT U331 ( .A(n581), .Y(n314) );
  INVX0_HVT U332 ( .A(n579), .Y(n315) );
  INVX0_HVT U333 ( .A(n577), .Y(n316) );
  INVX0_HVT U334 ( .A(n576), .Y(n317) );
  INVX0_HVT U335 ( .A(n574), .Y(n318) );
  INVX0_HVT U336 ( .A(n573), .Y(n319) );
  INVX0_HVT U337 ( .A(n570), .Y(n320) );
  INVX0_HVT U338 ( .A(n567), .Y(n322) );
  INVX0_HVT U339 ( .A(n566), .Y(n323) );
  INVX0_HVT U340 ( .A(n565), .Y(n324) );
  INVX0_HVT U341 ( .A(n564), .Y(n325) );
  INVX0_HVT U342 ( .A(n562), .Y(n326) );
  INVX0_HVT U343 ( .A(n560), .Y(n327) );
  INVX0_HVT U344 ( .A(n559), .Y(n328) );
  INVX0_HVT U345 ( .A(n557), .Y(n329) );
  INVX0_HVT U346 ( .A(n556), .Y(n330) );
  INVX0_HVT U347 ( .A(n555), .Y(n331) );
  INVX0_HVT U348 ( .A(n373), .Y(n332) );
  INVX0_HVT U349 ( .A(n554), .Y(n333) );
  INVX0_HVT U350 ( .A(n553), .Y(n334) );
  INVX0_HVT U351 ( .A(n551), .Y(n335) );
  INVX0_HVT U352 ( .A(n549), .Y(n336) );
  INVX0_HVT U353 ( .A(n548), .Y(n337) );
  INVX0_HVT U354 ( .A(n547), .Y(n338) );
  INVX0_HVT U355 ( .A(n546), .Y(n339) );
  INVX0_HVT U356 ( .A(n545), .Y(n340) );
  INVX0_HVT U357 ( .A(n544), .Y(n341) );
  INVX0_HVT U358 ( .A(n543), .Y(n342) );
  INVX0_HVT U359 ( .A(n514), .Y(n343) );
  INVX0_HVT U360 ( .A(n572), .Y(n344) );
  INVX0_HVT U361 ( .A(n474), .Y(n345) );
  INVX0_HVT U362 ( .A(n379), .Y(n346) );
  INVX0_HVT U363 ( .A(n530), .Y(n347) );
  INVX0_HVT U364 ( .A(n433), .Y(n348) );
  INVX0_HVT U365 ( .A(n378), .Y(n349) );
  INVX0_HVT U366 ( .A(n377), .Y(n350) );
  INVX0_HVT U367 ( .A(n375), .Y(n352) );
  INVX0_HVT U368 ( .A(n374), .Y(n353) );
  INVX0_HVT U369 ( .A(n493), .Y(n354) );
  INVX0_HVT U370 ( .A(n483), .Y(n355) );
  INVX0_HVT U371 ( .A(n372), .Y(n356) );
  INVX0_HVT U372 ( .A(n371), .Y(n357) );
  INVX0_HVT U373 ( .A(n370), .Y(n358) );
  INVX0_HVT U374 ( .A(n369), .Y(n359) );
  INVX0_HVT U375 ( .A(n368), .Y(n360) );
endmodule

