
module inv_Mix_Column ( in, out1 );
  input [127:0] in;
  output [127:0] out1;
  wire   n50, n51, n53, n54, n55, n57, n59, n60, n61, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n92, n93, n96, n97, n98, n99,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n122, n123, n124,
         n125, n126, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n159, n160, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n194, n195, n196, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n208, n209, n210, n212,
         n213, n214, n215, n216, n217, n218, n219, n221, n222, n224, n225,
         n226, n228, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n295, n296, n297,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n311,
         n312, n313, n314, n316, n317, n318, n319, n320, n321, n323, n324,
         n325, n326, n327, n328, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n350, n351, n354, n355, n356, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n386,
         n387, n388, n390, n391, n392, n393, n394, n395, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n410, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n433, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n450, n451, n452, n453, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n502, n503, n505, n506, n507, n509, n510, n511,
         n512, n513, n514, n515, n516, n518, n519, n520, n521, n523, n524,
         n525, n526, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n555, n556, n557, n558, n559, n560,
         n561, n563, n564, n565, n566, n567, n568, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n596, n597, n600, n601,
         n602, n603, n605, n606, n607, n608, n609, n610, n613, n614, n615,
         n617, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n52, n56, n58, n62, n73, n91, n94,
         n95, n100, n111, n121, n127, n142, n143, n144, n158, n161, n192, n193,
         n197, n207, n211, n220, n223, n227, n229, n247, n260, n261, n294,
         n298, n299, n310, n315, n322, n329, n349, n352, n353, n357, n384,
         n385, n389, n396, n409, n411, n432, n434, n449, n454, n466, n480,
         n490, n491, n501, n504, n508, n517, n522, n527, n553, n554, n562,
         n569, n570, n571, n594, n595, n598, n599, n604, n611, n612, n616,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550;

  XNOR3X1_HVT U506 ( .A1(n77), .A2(n78), .A3(n79), .Y(out1[95]) );
  XNOR3X1_HVT U534 ( .A1(n173), .A2(n174), .A3(n175), .Y(out1[80]) );
  XNOR3X1_HVT U537 ( .A1(n178), .A2(n179), .A3(n180), .Y(out1[7]) );
  XNOR3X1_HVT U539 ( .A1(n183), .A2(n184), .A3(n185), .Y(out1[79]) );
  XNOR3X1_HVT U554 ( .A1(n183), .A2(n213), .A3(n214), .Y(out1[71]) );
  XNOR3X1_HVT U569 ( .A1(n230), .A2(n165), .A3(n208), .Y(out1[65]) );
  XNOR3X1_HVT U572 ( .A1(n231), .A2(n128), .A3(n212), .Y(out1[64]) );
  XNOR3X1_HVT U592 ( .A1(n281), .A2(n282), .A3(n283), .Y(out1[55]) );
  XNOR3X1_HVT U605 ( .A1(n338), .A2(n339), .A3(n340), .Y(out1[48]) );
  XNOR3X1_HVT U609 ( .A1(n286), .A2(n1526), .A3(n280), .Y(n345) );
  XNOR3X1_HVT U621 ( .A1(n371), .A2(n342), .A3(n372), .Y(out1[40]) );
  XNOR3X1_HVT U625 ( .A1(n343), .A2(n379), .A3(n380), .Y(out1[39]) );
  XNOR3X1_HVT U641 ( .A1(n393), .A2(n284), .A3(n372), .Y(out1[32]) );
  XNOR3X1_HVT U653 ( .A1(n425), .A2(n426), .A3(n427), .Y(out1[26]) );
  XNOR3X1_HVT U657 ( .A1(n436), .A2(n437), .A3(n438), .Y(out1[24]) );
  XNOR3X1_HVT U670 ( .A1(n475), .A2(n476), .A3(n427), .Y(out1[18]) );
  XNOR3X1_HVT U674 ( .A1(n481), .A2(n181), .A3(n438), .Y(out1[16]) );
  XNOR3X1_HVT U677 ( .A1(n437), .A2(n484), .A3(n485), .Y(out1[15]) );
  XNOR3X1_HVT U685 ( .A1(n494), .A2(n495), .A3(n496), .Y(out1[127]) );
  XNOR3X1_HVT U698 ( .A1(n532), .A2(n533), .A3(n534), .Y(out1[120]) );
  XNOR3X1_HVT U702 ( .A1(n537), .A2(n538), .A3(n539), .Y(out1[119]) );
  XNOR3X1_HVT U715 ( .A1(n584), .A2(n585), .A3(n534), .Y(out1[112]) );
  XNOR3X1_HVT U743 ( .A1(n482), .A2(n440), .A3(n617), .Y(out1[0]) );
  INVX1_HVT U1 ( .A(in[39]), .Y(n1341) );
  INVX0_HVT U2 ( .A(n50), .Y(n1274) );
  INVX0_HVT U3 ( .A(n369), .Y(n1451) );
  XOR3X2_HVT U4 ( .A1(n1172), .A2(n1), .A3(n265), .Y(n658) );
  IBUFFX16_HVT U5 ( .A(n25), .Y(n1) );
  INVX0_HVT U6 ( .A(in[63]), .Y(n1452) );
  INVX0_HVT U7 ( .A(in[38]), .Y(n1193) );
  INVX1_HVT U8 ( .A(in[93]), .Y(n1287) );
  XNOR3X1_HVT U9 ( .A1(n205), .A2(n1035), .A3(n163), .Y(n933) );
  INVX0_HVT U10 ( .A(n515), .Y(n2) );
  INVX1_HVT U11 ( .A(n2), .Y(n3) );
  XOR3X2_HVT U12 ( .A1(n4), .A2(n5), .A3(n276), .Y(n367) );
  IBUFFX16_HVT U13 ( .A(n370), .Y(n4) );
  IBUFFX16_HVT U14 ( .A(n1401), .Y(n5) );
  INVX1_HVT U15 ( .A(n597), .Y(n1423) );
  XNOR2X1_HVT U16 ( .A1(n514), .A2(n768), .Y(n596) );
  INVX1_HVT U17 ( .A(in[118]), .Y(n1142) );
  INVX0_HVT U18 ( .A(n1155), .Y(n1167) );
  NBUFFX4_HVT U19 ( .A(in[118]), .Y(n1441) );
  IBUFFX2_HVT U20 ( .A(n560), .Y(n6) );
  INVX1_HVT U21 ( .A(n6), .Y(n7) );
  XOR3X2_HVT U22 ( .A1(n395), .A2(n1145), .A3(n401), .Y(n398) );
  INVX1_HVT U23 ( .A(n1007), .Y(n8) );
  INVX2_HVT U24 ( .A(n274), .Y(n1007) );
  NAND2X0_HVT U25 ( .A1(n647), .A2(n648), .Y(n9) );
  XOR2X2_HVT U26 ( .A1(n318), .A2(in[50]), .Y(n267) );
  INVX0_HVT U27 ( .A(n225), .Y(n1372) );
  INVX2_HVT U28 ( .A(in[15]), .Y(n991) );
  INVX0_HVT U29 ( .A(in[65]), .Y(n357) );
  IBUFFX2_HVT U30 ( .A(n1531), .Y(n11) );
  INVX0_HVT U31 ( .A(n1340), .Y(n10) );
  XOR3X2_HVT U32 ( .A1(n341), .A2(n11), .A3(n342), .Y(n279) );
  INVX1_HVT U33 ( .A(n141), .Y(n1104) );
  INVX0_HVT U34 ( .A(in[24]), .Y(n1321) );
  XNOR2X2_HVT U35 ( .A1(n709), .A2(n1521), .Y(n435) );
  IBUFFX2_HVT U36 ( .A(n1521), .Y(n992) );
  IBUFFX2_HVT U37 ( .A(in[104]), .Y(n1173) );
  NBUFFX4_HVT U38 ( .A(n938), .Y(n45) );
  INVX1_HVT U39 ( .A(n1374), .Y(n12) );
  INVX1_HVT U40 ( .A(n169), .Y(n1374) );
  INVX0_HVT U41 ( .A(n330), .Y(n1114) );
  INVX1_HVT U42 ( .A(n858), .Y(n13) );
  OR2X2_HVT U43 ( .A1(in[121]), .A2(in[126]), .Y(n1092) );
  INVX1_HVT U44 ( .A(n410), .Y(n1005) );
  INVX1_HVT U45 ( .A(n1324), .Y(n111) );
  INVX1_HVT U46 ( .A(n456), .Y(n1210) );
  XNOR2X2_HVT U47 ( .A1(n474), .A2(n473), .Y(n376) );
  NAND2X0_HVT U48 ( .A1(n194), .A2(n1426), .Y(n16) );
  NAND2X0_HVT U49 ( .A1(n14), .A2(n15), .Y(n17) );
  NAND2X0_HVT U50 ( .A1(n16), .A2(n17), .Y(n145) );
  INVX0_HVT U51 ( .A(n194), .Y(n14) );
  IBUFFX2_HVT U52 ( .A(n1426), .Y(n15) );
  INVX0_HVT U53 ( .A(n145), .Y(n1116) );
  XNOR3X1_HVT U54 ( .A1(n768), .A2(n561), .A3(n7), .Y(n1475) );
  IBUFFX2_HVT U55 ( .A(in[75]), .Y(n18) );
  INVX1_HVT U56 ( .A(n18), .Y(n19) );
  INVX1_HVT U57 ( .A(n1529), .Y(n247) );
  XOR3X2_HVT U58 ( .A1(n1465), .A2(n506), .A3(n507), .Y(n505) );
  INVX1_HVT U59 ( .A(in[117]), .Y(n1124) );
  XOR3X2_HVT U60 ( .A1(n1464), .A2(n550), .A3(n970), .Y(n549) );
  NBUFFX2_HVT U61 ( .A(n366), .Y(n20) );
  NAND2X0_HVT U62 ( .A1(n1477), .A2(n1476), .Y(n23) );
  NAND2X0_HVT U63 ( .A1(n21), .A2(n22), .Y(n24) );
  NAND2X0_HVT U64 ( .A1(n23), .A2(n24), .Y(out1[108]) );
  INVX0_HVT U65 ( .A(n1477), .Y(n21) );
  INVX0_HVT U66 ( .A(n1476), .Y(n22) );
  XOR3X2_HVT U67 ( .A1(n596), .A2(n1382), .A3(n601), .Y(n1477) );
  INVX1_HVT U68 ( .A(in[69]), .Y(n1201) );
  AND2X1_HVT U69 ( .A1(n260), .A2(n261), .Y(n25) );
  INVX0_HVT U70 ( .A(in[42]), .Y(n229) );
  INVX0_HVT U71 ( .A(in[46]), .Y(n1528) );
  XOR2X2_HVT U72 ( .A1(n326), .A2(in[12]), .Y(n399) );
  XNOR2X1_HVT U73 ( .A1(in[27]), .A2(n979), .Y(n326) );
  NBUFFX2_HVT U74 ( .A(n148), .Y(n26) );
  XOR2X2_HVT U75 ( .A1(n719), .A2(n1437), .Y(n416) );
  INVX1_HVT U76 ( .A(n408), .Y(n751) );
  XNOR2X1_HVT U77 ( .A1(n1357), .A2(in[61]), .Y(n275) );
  XNOR2X2_HVT U78 ( .A1(n1438), .A2(n1524), .Y(n433) );
  NBUFFX2_HVT U79 ( .A(n273), .Y(n27) );
  NAND2X0_HVT U80 ( .A1(n303), .A2(n1053), .Y(n30) );
  NAND2X0_HVT U81 ( .A1(n28), .A2(n29), .Y(n31) );
  NAND2X0_HVT U82 ( .A1(n30), .A2(n31), .Y(n293) );
  INVX0_HVT U83 ( .A(n303), .Y(n28) );
  INVX0_HVT U84 ( .A(n1053), .Y(n29) );
  INVX1_HVT U85 ( .A(n1359), .Y(n1053) );
  XNOR2X2_HVT U86 ( .A1(n148), .A2(in[92]), .Y(n89) );
  INVX0_HVT U87 ( .A(n228), .Y(n1164) );
  NBUFFX4_HVT U88 ( .A(n559), .Y(n768) );
  INVX1_HVT U89 ( .A(n1374), .Y(n39) );
  XOR3X1_HVT U90 ( .A1(n82), .A2(n32), .A3(n84), .Y(out1[94]) );
  IBUFFX16_HVT U91 ( .A(n83), .Y(n32) );
  NAND2X0_HVT U92 ( .A1(n537), .A2(n34), .Y(n35) );
  NAND2X0_HVT U93 ( .A1(n33), .A2(n494), .Y(n36) );
  NAND2X0_HVT U94 ( .A1(n35), .A2(n36), .Y(n588) );
  IBUFFX2_HVT U95 ( .A(n537), .Y(n33) );
  INVX0_HVT U96 ( .A(n494), .Y(n34) );
  XNOR2X2_HVT U97 ( .A1(in[124]), .A2(n1550), .Y(n537) );
  INVX1_HVT U98 ( .A(n798), .Y(n37) );
  INVX2_HVT U99 ( .A(n593), .Y(n798) );
  INVX1_HVT U100 ( .A(in[46]), .Y(n1244) );
  INVX1_HVT U101 ( .A(n979), .Y(n1247) );
  NAND2X0_HVT U102 ( .A1(n1211), .A2(n94), .Y(n38) );
  XOR3X2_HVT U103 ( .A1(n641), .A2(n39), .A3(n117), .Y(n167) );
  XNOR2X2_HVT U104 ( .A1(n1053), .A2(n40), .Y(n288) );
  IBUFFX16_HVT U105 ( .A(in[36]), .Y(n40) );
  INVX1_HVT U106 ( .A(in[45]), .Y(n1337) );
  INVX0_HVT U107 ( .A(n600), .Y(n1382) );
  IBUFFX2_HVT U108 ( .A(in[41]), .Y(n1400) );
  NAND2X0_HVT U109 ( .A1(in[41]), .A2(n1528), .Y(n43) );
  NAND2X0_HVT U110 ( .A1(n41), .A2(n42), .Y(n44) );
  NAND2X0_HVT U111 ( .A1(n43), .A2(n44), .Y(n362) );
  INVX0_HVT U112 ( .A(in[41]), .Y(n41) );
  INVX0_HVT U113 ( .A(n1528), .Y(n42) );
  INVX1_HVT U114 ( .A(in[126]), .Y(n858) );
  XNOR3X2_HVT U115 ( .A1(n45), .A2(n49), .A3(n235), .Y(n371) );
  INVX1_HVT U116 ( .A(in[47]), .Y(n1529) );
  XOR3X2_HVT U117 ( .A1(n966), .A2(n47), .A3(n46), .Y(n1350) );
  IBUFFX16_HVT U118 ( .A(n997), .Y(n46) );
  NAND2X0_HVT U119 ( .A1(n1249), .A2(n1243), .Y(n47) );
  INVX0_HVT U120 ( .A(n1425), .Y(n48) );
  INVX0_HVT U121 ( .A(n155), .Y(n1425) );
  INVX2_HVT U122 ( .A(n1090), .Y(n1315) );
  INVX0_HVT U123 ( .A(in[46]), .Y(n49) );
  XNOR2X2_HVT U124 ( .A1(n824), .A2(n628), .Y(n341) );
  INVX1_HVT U125 ( .A(n448), .Y(n52) );
  INVX1_HVT U126 ( .A(n52), .Y(n56) );
  XNOR2X1_HVT U127 ( .A1(in[112]), .A2(n695), .Y(n535) );
  INVX1_HVT U128 ( .A(n511), .Y(n1042) );
  INVX0_HVT U129 ( .A(in[45]), .Y(n878) );
  XOR3X2_HVT U130 ( .A1(n58), .A2(n62), .A3(n273), .Y(n332) );
  IBUFFX16_HVT U131 ( .A(n333), .Y(n58) );
  IBUFFX16_HVT U132 ( .A(n1401), .Y(n62) );
  IBUFFX2_HVT U133 ( .A(n581), .Y(n1128) );
  INVX1_HVT U134 ( .A(n1518), .Y(n197) );
  IBUFFX2_HVT U135 ( .A(in[8]), .Y(n73) );
  INVX1_HVT U136 ( .A(n73), .Y(n91) );
  IBUFFX2_HVT U137 ( .A(n226), .Y(n639) );
  XOR3X2_HVT U138 ( .A1(n301), .A2(n383), .A3(n928), .Y(n1450) );
  XNOR2X2_HVT U139 ( .A1(n154), .A2(in[83]), .Y(n101) );
  XNOR2X1_HVT U140 ( .A1(n525), .A2(n574), .Y(n528) );
  NAND2X0_HVT U141 ( .A1(n1101), .A2(n1100), .Y(n94) );
  XOR3X2_HVT U142 ( .A1(n497), .A2(n466), .A3(n609), .Y(out1[104]) );
  INVX2_HVT U143 ( .A(in[95]), .Y(n1541) );
  INVX2_HVT U144 ( .A(n1171), .Y(n942) );
  XNOR2X2_HVT U145 ( .A1(n96), .A2(n1324), .Y(n95) );
  INVX8_HVT U146 ( .A(n95), .Y(n82) );
  INVX0_HVT U147 ( .A(in[119]), .Y(n1549) );
  XOR3X2_HVT U148 ( .A1(n20), .A2(n1400), .A3(n270), .Y(n363) );
  XNOR2X2_HVT U149 ( .A1(n778), .A2(n274), .Y(n270) );
  NBUFFX4_HVT U150 ( .A(n1452), .Y(n1358) );
  NAND2X0_HVT U151 ( .A1(n745), .A2(n746), .Y(n100) );
  XOR3X2_HVT U152 ( .A1(n111), .A2(n80), .A3(n81), .Y(n79) );
  NBUFFX2_HVT U153 ( .A(in[110]), .Y(n121) );
  INVX0_HVT U154 ( .A(n1286), .Y(n807) );
  IBUFFX2_HVT U155 ( .A(n1096), .Y(n127) );
  INVX1_HVT U156 ( .A(n127), .Y(n142) );
  IBUFFX2_HVT U157 ( .A(n224), .Y(n143) );
  INVX0_HVT U158 ( .A(n143), .Y(n144) );
  IBUFFX2_HVT U159 ( .A(in[81]), .Y(n158) );
  INVX1_HVT U160 ( .A(n158), .Y(n161) );
  IBUFFX2_HVT U161 ( .A(n102), .Y(n1504) );
  INVX0_HVT U162 ( .A(in[2]), .Y(n1026) );
  XNOR2X2_HVT U163 ( .A1(n530), .A2(n1089), .Y(n579) );
  NAND2X0_HVT U164 ( .A1(n299), .A2(n310), .Y(n192) );
  XOR3X2_HVT U165 ( .A1(n1419), .A2(n89), .A3(n775), .Y(n88) );
  INVX1_HVT U166 ( .A(n251), .Y(n1359) );
  IBUFFX2_HVT U167 ( .A(n1097), .Y(n193) );
  INVX1_HVT U168 ( .A(in[100]), .Y(n1097) );
  INVX1_HVT U169 ( .A(n783), .Y(n1388) );
  XOR3X2_HVT U170 ( .A1(n197), .A2(n444), .A3(n182), .Y(n485) );
  NAND2X0_HVT U171 ( .A1(n352), .A2(n353), .Y(n207) );
  INVX0_HVT U172 ( .A(in[53]), .Y(n1530) );
  XNOR2X2_HVT U173 ( .A1(n1009), .A2(in[53]), .Y(n282) );
  INVX1_HVT U174 ( .A(in[53]), .Y(n1343) );
  XOR3X2_HVT U175 ( .A1(n220), .A2(n568), .A3(n211), .Y(n1469) );
  IBUFFX16_HVT U176 ( .A(n60), .Y(n211) );
  NAND2X0_HVT U177 ( .A1(n654), .A2(n655), .Y(n220) );
  XOR3X2_HVT U178 ( .A1(n223), .A2(n443), .A3(n394), .Y(n442) );
  IBUFFX16_HVT U179 ( .A(n1402), .Y(n223) );
  IBUFFX2_HVT U180 ( .A(n1283), .Y(n953) );
  INVX0_HVT U181 ( .A(n1248), .Y(n227) );
  NAND2X0_HVT U182 ( .A1(in[42]), .A2(n1529), .Y(n260) );
  NAND2X0_HVT U183 ( .A1(n229), .A2(n247), .Y(n261) );
  NAND2X0_HVT U184 ( .A1(n260), .A2(n261), .Y(n311) );
  NBUFFX16_HVT U185 ( .A(n414), .Y(n927) );
  INVX2_HVT U186 ( .A(in[71]), .Y(n1535) );
  XNOR2X2_HVT U187 ( .A1(n1300), .A2(n1543), .Y(n560) );
  IBUFFX2_HVT U188 ( .A(n1543), .Y(n1293) );
  XOR3X1_HVT U189 ( .A1(n741), .A2(n1500), .A3(n138), .Y(out1[85]) );
  INVX1_HVT U190 ( .A(n952), .Y(n737) );
  INVX1_HVT U191 ( .A(in[49]), .Y(n1012) );
  NAND2X0_HVT U192 ( .A1(n728), .A2(n727), .Y(n299) );
  NAND2X0_HVT U193 ( .A1(n294), .A2(n298), .Y(n310) );
  NAND2X0_HVT U194 ( .A1(n299), .A2(n310), .Y(n548) );
  INVX1_HVT U195 ( .A(n558), .Y(n294) );
  INVX0_HVT U196 ( .A(n727), .Y(n298) );
  IBUFFX2_HVT U197 ( .A(n1078), .Y(n727) );
  INVX1_HVT U198 ( .A(in[54]), .Y(n1314) );
  XOR3X2_HVT U199 ( .A1(n315), .A2(n181), .A3(n182), .Y(n180) );
  IBUFFX16_HVT U200 ( .A(n1277), .Y(n315) );
  INVX1_HVT U201 ( .A(n1242), .Y(n1550) );
  INVX1_HVT U202 ( .A(n1201), .Y(n1183) );
  INVX1_HVT U203 ( .A(n786), .Y(n322) );
  IBUFFX2_HVT U204 ( .A(n1108), .Y(n786) );
  INVX1_HVT U205 ( .A(n1535), .Y(n994) );
  NAND2X0_HVT U206 ( .A1(n1269), .A2(in[51]), .Y(n352) );
  NAND2X0_HVT U207 ( .A1(n329), .A2(n349), .Y(n353) );
  NAND2X0_HVT U208 ( .A1(n352), .A2(n353), .Y(n1275) );
  INVX1_HVT U209 ( .A(n1269), .Y(n329) );
  IBUFFX2_HVT U210 ( .A(in[51]), .Y(n349) );
  NAND2X0_HVT U211 ( .A1(in[65]), .A2(n396), .Y(n385) );
  NAND2X0_HVT U212 ( .A1(n357), .A2(n384), .Y(n389) );
  NAND2X0_HVT U213 ( .A1(n385), .A2(n389), .Y(n226) );
  INVX1_HVT U214 ( .A(in[70]), .Y(n384) );
  INVX0_HVT U215 ( .A(n384), .Y(n396) );
  INVX1_HVT U216 ( .A(n1527), .Y(n1342) );
  NAND2X0_HVT U217 ( .A1(n754), .A2(n755), .Y(n409) );
  NAND2X0_HVT U218 ( .A1(n409), .A2(n411), .Y(n1166) );
  AND2X1_HVT U219 ( .A1(n1116), .A2(n756), .Y(n411) );
  INVX0_HVT U220 ( .A(n777), .Y(n1172) );
  INVX1_HVT U221 ( .A(n1532), .Y(n1456) );
  INVX0_HVT U222 ( .A(n1532), .Y(n562) );
  NAND2X0_HVT U223 ( .A1(n509), .A2(n1261), .Y(n449) );
  NAND2X0_HVT U224 ( .A1(n432), .A2(n434), .Y(n454) );
  NAND2X0_HVT U225 ( .A1(n449), .A2(n454), .Y(out1[124]) );
  INVX0_HVT U226 ( .A(n509), .Y(n432) );
  INVX0_HVT U227 ( .A(n1261), .Y(n434) );
  XOR3X2_HVT U228 ( .A1(n511), .A2(n947), .A3(n512), .Y(n509) );
  XOR3X2_HVT U229 ( .A1(n1078), .A2(n759), .A3(n1079), .Y(n1261) );
  XOR2X2_HVT U230 ( .A1(in[44]), .A2(n1283), .Y(n344) );
  INVX2_HVT U231 ( .A(n1337), .Y(n1283) );
  INVX1_HVT U232 ( .A(n621), .Y(n423) );
  IBUFFX16_HVT U233 ( .A(n586), .Y(n466) );
  XNOR2X2_HVT U234 ( .A1(n9), .A2(n1418), .Y(n926) );
  XOR3X2_HVT U235 ( .A1(n1356), .A2(n242), .A3(n243), .Y(out1[61]) );
  XNOR2X2_HVT U236 ( .A1(n571), .A2(n1285), .Y(n241) );
  XNOR2X1_HVT U237 ( .A1(n12), .A2(n118), .Y(n110) );
  NAND2X0_HVT U238 ( .A1(n131), .A2(n95), .Y(n490) );
  NAND2X0_HVT U239 ( .A1(n480), .A2(n82), .Y(n491) );
  NAND2X0_HVT U240 ( .A1(n490), .A2(n491), .Y(n186) );
  INVX0_HVT U241 ( .A(n131), .Y(n480) );
  XNOR2X2_HVT U242 ( .A1(n825), .A2(n304), .Y(n350) );
  INVX1_HVT U243 ( .A(in[69]), .Y(n1170) );
  AND2X1_HVT U244 ( .A1(n934), .A2(n1146), .Y(n501) );
  INVX0_HVT U245 ( .A(in[85]), .Y(n672) );
  NAND2X0_HVT U246 ( .A1(n313), .A2(n1418), .Y(n517) );
  NAND2X0_HVT U247 ( .A1(n504), .A2(n508), .Y(n522) );
  NAND2X0_HVT U248 ( .A1(n517), .A2(n522), .Y(n303) );
  INVX1_HVT U249 ( .A(n313), .Y(n504) );
  INVX0_HVT U250 ( .A(n1418), .Y(n508) );
  NBUFFX2_HVT U251 ( .A(n1013), .Y(n1418) );
  XOR3X1_HVT U252 ( .A1(n527), .A2(n441), .A3(n442), .Y(out1[23]) );
  IBUFFX16_HVT U253 ( .A(n440), .Y(n527) );
  NAND2X0_HVT U254 ( .A1(n680), .A2(n681), .Y(n553) );
  XNOR2X2_HVT U255 ( .A1(in[50]), .A2(n1531), .Y(n554) );
  XOR3X2_HVT U256 ( .A1(n290), .A2(n562), .A3(n295), .Y(n381) );
  XNOR2X1_HVT U257 ( .A1(n1173), .A2(n10), .Y(n74) );
  INVX1_HVT U258 ( .A(n1128), .Y(n604) );
  AND2X1_HVT U259 ( .A1(n715), .A2(n716), .Y(n569) );
  XOR2X2_HVT U260 ( .A1(n1321), .A2(n1439), .Y(n483) );
  XNOR2X2_HVT U261 ( .A1(n1124), .A2(n1441), .Y(n582) );
  INVX1_HVT U262 ( .A(n1124), .Y(n1125) );
  NBUFFX2_HVT U263 ( .A(n500), .Y(n570) );
  XNOR2X2_HVT U264 ( .A1(n554), .A2(n1418), .Y(n571) );
  INVX1_HVT U265 ( .A(n1544), .Y(n885) );
  IBUFFX2_HVT U266 ( .A(in[88]), .Y(n594) );
  INVX1_HVT U267 ( .A(n594), .Y(n595) );
  AND2X1_HVT U268 ( .A1(n1242), .A2(in[120]), .Y(n598) );
  XOR3X2_HVT U269 ( .A1(n588), .A2(n599), .A3(n590), .Y(out1[111]) );
  IBUFFX16_HVT U270 ( .A(n589), .Y(n599) );
  XNOR2X1_HVT U271 ( .A1(n48), .A2(n1510), .Y(n97) );
  INVX1_HVT U272 ( .A(n854), .Y(n1176) );
  XOR3X2_HVT U273 ( .A1(n604), .A2(n611), .A3(n69), .Y(n608) );
  IBUFFX16_HVT U274 ( .A(n1129), .Y(n611) );
  NAND2X0_HVT U275 ( .A1(n1354), .A2(n1410), .Y(n612) );
  NAND2X0_HVT U276 ( .A1(n1377), .A2(n1495), .Y(n616) );
  INVX2_HVT U277 ( .A(n1428), .Y(n1200) );
  INVX1_HVT U278 ( .A(n929), .Y(n618) );
  XNOR2X1_HVT U279 ( .A1(n99), .A2(n1291), .Y(n131) );
  INVX0_HVT U280 ( .A(n247), .Y(n938) );
  INVX1_HVT U281 ( .A(n25), .Y(n671) );
  INVX0_HVT U282 ( .A(in[97]), .Y(n1225) );
  INVX0_HVT U283 ( .A(n118), .Y(n874) );
  IBUFFX2_HVT U284 ( .A(n571), .Y(n619) );
  INVX1_HVT U285 ( .A(n619), .Y(n620) );
  INVX1_HVT U286 ( .A(n1546), .Y(n771) );
  XOR3X2_HVT U287 ( .A1(n209), .A2(n1392), .A3(n170), .Y(n230) );
  XNOR2X2_HVT U288 ( .A1(n430), .A2(n1439), .Y(n621) );
  XOR3X2_HVT U289 ( .A1(n278), .A2(n622), .A3(n339), .Y(n372) );
  IBUFFX16_HVT U290 ( .A(n949), .Y(n622) );
  INVX0_HVT U291 ( .A(n583), .Y(n1306) );
  XOR2X2_HVT U292 ( .A1(n435), .A2(in[10]), .Y(n405) );
  IBUFFX2_HVT U293 ( .A(in[70]), .Y(n1390) );
  AND2X1_HVT U294 ( .A1(n835), .A2(n834), .Y(n623) );
  XNOR2X2_HVT U295 ( .A1(n1494), .A2(n1290), .Y(n80) );
  NAND2X0_HVT U296 ( .A1(n309), .A2(n625), .Y(n626) );
  NAND2X0_HVT U297 ( .A1(n624), .A2(n920), .Y(n627) );
  NAND2X0_HVT U298 ( .A1(n626), .A2(n627), .Y(out1[51]) );
  INVX0_HVT U299 ( .A(n309), .Y(n624) );
  INVX0_HVT U300 ( .A(n920), .Y(n625) );
  NBUFFX2_HVT U301 ( .A(in[40]), .Y(n628) );
  XNOR2X1_HVT U302 ( .A1(n308), .A2(n307), .Y(n920) );
  XNOR2X2_HVT U303 ( .A1(n629), .A2(n1431), .Y(n602) );
  NAND2X0_HVT U304 ( .A1(n1083), .A2(n1082), .Y(n629) );
  INVX0_HVT U305 ( .A(n1431), .Y(n820) );
  NAND2X0_HVT U306 ( .A1(n1107), .A2(n1108), .Y(n630) );
  NBUFFX2_HVT U307 ( .A(n191), .Y(n631) );
  INVX0_HVT U308 ( .A(in[102]), .Y(n1543) );
  XNOR2X2_HVT U309 ( .A1(n515), .A2(n867), .Y(n547) );
  XNOR2X1_HVT U310 ( .A1(n206), .A2(in[74]), .Y(n163) );
  XOR3X2_HVT U311 ( .A1(n106), .A2(n632), .A3(n108), .Y(out1[90]) );
  IBUFFX16_HVT U312 ( .A(n107), .Y(n632) );
  IBUFFX2_HVT U313 ( .A(n264), .Y(n633) );
  INVX1_HVT U314 ( .A(n633), .Y(n634) );
  INVX1_HVT U315 ( .A(n201), .Y(n854) );
  INVX2_HVT U316 ( .A(in[12]), .Y(n1519) );
  IBUFFX2_HVT U317 ( .A(in[91]), .Y(n635) );
  INVX1_HVT U318 ( .A(n635), .Y(n636) );
  NAND2X0_HVT U319 ( .A1(n903), .A2(n904), .Y(n637) );
  XOR3X2_HVT U320 ( .A1(n638), .A2(n1282), .A3(n156), .Y(n102) );
  AND2X1_HVT U321 ( .A1(n1190), .A2(n1191), .Y(n638) );
  XOR3X1_HVT U322 ( .A1(n784), .A2(n109), .A3(n110), .Y(n106) );
  INVX1_HVT U323 ( .A(n639), .Y(n640) );
  INVX0_HVT U324 ( .A(in[15]), .Y(n1521) );
  IBUFFX16_HVT U325 ( .A(n168), .Y(n641) );
  NBUFFX2_HVT U326 ( .A(n142), .Y(n642) );
  INVX0_HVT U327 ( .A(n171), .Y(n643) );
  INVX1_HVT U328 ( .A(n643), .Y(n644) );
  INVX2_HVT U329 ( .A(n1124), .Y(n695) );
  INVX1_HVT U330 ( .A(n435), .Y(n1301) );
  INVX1_HVT U331 ( .A(n1370), .Y(n664) );
  NAND2X0_HVT U332 ( .A1(in[51]), .A2(n646), .Y(n647) );
  NAND2X0_HVT U333 ( .A1(n645), .A2(n1328), .Y(n648) );
  NAND2X0_HVT U334 ( .A1(n647), .A2(n648), .Y(n251) );
  INVX0_HVT U335 ( .A(in[51]), .Y(n645) );
  INVX0_HVT U336 ( .A(n1328), .Y(n646) );
  INVX0_HVT U337 ( .A(n678), .Y(n649) );
  INVX0_HVT U338 ( .A(in[55]), .Y(n678) );
  INVX0_HVT U339 ( .A(n186), .Y(n650) );
  INVX1_HVT U340 ( .A(n650), .Y(n651) );
  IBUFFX2_HVT U341 ( .A(n472), .Y(n1370) );
  INVX0_HVT U342 ( .A(in[70]), .Y(n1534) );
  INVX1_HVT U343 ( .A(n1343), .Y(n1285) );
  IBUFFX2_HVT U344 ( .A(n1359), .Y(n1348) );
  NAND2X0_HVT U345 ( .A1(n1548), .A2(n576), .Y(n654) );
  NAND2X0_HVT U346 ( .A1(n652), .A2(n653), .Y(n655) );
  NAND2X0_HVT U347 ( .A1(n654), .A2(n655), .Y(n567) );
  INVX0_HVT U348 ( .A(n576), .Y(n652) );
  INVX4_HVT U349 ( .A(n1548), .Y(n653) );
  INVX4_HVT U350 ( .A(n695), .Y(n1548) );
  INVX2_HVT U351 ( .A(n729), .Y(n730) );
  NBUFFX2_HVT U352 ( .A(n362), .Y(n656) );
  INVX0_HVT U353 ( .A(n598), .Y(n657) );
  INVX1_HVT U354 ( .A(in[55]), .Y(n1531) );
  XOR3X2_HVT U355 ( .A1(n658), .A2(n659), .A3(n358), .Y(out1[43]) );
  NAND2X0_HVT U356 ( .A1(n1068), .A2(n1067), .Y(n659) );
  XNOR2X2_HVT U357 ( .A1(n205), .A2(n660), .Y(n164) );
  IBUFFX16_HVT U358 ( .A(in[66]), .Y(n660) );
  NBUFFX2_HVT U359 ( .A(n640), .Y(n661) );
  IBUFFX2_HVT U360 ( .A(in[36]), .Y(n1327) );
  INVX1_HVT U361 ( .A(in[59]), .Y(n1351) );
  XNOR3X1_HVT U362 ( .A1(n291), .A2(n1268), .A3(n244), .Y(n347) );
  INVX1_HVT U363 ( .A(n831), .Y(n829) );
  INVX1_HVT U364 ( .A(n610), .Y(n831) );
  AND2X1_HVT U365 ( .A1(n857), .A2(n856), .Y(n662) );
  XOR3X2_HVT U366 ( .A1(n663), .A2(n664), .A3(n375), .Y(n536) );
  IBUFFX16_HVT U367 ( .A(n470), .Y(n663) );
  XNOR2X2_HVT U368 ( .A1(n728), .A2(n1125), .Y(n503) );
  XOR2X1_HVT U369 ( .A1(n1342), .A2(in[38]), .Y(n365) );
  NAND2X0_HVT U370 ( .A1(n864), .A2(n865), .Y(n665) );
  XOR3X2_HVT U371 ( .A1(n1367), .A2(n1366), .A3(n669), .Y(out1[73]) );
  INVX1_HVT U372 ( .A(n669), .Y(n208) );
  NAND2X0_HVT U373 ( .A1(n1225), .A2(n1543), .Y(n666) );
  IBUFFX2_HVT U374 ( .A(n602), .Y(n674) );
  XOR2X2_HVT U375 ( .A1(n68), .A2(n1226), .Y(n580) );
  XNOR2X2_HVT U376 ( .A1(n820), .A2(n1081), .Y(n68) );
  AND2X1_HVT U377 ( .A1(n812), .A2(n668), .Y(n667) );
  NAND2X0_HVT U378 ( .A1(n810), .A2(n811), .Y(n668) );
  XOR3X2_HVT U379 ( .A1(n116), .A2(n670), .A3(n166), .Y(n669) );
  IBUFFX16_HVT U380 ( .A(n1252), .Y(n670) );
  XOR3X2_HVT U381 ( .A1(n1269), .A2(n671), .A3(n262), .Y(n309) );
  INVX0_HVT U382 ( .A(in[64]), .Y(n993) );
  INVX2_HVT U383 ( .A(n1520), .Y(n1402) );
  XNOR2X2_HVT U384 ( .A1(n1547), .A2(n1397), .Y(n494) );
  INVX2_HVT U385 ( .A(in[116]), .Y(n1547) );
  INVX1_HVT U386 ( .A(n552), .Y(n1333) );
  XOR3X1_HVT U387 ( .A1(n376), .A2(n1434), .A3(n378), .Y(n373) );
  XOR3X2_HVT U388 ( .A1(n268), .A2(n1077), .A3(n266), .Y(out1[58]) );
  INVX0_HVT U389 ( .A(n407), .Y(n750) );
  INVX2_HVT U390 ( .A(in[32]), .Y(n1030) );
  INVX1_HVT U391 ( .A(n672), .Y(n673) );
  INVX1_HVT U392 ( .A(n674), .Y(n675) );
  INVX2_HVT U393 ( .A(n1502), .Y(n1503) );
  INVX0_HVT U394 ( .A(n1480), .Y(n1002) );
  INVX0_HVT U395 ( .A(n1370), .Y(n676) );
  NAND2X0_HVT U396 ( .A1(n983), .A2(n984), .Y(n677) );
  NAND2X0_HVT U397 ( .A1(n649), .A2(n679), .Y(n680) );
  NAND2X0_HVT U398 ( .A1(n678), .A2(in[48]), .Y(n681) );
  NAND2X0_HVT U399 ( .A1(n680), .A2(n681), .Y(n336) );
  INVX0_HVT U400 ( .A(in[48]), .Y(n679) );
  INVX0_HVT U401 ( .A(n553), .Y(n989) );
  IBUFFX2_HVT U402 ( .A(n1063), .Y(n682) );
  INVX0_HVT U403 ( .A(n682), .Y(n683) );
  INVX1_HVT U404 ( .A(in[101]), .Y(n1542) );
  XOR3X2_HVT U405 ( .A1(n684), .A2(n97), .A3(n87), .Y(n1364) );
  IBUFFX16_HVT U406 ( .A(n1365), .Y(n684) );
  INVX2_HVT U407 ( .A(in[22]), .Y(n1522) );
  NAND2X0_HVT U408 ( .A1(n958), .A2(n1525), .Y(n685) );
  IBUFFX2_HVT U409 ( .A(n516), .Y(n957) );
  INVX1_HVT U410 ( .A(n478), .Y(n686) );
  INVX1_HVT U411 ( .A(n686), .Y(n687) );
  INVX1_HVT U412 ( .A(in[22]), .Y(n980) );
  INVX0_HVT U413 ( .A(n1317), .Y(n1318) );
  XOR3X1_HVT U414 ( .A1(n1426), .A2(n139), .A3(n90), .Y(n138) );
  XNOR2X1_HVT U415 ( .A1(n103), .A2(n1290), .Y(n779) );
  NAND2X0_HVT U416 ( .A1(n1485), .A2(n321), .Y(n690) );
  NAND2X0_HVT U417 ( .A1(n688), .A2(n689), .Y(n691) );
  NAND2X0_HVT U418 ( .A1(n690), .A2(n691), .Y(out1[4]) );
  INVX0_HVT U419 ( .A(n1485), .Y(n688) );
  INVX0_HVT U420 ( .A(n321), .Y(n689) );
  XOR3X2_HVT U421 ( .A1(n569), .A2(n1120), .A3(n325), .Y(n1485) );
  XOR2X1_HVT U422 ( .A1(n256), .A2(n968), .Y(n321) );
  INVX0_HVT U423 ( .A(n1209), .Y(n1208) );
  INVX2_HVT U424 ( .A(n980), .Y(n981) );
  NAND2X0_HVT U425 ( .A1(n423), .A2(n1371), .Y(n693) );
  NAND2X0_HVT U426 ( .A1(n621), .A2(n692), .Y(n694) );
  NAND2X0_HVT U427 ( .A1(n693), .A2(n694), .Y(n467) );
  INVX0_HVT U428 ( .A(n1371), .Y(n692) );
  IBUFFX2_HVT U429 ( .A(in[27]), .Y(n1371) );
  INVX0_HVT U430 ( .A(n467), .Y(n1317) );
  INVX0_HVT U431 ( .A(n59), .Y(n731) );
  NAND2X0_HVT U432 ( .A1(n492), .A2(n1296), .Y(n698) );
  NAND2X0_HVT U433 ( .A1(n696), .A2(n697), .Y(n699) );
  NAND2X0_HVT U434 ( .A1(n698), .A2(n699), .Y(n457) );
  INVX1_HVT U435 ( .A(n492), .Y(n696) );
  INVX0_HVT U436 ( .A(n1296), .Y(n697) );
  INVX0_HVT U437 ( .A(n457), .Y(n713) );
  NAND2X0_HVT U438 ( .A1(in[123]), .A2(n701), .Y(n702) );
  NAND2X0_HVT U439 ( .A1(n700), .A2(n1280), .Y(n703) );
  NAND2X0_HVT U440 ( .A1(n702), .A2(n703), .Y(n516) );
  INVX0_HVT U441 ( .A(in[123]), .Y(n700) );
  INVX0_HVT U442 ( .A(n1280), .Y(n701) );
  INVX0_HVT U443 ( .A(n1242), .Y(n1280) );
  XOR2X2_HVT U444 ( .A1(n516), .A2(n1090), .Y(n542) );
  INVX0_HVT U445 ( .A(n895), .Y(n704) );
  XNOR2X2_HVT U446 ( .A1(n1329), .A2(n1200), .Y(n705) );
  NAND2X0_HVT U447 ( .A1(n804), .A2(n805), .Y(n706) );
  XNOR2X2_HVT U448 ( .A1(in[91]), .A2(n1196), .Y(n99) );
  IBUFFX2_HVT U449 ( .A(n430), .Y(n1325) );
  XNOR2X1_HVT U450 ( .A1(n1022), .A2(n577), .Y(n66) );
  IBUFFX2_HVT U451 ( .A(in[48]), .Y(n914) );
  INVX2_HVT U452 ( .A(n565), .Y(n1323) );
  INVX0_HVT U453 ( .A(in[23]), .Y(n1221) );
  INVX0_HVT U454 ( .A(in[31]), .Y(n979) );
  INVX1_HVT U455 ( .A(in[1]), .Y(n1404) );
  IBUFFX2_HVT U456 ( .A(in[65]), .Y(n929) );
  NBUFFX2_HVT U457 ( .A(n419), .Y(n707) );
  INVX0_HVT U458 ( .A(in[89]), .Y(n802) );
  XNOR2X2_HVT U459 ( .A1(n710), .A2(n63), .Y(n72) );
  XNOR2X2_HVT U460 ( .A1(in[35]), .A2(n949), .Y(n708) );
  IBUFFX2_HVT U461 ( .A(n388), .Y(n852) );
  INVX0_HVT U462 ( .A(in[14]), .Y(n709) );
  INVX1_HVT U463 ( .A(n763), .Y(n710) );
  INVX1_HVT U464 ( .A(in[110]), .Y(n1546) );
  NAND2X0_HVT U465 ( .A1(n962), .A2(n963), .Y(n711) );
  XOR3X2_HVT U466 ( .A1(n446), .A2(n712), .A3(n258), .Y(n445) );
  IBUFFX16_HVT U467 ( .A(n1297), .Y(n712) );
  NAND2X0_HVT U468 ( .A1(n457), .A2(n1519), .Y(n715) );
  NAND2X0_HVT U469 ( .A1(n713), .A2(n714), .Y(n716) );
  NAND2X0_HVT U470 ( .A1(n715), .A2(n716), .Y(n323) );
  IBUFFX2_HVT U471 ( .A(n1519), .Y(n714) );
  INVX0_HVT U472 ( .A(n323), .Y(n1211) );
  INVX2_HVT U473 ( .A(n1539), .Y(n1284) );
  NBUFFX2_HVT U474 ( .A(n376), .Y(n717) );
  XOR3X2_HVT U475 ( .A1(n312), .A2(n787), .A3(n314), .Y(n262) );
  INVX2_HVT U476 ( .A(n858), .Y(n859) );
  IBUFFX2_HVT U477 ( .A(n708), .Y(n948) );
  XNOR2X1_HVT U478 ( .A1(n1228), .A2(n348), .Y(n383) );
  IBUFFX2_HVT U479 ( .A(n1244), .Y(n1245) );
  IBUFFX2_HVT U480 ( .A(n101), .Y(n884) );
  XOR3X2_HVT U481 ( .A1(n1111), .A2(n1112), .A3(n64), .Y(n607) );
  XNOR2X2_HVT U482 ( .A1(in[100]), .A2(n1507), .Y(n541) );
  XOR2X2_HVT U483 ( .A1(n1056), .A2(n815), .Y(n162) );
  XNOR2X2_HVT U484 ( .A1(in[24]), .A2(n979), .Y(n430) );
  INVX0_HVT U485 ( .A(n377), .Y(n718) );
  INVX1_HVT U486 ( .A(n718), .Y(n719) );
  XOR3X2_HVT U487 ( .A1(n402), .A2(n720), .A3(n404), .Y(out1[2]) );
  IBUFFX16_HVT U488 ( .A(n403), .Y(n720) );
  IBUFFX2_HVT U489 ( .A(n164), .Y(n772) );
  XOR3X2_HVT U490 ( .A1(n1192), .A2(n1168), .A3(n156), .Y(n1471) );
  NAND2X0_HVT U491 ( .A1(n1031), .A2(n1030), .Y(n721) );
  XOR3X2_HVT U492 ( .A1(n1052), .A2(n978), .A3(n250), .Y(n1481) );
  INVX1_HVT U493 ( .A(n1325), .Y(n722) );
  IBUFFX2_HVT U494 ( .A(in[96]), .Y(n723) );
  INVX1_HVT U495 ( .A(n723), .Y(n724) );
  XNOR3X1_HVT U496 ( .A1(n868), .A2(n734), .A3(n196), .Y(n222) );
  IBUFFX2_HVT U497 ( .A(in[14]), .Y(n1520) );
  NBUFFX2_HVT U498 ( .A(n595), .Y(n725) );
  INVX0_HVT U499 ( .A(n307), .Y(n1447) );
  INVX2_HVT U500 ( .A(in[85]), .Y(n1539) );
  XNOR2X2_HVT U501 ( .A1(n525), .A2(n844), .Y(n572) );
  INVX2_HVT U502 ( .A(in[84]), .Y(n1538) );
  INVX1_HVT U503 ( .A(in[18]), .Y(n1329) );
  NBUFFX2_HVT U504 ( .A(n405), .Y(n726) );
  INVX0_HVT U505 ( .A(n513), .Y(n1078) );
  XOR3X2_HVT U507 ( .A1(n346), .A2(n1453), .A3(n381), .Y(out1[38]) );
  XNOR2X2_HVT U508 ( .A1(n564), .A2(n1440), .Y(n728) );
  INVX1_HVT U509 ( .A(in[102]), .Y(n729) );
  INVX1_HVT U510 ( .A(in[112]), .Y(n890) );
  XOR3X2_HVT U511 ( .A1(n731), .A2(n732), .A3(n521), .Y(n1265) );
  AND2X1_HVT U512 ( .A1(n817), .A2(n683), .Y(n732) );
  INVX1_HVT U513 ( .A(in[34]), .Y(n1016) );
  NBUFFX2_HVT U514 ( .A(n144), .Y(n733) );
  XNOR2X2_HVT U515 ( .A1(n304), .A2(n1384), .Y(n290) );
  XNOR2X2_HVT U516 ( .A1(n673), .A2(n815), .Y(n168) );
  XNOR2X2_HVT U517 ( .A1(n157), .A2(n1324), .Y(n734) );
  XNOR2X2_HVT U518 ( .A1(n1196), .A2(n803), .Y(n109) );
  INVX1_HVT U519 ( .A(in[94]), .Y(n803) );
  XOR3X1_HVT U520 ( .A1(n1340), .A2(n538), .A3(n502), .Y(n544) );
  NBUFFX2_HVT U521 ( .A(n1195), .Y(n735) );
  XOR3X2_HVT U522 ( .A1(n736), .A2(n737), .A3(n102), .Y(n153) );
  IBUFFX16_HVT U523 ( .A(n1206), .Y(n736) );
  NAND2X0_HVT U524 ( .A1(n1194), .A2(n387), .Y(n738) );
  XNOR3X1_HVT U525 ( .A1(n418), .A2(n951), .A3(n707), .Y(n412) );
  XNOR2X2_HVT U526 ( .A1(n224), .A2(n673), .Y(n150) );
  XOR3X2_HVT U527 ( .A1(n739), .A2(n235), .A3(n236), .Y(n234) );
  IBUFFX16_HVT U528 ( .A(n1417), .Y(n739) );
  XOR3X2_HVT U529 ( .A1(n662), .A2(n1388), .A3(n1373), .Y(n92) );
  NBUFFX2_HVT U530 ( .A(n356), .Y(n740) );
  NBUFFX2_HVT U531 ( .A(n136), .Y(n741) );
  AND2X1_HVT U532 ( .A1(n905), .A2(n906), .Y(n742) );
  XNOR2X2_HVT U533 ( .A1(n155), .A2(n1510), .Y(n1363) );
  IBUFFX2_HVT U535 ( .A(n1510), .Y(n1511) );
  XNOR2X2_HVT U536 ( .A1(n1384), .A2(n1456), .Y(n280) );
  IBUFFX2_HVT U538 ( .A(n563), .Y(n1313) );
  NAND2X0_HVT U540 ( .A1(n547), .A2(n503), .Y(n745) );
  NAND2X0_HVT U541 ( .A1(n743), .A2(n744), .Y(n746) );
  NAND2X0_HVT U542 ( .A1(n745), .A2(n746), .Y(n597) );
  INVX0_HVT U543 ( .A(n547), .Y(n743) );
  INVX0_HVT U544 ( .A(n503), .Y(n744) );
  IBUFFX2_HVT U545 ( .A(n596), .Y(n1422) );
  IBUFFX2_HVT U546 ( .A(n407), .Y(n767) );
  NAND2X0_HVT U547 ( .A1(n959), .A2(n685), .Y(n747) );
  AND2X1_HVT U548 ( .A1(n721), .A2(n1032), .Y(n748) );
  XNOR2X2_HVT U549 ( .A1(n1287), .A2(n1291), .Y(n119) );
  NBUFFX2_HVT U550 ( .A(n543), .Y(n749) );
  XNOR2X2_HVT U551 ( .A1(n515), .A2(n788), .Y(n1079) );
  XOR3X2_HVT U552 ( .A1(n750), .A2(n751), .A3(n1483), .Y(out1[29]) );
  NAND2X0_HVT U553 ( .A1(n1336), .A2(n824), .Y(n752) );
  IBUFFX2_HVT U555 ( .A(in[121]), .Y(n1089) );
  INVX0_HVT U556 ( .A(in[126]), .Y(n1090) );
  IBUFFX2_HVT U557 ( .A(in[33]), .Y(n916) );
  INVX1_HVT U558 ( .A(in[87]), .Y(n1055) );
  NBUFFX2_HVT U559 ( .A(n302), .Y(n753) );
  INVX1_HVT U560 ( .A(n1247), .Y(n873) );
  NAND2X0_HVT U561 ( .A1(n195), .A2(n221), .Y(n756) );
  NAND2X0_HVT U562 ( .A1(n754), .A2(n755), .Y(n757) );
  NAND2X0_HVT U563 ( .A1(n757), .A2(n756), .Y(n1405) );
  INVX0_HVT U564 ( .A(n195), .Y(n754) );
  IBUFFX2_HVT U565 ( .A(n221), .Y(n755) );
  INVX0_HVT U566 ( .A(n784), .Y(n758) );
  XNOR2X2_HVT U567 ( .A1(n149), .A2(n188), .Y(n221) );
  INVX2_HVT U568 ( .A(n806), .Y(n784) );
  XOR2X2_HVT U570 ( .A1(n361), .A2(n656), .Y(n265) );
  NBUFFX2_HVT U571 ( .A(n514), .Y(n759) );
  IBUFFX2_HVT U573 ( .A(n103), .Y(n1168) );
  INVX0_HVT U574 ( .A(n1306), .Y(n760) );
  XOR2X2_HVT U575 ( .A1(n1328), .A2(n1417), .Y(n318) );
  INVX1_HVT U576 ( .A(n1300), .Y(n780) );
  INVX1_HVT U577 ( .A(n801), .Y(n1300) );
  NBUFFX2_HVT U578 ( .A(n69), .Y(n761) );
  XNOR2X2_HVT U579 ( .A1(n934), .A2(n1429), .Y(n418) );
  INVX2_HVT U580 ( .A(in[19]), .Y(n934) );
  XOR3X2_HVT U581 ( .A1(n1007), .A2(n275), .A3(n276), .Y(n271) );
  NBUFFX2_HVT U582 ( .A(n64), .Y(n762) );
  AND2X1_HVT U583 ( .A1(n1132), .A2(n1133), .Y(n763) );
  NBUFFX2_HVT U584 ( .A(n728), .Y(n764) );
  NBUFFX2_HVT U585 ( .A(n199), .Y(n765) );
  IBUFFX2_HVT U586 ( .A(n993), .Y(n766) );
  XOR3X1_HVT U587 ( .A1(n767), .A2(n484), .A3(n486), .Y(out1[14]) );
  INVX0_HVT U588 ( .A(n605), .Y(n769) );
  INVX0_HVT U589 ( .A(n769), .Y(n770) );
  XOR3X2_HVT U590 ( .A1(n821), .A2(n771), .A3(n75), .Y(n609) );
  XOR3X2_HVT U591 ( .A1(n203), .A2(n772), .A3(n204), .Y(out1[74]) );
  NBUFFX2_HVT U593 ( .A(n644), .Y(n773) );
  NAND2X0_HVT U594 ( .A1(n1015), .A2(n1014), .Y(n774) );
  NAND2X0_HVT U595 ( .A1(n1105), .A2(n1106), .Y(n775) );
  NBUFFX2_HVT U596 ( .A(n86), .Y(n776) );
  INVX0_HVT U597 ( .A(in[87]), .Y(n1540) );
  AND2X1_HVT U598 ( .A1(n1339), .A2(n1338), .Y(n777) );
  INVX0_HVT U599 ( .A(n1401), .Y(n778) );
  XNOR2X2_HVT U600 ( .A1(n1534), .A2(n781), .Y(n205) );
  XOR3X2_HVT U601 ( .A1(n568), .A2(n780), .A3(n521), .Y(n1299) );
  NBUFFX2_HVT U602 ( .A(in[71]), .Y(n781) );
  NAND2X0_HVT U603 ( .A1(n1405), .A2(n145), .Y(n782) );
  NAND2X0_HVT U604 ( .A1(n812), .A2(n813), .Y(n783) );
  XOR3X2_HVT U606 ( .A1(n503), .A2(n1079), .A3(n505), .Y(out1[125]) );
  XNOR2X1_HVT U607 ( .A1(n734), .A2(n96), .Y(n137) );
  XOR3X2_HVT U608 ( .A1(n687), .A2(n1041), .A3(n406), .Y(n475) );
  INVX2_HVT U610 ( .A(n1340), .Y(n1278) );
  NBUFFX2_HVT U611 ( .A(n218), .Y(n785) );
  XNOR2X2_HVT U612 ( .A1(n513), .A2(n786), .Y(n499) );
  XNOR3X2_HVT U613 ( .A1(n269), .A2(in[57]), .A3(n270), .Y(n266) );
  NBUFFX2_HVT U614 ( .A(n554), .Y(n787) );
  INVX0_HVT U615 ( .A(n957), .Y(n788) );
  INVX1_HVT U616 ( .A(n417), .Y(n832) );
  IBUFFX2_HVT U617 ( .A(n677), .Y(n1039) );
  IBUFFX2_HVT U618 ( .A(n51), .Y(n789) );
  INVX1_HVT U619 ( .A(n789), .Y(n790) );
  NAND2X0_HVT U620 ( .A1(n1037), .A2(n1522), .Y(n793) );
  NAND2X0_HVT U622 ( .A1(n791), .A2(n792), .Y(n794) );
  NAND2X0_HVT U623 ( .A1(n793), .A2(n794), .Y(n465) );
  INVX0_HVT U624 ( .A(n1037), .Y(n791) );
  INVX0_HVT U626 ( .A(n1522), .Y(n792) );
  INVX1_HVT U627 ( .A(n1031), .Y(n949) );
  INVX0_HVT U628 ( .A(in[39]), .Y(n1527) );
  NBUFFX2_HVT U629 ( .A(n293), .Y(n795) );
  XNOR2X1_HVT U630 ( .A1(n950), .A2(n56), .Y(n487) );
  INVX1_HVT U631 ( .A(n950), .Y(n951) );
  INVX1_HVT U632 ( .A(n330), .Y(n818) );
  IBUFFX2_HVT U633 ( .A(n705), .Y(n796) );
  INVX1_HVT U634 ( .A(n796), .Y(n797) );
  XOR3X2_HVT U635 ( .A1(n3), .A2(n798), .A3(n704), .Y(n1476) );
  IBUFFX2_HVT U636 ( .A(in[99]), .Y(n799) );
  INVX1_HVT U637 ( .A(n799), .Y(n800) );
  NAND2X0_HVT U638 ( .A1(n1180), .A2(n1181), .Y(n801) );
  XOR3X2_HVT U639 ( .A1(n945), .A2(n45), .A3(n279), .Y(n340) );
  NAND2X0_HVT U640 ( .A1(in[94]), .A2(in[89]), .Y(n804) );
  NAND2X0_HVT U642 ( .A1(n802), .A2(n803), .Y(n805) );
  NAND2X0_HVT U643 ( .A1(n805), .A2(n804), .Y(n201) );
  INVX1_HVT U644 ( .A(n802), .Y(n806) );
  XOR3X2_HVT U645 ( .A1(n545), .A2(n807), .A3(n550), .Y(n830) );
  IBUFFX2_HVT U646 ( .A(n566), .Y(n808) );
  INVX1_HVT U647 ( .A(n808), .Y(n809) );
  NAND2X0_HVT U648 ( .A1(n150), .A2(n1419), .Y(n812) );
  NAND2X0_HVT U649 ( .A1(n810), .A2(n811), .Y(n813) );
  INVX1_HVT U650 ( .A(n150), .Y(n810) );
  IBUFFX2_HVT U651 ( .A(n1419), .Y(n811) );
  IBUFFX2_HVT U652 ( .A(in[86]), .Y(n814) );
  INVX2_HVT U654 ( .A(n814), .Y(n815) );
  INVX0_HVT U655 ( .A(n1538), .Y(n1419) );
  XOR3X2_HVT U656 ( .A1(n763), .A2(n816), .A3(n66), .Y(n1060) );
  IBUFFX16_HVT U658 ( .A(in[105]), .Y(n816) );
  XOR3X2_HVT U659 ( .A1(n292), .A2(n795), .A3(n1395), .Y(out1[53]) );
  INVX0_HVT U660 ( .A(n519), .Y(n822) );
  XOR3X2_HVT U661 ( .A1(n882), .A2(n570), .A3(n1473), .Y(out1[126]) );
  NAND2X0_HVT U662 ( .A1(n867), .A2(n1062), .Y(n817) );
  XOR3X1_HVT U663 ( .A1(n818), .A2(n331), .A3(n332), .Y(out1[49]) );
  XNOR2X2_HVT U664 ( .A1(n577), .A2(n1542), .Y(n57) );
  XOR3X2_HVT U665 ( .A1(n543), .A2(n1199), .A3(n551), .Y(n613) );
  XOR3X2_HVT U666 ( .A1(n927), .A2(n1421), .A3(n1311), .Y(n413) );
  IBUFFX2_HVT U667 ( .A(n354), .Y(n1442) );
  XNOR2X2_HVT U668 ( .A1(n1281), .A2(n859), .Y(n525) );
  IBUFFX2_HVT U669 ( .A(in[109]), .Y(n1545) );
  XOR3X2_HVT U671 ( .A1(n67), .A2(n1020), .A3(n761), .Y(out1[97]) );
  XOR3X2_HVT U672 ( .A1(n190), .A2(n1375), .A3(n1143), .Y(n1488) );
  NAND2X0_HVT U673 ( .A1(n894), .A2(n895), .Y(n819) );
  INVX0_HVT U675 ( .A(in[101]), .Y(n1431) );
  NBUFFX2_HVT U676 ( .A(n1276), .Y(n821) );
  INVX1_HVT U678 ( .A(n822), .Y(n823) );
  XOR3X2_HVT U679 ( .A1(n623), .A2(n256), .A3(n257), .Y(out1[5]) );
  IBUFFX2_HVT U680 ( .A(n57), .Y(n1386) );
  INVX1_HVT U681 ( .A(n878), .Y(n824) );
  XNOR2X1_HVT U682 ( .A1(n560), .A2(n37), .Y(n614) );
  XNOR2X2_HVT U683 ( .A1(n478), .A2(n1202), .Y(n429) );
  NBUFFX2_HVT U684 ( .A(n252), .Y(n825) );
  INVX1_HVT U686 ( .A(n851), .Y(n840) );
  XNOR3X1_HVT U687 ( .A1(n132), .A2(n1234), .A3(n1368), .Y(n851) );
  XNOR2X2_HVT U688 ( .A1(n96), .A2(n1233), .Y(n132) );
  XNOR2X2_HVT U689 ( .A1(n705), .A2(n1506), .Y(n918) );
  INVX1_HVT U690 ( .A(n1528), .Y(n877) );
  XNOR2X2_HVT U691 ( .A1(n1507), .A2(n730), .Y(n63) );
  IBUFFX2_HVT U692 ( .A(in[26]), .Y(n826) );
  INVX1_HVT U693 ( .A(n826), .Y(n827) );
  INVX0_HVT U694 ( .A(in[31]), .Y(n1246) );
  NBUFFX2_HVT U695 ( .A(n1509), .Y(n828) );
  INVX0_HVT U696 ( .A(n471), .Y(n1509) );
  INVX2_HVT U697 ( .A(in[7]), .Y(n1027) );
  IBUFFX2_HVT U699 ( .A(in[6]), .Y(n1518) );
  XNOR2X2_HVT U700 ( .A1(n1523), .A2(n1439), .Y(n395) );
  XOR3X2_HVT U701 ( .A1(n591), .A2(n829), .A3(n830), .Y(out1[102]) );
  XNOR2X1_HVT U703 ( .A1(n492), .A2(n493), .Y(n421) );
  XNOR2X2_HVT U704 ( .A1(n410), .A2(n452), .Y(n259) );
  NAND2X0_HVT U705 ( .A1(n417), .A2(n1297), .Y(n834) );
  NAND2X0_HVT U706 ( .A1(n832), .A2(n833), .Y(n835) );
  NAND2X0_HVT U707 ( .A1(n835), .A2(n834), .Y(n255) );
  IBUFFX2_HVT U708 ( .A(n1297), .Y(n833) );
  INVX1_HVT U709 ( .A(in[23]), .Y(n1428) );
  NAND2X0_HVT U710 ( .A1(n1478), .A2(n615), .Y(n838) );
  NAND2X0_HVT U711 ( .A1(n836), .A2(n837), .Y(n839) );
  NAND2X0_HVT U712 ( .A1(n838), .A2(n839), .Y(out1[100]) );
  INVX0_HVT U713 ( .A(n1478), .Y(n836) );
  INVX0_HVT U714 ( .A(n615), .Y(n837) );
  INVX0_HVT U716 ( .A(in[98]), .Y(n1179) );
  IBUFFX2_HVT U717 ( .A(n1070), .Y(n1071) );
  XOR3X2_HVT U718 ( .A1(n191), .A2(n1267), .A3(n840), .Y(out1[69]) );
  NBUFFX2_HVT U719 ( .A(in[90]), .Y(n841) );
  INVX1_HVT U720 ( .A(n499), .Y(n846) );
  XNOR2X2_HVT U721 ( .A1(n1417), .A2(in[53]), .Y(n333) );
  IBUFFX2_HVT U722 ( .A(n1179), .Y(n842) );
  INVX0_HVT U723 ( .A(n417), .Y(n950) );
  IBUFFX2_HVT U724 ( .A(in[122]), .Y(n843) );
  INVX1_HVT U725 ( .A(n843), .Y(n844) );
  INVX0_HVT U726 ( .A(n547), .Y(n1430) );
  IBUFFX2_HVT U727 ( .A(in[123]), .Y(n1048) );
  NAND2X0_HVT U728 ( .A1(n542), .A2(n846), .Y(n847) );
  NAND2X0_HVT U729 ( .A1(n845), .A2(n499), .Y(n848) );
  NAND2X0_HVT U730 ( .A1(n847), .A2(n848), .Y(n591) );
  INVX0_HVT U731 ( .A(n542), .Y(n845) );
  XOR2X2_HVT U732 ( .A1(n867), .A2(n859), .Y(n530) );
  XOR3X2_HVT U733 ( .A1(n530), .A2(n940), .A3(n1127), .Y(n1175) );
  INVX1_HVT U734 ( .A(n1270), .Y(n1155) );
  INVX0_HVT U735 ( .A(n779), .Y(n849) );
  INVX1_HVT U736 ( .A(n849), .Y(n850) );
  INVX0_HVT U737 ( .A(n852), .Y(n853) );
  XOR2X2_HVT U738 ( .A1(n1499), .A2(n1436), .Y(n181) );
  NAND2X0_HVT U739 ( .A1(n870), .A2(n706), .Y(n856) );
  NAND2X0_HVT U740 ( .A1(n854), .A2(n855), .Y(n857) );
  NAND2X0_HVT U741 ( .A1(n857), .A2(n856), .Y(n93) );
  INVX0_HVT U742 ( .A(n870), .Y(n855) );
  INVX2_HVT U744 ( .A(in[37]), .Y(n1525) );
  XNOR2X2_HVT U745 ( .A1(n600), .A2(n1464), .Y(n860) );
  NAND2X0_HVT U746 ( .A1(n896), .A2(n819), .Y(n861) );
  NAND2X0_HVT U747 ( .A1(n943), .A2(n944), .Y(n862) );
  NAND2X0_HVT U748 ( .A1(n93), .A2(n1186), .Y(n864) );
  NAND2X0_HVT U749 ( .A1(n662), .A2(n863), .Y(n865) );
  NAND2X0_HVT U750 ( .A1(n865), .A2(n864), .Y(n1270) );
  INVX2_HVT U751 ( .A(n1186), .Y(n863) );
  INVX2_HVT U752 ( .A(n1234), .Y(n1186) );
  INVX1_HVT U753 ( .A(in[120]), .Y(n1094) );
  INVX1_HVT U754 ( .A(n334), .Y(n1336) );
  XNOR2X2_HVT U755 ( .A1(in[43]), .A2(n45), .Y(n304) );
  INVX2_HVT U756 ( .A(n555), .Y(n1043) );
  OR2X1_HVT U757 ( .A1(n246), .A2(n1481), .Y(n977) );
  XNOR2X2_HVT U758 ( .A1(n1195), .A2(n463), .Y(n1273) );
  INVX1_HVT U759 ( .A(n556), .Y(n894) );
  IBUFFX2_HVT U760 ( .A(n825), .Y(n1349) );
  XNOR2X2_HVT U761 ( .A1(n206), .A2(n109), .Y(n120) );
  INVX0_HVT U762 ( .A(in[125]), .Y(n866) );
  INVX1_HVT U763 ( .A(n866), .Y(n867) );
  NBUFFX2_HVT U764 ( .A(n99), .Y(n868) );
  XOR3X2_HVT U765 ( .A1(n869), .A2(n122), .A3(n123), .Y(out1[88]) );
  XOR3X2_HVT U766 ( .A1(n1196), .A2(n1291), .A3(n124), .Y(n869) );
  NBUFFX2_HVT U767 ( .A(in[93]), .Y(n870) );
  XOR3X2_HVT U768 ( .A1(n871), .A2(n177), .A3(n212), .Y(out1[72]) );
  XOR3X2_HVT U769 ( .A1(n1503), .A2(n1511), .A3(n80), .Y(n871) );
  XNOR3X1_HVT U770 ( .A1(n322), .A2(n883), .A3(n587), .Y(n584) );
  XNOR2X1_HVT U771 ( .A1(n1268), .A2(n1417), .Y(n284) );
  XNOR3X1_HVT U772 ( .A1(n1522), .A2(n991), .A3(n483), .Y(n481) );
  XNOR3X1_HVT U773 ( .A1(n74), .A2(n1397), .A3(n586), .Y(n534) );
  XOR3X2_HVT U774 ( .A1(n439), .A2(n872), .A3(n483), .Y(n113) );
  IBUFFX16_HVT U775 ( .A(n1224), .Y(n872) );
  INVX0_HVT U776 ( .A(in[107]), .Y(n1163) );
  XOR3X1_HVT U777 ( .A1(n1343), .A2(n233), .A3(n240), .Y(n239) );
  XOR2X2_HVT U778 ( .A1(in[52]), .A2(n1328), .Y(n232) );
  INVX1_HVT U779 ( .A(in[52]), .Y(n1009) );
  XOR3X2_HVT U780 ( .A1(n873), .A2(n1266), .A3(n439), .Y(n436) );
  INVX0_HVT U781 ( .A(n1507), .Y(n1257) );
  XOR3X2_HVT U782 ( .A1(n874), .A2(n119), .A3(n120), .Y(n115) );
  XOR3X2_HVT U783 ( .A1(n651), .A2(n875), .A3(n215), .Y(out1[70]) );
  IBUFFX16_HVT U784 ( .A(n213), .Y(n875) );
  INVX1_HVT U785 ( .A(in[38]), .Y(n1526) );
  INVX0_HVT U786 ( .A(n926), .Y(n237) );
  XNOR3X1_HVT U787 ( .A1(n343), .A2(n344), .A3(n345), .Y(out1[47]) );
  XOR3X2_HVT U788 ( .A1(n394), .A2(n395), .A3(n876), .Y(out1[31]) );
  XOR3X2_HVT U789 ( .A1(n114), .A2(n1506), .A3(n397), .Y(n876) );
  XNOR2X2_HVT U790 ( .A1(in[25]), .A2(n922), .Y(n493) );
  NAND2X0_HVT U791 ( .A1(n1132), .A2(n1133), .Y(n575) );
  INVX1_HVT U792 ( .A(n426), .Y(n1414) );
  XOR3X2_HVT U793 ( .A1(n877), .A2(n284), .A3(n236), .Y(n283) );
  XNOR2X2_HVT U794 ( .A1(n362), .A2(n878), .Y(n354) );
  INVX0_HVT U795 ( .A(n462), .Y(n1159) );
  INVX0_HVT U796 ( .A(n1532), .Y(n879) );
  XNOR2X2_HVT U797 ( .A1(n269), .A2(n880), .Y(n316) );
  IBUFFX16_HVT U798 ( .A(in[58]), .Y(n880) );
  XOR3X2_HVT U799 ( .A1(n316), .A2(n916), .A3(n267), .Y(n364) );
  INVX1_HVT U800 ( .A(n267), .Y(n1077) );
  INVX1_HVT U801 ( .A(n542), .Y(n921) );
  INVX0_HVT U802 ( .A(n118), .Y(n1392) );
  NAND2X0_HVT U803 ( .A1(n890), .A2(n891), .Y(n881) );
  INVX1_HVT U804 ( .A(n1549), .Y(n891) );
  NBUFFX2_HVT U805 ( .A(n499), .Y(n882) );
  XNOR3X1_HVT U806 ( .A1(n541), .A2(n1293), .A3(n533), .Y(n590) );
  NBUFFX2_HVT U807 ( .A(in[111]), .Y(n883) );
  XOR3X2_HVT U808 ( .A1(n1474), .A2(n884), .A3(n1504), .Y(out1[91]) );
  XNOR2X2_HVT U809 ( .A1(in[74]), .A2(n898), .Y(n155) );
  INVX0_HVT U810 ( .A(in[79]), .Y(n898) );
  INVX0_HVT U811 ( .A(in[72]), .Y(n886) );
  INVX1_HVT U812 ( .A(n886), .Y(n887) );
  XNOR3X1_HVT U813 ( .A1(n232), .A2(n233), .A3(n234), .Y(out1[63]) );
  NAND2X0_HVT U814 ( .A1(n892), .A2(n881), .Y(n888) );
  NAND2X0_HVT U815 ( .A1(n1082), .A2(n666), .Y(n889) );
  NAND2X0_HVT U816 ( .A1(n1034), .A2(in[112]), .Y(n892) );
  NAND2X0_HVT U817 ( .A1(n890), .A2(n891), .Y(n893) );
  NAND2X0_HVT U818 ( .A1(n892), .A2(n893), .Y(n576) );
  NAND2X0_HVT U819 ( .A1(n556), .A2(n557), .Y(n896) );
  NAND2X0_HVT U820 ( .A1(n894), .A2(n895), .Y(n897) );
  NAND2X0_HVT U821 ( .A1(n896), .A2(n897), .Y(n512) );
  INVX1_HVT U822 ( .A(n557), .Y(n895) );
  XNOR2X2_HVT U823 ( .A1(in[90]), .A2(n1541), .Y(n103) );
  INVX1_HVT U824 ( .A(n614), .Y(n1466) );
  XOR2X2_HVT U825 ( .A1(n365), .A2(n318), .Y(n330) );
  NAND2X0_HVT U826 ( .A1(n1448), .A2(n1449), .Y(n901) );
  NAND2X0_HVT U827 ( .A1(n899), .A2(n900), .Y(n902) );
  NAND2X0_HVT U828 ( .A1(n901), .A2(n902), .Y(out1[44]) );
  INVX0_HVT U829 ( .A(n1448), .Y(n899) );
  INVX0_HVT U830 ( .A(n1449), .Y(n900) );
  NAND2X0_HVT U831 ( .A1(n386), .A2(n1285), .Y(n905) );
  NAND2X0_HVT U832 ( .A1(n903), .A2(n904), .Y(n906) );
  NAND2X0_HVT U833 ( .A1(n905), .A2(n637), .Y(n306) );
  INVX0_HVT U834 ( .A(n386), .Y(n903) );
  INVX2_HVT U835 ( .A(n1285), .Y(n904) );
  XOR3X2_HVT U836 ( .A1(n1442), .A2(n1443), .A3(n355), .Y(n1448) );
  XOR3X2_HVT U837 ( .A1(n582), .A2(n1306), .A3(n72), .Y(n578) );
  XOR2X2_HVT U838 ( .A1(n296), .A2(n297), .Y(n245) );
  XOR2X1_HVT U839 ( .A1(n209), .A2(n618), .Y(n172) );
  XOR2X2_HVT U840 ( .A1(n129), .A2(n130), .Y(n81) );
  INVX0_HVT U841 ( .A(in[30]), .Y(n922) );
  XOR3X2_HVT U842 ( .A1(n1469), .A2(n1197), .A3(n1198), .Y(out1[115]) );
  NAND2X0_HVT U843 ( .A1(n1010), .A2(n1011), .Y(n907) );
  XOR3X2_HVT U844 ( .A1(n423), .A2(n1434), .A3(n1154), .Y(n420) );
  XNOR2X2_HVT U845 ( .A1(n1432), .A2(n908), .Y(n60) );
  AND2X1_HVT U846 ( .A1(n1109), .A2(n630), .Y(n908) );
  XNOR2X2_HVT U847 ( .A1(n883), .A2(n1546), .Y(n574) );
  NAND2X0_HVT U848 ( .A1(n1450), .A2(n1347), .Y(n911) );
  NAND2X0_HVT U849 ( .A1(n909), .A2(n910), .Y(n912) );
  NAND2X0_HVT U850 ( .A1(n911), .A2(n912), .Y(out1[36]) );
  INVX0_HVT U851 ( .A(n1450), .Y(n909) );
  INVX0_HVT U852 ( .A(n1347), .Y(n910) );
  XNOR3X1_HVT U853 ( .A1(n1358), .A2(n1526), .A3(n341), .Y(n393) );
  XNOR2X2_HVT U854 ( .A1(n915), .A2(n1530), .Y(n278) );
  INVX0_HVT U855 ( .A(n888), .Y(n1021) );
  INVX1_HVT U856 ( .A(n1274), .Y(n913) );
  IBUFFX2_HVT U857 ( .A(n614), .Y(n1051) );
  INVX1_HVT U858 ( .A(n914), .Y(n915) );
  XNOR2X2_HVT U859 ( .A1(n369), .A2(n916), .Y(n337) );
  XOR3X2_HVT U860 ( .A1(n1424), .A2(n1422), .A3(n1423), .Y(out1[109]) );
  XNOR2X2_HVT U861 ( .A1(in[35]), .A2(n949), .Y(n348) );
  XOR3X1_HVT U862 ( .A1(n1337), .A2(n282), .A3(n240), .Y(n289) );
  INVX1_HVT U863 ( .A(n249), .Y(n1052) );
  NAND2X0_HVT U864 ( .A1(n1211), .A2(n94), .Y(n917) );
  NBUFFX2_HVT U865 ( .A(n676), .Y(n919) );
  XOR3X2_HVT U866 ( .A1(n258), .A2(in[28]), .A3(n259), .Y(n257) );
  XOR2X2_HVT U867 ( .A1(n57), .A2(n800), .Y(n565) );
  XOR2X2_HVT U868 ( .A1(n444), .A2(n178), .Y(n394) );
  IBUFFX2_HVT U869 ( .A(n1394), .Y(n1324) );
  INVX2_HVT U870 ( .A(in[86]), .Y(n1394) );
  XOR3X1_HVT U871 ( .A1(n921), .A2(n749), .A3(n544), .Y(out1[118]) );
  XOR3X2_HVT U872 ( .A1(n469), .A2(n1435), .A3(n536), .Y(out1[11]) );
  INVX2_HVT U873 ( .A(n1428), .Y(n1429) );
  INVX1_HVT U874 ( .A(in[79]), .Y(n1537) );
  INVX1_HVT U875 ( .A(n989), .Y(n990) );
  INVX0_HVT U876 ( .A(n1280), .Y(n1281) );
  INVX1_HVT U877 ( .A(n1289), .Y(n1111) );
  INVX0_HVT U878 ( .A(n941), .Y(n1112) );
  INVX0_HVT U879 ( .A(n1182), .Y(n1161) );
  INVX1_HVT U880 ( .A(n151), .Y(n988) );
  XNOR2X1_HVT U881 ( .A1(n1251), .A2(in[20]), .Y(n219) );
  INVX0_HVT U882 ( .A(n1306), .Y(n1129) );
  INVX0_HVT U883 ( .A(n68), .Y(n1020) );
  INVX0_HVT U884 ( .A(n1165), .Y(n1252) );
  INVX1_HVT U885 ( .A(n1357), .Y(n1080) );
  INVX1_HVT U886 ( .A(n573), .Y(n1008) );
  INVX0_HVT U887 ( .A(in[11]), .Y(n1047) );
  INVX1_HVT U888 ( .A(n1313), .Y(n1023) );
  INVX1_HVT U889 ( .A(n165), .Y(n1102) );
  INVX0_HVT U890 ( .A(in[44]), .Y(n1126) );
  INVX1_HVT U891 ( .A(n408), .Y(n1421) );
  INVX1_HVT U892 ( .A(n1277), .Y(n1266) );
  INVX1_HVT U893 ( .A(n518), .Y(n1264) );
  INVX0_HVT U894 ( .A(n1313), .Y(n1197) );
  INVX0_HVT U895 ( .A(n589), .Y(n1065) );
  INVX1_HVT U896 ( .A(n528), .Y(n1158) );
  XOR3X1_HVT U897 ( .A1(n125), .A2(n126), .A3(n1271), .Y(out1[87]) );
  INVX0_HVT U898 ( .A(n131), .Y(n1098) );
  INVX0_HVT U899 ( .A(n154), .Y(n1206) );
  INVX0_HVT U900 ( .A(n184), .Y(n1238) );
  INVX0_HVT U901 ( .A(n758), .Y(n1035) );
  XOR3X1_HVT U902 ( .A1(n925), .A2(n316), .A3(n317), .Y(out1[50]) );
  INVX0_HVT U903 ( .A(n1418), .Y(n945) );
  INVX0_HVT U904 ( .A(n1420), .Y(n956) );
  INVX1_HVT U905 ( .A(n1320), .Y(n1259) );
  INVX0_HVT U906 ( .A(n441), .Y(n1113) );
  INVX1_HVT U907 ( .A(n1188), .Y(n1192) );
  INVX0_HVT U908 ( .A(n424), .Y(n1153) );
  INVX0_HVT U909 ( .A(n1400), .Y(n1140) );
  INVX1_HVT U910 ( .A(n140), .Y(n1103) );
  AND2X1_HVT U911 ( .A1(n1018), .A2(n985), .Y(n923) );
  INVX0_HVT U912 ( .A(n1479), .Y(n1303) );
  NAND2X0_HVT U913 ( .A1(n1169), .A2(n1190), .Y(n924) );
  XNOR2X2_HVT U914 ( .A1(n990), .A2(n1069), .Y(n925) );
  INVX1_HVT U915 ( .A(n1495), .Y(n1378) );
  INVX1_HVT U916 ( .A(in[105]), .Y(n941) );
  INVX0_HVT U917 ( .A(in[68]), .Y(n1233) );
  INVX1_HVT U918 ( .A(n1413), .Y(n1093) );
  INVX0_HVT U919 ( .A(n1131), .Y(n1224) );
  INVX0_HVT U920 ( .A(n1193), .Y(n1194) );
  INVX1_HVT U921 ( .A(n350), .Y(n1443) );
  INVX1_HVT U922 ( .A(n938), .Y(n939) );
  INVX1_HVT U923 ( .A(in[124]), .Y(n1199) );
  INVX0_HVT U924 ( .A(in[92]), .Y(n1234) );
  INVX1_HVT U925 ( .A(n1287), .Y(n1362) );
  INVX1_HVT U926 ( .A(n146), .Y(n1115) );
  INVX1_HVT U927 ( .A(in[28]), .Y(n1523) );
  INVX1_HVT U928 ( .A(n1325), .Y(n1160) );
  INVX0_HVT U929 ( .A(n1459), .Y(n1214) );
  INVX1_HVT U930 ( .A(n450), .Y(n1406) );
  XNOR2X1_HVT U931 ( .A1(n770), .A2(n862), .Y(n518) );
  INVX0_HVT U932 ( .A(n55), .Y(n1001) );
  INVX1_HVT U933 ( .A(n519), .Y(n1198) );
  NAND2X0_HVT U934 ( .A1(n1514), .A2(n1515), .Y(n928) );
  XOR3X2_HVT U935 ( .A1(n420), .A2(n1435), .A3(n422), .Y(out1[27]) );
  IBUFFX2_HVT U936 ( .A(n190), .Y(n1174) );
  XOR3X2_HVT U937 ( .A1(n107), .A2(n929), .A3(n160), .Y(n204) );
  XNOR2X2_HVT U938 ( .A1(n1516), .A2(in[5]), .Y(n179) );
  NBUFFX2_HVT U939 ( .A(n991), .Y(n930) );
  IBUFFX2_HVT U940 ( .A(in[106]), .Y(n931) );
  INVX1_HVT U941 ( .A(n931), .Y(n932) );
  INVX0_HVT U942 ( .A(in[37]), .Y(n1268) );
  XNOR2X2_HVT U943 ( .A1(n302), .A2(n301), .Y(n250) );
  XOR3X2_HVT U944 ( .A1(n933), .A2(n159), .A3(n204), .Y(out1[66]) );
  NAND2X0_HVT U945 ( .A1(n471), .A2(in[19]), .Y(n935) );
  NAND2X0_HVT U946 ( .A1(n501), .A2(n1147), .Y(n936) );
  NAND2X0_HVT U947 ( .A1(n935), .A2(n936), .Y(n424) );
  XNOR2X2_HVT U948 ( .A1(in[67]), .A2(n1535), .Y(n188) );
  XOR2X2_HVT U949 ( .A1(n53), .A2(n1088), .Y(n937) );
  XOR2X2_HVT U950 ( .A1(n459), .A2(n937), .Y(n431) );
  IBUFFX2_HVT U951 ( .A(n1262), .Y(n1088) );
  XOR3X1_HVT U952 ( .A1(n1272), .A2(n460), .A3(n431), .Y(out1[17]) );
  XNOR2X1_HVT U953 ( .A1(n1296), .A2(n1520), .Y(n54) );
  INVX1_HVT U954 ( .A(in[109]), .Y(n1340) );
  IBUFFX2_HVT U955 ( .A(in[3]), .Y(n1054) );
  NAND2X0_HVT U956 ( .A1(n642), .A2(n657), .Y(n940) );
  NAND2X0_HVT U957 ( .A1(in[105]), .A2(n1171), .Y(n943) );
  NAND2X0_HVT U958 ( .A1(n941), .A2(n942), .Y(n944) );
  NAND2X0_HVT U959 ( .A1(n943), .A2(n944), .Y(n606) );
  XNOR2X2_HVT U960 ( .A1(n311), .A2(n877), .Y(n252) );
  INVX1_HVT U961 ( .A(in[67]), .Y(n1232) );
  NAND2X0_HVT U962 ( .A1(n1045), .A2(n1044), .Y(n946) );
  AND2X1_HVT U963 ( .A1(n1074), .A2(n1075), .Y(n947) );
  XOR3X2_HVT U964 ( .A1(n1057), .A2(n948), .A3(n753), .Y(n1449) );
  XOR2X2_HVT U965 ( .A1(in[68]), .A2(n781), .Y(n130) );
  XOR3X1_HVT U966 ( .A1(n206), .A2(n1093), .A3(n110), .Y(n203) );
  XNOR2X2_HVT U967 ( .A1(in[11]), .A2(n992), .Y(n448) );
  INVX1_HVT U968 ( .A(n217), .Y(n967) );
  INVX1_HVT U969 ( .A(n1241), .Y(n1242) );
  INVX1_HVT U970 ( .A(in[5]), .Y(n1517) );
  INVX1_HVT U971 ( .A(n1425), .Y(n952) );
  XNOR2X2_HVT U972 ( .A1(n252), .A2(n953), .Y(n296) );
  XNOR2X2_HVT U973 ( .A1(n99), .A2(in[76]), .Y(n83) );
  IBUFFX2_HVT U974 ( .A(n564), .Y(n954) );
  INVX1_HVT U975 ( .A(n954), .Y(n955) );
  XNOR2X1_HVT U976 ( .A1(n328), .A2(n1251), .Y(n256) );
  INVX0_HVT U977 ( .A(n121), .Y(n1171) );
  XOR3X2_HVT U978 ( .A1(n956), .A2(n1005), .A3(n964), .Y(n1483) );
  XOR3X2_HVT U979 ( .A1(n675), .A2(n957), .A3(n764), .Y(n615) );
  NAND2X0_HVT U980 ( .A1(n1038), .A2(n390), .Y(n959) );
  NAND2X0_HVT U981 ( .A1(n958), .A2(n1525), .Y(n960) );
  NAND2X0_HVT U982 ( .A1(n960), .A2(n959), .Y(n1059) );
  INVX0_HVT U983 ( .A(n390), .Y(n958) );
  INVX0_HVT U984 ( .A(n1059), .Y(n359) );
  INVX1_HVT U985 ( .A(n241), .Y(n1356) );
  NAND2X0_HVT U986 ( .A1(n447), .A2(n967), .Y(n962) );
  NAND2X0_HVT U987 ( .A1(n961), .A2(n217), .Y(n963) );
  NAND2X0_HVT U988 ( .A1(n962), .A2(n963), .Y(n400) );
  INVX0_HVT U989 ( .A(n447), .Y(n961) );
  XOR3X1_HVT U990 ( .A1(n1548), .A2(n999), .A3(n502), .Y(n1473) );
  INVX0_HVT U991 ( .A(n495), .Y(n999) );
  XNOR2X1_HVT U992 ( .A1(n418), .A2(n1516), .Y(n258) );
  XNOR2X1_HVT U993 ( .A1(in[56]), .A2(in[61]), .Y(n339) );
  NAND2X0_HVT U994 ( .A1(n983), .A2(n984), .Y(n964) );
  INVX0_HVT U995 ( .A(n969), .Y(n965) );
  NBUFFX2_HVT U996 ( .A(n359), .Y(n966) );
  XOR3X2_HVT U997 ( .A1(n216), .A2(n967), .A3(n785), .Y(out1[6]) );
  XNOR2X2_HVT U998 ( .A1(in[0]), .A2(n1517), .Y(n112) );
  XOR3X2_HVT U999 ( .A1(n850), .A2(n188), .A3(n1115), .Y(n1487) );
  INVX0_HVT U1000 ( .A(n1385), .Y(n1041) );
  XNOR2X1_HVT U1001 ( .A1(n326), .A2(n918), .Y(n968) );
  AND2X1_HVT U1002 ( .A1(n1028), .A2(n1029), .Y(n969) );
  XNOR2X2_HVT U1003 ( .A1(n1251), .A2(n1518), .Y(n447) );
  XOR2X1_HVT U1004 ( .A1(n275), .A2(in[57]), .Y(n331) );
  NAND2X0_HVT U1005 ( .A1(n1334), .A2(n1335), .Y(n970) );
  XNOR3X1_HVT U1006 ( .A1(n112), .A2(n1429), .A3(n482), .Y(n438) );
  NAND2X0_HVT U1007 ( .A1(n923), .A2(n1193), .Y(n971) );
  NAND2X0_HVT U1008 ( .A1(n1016), .A2(n1017), .Y(n972) );
  NAND2X0_HVT U1009 ( .A1(n972), .A2(n973), .Y(n987) );
  AND2X1_HVT U1010 ( .A1(n1018), .A2(n1193), .Y(n973) );
  INVX1_HVT U1011 ( .A(n54), .Y(n1000) );
  NAND2X0_HVT U1012 ( .A1(n971), .A2(n738), .Y(n974) );
  IBUFFX2_HVT U1013 ( .A(n982), .Y(n975) );
  INVX1_HVT U1014 ( .A(n451), .Y(n982) );
  NAND2X0_HVT U1015 ( .A1(n246), .A2(n1481), .Y(n976) );
  NAND2X0_HVT U1016 ( .A1(n976), .A2(n977), .Y(out1[60]) );
  XOR3X2_HVT U1017 ( .A1(n1348), .A2(n1349), .A3(n242), .Y(n246) );
  AND2X1_HVT U1018 ( .A1(n1412), .A2(n1457), .Y(n978) );
  NAND2X0_HVT U1019 ( .A1(n451), .A2(n255), .Y(n983) );
  NAND2X0_HVT U1020 ( .A1(n982), .A2(n623), .Y(n984) );
  NAND2X0_HVT U1021 ( .A1(n1016), .A2(n1017), .Y(n985) );
  NAND2X0_HVT U1022 ( .A1(n387), .A2(n1194), .Y(n986) );
  NAND2X0_HVT U1023 ( .A1(n986), .A2(n987), .Y(n305) );
  XOR3X2_HVT U1024 ( .A1(n776), .A2(n1344), .A3(n88), .Y(out1[93]) );
  XOR3X1_HVT U1025 ( .A1(n988), .A2(n152), .A3(n153), .Y(out1[83]) );
  INVX0_HVT U1026 ( .A(in[16]), .Y(n1070) );
  XNOR2X2_HVT U1027 ( .A1(in[60]), .A2(n1358), .Y(n281) );
  INVX1_HVT U1028 ( .A(n1221), .Y(n998) );
  NAND2X0_HVT U1029 ( .A1(in[64]), .A2(n1535), .Y(n995) );
  NAND2X0_HVT U1030 ( .A1(n993), .A2(n994), .Y(n996) );
  NAND2X0_HVT U1031 ( .A1(n995), .A2(n996), .Y(n228) );
  NBUFFX2_HVT U1032 ( .A(n263), .Y(n997) );
  XOR3X2_HVT U1033 ( .A1(n53), .A2(n1000), .A3(n1001), .Y(n1472) );
  NAND2X0_HVT U1034 ( .A1(n1303), .A2(n1480), .Y(n1003) );
  NAND2X0_HVT U1035 ( .A1(n1002), .A2(n1479), .Y(n1004) );
  NAND2X0_HVT U1036 ( .A1(n1003), .A2(n1004), .Y(out1[52]) );
  XNOR2X2_HVT U1037 ( .A1(in[26]), .A2(n1246), .Y(n377) );
  INVX0_HVT U1038 ( .A(n974), .Y(n1227) );
  XNOR2X2_HVT U1039 ( .A1(n98), .A2(n1362), .Y(n136) );
  AND2X1_HVT U1040 ( .A1(n642), .A2(n657), .Y(n1006) );
  INVX1_HVT U1041 ( .A(n1142), .Y(n1108) );
  INVX1_HVT U1042 ( .A(in[61]), .Y(n1532) );
  XOR3X1_HVT U1043 ( .A1(n523), .A2(n1008), .A3(n607), .Y(out1[106]) );
  NAND2X0_HVT U1044 ( .A1(n1070), .A2(n998), .Y(n1223) );
  NAND2X0_HVT U1045 ( .A1(n1403), .A2(n306), .Y(n1010) );
  NAND2X0_HVT U1046 ( .A1(n742), .A2(n1009), .Y(n1011) );
  NAND2X0_HVT U1047 ( .A1(n1011), .A2(n1010), .Y(n249) );
  NAND2X0_HVT U1048 ( .A1(in[49]), .A2(n1314), .Y(n1014) );
  NAND2X0_HVT U1049 ( .A1(n1012), .A2(n1013), .Y(n1015) );
  NAND2X0_HVT U1050 ( .A1(n1015), .A2(n1014), .Y(n386) );
  INVX1_HVT U1051 ( .A(n1314), .Y(n1013) );
  XNOR2X2_HVT U1052 ( .A1(n365), .A2(n1016), .Y(n320) );
  NAND2X0_HVT U1053 ( .A1(in[34]), .A2(n1527), .Y(n1018) );
  NAND2X0_HVT U1054 ( .A1(n1016), .A2(n1017), .Y(n1019) );
  NAND2X0_HVT U1055 ( .A1(n1019), .A2(n1018), .Y(n387) );
  INVX0_HVT U1056 ( .A(n1341), .Y(n1017) );
  XOR3X2_HVT U1057 ( .A1(n373), .A2(n1058), .A3(n1148), .Y(out1[3]) );
  INVX1_HVT U1058 ( .A(n1021), .Y(n1022) );
  XOR3X2_HVT U1059 ( .A1(n809), .A2(n1023), .A3(n1299), .Y(n603) );
  XNOR2X2_HVT U1060 ( .A1(n1038), .A2(n1526), .Y(n369) );
  NAND2X0_HVT U1061 ( .A1(n1117), .A2(n1118), .Y(n1024) );
  INVX0_HVT U1062 ( .A(n1227), .Y(n1025) );
  INVX1_HVT U1063 ( .A(n1227), .Y(n1228) );
  NAND2X0_HVT U1064 ( .A1(in[2]), .A2(n1027), .Y(n1028) );
  NAND2X0_HVT U1065 ( .A1(n1026), .A2(in[7]), .Y(n1029) );
  NAND2X0_HVT U1066 ( .A1(n1028), .A2(n1029), .Y(n489) );
  NAND2X0_HVT U1067 ( .A1(in[32]), .A2(n1341), .Y(n1032) );
  NAND2X0_HVT U1068 ( .A1(n1031), .A2(n1030), .Y(n1033) );
  NAND2X0_HVT U1069 ( .A1(n1033), .A2(n1032), .Y(n390) );
  INVX1_HVT U1070 ( .A(n1341), .Y(n1031) );
  INVX0_HVT U1071 ( .A(in[119]), .Y(n1034) );
  XNOR2X2_HVT U1072 ( .A1(n1283), .A2(n1496), .Y(n235) );
  XNOR2X2_HVT U1073 ( .A1(in[14]), .A2(in[9]), .Y(n492) );
  INVX1_HVT U1074 ( .A(n923), .Y(n1073) );
  INVX0_HVT U1075 ( .A(in[21]), .Y(n1036) );
  INVX1_HVT U1076 ( .A(n1036), .Y(n1037) );
  XNOR3X1_HVT U1077 ( .A1(n304), .A2(n1025), .A3(n1307), .Y(n1479) );
  INVX1_HVT U1078 ( .A(n1525), .Y(n1038) );
  INVX0_HVT U1079 ( .A(n1039), .Y(n1040) );
  INVX0_HVT U1080 ( .A(in[7]), .Y(n1130) );
  NAND2X0_HVT U1081 ( .A1(n1043), .A2(n511), .Y(n1044) );
  NAND2X0_HVT U1082 ( .A1(n1042), .A2(n555), .Y(n1045) );
  NAND2X0_HVT U1083 ( .A1(n1045), .A2(n1044), .Y(n601) );
  NAND2X0_HVT U1084 ( .A1(n1109), .A2(n1110), .Y(n1046) );
  XNOR2X2_HVT U1085 ( .A1(n470), .A2(n1047), .Y(n378) );
  XNOR3X1_HVT U1086 ( .A1(n287), .A2(n288), .A3(n289), .Y(out1[54]) );
  XNOR2X2_HVT U1087 ( .A1(n1319), .A2(n1525), .Y(n342) );
  XOR3X2_HVT U1088 ( .A1(n1213), .A2(n179), .A3(n219), .Y(n216) );
  INVX0_HVT U1089 ( .A(n1438), .Y(n1213) );
  XNOR2X2_HVT U1090 ( .A1(n520), .A2(n1048), .Y(n568) );
  NBUFFX2_HVT U1091 ( .A(n1022), .Y(n1049) );
  XNOR2X2_HVT U1092 ( .A1(in[3]), .A2(n1130), .Y(n1251) );
  INVX1_HVT U1093 ( .A(n1130), .Y(n1131) );
  AND2X1_HVT U1094 ( .A1(n782), .A2(n222), .Y(n1050) );
  XOR3X2_HVT U1095 ( .A1(n613), .A2(n1051), .A3(n100), .Y(out1[101]) );
  XNOR2X2_HVT U1096 ( .A1(n264), .A2(n1352), .Y(n308) );
  XNOR2X2_HVT U1097 ( .A1(n374), .A2(n1054), .Y(n469) );
  INVX1_HVT U1098 ( .A(n1540), .Y(n1056) );
  INVX1_HVT U1099 ( .A(in[4]), .Y(n1516) );
  XOR3X2_HVT U1100 ( .A1(n435), .A2(n1385), .A3(n404), .Y(n1416) );
  IBUFFX2_HVT U1101 ( .A(n253), .Y(n1057) );
  XNOR2X2_HVT U1102 ( .A1(n168), .A2(n1182), .Y(n116) );
  IBUFFX2_HVT U1103 ( .A(n374), .Y(n1058) );
  INVX0_HVT U1104 ( .A(n221), .Y(n1267) );
  IBUFFX2_HVT U1105 ( .A(n1251), .Y(n1207) );
  XOR3X2_HVT U1106 ( .A1(n1060), .A2(n572), .A3(n524), .Y(out1[114]) );
  IBUFFX2_HVT U1107 ( .A(n719), .Y(n1434) );
  XOR3X2_HVT U1108 ( .A1(n1061), .A2(n523), .A3(n524), .Y(out1[122]) );
  XOR3X2_HVT U1109 ( .A1(n525), .A2(n1089), .A3(n526), .Y(n1061) );
  XNOR2X2_HVT U1110 ( .A1(n292), .A2(n241), .Y(n351) );
  XNOR2X2_HVT U1111 ( .A1(n1351), .A2(n1533), .Y(n254) );
  NAND2X0_HVT U1112 ( .A1(n866), .A2(n70), .Y(n1063) );
  NAND2X0_HVT U1113 ( .A1(n1062), .A2(n867), .Y(n1064) );
  NAND2X0_HVT U1114 ( .A1(n1064), .A2(n1063), .Y(n520) );
  INVX0_HVT U1115 ( .A(n70), .Y(n1062) );
  XOR3X2_HVT U1116 ( .A1(n591), .A2(n1065), .A3(n592), .Y(out1[110]) );
  NAND2X0_HVT U1117 ( .A1(n359), .A2(n1326), .Y(n1067) );
  NAND2X0_HVT U1118 ( .A1(n1066), .A2(n747), .Y(n1068) );
  NAND2X0_HVT U1119 ( .A1(n1067), .A2(n1068), .Y(n314) );
  INVX0_HVT U1120 ( .A(n1326), .Y(n1066) );
  INVX1_HVT U1121 ( .A(n748), .Y(n1069) );
  XNOR2X2_HVT U1122 ( .A1(n1071), .A2(n1499), .Y(n439) );
  XNOR3X1_HVT U1123 ( .A1(n1541), .A2(n1390), .A3(n176), .Y(n231) );
  INVX1_HVT U1124 ( .A(n1187), .Y(n1072) );
  INVX0_HVT U1125 ( .A(n889), .Y(n1432) );
  XOR3X2_HVT U1126 ( .A1(n1275), .A2(n1073), .A3(n308), .Y(n358) );
  NAND2X0_HVT U1127 ( .A1(n605), .A2(n1286), .Y(n1074) );
  NAND2X0_HVT U1128 ( .A1(n1076), .A2(n1091), .Y(n1075) );
  NAND2X0_HVT U1129 ( .A1(n1074), .A2(n1075), .Y(n510) );
  AND2X1_HVT U1130 ( .A1(n1092), .A2(n807), .Y(n1076) );
  XOR3X2_HVT U1131 ( .A1(n391), .A2(n925), .A3(n364), .Y(out1[34]) );
  IBUFFX2_HVT U1132 ( .A(n1294), .Y(n1150) );
  XNOR2X2_HVT U1133 ( .A1(n254), .A2(n1080), .Y(n287) );
  XNOR2X2_HVT U1134 ( .A1(n269), .A2(n20), .Y(n276) );
  INVX0_HVT U1135 ( .A(n117), .Y(n1501) );
  XOR3X2_HVT U1136 ( .A1(n588), .A2(n610), .A3(n1493), .Y(out1[103]) );
  NAND2X0_HVT U1137 ( .A1(in[97]), .A2(n730), .Y(n1082) );
  NAND2X0_HVT U1138 ( .A1(n1225), .A2(n1543), .Y(n1083) );
  INVX0_HVT U1139 ( .A(n730), .Y(n1081) );
  NAND2X0_HVT U1140 ( .A1(n415), .A2(n1214), .Y(n1084) );
  NAND2X0_HVT U1141 ( .A1(n1087), .A2(n1212), .Y(n1085) );
  NAND2X0_HVT U1142 ( .A1(n1084), .A2(n1085), .Y(n1427) );
  IBUFFX2_HVT U1143 ( .A(n1404), .Y(n1086) );
  AND2X1_HVT U1144 ( .A1(n917), .A2(n1459), .Y(n1087) );
  NAND2X0_HVT U1145 ( .A1(in[121]), .A2(n13), .Y(n1091) );
  NAND2X0_HVT U1146 ( .A1(n1092), .A2(n1091), .Y(n605) );
  XNOR2X2_HVT U1147 ( .A1(in[17]), .A2(n981), .Y(n473) );
  NAND2X0_HVT U1148 ( .A1(n1242), .A2(in[120]), .Y(n1095) );
  NAND2X0_HVT U1149 ( .A1(n1094), .A2(n1241), .Y(n1096) );
  NAND2X0_HVT U1150 ( .A1(n1095), .A2(n1096), .Y(n70) );
  XNOR2X2_HVT U1151 ( .A1(n513), .A2(n1097), .Y(n543) );
  XOR3X1_HVT U1152 ( .A1(n1098), .A2(n132), .A3(n133), .Y(out1[86]) );
  NAND2X0_HVT U1153 ( .A1(n1516), .A2(n324), .Y(n1100) );
  NAND2X0_HVT U1154 ( .A1(n1099), .A2(n1463), .Y(n1101) );
  NAND2X0_HVT U1155 ( .A1(n1101), .A2(n1100), .Y(n456) );
  INVX1_HVT U1156 ( .A(n324), .Y(n1099) );
  INVX0_HVT U1157 ( .A(in[127]), .Y(n1241) );
  XOR3X1_HVT U1158 ( .A1(n1102), .A2(n166), .A3(n167), .Y(out1[81]) );
  XNOR2X1_HVT U1159 ( .A1(n661), .A2(n733), .Y(n151) );
  XOR3X2_HVT U1160 ( .A1(n135), .A2(n1183), .A3(n89), .Y(n187) );
  NAND2X0_HVT U1161 ( .A1(n140), .A2(n1104), .Y(n1105) );
  NAND2X0_HVT U1162 ( .A1(n1103), .A2(n141), .Y(n1106) );
  NAND2X0_HVT U1163 ( .A1(n1105), .A2(n1106), .Y(n90) );
  XNOR2X2_HVT U1164 ( .A1(n1376), .A2(n1536), .Y(n206) );
  NAND2X0_HVT U1165 ( .A1(in[113]), .A2(n1142), .Y(n1109) );
  NAND2X0_HVT U1166 ( .A1(n1107), .A2(n1108), .Y(n1110) );
  INVX0_HVT U1167 ( .A(in[113]), .Y(n1107) );
  XOR3X1_HVT U1168 ( .A1(n1378), .A2(n126), .A3(n85), .Y(n133) );
  XNOR2X2_HVT U1169 ( .A1(n1363), .A2(n1378), .Y(n140) );
  INVX0_HVT U1170 ( .A(n1537), .Y(n1502) );
  INVX1_HVT U1171 ( .A(n163), .Y(n1162) );
  INVX1_HVT U1172 ( .A(n1258), .Y(n1144) );
  XOR3X2_HVT U1173 ( .A1(n400), .A2(n1113), .A3(n445), .Y(out1[22]) );
  XOR3X2_HVT U1174 ( .A1(n392), .A2(n1114), .A3(n368), .Y(out1[33]) );
  NAND2X0_HVT U1175 ( .A1(n146), .A2(n1116), .Y(n1117) );
  NAND2X0_HVT U1176 ( .A1(n1115), .A2(n145), .Y(n1118) );
  NAND2X0_HVT U1177 ( .A1(n1117), .A2(n1118), .Y(n1373) );
  INVX0_HVT U1178 ( .A(n1210), .Y(n1119) );
  INVX1_HVT U1179 ( .A(n1099), .Y(n1120) );
  NAND2X0_HVT U1180 ( .A1(n1150), .A2(n1317), .Y(n1121) );
  NAND2X0_HVT U1181 ( .A1(n1153), .A2(n969), .Y(n1122) );
  NAND2X0_HVT U1182 ( .A1(n1122), .A2(n1123), .Y(n1152) );
  AND2X1_HVT U1183 ( .A1(n1317), .A2(n1134), .Y(n1123) );
  XOR3X2_HVT U1184 ( .A1(n318), .A2(n1140), .A3(n268), .Y(n317) );
  XNOR2X2_HVT U1185 ( .A1(n354), .A2(n1126), .Y(n301) );
  XNOR2X2_HVT U1186 ( .A1(n463), .A2(n1187), .Y(n374) );
  INVX0_HVT U1187 ( .A(n531), .Y(n1127) );
  INVX0_HVT U1188 ( .A(n1427), .Y(n1235) );
  NAND2X0_HVT U1189 ( .A1(n1397), .A2(n1142), .Y(n1132) );
  NAND2X0_HVT U1190 ( .A1(n1034), .A2(n1440), .Y(n1133) );
  NAND2X0_HVT U1191 ( .A1(n965), .A2(n424), .Y(n1134) );
  NAND2X0_HVT U1192 ( .A1(n1153), .A2(n969), .Y(n1135) );
  NAND2X0_HVT U1193 ( .A1(n1135), .A2(n1134), .Y(n1294) );
  XNOR2X2_HVT U1194 ( .A1(n59), .A2(n1315), .Y(n515) );
  NAND2X0_HVT U1195 ( .A1(n1467), .A2(n1475), .Y(n1138) );
  NAND2X0_HVT U1196 ( .A1(n1136), .A2(n1137), .Y(n1139) );
  NAND2X0_HVT U1197 ( .A1(n1138), .A2(n1139), .Y(out1[116]) );
  INVX0_HVT U1198 ( .A(n1467), .Y(n1136) );
  INVX0_HVT U1199 ( .A(n1475), .Y(n1137) );
  XNOR2X2_HVT U1200 ( .A1(n1510), .A2(n1288), .Y(n124) );
  INVX1_HVT U1201 ( .A(n579), .Y(n1219) );
  NAND2X0_HVT U1202 ( .A1(n667), .A2(n1155), .Y(n1141) );
  NAND2X0_HVT U1203 ( .A1(n1156), .A2(n1141), .Y(n1143) );
  NAND2X0_HVT U1204 ( .A1(n1258), .A2(n1498), .Y(n1146) );
  NAND2X0_HVT U1205 ( .A1(n1144), .A2(n1145), .Y(n1147) );
  NAND2X0_HVT U1206 ( .A1(n1147), .A2(n1146), .Y(n471) );
  INVX0_HVT U1207 ( .A(n1499), .Y(n1145) );
  NAND2X0_HVT U1208 ( .A1(n1121), .A2(n1151), .Y(n1148) );
  INVX0_HVT U1209 ( .A(n479), .Y(n1258) );
  INVX1_HVT U1210 ( .A(n229), .Y(n1149) );
  NAND2X0_HVT U1211 ( .A1(n1294), .A2(n1318), .Y(n1151) );
  NAND2X0_HVT U1212 ( .A1(n1151), .A2(n1152), .Y(n375) );
  INVX1_HVT U1213 ( .A(n1153), .Y(n1154) );
  NAND2X0_HVT U1214 ( .A1(n783), .A2(n665), .Y(n1156) );
  NAND2X0_HVT U1215 ( .A1(n667), .A2(n1155), .Y(n1157) );
  NAND2X0_HVT U1216 ( .A1(n1156), .A2(n1157), .Y(n195) );
  XOR3X1_HVT U1217 ( .A1(n1158), .A2(n580), .A3(n608), .Y(out1[105]) );
  XNOR2X2_HVT U1218 ( .A1(n366), .A2(n1149), .Y(n319) );
  XOR3X1_HVT U1219 ( .A1(n1518), .A2(n1247), .A3(n113), .Y(n617) );
  XOR3X2_HVT U1220 ( .A1(n1159), .A2(n1160), .A3(n51), .Y(n461) );
  XNOR2X2_HVT U1221 ( .A1(n253), .A2(n1444), .Y(n242) );
  XOR3X2_HVT U1222 ( .A1(n1220), .A2(n460), .A3(n461), .Y(out1[1]) );
  XNOR2X2_HVT U1223 ( .A1(n253), .A2(n1456), .Y(n292) );
  XNOR2X2_HVT U1224 ( .A1(n1329), .A2(n1200), .Y(n468) );
  XOR3X2_HVT U1225 ( .A1(n164), .A2(n1161), .A3(n1162), .Y(n108) );
  XOR2X2_HVT U1226 ( .A1(n1176), .A2(n202), .Y(n105) );
  XNOR2X2_HVT U1227 ( .A1(n566), .A2(n1163), .Y(n61) );
  XNOR3X2_HVT U1228 ( .A1(n546), .A2(n1542), .A3(n506), .Y(n592) );
  INVX1_HVT U1229 ( .A(n1164), .Y(n1165) );
  NAND2X0_HVT U1230 ( .A1(n1166), .A2(n782), .Y(n1468) );
  XOR3X2_HVT U1231 ( .A1(n104), .A2(n1168), .A3(n105), .Y(n1474) );
  NAND2X0_HVT U1232 ( .A1(n1177), .A2(n1178), .Y(n1169) );
  XNOR2X2_HVT U1233 ( .A1(n149), .A2(n1170), .Y(n141) );
  XOR3X1_HVT U1234 ( .A1(n518), .A2(n1323), .A3(n603), .Y(out1[107]) );
  XNOR2X2_HVT U1235 ( .A1(n448), .A2(n1402), .Y(n217) );
  XOR2X2_HVT U1236 ( .A1(n779), .A2(n868), .Y(n87) );
  XOR3X2_HVT U1237 ( .A1(n189), .A2(n1174), .A3(n631), .Y(out1[77]) );
  XNOR2X2_HVT U1238 ( .A1(n188), .A2(n1390), .Y(n135) );
  XOR3X2_HVT U1239 ( .A1(n1175), .A2(n528), .A3(n529), .Y(out1[121]) );
  NAND2X0_HVT U1240 ( .A1(n1164), .A2(n1183), .Y(n1177) );
  NAND2X0_HVT U1241 ( .A1(n1177), .A2(n1178), .Y(n1191) );
  AND2X1_HVT U1242 ( .A1(n1184), .A2(n1189), .Y(n1178) );
  IBUFFX2_HVT U1243 ( .A(n1232), .Y(n1189) );
  NAND2X0_HVT U1244 ( .A1(in[98]), .A2(n1544), .Y(n1180) );
  NAND2X0_HVT U1245 ( .A1(n1179), .A2(n885), .Y(n1181) );
  NBUFFX2_HVT U1246 ( .A(n161), .Y(n1182) );
  IBUFFX2_HVT U1247 ( .A(n459), .Y(n1220) );
  NAND2X0_HVT U1248 ( .A1(n228), .A2(n1201), .Y(n1184) );
  NAND2X0_HVT U1249 ( .A1(n1164), .A2(n1183), .Y(n1185) );
  NAND2X0_HVT U1250 ( .A1(n1185), .A2(n1184), .Y(n199) );
  INVX0_HVT U1251 ( .A(n765), .Y(n1188) );
  IBUFFX2_HVT U1252 ( .A(n337), .Y(n1446) );
  XNOR2X2_HVT U1253 ( .A1(in[96]), .A2(n1544), .Y(n577) );
  XNOR2X1_HVT U1254 ( .A1(n853), .A2(n774), .Y(n307) );
  XNOR2X2_HVT U1255 ( .A1(n593), .A2(n1081), .Y(n546) );
  XNOR2X2_HVT U1256 ( .A1(n377), .A2(n1437), .Y(n1209) );
  INVX1_HVT U1257 ( .A(n1292), .Y(n1187) );
  INVX1_HVT U1258 ( .A(n1517), .Y(n1292) );
  NAND2X0_HVT U1259 ( .A1(n199), .A2(n1232), .Y(n1190) );
  XNOR3X1_HVT U1260 ( .A1(n237), .A2(n238), .A3(n239), .Y(out1[62]) );
  XNOR2X2_HVT U1261 ( .A1(n418), .A2(n1506), .Y(n401) );
  XNOR2X1_HVT U1262 ( .A1(n724), .A2(n1542), .Y(n586) );
  XOR3X2_HVT U1263 ( .A1(n1331), .A2(n1160), .A3(n431), .Y(out1[25]) );
  XNOR2X2_HVT U1264 ( .A1(n465), .A2(n1304), .Y(n1195) );
  IBUFFX2_HVT U1265 ( .A(n465), .Y(n1505) );
  NBUFFX2_HVT U1266 ( .A(in[95]), .Y(n1196) );
  XOR3X1_HVT U1267 ( .A1(n1539), .A2(n78), .A3(n85), .Y(n84) );
  INVX1_HVT U1268 ( .A(in[103]), .Y(n1544) );
  XNOR2X2_HVT U1269 ( .A1(n50), .A2(n1297), .Y(n470) );
  IBUFFX2_HVT U1270 ( .A(n1329), .Y(n1202) );
  NAND2X0_HVT U1271 ( .A1(n1316), .A2(n413), .Y(n1204) );
  NAND2X0_HVT U1272 ( .A1(n412), .A2(n1203), .Y(n1205) );
  NAND2X0_HVT U1273 ( .A1(n1204), .A2(n1205), .Y(out1[28]) );
  INVX0_HVT U1274 ( .A(n413), .Y(n1203) );
  XOR3X2_HVT U1275 ( .A1(n975), .A2(n1260), .A3(n488), .Y(out1[13]) );
  XNOR2X2_HVT U1276 ( .A1(n1131), .A2(n1518), .Y(n403) );
  INVX1_HVT U1277 ( .A(n477), .Y(n1415) );
  XNOR2X2_HVT U1278 ( .A1(in[33]), .A2(in[38]), .Y(n388) );
  XNOR2X1_HVT U1279 ( .A1(n918), .A2(n418), .Y(n450) );
  INVX1_HVT U1280 ( .A(in[30]), .Y(n1524) );
  XOR3X2_HVT U1281 ( .A1(n1207), .A2(n1208), .A3(n325), .Y(n1486) );
  XOR2X1_HVT U1282 ( .A1(n913), .A2(n722), .Y(n426) );
  INVX1_HVT U1283 ( .A(n1524), .Y(n1437) );
  XNOR2X2_HVT U1284 ( .A1(n1436), .A2(in[5]), .Y(n462) );
  XNOR2X2_HVT U1285 ( .A1(n1209), .A2(n1438), .Y(n452) );
  NAND2X0_HVT U1286 ( .A1(n1210), .A2(n323), .Y(n1212) );
  NAND2X0_HVT U1287 ( .A1(n1212), .A2(n38), .Y(n415) );
  INVX0_HVT U1288 ( .A(n415), .Y(n1310) );
  NAND2X0_HVT U1289 ( .A1(n1486), .A2(n1322), .Y(n1217) );
  NAND2X0_HVT U1290 ( .A1(n1215), .A2(n1216), .Y(n1218) );
  NAND2X0_HVT U1291 ( .A1(n1217), .A2(n1218), .Y(out1[12]) );
  INVX0_HVT U1292 ( .A(n1486), .Y(n1215) );
  INVX0_HVT U1293 ( .A(n1322), .Y(n1216) );
  XOR3X2_HVT U1294 ( .A1(n578), .A2(n1219), .A3(n529), .Y(out1[113]) );
  XNOR2X2_HVT U1295 ( .A1(n574), .A2(n932), .Y(n65) );
  XOR3X2_HVT U1296 ( .A1(n1466), .A2(n860), .A3(n946), .Y(n1478) );
  NAND2X0_HVT U1297 ( .A1(in[16]), .A2(n1221), .Y(n1222) );
  NAND2X0_HVT U1298 ( .A1(n1223), .A2(n1222), .Y(n479) );
  INVX1_HVT U1299 ( .A(n1225), .Y(n1226) );
  XNOR3X1_HVT U1300 ( .A1(n56), .A2(n328), .A3(n458), .Y(n453) );
  XNOR2X2_HVT U1301 ( .A1(n1283), .A2(n49), .Y(n370) );
  XNOR2X2_HVT U1302 ( .A1(in[99]), .A2(n1544), .Y(n593) );
  XOR2X2_HVT U1303 ( .A1(n125), .A2(n77), .Y(n183) );
  XNOR2X2_HVT U1304 ( .A1(n1538), .A2(n1056), .Y(n77) );
  NAND2X0_HVT U1305 ( .A1(n1235), .A2(n450), .Y(n1229) );
  NAND2X0_HVT U1306 ( .A1(n1230), .A2(n1229), .Y(n1399) );
  AND2X1_HVT U1307 ( .A1(n1236), .A2(n1231), .Y(n1230) );
  INVX0_HVT U1308 ( .A(n453), .Y(n1231) );
  XNOR2X2_HVT U1309 ( .A1(n516), .A2(in[108]), .Y(n500) );
  XNOR2X2_HVT U1310 ( .A1(in[0]), .A2(n1027), .Y(n463) );
  NAND2X0_HVT U1311 ( .A1(n1427), .A2(n1406), .Y(n1236) );
  NAND2X0_HVT U1312 ( .A1(n1235), .A2(n450), .Y(n1237) );
  NAND2X0_HVT U1313 ( .A1(n1237), .A2(n1236), .Y(n1484) );
  XNOR2X2_HVT U1314 ( .A1(n463), .A2(n1262), .Y(n406) );
  XNOR2X2_HVT U1315 ( .A1(n575), .A2(n1240), .Y(n526) );
  XOR3X2_HVT U1316 ( .A1(n186), .A2(n1238), .A3(n187), .Y(out1[78]) );
  XOR3X2_HVT U1317 ( .A1(n548), .A2(n1043), .A3(n861), .Y(n1467) );
  XOR3X2_HVT U1318 ( .A1(n1430), .A2(n192), .A3(n549), .Y(out1[117]) );
  IBUFFX2_HVT U1319 ( .A(in[114]), .Y(n1239) );
  INVX1_HVT U1320 ( .A(n1239), .Y(n1240) );
  XOR3X2_HVT U1321 ( .A1(n1463), .A2(n399), .A3(n259), .Y(n488) );
  NAND2X0_HVT U1322 ( .A1(n777), .A2(n1248), .Y(n1243) );
  XNOR2X2_HVT U1323 ( .A1(n583), .A2(n1278), .Y(n566) );
  INVX2_HVT U1324 ( .A(in[111]), .Y(n1276) );
  INVX1_HVT U1325 ( .A(n487), .Y(n1260) );
  IBUFFX2_HVT U1326 ( .A(n96), .Y(n1365) );
  XOR2X2_HVT U1327 ( .A1(n162), .A2(in[82]), .Y(n107) );
  XOR3X2_HVT U1328 ( .A1(n365), .A2(n319), .A3(n1346), .Y(n391) );
  NAND2X0_HVT U1329 ( .A1(n360), .A2(n227), .Y(n1249) );
  NAND2X0_HVT U1330 ( .A1(n777), .A2(n1248), .Y(n1250) );
  NAND2X0_HVT U1331 ( .A1(n1250), .A2(n1249), .Y(n312) );
  INVX0_HVT U1332 ( .A(in[43]), .Y(n1248) );
  XNOR2X2_HVT U1333 ( .A1(n336), .A2(n1343), .Y(n1269) );
  NAND2X0_HVT U1334 ( .A1(n1369), .A2(n1489), .Y(n1255) );
  NAND2X0_HVT U1335 ( .A1(n1253), .A2(n1254), .Y(n1256) );
  NAND2X0_HVT U1336 ( .A1(n1255), .A2(n1256), .Y(out1[84]) );
  INVX0_HVT U1337 ( .A(n1489), .Y(n1253) );
  INVX0_HVT U1338 ( .A(n1369), .Y(n1254) );
  IBUFFX2_HVT U1339 ( .A(n157), .Y(n1282) );
  INVX0_HVT U1340 ( .A(n137), .Y(n1500) );
  XOR3X2_HVT U1341 ( .A1(n535), .A2(n1257), .A3(n587), .Y(n75) );
  XNOR2X2_HVT U1342 ( .A1(n326), .A2(n1277), .Y(n446) );
  XOR3X2_HVT U1343 ( .A1(n398), .A2(n399), .A3(n711), .Y(out1[30]) );
  XNOR2X2_HVT U1344 ( .A1(n171), .A2(n1284), .Y(n154) );
  XOR3X2_HVT U1345 ( .A1(n1259), .A2(n428), .A3(n429), .Y(n425) );
  XNOR2X2_HVT U1346 ( .A1(n147), .A2(n1284), .Y(n86) );
  NBUFFX2_HVT U1347 ( .A(n1144), .Y(n1262) );
  IBUFFX2_HVT U1348 ( .A(n334), .Y(n1401) );
  NBUFFX2_HVT U1349 ( .A(in[113]), .Y(n1263) );
  XOR3X2_HVT U1350 ( .A1(n1265), .A2(n1264), .A3(n823), .Y(out1[123]) );
  XNOR2X2_HVT U1351 ( .A1(n582), .A2(n1263), .Y(n531) );
  XNOR2X2_HVT U1352 ( .A1(n305), .A2(n1268), .Y(n297) );
  INVX0_HVT U1353 ( .A(in[76]), .Y(n1426) );
  INVX0_HVT U1354 ( .A(n551), .Y(n1332) );
  INVX0_HVT U1355 ( .A(n1547), .Y(n1465) );
  INVX0_HVT U1356 ( .A(n1444), .Y(n1407) );
  INVX0_HVT U1357 ( .A(n1440), .Y(n1279) );
  INVX0_HVT U1358 ( .A(n1391), .Y(n1361) );
  INVX0_HVT U1359 ( .A(n162), .Y(n1391) );
  INVX1_HVT U1360 ( .A(n172), .Y(n1366) );
  INVX1_HVT U1361 ( .A(n222), .Y(n1460) );
  INVX0_HVT U1362 ( .A(n574), .Y(n1289) );
  XNOR3X1_HVT U1363 ( .A1(n129), .A2(n1290), .A3(n173), .Y(n214) );
  INVX0_HVT U1364 ( .A(n344), .Y(n1383) );
  INVX1_HVT U1365 ( .A(n379), .Y(n1453) );
  INVX0_HVT U1366 ( .A(n1516), .Y(n1463) );
  INVX1_HVT U1367 ( .A(n1536), .Y(n1510) );
  INVX1_HVT U1368 ( .A(n421), .Y(n1435) );
  INVX1_HVT U1369 ( .A(in[63]), .Y(n1533) );
  INVX0_HVT U1370 ( .A(in[60]), .Y(n1330) );
  INVX1_HVT U1371 ( .A(in[20]), .Y(n1420) );
  XNOR2X2_HVT U1372 ( .A1(n433), .A2(n1320), .Y(n464) );
  INVX0_HVT U1373 ( .A(n433), .Y(n1295) );
  XOR3X2_HVT U1374 ( .A1(n1511), .A2(n128), .A3(n81), .Y(n1271) );
  INVX1_HVT U1375 ( .A(n278), .Y(n1345) );
  XOR3X2_HVT U1376 ( .A1(n913), .A2(n1505), .A3(n464), .Y(n1272) );
  XNOR3X1_HVT U1377 ( .A1(n540), .A2(n1315), .A3(n585), .Y(n1493) );
  INVX1_HVT U1378 ( .A(n272), .Y(n1396) );
  XNOR2X2_HVT U1379 ( .A1(n333), .A2(n1309), .Y(n272) );
  XOR3X2_HVT U1380 ( .A1(n122), .A2(n994), .A3(n174), .Y(n212) );
  XNOR2X1_HVT U1381 ( .A1(n708), .A2(n1009), .Y(n295) );
  INVX0_HVT U1382 ( .A(n1009), .Y(n1403) );
  XOR3X2_HVT U1383 ( .A1(n1472), .A2(n1274), .A3(n790), .Y(out1[9]) );
  XNOR2X2_HVT U1384 ( .A1(in[80]), .A2(n1540), .Y(n171) );
  XNOR3X1_HVT U1385 ( .A1(n1281), .A2(n1315), .A3(n535), .Y(n532) );
  XNOR2X2_HVT U1386 ( .A1(n559), .A2(n942), .Y(n545) );
  XNOR2X2_HVT U1387 ( .A1(in[107]), .A2(n1276), .Y(n559) );
  XNOR2X2_HVT U1388 ( .A1(n1464), .A2(n821), .Y(n540) );
  INVX1_HVT U1389 ( .A(in[108]), .Y(n1464) );
  XOR2X2_HVT U1390 ( .A1(in[36]), .A2(n1342), .Y(n286) );
  XNOR3X1_HVT U1391 ( .A1(n942), .A2(n76), .A3(n498), .Y(n539) );
  INVX1_HVT U1392 ( .A(n1437), .Y(n1277) );
  XNOR2X2_HVT U1393 ( .A1(in[10]), .A2(n991), .Y(n472) );
  XOR3X2_HVT U1394 ( .A1(n930), .A2(n1520), .A3(n114), .Y(n1491) );
  XNOR2X2_HVT U1395 ( .A1(in[8]), .A2(n991), .Y(n50) );
  INVX0_HVT U1396 ( .A(n320), .Y(n1445) );
  INVX1_HVT U1397 ( .A(n87), .Y(n1344) );
  INVX1_HVT U1398 ( .A(n383), .Y(n1355) );
  XOR3X2_HVT U1399 ( .A1(n1279), .A2(n497), .A3(n498), .Y(n496) );
  XNOR2X2_HVT U1400 ( .A1(in[83]), .A2(n1055), .Y(n96) );
  XNOR2X2_HVT U1401 ( .A1(n514), .A2(n1545), .Y(n551) );
  XNOR2X2_HVT U1402 ( .A1(n103), .A2(n1290), .Y(n98) );
  INVX1_HVT U1403 ( .A(n412), .Y(n1316) );
  XNOR2X2_HVT U1404 ( .A1(n118), .A2(n870), .Y(n104) );
  NBUFFX2_HVT U1405 ( .A(in[125]), .Y(n1286) );
  INVX1_HVT U1406 ( .A(n1287), .Y(n1288) );
  IBUFFX2_HVT U1407 ( .A(in[35]), .Y(n1326) );
  NBUFFX2_HVT U1408 ( .A(in[94]), .Y(n1290) );
  NBUFFX2_HVT U1409 ( .A(in[94]), .Y(n1291) );
  XNOR2X2_HVT U1410 ( .A1(n328), .A2(n1072), .Y(n451) );
  XOR3X2_HVT U1411 ( .A1(n55), .A2(n1295), .A3(n735), .Y(n1331) );
  NBUFFX2_HVT U1412 ( .A(in[13]), .Y(n1296) );
  NBUFFX2_HVT U1413 ( .A(in[13]), .Y(n1297) );
  NBUFFX2_HVT U1414 ( .A(in[13]), .Y(n1298) );
  XNOR2X2_HVT U1415 ( .A1(n1301), .A2(n428), .Y(n55) );
  INVX1_HVT U1416 ( .A(n1094), .Y(n1302) );
  XOR3X2_HVT U1417 ( .A1(n612), .A2(n293), .A3(n250), .Y(n1480) );
  IBUFFX2_HVT U1418 ( .A(in[17]), .Y(n1304) );
  INVX1_HVT U1419 ( .A(n1304), .Y(n1305) );
  INVX1_HVT U1420 ( .A(n1310), .Y(n1311) );
  INVX1_HVT U1421 ( .A(n742), .Y(n1307) );
  IBUFFX2_HVT U1422 ( .A(in[49]), .Y(n1308) );
  INVX2_HVT U1423 ( .A(n1308), .Y(n1309) );
  XNOR2X2_HVT U1424 ( .A1(in[122]), .A2(n1550), .Y(n59) );
  XOR3X2_HVT U1425 ( .A1(n726), .A2(n1305), .A3(n477), .Y(n427) );
  XNOR2X2_HVT U1426 ( .A1(n1247), .A2(n1524), .Y(n428) );
  INVX1_HVT U1427 ( .A(n810), .Y(n1312) );
  XNOR2X2_HVT U1428 ( .A1(n560), .A2(n1431), .Y(n552) );
  INVX1_HVT U1429 ( .A(n1030), .Y(n1319) );
  XNOR2X2_HVT U1430 ( .A1(in[81]), .A2(n1394), .Y(n224) );
  XOR3X2_HVT U1431 ( .A1(n1167), .A2(n137), .A3(n1024), .Y(n1489) );
  XNOR2X2_HVT U1432 ( .A1(n157), .A2(n1324), .Y(n147) );
  NBUFFX2_HVT U1433 ( .A(in[25]), .Y(n1320) );
  XOR3X2_HVT U1434 ( .A1(n405), .A2(n1320), .A3(n406), .Y(n402) );
  XOR3X2_HVT U1435 ( .A1(n1119), .A2(n1512), .A3(n487), .Y(n1322) );
  XNOR2X2_HVT U1436 ( .A1(n348), .A2(n1526), .Y(n291) );
  XOR3X2_HVT U1437 ( .A1(n65), .A2(n1263), .A3(n573), .Y(n524) );
  XNOR2X2_HVT U1438 ( .A1(n600), .A2(n1464), .Y(n556) );
  XNOR2X2_HVT U1439 ( .A1(in[88]), .A2(n1541), .Y(n118) );
  XNOR2X2_HVT U1440 ( .A1(n1273), .A2(n464), .Y(n51) );
  XOR3X2_HVT U1441 ( .A1(n297), .A2(n1327), .A3(n238), .Y(n1353) );
  XNOR2X2_HVT U1442 ( .A1(n1429), .A2(n1522), .Y(n478) );
  XOR3X2_HVT U1443 ( .A1(n1072), .A2(n447), .A3(n218), .Y(n486) );
  NBUFFX2_HVT U1444 ( .A(in[55]), .Y(n1328) );
  XOR3X2_HVT U1445 ( .A1(n296), .A2(n1330), .A3(n288), .Y(n382) );
  NAND2X0_HVT U1446 ( .A1(n551), .A2(n1333), .Y(n1334) );
  NAND2X0_HVT U1447 ( .A1(n1332), .A2(n552), .Y(n1335) );
  NAND2X0_HVT U1448 ( .A1(n1334), .A2(n1335), .Y(n507) );
  NAND2X0_HVT U1449 ( .A1(n1337), .A2(n334), .Y(n1338) );
  NAND2X0_HVT U1450 ( .A1(n1336), .A2(n824), .Y(n1339) );
  NAND2X0_HVT U1451 ( .A1(n752), .A2(n1338), .Y(n360) );
  XNOR2X2_HVT U1452 ( .A1(n1363), .A2(n148), .Y(n190) );
  XNOR2X2_HVT U1453 ( .A1(in[114]), .A2(n1549), .Y(n564) );
  XNOR2X2_HVT U1454 ( .A1(n567), .A2(in[115]), .Y(n521) );
  XOR3X2_HVT U1455 ( .A1(n526), .A2(n1226), .A3(n572), .Y(n64) );
  XNOR2X2_HVT U1456 ( .A1(n564), .A2(n1440), .Y(n558) );
  XNOR2X1_HVT U1457 ( .A1(in[44]), .A2(n254), .Y(n238) );
  XNOR2X2_HVT U1458 ( .A1(n462), .A2(n1404), .Y(n53) );
  XOR3X2_HVT U1459 ( .A1(n1394), .A2(n1503), .A3(n123), .Y(n175) );
  XOR3X2_HVT U1460 ( .A1(n115), .A2(n116), .A3(n1501), .Y(out1[89]) );
  XOR3X2_HVT U1461 ( .A1(n277), .A2(n1345), .A3(n279), .Y(out1[56]) );
  IBUFFX2_HVT U1462 ( .A(in[57]), .Y(n1346) );
  XOR3X2_HVT U1463 ( .A1(n1407), .A2(n740), .A3(n620), .Y(n1347) );
  XOR3X2_HVT U1464 ( .A1(n1350), .A2(n1447), .A3(n358), .Y(out1[35]) );
  INVX1_HVT U1465 ( .A(n1497), .Y(n1357) );
  INVX1_HVT U1466 ( .A(n1351), .Y(n1352) );
  XOR3X2_HVT U1467 ( .A1(n1353), .A2(n1443), .A3(n351), .Y(out1[45]) );
  IBUFFX2_HVT U1468 ( .A(n254), .Y(n1444) );
  NAND2X0_HVT U1469 ( .A1(n1408), .A2(n1409), .Y(n1354) );
  XOR3X2_HVT U1470 ( .A1(n382), .A2(n1355), .A3(n351), .Y(out1[37]) );
  XNOR2X2_HVT U1471 ( .A1(n287), .A2(n926), .Y(n346) );
  NAND2X0_HVT U1472 ( .A1(n1354), .A2(n1410), .Y(n1360) );
  XNOR2X2_HVT U1473 ( .A1(n1330), .A2(n879), .Y(n233) );
  XOR3X2_HVT U1474 ( .A1(n1361), .A2(n1093), .A3(n108), .Y(n1482) );
  XOR3X2_HVT U1475 ( .A1(n134), .A2(n1362), .A3(n139), .Y(n215) );
  XNOR2X2_HVT U1476 ( .A1(n92), .A2(n1364), .Y(out1[92]) );
  INVX2_HVT U1477 ( .A(in[78]), .Y(n1536) );
  XOR3X2_HVT U1478 ( .A1(n210), .A2(n12), .A3(n120), .Y(n1367) );
  XOR3X2_HVT U1479 ( .A1(n1471), .A2(n988), .A3(n198), .Y(out1[67]) );
  INVX1_HVT U1480 ( .A(n1103), .Y(n1368) );
  XOR3X2_HVT U1481 ( .A1(n26), .A2(n1312), .A3(n149), .Y(n1369) );
  XNOR2X2_HVT U1482 ( .A1(n1358), .A2(n1497), .Y(n269) );
  XOR3X2_HVT U1483 ( .A1(n176), .A2(n1056), .A3(n177), .Y(n123) );
  XOR3X2_HVT U1484 ( .A1(n1490), .A2(n1406), .A3(n1040), .Y(out1[21]) );
  XNOR2X2_HVT U1485 ( .A1(n493), .A2(n1438), .Y(n419) );
  XOR3X2_HVT U1486 ( .A1(n101), .A2(n1372), .A3(n152), .Y(n198) );
  XNOR2X2_HVT U1487 ( .A1(n136), .A2(n86), .Y(n191) );
  XNOR2X2_HVT U1488 ( .A1(n148), .A2(n1510), .Y(n134) );
  INVX1_HVT U1489 ( .A(n202), .Y(n1377) );
  AND2X1_HVT U1490 ( .A1(n1379), .A2(n616), .Y(n1375) );
  XNOR2X2_HVT U1491 ( .A1(n200), .A2(n19), .Y(n156) );
  INVX1_HVT U1492 ( .A(n898), .Y(n1376) );
  NAND2X0_HVT U1493 ( .A1(n202), .A2(n1378), .Y(n1379) );
  NAND2X0_HVT U1494 ( .A1(n1377), .A2(n1495), .Y(n1380) );
  NAND2X0_HVT U1495 ( .A1(n1380), .A2(n1379), .Y(n194) );
  XNOR2X1_HVT U1496 ( .A1(n1494), .A2(n887), .Y(n176) );
  XOR3X2_HVT U1497 ( .A1(n1381), .A2(n924), .A3(n198), .Y(out1[75]) );
  XOR3X2_HVT U1498 ( .A1(n200), .A2(n952), .A3(n105), .Y(n1381) );
  XNOR2X2_HVT U1499 ( .A1(n1494), .A2(n1536), .Y(n210) );
  XNOR2X2_HVT U1500 ( .A1(n581), .A2(n941), .Y(n71) );
  XNOR2X2_HVT U1501 ( .A1(n1278), .A2(n1393), .Y(n581) );
  XOR3X2_HVT U1502 ( .A1(n1383), .A2(n346), .A3(n347), .Y(out1[46]) );
  XNOR2X2_HVT U1503 ( .A1(in[58]), .A2(n1533), .Y(n263) );
  NBUFFX2_HVT U1504 ( .A(n1245), .Y(n1384) );
  NBUFFX2_HVT U1505 ( .A(in[9]), .Y(n1385) );
  XOR3X2_HVT U1506 ( .A1(n1387), .A2(n1386), .A3(n1299), .Y(out1[99]) );
  XOR3X2_HVT U1507 ( .A1(n59), .A2(n60), .A3(n61), .Y(n1387) );
  XOR3X2_HVT U1508 ( .A1(n1233), .A2(n83), .A3(n141), .Y(n189) );
  XNOR2X2_HVT U1509 ( .A1(n225), .A2(n1389), .Y(n149) );
  INVX1_HVT U1510 ( .A(n1534), .Y(n1389) );
  NBUFFX2_HVT U1511 ( .A(n766), .Y(n1433) );
  XNOR2X2_HVT U1512 ( .A1(in[66]), .A2(n1535), .Y(n225) );
  INVX1_HVT U1513 ( .A(n1546), .Y(n1393) );
  XNOR2X2_HVT U1514 ( .A1(n196), .A2(in[68]), .Y(n146) );
  XNOR3X2_HVT U1515 ( .A1(n130), .A2(n1390), .A3(n124), .Y(n185) );
  XNOR2X2_HVT U1516 ( .A1(n290), .A2(n291), .Y(n240) );
  XOR3X2_HVT U1517 ( .A1(in[44]), .A2(n295), .A3(n245), .Y(n1395) );
  XNOR2X2_HVT U1518 ( .A1(n226), .A2(n1201), .Y(n196) );
  XNOR2X2_HVT U1519 ( .A1(n1034), .A2(in[115]), .Y(n513) );
  XOR3X2_HVT U1520 ( .A1(n271), .A2(n1396), .A3(n27), .Y(out1[57]) );
  XNOR2X2_HVT U1521 ( .A1(n1529), .A2(in[40]), .Y(n334) );
  NBUFFX2_HVT U1522 ( .A(in[119]), .Y(n1397) );
  NAND2X0_HVT U1523 ( .A1(n453), .A2(n1484), .Y(n1398) );
  NAND2X0_HVT U1524 ( .A1(n1398), .A2(n1399), .Y(out1[20]) );
  XNOR2X2_HVT U1525 ( .A1(n939), .A2(n1244), .Y(n366) );
  XOR3X2_HVT U1526 ( .A1(n244), .A2(n1403), .A3(n245), .Y(n243) );
  XOR3X2_HVT U1527 ( .A1(n452), .A2(n1519), .A3(n219), .Y(n1490) );
  XNOR2X2_HVT U1528 ( .A1(n1404), .A2(in[6]), .Y(n474) );
  NAND2X0_HVT U1529 ( .A1(n1330), .A2(n248), .Y(n1410) );
  NAND2X0_HVT U1530 ( .A1(n1408), .A2(n1409), .Y(n1411) );
  NAND2X0_HVT U1531 ( .A1(n1411), .A2(n1410), .Y(n300) );
  INVX0_HVT U1532 ( .A(n248), .Y(n1408) );
  INVX1_HVT U1533 ( .A(n1330), .Y(n1409) );
  NAND2X0_HVT U1534 ( .A1(n1532), .A2(n1455), .Y(n1412) );
  INVX0_HVT U1535 ( .A(n300), .Y(n1513) );
  XNOR2X2_HVT U1536 ( .A1(n210), .A2(n1413), .Y(n170) );
  NBUFFX2_HVT U1537 ( .A(in[73]), .Y(n1413) );
  XOR3X2_HVT U1538 ( .A1(n272), .A2(n748), .A3(n331), .Y(n368) );
  XOR3X1_HVT U1539 ( .A1(n1414), .A2(n1415), .A3(n1416), .Y(out1[10]) );
  NBUFFX2_HVT U1540 ( .A(in[54]), .Y(n1417) );
  XNOR2X2_HVT U1541 ( .A1(n455), .A2(n1420), .Y(n414) );
  XOR3X2_HVT U1542 ( .A1(n193), .A2(n500), .A3(n552), .Y(n1424) );
  XNOR2X2_HVT U1543 ( .A1(n458), .A2(n414), .Y(n325) );
  XOR3X2_HVT U1544 ( .A1(n170), .A2(n773), .A3(n172), .Y(n117) );
  XNOR2X2_HVT U1545 ( .A1(n169), .A2(n1378), .Y(n200) );
  IBUFFX2_HVT U1546 ( .A(n455), .Y(n1459) );
  XNOR2X2_HVT U1547 ( .A1(n1488), .A2(n1487), .Y(out1[76]) );
  IBUFFX2_HVT U1548 ( .A(in[103]), .Y(n1507) );
  XNOR2X2_HVT U1549 ( .A1(n1046), .A2(n1125), .Y(n561) );
  XOR3X2_HVT U1550 ( .A1(n531), .A2(n577), .A3(n579), .Y(n69) );
  XNOR2X2_HVT U1551 ( .A1(n327), .A2(n1498), .Y(n410) );
  XNOR2X2_HVT U1552 ( .A1(n388), .A2(n1525), .Y(n356) );
  XOR3X2_HVT U1553 ( .A1(n1550), .A2(n1293), .A3(n76), .Y(n1492) );
  NBUFFX2_HVT U1554 ( .A(in[6]), .Y(n1436) );
  XNOR2X2_HVT U1555 ( .A1(n602), .A2(in[100]), .Y(n557) );
  XOR2X2_HVT U1556 ( .A1(n54), .A2(n1385), .Y(n459) );
  NBUFFX2_HVT U1557 ( .A(in[29]), .Y(n1438) );
  NBUFFX2_HVT U1558 ( .A(in[29]), .Y(n1439) );
  XNOR2X2_HVT U1559 ( .A1(n489), .A2(n1436), .Y(n328) );
  XNOR2X2_HVT U1560 ( .A1(n474), .A2(n1517), .Y(n324) );
  XNOR2X2_HVT U1561 ( .A1(n419), .A2(n1523), .Y(n458) );
  XNOR2X2_HVT U1562 ( .A1(n1055), .A2(in[82]), .Y(n157) );
  XNOR2X2_HVT U1563 ( .A1(n472), .A2(n1402), .Y(n417) );
  NBUFFX2_HVT U1564 ( .A(in[118]), .Y(n1440) );
  XOR2X2_HVT U1565 ( .A1(n416), .A2(n326), .Y(n408) );
  XNOR2X2_HVT U1566 ( .A1(n561), .A2(in[116]), .Y(n511) );
  XNOR2X2_HVT U1567 ( .A1(n510), .A2(n1199), .Y(n555) );
  XOR3X2_HVT U1568 ( .A1(n363), .A2(n1445), .A3(n364), .Y(out1[42]) );
  XOR3X2_HVT U1569 ( .A1(n367), .A2(n1446), .A3(n368), .Y(out1[41]) );
  XOR3X2_HVT U1570 ( .A1(n1451), .A2(n8), .A3(n335), .Y(n392) );
  XOR3X2_HVT U1571 ( .A1(n1533), .A2(n1497), .A3(n280), .Y(n277) );
  XOR3X2_HVT U1572 ( .A1(n262), .A2(n207), .A3(n1454), .Y(out1[59]) );
  XOR3X2_HVT U1573 ( .A1(n265), .A2(n997), .A3(n634), .Y(n1454) );
  NAND2X0_HVT U1574 ( .A1(n1456), .A2(n361), .Y(n1457) );
  NAND2X0_HVT U1575 ( .A1(n1455), .A2(n1532), .Y(n1458) );
  NAND2X0_HVT U1576 ( .A1(n1458), .A2(n1457), .Y(n248) );
  INVX1_HVT U1577 ( .A(n361), .Y(n1455) );
  XNOR2X2_HVT U1578 ( .A1(n263), .A2(n1496), .Y(n253) );
  XNOR2X2_HVT U1579 ( .A1(n274), .A2(in[61]), .Y(n264) );
  XNOR2X2_HVT U1580 ( .A1(in[56]), .A2(n1452), .Y(n274) );
  XOR3X2_HVT U1581 ( .A1(n429), .A2(n1086), .A3(n476), .Y(n404) );
  NAND2X0_HVT U1582 ( .A1(n1166), .A2(n1050), .Y(n1461) );
  NAND2X0_HVT U1583 ( .A1(n1460), .A2(n1468), .Y(n1462) );
  NAND2X0_HVT U1584 ( .A1(n1461), .A2(n1462), .Y(out1[68]) );
  XOR3X2_HVT U1585 ( .A1(n378), .A2(n797), .A3(n469), .Y(n422) );
  XNOR2X2_HVT U1586 ( .A1(in[104]), .A2(n1276), .Y(n583) );
  XNOR2X2_HVT U1587 ( .A1(n563), .A2(n1393), .Y(n514) );
  XNOR2X2_HVT U1588 ( .A1(n606), .A2(n1545), .Y(n600) );
  XOR2X2_HVT U1589 ( .A1(n285), .A2(n286), .Y(n236) );
  XOR3X2_HVT U1590 ( .A1(n319), .A2(n1309), .A3(n320), .Y(n268) );
  XNOR2X2_HVT U1591 ( .A1(n370), .A2(n1140), .Y(n335) );
  XNOR2X2_HVT U1592 ( .A1(n356), .A2(in[36]), .Y(n302) );
  XOR2X2_HVT U1593 ( .A1(n397), .A2(n443), .Y(n182) );
  XOR2X2_HVT U1594 ( .A1(n281), .A2(n232), .Y(n343) );
  XOR3X2_HVT U1595 ( .A1(n335), .A2(n990), .A3(n337), .Y(n273) );
  XNOR2X2_HVT U1596 ( .A1(in[50]), .A2(n1531), .Y(n313) );
  XOR2X2_HVT U1597 ( .A1(n401), .A2(n446), .Y(n218) );
  XNOR2X2_HVT U1598 ( .A1(n468), .A2(n1506), .Y(n327) );
  XOR3X2_HVT U1599 ( .A1(n61), .A2(n955), .A3(n565), .Y(n519) );
  XOR3X2_HVT U1600 ( .A1(n65), .A2(n1089), .A3(n66), .Y(n1508) );
  XNOR2X2_HVT U1601 ( .A1(n473), .A2(n1498), .Y(n455) );
  XOR3X2_HVT U1602 ( .A1(n71), .A2(n1049), .A3(n580), .Y(n529) );
  XNOR2X2_HVT U1603 ( .A1(n545), .A2(n546), .Y(n502) );
  XNOR2X2_HVT U1604 ( .A1(n134), .A2(n135), .Y(n85) );
  XNOR2X2_HVT U1605 ( .A1(n540), .A2(n541), .Y(n498) );
  XNOR2X2_HVT U1606 ( .A1(in[106]), .A2(n1276), .Y(n563) );
  XNOR2X2_HVT U1607 ( .A1(in[73]), .A2(n1536), .Y(n202) );
  XOR3X2_HVT U1608 ( .A1(n1508), .A2(n63), .A3(n762), .Y(out1[98]) );
  XOR3X2_HVT U1609 ( .A1(n1470), .A2(n1318), .A3(n422), .Y(out1[19]) );
  XOR3X2_HVT U1610 ( .A1(n828), .A2(n919), .A3(n717), .Y(n1470) );
  XNOR2X2_HVT U1611 ( .A1(in[72]), .A2(n1537), .Y(n169) );
  XNOR2X2_HVT U1612 ( .A1(in[57]), .A2(in[62]), .Y(n361) );
  XOR3X2_HVT U1613 ( .A1(n71), .A2(n1006), .A3(n72), .Y(n67) );
  XNOR2X2_HVT U1614 ( .A1(in[75]), .A2(n1503), .Y(n148) );
  XOR2X1_HVT U1615 ( .A1(n687), .A2(n403), .Y(n460) );
  XNOR2X1_HVT U1616 ( .A1(n940), .A2(n760), .Y(n523) );
  XOR2X1_HVT U1617 ( .A1(n205), .A2(n162), .Y(n165) );
  XNOR2X1_HVT U1618 ( .A1(n188), .A2(n1538), .Y(n139) );
  XNOR2X1_HVT U1619 ( .A1(n593), .A2(n1547), .Y(n550) );
  XOR2X1_HVT U1620 ( .A1(n1165), .A2(n644), .Y(n159) );
  XNOR2X1_HVT U1621 ( .A1(n1390), .A2(n1539), .Y(n173) );
  XNOR2X1_HVT U1622 ( .A1(n1526), .A2(n1530), .Y(n338) );
  XOR3X1_HVT U1623 ( .A1(n159), .A2(n160), .A3(n1482), .Y(out1[82]) );
  XNOR2X1_HVT U1624 ( .A1(n559), .A2(in[124]), .Y(n506) );
  XNOR3X1_HVT U1625 ( .A1(n285), .A2(n1496), .A3(n338), .Y(n380) );
  XNOR3X1_HVT U1626 ( .A1(n1491), .A2(n112), .A3(n113), .Y(out1[8]) );
  XNOR2X1_HVT U1627 ( .A1(n304), .A2(in[60]), .Y(n244) );
  XNOR3X1_HVT U1628 ( .A1(n1492), .A2(n74), .A3(n75), .Y(out1[96]) );
  XOR2X1_HVT U1629 ( .A1(n428), .A2(n827), .Y(n476) );
  XNOR2X1_HVT U1630 ( .A1(in[69]), .A2(n1534), .Y(n209) );
  XNOR2X1_HVT U1631 ( .A1(n1522), .A2(n1292), .Y(n440) );
  XOR2X1_HVT U1632 ( .A1(n109), .A2(n841), .Y(n160) );
  XOR2X1_HVT U1633 ( .A1(in[101]), .A2(n1441), .Y(n76) );
  XOR2X1_HVT U1634 ( .A1(n119), .A2(n806), .Y(n166) );
  XOR2X1_HVT U1635 ( .A1(n63), .A2(n842), .Y(n573) );
  XNOR2X1_HVT U1636 ( .A1(n1199), .A2(n1286), .Y(n495) );
  XNOR2X1_HVT U1637 ( .A1(n1433), .A2(n1170), .Y(n177) );
  XNOR2X1_HVT U1638 ( .A1(n1302), .A2(n867), .Y(n587) );
  XNOR2X1_HVT U1639 ( .A1(n104), .A2(n636), .Y(n152) );
  XNOR2X1_HVT U1640 ( .A1(n1520), .A2(n1439), .Y(n437) );
  XNOR2X1_HVT U1641 ( .A1(n1298), .A2(n1266), .Y(n114) );
  XNOR2X1_HVT U1642 ( .A1(in[68]), .A2(n1170), .Y(n213) );
  XOR2X1_HVT U1643 ( .A1(n91), .A2(n1298), .Y(n482) );
  XNOR2X1_HVT U1644 ( .A1(in[92]), .A2(n1541), .Y(n125) );
  XNOR2X1_HVT U1645 ( .A1(n1547), .A2(n1125), .Y(n538) );
  XNOR2X1_HVT U1646 ( .A1(in[36]), .A2(n1268), .Y(n379) );
  XNOR2X1_HVT U1647 ( .A1(in[100]), .A2(n1542), .Y(n610) );
  XNOR2X1_HVT U1648 ( .A1(n1519), .A2(n1298), .Y(n484) );
  XNOR2X1_HVT U1649 ( .A1(n1234), .A2(n1288), .Y(n78) );
  XOR2X1_HVT U1650 ( .A1(n403), .A2(in[2]), .Y(n477) );
  XNOR2X1_HVT U1651 ( .A1(n448), .A2(in[28]), .Y(n407) );
  XNOR2X1_HVT U1652 ( .A1(n725), .A2(n1288), .Y(n174) );
  XNOR2X1_HVT U1653 ( .A1(in[80]), .A2(n1539), .Y(n122) );
  XNOR2X1_HVT U1654 ( .A1(in[4]), .A2(n1027), .Y(n444) );
  XNOR2X1_HVT U1655 ( .A1(n1538), .A2(n1284), .Y(n126) );
  XNOR2X1_HVT U1656 ( .A1(in[76]), .A2(n1376), .Y(n129) );
  XNOR2X1_HVT U1657 ( .A1(in[108]), .A2(n1545), .Y(n589) );
  XNOR2X1_HVT U1658 ( .A1(n1545), .A2(n1315), .Y(n497) );
  NBUFFX2_HVT U1659 ( .A(in[77]), .Y(n1494) );
  NBUFFX2_HVT U1660 ( .A(in[77]), .Y(n1495) );
  NBUFFX2_HVT U1661 ( .A(in[62]), .Y(n1496) );
  NBUFFX2_HVT U1662 ( .A(in[62]), .Y(n1497) );
  NBUFFX2_HVT U1663 ( .A(in[21]), .Y(n1498) );
  NBUFFX2_HVT U1664 ( .A(in[21]), .Y(n1499) );
  XOR2X1_HVT U1665 ( .A1(in[20]), .A2(n1498), .Y(n441) );
  XOR2X1_HVT U1666 ( .A1(in[76]), .A2(n1495), .Y(n184) );
  NBUFFX2_HVT U1667 ( .A(n981), .Y(n1506) );
  INVX1_HVT U1668 ( .A(n713), .Y(n1512) );
  XNOR2X1_HVT U1669 ( .A1(in[20]), .A2(n1429), .Y(n397) );
  XNOR2X1_HVT U1670 ( .A1(n1293), .A2(n1548), .Y(n585) );
  NAND2X0_HVT U1671 ( .A1(n1360), .A2(n1052), .Y(n1514) );
  NAND2X0_HVT U1672 ( .A1(n1513), .A2(n907), .Y(n1515) );
  NAND2X0_HVT U1673 ( .A1(n1515), .A2(n1514), .Y(n355) );
  XNOR2X1_HVT U1674 ( .A1(n1519), .A2(n992), .Y(n178) );
  XNOR2X1_HVT U1675 ( .A1(in[44]), .A2(n939), .Y(n285) );
  XOR2X1_HVT U1676 ( .A1(n1393), .A2(n1286), .Y(n533) );
  XNOR2X1_HVT U1677 ( .A1(n1523), .A2(n1247), .Y(n443) );
  XNOR2X1_HVT U1678 ( .A1(n1201), .A2(n1324), .Y(n128) );
endmodule

