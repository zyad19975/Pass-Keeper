
module inv_sbox_15 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n196, n197, n198, n199, n200, n201, n202, n208, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610;

  NAND2X0_HVT U1 ( .A1(n259), .A2(n201), .Y(n610) );
  NAND2X0_HVT U4 ( .A1(n279), .A2(n609), .Y(n607) );
  NAND2X0_HVT U5 ( .A1(n607), .A2(n322), .Y(n606) );
  NAND2X0_HVT U6 ( .A1(n328), .A2(n274), .Y(n604) );
  NAND2X0_HVT U7 ( .A1(n279), .A2(n323), .Y(n603) );
  NAND2X0_HVT U8 ( .A1(n280), .A2(n322), .Y(n602) );
  NAND2X0_HVT U9 ( .A1(n610), .A2(n602), .Y(n601) );
  NAND2X0_HVT U10 ( .A1(n274), .A2(n599), .Y(n600) );
  NAND2X0_HVT U11 ( .A1(n291), .A2(n327), .Y(n598) );
  NAND2X0_HVT U12 ( .A1(n328), .A2(n311), .Y(n597) );
  NAND2X0_HVT U13 ( .A1(n325), .A2(n602), .Y(n596) );
  NAND2X0_HVT U15 ( .A1(n319), .A2(n330), .Y(n594) );
  NAND2X0_HVT U19 ( .A1(n329), .A2(n399), .Y(n589) );
  NAND2X0_HVT U25 ( .A1(n292), .A2(n312), .Y(n605) );
  NAND2X0_HVT U32 ( .A1(n313), .A2(n218), .Y(n577) );
  NAND2X0_HVT U35 ( .A1(n602), .A2(n208), .Y(n574) );
  NAND2X0_HVT U38 ( .A1(n311), .A2(n239), .Y(n571) );
  NAND2X0_HVT U42 ( .A1(n604), .A2(n208), .Y(n567) );
  OA21X1_HVT U53 ( .A1(n338), .A2(n559), .A3(n366), .Y(n557) );
  NAND2X0_HVT U55 ( .A1(n324), .A2(n607), .Y(n555) );
  AO21X1_HVT U60 ( .A1(n549), .A2(n308), .A3(n588), .Y(n550) );
  MUX41X1_HVT U62 ( .A1(n548), .A3(n554), .A2(n552), .A4(n556), .S0(n318), 
        .S1(n257), .Y(n547) );
  MUX41X1_HVT U65 ( .A1(n358), .A3(n360), .A2(n359), .A4(n571), .S0(n304), 
        .S1(n335), .Y(n544) );
  NAND2X0_HVT U66 ( .A1(n330), .A2(n228), .Y(n543) );
  MUX41X1_HVT U67 ( .A1(n355), .A3(n382), .A2(n357), .A4(n543), .S0(n310), 
        .S1(n301), .Y(n542) );
  NAND2X0_HVT U72 ( .A1(n320), .A2(n603), .Y(n538) );
  MUX41X1_HVT U73 ( .A1(n582), .A3(n538), .A2(n383), .A4(n312), .S0(n309), 
        .S1(n300), .Y(n537) );
  MUX41X1_HVT U74 ( .A1(n600), .A3(n371), .A2(n370), .A4(n361), .S0(n304), 
        .S1(n334), .Y(n536) );
  MUX41X1_HVT U78 ( .A1(n533), .A3(n537), .A2(n536), .A4(n539), .S0(n318), 
        .S1(n257), .Y(n532) );
  MUX41X1_HVT U79 ( .A1(n367), .A3(n591), .A2(n369), .A4(n592), .S0(n304), 
        .S1(n334), .Y(n531) );
  MUX41X1_HVT U80 ( .A1(n385), .A3(n381), .A2(n601), .A4(n606), .S0(n303), 
        .S1(n336), .Y(n530) );
  NAND2X0_HVT U81 ( .A1(n327), .A2(n603), .Y(n529) );
  AND2X1_HVT U82 ( .A1(n241), .A2(n325), .Y(n528) );
  MUX41X1_HVT U83 ( .A1(n528), .A3(n368), .A2(n258), .A4(n529), .S0(n303), 
        .S1(n281), .Y(n527) );
  MUX41X1_HVT U84 ( .A1(n298), .A3(n367), .A2(n386), .A4(n243), .S0(n304), 
        .S1(n282), .Y(n526) );
  MUX41X1_HVT U85 ( .A1(n526), .A3(n530), .A2(n527), .A4(n531), .S0(n318), 
        .S1(n257), .Y(n525) );
  MUX41X1_HVT U88 ( .A1(n357), .A3(n342), .A2(n579), .A4(n563), .S0(n303), 
        .S1(n336), .Y(n523) );
  NAND2X0_HVT U89 ( .A1(n218), .A2(n227), .Y(n522) );
  MUX41X1_HVT U90 ( .A1(n272), .A3(n603), .A2(n562), .A4(n522), .S0(n303), 
        .S1(n334), .Y(n521) );
  MUX41X1_HVT U96 ( .A1(n382), .A3(n596), .A2(n365), .A4(n388), .S0(n304), 
        .S1(n281), .Y(n515) );
  MUX41X1_HVT U98 ( .A1(n514), .A3(n389), .A2(n373), .A4(n581), .S0(n304), 
        .S1(n282), .Y(n513) );
  MUX41X1_HVT U99 ( .A1(n577), .A3(n359), .A2(n561), .A4(n593), .S0(n282), 
        .S1(n301), .Y(n512) );
  NAND2X0_HVT U100 ( .A1(n291), .A2(n396), .Y(n511) );
  MUX41X1_HVT U101 ( .A1(n390), .A3(n597), .A2(n372), .A4(n511), .S0(n281), 
        .S1(n304), .Y(n510) );
  AND2X1_HVT U104 ( .A1(n603), .A2(n321), .Y(n508) );
  MUX41X1_HVT U107 ( .A1(n390), .A3(n324), .A2(n506), .A4(n348), .S0(n303), 
        .S1(n281), .Y(n505) );
  MUX41X1_HVT U108 ( .A1(n361), .A3(n319), .A2(n266), .A4(n326), .S0(n304), 
        .S1(n282), .Y(n504) );
  MUX41X1_HVT U109 ( .A1(n389), .A3(n342), .A2(n386), .A4(n379), .S0(n303), 
        .S1(n336), .Y(n503) );
  MUX41X1_HVT U110 ( .A1(n503), .A3(n505), .A2(n504), .A4(n507), .S0(in[5]), 
        .S1(n316), .Y(n502) );
  NAND2X0_HVT U114 ( .A1(n268), .A2(n603), .Y(n498) );
  MUX41X1_HVT U115 ( .A1(n498), .A3(n598), .A2(n375), .A4(n325), .S0(n281), 
        .S1(n301), .Y(n497) );
  MUX41X1_HVT U116 ( .A1(n374), .A3(n367), .A2(n342), .A4(n594), .S0(n302), 
        .S1(n336), .Y(n496) );
  NAND2X0_HVT U118 ( .A1(n239), .A2(n259), .Y(n494) );
  MUX41X1_HVT U119 ( .A1(n392), .A3(n495), .A2(n572), .A4(n494), .S0(n302), 
        .S1(n334), .Y(n493) );
  MUX41X1_HVT U122 ( .A1(n380), .A3(n293), .A2(n563), .A4(n384), .S0(n302), 
        .S1(n336), .Y(n491) );
  MUX41X1_HVT U124 ( .A1(n296), .A3(n490), .A2(n586), .A4(n290), .S0(n308), 
        .S1(n302), .Y(n489) );
  AOI21X1_HVT U127 ( .A1(n307), .A2(n485), .A3(n349), .Y(n486) );
  NAND2X0_HVT U129 ( .A1(n306), .A2(n268), .Y(n483) );
  MUX41X1_HVT U130 ( .A1(n483), .A3(n484), .A2(n487), .A4(n486), .S0(n310), 
        .S1(n316), .Y(n482) );
  AND2X1_HVT U131 ( .A1(n228), .A2(n291), .Y(n481) );
  MUX41X1_HVT U132 ( .A1(n346), .A3(n481), .A2(n394), .A4(n355), .S0(n309), 
        .S1(n300), .Y(n480) );
  MUX41X1_HVT U133 ( .A1(n395), .A3(n348), .A2(n555), .A4(n347), .S0(n308), 
        .S1(n300), .Y(n479) );
  MUX41X1_HVT U136 ( .A1(n560), .A3(n511), .A2(n477), .A4(n353), .S0(n306), 
        .S1(n282), .Y(n476) );
  MUX41X1_HVT U137 ( .A1(n602), .A3(n580), .A2(n243), .A4(n388), .S0(n310), 
        .S1(n304), .Y(n475) );
  MUX41X1_HVT U139 ( .A1(n474), .A3(n478), .A2(n482), .A4(n488), .S0(in[5]), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n370), .A3(n294), .A2(n364), .A4(n598), .S0(n309), 
        .S1(n301), .Y(n473) );
  NAND2X0_HVT U141 ( .A1(n319), .A2(n218), .Y(n472) );
  MUX41X1_HVT U142 ( .A1(n472), .A3(n570), .A2(n393), .A4(n364), .S0(n307), 
        .S1(n281), .Y(n471) );
  MUX41X1_HVT U143 ( .A1(n227), .A3(n376), .A2(n589), .A4(n586), .S0(n305), 
        .S1(n334), .Y(n470) );
  MUX41X1_HVT U145 ( .A1(n578), .A3(n391), .A2(n469), .A4(n529), .S0(n307), 
        .S1(n281), .Y(n468) );
  MUX41X1_HVT U146 ( .A1(n468), .A3(n470), .A2(n471), .A4(n473), .S0(in[1]), 
        .S1(n318), .Y(n467) );
  AO21X1_HVT U148 ( .A1(n310), .A2(n350), .A3(n396), .Y(n465) );
  MUX41X1_HVT U151 ( .A1(n258), .A3(n373), .A2(n362), .A4(n463), .S0(n308), 
        .S1(n300), .Y(n462) );
  MUX41X1_HVT U155 ( .A1(n364), .A3(n598), .A2(n590), .A4(n365), .S0(n305), 
        .S1(n282), .Y(n458) );
  MUX41X1_HVT U156 ( .A1(n458), .A3(n462), .A2(n459), .A4(n464), .S0(in[5]), 
        .S1(n316), .Y(n457) );
  NAND2X0_HVT U159 ( .A1(n454), .A2(n453), .Y(n455) );
  NAND2X0_HVT U163 ( .A1(n331), .A2(n397), .Y(n449) );
  NAND2X0_HVT U166 ( .A1(n599), .A2(n445), .Y(n446) );
  MUX41X1_HVT U170 ( .A1(n297), .A3(n295), .A2(n296), .A4(n442), .S0(n305), 
        .S1(n335), .Y(n441) );
  MUX41X1_HVT U172 ( .A1(n522), .A3(n440), .A2(n295), .A4(n587), .S0(n305), 
        .S1(n336), .Y(n439) );
  MUX41X1_HVT U173 ( .A1(n274), .A3(n271), .A2(n326), .A4(n573), .S0(n305), 
        .S1(n335), .Y(n438) );
  MUX41X1_HVT U174 ( .A1(n387), .A3(n555), .A2(n395), .A4(n208), .S0(n305), 
        .S1(n282), .Y(n437) );
  MUX41X1_HVT U175 ( .A1(n437), .A3(n438), .A2(n439), .A4(n441), .S0(n257), 
        .S1(n318), .Y(n436) );
  NAND2X0_HVT U177 ( .A1(n329), .A2(n259), .Y(n435) );
  AND2X1_HVT U179 ( .A1(n241), .A2(n321), .Y(n433) );
  MUX41X1_HVT U180 ( .A1(n577), .A3(n340), .A2(n433), .A4(n564), .S0(n305), 
        .S1(n335), .Y(n432) );
  MUX41X1_HVT U183 ( .A1(n376), .A3(n381), .A2(n361), .A4(n567), .S0(n308), 
        .S1(n300), .Y(n429) );
  AND2X1_HVT U185 ( .A1(n208), .A2(n218), .Y(n427) );
  NAND2X0_HVT U191 ( .A1(n338), .A2(n354), .Y(n421) );
  AND2X1_HVT U192 ( .A1(n371), .A2(n419), .Y(n420) );
  NAND2X0_HVT U194 ( .A1(n567), .A2(n419), .Y(n417) );
  NAND2X0_HVT U198 ( .A1(n280), .A2(n208), .Y(n599) );
  NAND2X0_HVT U200 ( .A1(n322), .A2(n229), .Y(n485) );
  NAND2X0_HVT U207 ( .A1(n291), .A2(n270), .Y(n549) );
  MUX21X2_HVT U2 ( .A1(n201), .A2(n400), .S0(n280), .Y(n573) );
  IBUFFX2_HVT U3 ( .A(n257), .Y(n233) );
  MUX41X1_HVT U14 ( .A1(n417), .A3(n418), .A2(n421), .A4(n420), .S0(n196), 
        .S1(n257), .Y(n416) );
  IBUFFX16_HVT U16 ( .A(n303), .Y(n196) );
  XOR2X2_HVT U17 ( .A1(n269), .A2(n250), .Y(n572) );
  MUX21X2_HVT U18 ( .A1(n555), .A2(n290), .S0(n197), .Y(n551) );
  IBUFFX16_HVT U20 ( .A(n309), .Y(n197) );
  MUX21X2_HVT U21 ( .A1(n568), .A2(n383), .S0(n339), .Y(n424) );
  IBUFFX2_HVT U22 ( .A(n339), .Y(n335) );
  XOR2X1_HVT U23 ( .A1(n314), .A2(in[3]), .Y(n593) );
  MUX41X1_HVT U24 ( .A1(n360), .A3(n377), .A2(n451), .A4(n574), .S0(n198), 
        .S1(n335), .Y(n450) );
  IBUFFX16_HVT U26 ( .A(n305), .Y(n198) );
  INVX0_HVT U27 ( .A(n268), .Y(n270) );
  INVX2_HVT U28 ( .A(n315), .Y(n257) );
  INVX0_HVT U29 ( .A(n315), .Y(n224) );
  IBUFFX2_HVT U30 ( .A(n315), .Y(n316) );
  NBUFFX2_HVT U31 ( .A(n401), .Y(n199) );
  AO21X1_HVT U33 ( .A1(n280), .A2(n396), .A3(n338), .Y(n419) );
  MUX21X2_HVT U34 ( .A1(n298), .A2(n584), .S0(n200), .Y(n461) );
  IBUFFX16_HVT U36 ( .A(n309), .Y(n200) );
  OA21X2_HVT U37 ( .A1(n343), .A2(n338), .A3(n352), .Y(n460) );
  NBUFFX2_HVT U39 ( .A(n401), .Y(n201) );
  OR2X2_HVT U40 ( .A1(n311), .A2(n199), .Y(n608) );
  NBUFFX2_HVT U41 ( .A(n199), .Y(n313) );
  INVX0_HVT U43 ( .A(n584), .Y(n364) );
  IBUFFX2_HVT U44 ( .A(n593), .Y(n400) );
  MUX21X2_HVT U45 ( .A1(n460), .A2(n461), .S0(n307), .Y(n459) );
  INVX2_HVT U46 ( .A(n588), .Y(n361) );
  MUX21X2_HVT U47 ( .A1(n320), .A2(n313), .S0(n279), .Y(n584) );
  MUX21X2_HVT U48 ( .A1(n319), .A2(n311), .S0(n331), .Y(n588) );
  INVX0_HVT U49 ( .A(n329), .Y(n229) );
  INVX0_HVT U50 ( .A(n279), .Y(n239) );
  IBUFFX2_HVT U51 ( .A(n573), .Y(n372) );
  MUX21X1_HVT U52 ( .A1(n201), .A2(n397), .S0(n280), .Y(n463) );
  INVX0_HVT U54 ( .A(n400), .Y(n202) );
  INVX1_HVT U56 ( .A(n202), .Y(n208) );
  NAND2X0_HVT U57 ( .A1(n324), .A2(n218), .Y(n219) );
  NAND2X0_HVT U58 ( .A1(n327), .A2(n329), .Y(n220) );
  NAND2X0_HVT U59 ( .A1(n219), .A2(n220), .Y(n591) );
  INVX0_HVT U61 ( .A(n329), .Y(n218) );
  NAND2X0_HVT U63 ( .A1(n532), .A2(n221), .Y(n222) );
  NAND2X0_HVT U64 ( .A1(n525), .A2(n225), .Y(n223) );
  NAND2X0_HVT U68 ( .A1(n222), .A2(n223), .Y(out[1]) );
  INVX0_HVT U69 ( .A(n225), .Y(n221) );
  INVX1_HVT U70 ( .A(n332), .Y(n329) );
  INVX0_HVT U71 ( .A(n591), .Y(n358) );
  INVX1_HVT U75 ( .A(n240), .Y(n225) );
  INVX0_HVT U76 ( .A(in[3]), .Y(n398) );
  MUX41X1_HVT U77 ( .A1(n444), .A3(n450), .A2(n448), .A4(n452), .S0(n318), 
        .S1(n224), .Y(n443) );
  INVX1_HVT U86 ( .A(n332), .Y(n330) );
  MUX21X2_HVT U87 ( .A1(n535), .A2(n534), .S0(n307), .Y(n533) );
  MUX21X2_HVT U91 ( .A1(n321), .A2(n325), .S0(n331), .Y(n451) );
  INVX1_HVT U92 ( .A(n332), .Y(n280) );
  INVX1_HVT U93 ( .A(n273), .Y(n268) );
  INVX1_HVT U94 ( .A(n235), .Y(n442) );
  INVX0_HVT U95 ( .A(n397), .Y(n226) );
  INVX1_HVT U97 ( .A(n226), .Y(n227) );
  NBUFFX2_HVT U102 ( .A(n292), .Y(n228) );
  MUX21X1_HVT U103 ( .A1(n397), .A2(n399), .S0(n229), .Y(n495) );
  NAND2X0_HVT U105 ( .A1(n492), .A2(n230), .Y(n231) );
  NAND2X0_HVT U106 ( .A1(n502), .A2(in[7]), .Y(n232) );
  NAND2X0_HVT U111 ( .A1(n231), .A2(n232), .Y(out[3]) );
  IBUFFX2_HVT U112 ( .A(in[7]), .Y(n230) );
  INVX0_HVT U113 ( .A(n605), .Y(n397) );
  IBUFFX2_HVT U117 ( .A(n401), .Y(n292) );
  MUX41X1_HVT U120 ( .A1(n426), .A3(n423), .A2(n425), .A4(n424), .S0(n233), 
        .S1(n234), .Y(n422) );
  IBUFFX16_HVT U121 ( .A(n300), .Y(n234) );
  MUX21X1_HVT U123 ( .A1(n268), .A2(n323), .S0(n249), .Y(n235) );
  NAND2X0_HVT U125 ( .A1(n327), .A2(n236), .Y(n237) );
  NAND2X0_HVT U126 ( .A1(n321), .A2(n239), .Y(n238) );
  NAND2X0_HVT U128 ( .A1(n237), .A2(n238), .Y(n403) );
  INVX0_HVT U134 ( .A(n239), .Y(n236) );
  INVX0_HVT U135 ( .A(n403), .Y(n394) );
  IBUFFX16_HVT U138 ( .A(n263), .Y(n240) );
  MUX21X2_HVT U144 ( .A1(n298), .A2(n561), .S0(n310), .Y(n425) );
  MUX21X2_HVT U147 ( .A1(n394), .A2(n346), .S0(n308), .Y(n466) );
  MUX21X2_HVT U149 ( .A1(n457), .A2(n467), .S0(in[7]), .Y(out[5]) );
  MUX21X1_HVT U150 ( .A1(n362), .A2(n607), .S0(n306), .Y(n546) );
  INVX0_HVT U152 ( .A(n332), .Y(n331) );
  INVX1_HVT U153 ( .A(n347), .Y(n241) );
  INVX0_HVT U154 ( .A(n584), .Y(n242) );
  INVX1_HVT U157 ( .A(n242), .Y(n243) );
  NAND2X0_HVT U158 ( .A1(n429), .A2(n244), .Y(n245) );
  NAND2X0_HVT U160 ( .A1(n430), .A2(n257), .Y(n246) );
  NAND2X0_HVT U161 ( .A1(n245), .A2(n246), .Y(n428) );
  IBUFFX2_HVT U162 ( .A(n257), .Y(n244) );
  MUX41X1_HVT U164 ( .A1(n270), .A3(n241), .A2(n351), .A4(n598), .S0(n247), 
        .S1(n336), .Y(n539) );
  IBUFFX16_HVT U165 ( .A(n303), .Y(n247) );
  INVX1_HVT U167 ( .A(n339), .Y(n337) );
  INVX1_HVT U168 ( .A(n610), .Y(n273) );
  INVX1_HVT U169 ( .A(n415), .Y(n381) );
  MUX21X2_HVT U171 ( .A1(n557), .A2(n558), .S0(n248), .Y(n556) );
  IBUFFX16_HVT U176 ( .A(n306), .Y(n248) );
  INVX1_HVT U178 ( .A(in[0]), .Y(n332) );
  MUX41X1_HVT U181 ( .A1(n497), .A3(n493), .A2(n499), .A4(n496), .S0(n317), 
        .S1(n316), .Y(n492) );
  AO21X2_HVT U182 ( .A1(n375), .A2(n309), .A3(n585), .Y(n500) );
  MUX21X2_HVT U184 ( .A1(n349), .A2(n568), .S0(n310), .Y(n501) );
  NBUFFX16_HVT U186 ( .A(n337), .Y(n310) );
  OA21X1_HVT U187 ( .A1(n367), .A2(n338), .A3(n549), .Y(n423) );
  NBUFFX2_HVT U188 ( .A(n279), .Y(n249) );
  NBUFFX2_HVT U189 ( .A(n279), .Y(n250) );
  NBUFFX2_HVT U190 ( .A(n279), .Y(n251) );
  IBUFFX2_HVT U193 ( .A(n332), .Y(n328) );
  MUX21X2_HVT U195 ( .A1(n365), .A2(n356), .S0(n310), .Y(n558) );
  INVX0_HVT U196 ( .A(n266), .Y(n583) );
  MUX41X1_HVT U197 ( .A1(n345), .A3(n298), .A2(n387), .A4(n266), .S0(n302), 
        .S1(n334), .Y(n524) );
  MUX21X1_HVT U199 ( .A1(n446), .A2(n447), .S0(n306), .Y(n444) );
  INVX0_HVT U201 ( .A(n566), .Y(n376) );
  INVX1_HVT U202 ( .A(n278), .Y(n568) );
  INVX1_HVT U203 ( .A(n339), .Y(n336) );
  INVX0_HVT U204 ( .A(n275), .Y(n559) );
  INVX1_HVT U205 ( .A(in[4]), .Y(n338) );
  INVX0_HVT U206 ( .A(n201), .Y(n267) );
  INVX1_HVT U208 ( .A(in[4]), .Y(n339) );
  NBUFFX2_HVT U209 ( .A(n401), .Y(n314) );
  INVX1_HVT U210 ( .A(in[1]), .Y(n315) );
  INVX1_HVT U211 ( .A(n398), .Y(n259) );
  INVX1_HVT U212 ( .A(in[7]), .Y(n263) );
  INVX1_HVT U213 ( .A(in[5]), .Y(n317) );
  INVX1_HVT U214 ( .A(n335), .Y(n256) );
  INVX1_HVT U215 ( .A(n306), .Y(n262) );
  MUX21X2_HVT U216 ( .A1(n500), .A2(n501), .S0(n307), .Y(n499) );
  NAND2X0_HVT U217 ( .A1(n455), .A2(n262), .Y(n252) );
  NAND2X0_HVT U218 ( .A1(n456), .A2(n307), .Y(n253) );
  NAND2X0_HVT U219 ( .A1(n252), .A2(n253), .Y(n452) );
  NAND2X0_HVT U220 ( .A1(n443), .A2(in[7]), .Y(n254) );
  NAND2X0_HVT U221 ( .A1(n436), .A2(n263), .Y(n255) );
  NAND2X0_HVT U222 ( .A1(n254), .A2(n255), .Y(out[6]) );
  MUX21X1_HVT U223 ( .A1(n566), .A2(n384), .S0(n309), .Y(n456) );
  MUX41X1_HVT U224 ( .A1(n572), .A3(n361), .A2(n601), .A4(n449), .S0(n302), 
        .S1(n256), .Y(n448) );
  OA21X1_HVT U225 ( .A1(n344), .A2(n338), .A3(n588), .Y(n534) );
  XOR2X2_HVT U226 ( .A1(n321), .A2(n249), .Y(n561) );
  MUX21X1_HVT U227 ( .A1(n259), .A2(n593), .S0(n330), .Y(n258) );
  NAND2X0_HVT U228 ( .A1(n324), .A2(n283), .Y(n260) );
  NAND2X0_HVT U229 ( .A1(n520), .A2(n291), .Y(n261) );
  NAND2X0_HVT U230 ( .A1(n260), .A2(n261), .Y(n519) );
  MUX21X2_HVT U231 ( .A1(n519), .A2(n518), .S0(n262), .Y(n517) );
  NAND2X2_HVT U232 ( .A1(n509), .A2(n263), .Y(n264) );
  NAND2X0_HVT U233 ( .A1(n516), .A2(in[7]), .Y(n265) );
  NAND2X0_HVT U234 ( .A1(n264), .A2(n265), .Y(out[2]) );
  MUX21X1_HVT U235 ( .A1(n311), .A2(n399), .S0(n328), .Y(n566) );
  MUX21X1_HVT U236 ( .A1(n267), .A2(n327), .S0(n328), .Y(n266) );
  INVX1_HVT U237 ( .A(n412), .Y(n384) );
  MUX41X1_HVT U238 ( .A1(n517), .A3(n521), .A2(n523), .A4(n524), .S0(n316), 
        .S1(n318), .Y(n516) );
  INVX1_HVT U239 ( .A(n273), .Y(n269) );
  INVX1_HVT U240 ( .A(n269), .Y(n271) );
  INVX1_HVT U241 ( .A(n269), .Y(n272) );
  INVX1_HVT U242 ( .A(n273), .Y(n274) );
  MUX21X1_HVT U243 ( .A1(n326), .A2(n324), .S0(n329), .Y(n275) );
  INVX1_HVT U244 ( .A(n326), .Y(n396) );
  INVX1_HVT U245 ( .A(n332), .Y(n279) );
  NAND2X0_HVT U246 ( .A1(n586), .A2(n282), .Y(n276) );
  NAND2X0_HVT U247 ( .A1(n583), .A2(n256), .Y(n277) );
  NAND2X0_HVT U248 ( .A1(n276), .A2(n277), .Y(n447) );
  MUX21X1_HVT U249 ( .A1(n323), .A2(n199), .S0(n332), .Y(n278) );
  INVX1_HVT U250 ( .A(n323), .Y(n399) );
  INVX1_HVT U251 ( .A(in[6]), .Y(n401) );
  NBUFFX2_HVT U252 ( .A(n398), .Y(n312) );
  INVX0_HVT U253 ( .A(n356), .Y(n289) );
  INVX0_HVT U254 ( .A(n595), .Y(n355) );
  AO21X1_HVT U255 ( .A1(n320), .A2(n607), .A3(n338), .Y(n445) );
  MUX21X1_HVT U256 ( .A1(n397), .A2(n272), .S0(n251), .Y(n565) );
  MUX21X1_HVT U257 ( .A1(n489), .A2(n491), .S0(n316), .Y(n488) );
  INVX0_HVT U258 ( .A(n565), .Y(n377) );
  INVX1_HVT U259 ( .A(n339), .Y(n281) );
  INVX1_HVT U260 ( .A(n339), .Y(n282) );
  MUX41X1_HVT U261 ( .A1(n508), .A3(n529), .A2(n391), .A4(n595), .S0(n262), 
        .S1(n256), .Y(n507) );
  INVX1_HVT U262 ( .A(n339), .Y(n334) );
  MUX41X1_HVT U263 ( .A1(n515), .A3(n512), .A2(n513), .A4(n510), .S0(n317), 
        .S1(n315), .Y(n509) );
  INVX1_HVT U264 ( .A(n582), .Y(n365) );
  NAND2X0_HVT U265 ( .A1(n398), .A2(n283), .Y(n284) );
  NAND2X0_HVT U266 ( .A1(n326), .A2(n291), .Y(n285) );
  NAND2X0_HVT U267 ( .A1(n284), .A2(n285), .Y(n290) );
  INVX0_HVT U268 ( .A(n291), .Y(n283) );
  MUX41X1_HVT U269 ( .A1(n555), .A3(n266), .A2(n593), .A4(n381), .S0(n262), 
        .S1(n338), .Y(n554) );
  INVX0_HVT U270 ( .A(n290), .Y(n586) );
  INVX1_HVT U271 ( .A(n288), .Y(n541) );
  MUX41X1_HVT U272 ( .A1(n348), .A3(n345), .A2(n607), .A4(n258), .S0(n334), 
        .S1(n302), .Y(n430) );
  MUX41X1_HVT U273 ( .A1(n431), .A3(n422), .A2(n428), .A4(n416), .S0(n263), 
        .S1(n317), .Y(out[7]) );
  INVX0_HVT U274 ( .A(n279), .Y(n291) );
  AO21X2_HVT U275 ( .A1(n239), .A2(n274), .A3(n338), .Y(n453) );
  NAND2X0_HVT U276 ( .A1(n432), .A2(n315), .Y(n286) );
  NAND2X0_HVT U277 ( .A1(n434), .A2(n316), .Y(n287) );
  NAND2X0_HVT U278 ( .A1(n286), .A2(n287), .Y(n431) );
  MUX41X1_HVT U279 ( .A1(n272), .A3(n289), .A2(n398), .A4(n595), .S0(n262), 
        .S1(n338), .Y(n288) );
  MUX21X2_HVT U280 ( .A1(n547), .A2(n540), .S0(n263), .Y(out[0]) );
  NBUFFX2_HVT U281 ( .A(n593), .Y(n319) );
  MUX41X1_HVT U282 ( .A1(n545), .A3(n542), .A2(n544), .A4(n541), .S0(n317), 
        .S1(n315), .Y(n540) );
  INVX2_HVT U283 ( .A(n317), .Y(n318) );
  MUX21X2_HVT U284 ( .A1(n361), .A2(n546), .S0(n299), .Y(n545) );
  INVX1_HVT U285 ( .A(n587), .Y(n362) );
  MUX41X1_HVT U286 ( .A1(n565), .A3(n271), .A2(n435), .A4(n297), .S0(n262), 
        .S1(n256), .Y(n434) );
  INVX1_HVT U287 ( .A(n413), .Y(n383) );
  MUX21X1_HVT U288 ( .A1(n384), .A2(n341), .S0(n310), .Y(n535) );
  MUX21X2_HVT U289 ( .A1(n551), .A2(n550), .S0(n306), .Y(n548) );
  NBUFFX2_HVT U290 ( .A(n609), .Y(n326) );
  NBUFFX2_HVT U291 ( .A(n609), .Y(n327) );
  AND2X1_HVT U292 ( .A1(n327), .A2(n594), .Y(n293) );
  MUX21X1_HVT U293 ( .A1(n378), .A2(n296), .S0(n308), .Y(n418) );
  MUX21X1_HVT U294 ( .A1(n400), .A2(n396), .S0(n330), .Y(n587) );
  MUX21X1_HVT U295 ( .A1(n396), .A2(n400), .S0(n328), .Y(n576) );
  MUX21X1_HVT U296 ( .A1(n319), .A2(n272), .S0(n328), .Y(n578) );
  MUX21X1_HVT U297 ( .A1(n271), .A2(n313), .S0(n251), .Y(n440) );
  NAND2X0_HVT U298 ( .A1(n398), .A2(n314), .Y(n609) );
  MUX21X1_HVT U299 ( .A1(n272), .A2(n320), .S0(n328), .Y(n409) );
  MUX21X1_HVT U300 ( .A1(n396), .A2(n313), .S0(n280), .Y(n413) );
  MUX21X1_HVT U301 ( .A1(n270), .A2(n397), .S0(n250), .Y(n581) );
  MUX21X1_HVT U302 ( .A1(n400), .A2(n312), .S0(n329), .Y(n570) );
  MUX21X1_HVT U303 ( .A1(n312), .A2(n396), .S0(n251), .Y(n579) );
  MUX21X1_HVT U304 ( .A1(n208), .A2(n313), .S0(n250), .Y(n404) );
  MUX21X1_HVT U305 ( .A1(n466), .A2(n465), .S0(n306), .Y(n464) );
  MUX21X1_HVT U306 ( .A1(n201), .A2(n327), .S0(n250), .Y(n506) );
  MUX21X1_HVT U307 ( .A1(n393), .A2(n294), .S0(n306), .Y(n487) );
  MUX21X1_HVT U308 ( .A1(n351), .A2(n319), .S0(n310), .Y(n518) );
  MUX21X1_HVT U309 ( .A1(n319), .A2(n201), .S0(n309), .Y(n520) );
  XOR2X1_HVT U310 ( .A1(n319), .A2(n250), .Y(n563) );
  MUX21X1_HVT U311 ( .A1(n399), .A2(n311), .S0(n251), .Y(n412) );
  MUX21X1_HVT U312 ( .A1(n320), .A2(n397), .S0(n331), .Y(n575) );
  MUX21X1_HVT U313 ( .A1(n201), .A2(n320), .S0(n331), .Y(n569) );
  MUX21X1_HVT U314 ( .A1(n311), .A2(n327), .S0(n280), .Y(n411) );
  XNOR2X1_HVT U315 ( .A1(n326), .A2(n330), .Y(n294) );
  MUX21X1_HVT U316 ( .A1(n274), .A2(n327), .S0(n279), .Y(n595) );
  MUX21X1_HVT U317 ( .A1(n576), .A2(n293), .S0(n307), .Y(n484) );
  XOR2X1_HVT U318 ( .A1(n324), .A2(n330), .Y(n562) );
  AND2X1_HVT U319 ( .A1(n604), .A2(n327), .Y(n295) );
  MUX21X1_HVT U320 ( .A1(n312), .A2(n313), .S0(n329), .Y(n564) );
  MUX21X1_HVT U321 ( .A1(n324), .A2(n312), .S0(n280), .Y(n590) );
  MUX21X1_HVT U322 ( .A1(n312), .A2(n324), .S0(n328), .Y(n406) );
  AND2X1_HVT U323 ( .A1(n330), .A2(n313), .Y(n296) );
  MUX21X1_HVT U324 ( .A1(n325), .A2(n201), .S0(n330), .Y(n490) );
  NBUFFX2_HVT U325 ( .A(n337), .Y(n309) );
  NBUFFX2_HVT U326 ( .A(n337), .Y(n308) );
  MUX21X1_HVT U327 ( .A1(n427), .A2(n385), .S0(n308), .Y(n426) );
  MUX21X1_HVT U328 ( .A1(n326), .A2(n322), .S0(n280), .Y(n469) );
  NBUFFX2_HVT U329 ( .A(n593), .Y(n320) );
  MUX21X1_HVT U330 ( .A1(n363), .A2(n553), .S0(n299), .Y(n552) );
  MUX21X1_HVT U331 ( .A1(n364), .A2(n606), .S0(n307), .Y(n553) );
  AND2X1_HVT U332 ( .A1(n399), .A2(n218), .Y(n297) );
  NBUFFX2_HVT U333 ( .A(n605), .Y(n321) );
  NBUFFX2_HVT U334 ( .A(n608), .Y(n323) );
  AND2X1_HVT U335 ( .A1(n325), .A2(n291), .Y(n298) );
  NBUFFX2_HVT U336 ( .A(n608), .Y(n325) );
  NBUFFX2_HVT U337 ( .A(n605), .Y(n322) );
  NBUFFX2_HVT U338 ( .A(n608), .Y(n324) );
  NBUFFX2_HVT U339 ( .A(n398), .Y(n311) );
  NBUFFX2_HVT U340 ( .A(n301), .Y(n305) );
  NBUFFX2_HVT U341 ( .A(n333), .Y(n307) );
  NBUFFX2_HVT U342 ( .A(in[2]), .Y(n306) );
  XNOR2X1_HVT U343 ( .A1(n338), .A2(n302), .Y(n299) );
  NBUFFX2_HVT U344 ( .A(n333), .Y(n302) );
  NBUFFX2_HVT U345 ( .A(n333), .Y(n304) );
  NBUFFX2_HVT U346 ( .A(n333), .Y(n303) );
  NBUFFX2_HVT U347 ( .A(n333), .Y(n300) );
  NBUFFX2_HVT U348 ( .A(n333), .Y(n301) );
  MUX21X1_HVT U349 ( .A1(n272), .A2(n259), .S0(n329), .Y(n402) );
  MUX21X1_HVT U350 ( .A1(n292), .A2(n271), .S0(n330), .Y(n585) );
  MUX21X1_HVT U351 ( .A1(n269), .A2(n259), .S0(n331), .Y(n454) );
  MUX21X1_HVT U352 ( .A1(n322), .A2(n259), .S0(n250), .Y(n514) );
  MUX21X1_HVT U353 ( .A1(n479), .A2(n480), .S0(n316), .Y(n478) );
  MUX21X1_HVT U354 ( .A1(n475), .A2(n476), .S0(in[1]), .Y(n474) );
  XOR2X1_HVT U355 ( .A1(n280), .A2(n228), .Y(n560) );
  MUX21X1_HVT U356 ( .A1(n396), .A2(n228), .S0(n329), .Y(n477) );
  MUX21X1_HVT U357 ( .A1(n292), .A2(n397), .S0(n331), .Y(n415) );
  MUX21X1_HVT U358 ( .A1(n322), .A2(n292), .S0(n331), .Y(n580) );
  MUX21X1_HVT U359 ( .A1(n313), .A2(n259), .S0(n249), .Y(n582) );
  MUX21X1_HVT U360 ( .A1(n259), .A2(n274), .S0(n331), .Y(n408) );
  MUX21X1_HVT U361 ( .A1(n259), .A2(n322), .S0(n249), .Y(n407) );
  MUX21X1_HVT U362 ( .A1(n228), .A2(n325), .S0(n251), .Y(n414) );
  MUX21X1_HVT U363 ( .A1(n325), .A2(n228), .S0(n283), .Y(n410) );
  MUX21X1_HVT U364 ( .A1(n312), .A2(n292), .S0(n330), .Y(n405) );
  NBUFFX2_HVT U365 ( .A(in[2]), .Y(n333) );
  MUX21X1_HVT U366 ( .A1(n292), .A2(n268), .S0(n328), .Y(n592) );
  INVX0_HVT U367 ( .A(n598), .Y(n340) );
  INVX0_HVT U368 ( .A(n577), .Y(n341) );
  INVX0_HVT U369 ( .A(n571), .Y(n342) );
  INVX0_HVT U370 ( .A(n511), .Y(n343) );
  INVX0_HVT U371 ( .A(n472), .Y(n344) );
  INVX0_HVT U372 ( .A(n607), .Y(n345) );
  INVX0_HVT U373 ( .A(n606), .Y(n346) );
  INVX0_HVT U374 ( .A(n604), .Y(n347) );
  INVX0_HVT U375 ( .A(n567), .Y(n348) );
  INVX0_HVT U376 ( .A(n603), .Y(n349) );
  INVX0_HVT U377 ( .A(n602), .Y(n350) );
  INVX0_HVT U378 ( .A(n574), .Y(n351) );
  INVX0_HVT U379 ( .A(n596), .Y(n352) );
  INVX0_HVT U380 ( .A(n601), .Y(n353) );
  INVX0_HVT U381 ( .A(n597), .Y(n354) );
  INVX0_HVT U382 ( .A(n594), .Y(n356) );
  INVX0_HVT U383 ( .A(n592), .Y(n357) );
  INVX0_HVT U384 ( .A(n590), .Y(n359) );
  INVX0_HVT U385 ( .A(n589), .Y(n360) );
  INVX0_HVT U386 ( .A(n585), .Y(n363) );
  INVX0_HVT U387 ( .A(n581), .Y(n366) );
  INVX0_HVT U388 ( .A(n580), .Y(n367) );
  INVX0_HVT U389 ( .A(n579), .Y(n368) );
  INVX0_HVT U390 ( .A(n578), .Y(n369) );
  INVX0_HVT U391 ( .A(n576), .Y(n370) );
  INVX0_HVT U392 ( .A(n575), .Y(n371) );
  INVX0_HVT U393 ( .A(n572), .Y(n373) );
  INVX0_HVT U394 ( .A(n570), .Y(n374) );
  INVX0_HVT U395 ( .A(n569), .Y(n375) );
  INVX0_HVT U396 ( .A(n564), .Y(n378) );
  INVX0_HVT U397 ( .A(n563), .Y(n379) );
  INVX0_HVT U398 ( .A(n600), .Y(n380) );
  INVX0_HVT U399 ( .A(n414), .Y(n382) );
  INVX0_HVT U400 ( .A(n411), .Y(n385) );
  INVX0_HVT U401 ( .A(n410), .Y(n386) );
  INVX0_HVT U402 ( .A(n409), .Y(n387) );
  INVX0_HVT U403 ( .A(n408), .Y(n388) );
  INVX0_HVT U404 ( .A(n407), .Y(n389) );
  INVX0_HVT U405 ( .A(n406), .Y(n390) );
  INVX0_HVT U406 ( .A(n405), .Y(n391) );
  INVX0_HVT U407 ( .A(n454), .Y(n392) );
  INVX0_HVT U408 ( .A(n404), .Y(n393) );
  INVX0_HVT U409 ( .A(n402), .Y(n395) );
endmodule

