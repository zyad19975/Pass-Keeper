
module sbox_0 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n119, n120, n121, n122, n123, n124, n125, n126, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n214, n215, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n233, n234, n235, n237, n239, n240,
         n241, n242, n244, n245, n246, n247, n248, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n260, n262, n263, n265, n266, n267,
         n268, n272, n274, n275, n276, n277, n278, n279, n281, n284, n285,
         n286, n287, n288, n290, n291, n292, n294, n295, n296, n298, n299,
         n300, n301, n302, n12, n18, n19, n23, n50, n78, n118, n127, n210,
         n211, n212, n213, n216, n217, n218, n219, n231, n232, n236, n238,
         n243, n249, n259, n261, n264, n269, n270, n271, n273, n280, n282,
         n283, n289, n293, n297, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472;

  NAND2X0_HVT U4 ( .A1(n448), .A2(n3), .Y(n4) );
  NAND2X0_HVT U5 ( .A1(n364), .A2(n442), .Y(n6) );
  NAND2X0_HVT U15 ( .A1(n3), .A2(n389), .Y(n16) );
  NAND2X0_HVT U21 ( .A1(n448), .A2(n461), .Y(n22) );
  NAND2X0_HVT U24 ( .A1(n436), .A2(n461), .Y(n25) );
  NAND2X0_HVT U33 ( .A1(n266), .A2(n461), .Y(n34) );
  NAND2X0_HVT U42 ( .A1(n457), .A2(n436), .Y(n43) );
  MUX41X1_HVT U51 ( .A1(n294), .A3(n260), .A2(n301), .A4(n291), .S0(n469), 
        .S1(n431), .Y(n52) );
  NAND2X0_HVT U56 ( .A1(n448), .A2(n59), .Y(n58) );
  NAND2X0_HVT U58 ( .A1(n454), .A2(n3), .Y(n61) );
  NAND2X0_HVT U62 ( .A1(n461), .A2(n450), .Y(n65) );
  AO21X1_HVT U66 ( .A1(n242), .A2(n466), .A3(n239), .Y(n69) );
  MUX41X1_HVT U68 ( .A1(n286), .A3(n69), .A2(n70), .A4(n68), .S0(n427), .S1(
        n470), .Y(n71) );
  NAND2X0_HVT U73 ( .A1(n446), .A2(n76), .Y(n75) );
  MUX41X1_HVT U74 ( .A1(n74), .A3(n27), .A2(n75), .A4(n25), .S0(n463), .S1(
        n470), .Y(n77) );
  MUX41X1_HVT U77 ( .A1(n9), .A3(n265), .A2(n79), .A4(n278), .S0(n432), .S1(
        n425), .Y(n80) );
  AND2X1_HVT U83 ( .A1(n457), .A2(n439), .Y(n87) );
  NAND2X0_HVT U85 ( .A1(n461), .A2(n346), .Y(n89) );
  MUX41X1_HVT U86 ( .A1(n247), .A3(n89), .A2(n418), .A4(n417), .S0(n427), .S1(
        n468), .Y(n90) );
  MUX41X1_HVT U96 ( .A1(n233), .A3(n420), .A2(n245), .A4(n99), .S0(n427), .S1(
        n382), .Y(n100) );
  MUX41X1_HVT U97 ( .A1(n244), .A3(n420), .A2(n402), .A4(n16), .S0(n427), .S1(
        n413), .Y(n101) );
  NAND2X0_HVT U101 ( .A1(n106), .A2(n107), .Y(n105) );
  MUX41X1_HVT U103 ( .A1(n3), .A3(n258), .A2(n272), .A4(n36), .S0(n427), .S1(
        n382), .Y(n109) );
  MUX41X1_HVT U105 ( .A1(n250), .A3(n49), .A2(n110), .A4(n262), .S0(n427), 
        .S1(n413), .Y(n111) );
  NAND2X0_HVT U110 ( .A1(n450), .A2(n116), .Y(n115) );
  AND2X1_HVT U115 ( .A1(n356), .A2(n392), .Y(n121) );
  MUX41X1_HVT U135 ( .A1(n279), .A3(n246), .A2(n6), .A4(n28), .S0(n428), .S1(
        n468), .Y(n142) );
  AND2X1_HVT U140 ( .A1(n330), .A2(n347), .Y(n147) );
  MUX41X1_HVT U141 ( .A1(n26), .A3(n339), .A2(n147), .A4(n212), .S0(n213), 
        .S1(n469), .Y(n148) );
  MUX41X1_HVT U142 ( .A1(n284), .A3(n390), .A2(n263), .A4(n445), .S0(n213), 
        .S1(n470), .Y(n149) );
  NAND2X0_HVT U146 ( .A1(n457), .A2(n455), .Y(n76) );
  MUX41X1_HVT U147 ( .A1(n295), .A3(n76), .A2(n244), .A4(n47), .S0(n315), .S1(
        n468), .Y(n153) );
  MUX41X1_HVT U153 ( .A1(n115), .A3(n415), .A2(n450), .A4(n256), .S0(n238), 
        .S1(n382), .Y(n159) );
  AND2X1_HVT U154 ( .A1(n434), .A2(n436), .Y(n160) );
  NAND2X0_HVT U158 ( .A1(n401), .A2(n346), .Y(n164) );
  MUX41X1_HVT U159 ( .A1(n365), .A3(n391), .A2(n164), .A4(n237), .S0(n426), 
        .S1(n413), .Y(n165) );
  AND2X1_HVT U162 ( .A1(n386), .A2(n76), .Y(n168) );
  MUX41X1_HVT U163 ( .A1(n320), .A3(n168), .A2(n419), .A4(n167), .S0(n426), 
        .S1(n413), .Y(n169) );
  NAND2X0_HVT U166 ( .A1(n454), .A2(n59), .Y(n172) );
  NAND2X0_HVT U167 ( .A1(n296), .A2(n461), .Y(n173) );
  MUX41X1_HVT U168 ( .A1(n277), .A3(n445), .A2(n173), .A4(n172), .S0(n426), 
        .S1(n469), .Y(n174) );
  NAND2X0_HVT U174 ( .A1(n23), .A2(n385), .Y(n14) );
  MUX41X1_HVT U176 ( .A1(n440), .A3(n179), .A2(n281), .A4(n14), .S0(n382), 
        .S1(n425), .Y(n180) );
  NAND2X0_HVT U177 ( .A1(n355), .A2(n441), .Y(n181) );
  MUX41X1_HVT U180 ( .A1(n287), .A3(n9), .A2(n365), .A4(n416), .S0(n432), .S1(
        n426), .Y(n184) );
  MUX41X1_HVT U189 ( .A1(n192), .A3(n14), .A2(n191), .A4(n262), .S0(n432), 
        .S1(n425), .Y(n193) );
  AO21X1_HVT U197 ( .A1(n418), .A2(n433), .A3(n248), .Y(n200) );
  MUX41X1_HVT U203 ( .A1(n37), .A3(n299), .A2(n309), .A4(n33), .S0(n426), .S1(
        n469), .Y(n206) );
  NAND2X0_HVT U208 ( .A1(n356), .A2(n449), .Y(n116) );
  NAND2X0_HVT U212 ( .A1(n393), .A2(n445), .Y(n59) );
  NAND2X0_HVT U214 ( .A1(n386), .A2(n461), .Y(n214) );
  NAND2X0_HVT U215 ( .A1(n116), .A2(n446), .Y(n215) );
  NAND2X0_HVT U218 ( .A1(n246), .A2(n457), .Y(n157) );
  NAND2X0_HVT U220 ( .A1(n433), .A2(n214), .Y(n84) );
  INVX0_HVT U241 ( .A(n25), .Y(n233) );
  INVX0_HVT U242 ( .A(n43), .Y(n234) );
  INVX0_HVT U245 ( .A(n6), .Y(n237) );
  INVX0_HVT U247 ( .A(n76), .Y(n239) );
  INVX0_HVT U256 ( .A(n157), .Y(n248) );
  INVX0_HVT U265 ( .A(n27), .Y(n257) );
  INVX0_HVT U268 ( .A(n22), .Y(n260) );
  INVX0_HVT U270 ( .A(n215), .Y(n262) );
  INVX0_HVT U283 ( .A(n13), .Y(n275) );
  INVX0_HVT U284 ( .A(n214), .Y(n276) );
  INVX0_HVT U289 ( .A(n107), .Y(n281) );
  INVX0_HVT U295 ( .A(n4), .Y(n287) );
  INVX0_HVT U296 ( .A(n16), .Y(n288) );
  INVX0_HVT U300 ( .A(n42), .Y(n292) );
  INVX0_HVT U302 ( .A(n220), .Y(n294) );
  INVX0_HVT U303 ( .A(n228), .Y(n295) );
  INVX0_HVT U306 ( .A(n173), .Y(n298) );
  INVX0_HVT U309 ( .A(n20), .Y(n301) );
  MUX21X1_HVT U1 ( .A1(n442), .A2(n439), .S0(n23), .Y(n31) );
  INVX0_HVT U2 ( .A(n465), .Y(n464) );
  INVX1_HVT U3 ( .A(n434), .Y(n303) );
  MUX21X1_HVT U6 ( .A1(n392), .A2(n442), .S0(n23), .Y(n17) );
  MUX21X1_HVT U7 ( .A1(n445), .A2(n21), .S0(n303), .Y(n82) );
  MUX21X1_HVT U8 ( .A1(n443), .A2(n350), .S0(n456), .Y(n41) );
  OA21X1_HVT U9 ( .A1(n422), .A2(n472), .A3(n32), .Y(n176) );
  INVX1_HVT U10 ( .A(n31), .Y(n251) );
  INVX1_HVT U11 ( .A(n387), .Y(n389) );
  INVX1_HVT U12 ( .A(n444), .Y(n246) );
  MUX21X1_HVT U13 ( .A1(n234), .A2(n253), .S0(n433), .Y(n199) );
  INVX1_HVT U14 ( .A(n212), .Y(n33) );
  INVX1_HVT U16 ( .A(n444), .Y(n406) );
  MUX21X1_HVT U17 ( .A1(n439), .A2(n346), .S0(n402), .Y(n37) );
  MUX21X1_HVT U18 ( .A1(n296), .A2(n312), .S0(n351), .Y(n349) );
  XOR2X1_HVT U19 ( .A1(n23), .A2(n424), .Y(n351) );
  AND3X1_HVT U20 ( .A1(n428), .A2(n461), .A3(n439), .Y(n136) );
  MUX21X1_HVT U22 ( .A1(n328), .A2(n212), .S0(n463), .Y(n138) );
  MUX21X1_HVT U23 ( .A1(n250), .A2(n31), .S0(n463), .Y(n135) );
  AO21X1_HVT U25 ( .A1(n434), .A2(n97), .A3(n248), .Y(n96) );
  INVX1_HVT U26 ( .A(n127), .Y(n3) );
  INVX1_HVT U27 ( .A(n30), .Y(n272) );
  INVX1_HVT U28 ( .A(n15), .Y(n290) );
  MUX21X1_HVT U29 ( .A1(n151), .A2(n150), .S0(n321), .Y(n152) );
  MUX21X1_HVT U30 ( .A1(n83), .A2(n82), .S0(n341), .Y(n85) );
  INVX1_HVT U31 ( .A(n431), .Y(n12) );
  INVX1_HVT U32 ( .A(n431), .Y(n231) );
  INVX1_HVT U34 ( .A(in[7]), .Y(n471) );
  INVX0_HVT U35 ( .A(n471), .Y(n413) );
  INVX0_HVT U36 ( .A(n471), .Y(n382) );
  INVX1_HVT U37 ( .A(n471), .Y(n470) );
  INVX1_HVT U38 ( .A(n471), .Y(n469) );
  MUX21X1_HVT U39 ( .A1(n31), .A2(n215), .S0(n432), .Y(n225) );
  MUX21X1_HVT U40 ( .A1(n415), .A2(n103), .S0(n48), .Y(n104) );
  NBUFFX2_HVT U41 ( .A(in[4]), .Y(n438) );
  INVX0_HVT U43 ( .A(n26), .Y(n300) );
  MUX41X1_HVT U44 ( .A1(n205), .A3(n207), .A2(n206), .A4(n208), .S0(n329), 
        .S1(n12), .Y(n209) );
  NAND2X0_HVT U45 ( .A1(n156), .A2(n270), .Y(n18) );
  NAND2X0_HVT U46 ( .A1(n155), .A2(n429), .Y(n19) );
  NAND2X0_HVT U47 ( .A1(n18), .A2(n19), .Y(n158) );
  MUX21X1_HVT U48 ( .A1(n409), .A2(n410), .S0(n413), .Y(n93) );
  XOR2X2_HVT U49 ( .A1(n451), .A2(n457), .Y(n51) );
  INVX1_HVT U50 ( .A(n363), .Y(n23) );
  INVX0_HVT U52 ( .A(in[1]), .Y(n363) );
  INVX1_HVT U53 ( .A(n224), .Y(n278) );
  INVX1_HVT U54 ( .A(n349), .Y(n119) );
  INVX1_HVT U55 ( .A(n17), .Y(n285) );
  INVX1_HVT U57 ( .A(n363), .Y(n458) );
  OR2X1_HVT U59 ( .A1(n439), .A2(n23), .Y(n36) );
  INVX1_HVT U60 ( .A(n456), .Y(n461) );
  INVX1_HVT U61 ( .A(n7), .Y(n383) );
  INVX0_HVT U63 ( .A(n36), .Y(n256) );
  INVX1_HVT U64 ( .A(in[4]), .Y(n255) );
  MUX21X2_HVT U65 ( .A1(n390), .A2(n266), .S0(n401), .Y(n99) );
  MUX21X1_HVT U67 ( .A1(n391), .A2(n346), .S0(n340), .Y(n167) );
  NAND2X0_HVT U69 ( .A1(n448), .A2(n50), .Y(n78) );
  NAND2X0_HVT U70 ( .A1(n386), .A2(n459), .Y(n118) );
  NAND2X0_HVT U71 ( .A1(n78), .A2(n118), .Y(n38) );
  INVX0_HVT U72 ( .A(n459), .Y(n50) );
  INVX1_HVT U75 ( .A(n460), .Y(n355) );
  AND2X1_HVT U76 ( .A1(n458), .A2(n2), .Y(n127) );
  IBUFFX2_HVT U78 ( .A(n471), .Y(n468) );
  NAND2X0_HVT U79 ( .A1(n96), .A2(n321), .Y(n210) );
  NAND2X0_HVT U80 ( .A1(n95), .A2(n429), .Y(n211) );
  NAND2X0_HVT U81 ( .A1(n210), .A2(n211), .Y(n98) );
  MUX21X1_HVT U82 ( .A1(n442), .A2(n441), .S0(n464), .Y(n312) );
  MUX21X1_HVT U84 ( .A1(n449), .A2(n441), .S0(n356), .Y(n212) );
  INVX1_HVT U87 ( .A(n449), .Y(n266) );
  OA21X1_HVT U88 ( .A1(n35), .A2(n472), .A3(n284), .Y(n188) );
  NAND2X0_HVT U89 ( .A1(n15), .A2(n213), .Y(n216) );
  NAND2X0_HVT U90 ( .A1(n405), .A2(n332), .Y(n217) );
  NAND2X0_HVT U91 ( .A1(n216), .A2(n217), .Y(n103) );
  INVX0_HVT U92 ( .A(n308), .Y(n213) );
  NAND2X0_HVT U93 ( .A1(n240), .A2(n50), .Y(n218) );
  NAND2X0_HVT U94 ( .A1(n406), .A2(n401), .Y(n219) );
  NAND2X0_HVT U95 ( .A1(n218), .A2(n219), .Y(n405) );
  MUX21X1_HVT U98 ( .A1(n451), .A2(n446), .S0(n364), .Y(n15) );
  INVX1_HVT U99 ( .A(n388), .Y(n392) );
  MUX41X1_HVT U100 ( .A1(n93), .A3(n100), .A2(n98), .A4(n101), .S0(n329), .S1(
        n231), .Y(n102) );
  MUX21X2_HVT U102 ( .A1(n132), .A2(n133), .S0(n231), .Y(n134) );
  INVX0_HVT U104 ( .A(n388), .Y(n391) );
  MUX21X2_HVT U106 ( .A1(n385), .A2(n440), .S0(n457), .Y(n79) );
  NBUFFX4_HVT U107 ( .A(in[3]), .Y(n437) );
  INVX0_HVT U108 ( .A(n37), .Y(n252) );
  INVX1_HVT U109 ( .A(n462), .Y(n424) );
  INVX1_HVT U111 ( .A(n424), .Y(n425) );
  INVX0_HVT U112 ( .A(n448), .Y(n282) );
  INVX0_HVT U113 ( .A(n424), .Y(n426) );
  MUX21X1_HVT U114 ( .A1(n447), .A2(n455), .S0(n402), .Y(n97) );
  INVX1_HVT U116 ( .A(n429), .Y(n308) );
  INVX1_HVT U117 ( .A(n11), .Y(n242) );
  INVX1_HVT U118 ( .A(n116), .Y(n263) );
  NAND2X0_HVT U119 ( .A1(n268), .A2(n413), .Y(n396) );
  INVX1_HVT U120 ( .A(n426), .Y(n341) );
  INVX1_HVT U121 ( .A(n426), .Y(n270) );
  AO21X1_HVT U122 ( .A1(n347), .A2(n246), .A3(n472), .Y(n106) );
  INVX1_HVT U123 ( .A(in[7]), .Y(n472) );
  INVX1_HVT U124 ( .A(n223), .Y(n247) );
  INVX1_HVT U125 ( .A(n432), .Y(n336) );
  INVX0_HVT U126 ( .A(n433), .Y(n398) );
  INVX0_HVT U127 ( .A(n460), .Y(n459) );
  INVX1_HVT U128 ( .A(n383), .Y(n388) );
  MUX21X1_HVT U129 ( .A1(n181), .A2(n328), .S0(n332), .Y(n380) );
  MUX21X1_HVT U130 ( .A1(n39), .A2(n253), .S0(n332), .Y(n381) );
  MUX41X1_HVT U131 ( .A1(n20), .A3(n277), .A2(n11), .A4(n58), .S0(n376), .S1(
        n466), .Y(n60) );
  MUX41X1_HVT U132 ( .A1(n3), .A3(n369), .A2(n405), .A4(n254), .S0(n270), .S1(
        n469), .Y(n208) );
  MUX21X1_HVT U133 ( .A1(n278), .A2(n246), .S0(n433), .Y(n155) );
  NAND2X0_HVT U134 ( .A1(n369), .A2(n235), .Y(n232) );
  INVX1_HVT U136 ( .A(n463), .Y(n321) );
  MUX21X1_HVT U137 ( .A1(n453), .A2(n452), .S0(n458), .Y(n191) );
  MUX41X1_HVT U138 ( .A1(n195), .A3(n51), .A2(n36), .A4(n43), .S0(n341), .S1(
        n338), .Y(n196) );
  INVX0_HVT U139 ( .A(n235), .Y(n236) );
  INVX1_HVT U143 ( .A(in[3]), .Y(n235) );
  MUX21X1_HVT U144 ( .A1(n447), .A2(n236), .S0(n458), .Y(n9) );
  INVX0_HVT U145 ( .A(n38), .Y(n274) );
  MUX41X1_HVT U148 ( .A1(n184), .A3(n182), .A2(n183), .A4(n180), .S0(n435), 
        .S1(n466), .Y(n185) );
  NBUFFX2_HVT U149 ( .A(n466), .Y(n430) );
  MUX41X1_HVT U150 ( .A1(n139), .A3(n126), .A2(n134), .A4(n120), .S0(n318), 
        .S1(n435), .Y(out[3]) );
  MUX41X1_HVT U151 ( .A1(n158), .A3(n159), .A2(n163), .A4(n165), .S0(n231), 
        .S1(n329), .Y(n166) );
  MUX21X1_HVT U152 ( .A1(n161), .A2(n162), .S0(n332), .Y(n163) );
  INVX1_HVT U155 ( .A(in[0]), .Y(n329) );
  OA21X1_HVT U156 ( .A1(n298), .A2(n472), .A3(n32), .Y(n151) );
  XOR2X2_HVT U157 ( .A1(n425), .A2(n467), .Y(n48) );
  MUX41X1_HVT U160 ( .A1(n300), .A3(n13), .A2(n32), .A4(n121), .S0(n376), .S1(
        n238), .Y(n122) );
  INVX1_HVT U161 ( .A(n332), .Y(n238) );
  INVX0_HVT U164 ( .A(n469), .Y(n376) );
  NAND2X0_HVT U165 ( .A1(n346), .A2(n50), .Y(n243) );
  NAND2X0_HVT U169 ( .A1(n442), .A2(n459), .Y(n249) );
  NAND2X0_HVT U170 ( .A1(n243), .A2(n249), .Y(n35) );
  INVX0_HVT U171 ( .A(n35), .Y(n241) );
  NAND2X0_HVT U172 ( .A1(n252), .A2(n308), .Y(n259) );
  NAND2X0_HVT U173 ( .A1(n3), .A2(n464), .Y(n261) );
  NAND2X0_HVT U175 ( .A1(n259), .A2(n261), .Y(n113) );
  MUX41X1_HVT U178 ( .A1(n171), .A3(n177), .A2(n169), .A4(n174), .S0(n329), 
        .S1(n430), .Y(n178) );
  NAND2X0_HVT U179 ( .A1(n39), .A2(n303), .Y(n264) );
  NAND2X0_HVT U181 ( .A1(n265), .A2(n432), .Y(n269) );
  NAND2X0_HVT U182 ( .A1(n264), .A2(n269), .Y(n162) );
  INVX0_HVT U183 ( .A(n339), .Y(n39) );
  MUX21X2_HVT U184 ( .A1(n200), .A2(n199), .S0(n308), .Y(n201) );
  XNOR2X2_HVT U185 ( .A1(n438), .A2(n437), .Y(n7) );
  INVX1_HVT U186 ( .A(n338), .Y(n333) );
  INVX1_HVT U187 ( .A(n97), .Y(n265) );
  MUX21X2_HVT U188 ( .A1(n124), .A2(n123), .S0(n433), .Y(n125) );
  INVX1_HVT U190 ( .A(n384), .Y(n386) );
  INVX0_HVT U191 ( .A(n383), .Y(n387) );
  MUX41X1_HVT U192 ( .A1(n37), .A3(n295), .A2(n34), .A4(n417), .S0(n270), .S1(
        n303), .Y(n143) );
  MUX21X1_HVT U193 ( .A1(n350), .A2(n386), .S0(n50), .Y(n26) );
  INVX0_HVT U194 ( .A(n29), .Y(n250) );
  MUX21X2_HVT U195 ( .A1(n256), .A2(n241), .S0(n429), .Y(n123) );
  MUX41X1_HVT U196 ( .A1(n365), .A3(n58), .A2(n24), .A4(n241), .S0(n270), .S1(
        n470), .Y(n207) );
  INVX1_HVT U198 ( .A(n9), .Y(n258) );
  INVX1_HVT U199 ( .A(n7), .Y(n384) );
  NAND2X0_HVT U200 ( .A1(n280), .A2(n12), .Y(n271) );
  NAND2X0_HVT U201 ( .A1(n461), .A2(n466), .Y(n273) );
  NAND2X0_HVT U202 ( .A1(n271), .A2(n273), .Y(n68) );
  MUX21X1_HVT U204 ( .A1(n282), .A2(n436), .S0(n401), .Y(n280) );
  INVX1_HVT U205 ( .A(n255), .Y(n369) );
  NAND2X0_HVT U206 ( .A1(n204), .A2(n270), .Y(n283) );
  NAND2X0_HVT U207 ( .A1(n203), .A2(n463), .Y(n289) );
  NAND2X0_HVT U209 ( .A1(n283), .A2(n289), .Y(n205) );
  MUX21X1_HVT U210 ( .A1(n17), .A2(n416), .S0(n432), .Y(n203) );
  MUX41X1_HVT U211 ( .A1(n201), .A3(n198), .A2(n197), .A4(n196), .S0(n431), 
        .S1(n435), .Y(n202) );
  MUX21X1_HVT U213 ( .A1(n128), .A2(n129), .S0(n468), .Y(n132) );
  INVX0_HVT U216 ( .A(n460), .Y(n401) );
  MUX41X1_HVT U217 ( .A1(n114), .A3(n117), .A2(n113), .A4(n119), .S0(n231), 
        .S1(n398), .Y(n120) );
  MUX21X2_HVT U219 ( .A1(n127), .A2(n30), .S0(n303), .Y(n150) );
  MUX41X1_HVT U221 ( .A1(n71), .A3(n63), .A2(n67), .A4(n57), .S0(n318), .S1(
        n435), .Y(out[0]) );
  NAND2X0_HVT U222 ( .A1(n56), .A2(n308), .Y(n293) );
  NAND2X0_HVT U223 ( .A1(n52), .A2(n428), .Y(n297) );
  NAND2X0_HVT U224 ( .A1(n293), .A2(n297), .Y(n57) );
  MUX21X1_HVT U225 ( .A1(n54), .A2(n53), .S0(n432), .Y(n56) );
  INVX0_HVT U226 ( .A(n450), .Y(n296) );
  NAND2X0_HVT U227 ( .A1(n255), .A2(n236), .Y(n2) );
  INVX1_HVT U228 ( .A(n337), .Y(n170) );
  MUX21X1_HVT U229 ( .A1(n442), .A2(n330), .S0(n331), .Y(n222) );
  INVX0_HVT U230 ( .A(n405), .Y(n32) );
  MUX21X2_HVT U231 ( .A1(n440), .A2(n266), .S0(n402), .Y(n30) );
  NBUFFX2_HVT U232 ( .A(n467), .Y(n434) );
  INVX0_HVT U233 ( .A(n364), .Y(n340) );
  NAND2X0_HVT U234 ( .A1(n115), .A2(n213), .Y(n304) );
  NAND2X0_HVT U235 ( .A1(n32), .A2(n308), .Y(n305) );
  NAND2X0_HVT U236 ( .A1(n304), .A2(n305), .Y(n117) );
  INVX0_HVT U237 ( .A(n355), .Y(n331) );
  NAND2X0_HVT U238 ( .A1(n4), .A2(n315), .Y(n306) );
  NAND2X0_HVT U239 ( .A1(n144), .A2(n308), .Y(n307) );
  NAND2X0_HVT U240 ( .A1(n306), .A2(n307), .Y(n145) );
  XOR2X1_HVT U243 ( .A1(n472), .A2(n28), .Y(n45) );
  NAND2X0_HVT U244 ( .A1(n55), .A2(n44), .Y(n54) );
  INVX0_HVT U246 ( .A(n280), .Y(n309) );
  INVX1_HVT U248 ( .A(n363), .Y(n456) );
  INVX0_HVT U249 ( .A(n453), .Y(n240) );
  INVX1_HVT U250 ( .A(in[1]), .Y(n460) );
  NAND2X0_HVT U251 ( .A1(n436), .A2(n12), .Y(n310) );
  NAND2X0_HVT U252 ( .A1(n36), .A2(n466), .Y(n311) );
  NAND2X0_HVT U253 ( .A1(n310), .A2(n311), .Y(n53) );
  INVX1_HVT U254 ( .A(in[2]), .Y(n465) );
  INVX0_HVT U255 ( .A(n40), .Y(n268) );
  INVX0_HVT U257 ( .A(n320), .Y(n328) );
  INVX1_HVT U258 ( .A(n384), .Y(n385) );
  INVX1_HVT U259 ( .A(n460), .Y(n402) );
  MUX41X1_HVT U260 ( .A1(n447), .A3(n268), .A2(n257), .A4(n292), .S0(n336), 
        .S1(n462), .Y(n186) );
  MUX41X1_HVT U261 ( .A1(n189), .A3(n186), .A2(n193), .A4(n190), .S0(n430), 
        .S1(n329), .Y(n194) );
  AND3X2_HVT U262 ( .A1(n450), .A2(n59), .A3(n84), .Y(n83) );
  NAND2X0_HVT U263 ( .A1(n89), .A2(n336), .Y(n313) );
  NAND2X0_HVT U264 ( .A1(n436), .A2(n433), .Y(n314) );
  NAND2X0_HVT U266 ( .A1(n313), .A2(n314), .Y(n187) );
  NAND2X0_HVT U267 ( .A1(n187), .A2(n315), .Y(n316) );
  NAND2X0_HVT U269 ( .A1(n188), .A2(n321), .Y(n317) );
  NAND2X0_HVT U271 ( .A1(n316), .A2(n317), .Y(n189) );
  INVX0_HVT U272 ( .A(n321), .Y(n315) );
  INVX1_HVT U273 ( .A(n377), .Y(n318) );
  INVX1_HVT U274 ( .A(in[6]), .Y(n377) );
  MUX41X1_HVT U275 ( .A1(n296), .A3(n300), .A2(n244), .A4(n247), .S0(n427), 
        .S1(n472), .Y(n319) );
  IBUFFX2_HVT U276 ( .A(n59), .Y(n244) );
  MUX21X1_HVT U277 ( .A1(n330), .A2(n441), .S0(n340), .Y(n320) );
  MUX21X2_HVT U278 ( .A1(n240), .A2(n350), .S0(n331), .Y(n28) );
  MUX21X1_HVT U279 ( .A1(n347), .A2(n3), .S0(n321), .Y(n131) );
  INVX0_HVT U280 ( .A(n359), .Y(n128) );
  NAND2X0_HVT U281 ( .A1(n266), .A2(n50), .Y(n322) );
  NAND2X0_HVT U282 ( .A1(n296), .A2(n459), .Y(n323) );
  NAND2X0_HVT U285 ( .A1(n322), .A2(n323), .Y(n179) );
  INVX0_HVT U286 ( .A(n452), .Y(n350) );
  INVX1_HVT U287 ( .A(n465), .Y(n463) );
  INVX1_HVT U288 ( .A(n453), .Y(n346) );
  INVX1_HVT U290 ( .A(n460), .Y(n457) );
  NAND2X0_HVT U291 ( .A1(n72), .A2(n315), .Y(n324) );
  NAND2X0_HVT U292 ( .A1(n45), .A2(n332), .Y(n325) );
  NAND2X0_HVT U293 ( .A1(n324), .A2(n325), .Y(n73) );
  INVX1_HVT U294 ( .A(n429), .Y(n332) );
  NBUFFX2_HVT U297 ( .A(n255), .Y(n441) );
  NAND2X0_HVT U298 ( .A1(n64), .A2(n315), .Y(n326) );
  NAND2X0_HVT U299 ( .A1(n66), .A2(n341), .Y(n327) );
  NAND2X0_HVT U301 ( .A1(n326), .A2(n327), .Y(n67) );
  MUX21X1_HVT U304 ( .A1(n419), .A2(n285), .S0(n428), .Y(n137) );
  NBUFFX2_HVT U305 ( .A(n10), .Y(n330) );
  MUX21X1_HVT U307 ( .A1(n346), .A2(n245), .S0(n434), .Y(n72) );
  INVX1_HVT U308 ( .A(n382), .Y(n338) );
  OA21X1_HVT U310 ( .A1(n274), .A2(n465), .A3(n352), .Y(n114) );
  NAND2X0_HVT U311 ( .A1(n302), .A2(n341), .Y(n334) );
  NAND2X0_HVT U312 ( .A1(n140), .A2(n428), .Y(n335) );
  NAND2X0_HVT U313 ( .A1(n334), .A2(n335), .Y(n141) );
  MUX21X1_HVT U314 ( .A1(n267), .A2(n330), .S0(n433), .Y(n140) );
  MUX41X1_HVT U315 ( .A1(n152), .A3(n148), .A2(n153), .A4(n149), .S0(n435), 
        .S1(n231), .Y(n154) );
  MUX41X1_HVT U316 ( .A1(n423), .A3(n22), .A2(n267), .A4(n286), .S0(n321), 
        .S1(n468), .Y(n133) );
  MUX21X1_HVT U317 ( .A1(n440), .A2(n266), .S0(n340), .Y(n226) );
  MUX21X1_HVT U318 ( .A1(n449), .A2(n454), .S0(n340), .Y(n339) );
  INVX1_HVT U319 ( .A(n227), .Y(n279) );
  INVX1_HVT U320 ( .A(n226), .Y(n267) );
  INVX0_HVT U321 ( .A(n41), .Y(n299) );
  MUX41X1_HVT U322 ( .A1(n28), .A3(n42), .A2(n446), .A4(n279), .S0(n336), .S1(
        n425), .Y(n197) );
  INVX1_HVT U323 ( .A(n222), .Y(n245) );
  NBUFFX2_HVT U324 ( .A(n232), .Y(n446) );
  MUX21X1_HVT U325 ( .A1(n294), .A2(n92), .S0(n464), .Y(n410) );
  MUX21X1_HVT U326 ( .A1(n451), .A2(n446), .S0(n347), .Y(n337) );
  MUX41X1_HVT U327 ( .A1(n170), .A3(n47), .A2(n251), .A4(n22), .S0(n338), .S1(
        n424), .Y(n171) );
  NAND2X0_HVT U328 ( .A1(n131), .A2(n130), .Y(n129) );
  MUX41X1_HVT U329 ( .A1(n245), .A3(n385), .A2(n38), .A4(n453), .S0(n341), 
        .S1(n470), .Y(n198) );
  NAND2X0_HVT U330 ( .A1(n176), .A2(n315), .Y(n342) );
  NAND2X0_HVT U331 ( .A1(n175), .A2(n270), .Y(n343) );
  NAND2X0_HVT U332 ( .A1(n342), .A2(n343), .Y(n177) );
  NAND2X0_HVT U333 ( .A1(n60), .A2(n315), .Y(n344) );
  NAND2X0_HVT U334 ( .A1(n62), .A2(n341), .Y(n345) );
  NAND2X0_HVT U335 ( .A1(n344), .A2(n345), .Y(n63) );
  NAND2X0_HVT U336 ( .A1(n350), .A2(n347), .Y(n348) );
  NAND2X0_HVT U337 ( .A1(n348), .A2(n394), .Y(n20) );
  INVX0_HVT U338 ( .A(n402), .Y(n347) );
  INVX1_HVT U339 ( .A(n221), .Y(n277) );
  NBUFFX2_HVT U340 ( .A(n235), .Y(n443) );
  MUX21X1_HVT U341 ( .A1(n446), .A2(n447), .S0(n393), .Y(n352) );
  NAND2X0_HVT U342 ( .A1(n125), .A2(n231), .Y(n353) );
  NAND2X0_HVT U343 ( .A1(n122), .A2(n430), .Y(n354) );
  NAND2X0_HVT U344 ( .A1(n353), .A2(n354), .Y(n126) );
  IBUFFX2_HVT U345 ( .A(n460), .Y(n356) );
  NAND2X0_HVT U346 ( .A1(n441), .A2(n331), .Y(n357) );
  NAND2X0_HVT U347 ( .A1(n443), .A2(n355), .Y(n358) );
  MUX21X1_HVT U348 ( .A1(n34), .A2(n360), .S0(n463), .Y(n359) );
  AND2X1_HVT U349 ( .A1(n357), .A2(n358), .Y(n360) );
  NAND2X0_HVT U350 ( .A1(n451), .A2(n366), .Y(n361) );
  NAND2X0_HVT U351 ( .A1(n94), .A2(n421), .Y(n362) );
  NAND2X0_HVT U352 ( .A1(n361), .A2(n362), .Y(n95) );
  MUX21X1_HVT U353 ( .A1(n436), .A2(n440), .S0(n434), .Y(n94) );
  INVX1_HVT U354 ( .A(n363), .Y(n364) );
  INVX0_HVT U355 ( .A(n421), .Y(n366) );
  NAND2X0_HVT U356 ( .A1(n14), .A2(n454), .Y(n365) );
  MUX41X1_HVT U357 ( .A1(n104), .A3(n109), .A2(n108), .A4(n111), .S0(n329), 
        .S1(n231), .Y(n112) );
  NAND2X0_HVT U358 ( .A1(n160), .A2(n366), .Y(n367) );
  NAND2X0_HVT U359 ( .A1(n450), .A2(n421), .Y(n368) );
  NAND2X0_HVT U360 ( .A1(n367), .A2(n368), .Y(n161) );
  NAND2X0_HVT U361 ( .A1(n14), .A2(n454), .Y(n13) );
  MUX41X1_HVT U362 ( .A1(n86), .A3(n90), .A2(n85), .A4(n88), .S0(n329), .S1(
        n430), .Y(n91) );
  XNOR2X1_HVT U363 ( .A1(n369), .A2(n401), .Y(n27) );
  MUX41X1_HVT U364 ( .A1(n389), .A3(n285), .A2(n320), .A4(n415), .S0(n336), 
        .S1(n12), .Y(n64) );
  INVX0_HVT U365 ( .A(n21), .Y(n291) );
  OA21X1_HVT U366 ( .A1(n8), .A2(n472), .A3(n339), .Y(n204) );
  NAND2X0_HVT U367 ( .A1(n146), .A2(n318), .Y(n370) );
  NAND2X0_HVT U368 ( .A1(n154), .A2(n377), .Y(n371) );
  NAND2X0_HVT U369 ( .A1(n370), .A2(n371), .Y(out[4]) );
  MUX41X1_HVT U370 ( .A1(n352), .A3(n422), .A2(n61), .A4(n423), .S0(n376), 
        .S1(n12), .Y(n62) );
  XNOR2X1_HVT U371 ( .A1(n384), .A2(n364), .Y(n47) );
  MUX41X1_HVT U372 ( .A1(n40), .A3(n420), .A2(n47), .A4(n76), .S0(n424), .S1(
        n333), .Y(n190) );
  OA21X1_HVT U373 ( .A1(n41), .A2(n472), .A3(n157), .Y(n156) );
  MUX41X1_HVT U374 ( .A1(n275), .A3(n290), .A2(n65), .A4(n288), .S0(n470), 
        .S1(n12), .Y(n66) );
  INVX1_HVT U375 ( .A(n471), .Y(n467) );
  MUX41X1_HVT U376 ( .A1(n276), .A3(n253), .A2(n29), .A4(n254), .S0(n464), 
        .S1(n398), .Y(n183) );
  INVX1_HVT U377 ( .A(n225), .Y(n302) );
  NAND2X0_HVT U378 ( .A1(n381), .A2(n413), .Y(n372) );
  NAND2X0_HVT U379 ( .A1(n380), .A2(n376), .Y(n373) );
  NAND2X0_HVT U380 ( .A1(n372), .A2(n373), .Y(n182) );
  AO21X1_HVT U381 ( .A1(n429), .A2(n446), .A3(n385), .Y(n124) );
  INVX1_HVT U382 ( .A(n230), .Y(n254) );
  NAND2X0_HVT U383 ( .A1(n43), .A2(n213), .Y(n374) );
  NAND2X0_HVT U384 ( .A1(n47), .A2(n332), .Y(n375) );
  NAND2X0_HVT U385 ( .A1(n374), .A2(n375), .Y(n409) );
  NAND2X0_HVT U386 ( .A1(n91), .A2(n377), .Y(n378) );
  NAND2X0_HVT U387 ( .A1(n81), .A2(n318), .Y(n379) );
  NAND2X0_HVT U388 ( .A1(n378), .A2(n379), .Y(out[1]) );
  NAND2X0_HVT U389 ( .A1(n194), .A2(n377), .Y(n399) );
  INVX1_HVT U390 ( .A(n229), .Y(n253) );
  INVX1_HVT U391 ( .A(n388), .Y(n390) );
  NAND2X0_HVT U392 ( .A1(n436), .A2(n393), .Y(n394) );
  NAND2X0_HVT U393 ( .A1(n390), .A2(n331), .Y(n395) );
  NAND2X0_HVT U394 ( .A1(n394), .A2(n395), .Y(n24) );
  INVX1_HVT U395 ( .A(n363), .Y(n393) );
  INVX0_HVT U396 ( .A(n24), .Y(n284) );
  NAND2X0_HVT U397 ( .A1(n178), .A2(n377), .Y(n403) );
  NBUFFX2_HVT U398 ( .A(in[4]), .Y(n439) );
  MUX41X1_HVT U399 ( .A1(n137), .A3(n135), .A2(n138), .A4(n136), .S0(n430), 
        .S1(n336), .Y(n139) );
  NBUFFX2_HVT U400 ( .A(n255), .Y(n440) );
  MUX41X1_HVT U401 ( .A1(n145), .A3(n143), .A2(n142), .A4(n141), .S0(n430), 
        .S1(n435), .Y(n146) );
  NAND2X0_HVT U402 ( .A1(n24), .A2(n398), .Y(n397) );
  NAND2X0_HVT U403 ( .A1(n396), .A2(n397), .Y(n144) );
  INVX1_HVT U404 ( .A(n8), .Y(n286) );
  MUX21X1_HVT U405 ( .A1(n389), .A2(n240), .S0(n457), .Y(n8) );
  NAND2X0_HVT U406 ( .A1(n185), .A2(in[6]), .Y(n400) );
  NAND2X0_HVT U407 ( .A1(n400), .A2(n399), .Y(out[6]) );
  MUX41X1_HVT U408 ( .A1(n87), .A3(n17), .A2(n386), .A4(n284), .S0(n321), .S1(
        n472), .Y(n88) );
  NAND2X0_HVT U409 ( .A1(n166), .A2(n318), .Y(n404) );
  NAND2X0_HVT U410 ( .A1(n404), .A2(n403), .Y(out[5]) );
  MUX41X1_HVT U411 ( .A1(n233), .A3(n15), .A2(n46), .A4(n291), .S0(n427), .S1(
        n472), .Y(n86) );
  MUX41X1_HVT U412 ( .A1(n73), .A3(n319), .A2(n77), .A4(n80), .S0(n329), .S1(
        n231), .Y(n81) );
  NAND2X0_HVT U413 ( .A1(n209), .A2(n377), .Y(n407) );
  NAND2X0_HVT U414 ( .A1(n202), .A2(n318), .Y(n408) );
  NAND2X0_HVT U415 ( .A1(n407), .A2(n408), .Y(out[7]) );
  NAND2X0_HVT U416 ( .A1(n112), .A2(n377), .Y(n411) );
  NAND2X0_HVT U417 ( .A1(n102), .A2(n318), .Y(n412) );
  NAND2X0_HVT U418 ( .A1(n411), .A2(n412), .Y(out[2]) );
  NBUFFX2_HVT U419 ( .A(n5), .Y(n447) );
  NBUFFX2_HVT U420 ( .A(n5), .Y(n448) );
  NBUFFX2_HVT U421 ( .A(n5), .Y(n449) );
  MUX21X1_HVT U422 ( .A1(n258), .A2(n246), .S0(n466), .Y(n70) );
  AND2X1_HVT U423 ( .A1(n454), .A2(n116), .Y(n415) );
  AND2X1_HVT U424 ( .A1(n391), .A2(n59), .Y(n416) );
  AND2X1_HVT U425 ( .A1(n450), .A2(n76), .Y(n417) );
  NAND2X0_HVT U426 ( .A1(n255), .A2(n235), .Y(n5) );
  MUX21X1_HVT U427 ( .A1(n330), .A2(n455), .S0(n428), .Y(n130) );
  MUX21X1_HVT U428 ( .A1(n443), .A2(n240), .S0(n364), .Y(n11) );
  MUX21X1_HVT U429 ( .A1(n452), .A2(n441), .S0(n393), .Y(n220) );
  MUX21X1_HVT U430 ( .A1(n452), .A2(n389), .S0(n355), .Y(n42) );
  MUX21X1_HVT U431 ( .A1(n392), .A2(n441), .S0(n401), .Y(n107) );
  MUX21X1_HVT U432 ( .A1(n442), .A2(n441), .S0(n457), .Y(n195) );
  XOR2X1_HVT U433 ( .A1(n356), .A2(n246), .Y(n46) );
  MUX21X1_HVT U434 ( .A1(n448), .A2(n330), .S0(n356), .Y(n92) );
  MUX21X1_HVT U435 ( .A1(n443), .A2(n455), .S0(n459), .Y(n192) );
  MUX21X1_HVT U436 ( .A1(n445), .A2(n440), .S0(n364), .Y(n74) );
  MUX21X1_HVT U437 ( .A1(n442), .A2(n386), .S0(n458), .Y(n224) );
  MUX21X1_HVT U438 ( .A1(n266), .A2(n346), .S0(n466), .Y(n55) );
  XOR2X1_HVT U439 ( .A1(n402), .A2(n431), .Y(n44) );
  MUX21X1_HVT U440 ( .A1(n385), .A2(n246), .S0(n393), .Y(n227) );
  XNOR2X1_HVT U441 ( .A1(n453), .A2(n459), .Y(n418) );
  XNOR2X1_HVT U442 ( .A1(n447), .A2(n459), .Y(n419) );
  MUX21X1_HVT U443 ( .A1(n451), .A2(n447), .S0(n355), .Y(n228) );
  NBUFFX2_HVT U444 ( .A(n10), .Y(n444) );
  AND2X1_HVT U445 ( .A1(n458), .A2(n296), .Y(n420) );
  NBUFFX2_HVT U446 ( .A(n232), .Y(n445) );
  NBUFFX2_HVT U447 ( .A(n1), .Y(n453) );
  NBUFFX2_HVT U448 ( .A(n2), .Y(n450) );
  NBUFFX2_HVT U449 ( .A(n2), .Y(n451) );
  NBUFFX2_HVT U450 ( .A(n235), .Y(n442) );
  NBUFFX2_HVT U451 ( .A(n2), .Y(n452) );
  NBUFFX2_HVT U452 ( .A(n1), .Y(n455) );
  NBUFFX2_HVT U453 ( .A(n1), .Y(n454) );
  NBUFFX2_HVT U454 ( .A(in[5]), .Y(n431) );
  NBUFFX2_HVT U455 ( .A(n467), .Y(n432) );
  NBUFFX2_HVT U456 ( .A(n467), .Y(n433) );
  NBUFFX2_HVT U457 ( .A(n464), .Y(n428) );
  NBUFFX2_HVT U458 ( .A(n464), .Y(n429) );
  NBUFFX2_HVT U459 ( .A(n463), .Y(n427) );
  MUX21X1_HVT U460 ( .A1(n439), .A2(n452), .S0(n393), .Y(n21) );
  MUX21X1_HVT U461 ( .A1(n439), .A2(n385), .S0(n393), .Y(n221) );
  MUX21X1_HVT U462 ( .A1(n436), .A2(n266), .S0(n355), .Y(n40) );
  MUX21X1_HVT U463 ( .A1(n455), .A2(n439), .S0(n23), .Y(n29) );
  MUX21X1_HVT U464 ( .A1(n439), .A2(n445), .S0(n401), .Y(n229) );
  MUX21X1_HVT U465 ( .A1(n105), .A2(n302), .S0(n428), .Y(n108) );
  XOR2X1_HVT U466 ( .A1(n402), .A2(n436), .Y(n49) );
  MUX21X1_HVT U467 ( .A1(n445), .A2(n391), .S0(n356), .Y(n110) );
  MUX21X1_HVT U468 ( .A1(n330), .A2(n245), .S0(n434), .Y(n175) );
  MUX21X1_HVT U469 ( .A1(n439), .A2(n454), .S0(n23), .Y(n230) );
  MUX21X1_HVT U470 ( .A1(n436), .A2(n246), .S0(n458), .Y(n223) );
  XNOR2X1_HVT U471 ( .A1(n471), .A2(n355), .Y(n421) );
  NAND2X0_HVT U472 ( .A1(n369), .A2(n235), .Y(n10) );
  AND2X1_HVT U473 ( .A1(n390), .A2(n461), .Y(n422) );
  NAND2X0_HVT U474 ( .A1(n438), .A2(n437), .Y(n1) );
  AND2X1_HVT U475 ( .A1(n443), .A2(n461), .Y(n423) );
  INVX1_HVT U476 ( .A(n465), .Y(n462) );
  NBUFFX2_HVT U477 ( .A(in[5]), .Y(n466) );
  NBUFFX2_HVT U478 ( .A(in[3]), .Y(n436) );
  NBUFFX2_HVT U479 ( .A(in[0]), .Y(n435) );
endmodule

