
module sbox_4 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n14, n23, n210, n211, n212, n213, n216, n217, n218, n219, n224, n226,
         n227, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605;

  NAND2X0_HVT U3 ( .A1(n252), .A2(n320), .Y(n603) );
  NAND2X0_HVT U4 ( .A1(n318), .A2(n603), .Y(n602) );
  NAND2X0_HVT U5 ( .A1(n252), .A2(n305), .Y(n600) );
  NAND2X0_HVT U13 ( .A1(n244), .A2(n323), .Y(n593) );
  NAND2X0_HVT U15 ( .A1(n603), .A2(n307), .Y(n591) );
  NAND2X0_HVT U21 ( .A1(n318), .A2(n264), .Y(n585) );
  NAND2X0_HVT U24 ( .A1(n313), .A2(n263), .Y(n583) );
  NAND2X0_HVT U33 ( .A1(n383), .A2(n264), .Y(n574) );
  NAND2X0_HVT U35 ( .A1(n311), .A2(n264), .Y(n572) );
  NAND2X0_HVT U42 ( .A1(n252), .A2(n313), .Y(n565) );
  NAND2X0_HVT U53 ( .A1(n553), .A2(n564), .Y(n554) );
  NAND2X0_HVT U56 ( .A1(n318), .A2(n549), .Y(n550) );
  MUX41X1_HVT U57 ( .A1(n375), .A3(n587), .A2(n550), .A4(n595), .S0(n331), 
        .S1(n299), .Y(n548) );
  NAND2X0_HVT U58 ( .A1(n323), .A2(n603), .Y(n547) );
  MUX41X1_HVT U59 ( .A1(n292), .A3(n547), .A2(n290), .A4(n350), .S0(n331), 
        .S1(n299), .Y(n546) );
  MUX41X1_HVT U61 ( .A1(n288), .A3(n349), .A2(n348), .A4(n306), .S0(n331), 
        .S1(n299), .Y(n544) );
  NAND2X0_HVT U62 ( .A1(n263), .A2(n321), .Y(n543) );
  MUX41X1_HVT U63 ( .A1(n543), .A3(n341), .A2(n369), .A4(n347), .S0(n331), 
        .S1(n299), .Y(n542) );
  AO21X1_HVT U66 ( .A1(n345), .A2(n301), .A3(n368), .Y(n539) );
  MUX41X1_HVT U68 ( .A1(n343), .A3(n539), .A2(n538), .A4(n540), .S0(n293), 
        .S1(n276), .Y(n537) );
  MUX41X1_HVT U69 ( .A1(n537), .A3(n545), .A2(n541), .A4(n551), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n315), .A2(n532), .Y(n533) );
  MUX41X1_HVT U74 ( .A1(n534), .A3(n581), .A2(n533), .A4(n583), .S0(n295), 
        .S1(n330), .Y(n531) );
  MUX41X1_HVT U75 ( .A1(n372), .A3(n377), .A2(n387), .A4(n354), .S0(n293), 
        .S1(n276), .Y(n530) );
  MUX41X1_HVT U77 ( .A1(n597), .A3(n378), .A2(n529), .A4(n261), .S0(n302), 
        .S1(n329), .Y(n528) );
  MUX41X1_HVT U78 ( .A1(n528), .A3(n531), .A2(n530), .A4(n535), .S0(in[0]), 
        .S1(n299), .Y(n527) );
  AND3X1_HVT U80 ( .A1(n320), .A2(n549), .A3(n524), .Y(n525) );
  AND2X1_HVT U83 ( .A1(n236), .A2(n245), .Y(n521) );
  NAND2X0_HVT U85 ( .A1(n264), .A2(n386), .Y(n519) );
  AO21X1_HVT U93 ( .A1(n304), .A2(n511), .A3(n373), .Y(n512) );
  MUX41X1_HVT U96 ( .A1(n336), .A3(n287), .A2(n376), .A4(n509), .S0(n293), 
        .S1(n238), .Y(n508) );
  MUX41X1_HVT U97 ( .A1(n372), .A3(n287), .A2(n236), .A4(n591), .S0(n293), 
        .S1(n238), .Y(n507) );
  NAND2X0_HVT U101 ( .A1(n502), .A2(n501), .Y(n503) );
  MUX41X1_HVT U103 ( .A1(n603), .A3(n344), .A2(n357), .A4(n572), .S0(n293), 
        .S1(n238), .Y(n499) );
  MUX41X1_HVT U105 ( .A1(n356), .A3(n559), .A2(n498), .A4(n371), .S0(n293), 
        .S1(n238), .Y(n497) );
  MUX41X1_HVT U106 ( .A1(n497), .A3(n500), .A2(n499), .A4(n504), .S0(in[0]), 
        .S1(in[5]), .Y(n496) );
  NAND2X0_HVT U110 ( .A1(n320), .A2(n492), .Y(n493) );
  AND2X1_HVT U115 ( .A1(n252), .A2(n306), .Y(n487) );
  NAND2X0_HVT U123 ( .A1(n478), .A2(n477), .Y(n479) );
  MUX41X1_HVT U125 ( .A1(n585), .A3(n292), .A2(n343), .A4(n246), .S0(n294), 
        .S1(n331), .Y(n475) );
  MUX41X1_HVT U131 ( .A1(n470), .A3(n472), .A2(n471), .A4(n473), .S0(n301), 
        .S1(n331), .Y(n469) );
  MUX41X1_HVT U136 ( .A1(n285), .A3(n574), .A2(n380), .A4(n571), .S0(n294), 
        .S1(n331), .Y(n465) );
  MUX41X1_HVT U139 ( .A1(n463), .A3(n466), .A2(n465), .A4(n467), .S0(n312), 
        .S1(n300), .Y(n462) );
  AND2X1_HVT U140 ( .A1(n314), .A2(n262), .Y(n461) );
  MUX41X1_HVT U141 ( .A1(n582), .A3(n255), .A2(n461), .A4(n361), .S0(n295), 
        .S1(n331), .Y(n460) );
  OA21X1_HVT U144 ( .A1(n338), .A2(n333), .A3(n576), .Y(n457) );
  NAND2X0_HVT U146 ( .A1(n252), .A2(n323), .Y(n532) );
  OA21X1_HVT U151 ( .A1(n567), .A2(n333), .A3(n451), .Y(n452) );
  AND2X1_HVT U154 ( .A1(n304), .A2(n313), .Y(n448) );
  NAND2X0_HVT U158 ( .A1(n236), .A2(n386), .Y(n444) );
  MUX41X1_HVT U159 ( .A1(n593), .A3(n306), .A2(n444), .A4(n273), .S0(n296), 
        .S1(n238), .Y(n443) );
  MUX41X1_HVT U160 ( .A1(n443), .A3(n449), .A2(n445), .A4(n450), .S0(n312), 
        .S1(n300), .Y(n442) );
  AND2X1_HVT U162 ( .A1(n250), .A2(n532), .Y(n440) );
  MUX41X1_HVT U163 ( .A1(n349), .A3(n440), .A2(n286), .A4(n441), .S0(n295), 
        .S1(n238), .Y(n439) );
  MUX41X1_HVT U165 ( .A1(n585), .A3(n358), .A2(n561), .A4(n438), .S0(n331), 
        .S1(n329), .Y(n437) );
  NAND2X0_HVT U166 ( .A1(n323), .A2(n549), .Y(n436) );
  NAND2X0_HVT U167 ( .A1(n387), .A2(n264), .Y(n435) );
  MUX41X1_HVT U168 ( .A1(n375), .A3(n314), .A2(n435), .A4(n436), .S0(n298), 
        .S1(n330), .Y(n434) );
  MUX41X1_HVT U176 ( .A1(n309), .A3(n429), .A2(n379), .A4(n244), .S0(n331), 
        .S1(n297), .Y(n428) );
  NAND2X0_HVT U177 ( .A1(n252), .A2(n310), .Y(n427) );
  MUX41X1_HVT U178 ( .A1(n589), .A3(n427), .A2(n381), .A4(n569), .S0(n295), 
        .S1(n330), .Y(n426) );
  MUX41X1_HVT U179 ( .A1(n579), .A3(n382), .A2(n339), .A4(n381), .S0(n329), 
        .S1(n276), .Y(n425) );
  MUX41X1_HVT U180 ( .A1(n342), .A3(n597), .A2(n593), .A4(n284), .S0(n302), 
        .S1(n329), .Y(n424) );
  MUX41X1_HVT U181 ( .A1(n424), .A3(n426), .A2(n425), .A4(n428), .S0(n312), 
        .S1(n300), .Y(n423) );
  MUX41X1_HVT U182 ( .A1(n364), .A3(n317), .A2(n366), .A4(n355), .S0(n331), 
        .S1(n329), .Y(n422) );
  OA21X1_HVT U184 ( .A1(n573), .A2(n333), .A3(n353), .Y(n420) );
  MUX41X1_HVT U189 ( .A1(n416), .A3(n244), .A2(n417), .A4(n371), .S0(n302), 
        .S1(n298), .Y(n415) );
  MUX41X1_HVT U193 ( .A1(n565), .A3(n572), .A2(n557), .A4(n413), .S0(n329), 
        .S1(n330), .Y(n412) );
  MUX41X1_HVT U194 ( .A1(n566), .A3(n580), .A2(n267), .A4(n314), .S0(n302), 
        .S1(n297), .Y(n411) );
  MUX41X1_HVT U195 ( .A1(n250), .A3(n376), .A2(n322), .A4(n570), .S0(n329), 
        .S1(n276), .Y(n410) );
  AO21X1_HVT U197 ( .A1(n289), .A2(n303), .A3(n373), .Y(n408) );
  OA21X1_HVT U201 ( .A1(n598), .A2(n333), .A3(n255), .Y(n404) );
  MUX41X1_HVT U203 ( .A1(n571), .A3(n365), .A2(n594), .A4(n575), .S0(n293), 
        .S1(n330), .Y(n402) );
  MUX41X1_HVT U204 ( .A1(n550), .A3(n593), .A2(n362), .A4(n584), .S0(n329), 
        .S1(n330), .Y(n401) );
  MUX41X1_HVT U205 ( .A1(n245), .A3(n603), .A2(n382), .A4(n360), .S0(n293), 
        .S1(n276), .Y(n400) );
  NAND2X0_HVT U208 ( .A1(n252), .A2(n318), .Y(n492) );
  NAND2X0_HVT U212 ( .A1(n252), .A2(n315), .Y(n549) );
  NAND2X0_HVT U214 ( .A1(n599), .A2(n263), .Y(n398) );
  NAND2X0_HVT U215 ( .A1(n492), .A2(n316), .Y(n397) );
  NAND2X0_HVT U218 ( .A1(n384), .A2(n324), .Y(n451) );
  NAND2X0_HVT U220 ( .A1(n303), .A2(n398), .Y(n524) );
  MUX21X2_HVT U1 ( .A1(n316), .A2(n586), .S0(n14), .Y(n526) );
  IBUFFX16_HVT U2 ( .A(n304), .Y(n14) );
  NAND2X0_HVT U6 ( .A1(n602), .A2(n23), .Y(n210) );
  NAND2X0_HVT U7 ( .A1(n464), .A2(n269), .Y(n211) );
  NAND2X0_HVT U8 ( .A1(n210), .A2(n211), .Y(n463) );
  IBUFFX2_HVT U9 ( .A(n269), .Y(n23) );
  MUX21X1_HVT U10 ( .A1(n364), .A2(n584), .S0(n270), .Y(n464) );
  INVX0_HVT U11 ( .A(n584), .Y(n353) );
  INVX2_HVT U12 ( .A(in[7]), .Y(n334) );
  MUX21X2_HVT U14 ( .A1(n457), .A2(n458), .S0(n212), .Y(n456) );
  IBUFFX16_HVT U16 ( .A(n297), .Y(n212) );
  MUX21X2_HVT U17 ( .A1(n512), .A2(n513), .S0(n298), .Y(n510) );
  INVX2_HVT U18 ( .A(n262), .Y(n324) );
  MUX21X1_HVT U19 ( .A1(n305), .A2(n315), .S0(n263), .Y(n394) );
  MUX21X1_HVT U20 ( .A1(n217), .A2(n216), .S0(n218), .Y(n213) );
  IBUFFX16_HVT U22 ( .A(n213), .Y(n535) );
  IBUFFX16_HVT U23 ( .A(n536), .Y(n216) );
  IBUFFX16_HVT U25 ( .A(n563), .Y(n217) );
  IBUFFX16_HVT U26 ( .A(n269), .Y(n218) );
  INVX1_HVT U27 ( .A(n263), .Y(n325) );
  NAND2X2_HVT U28 ( .A1(n226), .A2(n227), .Y(out[5]) );
  INVX2_HVT U29 ( .A(n262), .Y(n327) );
  MUX21X2_HVT U30 ( .A1(n386), .A2(n376), .S0(n304), .Y(n536) );
  INVX2_HVT U31 ( .A(in[1]), .Y(n262) );
  MUX21X1_HVT U32 ( .A1(n305), .A2(n386), .S0(n328), .Y(n573) );
  MUX21X2_HVT U34 ( .A1(n486), .A2(n483), .S0(n219), .Y(n482) );
  IBUFFX16_HVT U36 ( .A(n301), .Y(n219) );
  MUX21X2_HVT U37 ( .A1(n322), .A2(n315), .S0(n326), .Y(n576) );
  NAND2X0_HVT U38 ( .A1(n442), .A2(n224), .Y(n226) );
  NAND2X0_HVT U39 ( .A1(n430), .A2(n256), .Y(n227) );
  IBUFFX2_HVT U40 ( .A(n256), .Y(n224) );
  INVX0_HVT U41 ( .A(in[6]), .Y(n256) );
  MUX21X2_HVT U43 ( .A1(n484), .A2(n485), .S0(n303), .Y(n483) );
  INVX1_HVT U44 ( .A(n573), .Y(n362) );
  MUX21X2_HVT U45 ( .A1(n576), .A2(n493), .S0(n294), .Y(n491) );
  OA21X1_HVT U46 ( .A1(n290), .A2(n333), .A3(n576), .Y(n432) );
  MUX41X1_HVT U47 ( .A1(n523), .A3(n520), .A2(n522), .A4(n518), .S0(n231), 
        .S1(n232), .Y(n517) );
  IBUFFX16_HVT U48 ( .A(n312), .Y(n231) );
  IBUFFX16_HVT U49 ( .A(n300), .Y(n232) );
  IBUFFX2_HVT U50 ( .A(n578), .Y(n357) );
  MUX21X2_HVT U51 ( .A1(n578), .A2(n340), .S0(n304), .Y(n458) );
  INVX2_HVT U52 ( .A(n333), .Y(n330) );
  INVX4_HVT U54 ( .A(n235), .Y(n333) );
  INVX1_HVT U55 ( .A(in[1]), .Y(n263) );
  INVX2_HVT U60 ( .A(n328), .Y(n326) );
  NAND2X2_HVT U64 ( .A1(n257), .A2(n258), .Y(out[1]) );
  INVX2_HVT U65 ( .A(n332), .Y(n233) );
  IBUFFX2_HVT U67 ( .A(n334), .Y(n332) );
  INVX0_HVT U70 ( .A(in[7]), .Y(n234) );
  INVX1_HVT U71 ( .A(n234), .Y(n235) );
  NBUFFX2_HVT U72 ( .A(n332), .Y(n304) );
  INVX0_HVT U76 ( .A(n328), .Y(n236) );
  INVX1_HVT U79 ( .A(in[1]), .Y(n328) );
  MUX21X2_HVT U81 ( .A1(n462), .A2(n454), .S0(n237), .Y(out[4]) );
  IBUFFX16_HVT U82 ( .A(in[6]), .Y(n237) );
  NBUFFX4_HVT U84 ( .A(n235), .Y(n238) );
  MUX41X1_HVT U86 ( .A1(n519), .A3(n377), .A2(n285), .A4(n289), .S0(n239), 
        .S1(n238), .Y(n518) );
  IBUFFX16_HVT U87 ( .A(n293), .Y(n239) );
  MUX41X1_HVT U88 ( .A1(n474), .A3(n488), .A2(n469), .A4(n482), .S0(n240), 
        .S1(n274), .Y(out[3]) );
  IBUFFX16_HVT U89 ( .A(n256), .Y(n240) );
  MUX21X1_HVT U90 ( .A1(n305), .A2(n310), .S0(n263), .Y(n481) );
  MUX21X1_HVT U91 ( .A1(n242), .A2(n574), .S0(n243), .Y(n241) );
  IBUFFX16_HVT U92 ( .A(n241), .Y(n480) );
  IBUFFX16_HVT U94 ( .A(n481), .Y(n242) );
  IBUFFX16_HVT U95 ( .A(n295), .Y(n243) );
  INVX2_HVT U98 ( .A(n334), .Y(n331) );
  NBUFFX2_HVT U99 ( .A(n388), .Y(n309) );
  MUX21X1_HVT U100 ( .A1(n311), .A2(n383), .S0(n327), .Y(n578) );
  NBUFFX2_HVT U102 ( .A(n268), .Y(n308) );
  NBUFFX2_HVT U104 ( .A(in[5]), .Y(n301) );
  INVX0_HVT U107 ( .A(n310), .Y(n247) );
  MUX21X1_HVT U108 ( .A1(n308), .A2(n313), .S0(n327), .Y(n584) );
  MUX21X1_HVT U109 ( .A1(n319), .A2(n322), .S0(n252), .Y(n251) );
  MUX21X1_HVT U111 ( .A1(n305), .A2(n387), .S0(n326), .Y(n567) );
  MUX21X1_HVT U112 ( .A1(n246), .A2(n316), .S0(n303), .Y(n468) );
  NAND2X0_HVT U113 ( .A1(n253), .A2(n254), .Y(out[2]) );
  INVX0_HVT U114 ( .A(n259), .Y(n570) );
  MUX21X1_HVT U116 ( .A1(n318), .A2(n316), .S0(n326), .Y(n516) );
  INVX0_HVT U117 ( .A(n255), .Y(n569) );
  NAND2X0_HVT U118 ( .A1(n479), .A2(n302), .Y(n265) );
  INVX1_HVT U119 ( .A(n269), .Y(n329) );
  MUX21X1_HVT U120 ( .A1(n261), .A2(n384), .S0(n303), .Y(n453) );
  MUX21X1_HVT U121 ( .A1(n359), .A2(n468), .S0(n297), .Y(n467) );
  OR2X1_HVT U122 ( .A1(n264), .A2(n268), .Y(n244) );
  INVX0_HVT U124 ( .A(n600), .Y(n273) );
  INVX1_HVT U126 ( .A(n312), .Y(n274) );
  INVX1_HVT U127 ( .A(n262), .Y(n252) );
  INVX1_HVT U128 ( .A(in[3]), .Y(n385) );
  INVX0_HVT U129 ( .A(n298), .Y(n269) );
  NBUFFX2_HVT U130 ( .A(in[2]), .Y(n293) );
  INVX0_HVT U132 ( .A(n294), .Y(n275) );
  INVX1_HVT U133 ( .A(in[5]), .Y(n277) );
  INVX1_HVT U134 ( .A(n303), .Y(n270) );
  INVX1_HVT U135 ( .A(n309), .Y(n245) );
  MUX21X2_HVT U137 ( .A1(n452), .A2(n453), .S0(n298), .Y(n450) );
  MUX21X1_HVT U138 ( .A1(n247), .A2(n317), .S0(n262), .Y(n246) );
  INVX1_HVT U142 ( .A(n318), .Y(n260) );
  INVX1_HVT U143 ( .A(n251), .Y(n580) );
  NAND2X0_HVT U145 ( .A1(n284), .A2(n302), .Y(n248) );
  NAND2X0_HVT U147 ( .A1(n590), .A2(n270), .Y(n249) );
  NAND2X0_HVT U148 ( .A1(n248), .A2(n249), .Y(n405) );
  MUX21X1_HVT U149 ( .A1(n305), .A2(n307), .S0(n263), .Y(n590) );
  INVX0_HVT U150 ( .A(n590), .Y(n348) );
  MUX21X2_HVT U152 ( .A1(n386), .A2(n308), .S0(n328), .Y(n598) );
  INVX0_HVT U153 ( .A(n306), .Y(n250) );
  IBUFFX2_HVT U155 ( .A(n268), .Y(n599) );
  INVX1_HVT U156 ( .A(n319), .Y(n387) );
  XNOR2X1_HVT U157 ( .A1(n599), .A2(n262), .Y(n561) );
  MUX41X1_HVT U161 ( .A1(n561), .A3(n374), .A2(n565), .A4(n516), .S0(n238), 
        .S1(n294), .Y(n515) );
  NAND2X0_HVT U164 ( .A1(n496), .A2(n256), .Y(n253) );
  NAND2X0_HVT U169 ( .A1(n506), .A2(in[6]), .Y(n254) );
  MUX21X1_HVT U170 ( .A1(n552), .A2(n556), .S0(n297), .Y(n551) );
  MUX21X2_HVT U171 ( .A1(n546), .A2(n548), .S0(n296), .Y(n545) );
  MUX21X1_HVT U172 ( .A1(n317), .A2(n322), .S0(n328), .Y(n255) );
  MUX41X1_HVT U173 ( .A1(n403), .A3(n402), .A2(n401), .A4(n400), .S0(n277), 
        .S1(n274), .Y(n399) );
  MUX21X2_HVT U174 ( .A1(n423), .A2(n414), .S0(n256), .Y(out[6]) );
  INVX1_HVT U175 ( .A(n582), .Y(n354) );
  MUX21X1_HVT U183 ( .A1(n569), .A2(n378), .S0(n302), .Y(n446) );
  MUX21X1_HVT U185 ( .A1(n387), .A2(n599), .S0(n262), .Y(n582) );
  NAND2X0_HVT U186 ( .A1(n517), .A2(n256), .Y(n257) );
  NAND2X0_HVT U187 ( .A1(n527), .A2(in[6]), .Y(n258) );
  MUX21X1_HVT U188 ( .A1(n268), .A2(n260), .S0(n328), .Y(n259) );
  MUX41X1_HVT U190 ( .A1(n422), .A3(n419), .A2(n418), .A4(n415), .S0(n277), 
        .S1(n274), .Y(n414) );
  MUX41X1_HVT U191 ( .A1(n410), .A3(n412), .A2(n407), .A4(n411), .S0(in[0]), 
        .S1(n277), .Y(n406) );
  XOR2X2_HVT U192 ( .A1(n270), .A2(n580), .Y(n563) );
  NBUFFX4_HVT U196 ( .A(n388), .Y(n311) );
  MUX21X1_HVT U198 ( .A1(n268), .A2(n313), .S0(n263), .Y(n261) );
  MUX41X1_HVT U199 ( .A1(n576), .A3(n354), .A2(n487), .A4(n593), .S0(n275), 
        .S1(n233), .Y(n486) );
  MUX41X1_HVT U200 ( .A1(n561), .A3(n532), .A2(n568), .A4(n287), .S0(n275), 
        .S1(n270), .Y(n418) );
  MUX41X1_HVT U202 ( .A1(n353), .A3(n590), .A2(n250), .A4(n521), .S0(n238), 
        .S1(n293), .Y(n520) );
  MUX21X1_HVT U206 ( .A1(n311), .A2(n305), .S0(n264), .Y(n413) );
  INVX1_HVT U207 ( .A(n252), .Y(n264) );
  INVX1_HVT U209 ( .A(n394), .Y(n376) );
  NAND2X0_HVT U210 ( .A1(n480), .A2(n270), .Y(n266) );
  NAND2X0_HVT U211 ( .A1(n265), .A2(n266), .Y(n476) );
  MUX21X2_HVT U213 ( .A1(n476), .A2(n475), .S0(n277), .Y(n474) );
  MUX41X1_HVT U216 ( .A1(n314), .A3(n370), .A2(n306), .A4(n353), .S0(n275), 
        .S1(n233), .Y(n459) );
  INVX1_HVT U217 ( .A(n271), .Y(n466) );
  MUX41X1_HVT U219 ( .A1(n456), .A3(n460), .A2(n455), .A4(n459), .S0(in[0]), 
        .S1(n277), .Y(n454) );
  MUX21X2_HVT U221 ( .A1(n446), .A2(n447), .S0(n298), .Y(n445) );
  MUX41X1_HVT U222 ( .A1(n592), .A3(n336), .A2(n352), .A4(n562), .S0(n269), 
        .S1(n333), .Y(n522) );
  MUX41X1_HVT U223 ( .A1(n508), .A3(n515), .A2(n507), .A4(n510), .S0(n312), 
        .S1(n277), .Y(n506) );
  AO21X2_HVT U224 ( .A1(n263), .A2(n384), .A3(n333), .Y(n502) );
  MUX21X1_HVT U225 ( .A1(n268), .A2(n314), .S0(n325), .Y(n267) );
  XNOR2X2_HVT U226 ( .A1(n309), .A2(in[3]), .Y(n268) );
  INVX0_HVT U227 ( .A(n267), .Y(n272) );
  NBUFFX2_HVT U228 ( .A(n268), .Y(n307) );
  MUX41X1_HVT U229 ( .A1(n251), .A3(n273), .A2(n314), .A4(n272), .S0(n275), 
        .S1(n233), .Y(n271) );
  MUX41X1_HVT U230 ( .A1(n337), .A3(n319), .A2(n288), .A4(n493), .S0(n275), 
        .S1(n333), .Y(n449) );
  NBUFFX2_HVT U231 ( .A(n330), .Y(n276) );
  MUX41X1_HVT U232 ( .A1(n439), .A3(n434), .A2(n437), .A4(n431), .S0(n274), 
        .S1(n277), .Y(n430) );
  INVX0_HVT U233 ( .A(n295), .Y(n280) );
  OA21X1_HVT U234 ( .A1(n259), .A2(n275), .A3(n350), .Y(n494) );
  NAND2X0_HVT U235 ( .A1(n490), .A2(n281), .Y(n282) );
  NAND2X0_HVT U236 ( .A1(n406), .A2(in[6]), .Y(n278) );
  NAND2X0_HVT U237 ( .A1(n399), .A2(n256), .Y(n279) );
  NAND2X0_HVT U238 ( .A1(n278), .A2(n279), .Y(out[7]) );
  AND3X2_HVT U239 ( .A1(n297), .A2(n264), .A3(n245), .Y(n472) );
  AO21X2_HVT U240 ( .A1(n298), .A2(n314), .A3(n250), .Y(n484) );
  MUX21X2_HVT U241 ( .A1(n404), .A2(n405), .S0(n296), .Y(n403) );
  MUX41X1_HVT U242 ( .A1(n561), .A3(n372), .A2(n532), .A4(n380), .S0(n280), 
        .S1(n233), .Y(n455) );
  MUX41X1_HVT U243 ( .A1(n352), .A3(n351), .A2(n335), .A4(n374), .S0(n233), 
        .S1(n277), .Y(n556) );
  INVX1_HVT U244 ( .A(n558), .Y(n281) );
  XOR2X1_HVT U245 ( .A1(n280), .A2(n233), .Y(n560) );
  MUX41X1_HVT U246 ( .A1(n489), .A3(n491), .A2(n495), .A4(n494), .S0(n238), 
        .S1(n301), .Y(n488) );
  NAND2X0_HVT U247 ( .A1(n321), .A2(n558), .Y(n283) );
  NAND2X0_HVT U248 ( .A1(n282), .A2(n283), .Y(n489) );
  XOR2X1_HVT U249 ( .A1(n324), .A2(n296), .Y(n558) );
  NBUFFX2_HVT U250 ( .A(n332), .Y(n302) );
  XNOR2X1_HVT U251 ( .A1(n333), .A2(n324), .Y(n291) );
  MUX21X2_HVT U252 ( .A1(n367), .A2(n381), .S0(n303), .Y(n409) );
  MUX21X2_HVT U253 ( .A1(n542), .A2(n544), .S0(n296), .Y(n541) );
  MUX21X2_HVT U254 ( .A1(n288), .A2(n505), .S0(n560), .Y(n504) );
  MUX21X2_HVT U255 ( .A1(n360), .A2(n592), .S0(n298), .Y(n505) );
  INVX1_HVT U256 ( .A(n317), .Y(n383) );
  MUX21X1_HVT U257 ( .A1(n286), .A2(n348), .S0(n294), .Y(n471) );
  NBUFFX2_HVT U258 ( .A(n268), .Y(n306) );
  AND2X1_HVT U259 ( .A1(n308), .A2(n549), .Y(n284) );
  NBUFFX2_HVT U260 ( .A(n601), .Y(n317) );
  MUX21X1_HVT U261 ( .A1(n383), .A2(n386), .S0(n301), .Y(n553) );
  NBUFFX2_HVT U262 ( .A(n601), .Y(n318) );
  MUX21X1_HVT U263 ( .A1(n344), .A2(n384), .S0(n301), .Y(n538) );
  AND2X1_HVT U264 ( .A1(n320), .A2(n532), .Y(n285) );
  MUX21X1_HVT U265 ( .A1(n320), .A2(n307), .S0(n326), .Y(n566) );
  MUX21X1_HVT U266 ( .A1(n306), .A2(n311), .S0(n325), .Y(n501) );
  MUX21X1_HVT U267 ( .A1(n383), .A2(n387), .S0(n326), .Y(n429) );
  MUX21X1_HVT U268 ( .A1(n386), .A2(n307), .S0(n325), .Y(n441) );
  MUX21X1_HVT U269 ( .A1(n307), .A2(n383), .S0(n325), .Y(n509) );
  MUX21X1_HVT U270 ( .A1(n599), .A2(n311), .S0(n326), .Y(n529) );
  MUX21X1_HVT U271 ( .A1(n337), .A2(n362), .S0(n294), .Y(n485) );
  NAND2X0_HVT U272 ( .A1(n309), .A2(n385), .Y(n601) );
  NBUFFX2_HVT U273 ( .A(n604), .Y(n319) );
  INVX1_HVT U274 ( .A(n322), .Y(n386) );
  NBUFFX2_HVT U275 ( .A(n604), .Y(n320) );
  XOR2X1_HVT U276 ( .A1(n324), .A2(n384), .Y(n562) );
  MUX21X1_HVT U277 ( .A1(n385), .A2(n323), .S0(n325), .Y(n416) );
  MUX21X1_HVT U278 ( .A1(n322), .A2(n320), .S0(n325), .Y(n417) );
  MUX21X1_HVT U279 ( .A1(n384), .A2(n383), .S0(n327), .Y(n588) );
  INVX1_HVT U280 ( .A(n314), .Y(n384) );
  MUX21X1_HVT U281 ( .A1(n321), .A2(n315), .S0(n327), .Y(n592) );
  MUX21X1_HVT U282 ( .A1(n317), .A2(n323), .S0(n324), .Y(n511) );
  MUX21X1_HVT U283 ( .A1(n305), .A2(n386), .S0(n327), .Y(n595) );
  NBUFFX2_HVT U284 ( .A(n604), .Y(n321) );
  XOR2X1_HVT U285 ( .A1(n319), .A2(n324), .Y(n557) );
  MUX21X1_HVT U286 ( .A1(n319), .A2(n310), .S0(n325), .Y(n396) );
  XNOR2X1_HVT U287 ( .A1(n317), .A2(n324), .Y(n286) );
  AND2X1_HVT U288 ( .A1(n252), .A2(n387), .Y(n287) );
  MUX21X1_HVT U289 ( .A1(n318), .A2(n305), .S0(n327), .Y(n594) );
  AND2X1_HVT U290 ( .A1(n323), .A2(n492), .Y(n288) );
  MUX21X1_HVT U291 ( .A1(n319), .A2(n318), .S0(n324), .Y(n391) );
  XNOR2X1_HVT U292 ( .A1(n322), .A2(n324), .Y(n289) );
  MUX21X1_HVT U293 ( .A1(n316), .A2(n310), .S0(n326), .Y(n534) );
  MUX21X1_HVT U294 ( .A1(n316), .A2(n323), .S0(n297), .Y(n478) );
  XOR2X1_HVT U295 ( .A1(n309), .A2(n324), .Y(n581) );
  NBUFFX2_HVT U296 ( .A(n332), .Y(n303) );
  NBUFFX2_HVT U297 ( .A(n385), .Y(n305) );
  NBUFFX2_HVT U298 ( .A(in[2]), .Y(n294) );
  NBUFFX2_HVT U299 ( .A(in[2]), .Y(n295) );
  NBUFFX2_HVT U300 ( .A(in[5]), .Y(n300) );
  NBUFFX2_HVT U301 ( .A(in[2]), .Y(n297) );
  NBUFFX2_HVT U302 ( .A(in[2]), .Y(n298) );
  NBUFFX2_HVT U303 ( .A(in[2]), .Y(n296) );
  NBUFFX2_HVT U304 ( .A(in[5]), .Y(n299) );
  MUX21X1_HVT U305 ( .A1(n503), .A2(n359), .S0(n297), .Y(n500) );
  MUX21X1_HVT U306 ( .A1(n420), .A2(n421), .S0(n296), .Y(n419) );
  MUX21X1_HVT U307 ( .A1(n519), .A2(n313), .S0(n303), .Y(n421) );
  XOR2X1_HVT U308 ( .A1(n324), .A2(in[3]), .Y(n559) );
  MUX21X1_HVT U309 ( .A1(n315), .A2(n308), .S0(n326), .Y(n498) );
  MUX21X1_HVT U310 ( .A1(n526), .A2(n525), .S0(n298), .Y(n523) );
  MUX21X1_HVT U311 ( .A1(n433), .A2(n432), .S0(n297), .Y(n431) );
  MUX21X1_HVT U312 ( .A1(n316), .A2(n376), .S0(n304), .Y(n433) );
  MUX21X1_HVT U313 ( .A1(n384), .A2(n387), .S0(n325), .Y(n438) );
  AND2X1_HVT U314 ( .A1(n308), .A2(n264), .Y(n290) );
  MUX21X1_HVT U315 ( .A1(n313), .A2(n383), .S0(n326), .Y(n568) );
  MUX21X1_HVT U316 ( .A1(n448), .A2(n321), .S0(n291), .Y(n447) );
  MUX21X1_HVT U317 ( .A1(n589), .A2(n361), .S0(n295), .Y(n470) );
  NAND2X0_HVT U318 ( .A1(in[3]), .A2(n311), .Y(n604) );
  NBUFFX2_HVT U319 ( .A(n605), .Y(n322) );
  MUX21X1_HVT U320 ( .A1(n387), .A2(n313), .S0(n327), .Y(n587) );
  MUX21X1_HVT U321 ( .A1(n363), .A2(n603), .S0(n295), .Y(n495) );
  MUX21X1_HVT U322 ( .A1(n554), .A2(n555), .S0(n302), .Y(n552) );
  MUX21X1_HVT U323 ( .A1(n313), .A2(n572), .S0(n301), .Y(n555) );
  XOR2X1_HVT U324 ( .A1(n324), .A2(n300), .Y(n564) );
  MUX21X1_HVT U325 ( .A1(n603), .A2(n262), .S0(n296), .Y(n477) );
  NBUFFX2_HVT U326 ( .A(n596), .Y(n314) );
  MUX21X1_HVT U327 ( .A1(n313), .A2(n384), .S0(n325), .Y(n393) );
  MUX21X1_HVT U328 ( .A1(n577), .A2(n397), .S0(n302), .Y(n392) );
  MUX21X1_HVT U329 ( .A1(n318), .A2(n313), .S0(n327), .Y(n597) );
  MUX21X1_HVT U330 ( .A1(n346), .A2(n263), .S0(n301), .Y(n540) );
  NBUFFX2_HVT U331 ( .A(n596), .Y(n315) );
  MUX21X1_HVT U332 ( .A1(n356), .A2(n577), .S0(n295), .Y(n473) );
  MUX21X1_HVT U333 ( .A1(n321), .A2(n514), .S0(n291), .Y(n513) );
  MUX21X1_HVT U334 ( .A1(n313), .A2(n310), .S0(n304), .Y(n514) );
  NBUFFX2_HVT U335 ( .A(n605), .Y(n323) );
  NBUFFX2_HVT U336 ( .A(n388), .Y(n310) );
  NBUFFX2_HVT U337 ( .A(n596), .Y(n316) );
  AND2X1_HVT U338 ( .A1(n305), .A2(n264), .Y(n292) );
  MUX21X1_HVT U339 ( .A1(n409), .A2(n408), .S0(n296), .Y(n407) );
  INVX0_HVT U340 ( .A(in[4]), .Y(n388) );
  MUX21X1_HVT U341 ( .A1(n383), .A2(n245), .S0(n326), .Y(n575) );
  NAND2X0_HVT U342 ( .A1(in[3]), .A2(in[4]), .Y(n605) );
  MUX21X1_HVT U343 ( .A1(n245), .A2(n599), .S0(n325), .Y(n395) );
  MUX21X1_HVT U344 ( .A1(n245), .A2(n386), .S0(n326), .Y(n571) );
  MUX21X1_HVT U345 ( .A1(n245), .A2(n384), .S0(n327), .Y(n589) );
  NAND2X0_HVT U346 ( .A1(in[4]), .A2(n385), .Y(n596) );
  MUX21X1_HVT U347 ( .A1(n245), .A2(n321), .S0(n327), .Y(n586) );
  MUX21X1_HVT U348 ( .A1(n323), .A2(n245), .S0(n327), .Y(n579) );
  MUX21X1_HVT U349 ( .A1(n313), .A2(n245), .S0(n294), .Y(n490) );
  MUX21X1_HVT U350 ( .A1(n245), .A2(n315), .S0(n325), .Y(n390) );
  MUX21X1_HVT U351 ( .A1(n245), .A2(n323), .S0(n326), .Y(n389) );
  MUX21X1_HVT U352 ( .A1(n305), .A2(n245), .S0(n327), .Y(n577) );
  NBUFFX2_HVT U353 ( .A(in[3]), .Y(n313) );
  NBUFFX2_HVT U354 ( .A(in[0]), .Y(n312) );
  INVX0_HVT U355 ( .A(n585), .Y(n335) );
  INVX0_HVT U356 ( .A(n583), .Y(n336) );
  INVX0_HVT U357 ( .A(n572), .Y(n337) );
  INVX0_HVT U358 ( .A(n435), .Y(n338) );
  INVX0_HVT U359 ( .A(n398), .Y(n339) );
  INVX0_HVT U360 ( .A(n603), .Y(n340) );
  INVX0_HVT U361 ( .A(n591), .Y(n341) );
  INVX0_HVT U362 ( .A(n602), .Y(n342) );
  INVX0_HVT U363 ( .A(n598), .Y(n343) );
  INVX0_HVT U364 ( .A(n597), .Y(n344) );
  INVX0_HVT U365 ( .A(n595), .Y(n345) );
  INVX0_HVT U366 ( .A(n594), .Y(n346) );
  INVX0_HVT U367 ( .A(n592), .Y(n347) );
  INVX0_HVT U368 ( .A(n589), .Y(n349) );
  INVX0_HVT U369 ( .A(n588), .Y(n350) );
  INVX0_HVT U370 ( .A(n587), .Y(n351) );
  INVX0_HVT U371 ( .A(n586), .Y(n352) );
  INVX0_HVT U372 ( .A(n581), .Y(n355) );
  INVX0_HVT U373 ( .A(n579), .Y(n356) );
  INVX0_HVT U374 ( .A(n577), .Y(n358) );
  INVX0_HVT U375 ( .A(n392), .Y(n359) );
  INVX0_HVT U376 ( .A(n576), .Y(n360) );
  INVX0_HVT U377 ( .A(n575), .Y(n361) );
  INVX0_HVT U378 ( .A(n571), .Y(n363) );
  INVX0_HVT U379 ( .A(n568), .Y(n364) );
  INVX0_HVT U380 ( .A(n567), .Y(n365) );
  INVX0_HVT U381 ( .A(n566), .Y(n366) );
  INVX0_HVT U382 ( .A(n565), .Y(n367) );
  INVX0_HVT U383 ( .A(n532), .Y(n368) );
  INVX0_HVT U384 ( .A(n593), .Y(n369) );
  INVX0_HVT U385 ( .A(n492), .Y(n370) );
  INVX0_HVT U386 ( .A(n397), .Y(n371) );
  INVX0_HVT U387 ( .A(n549), .Y(n372) );
  INVX0_HVT U388 ( .A(n451), .Y(n373) );
  INVX0_HVT U389 ( .A(n396), .Y(n374) );
  INVX0_HVT U390 ( .A(n395), .Y(n375) );
  INVX0_HVT U391 ( .A(n393), .Y(n377) );
  INVX0_HVT U392 ( .A(n511), .Y(n378) );
  INVX0_HVT U393 ( .A(n501), .Y(n379) );
  INVX0_HVT U394 ( .A(n391), .Y(n380) );
  INVX0_HVT U395 ( .A(n390), .Y(n381) );
  INVX0_HVT U396 ( .A(n389), .Y(n382) );
endmodule

