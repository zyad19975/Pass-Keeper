
module Mix_Column ( in, out );
  input [127:0] in;
  output [127:0] out;
  wire   n16, n17, n19, n21, n22, n23, n24, n26, n27, n28, n29, n30, n31, n34,
         n35, n36, n38, n39, n40, n42, n43, n44, n46, n47, n48, n50, n51, n53,
         n55, n56, n57, n58, n60, n61, n63, n64, n65, n66, n67, n69, n71, n72,
         n74, n75, n78, n79, n80, n81, n82, n86, n87, n88, n89, n90, n93, n94,
         n95, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n110, n111, n114, n115, n117, n118, n119, n121, n122, n123, n124,
         n126, n127, n129, n130, n131, n133, n134, n135, n137, n138, n140,
         n141, n145, n146, n147, n148, n149, n150, n151, n152, n154, n157,
         n158, n159, n160, n161, n162, n163, n166, n169, n176, n177, n178,
         n179, n180, n181, n182, n184, n185, n187, n188, n189, n190, n193,
         n194, n197, n198, n199, n200, n201, n202, n209, n210, n213, n216,
         n218, n220, n221, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n18, n20, n32, n33, n37, n41, n45, n49, n52, n54, n59,
         n62, n68, n70, n73, n76, n77, n83, n84, n85, n91, n92, n96, n107,
         n109, n112, n113, n116, n120, n125, n128, n132, n136, n139, n142,
         n143, n144, n153, n155, n156, n164, n165, n167, n168, n170, n171,
         n172, n173, n174, n175, n183, n186, n191, n192, n195, n196, n203,
         n204, n205, n206, n207, n208, n211, n212, n214, n215, n217, n219,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587;

  XOR3X2_HVT U129 ( .A1(n178), .A2(n388), .A3(n179), .Y(out[126]) );
  XNOR3X1_HVT U225 ( .A1(n570), .A2(in[67]), .A3(n499), .Y(n69) );
  XOR2X2_HVT U1 ( .A1(in[28]), .A2(n480), .Y(n95) );
  XOR3X2_HVT U2 ( .A1(n154), .A2(n10), .A3(n394), .Y(out[13]) );
  IBUFFX2_HVT U3 ( .A(in[69]), .Y(n290) );
  XOR3X1_HVT U4 ( .A1(n113), .A2(n509), .A3(n538), .Y(n134) );
  XNOR2X2_HVT U5 ( .A1(n552), .A2(n561), .Y(n538) );
  XOR2X2_HVT U6 ( .A1(in[100]), .A2(in[108]), .Y(n184) );
  INVX2_HVT U7 ( .A(in[103]), .Y(n456) );
  XOR2X2_HVT U8 ( .A1(n356), .A2(n560), .Y(n157) );
  XOR2X2_HVT U9 ( .A1(in[76]), .A2(in[68]), .Y(n35) );
  XOR3X2_HVT U10 ( .A1(n547), .A2(in[83]), .A3(n35), .Y(n34) );
  XNOR2X2_HVT U11 ( .A1(n232), .A2(in[120]), .Y(n414) );
  INVX2_HVT U12 ( .A(n535), .Y(n401) );
  XOR2X1_HVT U13 ( .A1(in[126]), .A2(n576), .Y(n218) );
  XNOR2X2_HVT U14 ( .A1(in[88]), .A2(n582), .Y(n466) );
  INVX2_HVT U15 ( .A(n456), .Y(n457) );
  NBUFFX2_HVT U16 ( .A(n150), .Y(n1) );
  XOR2X2_HVT U17 ( .A1(in[99]), .A2(n578), .Y(n187) );
  XOR2X2_HVT U18 ( .A1(in[44]), .A2(in[52]), .Y(n108) );
  XOR2X2_HVT U19 ( .A1(in[52]), .A2(in[60]), .Y(n90) );
  XOR2X2_HVT U20 ( .A1(in[89]), .A2(in[65]), .Y(n58) );
  NAND2X0_HVT U21 ( .A1(n324), .A2(n325), .Y(n2) );
  XOR3X2_HVT U22 ( .A1(n84), .A2(n508), .A3(n85), .Y(n213) );
  INVX1_HVT U23 ( .A(n109), .Y(n84) );
  XNOR2X2_HVT U24 ( .A1(in[73]), .A2(in[65]), .Y(n44) );
  INVX1_HVT U25 ( .A(n28), .Y(n374) );
  XOR3X2_HVT U26 ( .A1(n42), .A2(n3), .A3(n368), .Y(out[8]) );
  IBUFFX16_HVT U27 ( .A(n530), .Y(n3) );
  IBUFFX2_HVT U28 ( .A(in[75]), .Y(n45) );
  XOR2X2_HVT U29 ( .A1(n573), .A2(n41), .Y(n46) );
  INVX1_HVT U30 ( .A(n259), .Y(n41) );
  XNOR2X2_HVT U31 ( .A1(n4), .A2(n5), .Y(n194) );
  XOR2X2_HVT U32 ( .A1(n551), .A2(n356), .Y(n4) );
  XNOR2X2_HVT U33 ( .A1(n509), .A2(in[27]), .Y(n5) );
  XOR3X2_HVT U34 ( .A1(n553), .A2(n480), .A3(n6), .Y(n248) );
  IBUFFX16_HVT U35 ( .A(n427), .Y(n6) );
  XOR2X2_HVT U36 ( .A1(in[21]), .A2(in[30]), .Y(n404) );
  INVX2_HVT U37 ( .A(in[2]), .Y(n509) );
  XOR3X2_HVT U38 ( .A1(n543), .A2(in[27]), .A3(n118), .Y(n117) );
  XNOR2X2_HVT U39 ( .A1(n32), .A2(in[6]), .Y(n147) );
  INVX2_HVT U40 ( .A(in[14]), .Y(n32) );
  XOR2X2_HVT U41 ( .A1(n519), .A2(n556), .Y(n328) );
  XOR3X2_HVT U42 ( .A1(n530), .A2(n379), .A3(n151), .Y(n176) );
  IBUFFX2_HVT U43 ( .A(in[1]), .Y(n454) );
  INVX1_HVT U44 ( .A(n280), .Y(n292) );
  XOR3X2_HVT U45 ( .A1(n542), .A2(in[3]), .A3(n7), .Y(n255) );
  IBUFFX16_HVT U46 ( .A(n562), .Y(n7) );
  INVX2_HVT U47 ( .A(n552), .Y(n542) );
  XOR3X2_HVT U48 ( .A1(n147), .A2(n142), .A3(n63), .Y(out[15]) );
  XNOR2X2_HVT U49 ( .A1(n9), .A2(n8), .Y(n66) );
  IBUFFX16_HVT U50 ( .A(n455), .Y(n8) );
  NAND2X0_HVT U51 ( .A1(n281), .A2(n282), .Y(n9) );
  NBUFFX2_HVT U52 ( .A(in[5]), .Y(n10) );
  XOR2X2_HVT U53 ( .A1(n360), .A2(in[126]), .Y(n198) );
  INVX1_HVT U54 ( .A(n66), .Y(n223) );
  XOR3X2_HVT U55 ( .A1(n48), .A2(n231), .A3(n374), .Y(out[87]) );
  XOR2X2_HVT U56 ( .A1(in[94]), .A2(in[86]), .Y(n65) );
  INVX1_HVT U57 ( .A(in[86]), .Y(n192) );
  INVX1_HVT U58 ( .A(n400), .Y(n168) );
  INVX0_HVT U59 ( .A(n94), .Y(n394) );
  XOR2X1_HVT U60 ( .A1(in[20]), .A2(in[12]), .Y(n118) );
  INVX1_HVT U61 ( .A(n228), .Y(n231) );
  XOR3X2_HVT U62 ( .A1(n162), .A2(n371), .A3(n163), .Y(out[24]) );
  INVX2_HVT U63 ( .A(n584), .Y(n513) );
  INVX2_HVT U64 ( .A(n424), .Y(n425) );
  XOR3X2_HVT U65 ( .A1(n159), .A2(n397), .A3(n161), .Y(out[25]) );
  INVX1_HVT U66 ( .A(in[27]), .Y(n537) );
  XOR2X2_HVT U67 ( .A1(in[28]), .A2(in[20]), .Y(n151) );
  XNOR2X2_HVT U68 ( .A1(in[3]), .A2(in[27]), .Y(n327) );
  INVX2_HVT U69 ( .A(n549), .Y(n550) );
  INVX1_HVT U70 ( .A(n514), .Y(n143) );
  XNOR2X1_HVT U71 ( .A1(in[56]), .A2(n536), .Y(n121) );
  XNOR2X1_HVT U72 ( .A1(in[61]), .A2(in[53]), .Y(n88) );
  INVX1_HVT U73 ( .A(n359), .Y(n360) );
  XOR2X1_HVT U74 ( .A1(in[121]), .A2(in[113]), .Y(n189) );
  OR2X1_HVT U75 ( .A1(n36), .A2(n315), .Y(n288) );
  XOR3X2_HVT U76 ( .A1(n372), .A2(n316), .A3(n38), .Y(n36) );
  INVX1_HVT U77 ( .A(n491), .Y(n492) );
  INVX0_HVT U78 ( .A(n442), .Y(n11) );
  INVX1_HVT U79 ( .A(in[104]), .Y(n442) );
  INVX2_HVT U80 ( .A(n570), .Y(n279) );
  INVX0_HVT U81 ( .A(n279), .Y(n52) );
  INVX1_HVT U82 ( .A(n458), .Y(n289) );
  INVX0_HVT U83 ( .A(n456), .Y(n458) );
  INVX0_HVT U84 ( .A(in[46]), .Y(n233) );
  IBUFFX2_HVT U85 ( .A(n210), .Y(n76) );
  XOR2X2_HVT U86 ( .A1(in[72]), .A2(n571), .Y(n61) );
  XOR2X2_HVT U87 ( .A1(in[94]), .A2(n571), .Y(n75) );
  XOR3X2_HVT U88 ( .A1(n12), .A2(n576), .A3(n23), .Y(out[104]) );
  XOR2X1_HVT U89 ( .A1(in[120]), .A2(n585), .Y(n12) );
  INVX1_HVT U90 ( .A(n512), .Y(n13) );
  INVX1_HVT U91 ( .A(in[82]), .Y(n512) );
  INVX1_HVT U92 ( .A(n210), .Y(n586) );
  NAND2X0_HVT U93 ( .A1(n334), .A2(n335), .Y(n14) );
  XOR3X2_HVT U94 ( .A1(n252), .A2(in[45]), .A3(n88), .Y(out[37]) );
  XOR2X1_HVT U95 ( .A1(in[97]), .A2(n336), .Y(n21) );
  INVX0_HVT U96 ( .A(in[77]), .Y(n460) );
  XOR2X1_HVT U97 ( .A1(in[33]), .A2(in[57]), .Y(n119) );
  XOR2X2_HVT U98 ( .A1(in[56]), .A2(in[48]), .Y(n420) );
  IBUFFX2_HVT U99 ( .A(n29), .Y(n54) );
  INVX0_HVT U100 ( .A(n204), .Y(n15) );
  XOR3X2_HVT U101 ( .A1(in[57]), .A2(n204), .A3(n361), .Y(n396) );
  XOR2X2_HVT U102 ( .A1(in[90]), .A2(in[82]), .Y(n71) );
  XNOR2X1_HVT U103 ( .A1(in[29]), .A2(in[5]), .Y(n504) );
  INVX1_HVT U104 ( .A(in[18]), .Y(n514) );
  INVX0_HVT U105 ( .A(in[127]), .Y(n18) );
  INVX1_HVT U106 ( .A(n18), .Y(n20) );
  XNOR2X2_HVT U107 ( .A1(n18), .A2(in[118]), .Y(n197) );
  INVX1_HVT U108 ( .A(n372), .Y(n496) );
  XOR3X1_HVT U109 ( .A1(n500), .A2(n381), .A3(n95), .Y(n418) );
  XOR3X2_HVT U110 ( .A1(n37), .A2(n32), .A3(n33), .Y(out[23]) );
  IBUFFX16_HVT U111 ( .A(n146), .Y(n33) );
  XOR2X1_HVT U112 ( .A1(in[22]), .A2(n561), .Y(n37) );
  INVX0_HVT U113 ( .A(n372), .Y(n373) );
  INVX1_HVT U114 ( .A(in[72]), .Y(n259) );
  INVX0_HVT U115 ( .A(n45), .Y(n49) );
  XOR3X2_HVT U116 ( .A1(n64), .A2(n52), .A3(n54), .Y(out[79]) );
  IBUFFX2_HVT U117 ( .A(n447), .Y(n109) );
  INVX0_HVT U118 ( .A(in[44]), .Y(n488) );
  INVX1_HVT U119 ( .A(n108), .Y(n521) );
  XOR3X2_HVT U120 ( .A1(n443), .A2(n442), .A3(n444), .Y(out[120]) );
  XOR2X2_HVT U121 ( .A1(n245), .A2(n579), .Y(n444) );
  XOR3X2_HVT U122 ( .A1(n59), .A2(n253), .A3(n62), .Y(n265) );
  IBUFFX16_HVT U123 ( .A(n447), .Y(n59) );
  XNOR2X1_HVT U124 ( .A1(n489), .A2(n579), .Y(n62) );
  XNOR2X2_HVT U125 ( .A1(n457), .A2(n575), .Y(n177) );
  XOR2X2_HVT U126 ( .A1(n395), .A2(n559), .Y(n163) );
  INVX0_HVT U127 ( .A(in[97]), .Y(n68) );
  INVX1_HVT U128 ( .A(n68), .Y(n70) );
  INVX0_HVT U130 ( .A(n429), .Y(n73) );
  XOR3X2_HVT U131 ( .A1(n180), .A2(n73), .A3(n76), .Y(out[110]) );
  INVX0_HVT U132 ( .A(n269), .Y(n77) );
  INVX0_HVT U133 ( .A(n77), .Y(n83) );
  INVX0_HVT U134 ( .A(in[20]), .Y(n453) );
  XOR2X1_HVT U135 ( .A1(in[99]), .A2(in[98]), .Y(n85) );
  XOR3X1_HVT U136 ( .A1(n100), .A2(n382), .A3(n131), .Y(out[41]) );
  INVX1_HVT U137 ( .A(n111), .Y(n252) );
  NAND2X0_HVT U138 ( .A1(n411), .A2(n412), .Y(n96) );
  NAND2X0_HVT U139 ( .A1(n91), .A2(n92), .Y(n107) );
  NAND2X0_HVT U140 ( .A1(n96), .A2(n107), .Y(out[27]) );
  INVX1_HVT U141 ( .A(n411), .Y(n91) );
  INVX0_HVT U142 ( .A(n412), .Y(n92) );
  INVX0_HVT U143 ( .A(in[9]), .Y(n284) );
  XNOR2X2_HVT U144 ( .A1(in[113]), .A2(in[105]), .Y(n24) );
  INVX0_HVT U145 ( .A(n537), .Y(n112) );
  INVX1_HVT U146 ( .A(n112), .Y(n113) );
  INVX1_HVT U147 ( .A(n507), .Y(n508) );
  XOR2X2_HVT U148 ( .A1(in[98]), .A2(in[106]), .Y(n188) );
  INVX0_HVT U149 ( .A(in[99]), .Y(n437) );
  INVX2_HVT U150 ( .A(in[19]), .Y(n549) );
  NBUFFX2_HVT U151 ( .A(in[113]), .Y(n116) );
  NAND2X0_HVT U152 ( .A1(n185), .A2(n125), .Y(n128) );
  NAND2X0_HVT U153 ( .A1(n120), .A2(n349), .Y(n132) );
  NAND2X0_HVT U154 ( .A1(n128), .A2(n132), .Y(out[123]) );
  INVX1_HVT U155 ( .A(n185), .Y(n120) );
  INVX0_HVT U156 ( .A(n349), .Y(n125) );
  XOR3X1_HVT U157 ( .A1(n493), .A2(n527), .A3(n187), .Y(n185) );
  XOR2X2_HVT U158 ( .A1(in[73]), .A2(in[81]), .Y(n57) );
  INVX2_HVT U159 ( .A(n464), .Y(n465) );
  XNOR2X1_HVT U160 ( .A1(in[114]), .A2(in[122]), .Y(n22) );
  INVX1_HVT U161 ( .A(n522), .Y(n498) );
  INVX1_HVT U162 ( .A(in[112]), .Y(n585) );
  INVX0_HVT U163 ( .A(n581), .Y(n371) );
  XNOR2X1_HVT U164 ( .A1(in[59]), .A2(n536), .Y(n114) );
  INVX1_HVT U165 ( .A(in[125]), .Y(n491) );
  XOR3X1_HVT U166 ( .A1(n487), .A2(n579), .A3(n437), .Y(n220) );
  INVX1_HVT U167 ( .A(n486), .Y(n487) );
  INVX1_HVT U168 ( .A(n533), .Y(n249) );
  INVX1_HVT U169 ( .A(n277), .Y(n278) );
  INVX1_HVT U170 ( .A(n258), .Y(n144) );
  INVX0_HVT U171 ( .A(in[38]), .Y(n405) );
  XOR3X1_HVT U172 ( .A1(n462), .A2(n460), .A3(n461), .Y(out[86]) );
  INVX0_HVT U173 ( .A(n22), .Y(n173) );
  INVX0_HVT U174 ( .A(n489), .Y(n172) );
  INVX1_HVT U175 ( .A(in[87]), .Y(n584) );
  INVX0_HVT U176 ( .A(n299), .Y(n283) );
  INVX1_HVT U177 ( .A(n122), .Y(n382) );
  INVX0_HVT U178 ( .A(n160), .Y(n397) );
  INVX1_HVT U179 ( .A(n553), .Y(n142) );
  INVX0_HVT U180 ( .A(n581), .Y(n402) );
  INVX0_HVT U181 ( .A(in[73]), .Y(n326) );
  INVX0_HVT U182 ( .A(in[39]), .Y(n398) );
  INVX1_HVT U183 ( .A(n572), .Y(n280) );
  INVX1_HVT U184 ( .A(in[26]), .Y(n535) );
  INVX1_HVT U185 ( .A(n290), .Y(n291) );
  INVX1_HVT U186 ( .A(n554), .Y(n530) );
  XOR2X2_HVT U187 ( .A1(n571), .A2(n496), .Y(n136) );
  INVX0_HVT U188 ( .A(n528), .Y(n347) );
  INVX1_HVT U189 ( .A(in[106]), .Y(n208) );
  INVX1_HVT U190 ( .A(in[105]), .Y(n274) );
  INVX1_HVT U191 ( .A(in[35]), .Y(n529) );
  INVX0_HVT U192 ( .A(n529), .Y(n322) );
  INVX1_HVT U193 ( .A(in[62]), .Y(n303) );
  XNOR2X1_HVT U194 ( .A1(in[92]), .A2(in[84]), .Y(n139) );
  XOR2X1_HVT U195 ( .A1(in[49]), .A2(in[57]), .Y(n100) );
  INVX1_HVT U196 ( .A(n101), .Y(n294) );
  INVX1_HVT U197 ( .A(in[6]), .Y(n470) );
  INVX1_HVT U198 ( .A(in[83]), .Y(n518) );
  INVX1_HVT U199 ( .A(n262), .Y(n494) );
  INVX1_HVT U200 ( .A(in[64]), .Y(n262) );
  INVX0_HVT U201 ( .A(in[67]), .Y(n331) );
  NBUFFX2_HVT U202 ( .A(in[39]), .Y(n563) );
  INVX1_HVT U203 ( .A(in[41]), .Y(n300) );
  INVX0_HVT U204 ( .A(n437), .Y(n348) );
  INVX1_HVT U205 ( .A(in[70]), .Y(n254) );
  INVX1_HVT U206 ( .A(in[48]), .Y(n332) );
  INVX1_HVT U207 ( .A(n90), .Y(n417) );
  INVX0_HVT U208 ( .A(in[54]), .Y(n205) );
  INVX0_HVT U209 ( .A(in[59]), .Y(n433) );
  INVX1_HVT U210 ( .A(in[87]), .Y(n372) );
  INVX0_HVT U211 ( .A(in[85]), .Y(n463) );
  INVX1_HVT U212 ( .A(n463), .Y(n362) );
  INVX0_HVT U213 ( .A(in[16]), .Y(n386) );
  XOR3X2_HVT U214 ( .A1(n271), .A2(n264), .A3(n482), .Y(n131) );
  IBUFFX2_HVT U215 ( .A(in[76]), .Y(n236) );
  IBUFFX2_HVT U216 ( .A(n147), .Y(n403) );
  XNOR2X1_HVT U217 ( .A1(n285), .A2(in[17]), .Y(n320) );
  NAND2X0_HVT U218 ( .A1(n258), .A2(n110), .Y(n155) );
  NAND2X0_HVT U219 ( .A1(n144), .A2(n153), .Y(n156) );
  NAND2X0_HVT U220 ( .A1(n155), .A2(n156), .Y(out[52]) );
  INVX1_HVT U221 ( .A(n110), .Y(n153) );
  INVX0_HVT U222 ( .A(in[17]), .Y(n422) );
  XOR3X1_HVT U223 ( .A1(n525), .A2(n565), .A3(n114), .Y(n501) );
  OR2X1_HVT U224 ( .A1(n423), .A2(in[61]), .Y(n234) );
  INVX1_HVT U226 ( .A(n361), .Y(n164) );
  INVX1_HVT U227 ( .A(in[56]), .Y(n361) );
  INVX0_HVT U228 ( .A(in[110]), .Y(n385) );
  XNOR2X2_HVT U229 ( .A1(n11), .A2(n577), .Y(n165) );
  XNOR2X2_HVT U230 ( .A1(n585), .A2(in[104]), .Y(n26) );
  INVX1_HVT U231 ( .A(in[75]), .Y(n455) );
  NAND2X0_HVT U232 ( .A1(n399), .A2(n400), .Y(n170) );
  NAND2X0_HVT U233 ( .A1(n167), .A2(n168), .Y(n171) );
  NAND2X0_HVT U234 ( .A1(n170), .A2(n171), .Y(out[19]) );
  INVX0_HVT U235 ( .A(n399), .Y(n167) );
  XNOR2X1_HVT U236 ( .A1(n328), .A2(n381), .Y(n400) );
  IBUFFX2_HVT U237 ( .A(in[109]), .Y(n440) );
  IBUFFX2_HVT U238 ( .A(in[8]), .Y(n270) );
  XOR3X2_HVT U239 ( .A1(n190), .A2(n172), .A3(n173), .Y(out[106]) );
  NAND2X0_HVT U240 ( .A1(n502), .A2(n501), .Y(n183) );
  NAND2X0_HVT U241 ( .A1(n174), .A2(n175), .Y(n186) );
  NAND2X0_HVT U242 ( .A1(n183), .A2(n186), .Y(out[51]) );
  INVX1_HVT U243 ( .A(n502), .Y(n174) );
  INVX0_HVT U244 ( .A(n501), .Y(n175) );
  NAND2X0_HVT U245 ( .A1(in[95]), .A2(n192), .Y(n195) );
  NAND2X0_HVT U246 ( .A1(n191), .A2(in[86]), .Y(n196) );
  NAND2X0_HVT U247 ( .A1(n195), .A2(n196), .Y(n48) );
  INVX1_HVT U248 ( .A(n573), .Y(n191) );
  XNOR2X2_HVT U249 ( .A1(n203), .A2(n127), .Y(out[43]) );
  XNOR2X2_HVT U250 ( .A1(n406), .A2(n529), .Y(n203) );
  INVX1_HVT U251 ( .A(in[107]), .Y(n256) );
  XOR3X2_HVT U252 ( .A1(n21), .A2(n193), .A3(n370), .Y(out[113]) );
  XOR2X1_HVT U253 ( .A1(in[108]), .A2(in[116]), .Y(n199) );
  INVX0_HVT U254 ( .A(in[108]), .Y(n449) );
  NAND2X0_HVT U255 ( .A1(n15), .A2(n205), .Y(n206) );
  NAND2X0_HVT U256 ( .A1(n204), .A2(in[54]), .Y(n207) );
  NAND2X0_HVT U257 ( .A1(n206), .A2(n207), .Y(n106) );
  INVX0_HVT U258 ( .A(in[63]), .Y(n204) );
  INVX0_HVT U259 ( .A(in[50]), .Y(n525) );
  XOR3X2_HVT U260 ( .A1(n35), .A2(n291), .A3(n428), .Y(out[77]) );
  XOR3X2_HVT U261 ( .A1(n575), .A2(n256), .A3(n208), .Y(n247) );
  NAND2X0_HVT U262 ( .A1(in[49]), .A2(n300), .Y(n212) );
  NAND2X0_HVT U263 ( .A1(n211), .A2(in[41]), .Y(n214) );
  NAND2X0_HVT U264 ( .A1(n212), .A2(n214), .Y(n115) );
  IBUFFX2_HVT U265 ( .A(in[49]), .Y(n211) );
  NAND2X0_HVT U266 ( .A1(n221), .A2(n217), .Y(n219) );
  NAND2X0_HVT U267 ( .A1(n215), .A2(n220), .Y(n222) );
  NAND2X0_HVT U268 ( .A1(n219), .A2(n222), .Y(out[100]) );
  INVX1_HVT U269 ( .A(n221), .Y(n215) );
  INVX0_HVT U270 ( .A(n220), .Y(n217) );
  NAND2X0_HVT U271 ( .A1(n66), .A2(n224), .Y(n225) );
  NAND2X0_HVT U272 ( .A1(n223), .A2(n67), .Y(n226) );
  NAND2X0_HVT U273 ( .A1(n225), .A2(n226), .Y(out[76]) );
  INVX0_HVT U274 ( .A(n67), .Y(n224) );
  XNOR2X2_HVT U275 ( .A1(n243), .A2(in[35]), .Y(n548) );
  INVX0_HVT U276 ( .A(in[58]), .Y(n380) );
  NAND2X0_HVT U277 ( .A1(in[93]), .A2(n228), .Y(n229) );
  NAND2X0_HVT U278 ( .A1(n227), .A2(in[78]), .Y(n230) );
  NAND2X0_HVT U279 ( .A1(n229), .A2(n230), .Y(n263) );
  INVX0_HVT U280 ( .A(in[93]), .Y(n227) );
  INVX1_HVT U281 ( .A(in[78]), .Y(n228) );
  INVX1_HVT U282 ( .A(n244), .Y(n232) );
  INVX1_HVT U283 ( .A(in[96]), .Y(n244) );
  XOR3X2_HVT U284 ( .A1(n260), .A2(n333), .A3(n540), .Y(n258) );
  NAND2X0_HVT U285 ( .A1(n233), .A2(in[61]), .Y(n235) );
  NAND2X0_HVT U286 ( .A1(n234), .A2(n235), .Y(n138) );
  XOR3X2_HVT U287 ( .A1(in[68]), .A2(in[67]), .A3(n139), .Y(n67) );
  XOR3X2_HVT U288 ( .A1(n26), .A2(n445), .A3(n27), .Y(out[96]) );
  XOR3X2_HVT U289 ( .A1(n236), .A2(n455), .A3(n257), .Y(n409) );
  NAND2X0_HVT U290 ( .A1(n90), .A2(n347), .Y(n237) );
  NAND2X0_HVT U291 ( .A1(n417), .A2(n528), .Y(n238) );
  NAND2X0_HVT U292 ( .A1(n237), .A2(n238), .Y(n468) );
  INVX0_HVT U293 ( .A(n468), .Y(n323) );
  NAND2X0_HVT U294 ( .A1(n438), .A2(n348), .Y(n240) );
  NAND2X0_HVT U295 ( .A1(n239), .A2(n437), .Y(n241) );
  NAND2X0_HVT U296 ( .A1(n240), .A2(n241), .Y(n531) );
  INVX1_HVT U297 ( .A(n438), .Y(n239) );
  INVX0_HVT U298 ( .A(in[50]), .Y(n242) );
  INVX1_HVT U299 ( .A(n242), .Y(n243) );
  XOR3X2_HVT U300 ( .A1(n189), .A2(n165), .A3(n216), .Y(out[105]) );
  INVX1_HVT U301 ( .A(n244), .Y(n245) );
  INVX0_HVT U302 ( .A(n201), .Y(n364) );
  INVX2_HVT U303 ( .A(in[42]), .Y(n337) );
  INVX1_HVT U304 ( .A(n50), .Y(n476) );
  XNOR3X1_HVT U305 ( .A1(n578), .A2(in[121]), .A3(n459), .Y(n251) );
  INVX0_HVT U306 ( .A(n493), .Y(n253) );
  XNOR2X2_HVT U307 ( .A1(n545), .A2(in[26]), .Y(n503) );
  XNOR2X2_HVT U308 ( .A1(n246), .A2(n247), .Y(out[115]) );
  XOR3X2_HVT U309 ( .A1(n534), .A2(n510), .A3(n511), .Y(n246) );
  INVX1_HVT U310 ( .A(in[33]), .Y(n264) );
  XNOR2X2_HVT U311 ( .A1(n176), .A2(n248), .Y(out[12]) );
  INVX1_HVT U312 ( .A(n527), .Y(n510) );
  INVX0_HVT U313 ( .A(n545), .Y(n379) );
  INVX0_HVT U314 ( .A(in[28]), .Y(n543) );
  XNOR2X2_HVT U315 ( .A1(n488), .A2(in[36]), .Y(n93) );
  XNOR2X2_HVT U316 ( .A1(in[45]), .A2(in[37]), .Y(n89) );
  INVX1_HVT U317 ( .A(in[51]), .Y(n260) );
  XOR3X2_HVT U318 ( .A1(n557), .A2(n422), .A3(n395), .Y(n161) );
  XOR2X2_HVT U319 ( .A1(in[58]), .A2(n568), .Y(n98) );
  XNOR2X1_HVT U320 ( .A1(n164), .A2(n568), .Y(n101) );
  INVX1_HVT U321 ( .A(in[114]), .Y(n534) );
  INVX0_HVT U322 ( .A(n40), .Y(n250) );
  XOR3X2_HVT U323 ( .A1(n249), .A2(n256), .A3(n445), .Y(n19) );
  INVX0_HVT U324 ( .A(n39), .Y(n318) );
  INVX0_HVT U325 ( .A(in[34]), .Y(n516) );
  XOR3X2_HVT U326 ( .A1(n39), .A2(n13), .A3(n250), .Y(out[90]) );
  XOR2X2_HVT U327 ( .A1(in[116]), .A2(in[124]), .Y(n181) );
  XNOR2X2_HVT U328 ( .A1(n299), .A2(n567), .Y(n104) );
  XNOR2X2_HVT U329 ( .A1(n256), .A2(n520), .Y(n438) );
  INVX0_HVT U330 ( .A(in[4]), .Y(n479) );
  XOR3X2_HVT U331 ( .A1(n23), .A2(n24), .A3(n251), .Y(out[97]) );
  INVX1_HVT U332 ( .A(in[115]), .Y(n507) );
  INVX0_HVT U333 ( .A(in[115]), .Y(n533) );
  XOR3X2_HVT U334 ( .A1(n31), .A2(in[93]), .A3(n476), .Y(out[85]) );
  XOR3X2_HVT U335 ( .A1(n31), .A2(n254), .A3(n65), .Y(out[78]) );
  XNOR2X2_HVT U336 ( .A1(n117), .A2(n255), .Y(out[4]) );
  XNOR2X1_HVT U337 ( .A1(in[112]), .A2(n587), .Y(n193) );
  XOR3X1_HVT U338 ( .A1(n544), .A2(n260), .A3(n93), .Y(n408) );
  INVX1_HVT U339 ( .A(n53), .Y(n257) );
  XOR3X2_HVT U340 ( .A1(n447), .A2(n457), .A3(n199), .Y(n221) );
  INVX1_HVT U341 ( .A(in[40]), .Y(n299) );
  INVX0_HVT U342 ( .A(in[25]), .Y(n505) );
  XOR2X1_HVT U343 ( .A1(in[94]), .A2(in[85]), .Y(n462) );
  XOR3X2_HVT U344 ( .A1(n259), .A2(n326), .A3(n292), .Y(n451) );
  INVX1_HVT U345 ( .A(n386), .Y(n395) );
  XOR3X2_HVT U346 ( .A1(n380), .A2(n260), .A3(n261), .Y(n141) );
  XNOR2X1_HVT U347 ( .A1(n568), .A2(in[59]), .Y(n261) );
  XOR3X2_HVT U348 ( .A1(n569), .A2(n262), .A3(in[65]), .Y(n72) );
  INVX1_HVT U349 ( .A(in[124]), .Y(n486) );
  XOR3X2_HVT U350 ( .A1(in[43]), .A2(n337), .A3(n529), .Y(n502) );
  INVX0_HVT U351 ( .A(n337), .Y(n338) );
  XOR3X2_HVT U352 ( .A1(n263), .A2(n291), .A3(n65), .Y(out[70]) );
  XNOR2X2_HVT U353 ( .A1(n265), .A2(n19), .Y(out[99]) );
  XOR3X2_HVT U354 ( .A1(n537), .A2(n562), .A3(n559), .Y(n152) );
  XNOR2X2_HVT U355 ( .A1(n408), .A2(n266), .Y(out[60]) );
  XOR3X2_HVT U356 ( .A1(n568), .A2(n433), .A3(n333), .Y(n266) );
  INVX0_HVT U357 ( .A(in[30]), .Y(n267) );
  INVX1_HVT U358 ( .A(n267), .Y(n268) );
  XOR2X2_HVT U359 ( .A1(n270), .A2(n555), .Y(n269) );
  NAND2X0_HVT U360 ( .A1(in[32]), .A2(n271), .Y(n272) );
  NAND2X0_HVT U361 ( .A1(n482), .A2(n563), .Y(n273) );
  NAND2X0_HVT U362 ( .A1(n272), .A2(n273), .Y(n133) );
  INVX1_HVT U363 ( .A(in[39]), .Y(n271) );
  INVX1_HVT U364 ( .A(n479), .Y(n480) );
  XNOR2X2_HVT U365 ( .A1(n61), .A2(n40), .Y(n277) );
  XOR3X2_HVT U366 ( .A1(n453), .A2(n549), .A3(n154), .Y(n452) );
  XOR2X2_HVT U367 ( .A1(in[4]), .A2(in[12]), .Y(n154) );
  INVX0_HVT U368 ( .A(n398), .Y(n275) );
  INVX1_HVT U369 ( .A(n276), .Y(out[31]) );
  XOR3X2_HVT U370 ( .A1(n146), .A2(n557), .A3(n78), .Y(n276) );
  XNOR2X2_HVT U371 ( .A1(n278), .A2(n72), .Y(out[73]) );
  XOR2X2_HVT U372 ( .A1(in[72]), .A2(n582), .Y(n295) );
  NAND2X0_HVT U373 ( .A1(n570), .A2(n280), .Y(n281) );
  NAND2X0_HVT U374 ( .A1(n279), .A2(n572), .Y(n282) );
  XOR3X2_HVT U375 ( .A1(n565), .A2(n301), .A3(n283), .Y(n434) );
  INVX1_HVT U376 ( .A(n284), .Y(n285) );
  INVX0_HVT U377 ( .A(n442), .Y(n286) );
  XOR2X2_HVT U378 ( .A1(n494), .A2(n569), .Y(n74) );
  XOR3X2_HVT U379 ( .A1(n31), .A2(n362), .A3(n139), .Y(out[93]) );
  XOR3X2_HVT U380 ( .A1(n188), .A2(n493), .A3(n24), .Y(out[114]) );
  INVX1_HVT U381 ( .A(in[46]), .Y(n423) );
  NAND2X0_HVT U382 ( .A1(n36), .A2(n315), .Y(n287) );
  NAND2X0_HVT U383 ( .A1(n287), .A2(n288), .Y(out[91]) );
  INVX1_HVT U384 ( .A(in[98]), .Y(n489) );
  XOR3X2_HVT U385 ( .A1(n70), .A2(n289), .A3(in[96]), .Y(n216) );
  XNOR3X1_HVT U386 ( .A1(n93), .A2(n435), .A3(n88), .Y(out[45]) );
  XOR3X2_HVT U387 ( .A1(n292), .A2(n450), .A3(n293), .Y(n515) );
  XNOR2X1_HVT U388 ( .A1(n522), .A2(in[83]), .Y(n293) );
  INVX1_HVT U389 ( .A(n378), .Y(n369) );
  XOR3X2_HVT U390 ( .A1(n513), .A2(in[81]), .A3(in[80]), .Y(n383) );
  XOR3X2_HVT U391 ( .A1(n102), .A2(n294), .A3(n103), .Y(out[57]) );
  XOR3X2_HVT U392 ( .A1(n160), .A2(n509), .A3(n149), .Y(out[10]) );
  INVX1_HVT U393 ( .A(n159), .Y(n357) );
  XOR3X2_HVT U394 ( .A1(n484), .A2(n563), .A3(n516), .Y(n541) );
  XOR3X1_HVT U395 ( .A1(n512), .A2(n280), .A3(n56), .Y(n524) );
  INVX1_HVT U396 ( .A(n518), .Y(n316) );
  XOR3X2_HVT U397 ( .A1(n295), .A2(n569), .A3(n43), .Y(out[64]) );
  NAND2X0_HVT U398 ( .A1(n330), .A2(in[67]), .Y(n297) );
  NAND2X0_HVT U399 ( .A1(n296), .A2(n331), .Y(n298) );
  NAND2X0_HVT U400 ( .A1(n297), .A2(n298), .Y(n80) );
  INVX0_HVT U401 ( .A(n330), .Y(n296) );
  INVX0_HVT U402 ( .A(n80), .Y(n473) );
  IBUFFX2_HVT U403 ( .A(in[52]), .Y(n544) );
  INVX1_HVT U404 ( .A(n566), .Y(n540) );
  XOR3X2_HVT U405 ( .A1(n145), .A2(n275), .A3(n294), .Y(out[32]) );
  XNOR2X2_HVT U406 ( .A1(in[66]), .A2(n450), .Y(n39) );
  INVX1_HVT U407 ( .A(n300), .Y(n301) );
  XOR3X2_HVT U408 ( .A1(n378), .A2(n518), .A3(n302), .Y(n81) );
  XNOR2X1_HVT U409 ( .A1(n574), .A2(in[91]), .Y(n302) );
  XNOR3X1_HVT U410 ( .A1(in[95]), .A2(in[92]), .A3(n498), .Y(n79) );
  INVX1_HVT U411 ( .A(in[91]), .Y(n522) );
  NAND2X0_HVT U412 ( .A1(in[62]), .A2(n304), .Y(n305) );
  NAND2X0_HVT U413 ( .A1(n303), .A2(in[53]), .Y(n306) );
  NAND2X0_HVT U414 ( .A1(n305), .A2(n306), .Y(n407) );
  INVX1_HVT U415 ( .A(in[53]), .Y(n304) );
  INVX0_HVT U416 ( .A(in[55]), .Y(n539) );
  XOR3X2_HVT U417 ( .A1(n119), .A2(n105), .A3(n434), .Y(out[49]) );
  INVX1_HVT U418 ( .A(n89), .Y(n416) );
  NBUFFX2_HVT U419 ( .A(in[47]), .Y(n565) );
  XNOR2X2_HVT U420 ( .A1(n422), .A2(in[25]), .Y(n16) );
  XNOR2X2_HVT U421 ( .A1(n332), .A2(in[40]), .Y(n145) );
  INVX1_HVT U422 ( .A(n558), .Y(n317) );
  NAND2X0_HVT U423 ( .A1(n134), .A2(n308), .Y(n309) );
  NAND2X0_HVT U424 ( .A1(n307), .A2(n135), .Y(n310) );
  NAND2X0_HVT U425 ( .A1(n309), .A2(n310), .Y(out[3]) );
  INVX0_HVT U426 ( .A(n134), .Y(n307) );
  INVX0_HVT U427 ( .A(n135), .Y(n308) );
  XOR3X2_HVT U428 ( .A1(n550), .A2(n546), .A3(n514), .Y(n412) );
  NAND2X0_HVT U429 ( .A1(n55), .A2(n524), .Y(n313) );
  NAND2X0_HVT U430 ( .A1(n311), .A2(n312), .Y(n314) );
  NAND2X0_HVT U431 ( .A1(n313), .A2(n314), .Y(out[83]) );
  INVX1_HVT U432 ( .A(n524), .Y(n311) );
  INVX0_HVT U433 ( .A(n55), .Y(n312) );
  XNOR3X1_HVT U434 ( .A1(n539), .A2(in[51]), .A3(n98), .Y(n485) );
  XOR3X2_HVT U435 ( .A1(n13), .A2(in[67]), .A3(n49), .Y(n315) );
  XOR3X2_HVT U436 ( .A1(n530), .A2(n549), .A3(n317), .Y(n166) );
  XOR3X2_HVT U437 ( .A1(n57), .A2(n369), .A3(n318), .Y(out[82]) );
  XOR3X2_HVT U438 ( .A1(n550), .A2(n554), .A3(in[10]), .Y(n319) );
  XOR3X2_HVT U439 ( .A1(n586), .A2(n413), .A3(n177), .Y(out[127]) );
  INVX0_HVT U440 ( .A(n587), .Y(n413) );
  INVX1_HVT U441 ( .A(n321), .Y(out[39]) );
  XOR3X2_HVT U442 ( .A1(n137), .A2(in[38]), .A3(n123), .Y(n321) );
  NAND2X0_HVT U443 ( .A1(n529), .A2(n468), .Y(n324) );
  NAND2X0_HVT U444 ( .A1(n322), .A2(n323), .Y(n325) );
  NAND2X0_HVT U445 ( .A1(n324), .A2(n325), .Y(n126) );
  INVX0_HVT U446 ( .A(n126), .Y(n390) );
  XNOR2X2_HVT U447 ( .A1(n275), .A2(n565), .Y(n86) );
  XOR3X2_HVT U448 ( .A1(n559), .A2(n143), .A3(n327), .Y(n399) );
  NBUFFX2_HVT U449 ( .A(in[116]), .Y(n329) );
  NAND2X0_HVT U450 ( .A1(n478), .A2(n477), .Y(n330) );
  XNOR2X1_HVT U451 ( .A1(in[18]), .A2(in[26]), .Y(n149) );
  NAND2X0_HVT U452 ( .A1(in[48]), .A2(n539), .Y(n334) );
  NAND2X0_HVT U453 ( .A1(n332), .A2(n333), .Y(n335) );
  NAND2X0_HVT U454 ( .A1(n334), .A2(n335), .Y(n105) );
  INVX0_HVT U455 ( .A(n539), .Y(n333) );
  XOR3X2_HVT U456 ( .A1(n564), .A2(n337), .A3(n129), .Y(n127) );
  XOR3X2_HVT U457 ( .A1(n42), .A2(n320), .A3(n169), .Y(out[1]) );
  INVX1_HVT U458 ( .A(n497), .Y(n336) );
  INVX1_HVT U459 ( .A(in[121]), .Y(n497) );
  XNOR2X2_HVT U460 ( .A1(n359), .A2(n491), .Y(n179) );
  INVX1_HVT U461 ( .A(in[55]), .Y(n536) );
  NAND2X0_HVT U462 ( .A1(n81), .A2(n340), .Y(n341) );
  NAND2X0_HVT U463 ( .A1(n339), .A2(n82), .Y(n342) );
  NAND2X0_HVT U464 ( .A1(n341), .A2(n342), .Y(out[67]) );
  INVX0_HVT U465 ( .A(n81), .Y(n339) );
  INVX1_HVT U466 ( .A(n82), .Y(n340) );
  XNOR2X1_HVT U467 ( .A1(in[33]), .A2(n301), .Y(n102) );
  XNOR2X1_HVT U468 ( .A1(in[110]), .A2(n492), .Y(n439) );
  XOR3X2_HVT U469 ( .A1(in[75]), .A2(n279), .A3(n499), .Y(n82) );
  NAND2X0_HVT U470 ( .A1(n485), .A2(n97), .Y(n345) );
  NAND2X0_HVT U471 ( .A1(n343), .A2(n344), .Y(n346) );
  NAND2X0_HVT U472 ( .A1(n345), .A2(n346), .Y(out[59]) );
  INVX0_HVT U473 ( .A(n485), .Y(n343) );
  INVX0_HVT U474 ( .A(n97), .Y(n344) );
  XOR2X2_HVT U475 ( .A1(in[36]), .A2(in[60]), .Y(n111) );
  XNOR2X1_HVT U476 ( .A1(n232), .A2(n458), .Y(n23) );
  XOR2X2_HVT U477 ( .A1(in[1]), .A2(in[25]), .Y(n148) );
  XOR3X2_HVT U478 ( .A1(n95), .A2(n467), .A3(n94), .Y(out[5]) );
  XNOR2X2_HVT U479 ( .A1(n274), .A2(in[97]), .Y(n190) );
  INVX0_HVT U480 ( .A(in[84]), .Y(n547) );
  XOR3X2_HVT U481 ( .A1(n507), .A2(n534), .A3(n256), .Y(n349) );
  XOR2X2_HVT U482 ( .A1(in[81]), .A2(in[89]), .Y(n40) );
  NAND2X0_HVT U483 ( .A1(n182), .A2(n415), .Y(n352) );
  NAND2X0_HVT U484 ( .A1(n350), .A2(n351), .Y(n353) );
  NAND2X0_HVT U485 ( .A1(n352), .A2(n353), .Y(out[124]) );
  INVX1_HVT U486 ( .A(n415), .Y(n350) );
  INVX0_HVT U487 ( .A(n182), .Y(n351) );
  XOR3X2_HVT U488 ( .A1(n329), .A2(n508), .A3(n184), .Y(n415) );
  XOR3X2_HVT U489 ( .A1(n179), .A2(n440), .A3(n202), .Y(out[101]) );
  INVX1_HVT U490 ( .A(in[88]), .Y(n354) );
  INVX1_HVT U491 ( .A(n354), .Y(n355) );
  INVX1_HVT U492 ( .A(n427), .Y(n356) );
  INVX1_HVT U493 ( .A(in[3]), .Y(n427) );
  XOR3X2_HVT U494 ( .A1(n358), .A2(n386), .A3(n357), .Y(out[0]) );
  XOR2X2_HVT U495 ( .A1(n465), .A2(n551), .Y(n358) );
  INVX1_HVT U496 ( .A(in[119]), .Y(n587) );
  XOR3X2_HVT U497 ( .A1(n124), .A2(n435), .A3(n138), .Y(out[38]) );
  INVX1_HVT U498 ( .A(in[90]), .Y(n378) );
  XNOR2X2_HVT U499 ( .A1(n498), .A2(n372), .Y(n56) );
  INVX1_HVT U500 ( .A(in[117]), .Y(n359) );
  INVX1_HVT U501 ( .A(n546), .Y(n381) );
  INVX1_HVT U502 ( .A(n545), .Y(n546) );
  XOR3X2_HVT U503 ( .A1(n320), .A2(n401), .A3(n158), .Y(out[18]) );
  XOR2X2_HVT U504 ( .A1(n574), .A2(n369), .Y(n38) );
  INVX1_HVT U505 ( .A(in[21]), .Y(n424) );
  XNOR2X2_HVT U506 ( .A1(n496), .A2(n573), .Y(n64) );
  INVX1_HVT U507 ( .A(n29), .Y(n461) );
  XNOR2X2_HVT U508 ( .A1(n362), .A2(in[93]), .Y(n30) );
  INVX0_HVT U509 ( .A(in[36]), .Y(n528) );
  XNOR2X2_HVT U510 ( .A1(n495), .A2(n322), .Y(n363) );
  NAND2X0_HVT U511 ( .A1(n201), .A2(n365), .Y(n366) );
  NAND2X0_HVT U512 ( .A1(n364), .A2(n200), .Y(n367) );
  NAND2X0_HVT U513 ( .A1(n366), .A2(n367), .Y(out[116]) );
  INVX1_HVT U514 ( .A(n200), .Y(n365) );
  XOR3X2_HVT U515 ( .A1(n527), .A2(n507), .A3(n577), .Y(n200) );
  XOR3X2_HVT U516 ( .A1(n449), .A2(in[107]), .A3(n202), .Y(n201) );
  XNOR2X2_HVT U517 ( .A1(n580), .A2(in[16]), .Y(n368) );
  NBUFFX2_HVT U518 ( .A(in[37]), .Y(n435) );
  XOR3X2_HVT U519 ( .A1(n576), .A2(in[105]), .A3(n286), .Y(n370) );
  NAND2X0_HVT U520 ( .A1(n140), .A2(n384), .Y(n376) );
  NAND2X0_HVT U521 ( .A1(n375), .A2(n363), .Y(n377) );
  NAND2X0_HVT U522 ( .A1(n377), .A2(n376), .Y(out[36]) );
  INVX0_HVT U523 ( .A(n384), .Y(n375) );
  XOR2X2_HVT U524 ( .A1(in[58]), .A2(in[50]), .Y(n130) );
  XOR2X2_HVT U525 ( .A1(in[1]), .A2(n285), .Y(n160) );
  XOR3X2_HVT U526 ( .A1(n115), .A2(n380), .A3(n99), .Y(out[50]) );
  XOR2X1_HVT U527 ( .A1(in[51]), .A2(in[59]), .Y(n129) );
  XOR3X2_HVT U528 ( .A1(n43), .A2(n44), .A3(n383), .Y(out[89]) );
  XOR3X2_HVT U529 ( .A1(in[49]), .A2(n333), .A3(n332), .Y(n103) );
  XOR3X2_HVT U530 ( .A1(n567), .A2(in[60]), .A3(in[59]), .Y(n384) );
  XOR3X2_HVT U531 ( .A1(n197), .A2(n385), .A3(n177), .Y(out[119]) );
  INVX0_HVT U532 ( .A(in[22]), .Y(n426) );
  IBUFFX2_HVT U533 ( .A(in[118]), .Y(n387) );
  INVX1_HVT U534 ( .A(n387), .Y(n388) );
  NAND2X0_HVT U535 ( .A1(n2), .A2(n483), .Y(n391) );
  NAND2X0_HVT U536 ( .A1(n389), .A2(n390), .Y(n392) );
  NAND2X0_HVT U537 ( .A1(n391), .A2(n392), .Y(out[44]) );
  INVX1_HVT U538 ( .A(n483), .Y(n389) );
  XOR3X2_HVT U539 ( .A1(n269), .A2(n402), .A3(n393), .Y(out[16]) );
  XOR2X2_HVT U540 ( .A1(n580), .A2(n558), .Y(n393) );
  XOR3X2_HVT U541 ( .A1(n115), .A2(n396), .A3(n133), .Y(out[33]) );
  XNOR2X2_HVT U542 ( .A1(n557), .A2(n560), .Y(n63) );
  XOR3X2_HVT U543 ( .A1(n16), .A2(n83), .A3(n17), .Y(out[9]) );
  XNOR2X2_HVT U544 ( .A1(n271), .A2(n521), .Y(n495) );
  XOR3X2_HVT U545 ( .A1(n401), .A2(n558), .A3(n157), .Y(n411) );
  XOR3X2_HVT U546 ( .A1(n404), .A2(n467), .A3(n403), .Y(out[22]) );
  XOR3X2_HVT U547 ( .A1(n124), .A2(n405), .A3(n89), .Y(out[46]) );
  XNOR2X1_HVT U548 ( .A1(in[99]), .A2(in[123]), .Y(n511) );
  INVX0_HVT U549 ( .A(n578), .Y(n410) );
  INVX1_HVT U550 ( .A(n519), .Y(n506) );
  INVX1_HVT U551 ( .A(in[43]), .Y(n484) );
  INVX1_HVT U552 ( .A(in[32]), .Y(n482) );
  INVX1_HVT U553 ( .A(n289), .Y(n445) );
  XOR2X2_HVT U554 ( .A1(in[34]), .A2(n563), .Y(n406) );
  INVX1_HVT U555 ( .A(n79), .Y(n481) );
  INVX1_HVT U556 ( .A(in[122]), .Y(n493) );
  INVX1_HVT U557 ( .A(in[74]), .Y(n526) );
  INVX0_HVT U558 ( .A(in[102]), .Y(n429) );
  INVX1_HVT U559 ( .A(n65), .Y(n583) );
  XNOR2X1_HVT U560 ( .A1(in[88]), .A2(n584), .Y(n60) );
  XOR3X2_HVT U561 ( .A1(n407), .A2(in[45]), .A3(n87), .Y(out[54]) );
  INVX1_HVT U562 ( .A(n419), .Y(out[53]) );
  INVX1_HVT U563 ( .A(n180), .Y(n436) );
  XOR3X2_HVT U564 ( .A1(n53), .A2(n460), .A3(n30), .Y(out[69]) );
  XOR2X2_HVT U565 ( .A1(n51), .A2(n409), .Y(out[84]) );
  XNOR2X1_HVT U566 ( .A1(n587), .A2(n410), .Y(n209) );
  XOR3X2_HVT U567 ( .A1(n414), .A2(n413), .A3(n165), .Y(out[112]) );
  XNOR2X2_HVT U568 ( .A1(in[38]), .A2(n423), .Y(n87) );
  INVX1_HVT U569 ( .A(in[123]), .Y(n447) );
  XOR3X2_HVT U570 ( .A1(n416), .A2(n304), .A3(n417), .Y(out[61]) );
  XNOR2X2_HVT U571 ( .A1(in[22]), .A2(n268), .Y(n78) );
  INVX0_HVT U572 ( .A(n87), .Y(n441) );
  XNOR2X2_HVT U573 ( .A1(n418), .A2(n166), .Y(out[20]) );
  INVX0_HVT U574 ( .A(in[12]), .Y(n500) );
  XNOR2X2_HVT U575 ( .A1(n425), .A2(in[29]), .Y(n94) );
  XNOR2X1_HVT U576 ( .A1(n569), .A2(n572), .Y(n28) );
  INVX1_HVT U577 ( .A(in[120]), .Y(n459) );
  INVX1_HVT U578 ( .A(n517), .Y(n499) );
  XOR3X2_HVT U579 ( .A1(n108), .A2(in[61]), .A3(n89), .Y(n419) );
  XOR2X1_HVT U580 ( .A1(in[100]), .A2(in[124]), .Y(n202) );
  INVX0_HVT U581 ( .A(n30), .Y(n428) );
  IBUFFX2_HVT U582 ( .A(n193), .Y(n443) );
  XOR3X2_HVT U583 ( .A1(n124), .A2(n536), .A3(n86), .Y(out[63]) );
  XOR3X2_HVT U584 ( .A1(n420), .A2(n564), .A3(n133), .Y(out[40]) );
  XNOR2X2_HVT U585 ( .A1(in[102]), .A2(in[110]), .Y(n178) );
  XOR3X2_HVT U586 ( .A1(n421), .A2(n148), .A3(n163), .Y(out[17]) );
  XOR3X2_HVT U587 ( .A1(in[9]), .A2(n465), .A3(n556), .Y(n421) );
  XNOR2X2_HVT U588 ( .A1(in[30]), .A2(n471), .Y(n490) );
  XOR3X2_HVT U589 ( .A1(n106), .A2(n423), .A3(n86), .Y(out[55]) );
  XOR3X2_HVT U590 ( .A1(n104), .A2(in[32]), .A3(n14), .Y(out[56]) );
  XOR3X2_HVT U591 ( .A1(n150), .A2(n470), .A3(n78), .Y(out[14]) );
  XOR3X2_HVT U592 ( .A1(n147), .A2(n426), .A3(n94), .Y(out[30]) );
  INVX1_HVT U593 ( .A(n469), .Y(n472) );
  XOR2X2_HVT U594 ( .A1(in[126]), .A2(in[118]), .Y(n210) );
  XOR3X2_HVT U595 ( .A1(n74), .A2(n57), .A3(n430), .Y(out[65]) );
  XOR3X2_HVT U596 ( .A1(n573), .A2(in[89]), .A3(n355), .Y(n430) );
  XOR3X2_HVT U597 ( .A1(n121), .A2(in[32]), .A3(n122), .Y(out[48]) );
  XNOR2X2_HVT U598 ( .A1(n213), .A2(n431), .Y(out[107]) );
  XOR3X2_HVT U599 ( .A1(n577), .A2(in[106]), .A3(n457), .Y(n431) );
  INVX1_HVT U600 ( .A(n303), .Y(n432) );
  XOR2X2_HVT U601 ( .A1(in[76]), .A2(in[84]), .Y(n50) );
  XOR3X2_HVT U602 ( .A1(n436), .A2(n492), .A3(n199), .Y(out[117]) );
  XNOR2X2_HVT U603 ( .A1(n136), .A2(n316), .Y(n51) );
  XOR3X2_HVT U604 ( .A1(n439), .A2(n469), .A3(n586), .Y(out[102]) );
  XOR3X2_HVT U605 ( .A1(n198), .A2(n440), .A3(n178), .Y(out[118]) );
  XOR3X2_HVT U606 ( .A1(n123), .A2(n275), .A3(n441), .Y(out[47]) );
  XOR3X2_HVT U607 ( .A1(n566), .A2(n398), .A3(n484), .Y(n483) );
  INVX1_HVT U608 ( .A(n181), .Y(n448) );
  XNOR3X1_HVT U609 ( .A1(n181), .A2(n360), .A3(n180), .Y(out[125]) );
  XOR3X2_HVT U610 ( .A1(n178), .A2(n445), .A3(n209), .Y(out[111]) );
  XOR3X2_HVT U611 ( .A1(n27), .A2(n190), .A3(n446), .Y(out[121]) );
  XOR3X2_HVT U612 ( .A1(n587), .A2(n585), .A3(n116), .Y(n446) );
  XOR3X2_HVT U613 ( .A1(n578), .A2(n527), .A3(n447), .Y(n182) );
  XOR3X2_HVT U614 ( .A1(n457), .A2(in[100]), .A3(n448), .Y(n532) );
  XOR2X2_HVT U615 ( .A1(in[0]), .A2(n552), .Y(n42) );
  XOR2X2_HVT U616 ( .A1(n432), .A2(n566), .Y(n137) );
  XOR2X2_HVT U617 ( .A1(n555), .A2(n553), .Y(n146) );
  INVX1_HVT U618 ( .A(n526), .Y(n450) );
  XOR3X2_HVT U619 ( .A1(n60), .A2(n494), .A3(n61), .Y(out[80]) );
  NBUFFX2_HVT U620 ( .A(in[15]), .Y(n555) );
  INVX1_HVT U621 ( .A(n575), .Y(n520) );
  NBUFFX2_HVT U622 ( .A(in[7]), .Y(n551) );
  XOR2X2_HVT U623 ( .A1(in[120]), .A2(n20), .Y(n27) );
  XOR3X2_HVT U624 ( .A1(n58), .A2(n47), .A3(n451), .Y(out[81]) );
  XOR3X2_HVT U625 ( .A1(n551), .A2(n454), .A3(in[0]), .Y(n17) );
  XOR2X2_HVT U626 ( .A1(in[24]), .A2(n561), .Y(n159) );
  INVX1_HVT U627 ( .A(in[24]), .Y(n580) );
  NBUFFX2_HVT U628 ( .A(in[23]), .Y(n559) );
  XOR2X2_HVT U629 ( .A1(n536), .A2(n567), .Y(n123) );
  XOR2X2_HVT U630 ( .A1(in[68]), .A2(in[92]), .Y(n53) );
  XOR3X2_HVT U631 ( .A1(n75), .A2(n254), .A3(n64), .Y(out[71]) );
  XNOR2X2_HVT U632 ( .A1(n355), .A2(n574), .Y(n43) );
  NBUFFX2_HVT U633 ( .A(in[71]), .Y(n569) );
  INVX1_HVT U634 ( .A(in[8]), .Y(n464) );
  XOR3X2_HVT U635 ( .A1(n466), .A2(n572), .A3(n74), .Y(out[72]) );
  INVX1_HVT U636 ( .A(in[13]), .Y(n467) );
  XNOR2X2_HVT U637 ( .A1(n548), .A2(n484), .Y(n97) );
  NBUFFX2_HVT U638 ( .A(in[101]), .Y(n469) );
  XNOR2X2_HVT U639 ( .A1(in[109]), .A2(in[101]), .Y(n180) );
  INVX1_HVT U640 ( .A(n470), .Y(n471) );
  XOR3X2_HVT U641 ( .A1(n179), .A2(n472), .A3(n184), .Y(out[109]) );
  NAND2X0_HVT U642 ( .A1(n481), .A2(n80), .Y(n474) );
  NAND2X0_HVT U643 ( .A1(n79), .A2(n473), .Y(n475) );
  NAND2X0_HVT U644 ( .A1(n475), .A2(n474), .Y(out[68]) );
  INVX1_HVT U645 ( .A(in[80]), .Y(n582) );
  NAND2X0_HVT U646 ( .A1(n50), .A2(n279), .Y(n477) );
  NAND2X0_HVT U647 ( .A1(n476), .A2(in[71]), .Y(n478) );
  XOR3X2_HVT U648 ( .A1(n30), .A2(n192), .A3(n29), .Y(out[94]) );
  XOR3X2_HVT U649 ( .A1(n488), .A2(n111), .A3(in[43]), .Y(n110) );
  XOR3X2_HVT U650 ( .A1(n218), .A2(n429), .A3(n209), .Y(out[103]) );
  XOR3X2_HVT U651 ( .A1(n22), .A2(n208), .A3(n21), .Y(out[98]) );
  XOR3X2_HVT U652 ( .A1(n490), .A2(n556), .A3(n63), .Y(out[7]) );
  XOR3X2_HVT U653 ( .A1(n47), .A2(n494), .A3(n46), .Y(out[88]) );
  XNOR2X2_HVT U654 ( .A1(n495), .A2(n529), .Y(n140) );
  XOR3X2_HVT U655 ( .A1(n88), .A2(n205), .A3(n87), .Y(out[62]) );
  XOR3X2_HVT U656 ( .A1(n583), .A2(n373), .A3(n28), .Y(out[95]) );
  XOR2X2_HVT U657 ( .A1(in[80]), .A2(n513), .Y(n47) );
  INVX1_HVT U658 ( .A(in[11]), .Y(n545) );
  XOR2X2_HVT U659 ( .A1(in[70]), .A2(n231), .Y(n29) );
  INVX1_HVT U660 ( .A(in[66]), .Y(n517) );
  XNOR2X2_HVT U661 ( .A1(in[77]), .A2(in[69]), .Y(n31) );
  XOR3X2_HVT U662 ( .A1(n151), .A2(n425), .A3(n1), .Y(out[29]) );
  XOR3X2_HVT U663 ( .A1(n150), .A2(in[29]), .A3(n118), .Y(out[21]) );
  XOR2X2_HVT U664 ( .A1(in[13]), .A2(in[5]), .Y(n150) );
  XOR2X2_HVT U665 ( .A1(n564), .A2(in[40]), .Y(n122) );
  XOR3X2_HVT U666 ( .A1(n504), .A2(in[14]), .A3(n78), .Y(out[6]) );
  XOR3X2_HVT U667 ( .A1(n560), .A2(n505), .A3(in[24]), .Y(n169) );
  XNOR2X2_HVT U668 ( .A1(n452), .A2(n152), .Y(out[28]) );
  XOR2X2_HVT U669 ( .A1(n465), .A2(n562), .Y(n162) );
  XNOR2X2_HVT U670 ( .A1(n194), .A2(n319), .Y(out[11]) );
  XOR3X2_HVT U671 ( .A1(n148), .A2(n506), .A3(n149), .Y(out[2]) );
  XNOR2X2_HVT U672 ( .A1(n503), .A2(n550), .Y(n135) );
  XNOR2X2_HVT U673 ( .A1(in[34]), .A2(in[42]), .Y(n99) );
  XOR3X2_HVT U674 ( .A1(n158), .A2(n514), .A3(n16), .Y(out[26]) );
  XNOR2X2_HVT U675 ( .A1(in[2]), .A2(in[10]), .Y(n158) );
  XNOR2X2_HVT U676 ( .A1(n515), .A2(n69), .Y(out[75]) );
  XOR2X2_HVT U677 ( .A1(in[62]), .A2(in[54]), .Y(n124) );
  XOR3X2_HVT U678 ( .A1(n130), .A2(n516), .A3(n102), .Y(out[42]) );
  XOR3X2_HVT U679 ( .A1(n71), .A2(n517), .A3(n44), .Y(out[74]) );
  NBUFFX2_HVT U680 ( .A(in[10]), .Y(n519) );
  XNOR2X2_HVT U681 ( .A1(n523), .A2(n34), .Y(out[92]) );
  XOR3X2_HVT U682 ( .A1(n574), .A2(n498), .A3(n373), .Y(n523) );
  XOR3X2_HVT U683 ( .A1(n99), .A2(n525), .A3(n100), .Y(out[58]) );
  XOR3X2_HVT U684 ( .A1(n45), .A2(n331), .A3(n526), .Y(n55) );
  XOR3X2_HVT U685 ( .A1(n71), .A2(n450), .A3(n58), .Y(out[66]) );
  XOR3X2_HVT U686 ( .A1(n130), .A2(n338), .A3(n119), .Y(out[34]) );
  NBUFFX2_HVT U687 ( .A(in[119]), .Y(n527) );
  XNOR2X2_HVT U688 ( .A1(n531), .A2(n532), .Y(out[108]) );
  XOR3X2_HVT U689 ( .A1(n189), .A2(in[114]), .A3(n188), .Y(out[122]) );
  XNOR2X2_HVT U690 ( .A1(n141), .A2(n541), .Y(out[35]) );
  NBUFFX2_HVT U691 ( .A(in[15]), .Y(n556) );
  NBUFFX2_HVT U692 ( .A(in[71]), .Y(n570) );
  NBUFFX2_HVT U693 ( .A(in[63]), .Y(n568) );
  NBUFFX2_HVT U694 ( .A(in[95]), .Y(n574) );
  NBUFFX2_HVT U695 ( .A(in[111]), .Y(n577) );
  NBUFFX2_HVT U696 ( .A(in[47]), .Y(n566) );
  NBUFFX2_HVT U697 ( .A(in[31]), .Y(n562) );
  NBUFFX2_HVT U698 ( .A(in[79]), .Y(n572) );
  NBUFFX2_HVT U699 ( .A(in[111]), .Y(n576) );
  NBUFFX2_HVT U700 ( .A(in[7]), .Y(n553) );
  NBUFFX2_HVT U701 ( .A(in[63]), .Y(n567) );
  NBUFFX2_HVT U702 ( .A(in[95]), .Y(n573) );
  NBUFFX2_HVT U703 ( .A(in[7]), .Y(n552) );
  NBUFFX2_HVT U704 ( .A(in[23]), .Y(n558) );
  NBUFFX2_HVT U705 ( .A(in[111]), .Y(n575) );
  NBUFFX2_HVT U706 ( .A(in[31]), .Y(n561) );
  NBUFFX2_HVT U707 ( .A(in[127]), .Y(n579) );
  NBUFFX2_HVT U708 ( .A(in[23]), .Y(n557) );
  NBUFFX2_HVT U709 ( .A(in[15]), .Y(n554) );
  NBUFFX2_HVT U710 ( .A(in[127]), .Y(n578) );
  NBUFFX2_HVT U711 ( .A(in[31]), .Y(n560) );
  NBUFFX2_HVT U712 ( .A(in[47]), .Y(n564) );
  NBUFFX2_HVT U713 ( .A(in[79]), .Y(n571) );
  INVX0_HVT U714 ( .A(in[0]), .Y(n581) );
endmodule

