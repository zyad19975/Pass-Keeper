
module add_round_keys_1 ( state, subkey, out );
  input [127:0] state;
  input [127:0] subkey;
  output [127:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538;

  INVX0_HVT U1 ( .A(subkey[114]), .Y(n244) );
  INVX0_HVT U2 ( .A(state[58]), .Y(n225) );
  INVX1_HVT U3 ( .A(state[25]), .Y(n448) );
  INVX1_HVT U4 ( .A(subkey[27]), .Y(n473) );
  INVX1_HVT U5 ( .A(state[73]), .Y(n167) );
  INVX1_HVT U6 ( .A(state[17]), .Y(n275) );
  INVX1_HVT U7 ( .A(subkey[71]), .Y(n445) );
  INVX1_HVT U8 ( .A(subkey[29]), .Y(n151) );
  INVX0_HVT U9 ( .A(state[41]), .Y(n339) );
  INVX0_HVT U10 ( .A(subkey[11]), .Y(n272) );
  INVX1_HVT U11 ( .A(state[22]), .Y(n198) );
  INVX0_HVT U12 ( .A(state[95]), .Y(n119) );
  INVX1_HVT U13 ( .A(subkey[125]), .Y(n64) );
  INVX1_HVT U14 ( .A(state[9]), .Y(n130) );
  INVX0_HVT U15 ( .A(subkey[124]), .Y(n372) );
  INVX0_HVT U16 ( .A(n517), .Y(n1) );
  INVX1_HVT U17 ( .A(subkey[95]), .Y(n118) );
  INVX1_HVT U18 ( .A(subkey[50]), .Y(n409) );
  INVX0_HVT U19 ( .A(n513), .Y(n2) );
  INVX1_HVT U20 ( .A(state[49]), .Y(n413) );
  INVX1_HVT U21 ( .A(subkey[1]), .Y(n487) );
  INVX1_HVT U22 ( .A(n50), .Y(n18) );
  INVX0_HVT U23 ( .A(subkey[2]), .Y(n50) );
  INVX1_HVT U24 ( .A(subkey[108]), .Y(n364) );
  INVX1_HVT U25 ( .A(subkey[57]), .Y(n299) );
  INVX1_HVT U26 ( .A(subkey[96]), .Y(n334) );
  INVX0_HVT U27 ( .A(subkey[99]), .Y(n483) );
  INVX1_HVT U28 ( .A(subkey[101]), .Y(n253) );
  INVX0_HVT U29 ( .A(subkey[107]), .Y(n383) );
  INVX1_HVT U30 ( .A(subkey[113]), .Y(n300) );
  INVX1_HVT U31 ( .A(subkey[88]), .Y(n40) );
  INVX1_HVT U32 ( .A(subkey[105]), .Y(n501) );
  INVX1_HVT U33 ( .A(n244), .Y(n210) );
  INVX1_HVT U34 ( .A(subkey[116]), .Y(n480) );
  INVX1_HVT U35 ( .A(subkey[120]), .Y(n493) );
  INVX1_HVT U36 ( .A(subkey[100]), .Y(n110) );
  INVX1_HVT U37 ( .A(subkey[115]), .Y(n263) );
  INVX1_HVT U38 ( .A(subkey[112]), .Y(n477) );
  INVX0_HVT U39 ( .A(subkey[61]), .Y(n139) );
  INVX1_HVT U40 ( .A(subkey[106]), .Y(n344) );
  INVX1_HVT U41 ( .A(subkey[104]), .Y(n27) );
  INVX1_HVT U42 ( .A(subkey[118]), .Y(n488) );
  INVX1_HVT U43 ( .A(subkey[97]), .Y(n279) );
  INVX1_HVT U44 ( .A(subkey[126]), .Y(n348) );
  INVX1_HVT U45 ( .A(subkey[117]), .Y(n284) );
  INVX1_HVT U46 ( .A(subkey[109]), .Y(n321) );
  INVX0_HVT U47 ( .A(n281), .Y(n3) );
  INVX0_HVT U48 ( .A(n193), .Y(n4) );
  INVX1_HVT U49 ( .A(subkey[102]), .Y(n96) );
  INVX0_HVT U50 ( .A(n305), .Y(n5) );
  OR2X1_HVT U51 ( .A1(subkey[119]), .A2(n245), .Y(n246) );
  INVX0_HVT U52 ( .A(n465), .Y(n37) );
  INVX0_HVT U53 ( .A(n222), .Y(n6) );
  INVX0_HVT U54 ( .A(n394), .Y(n54) );
  INVX0_HVT U55 ( .A(subkey[10]), .Y(n174) );
  INVX0_HVT U56 ( .A(n187), .Y(n7) );
  INVX0_HVT U57 ( .A(n424), .Y(n8) );
  INVX0_HVT U58 ( .A(n535), .Y(n9) );
  INVX0_HVT U59 ( .A(subkey[75]), .Y(n535) );
  INVX1_HVT U60 ( .A(state[111]), .Y(n111) );
  NAND2X0_HVT U61 ( .A1(state[118]), .A2(n488), .Y(n11) );
  NAND2X0_HVT U62 ( .A1(subkey[118]), .A2(n10), .Y(n12) );
  NAND2X0_HVT U63 ( .A1(n11), .A2(n12), .Y(out[118]) );
  INVX0_HVT U64 ( .A(state[118]), .Y(n10) );
  OR2X1_HVT U65 ( .A1(subkey[54]), .A2(n317), .Y(n319) );
  NAND2X0_HVT U66 ( .A1(state[106]), .A2(n344), .Y(n14) );
  NAND2X0_HVT U67 ( .A1(n13), .A2(subkey[106]), .Y(n15) );
  NAND2X0_HVT U68 ( .A1(n14), .A2(n15), .Y(out[106]) );
  INVX0_HVT U69 ( .A(state[106]), .Y(n13) );
  INVX0_HVT U70 ( .A(subkey[25]), .Y(n449) );
  INVX0_HVT U71 ( .A(n532), .Y(n32) );
  OR2X1_HVT U72 ( .A1(subkey[98]), .A2(n327), .Y(n329) );
  OR2X1_HVT U73 ( .A1(subkey[46]), .A2(n324), .Y(n325) );
  INVX1_HVT U74 ( .A(n371), .Y(n21) );
  OR2X1_HVT U75 ( .A1(subkey[31]), .A2(n421), .Y(n422) );
  INVX0_HVT U76 ( .A(n126), .Y(n16) );
  NAND2X0_HVT U77 ( .A1(state[2]), .A2(n50), .Y(n19) );
  NAND2X0_HVT U78 ( .A1(n18), .A2(n17), .Y(n20) );
  NAND2X0_HVT U79 ( .A1(n19), .A2(n20), .Y(out[2]) );
  INVX0_HVT U80 ( .A(state[2]), .Y(n17) );
  INVX0_HVT U81 ( .A(subkey[14]), .Y(n301) );
  INVX0_HVT U82 ( .A(state[42]), .Y(n182) );
  INVX0_HVT U83 ( .A(subkey[103]), .Y(n218) );
  INVX0_HVT U84 ( .A(subkey[91]), .Y(n457) );
  NAND2X0_HVT U85 ( .A1(state[104]), .A2(n27), .Y(n23) );
  NAND2X0_HVT U86 ( .A1(n22), .A2(subkey[104]), .Y(n24) );
  NAND2X0_HVT U87 ( .A1(n23), .A2(n24), .Y(out[104]) );
  INVX0_HVT U88 ( .A(state[104]), .Y(n22) );
  INVX0_HVT U89 ( .A(subkey[59]), .Y(n368) );
  INVX0_HVT U90 ( .A(subkey[58]), .Y(n226) );
  INVX0_HVT U91 ( .A(subkey[123]), .Y(n314) );
  INVX0_HVT U92 ( .A(subkey[64]), .Y(n236) );
  OR2X1_HVT U93 ( .A1(subkey[111]), .A2(n111), .Y(n113) );
  INVX0_HVT U94 ( .A(subkey[4]), .Y(n500) );
  INVX0_HVT U95 ( .A(n461), .Y(n25) );
  INVX0_HVT U96 ( .A(subkey[74]), .Y(n68) );
  INVX0_HVT U97 ( .A(subkey[73]), .Y(n166) );
  INVX0_HVT U98 ( .A(state[86]), .Y(n71) );
  INVX0_HVT U99 ( .A(subkey[28]), .Y(n26) );
  INVX0_HVT U100 ( .A(n151), .Y(n28) );
  INVX0_HVT U101 ( .A(subkey[65]), .Y(n233) );
  INVX0_HVT U102 ( .A(n118), .Y(n29) );
  INVX0_HVT U103 ( .A(n186), .Y(n30) );
  OR2X1_HVT U104 ( .A1(n345), .A2(subkey[79]), .Y(n347) );
  INVX0_HVT U105 ( .A(subkey[32]), .Y(n260) );
  INVX0_HVT U106 ( .A(state[82]), .Y(n330) );
  INVX0_HVT U107 ( .A(subkey[39]), .Y(n399) );
  INVX0_HVT U108 ( .A(n448), .Y(n31) );
  NAND2X0_HVT U109 ( .A1(n104), .A2(state[76]), .Y(n105) );
  INVX0_HVT U110 ( .A(n237), .Y(n33) );
  INVX0_HVT U111 ( .A(n473), .Y(n34) );
  INVX0_HVT U112 ( .A(n167), .Y(n35) );
  INVX0_HVT U113 ( .A(n232), .Y(n36) );
  INVX0_HVT U114 ( .A(state[122]), .Y(n59) );
  INVX0_HVT U115 ( .A(n206), .Y(n38) );
  INVX0_HVT U116 ( .A(state[36]), .Y(n379) );
  OR2X1_HVT U117 ( .A1(subkey[40]), .A2(n288), .Y(n289) );
  INVX0_HVT U118 ( .A(subkey[3]), .Y(n461) );
  INVX0_HVT U119 ( .A(subkey[72]), .Y(n187) );
  NAND2X0_HVT U120 ( .A1(state[88]), .A2(n40), .Y(n41) );
  NAND2X0_HVT U121 ( .A1(n39), .A2(subkey[88]), .Y(n42) );
  NAND2X0_HVT U122 ( .A1(n41), .A2(n42), .Y(out[88]) );
  INVX0_HVT U123 ( .A(state[88]), .Y(n39) );
  OR2X1_HVT U124 ( .A1(n229), .A2(state[51]), .Y(n231) );
  INVX0_HVT U125 ( .A(n436), .Y(n43) );
  INVX0_HVT U126 ( .A(n432), .Y(n44) );
  INVX0_HVT U127 ( .A(subkey[33]), .Y(n441) );
  INVX0_HVT U128 ( .A(subkey[69]), .Y(n432) );
  INVX0_HVT U129 ( .A(subkey[42]), .Y(n183) );
  INVX0_HVT U130 ( .A(subkey[6]), .Y(n375) );
  INVX0_HVT U131 ( .A(subkey[44]), .Y(n163) );
  INVX0_HVT U132 ( .A(subkey[36]), .Y(n478) );
  INVX0_HVT U133 ( .A(state[11]), .Y(n271) );
  INVX0_HVT U134 ( .A(n130), .Y(n45) );
  INVX0_HVT U135 ( .A(subkey[18]), .Y(n49) );
  INVX0_HVT U136 ( .A(state[47]), .Y(n114) );
  INVX0_HVT U137 ( .A(state[29]), .Y(n150) );
  INVX0_HVT U138 ( .A(n217), .Y(n46) );
  INVX0_HVT U139 ( .A(n95), .Y(n47) );
  INVX0_HVT U140 ( .A(n198), .Y(n48) );
  OR2X1_HVT U141 ( .A1(n49), .A2(state[18]), .Y(n342) );
  INVX0_HVT U142 ( .A(n275), .Y(n51) );
  NAND2X0_HVT U143 ( .A1(n177), .A2(n176), .Y(out[10]) );
  INVX0_HVT U144 ( .A(state[32]), .Y(n259) );
  INVX0_HVT U145 ( .A(subkey[87]), .Y(n489) );
  INVX0_HVT U146 ( .A(state[68]), .Y(n158) );
  INVX0_HVT U147 ( .A(state[76]), .Y(n103) );
  INVX0_HVT U148 ( .A(state[84]), .Y(n387) );
  INVX1_HVT U149 ( .A(n313), .Y(n52) );
  INVX0_HVT U150 ( .A(n413), .Y(n53) );
  INVX0_HVT U151 ( .A(subkey[21]), .Y(n281) );
  INVX0_HVT U152 ( .A(subkey[24]), .Y(n452) );
  INVX1_HVT U153 ( .A(subkey[0]), .Y(n170) );
  NAND2X0_HVT U154 ( .A1(state[7]), .A2(n56), .Y(n57) );
  NAND2X0_HVT U155 ( .A1(n55), .A2(subkey[7]), .Y(n58) );
  NAND2X0_HVT U156 ( .A1(n57), .A2(n58), .Y(out[7]) );
  INVX0_HVT U157 ( .A(state[7]), .Y(n55) );
  INVX0_HVT U158 ( .A(subkey[7]), .Y(n56) );
  INVX0_HVT U159 ( .A(state[14]), .Y(n302) );
  INVX0_HVT U160 ( .A(state[110]), .Y(n99) );
  INVX0_HVT U161 ( .A(state[94]), .Y(n268) );
  INVX0_HVT U162 ( .A(subkey[43]), .Y(n476) );
  NAND2X0_HVT U163 ( .A1(state[122]), .A2(n60), .Y(n61) );
  NAND2X0_HVT U164 ( .A1(n59), .A2(subkey[122]), .Y(n62) );
  NAND2X0_HVT U165 ( .A1(n61), .A2(n62), .Y(out[122]) );
  INVX0_HVT U166 ( .A(subkey[122]), .Y(n60) );
  NAND2X0_HVT U167 ( .A1(state[125]), .A2(n64), .Y(n65) );
  NAND2X0_HVT U168 ( .A1(n63), .A2(subkey[125]), .Y(n66) );
  NAND2X0_HVT U169 ( .A1(n65), .A2(n66), .Y(out[125]) );
  INVX0_HVT U170 ( .A(state[125]), .Y(n63) );
  INVX0_HVT U171 ( .A(subkey[45]), .Y(n309) );
  NAND2X0_HVT U172 ( .A1(state[74]), .A2(n68), .Y(n69) );
  NAND2X0_HVT U173 ( .A1(subkey[74]), .A2(n67), .Y(n70) );
  NAND2X0_HVT U174 ( .A1(n69), .A2(n70), .Y(out[74]) );
  INVX0_HVT U175 ( .A(state[74]), .Y(n67) );
  INVX0_HVT U176 ( .A(subkey[19]), .Y(n527) );
  INVX0_HVT U177 ( .A(subkey[34]), .Y(n296) );
  NAND2X0_HVT U178 ( .A1(state[86]), .A2(n72), .Y(n73) );
  NAND2X0_HVT U179 ( .A1(n71), .A2(subkey[86]), .Y(n74) );
  NAND2X0_HVT U180 ( .A1(n73), .A2(n74), .Y(out[86]) );
  INVX1_HVT U181 ( .A(subkey[86]), .Y(n72) );
  INVX0_HVT U182 ( .A(state[16]), .Y(n202) );
  INVX0_HVT U183 ( .A(state[71]), .Y(n444) );
  INVX0_HVT U184 ( .A(state[85]), .Y(n292) );
  INVX0_HVT U185 ( .A(state[10]), .Y(n175) );
  INVX0_HVT U186 ( .A(state[72]), .Y(n186) );
  INVX0_HVT U187 ( .A(subkey[63]), .Y(n468) );
  INVX0_HVT U188 ( .A(state[23]), .Y(n214) );
  INVX0_HVT U189 ( .A(state[77]), .Y(n155) );
  NAND2X0_HVT U190 ( .A1(subkey[5]), .A2(n76), .Y(n77) );
  NAND2X0_HVT U191 ( .A1(n75), .A2(state[5]), .Y(n78) );
  NAND2X0_HVT U192 ( .A1(n78), .A2(n77), .Y(out[5]) );
  INVX0_HVT U193 ( .A(subkey[5]), .Y(n75) );
  INVX0_HVT U194 ( .A(state[5]), .Y(n76) );
  INVX0_HVT U195 ( .A(state[103]), .Y(n217) );
  INVX1_HVT U196 ( .A(state[102]), .Y(n95) );
  NAND2X0_HVT U197 ( .A1(state[70]), .A2(n80), .Y(n81) );
  NAND2X0_HVT U198 ( .A1(n79), .A2(subkey[70]), .Y(n82) );
  NAND2X0_HVT U199 ( .A1(n81), .A2(n82), .Y(out[70]) );
  INVX0_HVT U200 ( .A(state[70]), .Y(n79) );
  INVX0_HVT U201 ( .A(subkey[70]), .Y(n80) );
  NAND2X0_HVT U202 ( .A1(n84), .A2(state[38]), .Y(n85) );
  NAND2X0_HVT U203 ( .A1(n83), .A2(subkey[38]), .Y(n86) );
  NAND2X0_HVT U204 ( .A1(n85), .A2(n86), .Y(out[38]) );
  INVX0_HVT U205 ( .A(state[38]), .Y(n83) );
  INVX0_HVT U206 ( .A(subkey[38]), .Y(n84) );
  INVX0_HVT U207 ( .A(state[66]), .Y(n306) );
  INVX0_HVT U208 ( .A(n174), .Y(n87) );
  INVX0_HVT U209 ( .A(state[93]), .Y(n391) );
  NAND2X0_HVT U210 ( .A1(n89), .A2(state[62]), .Y(n90) );
  NAND2X0_HVT U211 ( .A1(subkey[62]), .A2(n88), .Y(n91) );
  NAND2X0_HVT U212 ( .A1(n90), .A2(n91), .Y(out[62]) );
  INVX0_HVT U213 ( .A(state[62]), .Y(n88) );
  INVX0_HVT U214 ( .A(subkey[62]), .Y(n89) );
  INVX0_HVT U215 ( .A(state[83]), .Y(n437) );
  INVX0_HVT U216 ( .A(state[127]), .Y(n206) );
  NAND2X0_HVT U217 ( .A1(state[1]), .A2(n487), .Y(n93) );
  NAND2X0_HVT U218 ( .A1(n92), .A2(subkey[1]), .Y(n94) );
  NAND2X0_HVT U219 ( .A1(n93), .A2(n94), .Y(out[1]) );
  INVX0_HVT U220 ( .A(state[1]), .Y(n92) );
  NAND2X0_HVT U221 ( .A1(n47), .A2(n96), .Y(n97) );
  NAND2X0_HVT U222 ( .A1(n95), .A2(subkey[102]), .Y(n98) );
  NAND2X0_HVT U223 ( .A1(n97), .A2(n98), .Y(out[102]) );
  INVX0_HVT U224 ( .A(state[40]), .Y(n288) );
  INVX0_HVT U225 ( .A(state[8]), .Y(n146) );
  NAND2X0_HVT U226 ( .A1(state[110]), .A2(n100), .Y(n101) );
  NAND2X0_HVT U227 ( .A1(subkey[110]), .A2(n99), .Y(n102) );
  NAND2X0_HVT U228 ( .A1(n102), .A2(n101), .Y(out[110]) );
  INVX0_HVT U229 ( .A(subkey[110]), .Y(n100) );
  INVX0_HVT U230 ( .A(state[34]), .Y(n295) );
  INVX0_HVT U231 ( .A(state[61]), .Y(n138) );
  NAND2X0_HVT U232 ( .A1(n103), .A2(subkey[76]), .Y(n106) );
  NAND2X0_HVT U233 ( .A1(n105), .A2(n106), .Y(out[76]) );
  INVX0_HVT U234 ( .A(subkey[76]), .Y(n104) );
  NAND2X0_HVT U235 ( .A1(n263), .A2(state[115]), .Y(n108) );
  NAND2X0_HVT U236 ( .A1(n107), .A2(subkey[115]), .Y(n109) );
  NAND2X0_HVT U237 ( .A1(n108), .A2(n109), .Y(out[115]) );
  INVX0_HVT U238 ( .A(state[115]), .Y(n107) );
  OR2X1_HVT U239 ( .A1(n110), .A2(state[100]), .Y(n521) );
  NAND2X0_HVT U240 ( .A1(subkey[111]), .A2(n111), .Y(n112) );
  NAND2X0_HVT U241 ( .A1(n113), .A2(n112), .Y(out[111]) );
  INVX0_HVT U242 ( .A(state[0]), .Y(n171) );
  INVX0_HVT U243 ( .A(state[21]), .Y(n280) );
  NAND2X0_HVT U244 ( .A1(n115), .A2(state[47]), .Y(n116) );
  NAND2X0_HVT U245 ( .A1(subkey[47]), .A2(n114), .Y(n117) );
  NAND2X0_HVT U246 ( .A1(n116), .A2(n117), .Y(out[47]) );
  INVX0_HVT U247 ( .A(subkey[47]), .Y(n115) );
  NAND2X0_HVT U248 ( .A1(n29), .A2(n119), .Y(n120) );
  NAND2X0_HVT U249 ( .A1(state[95]), .A2(n118), .Y(n121) );
  NAND2X0_HVT U250 ( .A1(n120), .A2(n121), .Y(out[95]) );
  INVX0_HVT U251 ( .A(state[45]), .Y(n310) );
  NAND2X0_HVT U252 ( .A1(state[13]), .A2(n123), .Y(n124) );
  NAND2X0_HVT U253 ( .A1(n122), .A2(subkey[13]), .Y(n125) );
  NAND2X0_HVT U254 ( .A1(n124), .A2(n125), .Y(out[13]) );
  INVX0_HVT U255 ( .A(state[13]), .Y(n122) );
  INVX0_HVT U256 ( .A(subkey[13]), .Y(n123) );
  NAND2X0_HVT U257 ( .A1(n16), .A2(n127), .Y(n128) );
  NAND2X0_HVT U258 ( .A1(subkey[78]), .A2(n126), .Y(n129) );
  NAND2X0_HVT U259 ( .A1(n128), .A2(n129), .Y(out[78]) );
  INVX0_HVT U260 ( .A(state[78]), .Y(n126) );
  INVX0_HVT U261 ( .A(subkey[78]), .Y(n127) );
  INVX0_HVT U262 ( .A(state[37]), .Y(n353) );
  INVX0_HVT U263 ( .A(state[50]), .Y(n410) );
  INVX0_HVT U264 ( .A(state[52]), .Y(n465) );
  INVX0_HVT U265 ( .A(subkey[121]), .Y(n513) );
  NAND2X0_HVT U266 ( .A1(n45), .A2(n131), .Y(n132) );
  NAND2X0_HVT U267 ( .A1(subkey[9]), .A2(n130), .Y(n133) );
  NAND2X0_HVT U268 ( .A1(n132), .A2(n133), .Y(out[9]) );
  INVX0_HVT U269 ( .A(subkey[9]), .Y(n131) );
  NAND2X0_HVT U270 ( .A1(subkey[30]), .A2(n135), .Y(n136) );
  NAND2X0_HVT U271 ( .A1(state[30]), .A2(n134), .Y(n137) );
  NAND2X0_HVT U272 ( .A1(n137), .A2(n136), .Y(out[30]) );
  INVX0_HVT U273 ( .A(subkey[30]), .Y(n134) );
  INVX0_HVT U274 ( .A(state[30]), .Y(n135) );
  NAND2X0_HVT U275 ( .A1(n139), .A2(state[61]), .Y(n140) );
  NAND2X0_HVT U276 ( .A1(n138), .A2(subkey[61]), .Y(n141) );
  NAND2X0_HVT U277 ( .A1(n140), .A2(n141), .Y(out[61]) );
  INVX0_HVT U278 ( .A(state[15]), .Y(n425) );
  NAND2X0_HVT U279 ( .A1(state[26]), .A2(n143), .Y(n144) );
  NAND2X0_HVT U280 ( .A1(n142), .A2(subkey[26]), .Y(n145) );
  NAND2X0_HVT U281 ( .A1(n145), .A2(n144), .Y(out[26]) );
  INVX0_HVT U282 ( .A(state[26]), .Y(n142) );
  INVX0_HVT U283 ( .A(subkey[26]), .Y(n143) );
  INVX0_HVT U284 ( .A(state[87]), .Y(n490) );
  INVX0_HVT U285 ( .A(subkey[16]), .Y(n201) );
  INVX1_HVT U286 ( .A(subkey[20]), .Y(n531) );
  INVX0_HVT U287 ( .A(subkey[93]), .Y(n390) );
  NAND2X0_HVT U288 ( .A1(n147), .A2(state[8]), .Y(n148) );
  NAND2X0_HVT U289 ( .A1(n146), .A2(subkey[8]), .Y(n149) );
  NAND2X0_HVT U290 ( .A1(n148), .A2(n149), .Y(out[8]) );
  INVX0_HVT U291 ( .A(subkey[8]), .Y(n147) );
  NAND2X0_HVT U292 ( .A1(state[29]), .A2(n151), .Y(n152) );
  NAND2X0_HVT U293 ( .A1(n28), .A2(n150), .Y(n153) );
  NAND2X0_HVT U294 ( .A1(n152), .A2(n153), .Y(out[29]) );
  INVX0_HVT U295 ( .A(state[65]), .Y(n232) );
  NAND2X0_HVT U296 ( .A1(n155), .A2(subkey[77]), .Y(n156) );
  NAND2X0_HVT U297 ( .A1(state[77]), .A2(n154), .Y(n157) );
  NAND2X0_HVT U298 ( .A1(n157), .A2(n156), .Y(out[77]) );
  INVX0_HVT U299 ( .A(subkey[77]), .Y(n154) );
  INVX0_HVT U300 ( .A(state[64]), .Y(n237) );
  INVX0_HVT U301 ( .A(state[80]), .Y(n524) );
  INVX0_HVT U302 ( .A(state[114]), .Y(n209) );
  NAND2X0_HVT U303 ( .A1(state[68]), .A2(n159), .Y(n160) );
  NAND2X0_HVT U304 ( .A1(subkey[68]), .A2(n158), .Y(n161) );
  NAND2X0_HVT U305 ( .A1(n161), .A2(n160), .Y(out[68]) );
  INVX0_HVT U306 ( .A(subkey[68]), .Y(n159) );
  INVX0_HVT U307 ( .A(state[92]), .Y(n394) );
  NAND2X0_HVT U308 ( .A1(state[44]), .A2(n163), .Y(n164) );
  NAND2X0_HVT U309 ( .A1(n162), .A2(subkey[44]), .Y(n165) );
  NAND2X0_HVT U310 ( .A1(n164), .A2(n165), .Y(out[44]) );
  INVX0_HVT U311 ( .A(state[44]), .Y(n162) );
  NAND2X0_HVT U312 ( .A1(subkey[73]), .A2(n167), .Y(n168) );
  NAND2X0_HVT U313 ( .A1(n35), .A2(n166), .Y(n169) );
  NAND2X0_HVT U314 ( .A1(n169), .A2(n168), .Y(out[73]) );
  NAND2X0_HVT U315 ( .A1(n171), .A2(subkey[0]), .Y(n172) );
  NAND2X0_HVT U316 ( .A1(n170), .A2(state[0]), .Y(n173) );
  NAND2X0_HVT U317 ( .A1(n173), .A2(n172), .Y(out[0]) );
  NAND2X0_HVT U318 ( .A1(n87), .A2(n175), .Y(n176) );
  NAND2X0_HVT U319 ( .A1(state[10]), .A2(n174), .Y(n177) );
  INVX0_HVT U320 ( .A(state[59]), .Y(n367) );
  INVX0_HVT U321 ( .A(state[39]), .Y(n398) );
  NAND2X0_HVT U322 ( .A1(state[60]), .A2(n179), .Y(n180) );
  NAND2X0_HVT U323 ( .A1(subkey[60]), .A2(n178), .Y(n181) );
  NAND2X0_HVT U324 ( .A1(n180), .A2(n181), .Y(out[60]) );
  INVX0_HVT U325 ( .A(state[60]), .Y(n178) );
  INVX0_HVT U326 ( .A(subkey[60]), .Y(n179) );
  INVX0_HVT U327 ( .A(subkey[66]), .Y(n305) );
  NAND2X0_HVT U328 ( .A1(state[42]), .A2(n183), .Y(n184) );
  NAND2X0_HVT U329 ( .A1(subkey[42]), .A2(n182), .Y(n185) );
  NAND2X0_HVT U330 ( .A1(n184), .A2(n185), .Y(out[42]) );
  INVX0_HVT U331 ( .A(subkey[89]), .Y(n517) );
  INVX0_HVT U332 ( .A(state[54]), .Y(n317) );
  INVX0_HVT U333 ( .A(subkey[85]), .Y(n291) );
  NAND2X0_HVT U334 ( .A1(n30), .A2(n187), .Y(n188) );
  NAND2X0_HVT U335 ( .A1(n186), .A2(n7), .Y(n189) );
  NAND2X0_HVT U336 ( .A1(n188), .A2(n189), .Y(out[72]) );
  INVX0_HVT U337 ( .A(state[33]), .Y(n440) );
  NAND2X0_HVT U338 ( .A1(state[4]), .A2(n500), .Y(n191) );
  NAND2X0_HVT U339 ( .A1(subkey[4]), .A2(n190), .Y(n192) );
  NAND2X0_HVT U340 ( .A1(n191), .A2(n192), .Y(out[4]) );
  INVX0_HVT U341 ( .A(state[4]), .Y(n190) );
  NAND2X0_HVT U342 ( .A1(n194), .A2(n4), .Y(n195) );
  NAND2X0_HVT U343 ( .A1(n193), .A2(state[56]), .Y(n196) );
  NAND2X0_HVT U344 ( .A1(n196), .A2(n195), .Y(out[56]) );
  INVX0_HVT U345 ( .A(subkey[56]), .Y(n193) );
  INVX0_HVT U346 ( .A(state[56]), .Y(n194) );
  NAND2X0_HVT U347 ( .A1(subkey[22]), .A2(n198), .Y(n199) );
  NAND2X0_HVT U348 ( .A1(n48), .A2(n197), .Y(n200) );
  NAND2X0_HVT U349 ( .A1(n200), .A2(n199), .Y(out[22]) );
  INVX0_HVT U350 ( .A(subkey[22]), .Y(n197) );
  NAND2X0_HVT U351 ( .A1(subkey[16]), .A2(n202), .Y(n203) );
  NAND2X0_HVT U352 ( .A1(state[16]), .A2(n201), .Y(n204) );
  NAND2X0_HVT U353 ( .A1(n204), .A2(n203), .Y(out[16]) );
  NAND2X0_HVT U354 ( .A1(subkey[127]), .A2(n206), .Y(n207) );
  NAND2X0_HVT U355 ( .A1(n38), .A2(n205), .Y(n208) );
  NAND2X0_HVT U356 ( .A1(n208), .A2(n207), .Y(out[127]) );
  INVX0_HVT U357 ( .A(subkey[127]), .Y(n205) );
  INVX0_HVT U358 ( .A(state[35]), .Y(n506) );
  INVX0_HVT U359 ( .A(state[55]), .Y(n360) );
  INVX0_HVT U360 ( .A(state[24]), .Y(n453) );
  NAND2X0_HVT U361 ( .A1(state[114]), .A2(n244), .Y(n211) );
  NAND2X0_HVT U362 ( .A1(n209), .A2(n210), .Y(n212) );
  NAND2X0_HVT U363 ( .A1(n211), .A2(n212), .Y(out[114]) );
  NAND2X0_HVT U364 ( .A1(subkey[23]), .A2(n214), .Y(n215) );
  NAND2X0_HVT U365 ( .A1(state[23]), .A2(n213), .Y(n216) );
  NAND2X0_HVT U366 ( .A1(n216), .A2(n215), .Y(out[23]) );
  INVX0_HVT U367 ( .A(subkey[23]), .Y(n213) );
  INVX0_HVT U368 ( .A(state[109]), .Y(n320) );
  INVX0_HVT U369 ( .A(subkey[48]), .Y(n248) );
  INVX0_HVT U370 ( .A(state[90]), .Y(n221) );
  NAND2X0_HVT U371 ( .A1(n46), .A2(n218), .Y(n219) );
  NAND2X0_HVT U372 ( .A1(n217), .A2(subkey[103]), .Y(n220) );
  NAND2X0_HVT U373 ( .A1(n219), .A2(n220), .Y(out[103]) );
  NAND2X0_HVT U374 ( .A1(n222), .A2(state[90]), .Y(n223) );
  NAND2X0_HVT U375 ( .A1(n221), .A2(n6), .Y(n224) );
  NAND2X0_HVT U376 ( .A1(n223), .A2(n224), .Y(out[90]) );
  INVX0_HVT U377 ( .A(subkey[90]), .Y(n222) );
  NAND2X0_HVT U378 ( .A1(state[58]), .A2(n226), .Y(n227) );
  NAND2X0_HVT U379 ( .A1(subkey[58]), .A2(n225), .Y(n228) );
  NAND2X0_HVT U380 ( .A1(n227), .A2(n228), .Y(out[58]) );
  NAND2X0_HVT U381 ( .A1(n229), .A2(state[51]), .Y(n230) );
  NAND2X0_HVT U382 ( .A1(n231), .A2(n230), .Y(out[51]) );
  INVX0_HVT U383 ( .A(subkey[51]), .Y(n229) );
  NAND2X0_HVT U384 ( .A1(n36), .A2(n233), .Y(n234) );
  NAND2X0_HVT U385 ( .A1(subkey[65]), .A2(n232), .Y(n235) );
  NAND2X0_HVT U386 ( .A1(n234), .A2(n235), .Y(out[65]) );
  NAND2X0_HVT U387 ( .A1(subkey[64]), .A2(n237), .Y(n238) );
  NAND2X0_HVT U388 ( .A1(n33), .A2(n236), .Y(n239) );
  NAND2X0_HVT U389 ( .A1(n239), .A2(n238), .Y(out[64]) );
  INVX0_HVT U390 ( .A(state[46]), .Y(n324) );
  INVX0_HVT U391 ( .A(subkey[35]), .Y(n505) );
  NAND2X0_HVT U392 ( .A1(state[57]), .A2(n299), .Y(n242) );
  NAND2X0_HVT U393 ( .A1(n241), .A2(n240), .Y(n243) );
  NAND2X0_HVT U394 ( .A1(n242), .A2(n243), .Y(out[57]) );
  INVX0_HVT U395 ( .A(state[57]), .Y(n240) );
  INVX0_HVT U396 ( .A(n299), .Y(n241) );
  INVX0_HVT U397 ( .A(state[126]), .Y(n349) );
  NAND2X0_HVT U398 ( .A1(n245), .A2(subkey[119]), .Y(n247) );
  NAND2X0_HVT U399 ( .A1(n246), .A2(n247), .Y(out[119]) );
  INVX0_HVT U400 ( .A(state[119]), .Y(n245) );
  NAND2X0_HVT U401 ( .A1(subkey[48]), .A2(n249), .Y(n250) );
  NAND2X0_HVT U402 ( .A1(state[48]), .A2(n248), .Y(n251) );
  NAND2X0_HVT U403 ( .A1(n251), .A2(n250), .Y(out[48]) );
  INVX0_HVT U404 ( .A(state[48]), .Y(n249) );
  INVX0_HVT U405 ( .A(state[75]), .Y(n536) );
  NAND2X0_HVT U406 ( .A1(n253), .A2(state[101]), .Y(n254) );
  NAND2X0_HVT U407 ( .A1(n252), .A2(subkey[101]), .Y(n255) );
  NAND2X0_HVT U408 ( .A1(n254), .A2(n255), .Y(out[101]) );
  INVX0_HVT U409 ( .A(state[101]), .Y(n252) );
  INVX0_HVT U410 ( .A(state[6]), .Y(n376) );
  NAND2X0_HVT U411 ( .A1(n300), .A2(state[113]), .Y(n257) );
  NAND2X0_HVT U412 ( .A1(n256), .A2(subkey[113]), .Y(n258) );
  NAND2X0_HVT U413 ( .A1(n257), .A2(n258), .Y(out[113]) );
  INVX0_HVT U414 ( .A(state[113]), .Y(n256) );
  INVX0_HVT U415 ( .A(state[108]), .Y(n363) );
  NAND2X0_HVT U416 ( .A1(state[32]), .A2(n260), .Y(n261) );
  NAND2X0_HVT U417 ( .A1(n259), .A2(subkey[32]), .Y(n262) );
  NAND2X0_HVT U418 ( .A1(n261), .A2(n262), .Y(out[32]) );
  NAND2X0_HVT U419 ( .A1(n279), .A2(state[97]), .Y(n265) );
  NAND2X0_HVT U420 ( .A1(n264), .A2(subkey[97]), .Y(n266) );
  NAND2X0_HVT U421 ( .A1(n265), .A2(n266), .Y(out[97]) );
  INVX0_HVT U422 ( .A(state[97]), .Y(n264) );
  INVX0_HVT U423 ( .A(state[123]), .Y(n313) );
  INVX0_HVT U424 ( .A(subkey[92]), .Y(n395) );
  NAND2X0_HVT U425 ( .A1(subkey[94]), .A2(n268), .Y(n269) );
  NAND2X0_HVT U426 ( .A1(state[94]), .A2(n267), .Y(n270) );
  NAND2X0_HVT U427 ( .A1(n270), .A2(n269), .Y(out[94]) );
  INVX0_HVT U428 ( .A(subkey[94]), .Y(n267) );
  NAND2X0_HVT U429 ( .A1(n272), .A2(state[11]), .Y(n273) );
  NAND2X0_HVT U430 ( .A1(subkey[11]), .A2(n271), .Y(n274) );
  NAND2X0_HVT U431 ( .A1(n273), .A2(n274), .Y(out[11]) );
  INVX0_HVT U432 ( .A(state[98]), .Y(n327) );
  NAND2X0_HVT U433 ( .A1(n51), .A2(n276), .Y(n277) );
  NAND2X0_HVT U434 ( .A1(subkey[17]), .A2(n275), .Y(n278) );
  NAND2X0_HVT U435 ( .A1(n277), .A2(n278), .Y(out[17]) );
  INVX0_HVT U436 ( .A(subkey[17]), .Y(n276) );
  NAND2X0_HVT U437 ( .A1(state[21]), .A2(n281), .Y(n282) );
  NAND2X0_HVT U438 ( .A1(n280), .A2(n3), .Y(n283) );
  NAND2X0_HVT U439 ( .A1(n282), .A2(n283), .Y(out[21]) );
  NAND2X0_HVT U440 ( .A1(n285), .A2(subkey[117]), .Y(n286) );
  NAND2X0_HVT U441 ( .A1(state[117]), .A2(n284), .Y(n287) );
  NAND2X0_HVT U442 ( .A1(n287), .A2(n286), .Y(out[117]) );
  INVX0_HVT U443 ( .A(state[117]), .Y(n285) );
  NAND2X0_HVT U444 ( .A1(subkey[40]), .A2(n288), .Y(n290) );
  NAND2X0_HVT U445 ( .A1(n289), .A2(n290), .Y(out[40]) );
  INVX0_HVT U446 ( .A(state[121]), .Y(n514) );
  NAND2X0_HVT U447 ( .A1(n292), .A2(subkey[85]), .Y(n293) );
  NAND2X0_HVT U448 ( .A1(state[85]), .A2(n291), .Y(n294) );
  NAND2X0_HVT U449 ( .A1(n294), .A2(n293), .Y(out[85]) );
  NAND2X0_HVT U450 ( .A1(state[34]), .A2(n296), .Y(n297) );
  NAND2X0_HVT U451 ( .A1(n295), .A2(subkey[34]), .Y(n298) );
  NAND2X0_HVT U452 ( .A1(n297), .A2(n298), .Y(out[34]) );
  INVX0_HVT U453 ( .A(state[69]), .Y(n433) );
  NAND2X0_HVT U454 ( .A1(n302), .A2(subkey[14]), .Y(n303) );
  NAND2X0_HVT U455 ( .A1(n301), .A2(state[14]), .Y(n304) );
  NAND2X0_HVT U456 ( .A1(n304), .A2(n303), .Y(out[14]) );
  INVX0_HVT U457 ( .A(state[53]), .Y(n406) );
  INVX0_HVT U458 ( .A(state[96]), .Y(n335) );
  NAND2X0_HVT U459 ( .A1(n306), .A2(n5), .Y(n307) );
  NAND2X0_HVT U460 ( .A1(state[66]), .A2(n305), .Y(n308) );
  NAND2X0_HVT U461 ( .A1(n308), .A2(n307), .Y(out[66]) );
  NAND2X0_HVT U462 ( .A1(n310), .A2(subkey[45]), .Y(n311) );
  NAND2X0_HVT U463 ( .A1(state[45]), .A2(n309), .Y(n312) );
  NAND2X0_HVT U464 ( .A1(n312), .A2(n311), .Y(out[45]) );
  INVX0_HVT U465 ( .A(state[89]), .Y(n518) );
  INVX0_HVT U466 ( .A(state[19]), .Y(n528) );
  NAND2X0_HVT U467 ( .A1(n52), .A2(n314), .Y(n315) );
  NAND2X0_HVT U468 ( .A1(n313), .A2(subkey[123]), .Y(n316) );
  NAND2X0_HVT U469 ( .A1(n315), .A2(n316), .Y(out[123]) );
  NAND2X0_HVT U470 ( .A1(subkey[54]), .A2(n317), .Y(n318) );
  NAND2X0_HVT U471 ( .A1(n319), .A2(n318), .Y(out[54]) );
  INVX0_HVT U472 ( .A(state[79]), .Y(n345) );
  NAND2X0_HVT U473 ( .A1(state[109]), .A2(n321), .Y(n322) );
  NAND2X0_HVT U474 ( .A1(n320), .A2(subkey[109]), .Y(n323) );
  NAND2X0_HVT U475 ( .A1(n322), .A2(n323), .Y(out[109]) );
  NAND2X0_HVT U476 ( .A1(n324), .A2(subkey[46]), .Y(n326) );
  NAND2X0_HVT U477 ( .A1(n325), .A2(n326), .Y(out[46]) );
  INVX0_HVT U478 ( .A(state[107]), .Y(n382) );
  NAND2X0_HVT U479 ( .A1(n327), .A2(subkey[98]), .Y(n328) );
  NAND2X0_HVT U480 ( .A1(n329), .A2(n328), .Y(out[98]) );
  INVX0_HVT U481 ( .A(state[91]), .Y(n456) );
  INVX0_HVT U482 ( .A(subkey[52]), .Y(n464) );
  INVX0_HVT U483 ( .A(state[124]), .Y(n371) );
  INVX1_HVT U484 ( .A(subkey[55]), .Y(n359) );
  NAND2X0_HVT U485 ( .A1(n331), .A2(state[82]), .Y(n332) );
  NAND2X0_HVT U486 ( .A1(n330), .A2(subkey[82]), .Y(n333) );
  NAND2X0_HVT U487 ( .A1(n333), .A2(n332), .Y(out[82]) );
  INVX0_HVT U488 ( .A(subkey[82]), .Y(n331) );
  NAND2X0_HVT U489 ( .A1(subkey[96]), .A2(n335), .Y(n336) );
  NAND2X0_HVT U490 ( .A1(state[96]), .A2(n334), .Y(n337) );
  NAND2X0_HVT U491 ( .A1(n337), .A2(n336), .Y(out[96]) );
  NAND2X0_HVT U492 ( .A1(n339), .A2(subkey[41]), .Y(n340) );
  NAND2X0_HVT U493 ( .A1(state[41]), .A2(n338), .Y(n341) );
  NAND2X0_HVT U494 ( .A1(n341), .A2(n340), .Y(out[41]) );
  INVX0_HVT U495 ( .A(subkey[41]), .Y(n338) );
  NAND2X0_HVT U496 ( .A1(n49), .A2(state[18]), .Y(n343) );
  NAND2X0_HVT U497 ( .A1(n342), .A2(n343), .Y(out[18]) );
  INVX0_HVT U498 ( .A(state[31]), .Y(n421) );
  NAND2X0_HVT U499 ( .A1(subkey[79]), .A2(n345), .Y(n346) );
  NAND2X0_HVT U500 ( .A1(n346), .A2(n347), .Y(out[79]) );
  NAND2X0_HVT U501 ( .A1(subkey[126]), .A2(n349), .Y(n350) );
  NAND2X0_HVT U502 ( .A1(state[126]), .A2(n348), .Y(n351) );
  NAND2X0_HVT U503 ( .A1(n351), .A2(n350), .Y(out[126]) );
  NAND2X0_HVT U504 ( .A1(subkey[37]), .A2(n353), .Y(n354) );
  NAND2X0_HVT U505 ( .A1(n352), .A2(state[37]), .Y(n355) );
  NAND2X0_HVT U506 ( .A1(n355), .A2(n354), .Y(out[37]) );
  INVX0_HVT U507 ( .A(subkey[37]), .Y(n352) );
  NAND2X0_HVT U508 ( .A1(state[112]), .A2(n477), .Y(n357) );
  NAND2X0_HVT U509 ( .A1(n356), .A2(subkey[112]), .Y(n358) );
  NAND2X0_HVT U510 ( .A1(n357), .A2(n358), .Y(out[112]) );
  INVX0_HVT U511 ( .A(state[112]), .Y(n356) );
  INVX0_HVT U512 ( .A(state[116]), .Y(n479) );
  NAND2X0_HVT U513 ( .A1(n360), .A2(subkey[55]), .Y(n361) );
  NAND2X0_HVT U514 ( .A1(state[55]), .A2(n359), .Y(n362) );
  NAND2X0_HVT U515 ( .A1(n362), .A2(n361), .Y(out[55]) );
  NAND2X0_HVT U516 ( .A1(state[108]), .A2(n364), .Y(n365) );
  NAND2X0_HVT U517 ( .A1(n363), .A2(subkey[108]), .Y(n366) );
  NAND2X0_HVT U518 ( .A1(n365), .A2(n366), .Y(out[108]) );
  INVX0_HVT U519 ( .A(state[28]), .Y(n497) );
  NAND2X0_HVT U520 ( .A1(state[59]), .A2(n368), .Y(n369) );
  NAND2X0_HVT U521 ( .A1(n367), .A2(subkey[59]), .Y(n370) );
  NAND2X0_HVT U522 ( .A1(n369), .A2(n370), .Y(out[59]) );
  NAND2X0_HVT U523 ( .A1(n21), .A2(n372), .Y(n373) );
  NAND2X0_HVT U524 ( .A1(n371), .A2(subkey[124]), .Y(n374) );
  NAND2X0_HVT U525 ( .A1(n373), .A2(n374), .Y(out[124]) );
  NAND2X0_HVT U526 ( .A1(subkey[6]), .A2(n376), .Y(n377) );
  NAND2X0_HVT U527 ( .A1(state[6]), .A2(n375), .Y(n378) );
  NAND2X0_HVT U528 ( .A1(n378), .A2(n377), .Y(out[6]) );
  NAND2X0_HVT U529 ( .A1(n478), .A2(state[36]), .Y(n380) );
  NAND2X0_HVT U530 ( .A1(n379), .A2(subkey[36]), .Y(n381) );
  NAND2X0_HVT U531 ( .A1(n380), .A2(n381), .Y(out[36]) );
  NAND2X0_HVT U532 ( .A1(state[107]), .A2(n383), .Y(n384) );
  NAND2X0_HVT U533 ( .A1(subkey[107]), .A2(n382), .Y(n385) );
  NAND2X0_HVT U534 ( .A1(n385), .A2(n384), .Y(out[107]) );
  INVX0_HVT U535 ( .A(subkey[15]), .Y(n424) );
  NAND2X0_HVT U536 ( .A1(n387), .A2(subkey[84]), .Y(n388) );
  NAND2X0_HVT U537 ( .A1(state[84]), .A2(n386), .Y(n389) );
  NAND2X0_HVT U538 ( .A1(n389), .A2(n388), .Y(out[84]) );
  INVX0_HVT U539 ( .A(subkey[84]), .Y(n386) );
  INVX0_HVT U540 ( .A(state[120]), .Y(n494) );
  NAND2X0_HVT U541 ( .A1(subkey[93]), .A2(n391), .Y(n392) );
  NAND2X0_HVT U542 ( .A1(state[93]), .A2(n390), .Y(n393) );
  NAND2X0_HVT U543 ( .A1(n392), .A2(n393), .Y(out[93]) );
  NAND2X0_HVT U544 ( .A1(n54), .A2(n395), .Y(n396) );
  NAND2X0_HVT U545 ( .A1(n394), .A2(subkey[92]), .Y(n397) );
  NAND2X0_HVT U546 ( .A1(n396), .A2(n397), .Y(out[92]) );
  NAND2X0_HVT U547 ( .A1(n399), .A2(state[39]), .Y(n400) );
  NAND2X0_HVT U548 ( .A1(n398), .A2(subkey[39]), .Y(n401) );
  NAND2X0_HVT U549 ( .A1(n400), .A2(n401), .Y(out[39]) );
  NAND2X0_HVT U550 ( .A1(state[43]), .A2(n476), .Y(n403) );
  NAND2X0_HVT U551 ( .A1(n402), .A2(subkey[43]), .Y(n404) );
  NAND2X0_HVT U552 ( .A1(n404), .A2(n403), .Y(out[43]) );
  INVX0_HVT U553 ( .A(state[43]), .Y(n402) );
  INVX0_HVT U554 ( .A(subkey[53]), .Y(n405) );
  NAND2X0_HVT U555 ( .A1(n406), .A2(subkey[53]), .Y(n407) );
  NAND2X0_HVT U556 ( .A1(n405), .A2(state[53]), .Y(n408) );
  NAND2X0_HVT U557 ( .A1(n408), .A2(n407), .Y(out[53]) );
  NAND2X0_HVT U558 ( .A1(subkey[50]), .A2(n410), .Y(n411) );
  NAND2X0_HVT U559 ( .A1(state[50]), .A2(n409), .Y(n412) );
  NAND2X0_HVT U560 ( .A1(n411), .A2(n412), .Y(out[50]) );
  INVX0_HVT U561 ( .A(state[67]), .Y(n509) );
  NAND2X0_HVT U562 ( .A1(n53), .A2(n414), .Y(n415) );
  NAND2X0_HVT U563 ( .A1(subkey[49]), .A2(n413), .Y(n416) );
  NAND2X0_HVT U564 ( .A1(n415), .A2(n416), .Y(out[49]) );
  INVX0_HVT U565 ( .A(subkey[49]), .Y(n414) );
  NAND2X0_HVT U566 ( .A1(state[12]), .A2(n418), .Y(n419) );
  NAND2X0_HVT U567 ( .A1(subkey[12]), .A2(n417), .Y(n420) );
  NAND2X0_HVT U568 ( .A1(n419), .A2(n420), .Y(out[12]) );
  INVX0_HVT U569 ( .A(state[12]), .Y(n417) );
  INVX0_HVT U570 ( .A(subkey[12]), .Y(n418) );
  INVX0_HVT U571 ( .A(subkey[80]), .Y(n523) );
  INVX0_HVT U572 ( .A(subkey[67]), .Y(n510) );
  INVX0_HVT U573 ( .A(subkey[83]), .Y(n436) );
  NAND2X0_HVT U574 ( .A1(subkey[31]), .A2(n421), .Y(n423) );
  NAND2X0_HVT U575 ( .A1(n422), .A2(n423), .Y(out[31]) );
  INVX0_HVT U576 ( .A(state[27]), .Y(n472) );
  NAND2X0_HVT U577 ( .A1(n8), .A2(n425), .Y(n426) );
  NAND2X0_HVT U578 ( .A1(state[15]), .A2(n424), .Y(n427) );
  NAND2X0_HVT U579 ( .A1(n427), .A2(n426), .Y(out[15]) );
  INVX0_HVT U580 ( .A(state[105]), .Y(n502) );
  INVX0_HVT U581 ( .A(state[3]), .Y(n460) );
  NAND2X0_HVT U582 ( .A1(subkey[81]), .A2(n429), .Y(n430) );
  NAND2X0_HVT U583 ( .A1(n428), .A2(state[81]), .Y(n431) );
  NAND2X0_HVT U584 ( .A1(n431), .A2(n430), .Y(out[81]) );
  INVX0_HVT U585 ( .A(subkey[81]), .Y(n428) );
  INVX0_HVT U586 ( .A(state[81]), .Y(n429) );
  NAND2X0_HVT U587 ( .A1(n44), .A2(n433), .Y(n434) );
  NAND2X0_HVT U588 ( .A1(state[69]), .A2(n432), .Y(n435) );
  NAND2X0_HVT U589 ( .A1(n435), .A2(n434), .Y(out[69]) );
  NAND2X0_HVT U590 ( .A1(n43), .A2(n437), .Y(n438) );
  NAND2X0_HVT U591 ( .A1(state[83]), .A2(n436), .Y(n439) );
  NAND2X0_HVT U592 ( .A1(n439), .A2(n438), .Y(out[83]) );
  NAND2X0_HVT U593 ( .A1(state[33]), .A2(n441), .Y(n442) );
  NAND2X0_HVT U594 ( .A1(n440), .A2(subkey[33]), .Y(n443) );
  NAND2X0_HVT U595 ( .A1(n442), .A2(n443), .Y(out[33]) );
  NAND2X0_HVT U596 ( .A1(state[71]), .A2(n445), .Y(n446) );
  NAND2X0_HVT U597 ( .A1(subkey[71]), .A2(n444), .Y(n447) );
  NAND2X0_HVT U598 ( .A1(n446), .A2(n447), .Y(out[71]) );
  NAND2X0_HVT U599 ( .A1(n31), .A2(n449), .Y(n450) );
  NAND2X0_HVT U600 ( .A1(n448), .A2(subkey[25]), .Y(n451) );
  NAND2X0_HVT U601 ( .A1(n450), .A2(n451), .Y(out[25]) );
  NAND2X0_HVT U602 ( .A1(subkey[24]), .A2(n453), .Y(n454) );
  NAND2X0_HVT U603 ( .A1(state[24]), .A2(n452), .Y(n455) );
  NAND2X0_HVT U604 ( .A1(n455), .A2(n454), .Y(out[24]) );
  INVX0_HVT U605 ( .A(state[99]), .Y(n484) );
  NAND2X0_HVT U606 ( .A1(state[91]), .A2(n457), .Y(n458) );
  NAND2X0_HVT U607 ( .A1(n456), .A2(subkey[91]), .Y(n459) );
  NAND2X0_HVT U608 ( .A1(n458), .A2(n459), .Y(out[91]) );
  NAND2X0_HVT U609 ( .A1(state[3]), .A2(n461), .Y(n462) );
  NAND2X0_HVT U610 ( .A1(n25), .A2(n460), .Y(n463) );
  NAND2X0_HVT U611 ( .A1(n462), .A2(n463), .Y(out[3]) );
  NAND2X0_HVT U612 ( .A1(subkey[52]), .A2(n465), .Y(n466) );
  NAND2X0_HVT U613 ( .A1(n37), .A2(n464), .Y(n467) );
  NAND2X0_HVT U614 ( .A1(n467), .A2(n466), .Y(out[52]) );
  NAND2X0_HVT U615 ( .A1(subkey[63]), .A2(n469), .Y(n470) );
  NAND2X0_HVT U616 ( .A1(state[63]), .A2(n468), .Y(n471) );
  NAND2X0_HVT U617 ( .A1(n471), .A2(n470), .Y(out[63]) );
  INVX0_HVT U618 ( .A(state[63]), .Y(n469) );
  NAND2X0_HVT U619 ( .A1(state[27]), .A2(n473), .Y(n474) );
  NAND2X0_HVT U620 ( .A1(n34), .A2(n472), .Y(n475) );
  NAND2X0_HVT U621 ( .A1(n474), .A2(n475), .Y(out[27]) );
  NAND2X0_HVT U622 ( .A1(state[116]), .A2(n480), .Y(n481) );
  NAND2X0_HVT U623 ( .A1(subkey[116]), .A2(n479), .Y(n482) );
  NAND2X0_HVT U624 ( .A1(n481), .A2(n482), .Y(out[116]) );
  NAND2X0_HVT U625 ( .A1(subkey[99]), .A2(n484), .Y(n485) );
  NAND2X0_HVT U626 ( .A1(n483), .A2(state[99]), .Y(n486) );
  NAND2X0_HVT U627 ( .A1(n486), .A2(n485), .Y(out[99]) );
  NAND2X0_HVT U628 ( .A1(subkey[87]), .A2(n490), .Y(n491) );
  NAND2X0_HVT U629 ( .A1(state[87]), .A2(n489), .Y(n492) );
  NAND2X0_HVT U630 ( .A1(n492), .A2(n491), .Y(out[87]) );
  NAND2X0_HVT U631 ( .A1(subkey[120]), .A2(n494), .Y(n495) );
  NAND2X0_HVT U632 ( .A1(state[120]), .A2(n493), .Y(n496) );
  NAND2X0_HVT U633 ( .A1(n496), .A2(n495), .Y(out[120]) );
  NAND2X0_HVT U634 ( .A1(n497), .A2(subkey[28]), .Y(n498) );
  NAND2X0_HVT U635 ( .A1(n26), .A2(state[28]), .Y(n499) );
  NAND2X0_HVT U636 ( .A1(n499), .A2(n498), .Y(out[28]) );
  NAND2X0_HVT U637 ( .A1(subkey[105]), .A2(n502), .Y(n503) );
  NAND2X0_HVT U638 ( .A1(state[105]), .A2(n501), .Y(n504) );
  NAND2X0_HVT U639 ( .A1(n504), .A2(n503), .Y(out[105]) );
  NAND2X0_HVT U640 ( .A1(subkey[35]), .A2(n506), .Y(n507) );
  NAND2X0_HVT U641 ( .A1(n505), .A2(state[35]), .Y(n508) );
  NAND2X0_HVT U642 ( .A1(n508), .A2(n507), .Y(out[35]) );
  NAND2X0_HVT U643 ( .A1(state[67]), .A2(n510), .Y(n511) );
  NAND2X0_HVT U644 ( .A1(n509), .A2(subkey[67]), .Y(n512) );
  NAND2X0_HVT U645 ( .A1(n511), .A2(n512), .Y(out[67]) );
  NAND2X0_HVT U646 ( .A1(n2), .A2(n514), .Y(n515) );
  NAND2X0_HVT U647 ( .A1(state[121]), .A2(n513), .Y(n516) );
  NAND2X0_HVT U648 ( .A1(n516), .A2(n515), .Y(out[121]) );
  NAND2X0_HVT U649 ( .A1(n1), .A2(n518), .Y(n519) );
  NAND2X0_HVT U650 ( .A1(state[89]), .A2(n517), .Y(n520) );
  NAND2X0_HVT U651 ( .A1(n520), .A2(n519), .Y(out[89]) );
  INVX0_HVT U652 ( .A(state[20]), .Y(n532) );
  NAND2X0_HVT U653 ( .A1(n110), .A2(state[100]), .Y(n522) );
  NAND2X0_HVT U654 ( .A1(n521), .A2(n522), .Y(out[100]) );
  NAND2X0_HVT U655 ( .A1(subkey[80]), .A2(n524), .Y(n525) );
  NAND2X0_HVT U656 ( .A1(n523), .A2(state[80]), .Y(n526) );
  NAND2X0_HVT U657 ( .A1(n526), .A2(n525), .Y(out[80]) );
  NAND2X0_HVT U658 ( .A1(subkey[19]), .A2(n528), .Y(n529) );
  NAND2X0_HVT U659 ( .A1(n527), .A2(state[19]), .Y(n530) );
  NAND2X0_HVT U660 ( .A1(n530), .A2(n529), .Y(out[19]) );
  NAND2X0_HVT U661 ( .A1(subkey[20]), .A2(n532), .Y(n533) );
  NAND2X0_HVT U662 ( .A1(n32), .A2(n531), .Y(n534) );
  NAND2X0_HVT U663 ( .A1(n534), .A2(n533), .Y(out[20]) );
  NAND2X0_HVT U664 ( .A1(n536), .A2(n9), .Y(n537) );
  NAND2X0_HVT U665 ( .A1(state[75]), .A2(n535), .Y(n538) );
  NAND2X0_HVT U666 ( .A1(n538), .A2(n537), .Y(out[75]) );
endmodule

