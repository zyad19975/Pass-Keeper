
module sbox_3 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n19, n23, n48, n50, n210, n211, n212, n213, n216, n217, n218, n219,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631;

  NAND2X0_HVT U4 ( .A1(n339), .A2(n271), .Y(n628) );
  NAND2X0_HVT U5 ( .A1(n346), .A2(n293), .Y(n626) );
  NAND2X0_HVT U13 ( .A1(n618), .A2(n344), .Y(n619) );
  NAND2X0_HVT U21 ( .A1(n338), .A2(n350), .Y(n611) );
  NAND2X0_HVT U24 ( .A1(n335), .A2(n350), .Y(n609) );
  NAND2X0_HVT U33 ( .A1(n408), .A2(n350), .Y(n600) );
  NAND2X0_HVT U35 ( .A1(n333), .A2(n350), .Y(n598) );
  NAND2X0_HVT U42 ( .A1(n347), .A2(n335), .Y(n591) );
  NAND2X0_HVT U53 ( .A1(n581), .A2(n590), .Y(n582) );
  NAND2X0_HVT U56 ( .A1(n339), .A2(n577), .Y(n578) );
  MUX41X1_HVT U57 ( .A1(n397), .A3(n613), .A2(n578), .A4(n621), .S0(n353), 
        .S1(n352), .Y(n576) );
  NAND2X0_HVT U58 ( .A1(n344), .A2(n272), .Y(n575) );
  MUX41X1_HVT U59 ( .A1(n319), .A3(n575), .A2(n317), .A4(n304), .S0(n353), 
        .S1(in[5]), .Y(n574) );
  MUX41X1_HVT U61 ( .A1(n316), .A3(n372), .A2(n371), .A4(n330), .S0(n353), 
        .S1(in[5]), .Y(n572) );
  NAND2X0_HVT U62 ( .A1(n350), .A2(n342), .Y(n571) );
  MUX41X1_HVT U63 ( .A1(n571), .A3(n260), .A2(n391), .A4(n370), .S0(n353), 
        .S1(in[5]), .Y(n570) );
  AO21X1_HVT U66 ( .A1(n368), .A2(n326), .A3(n390), .Y(n567) );
  MUX41X1_HVT U68 ( .A1(n366), .A3(n567), .A2(n566), .A4(n568), .S0(n320), 
        .S1(n328), .Y(n565) );
  MUX41X1_HVT U69 ( .A1(n565), .A3(n573), .A2(n569), .A4(n579), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n336), .A2(n560), .Y(n561) );
  MUX41X1_HVT U74 ( .A1(n562), .A3(n607), .A2(n561), .A4(n609), .S0(n322), 
        .S1(n354), .Y(n559) );
  MUX41X1_HVT U75 ( .A1(n394), .A3(n399), .A2(n412), .A4(n375), .S0(n320), 
        .S1(n327), .Y(n558) );
  MUX41X1_HVT U77 ( .A1(n623), .A3(n401), .A2(n557), .A4(n400), .S0(n327), 
        .S1(n351), .Y(n556) );
  MUX41X1_HVT U78 ( .A1(n556), .A3(n559), .A2(n558), .A4(n563), .S0(in[0]), 
        .S1(n352), .Y(n555) );
  AND3X1_HVT U80 ( .A1(n341), .A2(n577), .A3(n552), .Y(n553) );
  AND2X1_HVT U83 ( .A1(n278), .A2(n251), .Y(n549) );
  MUX41X1_HVT U84 ( .A1(n374), .A3(n625), .A2(n615), .A4(n549), .S0(n320), 
        .S1(n255), .Y(n548) );
  NAND2X0_HVT U85 ( .A1(n350), .A2(n411), .Y(n547) );
  MUX41X1_HVT U86 ( .A1(n399), .A3(n547), .A2(n314), .A4(n312), .S0(n320), 
        .S1(n255), .Y(n546) );
  AO21X1_HVT U93 ( .A1(n329), .A2(n539), .A3(n395), .Y(n540) );
  MUX41X1_HVT U96 ( .A1(n358), .A3(n315), .A2(n398), .A4(n537), .S0(n320), 
        .S1(n255), .Y(n536) );
  MUX41X1_HVT U97 ( .A1(n394), .A3(n315), .A2(n346), .A4(n616), .S0(n320), 
        .S1(n255), .Y(n535) );
  MUX41X1_HVT U98 ( .A1(n535), .A3(n538), .A2(n536), .A4(n543), .S0(in[0]), 
        .S1(n352), .Y(n534) );
  NAND2X0_HVT U101 ( .A1(n530), .A2(n529), .Y(n531) );
  MUX41X1_HVT U103 ( .A1(n271), .A3(n367), .A2(n378), .A4(n598), .S0(n320), 
        .S1(n255), .Y(n527) );
  MUX41X1_HVT U105 ( .A1(n377), .A3(n586), .A2(n526), .A4(n393), .S0(n320), 
        .S1(n255), .Y(n525) );
  OA21X1_HVT U109 ( .A1(n385), .A2(n263), .A3(n304), .Y(n522) );
  NAND2X0_HVT U110 ( .A1(n341), .A2(n520), .Y(n521) );
  MUX41X1_HVT U114 ( .A1(n517), .A3(n523), .A2(n519), .A4(n522), .S0(n326), 
        .S1(n255), .Y(n516) );
  AND2X1_HVT U115 ( .A1(n346), .A2(n330), .Y(n515) );
  MUX41X1_HVT U116 ( .A1(n619), .A3(n515), .A2(n375), .A4(n602), .S0(n321), 
        .S1(n353), .Y(n514) );
  NAND2X0_HVT U123 ( .A1(n506), .A2(n505), .Y(n507) );
  MUX41X1_HVT U125 ( .A1(n611), .A3(n319), .A2(n366), .A4(n403), .S0(n321), 
        .S1(n353), .Y(n503) );
  MUX41X1_HVT U131 ( .A1(n498), .A3(n500), .A2(n499), .A4(n501), .S0(n326), 
        .S1(n353), .Y(n497) );
  MUX41X1_HVT U136 ( .A1(n312), .A3(n600), .A2(n405), .A4(n597), .S0(n321), 
        .S1(n353), .Y(n493) );
  AND2X1_HVT U140 ( .A1(n336), .A2(n349), .Y(n489) );
  MUX41X1_HVT U141 ( .A1(n608), .A3(n386), .A2(n489), .A4(n382), .S0(n322), 
        .S1(n353), .Y(n488) );
  MUX41X1_HVT U142 ( .A1(n374), .A3(n330), .A2(n392), .A4(n622), .S0(n321), 
        .S1(n353), .Y(n487) );
  OA21X1_HVT U144 ( .A1(n361), .A2(n231), .A3(n602), .Y(n485) );
  NAND2X0_HVT U146 ( .A1(n249), .A2(n344), .Y(n560) );
  MUX41X1_HVT U147 ( .A1(n405), .A3(n560), .A2(n394), .A4(n587), .S0(n322), 
        .S1(n353), .Y(n483) );
  MUX41X1_HVT U148 ( .A1(n483), .A3(n487), .A2(n484), .A4(n488), .S0(in[0]), 
        .S1(in[5]), .Y(n482) );
  OA21X1_HVT U151 ( .A1(n593), .A2(n231), .A3(n479), .Y(n480) );
  MUX41X1_HVT U153 ( .A1(n521), .A3(n316), .A2(n340), .A4(n360), .S0(n321), 
        .S1(n255), .Y(n477) );
  AND2X1_HVT U154 ( .A1(n329), .A2(n335), .Y(n476) );
  NAND2X0_HVT U158 ( .A1(n346), .A2(n411), .Y(n472) );
  MUX41X1_HVT U159 ( .A1(n619), .A3(n330), .A2(n472), .A4(n365), .S0(n248), 
        .S1(n255), .Y(n471) );
  AND2X1_HVT U162 ( .A1(n625), .A2(n560), .Y(n468) );
  MUX41X1_HVT U163 ( .A1(n372), .A3(n468), .A2(n313), .A4(n469), .S0(n248), 
        .S1(n255), .Y(n467) );
  NAND2X0_HVT U166 ( .A1(n344), .A2(n577), .Y(n464) );
  NAND2X0_HVT U167 ( .A1(n412), .A2(n350), .Y(n463) );
  MUX41X1_HVT U168 ( .A1(n397), .A3(n622), .A2(n463), .A4(n464), .S0(n248), 
        .S1(n354), .Y(n462) );
  OA21X1_HVT U170 ( .A1(n317), .A2(n219), .A3(n602), .Y(n460) );
  NAND2X0_HVT U174 ( .A1(n347), .A2(n625), .Y(n618) );
  NAND2X0_HVT U177 ( .A1(n348), .A2(n332), .Y(n455) );
  MUX41X1_HVT U178 ( .A1(n614), .A3(n455), .A2(n406), .A4(n595), .S0(n322), 
        .S1(n327), .Y(n454) );
  MUX41X1_HVT U179 ( .A1(n605), .A3(n407), .A2(n362), .A4(n406), .S0(n248), 
        .S1(n354), .Y(n453) );
  MUX41X1_HVT U180 ( .A1(n364), .A3(n623), .A2(n619), .A4(n311), .S0(n327), 
        .S1(n351), .Y(n452) );
  MUX41X1_HVT U181 ( .A1(n452), .A3(n454), .A2(n453), .A4(n456), .S0(in[0]), 
        .S1(n325), .Y(n451) );
  OA21X1_HVT U184 ( .A1(n599), .A2(n231), .A3(n374), .Y(n448) );
  MUX41X1_HVT U189 ( .A1(n444), .A3(n618), .A2(n445), .A4(n393), .S0(n327), 
        .S1(n351), .Y(n443) );
  MUX41X1_HVT U193 ( .A1(n591), .A3(n598), .A2(n585), .A4(n441), .S0(n351), 
        .S1(n354), .Y(n440) );
  MUX41X1_HVT U195 ( .A1(n625), .A3(n398), .A2(n343), .A4(n596), .S0(n248), 
        .S1(n329), .Y(n438) );
  AO21X1_HVT U197 ( .A1(n314), .A2(n328), .A3(n395), .Y(n436) );
  OA21X1_HVT U201 ( .A1(n624), .A2(n219), .A3(n386), .Y(n432) );
  MUX41X1_HVT U203 ( .A1(n597), .A3(n264), .A2(n620), .A4(n601), .S0(n351), 
        .S1(n328), .Y(n430) );
  MUX41X1_HVT U205 ( .A1(n256), .A3(n271), .A2(n407), .A4(n381), .S0(n351), 
        .S1(n354), .Y(n428) );
  NAND2X0_HVT U208 ( .A1(n347), .A2(n338), .Y(n520) );
  NAND2X0_HVT U212 ( .A1(n345), .A2(n336), .Y(n577) );
  NAND2X0_HVT U214 ( .A1(n625), .A2(n350), .Y(n426) );
  NAND2X0_HVT U215 ( .A1(n520), .A2(n337), .Y(n425) );
  AO21X1_HVT U216 ( .A1(n349), .A2(n409), .A3(n231), .Y(n530) );
  NAND2X0_HVT U218 ( .A1(n409), .A2(n348), .Y(n479) );
  NAND2X0_HVT U220 ( .A1(n328), .A2(n426), .Y(n552) );
  MUX41X1_HVT U1 ( .A1(n473), .A3(n478), .A2(n471), .A4(n477), .S0(in[0]), 
        .S1(n19), .Y(n470) );
  IBUFFX16_HVT U2 ( .A(n325), .Y(n19) );
  DELLN1X2_HVT U3 ( .A(in[2]), .Y(n320) );
  MUX21X1_HVT U6 ( .A1(n474), .A2(n475), .S0(n324), .Y(n473) );
  INVX1_HVT U7 ( .A(n322), .Y(n246) );
  NBUFFX16_HVT U8 ( .A(n354), .Y(n328) );
  NAND2X0_HVT U9 ( .A1(n504), .A2(n23), .Y(n48) );
  NAND2X0_HVT U10 ( .A1(n503), .A2(n213), .Y(n50) );
  NAND2X0_HVT U11 ( .A1(n48), .A2(n50), .Y(n502) );
  INVX0_HVT U12 ( .A(n213), .Y(n23) );
  MUX21X1_HVT U14 ( .A1(n507), .A2(n508), .S0(n254), .Y(n504) );
  IBUFFX2_HVT U15 ( .A(n326), .Y(n213) );
  NAND2X1_HVT U16 ( .A1(n458), .A2(n210), .Y(n211) );
  NAND2X0_HVT U17 ( .A1(n470), .A2(in[6]), .Y(n212) );
  NAND2X0_HVT U18 ( .A1(n211), .A2(n212), .Y(out[5]) );
  IBUFFX2_HVT U19 ( .A(in[6]), .Y(n210) );
  INVX2_HVT U20 ( .A(in[7]), .Y(n356) );
  NBUFFX2_HVT U22 ( .A(in[7]), .Y(n255) );
  MUX21X2_HVT U23 ( .A1(n480), .A2(n481), .S0(n324), .Y(n478) );
  MUX41X1_HVT U25 ( .A1(n435), .A3(n439), .A2(n438), .A4(n440), .S0(in[0]), 
        .S1(n216), .Y(n434) );
  IBUFFX16_HVT U26 ( .A(n217), .Y(n216) );
  IBUFFX16_HVT U27 ( .A(n325), .Y(n217) );
  INVX2_HVT U28 ( .A(n355), .Y(n218) );
  INVX2_HVT U29 ( .A(n218), .Y(n219) );
  IBUFFX2_HVT U30 ( .A(n218), .Y(n231) );
  MUX21X2_HVT U31 ( .A1(n476), .A2(n342), .S0(n318), .Y(n475) );
  NAND2X1_HVT U32 ( .A1(n540), .A2(n232), .Y(n233) );
  NAND2X0_HVT U34 ( .A1(n541), .A2(n324), .Y(n234) );
  NAND2X0_HVT U36 ( .A1(n233), .A2(n234), .Y(n538) );
  IBUFFX2_HVT U37 ( .A(n324), .Y(n232) );
  NAND2X1_HVT U38 ( .A1(n524), .A2(n235), .Y(n236) );
  NAND2X0_HVT U39 ( .A1(n534), .A2(n244), .Y(n237) );
  NAND2X0_HVT U40 ( .A1(n236), .A2(n237), .Y(out[2]) );
  INVX1_HVT U41 ( .A(n244), .Y(n235) );
  MUX21X1_HVT U43 ( .A1(n342), .A2(n542), .S0(n318), .Y(n541) );
  IBUFFX2_HVT U44 ( .A(n303), .Y(n244) );
  IBUFFX4_HVT U45 ( .A(n356), .Y(n353) );
  INVX4_HVT U46 ( .A(n356), .Y(n354) );
  INVX0_HVT U47 ( .A(n354), .Y(n305) );
  XNOR2X2_HVT U48 ( .A1(n219), .A2(n278), .Y(n318) );
  NAND2X0_HVT U49 ( .A1(n380), .A2(n238), .Y(n239) );
  NAND2X0_HVT U50 ( .A1(n496), .A2(n274), .Y(n240) );
  NAND2X0_HVT U51 ( .A1(n239), .A2(n240), .Y(n495) );
  IBUFFX2_HVT U52 ( .A(n274), .Y(n238) );
  NAND2X0_HVT U54 ( .A1(n482), .A2(n241), .Y(n242) );
  NAND2X0_HVT U55 ( .A1(n490), .A2(n245), .Y(n243) );
  NAND2X2_HVT U60 ( .A1(n242), .A2(n243), .Y(out[4]) );
  INVX1_HVT U64 ( .A(n245), .Y(n241) );
  INVX1_HVT U65 ( .A(n419), .Y(n380) );
  INVX0_HVT U67 ( .A(n263), .Y(n274) );
  IBUFFX2_HVT U70 ( .A(n303), .Y(n245) );
  IBUFFX2_HVT U71 ( .A(in[7]), .Y(n355) );
  MUX41X1_HVT U72 ( .A1(n606), .A3(n626), .A2(n409), .A4(n404), .S0(n246), 
        .S1(n355), .Y(n494) );
  INVX1_HVT U76 ( .A(n286), .Y(n247) );
  INVX0_HVT U79 ( .A(n323), .Y(n263) );
  INVX1_HVT U81 ( .A(n262), .Y(n248) );
  INVX0_HVT U82 ( .A(n324), .Y(n262) );
  INVX1_HVT U87 ( .A(n329), .Y(n254) );
  MUX21X1_HVT U88 ( .A1(n595), .A2(n401), .S0(n327), .Y(n474) );
  INVX0_HVT U89 ( .A(n305), .Y(n267) );
  INVX0_HVT U90 ( .A(n349), .Y(n249) );
  INVX0_HVT U91 ( .A(n349), .Y(n250) );
  INVX0_HVT U92 ( .A(n349), .Y(n345) );
  IBUFFX16_HVT U94 ( .A(n349), .Y(n347) );
  MUX21X1_HVT U95 ( .A1(n341), .A2(n331), .S0(n249), .Y(n592) );
  INVX1_HVT U99 ( .A(n413), .Y(n251) );
  INVX0_HVT U100 ( .A(in[4]), .Y(n252) );
  INVX2_HVT U102 ( .A(in[4]), .Y(n413) );
  INVX0_HVT U104 ( .A(n266), .Y(n253) );
  INVX0_HVT U106 ( .A(n345), .Y(n266) );
  INVX2_HVT U107 ( .A(in[1]), .Y(n349) );
  INVX1_HVT U108 ( .A(n349), .Y(n346) );
  INVX0_HVT U111 ( .A(n413), .Y(n256) );
  INVX1_HVT U112 ( .A(n273), .Y(n606) );
  NAND2X1_HVT U113 ( .A1(n564), .A2(n257), .Y(n258) );
  NAND2X0_HVT U117 ( .A1(n589), .A2(n263), .Y(n259) );
  NAND2X0_HVT U118 ( .A1(n258), .A2(n259), .Y(n563) );
  INVX1_HVT U119 ( .A(n263), .Y(n257) );
  MUX21X1_HVT U120 ( .A1(n340), .A2(n344), .S0(n253), .Y(n273) );
  XOR2X1_HVT U121 ( .A1(n219), .A2(n606), .Y(n589) );
  AND2X1_HVT U122 ( .A1(n272), .A2(n331), .Y(n260) );
  IBUFFX4_HVT U124 ( .A(n260), .Y(n616) );
  MUX41X1_HVT U126 ( .A1(n548), .A3(n551), .A2(n546), .A4(n550), .S0(in[0]), 
        .S1(n261), .Y(n545) );
  IBUFFX16_HVT U127 ( .A(n325), .Y(n261) );
  MUX21X2_HVT U128 ( .A1(n612), .A2(n337), .S0(n329), .Y(n554) );
  INVX0_HVT U129 ( .A(n264), .Y(n593) );
  MUX21X2_HVT U130 ( .A1(n553), .A2(n554), .S0(n262), .Y(n551) );
  NBUFFX4_HVT U132 ( .A(n270), .Y(n342) );
  NBUFFX4_HVT U133 ( .A(n270), .Y(n341) );
  MUX21X1_HVT U134 ( .A1(n342), .A2(n265), .S0(n266), .Y(n264) );
  IBUFFX16_HVT U135 ( .A(n293), .Y(n265) );
  INVX0_HVT U137 ( .A(n340), .Y(n412) );
  MUX41X1_HVT U138 ( .A1(n292), .A3(n373), .A2(n396), .A4(n357), .S0(n267), 
        .S1(n268), .Y(n584) );
  IBUFFX16_HVT U139 ( .A(in[5]), .Y(n268) );
  INVX0_HVT U143 ( .A(n292), .Y(n613) );
  INVX0_HVT U145 ( .A(n630), .Y(n269) );
  INVX0_HVT U149 ( .A(n269), .Y(n270) );
  NBUFFX2_HVT U150 ( .A(n629), .Y(n271) );
  NBUFFX2_HVT U152 ( .A(n629), .Y(n272) );
  NAND2X0_HVT U155 ( .A1(n250), .A2(n341), .Y(n629) );
  INVX0_HVT U156 ( .A(n351), .Y(n286) );
  MUX21X1_HVT U157 ( .A1(n492), .A2(n628), .S0(n324), .Y(n491) );
  INVX0_HVT U160 ( .A(n335), .Y(n293) );
  INVX1_HVT U161 ( .A(n281), .Y(n278) );
  INVX0_HVT U164 ( .A(in[6]), .Y(n303) );
  INVX1_HVT U165 ( .A(in[5]), .Y(n287) );
  NBUFFX2_HVT U169 ( .A(n352), .Y(n325) );
  INVX1_HVT U171 ( .A(in[0]), .Y(n291) );
  INVX1_HVT U172 ( .A(n263), .Y(n294) );
  INVX0_HVT U173 ( .A(n323), .Y(n288) );
  XOR2X1_HVT U175 ( .A1(n277), .A2(n281), .Y(n587) );
  MUX41X1_HVT U176 ( .A1(n587), .A3(n560), .A2(n594), .A4(n315), .S0(n263), 
        .S1(n305), .Y(n446) );
  INVX1_HVT U182 ( .A(n277), .Y(n625) );
  NAND2X0_HVT U183 ( .A1(n576), .A2(n274), .Y(n275) );
  NAND2X0_HVT U185 ( .A1(n574), .A2(n262), .Y(n276) );
  NAND2X0_HVT U186 ( .A1(n275), .A2(n276), .Y(n573) );
  IBUFFX2_HVT U187 ( .A(n592), .Y(n388) );
  MUX21X2_HVT U188 ( .A1(n511), .A2(n514), .S0(n326), .Y(n510) );
  MUX41X1_HVT U190 ( .A1(n617), .A3(n358), .A2(n373), .A4(n588), .S0(n288), 
        .S1(n231), .Y(n550) );
  INVX1_HVT U191 ( .A(n423), .Y(n397) );
  XNOR2X1_HVT U192 ( .A1(n413), .A2(n334), .Y(n277) );
  MUX21X1_HVT U194 ( .A1(n311), .A2(n615), .S0(n305), .Y(n433) );
  MUX21X1_HVT U196 ( .A1(n331), .A2(n411), .S0(n249), .Y(n624) );
  NAND2X0_HVT U198 ( .A1(n427), .A2(n303), .Y(n297) );
  MUX21X1_HVT U199 ( .A1(n333), .A2(n330), .S0(n281), .Y(n529) );
  MUX41X1_HVT U200 ( .A1(n333), .A3(n457), .A2(n402), .A4(n618), .S0(n327), 
        .S1(n247), .Y(n456) );
  NAND2X0_HVT U202 ( .A1(n410), .A2(n278), .Y(n279) );
  NAND2X0_HVT U204 ( .A1(n331), .A2(n281), .Y(n280) );
  NAND2X0_HVT U206 ( .A1(n279), .A2(n280), .Y(n615) );
  IBUFFX2_HVT U207 ( .A(in[1]), .Y(n281) );
  INVX0_HVT U209 ( .A(n615), .Y(n371) );
  NAND2X0_HVT U210 ( .A1(n335), .A2(n278), .Y(n282) );
  NAND2X0_HVT U211 ( .A1(n330), .A2(n350), .Y(n283) );
  NAND2X0_HVT U213 ( .A1(n282), .A2(n283), .Y(n610) );
  MUX21X1_HVT U217 ( .A1(n610), .A2(n387), .S0(n328), .Y(n492) );
  NAND2X0_HVT U219 ( .A1(n580), .A2(n288), .Y(n284) );
  NAND2X0_HVT U221 ( .A1(n584), .A2(n294), .Y(n285) );
  NAND2X0_HVT U222 ( .A1(n284), .A2(n285), .Y(n579) );
  MUX41X1_HVT U223 ( .A1(n610), .A3(n383), .A2(n619), .A4(n578), .S0(n286), 
        .S1(n219), .Y(n429) );
  MUX41X1_HVT U224 ( .A1(n493), .A3(n495), .A2(n491), .A4(n494), .S0(in[0]), 
        .S1(n287), .Y(n490) );
  NAND2X0_HVT U225 ( .A1(n448), .A2(n288), .Y(n289) );
  NAND2X0_HVT U226 ( .A1(n449), .A2(n323), .Y(n290) );
  NAND2X0_HVT U227 ( .A1(n289), .A2(n290), .Y(n447) );
  MUX41X1_HVT U228 ( .A1(n447), .A3(n450), .A2(n443), .A4(n446), .S0(n325), 
        .S1(n291), .Y(n442) );
  MUX21X1_HVT U229 ( .A1(n293), .A2(n340), .S0(n349), .Y(n292) );
  NAND2X0_HVT U230 ( .A1(n436), .A2(n294), .Y(n295) );
  NAND2X0_HVT U231 ( .A1(n437), .A2(n263), .Y(n296) );
  NAND2X0_HVT U232 ( .A1(n296), .A2(n295), .Y(n435) );
  NAND2X0_HVT U233 ( .A1(n434), .A2(in[6]), .Y(n298) );
  NAND2X0_HVT U234 ( .A1(n298), .A2(n297), .Y(out[7]) );
  NAND2X0_HVT U235 ( .A1(n570), .A2(n263), .Y(n299) );
  NAND2X0_HVT U236 ( .A1(n572), .A2(n323), .Y(n300) );
  NAND2X0_HVT U237 ( .A1(n299), .A2(n300), .Y(n569) );
  NAND2X0_HVT U238 ( .A1(n432), .A2(n262), .Y(n301) );
  NAND2X0_HVT U239 ( .A1(n433), .A2(n323), .Y(n302) );
  NAND2X0_HVT U240 ( .A1(n301), .A2(n302), .Y(n431) );
  NBUFFX2_HVT U241 ( .A(n277), .Y(n331) );
  XNOR2X1_HVT U242 ( .A1(n349), .A2(n288), .Y(n310) );
  AO21X2_HVT U243 ( .A1(n324), .A2(n336), .A3(n625), .Y(n512) );
  MUX41X1_HVT U244 ( .A1(n544), .A3(n396), .A2(n591), .A4(n587), .S0(n262), 
        .S1(n231), .Y(n543) );
  XNOR2X1_HVT U245 ( .A1(n263), .A2(n305), .Y(n309) );
  INVX2_HVT U246 ( .A(n288), .Y(n351) );
  MUX21X2_HVT U247 ( .A1(n533), .A2(n316), .S0(n309), .Y(n532) );
  MUX41X1_HVT U248 ( .A1(n428), .A3(n429), .A2(n430), .A4(n431), .S0(n325), 
        .S1(in[0]), .Y(n427) );
  NBUFFX2_HVT U249 ( .A(n413), .Y(n332) );
  AND3X2_HVT U250 ( .A1(n294), .A2(n350), .A3(n251), .Y(n500) );
  NBUFFX2_HVT U251 ( .A(n252), .Y(n333) );
  NBUFFX2_HVT U252 ( .A(in[2]), .Y(n321) );
  MUX21X1_HVT U253 ( .A1(n337), .A2(n339), .S0(n249), .Y(n304) );
  MUX41X1_HVT U254 ( .A1(n466), .A3(n587), .A2(n379), .A4(n611), .S0(n231), 
        .S1(n262), .Y(n465) );
  MUX41X1_HVT U255 ( .A1(n467), .A3(n462), .A2(n465), .A4(n459), .S0(n291), 
        .S1(n287), .Y(n458) );
  MUX41X1_HVT U256 ( .A1(n376), .A3(n388), .A2(n627), .A4(n387), .S0(n231), 
        .S1(n262), .Y(n450) );
  MUX41X1_HVT U257 ( .A1(n516), .A3(n502), .A2(n510), .A4(n497), .S0(n303), 
        .S1(n291), .Y(out[3]) );
  MUX41X1_HVT U258 ( .A1(n532), .A3(n527), .A2(n528), .A4(n525), .S0(n291), 
        .S1(n287), .Y(n524) );
  MUX41X1_HVT U259 ( .A1(n622), .A3(n404), .A2(n606), .A4(n592), .S0(n305), 
        .S1(n263), .Y(n439) );
  NAND2X0_HVT U260 ( .A1(n342), .A2(n306), .Y(n307) );
  NAND2X0_HVT U261 ( .A1(n518), .A2(n310), .Y(n308) );
  NAND2X0_HVT U262 ( .A1(n307), .A2(n308), .Y(n517) );
  INVX0_HVT U263 ( .A(n310), .Y(n306) );
  INVX0_HVT U264 ( .A(n349), .Y(n348) );
  INVX0_HVT U265 ( .A(n334), .Y(n410) );
  MUX21X2_HVT U266 ( .A1(n442), .A2(n451), .S0(in[6]), .Y(out[6]) );
  MUX21X2_HVT U267 ( .A1(n545), .A2(n555), .S0(in[6]), .Y(out[1]) );
  INVX1_HVT U268 ( .A(n627), .Y(n408) );
  AND2X1_HVT U269 ( .A1(n331), .A2(n577), .Y(n311) );
  MUX21X1_HVT U270 ( .A1(n313), .A2(n371), .S0(n321), .Y(n499) );
  NBUFFX2_HVT U271 ( .A(n277), .Y(n330) );
  NBUFFX2_HVT U272 ( .A(n627), .Y(n338) );
  NBUFFX2_HVT U273 ( .A(n627), .Y(n339) );
  MUX21X1_HVT U274 ( .A1(n408), .A2(n411), .S0(n326), .Y(n581) );
  MUX21X1_HVT U275 ( .A1(n602), .A2(n521), .S0(n321), .Y(n519) );
  MUX21X1_HVT U276 ( .A1(n367), .A2(n409), .S0(n326), .Y(n566) );
  AND2X1_HVT U277 ( .A1(n341), .A2(n560), .Y(n312) );
  MUX21X1_HVT U278 ( .A1(n339), .A2(n625), .S0(n347), .Y(n596) );
  MUX21X1_HVT U279 ( .A1(n408), .A2(n412), .S0(n249), .Y(n457) );
  MUX21X1_HVT U280 ( .A1(n411), .A2(n408), .S0(n345), .Y(n595) );
  MUX21X1_HVT U281 ( .A1(n331), .A2(n408), .S0(n278), .Y(n537) );
  NAND2X0_HVT U282 ( .A1(n332), .A2(n410), .Y(n627) );
  MUX21X1_HVT U283 ( .A1(n625), .A2(n409), .S0(n346), .Y(n417) );
  NBUFFX2_HVT U284 ( .A(n630), .Y(n340) );
  MUX21X1_HVT U285 ( .A1(n625), .A2(n412), .S0(n249), .Y(n608) );
  MUX21X1_HVT U286 ( .A1(n411), .A2(n331), .S0(n347), .Y(n469) );
  MUX21X1_HVT U287 ( .A1(n338), .A2(n337), .S0(n348), .Y(n544) );
  MUX21X1_HVT U288 ( .A1(n625), .A2(n332), .S0(n348), .Y(n557) );
  INVX1_HVT U289 ( .A(n622), .Y(n409) );
  INVX1_HVT U290 ( .A(n343), .Y(n411) );
  MUX21X1_HVT U291 ( .A1(n411), .A2(n293), .S0(n249), .Y(n599) );
  MUX21X1_HVT U292 ( .A1(n333), .A2(n408), .S0(n348), .Y(n604) );
  MUX21X1_HVT U293 ( .A1(n403), .A2(n337), .S0(n328), .Y(n496) );
  MUX21X1_HVT U294 ( .A1(n512), .A2(n513), .S0(n328), .Y(n511) );
  MUX21X1_HVT U295 ( .A1(n360), .A2(n383), .S0(n321), .Y(n513) );
  MUX21X1_HVT U296 ( .A1(n410), .A2(n332), .S0(n345), .Y(n441) );
  XOR2X1_HVT U297 ( .A1(n340), .A2(n250), .Y(n585) );
  MUX21X1_HVT U298 ( .A1(n408), .A2(n333), .S0(n250), .Y(n418) );
  MUX21X1_HVT U299 ( .A1(n293), .A2(n625), .S0(n250), .Y(n420) );
  MUX21X1_HVT U300 ( .A1(n338), .A2(n293), .S0(n250), .Y(n620) );
  MUX21X1_HVT U301 ( .A1(n359), .A2(n509), .S0(n322), .Y(n508) );
  MUX21X1_HVT U302 ( .A1(n332), .A2(n293), .S0(n250), .Y(n509) );
  MUX21X1_HVT U303 ( .A1(n293), .A2(n344), .S0(n348), .Y(n444) );
  MUX21X1_HVT U304 ( .A1(n343), .A2(n341), .S0(n347), .Y(n445) );
  MUX21X1_HVT U305 ( .A1(n343), .A2(n336), .S0(n345), .Y(n602) );
  MUX21X1_HVT U306 ( .A1(n342), .A2(n336), .S0(n345), .Y(n617) );
  MUX21X1_HVT U307 ( .A1(n627), .A2(n344), .S0(n278), .Y(n539) );
  MUX21X1_HVT U308 ( .A1(n293), .A2(n411), .S0(n345), .Y(n621) );
  MUX21X1_HVT U309 ( .A1(n381), .A2(n617), .S0(n324), .Y(n533) );
  XOR2X1_HVT U310 ( .A1(n278), .A2(n409), .Y(n588) );
  XNOR2X1_HVT U311 ( .A1(n339), .A2(n346), .Y(n313) );
  XNOR2X1_HVT U312 ( .A1(n343), .A2(n278), .Y(n314) );
  AND2X1_HVT U313 ( .A1(n278), .A2(n412), .Y(n315) );
  MUX21X1_HVT U314 ( .A1(n336), .A2(n410), .S0(n249), .Y(n422) );
  AND2X1_HVT U315 ( .A1(n344), .A2(n520), .Y(n316) );
  MUX21X1_HVT U316 ( .A1(n340), .A2(n333), .S0(n249), .Y(n424) );
  MUX21X1_HVT U317 ( .A1(n340), .A2(n338), .S0(n346), .Y(n416) );
  MUX21X1_HVT U318 ( .A1(n337), .A2(n333), .S0(n348), .Y(n562) );
  MUX21X1_HVT U319 ( .A1(n337), .A2(n344), .S0(n324), .Y(n506) );
  XOR2X1_HVT U320 ( .A1(n332), .A2(n250), .Y(n607) );
  NBUFFX2_HVT U321 ( .A(n354), .Y(n327) );
  NBUFFX2_HVT U322 ( .A(n354), .Y(n329) );
  NBUFFX2_HVT U323 ( .A(n352), .Y(n326) );
  NBUFFX2_HVT U324 ( .A(in[2]), .Y(n323) );
  NBUFFX2_HVT U325 ( .A(in[2]), .Y(n322) );
  NBUFFX2_HVT U326 ( .A(in[2]), .Y(n324) );
  MUX21X1_HVT U327 ( .A1(n531), .A2(n380), .S0(n320), .Y(n528) );
  MUX21X1_HVT U328 ( .A1(n547), .A2(n335), .S0(n328), .Y(n449) );
  XOR2X1_HVT U329 ( .A1(n347), .A2(n334), .Y(n586) );
  MUX21X1_HVT U330 ( .A1(n336), .A2(n330), .S0(n278), .Y(n526) );
  NAND2X0_HVT U331 ( .A1(n334), .A2(n333), .Y(n630) );
  AND2X1_HVT U332 ( .A1(n330), .A2(n350), .Y(n317) );
  NBUFFX2_HVT U333 ( .A(n631), .Y(n343) );
  MUX21X1_HVT U334 ( .A1(n335), .A2(n408), .S0(n278), .Y(n594) );
  MUX21X1_HVT U335 ( .A1(n411), .A2(n398), .S0(n329), .Y(n564) );
  MUX21X1_HVT U336 ( .A1(n461), .A2(n460), .S0(n274), .Y(n459) );
  MUX21X1_HVT U337 ( .A1(n337), .A2(n398), .S0(n329), .Y(n461) );
  MUX21X1_HVT U338 ( .A1(n486), .A2(n485), .S0(n274), .Y(n484) );
  MUX21X1_HVT U339 ( .A1(n604), .A2(n363), .S0(n329), .Y(n486) );
  MUX21X1_HVT U340 ( .A1(n400), .A2(n409), .S0(n328), .Y(n481) );
  MUX21X1_HVT U341 ( .A1(n384), .A2(n272), .S0(n322), .Y(n523) );
  MUX21X1_HVT U342 ( .A1(n614), .A2(n382), .S0(n322), .Y(n498) );
  MUX21X1_HVT U343 ( .A1(n271), .A2(n349), .S0(n323), .Y(n505) );
  MUX21X1_HVT U344 ( .A1(n409), .A2(n412), .S0(n250), .Y(n466) );
  NBUFFX2_HVT U345 ( .A(n622), .Y(n336) );
  MUX21X1_HVT U346 ( .A1(n582), .A2(n583), .S0(n327), .Y(n580) );
  MUX21X1_HVT U347 ( .A1(n335), .A2(n598), .S0(n326), .Y(n583) );
  XOR2X1_HVT U348 ( .A1(n348), .A2(n325), .Y(n590) );
  MUX21X1_HVT U349 ( .A1(n389), .A2(n406), .S0(n328), .Y(n437) );
  MUX21X1_HVT U350 ( .A1(n335), .A2(n409), .S0(n348), .Y(n421) );
  NBUFFX2_HVT U351 ( .A(n631), .Y(n344) );
  MUX21X1_HVT U352 ( .A1(n603), .A2(n425), .S0(n327), .Y(n419) );
  MUX21X1_HVT U353 ( .A1(n339), .A2(n335), .S0(n278), .Y(n623) );
  MUX21X1_HVT U354 ( .A1(n377), .A2(n603), .S0(n322), .Y(n501) );
  MUX21X1_HVT U355 ( .A1(n369), .A2(n350), .S0(n326), .Y(n568) );
  MUX21X1_HVT U356 ( .A1(n335), .A2(n332), .S0(n329), .Y(n542) );
  NBUFFX2_HVT U357 ( .A(n622), .Y(n337) );
  AND2X1_HVT U358 ( .A1(n410), .A2(n350), .Y(n319) );
  NBUFFX2_HVT U359 ( .A(in[5]), .Y(n352) );
  MUX21X1_HVT U360 ( .A1(n408), .A2(n251), .S0(n346), .Y(n601) );
  NAND2X0_HVT U361 ( .A1(in[4]), .A2(n410), .Y(n622) );
  NAND2X0_HVT U362 ( .A1(n334), .A2(in[4]), .Y(n631) );
  MUX21X1_HVT U363 ( .A1(n251), .A2(n411), .S0(n348), .Y(n597) );
  MUX21X1_HVT U364 ( .A1(n251), .A2(n625), .S0(n346), .Y(n423) );
  MUX21X1_HVT U365 ( .A1(n251), .A2(n409), .S0(n278), .Y(n614) );
  MUX21X1_HVT U366 ( .A1(n251), .A2(n342), .S0(n347), .Y(n612) );
  MUX21X1_HVT U367 ( .A1(n251), .A2(n336), .S0(n347), .Y(n415) );
  MUX21X1_HVT U368 ( .A1(n251), .A2(n344), .S0(n346), .Y(n414) );
  MUX21X1_HVT U369 ( .A1(n344), .A2(n251), .S0(n250), .Y(n605) );
  MUX21X1_HVT U370 ( .A1(n335), .A2(n251), .S0(n321), .Y(n518) );
  MUX21X1_HVT U371 ( .A1(n293), .A2(n251), .S0(n345), .Y(n603) );
  NBUFFX2_HVT U372 ( .A(in[3]), .Y(n334) );
  INVX0_HVT U373 ( .A(in[1]), .Y(n350) );
  NBUFFX2_HVT U374 ( .A(in[3]), .Y(n335) );
  INVX0_HVT U375 ( .A(n611), .Y(n357) );
  INVX0_HVT U376 ( .A(n609), .Y(n358) );
  INVX0_HVT U377 ( .A(n600), .Y(n359) );
  INVX0_HVT U378 ( .A(n598), .Y(n360) );
  INVX0_HVT U379 ( .A(n463), .Y(n361) );
  INVX0_HVT U380 ( .A(n426), .Y(n362) );
  INVX0_HVT U381 ( .A(n271), .Y(n363) );
  INVX0_HVT U382 ( .A(n628), .Y(n364) );
  INVX0_HVT U383 ( .A(n626), .Y(n365) );
  INVX0_HVT U384 ( .A(n624), .Y(n366) );
  INVX0_HVT U385 ( .A(n623), .Y(n367) );
  INVX0_HVT U386 ( .A(n621), .Y(n368) );
  INVX0_HVT U387 ( .A(n620), .Y(n369) );
  INVX0_HVT U388 ( .A(n617), .Y(n370) );
  INVX0_HVT U389 ( .A(n614), .Y(n372) );
  INVX0_HVT U390 ( .A(n612), .Y(n373) );
  INVX0_HVT U391 ( .A(n610), .Y(n374) );
  INVX0_HVT U392 ( .A(n608), .Y(n375) );
  INVX0_HVT U393 ( .A(n607), .Y(n376) );
  INVX0_HVT U394 ( .A(n605), .Y(n377) );
  INVX0_HVT U395 ( .A(n604), .Y(n378) );
  INVX0_HVT U396 ( .A(n603), .Y(n379) );
  INVX0_HVT U397 ( .A(n602), .Y(n381) );
  INVX0_HVT U398 ( .A(n601), .Y(n382) );
  INVX0_HVT U399 ( .A(n599), .Y(n383) );
  INVX0_HVT U400 ( .A(n597), .Y(n384) );
  INVX0_HVT U401 ( .A(n596), .Y(n385) );
  INVX0_HVT U402 ( .A(n595), .Y(n386) );
  INVX0_HVT U403 ( .A(n594), .Y(n387) );
  INVX0_HVT U404 ( .A(n591), .Y(n389) );
  INVX0_HVT U405 ( .A(n560), .Y(n390) );
  INVX0_HVT U406 ( .A(n619), .Y(n391) );
  INVX0_HVT U407 ( .A(n520), .Y(n392) );
  INVX0_HVT U408 ( .A(n425), .Y(n393) );
  INVX0_HVT U409 ( .A(n577), .Y(n394) );
  INVX0_HVT U410 ( .A(n479), .Y(n395) );
  INVX0_HVT U411 ( .A(n424), .Y(n396) );
  INVX0_HVT U412 ( .A(n422), .Y(n398) );
  INVX0_HVT U413 ( .A(n421), .Y(n399) );
  INVX0_HVT U414 ( .A(n420), .Y(n400) );
  INVX0_HVT U415 ( .A(n539), .Y(n401) );
  INVX0_HVT U416 ( .A(n529), .Y(n402) );
  INVX0_HVT U417 ( .A(n418), .Y(n403) );
  INVX0_HVT U418 ( .A(n417), .Y(n404) );
  INVX0_HVT U419 ( .A(n416), .Y(n405) );
  INVX0_HVT U420 ( .A(n415), .Y(n406) );
  INVX0_HVT U421 ( .A(n414), .Y(n407) );
endmodule

