
module round ( in, round_num, keyin, keyout, out );
  input [127:0] in;
  input [3:0] round_num;
  input [127:0] keyin;
  output [127:0] keyout;
  output [127:0] out;
  wire   n130, n131, n132, \_0_net_[127] , \_0_net_[126] , \_0_net_[125] ,
         \_0_net_[124] , \_0_net_[123] , \_0_net_[122] , \_0_net_[121] ,
         \_0_net_[120] , \_0_net_[119] , \_0_net_[118] , \_0_net_[117] ,
         \_0_net_[116] , \_0_net_[115] , \_0_net_[114] , \_0_net_[113] ,
         \_0_net_[112] , \_0_net_[111] , \_0_net_[110] , \_0_net_[109] ,
         \_0_net_[108] , \_0_net_[107] , \_0_net_[106] , \_0_net_[105] ,
         \_0_net_[104] , \_0_net_[103] , \_0_net_[102] , \_0_net_[101] ,
         \_0_net_[100] , \_0_net_[99] , \_0_net_[98] , \_0_net_[97] ,
         \_0_net_[96] , \_0_net_[95] , \_0_net_[94] , \_0_net_[93] ,
         \_0_net_[92] , \_0_net_[91] , \_0_net_[90] , \_0_net_[89] ,
         \_0_net_[88] , \_0_net_[87] , \_0_net_[86] , \_0_net_[85] ,
         \_0_net_[84] , \_0_net_[83] , \_0_net_[82] , \_0_net_[81] ,
         \_0_net_[80] , \_0_net_[79] , \_0_net_[78] , \_0_net_[77] ,
         \_0_net_[76] , \_0_net_[75] , \_0_net_[74] , \_0_net_[73] ,
         \_0_net_[72] , \_0_net_[71] , \_0_net_[70] , \_0_net_[69] ,
         \_0_net_[68] , \_0_net_[67] , \_0_net_[66] , \_0_net_[65] ,
         \_0_net_[64] , \_0_net_[63] , \_0_net_[62] , \_0_net_[61] ,
         \_0_net_[60] , \_0_net_[59] , \_0_net_[58] , \_0_net_[57] ,
         \_0_net_[56] , \_0_net_[55] , \_0_net_[54] , \_0_net_[53] ,
         \_0_net_[52] , \_0_net_[51] , \_0_net_[50] , \_0_net_[49] ,
         \_0_net_[48] , \_0_net_[47] , \_0_net_[46] , \_0_net_[45] ,
         \_0_net_[44] , \_0_net_[43] , \_0_net_[42] , \_0_net_[41] ,
         \_0_net_[40] , \_0_net_[39] , \_0_net_[38] , \_0_net_[37] ,
         \_0_net_[36] , \_0_net_[35] , \_0_net_[34] , \_0_net_[33] ,
         \_0_net_[32] , \_0_net_[31] , \_0_net_[30] , \_0_net_[29] ,
         \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , \_0_net_[25] ,
         \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , \_0_net_[21] ,
         \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , \_0_net_[17] ,
         \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , \_0_net_[13] ,
         \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , \_0_net_[9] ,
         \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] ,
         \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_0_net_[0] , n2, n3, n1,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129;
  wire   [127:0] sb_out;
  wire   [127:0] sr_out;
  wire   [127:0] mc_out;

  AO22X1_HVT U2 ( .A1(mc_out[9]), .A2(n116), .A3(n90), .A4(n119), .Y(
        \_0_net_[9] ) );
  AO22X1_HVT U3 ( .A1(mc_out[99]), .A2(n116), .A3(sr_out[99]), .A4(n119), .Y(
        \_0_net_[99] ) );
  AO22X1_HVT U4 ( .A1(mc_out[98]), .A2(n116), .A3(n15), .A4(n119), .Y(
        \_0_net_[98] ) );
  AO22X1_HVT U5 ( .A1(mc_out[97]), .A2(n116), .A3(sr_out[97]), .A4(n119), .Y(
        \_0_net_[97] ) );
  AO22X1_HVT U6 ( .A1(mc_out[96]), .A2(n115), .A3(n6), .A4(n119), .Y(
        \_0_net_[96] ) );
  AO22X1_HVT U7 ( .A1(mc_out[95]), .A2(n115), .A3(n91), .A4(n119), .Y(
        \_0_net_[95] ) );
  AO22X1_HVT U8 ( .A1(n115), .A2(mc_out[94]), .A3(sr_out[94]), .A4(n119), .Y(
        \_0_net_[94] ) );
  AO22X1_HVT U9 ( .A1(n115), .A2(mc_out[93]), .A3(sr_out[93]), .A4(n119), .Y(
        \_0_net_[93] ) );
  AO22X1_HVT U11 ( .A1(mc_out[91]), .A2(n115), .A3(sr_out[91]), .A4(n119), .Y(
        \_0_net_[91] ) );
  AO22X1_HVT U12 ( .A1(mc_out[90]), .A2(n115), .A3(n22), .A4(n119), .Y(
        \_0_net_[90] ) );
  AO22X1_HVT U13 ( .A1(mc_out[8]), .A2(n115), .A3(sr_out[8]), .A4(n119), .Y(
        \_0_net_[8] ) );
  AO22X1_HVT U15 ( .A1(mc_out[88]), .A2(n115), .A3(sr_out[88]), .A4(n120), .Y(
        \_0_net_[88] ) );
  AO22X1_HVT U16 ( .A1(n115), .A2(mc_out[87]), .A3(sr_out[87]), .A4(n120), .Y(
        \_0_net_[87] ) );
  AO22X1_HVT U17 ( .A1(mc_out[86]), .A2(n115), .A3(n56), .A4(n120), .Y(
        \_0_net_[86] ) );
  AO22X1_HVT U18 ( .A1(mc_out[85]), .A2(n115), .A3(n60), .A4(n120), .Y(
        \_0_net_[85] ) );
  AO22X1_HVT U19 ( .A1(mc_out[84]), .A2(n115), .A3(sr_out[84]), .A4(n120), .Y(
        \_0_net_[84] ) );
  AO22X1_HVT U20 ( .A1(mc_out[83]), .A2(n115), .A3(n31), .A4(n120), .Y(
        \_0_net_[83] ) );
  AO22X1_HVT U21 ( .A1(mc_out[82]), .A2(n114), .A3(n13), .A4(n120), .Y(
        \_0_net_[82] ) );
  AO22X1_HVT U22 ( .A1(mc_out[81]), .A2(n114), .A3(n43), .A4(n120), .Y(
        \_0_net_[81] ) );
  AO22X1_HVT U23 ( .A1(mc_out[80]), .A2(n114), .A3(sr_out[80]), .A4(n120), .Y(
        \_0_net_[80] ) );
  AO22X1_HVT U24 ( .A1(mc_out[7]), .A2(n114), .A3(n99), .A4(n120), .Y(
        \_0_net_[7] ) );
  AO22X1_HVT U25 ( .A1(mc_out[79]), .A2(n114), .A3(sr_out[79]), .A4(n120), .Y(
        \_0_net_[79] ) );
  AO22X1_HVT U26 ( .A1(mc_out[78]), .A2(n114), .A3(sr_out[78]), .A4(n121), .Y(
        \_0_net_[78] ) );
  AO22X1_HVT U27 ( .A1(n114), .A2(mc_out[77]), .A3(sr_out[77]), .A4(n121), .Y(
        \_0_net_[77] ) );
  AO22X1_HVT U30 ( .A1(mc_out[74]), .A2(n114), .A3(sr_out[74]), .A4(n121), .Y(
        \_0_net_[74] ) );
  AO22X1_HVT U31 ( .A1(mc_out[73]), .A2(n114), .A3(sr_out[73]), .A4(n121), .Y(
        \_0_net_[73] ) );
  AO22X1_HVT U32 ( .A1(mc_out[72]), .A2(n114), .A3(sr_out[72]), .A4(n121), .Y(
        \_0_net_[72] ) );
  AO22X1_HVT U33 ( .A1(mc_out[71]), .A2(n114), .A3(sr_out[71]), .A4(n121), .Y(
        \_0_net_[71] ) );
  AO22X1_HVT U34 ( .A1(mc_out[70]), .A2(n114), .A3(sr_out[70]), .A4(n121), .Y(
        \_0_net_[70] ) );
  AO22X1_HVT U35 ( .A1(mc_out[6]), .A2(n114), .A3(n46), .A4(n121), .Y(
        \_0_net_[6] ) );
  AO22X1_HVT U36 ( .A1(mc_out[69]), .A2(n113), .A3(n74), .A4(n121), .Y(
        \_0_net_[69] ) );
  AO22X1_HVT U37 ( .A1(mc_out[68]), .A2(n113), .A3(sr_out[68]), .A4(n121), .Y(
        \_0_net_[68] ) );
  AO22X1_HVT U38 ( .A1(mc_out[67]), .A2(n113), .A3(n82), .A4(n122), .Y(
        \_0_net_[67] ) );
  AO22X1_HVT U39 ( .A1(mc_out[66]), .A2(n113), .A3(sr_out[66]), .A4(n122), .Y(
        \_0_net_[66] ) );
  AO22X1_HVT U40 ( .A1(mc_out[65]), .A2(n113), .A3(sr_out[65]), .A4(n122), .Y(
        \_0_net_[65] ) );
  AO22X1_HVT U41 ( .A1(n113), .A2(mc_out[64]), .A3(sr_out[64]), .A4(n122), .Y(
        \_0_net_[64] ) );
  AO22X1_HVT U43 ( .A1(mc_out[62]), .A2(n113), .A3(n70), .A4(n122), .Y(
        \_0_net_[62] ) );
  AO22X1_HVT U44 ( .A1(mc_out[61]), .A2(n113), .A3(sr_out[61]), .A4(n122), .Y(
        \_0_net_[61] ) );
  AO22X1_HVT U46 ( .A1(mc_out[5]), .A2(n113), .A3(n68), .A4(n122), .Y(
        \_0_net_[5] ) );
  AO22X1_HVT U47 ( .A1(mc_out[59]), .A2(n113), .A3(n23), .A4(n122), .Y(
        \_0_net_[59] ) );
  AO22X1_HVT U48 ( .A1(mc_out[58]), .A2(n113), .A3(sr_out[58]), .A4(n122), .Y(
        \_0_net_[58] ) );
  AO22X1_HVT U49 ( .A1(mc_out[57]), .A2(n113), .A3(sr_out[57]), .A4(n122), .Y(
        \_0_net_[57] ) );
  AO22X1_HVT U50 ( .A1(mc_out[56]), .A2(n113), .A3(sr_out[56]), .A4(n123), .Y(
        \_0_net_[56] ) );
  AO22X1_HVT U52 ( .A1(mc_out[54]), .A2(n112), .A3(n81), .A4(n123), .Y(
        \_0_net_[54] ) );
  AO22X1_HVT U56 ( .A1(mc_out[50]), .A2(n112), .A3(n123), .A4(sr_out[50]), .Y(
        \_0_net_[50] ) );
  AO22X1_HVT U57 ( .A1(mc_out[4]), .A2(n112), .A3(sr_out[4]), .A4(n123), .Y(
        \_0_net_[4] ) );
  AO22X1_HVT U58 ( .A1(mc_out[49]), .A2(n112), .A3(n123), .A4(sr_out[49]), .Y(
        \_0_net_[49] ) );
  AO22X1_HVT U59 ( .A1(mc_out[48]), .A2(n112), .A3(n75), .A4(n123), .Y(
        \_0_net_[48] ) );
  AO22X1_HVT U60 ( .A1(mc_out[47]), .A2(n112), .A3(n69), .A4(n123), .Y(
        \_0_net_[47] ) );
  AO22X1_HVT U61 ( .A1(mc_out[46]), .A2(n112), .A3(sr_out[46]), .A4(n123), .Y(
        \_0_net_[46] ) );
  AO22X1_HVT U62 ( .A1(mc_out[45]), .A2(n112), .A3(sr_out[45]), .A4(n124), .Y(
        \_0_net_[45] ) );
  AO22X1_HVT U63 ( .A1(mc_out[44]), .A2(n112), .A3(n78), .A4(n124), .Y(
        \_0_net_[44] ) );
  AO22X1_HVT U65 ( .A1(mc_out[42]), .A2(n112), .A3(n16), .A4(n124), .Y(
        \_0_net_[42] ) );
  AO22X1_HVT U67 ( .A1(mc_out[40]), .A2(n111), .A3(sr_out[40]), .A4(n124), .Y(
        \_0_net_[40] ) );
  AO22X1_HVT U68 ( .A1(mc_out[3]), .A2(n111), .A3(sr_out[3]), .A4(n124), .Y(
        \_0_net_[3] ) );
  AO22X1_HVT U70 ( .A1(mc_out[38]), .A2(n111), .A3(sr_out[38]), .A4(n124), .Y(
        \_0_net_[38] ) );
  AO22X1_HVT U71 ( .A1(mc_out[37]), .A2(n111), .A3(n12), .A4(n124), .Y(
        \_0_net_[37] ) );
  AO22X1_HVT U72 ( .A1(mc_out[36]), .A2(n111), .A3(sr_out[36]), .A4(n124), .Y(
        \_0_net_[36] ) );
  AO22X1_HVT U75 ( .A1(mc_out[33]), .A2(n111), .A3(sr_out[33]), .A4(n125), .Y(
        \_0_net_[33] ) );
  AO22X1_HVT U76 ( .A1(mc_out[32]), .A2(n111), .A3(sr_out[32]), .A4(n125), .Y(
        \_0_net_[32] ) );
  AO22X1_HVT U77 ( .A1(mc_out[31]), .A2(n111), .A3(n84), .A4(n125), .Y(
        \_0_net_[31] ) );
  AO22X1_HVT U78 ( .A1(mc_out[30]), .A2(n111), .A3(sr_out[30]), .A4(n125), .Y(
        \_0_net_[30] ) );
  AO22X1_HVT U79 ( .A1(mc_out[2]), .A2(n111), .A3(sr_out[2]), .A4(n125), .Y(
        \_0_net_[2] ) );
  AO22X1_HVT U80 ( .A1(mc_out[29]), .A2(n111), .A3(n24), .A4(n125), .Y(
        \_0_net_[29] ) );
  AO22X1_HVT U82 ( .A1(mc_out[27]), .A2(n110), .A3(n72), .A4(n125), .Y(
        \_0_net_[27] ) );
  AO22X1_HVT U83 ( .A1(mc_out[26]), .A2(n110), .A3(sr_out[26]), .A4(n125), .Y(
        \_0_net_[26] ) );
  AO22X1_HVT U84 ( .A1(mc_out[25]), .A2(n110), .A3(sr_out[25]), .A4(n125), .Y(
        \_0_net_[25] ) );
  AO22X1_HVT U85 ( .A1(mc_out[24]), .A2(n110), .A3(n96), .A4(n125), .Y(
        \_0_net_[24] ) );
  AO22X1_HVT U86 ( .A1(mc_out[23]), .A2(n110), .A3(n55), .A4(n126), .Y(
        \_0_net_[23] ) );
  AO22X1_HVT U87 ( .A1(mc_out[22]), .A2(n110), .A3(n7), .A4(n126), .Y(
        \_0_net_[22] ) );
  AO22X1_HVT U88 ( .A1(mc_out[21]), .A2(n110), .A3(sr_out[21]), .A4(n126), .Y(
        \_0_net_[21] ) );
  AO22X1_HVT U90 ( .A1(mc_out[1]), .A2(n110), .A3(sr_out[1]), .A4(n126), .Y(
        \_0_net_[1] ) );
  AO22X1_HVT U92 ( .A1(mc_out[18]), .A2(n110), .A3(sr_out[18]), .A4(n126), .Y(
        \_0_net_[18] ) );
  AO22X1_HVT U93 ( .A1(mc_out[17]), .A2(n110), .A3(sr_out[17]), .A4(n126), .Y(
        \_0_net_[17] ) );
  AO22X1_HVT U94 ( .A1(mc_out[16]), .A2(n110), .A3(sr_out[16]), .A4(n126), .Y(
        \_0_net_[16] ) );
  AO22X1_HVT U95 ( .A1(mc_out[15]), .A2(n110), .A3(n101), .A4(n126), .Y(
        \_0_net_[15] ) );
  AO22X1_HVT U96 ( .A1(mc_out[14]), .A2(n109), .A3(sr_out[14]), .A4(n126), .Y(
        \_0_net_[14] ) );
  AO22X1_HVT U97 ( .A1(mc_out[13]), .A2(n109), .A3(sr_out[13]), .A4(n126), .Y(
        \_0_net_[13] ) );
  AO22X1_HVT U98 ( .A1(mc_out[12]), .A2(n109), .A3(n42), .A4(n127), .Y(
        \_0_net_[12] ) );
  AO22X1_HVT U99 ( .A1(mc_out[127]), .A2(n109), .A3(n100), .A4(n127), .Y(
        \_0_net_[127] ) );
  AO22X1_HVT U100 ( .A1(mc_out[126]), .A2(n109), .A3(n9), .A4(n127), .Y(
        \_0_net_[126] ) );
  AO22X1_HVT U101 ( .A1(mc_out[125]), .A2(n109), .A3(sr_out[125]), .A4(n127), 
        .Y(\_0_net_[125] ) );
  AO22X1_HVT U102 ( .A1(mc_out[124]), .A2(n109), .A3(sr_out[124]), .A4(n127), 
        .Y(\_0_net_[124] ) );
  AO22X1_HVT U103 ( .A1(mc_out[123]), .A2(n109), .A3(sr_out[123]), .A4(n127), 
        .Y(\_0_net_[123] ) );
  AO22X1_HVT U104 ( .A1(mc_out[122]), .A2(n109), .A3(sr_out[122]), .A4(n127), 
        .Y(\_0_net_[122] ) );
  AO22X1_HVT U105 ( .A1(mc_out[121]), .A2(n109), .A3(sr_out[121]), .A4(n127), 
        .Y(\_0_net_[121] ) );
  AO22X1_HVT U106 ( .A1(mc_out[120]), .A2(n109), .A3(sr_out[120]), .A4(n127), 
        .Y(\_0_net_[120] ) );
  AO22X1_HVT U108 ( .A1(mc_out[119]), .A2(n109), .A3(sr_out[119]), .A4(n127), 
        .Y(\_0_net_[119] ) );
  AO22X1_HVT U109 ( .A1(mc_out[118]), .A2(n109), .A3(sr_out[118]), .A4(n127), 
        .Y(\_0_net_[118] ) );
  AO22X1_HVT U110 ( .A1(n109), .A2(mc_out[117]), .A3(sr_out[117]), .A4(n128), 
        .Y(\_0_net_[117] ) );
  AO22X1_HVT U111 ( .A1(mc_out[116]), .A2(n108), .A3(n83), .A4(n128), .Y(
        \_0_net_[116] ) );
  AO22X1_HVT U112 ( .A1(mc_out[115]), .A2(n108), .A3(sr_out[115]), .A4(n128), 
        .Y(\_0_net_[115] ) );
  AO22X1_HVT U113 ( .A1(mc_out[114]), .A2(n108), .A3(sr_out[114]), .A4(n128), 
        .Y(\_0_net_[114] ) );
  AO22X1_HVT U114 ( .A1(mc_out[113]), .A2(n108), .A3(n87), .A4(n128), .Y(
        \_0_net_[113] ) );
  AO22X1_HVT U115 ( .A1(mc_out[112]), .A2(n108), .A3(sr_out[112]), .A4(n128), 
        .Y(\_0_net_[112] ) );
  AO22X1_HVT U116 ( .A1(mc_out[111]), .A2(n108), .A3(n21), .A4(n128), .Y(
        \_0_net_[111] ) );
  AO22X1_HVT U117 ( .A1(mc_out[110]), .A2(n108), .A3(sr_out[110]), .A4(n128), 
        .Y(\_0_net_[110] ) );
  AO22X1_HVT U118 ( .A1(mc_out[10]), .A2(n108), .A3(sr_out[10]), .A4(n128), 
        .Y(\_0_net_[10] ) );
  AO22X1_HVT U119 ( .A1(mc_out[109]), .A2(n108), .A3(sr_out[109]), .A4(n128), 
        .Y(\_0_net_[109] ) );
  AO22X1_HVT U120 ( .A1(mc_out[108]), .A2(n108), .A3(sr_out[108]), .A4(n128), 
        .Y(\_0_net_[108] ) );
  AO22X1_HVT U121 ( .A1(mc_out[107]), .A2(n108), .A3(sr_out[107]), .A4(n128), 
        .Y(\_0_net_[107] ) );
  AO22X1_HVT U122 ( .A1(mc_out[106]), .A2(n108), .A3(n54), .A4(n129), .Y(
        \_0_net_[106] ) );
  AO22X1_HVT U123 ( .A1(mc_out[105]), .A2(n108), .A3(n5), .A4(n129), .Y(
        \_0_net_[105] ) );
  AO22X1_HVT U124 ( .A1(mc_out[104]), .A2(n108), .A3(sr_out[104]), .A4(n129), 
        .Y(\_0_net_[104] ) );
  AO22X1_HVT U125 ( .A1(mc_out[103]), .A2(n108), .A3(sr_out[103]), .A4(n129), 
        .Y(\_0_net_[103] ) );
  AO22X1_HVT U126 ( .A1(mc_out[102]), .A2(n107), .A3(sr_out[102]), .A4(n129), 
        .Y(\_0_net_[102] ) );
  AO22X1_HVT U127 ( .A1(mc_out[101]), .A2(n107), .A3(n67), .A4(n129), .Y(
        \_0_net_[101] ) );
  AO22X1_HVT U128 ( .A1(mc_out[100]), .A2(n107), .A3(sr_out[100]), .A4(n129), 
        .Y(\_0_net_[100] ) );
  AO22X1_HVT U129 ( .A1(mc_out[0]), .A2(n106), .A3(sr_out[0]), .A4(n129), .Y(
        \_0_net_[0] ) );
  OR3X1_HVT U130 ( .A1(round_num[2]), .A2(round_num[0]), .A3(n3), .Y(n2) );
  NAND2X0_HVT U131 ( .A1(round_num[3]), .A2(round_num[1]), .Y(n3) );
  keygen_0 x ( .round_num(round_num), .keyin({keyin[127:8], n103, keyin[6:0]}), 
        .keyout({keyout[127:95], n130, keyout[93:91], n131, keyout[89:26], 
        n132, keyout[24:0]}) );
  subbytes sb ( .in(in), .out(sb_out) );
  shift_rows sr ( .in(sb_out), .out(sr_out) );
  Mix_Column mc ( .in({sr_out[127:116], n86, sr_out[114:88], n102, 
        sr_out[86:85], n49, sr_out[83:0]}), .out(mc_out) );
  add_round_keys_1 adk ( .state({\_0_net_[127] , \_0_net_[126] , 
        \_0_net_[125] , \_0_net_[124] , \_0_net_[123] , \_0_net_[122] , 
        \_0_net_[121] , \_0_net_[120] , \_0_net_[119] , \_0_net_[118] , 
        \_0_net_[117] , \_0_net_[116] , \_0_net_[115] , \_0_net_[114] , 
        \_0_net_[113] , \_0_net_[112] , \_0_net_[111] , \_0_net_[110] , 
        \_0_net_[109] , \_0_net_[108] , \_0_net_[107] , \_0_net_[106] , 
        \_0_net_[105] , \_0_net_[104] , \_0_net_[103] , \_0_net_[102] , 
        \_0_net_[101] , \_0_net_[100] , \_0_net_[99] , \_0_net_[98] , 
        \_0_net_[97] , \_0_net_[96] , \_0_net_[95] , \_0_net_[94] , 
        \_0_net_[93] , \_0_net_[92] , \_0_net_[91] , \_0_net_[90] , 
        \_0_net_[89] , \_0_net_[88] , \_0_net_[87] , \_0_net_[86] , 
        \_0_net_[85] , \_0_net_[84] , \_0_net_[83] , \_0_net_[82] , 
        \_0_net_[81] , \_0_net_[80] , \_0_net_[79] , \_0_net_[78] , 
        \_0_net_[77] , \_0_net_[76] , \_0_net_[75] , \_0_net_[74] , 
        \_0_net_[73] , \_0_net_[72] , \_0_net_[71] , \_0_net_[70] , 
        \_0_net_[69] , \_0_net_[68] , \_0_net_[67] , \_0_net_[66] , 
        \_0_net_[65] , \_0_net_[64] , \_0_net_[63] , \_0_net_[62] , 
        \_0_net_[61] , \_0_net_[60] , \_0_net_[59] , \_0_net_[58] , 
        \_0_net_[57] , \_0_net_[56] , \_0_net_[55] , \_0_net_[54] , 
        \_0_net_[53] , \_0_net_[52] , \_0_net_[51] , \_0_net_[50] , 
        \_0_net_[49] , \_0_net_[48] , \_0_net_[47] , \_0_net_[46] , 
        \_0_net_[45] , \_0_net_[44] , \_0_net_[43] , \_0_net_[42] , 
        \_0_net_[41] , \_0_net_[40] , \_0_net_[39] , \_0_net_[38] , 
        \_0_net_[37] , \_0_net_[36] , \_0_net_[35] , \_0_net_[34] , 
        \_0_net_[33] , \_0_net_[32] , \_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_0_net_[0] }), 
        .subkey({keyout[127:95], n130, keyout[93:91], n131, keyout[89:26], 
        n132, keyout[24:0]}), .out(out) );
  IBUFFX2_HVT U1 ( .A(n132), .Y(n1) );
  INVX0_HVT U10 ( .A(n1), .Y(keyout[25]) );
  DELLN2X2_HVT U14 ( .A(sr_out[105]), .Y(n5) );
  DELLN2X2_HVT U28 ( .A(sr_out[81]), .Y(n43) );
  NBUFFX2_HVT U29 ( .A(sr_out[106]), .Y(n52) );
  DELLN2X2_HVT U42 ( .A(sr_out[96]), .Y(n6) );
  DELLN2X2_HVT U45 ( .A(sr_out[22]), .Y(n7) );
  DELLN2X2_HVT U51 ( .A(sr_out[39]), .Y(n95) );
  DELLN1X2_HVT U53 ( .A(sr_out[35]), .Y(n8) );
  DELLN2X2_HVT U54 ( .A(sr_out[83]), .Y(n31) );
  DELLN2X2_HVT U55 ( .A(sr_out[126]), .Y(n9) );
  NBUFFX2_HVT U64 ( .A(sr_out[9]), .Y(n90) );
  NAND2X0_HVT U66 ( .A1(mc_out[76]), .A2(n114), .Y(n10) );
  NAND2X1_HVT U69 ( .A1(n71), .A2(n121), .Y(n11) );
  NAND2X0_HVT U73 ( .A1(n10), .A2(n11), .Y(\_0_net_[76] ) );
  IBUFFX16_HVT U74 ( .A(n117), .Y(n114) );
  DELLN1X2_HVT U81 ( .A(sr_out[76]), .Y(n71) );
  INVX1_HVT U89 ( .A(n107), .Y(n121) );
  DELLN2X2_HVT U91 ( .A(sr_out[37]), .Y(n12) );
  DELLN2X2_HVT U107 ( .A(sr_out[86]), .Y(n56) );
  DELLN1X2_HVT U132 ( .A(sr_out[82]), .Y(n13) );
  DELLN2X2_HVT U133 ( .A(sr_out[20]), .Y(n14) );
  NAND2X0_HVT U134 ( .A1(n126), .A2(n14), .Y(n45) );
  NBUFFX2_HVT U135 ( .A(sr_out[12]), .Y(n42) );
  NBUFFX2_HVT U136 ( .A(sr_out[44]), .Y(n78) );
  DELLN1X2_HVT U137 ( .A(sr_out[98]), .Y(n15) );
  DELLN2X2_HVT U138 ( .A(sr_out[42]), .Y(n16) );
  NAND2X0_HVT U139 ( .A1(sr_out[34]), .A2(n125), .Y(n48) );
  NAND2X0_HVT U140 ( .A1(mc_out[92]), .A2(n115), .Y(n17) );
  NAND2X1_HVT U141 ( .A1(sr_out[92]), .A2(n119), .Y(n18) );
  NAND2X0_HVT U142 ( .A1(n17), .A2(n18), .Y(\_0_net_[92] ) );
  INVX2_HVT U143 ( .A(n117), .Y(n115) );
  NAND2X0_HVT U144 ( .A1(mc_out[28]), .A2(n110), .Y(n19) );
  NAND2X0_HVT U145 ( .A1(sr_out[28]), .A2(n125), .Y(n20) );
  NAND2X0_HVT U146 ( .A1(n19), .A2(n20), .Y(\_0_net_[28] ) );
  INVX1_HVT U147 ( .A(n118), .Y(n110) );
  DELLN2X2_HVT U148 ( .A(sr_out[111]), .Y(n21) );
  NBUFFX2_HVT U149 ( .A(sr_out[90]), .Y(n22) );
  DELLN2X2_HVT U150 ( .A(sr_out[55]), .Y(n61) );
  DELLN2X2_HVT U151 ( .A(sr_out[59]), .Y(n23) );
  DELLN1X2_HVT U152 ( .A(sr_out[101]), .Y(n41) );
  DELLN2X2_HVT U153 ( .A(sr_out[29]), .Y(n24) );
  NAND2X0_HVT U154 ( .A1(mc_out[55]), .A2(n112), .Y(n25) );
  NAND2X1_HVT U155 ( .A1(n61), .A2(n123), .Y(n26) );
  NAND2X0_HVT U156 ( .A1(n25), .A2(n26), .Y(\_0_net_[55] ) );
  DELLN2X2_HVT U157 ( .A(sr_out[63]), .Y(n50) );
  NAND2X0_HVT U158 ( .A1(mc_out[39]), .A2(n111), .Y(n27) );
  NAND2X0_HVT U159 ( .A1(n95), .A2(n124), .Y(n28) );
  NAND2X0_HVT U160 ( .A1(n27), .A2(n28), .Y(\_0_net_[39] ) );
  NAND2X0_HVT U161 ( .A1(mc_out[19]), .A2(n110), .Y(n29) );
  NAND2X0_HVT U162 ( .A1(sr_out[19]), .A2(n126), .Y(n30) );
  NAND2X0_HVT U163 ( .A1(n29), .A2(n30), .Y(\_0_net_[19] ) );
  NAND2X0_HVT U164 ( .A1(sr_out[75]), .A2(n121), .Y(n77) );
  NAND2X0_HVT U165 ( .A1(mc_out[89]), .A2(n115), .Y(n32) );
  NAND2X0_HVT U166 ( .A1(sr_out[89]), .A2(n120), .Y(n33) );
  NAND2X0_HVT U167 ( .A1(n32), .A2(n33), .Y(\_0_net_[89] ) );
  NAND2X0_HVT U168 ( .A1(mc_out[63]), .A2(n113), .Y(n34) );
  NAND2X0_HVT U169 ( .A1(n50), .A2(n122), .Y(n35) );
  NAND2X0_HVT U170 ( .A1(n34), .A2(n35), .Y(\_0_net_[63] ) );
  NAND2X0_HVT U171 ( .A1(mc_out[53]), .A2(n112), .Y(n36) );
  NAND2X0_HVT U172 ( .A1(sr_out[53]), .A2(n123), .Y(n37) );
  NAND2X0_HVT U173 ( .A1(n36), .A2(n37), .Y(\_0_net_[53] ) );
  NAND2X0_HVT U174 ( .A1(mc_out[11]), .A2(n109), .Y(n38) );
  NAND2X0_HVT U175 ( .A1(sr_out[11]), .A2(n127), .Y(n39) );
  NAND2X0_HVT U176 ( .A1(n38), .A2(n39), .Y(\_0_net_[11] ) );
  DELLN2X2_HVT U177 ( .A(sr_out[41]), .Y(n40) );
  NBUFFX2_HVT U178 ( .A(sr_out[84]), .Y(n49) );
  IBUFFX2_HVT U179 ( .A(n41), .Y(n66) );
  NAND2X0_HVT U180 ( .A1(mc_out[20]), .A2(n110), .Y(n44) );
  NAND2X0_HVT U181 ( .A1(n44), .A2(n45), .Y(\_0_net_[20] ) );
  INVX0_HVT U182 ( .A(n106), .Y(n126) );
  DELLN2X2_HVT U183 ( .A(sr_out[6]), .Y(n46) );
  NAND2X0_HVT U184 ( .A1(mc_out[34]), .A2(n111), .Y(n47) );
  NAND2X0_HVT U185 ( .A1(n47), .A2(n48), .Y(\_0_net_[34] ) );
  INVX0_HVT U186 ( .A(n106), .Y(n125) );
  DELLN2X2_HVT U187 ( .A(sr_out[15]), .Y(n101) );
  DELLN1X2_HVT U188 ( .A(sr_out[85]), .Y(n51) );
  DELLN1X2_HVT U189 ( .A(sr_out[62]), .Y(n70) );
  IBUFFX2_HVT U190 ( .A(n52), .Y(n53) );
  INVX1_HVT U191 ( .A(n53), .Y(n54) );
  DELLN2X2_HVT U192 ( .A(sr_out[31]), .Y(n84) );
  DELLN2X2_HVT U193 ( .A(sr_out[23]), .Y(n55) );
  DELLN1X2_HVT U194 ( .A(sr_out[5]), .Y(n68) );
  NBUFFX2_HVT U195 ( .A(sr_out[113]), .Y(n87) );
  NBUFFX2_HVT U196 ( .A(sr_out[60]), .Y(n94) );
  IBUFFX2_HVT U197 ( .A(n130), .Y(n57) );
  INVX0_HVT U198 ( .A(n57), .Y(keyout[94]) );
  IBUFFX2_HVT U199 ( .A(n51), .Y(n59) );
  INVX1_HVT U200 ( .A(n59), .Y(n60) );
  NAND2X0_HVT U201 ( .A1(mc_out[41]), .A2(n111), .Y(n62) );
  NAND2X0_HVT U202 ( .A1(n40), .A2(n124), .Y(n63) );
  NAND2X0_HVT U203 ( .A1(n62), .A2(n63), .Y(\_0_net_[41] ) );
  INVX1_HVT U204 ( .A(n117), .Y(n111) );
  NAND2X0_HVT U205 ( .A1(mc_out[51]), .A2(n112), .Y(n64) );
  NAND2X0_HVT U206 ( .A1(n123), .A2(sr_out[51]), .Y(n65) );
  NAND2X0_HVT U207 ( .A1(n64), .A2(n65), .Y(\_0_net_[51] ) );
  INVX1_HVT U208 ( .A(n107), .Y(n123) );
  INVX1_HVT U209 ( .A(n66), .Y(n67) );
  DELLN2X2_HVT U210 ( .A(sr_out[47]), .Y(n69) );
  DELLN2X2_HVT U211 ( .A(sr_out[27]), .Y(n72) );
  IBUFFX2_HVT U212 ( .A(sr_out[69]), .Y(n73) );
  INVX1_HVT U213 ( .A(n73), .Y(n74) );
  DELLN2X2_HVT U214 ( .A(sr_out[48]), .Y(n75) );
  NAND2X0_HVT U215 ( .A1(mc_out[75]), .A2(n114), .Y(n76) );
  NAND2X0_HVT U216 ( .A1(n76), .A2(n77), .Y(\_0_net_[75] ) );
  NAND2X0_HVT U217 ( .A1(n8), .A2(n124), .Y(n89) );
  NAND2X0_HVT U218 ( .A1(mc_out[52]), .A2(n112), .Y(n79) );
  NAND2X0_HVT U219 ( .A1(sr_out[52]), .A2(n123), .Y(n80) );
  NAND2X0_HVT U220 ( .A1(n79), .A2(n80), .Y(\_0_net_[52] ) );
  INVX1_HVT U221 ( .A(n117), .Y(n112) );
  DELLN2X2_HVT U222 ( .A(sr_out[54]), .Y(n81) );
  DELLN2X2_HVT U223 ( .A(sr_out[67]), .Y(n82) );
  DELLN2X2_HVT U224 ( .A(sr_out[116]), .Y(n83) );
  INVX1_HVT U225 ( .A(sr_out[115]), .Y(n85) );
  INVX2_HVT U226 ( .A(n85), .Y(n86) );
  NBUFFX2_HVT U227 ( .A(sr_out[87]), .Y(n102) );
  NAND2X0_HVT U228 ( .A1(n111), .A2(mc_out[35]), .Y(n88) );
  NAND2X0_HVT U229 ( .A1(n88), .A2(n89), .Y(\_0_net_[35] ) );
  DELLN2X2_HVT U230 ( .A(sr_out[95]), .Y(n91) );
  NAND2X0_HVT U231 ( .A1(mc_out[60]), .A2(n113), .Y(n92) );
  NAND2X0_HVT U232 ( .A1(n94), .A2(n122), .Y(n93) );
  NAND2X0_HVT U233 ( .A1(n92), .A2(n93), .Y(\_0_net_[60] ) );
  DELLN2X2_HVT U234 ( .A(sr_out[24]), .Y(n96) );
  NAND2X0_HVT U235 ( .A1(mc_out[43]), .A2(n112), .Y(n97) );
  NAND2X0_HVT U236 ( .A1(sr_out[43]), .A2(n124), .Y(n98) );
  NAND2X0_HVT U237 ( .A1(n97), .A2(n98), .Y(\_0_net_[43] ) );
  DELLN2X2_HVT U238 ( .A(sr_out[7]), .Y(n99) );
  DELLN2X2_HVT U239 ( .A(sr_out[127]), .Y(n100) );
  NBUFFX16_HVT U240 ( .A(keyin[7]), .Y(n103) );
  IBUFFX2_HVT U241 ( .A(n131), .Y(n104) );
  INVX1_HVT U242 ( .A(n104), .Y(keyout[90]) );
  INVX0_HVT U243 ( .A(n107), .Y(n119) );
  INVX0_HVT U244 ( .A(n118), .Y(n107) );
  INVX0_HVT U245 ( .A(n118), .Y(n106) );
  INVX0_HVT U246 ( .A(n117), .Y(n116) );
  INVX1_HVT U247 ( .A(n2), .Y(n117) );
  INVX1_HVT U248 ( .A(n107), .Y(n122) );
  INVX1_HVT U249 ( .A(n107), .Y(n120) );
  INVX1_HVT U250 ( .A(n106), .Y(n124) );
  INVX1_HVT U251 ( .A(n106), .Y(n127) );
  INVX1_HVT U252 ( .A(n106), .Y(n128) );
  INVX1_HVT U253 ( .A(n106), .Y(n129) );
  INVX1_HVT U254 ( .A(n117), .Y(n113) );
  INVX1_HVT U255 ( .A(n118), .Y(n109) );
  INVX1_HVT U256 ( .A(n118), .Y(n108) );
  INVX0_HVT U257 ( .A(n2), .Y(n118) );
endmodule

