
module add_round_keys_1 ( state, subkey, out );
  input [127:0] state;
  input [127:0] subkey;
  output [127:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310;

  XOR2X2_HVT U3 ( .A1(subkey[98]), .A2(state[98]), .Y(out[98]) );
  XOR2X2_HVT U12 ( .A1(subkey[8]), .A2(state[8]), .Y(out[8]) );
  XOR2X2_HVT U14 ( .A1(subkey[88]), .A2(state[88]), .Y(out[88]) );
  XOR2X2_HVT U15 ( .A1(subkey[87]), .A2(state[87]), .Y(out[87]) );
  XOR2X2_HVT U20 ( .A1(subkey[82]), .A2(state[82]), .Y(out[82]) );
  XOR2X2_HVT U22 ( .A1(subkey[80]), .A2(state[80]), .Y(out[80]) );
  XOR2X2_HVT U23 ( .A1(subkey[7]), .A2(state[7]), .Y(out[7]) );
  XOR2X2_HVT U29 ( .A1(subkey[74]), .A2(state[74]), .Y(out[74]) );
  XOR2X2_HVT U31 ( .A1(subkey[72]), .A2(state[72]), .Y(out[72]) );
  XOR2X2_HVT U33 ( .A1(subkey[70]), .A2(state[70]), .Y(out[70]) );
  XOR2X2_HVT U34 ( .A1(state[6]), .A2(subkey[6]), .Y(out[6]) );
  XOR2X2_HVT U35 ( .A1(state[69]), .A2(subkey[69]), .Y(out[69]) );
  XOR2X2_HVT U40 ( .A1(subkey[64]), .A2(state[64]), .Y(out[64]) );
  XOR2X2_HVT U50 ( .A1(subkey[55]), .A2(state[55]), .Y(out[55]) );
  XOR2X2_HVT U51 ( .A1(subkey[54]), .A2(state[54]), .Y(out[54]) );
  XOR2X2_HVT U57 ( .A1(state[49]), .A2(subkey[49]), .Y(out[49]) );
  XOR2X2_HVT U58 ( .A1(subkey[48]), .A2(state[48]), .Y(out[48]) );
  XOR2X2_HVT U59 ( .A1(state[47]), .A2(subkey[47]), .Y(out[47]) );
  XOR2X2_HVT U62 ( .A1(state[44]), .A2(subkey[44]), .Y(out[44]) );
  XOR2X2_HVT U64 ( .A1(state[42]), .A2(subkey[42]), .Y(out[42]) );
  XOR2X2_HVT U66 ( .A1(state[40]), .A2(subkey[40]), .Y(out[40]) );
  XOR2X2_HVT U70 ( .A1(state[37]), .A2(subkey[37]), .Y(out[37]) );
  XOR2X2_HVT U77 ( .A1(state[30]), .A2(subkey[30]), .Y(out[30]) );
  XOR2X2_HVT U78 ( .A1(subkey[2]), .A2(state[2]), .Y(out[2]) );
  XOR2X2_HVT U79 ( .A1(subkey[29]), .A2(state[29]), .Y(out[29]) );
  XOR2X2_HVT U82 ( .A1(subkey[26]), .A2(state[26]), .Y(out[26]) );
  XOR2X2_HVT U87 ( .A1(subkey[21]), .A2(state[21]), .Y(out[21]) );
  XOR2X2_HVT U92 ( .A1(state[17]), .A2(subkey[17]), .Y(out[17]) );
  XOR2X2_HVT U93 ( .A1(subkey[16]), .A2(state[16]), .Y(out[16]) );
  XOR2X2_HVT U95 ( .A1(subkey[14]), .A2(state[14]), .Y(out[14]) );
  XOR2X2_HVT U96 ( .A1(subkey[13]), .A2(state[13]), .Y(out[13]) );
  XOR2X2_HVT U103 ( .A1(subkey[122]), .A2(state[122]), .Y(out[122]) );
  XOR2X2_HVT U107 ( .A1(subkey[119]), .A2(state[119]), .Y(out[119]) );
  XOR2X2_HVT U114 ( .A1(subkey[112]), .A2(state[112]), .Y(out[112]) );
  XOR2X2_HVT U117 ( .A1(subkey[10]), .A2(state[10]), .Y(out[10]) );
  XOR2X2_HVT U123 ( .A1(subkey[104]), .A2(state[104]), .Y(out[104]) );
  XOR2X2_HVT U126 ( .A1(state[101]), .A2(subkey[101]), .Y(out[101]) );
  XOR2X2_HVT U128 ( .A1(subkey[0]), .A2(state[0]), .Y(out[0]) );
  XOR2X1_HVT U1 ( .A1(state[120]), .A2(subkey[120]), .Y(out[120]) );
  NAND2X0_HVT U2 ( .A1(state[76]), .A2(n6), .Y(n3) );
  NAND2X0_HVT U4 ( .A1(n1), .A2(n2), .Y(n4) );
  NAND2X0_HVT U5 ( .A1(n3), .A2(n4), .Y(out[76]) );
  INVX0_HVT U6 ( .A(state[76]), .Y(n1) );
  INVX16_HVT U7 ( .A(n6), .Y(n2) );
  OR2X1_HVT U8 ( .A1(n5), .A2(state[68]), .Y(n273) );
  IBUFFX16_HVT U9 ( .A(subkey[68]), .Y(n5) );
  IBUFFX16_HVT U10 ( .A(subkey[76]), .Y(n6) );
  INVX1_HVT U11 ( .A(state[4]), .Y(n195) );
  NAND2X0_HVT U13 ( .A1(state[28]), .A2(n206), .Y(n9) );
  NAND2X0_HVT U16 ( .A1(n7), .A2(n8), .Y(n10) );
  NAND2X0_HVT U17 ( .A1(n10), .A2(n9), .Y(out[28]) );
  INVX0_HVT U18 ( .A(state[28]), .Y(n7) );
  INVX0_HVT U19 ( .A(n206), .Y(n8) );
  IBUFFX2_HVT U21 ( .A(subkey[28]), .Y(n206) );
  INVX0_HVT U24 ( .A(subkey[103]), .Y(n37) );
  INVX0_HVT U25 ( .A(subkey[52]), .Y(n20) );
  XOR2X2_HVT U26 ( .A1(state[15]), .A2(subkey[15]), .Y(out[15]) );
  XOR2X2_HVT U27 ( .A1(subkey[127]), .A2(state[127]), .Y(out[127]) );
  NAND2X0_HVT U28 ( .A1(state[107]), .A2(n89), .Y(n13) );
  NAND2X0_HVT U30 ( .A1(n11), .A2(n12), .Y(n14) );
  NAND2X0_HVT U32 ( .A1(n13), .A2(n14), .Y(out[107]) );
  INVX0_HVT U36 ( .A(state[107]), .Y(n11) );
  INVX0_HVT U37 ( .A(n89), .Y(n12) );
  IBUFFX2_HVT U38 ( .A(subkey[107]), .Y(n89) );
  NAND2X0_HVT U39 ( .A1(state[105]), .A2(n19), .Y(n17) );
  NAND2X0_HVT U41 ( .A1(n15), .A2(n16), .Y(n18) );
  NAND2X0_HVT U42 ( .A1(n17), .A2(n18), .Y(out[105]) );
  INVX0_HVT U43 ( .A(state[105]), .Y(n15) );
  INVX16_HVT U44 ( .A(n19), .Y(n16) );
  IBUFFX16_HVT U45 ( .A(subkey[105]), .Y(n19) );
  OR2X1_HVT U46 ( .A1(n20), .A2(state[52]), .Y(n242) );
  INVX0_HVT U47 ( .A(subkey[116]), .Y(n151) );
  INVX0_HVT U48 ( .A(subkey[121]), .Y(n81) );
  INVX1_HVT U49 ( .A(subkey[100]), .Y(n122) );
  INVX0_HVT U52 ( .A(subkey[90]), .Y(n85) );
  INVX0_HVT U53 ( .A(subkey[85]), .Y(n21) );
  INVX0_HVT U54 ( .A(subkey[43]), .Y(n285) );
  INVX0_HVT U55 ( .A(subkey[39]), .Y(n245) );
  INVX0_HVT U56 ( .A(subkey[38]), .Y(n29) );
  INVX1_HVT U60 ( .A(subkey[20]), .Y(n228) );
  INVX1_HVT U61 ( .A(subkey[18]), .Y(n25) );
  INVX1_HVT U63 ( .A(subkey[1]), .Y(n131) );
  INVX0_HVT U65 ( .A(subkey[114]), .Y(n45) );
  INVX0_HVT U67 ( .A(subkey[96]), .Y(n146) );
  INVX1_HVT U68 ( .A(subkey[23]), .Y(n250) );
  INVX0_HVT U69 ( .A(subkey[35]), .Y(n244) );
  OR2X1_HVT U71 ( .A1(n267), .A2(state[75]), .Y(n180) );
  NAND2X0_HVT U72 ( .A1(subkey[85]), .A2(n22), .Y(n23) );
  NAND2X0_HVT U73 ( .A1(n21), .A2(state[85]), .Y(n24) );
  NAND2X0_HVT U74 ( .A1(n23), .A2(n24), .Y(out[85]) );
  INVX0_HVT U75 ( .A(state[85]), .Y(n22) );
  NAND2X0_HVT U76 ( .A1(subkey[18]), .A2(n26), .Y(n27) );
  NAND2X0_HVT U80 ( .A1(n25), .A2(state[18]), .Y(n28) );
  NAND2X0_HVT U81 ( .A1(n27), .A2(n28), .Y(out[18]) );
  INVX0_HVT U83 ( .A(state[18]), .Y(n26) );
  NAND2X0_HVT U84 ( .A1(subkey[38]), .A2(n30), .Y(n31) );
  NAND2X0_HVT U85 ( .A1(n29), .A2(state[38]), .Y(n32) );
  NAND2X0_HVT U86 ( .A1(n31), .A2(n32), .Y(out[38]) );
  INVX0_HVT U88 ( .A(state[38]), .Y(n30) );
  XOR2X2_HVT U89 ( .A1(subkey[118]), .A2(state[118]), .Y(out[118]) );
  INVX1_HVT U90 ( .A(subkey[75]), .Y(n267) );
  NAND2X0_HVT U91 ( .A1(subkey[126]), .A2(n34), .Y(n35) );
  NAND2X0_HVT U94 ( .A1(n33), .A2(state[126]), .Y(n36) );
  NAND2X0_HVT U97 ( .A1(n35), .A2(n36), .Y(out[126]) );
  IBUFFX2_HVT U98 ( .A(subkey[126]), .Y(n33) );
  INVX0_HVT U99 ( .A(state[126]), .Y(n34) );
  NAND2X0_HVT U100 ( .A1(subkey[103]), .A2(n38), .Y(n39) );
  NAND2X0_HVT U101 ( .A1(n37), .A2(state[103]), .Y(n40) );
  NAND2X0_HVT U102 ( .A1(n39), .A2(n40), .Y(out[103]) );
  INVX0_HVT U104 ( .A(state[103]), .Y(n38) );
  NAND2X0_HVT U105 ( .A1(subkey[106]), .A2(n42), .Y(n43) );
  NAND2X0_HVT U106 ( .A1(state[106]), .A2(n41), .Y(n44) );
  NAND2X0_HVT U108 ( .A1(n43), .A2(n44), .Y(out[106]) );
  IBUFFX2_HVT U109 ( .A(subkey[106]), .Y(n41) );
  INVX0_HVT U110 ( .A(state[106]), .Y(n42) );
  XNOR2X2_HVT U111 ( .A1(state[114]), .A2(n45), .Y(out[114]) );
  NAND2X0_HVT U112 ( .A1(subkey[111]), .A2(n47), .Y(n48) );
  NAND2X0_HVT U113 ( .A1(n46), .A2(state[111]), .Y(n49) );
  NAND2X0_HVT U115 ( .A1(n48), .A2(n49), .Y(out[111]) );
  IBUFFX2_HVT U116 ( .A(subkey[111]), .Y(n46) );
  INVX0_HVT U118 ( .A(state[111]), .Y(n47) );
  NAND2X0_HVT U119 ( .A1(subkey[93]), .A2(n51), .Y(n52) );
  NAND2X0_HVT U120 ( .A1(n50), .A2(state[93]), .Y(n53) );
  NAND2X0_HVT U121 ( .A1(n52), .A2(n53), .Y(out[93]) );
  INVX0_HVT U122 ( .A(subkey[93]), .Y(n50) );
  INVX0_HVT U124 ( .A(state[93]), .Y(n51) );
  NAND2X0_HVT U125 ( .A1(state[33]), .A2(n55), .Y(n56) );
  NAND2X0_HVT U127 ( .A1(n54), .A2(subkey[33]), .Y(n57) );
  NAND2X0_HVT U129 ( .A1(n56), .A2(n57), .Y(out[33]) );
  INVX0_HVT U130 ( .A(state[33]), .Y(n54) );
  INVX0_HVT U131 ( .A(subkey[33]), .Y(n55) );
  NAND2X0_HVT U132 ( .A1(subkey[102]), .A2(n59), .Y(n60) );
  NAND2X0_HVT U133 ( .A1(n58), .A2(state[102]), .Y(n61) );
  NAND2X0_HVT U134 ( .A1(n60), .A2(n61), .Y(out[102]) );
  IBUFFX2_HVT U135 ( .A(subkey[102]), .Y(n58) );
  INVX0_HVT U136 ( .A(state[102]), .Y(n59) );
  NAND2X0_HVT U137 ( .A1(subkey[9]), .A2(n63), .Y(n64) );
  NAND2X0_HVT U138 ( .A1(n62), .A2(state[9]), .Y(n65) );
  NAND2X0_HVT U139 ( .A1(n64), .A2(n65), .Y(out[9]) );
  INVX0_HVT U140 ( .A(subkey[9]), .Y(n62) );
  INVX0_HVT U141 ( .A(state[9]), .Y(n63) );
  INVX1_HVT U142 ( .A(subkey[51]), .Y(n277) );
  NAND2X0_HVT U143 ( .A1(n250), .A2(state[23]), .Y(n67) );
  NAND2X0_HVT U144 ( .A1(subkey[23]), .A2(n66), .Y(n68) );
  NAND2X0_HVT U145 ( .A1(n67), .A2(n68), .Y(out[23]) );
  INVX0_HVT U146 ( .A(state[23]), .Y(n66) );
  NAND2X0_HVT U147 ( .A1(subkey[117]), .A2(n70), .Y(n71) );
  NAND2X0_HVT U148 ( .A1(n69), .A2(state[117]), .Y(n72) );
  NAND2X0_HVT U149 ( .A1(n71), .A2(n72), .Y(out[117]) );
  IBUFFX2_HVT U150 ( .A(subkey[117]), .Y(n69) );
  INVX0_HVT U151 ( .A(state[117]), .Y(n70) );
  NAND2X0_HVT U152 ( .A1(state[50]), .A2(n74), .Y(n75) );
  NAND2X0_HVT U153 ( .A1(n73), .A2(subkey[50]), .Y(n76) );
  NAND2X0_HVT U154 ( .A1(n75), .A2(n76), .Y(out[50]) );
  INVX0_HVT U155 ( .A(state[50]), .Y(n73) );
  INVX0_HVT U156 ( .A(subkey[50]), .Y(n74) );
  NAND2X0_HVT U157 ( .A1(state[25]), .A2(n78), .Y(n79) );
  NAND2X0_HVT U158 ( .A1(n77), .A2(subkey[25]), .Y(n80) );
  NAND2X0_HVT U159 ( .A1(n79), .A2(n80), .Y(out[25]) );
  INVX0_HVT U160 ( .A(state[25]), .Y(n77) );
  INVX0_HVT U161 ( .A(subkey[25]), .Y(n78) );
  NAND2X0_HVT U162 ( .A1(subkey[121]), .A2(n82), .Y(n83) );
  NAND2X0_HVT U163 ( .A1(n81), .A2(state[121]), .Y(n84) );
  NAND2X0_HVT U164 ( .A1(n83), .A2(n84), .Y(out[121]) );
  INVX0_HVT U165 ( .A(state[121]), .Y(n82) );
  NAND2X0_HVT U166 ( .A1(subkey[90]), .A2(n86), .Y(n87) );
  NAND2X0_HVT U167 ( .A1(n85), .A2(state[90]), .Y(n88) );
  NAND2X0_HVT U168 ( .A1(n87), .A2(n88), .Y(out[90]) );
  INVX0_HVT U169 ( .A(state[90]), .Y(n86) );
  NAND2X0_HVT U170 ( .A1(subkey[32]), .A2(n91), .Y(n92) );
  NAND2X0_HVT U171 ( .A1(n90), .A2(state[32]), .Y(n93) );
  NAND2X0_HVT U172 ( .A1(n92), .A2(n93), .Y(out[32]) );
  INVX0_HVT U173 ( .A(subkey[32]), .Y(n90) );
  INVX0_HVT U174 ( .A(state[32]), .Y(n91) );
  NAND2X0_HVT U175 ( .A1(state[60]), .A2(n95), .Y(n96) );
  NAND2X0_HVT U176 ( .A1(n94), .A2(subkey[60]), .Y(n97) );
  NAND2X0_HVT U177 ( .A1(n96), .A2(n97), .Y(out[60]) );
  INVX0_HVT U178 ( .A(state[60]), .Y(n94) );
  INVX0_HVT U179 ( .A(subkey[60]), .Y(n95) );
  INVX0_HVT U180 ( .A(subkey[67]), .Y(n207) );
  NAND2X0_HVT U181 ( .A1(subkey[24]), .A2(n99), .Y(n100) );
  NAND2X0_HVT U182 ( .A1(n98), .A2(state[24]), .Y(n101) );
  NAND2X0_HVT U183 ( .A1(n100), .A2(n101), .Y(out[24]) );
  INVX0_HVT U184 ( .A(subkey[24]), .Y(n98) );
  INVX0_HVT U185 ( .A(state[24]), .Y(n99) );
  INVX0_HVT U186 ( .A(subkey[83]), .Y(n176) );
  NAND2X0_HVT U187 ( .A1(subkey[22]), .A2(n103), .Y(n104) );
  NAND2X0_HVT U188 ( .A1(n102), .A2(state[22]), .Y(n105) );
  NAND2X0_HVT U189 ( .A1(n104), .A2(n105), .Y(out[22]) );
  INVX0_HVT U190 ( .A(subkey[22]), .Y(n102) );
  INVX0_HVT U191 ( .A(state[22]), .Y(n103) );
  NAND2X0_HVT U192 ( .A1(state[124]), .A2(n107), .Y(n108) );
  NAND2X0_HVT U193 ( .A1(n106), .A2(subkey[124]), .Y(n109) );
  NAND2X0_HVT U194 ( .A1(n108), .A2(n109), .Y(out[124]) );
  INVX0_HVT U195 ( .A(state[124]), .Y(n106) );
  INVX0_HVT U196 ( .A(subkey[124]), .Y(n107) );
  NAND2X0_HVT U197 ( .A1(subkey[56]), .A2(n111), .Y(n112) );
  NAND2X0_HVT U198 ( .A1(n110), .A2(state[56]), .Y(n113) );
  NAND2X0_HVT U199 ( .A1(n112), .A2(n113), .Y(out[56]) );
  INVX0_HVT U200 ( .A(subkey[56]), .Y(n110) );
  INVX0_HVT U201 ( .A(state[56]), .Y(n111) );
  NAND2X0_HVT U202 ( .A1(subkey[81]), .A2(n115), .Y(n116) );
  NAND2X0_HVT U203 ( .A1(n114), .A2(state[81]), .Y(n117) );
  NAND2X0_HVT U204 ( .A1(n116), .A2(n117), .Y(out[81]) );
  INVX0_HVT U205 ( .A(subkey[81]), .Y(n114) );
  INVX0_HVT U206 ( .A(state[81]), .Y(n115) );
  NAND2X0_HVT U207 ( .A1(state[20]), .A2(n228), .Y(n120) );
  NAND2X0_HVT U208 ( .A1(n118), .A2(n119), .Y(n121) );
  NAND2X0_HVT U209 ( .A1(n120), .A2(n121), .Y(out[20]) );
  INVX0_HVT U210 ( .A(state[20]), .Y(n118) );
  INVX0_HVT U211 ( .A(n228), .Y(n119) );
  NAND2X0_HVT U212 ( .A1(subkey[100]), .A2(n123), .Y(n124) );
  NAND2X0_HVT U213 ( .A1(n122), .A2(state[100]), .Y(n125) );
  NAND2X0_HVT U214 ( .A1(n124), .A2(n125), .Y(out[100]) );
  INVX0_HVT U215 ( .A(state[100]), .Y(n123) );
  INVX1_HVT U216 ( .A(state[41]), .Y(n282) );
  NAND2X0_HVT U217 ( .A1(subkey[65]), .A2(n127), .Y(n128) );
  NAND2X0_HVT U218 ( .A1(n126), .A2(state[65]), .Y(n129) );
  NAND2X0_HVT U219 ( .A1(n128), .A2(n129), .Y(out[65]) );
  INVX0_HVT U220 ( .A(subkey[65]), .Y(n126) );
  INVX0_HVT U221 ( .A(state[65]), .Y(n127) );
  NAND2X0_HVT U222 ( .A1(state[1]), .A2(n131), .Y(n132) );
  NAND2X0_HVT U223 ( .A1(n130), .A2(subkey[1]), .Y(n133) );
  NAND2X0_HVT U224 ( .A1(n132), .A2(n133), .Y(out[1]) );
  INVX0_HVT U225 ( .A(state[1]), .Y(n130) );
  NAND2X0_HVT U226 ( .A1(subkey[86]), .A2(n135), .Y(n136) );
  NAND2X0_HVT U227 ( .A1(n134), .A2(state[86]), .Y(n137) );
  NAND2X0_HVT U228 ( .A1(n136), .A2(n137), .Y(out[86]) );
  INVX0_HVT U229 ( .A(subkey[86]), .Y(n134) );
  INVX0_HVT U230 ( .A(state[86]), .Y(n135) );
  NAND2X0_HVT U231 ( .A1(subkey[109]), .A2(n139), .Y(n140) );
  NAND2X0_HVT U232 ( .A1(n138), .A2(state[109]), .Y(n141) );
  NAND2X0_HVT U233 ( .A1(n140), .A2(n141), .Y(out[109]) );
  INVX0_HVT U234 ( .A(subkey[109]), .Y(n138) );
  INVX0_HVT U235 ( .A(state[109]), .Y(n139) );
  NAND2X0_HVT U236 ( .A1(subkey[34]), .A2(n143), .Y(n144) );
  NAND2X0_HVT U237 ( .A1(n142), .A2(state[34]), .Y(n145) );
  NAND2X0_HVT U238 ( .A1(n144), .A2(n145), .Y(out[34]) );
  INVX0_HVT U239 ( .A(subkey[34]), .Y(n142) );
  INVX0_HVT U240 ( .A(state[34]), .Y(n143) );
  XNOR2X2_HVT U241 ( .A1(state[96]), .A2(n146), .Y(out[96]) );
  NAND2X0_HVT U242 ( .A1(state[108]), .A2(n148), .Y(n149) );
  NAND2X0_HVT U243 ( .A1(n147), .A2(subkey[108]), .Y(n150) );
  NAND2X0_HVT U244 ( .A1(n149), .A2(n150), .Y(out[108]) );
  INVX0_HVT U245 ( .A(state[108]), .Y(n147) );
  INVX0_HVT U246 ( .A(subkey[108]), .Y(n148) );
  XNOR2X2_HVT U247 ( .A1(state[116]), .A2(n151), .Y(out[116]) );
  NAND2X0_HVT U248 ( .A1(subkey[58]), .A2(n153), .Y(n154) );
  NAND2X0_HVT U249 ( .A1(n152), .A2(state[58]), .Y(n155) );
  NAND2X0_HVT U250 ( .A1(n154), .A2(n155), .Y(out[58]) );
  INVX0_HVT U251 ( .A(subkey[58]), .Y(n152) );
  INVX0_HVT U252 ( .A(state[58]), .Y(n153) );
  INVX0_HVT U253 ( .A(state[59]), .Y(n291) );
  NAND2X0_HVT U254 ( .A1(subkey[71]), .A2(n157), .Y(n158) );
  NAND2X0_HVT U255 ( .A1(n156), .A2(state[71]), .Y(n159) );
  NAND2X0_HVT U256 ( .A1(n158), .A2(n159), .Y(out[71]) );
  INVX0_HVT U257 ( .A(subkey[71]), .Y(n156) );
  INVX0_HVT U258 ( .A(state[71]), .Y(n157) );
  INVX1_HVT U259 ( .A(subkey[36]), .Y(n220) );
  INVX0_HVT U260 ( .A(subkey[19]), .Y(n249) );
  NAND2X0_HVT U261 ( .A1(state[99]), .A2(n161), .Y(n162) );
  NAND2X0_HVT U262 ( .A1(n160), .A2(subkey[99]), .Y(n163) );
  NAND2X0_HVT U263 ( .A1(n162), .A2(n163), .Y(out[99]) );
  INVX0_HVT U264 ( .A(state[99]), .Y(n160) );
  IBUFFX2_HVT U265 ( .A(subkey[99]), .Y(n161) );
  NAND2X0_HVT U266 ( .A1(state[35]), .A2(n244), .Y(n165) );
  NAND2X0_HVT U267 ( .A1(n164), .A2(subkey[35]), .Y(n166) );
  NAND2X0_HVT U268 ( .A1(n165), .A2(n166), .Y(out[35]) );
  INVX0_HVT U269 ( .A(state[35]), .Y(n164) );
  NAND2X0_HVT U270 ( .A1(subkey[62]), .A2(n168), .Y(n169) );
  NAND2X0_HVT U271 ( .A1(n167), .A2(state[62]), .Y(n170) );
  NAND2X0_HVT U272 ( .A1(n169), .A2(n170), .Y(out[62]) );
  INVX0_HVT U273 ( .A(subkey[62]), .Y(n167) );
  INVX0_HVT U274 ( .A(state[62]), .Y(n168) );
  NAND2X0_HVT U275 ( .A1(subkey[46]), .A2(n172), .Y(n173) );
  NAND2X0_HVT U276 ( .A1(n171), .A2(state[46]), .Y(n174) );
  NAND2X0_HVT U277 ( .A1(n173), .A2(n174), .Y(out[46]) );
  INVX0_HVT U278 ( .A(subkey[46]), .Y(n171) );
  INVX0_HVT U279 ( .A(state[46]), .Y(n172) );
  INVX1_HVT U280 ( .A(subkey[66]), .Y(n193) );
  NAND2X0_HVT U281 ( .A1(state[83]), .A2(n176), .Y(n177) );
  NAND2X0_HVT U282 ( .A1(n175), .A2(subkey[83]), .Y(n178) );
  NAND2X0_HVT U283 ( .A1(n177), .A2(n178), .Y(out[83]) );
  INVX0_HVT U284 ( .A(state[83]), .Y(n175) );
  NAND2X0_HVT U285 ( .A1(state[75]), .A2(n267), .Y(n179) );
  NAND2X0_HVT U286 ( .A1(n180), .A2(n179), .Y(out[75]) );
  NAND2X0_HVT U287 ( .A1(subkey[61]), .A2(n182), .Y(n183) );
  NAND2X0_HVT U288 ( .A1(n181), .A2(state[61]), .Y(n184) );
  NAND2X0_HVT U289 ( .A1(n183), .A2(n184), .Y(out[61]) );
  INVX0_HVT U290 ( .A(subkey[61]), .Y(n181) );
  INVX0_HVT U291 ( .A(state[61]), .Y(n182) );
  NAND2X0_HVT U292 ( .A1(state[45]), .A2(n186), .Y(n187) );
  NAND2X0_HVT U293 ( .A1(n185), .A2(subkey[45]), .Y(n188) );
  NAND2X0_HVT U294 ( .A1(n187), .A2(n188), .Y(out[45]) );
  INVX0_HVT U295 ( .A(state[45]), .Y(n185) );
  INVX0_HVT U296 ( .A(subkey[45]), .Y(n186) );
  NAND2X0_HVT U297 ( .A1(state[84]), .A2(n190), .Y(n191) );
  NAND2X0_HVT U298 ( .A1(n189), .A2(subkey[84]), .Y(n192) );
  NAND2X0_HVT U299 ( .A1(n191), .A2(n192), .Y(out[84]) );
  INVX0_HVT U300 ( .A(state[84]), .Y(n189) );
  INVX0_HVT U301 ( .A(subkey[84]), .Y(n190) );
  XNOR2X2_HVT U302 ( .A1(state[66]), .A2(n193), .Y(out[66]) );
  NAND2X0_HVT U303 ( .A1(subkey[4]), .A2(n195), .Y(n196) );
  NAND2X0_HVT U304 ( .A1(n194), .A2(state[4]), .Y(n197) );
  NAND2X0_HVT U305 ( .A1(n196), .A2(n197), .Y(out[4]) );
  INVX0_HVT U306 ( .A(subkey[4]), .Y(n194) );
  NAND2X0_HVT U307 ( .A1(subkey[79]), .A2(n199), .Y(n200) );
  NAND2X0_HVT U308 ( .A1(n198), .A2(state[79]), .Y(n201) );
  NAND2X0_HVT U309 ( .A1(n200), .A2(n201), .Y(out[79]) );
  INVX0_HVT U310 ( .A(subkey[79]), .Y(n198) );
  INVX0_HVT U311 ( .A(state[79]), .Y(n199) );
  INVX0_HVT U312 ( .A(subkey[27]), .Y(n289) );
  NAND2X0_HVT U313 ( .A1(state[12]), .A2(n203), .Y(n204) );
  NAND2X0_HVT U314 ( .A1(n202), .A2(subkey[12]), .Y(n205) );
  NAND2X0_HVT U315 ( .A1(n204), .A2(n205), .Y(out[12]) );
  INVX0_HVT U316 ( .A(state[12]), .Y(n202) );
  INVX0_HVT U317 ( .A(subkey[12]), .Y(n203) );
  XNOR2X2_HVT U318 ( .A1(n207), .A2(state[67]), .Y(out[67]) );
  NAND2X0_HVT U319 ( .A1(subkey[113]), .A2(n209), .Y(n210) );
  NAND2X0_HVT U320 ( .A1(n208), .A2(state[113]), .Y(n211) );
  NAND2X0_HVT U321 ( .A1(n210), .A2(n211), .Y(out[113]) );
  IBUFFX2_HVT U322 ( .A(subkey[113]), .Y(n208) );
  INVX0_HVT U323 ( .A(state[113]), .Y(n209) );
  NAND2X0_HVT U324 ( .A1(subkey[94]), .A2(n213), .Y(n214) );
  NAND2X0_HVT U325 ( .A1(n212), .A2(state[94]), .Y(n215) );
  NAND2X0_HVT U326 ( .A1(n214), .A2(n215), .Y(out[94]) );
  INVX0_HVT U327 ( .A(subkey[94]), .Y(n212) );
  INVX0_HVT U328 ( .A(state[94]), .Y(n213) );
  INVX0_HVT U329 ( .A(state[57]), .Y(n260) );
  NAND2X0_HVT U330 ( .A1(subkey[77]), .A2(n217), .Y(n218) );
  NAND2X0_HVT U331 ( .A1(n216), .A2(state[77]), .Y(n219) );
  NAND2X0_HVT U332 ( .A1(n218), .A2(n219), .Y(out[77]) );
  INVX0_HVT U333 ( .A(subkey[77]), .Y(n216) );
  INVX0_HVT U334 ( .A(state[77]), .Y(n217) );
  OR2X1_HVT U335 ( .A1(n220), .A2(state[36]), .Y(n275) );
  NAND2X0_HVT U336 ( .A1(subkey[31]), .A2(n222), .Y(n223) );
  NAND2X0_HVT U337 ( .A1(n221), .A2(state[31]), .Y(n224) );
  NAND2X0_HVT U338 ( .A1(n223), .A2(n224), .Y(out[31]) );
  IBUFFX2_HVT U339 ( .A(subkey[31]), .Y(n221) );
  INVX0_HVT U340 ( .A(state[31]), .Y(n222) );
  NAND2X0_HVT U341 ( .A1(state[27]), .A2(n289), .Y(n226) );
  NAND2X0_HVT U342 ( .A1(n225), .A2(subkey[27]), .Y(n227) );
  NAND2X0_HVT U343 ( .A1(n226), .A2(n227), .Y(out[27]) );
  INVX0_HVT U344 ( .A(state[27]), .Y(n225) );
  XOR2X2_HVT U345 ( .A1(subkey[110]), .A2(state[110]), .Y(out[110]) );
  NAND2X0_HVT U346 ( .A1(subkey[89]), .A2(n230), .Y(n231) );
  NAND2X0_HVT U347 ( .A1(state[89]), .A2(n229), .Y(n232) );
  NAND2X0_HVT U348 ( .A1(n231), .A2(n232), .Y(out[89]) );
  INVX0_HVT U349 ( .A(subkey[89]), .Y(n229) );
  INVX0_HVT U350 ( .A(state[89]), .Y(n230) );
  NAND2X0_HVT U351 ( .A1(subkey[73]), .A2(n234), .Y(n235) );
  NAND2X0_HVT U352 ( .A1(n233), .A2(state[73]), .Y(n236) );
  NAND2X0_HVT U353 ( .A1(n235), .A2(n236), .Y(out[73]) );
  INVX0_HVT U354 ( .A(subkey[73]), .Y(n233) );
  INVX0_HVT U355 ( .A(state[73]), .Y(n234) );
  NAND2X0_HVT U356 ( .A1(state[123]), .A2(n238), .Y(n239) );
  NAND2X0_HVT U357 ( .A1(n237), .A2(subkey[123]), .Y(n240) );
  NAND2X0_HVT U358 ( .A1(n239), .A2(n240), .Y(out[123]) );
  INVX0_HVT U359 ( .A(state[123]), .Y(n237) );
  INVX0_HVT U360 ( .A(subkey[123]), .Y(n238) );
  NAND2X0_HVT U361 ( .A1(n241), .A2(state[52]), .Y(n243) );
  NAND2X0_HVT U362 ( .A1(n242), .A2(n243), .Y(out[52]) );
  IBUFFX2_HVT U363 ( .A(subkey[52]), .Y(n241) );
  NAND2X0_HVT U364 ( .A1(subkey[39]), .A2(n246), .Y(n247) );
  NAND2X0_HVT U365 ( .A1(state[39]), .A2(n245), .Y(n248) );
  NAND2X0_HVT U366 ( .A1(n247), .A2(n248), .Y(out[39]) );
  INVX0_HVT U367 ( .A(state[39]), .Y(n246) );
  XNOR2X2_HVT U368 ( .A1(state[19]), .A2(n249), .Y(out[19]) );
  INVX0_HVT U369 ( .A(subkey[92]), .Y(n298) );
  INVX1_HVT U370 ( .A(subkey[3]), .Y(n302) );
  INVX0_HVT U371 ( .A(subkey[68]), .Y(n274) );
  INVX0_HVT U372 ( .A(subkey[11]), .Y(n255) );
  INVX0_HVT U373 ( .A(subkey[91]), .Y(n268) );
  INVX0_HVT U374 ( .A(subkey[97]), .Y(n294) );
  INVX0_HVT U375 ( .A(subkey[125]), .Y(n251) );
  INVX0_HVT U376 ( .A(subkey[41]), .Y(n281) );
  INVX0_HVT U377 ( .A(subkey[95]), .Y(n263) );
  NAND2X0_HVT U378 ( .A1(subkey[125]), .A2(n252), .Y(n253) );
  NAND2X0_HVT U379 ( .A1(state[125]), .A2(n251), .Y(n254) );
  NAND2X0_HVT U380 ( .A1(n253), .A2(n254), .Y(out[125]) );
  INVX0_HVT U381 ( .A(state[125]), .Y(n252) );
  NAND2X0_HVT U382 ( .A1(subkey[11]), .A2(n256), .Y(n257) );
  NAND2X0_HVT U383 ( .A1(n255), .A2(state[11]), .Y(n258) );
  NAND2X0_HVT U384 ( .A1(n257), .A2(n258), .Y(out[11]) );
  INVX0_HVT U385 ( .A(state[11]), .Y(n256) );
  NAND2X0_HVT U386 ( .A1(subkey[57]), .A2(n260), .Y(n261) );
  NAND2X0_HVT U387 ( .A1(state[57]), .A2(n259), .Y(n262) );
  NAND2X0_HVT U388 ( .A1(n261), .A2(n262), .Y(out[57]) );
  INVX0_HVT U389 ( .A(subkey[57]), .Y(n259) );
  XOR2X2_HVT U390 ( .A1(state[78]), .A2(subkey[78]), .Y(out[78]) );
  NAND2X0_HVT U391 ( .A1(subkey[95]), .A2(n264), .Y(n265) );
  NAND2X0_HVT U392 ( .A1(n263), .A2(state[95]), .Y(n266) );
  NAND2X0_HVT U393 ( .A1(n265), .A2(n266), .Y(out[95]) );
  INVX0_HVT U394 ( .A(state[95]), .Y(n264) );
  NAND2X0_HVT U395 ( .A1(subkey[91]), .A2(n269), .Y(n270) );
  NAND2X0_HVT U396 ( .A1(state[91]), .A2(n268), .Y(n271) );
  NAND2X0_HVT U397 ( .A1(n270), .A2(n271), .Y(out[91]) );
  INVX0_HVT U398 ( .A(state[91]), .Y(n269) );
  NAND2X0_HVT U399 ( .A1(n274), .A2(state[68]), .Y(n272) );
  NAND2X0_HVT U400 ( .A1(n272), .A2(n273), .Y(out[68]) );
  XOR2X2_HVT U401 ( .A1(subkey[63]), .A2(state[63]), .Y(out[63]) );
  NAND2X0_HVT U402 ( .A1(n220), .A2(state[36]), .Y(n276) );
  NAND2X0_HVT U403 ( .A1(n276), .A2(n275), .Y(out[36]) );
  INVX1_HVT U404 ( .A(state[53]), .Y(n310) );
  NAND2X0_HVT U405 ( .A1(subkey[51]), .A2(n278), .Y(n279) );
  NAND2X0_HVT U406 ( .A1(state[51]), .A2(n277), .Y(n280) );
  NAND2X0_HVT U407 ( .A1(n279), .A2(n280), .Y(out[51]) );
  INVX0_HVT U408 ( .A(state[51]), .Y(n278) );
  INVX0_HVT U409 ( .A(subkey[59]), .Y(n290) );
  NAND2X0_HVT U410 ( .A1(subkey[41]), .A2(n282), .Y(n283) );
  NAND2X0_HVT U411 ( .A1(state[41]), .A2(n281), .Y(n284) );
  NAND2X0_HVT U412 ( .A1(n284), .A2(n283), .Y(out[41]) );
  NAND2X0_HVT U413 ( .A1(subkey[43]), .A2(n286), .Y(n287) );
  NAND2X0_HVT U414 ( .A1(state[43]), .A2(n285), .Y(n288) );
  NAND2X0_HVT U415 ( .A1(n287), .A2(n288), .Y(out[43]) );
  INVX0_HVT U416 ( .A(state[43]), .Y(n286) );
  XOR2X2_HVT U417 ( .A1(state[5]), .A2(subkey[5]), .Y(out[5]) );
  INVX1_HVT U418 ( .A(state[3]), .Y(n303) );
  NAND2X0_HVT U419 ( .A1(subkey[59]), .A2(n291), .Y(n292) );
  NAND2X0_HVT U420 ( .A1(n290), .A2(state[59]), .Y(n293) );
  NAND2X0_HVT U421 ( .A1(n292), .A2(n293), .Y(out[59]) );
  NAND2X0_HVT U422 ( .A1(subkey[97]), .A2(n295), .Y(n296) );
  NAND2X0_HVT U423 ( .A1(n294), .A2(state[97]), .Y(n297) );
  NAND2X0_HVT U424 ( .A1(n296), .A2(n297), .Y(out[97]) );
  INVX0_HVT U425 ( .A(state[97]), .Y(n295) );
  NAND2X0_HVT U426 ( .A1(subkey[92]), .A2(n299), .Y(n300) );
  NAND2X0_HVT U427 ( .A1(n298), .A2(state[92]), .Y(n301) );
  NAND2X0_HVT U428 ( .A1(n300), .A2(n301), .Y(out[92]) );
  INVX0_HVT U429 ( .A(state[92]), .Y(n299) );
  NAND2X0_HVT U430 ( .A1(subkey[3]), .A2(n303), .Y(n304) );
  NAND2X0_HVT U431 ( .A1(n302), .A2(state[3]), .Y(n305) );
  NAND2X0_HVT U432 ( .A1(n304), .A2(n305), .Y(out[3]) );
  NAND2X0_HVT U433 ( .A1(subkey[115]), .A2(n307), .Y(n308) );
  NAND2X0_HVT U434 ( .A1(n306), .A2(state[115]), .Y(n309) );
  NAND2X0_HVT U435 ( .A1(n309), .A2(n308), .Y(out[115]) );
  INVX0_HVT U436 ( .A(subkey[115]), .Y(n306) );
  INVX0_HVT U437 ( .A(state[115]), .Y(n307) );
  XNOR2X2_HVT U438 ( .A1(subkey[53]), .A2(n310), .Y(out[53]) );
endmodule

