
module inv_sbox_8 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n1, n52, n58, n83, n196, n197, n198, n199, n200, n201, n202, n205,
         n208, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624;

  NAND2X0_HVT U4 ( .A1(n312), .A2(n351), .Y(n622) );
  NAND2X0_HVT U5 ( .A1(n622), .A2(n302), .Y(n621) );
  NAND2X0_HVT U6 ( .A1(n354), .A2(n236), .Y(n619) );
  NAND2X0_HVT U8 ( .A1(n353), .A2(n303), .Y(n617) );
  NAND2X0_HVT U9 ( .A1(n237), .A2(n617), .Y(n616) );
  NAND2X0_HVT U10 ( .A1(n236), .A2(n614), .Y(n615) );
  NAND2X0_HVT U11 ( .A1(n264), .A2(n352), .Y(n613) );
  NAND2X0_HVT U12 ( .A1(n281), .A2(n341), .Y(n612) );
  NAND2X0_HVT U13 ( .A1(n349), .A2(n267), .Y(n611) );
  NAND2X0_HVT U15 ( .A1(n315), .A2(n353), .Y(n609) );
  NAND2X0_HVT U19 ( .A1(n356), .A2(n419), .Y(n604) );
  NAND2X0_HVT U32 ( .A1(n318), .A2(n358), .Y(n592) );
  NAND2X0_HVT U35 ( .A1(n617), .A2(n420), .Y(n589) );
  NAND2X0_HVT U38 ( .A1(n341), .A2(n264), .Y(n586) );
  NAND2X0_HVT U42 ( .A1(n619), .A2(n420), .Y(n582) );
  NAND2X0_HVT U55 ( .A1(n349), .A2(n622), .Y(n571) );
  MUX41X1_HVT U56 ( .A1(n402), .A3(n315), .A2(n389), .A4(n571), .S0(n334), 
        .S1(n363), .Y(n570) );
  AO21X1_HVT U60 ( .A1(n566), .A2(n337), .A3(n603), .Y(n567) );
  NAND2X0_HVT U66 ( .A1(n353), .A2(n306), .Y(n560) );
  MUX41X1_HVT U67 ( .A1(n381), .A3(n403), .A2(n383), .A4(n560), .S0(n339), 
        .S1(n359), .Y(n559) );
  MUX41X1_HVT U69 ( .A1(n558), .A3(n561), .A2(n559), .A4(n562), .S0(in[5]), 
        .S1(n344), .Y(n557) );
  MUX41X1_HVT U71 ( .A1(n288), .A3(n241), .A2(n613), .A4(n377), .S0(n333), 
        .S1(n279), .Y(n556) );
  NAND2X0_HVT U72 ( .A1(n347), .A2(n618), .Y(n555) );
  MUX41X1_HVT U73 ( .A1(n597), .A3(n555), .A2(n307), .A4(n340), .S0(n338), 
        .S1(n331), .Y(n554) );
  MUX41X1_HVT U74 ( .A1(n615), .A3(n393), .A2(n392), .A4(n387), .S0(n334), 
        .S1(n362), .Y(n553) );
  OA21X1_HVT U76 ( .A1(n370), .A2(n364), .A3(n603), .Y(n551) );
  MUX41X1_HVT U80 ( .A1(n405), .A3(n402), .A2(n616), .A4(n621), .S0(n333), 
        .S1(n363), .Y(n547) );
  NAND2X0_HVT U81 ( .A1(n352), .A2(n618), .Y(n546) );
  MUX41X1_HVT U84 ( .A1(n329), .A3(n391), .A2(n406), .A4(n599), .S0(n334), 
        .S1(n362), .Y(n544) );
  MUX41X1_HVT U87 ( .A1(n371), .A3(n329), .A2(n407), .A4(n389), .S0(n332), 
        .S1(n363), .Y(n542) );
  MUX41X1_HVT U88 ( .A1(n383), .A3(n368), .A2(n594), .A4(n578), .S0(n333), 
        .S1(n278), .Y(n541) );
  NAND2X0_HVT U89 ( .A1(n264), .A2(n300), .Y(n540) );
  MUX41X1_HVT U90 ( .A1(n242), .A3(n618), .A2(n577), .A4(n540), .S0(n333), 
        .S1(n363), .Y(n539) );
  MUX41X1_HVT U95 ( .A1(n535), .A3(n541), .A2(n539), .A4(n542), .S0(in[5]), 
        .S1(n345), .Y(n534) );
  MUX41X1_HVT U96 ( .A1(n403), .A3(n611), .A2(n390), .A4(n408), .S0(n334), 
        .S1(n278), .Y(n533) );
  MUX41X1_HVT U98 ( .A1(n532), .A3(n409), .A2(n395), .A4(n596), .S0(n334), 
        .S1(n278), .Y(n531) );
  MUX41X1_HVT U99 ( .A1(n592), .A3(n385), .A2(n576), .A4(n347), .S0(n361), 
        .S1(n359), .Y(n530) );
  NAND2X0_HVT U100 ( .A1(n358), .A2(n416), .Y(n529) );
  MUX41X1_HVT U101 ( .A1(n410), .A3(n612), .A2(n394), .A4(n529), .S0(n363), 
        .S1(n359), .Y(n528) );
  MUX41X1_HVT U102 ( .A1(n528), .A3(n531), .A2(n530), .A4(n533), .S0(n295), 
        .S1(n344), .Y(n527) );
  AND2X1_HVT U104 ( .A1(n618), .A2(n302), .Y(n526) );
  MUX41X1_HVT U105 ( .A1(n610), .A3(n411), .A2(n546), .A4(n526), .S0(n334), 
        .S1(n362), .Y(n525) );
  MUX41X1_HVT U107 ( .A1(n410), .A3(n623), .A2(n524), .A4(n199), .S0(n333), 
        .S1(n279), .Y(n523) );
  MUX41X1_HVT U109 ( .A1(n409), .A3(n368), .A2(n406), .A4(n400), .S0(n333), 
        .S1(n363), .Y(n521) );
  MUX41X1_HVT U110 ( .A1(n521), .A3(n523), .A2(n522), .A4(n525), .S0(n295), 
        .S1(n345), .Y(n520) );
  NAND2X0_HVT U114 ( .A1(n237), .A2(n618), .Y(n516) );
  MUX41X1_HVT U115 ( .A1(n516), .A3(n613), .A2(n397), .A4(n623), .S0(n278), 
        .S1(n359), .Y(n515) );
  MUX41X1_HVT U116 ( .A1(n396), .A3(n391), .A2(n368), .A4(n609), .S0(n332), 
        .S1(n363), .Y(n514) );
  NAND2X0_HVT U118 ( .A1(n264), .A2(n296), .Y(n512) );
  MUX41X1_HVT U119 ( .A1(n412), .A3(n513), .A2(n587), .A4(n512), .S0(n332), 
        .S1(n278), .Y(n511) );
  MUX41X1_HVT U120 ( .A1(n511), .A3(n515), .A2(n514), .A4(n517), .S0(n295), 
        .S1(n345), .Y(n510) );
  MUX41X1_HVT U122 ( .A1(n401), .A3(n325), .A2(n578), .A4(n404), .S0(n332), 
        .S1(n279), .Y(n509) );
  MUX41X1_HVT U124 ( .A1(n327), .A3(n508), .A2(n601), .A4(n314), .S0(n337), 
        .S1(n332), .Y(n507) );
  AOI21X1_HVT U127 ( .A1(n336), .A2(n503), .A3(n375), .Y(n504) );
  NAND2X0_HVT U129 ( .A1(n334), .A2(n236), .Y(n501) );
  MUX41X1_HVT U130 ( .A1(n501), .A3(n502), .A2(n505), .A4(n504), .S0(n339), 
        .S1(n345), .Y(n500) );
  AND2X1_HVT U131 ( .A1(n306), .A2(n264), .Y(n499) );
  MUX41X1_HVT U132 ( .A1(n372), .A3(n499), .A2(n414), .A4(n381), .S0(n338), 
        .S1(n331), .Y(n498) );
  MUX41X1_HVT U133 ( .A1(n415), .A3(n199), .A2(n571), .A4(n373), .S0(n337), 
        .S1(n331), .Y(n497) );
  MUX41X1_HVT U136 ( .A1(n575), .A3(n529), .A2(n495), .A4(n379), .S0(n359), 
        .S1(n279), .Y(n494) );
  MUX41X1_HVT U137 ( .A1(n267), .A3(n595), .A2(n599), .A4(n408), .S0(n339), 
        .S1(n336), .Y(n493) );
  MUX41X1_HVT U139 ( .A1(n492), .A3(n496), .A2(n500), .A4(n506), .S0(n295), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n392), .A3(n326), .A2(n388), .A4(n613), .S0(n338), 
        .S1(n359), .Y(n491) );
  NAND2X0_HVT U141 ( .A1(n315), .A2(n358), .Y(n490) );
  MUX41X1_HVT U143 ( .A1(n299), .A3(n289), .A2(n604), .A4(n601), .S0(n335), 
        .S1(n279), .Y(n488) );
  MUX41X1_HVT U145 ( .A1(n593), .A3(n411), .A2(n487), .A4(n546), .S0(n336), 
        .S1(n279), .Y(n486) );
  MUX41X1_HVT U146 ( .A1(n486), .A3(n488), .A2(n489), .A4(n491), .S0(n344), 
        .S1(n295), .Y(n485) );
  AO21X1_HVT U148 ( .A1(n339), .A2(n376), .A3(n416), .Y(n483) );
  MUX41X1_HVT U151 ( .A1(n313), .A3(n395), .A2(n304), .A4(n481), .S0(n337), 
        .S1(n335), .Y(n480) );
  MUX41X1_HVT U155 ( .A1(n388), .A3(n613), .A2(n605), .A4(n390), .S0(n335), 
        .S1(n362), .Y(n476) );
  MUX41X1_HVT U156 ( .A1(n476), .A3(n480), .A2(n477), .A4(n482), .S0(n295), 
        .S1(n345), .Y(n475) );
  NAND2X0_HVT U159 ( .A1(n472), .A2(n471), .Y(n473) );
  NAND2X0_HVT U163 ( .A1(n284), .A2(n300), .Y(n467) );
  MUX41X1_HVT U164 ( .A1(n616), .A3(n467), .A2(n587), .A4(n387), .S0(n332), 
        .S1(n362), .Y(n466) );
  NAND2X0_HVT U166 ( .A1(n614), .A2(n463), .Y(n464) );
  MUX41X1_HVT U170 ( .A1(n328), .A3(n324), .A2(n327), .A4(n460), .S0(n335), 
        .S1(n279), .Y(n459) );
  MUX41X1_HVT U172 ( .A1(n540), .A3(n458), .A2(n324), .A4(n602), .S0(n335), 
        .S1(n278), .Y(n457) );
  MUX41X1_HVT U174 ( .A1(n407), .A3(n571), .A2(n415), .A4(n420), .S0(n335), 
        .S1(n362), .Y(n455) );
  NAND2X0_HVT U177 ( .A1(n355), .A2(n296), .Y(n453) );
  AND2X1_HVT U179 ( .A1(n288), .A2(n303), .Y(n451) );
  MUX41X1_HVT U180 ( .A1(n592), .A3(n366), .A2(n451), .A4(n579), .S0(n335), 
        .S1(n278), .Y(n450) );
  MUX41X1_HVT U182 ( .A1(n374), .A3(n622), .A2(n371), .A4(n313), .S0(n332), 
        .S1(n362), .Y(n448) );
  MUX41X1_HVT U183 ( .A1(n289), .A3(n402), .A2(n387), .A4(n201), .S0(n337), 
        .S1(n331), .Y(n447) );
  AND2X1_HVT U185 ( .A1(n420), .A2(n264), .Y(n445) );
  OA21X1_HVT U189 ( .A1(n391), .A2(n364), .A3(n566), .Y(n441) );
  NAND2X0_HVT U191 ( .A1(n364), .A2(n380), .Y(n439) );
  AND2X1_HVT U192 ( .A1(n393), .A2(n437), .Y(n438) );
  NAND2X0_HVT U194 ( .A1(n201), .A2(n437), .Y(n435) );
  NAND2X0_HVT U198 ( .A1(n355), .A2(n420), .Y(n614) );
  NAND2X0_HVT U200 ( .A1(n303), .A2(n264), .Y(n503) );
  AO21X1_HVT U204 ( .A1(n347), .A2(n622), .A3(n364), .Y(n463) );
  NAND2X0_HVT U207 ( .A1(n264), .A2(n242), .Y(n566) );
  MUX21X1_HVT U1 ( .A1(n58), .A2(n52), .S0(n83), .Y(n1) );
  IBUFFX16_HVT U2 ( .A(n416), .Y(n52) );
  IBUFFX16_HVT U3 ( .A(n419), .Y(n58) );
  IBUFFX16_HVT U7 ( .A(n285), .Y(n83) );
  MUX21X2_HVT U14 ( .A1(n510), .A2(n520), .S0(n196), .Y(out[3]) );
  IBUFFX16_HVT U16 ( .A(n297), .Y(n196) );
  MUX41X1_HVT U17 ( .A1(n315), .A3(n387), .A2(n350), .A4(n389), .S0(n197), 
        .S1(n278), .Y(n522) );
  IBUFFX16_HVT U18 ( .A(n334), .Y(n197) );
  INVX1_HVT U20 ( .A(n374), .Y(n198) );
  INVX1_HVT U21 ( .A(n198), .Y(n199) );
  INVX0_HVT U22 ( .A(n582), .Y(n200) );
  INVX0_HVT U23 ( .A(n200), .Y(n201) );
  NAND2X0_HVT U24 ( .A1(n448), .A2(n202), .Y(n205) );
  NAND2X0_HVT U25 ( .A1(n447), .A2(n294), .Y(n208) );
  NAND2X0_HVT U26 ( .A1(n205), .A2(n208), .Y(n446) );
  IBUFFX2_HVT U27 ( .A(n294), .Y(n202) );
  INVX0_HVT U28 ( .A(in[1]), .Y(n294) );
  MUX21X2_HVT U29 ( .A1(n567), .A2(n568), .S0(n218), .Y(n565) );
  IBUFFX16_HVT U30 ( .A(n334), .Y(n218) );
  MUX21X1_HVT U31 ( .A1(n414), .A2(n372), .S0(n337), .Y(n484) );
  NAND2X0_HVT U33 ( .A1(n551), .A2(n219), .Y(n220) );
  NAND2X0_HVT U34 ( .A1(n552), .A2(n266), .Y(n221) );
  NAND2X0_HVT U36 ( .A1(n220), .A2(n221), .Y(n550) );
  INVX0_HVT U37 ( .A(n266), .Y(n219) );
  NAND2X0_HVT U39 ( .A1(n549), .A2(n222), .Y(n223) );
  NAND2X0_HVT U40 ( .A1(n543), .A2(n230), .Y(n224) );
  NAND2X0_HVT U41 ( .A1(n223), .A2(n224), .Y(out[1]) );
  INVX1_HVT U43 ( .A(n230), .Y(n222) );
  IBUFFX2_HVT U44 ( .A(n336), .Y(n266) );
  IBUFFX2_HVT U45 ( .A(in[7]), .Y(n230) );
  NBUFFX4_HVT U46 ( .A(n608), .Y(n347) );
  INVX0_HVT U47 ( .A(n295), .Y(n248) );
  INVX2_HVT U48 ( .A(n322), .Y(n608) );
  MUX21X2_HVT U49 ( .A1(n296), .A2(n349), .S0(n312), .Y(n289) );
  INVX0_HVT U50 ( .A(n361), .Y(n320) );
  INVX0_HVT U51 ( .A(n365), .Y(n361) );
  IBUFFX16_HVT U52 ( .A(n365), .Y(n362) );
  INVX1_HVT U53 ( .A(n322), .Y(n315) );
  NBUFFX4_HVT U54 ( .A(n417), .Y(n340) );
  INVX1_HVT U57 ( .A(n357), .Y(n354) );
  MUX21X2_HVT U58 ( .A1(n343), .A2(n420), .S0(n355), .Y(n588) );
  MUX41X1_HVT U59 ( .A1(n469), .A3(n589), .A2(n386), .A4(n398), .S0(n225), 
        .S1(n320), .Y(n468) );
  IBUFFX16_HVT U61 ( .A(n335), .Y(n225) );
  NAND2X0_HVT U62 ( .A1(n518), .A2(n226), .Y(n227) );
  NAND2X0_HVT U63 ( .A1(n519), .A2(n336), .Y(n228) );
  NAND2X0_HVT U64 ( .A1(n227), .A2(n228), .Y(n517) );
  IBUFFX2_HVT U65 ( .A(n336), .Y(n226) );
  AO21X1_HVT U68 ( .A1(n397), .A2(n338), .A3(n600), .Y(n518) );
  MUX21X1_HVT U70 ( .A1(n375), .A2(n583), .S0(n339), .Y(n519) );
  MUX21X1_HVT U75 ( .A1(n387), .A2(n563), .S0(n330), .Y(n562) );
  INVX1_HVT U77 ( .A(n330), .Y(n259) );
  MUX21X1_HVT U78 ( .A1(n478), .A2(n479), .S0(n336), .Y(n477) );
  MUX41X1_HVT U79 ( .A1(n440), .A3(n449), .A2(n434), .A4(n446), .S0(n229), 
        .S1(n346), .Y(out[7]) );
  IBUFFX16_HVT U82 ( .A(n297), .Y(n229) );
  INVX1_HVT U83 ( .A(n583), .Y(n311) );
  MUX21X2_HVT U85 ( .A1(n306), .A2(n419), .S0(n312), .Y(n583) );
  NAND2X0_HVT U86 ( .A1(n231), .A2(n341), .Y(n620) );
  IBUFFX16_HVT U91 ( .A(n318), .Y(n231) );
  IBUFFX2_HVT U92 ( .A(n341), .Y(n296) );
  NAND2X0_HVT U93 ( .A1(n352), .A2(n232), .Y(n233) );
  NAND2X0_HVT U94 ( .A1(n303), .A2(n235), .Y(n234) );
  NAND2X0_HVT U97 ( .A1(n233), .A2(n234), .Y(n422) );
  INVX4_HVT U103 ( .A(n235), .Y(n232) );
  IBUFFX2_HVT U106 ( .A(n284), .Y(n235) );
  INVX0_HVT U108 ( .A(n422), .Y(n414) );
  INVX2_HVT U111 ( .A(n298), .Y(n299) );
  INVX1_HVT U112 ( .A(n243), .Y(n236) );
  INVX1_HVT U113 ( .A(n243), .Y(n237) );
  INVX0_HVT U117 ( .A(n243), .Y(n238) );
  INVX0_HVT U121 ( .A(n418), .Y(n239) );
  INVX0_HVT U123 ( .A(n418), .Y(n240) );
  INVX1_HVT U125 ( .A(n239), .Y(n241) );
  INVX1_HVT U126 ( .A(n240), .Y(n242) );
  AND2X1_HVT U128 ( .A1(n265), .A2(n275), .Y(n243) );
  INVX2_HVT U134 ( .A(n608), .Y(n420) );
  INVX0_HVT U135 ( .A(n298), .Y(n300) );
  INVX1_HVT U138 ( .A(n346), .Y(n295) );
  IBUFFX2_HVT U142 ( .A(n365), .Y(n363) );
  IBUFFX2_HVT U144 ( .A(n319), .Y(n593) );
  MUX21X1_HVT U147 ( .A1(n314), .A2(n571), .S0(n338), .Y(n568) );
  MUX21X2_HVT U149 ( .A1(n260), .A2(n600), .S0(n259), .Y(n258) );
  MUX21X2_HVT U150 ( .A1(n306), .A2(n242), .S0(n356), .Y(n600) );
  MUX21X2_HVT U152 ( .A1(n534), .A2(n527), .S0(n244), .Y(out[2]) );
  IBUFFX16_HVT U153 ( .A(n254), .Y(n244) );
  MUX21X2_HVT U154 ( .A1(n238), .A2(n420), .S0(n358), .Y(n319) );
  NAND2X0_HVT U157 ( .A1(n329), .A2(n245), .Y(n246) );
  NAND2X0_HVT U158 ( .A1(n576), .A2(n339), .Y(n247) );
  NAND2X0_HVT U160 ( .A1(n246), .A2(n247), .Y(n443) );
  IBUFFX2_HVT U161 ( .A(n339), .Y(n245) );
  XOR2X1_HVT U162 ( .A1(n302), .A2(n312), .Y(n576) );
  MUX41X1_HVT U165 ( .A1(n457), .A3(n455), .A2(n459), .A4(n456), .S0(n248), 
        .S1(n249), .Y(n454) );
  IBUFFX16_HVT U167 ( .A(n294), .Y(n249) );
  NAND2X0_HVT U168 ( .A1(n315), .A2(n250), .Y(n251) );
  NAND2X0_HVT U169 ( .A1(n343), .A2(n338), .Y(n252) );
  NAND2X0_HVT U171 ( .A1(n251), .A2(n252), .Y(n538) );
  INVX0_HVT U173 ( .A(n338), .Y(n250) );
  MUX21X1_HVT U175 ( .A1(n538), .A2(n348), .S0(n284), .Y(n537) );
  MUX21X2_HVT U176 ( .A1(n241), .A2(n300), .S0(n285), .Y(n596) );
  MUX41X1_HVT U178 ( .A1(n443), .A3(n442), .A2(n444), .A4(n441), .S0(n274), 
        .S1(n331), .Y(n440) );
  MUX41X1_HVT U181 ( .A1(n468), .A3(n462), .A2(n470), .A4(n466), .S0(n346), 
        .S1(n253), .Y(n461) );
  IBUFFX16_HVT U184 ( .A(n294), .Y(n253) );
  INVX0_HVT U186 ( .A(n339), .Y(n269) );
  MUX21X2_HVT U187 ( .A1(n303), .A2(n348), .S0(n353), .Y(n469) );
  IBUFFX16_HVT U188 ( .A(n297), .Y(n254) );
  INVX2_HVT U190 ( .A(n620), .Y(n301) );
  INVX0_HVT U193 ( .A(n346), .Y(n262) );
  MUX21X2_HVT U195 ( .A1(n536), .A2(n537), .S0(n334), .Y(n535) );
  INVX1_HVT U196 ( .A(n595), .Y(n391) );
  XOR2X2_HVT U197 ( .A1(n275), .A2(n340), .Y(n322) );
  AOI21X2_HVT U199 ( .A1(n361), .A2(n1), .A3(n596), .Y(n573) );
  IBUFFX2_HVT U201 ( .A(in[4]), .Y(n364) );
  NBUFFX4_HVT U202 ( .A(n417), .Y(n341) );
  IBUFFX16_HVT U203 ( .A(n365), .Y(n278) );
  INVX1_HVT U205 ( .A(n258), .Y(n569) );
  MUX21X2_HVT U206 ( .A1(n574), .A2(n573), .S0(n335), .Y(n572) );
  NAND2X0_HVT U208 ( .A1(n621), .A2(n255), .Y(n256) );
  NAND2X0_HVT U209 ( .A1(n388), .A2(n273), .Y(n257) );
  INVX1_HVT U210 ( .A(n273), .Y(n255) );
  AND2X1_HVT U211 ( .A1(n256), .A2(n257), .Y(n260) );
  IBUFFX2_HVT U212 ( .A(n336), .Y(n273) );
  MUX41X1_HVT U213 ( .A1(n435), .A3(n436), .A2(n439), .A4(n438), .S0(n261), 
        .S1(n344), .Y(n434) );
  IBUFFX16_HVT U214 ( .A(n333), .Y(n261) );
  MUX41X1_HVT U215 ( .A1(n550), .A3(n554), .A2(n553), .A4(n556), .S0(n262), 
        .S1(n263), .Y(n549) );
  IBUFFX16_HVT U216 ( .A(n294), .Y(n263) );
  INVX1_HVT U217 ( .A(n599), .Y(n388) );
  OA21X1_HVT U218 ( .A1(n369), .A2(n364), .A3(n378), .Y(n478) );
  INVX1_HVT U219 ( .A(n268), .Y(n574) );
  INVX0_HVT U220 ( .A(in[0]), .Y(n264) );
  INVX0_HVT U221 ( .A(in[0]), .Y(n357) );
  INVX0_HVT U222 ( .A(n342), .Y(n265) );
  INVX1_HVT U223 ( .A(in[3]), .Y(n417) );
  IBUFFX2_HVT U224 ( .A(n357), .Y(n355) );
  INVX0_HVT U225 ( .A(n376), .Y(n267) );
  MUX21X1_HVT U226 ( .A1(n609), .A2(n597), .S0(n269), .Y(n268) );
  IBUFFX2_HVT U227 ( .A(n609), .Y(n382) );
  IBUFFX2_HVT U228 ( .A(n597), .Y(n390) );
  NAND2X0_HVT U229 ( .A1(n350), .A2(n270), .Y(n271) );
  NAND2X0_HVT U230 ( .A1(n608), .A2(n280), .Y(n272) );
  NAND2X0_HVT U231 ( .A1(n271), .A2(n272), .Y(n304) );
  INVX0_HVT U232 ( .A(n280), .Y(n270) );
  MUX21X1_HVT U233 ( .A1(n622), .A2(n304), .S0(n305), .Y(n563) );
  IBUFFX2_HVT U234 ( .A(n357), .Y(n353) );
  IBUFFX16_HVT U235 ( .A(n344), .Y(n274) );
  MUX21X1_HVT U236 ( .A1(n343), .A2(n416), .S0(n354), .Y(n598) );
  INVX1_HVT U237 ( .A(n276), .Y(n313) );
  INVX0_HVT U238 ( .A(n280), .Y(n281) );
  MUX21X1_HVT U239 ( .A1(n598), .A2(n601), .S0(n337), .Y(n465) );
  INVX0_HVT U240 ( .A(n315), .Y(n277) );
  INVX1_HVT U241 ( .A(n598), .Y(n389) );
  MUX21X1_HVT U242 ( .A1(n599), .A2(n329), .S0(n338), .Y(n479) );
  INVX0_HVT U243 ( .A(n333), .Y(n290) );
  NBUFFX2_HVT U244 ( .A(in[2]), .Y(n359) );
  INVX0_HVT U245 ( .A(n582), .Y(n374) );
  MUX21X1_HVT U246 ( .A1(n350), .A2(n342), .S0(n312), .Y(n314) );
  INVX0_HVT U247 ( .A(n357), .Y(n356) );
  INVX0_HVT U248 ( .A(n294), .Y(n345) );
  INVX0_HVT U249 ( .A(in[7]), .Y(n297) );
  INVX1_HVT U250 ( .A(in[6]), .Y(n275) );
  OR2X1_HVT U251 ( .A1(n341), .A2(n275), .Y(n623) );
  MUX21X1_HVT U252 ( .A1(n277), .A2(n340), .S0(n264), .Y(n276) );
  IBUFFX2_HVT U253 ( .A(n357), .Y(n312) );
  IBUFFX2_HVT U254 ( .A(n365), .Y(n279) );
  INVX1_HVT U255 ( .A(n357), .Y(n284) );
  INVX1_HVT U256 ( .A(n284), .Y(n280) );
  INVX0_HVT U257 ( .A(n314), .Y(n601) );
  IBUFFX2_HVT U258 ( .A(n357), .Y(n285) );
  INVX1_HVT U259 ( .A(n318), .Y(n306) );
  NAND2X0_HVT U260 ( .A1(n461), .A2(in[7]), .Y(n282) );
  NAND2X0_HVT U261 ( .A1(n454), .A2(n297), .Y(n283) );
  NAND2X0_HVT U262 ( .A1(n282), .A2(n283), .Y(out[6]) );
  MUX21X2_HVT U263 ( .A1(n483), .A2(n484), .S0(n290), .Y(n482) );
  INVX1_HVT U264 ( .A(n623), .Y(n419) );
  INVX1_HVT U265 ( .A(n431), .Y(n404) );
  IBUFFX2_HVT U266 ( .A(n622), .Y(n371) );
  NAND2X0_HVT U267 ( .A1(n464), .A2(n290), .Y(n286) );
  NAND2X0_HVT U268 ( .A1(n465), .A2(n333), .Y(n287) );
  NAND2X0_HVT U269 ( .A1(n286), .A2(n287), .Y(n462) );
  INVX1_HVT U270 ( .A(n373), .Y(n288) );
  MUX21X1_HVT U271 ( .A1(n473), .A2(n474), .S0(n336), .Y(n470) );
  MUX21X1_HVT U272 ( .A1(n581), .A2(n404), .S0(n338), .Y(n474) );
  INVX0_HVT U273 ( .A(n289), .Y(n581) );
  MUX21X1_HVT U274 ( .A1(n318), .A2(n347), .S0(n280), .Y(n599) );
  MUX41X1_HVT U275 ( .A1(n607), .A3(n319), .A2(n606), .A4(n391), .S0(n305), 
        .S1(n364), .Y(n548) );
  NAND2X0_HVT U276 ( .A1(n285), .A2(n348), .Y(n618) );
  INVX1_HVT U277 ( .A(n291), .Y(n545) );
  MUX41X1_HVT U278 ( .A1(n238), .A3(n382), .A2(n296), .A4(n381), .S0(n290), 
        .S1(n364), .Y(n558) );
  INVX0_HVT U279 ( .A(n546), .Y(n292) );
  MUX41X1_HVT U280 ( .A1(n292), .A3(n276), .A2(n594), .A4(n293), .S0(n290), 
        .S1(n364), .Y(n291) );
  NAND2X0_HVT U281 ( .A1(n288), .A2(n623), .Y(n293) );
  MUX41X1_HVT U282 ( .A1(n544), .A3(n545), .A2(n547), .A4(n548), .S0(in[1]), 
        .S1(in[5]), .Y(n543) );
  MUX41X1_HVT U283 ( .A1(n572), .A3(n569), .A2(n570), .A4(n565), .S0(n346), 
        .S1(n294), .Y(n564) );
  INVX0_HVT U284 ( .A(n323), .Y(n460) );
  INVX1_HVT U285 ( .A(n321), .Y(n458) );
  INVX0_HVT U286 ( .A(n304), .Y(n602) );
  INVX1_HVT U287 ( .A(n360), .Y(n305) );
  INVX1_HVT U288 ( .A(in[5]), .Y(n346) );
  INVX1_HVT U289 ( .A(n343), .Y(n308) );
  INVX1_HVT U290 ( .A(n294), .Y(n344) );
  MUX21X1_HVT U291 ( .A1(n299), .A2(n241), .S0(n285), .Y(n580) );
  IBUFFX2_HVT U292 ( .A(in[0]), .Y(n358) );
  MUX41X1_HVT U293 ( .A1(n586), .A3(n385), .A2(n386), .A4(n384), .S0(n305), 
        .S1(n364), .Y(n561) );
  MUX21X2_HVT U294 ( .A1(n557), .A2(n564), .S0(in[7]), .Y(out[0]) );
  INVX1_HVT U295 ( .A(in[4]), .Y(n365) );
  AO21X2_HVT U296 ( .A1(n358), .A2(n238), .A3(n365), .Y(n471) );
  AO21X2_HVT U297 ( .A1(n312), .A2(n416), .A3(n365), .Y(n437) );
  MUX41X1_HVT U298 ( .A1(n388), .A3(n413), .A2(n585), .A4(n490), .S0(n305), 
        .S1(n364), .Y(n489) );
  MUX21X2_HVT U299 ( .A1(n485), .A2(n475), .S0(n297), .Y(out[5]) );
  INVX0_HVT U300 ( .A(n301), .Y(n298) );
  INVX1_HVT U301 ( .A(n301), .Y(n302) );
  INVX1_HVT U302 ( .A(n301), .Y(n303) );
  INVX1_HVT U303 ( .A(n433), .Y(n402) );
  INVX1_HVT U304 ( .A(n350), .Y(n416) );
  INVX0_HVT U305 ( .A(n307), .Y(n310) );
  INVX1_HVT U306 ( .A(n309), .Y(n442) );
  NBUFFX2_HVT U307 ( .A(n275), .Y(n318) );
  MUX21X1_HVT U308 ( .A1(n308), .A2(n350), .S0(n264), .Y(n307) );
  MUX21X1_HVT U309 ( .A1(n311), .A2(n310), .S0(n320), .Y(n309) );
  NBUFFX2_HVT U310 ( .A(n275), .Y(n343) );
  INVX1_HVT U311 ( .A(n603), .Y(n387) );
  MUX21X1_HVT U312 ( .A1(n315), .A2(n341), .S0(n354), .Y(n603) );
  NAND2X0_HVT U313 ( .A1(n450), .A2(n294), .Y(n316) );
  NAND2X0_HVT U314 ( .A1(n452), .A2(n345), .Y(n317) );
  NAND2X0_HVT U315 ( .A1(n316), .A2(n317), .Y(n449) );
  MUX41X1_HVT U316 ( .A1(n588), .A3(n350), .A2(n242), .A4(n238), .S0(n305), 
        .S1(n320), .Y(n456) );
  MUX41X1_HVT U317 ( .A1(n580), .A3(n453), .A2(n241), .A4(n328), .S0(n320), 
        .S1(n305), .Y(n452) );
  MUX21X1_HVT U318 ( .A1(n308), .A2(n237), .S0(n358), .Y(n321) );
  INVX0_HVT U319 ( .A(n580), .Y(n398) );
  MUX21X1_HVT U320 ( .A1(n348), .A2(n236), .S0(n280), .Y(n323) );
  INVX1_HVT U321 ( .A(n237), .Y(n418) );
  NBUFFX2_HVT U322 ( .A(n624), .Y(n350) );
  NBUFFX2_HVT U323 ( .A(n624), .Y(n351) );
  AND2X1_HVT U324 ( .A1(n619), .A2(n351), .Y(n324) );
  NBUFFX2_HVT U325 ( .A(n624), .Y(n352) );
  MUX21X1_HVT U326 ( .A1(n399), .A2(n327), .S0(n337), .Y(n436) );
  AND2X1_HVT U327 ( .A1(n351), .A2(n609), .Y(n325) );
  MUX21X1_HVT U328 ( .A1(n241), .A2(n347), .S0(n281), .Y(n428) );
  NAND2X0_HVT U329 ( .A1(n340), .A2(n275), .Y(n624) );
  MUX21X1_HVT U330 ( .A1(n416), .A2(n420), .S0(n281), .Y(n591) );
  MUX21X1_HVT U331 ( .A1(n318), .A2(n300), .S0(n356), .Y(n481) );
  MUX21X1_HVT U332 ( .A1(n420), .A2(n342), .S0(n281), .Y(n585) );
  MUX21X1_HVT U333 ( .A1(n342), .A2(n416), .S0(n353), .Y(n594) );
  XOR2X1_HVT U334 ( .A1(n237), .A2(n355), .Y(n587) );
  MUX21X1_HVT U335 ( .A1(n420), .A2(n318), .S0(n285), .Y(n423) );
  MUX21X1_HVT U336 ( .A1(n343), .A2(n352), .S0(n284), .Y(n524) );
  MUX21X1_HVT U337 ( .A1(n419), .A2(n341), .S0(n355), .Y(n431) );
  MUX21X1_HVT U338 ( .A1(n413), .A2(n326), .S0(n335), .Y(n505) );
  XOR2X1_HVT U339 ( .A1(n347), .A2(n355), .Y(n578) );
  XNOR2X1_HVT U340 ( .A1(n350), .A2(n353), .Y(n326) );
  MUX21X1_HVT U341 ( .A1(n347), .A2(n299), .S0(n354), .Y(n590) );
  MUX21X1_HVT U342 ( .A1(n343), .A2(n347), .S0(n355), .Y(n584) );
  MUX21X1_HVT U343 ( .A1(n236), .A2(n352), .S0(n284), .Y(n610) );
  MUX21X1_HVT U344 ( .A1(n349), .A2(n351), .S0(n356), .Y(n606) );
  MUX21X1_HVT U345 ( .A1(n591), .A2(n325), .S0(n336), .Y(n502) );
  MUX21X1_HVT U346 ( .A1(n377), .A2(n315), .S0(n339), .Y(n536) );
  MUX21X1_HVT U347 ( .A1(n341), .A2(n351), .S0(n356), .Y(n430) );
  XOR2X1_HVT U348 ( .A1(n623), .A2(n356), .Y(n577) );
  MUX21X1_HVT U349 ( .A1(n348), .A2(n342), .S0(n356), .Y(n605) );
  MUX21X1_HVT U350 ( .A1(n342), .A2(n343), .S0(n285), .Y(n579) );
  AND2X1_HVT U351 ( .A1(n353), .A2(n343), .Y(n327) );
  MUX21X1_HVT U352 ( .A1(n340), .A2(n348), .S0(n284), .Y(n425) );
  MUX21X1_HVT U353 ( .A1(n349), .A2(n343), .S0(n285), .Y(n508) );
  NBUFFX2_HVT U354 ( .A(n361), .Y(n338) );
  NBUFFX2_HVT U355 ( .A(n361), .Y(n337) );
  NBUFFX2_HVT U356 ( .A(n361), .Y(n339) );
  MUX21X1_HVT U357 ( .A1(n445), .A2(n405), .S0(n337), .Y(n444) );
  MUX21X1_HVT U358 ( .A1(n350), .A2(n302), .S0(n353), .Y(n487) );
  AND2X1_HVT U359 ( .A1(n419), .A2(n358), .Y(n328) );
  MUX21X1_HVT U360 ( .A1(n507), .A2(n509), .S0(n344), .Y(n506) );
  MUX21X1_HVT U361 ( .A1(n404), .A2(n367), .S0(n339), .Y(n552) );
  AND2X1_HVT U362 ( .A1(n349), .A2(n358), .Y(n329) );
  NBUFFX2_HVT U363 ( .A(n623), .Y(n348) );
  NBUFFX2_HVT U364 ( .A(n623), .Y(n349) );
  NBUFFX2_HVT U365 ( .A(n417), .Y(n342) );
  NBUFFX2_HVT U366 ( .A(n360), .Y(n335) );
  NBUFFX2_HVT U367 ( .A(n360), .Y(n336) );
  NBUFFX2_HVT U368 ( .A(n360), .Y(n332) );
  XNOR2X1_HVT U369 ( .A1(n365), .A2(n332), .Y(n330) );
  NBUFFX2_HVT U370 ( .A(n360), .Y(n334) );
  NBUFFX2_HVT U371 ( .A(n359), .Y(n331) );
  NBUFFX2_HVT U372 ( .A(n360), .Y(n333) );
  MUX21X1_HVT U373 ( .A1(n242), .A2(n296), .S0(n285), .Y(n421) );
  MUX21X1_HVT U374 ( .A1(n303), .A2(n296), .S0(n353), .Y(n532) );
  MUX21X1_HVT U375 ( .A1(n236), .A2(n296), .S0(n355), .Y(n472) );
  MUX21X1_HVT U376 ( .A1(n497), .A2(n498), .S0(n345), .Y(n496) );
  MUX21X1_HVT U377 ( .A1(n493), .A2(n494), .S0(n344), .Y(n492) );
  MUX21X1_HVT U378 ( .A1(n419), .A2(n299), .S0(n356), .Y(n513) );
  MUX21X1_HVT U379 ( .A1(n318), .A2(n296), .S0(n353), .Y(n597) );
  MUX21X1_HVT U380 ( .A1(n296), .A2(n238), .S0(n281), .Y(n427) );
  MUX21X1_HVT U381 ( .A1(n296), .A2(n302), .S0(n354), .Y(n426) );
  NBUFFX2_HVT U382 ( .A(in[2]), .Y(n360) );
  MUX21X1_HVT U383 ( .A1(n340), .A2(n306), .S0(n285), .Y(n424) );
  MUX21X1_HVT U384 ( .A1(n348), .A2(n306), .S0(n355), .Y(n429) );
  MUX21X1_HVT U385 ( .A1(n306), .A2(n349), .S0(n284), .Y(n432) );
  MUX21X1_HVT U386 ( .A1(n306), .A2(n299), .S0(n356), .Y(n433) );
  MUX21X1_HVT U387 ( .A1(n416), .A2(n306), .S0(n354), .Y(n495) );
  XOR2X1_HVT U388 ( .A1(n354), .A2(n306), .Y(n575) );
  MUX21X1_HVT U389 ( .A1(n302), .A2(n306), .S0(n354), .Y(n595) );
  MUX21X1_HVT U390 ( .A1(n306), .A2(n237), .S0(n354), .Y(n607) );
  INVX0_HVT U391 ( .A(n613), .Y(n366) );
  INVX0_HVT U392 ( .A(n592), .Y(n367) );
  INVX0_HVT U393 ( .A(n586), .Y(n368) );
  INVX0_HVT U394 ( .A(n529), .Y(n369) );
  INVX0_HVT U395 ( .A(n490), .Y(n370) );
  INVX0_HVT U396 ( .A(n621), .Y(n372) );
  INVX0_HVT U397 ( .A(n619), .Y(n373) );
  INVX0_HVT U398 ( .A(n618), .Y(n375) );
  INVX0_HVT U399 ( .A(n617), .Y(n376) );
  INVX0_HVT U400 ( .A(n589), .Y(n377) );
  INVX0_HVT U401 ( .A(n611), .Y(n378) );
  INVX0_HVT U402 ( .A(n616), .Y(n379) );
  INVX0_HVT U403 ( .A(n612), .Y(n380) );
  INVX0_HVT U404 ( .A(n610), .Y(n381) );
  INVX0_HVT U405 ( .A(n607), .Y(n383) );
  INVX0_HVT U406 ( .A(n606), .Y(n384) );
  INVX0_HVT U407 ( .A(n605), .Y(n385) );
  INVX0_HVT U408 ( .A(n604), .Y(n386) );
  INVX0_HVT U409 ( .A(n591), .Y(n392) );
  INVX0_HVT U410 ( .A(n590), .Y(n393) );
  INVX0_HVT U411 ( .A(n588), .Y(n394) );
  INVX0_HVT U412 ( .A(n587), .Y(n395) );
  INVX0_HVT U413 ( .A(n585), .Y(n396) );
  INVX0_HVT U414 ( .A(n584), .Y(n397) );
  INVX0_HVT U415 ( .A(n579), .Y(n399) );
  INVX0_HVT U416 ( .A(n578), .Y(n400) );
  INVX0_HVT U417 ( .A(n615), .Y(n401) );
  INVX0_HVT U418 ( .A(n432), .Y(n403) );
  INVX0_HVT U419 ( .A(n430), .Y(n405) );
  INVX0_HVT U420 ( .A(n429), .Y(n406) );
  INVX0_HVT U421 ( .A(n428), .Y(n407) );
  INVX0_HVT U422 ( .A(n427), .Y(n408) );
  INVX0_HVT U423 ( .A(n426), .Y(n409) );
  INVX0_HVT U424 ( .A(n425), .Y(n410) );
  INVX0_HVT U425 ( .A(n424), .Y(n411) );
  INVX0_HVT U426 ( .A(n472), .Y(n412) );
  INVX0_HVT U427 ( .A(n423), .Y(n413) );
  INVX0_HVT U428 ( .A(n421), .Y(n415) );
endmodule

