
module inv_round ( in, last, keyin, out );
  input [127:0] in;
  input [127:0] keyin;
  output [127:0] out;
  input last;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88;
  wire   [127:0] sr_out;
  wire   [127:0] sb_out;
  wire   [127:0] oout;
  wire   [127:0] mc_out;

  AO22X1_HVT U2 ( .A1(oout[9]), .A2(n65), .A3(mc_out[9]), .A4(n78), .Y(out[9])
         );
  AO22X1_HVT U3 ( .A1(n47), .A2(n66), .A3(mc_out[99]), .A4(n78), .Y(out[99])
         );
  AO22X1_HVT U4 ( .A1(oout[98]), .A2(n66), .A3(mc_out[98]), .A4(n78), .Y(
        out[98]) );
  AO22X1_HVT U5 ( .A1(oout[97]), .A2(n66), .A3(mc_out[97]), .A4(n78), .Y(
        out[97]) );
  AO22X1_HVT U6 ( .A1(n59), .A2(n67), .A3(mc_out[96]), .A4(n78), .Y(out[96])
         );
  AO22X1_HVT U7 ( .A1(n13), .A2(n67), .A3(mc_out[95]), .A4(n78), .Y(out[95])
         );
  AO22X1_HVT U8 ( .A1(n17), .A2(n67), .A3(mc_out[94]), .A4(n78), .Y(out[94])
         );
  AO22X1_HVT U9 ( .A1(oout[93]), .A2(n67), .A3(mc_out[93]), .A4(n78), .Y(
        out[93]) );
  AO22X1_HVT U10 ( .A1(oout[92]), .A2(n67), .A3(mc_out[92]), .A4(n78), .Y(
        out[92]) );
  AO22X1_HVT U11 ( .A1(n21), .A2(n67), .A3(mc_out[91]), .A4(n78), .Y(out[91])
         );
  AO22X1_HVT U12 ( .A1(n19), .A2(n67), .A3(mc_out[90]), .A4(n78), .Y(out[90])
         );
  AO22X1_HVT U13 ( .A1(n18), .A2(n67), .A3(mc_out[8]), .A4(n78), .Y(out[8]) );
  AO22X1_HVT U14 ( .A1(oout[89]), .A2(n67), .A3(mc_out[89]), .A4(n79), .Y(
        out[89]) );
  AO22X1_HVT U15 ( .A1(oout[88]), .A2(n67), .A3(mc_out[88]), .A4(n79), .Y(
        out[88]) );
  AO22X1_HVT U16 ( .A1(oout[87]), .A2(n67), .A3(mc_out[87]), .A4(n79), .Y(
        out[87]) );
  AO22X1_HVT U17 ( .A1(n12), .A2(n67), .A3(mc_out[86]), .A4(n79), .Y(out[86])
         );
  AO22X1_HVT U18 ( .A1(n15), .A2(n67), .A3(mc_out[85]), .A4(n79), .Y(out[85])
         );
  AO22X1_HVT U19 ( .A1(oout[84]), .A2(n67), .A3(mc_out[84]), .A4(n79), .Y(
        out[84]) );
  AO22X1_HVT U20 ( .A1(oout[83]), .A2(n67), .A3(mc_out[83]), .A4(n79), .Y(
        out[83]) );
  AO22X1_HVT U21 ( .A1(oout[82]), .A2(n68), .A3(mc_out[82]), .A4(n79), .Y(
        out[82]) );
  AO22X1_HVT U22 ( .A1(oout[81]), .A2(n68), .A3(mc_out[81]), .A4(n79), .Y(
        out[81]) );
  AO22X1_HVT U23 ( .A1(n68), .A2(n11), .A3(mc_out[80]), .A4(n79), .Y(out[80])
         );
  AO22X1_HVT U24 ( .A1(n54), .A2(n68), .A3(mc_out[7]), .A4(n79), .Y(out[7]) );
  AO22X1_HVT U25 ( .A1(n5), .A2(n68), .A3(mc_out[79]), .A4(n79), .Y(out[79])
         );
  AO22X1_HVT U26 ( .A1(oout[78]), .A2(n68), .A3(mc_out[78]), .A4(n80), .Y(
        out[78]) );
  AO22X1_HVT U27 ( .A1(oout[77]), .A2(n68), .A3(mc_out[77]), .A4(n80), .Y(
        out[77]) );
  AO22X1_HVT U28 ( .A1(oout[76]), .A2(n68), .A3(mc_out[76]), .A4(n80), .Y(
        out[76]) );
  AO22X1_HVT U29 ( .A1(oout[75]), .A2(n68), .A3(mc_out[75]), .A4(n80), .Y(
        out[75]) );
  AO22X1_HVT U30 ( .A1(oout[74]), .A2(n68), .A3(mc_out[74]), .A4(n80), .Y(
        out[74]) );
  AO22X1_HVT U31 ( .A1(n68), .A2(n31), .A3(mc_out[73]), .A4(n80), .Y(out[73])
         );
  AO22X1_HVT U32 ( .A1(n6), .A2(n68), .A3(mc_out[72]), .A4(n80), .Y(out[72])
         );
  AO22X1_HVT U33 ( .A1(n56), .A2(n68), .A3(mc_out[71]), .A4(n80), .Y(out[71])
         );
  AO22X1_HVT U34 ( .A1(n50), .A2(n68), .A3(mc_out[70]), .A4(n80), .Y(out[70])
         );
  AO22X1_HVT U35 ( .A1(n4), .A2(n68), .A3(mc_out[6]), .A4(n80), .Y(out[6]) );
  AO22X1_HVT U36 ( .A1(oout[69]), .A2(n69), .A3(mc_out[69]), .A4(n80), .Y(
        out[69]) );
  AO22X1_HVT U37 ( .A1(oout[68]), .A2(n69), .A3(mc_out[68]), .A4(n80), .Y(
        out[68]) );
  AO22X1_HVT U38 ( .A1(oout[67]), .A2(n69), .A3(mc_out[67]), .A4(n81), .Y(
        out[67]) );
  AO22X1_HVT U39 ( .A1(n60), .A2(n69), .A3(mc_out[66]), .A4(n81), .Y(out[66])
         );
  AO22X1_HVT U40 ( .A1(n69), .A2(oout[65]), .A3(mc_out[65]), .A4(n81), .Y(
        out[65]) );
  AO22X1_HVT U41 ( .A1(oout[64]), .A2(n69), .A3(mc_out[64]), .A4(n81), .Y(
        out[64]) );
  AO22X1_HVT U42 ( .A1(n63), .A2(n69), .A3(mc_out[63]), .A4(n81), .Y(out[63])
         );
  AO22X1_HVT U43 ( .A1(n9), .A2(n69), .A3(mc_out[62]), .A4(n81), .Y(out[62])
         );
  AO22X1_HVT U44 ( .A1(n30), .A2(n69), .A3(mc_out[61]), .A4(n81), .Y(out[61])
         );
  AO22X1_HVT U45 ( .A1(oout[60]), .A2(n69), .A3(mc_out[60]), .A4(n81), .Y(
        out[60]) );
  AO22X1_HVT U46 ( .A1(oout[5]), .A2(n69), .A3(mc_out[5]), .A4(n81), .Y(out[5]) );
  AO22X1_HVT U47 ( .A1(n10), .A2(n69), .A3(mc_out[59]), .A4(n81), .Y(out[59])
         );
  AO22X1_HVT U48 ( .A1(n53), .A2(n69), .A3(mc_out[58]), .A4(n81), .Y(out[58])
         );
  AO22X1_HVT U49 ( .A1(n33), .A2(n69), .A3(mc_out[57]), .A4(n81), .Y(out[57])
         );
  AO22X1_HVT U50 ( .A1(n38), .A2(n69), .A3(n82), .A4(mc_out[56]), .Y(out[56])
         );
  AO22X1_HVT U51 ( .A1(oout[55]), .A2(n70), .A3(mc_out[55]), .A4(n82), .Y(
        out[55]) );
  AO22X1_HVT U52 ( .A1(n35), .A2(n70), .A3(mc_out[54]), .A4(n82), .Y(out[54])
         );
  AO22X1_HVT U53 ( .A1(n62), .A2(n70), .A3(mc_out[53]), .A4(n82), .Y(out[53])
         );
  AO22X1_HVT U54 ( .A1(n70), .A2(oout[52]), .A3(mc_out[52]), .A4(n82), .Y(
        out[52]) );
  AO22X1_HVT U55 ( .A1(n61), .A2(n70), .A3(mc_out[51]), .A4(n82), .Y(out[51])
         );
  AO22X1_HVT U56 ( .A1(oout[50]), .A2(n70), .A3(mc_out[50]), .A4(n82), .Y(
        out[50]) );
  AO22X1_HVT U57 ( .A1(oout[4]), .A2(n70), .A3(mc_out[4]), .A4(n82), .Y(out[4]) );
  AO22X1_HVT U58 ( .A1(oout[49]), .A2(n70), .A3(mc_out[49]), .A4(n82), .Y(
        out[49]) );
  AO22X1_HVT U59 ( .A1(oout[48]), .A2(n70), .A3(mc_out[48]), .A4(n82), .Y(
        out[48]) );
  AO22X1_HVT U60 ( .A1(n52), .A2(n70), .A3(mc_out[47]), .A4(n82), .Y(out[47])
         );
  AO22X1_HVT U61 ( .A1(oout[46]), .A2(n70), .A3(mc_out[46]), .A4(n82), .Y(
        out[46]) );
  AO22X1_HVT U62 ( .A1(oout[45]), .A2(n70), .A3(mc_out[45]), .A4(n83), .Y(
        out[45]) );
  AO22X1_HVT U63 ( .A1(oout[44]), .A2(n70), .A3(mc_out[44]), .A4(n83), .Y(
        out[44]) );
  AO22X1_HVT U64 ( .A1(oout[43]), .A2(n70), .A3(mc_out[43]), .A4(n83), .Y(
        out[43]) );
  AO22X1_HVT U65 ( .A1(oout[42]), .A2(n70), .A3(mc_out[42]), .A4(n83), .Y(
        out[42]) );
  AO22X1_HVT U66 ( .A1(n71), .A2(oout[41]), .A3(mc_out[41]), .A4(n83), .Y(
        out[41]) );
  AO22X1_HVT U67 ( .A1(n71), .A2(oout[40]), .A3(mc_out[40]), .A4(n83), .Y(
        out[40]) );
  AO22X1_HVT U68 ( .A1(n40), .A2(n71), .A3(mc_out[3]), .A4(n83), .Y(out[3]) );
  AO22X1_HVT U69 ( .A1(oout[39]), .A2(n71), .A3(mc_out[39]), .A4(n83), .Y(
        out[39]) );
  AO22X1_HVT U70 ( .A1(oout[38]), .A2(n71), .A3(n83), .A4(mc_out[38]), .Y(
        out[38]) );
  AO22X1_HVT U71 ( .A1(oout[37]), .A2(n71), .A3(mc_out[37]), .A4(n83), .Y(
        out[37]) );
  AO22X1_HVT U72 ( .A1(oout[36]), .A2(n71), .A3(mc_out[36]), .A4(n83), .Y(
        out[36]) );
  AO22X1_HVT U73 ( .A1(oout[35]), .A2(n71), .A3(mc_out[35]), .A4(n83), .Y(
        out[35]) );
  AO22X1_HVT U74 ( .A1(n16), .A2(n71), .A3(mc_out[34]), .A4(n84), .Y(out[34])
         );
  AO22X1_HVT U75 ( .A1(oout[33]), .A2(n71), .A3(mc_out[33]), .A4(n84), .Y(
        out[33]) );
  AO22X1_HVT U76 ( .A1(n24), .A2(n71), .A3(mc_out[32]), .A4(n84), .Y(out[32])
         );
  AO22X1_HVT U77 ( .A1(n20), .A2(n71), .A3(mc_out[31]), .A4(n84), .Y(out[31])
         );
  AO22X1_HVT U78 ( .A1(n71), .A2(n29), .A3(mc_out[30]), .A4(n84), .Y(out[30])
         );
  AO22X1_HVT U79 ( .A1(n49), .A2(n71), .A3(mc_out[2]), .A4(n84), .Y(out[2]) );
  AO22X1_HVT U80 ( .A1(oout[29]), .A2(n71), .A3(mc_out[29]), .A4(n84), .Y(
        out[29]) );
  AO22X1_HVT U81 ( .A1(oout[28]), .A2(n72), .A3(mc_out[28]), .A4(n84), .Y(
        out[28]) );
  AO22X1_HVT U82 ( .A1(n23), .A2(n72), .A3(mc_out[27]), .A4(n84), .Y(out[27])
         );
  AO22X1_HVT U83 ( .A1(n72), .A2(n26), .A3(mc_out[26]), .A4(n84), .Y(out[26])
         );
  AO22X1_HVT U84 ( .A1(n41), .A2(n72), .A3(mc_out[25]), .A4(n84), .Y(out[25])
         );
  AO22X1_HVT U85 ( .A1(n1), .A2(n72), .A3(mc_out[24]), .A4(n84), .Y(out[24])
         );
  AO22X1_HVT U86 ( .A1(n72), .A2(n7), .A3(mc_out[23]), .A4(n85), .Y(out[23])
         );
  AO22X1_HVT U87 ( .A1(n28), .A2(n72), .A3(mc_out[22]), .A4(n85), .Y(out[22])
         );
  AO22X1_HVT U88 ( .A1(oout[21]), .A2(n72), .A3(mc_out[21]), .A4(n85), .Y(
        out[21]) );
  AO22X1_HVT U89 ( .A1(oout[20]), .A2(n72), .A3(mc_out[20]), .A4(n85), .Y(
        out[20]) );
  AO22X1_HVT U90 ( .A1(oout[1]), .A2(n72), .A3(mc_out[1]), .A4(n85), .Y(out[1]) );
  AO22X1_HVT U91 ( .A1(n43), .A2(n72), .A3(mc_out[19]), .A4(n85), .Y(out[19])
         );
  AO22X1_HVT U92 ( .A1(n51), .A2(n72), .A3(mc_out[18]), .A4(n85), .Y(out[18])
         );
  AO22X1_HVT U93 ( .A1(n42), .A2(n72), .A3(mc_out[17]), .A4(n85), .Y(out[17])
         );
  AO22X1_HVT U94 ( .A1(oout[16]), .A2(n72), .A3(mc_out[16]), .A4(n85), .Y(
        out[16]) );
  AO22X1_HVT U95 ( .A1(oout[15]), .A2(n72), .A3(mc_out[15]), .A4(n85), .Y(
        out[15]) );
  AO22X1_HVT U96 ( .A1(n8), .A2(n73), .A3(mc_out[14]), .A4(n85), .Y(out[14])
         );
  AO22X1_HVT U97 ( .A1(oout[13]), .A2(n73), .A3(mc_out[13]), .A4(n85), .Y(
        out[13]) );
  AO22X1_HVT U98 ( .A1(oout[12]), .A2(n73), .A3(mc_out[12]), .A4(n86), .Y(
        out[12]) );
  AO22X1_HVT U99 ( .A1(n45), .A2(n73), .A3(mc_out[127]), .A4(n86), .Y(out[127]) );
  AO22X1_HVT U100 ( .A1(n55), .A2(n73), .A3(mc_out[126]), .A4(n86), .Y(
        out[126]) );
  AO22X1_HVT U101 ( .A1(n48), .A2(n73), .A3(mc_out[125]), .A4(n86), .Y(
        out[125]) );
  AO22X1_HVT U102 ( .A1(oout[124]), .A2(n73), .A3(mc_out[124]), .A4(n86), .Y(
        out[124]) );
  AO22X1_HVT U103 ( .A1(oout[123]), .A2(n73), .A3(mc_out[123]), .A4(n86), .Y(
        out[123]) );
  AO22X1_HVT U104 ( .A1(oout[122]), .A2(n73), .A3(mc_out[122]), .A4(n86), .Y(
        out[122]) );
  AO22X1_HVT U105 ( .A1(n73), .A2(n34), .A3(mc_out[121]), .A4(n86), .Y(
        out[121]) );
  AO22X1_HVT U106 ( .A1(oout[120]), .A2(n73), .A3(mc_out[120]), .A4(n86), .Y(
        out[120]) );
  AO22X1_HVT U107 ( .A1(oout[11]), .A2(n73), .A3(mc_out[11]), .A4(n86), .Y(
        out[11]) );
  AO22X1_HVT U108 ( .A1(n46), .A2(n73), .A3(mc_out[119]), .A4(n86), .Y(
        out[119]) );
  AO22X1_HVT U109 ( .A1(oout[118]), .A2(n73), .A3(mc_out[118]), .A4(n86), .Y(
        out[118]) );
  AO22X1_HVT U110 ( .A1(n3), .A2(n73), .A3(mc_out[117]), .A4(n87), .Y(out[117]) );
  AO22X1_HVT U111 ( .A1(oout[116]), .A2(n74), .A3(mc_out[116]), .A4(n87), .Y(
        out[116]) );
  AO22X1_HVT U112 ( .A1(n44), .A2(n74), .A3(mc_out[115]), .A4(n87), .Y(
        out[115]) );
  AO22X1_HVT U113 ( .A1(oout[114]), .A2(n74), .A3(mc_out[114]), .A4(n87), .Y(
        out[114]) );
  AO22X1_HVT U114 ( .A1(oout[113]), .A2(n74), .A3(mc_out[113]), .A4(n87), .Y(
        out[113]) );
  AO22X1_HVT U115 ( .A1(oout[112]), .A2(n74), .A3(mc_out[112]), .A4(n87), .Y(
        out[112]) );
  AO22X1_HVT U116 ( .A1(n64), .A2(n74), .A3(mc_out[111]), .A4(n87), .Y(
        out[111]) );
  AO22X1_HVT U117 ( .A1(n36), .A2(n74), .A3(mc_out[110]), .A4(n87), .Y(
        out[110]) );
  AO22X1_HVT U118 ( .A1(oout[10]), .A2(n74), .A3(mc_out[10]), .A4(n87), .Y(
        out[10]) );
  AO22X1_HVT U119 ( .A1(n37), .A2(n74), .A3(mc_out[109]), .A4(n87), .Y(
        out[109]) );
  AO22X1_HVT U120 ( .A1(oout[108]), .A2(n74), .A3(mc_out[108]), .A4(n87), .Y(
        out[108]) );
  AO22X1_HVT U121 ( .A1(n27), .A2(n74), .A3(mc_out[107]), .A4(n87), .Y(
        out[107]) );
  AO22X1_HVT U122 ( .A1(n39), .A2(n74), .A3(mc_out[106]), .A4(n88), .Y(
        out[106]) );
  AO22X1_HVT U123 ( .A1(n2), .A2(n74), .A3(mc_out[105]), .A4(n88), .Y(out[105]) );
  AO22X1_HVT U124 ( .A1(n74), .A2(n14), .A3(mc_out[104]), .A4(n88), .Y(
        out[104]) );
  AO22X1_HVT U125 ( .A1(oout[103]), .A2(n74), .A3(mc_out[103]), .A4(n88), .Y(
        out[103]) );
  AO22X1_HVT U126 ( .A1(n32), .A2(n75), .A3(mc_out[102]), .A4(n88), .Y(
        out[102]) );
  AO22X1_HVT U127 ( .A1(oout[101]), .A2(n75), .A3(mc_out[101]), .A4(n88), .Y(
        out[101]) );
  AO22X1_HVT U128 ( .A1(oout[100]), .A2(n75), .A3(mc_out[100]), .A4(n88), .Y(
        out[100]) );
  AO22X1_HVT U129 ( .A1(oout[0]), .A2(n75), .A3(mc_out[0]), .A4(n88), .Y(
        out[0]) );
  inv_shift_rows sr ( .in({in[127:80], n58, in[78:0]}), .out(sr_out) );
  inv_subbytes sb ( .in(sr_out), .out(sb_out) );
  inv_add_round_keys adk ( .state(sb_out), .subkey(keyin), .out(oout) );
  inv_Mix_Column mc ( .in(oout), .out1(mc_out) );
  DELLN2X2_HVT U1 ( .A(oout[24]), .Y(n1) );
  DELLN2X2_HVT U130 ( .A(oout[105]), .Y(n2) );
  DELLN2X2_HVT U131 ( .A(oout[117]), .Y(n3) );
  DELLN2X2_HVT U132 ( .A(oout[31]), .Y(n20) );
  DELLN2X2_HVT U133 ( .A(oout[109]), .Y(n37) );
  DELLN2X2_HVT U134 ( .A(oout[6]), .Y(n4) );
  DELLN2X2_HVT U135 ( .A(oout[79]), .Y(n5) );
  DELLN2X2_HVT U136 ( .A(oout[72]), .Y(n6) );
  DELLN2X2_HVT U137 ( .A(oout[23]), .Y(n7) );
  DELLN2X2_HVT U138 ( .A(oout[14]), .Y(n8) );
  DELLN2X2_HVT U139 ( .A(oout[62]), .Y(n9) );
  DELLN2X2_HVT U140 ( .A(oout[59]), .Y(n10) );
  NBUFFX2_HVT U141 ( .A(oout[111]), .Y(n64) );
  DELLN2X2_HVT U142 ( .A(oout[80]), .Y(n11) );
  DELLN2X2_HVT U143 ( .A(oout[86]), .Y(n12) );
  DELLN2X2_HVT U144 ( .A(oout[95]), .Y(n13) );
  NBUFFX2_HVT U145 ( .A(oout[34]), .Y(n16) );
  DELLN2X2_HVT U146 ( .A(oout[126]), .Y(n55) );
  DELLN2X2_HVT U147 ( .A(oout[104]), .Y(n14) );
  DELLN2X2_HVT U148 ( .A(oout[85]), .Y(n15) );
  DELLN2X2_HVT U149 ( .A(oout[94]), .Y(n17) );
  DELLN2X2_HVT U150 ( .A(oout[8]), .Y(n18) );
  DELLN2X2_HVT U151 ( .A(oout[47]), .Y(n52) );
  DELLN2X2_HVT U152 ( .A(oout[90]), .Y(n19) );
  DELLN2X2_HVT U153 ( .A(oout[91]), .Y(n21) );
  DELLN2X2_HVT U154 ( .A(oout[26]), .Y(n22) );
  DELLN2X2_HVT U155 ( .A(oout[27]), .Y(n23) );
  DELLN2X2_HVT U156 ( .A(oout[32]), .Y(n24) );
  IBUFFX2_HVT U157 ( .A(n22), .Y(n25) );
  INVX1_HVT U158 ( .A(n25), .Y(n26) );
  NBUFFX2_HVT U159 ( .A(oout[107]), .Y(n27) );
  DELLN2X2_HVT U160 ( .A(oout[22]), .Y(n28) );
  DELLN2X2_HVT U161 ( .A(oout[2]), .Y(n49) );
  DELLN2X2_HVT U162 ( .A(oout[30]), .Y(n29) );
  DELLN2X2_HVT U163 ( .A(oout[61]), .Y(n30) );
  DELLN2X2_HVT U164 ( .A(oout[19]), .Y(n43) );
  DELLN2X2_HVT U165 ( .A(oout[73]), .Y(n31) );
  DELLN2X2_HVT U166 ( .A(oout[125]), .Y(n48) );
  DELLN2X2_HVT U167 ( .A(oout[102]), .Y(n32) );
  DELLN2X2_HVT U168 ( .A(oout[57]), .Y(n33) );
  DELLN2X2_HVT U169 ( .A(oout[121]), .Y(n34) );
  DELLN2X2_HVT U170 ( .A(oout[54]), .Y(n35) );
  DELLN2X2_HVT U171 ( .A(oout[110]), .Y(n36) );
  DELLN1X2_HVT U172 ( .A(oout[119]), .Y(n46) );
  DELLN2X2_HVT U173 ( .A(oout[56]), .Y(n38) );
  DELLN2X2_HVT U174 ( .A(oout[106]), .Y(n39) );
  DELLN2X2_HVT U175 ( .A(oout[3]), .Y(n40) );
  DELLN2X2_HVT U176 ( .A(oout[25]), .Y(n41) );
  DELLN2X2_HVT U177 ( .A(oout[17]), .Y(n42) );
  DELLN2X2_HVT U178 ( .A(oout[115]), .Y(n44) );
  DELLN2X2_HVT U179 ( .A(oout[127]), .Y(n45) );
  INVX1_HVT U180 ( .A(n57), .Y(n58) );
  DELLN2X2_HVT U181 ( .A(oout[71]), .Y(n56) );
  DELLN2X2_HVT U182 ( .A(oout[99]), .Y(n47) );
  DELLN2X2_HVT U183 ( .A(oout[70]), .Y(n50) );
  DELLN2X2_HVT U184 ( .A(oout[18]), .Y(n51) );
  DELLN2X2_HVT U185 ( .A(oout[58]), .Y(n53) );
  DELLN2X2_HVT U186 ( .A(oout[7]), .Y(n54) );
  INVX1_HVT U187 ( .A(in[79]), .Y(n57) );
  DELLN2X2_HVT U188 ( .A(oout[96]), .Y(n59) );
  DELLN2X2_HVT U189 ( .A(oout[66]), .Y(n60) );
  DELLN2X2_HVT U190 ( .A(oout[51]), .Y(n61) );
  DELLN2X2_HVT U191 ( .A(oout[53]), .Y(n62) );
  DELLN2X2_HVT U192 ( .A(oout[63]), .Y(n63) );
  INVX0_HVT U193 ( .A(last), .Y(n76) );
  INVX1_HVT U194 ( .A(n66), .Y(n82) );
  INVX1_HVT U195 ( .A(n66), .Y(n81) );
  INVX1_HVT U196 ( .A(n66), .Y(n80) );
  INVX1_HVT U197 ( .A(n66), .Y(n78) );
  INVX1_HVT U198 ( .A(n66), .Y(n79) );
  INVX1_HVT U199 ( .A(n65), .Y(n84) );
  INVX1_HVT U200 ( .A(n65), .Y(n83) );
  INVX1_HVT U201 ( .A(n65), .Y(n85) );
  INVX1_HVT U202 ( .A(n65), .Y(n87) );
  INVX1_HVT U203 ( .A(n65), .Y(n86) );
  INVX1_HVT U204 ( .A(n65), .Y(n88) );
  INVX1_HVT U205 ( .A(n77), .Y(n68) );
  INVX1_HVT U206 ( .A(n77), .Y(n67) );
  INVX1_HVT U207 ( .A(n76), .Y(n70) );
  INVX1_HVT U208 ( .A(n76), .Y(n72) );
  INVX1_HVT U209 ( .A(n76), .Y(n71) );
  INVX1_HVT U210 ( .A(n76), .Y(n73) );
  INVX1_HVT U211 ( .A(n76), .Y(n74) );
  INVX1_HVT U212 ( .A(n77), .Y(n69) );
  INVX1_HVT U213 ( .A(n77), .Y(n66) );
  INVX1_HVT U214 ( .A(n77), .Y(n65) );
  INVX1_HVT U215 ( .A(n76), .Y(n75) );
  INVX0_HVT U216 ( .A(last), .Y(n77) );
endmodule

