
module inv_sbox_9 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n187, n196, n197, n198, n199, n200, n201, n202, n205, n208, n210,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605;

  NAND2X0_HVT U1 ( .A1(n277), .A2(n319), .Y(n605) );
  NAND2X0_HVT U5 ( .A1(n602), .A2(n327), .Y(n601) );
  NAND2X0_HVT U6 ( .A1(n335), .A2(n303), .Y(n599) );
  NAND2X0_HVT U9 ( .A1(n331), .A2(n597), .Y(n596) );
  NAND2X0_HVT U10 ( .A1(n303), .A2(n594), .Y(n595) );
  NAND2X0_HVT U11 ( .A1(n338), .A2(n278), .Y(n593) );
  NAND2X0_HVT U12 ( .A1(n259), .A2(n316), .Y(n592) );
  NAND2X0_HVT U13 ( .A1(n328), .A2(n597), .Y(n591) );
  NAND2X0_HVT U15 ( .A1(n325), .A2(n332), .Y(n589) );
  NAND2X0_HVT U19 ( .A1(n336), .A2(n238), .Y(n584) );
  NAND2X0_HVT U25 ( .A1(n281), .A2(n317), .Y(n600) );
  NAND2X0_HVT U32 ( .A1(n319), .A2(n338), .Y(n572) );
  NAND2X0_HVT U38 ( .A1(n316), .A2(n338), .Y(n566) );
  NAND2X0_HVT U42 ( .A1(n599), .A2(n399), .Y(n562) );
  OA21X1_HVT U53 ( .A1(n344), .A2(n554), .A3(n371), .Y(n552) );
  NAND2X0_HVT U55 ( .A1(n328), .A2(n602), .Y(n550) );
  MUX41X1_HVT U56 ( .A1(n383), .A3(n324), .A2(n369), .A4(n550), .S0(n308), 
        .S1(n271), .Y(n549) );
  AO21X1_HVT U60 ( .A1(n544), .A2(n312), .A3(n583), .Y(n545) );
  MUX41X1_HVT U62 ( .A1(n543), .A3(n549), .A2(n547), .A4(n551), .S0(in[5]), 
        .S1(n266), .Y(n542) );
  MUX41X1_HVT U65 ( .A1(n362), .A3(n364), .A2(n363), .A4(n566), .S0(n308), 
        .S1(n341), .Y(n539) );
  NAND2X0_HVT U66 ( .A1(n336), .A2(n222), .Y(n538) );
  MUX41X1_HVT U67 ( .A1(n359), .A3(n384), .A2(n361), .A4(n538), .S0(n314), 
        .S1(n275), .Y(n537) );
  MUX41X1_HVT U71 ( .A1(n248), .A3(n398), .A2(n593), .A4(n355), .S0(n307), 
        .S1(n247), .Y(n534) );
  NAND2X0_HVT U72 ( .A1(n325), .A2(n598), .Y(n533) );
  MUX41X1_HVT U73 ( .A1(n577), .A3(n533), .A2(n286), .A4(n315), .S0(n313), 
        .S1(n305), .Y(n532) );
  MUX41X1_HVT U74 ( .A1(n595), .A3(n375), .A2(n374), .A4(n365), .S0(n308), 
        .S1(n341), .Y(n531) );
  MUX41X1_HVT U78 ( .A1(n528), .A3(n532), .A2(n531), .A4(n534), .S0(n249), 
        .S1(n322), .Y(n527) );
  MUX41X1_HVT U80 ( .A1(n386), .A3(n383), .A2(n596), .A4(n601), .S0(n307), 
        .S1(n247), .Y(n525) );
  NAND2X0_HVT U81 ( .A1(n278), .A2(n598), .Y(n524) );
  AND2X1_HVT U82 ( .A1(n248), .A2(n328), .Y(n523) );
  MUX41X1_HVT U83 ( .A1(n523), .A3(n373), .A2(n202), .A4(n524), .S0(n307), 
        .S1(n340), .Y(n522) );
  MUX41X1_HVT U84 ( .A1(n300), .A3(n372), .A2(n387), .A4(n579), .S0(n308), 
        .S1(n340), .Y(n521) );
  MUX41X1_HVT U85 ( .A1(n521), .A3(n525), .A2(n522), .A4(n526), .S0(n249), 
        .S1(n322), .Y(n520) );
  MUX41X1_HVT U88 ( .A1(n361), .A3(n347), .A2(n574), .A4(n558), .S0(n307), 
        .S1(n271), .Y(n518) );
  NAND2X0_HVT U89 ( .A1(n338), .A2(n397), .Y(n517) );
  MUX41X1_HVT U96 ( .A1(n384), .A3(n591), .A2(n370), .A4(n388), .S0(n308), 
        .S1(n341), .Y(n510) );
  MUX41X1_HVT U99 ( .A1(n572), .A3(n363), .A2(n556), .A4(n324), .S0(n341), 
        .S1(n306), .Y(n507) );
  NAND2X0_HVT U100 ( .A1(n338), .A2(n396), .Y(n506) );
  AND2X1_HVT U104 ( .A1(n598), .A2(n326), .Y(n503) );
  MUX41X1_HVT U105 ( .A1(n590), .A3(n391), .A2(n524), .A4(n503), .S0(n308), 
        .S1(n314), .Y(n502) );
  MUX41X1_HVT U108 ( .A1(n365), .A3(n324), .A2(n369), .A4(n329), .S0(n308), 
        .S1(n271), .Y(n499) );
  MUX41X1_HVT U109 ( .A1(n389), .A3(n347), .A2(n387), .A4(n381), .S0(n307), 
        .S1(n271), .Y(n498) );
  MUX41X1_HVT U110 ( .A1(n498), .A3(n500), .A2(n499), .A4(n502), .S0(in[5]), 
        .S1(n322), .Y(n497) );
  AO21X1_HVT U112 ( .A1(n378), .A2(n313), .A3(n580), .Y(n495) );
  NAND2X0_HVT U114 ( .A1(n331), .A2(n598), .Y(n493) );
  MUX41X1_HVT U115 ( .A1(n493), .A3(n593), .A2(n378), .A4(n328), .S0(n271), 
        .S1(n305), .Y(n492) );
  MUX41X1_HVT U116 ( .A1(n377), .A3(n372), .A2(n347), .A4(n589), .S0(n306), 
        .S1(n271), .Y(n491) );
  NAND2X0_HVT U118 ( .A1(n338), .A2(n277), .Y(n489) );
  MUX41X1_HVT U119 ( .A1(n392), .A3(n490), .A2(n567), .A4(n489), .S0(n306), 
        .S1(n271), .Y(n488) );
  MUX41X1_HVT U120 ( .A1(n488), .A3(n492), .A2(n491), .A4(n494), .S0(n249), 
        .S1(n322), .Y(n487) );
  MUX41X1_HVT U122 ( .A1(n382), .A3(n296), .A2(n558), .A4(n385), .S0(n306), 
        .S1(n341), .Y(n486) );
  MUX41X1_HVT U124 ( .A1(n299), .A3(n485), .A2(n581), .A4(n295), .S0(n312), 
        .S1(n306), .Y(n484) );
  AOI21X1_HVT U127 ( .A1(n311), .A2(n480), .A3(n354), .Y(n481) );
  NAND2X0_HVT U129 ( .A1(n310), .A2(n605), .Y(n478) );
  MUX41X1_HVT U130 ( .A1(n478), .A3(n479), .A2(n482), .A4(n481), .S0(n314), 
        .S1(n322), .Y(n477) );
  AND2X1_HVT U131 ( .A1(n222), .A2(n224), .Y(n476) );
  MUX41X1_HVT U132 ( .A1(n351), .A3(n476), .A2(n394), .A4(n359), .S0(n313), 
        .S1(n305), .Y(n475) );
  MUX41X1_HVT U133 ( .A1(n395), .A3(n353), .A2(n550), .A4(n352), .S0(n312), 
        .S1(n304), .Y(n474) );
  MUX41X1_HVT U136 ( .A1(n555), .A3(n506), .A2(n472), .A4(n357), .S0(n310), 
        .S1(n340), .Y(n471) );
  MUX41X1_HVT U137 ( .A1(n597), .A3(n575), .A2(n579), .A4(n388), .S0(n314), 
        .S1(n304), .Y(n470) );
  MUX41X1_HVT U140 ( .A1(n374), .A3(n297), .A2(n368), .A4(n593), .S0(n313), 
        .S1(n275), .Y(n468) );
  NAND2X0_HVT U141 ( .A1(n325), .A2(n338), .Y(n467) );
  MUX41X1_HVT U142 ( .A1(n467), .A3(n565), .A2(n393), .A4(n368), .S0(n311), 
        .S1(n247), .Y(n466) );
  MUX41X1_HVT U145 ( .A1(n573), .A3(n391), .A2(n464), .A4(n524), .S0(n311), 
        .S1(n262), .Y(n463) );
  MUX41X1_HVT U151 ( .A1(n202), .A3(n376), .A2(n366), .A4(n458), .S0(n312), 
        .S1(n304), .Y(n457) );
  MUX41X1_HVT U155 ( .A1(n368), .A3(n593), .A2(n585), .A4(n370), .S0(n309), 
        .S1(n262), .Y(n453) );
  MUX41X1_HVT U156 ( .A1(n453), .A3(n457), .A2(n454), .A4(n459), .S0(n249), 
        .S1(n322), .Y(n452) );
  NAND2X0_HVT U159 ( .A1(n449), .A2(n448), .Y(n450) );
  MUX41X1_HVT U162 ( .A1(n289), .A3(n364), .A2(n569), .A4(n446), .S0(n309), 
        .S1(n340), .Y(n445) );
  NAND2X0_HVT U163 ( .A1(n336), .A2(n397), .Y(n444) );
  MUX41X1_HVT U164 ( .A1(n596), .A3(n444), .A2(n567), .A4(n365), .S0(n306), 
        .S1(n262), .Y(n443) );
  NAND2X0_HVT U166 ( .A1(n594), .A2(n440), .Y(n441) );
  MUX41X1_HVT U172 ( .A1(n517), .A3(n435), .A2(n298), .A4(n582), .S0(n309), 
        .S1(n262), .Y(n434) );
  MUX41X1_HVT U173 ( .A1(n331), .A3(n398), .A2(n329), .A4(n568), .S0(n309), 
        .S1(n262), .Y(n433) );
  MUX41X1_HVT U174 ( .A1(n283), .A3(n550), .A2(n395), .A4(n399), .S0(n309), 
        .S1(n262), .Y(n432) );
  NAND2X0_HVT U177 ( .A1(n332), .A2(n277), .Y(n430) );
  MUX41X1_HVT U178 ( .A1(n301), .A3(n430), .A2(n398), .A4(n560), .S0(n309), 
        .S1(n262), .Y(n429) );
  AND2X1_HVT U179 ( .A1(n248), .A2(n326), .Y(n428) );
  MUX41X1_HVT U183 ( .A1(n379), .A3(n383), .A2(n365), .A4(n562), .S0(n312), 
        .S1(n305), .Y(n424) );
  AND2X1_HVT U185 ( .A1(n399), .A2(n224), .Y(n422) );
  NAND2X0_HVT U191 ( .A1(n343), .A2(n358), .Y(n417) );
  AND2X1_HVT U192 ( .A1(n375), .A2(n415), .Y(n416) );
  NAND2X0_HVT U194 ( .A1(n562), .A2(n415), .Y(n413) );
  MUX41X1_HVT U195 ( .A1(n414), .A3(n413), .A2(n416), .A4(n417), .S0(n307), 
        .S1(n321), .Y(n412) );
  NAND2X0_HVT U198 ( .A1(n336), .A2(n399), .Y(n594) );
  NAND2X0_HVT U200 ( .A1(n327), .A2(n338), .Y(n480) );
  NAND2X0_HVT U207 ( .A1(n338), .A2(n398), .Y(n544) );
  MUX41X1_HVT U2 ( .A1(n512), .A3(n518), .A2(n516), .A4(n519), .S0(n187), .S1(
        n266), .Y(n511) );
  IBUFFX16_HVT U3 ( .A(n197), .Y(n187) );
  MUX21X1_HVT U4 ( .A1(n325), .A2(n355), .S0(n279), .Y(n513) );
  MUX21X2_HVT U7 ( .A1(n286), .A2(n563), .S0(n247), .Y(n246) );
  INVX2_HVT U8 ( .A(n279), .Y(n247) );
  INVX2_HVT U14 ( .A(n343), .Y(n271) );
  MUX41X1_HVT U16 ( .A1(n517), .A3(n557), .A2(n598), .A4(n398), .S0(n196), 
        .S1(n225), .Y(n516) );
  IBUFFX16_HVT U17 ( .A(n307), .Y(n196) );
  IBUFFX4_HVT U18 ( .A(n313), .Y(n225) );
  IBUFFX16_HVT U20 ( .A(n249), .Y(n197) );
  MUX21X2_HVT U21 ( .A1(n484), .A2(n486), .S0(n198), .Y(n483) );
  IBUFFX16_HVT U22 ( .A(n228), .Y(n198) );
  MUX21X1_HVT U23 ( .A1(n299), .A2(n380), .S0(n227), .Y(n414) );
  IBUFFX2_HVT U24 ( .A(n312), .Y(n227) );
  OR2X4_HVT U26 ( .A1(n285), .A2(n324), .Y(n569) );
  MUX41X1_HVT U27 ( .A1(n540), .A3(n537), .A2(n539), .A4(n536), .S0(n199), 
        .S1(n200), .Y(n535) );
  IBUFFX16_HVT U28 ( .A(n249), .Y(n199) );
  IBUFFX16_HVT U29 ( .A(n266), .Y(n200) );
  INVX0_HVT U30 ( .A(n562), .Y(n353) );
  MUX21X2_HVT U31 ( .A1(n325), .A2(n319), .S0(n267), .Y(n579) );
  MUX21X2_HVT U33 ( .A1(n513), .A2(n514), .S0(n201), .Y(n512) );
  IBUFFX16_HVT U34 ( .A(n260), .Y(n201) );
  MUX21X1_HVT U35 ( .A1(n300), .A2(n579), .S0(n225), .Y(n456) );
  MUX21X1_HVT U36 ( .A1(n205), .A2(n324), .S0(n332), .Y(n202) );
  IBUFFX16_HVT U37 ( .A(n315), .Y(n205) );
  MUX41X1_HVT U39 ( .A1(n350), .A3(n202), .A2(n353), .A4(n235), .S0(n208), 
        .S1(n279), .Y(n425) );
  IBUFFX16_HVT U40 ( .A(n245), .Y(n208) );
  INVX2_HVT U41 ( .A(n342), .Y(n343) );
  INVX1_HVT U43 ( .A(n582), .Y(n366) );
  INVX0_HVT U44 ( .A(n325), .Y(n284) );
  MUX21X1_HVT U45 ( .A1(n396), .A2(n399), .S0(n210), .Y(n582) );
  IBUFFX16_HVT U46 ( .A(n334), .Y(n210) );
  MUX21X2_HVT U47 ( .A1(n515), .A2(n603), .S0(n334), .Y(n514) );
  NBUFFX4_HVT U48 ( .A(n276), .Y(n317) );
  MUX21X2_HVT U49 ( .A1(n366), .A2(n235), .S0(n310), .Y(n541) );
  NAND2X0_HVT U50 ( .A1(n462), .A2(n263), .Y(n252) );
  MUX21X1_HVT U51 ( .A1(n605), .A2(n219), .S0(n336), .Y(n218) );
  IBUFFX16_HVT U52 ( .A(n218), .Y(n437) );
  IBUFFX16_HVT U54 ( .A(n238), .Y(n219) );
  MUX41X1_HVT U57 ( .A1(n437), .A3(n299), .A2(n298), .A4(n301), .S0(n220), 
        .S1(n261), .Y(n436) );
  IBUFFX16_HVT U58 ( .A(n309), .Y(n220) );
  MUX21X2_HVT U59 ( .A1(n281), .A2(n398), .S0(n268), .Y(n580) );
  MUX21X1_HVT U61 ( .A1(n495), .A2(n496), .S0(n311), .Y(n494) );
  IBUFFX2_HVT U63 ( .A(n565), .Y(n377) );
  INVX0_HVT U64 ( .A(n281), .Y(n221) );
  INVX1_HVT U68 ( .A(n221), .Y(n222) );
  INVX0_HVT U69 ( .A(n337), .Y(n223) );
  INVX1_HVT U70 ( .A(n223), .Y(n224) );
  INVX1_HVT U75 ( .A(in[0]), .Y(n337) );
  IBUFFX2_HVT U76 ( .A(n337), .Y(n334) );
  IBUFFX2_HVT U77 ( .A(n337), .Y(n335) );
  INVX0_HVT U79 ( .A(n337), .Y(n332) );
  INVX0_HVT U86 ( .A(n337), .Y(n333) );
  INVX0_HVT U87 ( .A(n224), .Y(n268) );
  MUX21X2_HVT U90 ( .A1(n552), .A2(n553), .S0(n226), .Y(n551) );
  IBUFFX16_HVT U91 ( .A(n310), .Y(n226) );
  IBUFFX16_HVT U92 ( .A(n321), .Y(n228) );
  INVX1_HVT U93 ( .A(n577), .Y(n370) );
  XOR2X1_HVT U94 ( .A1(n326), .A2(n258), .Y(n229) );
  IBUFFX16_HVT U95 ( .A(n229), .Y(n556) );
  MUX41X1_HVT U97 ( .A1(n421), .A3(n420), .A2(n419), .A4(n246), .S0(n230), 
        .S1(n231), .Y(n418) );
  IBUFFX16_HVT U98 ( .A(n305), .Y(n230) );
  IBUFFX16_HVT U101 ( .A(n266), .Y(n231) );
  MUX21X2_HVT U102 ( .A1(n385), .A2(n561), .S0(n232), .Y(n451) );
  IBUFFX16_HVT U103 ( .A(n313), .Y(n232) );
  MUX21X1_HVT U106 ( .A1(n303), .A2(n284), .S0(n333), .Y(n283) );
  MUX41X1_HVT U107 ( .A1(n350), .A3(n300), .A2(n283), .A4(n369), .S0(n233), 
        .S1(n234), .Y(n519) );
  IBUFFX16_HVT U111 ( .A(n245), .Y(n233) );
  IBUFFX16_HVT U113 ( .A(n344), .Y(n234) );
  INVX1_HVT U117 ( .A(n333), .Y(n338) );
  MUX21X2_HVT U121 ( .A1(n300), .A2(n556), .S0(n314), .Y(n420) );
  OA21X1_HVT U123 ( .A1(n348), .A2(n343), .A3(n356), .Y(n455) );
  INVX1_HVT U125 ( .A(n350), .Y(n235) );
  IBUFFX2_HVT U126 ( .A(n337), .Y(n267) );
  INVX0_HVT U128 ( .A(n602), .Y(n350) );
  MUX21X1_HVT U134 ( .A1(n281), .A2(n238), .S0(n333), .Y(n563) );
  INVX1_HVT U135 ( .A(n575), .Y(n372) );
  NAND2X0_HVT U138 ( .A1(n336), .A2(n330), .Y(n602) );
  INVX1_HVT U139 ( .A(n256), .Y(n261) );
  INVX0_HVT U143 ( .A(n327), .Y(n257) );
  INVX1_HVT U144 ( .A(n401), .Y(n394) );
  OA21X1_HVT U146 ( .A1(n372), .A2(n344), .A3(n544), .Y(n419) );
  MUX21X1_HVT U147 ( .A1(n354), .A2(n563), .S0(n314), .Y(n496) );
  OA21X1_HVT U148 ( .A1(n349), .A2(n343), .A3(n583), .Y(n529) );
  INVX1_HVT U149 ( .A(in[5]), .Y(n323) );
  INVX1_HVT U150 ( .A(n323), .Y(n249) );
  INVX0_HVT U152 ( .A(n302), .Y(n239) );
  INVX0_HVT U153 ( .A(n601), .Y(n351) );
  INVX1_HVT U154 ( .A(n603), .Y(n238) );
  INVX1_HVT U157 ( .A(n292), .Y(n263) );
  INVX1_HVT U158 ( .A(in[7]), .Y(n292) );
  INVX1_HVT U160 ( .A(n260), .Y(n275) );
  INVX1_HVT U161 ( .A(n310), .Y(n260) );
  INVX1_HVT U165 ( .A(n304), .Y(n245) );
  INVX1_HVT U167 ( .A(n322), .Y(n242) );
  INVX1_HVT U168 ( .A(n321), .Y(n272) );
  INVX1_HVT U169 ( .A(in[1]), .Y(n320) );
  INVX1_HVT U170 ( .A(n272), .Y(n266) );
  INVX0_HVT U171 ( .A(n342), .Y(n279) );
  INVX1_HVT U175 ( .A(in[4]), .Y(n344) );
  INVX0_HVT U176 ( .A(n344), .Y(n256) );
  INVX1_HVT U180 ( .A(n344), .Y(n342) );
  INVX1_HVT U181 ( .A(n343), .Y(n340) );
  NAND2X0_HVT U182 ( .A1(n279), .A2(n295), .Y(n236) );
  NAND2X0_HVT U184 ( .A1(n550), .A2(n313), .Y(n237) );
  NAND2X0_HVT U186 ( .A1(n236), .A2(n237), .Y(n546) );
  MUX21X1_HVT U187 ( .A1(n546), .A2(n545), .S0(n310), .Y(n543) );
  OR2X1_HVT U188 ( .A1(n258), .A2(n238), .Y(n598) );
  OR2X1_HVT U189 ( .A1(n276), .A2(n280), .Y(n603) );
  INVX1_HVT U190 ( .A(n280), .Y(n281) );
  MUX21X2_HVT U193 ( .A1(n530), .A2(n529), .S0(n311), .Y(n528) );
  NAND2X0_HVT U196 ( .A1(n367), .A2(n239), .Y(n240) );
  NAND2X0_HVT U197 ( .A1(n548), .A2(n302), .Y(n241) );
  NAND2X0_HVT U199 ( .A1(n240), .A2(n241), .Y(n547) );
  MUX21X1_HVT U201 ( .A1(n368), .A2(n601), .S0(n311), .Y(n548) );
  NAND2X0_HVT U202 ( .A1(n427), .A2(n242), .Y(n243) );
  NAND2X0_HVT U203 ( .A1(n429), .A2(n322), .Y(n244) );
  NAND2X0_HVT U204 ( .A1(n243), .A2(n244), .Y(n426) );
  MUX21X2_HVT U205 ( .A1(n497), .A2(n487), .S0(n292), .Y(out[3]) );
  MUX41X1_HVT U206 ( .A1(n282), .A3(n506), .A2(n390), .A4(n592), .S0(n340), 
        .S1(n245), .Y(n505) );
  INVX4_HVT U208 ( .A(n261), .Y(n262) );
  INVX1_HVT U209 ( .A(n337), .Y(n336) );
  MUX21X1_HVT U210 ( .A1(n329), .A2(n287), .S0(n333), .Y(n286) );
  INVX1_HVT U211 ( .A(n352), .Y(n248) );
  INVX0_HVT U212 ( .A(n599), .Y(n352) );
  NAND2X0_HVT U213 ( .A1(n460), .A2(n308), .Y(n250) );
  NAND2X0_HVT U214 ( .A1(n461), .A2(n260), .Y(n251) );
  NAND2X0_HVT U215 ( .A1(n250), .A2(n251), .Y(n459) );
  NAND2X0_HVT U216 ( .A1(n452), .A2(n292), .Y(n253) );
  NAND2X0_HVT U217 ( .A1(n252), .A2(n253), .Y(out[5]) );
  AO21X1_HVT U218 ( .A1(n314), .A2(n285), .A3(n396), .Y(n460) );
  MUX21X1_HVT U219 ( .A1(n394), .A2(n351), .S0(n312), .Y(n461) );
  NAND2X0_HVT U220 ( .A1(n438), .A2(n263), .Y(n254) );
  NAND2X0_HVT U221 ( .A1(n431), .A2(n292), .Y(n255) );
  NAND2X0_HVT U222 ( .A1(n254), .A2(n255), .Y(out[6]) );
  MUX21X1_HVT U223 ( .A1(n316), .A2(n238), .S0(n336), .Y(n561) );
  MUX21X1_HVT U224 ( .A1(n284), .A2(n303), .S0(n334), .Y(n288) );
  MUX41X1_HVT U225 ( .A1(n372), .A3(n586), .A2(n288), .A4(n587), .S0(n307), 
        .S1(n256), .Y(n526) );
  IBUFFX2_HVT U226 ( .A(n343), .Y(n341) );
  NAND2X0_HVT U227 ( .A1(n542), .A2(in[7]), .Y(n269) );
  OR2X1_HVT U228 ( .A1(n258), .A2(n257), .Y(n597) );
  INVX1_HVT U229 ( .A(n569), .Y(n355) );
  MUX41X1_HVT U230 ( .A1(n390), .A3(n501), .A2(n328), .A4(n353), .S0(n341), 
        .S1(n307), .Y(n500) );
  MUX41X1_HVT U231 ( .A1(n447), .A3(n443), .A2(n445), .A4(n439), .S0(n323), 
        .S1(n242), .Y(n438) );
  INVX1_HVT U232 ( .A(n333), .Y(n258) );
  INVX2_HVT U233 ( .A(n258), .Y(n259) );
  AO21X1_HVT U234 ( .A1(n588), .A2(n235), .A3(n343), .Y(n440) );
  IBUFFX2_HVT U235 ( .A(n288), .Y(n573) );
  MUX41X1_HVT U236 ( .A1(n376), .A3(n509), .A2(n576), .A4(n389), .S0(n279), 
        .S1(n275), .Y(n508) );
  NAND2X0_HVT U237 ( .A1(n511), .A2(n263), .Y(n264) );
  NAND2X0_HVT U238 ( .A1(n504), .A2(n292), .Y(n265) );
  NAND2X0_HVT U239 ( .A1(n264), .A2(n265), .Y(out[2]) );
  MUX21X1_HVT U240 ( .A1(n422), .A2(n386), .S0(n312), .Y(n421) );
  MUX41X1_HVT U241 ( .A1(n418), .A3(n412), .A2(n426), .A4(n423), .S0(n323), 
        .S1(n263), .Y(out[7]) );
  NAND2X0_HVT U242 ( .A1(n535), .A2(n292), .Y(n270) );
  NAND2X0_HVT U243 ( .A1(n269), .A2(n270), .Y(out[0]) );
  MUX41X1_HVT U244 ( .A1(n277), .A3(n359), .A2(n331), .A4(n360), .S0(n245), 
        .S1(n340), .Y(n536) );
  MUX41X1_HVT U245 ( .A1(n469), .A3(n477), .A2(n473), .A4(n483), .S0(n263), 
        .S1(n249), .Y(out[4]) );
  MUX21X2_HVT U246 ( .A1(n470), .A2(n471), .S0(n321), .Y(n469) );
  INVX1_HVT U247 ( .A(n320), .Y(n321) );
  IBUFFX2_HVT U248 ( .A(n561), .Y(n379) );
  MUX21X2_HVT U249 ( .A1(n450), .A2(n451), .S0(n311), .Y(n447) );
  INVX1_HVT U250 ( .A(n605), .Y(n398) );
  INVX0_HVT U251 ( .A(n282), .Y(n568) );
  INVX0_HVT U252 ( .A(n289), .Y(n560) );
  INVX0_HVT U253 ( .A(n295), .Y(n581) );
  NAND2X0_HVT U254 ( .A1(n365), .A2(n239), .Y(n290) );
  INVX1_HVT U255 ( .A(n276), .Y(n277) );
  INVX1_HVT U256 ( .A(in[6]), .Y(n280) );
  INVX1_HVT U257 ( .A(in[3]), .Y(n276) );
  INVX0_HVT U258 ( .A(n319), .Y(n287) );
  AO21X2_HVT U259 ( .A1(n224), .A2(n331), .A3(n343), .Y(n448) );
  MUX41X1_HVT U260 ( .A1(n559), .A3(n428), .A2(n345), .A4(n572), .S0(n245), 
        .S1(n344), .Y(n427) );
  MUX41X1_HVT U261 ( .A1(n468), .A3(n466), .A2(n465), .A4(n463), .S0(n320), 
        .S1(n323), .Y(n462) );
  NAND2X0_HVT U262 ( .A1(n424), .A2(n242), .Y(n273) );
  NAND2X0_HVT U263 ( .A1(n425), .A2(n321), .Y(n274) );
  NAND2X0_HVT U264 ( .A1(n274), .A2(n273), .Y(n423) );
  MUX41X1_HVT U265 ( .A1(n510), .A3(n507), .A2(n508), .A4(n505), .S0(n323), 
        .S1(n242), .Y(n504) );
  MUX21X2_HVT U266 ( .A1(n520), .A2(n527), .S0(n263), .Y(out[1]) );
  AO21X2_HVT U267 ( .A1(n336), .A2(n396), .A3(n343), .Y(n415) );
  NAND2X0_HVT U268 ( .A1(n315), .A2(n318), .Y(n278) );
  INVX0_HVT U269 ( .A(n597), .Y(n285) );
  MUX41X1_HVT U270 ( .A1(n434), .A3(n436), .A2(n432), .A4(n433), .S0(n321), 
        .S1(n323), .Y(n431) );
  MUX21X1_HVT U271 ( .A1(n324), .A2(n287), .S0(n258), .Y(n282) );
  INVX1_HVT U272 ( .A(n324), .Y(n399) );
  NBUFFX2_HVT U273 ( .A(n605), .Y(n331) );
  XNOR2X2_HVT U274 ( .A1(n318), .A2(n317), .Y(n588) );
  MUX21X1_HVT U275 ( .A1(n278), .A2(n331), .S0(n224), .Y(n590) );
  MUX21X1_HVT U276 ( .A1(n303), .A2(n326), .S0(n224), .Y(n289) );
  NAND2X0_HVT U277 ( .A1(n541), .A2(n302), .Y(n291) );
  NAND2X0_HVT U278 ( .A1(n290), .A2(n291), .Y(n540) );
  INVX1_HVT U279 ( .A(n583), .Y(n365) );
  NAND2X0_HVT U280 ( .A1(n441), .A2(n260), .Y(n293) );
  NAND2X0_HVT U281 ( .A1(n442), .A2(n310), .Y(n294) );
  NAND2X0_HVT U282 ( .A1(n293), .A2(n294), .Y(n439) );
  MUX21X1_HVT U283 ( .A1(n329), .A2(n276), .S0(n334), .Y(n295) );
  MUX21X1_HVT U284 ( .A1(n578), .A2(n581), .S0(n312), .Y(n442) );
  INVX1_HVT U285 ( .A(n329), .Y(n396) );
  MUX41X1_HVT U286 ( .A1(n581), .A3(n584), .A2(n379), .A4(n397), .S0(n260), 
        .S1(n279), .Y(n465) );
  MUX21X2_HVT U287 ( .A1(n455), .A2(n456), .S0(n311), .Y(n454) );
  NBUFFX2_HVT U288 ( .A(n604), .Y(n329) );
  NBUFFX2_HVT U289 ( .A(n604), .Y(n330) );
  AND2X1_HVT U290 ( .A1(n330), .A2(n589), .Y(n296) );
  MUX21X1_HVT U291 ( .A1(n396), .A2(n399), .S0(n335), .Y(n571) );
  MUX21X1_HVT U292 ( .A1(n318), .A2(n397), .S0(n335), .Y(n458) );
  MUX21X1_HVT U293 ( .A1(n399), .A2(n317), .S0(n336), .Y(n565) );
  MUX21X1_HVT U294 ( .A1(n318), .A2(n396), .S0(n268), .Y(n578) );
  MUX21X1_HVT U295 ( .A1(n326), .A2(n603), .S0(n334), .Y(n446) );
  MUX21X1_HVT U296 ( .A1(n398), .A2(n319), .S0(n336), .Y(n435) );
  NAND2X0_HVT U297 ( .A1(n315), .A2(n318), .Y(n604) );
  MUX21X1_HVT U298 ( .A1(n399), .A2(n319), .S0(n334), .Y(n402) );
  MUX21X1_HVT U299 ( .A1(n325), .A2(n316), .S0(n332), .Y(n583) );
  MUX21X1_HVT U300 ( .A1(n398), .A2(n397), .S0(n335), .Y(n576) );
  MUX21X1_HVT U301 ( .A1(n317), .A2(n396), .S0(n334), .Y(n574) );
  MUX21X1_HVT U302 ( .A1(n393), .A2(n297), .S0(n310), .Y(n482) );
  MUX21X1_HVT U303 ( .A1(n325), .A2(n319), .S0(n313), .Y(n515) );
  INVX1_HVT U304 ( .A(n326), .Y(n397) );
  MUX21X1_HVT U305 ( .A1(n571), .A2(n296), .S0(n311), .Y(n479) );
  MUX21X1_HVT U306 ( .A1(n326), .A2(n278), .S0(n335), .Y(n401) );
  XNOR2X1_HVT U307 ( .A1(n329), .A2(n268), .Y(n297) );
  MUX21X1_HVT U308 ( .A1(n325), .A2(n397), .S0(n268), .Y(n570) );
  MUX21X1_HVT U309 ( .A1(n316), .A2(n330), .S0(n267), .Y(n408) );
  MUX21X1_HVT U310 ( .A1(n318), .A2(n278), .S0(n332), .Y(n501) );
  XOR2X1_HVT U311 ( .A1(n324), .A2(n267), .Y(n558) );
  MUX21X1_HVT U312 ( .A1(n238), .A2(n316), .S0(n267), .Y(n409) );
  MUX21X1_HVT U313 ( .A1(n328), .A2(n330), .S0(n335), .Y(n586) );
  XOR2X1_HVT U314 ( .A1(n328), .A2(n267), .Y(n557) );
  MUX21X1_HVT U315 ( .A1(n319), .A2(n325), .S0(n259), .Y(n564) );
  MUX21X1_HVT U316 ( .A1(n603), .A2(n317), .S0(n259), .Y(n585) );
  MUX21X1_HVT U317 ( .A1(n317), .A2(n318), .S0(n334), .Y(n559) );
  AND2X1_HVT U318 ( .A1(n248), .A2(n330), .Y(n298) );
  MUX21X1_HVT U319 ( .A1(n328), .A2(n318), .S0(n259), .Y(n485) );
  MUX21X1_HVT U320 ( .A1(n315), .A2(n603), .S0(n335), .Y(n404) );
  AND2X1_HVT U321 ( .A1(n267), .A2(n319), .Y(n299) );
  NBUFFX2_HVT U322 ( .A(n342), .Y(n314) );
  NBUFFX2_HVT U323 ( .A(n342), .Y(n313) );
  NBUFFX2_HVT U324 ( .A(n342), .Y(n312) );
  NBUFFX2_HVT U325 ( .A(n280), .Y(n318) );
  NBUFFX2_HVT U326 ( .A(n588), .Y(n324) );
  NBUFFX2_HVT U327 ( .A(n276), .Y(n315) );
  NBUFFX2_HVT U328 ( .A(n588), .Y(n325) );
  MUX21X1_HVT U329 ( .A1(n370), .A2(n360), .S0(n314), .Y(n553) );
  MUX21X1_HVT U330 ( .A1(n396), .A2(n238), .S0(n268), .Y(n554) );
  MUX21X1_HVT U331 ( .A1(n329), .A2(n327), .S0(n334), .Y(n464) );
  NBUFFX2_HVT U332 ( .A(n600), .Y(n326) );
  AND2X1_HVT U333 ( .A1(n328), .A2(n338), .Y(n300) );
  AND2X1_HVT U334 ( .A1(n238), .A2(n338), .Y(n301) );
  MUX21X1_HVT U335 ( .A1(n385), .A2(n346), .S0(n314), .Y(n530) );
  XOR2X1_HVT U336 ( .A1(n605), .A2(n335), .Y(n567) );
  NBUFFX2_HVT U337 ( .A(n600), .Y(n327) );
  NBUFFX2_HVT U338 ( .A(n603), .Y(n328) );
  NBUFFX2_HVT U339 ( .A(n280), .Y(n319) );
  NBUFFX2_HVT U340 ( .A(n276), .Y(n316) );
  NBUFFX2_HVT U341 ( .A(n305), .Y(n309) );
  NBUFFX2_HVT U342 ( .A(n339), .Y(n311) );
  NBUFFX2_HVT U343 ( .A(n339), .Y(n310) );
  XNOR2X1_HVT U344 ( .A1(n344), .A2(n306), .Y(n302) );
  NBUFFX2_HVT U345 ( .A(n339), .Y(n306) );
  NBUFFX2_HVT U346 ( .A(n304), .Y(n308) );
  NBUFFX2_HVT U347 ( .A(n339), .Y(n304) );
  NBUFFX2_HVT U348 ( .A(n339), .Y(n305) );
  NBUFFX2_HVT U349 ( .A(n339), .Y(n307) );
  INVX1_HVT U350 ( .A(n320), .Y(n322) );
  MUX21X1_HVT U351 ( .A1(n398), .A2(n277), .S0(n259), .Y(n400) );
  MUX21X1_HVT U352 ( .A1(n331), .A2(n277), .S0(n268), .Y(n449) );
  MUX21X1_HVT U353 ( .A1(n474), .A2(n475), .S0(n322), .Y(n473) );
  MUX21X1_HVT U354 ( .A1(n327), .A2(n277), .S0(n268), .Y(n509) );
  XOR2X1_HVT U355 ( .A1(n332), .A2(n222), .Y(n555) );
  MUX21X1_HVT U356 ( .A1(n396), .A2(n222), .S0(n267), .Y(n472) );
  MUX21X1_HVT U357 ( .A1(n281), .A2(n397), .S0(n259), .Y(n411) );
  MUX21X1_HVT U358 ( .A1(n238), .A2(n397), .S0(n268), .Y(n490) );
  MUX21X1_HVT U359 ( .A1(n327), .A2(n281), .S0(n332), .Y(n575) );
  MUX21X1_HVT U360 ( .A1(n281), .A2(n303), .S0(n332), .Y(n587) );
  MUX21X1_HVT U361 ( .A1(n277), .A2(n331), .S0(n267), .Y(n406) );
  MUX21X1_HVT U362 ( .A1(n277), .A2(n327), .S0(n267), .Y(n405) );
  MUX21X1_HVT U363 ( .A1(n319), .A2(n277), .S0(n335), .Y(n577) );
  MUX21X1_HVT U364 ( .A1(n315), .A2(n222), .S0(n259), .Y(n403) );
  MUX21X1_HVT U365 ( .A1(n222), .A2(n328), .S0(n332), .Y(n410) );
  MUX21X1_HVT U366 ( .A1(n603), .A2(n222), .S0(n336), .Y(n407) );
  NBUFFX2_HVT U367 ( .A(in[2]), .Y(n339) );
  NAND2X0_HVT U368 ( .A1(n277), .A2(n319), .Y(n303) );
  INVX0_HVT U369 ( .A(n593), .Y(n345) );
  INVX0_HVT U370 ( .A(n572), .Y(n346) );
  INVX0_HVT U371 ( .A(n566), .Y(n347) );
  INVX0_HVT U372 ( .A(n506), .Y(n348) );
  INVX0_HVT U373 ( .A(n467), .Y(n349) );
  INVX0_HVT U374 ( .A(n598), .Y(n354) );
  INVX0_HVT U375 ( .A(n591), .Y(n356) );
  INVX0_HVT U376 ( .A(n596), .Y(n357) );
  INVX0_HVT U377 ( .A(n592), .Y(n358) );
  INVX0_HVT U378 ( .A(n590), .Y(n359) );
  INVX0_HVT U379 ( .A(n589), .Y(n360) );
  INVX0_HVT U380 ( .A(n587), .Y(n361) );
  INVX0_HVT U381 ( .A(n586), .Y(n362) );
  INVX0_HVT U382 ( .A(n585), .Y(n363) );
  INVX0_HVT U383 ( .A(n584), .Y(n364) );
  INVX0_HVT U384 ( .A(n580), .Y(n367) );
  INVX0_HVT U385 ( .A(n579), .Y(n368) );
  INVX0_HVT U386 ( .A(n578), .Y(n369) );
  INVX0_HVT U387 ( .A(n576), .Y(n371) );
  INVX0_HVT U388 ( .A(n574), .Y(n373) );
  INVX0_HVT U389 ( .A(n571), .Y(n374) );
  INVX0_HVT U390 ( .A(n570), .Y(n375) );
  INVX0_HVT U391 ( .A(n567), .Y(n376) );
  INVX0_HVT U392 ( .A(n564), .Y(n378) );
  INVX0_HVT U393 ( .A(n559), .Y(n380) );
  INVX0_HVT U394 ( .A(n558), .Y(n381) );
  INVX0_HVT U395 ( .A(n595), .Y(n382) );
  INVX0_HVT U396 ( .A(n411), .Y(n383) );
  INVX0_HVT U397 ( .A(n410), .Y(n384) );
  INVX0_HVT U398 ( .A(n409), .Y(n385) );
  INVX0_HVT U399 ( .A(n408), .Y(n386) );
  INVX0_HVT U400 ( .A(n407), .Y(n387) );
  INVX0_HVT U401 ( .A(n406), .Y(n388) );
  INVX0_HVT U402 ( .A(n405), .Y(n389) );
  INVX0_HVT U403 ( .A(n404), .Y(n390) );
  INVX0_HVT U404 ( .A(n403), .Y(n391) );
  INVX0_HVT U405 ( .A(n449), .Y(n392) );
  INVX0_HVT U406 ( .A(n402), .Y(n393) );
  INVX0_HVT U407 ( .A(n400), .Y(n395) );
endmodule

