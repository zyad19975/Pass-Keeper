
module sbox_0 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n214, n215,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n23,
         n48, n210, n211, n212, n213, n216, n217, n218, n219, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357;

  NAND2X0_HVT U3 ( .A1(n285), .A2(n282), .Y(n3) );
  NAND2X0_HVT U4 ( .A1(n281), .A2(n3), .Y(n4) );
  NAND2X0_HVT U5 ( .A1(n289), .A2(n269), .Y(n6) );
  NAND2X0_HVT U13 ( .A1(n14), .A2(n284), .Y(n13) );
  NAND2X0_HVT U15 ( .A1(n3), .A2(n271), .Y(n16) );
  NAND2X0_HVT U21 ( .A1(n280), .A2(n291), .Y(n22) );
  NAND2X0_HVT U24 ( .A1(n277), .A2(n291), .Y(n25) );
  NAND2X0_HVT U33 ( .A1(n352), .A2(n291), .Y(n34) );
  NAND2X0_HVT U35 ( .A1(n275), .A2(n290), .Y(n36) );
  NAND2X0_HVT U42 ( .A1(n233), .A2(n277), .Y(n43) );
  MUX41X1_HVT U51 ( .A1(n340), .A3(n298), .A2(n315), .A4(n316), .S0(n236), 
        .S1(n293), .Y(n52) );
  NAND2X0_HVT U53 ( .A1(n55), .A2(n44), .Y(n54) );
  NAND2X0_HVT U56 ( .A1(n281), .A2(n59), .Y(n58) );
  MUX41X1_HVT U57 ( .A1(n341), .A3(n20), .A2(n58), .A4(n11), .S0(n217), .S1(
        n293), .Y(n60) );
  NAND2X0_HVT U58 ( .A1(n284), .A2(n3), .Y(n61) );
  MUX41X1_HVT U59 ( .A1(n258), .A3(n61), .A2(n256), .A4(n314), .S0(n236), .S1(
        n293), .Y(n62) );
  MUX41X1_HVT U61 ( .A1(n254), .A3(n313), .A2(n312), .A4(n270), .S0(n218), 
        .S1(n293), .Y(n64) );
  NAND2X0_HVT U62 ( .A1(n291), .A2(n283), .Y(n65) );
  MUX41X1_HVT U63 ( .A1(n65), .A3(n305), .A2(n335), .A4(n311), .S0(n236), .S1(
        n293), .Y(n66) );
  AO21X1_HVT U66 ( .A1(n309), .A2(n266), .A3(n334), .Y(n69) );
  MUX41X1_HVT U68 ( .A1(n307), .A3(n69), .A2(n70), .A4(n68), .S0(n259), .S1(
        n236), .Y(n71) );
  MUX41X1_HVT U69 ( .A1(n71), .A3(n63), .A2(n67), .A4(n57), .S0(in[6]), .S1(
        n276), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n278), .A2(n76), .Y(n75) );
  MUX41X1_HVT U74 ( .A1(n74), .A3(n27), .A2(n75), .A4(n25), .S0(n261), .S1(
        n218), .Y(n77) );
  MUX41X1_HVT U75 ( .A1(n338), .A3(n343), .A2(n356), .A4(n318), .S0(n259), 
        .S1(n218), .Y(n78) );
  MUX41X1_HVT U77 ( .A1(n9), .A3(n345), .A2(n79), .A4(n344), .S0(n267), .S1(
        n264), .Y(n80) );
  MUX41X1_HVT U78 ( .A1(n80), .A3(n77), .A2(n78), .A4(n73), .S0(n276), .S1(
        in[5]), .Y(n81) );
  AND3X1_HVT U80 ( .A1(n282), .A2(n59), .A3(n84), .Y(n83) );
  MUX41X1_HVT U82 ( .A1(n46), .A3(n316), .A2(n299), .A4(n15), .S0(n259), .S1(
        n267), .Y(n86) );
  AND2X1_HVT U83 ( .A1(n287), .A2(n237), .Y(n87) );
  MUX41X1_HVT U84 ( .A1(n317), .A3(n7), .A2(n17), .A4(n87), .S0(n259), .S1(
        n294), .Y(n88) );
  NAND2X0_HVT U85 ( .A1(n291), .A2(n355), .Y(n89) );
  MUX41X1_HVT U86 ( .A1(n343), .A3(n89), .A2(n255), .A4(n251), .S0(n259), .S1(
        n217), .Y(n90) );
  MUX41X1_HVT U87 ( .A1(n90), .A3(n86), .A2(n88), .A4(n85), .S0(in[0]), .S1(
        n265), .Y(n91) );
  MUX41X1_HVT U90 ( .A1(n47), .A3(n43), .A2(n340), .A4(n92), .S0(n260), .S1(
        n294), .Y(n93) );
  AO21X1_HVT U93 ( .A1(n268), .A2(n97), .A3(n339), .Y(n96) );
  MUX41X1_HVT U96 ( .A1(n299), .A3(n253), .A2(n342), .A4(n99), .S0(n259), .S1(
        n236), .Y(n100) );
  MUX41X1_HVT U97 ( .A1(n338), .A3(n253), .A2(n234), .A4(n16), .S0(n259), .S1(
        n267), .Y(n101) );
  MUX41X1_HVT U98 ( .A1(n101), .A3(n98), .A2(n100), .A4(n93), .S0(n276), .S1(
        n265), .Y(n102) );
  NAND2X0_HVT U101 ( .A1(n106), .A2(n107), .Y(n105) );
  MUX41X1_HVT U103 ( .A1(n3), .A3(n308), .A2(n321), .A4(n36), .S0(n259), .S1(
        n241), .Y(n109) );
  MUX41X1_HVT U105 ( .A1(n320), .A3(n49), .A2(n110), .A4(n337), .S0(n259), 
        .S1(n295), .Y(n111) );
  NAND2X0_HVT U110 ( .A1(n282), .A2(n116), .Y(n115) );
  MUX41X1_HVT U114 ( .A1(n119), .A3(n113), .A2(n117), .A4(n114), .S0(n266), 
        .S1(n217), .Y(n120) );
  AND2X1_HVT U115 ( .A1(n288), .A2(n270), .Y(n121) );
  MUX41X1_HVT U116 ( .A1(n13), .A3(n121), .A2(n318), .A4(n32), .S0(n260), .S1(
        n218), .Y(n122) );
  NAND2X0_HVT U123 ( .A1(n130), .A2(n131), .Y(n129) );
  MUX41X1_HVT U125 ( .A1(n22), .A3(n258), .A2(n307), .A4(n347), .S0(n260), 
        .S1(n294), .Y(n133) );
  AND3X1_HVT U128 ( .A1(n263), .A2(n291), .A3(n237), .Y(n136) );
  MUX41X1_HVT U131 ( .A1(n138), .A3(n136), .A2(n137), .A4(n135), .S0(n266), 
        .S1(n236), .Y(n139) );
  MUX41X1_HVT U132 ( .A1(n139), .A3(n126), .A2(n134), .A4(n120), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  MUX41X1_HVT U136 ( .A1(n251), .A3(n34), .A2(n349), .A4(n37), .S0(n260), .S1(
        n217), .Y(n143) );
  MUX41X1_HVT U139 ( .A1(n145), .A3(n142), .A2(n143), .A4(n141), .S0(n276), 
        .S1(n293), .Y(n146) );
  AND2X1_HVT U140 ( .A1(n279), .A2(n291), .Y(n147) );
  MUX41X1_HVT U141 ( .A1(n26), .A3(n329), .A2(n147), .A4(n325), .S0(n261), 
        .S1(n294), .Y(n148) );
  NAND2X0_HVT U146 ( .A1(n234), .A2(n284), .Y(n76) );
  MUX41X1_HVT U147 ( .A1(n349), .A3(n76), .A2(n338), .A4(n47), .S0(n261), .S1(
        n295), .Y(n153) );
  MUX41X1_HVT U153 ( .A1(n115), .A3(n254), .A2(n2), .A4(n301), .S0(n260), .S1(
        n294), .Y(n159) );
  AND2X1_HVT U154 ( .A1(n268), .A2(n277), .Y(n160) );
  NAND2X0_HVT U158 ( .A1(n286), .A2(n355), .Y(n164) );
  MUX41X1_HVT U159 ( .A1(n13), .A3(n270), .A2(n164), .A4(n248), .S0(n262), 
        .S1(n217), .Y(n165) );
  MUX41X1_HVT U160 ( .A1(n165), .A3(n159), .A2(n163), .A4(n158), .S0(n276), 
        .S1(n265), .Y(n166) );
  AND2X1_HVT U162 ( .A1(n7), .A2(n76), .Y(n168) );
  MUX41X1_HVT U165 ( .A1(n22), .A3(n322), .A2(n47), .A4(n170), .S0(n218), .S1(
        n262), .Y(n171) );
  NAND2X0_HVT U166 ( .A1(n284), .A2(n59), .Y(n172) );
  NAND2X0_HVT U167 ( .A1(n356), .A2(n291), .Y(n173) );
  MUX41X1_HVT U168 ( .A1(n341), .A3(n279), .A2(n173), .A4(n172), .S0(n262), 
        .S1(n218), .Y(n174) );
  NAND2X0_HVT U174 ( .A1(n288), .A2(n7), .Y(n14) );
  NAND2X0_HVT U177 ( .A1(n285), .A2(n274), .Y(n181) );
  MUX41X1_HVT U178 ( .A1(n18), .A3(n181), .A2(n350), .A4(n39), .S0(n261), .S1(
        n218), .Y(n182) );
  MUX41X1_HVT U179 ( .A1(n29), .A3(n351), .A2(n303), .A4(n350), .S0(n259), 
        .S1(n294), .Y(n183) );
  MUX41X1_HVT U181 ( .A1(n184), .A3(n182), .A2(n183), .A4(n180), .S0(n276), 
        .S1(n265), .Y(n185) );
  MUX41X1_HVT U186 ( .A1(n253), .A3(n40), .A2(n76), .A4(n47), .S0(n259), .S1(
        n217), .Y(n190) );
  MUX41X1_HVT U195 ( .A1(n7), .A3(n342), .A2(n1), .A4(n38), .S0(n262), .S1(
        n295), .Y(n198) );
  AO21X1_HVT U197 ( .A1(n255), .A2(n268), .A3(n339), .Y(n200) );
  MUX41X1_HVT U204 ( .A1(n58), .A3(n13), .A2(n326), .A4(n24), .S0(n259), .S1(
        n295), .Y(n207) );
  MUX41X1_HVT U205 ( .A1(n237), .A3(n3), .A2(n351), .A4(n324), .S0(n264), .S1(
        n241), .Y(n208) );
  MUX41X1_HVT U206 ( .A1(n208), .A3(n206), .A2(n207), .A4(n205), .S0(n276), 
        .S1(n265), .Y(n209) );
  NAND2X0_HVT U208 ( .A1(n287), .A2(n280), .Y(n116) );
  NAND2X0_HVT U212 ( .A1(n234), .A2(n278), .Y(n59) );
  NAND2X0_HVT U214 ( .A1(n7), .A2(n291), .Y(n214) );
  NAND2X0_HVT U215 ( .A1(n116), .A2(n279), .Y(n215) );
  NAND2X0_HVT U218 ( .A1(n353), .A2(n285), .Y(n157) );
  NAND2X0_HVT U220 ( .A1(n294), .A2(n214), .Y(n84) );
  XNOR2X2_HVT U1 ( .A1(n273), .A2(in[3]), .Y(n23) );
  INVX8_HVT U2 ( .A(n23), .Y(n7) );
  MUX41X1_HVT U6 ( .A1(n346), .A3(n14), .A2(n273), .A4(n179), .S0(n48), .S1(
        n292), .Y(n180) );
  IBUFFX16_HVT U7 ( .A(n297), .Y(n48) );
  AO21X2_HVT U8 ( .A1(n264), .A2(n279), .A3(n7), .Y(n124) );
  MUX21X2_HVT U9 ( .A1(n66), .A2(n64), .S0(n262), .Y(n67) );
  NBUFFX4_HVT U10 ( .A(n357), .Y(n273) );
  MUX21X2_HVT U11 ( .A1(n282), .A2(n271), .S0(n287), .Y(n42) );
  INVX1_HVT U12 ( .A(n17), .Y(n312) );
  MUX21X1_HVT U14 ( .A1(n271), .A2(n355), .S0(n210), .Y(n167) );
  IBUFFX16_HVT U16 ( .A(n288), .Y(n210) );
  MUX41X1_HVT U17 ( .A1(n167), .A3(n252), .A2(n168), .A4(n313), .S0(n211), 
        .S1(n212), .Y(n169) );
  IBUFFX16_HVT U18 ( .A(n260), .Y(n211) );
  IBUFFX16_HVT U19 ( .A(n218), .Y(n212) );
  INVX0_HVT U20 ( .A(in[4]), .Y(n213) );
  INVX0_HVT U22 ( .A(in[4]), .Y(n357) );
  INVX0_HVT U23 ( .A(n290), .Y(n286) );
  INVX0_HVT U25 ( .A(n290), .Y(n285) );
  INVX0_HVT U26 ( .A(n290), .Y(n287) );
  AO21X1_HVT U27 ( .A1(n291), .A2(n353), .A3(n297), .Y(n106) );
  NBUFFX2_HVT U28 ( .A(in[4]), .Y(n216) );
  INVX0_HVT U29 ( .A(n213), .Y(n237) );
  INVX0_HVT U30 ( .A(in[7]), .Y(n297) );
  INVX1_HVT U31 ( .A(n296), .Y(n217) );
  INVX1_HVT U32 ( .A(in[7]), .Y(n296) );
  OA21X1_HVT U34 ( .A1(n256), .A2(n297), .A3(n32), .Y(n176) );
  INVX1_HVT U36 ( .A(in[2]), .Y(n292) );
  INVX1_HVT U37 ( .A(in[6]), .Y(n232) );
  NBUFFX2_HVT U38 ( .A(in[7]), .Y(n267) );
  INVX1_HVT U39 ( .A(n296), .Y(n294) );
  INVX1_HVT U40 ( .A(n246), .Y(n241) );
  INVX1_HVT U41 ( .A(n264), .Y(n235) );
  INVX1_HVT U43 ( .A(n293), .Y(n231) );
  INVX1_HVT U44 ( .A(in[0]), .Y(n219) );
  INVX2_HVT U45 ( .A(n296), .Y(n218) );
  MUX41X1_HVT U46 ( .A1(n306), .A3(n13), .A2(n9), .A4(n250), .S0(n264), .S1(
        n267), .Y(n184) );
  MUX41X1_HVT U47 ( .A1(n169), .A3(n174), .A2(n171), .A4(n177), .S0(n219), 
        .S1(n231), .Y(n178) );
  MUX21X2_HVT U48 ( .A1(n133), .A2(n132), .S0(n266), .Y(n134) );
  MUX21X2_HVT U49 ( .A1(n128), .A2(n129), .S0(n268), .Y(n132) );
  MUX21X2_HVT U50 ( .A1(n91), .A2(n81), .S0(in[6]), .Y(out[1]) );
  INVX2_HVT U52 ( .A(n296), .Y(n295) );
  MUX21X2_HVT U54 ( .A1(n202), .A2(n209), .S0(n232), .Y(out[7]) );
  IBUFFX2_HVT U55 ( .A(n290), .Y(n233) );
  INVX0_HVT U60 ( .A(n290), .Y(n234) );
  IBUFFX2_HVT U64 ( .A(n37), .Y(n327) );
  MUX41X1_HVT U65 ( .A1(n201), .A3(n198), .A2(n197), .A4(n196), .S0(n293), 
        .S1(in[0]), .Y(n202) );
  IBUFFX2_HVT U67 ( .A(n38), .Y(n328) );
  MUX21X2_HVT U70 ( .A1(n103), .A2(n254), .S0(n238), .Y(n104) );
  MUX41X1_HVT U71 ( .A1(n195), .A3(n51), .A2(n36), .A4(n43), .S0(n235), .S1(
        n246), .Y(n196) );
  INVX1_HVT U72 ( .A(n267), .Y(n246) );
  MUX21X2_HVT U76 ( .A1(n150), .A2(n151), .S0(n263), .Y(n152) );
  INVX1_HVT U79 ( .A(n229), .Y(n350) );
  MUX41X1_HVT U81 ( .A1(n337), .A3(n191), .A2(n14), .A4(n192), .S0(n246), .S1(
        n292), .Y(n193) );
  MUX21X2_HVT U88 ( .A1(n333), .A2(n350), .S0(n268), .Y(n199) );
  MUX21X2_HVT U89 ( .A1(n185), .A2(n194), .S0(n232), .Y(out[6]) );
  OA21X2_HVT U91 ( .A1(n328), .A2(n292), .A3(n314), .Y(n114) );
  NBUFFX2_HVT U92 ( .A(in[2]), .Y(n262) );
  MUX21X1_HVT U94 ( .A1(n118), .A2(n283), .S0(n50), .Y(n119) );
  MUX21X2_HVT U95 ( .A1(n156), .A2(n155), .S0(n264), .Y(n158) );
  INVX1_HVT U99 ( .A(n224), .Y(n344) );
  INVX1_HVT U100 ( .A(n222), .Y(n342) );
  MUX21X2_HVT U102 ( .A1(n161), .A2(n162), .S0(n235), .Y(n163) );
  NBUFFX2_HVT U104 ( .A(n295), .Y(n236) );
  IBUFFX2_HVT U106 ( .A(in[1]), .Y(n291) );
  IBUFFX2_HVT U107 ( .A(n39), .Y(n329) );
  MUX21X2_HVT U108 ( .A1(n39), .A2(n345), .S0(n267), .Y(n162) );
  OA21X1_HVT U109 ( .A1(n302), .A2(n297), .A3(n32), .Y(n151) );
  INVX0_HVT U111 ( .A(n28), .Y(n249) );
  MUX21X1_HVT U112 ( .A1(n324), .A2(n15), .S0(n264), .Y(n103) );
  OA21X1_HVT U113 ( .A1(n41), .A2(n297), .A3(n157), .Y(n156) );
  INVX0_HVT U117 ( .A(n227), .Y(n348) );
  INVX0_HVT U118 ( .A(n6), .Y(n248) );
  MUX41X1_HVT U119 ( .A1(n10), .A3(n336), .A2(n270), .A4(n317), .S0(n235), 
        .S1(n296), .Y(n149) );
  MUX41X1_HVT U120 ( .A1(n148), .A3(n152), .A2(n149), .A4(n153), .S0(n219), 
        .S1(n231), .Y(n154) );
  XNOR2X1_HVT U121 ( .A1(n292), .A2(n296), .Y(n238) );
  OA21X1_HVT U122 ( .A1(n35), .A2(n297), .A3(n317), .Y(n188) );
  MUX21X1_HVT U124 ( .A1(n144), .A2(n4), .S0(n264), .Y(n145) );
  NBUFFX2_HVT U126 ( .A(n23), .Y(n271) );
  NAND2X0_HVT U127 ( .A1(n277), .A2(n233), .Y(n239) );
  NAND2X0_HVT U129 ( .A1(n272), .A2(n291), .Y(n240) );
  NAND2X0_HVT U130 ( .A1(n239), .A2(n240), .Y(n24) );
  INVX2_HVT U133 ( .A(in[1]), .Y(n290) );
  INVX0_HVT U134 ( .A(n24), .Y(n317) );
  NAND2X0_HVT U135 ( .A1(n250), .A2(n241), .Y(n242) );
  NAND2X0_HVT U137 ( .A1(n17), .A2(n246), .Y(n243) );
  NAND2X0_HVT U138 ( .A1(n242), .A2(n243), .Y(n203) );
  NAND2X0_HVT U142 ( .A1(n204), .A2(n235), .Y(n244) );
  NAND2X0_HVT U143 ( .A1(n203), .A2(n262), .Y(n245) );
  NAND2X0_HVT U144 ( .A1(n244), .A2(n245), .Y(n205) );
  MUX21X1_HVT U145 ( .A1(n269), .A2(n271), .S0(n291), .Y(n17) );
  IBUFFX2_HVT U148 ( .A(n290), .Y(n288) );
  OA21X1_HVT U149 ( .A1(n8), .A2(n297), .A3(n329), .Y(n204) );
  INVX1_HVT U150 ( .A(n247), .Y(n142) );
  MUX41X1_HVT U151 ( .A1(n331), .A3(n37), .A2(n33), .A4(n12), .S0(n292), .S1(
        n295), .Y(n206) );
  MUX41X1_HVT U152 ( .A1(n190), .A3(n193), .A2(n186), .A4(n189), .S0(n231), 
        .S1(in[0]), .Y(n194) );
  MUX21X2_HVT U155 ( .A1(n166), .A2(n178), .S0(n232), .Y(out[5]) );
  MUX41X1_HVT U156 ( .A1(n319), .A3(n332), .A2(n281), .A4(n330), .S0(n297), 
        .S1(n292), .Y(n186) );
  MUX41X1_HVT U157 ( .A1(n249), .A3(n248), .A2(n10), .A4(n227), .S0(n235), 
        .S1(n297), .Y(n247) );
  MUX21X2_HVT U161 ( .A1(n146), .A2(n154), .S0(n232), .Y(out[4]) );
  MUX41X1_HVT U163 ( .A1(n278), .A3(n348), .A2(n28), .A4(n42), .S0(n246), .S1(
        n292), .Y(n197) );
  MUX41X1_HVT U164 ( .A1(n104), .A3(n109), .A2(n108), .A4(n111), .S0(n219), 
        .S1(n231), .Y(n112) );
  MUX21X2_HVT U169 ( .A1(n112), .A2(n102), .S0(in[6]), .Y(out[2]) );
  XOR2X1_HVT U170 ( .A1(n290), .A2(n292), .Y(n50) );
  INVX0_HVT U171 ( .A(n290), .Y(n289) );
  INVX0_HVT U172 ( .A(in[3]), .Y(n354) );
  INVX1_HVT U173 ( .A(n5), .Y(n352) );
  MUX21X1_HVT U175 ( .A1(n252), .A2(n312), .S0(n260), .Y(n137) );
  NBUFFX2_HVT U176 ( .A(n23), .Y(n272) );
  NBUFFX2_HVT U180 ( .A(n23), .Y(n270) );
  AND2X1_HVT U182 ( .A1(n272), .A2(n59), .Y(n250) );
  INVX1_HVT U183 ( .A(n2), .Y(n356) );
  MUX21X1_HVT U184 ( .A1(n352), .A2(n355), .S0(n266), .Y(n55) );
  NBUFFX2_HVT U185 ( .A(n5), .Y(n280) );
  MUX21X1_HVT U187 ( .A1(n32), .A2(n115), .S0(n260), .Y(n117) );
  NBUFFX2_HVT U188 ( .A(n5), .Y(n281) );
  MUX21X1_HVT U189 ( .A1(n308), .A2(n353), .S0(n266), .Y(n70) );
  AND2X1_HVT U190 ( .A1(n282), .A2(n76), .Y(n251) );
  MUX21X1_HVT U191 ( .A1(n272), .A2(n355), .S0(n289), .Y(n8) );
  MUX21X1_HVT U192 ( .A1(n270), .A2(n275), .S0(n234), .Y(n107) );
  MUX21X1_HVT U193 ( .A1(n24), .A2(n330), .S0(n267), .Y(n144) );
  MUX21X1_HVT U194 ( .A1(n352), .A2(n356), .S0(n234), .Y(n179) );
  MUX21X1_HVT U196 ( .A1(n271), .A2(n352), .S0(n233), .Y(n99) );
  MUX21X1_HVT U198 ( .A1(n281), .A2(n7), .S0(n286), .Y(n38) );
  MUX21X1_HVT U199 ( .A1(n7), .A2(n353), .S0(n287), .Y(n227) );
  MUX21X1_HVT U200 ( .A1(n7), .A2(n356), .S0(n233), .Y(n26) );
  MUX21X1_HVT U201 ( .A1(n280), .A2(n279), .S0(n233), .Y(n92) );
  MUX21X1_HVT U202 ( .A1(n7), .A2(n275), .S0(n233), .Y(n79) );
  XOR2X1_HVT U203 ( .A1(n7), .A2(n289), .Y(n47) );
  MUX21X1_HVT U207 ( .A1(n356), .A2(n355), .S0(n289), .Y(n28) );
  MUX21X1_HVT U209 ( .A1(n355), .A2(n352), .S0(n288), .Y(n39) );
  MUX21X1_HVT U210 ( .A1(n355), .A2(n269), .S0(n288), .Y(n35) );
  MUX21X1_HVT U211 ( .A1(n269), .A2(n356), .S0(n289), .Y(n41) );
  MUX21X1_HVT U213 ( .A1(n275), .A2(n352), .S0(n289), .Y(n30) );
  MUX21X1_HVT U216 ( .A1(n124), .A2(n123), .S0(n241), .Y(n125) );
  MUX21X1_HVT U217 ( .A1(n301), .A2(n326), .S0(n260), .Y(n123) );
  MUX21X1_HVT U219 ( .A1(n323), .A2(n140), .S0(n263), .Y(n141) );
  MUX21X1_HVT U221 ( .A1(n347), .A2(n279), .S0(n268), .Y(n140) );
  NAND2X0_HVT U222 ( .A1(n273), .A2(n354), .Y(n5) );
  MUX21X1_HVT U223 ( .A1(n352), .A2(n274), .S0(n288), .Y(n226) );
  MUX21X1_HVT U224 ( .A1(n269), .A2(n7), .S0(n289), .Y(n224) );
  INVX1_HVT U225 ( .A(n10), .Y(n353) );
  INVX1_HVT U226 ( .A(n1), .Y(n355) );
  MUX21X1_HVT U227 ( .A1(n283), .A2(n278), .S0(n234), .Y(n15) );
  MUX21X1_HVT U228 ( .A1(n300), .A2(n127), .S0(n261), .Y(n128) );
  MUX21X1_HVT U229 ( .A1(n274), .A2(n269), .S0(n286), .Y(n127) );
  NBUFFX2_HVT U230 ( .A(n2), .Y(n282) );
  NBUFFX2_HVT U231 ( .A(n2), .Y(n283) );
  XOR2X1_HVT U232 ( .A1(n286), .A2(n353), .Y(n46) );
  MUX21X1_HVT U233 ( .A1(n354), .A2(n284), .S0(n287), .Y(n192) );
  MUX21X1_HVT U234 ( .A1(n1), .A2(n282), .S0(n287), .Y(n191) );
  MUX21X1_HVT U235 ( .A1(n353), .A2(n352), .S0(n234), .Y(n19) );
  MUX21X1_HVT U236 ( .A1(n281), .A2(n284), .S0(n287), .Y(n97) );
  MUX21X1_HVT U237 ( .A1(n269), .A2(n355), .S0(n288), .Y(n11) );
  MUX21X1_HVT U238 ( .A1(n280), .A2(n269), .S0(n288), .Y(n12) );
  MUX21X1_HVT U239 ( .A1(n269), .A2(n275), .S0(n286), .Y(n195) );
  XOR2X1_HVT U240 ( .A1(n283), .A2(n233), .Y(n51) );
  MUX21X1_HVT U241 ( .A1(n283), .A2(n274), .S0(n234), .Y(n220) );
  XNOR2X1_HVT U242 ( .A1(n280), .A2(n233), .Y(n252) );
  AND2X1_HVT U243 ( .A1(n289), .A2(n356), .Y(n253) );
  MUX21X1_HVT U244 ( .A1(n284), .A2(n278), .S0(n285), .Y(n32) );
  MUX21X1_HVT U245 ( .A1(n2), .A2(n280), .S0(n233), .Y(n228) );
  AND2X1_HVT U246 ( .A1(n284), .A2(n116), .Y(n254) );
  XNOR2X1_HVT U247 ( .A1(n1), .A2(n285), .Y(n255) );
  MUX21X1_HVT U248 ( .A1(n278), .A2(n269), .S0(n285), .Y(n222) );
  MUX21X1_HVT U249 ( .A1(n279), .A2(n274), .S0(n288), .Y(n74) );
  MUX21X1_HVT U250 ( .A1(n279), .A2(n284), .S0(n263), .Y(n130) );
  XOR2X1_HVT U251 ( .A1(n273), .A2(n289), .Y(n27) );
  NBUFFX2_HVT U252 ( .A(in[7]), .Y(n268) );
  NBUFFX2_HVT U253 ( .A(n354), .Y(n269) );
  NBUFFX2_HVT U254 ( .A(in[2]), .Y(n260) );
  NBUFFX2_HVT U255 ( .A(in[5]), .Y(n266) );
  NBUFFX2_HVT U256 ( .A(in[2]), .Y(n261) );
  NBUFFX2_HVT U257 ( .A(in[5]), .Y(n265) );
  NBUFFX2_HVT U258 ( .A(n261), .Y(n263) );
  NBUFFX2_HVT U259 ( .A(in[2]), .Y(n264) );
  NBUFFX2_HVT U260 ( .A(in[2]), .Y(n259) );
  MUX21X1_HVT U261 ( .A1(n105), .A2(n323), .S0(n263), .Y(n108) );
  MUX21X1_HVT U262 ( .A1(n188), .A2(n187), .S0(n262), .Y(n189) );
  MUX21X1_HVT U263 ( .A1(n89), .A2(n277), .S0(n217), .Y(n187) );
  XOR2X1_HVT U264 ( .A1(n288), .A2(n277), .Y(n49) );
  MUX21X1_HVT U265 ( .A1(n278), .A2(n272), .S0(n234), .Y(n110) );
  MUX21X1_HVT U266 ( .A1(n82), .A2(n83), .S0(n264), .Y(n85) );
  MUX21X1_HVT U267 ( .A1(n21), .A2(n279), .S0(n268), .Y(n82) );
  MUX21X1_HVT U268 ( .A1(n175), .A2(n176), .S0(n263), .Y(n177) );
  MUX21X1_HVT U269 ( .A1(n279), .A2(n342), .S0(n268), .Y(n175) );
  AND2X1_HVT U270 ( .A1(n272), .A2(n291), .Y(n256) );
  MUX21X1_HVT U271 ( .A1(n277), .A2(n352), .S0(n285), .Y(n40) );
  MUX21X1_HVT U272 ( .A1(n45), .A2(n72), .S0(n262), .Y(n73) );
  MUX21X1_HVT U273 ( .A1(n355), .A2(n342), .S0(n268), .Y(n72) );
  XOR2X1_HVT U274 ( .A1(n297), .A2(n28), .Y(n45) );
  MUX21X1_HVT U275 ( .A1(n30), .A2(n304), .S0(n268), .Y(n150) );
  MUX21X1_HVT U276 ( .A1(n18), .A2(n325), .S0(n261), .Y(n138) );
  MUX21X1_HVT U277 ( .A1(n344), .A2(n353), .S0(n295), .Y(n155) );
  MUX21X1_HVT U278 ( .A1(n353), .A2(n356), .S0(n287), .Y(n170) );
  NAND2X0_HVT U279 ( .A1(in[3]), .A2(n275), .Y(n2) );
  NBUFFX2_HVT U280 ( .A(n357), .Y(n275) );
  MUX21X1_HVT U281 ( .A1(n356), .A2(n277), .S0(n285), .Y(n20) );
  MUX21X1_HVT U282 ( .A1(n327), .A2(n3), .S0(n261), .Y(n113) );
  MUX21X1_HVT U283 ( .A1(n160), .A2(n283), .S0(n257), .Y(n161) );
  MUX21X1_HVT U284 ( .A1(n54), .A2(n53), .S0(n267), .Y(n56) );
  MUX21X1_HVT U285 ( .A1(n277), .A2(n36), .S0(n266), .Y(n53) );
  XOR2X1_HVT U286 ( .A1(n234), .A2(n265), .Y(n44) );
  MUX21X1_HVT U287 ( .A1(n3), .A2(n291), .S0(n262), .Y(n131) );
  MUX21X1_HVT U288 ( .A1(n277), .A2(n353), .S0(n234), .Y(n223) );
  MUX21X1_HVT U289 ( .A1(n31), .A2(n215), .S0(n267), .Y(n225) );
  MUX21X1_HVT U290 ( .A1(n281), .A2(n277), .S0(n289), .Y(n9) );
  MUX21X1_HVT U291 ( .A1(n310), .A2(n291), .S0(n266), .Y(n68) );
  NBUFFX2_HVT U292 ( .A(n10), .Y(n278) );
  MUX21X1_HVT U293 ( .A1(n320), .A2(n31), .S0(n261), .Y(n135) );
  MUX21X1_HVT U294 ( .A1(n283), .A2(n94), .S0(n257), .Y(n95) );
  MUX21X1_HVT U295 ( .A1(n277), .A2(n274), .S0(n268), .Y(n94) );
  NBUFFX2_HVT U296 ( .A(n1), .Y(n284) );
  NBUFFX2_HVT U297 ( .A(n213), .Y(n274) );
  NBUFFX2_HVT U298 ( .A(n10), .Y(n279) );
  XNOR2X1_HVT U299 ( .A1(n297), .A2(n286), .Y(n257) );
  AND2X1_HVT U300 ( .A1(n269), .A2(n291), .Y(n258) );
  NBUFFX2_HVT U301 ( .A(in[5]), .Y(n293) );
  MUX21X1_HVT U302 ( .A1(n199), .A2(n200), .S0(n262), .Y(n201) );
  MUX21X1_HVT U303 ( .A1(n125), .A2(n122), .S0(n266), .Y(n126) );
  MUX21X1_HVT U304 ( .A1(n96), .A2(n95), .S0(n264), .Y(n98) );
  MUX21X1_HVT U305 ( .A1(n56), .A2(n52), .S0(n263), .Y(n57) );
  MUX21X1_HVT U306 ( .A1(n62), .A2(n60), .S0(n262), .Y(n63) );
  MUX21X1_HVT U307 ( .A1(n352), .A2(n237), .S0(n287), .Y(n33) );
  NAND2X0_HVT U308 ( .A1(n216), .A2(n354), .Y(n10) );
  NAND2X0_HVT U309 ( .A1(in[3]), .A2(n216), .Y(n1) );
  MUX21X1_HVT U310 ( .A1(n237), .A2(n7), .S0(n287), .Y(n221) );
  MUX21X1_HVT U311 ( .A1(n237), .A2(n355), .S0(n286), .Y(n37) );
  MUX21X1_HVT U312 ( .A1(n237), .A2(n353), .S0(n285), .Y(n18) );
  MUX21X1_HVT U313 ( .A1(n237), .A2(n283), .S0(n285), .Y(n21) );
  MUX21X1_HVT U314 ( .A1(n237), .A2(n278), .S0(n286), .Y(n229) );
  MUX21X1_HVT U315 ( .A1(n284), .A2(n237), .S0(n233), .Y(n29) );
  MUX21X1_HVT U316 ( .A1(n277), .A2(n237), .S0(n260), .Y(n118) );
  MUX21X1_HVT U317 ( .A1(n237), .A2(n284), .S0(n286), .Y(n230) );
  MUX21X1_HVT U318 ( .A1(n269), .A2(n237), .S0(n286), .Y(n31) );
  NBUFFX2_HVT U319 ( .A(in[3]), .Y(n277) );
  NBUFFX2_HVT U320 ( .A(in[0]), .Y(n276) );
  INVX0_HVT U321 ( .A(n22), .Y(n298) );
  INVX0_HVT U322 ( .A(n25), .Y(n299) );
  INVX0_HVT U323 ( .A(n34), .Y(n300) );
  INVX0_HVT U324 ( .A(n36), .Y(n301) );
  INVX0_HVT U325 ( .A(n173), .Y(n302) );
  INVX0_HVT U326 ( .A(n214), .Y(n303) );
  INVX0_HVT U327 ( .A(n3), .Y(n304) );
  INVX0_HVT U328 ( .A(n16), .Y(n305) );
  INVX0_HVT U329 ( .A(n4), .Y(n306) );
  INVX0_HVT U330 ( .A(n8), .Y(n307) );
  INVX0_HVT U331 ( .A(n9), .Y(n308) );
  INVX0_HVT U332 ( .A(n11), .Y(n309) );
  INVX0_HVT U333 ( .A(n12), .Y(n310) );
  INVX0_HVT U334 ( .A(n15), .Y(n311) );
  INVX0_HVT U335 ( .A(n18), .Y(n313) );
  INVX0_HVT U336 ( .A(n19), .Y(n314) );
  INVX0_HVT U337 ( .A(n20), .Y(n315) );
  INVX0_HVT U338 ( .A(n21), .Y(n316) );
  INVX0_HVT U339 ( .A(n26), .Y(n318) );
  INVX0_HVT U340 ( .A(n27), .Y(n319) );
  INVX0_HVT U341 ( .A(n29), .Y(n320) );
  INVX0_HVT U342 ( .A(n30), .Y(n321) );
  INVX0_HVT U343 ( .A(n31), .Y(n322) );
  INVX0_HVT U344 ( .A(n225), .Y(n323) );
  INVX0_HVT U345 ( .A(n32), .Y(n324) );
  INVX0_HVT U346 ( .A(n33), .Y(n325) );
  INVX0_HVT U347 ( .A(n35), .Y(n326) );
  INVX0_HVT U348 ( .A(n40), .Y(n330) );
  INVX0_HVT U349 ( .A(n41), .Y(n331) );
  INVX0_HVT U350 ( .A(n42), .Y(n332) );
  INVX0_HVT U351 ( .A(n43), .Y(n333) );
  INVX0_HVT U352 ( .A(n76), .Y(n334) );
  INVX0_HVT U353 ( .A(n13), .Y(n335) );
  INVX0_HVT U354 ( .A(n116), .Y(n336) );
  INVX0_HVT U355 ( .A(n215), .Y(n337) );
  INVX0_HVT U356 ( .A(n59), .Y(n338) );
  INVX0_HVT U357 ( .A(n157), .Y(n339) );
  INVX0_HVT U358 ( .A(n220), .Y(n340) );
  INVX0_HVT U359 ( .A(n221), .Y(n341) );
  INVX0_HVT U360 ( .A(n223), .Y(n343) );
  INVX0_HVT U361 ( .A(n97), .Y(n345) );
  INVX0_HVT U362 ( .A(n107), .Y(n346) );
  INVX0_HVT U363 ( .A(n226), .Y(n347) );
  INVX0_HVT U364 ( .A(n228), .Y(n349) );
  INVX0_HVT U365 ( .A(n230), .Y(n351) );
endmodule

