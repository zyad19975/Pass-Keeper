
module sbox_8 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n19, n23, n35, n38, n50, n87, n95, n96, n98, n118, n119, n210, n211,
         n212, n213, n216, n217, n218, n219, n220, n224, n225, n231, n232,
         n236, n238, n241, n246, n261, n264, n272, n273, n274, n278, n280,
         n282, n283, n284, n289, n293, n294, n297, n300, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776;

  NAND2X0_HVT U4 ( .A1(n391), .A2(n774), .Y(n773) );
  NAND2X0_HVT U5 ( .A1(n410), .A2(n502), .Y(n771) );
  NAND2X0_HVT U13 ( .A1(n763), .A2(n374), .Y(n764) );
  NAND2X0_HVT U21 ( .A1(n393), .A2(n509), .Y(n756) );
  NAND2X0_HVT U24 ( .A1(n398), .A2(n447), .Y(n754) );
  NAND2X0_HVT U33 ( .A1(n297), .A2(n509), .Y(n745) );
  NAND2X0_HVT U42 ( .A1(n356), .A2(n497), .Y(n738) );
  MUX41X1_HVT U51 ( .A1(n213), .A3(n545), .A2(n519), .A4(n525), .S0(n493), 
        .S1(n492), .Y(n730) );
  NAND2X0_HVT U53 ( .A1(n727), .A2(n737), .Y(n728) );
  NAND2X0_HVT U56 ( .A1(n392), .A2(n723), .Y(n724) );
  NAND2X0_HVT U58 ( .A1(n374), .A2(n774), .Y(n721) );
  MUX41X1_HVT U61 ( .A1(n481), .A3(n556), .A2(n530), .A4(n498), .S0(n349), 
        .S1(n492), .Y(n718) );
  NAND2X0_HVT U62 ( .A1(n447), .A2(n504), .Y(n717) );
  AO21X1_HVT U66 ( .A1(n562), .A2(n513), .A3(n564), .Y(n713) );
  NAND2X0_HVT U73 ( .A1(n272), .A2(n330), .Y(n707) );
  MUX41X1_HVT U74 ( .A1(n708), .A3(n752), .A2(n707), .A4(n754), .S0(n490), 
        .S1(n515), .Y(n705) );
  NAND2X0_HVT U85 ( .A1(n509), .A2(n563), .Y(n694) );
  MUX41X1_HVT U86 ( .A1(n558), .A3(n694), .A2(n482), .A4(n478), .S0(n433), 
        .S1(n515), .Y(n693) );
  MUX41X1_HVT U96 ( .A1(n568), .A3(n480), .A2(n559), .A4(n687), .S0(n433), 
        .S1(n516), .Y(n686) );
  NAND2X0_HVT U101 ( .A1(n680), .A2(n679), .Y(n681) );
  NAND2X0_HVT U110 ( .A1(n504), .A2(n670), .Y(n671) );
  AND2X1_HVT U115 ( .A1(n396), .A2(n498), .Y(n667) );
  MUX41X1_HVT U116 ( .A1(n470), .A3(n667), .A2(n472), .A4(n747), .S0(n377), 
        .S1(n349), .Y(n666) );
  NAND2X0_HVT U123 ( .A1(n658), .A2(n657), .Y(n659) );
  MUX41X1_HVT U125 ( .A1(n756), .A3(n485), .A2(n529), .A4(n540), .S0(n377), 
        .S1(n493), .Y(n655) );
  MUX41X1_HVT U136 ( .A1(n478), .A3(n745), .A2(n523), .A4(n743), .S0(n377), 
        .S1(n349), .Y(n645) );
  AND2X1_HVT U140 ( .A1(n430), .A2(n316), .Y(n641) );
  NAND2X0_HVT U146 ( .A1(n218), .A2(n373), .Y(n706) );
  AND2X1_HVT U154 ( .A1(n495), .A2(n398), .Y(n628) );
  NAND2X0_HVT U158 ( .A1(n395), .A2(n563), .Y(n624) );
  MUX41X1_HVT U159 ( .A1(n470), .A3(n498), .A2(n624), .A4(n565), .S0(n313), 
        .S1(n431), .Y(n623) );
  AND2X1_HVT U162 ( .A1(n706), .A2(n346), .Y(n620) );
  NAND2X0_HVT U166 ( .A1(n374), .A2(n723), .Y(n616) );
  NAND2X0_HVT U167 ( .A1(n371), .A2(n509), .Y(n615) );
  MUX41X1_HVT U168 ( .A1(n533), .A3(n430), .A2(n615), .A4(n616), .S0(n362), 
        .S1(n476), .Y(n614) );
  NAND2X0_HVT U174 ( .A1(n403), .A2(n220), .Y(n763) );
  MUX41X1_HVT U176 ( .A1(n212), .A3(n609), .A2(n531), .A4(n763), .S0(n304), 
        .S1(n453), .Y(n608) );
  NAND2X0_HVT U177 ( .A1(n507), .A2(n212), .Y(n607) );
  MUX41X1_HVT U179 ( .A1(n750), .A3(n551), .A2(n534), .A4(n552), .S0(n458), 
        .S1(n494), .Y(n605) );
  MUX41X1_HVT U180 ( .A1(n528), .A3(n768), .A2(n470), .A4(n23), .S0(n493), 
        .S1(n362), .Y(n604) );
  MUX41X1_HVT U182 ( .A1(n539), .A3(n772), .A2(n524), .A4(n548), .S0(n514), 
        .S1(n458), .Y(n602) );
  MUX41X1_HVT U189 ( .A1(n596), .A3(n763), .A2(n597), .A4(n544), .S0(n493), 
        .S1(n362), .Y(n595) );
  MUX41X1_HVT U190 ( .A1(n595), .A3(n598), .A2(n599), .A4(n602), .S0(n513), 
        .S1(n496), .Y(n594) );
  AO21X1_HVT U197 ( .A1(n482), .A2(n494), .A3(n557), .Y(n588) );
  NAND2X0_HVT U208 ( .A1(n440), .A2(n393), .Y(n670) );
  NAND2X0_HVT U212 ( .A1(n506), .A2(n321), .Y(n723) );
  NAND2X0_HVT U214 ( .A1(n381), .A2(n447), .Y(n578) );
  NAND2X0_HVT U215 ( .A1(n670), .A2(n272), .Y(n577) );
  NAND2X0_HVT U218 ( .A1(n428), .A2(n507), .Y(n631) );
  NAND2X0_HVT U220 ( .A1(n494), .A2(n578), .Y(n698) );
  INVX0_HVT U241 ( .A(n754), .Y(n568) );
  INVX0_HVT U245 ( .A(n771), .Y(n565) );
  INVX0_HVT U247 ( .A(n706), .Y(n564) );
  INVX0_HVT U250 ( .A(n766), .Y(n562) );
  INVX0_HVT U256 ( .A(n631), .Y(n557) );
  INVX0_HVT U260 ( .A(n743), .Y(n553) );
  INVX0_HVT U264 ( .A(n744), .Y(n549) );
  INVX0_HVT U265 ( .A(n752), .Y(n548) );
  INVX0_HVT U268 ( .A(n756), .Y(n545) );
  INVX0_HVT U270 ( .A(n577), .Y(n544) );
  INVX0_HVT U276 ( .A(n741), .Y(n539) );
  INVX0_HVT U278 ( .A(n745), .Y(n537) );
  INVX0_HVT U284 ( .A(n578), .Y(n534) );
  INVX0_HVT U289 ( .A(n679), .Y(n531) );
  INVX0_HVT U295 ( .A(n773), .Y(n528) );
  INVX0_HVT U296 ( .A(n761), .Y(n527) );
  INVX0_HVT U298 ( .A(n762), .Y(n526) );
  INVX0_HVT U306 ( .A(n615), .Y(n521) );
  INVX0_HVT U309 ( .A(n758), .Y(n519) );
  AOI21X1_HVT U1 ( .A1(n495), .A2(n688), .A3(n557), .Y(n402) );
  INVX1_HVT U2 ( .A(n372), .Y(n374) );
  NBUFFX2_HVT U3 ( .A(n566), .Y(n502) );
  INVX1_HVT U6 ( .A(n776), .Y(n475) );
  MUX21X1_HVT U7 ( .A1(n547), .A2(n428), .S0(n513), .Y(n712) );
  MUX21X1_HVT U8 ( .A1(n655), .A2(n656), .S0(n492), .Y(n654) );
  INVX0_HVT U9 ( .A(n518), .Y(n514) );
  INVX1_HVT U10 ( .A(n518), .Y(n304) );
  INVX0_HVT U11 ( .A(n490), .Y(n317) );
  INVX1_HVT U12 ( .A(n490), .Y(n35) );
  AND2X1_HVT U14 ( .A1(n334), .A2(n335), .Y(n19) );
  INVX1_HVT U15 ( .A(n541), .Y(n393) );
  AND2X1_HVT U16 ( .A1(n498), .A2(n723), .Y(n23) );
  INVX0_HVT U17 ( .A(n768), .Y(n547) );
  NAND2X0_HVT U18 ( .A1(n119), .A2(n35), .Y(n38) );
  NAND2X0_HVT U19 ( .A1(n648), .A2(n490), .Y(n50) );
  NAND2X0_HVT U20 ( .A1(n38), .A2(n50), .Y(n647) );
  MUX21X1_HVT U22 ( .A1(n430), .A2(n540), .S0(n427), .Y(n648) );
  XOR2X2_HVT U23 ( .A1(n499), .A2(n356), .Y(n752) );
  INVX1_HVT U25 ( .A(n770), .Y(n418) );
  MUX41X1_HVT U26 ( .A1(n118), .A3(n703), .A2(n542), .A4(n768), .S0(n350), 
        .S1(n35), .Y(n702) );
  NAND2X0_HVT U27 ( .A1(n391), .A2(n473), .Y(n87) );
  NAND2X0_HVT U28 ( .A1(n497), .A2(n506), .Y(n95) );
  NAND2X0_HVT U29 ( .A1(n87), .A2(n95), .Y(n768) );
  NAND2X0_HVT U30 ( .A1(n555), .A2(n284), .Y(n96) );
  NAND2X0_HVT U31 ( .A1(n748), .A2(n488), .Y(n98) );
  NAND2X0_HVT U32 ( .A1(n96), .A2(n98), .Y(n653) );
  MUX21X1_HVT U34 ( .A1(n469), .A2(n312), .S0(n352), .Y(n748) );
  INVX1_HVT U35 ( .A(n508), .Y(n410) );
  NBUFFX2_HVT U36 ( .A(n385), .Y(n505) );
  NBUFFX2_HVT U37 ( .A(n385), .Y(n504) );
  MUX21X2_HVT U38 ( .A1(n505), .A2(n767), .S0(n403), .Y(n762) );
  MUX21X1_HVT U39 ( .A1(n392), .A2(n374), .S0(n432), .Y(n688) );
  MUX21X1_HVT U40 ( .A1(n394), .A2(n549), .S0(n317), .Y(n665) );
  INVX1_HVT U41 ( .A(n511), .Y(n510) );
  INVX1_HVT U43 ( .A(n518), .Y(n515) );
  INVX1_HVT U44 ( .A(n738), .Y(n567) );
  XOR2X1_HVT U45 ( .A1(n280), .A2(n512), .Y(n737) );
  INVX1_HVT U46 ( .A(n493), .Y(n216) );
  INVX1_HVT U47 ( .A(n494), .Y(n427) );
  XOR2X1_HVT U48 ( .A1(n488), .A2(n495), .Y(n733) );
  INVX1_HVT U49 ( .A(n750), .Y(n555) );
  INVX1_HVT U50 ( .A(n488), .Y(n415) );
  INVX1_HVT U52 ( .A(n445), .Y(n749) );
  OA21X1_HVT U54 ( .A1(n521), .A2(n309), .A3(n337), .Y(n637) );
  NAND2X0_HVT U55 ( .A1(n542), .A2(n304), .Y(n375) );
  OA21X1_HVT U57 ( .A1(n483), .A2(n309), .A3(n747), .Y(n612) );
  XNOR2X1_HVT U59 ( .A1(n392), .A2(n432), .Y(n479) );
  INVX1_HVT U60 ( .A(n384), .Y(n385) );
  INVX1_HVT U63 ( .A(n323), .Y(n356) );
  NAND2X0_HVT U64 ( .A1(n23), .A2(n304), .Y(n344) );
  INVX1_HVT U65 ( .A(n493), .Y(n224) );
  NAND2X0_HVT U67 ( .A1(n664), .A2(n224), .Y(n451) );
  INVX1_HVT U68 ( .A(n670), .Y(n543) );
  XNOR2X1_HVT U69 ( .A1(n411), .A2(n356), .Y(n734) );
  INVX1_HVT U70 ( .A(n518), .Y(n516) );
  NBUFFX2_HVT U71 ( .A(in[5]), .Y(n513) );
  INVX1_HVT U72 ( .A(n518), .Y(n476) );
  MUX21X1_HVT U75 ( .A1(n499), .A2(n220), .S0(n390), .Y(n703) );
  NBUFFX2_HVT U76 ( .A(n510), .Y(n488) );
  NBUFFX2_HVT U77 ( .A(n514), .Y(n493) );
  INVX1_HVT U78 ( .A(n515), .Y(n336) );
  INVX1_HVT U79 ( .A(n323), .Y(n507) );
  INVX1_HVT U80 ( .A(n323), .Y(n396) );
  INVX1_HVT U81 ( .A(n323), .Y(n218) );
  INVX0_HVT U82 ( .A(n506), .Y(n316) );
  INVX1_HVT U83 ( .A(n489), .Y(n284) );
  INVX1_HVT U84 ( .A(n513), .Y(n387) );
  INVX1_HVT U87 ( .A(n514), .Y(n486) );
  INVX1_HVT U88 ( .A(n429), .Y(n342) );
  NBUFFX2_HVT U89 ( .A(n514), .Y(n495) );
  INVX1_HVT U90 ( .A(n304), .Y(n517) );
  NBUFFX2_HVT U91 ( .A(in[0]), .Y(n496) );
  INVX1_HVT U92 ( .A(n772), .Y(n541) );
  INVX0_HVT U93 ( .A(n391), .Y(n389) );
  INVX1_HVT U94 ( .A(n760), .Y(n530) );
  AND2X1_HVT U95 ( .A1(n319), .A2(n320), .Y(n118) );
  AND2X1_HVT U97 ( .A1(n365), .A2(n366), .Y(n119) );
  INVX1_HVT U98 ( .A(n380), .Y(n381) );
  AND2X1_HVT U99 ( .A1(n436), .A2(n437), .Y(n210) );
  AND2X1_HVT U100 ( .A1(n433), .A2(n400), .Y(n211) );
  INVX1_HVT U102 ( .A(n776), .Y(n372) );
  INVX1_HVT U103 ( .A(n500), .Y(n446) );
  MUX21X1_HVT U104 ( .A1(n393), .A2(n767), .S0(n322), .Y(n691) );
  INVX1_HVT U105 ( .A(n322), .Y(n323) );
  INVX1_HVT U106 ( .A(n397), .Y(n212) );
  AND2X1_HVT U107 ( .A1(n305), .A2(n306), .Y(n213) );
  MUX41X1_HVT U108 ( .A1(n527), .A3(n717), .A2(n526), .A4(n535), .S0(n216), 
        .S1(n492), .Y(n716) );
  INVX0_HVT U109 ( .A(n508), .Y(n395) );
  INVX1_HVT U111 ( .A(n550), .Y(n318) );
  INVX1_HVT U112 ( .A(n499), .Y(n397) );
  INVX0_HVT U113 ( .A(n440), .Y(n352) );
  INVX1_HVT U114 ( .A(n541), .Y(n391) );
  INVX0_HVT U117 ( .A(n323), .Y(n217) );
  INVX0_HVT U118 ( .A(n776), .Y(n563) );
  MUX21X1_HVT U119 ( .A1(n502), .A2(n371), .S0(n217), .Y(n740) );
  INVX1_HVT U120 ( .A(n522), .Y(n219) );
  INVX1_HVT U121 ( .A(n503), .Y(n522) );
  MUX21X1_HVT U122 ( .A1(n219), .A2(n418), .S0(n473), .Y(n472) );
  INVX0_HVT U124 ( .A(n477), .Y(n220) );
  INVX0_HVT U126 ( .A(n477), .Y(n770) );
  MUX21X1_HVT U127 ( .A1(n393), .A2(n219), .S0(n289), .Y(n571) );
  MUX41X1_HVT U128 ( .A1(n721), .A3(n485), .A2(n438), .A4(n483), .S0(n224), 
        .S1(n492), .Y(n720) );
  INVX1_HVT U129 ( .A(n356), .Y(n447) );
  INVX1_HVT U130 ( .A(n440), .Y(n390) );
  INVX1_HVT U131 ( .A(n372), .Y(n373) );
  INVX1_HVT U132 ( .A(n486), .Y(n349) );
  INVX0_HVT U133 ( .A(n742), .Y(n538) );
  INVX1_HVT U134 ( .A(n571), .Y(n523) );
  MUX21X2_HVT U135 ( .A1(n736), .A2(n710), .S0(n488), .Y(n709) );
  NAND2X0_HVT U137 ( .A1(n632), .A2(n412), .Y(n347) );
  MUX41X1_HVT U138 ( .A1(n210), .A3(n669), .A2(n673), .A4(n672), .S0(n516), 
        .S1(n491), .Y(n668) );
  INVX1_HVT U139 ( .A(n318), .Y(n307) );
  NBUFFX2_HVT U141 ( .A(n322), .Y(n432) );
  INVX0_HVT U142 ( .A(n769), .Y(n529) );
  INVX1_HVT U143 ( .A(n390), .Y(n280) );
  MUX41X1_HVT U144 ( .A1(n529), .A3(n713), .A2(n712), .A4(n714), .S0(n362), 
        .S1(n431), .Y(n711) );
  NAND2X0_HVT U145 ( .A1(n469), .A2(n352), .Y(n225) );
  NAND2X0_HVT U147 ( .A1(n475), .A2(n218), .Y(n231) );
  NAND2X0_HVT U148 ( .A1(n225), .A2(n231), .Y(n743) );
  INVX0_HVT U149 ( .A(n566), .Y(n361) );
  INVX1_HVT U150 ( .A(n740), .Y(n520) );
  MUX41X1_HVT U151 ( .A1(n591), .A3(n587), .A2(n592), .A4(n590), .S0(n368), 
        .S1(n512), .Y(n586) );
  NAND2X0_HVT U152 ( .A1(n303), .A2(n302), .Y(n232) );
  INVX0_HVT U153 ( .A(n278), .Y(n767) );
  NAND2X0_HVT U155 ( .A1(n728), .A2(n224), .Y(n236) );
  NAND2X0_HVT U156 ( .A1(n729), .A2(n493), .Y(n238) );
  NAND2X0_HVT U157 ( .A1(n236), .A2(n238), .Y(n726) );
  NAND2X0_HVT U160 ( .A1(n393), .A2(n509), .Y(n241) );
  NAND2X0_HVT U161 ( .A1(n502), .A2(n395), .Y(n246) );
  NAND2X0_HVT U163 ( .A1(n241), .A2(n246), .Y(n765) );
  NAND2X0_HVT U164 ( .A1(n505), .A2(n507), .Y(n261) );
  NAND2X0_HVT U165 ( .A1(n469), .A2(n352), .Y(n264) );
  NAND2X0_HVT U169 ( .A1(n261), .A2(n264), .Y(n757) );
  INVX0_HVT U170 ( .A(n757), .Y(n525) );
  XOR2X1_HVT U171 ( .A1(n217), .A2(n511), .Y(n487) );
  INVX1_HVT U172 ( .A(n220), .Y(n380) );
  INVX1_HVT U173 ( .A(n411), .Y(n346) );
  INVX0_HVT U175 ( .A(n429), .Y(n272) );
  INVX1_HVT U178 ( .A(n429), .Y(n430) );
  INVX0_HVT U181 ( .A(n321), .Y(n429) );
  INVX0_HVT U183 ( .A(n342), .Y(n428) );
  INVX0_HVT U184 ( .A(in[1]), .Y(n439) );
  XOR2X1_HVT U185 ( .A1(n503), .A2(n440), .Y(n731) );
  MUX21X1_HVT U186 ( .A1(n278), .A2(n371), .S0(n506), .Y(n618) );
  XOR2X1_HVT U187 ( .A1(n410), .A2(n278), .Y(n735) );
  INVX0_HVT U188 ( .A(n748), .Y(n554) );
  INVX0_HVT U191 ( .A(n343), .Y(n394) );
  NAND2X0_HVT U192 ( .A1(n428), .A2(n514), .Y(n273) );
  NAND2X0_HVT U193 ( .A1(n118), .A2(n427), .Y(n274) );
  NAND2X0_HVT U194 ( .A1(n273), .A2(n274), .Y(n633) );
  AND2X1_HVT U195 ( .A1(n446), .A2(n501), .Y(n278) );
  INVX0_HVT U196 ( .A(n765), .Y(n546) );
  INVX1_HVT U198 ( .A(n770), .Y(n411) );
  INVX1_HVT U199 ( .A(n576), .Y(n533) );
  NAND2X0_HVT U200 ( .A1(n418), .A2(n280), .Y(n282) );
  NAND2X0_HVT U201 ( .A1(n389), .A2(n390), .Y(n283) );
  NAND2X0_HVT U202 ( .A1(n282), .A2(n283), .Y(n388) );
  AND3X1_HVT U203 ( .A1(n510), .A2(n447), .A3(n397), .Y(n652) );
  MUX21X1_HVT U204 ( .A1(n699), .A2(n700), .S0(n317), .Y(n697) );
  AND3X1_HVT U205 ( .A1(n504), .A2(n723), .A3(n698), .Y(n699) );
  MUX41X1_HVT U206 ( .A1(n558), .A3(n560), .A2(n472), .A4(n371), .S0(n284), 
        .S1(n515), .Y(n704) );
  INVX1_HVT U207 ( .A(n759), .Y(n556) );
  INVX0_HVT U209 ( .A(n472), .Y(n753) );
  MUX41X1_HVT U210 ( .A1(n556), .A3(n620), .A2(n479), .A4(n621), .S0(n458), 
        .S1(n516), .Y(n619) );
  MUX41X1_HVT U211 ( .A1(n704), .A3(n702), .A2(n709), .A4(n705), .S0(n441), 
        .S1(n496), .Y(n701) );
  OA21X1_HVT U213 ( .A1(n343), .A2(n309), .A3(n308), .Y(n600) );
  NAND2X0_HVT U216 ( .A1(n505), .A2(n289), .Y(n293) );
  NAND2X0_HVT U217 ( .A1(n232), .A2(n410), .Y(n294) );
  NAND2X0_HVT U219 ( .A1(n293), .A2(n294), .Y(n739) );
  INVX0_HVT U221 ( .A(n395), .Y(n289) );
  INVX1_HVT U222 ( .A(n739), .Y(n524) );
  MUX21X2_HVT U223 ( .A1(n475), .A2(n559), .S0(n495), .Y(n710) );
  AND2X1_HVT U224 ( .A1(n501), .A2(n500), .Y(n297) );
  NAND2X0_HVT U225 ( .A1(n500), .A2(n361), .Y(n302) );
  NAND2X0_HVT U226 ( .A1(n318), .A2(n300), .Y(n303) );
  NAND2X0_HVT U227 ( .A1(n302), .A2(n303), .Y(n477) );
  INVX0_HVT U228 ( .A(n324), .Y(n300) );
  INVX1_HVT U229 ( .A(n471), .Y(n473) );
  MUX21X1_HVT U230 ( .A1(n446), .A2(n393), .S0(n471), .Y(n445) );
  MUX41X1_HVT U231 ( .A1(n618), .A3(n734), .A2(n554), .A4(n756), .S0(n224), 
        .S1(n35), .Y(n617) );
  INVX0_HVT U232 ( .A(n307), .Y(n469) );
  NAND2X0_HVT U233 ( .A1(n219), .A2(n289), .Y(n305) );
  NAND2X0_HVT U234 ( .A1(n499), .A2(n403), .Y(n306) );
  MUX41X1_HVT U235 ( .A1(n430), .A3(n532), .A2(n751), .A4(n739), .S0(n216), 
        .S1(n35), .Y(n591) );
  MUX21X1_HVT U236 ( .A1(n522), .A2(n563), .S0(n410), .Y(n751) );
  INVX1_HVT U237 ( .A(in[7]), .Y(n518) );
  MUX21X1_HVT U238 ( .A1(n499), .A2(n502), .S0(n390), .Y(n593) );
  NAND2X0_HVT U239 ( .A1(n363), .A2(n364), .Y(n678) );
  MUX41X1_HVT U240 ( .A1(n744), .A3(n738), .A2(n593), .A4(n731), .S0(n367), 
        .S1(n516), .Y(n592) );
  INVX1_HVT U242 ( .A(n367), .Y(n362) );
  AND2X1_HVT U243 ( .A1(n404), .A2(n358), .Y(n308) );
  INVX1_HVT U244 ( .A(n331), .Y(n438) );
  MUX41X1_HVT U246 ( .A1(n744), .A3(n445), .A2(n547), .A4(n774), .S0(n412), 
        .S1(n336), .Y(n677) );
  INVX1_HVT U248 ( .A(n473), .Y(n403) );
  NBUFFX2_HVT U249 ( .A(n517), .Y(n309) );
  NAND2X0_HVT U251 ( .A1(n613), .A2(n284), .Y(n310) );
  NAND2X0_HVT U252 ( .A1(n612), .A2(n453), .Y(n311) );
  NAND2X0_HVT U253 ( .A1(n310), .A2(n311), .Y(n611) );
  MUX21X1_HVT U254 ( .A1(n272), .A2(n559), .S0(n495), .Y(n613) );
  OR2X1_HVT U255 ( .A1(n397), .A2(n410), .Y(n744) );
  XOR2X2_HVT U257 ( .A1(n751), .A2(n517), .Y(n736) );
  NBUFFX2_HVT U258 ( .A(n300), .Y(n312) );
  NBUFFX2_HVT U259 ( .A(n566), .Y(n501) );
  INVX0_HVT U261 ( .A(n502), .Y(n398) );
  NAND2X0_HVT U262 ( .A1(n536), .A2(n313), .Y(n314) );
  NAND2X0_HVT U263 ( .A1(n415), .A2(n759), .Y(n315) );
  NAND2X0_HVT U266 ( .A1(n314), .A2(n315), .Y(n650) );
  INVX0_HVT U267 ( .A(n415), .Y(n313) );
  INVX0_HVT U269 ( .A(n746), .Y(n536) );
  INVX1_HVT U271 ( .A(n517), .Y(n431) );
  AO21X1_HVT U272 ( .A1(n316), .A2(n428), .A3(n517), .Y(n680) );
  INVX0_HVT U273 ( .A(n508), .Y(n506) );
  MUX21X1_HVT U274 ( .A1(n469), .A2(n278), .S0(n396), .Y(n759) );
  INVX1_HVT U275 ( .A(n688), .Y(n542) );
  NBUFFX2_HVT U277 ( .A(n510), .Y(n489) );
  INVX1_HVT U279 ( .A(n367), .Y(n453) );
  OA21X1_HVT U280 ( .A1(n309), .A2(n740), .A3(n631), .Y(n632) );
  INVX1_HVT U281 ( .A(in[3]), .Y(n566) );
  INVX1_HVT U282 ( .A(n508), .Y(n440) );
  NAND2X0_HVT U283 ( .A1(n502), .A2(n316), .Y(n319) );
  NAND2X0_HVT U285 ( .A1(n381), .A2(n396), .Y(n320) );
  MUX41X1_HVT U286 ( .A1(n481), .A3(n671), .A2(n549), .A4(n219), .S0(n448), 
        .S1(n515), .Y(n629) );
  NAND2X0_HVT U287 ( .A1(n446), .A2(n501), .Y(n321) );
  MUX41X1_HVT U288 ( .A1(n611), .A3(n614), .A2(n617), .A4(n619), .S0(n491), 
        .S1(n496), .Y(n610) );
  INVX1_HVT U290 ( .A(n439), .Y(n322) );
  INVX0_HVT U291 ( .A(in[1]), .Y(n508) );
  INVX0_HVT U292 ( .A(n747), .Y(n561) );
  INVX0_HVT U293 ( .A(n566), .Y(n324) );
  NAND2X0_HVT U294 ( .A1(n563), .A2(n289), .Y(n325) );
  NAND2X0_HVT U297 ( .A1(n380), .A2(n471), .Y(n326) );
  NAND2X0_HVT U299 ( .A1(n325), .A2(n326), .Y(n621) );
  INVX1_HVT U300 ( .A(n351), .Y(n327) );
  NAND2X0_HVT U301 ( .A1(n684), .A2(n327), .Y(n328) );
  NAND2X0_HVT U302 ( .A1(n674), .A2(n351), .Y(n329) );
  NAND2X0_HVT U303 ( .A1(n328), .A2(n329), .Y(out[2]) );
  INVX1_HVT U304 ( .A(in[6]), .Y(n351) );
  MUX41X1_HVT U305 ( .A1(n213), .A3(n691), .A2(n734), .A4(n738), .S0(n453), 
        .S1(n350), .Y(n690) );
  INVX1_HVT U307 ( .A(n564), .Y(n330) );
  MUX41X1_HVT U308 ( .A1(n544), .A3(n676), .A2(n732), .A4(n555), .S0(n412), 
        .S1(n350), .Y(n675) );
  INVX1_HVT U310 ( .A(n448), .Y(n433) );
  MUX21X1_HVT U311 ( .A1(n429), .A2(n389), .S0(n218), .Y(n331) );
  MUX41X1_HVT U312 ( .A1(n647), .A3(n646), .A2(n645), .A4(n643), .S0(n441), 
        .S1(n368), .Y(n642) );
  INVX1_HVT U313 ( .A(in[0]), .Y(n368) );
  NAND2X0_HVT U314 ( .A1(n272), .A2(n316), .Y(n332) );
  NAND2X0_HVT U315 ( .A1(n418), .A2(n217), .Y(n333) );
  NAND2X0_HVT U316 ( .A1(n332), .A2(n333), .Y(n676) );
  MUX41X1_HVT U317 ( .A1(n719), .A3(n711), .A2(n725), .A4(n715), .S0(n351), 
        .S1(n496), .Y(out[0]) );
  MUX41X1_HVT U318 ( .A1(n774), .A3(n397), .A2(n561), .A4(n551), .S0(n415), 
        .S1(n431), .Y(n580) );
  MUX21X2_HVT U319 ( .A1(n726), .A2(n730), .S0(n490), .Y(n725) );
  NAND2X0_HVT U320 ( .A1(n211), .A2(n401), .Y(n334) );
  NAND2X0_HVT U321 ( .A1(n402), .A2(n284), .Y(n335) );
  INVX0_HVT U322 ( .A(n561), .Y(n337) );
  MUX21X1_HVT U323 ( .A1(n600), .A2(n601), .S0(n489), .Y(n599) );
  MUX21X1_HVT U324 ( .A1(n372), .A2(n312), .S0(n440), .Y(n343) );
  NAND2X0_HVT U325 ( .A1(n638), .A2(n284), .Y(n338) );
  NAND2X0_HVT U326 ( .A1(n637), .A2(n489), .Y(n339) );
  NAND2X0_HVT U327 ( .A1(n338), .A2(n339), .Y(n636) );
  MUX21X1_HVT U328 ( .A1(n405), .A2(n749), .S0(n336), .Y(n638) );
  MUX21X1_HVT U329 ( .A1(n297), .A2(n469), .S0(n432), .Y(n746) );
  NAND2X0_HVT U330 ( .A1(n589), .A2(n415), .Y(n340) );
  NAND2X0_HVT U331 ( .A1(n588), .A2(n453), .Y(n341) );
  NAND2X0_HVT U332 ( .A1(n340), .A2(n341), .Y(n587) );
  INVX1_HVT U333 ( .A(in[4]), .Y(n550) );
  OR2X1_HVT U334 ( .A1(n381), .A2(n405), .Y(n761) );
  INVX1_HVT U335 ( .A(n405), .Y(n774) );
  OA21X1_HVT U336 ( .A1(n388), .A2(n448), .A3(n438), .Y(n672) );
  INVX1_HVT U337 ( .A(in[2]), .Y(n511) );
  NAND2X0_HVT U338 ( .A1(n760), .A2(n350), .Y(n345) );
  NAND2X0_HVT U339 ( .A1(n344), .A2(n345), .Y(n585) );
  MUX21X1_HVT U340 ( .A1(n232), .A2(n312), .S0(n471), .Y(n760) );
  NAND2X0_HVT U341 ( .A1(n633), .A2(n489), .Y(n348) );
  NAND2X0_HVT U342 ( .A1(n347), .A2(n348), .Y(n630) );
  INVX1_HVT U343 ( .A(n516), .Y(n350) );
  NBUFFX2_HVT U344 ( .A(n514), .Y(n494) );
  NBUFFX2_HVT U345 ( .A(n380), .Y(n498) );
  INVX0_HVT U346 ( .A(n723), .Y(n560) );
  MUX41X1_HVT U347 ( .A1(n677), .A3(n682), .A2(n675), .A4(n678), .S0(n496), 
        .S1(n441), .Y(n674) );
  NAND2X0_HVT U348 ( .A1(n767), .A2(n352), .Y(n353) );
  NAND2X0_HVT U349 ( .A1(n353), .A2(n246), .Y(n575) );
  NBUFFX2_HVT U350 ( .A(n550), .Y(n499) );
  INVX1_HVT U351 ( .A(n574), .Y(n558) );
  NAND2X0_HVT U352 ( .A1(n603), .A2(n327), .Y(n354) );
  NAND2X0_HVT U353 ( .A1(n594), .A2(n351), .Y(n355) );
  NAND2X0_HVT U354 ( .A1(n354), .A2(n355), .Y(out[6]) );
  NAND2X0_HVT U355 ( .A1(n297), .A2(n356), .Y(n357) );
  NAND2X0_HVT U356 ( .A1(n352), .A2(n232), .Y(n358) );
  NAND2X0_HVT U357 ( .A1(n357), .A2(n358), .Y(n687) );
  NBUFFX2_HVT U358 ( .A(n510), .Y(n490) );
  NAND2X0_HVT U359 ( .A1(n212), .A2(n396), .Y(n359) );
  NAND2X0_HVT U360 ( .A1(n498), .A2(n316), .Y(n360) );
  NAND2X0_HVT U361 ( .A1(n359), .A2(n360), .Y(n679) );
  MUX21X1_HVT U362 ( .A1(n479), .A2(n530), .S0(n488), .Y(n651) );
  MUX41X1_HVT U363 ( .A1(n520), .A3(n743), .A2(n746), .A4(n765), .S0(n412), 
        .S1(n476), .Y(n582) );
  NAND2X0_HVT U364 ( .A1(n119), .A2(n362), .Y(n363) );
  NAND2X0_HVT U365 ( .A1(n681), .A2(n367), .Y(n364) );
  NAND2X0_HVT U366 ( .A1(n748), .A2(n336), .Y(n365) );
  NAND2X0_HVT U367 ( .A1(n577), .A2(n493), .Y(n366) );
  INVX1_HVT U368 ( .A(n489), .Y(n367) );
  INVX0_HVT U369 ( .A(n575), .Y(n559) );
  MUX41X1_HVT U370 ( .A1(n480), .A3(n741), .A2(n330), .A4(n734), .S0(n377), 
        .S1(n516), .Y(n598) );
  INVX1_HVT U371 ( .A(n439), .Y(n471) );
  MUX21X2_HVT U372 ( .A1(n373), .A2(n321), .S0(n432), .Y(n747) );
  NAND2X0_HVT U373 ( .A1(n448), .A2(n561), .Y(n369) );
  NAND2X0_HVT U374 ( .A1(n762), .A2(n433), .Y(n370) );
  NAND2X0_HVT U375 ( .A1(n369), .A2(n370), .Y(n683) );
  INVX1_HVT U376 ( .A(n385), .Y(n371) );
  MUX41X1_HVT U377 ( .A1(n654), .A3(n649), .A2(n668), .A4(n662), .S0(n368), 
        .S1(n327), .Y(out[3]) );
  NAND2X0_HVT U378 ( .A1(n742), .A2(n224), .Y(n376) );
  NAND2X0_HVT U379 ( .A1(n375), .A2(n376), .Y(n626) );
  NAND2X0_HVT U380 ( .A1(n627), .A2(n377), .Y(n378) );
  NAND2X0_HVT U381 ( .A1(n626), .A2(n284), .Y(n379) );
  NAND2X0_HVT U382 ( .A1(n378), .A2(n379), .Y(n625) );
  INVX0_HVT U383 ( .A(n317), .Y(n377) );
  NBUFFX2_HVT U384 ( .A(n550), .Y(n500) );
  NAND2X0_HVT U385 ( .A1(n447), .A2(n491), .Y(n382) );
  NAND2X0_HVT U386 ( .A1(n546), .A2(n387), .Y(n383) );
  NAND2X0_HVT U387 ( .A1(n382), .A2(n383), .Y(n714) );
  INVX0_HVT U388 ( .A(n775), .Y(n384) );
  INVX1_HVT U389 ( .A(n488), .Y(n412) );
  NAND2X0_HVT U390 ( .A1(n416), .A2(n386), .Y(n437) );
  AND2X1_HVT U391 ( .A1(n417), .A2(n487), .Y(n386) );
  NAND2X0_HVT U392 ( .A1(n610), .A2(n351), .Y(n419) );
  INVX1_HVT U393 ( .A(n474), .Y(n590) );
  MUX41X1_HVT U394 ( .A1(n582), .A3(n583), .A2(n580), .A4(n581), .S0(n512), 
        .S1(n368), .Y(n579) );
  MUX21X1_HVT U395 ( .A1(n297), .A2(n371), .S0(n280), .Y(n609) );
  INVX1_HVT U396 ( .A(n572), .Y(n532) );
  XNOR2X1_HVT U397 ( .A1(n373), .A2(n217), .Y(n482) );
  INVX0_HVT U398 ( .A(n541), .Y(n392) );
  INVX0_HVT U399 ( .A(n410), .Y(n509) );
  MUX21X1_HVT U400 ( .A1(n475), .A2(n297), .S0(n280), .Y(n742) );
  INVX1_HVT U401 ( .A(n569), .Y(n551) );
  NAND2X0_HVT U402 ( .A1(n504), .A2(n399), .Y(n400) );
  NAND2X0_HVT U403 ( .A1(n689), .A2(n484), .Y(n401) );
  INVX0_HVT U404 ( .A(n484), .Y(n399) );
  MUX41X1_HVT U405 ( .A1(n606), .A3(n604), .A2(n608), .A4(n605), .S0(n368), 
        .S1(n513), .Y(n603) );
  NAND2X0_HVT U406 ( .A1(n497), .A2(n403), .Y(n404) );
  NAND2X0_HVT U407 ( .A1(n404), .A2(n358), .Y(n755) );
  MUX41X1_HVT U408 ( .A1(n19), .A3(n685), .A2(n690), .A4(n686), .S0(n368), 
        .S1(n491), .Y(n684) );
  AND2X1_HVT U409 ( .A1(n403), .A2(n505), .Y(n405) );
  NAND2X0_HVT U410 ( .A1(n722), .A2(n433), .Y(n406) );
  NAND2X0_HVT U411 ( .A1(n720), .A2(n415), .Y(n407) );
  NAND2X0_HVT U412 ( .A1(n407), .A2(n406), .Y(n719) );
  NAND2X0_HVT U413 ( .A1(n342), .A2(n304), .Y(n408) );
  NAND2X0_HVT U414 ( .A1(n757), .A2(n309), .Y(n409) );
  NAND2X0_HVT U415 ( .A1(n408), .A2(n409), .Y(n700) );
  MUX41X1_HVT U416 ( .A1(n480), .A3(n560), .A2(n761), .A4(n218), .S0(n448), 
        .S1(n431), .Y(n685) );
  MUX41X1_HVT U417 ( .A1(n428), .A3(n532), .A2(n751), .A4(n771), .S0(n412), 
        .S1(n349), .Y(n646) );
  MUX41X1_HVT U418 ( .A1(n651), .A3(n653), .A2(n650), .A4(n652), .S0(n512), 
        .S1(n309), .Y(n649) );
  OR2X1_HVT U419 ( .A1(n504), .A2(n487), .Y(n436) );
  OA21X1_HVT U420 ( .A1(n309), .A2(n769), .A3(n538), .Y(n584) );
  NAND2X0_HVT U421 ( .A1(n567), .A2(n216), .Y(n413) );
  NAND2X0_HVT U422 ( .A1(n552), .A2(n494), .Y(n414) );
  NAND2X0_HVT U423 ( .A1(n413), .A2(n414), .Y(n589) );
  MUX41X1_HVT U424 ( .A1(n308), .A3(n498), .A2(n543), .A4(n430), .S0(n377), 
        .S1(n349), .Y(n639) );
  NAND2X0_HVT U425 ( .A1(n398), .A2(n415), .Y(n416) );
  NAND2X0_HVT U426 ( .A1(n397), .A2(n488), .Y(n417) );
  INVX1_HVT U427 ( .A(n467), .Y(n695) );
  INVX1_HVT U428 ( .A(n764), .Y(n535) );
  MUX41X1_HVT U429 ( .A1(n625), .A3(n623), .A2(n630), .A4(n629), .S0(n441), 
        .S1(n496), .Y(n622) );
  NAND2X0_HVT U430 ( .A1(n622), .A2(n327), .Y(n420) );
  NAND2X0_HVT U431 ( .A1(n419), .A2(n420), .Y(out[5]) );
  INVX1_HVT U432 ( .A(n570), .Y(n552) );
  NAND2X0_HVT U433 ( .A1(n660), .A2(n309), .Y(n421) );
  NAND2X0_HVT U434 ( .A1(n659), .A2(n495), .Y(n422) );
  NAND2X0_HVT U435 ( .A1(n421), .A2(n422), .Y(n656) );
  NAND2X0_HVT U436 ( .A1(n718), .A2(n453), .Y(n423) );
  NAND2X0_HVT U437 ( .A1(n716), .A2(n284), .Y(n424) );
  NAND2X0_HVT U438 ( .A1(n423), .A2(n424), .Y(n715) );
  MUX41X1_HVT U439 ( .A1(n636), .A3(n640), .A2(n635), .A4(n639), .S0(n496), 
        .S1(n441), .Y(n634) );
  NAND2X0_HVT U440 ( .A1(n642), .A2(n327), .Y(n425) );
  NAND2X0_HVT U441 ( .A1(n634), .A2(n351), .Y(n426) );
  NAND2X0_HVT U442 ( .A1(n425), .A2(n426), .Y(out[4]) );
  INVX1_HVT U443 ( .A(n491), .Y(n441) );
  INVX1_HVT U444 ( .A(n535), .Y(n470) );
  MUX41X1_HVT U445 ( .A1(n380), .A3(n755), .A2(n468), .A4(n530), .S0(n448), 
        .S1(n476), .Y(n467) );
  MUX41X1_HVT U446 ( .A1(n697), .A3(n695), .A2(n696), .A4(n693), .S0(n368), 
        .S1(n441), .Y(n692) );
  NAND2X0_HVT U447 ( .A1(n773), .A2(n433), .Y(n434) );
  NAND2X0_HVT U448 ( .A1(n644), .A2(n448), .Y(n435) );
  NAND2X0_HVT U449 ( .A1(n434), .A2(n435), .Y(n643) );
  MUX21X1_HVT U450 ( .A1(n539), .A2(n755), .S0(n486), .Y(n644) );
  INVX1_HVT U451 ( .A(n490), .Y(n448) );
  MUX41X1_HVT U452 ( .A1(n525), .A3(n735), .A2(n762), .A4(n568), .S0(n415), 
        .S1(n476), .Y(n696) );
  NAND2X0_HVT U453 ( .A1(n459), .A2(n460), .Y(n669) );
  NBUFFX2_HVT U454 ( .A(n512), .Y(n491) );
  MUX41X1_HVT U455 ( .A1(n753), .A3(n538), .A2(n641), .A4(n536), .S0(n490), 
        .S1(n431), .Y(n640) );
  INVX1_HVT U456 ( .A(n573), .Y(n540) );
  NAND2X0_HVT U457 ( .A1(n481), .A2(n442), .Y(n443) );
  NAND2X0_HVT U458 ( .A1(n683), .A2(n733), .Y(n444) );
  NAND2X0_HVT U459 ( .A1(n444), .A2(n443), .Y(n682) );
  INVX0_HVT U460 ( .A(n733), .Y(n442) );
  MUX41X1_HVT U461 ( .A1(n766), .A3(n724), .A2(n758), .A4(n533), .S0(n486), 
        .S1(n387), .Y(n722) );
  NAND2X0_HVT U462 ( .A1(n456), .A2(n457), .Y(out[1]) );
  MUX41X1_HVT U463 ( .A1(n607), .A3(n759), .A2(n742), .A4(n552), .S0(n412), 
        .S1(n476), .Y(n606) );
  MUX21X1_HVT U464 ( .A1(n553), .A2(n774), .S0(n489), .Y(n673) );
  NAND2X0_HVT U465 ( .A1(n586), .A2(n327), .Y(n449) );
  NAND2X0_HVT U466 ( .A1(n579), .A2(n351), .Y(n450) );
  NAND2X0_HVT U467 ( .A1(n450), .A2(n449), .Y(out[7]) );
  NAND2X0_HVT U468 ( .A1(n665), .A2(n494), .Y(n452) );
  NAND2X0_HVT U469 ( .A1(n451), .A2(n452), .Y(n663) );
  AO21X1_HVT U470 ( .A1(n489), .A2(n430), .A3(n381), .Y(n664) );
  NAND2X0_HVT U471 ( .A1(n661), .A2(n453), .Y(n454) );
  NAND2X0_HVT U472 ( .A1(n537), .A2(n317), .Y(n455) );
  NAND2X0_HVT U473 ( .A1(n454), .A2(n455), .Y(n660) );
  NAND2X0_HVT U474 ( .A1(n701), .A2(in[6]), .Y(n456) );
  NAND2X0_HVT U475 ( .A1(n692), .A2(n351), .Y(n457) );
  NAND2X0_HVT U476 ( .A1(n458), .A2(n671), .Y(n459) );
  NAND2X0_HVT U477 ( .A1(n35), .A2(n747), .Y(n460) );
  INVX0_HVT U478 ( .A(n317), .Y(n458) );
  NAND2X0_HVT U479 ( .A1(n398), .A2(n387), .Y(n461) );
  NAND2X0_HVT U480 ( .A1(n744), .A2(n513), .Y(n462) );
  NAND2X0_HVT U481 ( .A1(n461), .A2(n462), .Y(n729) );
  NAND2X0_HVT U482 ( .A1(n584), .A2(n317), .Y(n463) );
  NAND2X0_HVT U483 ( .A1(n585), .A2(n488), .Y(n464) );
  NAND2X0_HVT U484 ( .A1(n464), .A2(n463), .Y(n583) );
  NAND2X0_HVT U485 ( .A1(n666), .A2(n513), .Y(n465) );
  NAND2X0_HVT U486 ( .A1(n663), .A2(n441), .Y(n466) );
  NAND2X0_HVT U487 ( .A1(n465), .A2(n466), .Y(n662) );
  NAND2X0_HVT U488 ( .A1(n217), .A2(n397), .Y(n468) );
  MUX21X1_HVT U489 ( .A1(n418), .A2(n475), .S0(n395), .Y(n769) );
  MUX41X1_HVT U490 ( .A1(n388), .A3(n475), .A2(n575), .A4(n418), .S0(n367), 
        .S1(n427), .Y(n474) );
  MUX41X1_HVT U491 ( .A1(n764), .A3(n724), .A2(n755), .A4(n394), .S0(n284), 
        .S1(n476), .Y(n581) );
  MUX41X1_HVT U492 ( .A1(n734), .A3(n560), .A2(n330), .A4(n523), .S0(n412), 
        .S1(n336), .Y(n635) );
  MUX21X1_HVT U493 ( .A1(n297), .A2(n563), .S0(n513), .Y(n727) );
  AND2X1_HVT U494 ( .A1(n706), .A2(n505), .Y(n478) );
  MUX21X1_HVT U495 ( .A1(n346), .A2(n429), .S0(n396), .Y(n572) );
  NAND2X0_HVT U496 ( .A1(n501), .A2(n500), .Y(n772) );
  MUX21X1_HVT U497 ( .A1(n297), .A2(n499), .S0(n395), .Y(n573) );
  NBUFFX2_HVT U498 ( .A(n775), .Y(n503) );
  MUX21X1_HVT U499 ( .A1(n499), .A2(n502), .S0(n507), .Y(n661) );
  MUX21X1_HVT U500 ( .A1(n502), .A2(n374), .S0(n506), .Y(n596) );
  MUX21X1_HVT U501 ( .A1(n374), .A2(n504), .S0(n410), .Y(n597) );
  MUX21X1_HVT U502 ( .A1(n502), .A2(n475), .S0(n396), .Y(n766) );
  AND2X1_HVT U503 ( .A1(n506), .A2(n371), .Y(n480) );
  AND2X1_HVT U504 ( .A1(n374), .A2(n670), .Y(n481) );
  MUX21X1_HVT U505 ( .A1(n272), .A2(n374), .S0(n489), .Y(n658) );
  MUX21X1_HVT U506 ( .A1(n767), .A2(n499), .S0(n507), .Y(n708) );
  NBUFFX2_HVT U507 ( .A(n512), .Y(n492) );
  MUX21X1_HVT U508 ( .A1(n694), .A2(n398), .S0(n494), .Y(n601) );
  XOR2X1_HVT U509 ( .A1(n218), .A2(n497), .Y(n732) );
  NAND2X0_HVT U510 ( .A1(n307), .A2(n361), .Y(n775) );
  AND2X1_HVT U511 ( .A1(n411), .A2(n447), .Y(n483) );
  MUX21X1_HVT U512 ( .A1(n497), .A2(n297), .S0(n218), .Y(n741) );
  MUX21X1_HVT U513 ( .A1(n371), .A2(n497), .S0(n432), .Y(n758) );
  MUX21X1_HVT U514 ( .A1(n628), .A2(n504), .S0(n484), .Y(n627) );
  MUX21X1_HVT U515 ( .A1(n774), .A2(n316), .S0(n488), .Y(n657) );
  MUX21X1_HVT U516 ( .A1(n497), .A2(n429), .S0(n506), .Y(n574) );
  MUX21X1_HVT U517 ( .A1(n497), .A2(n212), .S0(n495), .Y(n689) );
  XNOR2X1_HVT U518 ( .A1(n517), .A2(n471), .Y(n484) );
  AND2X1_HVT U519 ( .A1(n502), .A2(n447), .Y(n485) );
  NBUFFX2_HVT U520 ( .A(in[5]), .Y(n512) );
  NAND2X0_HVT U521 ( .A1(n318), .A2(n324), .Y(n776) );
  MUX21X1_HVT U522 ( .A1(n469), .A2(n346), .S0(n403), .Y(n576) );
  MUX21X1_HVT U523 ( .A1(n469), .A2(n342), .S0(n395), .Y(n570) );
  MUX21X1_HVT U524 ( .A1(n373), .A2(n469), .S0(n395), .Y(n750) );
  MUX21X1_HVT U525 ( .A1(n469), .A2(n373), .S0(n507), .Y(n569) );
  NBUFFX2_HVT U526 ( .A(n361), .Y(n497) );
endmodule

