
module sbox_7 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342;

  MUX21X1_HVT U1 ( .A1(n1), .A2(n2), .S0(in[6]), .Y(out[7]) );
  AO221X1_HVT U2 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .A5(n7), .Y(n2) );
  AO22X1_HVT U3 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .Y(n7) );
  AO221X1_HVT U4 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .A5(n16), .Y(n11)
         );
  AO221X1_HVT U5 ( .A1(n17), .A2(n18), .A3(n19), .A4(n20), .A5(n21), .Y(n16)
         );
  AO221X1_HVT U6 ( .A1(n13), .A2(n22), .A3(n14), .A4(n23), .A5(n24), .Y(n9) );
  AO22X1_HVT U7 ( .A1(n20), .A2(n25), .A3(n17), .A4(n26), .Y(n24) );
  NAND2X0_HVT U8 ( .A1(n27), .A2(n28), .Y(n23) );
  NAND2X0_HVT U9 ( .A1(n29), .A2(n30), .Y(n22) );
  AO221X1_HVT U10 ( .A1(n31), .A2(n14), .A3(n32), .A4(in[2]), .A5(n33), .Y(n6)
         );
  OAI22X1_HVT U11 ( .A1(n34), .A2(n35), .A3(n26), .A4(n36), .Y(n33) );
  AO221X1_HVT U12 ( .A1(n20), .A2(n37), .A3(n14), .A4(n38), .A5(n39), .Y(n4)
         );
  AO21X1_HVT U13 ( .A1(n17), .A2(n40), .A3(n41), .Y(n39) );
  AO221X1_HVT U14 ( .A1(n3), .A2(n42), .A3(n10), .A4(n43), .A5(n44), .Y(n1) );
  AO22X1_HVT U15 ( .A1(n8), .A2(n45), .A3(n5), .A4(n46), .Y(n44) );
  AO221X1_HVT U16 ( .A1(n47), .A2(n13), .A3(n48), .A4(n14), .A5(n49), .Y(n46)
         );
  AO22X1_HVT U17 ( .A1(n20), .A2(n50), .A3(n17), .A4(in[4]), .Y(n49) );
  AO221X1_HVT U18 ( .A1(n51), .A2(n52), .A3(n20), .A4(n53), .A5(n54), .Y(n45)
         );
  INVX0_HVT U19 ( .A(n55), .Y(n54) );
  AO21X1_HVT U20 ( .A1(n56), .A2(n57), .A3(n17), .Y(n52) );
  AO221X1_HVT U21 ( .A1(n13), .A2(n58), .A3(n59), .A4(n14), .A5(n60), .Y(n43)
         );
  OAI221X1_HVT U22 ( .A1(n61), .A2(n36), .A3(n62), .A4(n63), .A5(n64), .Y(n60)
         );
  AO221X1_HVT U23 ( .A1(n20), .A2(n65), .A3(n14), .A4(n66), .A5(n67), .Y(n42)
         );
  AO22X1_HVT U24 ( .A1(n13), .A2(n68), .A3(n17), .A4(n69), .Y(n67) );
  NAND2X0_HVT U25 ( .A1(n70), .A2(n71), .Y(n66) );
  NAND2X0_HVT U26 ( .A1(n50), .A2(n72), .Y(n65) );
  MUX21X1_HVT U27 ( .A1(n73), .A2(n74), .S0(in[6]), .Y(out[6]) );
  AO221X1_HVT U28 ( .A1(n10), .A2(n75), .A3(n5), .A4(n76), .A5(n77), .Y(n74)
         );
  AO22X1_HVT U29 ( .A1(n8), .A2(n78), .A3(n3), .A4(n79), .Y(n77) );
  AO221X1_HVT U30 ( .A1(n13), .A2(n80), .A3(n31), .A4(n14), .A5(n81), .Y(n79)
         );
  AO22X1_HVT U31 ( .A1(n17), .A2(n82), .A3(n20), .A4(n29), .Y(n81) );
  AO221X1_HVT U32 ( .A1(n14), .A2(n83), .A3(n20), .A4(n84), .A5(n85), .Y(n78)
         );
  AO22X1_HVT U33 ( .A1(n13), .A2(n86), .A3(n17), .A4(n87), .Y(n85) );
  NAND2X0_HVT U34 ( .A1(n88), .A2(n28), .Y(n83) );
  NAND3X0_HVT U35 ( .A1(n89), .A2(n55), .A3(n90), .Y(n76) );
  OA22X1_HVT U36 ( .A1(n63), .A2(n62), .A3(n91), .A4(n92), .Y(n90) );
  NAND3X0_HVT U37 ( .A1(n13), .A2(n93), .A3(n94), .Y(n55) );
  NAND3X0_HVT U38 ( .A1(n50), .A2(n61), .A3(n17), .Y(n89) );
  AO221X1_HVT U39 ( .A1(n48), .A2(n20), .A3(n31), .A4(n13), .A5(n95), .Y(n75)
         );
  OAI22X1_HVT U40 ( .A1(n36), .A2(n96), .A3(n97), .A4(n92), .Y(n95) );
  AND2X1_HVT U41 ( .A1(n93), .A2(n98), .Y(n31) );
  AND2X1_HVT U42 ( .A1(n99), .A2(n98), .Y(n48) );
  AO221X1_HVT U43 ( .A1(n3), .A2(n100), .A3(n5), .A4(n101), .A5(n102), .Y(n73)
         );
  AO22X1_HVT U44 ( .A1(n8), .A2(n103), .A3(n10), .A4(n104), .Y(n102) );
  AO221X1_HVT U45 ( .A1(n105), .A2(n17), .A3(n20), .A4(n106), .A5(n107), .Y(
        n104) );
  AO22X1_HVT U46 ( .A1(n14), .A2(n99), .A3(n13), .A4(n108), .Y(n107) );
  AO221X1_HVT U47 ( .A1(n109), .A2(n17), .A3(n110), .A4(n20), .A5(n111), .Y(
        n103) );
  AO22X1_HVT U48 ( .A1(n14), .A2(n61), .A3(n112), .A4(n13), .Y(n111) );
  INVX0_HVT U49 ( .A(n40), .Y(n110) );
  NAND2X0_HVT U50 ( .A1(n27), .A2(n113), .Y(n40) );
  NAND4X0_HVT U51 ( .A1(n114), .A2(n115), .A3(n116), .A4(n117), .Y(n101) );
  OA22X1_HVT U52 ( .A1(n62), .A2(n50), .A3(n12), .A4(n92), .Y(n117) );
  INVX0_HVT U53 ( .A(n86), .Y(n12) );
  NAND3X0_HVT U54 ( .A1(n15), .A2(n118), .A3(n119), .Y(n116) );
  AO221X1_HVT U55 ( .A1(n20), .A2(n120), .A3(in[3]), .A4(n13), .A5(n121), .Y(
        n100) );
  OAI21X1_HVT U56 ( .A1(n59), .A2(in[2]), .A3(n122), .Y(n121) );
  MUX21X1_HVT U57 ( .A1(n123), .A2(n124), .S0(in[6]), .Y(out[5]) );
  AO221X1_HVT U58 ( .A1(n5), .A2(n125), .A3(n8), .A4(n126), .A5(n127), .Y(n124) );
  AO22X1_HVT U59 ( .A1(n3), .A2(n128), .A3(n10), .A4(n129), .Y(n127) );
  OAI221X1_HVT U60 ( .A1(n51), .A2(n36), .A3(n92), .A4(n130), .A5(n131), .Y(
        n129) );
  MUX21X1_HVT U61 ( .A1(n132), .A2(n133), .S0(n134), .Y(n131) );
  NAND2X0_HVT U62 ( .A1(in[2]), .A2(n135), .Y(n133) );
  NAND2X0_HVT U63 ( .A1(in[3]), .A2(n13), .Y(n132) );
  AO221X1_HVT U64 ( .A1(n17), .A2(n136), .A3(n137), .A4(n20), .A5(n138), .Y(
        n128) );
  AO22X1_HVT U65 ( .A1(n14), .A2(n135), .A3(n139), .A4(n13), .Y(n138) );
  AO222X1_HVT U66 ( .A1(n140), .A2(n20), .A3(n141), .A4(n142), .A5(n143), .A6(
        n13), .Y(n126) );
  AO21X1_HVT U67 ( .A1(n144), .A2(n57), .A3(n17), .Y(n141) );
  NAND2X0_HVT U68 ( .A1(n28), .A2(n30), .Y(n144) );
  AO221X1_HVT U69 ( .A1(n14), .A2(n145), .A3(n146), .A4(n13), .A5(n147), .Y(
        n125) );
  AO22X1_HVT U70 ( .A1(n20), .A2(n94), .A3(n17), .A4(n148), .Y(n147) );
  INVX0_HVT U71 ( .A(n71), .Y(n146) );
  AO221X1_HVT U72 ( .A1(n10), .A2(n149), .A3(n8), .A4(n150), .A5(n151), .Y(
        n123) );
  AO22X1_HVT U73 ( .A1(n3), .A2(n152), .A3(n5), .A4(n153), .Y(n151) );
  AO222X1_HVT U74 ( .A1(n17), .A2(n154), .A3(n155), .A4(n156), .A5(n19), .A6(
        n14), .Y(n153) );
  AO21X1_HVT U75 ( .A1(n157), .A2(in[2]), .A3(n20), .Y(n155) );
  AO221X1_HVT U76 ( .A1(n13), .A2(n158), .A3(n17), .A4(n70), .A5(n159), .Y(
        n152) );
  AO22X1_HVT U77 ( .A1(n160), .A2(n14), .A3(n20), .A4(n108), .Y(n159) );
  NAND2X0_HVT U78 ( .A1(n28), .A2(n161), .Y(n158) );
  NAND3X0_HVT U79 ( .A1(n162), .A2(n163), .A3(n164), .Y(n150) );
  OA22X1_HVT U80 ( .A1(n36), .A2(n82), .A3(n92), .A4(n165), .Y(n164) );
  NAND3X0_HVT U81 ( .A1(n99), .A2(n18), .A3(n20), .Y(n163) );
  AO21X1_HVT U82 ( .A1(n113), .A2(n120), .A3(n35), .Y(n162) );
  AO221X1_HVT U83 ( .A1(n20), .A2(n154), .A3(n14), .A4(n135), .A5(n166), .Y(
        n149) );
  AO221X1_HVT U84 ( .A1(n13), .A2(n167), .A3(n168), .A4(n17), .A5(n169), .Y(
        n166) );
  INVX0_HVT U85 ( .A(n170), .Y(n169) );
  NAND2X0_HVT U86 ( .A1(n15), .A2(n93), .Y(n167) );
  MUX21X1_HVT U87 ( .A1(n171), .A2(n172), .S0(in[6]), .Y(out[4]) );
  AO221X1_HVT U88 ( .A1(n5), .A2(n173), .A3(n8), .A4(n174), .A5(n175), .Y(n172) );
  AO22X1_HVT U89 ( .A1(n10), .A2(n176), .A3(n3), .A4(n177), .Y(n175) );
  AO221X1_HVT U90 ( .A1(n14), .A2(n71), .A3(n37), .A4(n17), .A5(n178), .Y(n177) );
  AO22X1_HVT U91 ( .A1(n13), .A2(n38), .A3(n20), .A4(n143), .Y(n178) );
  AND2X1_HVT U92 ( .A1(n142), .A2(n97), .Y(n37) );
  AO221X1_HVT U93 ( .A1(n13), .A2(n69), .A3(n179), .A4(n14), .A5(n180), .Y(
        n176) );
  AO22X1_HVT U94 ( .A1(n20), .A2(n88), .A3(n181), .A4(n17), .Y(n180) );
  AND2X1_HVT U95 ( .A1(n99), .A2(n135), .Y(n181) );
  AO221X1_HVT U96 ( .A1(n182), .A2(n20), .A3(n183), .A4(n14), .A5(n184), .Y(
        n174) );
  AO21X1_HVT U97 ( .A1(n160), .A2(n17), .A3(n41), .Y(n184) );
  INVX0_HVT U98 ( .A(n185), .Y(n41) );
  AO222X1_HVT U99 ( .A1(n17), .A2(n58), .A3(in[2]), .A4(n186), .A5(n109), .A6(
        n14), .Y(n173) );
  INVX0_HVT U100 ( .A(n106), .Y(n109) );
  NAND2X0_HVT U101 ( .A1(n187), .A2(n72), .Y(n106) );
  NAND2X0_HVT U102 ( .A1(n61), .A2(n50), .Y(n186) );
  AO221X1_HVT U103 ( .A1(n8), .A2(n188), .A3(n10), .A4(n189), .A5(n190), .Y(
        n171) );
  AO22X1_HVT U104 ( .A1(n5), .A2(n191), .A3(n3), .A4(n192), .Y(n190) );
  NAND3X0_HVT U105 ( .A1(n185), .A2(n122), .A3(n193), .Y(n192) );
  OA22X1_HVT U106 ( .A1(n92), .A2(n194), .A3(n18), .A4(n62), .Y(n193) );
  NAND2X0_HVT U107 ( .A1(n13), .A2(n154), .Y(n185) );
  AO221X1_HVT U108 ( .A1(n179), .A2(n17), .A3(n20), .A4(n99), .A5(n195), .Y(
        n191) );
  AO22X1_HVT U109 ( .A1(n196), .A2(n14), .A3(n13), .A4(n108), .Y(n195) );
  AND2X1_HVT U110 ( .A1(n27), .A2(n194), .Y(n179) );
  AO221X1_HVT U111 ( .A1(n17), .A2(n197), .A3(n198), .A4(n156), .A5(n199), .Y(
        n189) );
  INVX0_HVT U112 ( .A(n200), .Y(n199) );
  OAI21X1_HVT U113 ( .A1(n201), .A2(n57), .A3(n62), .Y(n198) );
  NAND2X0_HVT U114 ( .A1(n25), .A2(n187), .Y(n197) );
  AO221X1_HVT U115 ( .A1(n202), .A2(n203), .A3(n17), .A4(n204), .A5(n205), .Y(
        n188) );
  AO22X1_HVT U116 ( .A1(n206), .A2(n13), .A3(n51), .A4(n20), .Y(n205) );
  INVX0_HVT U117 ( .A(n80), .Y(n51) );
  NAND2X0_HVT U118 ( .A1(n187), .A2(n120), .Y(n80) );
  MUX21X1_HVT U119 ( .A1(n207), .A2(n208), .S0(in[6]), .Y(out[3]) );
  MUX41X1_HVT U120 ( .A1(n209), .A3(n210), .A2(n211), .A4(n212), .S0(in[0]), 
        .S1(in[5]), .Y(n208) );
  AO222X1_HVT U121 ( .A1(n213), .A2(n17), .A3(n214), .A4(n215), .A5(n20), .A6(
        n50), .Y(n212) );
  AO21X1_HVT U122 ( .A1(in[7]), .A2(n216), .A3(n14), .Y(n215) );
  NAND2X0_HVT U123 ( .A1(n88), .A2(n113), .Y(n216) );
  INVX0_HVT U124 ( .A(n69), .Y(n213) );
  NAND2X0_HVT U125 ( .A1(n98), .A2(n145), .Y(n69) );
  AO221X1_HVT U126 ( .A1(n217), .A2(n20), .A3(n17), .A4(n148), .A5(n218), .Y(
        n211) );
  AO22X1_HVT U127 ( .A1(n219), .A2(n14), .A3(n13), .A4(n156), .Y(n218) );
  AO221X1_HVT U128 ( .A1(n13), .A2(n136), .A3(n14), .A4(n156), .A5(n220), .Y(
        n210) );
  MUX21X1_HVT U129 ( .A1(n221), .A2(n222), .S0(n119), .Y(n220) );
  XOR2X1_HVT U130 ( .A1(in[2]), .A2(in[1]), .Y(n119) );
  AND2X1_HVT U131 ( .A1(n135), .A2(n118), .Y(n222) );
  AO22X1_HVT U132 ( .A1(n20), .A2(in[4]), .A3(n17), .A4(in[3]), .Y(n221) );
  NAND2X0_HVT U133 ( .A1(n135), .A2(n194), .Y(n136) );
  AO221X1_HVT U134 ( .A1(n139), .A2(n14), .A3(n18), .A4(n118), .A5(n223), .Y(
        n209) );
  AO22X1_HVT U135 ( .A1(n59), .A2(n13), .A3(n20), .A4(n154), .Y(n223) );
  AND2X1_HVT U136 ( .A1(n71), .A2(n120), .Y(n59) );
  INVX0_HVT U137 ( .A(n25), .Y(n139) );
  MUX41X1_HVT U138 ( .A1(n224), .A3(n225), .A2(n226), .A4(n227), .S0(in[0]), 
        .S1(in[5]), .Y(n207) );
  NAND3X0_HVT U139 ( .A1(n228), .A2(n229), .A3(n230), .Y(n227) );
  OA221X1_HVT U140 ( .A1(n36), .A2(n88), .A3(n57), .A4(n71), .A5(n200), .Y(
        n230) );
  OA22X1_HVT U141 ( .A1(n62), .A2(n25), .A3(n35), .A4(n15), .Y(n228) );
  OAI222X1_HVT U142 ( .A1(n35), .A2(n160), .A3(n98), .A4(n62), .A5(n231), .A6(
        n92), .Y(n226) );
  AO221X1_HVT U143 ( .A1(n182), .A2(n13), .A3(n232), .A4(n14), .A5(n233), .Y(
        n225) );
  AO22X1_HVT U144 ( .A1(n17), .A2(n70), .A3(n234), .A4(n20), .Y(n233) );
  AND2X1_HVT U145 ( .A1(n88), .A2(n29), .Y(n182) );
  AO221X1_HVT U146 ( .A1(n235), .A2(n13), .A3(n236), .A4(n14), .A5(n237), .Y(
        n224) );
  AO22X1_HVT U147 ( .A1(n206), .A2(n20), .A3(n17), .A4(n82), .Y(n237) );
  INVX0_HVT U148 ( .A(n68), .Y(n206) );
  NAND2X0_HVT U149 ( .A1(n238), .A2(n88), .Y(n68) );
  INVX0_HVT U150 ( .A(n165), .Y(n236) );
  NAND2X0_HVT U151 ( .A1(n70), .A2(n187), .Y(n165) );
  MUX21X1_HVT U152 ( .A1(n239), .A2(n240), .S0(in[6]), .Y(out[2]) );
  AO221X1_HVT U153 ( .A1(n5), .A2(n241), .A3(n8), .A4(n242), .A5(n243), .Y(
        n240) );
  AO22X1_HVT U154 ( .A1(n10), .A2(n244), .A3(n3), .A4(n245), .Y(n243) );
  AO221X1_HVT U155 ( .A1(n14), .A2(n130), .A3(n134), .A4(n246), .A5(n247), .Y(
        n245) );
  MUX21X1_HVT U156 ( .A1(n32), .A2(n248), .S0(in[2]), .Y(n247) );
  NOR2X0_HVT U157 ( .A1(n134), .A2(n249), .Y(n248) );
  INVX0_HVT U158 ( .A(n142), .Y(n32) );
  AO22X1_HVT U159 ( .A1(n13), .A2(n87), .A3(n20), .A4(in[3]), .Y(n246) );
  XNOR2X1_HVT U160 ( .A1(n118), .A2(in[1]), .Y(n134) );
  NAND3X0_HVT U161 ( .A1(n250), .A2(n251), .A3(n252), .Y(n244) );
  AOI22X1_HVT U162 ( .A1(n17), .A2(n253), .A3(n14), .A4(n19), .Y(n252) );
  AO21X1_HVT U163 ( .A1(n187), .A2(n254), .A3(n35), .Y(n250) );
  AO221X1_HVT U164 ( .A1(n196), .A2(n13), .A3(n255), .A4(n14), .A5(n256), .Y(
        n242) );
  AO221X1_HVT U165 ( .A1(n17), .A2(n108), .A3(n20), .A4(n26), .A5(n21), .Y(
        n256) );
  NAND2X0_HVT U166 ( .A1(n97), .A2(n113), .Y(n108) );
  NAND4X0_HVT U167 ( .A1(n257), .A2(n251), .A3(n170), .A4(n64), .Y(n241) );
  NAND2X0_HVT U168 ( .A1(n14), .A2(in[1]), .Y(n170) );
  NAND2X0_HVT U169 ( .A1(n105), .A2(n20), .Y(n251) );
  INVX0_HVT U170 ( .A(n28), .Y(n105) );
  AO21X1_HVT U171 ( .A1(n94), .A2(n50), .A3(n35), .Y(n257) );
  AO221X1_HVT U172 ( .A1(n10), .A2(n258), .A3(n5), .A4(n259), .A5(n260), .Y(
        n239) );
  AO22X1_HVT U173 ( .A1(n3), .A2(n261), .A3(n262), .A4(n8), .Y(n260) );
  MUX21X1_HVT U174 ( .A1(n263), .A2(n137), .S0(n264), .Y(n262) );
  AND2X1_HVT U175 ( .A1(n92), .A2(n62), .Y(n264) );
  MUX21X1_HVT U176 ( .A1(n47), .A2(n265), .S0(in[2]), .Y(n263) );
  INVX0_HVT U177 ( .A(n156), .Y(n47) );
  NAND2X0_HVT U178 ( .A1(n93), .A2(n266), .Y(n156) );
  NAND3X0_HVT U179 ( .A1(n115), .A2(n267), .A3(n268), .Y(n261) );
  AOI22X1_HVT U180 ( .A1(n57), .A2(n84), .A3(n20), .A4(n160), .Y(n268) );
  AND2X1_HVT U181 ( .A1(n238), .A2(n30), .Y(n160) );
  NAND2X0_HVT U182 ( .A1(n97), .A2(n238), .Y(n84) );
  AO221X1_HVT U183 ( .A1(n217), .A2(n14), .A3(n96), .A4(n17), .A5(n269), .Y(
        n259) );
  AO221X1_HVT U184 ( .A1(n20), .A2(n270), .A3(n202), .A4(n203), .A5(n271), .Y(
        n269) );
  INVX0_HVT U185 ( .A(n115), .Y(n271) );
  NAND2X0_HVT U186 ( .A1(n183), .A2(n13), .Y(n115) );
  AND2X1_HVT U187 ( .A1(n154), .A2(n194), .Y(n183) );
  INVX0_HVT U188 ( .A(n267), .Y(n202) );
  NAND2X0_HVT U189 ( .A1(n71), .A2(n72), .Y(n270) );
  INVX0_HVT U190 ( .A(n231), .Y(n96) );
  NAND2X0_HVT U191 ( .A1(n238), .A2(n266), .Y(n231) );
  INVX0_HVT U192 ( .A(n113), .Y(n217) );
  NAND2X0_HVT U193 ( .A1(in[1]), .A2(n94), .Y(n113) );
  AO221X1_HVT U194 ( .A1(n14), .A2(n272), .A3(n17), .A4(n50), .A5(n273), .Y(
        n258) );
  AO22X1_HVT U195 ( .A1(n13), .A2(n25), .A3(n91), .A4(n20), .Y(n273) );
  INVX0_HVT U196 ( .A(n274), .Y(n91) );
  NAND2X0_HVT U197 ( .A1(n98), .A2(n194), .Y(n272) );
  MUX21X1_HVT U198 ( .A1(n275), .A2(n276), .S0(in[6]), .Y(out[1]) );
  AO221X1_HVT U199 ( .A1(n3), .A2(n277), .A3(n5), .A4(n278), .A5(n279), .Y(
        n276) );
  AO22X1_HVT U200 ( .A1(n8), .A2(n280), .A3(n10), .A4(n281), .Y(n279) );
  AO221X1_HVT U201 ( .A1(n219), .A2(n13), .A3(n14), .A4(n249), .A5(n282), .Y(
        n281) );
  OAI21X1_HVT U202 ( .A1(n283), .A2(n62), .A3(n64), .Y(n282) );
  INVX0_HVT U203 ( .A(n204), .Y(n219) );
  NAND2X0_HVT U204 ( .A1(n97), .A2(n28), .Y(n204) );
  NAND2X0_HVT U205 ( .A1(n249), .A2(in[1]), .Y(n28) );
  INVX0_HVT U206 ( .A(n284), .Y(n10) );
  AO221X1_HVT U207 ( .A1(n285), .A2(n20), .A3(n19), .A4(n13), .A5(n286), .Y(
        n280) );
  MUX21X1_HVT U208 ( .A1(n17), .A2(n14), .S0(n38), .Y(n286) );
  NAND2X0_HVT U209 ( .A1(n145), .A2(n201), .Y(n38) );
  OA21X1_HVT U210 ( .A1(n143), .A2(in[1]), .A3(n71), .Y(n19) );
  INVX0_HVT U211 ( .A(n287), .Y(n8) );
  AO221X1_HVT U212 ( .A1(n140), .A2(n13), .A3(n288), .A4(n14), .A5(n289), .Y(
        n278) );
  AO22X1_HVT U213 ( .A1(n17), .A2(n274), .A3(n20), .A4(n290), .Y(n289) );
  NAND2X0_HVT U214 ( .A1(n97), .A2(n29), .Y(n290) );
  INVX0_HVT U215 ( .A(n130), .Y(n288) );
  NAND2X0_HVT U216 ( .A1(n99), .A2(n70), .Y(n130) );
  AND2X1_HVT U217 ( .A1(n86), .A2(n30), .Y(n140) );
  INVX0_HVT U218 ( .A(n291), .Y(n5) );
  NAND3X0_HVT U219 ( .A1(n229), .A2(n292), .A3(n293), .Y(n277) );
  OA222X1_HVT U220 ( .A1(in[3]), .A2(n35), .A3(n294), .A4(n36), .A5(n112), 
        .A6(n62), .Y(n293) );
  AND2X1_HVT U221 ( .A1(n25), .A2(n238), .Y(n112) );
  OA21X1_HVT U222 ( .A1(in[1]), .A2(n143), .A3(n29), .Y(n294) );
  NAND2X0_HVT U223 ( .A1(n295), .A2(n14), .Y(n292) );
  OA22X1_HVT U224 ( .A1(n92), .A2(n154), .A3(n203), .A4(n35), .Y(n229) );
  INVX0_HVT U225 ( .A(n296), .Y(n3) );
  OAI221X1_HVT U226 ( .A1(n297), .A2(n296), .A3(n298), .A4(n291), .A5(n299), 
        .Y(n275) );
  OA22X1_HVT U227 ( .A1(n300), .A2(n287), .A3(n301), .A4(n284), .Y(n299) );
  NAND2X0_HVT U228 ( .A1(in[5]), .A2(n302), .Y(n284) );
  OA221X1_HVT U229 ( .A1(n235), .A2(n92), .A3(n94), .A4(n62), .A5(n303), .Y(
        n301) );
  OA21X1_HVT U230 ( .A1(n35), .A2(n238), .A3(n122), .Y(n303) );
  OR2X1_HVT U231 ( .A1(n58), .A2(n36), .Y(n122) );
  NAND2X0_HVT U232 ( .A1(n26), .A2(n254), .Y(n58) );
  NAND2X0_HVT U233 ( .A1(in[1]), .A2(in[4]), .Y(n238) );
  NAND2X0_HVT U234 ( .A1(in[5]), .A2(in[0]), .Y(n287) );
  OA221X1_HVT U235 ( .A1(n304), .A2(n36), .A3(n305), .A4(n306), .A5(n267), .Y(
        n300) );
  NAND2X0_HVT U236 ( .A1(n14), .A2(n154), .Y(n267) );
  NAND2X0_HVT U237 ( .A1(n93), .A2(n135), .Y(n306) );
  OA21X1_HVT U238 ( .A1(n57), .A2(n97), .A3(n62), .Y(n305) );
  NAND2X0_HVT U239 ( .A1(n18), .A2(n203), .Y(n97) );
  NAND2X0_HVT U240 ( .A1(n302), .A2(n307), .Y(n291) );
  INVX0_HVT U241 ( .A(in[0]), .Y(n302) );
  OA221X1_HVT U242 ( .A1(n92), .A2(n34), .A3(n36), .A4(n283), .A5(n308), .Y(
        n298) );
  OA22X1_HVT U243 ( .A1(n35), .A2(n309), .A3(n310), .A4(n62), .Y(n308) );
  INVX0_HVT U244 ( .A(n120), .Y(n310) );
  NAND2X0_HVT U245 ( .A1(n99), .A2(n135), .Y(n309) );
  NAND2X0_HVT U246 ( .A1(n142), .A2(n72), .Y(n283) );
  NAND2X0_HVT U247 ( .A1(n145), .A2(n266), .Y(n34) );
  NAND2X0_HVT U248 ( .A1(n15), .A2(n203), .Y(n266) );
  NAND2X0_HVT U249 ( .A1(in[0]), .A2(n307), .Y(n296) );
  INVX0_HVT U250 ( .A(in[5]), .Y(n307) );
  OA221X1_HVT U251 ( .A1(n311), .A2(n35), .A3(n62), .A4(n312), .A5(n313), .Y(
        n297) );
  OA221X1_HVT U252 ( .A1(n92), .A2(n72), .A3(n36), .A4(n161), .A5(n64), .Y(
        n313) );
  NAND2X0_HVT U253 ( .A1(n196), .A2(n17), .Y(n64) );
  INVX0_HVT U254 ( .A(n93), .Y(n196) );
  MUX41X1_HVT U255 ( .A1(n314), .A3(n315), .A2(n316), .A4(n317), .S0(in[0]), 
        .S1(in[6]), .Y(out[0]) );
  MUX21X1_HVT U256 ( .A1(n318), .A2(n319), .S0(in[5]), .Y(n317) );
  AO221X1_HVT U257 ( .A1(n304), .A2(n13), .A3(n14), .A4(n25), .A5(n320), .Y(
        n319) );
  AO22X1_HVT U258 ( .A1(n321), .A2(n20), .A3(n17), .A4(n120), .Y(n320) );
  NAND2X0_HVT U259 ( .A1(n285), .A2(n203), .Y(n120) );
  NAND2X0_HVT U260 ( .A1(n87), .A2(n203), .Y(n25) );
  INVX0_HVT U261 ( .A(n312), .Y(n304) );
  NAND2X0_HVT U262 ( .A1(n50), .A2(n98), .Y(n312) );
  AO221X1_HVT U263 ( .A1(n255), .A2(n20), .A3(n14), .A4(in[3]), .A5(n322), .Y(
        n318) );
  AO21X1_HVT U264 ( .A1(n17), .A2(n187), .A3(n21), .Y(n322) );
  NOR2X0_HVT U265 ( .A1(n70), .A2(n35), .Y(n21) );
  AND2X1_HVT U266 ( .A1(n27), .A2(n29), .Y(n255) );
  NAND2X0_HVT U267 ( .A1(in[1]), .A2(n87), .Y(n29) );
  MUX21X1_HVT U268 ( .A1(n323), .A2(n324), .S0(in[5]), .Y(n316) );
  AO221X1_HVT U269 ( .A1(n20), .A2(n325), .A3(n13), .A4(n326), .A5(n327), .Y(
        n324) );
  AO22X1_HVT U270 ( .A1(n214), .A2(n14), .A3(n157), .A4(n17), .Y(n327) );
  INVX0_HVT U271 ( .A(n254), .Y(n157) );
  AND2X1_HVT U272 ( .A1(n187), .A2(n161), .Y(n214) );
  NAND2X0_HVT U273 ( .A1(n143), .A2(n203), .Y(n161) );
  NAND2X0_HVT U274 ( .A1(n328), .A2(in[1]), .Y(n187) );
  NAND2X0_HVT U275 ( .A1(n145), .A2(n30), .Y(n326) );
  NAND2X0_HVT U276 ( .A1(n61), .A2(n93), .Y(n325) );
  NAND4X0_HVT U277 ( .A1(n114), .A2(n200), .A3(n329), .A4(n330), .Y(n323) );
  OA22X1_HVT U278 ( .A1(n321), .A2(n35), .A3(n15), .A4(n92), .Y(n330) );
  AND2X1_HVT U279 ( .A1(n26), .A2(n201), .Y(n321) );
  NAND2X0_HVT U280 ( .A1(n249), .A2(n203), .Y(n201) );
  INVX0_HVT U281 ( .A(n135), .Y(n249) );
  NAND2X0_HVT U282 ( .A1(n168), .A2(n20), .Y(n329) );
  AND2X1_HVT U283 ( .A1(n86), .A2(n98), .Y(n168) );
  OR2X1_HVT U284 ( .A1(n50), .A2(n92), .Y(n200) );
  NAND2X0_HVT U285 ( .A1(n234), .A2(n17), .Y(n114) );
  INVX0_HVT U286 ( .A(n30), .Y(n234) );
  NAND2X0_HVT U287 ( .A1(n203), .A2(n331), .Y(n30) );
  MUX21X1_HVT U288 ( .A1(n332), .A2(n333), .S0(in[5]), .Y(n315) );
  AO221X1_HVT U289 ( .A1(n63), .A2(n17), .A3(n235), .A4(n20), .A5(n334), .Y(
        n333) );
  AO22X1_HVT U290 ( .A1(n311), .A2(n14), .A3(n94), .A4(n13), .Y(n334) );
  INVX0_HVT U291 ( .A(n265), .Y(n311) );
  NAND2X0_HVT U292 ( .A1(n93), .A2(n27), .Y(n265) );
  NAND2X0_HVT U293 ( .A1(in[1]), .A2(n154), .Y(n93) );
  INVX0_HVT U294 ( .A(n53), .Y(n235) );
  NAND2X0_HVT U295 ( .A1(n71), .A2(n254), .Y(n53) );
  NAND2X0_HVT U296 ( .A1(in[1]), .A2(n331), .Y(n71) );
  INVX0_HVT U297 ( .A(n148), .Y(n63) );
  NAND2X0_HVT U298 ( .A1(n15), .A2(n86), .Y(n148) );
  NAND2X0_HVT U299 ( .A1(in[1]), .A2(n18), .Y(n86) );
  AO221X1_HVT U300 ( .A1(n335), .A2(n14), .A3(n17), .A4(n27), .A5(n336), .Y(
        n332) );
  AO22X1_HVT U301 ( .A1(n337), .A2(n13), .A3(n137), .A4(n20), .Y(n336) );
  AND2X1_HVT U302 ( .A1(n15), .A2(n194), .Y(n137) );
  NAND2X0_HVT U303 ( .A1(in[1]), .A2(n61), .Y(n194) );
  INVX0_HVT U304 ( .A(n82), .Y(n337) );
  NAND2X0_HVT U305 ( .A1(n142), .A2(n98), .Y(n82) );
  NAND2X0_HVT U306 ( .A1(in[4]), .A2(n203), .Y(n98) );
  NAND2X0_HVT U307 ( .A1(n143), .A2(in[1]), .Y(n142) );
  NAND2X0_HVT U308 ( .A1(n135), .A2(n203), .Y(n27) );
  AND2X1_HVT U309 ( .A1(n94), .A2(n50), .Y(n335) );
  NAND2X0_HVT U310 ( .A1(in[1]), .A2(n135), .Y(n50) );
  NAND2X0_HVT U311 ( .A1(in[3]), .A2(n87), .Y(n135) );
  AO221X1_HVT U312 ( .A1(n338), .A2(n13), .A3(n232), .A4(n17), .A5(n339), .Y(
        n314) );
  AO21X1_HVT U313 ( .A1(n295), .A2(n20), .A3(n340), .Y(n339) );
  MUX21X1_HVT U314 ( .A1(n341), .A2(n342), .S0(in[5]), .Y(n340) );
  AO222X1_HVT U315 ( .A1(n13), .A2(n203), .A3(n253), .A4(in[2]), .A5(n14), 
        .A6(n143), .Y(n342) );
  INVX0_HVT U316 ( .A(n154), .Y(n143) );
  NAND2X0_HVT U317 ( .A1(in[4]), .A2(n331), .Y(n154) );
  INVX0_HVT U318 ( .A(n92), .Y(n14) );
  INVX0_HVT U319 ( .A(n72), .Y(n253) );
  NAND2X0_HVT U320 ( .A1(in[3]), .A2(n203), .Y(n72) );
  OAI22X1_HVT U321 ( .A1(n274), .A2(n92), .A3(n26), .A4(n35), .Y(n341) );
  NAND2X0_HVT U322 ( .A1(in[7]), .A2(n57), .Y(n92) );
  NAND2X0_HVT U323 ( .A1(n70), .A2(n26), .Y(n274) );
  NAND2X0_HVT U324 ( .A1(in[1]), .A2(in[3]), .Y(n26) );
  NAND2X0_HVT U325 ( .A1(n203), .A2(n61), .Y(n70) );
  INVX0_HVT U326 ( .A(n62), .Y(n20) );
  NAND2X0_HVT U327 ( .A1(in[2]), .A2(n118), .Y(n62) );
  INVX0_HVT U328 ( .A(n99), .Y(n295) );
  NAND2X0_HVT U329 ( .A1(in[1]), .A2(n15), .Y(n99) );
  INVX0_HVT U330 ( .A(n36), .Y(n17) );
  NAND2X0_HVT U331 ( .A1(n57), .A2(n118), .Y(n36) );
  INVX0_HVT U332 ( .A(in[7]), .Y(n118) );
  INVX0_HVT U333 ( .A(in[2]), .Y(n57) );
  INVX0_HVT U334 ( .A(n56), .Y(n232) );
  NAND2X0_HVT U335 ( .A1(n254), .A2(n145), .Y(n56) );
  NAND2X0_HVT U336 ( .A1(n285), .A2(in[1]), .Y(n145) );
  INVX0_HVT U337 ( .A(n15), .Y(n285) );
  NAND2X0_HVT U338 ( .A1(n94), .A2(n203), .Y(n254) );
  INVX0_HVT U339 ( .A(n18), .Y(n94) );
  NAND2X0_HVT U340 ( .A1(n15), .A2(n61), .Y(n18) );
  NAND2X0_HVT U341 ( .A1(in[3]), .A2(in[4]), .Y(n15) );
  INVX0_HVT U342 ( .A(n35), .Y(n13) );
  NAND2X0_HVT U343 ( .A1(in[7]), .A2(in[2]), .Y(n35) );
  INVX0_HVT U344 ( .A(n88), .Y(n338) );
  NAND2X0_HVT U345 ( .A1(n328), .A2(n203), .Y(n88) );
  INVX0_HVT U346 ( .A(in[1]), .Y(n203) );
  INVX0_HVT U347 ( .A(n61), .Y(n328) );
  NAND2X0_HVT U348 ( .A1(n87), .A2(n331), .Y(n61) );
  INVX0_HVT U349 ( .A(in[3]), .Y(n331) );
  INVX0_HVT U350 ( .A(in[4]), .Y(n87) );
endmodule

