
module inv_sbox_4 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n196, n197, n198, n199, n200, n201, n202, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649;

  NAND2X0_HVT U1 ( .A1(n302), .A2(n361), .Y(n649) );
  NAND2X0_HVT U3 ( .A1(n302), .A2(n336), .Y(n647) );
  NAND2X0_HVT U4 ( .A1(n648), .A2(n273), .Y(n646) );
  NAND2X0_HVT U5 ( .A1(n646), .A2(n368), .Y(n645) );
  NAND2X0_HVT U8 ( .A1(n273), .A2(n321), .Y(n641) );
  NAND2X0_HVT U9 ( .A1(n349), .A2(n641), .Y(n640) );
  NAND2X0_HVT U10 ( .A1(n323), .A2(n638), .Y(n639) );
  NAND2X0_HVT U11 ( .A1(n262), .A2(n328), .Y(n637) );
  NAND2X0_HVT U12 ( .A1(n375), .A2(n359), .Y(n636) );
  NAND2X0_HVT U13 ( .A1(n371), .A2(n641), .Y(n635) );
  NAND2X0_HVT U15 ( .A1(n366), .A2(n276), .Y(n633) );
  NAND2X0_HVT U19 ( .A1(n276), .A2(n438), .Y(n628) );
  NAND2X0_HVT U25 ( .A1(n336), .A2(n301), .Y(n644) );
  NAND2X0_HVT U32 ( .A1(n361), .A2(n378), .Y(n616) );
  NAND2X0_HVT U35 ( .A1(n641), .A2(n439), .Y(n613) );
  NAND2X0_HVT U38 ( .A1(n360), .A2(n262), .Y(n610) );
  NAND2X0_HVT U42 ( .A1(n643), .A2(n327), .Y(n606) );
  OA21X1_HVT U53 ( .A1(n382), .A2(n598), .A3(n409), .Y(n596) );
  MUX41X1_HVT U56 ( .A1(n421), .A3(n312), .A2(n407), .A4(n594), .S0(n353), 
        .S1(n300), .Y(n593) );
  MUX41X1_HVT U62 ( .A1(n587), .A3(n593), .A2(n591), .A4(n595), .S0(n281), 
        .S1(n364), .Y(n586) );
  MUX41X1_HVT U65 ( .A1(n401), .A3(n403), .A2(n402), .A4(n610), .S0(n353), 
        .S1(n357), .Y(n583) );
  NAND2X0_HVT U66 ( .A1(n375), .A2(n254), .Y(n582) );
  MUX41X1_HVT U67 ( .A1(n398), .A3(n422), .A2(n400), .A4(n582), .S0(n357), 
        .S1(n354), .Y(n581) );
  MUX41X1_HVT U68 ( .A1(n398), .A3(n302), .A2(n399), .A4(n348), .S0(n352), 
        .S1(n332), .Y(n580) );
  MUX41X1_HVT U71 ( .A1(n643), .A3(n346), .A2(n637), .A4(n394), .S0(n352), 
        .S1(n381), .Y(n578) );
  NAND2X0_HVT U72 ( .A1(n221), .A2(n642), .Y(n577) );
  MUX41X1_HVT U73 ( .A1(n621), .A3(n577), .A2(n423), .A4(n359), .S0(n357), 
        .S1(n292), .Y(n576) );
  MUX41X1_HVT U74 ( .A1(n639), .A3(n412), .A2(n314), .A4(n268), .S0(n353), 
        .S1(n381), .Y(n575) );
  MUX41X1_HVT U78 ( .A1(n572), .A3(n576), .A2(n575), .A4(n578), .S0(n281), 
        .S1(n364), .Y(n571) );
  MUX41X1_HVT U79 ( .A1(n410), .A3(n630), .A2(n318), .A4(n631), .S0(n353), 
        .S1(n380), .Y(n570) );
  MUX41X1_HVT U80 ( .A1(n425), .A3(n421), .A2(n640), .A4(n316), .S0(n352), 
        .S1(n358), .Y(n569) );
  NAND2X0_HVT U81 ( .A1(n328), .A2(n642), .Y(n568) );
  AND2X1_HVT U82 ( .A1(n643), .A2(n369), .Y(n567) );
  MUX41X1_HVT U83 ( .A1(n567), .A3(n411), .A2(n315), .A4(n568), .S0(n352), 
        .S1(n332), .Y(n566) );
  MUX41X1_HVT U84 ( .A1(n343), .A3(n410), .A2(n426), .A4(n623), .S0(n353), 
        .S1(n381), .Y(n565) );
  MUX41X1_HVT U85 ( .A1(n565), .A3(n569), .A2(n566), .A4(n570), .S0(n281), 
        .S1(n364), .Y(n564) );
  MUX41X1_HVT U88 ( .A1(n400), .A3(n385), .A2(n618), .A4(n602), .S0(n352), 
        .S1(n381), .Y(n562) );
  NAND2X0_HVT U89 ( .A1(n262), .A2(n437), .Y(n561) );
  MUX41X1_HVT U90 ( .A1(n345), .A3(n642), .A2(n601), .A4(n561), .S0(n352), 
        .S1(n380), .Y(n560) );
  NAND2X0_HVT U100 ( .A1(n262), .A2(n436), .Y(n550) );
  MUX41X1_HVT U101 ( .A1(n430), .A3(n636), .A2(n413), .A4(n550), .S0(n358), 
        .S1(n350), .Y(n549) );
  AND2X1_HVT U104 ( .A1(n642), .A2(n368), .Y(n547) );
  MUX41X1_HVT U105 ( .A1(n634), .A3(n431), .A2(n568), .A4(n547), .S0(n353), 
        .S1(n380), .Y(n546) );
  MUX41X1_HVT U107 ( .A1(n430), .A3(n369), .A2(n545), .A4(n391), .S0(n352), 
        .S1(n381), .Y(n544) );
  MUX41X1_HVT U108 ( .A1(n268), .A3(n221), .A2(n407), .A4(n303), .S0(n353), 
        .S1(n380), .Y(n543) );
  MUX41X1_HVT U109 ( .A1(n429), .A3(n385), .A2(n426), .A4(n419), .S0(n352), 
        .S1(n380), .Y(n542) );
  MUX41X1_HVT U110 ( .A1(n542), .A3(n544), .A2(n543), .A4(n546), .S0(n281), 
        .S1(n238), .Y(n541) );
  AO21X1_HVT U112 ( .A1(n416), .A2(n358), .A3(n624), .Y(n539) );
  NAND2X0_HVT U114 ( .A1(n349), .A2(n642), .Y(n537) );
  MUX41X1_HVT U115 ( .A1(n537), .A3(n637), .A2(n416), .A4(n369), .S0(n357), 
        .S1(n296), .Y(n536) );
  MUX41X1_HVT U116 ( .A1(n415), .A3(n410), .A2(n385), .A4(n633), .S0(n351), 
        .S1(n381), .Y(n535) );
  NAND2X0_HVT U118 ( .A1(n378), .A2(n302), .Y(n533) );
  MUX41X1_HVT U119 ( .A1(n432), .A3(n534), .A2(n285), .A4(n533), .S0(n351), 
        .S1(n381), .Y(n532) );
  MUX41X1_HVT U122 ( .A1(n420), .A3(n339), .A2(n602), .A4(n424), .S0(n351), 
        .S1(n380), .Y(n530) );
  MUX41X1_HVT U124 ( .A1(n341), .A3(n529), .A2(n625), .A4(n337), .S0(n358), 
        .S1(n351), .Y(n528) );
  AOI21X1_HVT U127 ( .A1(n356), .A2(n524), .A3(n392), .Y(n525) );
  NAND2X0_HVT U129 ( .A1(n355), .A2(n348), .Y(n522) );
  MUX41X1_HVT U130 ( .A1(n522), .A3(n523), .A2(n526), .A4(n525), .S0(n357), 
        .S1(n238), .Y(n521) );
  AND2X1_HVT U131 ( .A1(n254), .A2(n378), .Y(n520) );
  MUX41X1_HVT U132 ( .A1(n389), .A3(n520), .A2(n434), .A4(n398), .S0(n357), 
        .S1(n292), .Y(n519) );
  MUX41X1_HVT U133 ( .A1(n435), .A3(n391), .A2(n594), .A4(n390), .S0(n358), 
        .S1(n350), .Y(n518) );
  MUX41X1_HVT U136 ( .A1(n599), .A3(n550), .A2(n516), .A4(n396), .S0(n355), 
        .S1(n380), .Y(n515) );
  MUX41X1_HVT U137 ( .A1(n641), .A3(n619), .A2(n623), .A4(n428), .S0(n358), 
        .S1(n350), .Y(n514) );
  MUX41X1_HVT U139 ( .A1(n513), .A3(n517), .A2(n521), .A4(n527), .S0(n281), 
        .S1(n282), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n314), .A3(n340), .A2(n406), .A4(n637), .S0(n358), 
        .S1(n296), .Y(n512) );
  NAND2X0_HVT U141 ( .A1(n366), .A2(n378), .Y(n511) );
  MUX41X1_HVT U143 ( .A1(n437), .A3(n417), .A2(n628), .A4(n625), .S0(n354), 
        .S1(n297), .Y(n509) );
  MUX41X1_HVT U145 ( .A1(n617), .A3(n431), .A2(n508), .A4(n568), .S0(n356), 
        .S1(n297), .Y(n507) );
  OA21X1_HVT U153 ( .A1(n386), .A2(n259), .A3(n395), .Y(n499) );
  MUX41X1_HVT U155 ( .A1(n406), .A3(n637), .A2(n629), .A4(n408), .S0(n354), 
        .S1(n297), .Y(n497) );
  NAND2X0_HVT U159 ( .A1(n493), .A2(n492), .Y(n494) );
  NAND2X0_HVT U163 ( .A1(n375), .A2(n437), .Y(n488) );
  NAND2X0_HVT U166 ( .A1(n638), .A2(n484), .Y(n485) );
  MUX41X1_HVT U172 ( .A1(n561), .A3(n479), .A2(n338), .A4(n626), .S0(n354), 
        .S1(n297), .Y(n478) );
  MUX41X1_HVT U174 ( .A1(n427), .A3(n594), .A2(n435), .A4(n327), .S0(n354), 
        .S1(n297), .Y(n476) );
  NAND2X0_HVT U177 ( .A1(n272), .A2(n302), .Y(n474) );
  MUX41X1_HVT U178 ( .A1(n342), .A3(n474), .A2(n346), .A4(n604), .S0(n354), 
        .S1(n297), .Y(n473) );
  AND2X1_HVT U179 ( .A1(n643), .A2(n367), .Y(n472) );
  AND2X1_HVT U185 ( .A1(n439), .A2(n378), .Y(n466) );
  OA21X1_HVT U189 ( .A1(n410), .A2(n291), .A3(n588), .Y(n462) );
  NAND2X0_HVT U191 ( .A1(n259), .A2(n397), .Y(n460) );
  AND2X1_HVT U192 ( .A1(n412), .A2(n458), .Y(n459) );
  NAND2X0_HVT U194 ( .A1(n606), .A2(n458), .Y(n456) );
  NAND2X0_HVT U198 ( .A1(n375), .A2(n439), .Y(n638) );
  NAND2X0_HVT U200 ( .A1(n367), .A2(n378), .Y(n524) );
  AO21X1_HVT U204 ( .A1(n221), .A2(n324), .A3(n259), .Y(n484) );
  NAND2X0_HVT U207 ( .A1(n262), .A2(n346), .Y(n588) );
  NAND2X0_HVT U2 ( .A1(n408), .A2(n196), .Y(n197) );
  NAND2X0_HVT U6 ( .A1(n399), .A2(n358), .Y(n198) );
  NAND2X0_HVT U7 ( .A1(n197), .A2(n198), .Y(n597) );
  INVX0_HVT U14 ( .A(n358), .Y(n196) );
  INVX1_HVT U16 ( .A(n621), .Y(n408) );
  MUX21X2_HVT U17 ( .A1(n589), .A2(n590), .S0(n199), .Y(n587) );
  IBUFFX16_HVT U18 ( .A(n355), .Y(n199) );
  OR2X2_HVT U20 ( .A1(n310), .A2(n388), .Y(n594) );
  NAND2X0_HVT U21 ( .A1(n564), .A2(n256), .Y(n257) );
  MUX41X1_HVT U22 ( .A1(n583), .A3(n580), .A2(n584), .A4(n581), .S0(n365), 
        .S1(n364), .Y(n579) );
  NAND2X0_HVT U23 ( .A1(n548), .A2(n200), .Y(n201) );
  NAND2X0_HVT U24 ( .A1(n555), .A2(n222), .Y(n202) );
  NAND2X0_HVT U26 ( .A1(n201), .A2(n202), .Y(out[2]) );
  INVX0_HVT U27 ( .A(n222), .Y(n200) );
  INVX1_HVT U28 ( .A(n236), .Y(n222) );
  NAND2X0_HVT U29 ( .A1(n359), .A2(n218), .Y(n219) );
  NAND2X0_HVT U30 ( .A1(n366), .A2(n262), .Y(n220) );
  NAND2X0_HVT U31 ( .A1(n219), .A2(n220), .Y(n627) );
  IBUFFX2_HVT U33 ( .A(n262), .Y(n218) );
  INVX1_HVT U34 ( .A(n250), .Y(n262) );
  INVX0_HVT U36 ( .A(n627), .Y(n268) );
  AO21X1_HVT U37 ( .A1(n588), .A2(n357), .A3(n627), .Y(n589) );
  OA21X1_HVT U39 ( .A1(n387), .A2(n291), .A3(n627), .Y(n573) );
  MUX21X1_HVT U40 ( .A1(n418), .A2(n341), .S0(n297), .Y(n457) );
  NBUFFX8_HVT U41 ( .A(n300), .Y(n297) );
  MUX21X2_HVT U43 ( .A1(n372), .A2(n360), .S0(n276), .Y(n337) );
  INVX1_HVT U44 ( .A(n337), .Y(n625) );
  NBUFFX2_HVT U45 ( .A(n312), .Y(n221) );
  INVX0_HVT U46 ( .A(n311), .Y(n312) );
  NBUFFX16_HVT U47 ( .A(n335), .Y(n362) );
  MUX21X1_HVT U48 ( .A1(n346), .A2(n362), .S0(n375), .Y(n479) );
  INVX1_HVT U49 ( .A(in[5]), .Y(n224) );
  MUX21X1_HVT U50 ( .A1(n405), .A2(n592), .S0(n344), .Y(n591) );
  MUX21X2_HVT U51 ( .A1(n594), .A2(n337), .S0(n278), .Y(n590) );
  IBUFFX2_HVT U52 ( .A(n347), .Y(n348) );
  INVX1_HVT U54 ( .A(n382), .Y(n300) );
  INVX0_HVT U55 ( .A(n347), .Y(n349) );
  MUX41X1_HVT U57 ( .A1(n510), .A3(n512), .A2(n507), .A4(n509), .S0(n223), 
        .S1(n224), .Y(n506) );
  IBUFFX16_HVT U58 ( .A(n363), .Y(n223) );
  NAND2X0_HVT U59 ( .A1(n558), .A2(n225), .Y(n226) );
  NAND2X0_HVT U60 ( .A1(n557), .A2(n235), .Y(n227) );
  NAND2X0_HVT U61 ( .A1(n226), .A2(n227), .Y(n556) );
  INVX0_HVT U63 ( .A(n235), .Y(n225) );
  MUX21X1_HVT U64 ( .A1(n394), .A2(n366), .S0(n293), .Y(n557) );
  IBUFFX2_HVT U69 ( .A(n355), .Y(n235) );
  NAND2X0_HVT U70 ( .A1(n231), .A2(n228), .Y(n229) );
  NAND2X0_HVT U75 ( .A1(n369), .A2(n272), .Y(n230) );
  NAND2X0_HVT U76 ( .A1(n229), .A2(n230), .Y(n269) );
  IBUFFX2_HVT U77 ( .A(n272), .Y(n228) );
  INVX1_HVT U86 ( .A(n377), .Y(n272) );
  INVX0_HVT U87 ( .A(n269), .Y(n607) );
  INVX2_HVT U91 ( .A(n278), .Y(n293) );
  INVX0_HVT U92 ( .A(n326), .Y(n231) );
  IBUFFX2_HVT U93 ( .A(n361), .Y(n326) );
  INVX2_HVT U94 ( .A(n372), .Y(n313) );
  INVX1_HVT U95 ( .A(n632), .Y(n311) );
  AO21X1_HVT U96 ( .A1(n373), .A2(n313), .A3(n259), .Y(n458) );
  MUX21X1_HVT U97 ( .A1(n607), .A2(n423), .S0(n278), .Y(n463) );
  NAND2X0_HVT U98 ( .A1(n370), .A2(n232), .Y(n233) );
  NAND2X0_HVT U99 ( .A1(n559), .A2(n239), .Y(n234) );
  NAND2X0_HVT U102 ( .A1(n233), .A2(n234), .Y(n558) );
  INVX0_HVT U103 ( .A(n239), .Y(n232) );
  IBUFFX16_HVT U106 ( .A(n282), .Y(n236) );
  IBUFFX2_HVT U111 ( .A(n276), .Y(n239) );
  MUX21X1_HVT U113 ( .A1(n310), .A2(n345), .S0(n237), .Y(n481) );
  IBUFFX16_HVT U117 ( .A(n275), .Y(n237) );
  INVX1_HVT U120 ( .A(n614), .Y(n412) );
  NBUFFX2_HVT U121 ( .A(n265), .Y(n238) );
  MUX41X1_HVT U123 ( .A1(n456), .A3(n460), .A2(n457), .A4(n459), .S0(n265), 
        .S1(n240), .Y(n455) );
  MUX41X1_HVT U125 ( .A1(n455), .A3(n467), .A2(n461), .A4(n470), .S0(n282), 
        .S1(n281), .Y(out[7]) );
  INVX0_HVT U126 ( .A(n363), .Y(n265) );
  IBUFFX2_HVT U128 ( .A(n352), .Y(n240) );
  NAND2X2_HVT U134 ( .A1(n373), .A2(n370), .Y(n642) );
  XNOR2X2_HVT U135 ( .A1(n345), .A2(n273), .Y(n611) );
  IBUFFX2_HVT U138 ( .A(n363), .Y(n364) );
  INVX2_HVT U142 ( .A(n382), .Y(n380) );
  MUX41X1_HVT U144 ( .A1(n616), .A3(n402), .A2(n600), .A4(n312), .S0(n380), 
        .S1(n355), .Y(n551) );
  MUX41X1_HVT U146 ( .A1(n422), .A3(n408), .A2(n635), .A4(n428), .S0(n380), 
        .S1(n353), .Y(n554) );
  INVX1_HVT U147 ( .A(n453), .Y(n422) );
  NAND2X0_HVT U148 ( .A1(n541), .A2(n241), .Y(n242) );
  NAND2X0_HVT U149 ( .A1(n531), .A2(n244), .Y(n243) );
  NAND2X0_HVT U150 ( .A1(n242), .A2(n243), .Y(out[3]) );
  INVX8_HVT U151 ( .A(n244), .Y(n241) );
  INVX2_HVT U152 ( .A(n251), .Y(n244) );
  MUX41X1_HVT U154 ( .A1(n345), .A3(n349), .A2(n612), .A4(n328), .S0(n245), 
        .S1(n299), .Y(n477) );
  IBUFFX16_HVT U156 ( .A(n354), .Y(n245) );
  MUX21X2_HVT U157 ( .A1(n540), .A2(n539), .S0(n246), .Y(n538) );
  IBUFFX16_HVT U158 ( .A(n356), .Y(n246) );
  MUX41X1_HVT U160 ( .A1(n429), .A3(n553), .A2(n620), .A4(n414), .S0(n247), 
        .S1(n381), .Y(n552) );
  IBUFFX16_HVT U161 ( .A(n353), .Y(n247) );
  MUX21X1_HVT U162 ( .A1(n360), .A2(n310), .S0(n376), .Y(n605) );
  INVX2_HVT U164 ( .A(n301), .Y(n302) );
  MUX41X1_HVT U165 ( .A1(n552), .A3(n554), .A2(n549), .A4(n551), .S0(n364), 
        .S1(n365), .Y(n548) );
  IBUFFX2_HVT U167 ( .A(n612), .Y(n413) );
  NBUFFX16_HVT U168 ( .A(n296), .Y(n351) );
  INVX2_HVT U169 ( .A(n298), .Y(n296) );
  INVX2_HVT U170 ( .A(n379), .Y(n298) );
  INVX0_HVT U171 ( .A(n369), .Y(n438) );
  MUX21X1_HVT U173 ( .A1(n437), .A2(n438), .S0(n248), .Y(n534) );
  IBUFFX16_HVT U175 ( .A(n273), .Y(n248) );
  MUX21X2_HVT U176 ( .A1(n346), .A2(n437), .S0(n277), .Y(n620) );
  INVX1_HVT U180 ( .A(n349), .Y(n346) );
  INVX0_HVT U181 ( .A(n451), .Y(n424) );
  INVX1_HVT U182 ( .A(n605), .Y(n417) );
  IBUFFX16_HVT U183 ( .A(in[1]), .Y(n363) );
  MUX41X1_HVT U184 ( .A1(n388), .A3(n343), .A2(n427), .A4(n407), .S0(n351), 
        .S1(n332), .Y(n563) );
  INVX1_HVT U186 ( .A(n447), .Y(n427) );
  INVX1_HVT U187 ( .A(n622), .Y(n407) );
  INVX0_HVT U188 ( .A(n632), .Y(n439) );
  INVX0_HVT U190 ( .A(n632), .Y(n327) );
  XNOR2X2_HVT U193 ( .A1(n362), .A2(n301), .Y(n632) );
  MUX21X1_HVT U195 ( .A1(n519), .A2(n518), .S0(n363), .Y(n517) );
  MUX41X1_HVT U196 ( .A1(n556), .A3(n560), .A2(n562), .A4(n563), .S0(n364), 
        .S1(n281), .Y(n555) );
  IBUFFX2_HVT U197 ( .A(n382), .Y(n381) );
  INVX0_HVT U199 ( .A(in[0]), .Y(n249) );
  INVX1_HVT U201 ( .A(n249), .Y(n250) );
  IBUFFX16_HVT U202 ( .A(n331), .Y(n251) );
  INVX2_HVT U203 ( .A(n274), .Y(n275) );
  MUX21X2_HVT U205 ( .A1(n316), .A2(n406), .S0(n252), .Y(n592) );
  IBUFFX16_HVT U206 ( .A(n356), .Y(n252) );
  MUX21X2_HVT U208 ( .A1(n268), .A2(n585), .S0(n344), .Y(n584) );
  INVX0_HVT U209 ( .A(n451), .Y(n253) );
  MUX21X1_HVT U210 ( .A1(n253), .A2(n384), .S0(n293), .Y(n574) );
  INVX1_HVT U211 ( .A(n274), .Y(n277) );
  INVX1_HVT U212 ( .A(n274), .Y(n276) );
  INVX2_HVT U213 ( .A(n374), .Y(n274) );
  INVX1_HVT U214 ( .A(n377), .Y(n273) );
  NBUFFX2_HVT U215 ( .A(n336), .Y(n254) );
  INVX1_HVT U216 ( .A(n335), .Y(n336) );
  INVX1_HVT U217 ( .A(n331), .Y(n282) );
  OR2X1_HVT U218 ( .A1(n274), .A2(n347), .Y(n643) );
  INVX1_HVT U219 ( .A(n377), .Y(n373) );
  MUX41X1_HVT U220 ( .A1(n388), .A3(n315), .A2(n391), .A4(n324), .S0(n255), 
        .S1(n286), .Y(n469) );
  IBUFFX16_HVT U221 ( .A(n289), .Y(n255) );
  NAND2X0_HVT U222 ( .A1(n571), .A2(n282), .Y(n258) );
  NAND2X0_HVT U223 ( .A1(n257), .A2(n258), .Y(out[1]) );
  IBUFFX2_HVT U224 ( .A(n282), .Y(n256) );
  INVX0_HVT U225 ( .A(n606), .Y(n391) );
  MUX41X1_HVT U226 ( .A1(n489), .A3(n483), .A2(n491), .A4(n487), .S0(n365), 
        .S1(n238), .Y(n482) );
  INVX2_HVT U227 ( .A(n365), .Y(n281) );
  IBUFFX2_HVT U228 ( .A(n377), .Y(n375) );
  INVX0_HVT U229 ( .A(n377), .Y(n374) );
  INVX0_HVT U230 ( .A(in[0]), .Y(n377) );
  MUX21X1_HVT U231 ( .A1(n360), .A2(n327), .S0(n262), .Y(n609) );
  AO21X1_HVT U232 ( .A1(n262), .A2(n323), .A3(n259), .Y(n492) );
  INVX0_HVT U233 ( .A(n298), .Y(n264) );
  INVX0_HVT U234 ( .A(n321), .Y(n290) );
  INVX0_HVT U235 ( .A(n603), .Y(n418) );
  INVX1_HVT U236 ( .A(in[5]), .Y(n365) );
  INVX1_HVT U237 ( .A(n351), .Y(n263) );
  INVX0_HVT U238 ( .A(n351), .Y(n289) );
  INVX0_HVT U239 ( .A(n637), .Y(n383) );
  INVX1_HVT U240 ( .A(n347), .Y(n323) );
  INVX1_HVT U241 ( .A(n649), .Y(n347) );
  INVX1_HVT U242 ( .A(n299), .Y(n278) );
  INVX1_HVT U243 ( .A(n299), .Y(n259) );
  INVX1_HVT U244 ( .A(n286), .Y(n332) );
  NBUFFX2_HVT U245 ( .A(n300), .Y(n299) );
  INVX1_HVT U246 ( .A(n299), .Y(n286) );
  INVX0_HVT U247 ( .A(n357), .Y(n291) );
  MUX21X2_HVT U248 ( .A1(n424), .A2(n605), .S0(n259), .Y(n495) );
  MUX21X1_HVT U249 ( .A1(n359), .A2(n438), .S0(n378), .Y(n451) );
  MUX21X2_HVT U250 ( .A1(n573), .A2(n574), .S0(n263), .Y(n572) );
  MUX41X1_HVT U251 ( .A1(n535), .A3(n538), .A2(n532), .A4(n536), .S0(n281), 
        .S1(n363), .Y(n531) );
  MUX21X2_HVT U252 ( .A1(n500), .A2(n499), .S0(n263), .Y(n498) );
  NAND2X0_HVT U253 ( .A1(n466), .A2(n291), .Y(n260) );
  NAND2X0_HVT U254 ( .A1(n425), .A2(n293), .Y(n261) );
  NAND2X0_HVT U255 ( .A1(n260), .A2(n261), .Y(n465) );
  INVX1_HVT U256 ( .A(n450), .Y(n425) );
  IBUFFX2_HVT U257 ( .A(n250), .Y(n378) );
  MUX41X1_HVT U258 ( .A1(n268), .A3(n611), .A2(n488), .A4(n640), .S0(n263), 
        .S1(n286), .Y(n487) );
  MUX41X1_HVT U259 ( .A1(n417), .A3(n421), .A2(n268), .A4(n606), .S0(n358), 
        .S1(n264), .Y(n468) );
  NAND2X0_HVT U260 ( .A1(n473), .A2(n265), .Y(n266) );
  NAND2X0_HVT U261 ( .A1(n471), .A2(n363), .Y(n267) );
  NAND2X0_HVT U262 ( .A1(n266), .A2(n267), .Y(n470) );
  MUX41X1_HVT U263 ( .A1(n463), .A3(n464), .A2(n462), .A4(n465), .S0(in[1]), 
        .S1(n296), .Y(n461) );
  NAND2X0_HVT U264 ( .A1(n468), .A2(n363), .Y(n270) );
  NAND2X0_HVT U265 ( .A1(n469), .A2(n265), .Y(n271) );
  NAND2X0_HVT U266 ( .A1(n270), .A2(n271), .Y(n467) );
  INVX1_HVT U267 ( .A(n289), .Y(n292) );
  MUX21X1_HVT U268 ( .A1(n367), .A2(n323), .S0(n250), .Y(n322) );
  INVX0_HVT U269 ( .A(n322), .Y(n604) );
  MUX41X1_HVT U270 ( .A1(n490), .A3(n613), .A2(n403), .A4(n322), .S0(n263), 
        .S1(n259), .Y(n489) );
  MUX41X1_HVT U271 ( .A1(n603), .A3(n472), .A2(n383), .A4(n616), .S0(n263), 
        .S1(n278), .Y(n471) );
  XNOR2X1_HVT U272 ( .A1(n327), .A2(n276), .Y(n602) );
  INVX1_HVT U273 ( .A(n449), .Y(n315) );
  IBUFFX2_HVT U274 ( .A(n602), .Y(n419) );
  NAND2X0_HVT U275 ( .A1(n475), .A2(n331), .Y(n279) );
  NAND2X0_HVT U276 ( .A1(n482), .A2(n282), .Y(n280) );
  NAND2X0_HVT U277 ( .A1(n279), .A2(n280), .Y(out[6]) );
  INVX1_HVT U278 ( .A(n452), .Y(n423) );
  MUX41X1_HVT U279 ( .A1(n478), .A3(n480), .A2(n476), .A4(n477), .S0(n238), 
        .S1(n365), .Y(n475) );
  NAND2X0_HVT U280 ( .A1(n494), .A2(n263), .Y(n283) );
  NAND2X0_HVT U281 ( .A1(n495), .A2(n356), .Y(n284) );
  NAND2X0_HVT U282 ( .A1(n283), .A2(n284), .Y(n491) );
  INVX0_HVT U283 ( .A(n414), .Y(n285) );
  INVX1_HVT U284 ( .A(n611), .Y(n414) );
  IBUFFX2_HVT U285 ( .A(n377), .Y(n376) );
  NAND2X0_HVT U286 ( .A1(n343), .A2(n259), .Y(n287) );
  NAND2X0_HVT U287 ( .A1(n600), .A2(n293), .Y(n288) );
  NAND2X0_HVT U288 ( .A1(n287), .A2(n288), .Y(n464) );
  XNOR2X1_HVT U289 ( .A1(n290), .A2(n273), .Y(n600) );
  MUX41X1_HVT U290 ( .A1(n414), .A3(n315), .A2(n502), .A4(n404), .S0(n291), 
        .S1(n292), .Y(n501) );
  NBUFFX2_HVT U291 ( .A(n632), .Y(n366) );
  NAND2X0_HVT U292 ( .A1(n343), .A2(n332), .Y(n333) );
  NAND2X0_HVT U293 ( .A1(n596), .A2(n356), .Y(n294) );
  INVX0_HVT U294 ( .A(n371), .Y(n310) );
  MUX21X1_HVT U295 ( .A1(n362), .A2(n439), .S0(n275), .Y(n612) );
  NAND2X0_HVT U296 ( .A1(n485), .A2(n289), .Y(n319) );
  MUX21X1_HVT U297 ( .A1(n632), .A2(n362), .S0(n373), .Y(n623) );
  INVX1_HVT U298 ( .A(in[7]), .Y(n331) );
  INVX1_HVT U299 ( .A(n615), .Y(n314) );
  INVX1_HVT U300 ( .A(n454), .Y(n421) );
  INVX1_HVT U301 ( .A(in[3]), .Y(n301) );
  INVX1_HVT U302 ( .A(in[6]), .Y(n335) );
  MUX21X1_HVT U303 ( .A1(n366), .A2(n362), .S0(n299), .Y(n559) );
  NAND2X0_HVT U304 ( .A1(n597), .A2(n289), .Y(n295) );
  NAND2X0_HVT U305 ( .A1(n294), .A2(n295), .Y(n595) );
  INVX1_HVT U306 ( .A(in[4]), .Y(n382) );
  MUX41X1_HVT U307 ( .A1(n338), .A3(n342), .A2(n481), .A4(n341), .S0(n298), 
        .S1(n299), .Y(n480) );
  AO21X2_HVT U308 ( .A1(n332), .A2(n393), .A3(n313), .Y(n504) );
  NAND2X0_HVT U309 ( .A1(n586), .A2(n282), .Y(n329) );
  INVX1_HVT U310 ( .A(n436), .Y(n303) );
  NAND2X0_HVT U311 ( .A1(n434), .A2(n291), .Y(n304) );
  NAND2X0_HVT U312 ( .A1(n389), .A2(n358), .Y(n305) );
  NAND2X0_HVT U313 ( .A1(n304), .A2(n305), .Y(n505) );
  NAND2X0_HVT U314 ( .A1(n504), .A2(n355), .Y(n306) );
  NAND2X0_HVT U315 ( .A1(n505), .A2(n263), .Y(n307) );
  NAND2X0_HVT U316 ( .A1(n306), .A2(n307), .Y(n503) );
  NAND2X0_HVT U317 ( .A1(n506), .A2(n282), .Y(n308) );
  NAND2X0_HVT U318 ( .A1(n496), .A2(n331), .Y(n309) );
  NAND2X0_HVT U319 ( .A1(n308), .A2(n309), .Y(out[5]) );
  INVX0_HVT U320 ( .A(n644), .Y(n437) );
  INVX0_HVT U321 ( .A(n648), .Y(n436) );
  INVX0_HVT U322 ( .A(n645), .Y(n389) );
  MUX21X1_HVT U323 ( .A1(n404), .A2(n324), .S0(n355), .Y(n585) );
  INVX0_HVT U324 ( .A(n389), .Y(n316) );
  INVX0_HVT U325 ( .A(n318), .Y(n617) );
  INVX0_HVT U326 ( .A(n313), .Y(n317) );
  INVX1_HVT U327 ( .A(n325), .Y(n502) );
  MUX21X1_HVT U328 ( .A1(n349), .A2(n439), .S0(n378), .Y(n318) );
  INVX1_HVT U329 ( .A(n441), .Y(n434) );
  MUX41X1_HVT U330 ( .A1(n406), .A3(n433), .A2(n609), .A4(n511), .S0(n263), 
        .S1(n278), .Y(n510) );
  NAND2X0_HVT U331 ( .A1(n486), .A2(n355), .Y(n320) );
  NAND2X0_HVT U332 ( .A1(n319), .A2(n320), .Y(n483) );
  MUX21X1_HVT U333 ( .A1(n622), .A2(n625), .S0(n293), .Y(n486) );
  MUX21X1_HVT U334 ( .A1(n361), .A2(n313), .S0(n272), .Y(n622) );
  MUX21X1_HVT U335 ( .A1(n327), .A2(n436), .S0(n378), .Y(n615) );
  NBUFFX2_HVT U336 ( .A(n644), .Y(n321) );
  NBUFFX2_HVT U337 ( .A(n301), .Y(n359) );
  INVX1_HVT U338 ( .A(n623), .Y(n406) );
  INVX1_HVT U339 ( .A(n388), .Y(n324) );
  MUX21X1_HVT U340 ( .A1(n367), .A2(n326), .S0(n262), .Y(n325) );
  NAND2X0_HVT U341 ( .A1(n359), .A2(n362), .Y(n328) );
  NAND2X0_HVT U342 ( .A1(n579), .A2(n331), .Y(n330) );
  NAND2X0_HVT U343 ( .A1(n329), .A2(n330), .Y(out[0]) );
  NAND2X0_HVT U344 ( .A1(n623), .A2(n382), .Y(n334) );
  NAND2X0_HVT U345 ( .A1(n333), .A2(n334), .Y(n500) );
  INVX1_HVT U346 ( .A(n626), .Y(n404) );
  MUX41X1_HVT U347 ( .A1(n498), .A3(n503), .A2(n497), .A4(n501), .S0(n281), 
        .S1(n363), .Y(n496) );
  NBUFFX2_HVT U348 ( .A(n328), .Y(n372) );
  AND2X1_HVT U349 ( .A1(n643), .A2(n303), .Y(n338) );
  AND2X1_HVT U350 ( .A1(n317), .A2(n633), .Y(n339) );
  NAND2X0_HVT U351 ( .A1(n359), .A2(n361), .Y(n648) );
  MUX21X1_HVT U352 ( .A1(n311), .A2(n436), .S0(n272), .Y(n626) );
  MUX21X1_HVT U353 ( .A1(n360), .A2(n313), .S0(n373), .Y(n618) );
  MUX21X1_HVT U354 ( .A1(n439), .A2(n362), .S0(n272), .Y(n442) );
  MUX21X1_HVT U355 ( .A1(n436), .A2(n438), .S0(n275), .Y(n598) );
  MUX21X1_HVT U356 ( .A1(n312), .A2(n437), .S0(n375), .Y(n614) );
  MUX21X1_HVT U357 ( .A1(n360), .A2(n303), .S0(n275), .Y(n450) );
  MUX21X1_HVT U358 ( .A1(n368), .A2(n370), .S0(n273), .Y(n490) );
  MUX21X1_HVT U359 ( .A1(n345), .A2(n312), .S0(n376), .Y(n447) );
  MUX21X1_HVT U360 ( .A1(n321), .A2(n372), .S0(n277), .Y(n441) );
  MUX21X1_HVT U361 ( .A1(n615), .A2(n339), .S0(n356), .Y(n523) );
  MUX21X1_HVT U362 ( .A1(n362), .A2(n317), .S0(n275), .Y(n545) );
  MUX21X1_HVT U363 ( .A1(n433), .A2(n340), .S0(n355), .Y(n526) );
  MUX21X1_HVT U364 ( .A1(n361), .A2(n312), .S0(n373), .Y(n608) );
  XNOR2X1_HVT U365 ( .A1(n303), .A2(n273), .Y(n340) );
  MUX21X1_HVT U366 ( .A1(n323), .A2(n648), .S0(n275), .Y(n634) );
  MUX21X1_HVT U367 ( .A1(n371), .A2(n303), .S0(n275), .Y(n630) );
  MUX21X1_HVT U368 ( .A1(n360), .A2(n361), .S0(n272), .Y(n603) );
  XOR2X1_HVT U369 ( .A1(n369), .A2(n375), .Y(n601) );
  MUX21X1_HVT U370 ( .A1(n370), .A2(n359), .S0(n277), .Y(n629) );
  AND2X1_HVT U371 ( .A1(n277), .A2(n362), .Y(n341) );
  MUX21X1_HVT U372 ( .A1(n360), .A2(n370), .S0(n373), .Y(n444) );
  MUX21X1_HVT U373 ( .A1(n371), .A2(n361), .S0(n376), .Y(n529) );
  NBUFFX2_HVT U374 ( .A(n300), .Y(n357) );
  NBUFFX2_HVT U375 ( .A(n300), .Y(n358) );
  AND2X1_HVT U376 ( .A1(n438), .A2(n378), .Y(n342) );
  NBUFFX2_HVT U377 ( .A(n335), .Y(n361) );
  NBUFFX2_HVT U378 ( .A(n644), .Y(n367) );
  NBUFFX2_HVT U379 ( .A(n647), .Y(n369) );
  AND2X1_HVT U380 ( .A1(n371), .A2(n262), .Y(n343) );
  MUX21X1_HVT U381 ( .A1(n328), .A2(n367), .S0(n373), .Y(n508) );
  NBUFFX2_HVT U382 ( .A(n647), .Y(n371) );
  MUX21X1_HVT U383 ( .A1(n392), .A2(n607), .S0(n357), .Y(n540) );
  MUX21X1_HVT U384 ( .A1(n528), .A2(n530), .S0(n364), .Y(n527) );
  NBUFFX2_HVT U385 ( .A(n644), .Y(n368) );
  NBUFFX2_HVT U386 ( .A(n647), .Y(n370) );
  NBUFFX2_HVT U387 ( .A(n301), .Y(n360) );
  NBUFFX2_HVT U388 ( .A(n350), .Y(n354) );
  NBUFFX2_HVT U389 ( .A(n379), .Y(n356) );
  NBUFFX2_HVT U390 ( .A(n379), .Y(n355) );
  XNOR2X1_HVT U391 ( .A1(n286), .A2(n351), .Y(n344) );
  NBUFFX2_HVT U392 ( .A(n356), .Y(n352) );
  NBUFFX2_HVT U393 ( .A(n350), .Y(n353) );
  NBUFFX2_HVT U394 ( .A(n379), .Y(n350) );
  MUX21X1_HVT U395 ( .A1(n336), .A2(n437), .S0(n375), .Y(n454) );
  MUX21X1_HVT U396 ( .A1(n367), .A2(n302), .S0(n375), .Y(n553) );
  MUX21X1_HVT U397 ( .A1(n514), .A2(n515), .S0(in[1]), .Y(n513) );
  MUX21X1_HVT U398 ( .A1(n345), .A2(n302), .S0(n276), .Y(n440) );
  MUX21X1_HVT U399 ( .A1(n336), .A2(n348), .S0(n275), .Y(n631) );
  MUX21X1_HVT U400 ( .A1(n348), .A2(n302), .S0(n375), .Y(n493) );
  MUX21X1_HVT U401 ( .A1(n368), .A2(n336), .S0(n376), .Y(n619) );
  XOR2X1_HVT U402 ( .A1(n376), .A2(n254), .Y(n599) );
  MUX21X1_HVT U403 ( .A1(n313), .A2(n254), .S0(n376), .Y(n516) );
  MUX21X1_HVT U404 ( .A1(n302), .A2(n348), .S0(n376), .Y(n446) );
  MUX21X1_HVT U405 ( .A1(n254), .A2(n346), .S0(n272), .Y(n624) );
  MUX21X1_HVT U406 ( .A1(n362), .A2(n302), .S0(n373), .Y(n621) );
  MUX21X1_HVT U407 ( .A1(n302), .A2(n368), .S0(n273), .Y(n445) );
  MUX21X1_HVT U408 ( .A1(n254), .A2(n371), .S0(n277), .Y(n453) );
  MUX21X1_HVT U409 ( .A1(n370), .A2(n254), .S0(n272), .Y(n448) );
  MUX21X1_HVT U410 ( .A1(n360), .A2(n254), .S0(n376), .Y(n443) );
  NBUFFX2_HVT U411 ( .A(in[2]), .Y(n379) );
  MUX21X1_HVT U412 ( .A1(n436), .A2(n361), .S0(n277), .Y(n452) );
  MUX21X1_HVT U413 ( .A1(n360), .A2(n327), .S0(n373), .Y(n449) );
  INVX1_HVT U414 ( .A(n323), .Y(n345) );
  INVX0_HVT U415 ( .A(n616), .Y(n384) );
  INVX0_HVT U416 ( .A(n610), .Y(n385) );
  INVX0_HVT U417 ( .A(n550), .Y(n386) );
  INVX0_HVT U418 ( .A(n511), .Y(n387) );
  INVX0_HVT U419 ( .A(n646), .Y(n388) );
  INVX0_HVT U420 ( .A(n643), .Y(n390) );
  INVX0_HVT U421 ( .A(n642), .Y(n392) );
  INVX0_HVT U422 ( .A(n641), .Y(n393) );
  INVX0_HVT U423 ( .A(n613), .Y(n394) );
  INVX0_HVT U424 ( .A(n635), .Y(n395) );
  INVX0_HVT U425 ( .A(n640), .Y(n396) );
  INVX0_HVT U426 ( .A(n636), .Y(n397) );
  INVX0_HVT U427 ( .A(n634), .Y(n398) );
  INVX0_HVT U428 ( .A(n633), .Y(n399) );
  INVX0_HVT U429 ( .A(n631), .Y(n400) );
  INVX0_HVT U430 ( .A(n630), .Y(n401) );
  INVX0_HVT U431 ( .A(n629), .Y(n402) );
  INVX0_HVT U432 ( .A(n628), .Y(n403) );
  INVX0_HVT U433 ( .A(n624), .Y(n405) );
  INVX0_HVT U434 ( .A(n620), .Y(n409) );
  INVX0_HVT U435 ( .A(n619), .Y(n410) );
  INVX0_HVT U436 ( .A(n618), .Y(n411) );
  INVX0_HVT U437 ( .A(n609), .Y(n415) );
  INVX0_HVT U438 ( .A(n608), .Y(n416) );
  INVX0_HVT U439 ( .A(n639), .Y(n420) );
  INVX0_HVT U440 ( .A(n448), .Y(n426) );
  INVX0_HVT U441 ( .A(n446), .Y(n428) );
  INVX0_HVT U442 ( .A(n445), .Y(n429) );
  INVX0_HVT U443 ( .A(n444), .Y(n430) );
  INVX0_HVT U444 ( .A(n443), .Y(n431) );
  INVX0_HVT U445 ( .A(n493), .Y(n432) );
  INVX0_HVT U446 ( .A(n442), .Y(n433) );
  INVX0_HVT U447 ( .A(n440), .Y(n435) );
endmodule

