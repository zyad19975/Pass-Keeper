
module sbox_6 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n50, n210, n211, n212, n213, n216, n217, n218, n219, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580;

  NAND2X0_HVT U3 ( .A1(n290), .A2(n283), .Y(n578) );
  NAND2X0_HVT U4 ( .A1(n281), .A2(n578), .Y(n577) );
  NAND2X0_HVT U5 ( .A1(n288), .A2(n270), .Y(n575) );
  NAND2X0_HVT U13 ( .A1(n567), .A2(n285), .Y(n568) );
  NAND2X0_HVT U15 ( .A1(n578), .A2(n272), .Y(n565) );
  NAND2X0_HVT U21 ( .A1(n280), .A2(n292), .Y(n559) );
  NAND2X0_HVT U24 ( .A1(n277), .A2(n292), .Y(n557) );
  NAND2X0_HVT U33 ( .A1(n356), .A2(n292), .Y(n548) );
  NAND2X0_HVT U35 ( .A1(n275), .A2(n292), .Y(n546) );
  NAND2X0_HVT U42 ( .A1(n286), .A2(n277), .Y(n539) );
  MUX41X1_HVT U51 ( .A1(n344), .A3(n302), .A2(n319), .A4(n320), .S0(n297), 
        .S1(n264), .Y(n532) );
  NAND2X0_HVT U53 ( .A1(n529), .A2(n538), .Y(n530) );
  NAND2X0_HVT U56 ( .A1(n281), .A2(n525), .Y(n526) );
  MUX41X1_HVT U57 ( .A1(n345), .A3(n561), .A2(n526), .A4(n570), .S0(n299), 
        .S1(n264), .Y(n524) );
  NAND2X0_HVT U58 ( .A1(n285), .A2(n578), .Y(n523) );
  MUX41X1_HVT U59 ( .A1(n258), .A3(n523), .A2(n256), .A4(n318), .S0(n296), 
        .S1(n264), .Y(n522) );
  MUX41X1_HVT U61 ( .A1(n254), .A3(n317), .A2(n316), .A4(n271), .S0(n296), 
        .S1(n264), .Y(n520) );
  NAND2X0_HVT U62 ( .A1(n292), .A2(n283), .Y(n519) );
  MUX41X1_HVT U63 ( .A1(n519), .A3(n309), .A2(n339), .A4(n315), .S0(n296), 
        .S1(n264), .Y(n518) );
  AO21X1_HVT U66 ( .A1(n313), .A2(n266), .A3(n338), .Y(n515) );
  MUX41X1_HVT U68 ( .A1(n311), .A3(n515), .A2(n514), .A4(n516), .S0(n259), 
        .S1(n241), .Y(n513) );
  MUX41X1_HVT U69 ( .A1(n513), .A3(n521), .A2(n517), .A4(n527), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n278), .A2(n508), .Y(n509) );
  MUX41X1_HVT U74 ( .A1(n510), .A3(n555), .A2(n509), .A4(n557), .S0(n261), 
        .S1(n299), .Y(n507) );
  MUX41X1_HVT U77 ( .A1(n572), .A3(n349), .A2(n505), .A4(n348), .S0(n267), 
        .S1(n293), .Y(n504) );
  MUX41X1_HVT U78 ( .A1(n504), .A3(n507), .A2(n506), .A4(n511), .S0(in[0]), 
        .S1(n264), .Y(n503) );
  AND3X1_HVT U80 ( .A1(n283), .A2(n525), .A3(n500), .Y(n501) );
  MUX41X1_HVT U82 ( .A1(n536), .A3(n320), .A2(n303), .A4(n566), .S0(n259), 
        .S1(n296), .Y(n498) );
  AND2X1_HVT U83 ( .A1(n287), .A2(n242), .Y(n497) );
  MUX41X1_HVT U84 ( .A1(n321), .A3(n574), .A2(n564), .A4(n497), .S0(n259), 
        .S1(n297), .Y(n496) );
  NAND2X0_HVT U85 ( .A1(n292), .A2(n359), .Y(n495) );
  MUX41X1_HVT U86 ( .A1(n347), .A3(n495), .A2(n255), .A4(n251), .S0(n259), 
        .S1(n299), .Y(n494) );
  MUX41X1_HVT U87 ( .A1(n494), .A3(n498), .A2(n496), .A4(n499), .S0(in[0]), 
        .S1(n295), .Y(n493) );
  AO21X1_HVT U93 ( .A1(n269), .A2(n487), .A3(n343), .Y(n488) );
  MUX41X1_HVT U96 ( .A1(n303), .A3(n253), .A2(n346), .A4(n485), .S0(n259), 
        .S1(n296), .Y(n484) );
  MUX41X1_HVT U97 ( .A1(n342), .A3(n253), .A2(n290), .A4(n565), .S0(n259), 
        .S1(n299), .Y(n483) );
  NAND2X0_HVT U101 ( .A1(n478), .A2(n477), .Y(n479) );
  MUX41X1_HVT U103 ( .A1(n578), .A3(n312), .A2(n325), .A4(n546), .S0(n259), 
        .S1(n297), .Y(n475) );
  MUX41X1_HVT U105 ( .A1(n324), .A3(n534), .A2(n474), .A4(n341), .S0(n259), 
        .S1(n297), .Y(n473) );
  OA21X1_HVT U109 ( .A1(n332), .A2(n294), .A3(n318), .Y(n470) );
  NAND2X0_HVT U110 ( .A1(n283), .A2(n468), .Y(n469) );
  AND2X1_HVT U115 ( .A1(n286), .A2(n271), .Y(n463) );
  MUX41X1_HVT U116 ( .A1(n568), .A3(n463), .A2(n322), .A4(n550), .S0(n260), 
        .S1(n298), .Y(n462) );
  NAND2X0_HVT U123 ( .A1(n454), .A2(n453), .Y(n455) );
  MUX41X1_HVT U125 ( .A1(n559), .A3(n258), .A2(n311), .A4(n351), .S0(n260), 
        .S1(n298), .Y(n451) );
  AND3X1_HVT U128 ( .A1(n263), .A2(n292), .A3(n242), .Y(n448) );
  MUX41X1_HVT U131 ( .A1(n446), .A3(n448), .A2(n447), .A4(n449), .S0(n266), 
        .S1(n296), .Y(n445) );
  MUX41X1_HVT U132 ( .A1(n445), .A3(n458), .A2(n450), .A4(n464), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  MUX41X1_HVT U136 ( .A1(n251), .A3(n548), .A2(n353), .A4(n545), .S0(n260), 
        .S1(n297), .Y(n441) );
  MUX41X1_HVT U139 ( .A1(n439), .A3(n442), .A2(n441), .A4(n443), .S0(n276), 
        .S1(n295), .Y(n438) );
  AND2X1_HVT U140 ( .A1(n279), .A2(n291), .Y(n437) );
  OA21X1_HVT U144 ( .A1(n306), .A2(n301), .A3(n550), .Y(n433) );
  NAND2X0_HVT U146 ( .A1(n286), .A2(n285), .Y(n508) );
  OA21X1_HVT U151 ( .A1(n541), .A2(n301), .A3(n427), .Y(n428) );
  MUX41X1_HVT U153 ( .A1(n469), .A3(n254), .A2(n282), .A4(n305), .S0(n260), 
        .S1(n297), .Y(n425) );
  AND2X1_HVT U154 ( .A1(n269), .A2(n277), .Y(n424) );
  NAND2X0_HVT U158 ( .A1(n289), .A2(n359), .Y(n420) );
  MUX41X1_HVT U159 ( .A1(n568), .A3(n271), .A2(n420), .A4(n233), .S0(n261), 
        .S1(n296), .Y(n419) );
  MUX41X1_HVT U160 ( .A1(n419), .A3(n425), .A2(n421), .A4(n426), .S0(n276), 
        .S1(n265), .Y(n418) );
  AND2X1_HVT U162 ( .A1(n574), .A2(n508), .Y(n416) );
  MUX41X1_HVT U163 ( .A1(n317), .A3(n416), .A2(n252), .A4(n417), .S0(n262), 
        .S1(n296), .Y(n415) );
  MUX41X1_HVT U165 ( .A1(n559), .A3(n326), .A2(n535), .A4(n414), .S0(n299), 
        .S1(n261), .Y(n413) );
  NAND2X0_HVT U166 ( .A1(n285), .A2(n525), .Y(n412) );
  NAND2X0_HVT U167 ( .A1(n360), .A2(n292), .Y(n411) );
  MUX41X1_HVT U168 ( .A1(n345), .A3(n279), .A2(n411), .A4(n412), .S0(n293), 
        .S1(n297), .Y(n410) );
  OA21X1_HVT U170 ( .A1(n256), .A2(n301), .A3(n550), .Y(n408) );
  MUX41X1_HVT U172 ( .A1(n407), .A3(n413), .A2(n410), .A4(n415), .S0(in[0]), 
        .S1(in[5]), .Y(n406) );
  NAND2X0_HVT U174 ( .A1(n236), .A2(n574), .Y(n567) );
  MUX41X1_HVT U176 ( .A1(n274), .A3(n405), .A2(n350), .A4(n567), .S0(n299), 
        .S1(n293), .Y(n404) );
  NAND2X0_HVT U177 ( .A1(n237), .A2(n274), .Y(n403) );
  MUX41X1_HVT U178 ( .A1(n563), .A3(n403), .A2(n354), .A4(n543), .S0(n261), 
        .S1(n241), .Y(n402) );
  MUX41X1_HVT U179 ( .A1(n553), .A3(n355), .A2(n307), .A4(n354), .S0(n293), 
        .S1(n241), .Y(n401) );
  MUX41X1_HVT U180 ( .A1(n310), .A3(n572), .A2(n568), .A4(n250), .S0(n267), 
        .S1(n293), .Y(n400) );
  MUX41X1_HVT U181 ( .A1(n400), .A3(n402), .A2(n401), .A4(n404), .S0(n276), 
        .S1(n265), .Y(n399) );
  MUX41X1_HVT U182 ( .A1(n334), .A3(n280), .A2(n336), .A4(n323), .S0(n297), 
        .S1(n293), .Y(n398) );
  OA21X1_HVT U184 ( .A1(n547), .A2(n301), .A3(n321), .Y(n396) );
  MUX41X1_HVT U186 ( .A1(n253), .A3(n542), .A2(n508), .A4(n535), .S0(n293), 
        .S1(n241), .Y(n394) );
  MUX41X1_HVT U189 ( .A1(n392), .A3(n567), .A2(n393), .A4(n341), .S0(n267), 
        .S1(n261), .Y(n391) );
  MUX41X1_HVT U190 ( .A1(n391), .A3(n394), .A2(n395), .A4(n398), .S0(n265), 
        .S1(in[0]), .Y(n390) );
  MUX41X1_HVT U193 ( .A1(n539), .A3(n546), .A2(n533), .A4(n389), .S0(n293), 
        .S1(n298), .Y(n388) );
  MUX41X1_HVT U194 ( .A1(n540), .A3(n554), .A2(n352), .A4(n279), .S0(n267), 
        .S1(n262), .Y(n387) );
  MUX41X1_HVT U195 ( .A1(n574), .A3(n346), .A2(n284), .A4(n544), .S0(n259), 
        .S1(n241), .Y(n386) );
  AO21X1_HVT U197 ( .A1(n255), .A2(n268), .A3(n343), .Y(n384) );
  MUX41X1_HVT U199 ( .A1(n383), .A3(n387), .A2(n386), .A4(n388), .S0(n276), 
        .S1(n265), .Y(n382) );
  MUX41X1_HVT U203 ( .A1(n545), .A3(n335), .A2(n569), .A4(n549), .S0(n263), 
        .S1(n299), .Y(n378) );
  MUX41X1_HVT U204 ( .A1(n526), .A3(n568), .A2(n330), .A4(n558), .S0(n293), 
        .S1(n297), .Y(n377) );
  NAND2X0_HVT U208 ( .A1(n289), .A2(n280), .Y(n468) );
  NAND2X0_HVT U212 ( .A1(n289), .A2(n278), .Y(n525) );
  NAND2X0_HVT U214 ( .A1(n574), .A2(n292), .Y(n374) );
  NAND2X0_HVT U215 ( .A1(n468), .A2(n279), .Y(n373) );
  NAND2X0_HVT U218 ( .A1(n357), .A2(n286), .Y(n427) );
  NAND2X0_HVT U220 ( .A1(n268), .A2(n374), .Y(n500) );
  XOR2X2_HVT U1 ( .A1(n301), .A2(n554), .Y(n537) );
  XOR2X1_HVT U2 ( .A1(n294), .A2(n301), .Y(n245) );
  AO21X2_HVT U6 ( .A1(n291), .A2(n357), .A3(n301), .Y(n478) );
  INVX4_HVT U7 ( .A(in[7]), .Y(n301) );
  IBUFFX2_HVT U8 ( .A(n291), .Y(n289) );
  XNOR2X2_HVT U9 ( .A1(n361), .A2(in[3]), .Y(n23) );
  INVX8_HVT U10 ( .A(n23), .Y(n574) );
  AO21X2_HVT U11 ( .A1(n262), .A2(n279), .A3(n574), .Y(n460) );
  MUX21X2_HVT U12 ( .A1(n558), .A2(n334), .S0(n268), .Y(n440) );
  MUX21X2_HVT U14 ( .A1(n397), .A2(n396), .S0(n48), .Y(n395) );
  IBUFFX16_HVT U16 ( .A(n262), .Y(n48) );
  NBUFFX2_HVT U17 ( .A(n23), .Y(n273) );
  INVX1_HVT U18 ( .A(n558), .Y(n321) );
  MUX21X2_HVT U19 ( .A1(n577), .A2(n440), .S0(n50), .Y(n439) );
  IBUFFX16_HVT U20 ( .A(n259), .Y(n50) );
  INVX1_HVT U22 ( .A(n291), .Y(n290) );
  MUX21X2_HVT U23 ( .A1(n277), .A2(n273), .S0(n210), .Y(n558) );
  IBUFFX16_HVT U25 ( .A(n236), .Y(n210) );
  NAND2X0_HVT U26 ( .A1(n380), .A2(n211), .Y(n212) );
  NAND2X0_HVT U27 ( .A1(n381), .A2(n262), .Y(n213) );
  NAND2X0_HVT U28 ( .A1(n212), .A2(n213), .Y(n379) );
  IBUFFX2_HVT U29 ( .A(n262), .Y(n211) );
  OA21X2_HVT U30 ( .A1(n573), .A2(n301), .A3(n333), .Y(n380) );
  MUX21X1_HVT U31 ( .A1(n564), .A2(n250), .S0(n267), .Y(n381) );
  IBUFFX2_HVT U32 ( .A(n300), .Y(n296) );
  IBUFFX2_HVT U34 ( .A(n300), .Y(n297) );
  INVX1_HVT U36 ( .A(n300), .Y(n299) );
  MUX21X1_HVT U37 ( .A1(n539), .A2(n535), .S0(n218), .Y(n216) );
  MUX21X1_HVT U38 ( .A1(n492), .A2(n344), .S0(n218), .Y(n217) );
  MUX21X1_HVT U39 ( .A1(n216), .A2(n217), .S0(n299), .Y(n491) );
  IBUFFX2_HVT U40 ( .A(n260), .Y(n218) );
  MUX21X2_HVT U41 ( .A1(n430), .A2(n438), .S0(in[6]), .Y(out[4]) );
  MUX21X2_HVT U43 ( .A1(n390), .A2(n399), .S0(in[6]), .Y(out[6]) );
  NBUFFX4_HVT U44 ( .A(n298), .Y(n241) );
  INVX2_HVT U45 ( .A(in[7]), .Y(n300) );
  INVX2_HVT U46 ( .A(n300), .Y(n298) );
  MUX21X2_HVT U47 ( .A1(n459), .A2(n462), .S0(n266), .Y(n458) );
  MUX41X1_HVT U48 ( .A1(n342), .A3(n360), .A2(n347), .A4(n322), .S0(n299), 
        .S1(n259), .Y(n506) );
  MUX21X2_HVT U49 ( .A1(n418), .A2(n406), .S0(n219), .Y(out[5]) );
  IBUFFX16_HVT U50 ( .A(in[6]), .Y(n219) );
  MUX41X1_HVT U52 ( .A1(n484), .A3(n491), .A2(n483), .A4(n486), .S0(n276), 
        .S1(n231), .Y(n482) );
  IBUFFX16_HVT U54 ( .A(n295), .Y(n231) );
  NBUFFX2_HVT U55 ( .A(in[5]), .Y(n266) );
  INVX0_HVT U60 ( .A(n232), .Y(n442) );
  INVX0_HVT U64 ( .A(n554), .Y(n234) );
  INVX1_HVT U65 ( .A(n291), .Y(n287) );
  INVX0_HVT U67 ( .A(n575), .Y(n233) );
  INVX0_HVT U70 ( .A(n261), .Y(n235) );
  INVX1_HVT U71 ( .A(in[4]), .Y(n361) );
  MUX41X1_HVT U72 ( .A1(n234), .A3(n233), .A2(n278), .A4(n365), .S0(n235), 
        .S1(n301), .Y(n232) );
  IBUFFX2_HVT U75 ( .A(n291), .Y(n236) );
  IBUFFX2_HVT U76 ( .A(n291), .Y(n237) );
  MUX21X1_HVT U79 ( .A1(n275), .A2(n270), .S0(n292), .Y(n389) );
  NAND2X0_HVT U81 ( .A1(n375), .A2(n238), .Y(n239) );
  NAND2X0_HVT U88 ( .A1(n382), .A2(in[6]), .Y(n240) );
  NAND2X0_HVT U89 ( .A1(n239), .A2(n240), .Y(out[7]) );
  IBUFFX2_HVT U90 ( .A(in[6]), .Y(n238) );
  MUX41X1_HVT U91 ( .A1(n578), .A3(n242), .A2(n328), .A4(n355), .S0(n294), 
        .S1(n299), .Y(n376) );
  IBUFFX2_HVT U92 ( .A(n291), .Y(n288) );
  MUX21X2_HVT U94 ( .A1(n254), .A2(n481), .S0(n245), .Y(n480) );
  INVX2_HVT U95 ( .A(in[1]), .Y(n291) );
  MUX41X1_HVT U98 ( .A1(n535), .A3(n342), .A2(n508), .A4(n353), .S0(n235), 
        .S1(n301), .Y(n431) );
  MUX21X2_HVT U99 ( .A1(n493), .A2(n503), .S0(in[6]), .Y(out[1]) );
  INVX1_HVT U100 ( .A(in[2]), .Y(n294) );
  NBUFFX2_HVT U102 ( .A(n23), .Y(n272) );
  MUX21X1_HVT U104 ( .A1(n272), .A2(n270), .S0(n290), .Y(n564) );
  INVX1_HVT U106 ( .A(n276), .Y(n243) );
  INVX1_HVT U107 ( .A(n295), .Y(n244) );
  INVX1_HVT U108 ( .A(n275), .Y(n242) );
  MUX41X1_HVT U111 ( .A1(n379), .A3(n377), .A2(n378), .A4(n376), .S0(n243), 
        .S1(n244), .Y(n375) );
  MUX41X1_HVT U112 ( .A1(n278), .A3(n340), .A2(n271), .A4(n321), .S0(n235), 
        .S1(n301), .Y(n435) );
  MUX41X1_HVT U113 ( .A1(n436), .A3(n432), .A2(n435), .A4(n431), .S0(n243), 
        .S1(n244), .Y(n430) );
  MUX41X1_HVT U114 ( .A1(n329), .A3(n437), .A2(n333), .A4(n556), .S0(n235), 
        .S1(n301), .Y(n436) );
  MUX41X1_HVT U117 ( .A1(n473), .A3(n476), .A2(n475), .A4(n480), .S0(in[0]), 
        .S1(n265), .Y(n472) );
  MUX41X1_HVT U118 ( .A1(n465), .A3(n467), .A2(n471), .A4(n470), .S0(n296), 
        .S1(n266), .Y(n464) );
  NAND2X0_HVT U119 ( .A1(n579), .A2(n246), .Y(n247) );
  NAND2X0_HVT U120 ( .A1(n466), .A2(n249), .Y(n248) );
  NAND2X0_HVT U121 ( .A1(n247), .A2(n248), .Y(n465) );
  INVX0_HVT U122 ( .A(n249), .Y(n246) );
  XNOR2X1_HVT U124 ( .A1(n289), .A2(n263), .Y(n249) );
  MUX21X2_HVT U126 ( .A1(n472), .A2(n482), .S0(in[6]), .Y(out[2]) );
  MUX21X2_HVT U127 ( .A1(n337), .A2(n354), .S0(n268), .Y(n385) );
  INVX0_HVT U129 ( .A(n291), .Y(n286) );
  INVX0_HVT U130 ( .A(in[3]), .Y(n358) );
  INVX0_HVT U133 ( .A(n294), .Y(n293) );
  INVX1_HVT U134 ( .A(n576), .Y(n356) );
  MUX21X1_HVT U135 ( .A1(n252), .A2(n316), .S0(n260), .Y(n447) );
  NBUFFX2_HVT U137 ( .A(n23), .Y(n271) );
  AND2X1_HVT U138 ( .A1(n273), .A2(n525), .Y(n250) );
  INVX1_HVT U141 ( .A(n282), .Y(n360) );
  MUX21X1_HVT U142 ( .A1(n356), .A2(n359), .S0(n266), .Y(n529) );
  NBUFFX2_HVT U143 ( .A(n576), .Y(n280) );
  MUX21X1_HVT U145 ( .A1(n550), .A2(n469), .S0(n260), .Y(n467) );
  NBUFFX2_HVT U147 ( .A(n576), .Y(n281) );
  MUX21X1_HVT U148 ( .A1(n312), .A2(n357), .S0(n266), .Y(n514) );
  AND2X1_HVT U149 ( .A1(n283), .A2(n508), .Y(n251) );
  MUX21X1_HVT U150 ( .A1(n273), .A2(n359), .S0(n286), .Y(n573) );
  MUX21X1_HVT U152 ( .A1(n451), .A2(n452), .S0(n266), .Y(n450) );
  MUX21X1_HVT U155 ( .A1(n456), .A2(n455), .S0(n269), .Y(n452) );
  MUX21X1_HVT U156 ( .A1(n283), .A2(n272), .S0(n288), .Y(n540) );
  MUX21X1_HVT U157 ( .A1(n271), .A2(n275), .S0(n290), .Y(n477) );
  MUX21X1_HVT U161 ( .A1(n272), .A2(n356), .S0(n286), .Y(n485) );
  MUX21X1_HVT U164 ( .A1(n281), .A2(n574), .S0(n237), .Y(n544) );
  MUX21X1_HVT U169 ( .A1(n356), .A2(n360), .S0(n286), .Y(n405) );
  MUX21X1_HVT U171 ( .A1(n359), .A2(n272), .S0(n290), .Y(n417) );
  MUX21X1_HVT U173 ( .A1(n574), .A2(n357), .S0(n236), .Y(n365) );
  MUX21X1_HVT U175 ( .A1(n574), .A2(n360), .S0(n290), .Y(n556) );
  MUX21X1_HVT U183 ( .A1(n280), .A2(n279), .S0(n236), .Y(n492) );
  MUX21X1_HVT U185 ( .A1(n574), .A2(n275), .S0(n288), .Y(n505) );
  XOR2X1_HVT U187 ( .A1(n574), .A2(n286), .Y(n535) );
  MUX21X1_HVT U188 ( .A1(n270), .A2(n574), .S0(n289), .Y(n368) );
  MUX21X1_HVT U191 ( .A1(n360), .A2(n359), .S0(n290), .Y(n554) );
  MUX21X1_HVT U192 ( .A1(n359), .A2(n356), .S0(n237), .Y(n543) );
  MUX21X1_HVT U196 ( .A1(n270), .A2(n360), .S0(n287), .Y(n541) );
  MUX21X1_HVT U198 ( .A1(n275), .A2(n356), .S0(n237), .Y(n552) );
  MUX21X1_HVT U200 ( .A1(n327), .A2(n444), .S0(n263), .Y(n443) );
  MUX21X1_HVT U201 ( .A1(n351), .A2(n279), .S0(n268), .Y(n444) );
  MUX21X1_HVT U202 ( .A1(n460), .A2(n461), .S0(n268), .Y(n459) );
  MUX21X1_HVT U205 ( .A1(n305), .A2(n330), .S0(n260), .Y(n461) );
  NAND2X0_HVT U206 ( .A1(n274), .A2(n358), .Y(n576) );
  MUX21X1_HVT U207 ( .A1(n356), .A2(n274), .S0(n288), .Y(n366) );
  NBUFFX2_HVT U209 ( .A(n579), .Y(n282) );
  MUX21X1_HVT U210 ( .A1(n283), .A2(n278), .S0(n288), .Y(n566) );
  MUX21X1_HVT U211 ( .A1(n359), .A2(n270), .S0(n287), .Y(n547) );
  MUX21X1_HVT U213 ( .A1(n357), .A2(n356), .S0(n287), .Y(n562) );
  MUX21X1_HVT U216 ( .A1(n328), .A2(n566), .S0(n263), .Y(n481) );
  MUX21X1_HVT U217 ( .A1(n304), .A2(n457), .S0(n261), .Y(n456) );
  MUX21X1_HVT U219 ( .A1(n274), .A2(n270), .S0(n288), .Y(n457) );
  NBUFFX2_HVT U221 ( .A(n579), .Y(n283) );
  MUX21X1_HVT U222 ( .A1(n270), .A2(n285), .S0(n237), .Y(n392) );
  MUX21X1_HVT U223 ( .A1(n284), .A2(n283), .S0(n290), .Y(n393) );
  INVX1_HVT U224 ( .A(n571), .Y(n357) );
  INVX1_HVT U225 ( .A(n284), .Y(n359) );
  MUX21X1_HVT U226 ( .A1(n281), .A2(n285), .S0(n236), .Y(n487) );
  MUX21X1_HVT U227 ( .A1(n270), .A2(n359), .S0(n287), .Y(n570) );
  XOR2X1_HVT U228 ( .A1(n287), .A2(n357), .Y(n536) );
  XOR2X1_HVT U229 ( .A1(n282), .A2(n289), .Y(n533) );
  MUX21X1_HVT U230 ( .A1(n282), .A2(n274), .S0(n237), .Y(n372) );
  XNOR2X1_HVT U231 ( .A1(n281), .A2(n236), .Y(n252) );
  AND2X1_HVT U232 ( .A1(n290), .A2(n360), .Y(n253) );
  MUX21X1_HVT U233 ( .A1(n284), .A2(n278), .S0(n286), .Y(n550) );
  MUX21X1_HVT U234 ( .A1(n280), .A2(n270), .S0(n236), .Y(n569) );
  MUX21X1_HVT U235 ( .A1(n282), .A2(n280), .S0(n288), .Y(n364) );
  AND2X1_HVT U236 ( .A1(n285), .A2(n468), .Y(n254) );
  XNOR2X1_HVT U237 ( .A1(n284), .A2(n287), .Y(n255) );
  MUX21X1_HVT U238 ( .A1(n278), .A2(n270), .S0(n237), .Y(n370) );
  MUX21X1_HVT U239 ( .A1(n279), .A2(n274), .S0(n286), .Y(n510) );
  MUX21X1_HVT U240 ( .A1(n279), .A2(n285), .S0(n263), .Y(n454) );
  XOR2X1_HVT U241 ( .A1(n274), .A2(n289), .Y(n555) );
  NBUFFX2_HVT U242 ( .A(n298), .Y(n269) );
  NBUFFX2_HVT U243 ( .A(n298), .Y(n267) );
  NBUFFX2_HVT U244 ( .A(n298), .Y(n268) );
  NBUFFX2_HVT U245 ( .A(n358), .Y(n270) );
  NBUFFX2_HVT U246 ( .A(in[2]), .Y(n260) );
  NBUFFX2_HVT U247 ( .A(in[2]), .Y(n261) );
  NBUFFX2_HVT U248 ( .A(in[5]), .Y(n265) );
  NBUFFX2_HVT U249 ( .A(in[2]), .Y(n263) );
  NBUFFX2_HVT U250 ( .A(in[2]), .Y(n262) );
  NBUFFX2_HVT U251 ( .A(n295), .Y(n264) );
  NBUFFX2_HVT U252 ( .A(in[2]), .Y(n259) );
  MUX21X1_HVT U253 ( .A1(n479), .A2(n327), .S0(n263), .Y(n476) );
  MUX21X1_HVT U254 ( .A1(n495), .A2(n277), .S0(n268), .Y(n397) );
  MUX21X1_HVT U255 ( .A1(n518), .A2(n520), .S0(n262), .Y(n517) );
  XOR2X1_HVT U256 ( .A1(n236), .A2(n277), .Y(n534) );
  MUX21X1_HVT U257 ( .A1(n278), .A2(n273), .S0(n236), .Y(n474) );
  MUX21X1_HVT U258 ( .A1(n502), .A2(n501), .S0(n260), .Y(n499) );
  MUX21X1_HVT U259 ( .A1(n560), .A2(n279), .S0(n269), .Y(n502) );
  MUX21X1_HVT U260 ( .A1(n409), .A2(n408), .S0(n263), .Y(n407) );
  MUX21X1_HVT U261 ( .A1(n279), .A2(n346), .S0(n269), .Y(n409) );
  MUX21X1_HVT U262 ( .A1(n428), .A2(n429), .S0(n262), .Y(n426) );
  MUX21X1_HVT U263 ( .A1(n348), .A2(n357), .S0(n268), .Y(n429) );
  MUX21X1_HVT U264 ( .A1(n357), .A2(n360), .S0(n289), .Y(n414) );
  AND2X1_HVT U265 ( .A1(n273), .A2(n292), .Y(n256) );
  MUX21X1_HVT U266 ( .A1(n277), .A2(n356), .S0(n237), .Y(n542) );
  MUX21X1_HVT U267 ( .A1(n537), .A2(n512), .S0(n262), .Y(n511) );
  MUX21X1_HVT U268 ( .A1(n359), .A2(n346), .S0(n269), .Y(n512) );
  MUX21X1_HVT U269 ( .A1(n434), .A2(n433), .S0(n263), .Y(n432) );
  MUX21X1_HVT U270 ( .A1(n552), .A2(n308), .S0(n269), .Y(n434) );
  NAND2X0_HVT U271 ( .A1(in[3]), .A2(n275), .Y(n579) );
  NBUFFX2_HVT U272 ( .A(n361), .Y(n275) );
  MUX21X1_HVT U273 ( .A1(n360), .A2(n277), .S0(n288), .Y(n561) );
  MUX21X1_HVT U274 ( .A1(n331), .A2(n578), .S0(n261), .Y(n471) );
  MUX21X1_HVT U275 ( .A1(n422), .A2(n423), .S0(n259), .Y(n421) );
  MUX21X1_HVT U276 ( .A1(n424), .A2(n283), .S0(n257), .Y(n423) );
  MUX21X1_HVT U277 ( .A1(n543), .A2(n349), .S0(n267), .Y(n422) );
  MUX21X1_HVT U278 ( .A1(n563), .A2(n329), .S0(n261), .Y(n446) );
  MUX21X1_HVT U279 ( .A1(n530), .A2(n531), .S0(n267), .Y(n528) );
  MUX21X1_HVT U280 ( .A1(n277), .A2(n546), .S0(n266), .Y(n531) );
  XOR2X1_HVT U281 ( .A1(n288), .A2(n265), .Y(n538) );
  MUX21X1_HVT U282 ( .A1(n578), .A2(n291), .S0(n262), .Y(n453) );
  NBUFFX2_HVT U283 ( .A(n580), .Y(n284) );
  MUX21X1_HVT U284 ( .A1(n277), .A2(n357), .S0(n236), .Y(n369) );
  MUX21X1_HVT U285 ( .A1(n551), .A2(n373), .S0(n267), .Y(n367) );
  MUX21X1_HVT U286 ( .A1(n281), .A2(n277), .S0(n287), .Y(n572) );
  MUX21X1_HVT U287 ( .A1(n314), .A2(n292), .S0(n266), .Y(n516) );
  NBUFFX2_HVT U288 ( .A(n571), .Y(n278) );
  MUX21X1_HVT U289 ( .A1(n324), .A2(n551), .S0(n261), .Y(n449) );
  MUX21X1_HVT U290 ( .A1(n283), .A2(n490), .S0(n257), .Y(n489) );
  MUX21X1_HVT U291 ( .A1(n277), .A2(n274), .S0(n269), .Y(n490) );
  NBUFFX2_HVT U292 ( .A(n580), .Y(n285) );
  NBUFFX2_HVT U293 ( .A(n361), .Y(n274) );
  NBUFFX2_HVT U294 ( .A(n571), .Y(n279) );
  XNOR2X1_HVT U295 ( .A1(n300), .A2(n289), .Y(n257) );
  AND2X1_HVT U296 ( .A1(n270), .A2(n292), .Y(n258) );
  NBUFFX2_HVT U297 ( .A(in[5]), .Y(n295) );
  MUX21X1_HVT U298 ( .A1(n385), .A2(n384), .S0(n262), .Y(n383) );
  MUX21X1_HVT U299 ( .A1(n488), .A2(n489), .S0(n263), .Y(n486) );
  MUX21X1_HVT U300 ( .A1(n528), .A2(n532), .S0(n263), .Y(n527) );
  MUX21X1_HVT U301 ( .A1(n522), .A2(n524), .S0(n262), .Y(n521) );
  MUX21X1_HVT U302 ( .A1(n356), .A2(n242), .S0(n288), .Y(n549) );
  MUX21X1_HVT U303 ( .A1(n242), .A2(n574), .S0(n287), .Y(n371) );
  MUX21X1_HVT U304 ( .A1(n242), .A2(n359), .S0(n290), .Y(n545) );
  MUX21X1_HVT U305 ( .A1(n242), .A2(n357), .S0(n289), .Y(n563) );
  NAND2X0_HVT U306 ( .A1(in[4]), .A2(n358), .Y(n571) );
  NAND2X0_HVT U307 ( .A1(in[3]), .A2(in[4]), .Y(n580) );
  MUX21X1_HVT U308 ( .A1(n242), .A2(n283), .S0(n237), .Y(n560) );
  MUX21X1_HVT U309 ( .A1(n285), .A2(n242), .S0(n289), .Y(n553) );
  MUX21X1_HVT U310 ( .A1(n277), .A2(n242), .S0(n260), .Y(n466) );
  MUX21X1_HVT U311 ( .A1(n242), .A2(n278), .S0(n290), .Y(n363) );
  MUX21X1_HVT U312 ( .A1(n242), .A2(n285), .S0(n286), .Y(n362) );
  MUX21X1_HVT U313 ( .A1(n270), .A2(n242), .S0(n237), .Y(n551) );
  INVX0_HVT U314 ( .A(in[1]), .Y(n292) );
  NBUFFX2_HVT U315 ( .A(in[3]), .Y(n277) );
  NBUFFX2_HVT U316 ( .A(in[0]), .Y(n276) );
  INVX0_HVT U317 ( .A(n559), .Y(n302) );
  INVX0_HVT U318 ( .A(n557), .Y(n303) );
  INVX0_HVT U319 ( .A(n548), .Y(n304) );
  INVX0_HVT U320 ( .A(n546), .Y(n305) );
  INVX0_HVT U321 ( .A(n411), .Y(n306) );
  INVX0_HVT U322 ( .A(n374), .Y(n307) );
  INVX0_HVT U323 ( .A(n578), .Y(n308) );
  INVX0_HVT U324 ( .A(n565), .Y(n309) );
  INVX0_HVT U325 ( .A(n577), .Y(n310) );
  INVX0_HVT U326 ( .A(n573), .Y(n311) );
  INVX0_HVT U327 ( .A(n572), .Y(n312) );
  INVX0_HVT U328 ( .A(n570), .Y(n313) );
  INVX0_HVT U329 ( .A(n569), .Y(n314) );
  INVX0_HVT U330 ( .A(n566), .Y(n315) );
  INVX0_HVT U331 ( .A(n564), .Y(n316) );
  INVX0_HVT U332 ( .A(n563), .Y(n317) );
  INVX0_HVT U333 ( .A(n562), .Y(n318) );
  INVX0_HVT U334 ( .A(n561), .Y(n319) );
  INVX0_HVT U335 ( .A(n560), .Y(n320) );
  INVX0_HVT U336 ( .A(n556), .Y(n322) );
  INVX0_HVT U337 ( .A(n555), .Y(n323) );
  INVX0_HVT U338 ( .A(n553), .Y(n324) );
  INVX0_HVT U339 ( .A(n552), .Y(n325) );
  INVX0_HVT U340 ( .A(n551), .Y(n326) );
  INVX0_HVT U341 ( .A(n367), .Y(n327) );
  INVX0_HVT U342 ( .A(n550), .Y(n328) );
  INVX0_HVT U343 ( .A(n549), .Y(n329) );
  INVX0_HVT U344 ( .A(n547), .Y(n330) );
  INVX0_HVT U345 ( .A(n545), .Y(n331) );
  INVX0_HVT U346 ( .A(n544), .Y(n332) );
  INVX0_HVT U347 ( .A(n543), .Y(n333) );
  INVX0_HVT U348 ( .A(n542), .Y(n334) );
  INVX0_HVT U349 ( .A(n541), .Y(n335) );
  INVX0_HVT U350 ( .A(n540), .Y(n336) );
  INVX0_HVT U351 ( .A(n539), .Y(n337) );
  INVX0_HVT U352 ( .A(n508), .Y(n338) );
  INVX0_HVT U353 ( .A(n568), .Y(n339) );
  INVX0_HVT U354 ( .A(n468), .Y(n340) );
  INVX0_HVT U355 ( .A(n373), .Y(n341) );
  INVX0_HVT U356 ( .A(n525), .Y(n342) );
  INVX0_HVT U357 ( .A(n427), .Y(n343) );
  INVX0_HVT U358 ( .A(n372), .Y(n344) );
  INVX0_HVT U359 ( .A(n371), .Y(n345) );
  INVX0_HVT U360 ( .A(n370), .Y(n346) );
  INVX0_HVT U361 ( .A(n369), .Y(n347) );
  INVX0_HVT U362 ( .A(n368), .Y(n348) );
  INVX0_HVT U363 ( .A(n487), .Y(n349) );
  INVX0_HVT U364 ( .A(n477), .Y(n350) );
  INVX0_HVT U365 ( .A(n366), .Y(n351) );
  INVX0_HVT U366 ( .A(n365), .Y(n352) );
  INVX0_HVT U367 ( .A(n364), .Y(n353) );
  INVX0_HVT U368 ( .A(n363), .Y(n354) );
  INVX0_HVT U369 ( .A(n362), .Y(n355) );
endmodule

