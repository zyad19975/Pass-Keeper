
module sbox_4 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n50, n121, n168, n210, n211, n212, n213, n216, n217, n218,
         n219, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597;

  NAND2X0_HVT U4 ( .A1(n302), .A2(n595), .Y(n594) );
  NAND2X0_HVT U5 ( .A1(n311), .A2(n291), .Y(n592) );
  NAND2X0_HVT U13 ( .A1(n584), .A2(n306), .Y(n585) );
  NAND2X0_HVT U15 ( .A1(n595), .A2(n293), .Y(n582) );
  NAND2X0_HVT U21 ( .A1(n302), .A2(n313), .Y(n576) );
  NAND2X0_HVT U24 ( .A1(n297), .A2(n313), .Y(n574) );
  NAND2X0_HVT U33 ( .A1(n375), .A2(n313), .Y(n565) );
  NAND2X0_HVT U35 ( .A1(n295), .A2(n313), .Y(n563) );
  NAND2X0_HVT U42 ( .A1(n50), .A2(n297), .Y(n556) );
  MUX41X1_HVT U51 ( .A1(n363), .A3(n323), .A2(n340), .A4(n341), .S0(n255), 
        .S1(n317), .Y(n549) );
  NAND2X0_HVT U53 ( .A1(n546), .A2(n555), .Y(n547) );
  NAND2X0_HVT U56 ( .A1(n302), .A2(n542), .Y(n543) );
  MUX41X1_HVT U57 ( .A1(n364), .A3(n578), .A2(n543), .A4(n587), .S0(n255), 
        .S1(n317), .Y(n541) );
  NAND2X0_HVT U58 ( .A1(n306), .A2(n595), .Y(n540) );
  MUX41X1_HVT U59 ( .A1(n280), .A3(n540), .A2(n278), .A4(n339), .S0(n254), 
        .S1(n317), .Y(n539) );
  MUX41X1_HVT U61 ( .A1(n276), .A3(n338), .A2(n337), .A4(n293), .S0(n255), 
        .S1(n317), .Y(n537) );
  NAND2X0_HVT U62 ( .A1(n313), .A2(n305), .Y(n536) );
  AO21X1_HVT U66 ( .A1(n334), .A2(n318), .A3(n358), .Y(n532) );
  MUX41X1_HVT U68 ( .A1(n332), .A3(n532), .A2(n531), .A4(n533), .S0(n281), 
        .S1(n254), .Y(n530) );
  MUX41X1_HVT U69 ( .A1(n530), .A3(n538), .A2(n534), .A4(n544), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n299), .A2(n525), .Y(n526) );
  MUX41X1_HVT U74 ( .A1(n527), .A3(n572), .A2(n526), .A4(n574), .S0(n283), 
        .S1(n320), .Y(n524) );
  MUX41X1_HVT U75 ( .A1(n361), .A3(n366), .A2(n379), .A4(n343), .S0(n281), 
        .S1(n255), .Y(n523) );
  MUX41X1_HVT U77 ( .A1(n589), .A3(n368), .A2(n522), .A4(n367), .S0(n288), 
        .S1(n315), .Y(n521) );
  MUX41X1_HVT U78 ( .A1(n521), .A3(n524), .A2(n523), .A4(n528), .S0(in[0]), 
        .S1(n317), .Y(n520) );
  AND3X1_HVT U80 ( .A1(n304), .A2(n542), .A3(n517), .Y(n518) );
  MUX41X1_HVT U82 ( .A1(n553), .A3(n341), .A2(n324), .A4(n583), .S0(n281), 
        .S1(n320), .Y(n515) );
  AND2X1_HVT U83 ( .A1(n310), .A2(n262), .Y(n514) );
  MUX41X1_HVT U84 ( .A1(n342), .A3(n591), .A2(n581), .A4(n514), .S0(n281), 
        .S1(n320), .Y(n513) );
  NAND2X0_HVT U85 ( .A1(n313), .A2(n378), .Y(n512) );
  MUX41X1_HVT U86 ( .A1(n366), .A3(n512), .A2(n277), .A4(n273), .S0(n281), 
        .S1(n319), .Y(n511) );
  MUX41X1_HVT U87 ( .A1(n511), .A3(n515), .A2(n513), .A4(n516), .S0(in[0]), 
        .S1(n286), .Y(n510) );
  MUX41X1_HVT U90 ( .A1(n552), .A3(n556), .A2(n363), .A4(n509), .S0(n282), 
        .S1(n254), .Y(n508) );
  AO21X1_HVT U93 ( .A1(n290), .A2(n504), .A3(n362), .Y(n505) );
  MUX41X1_HVT U96 ( .A1(n324), .A3(n275), .A2(n365), .A4(n502), .S0(n281), 
        .S1(n319), .Y(n501) );
  MUX41X1_HVT U97 ( .A1(n361), .A3(n275), .A2(n310), .A4(n582), .S0(n281), 
        .S1(n254), .Y(n500) );
  MUX41X1_HVT U98 ( .A1(n500), .A3(n503), .A2(n501), .A4(n508), .S0(n296), 
        .S1(n286), .Y(n499) );
  NAND2X0_HVT U101 ( .A1(n495), .A2(n494), .Y(n496) );
  MUX41X1_HVT U103 ( .A1(n595), .A3(n333), .A2(n346), .A4(n563), .S0(n281), 
        .S1(n320), .Y(n492) );
  MUX41X1_HVT U105 ( .A1(n345), .A3(n551), .A2(n491), .A4(n360), .S0(n281), 
        .S1(n255), .Y(n490) );
  NAND2X0_HVT U110 ( .A1(n304), .A2(n485), .Y(n486) );
  AO21X1_HVT U118 ( .A1(n285), .A2(n298), .A3(n591), .Y(n478) );
  NAND2X0_HVT U123 ( .A1(n472), .A2(n471), .Y(n473) );
  MUX41X1_HVT U125 ( .A1(n576), .A3(n280), .A2(n332), .A4(n370), .S0(n282), 
        .S1(n255), .Y(n469) );
  AND3X1_HVT U128 ( .A1(n285), .A2(n313), .A3(n262), .Y(n466) );
  MUX41X1_HVT U131 ( .A1(n464), .A3(n466), .A2(n465), .A4(n467), .S0(n318), 
        .S1(n320), .Y(n463) );
  MUX41X1_HVT U132 ( .A1(n463), .A3(n476), .A2(n468), .A4(n481), .S0(in[6]), 
        .S1(n296), .Y(out[3]) );
  MUX41X1_HVT U135 ( .A1(n371), .A3(n376), .A2(n592), .A4(n571), .S0(n283), 
        .S1(n254), .Y(n460) );
  MUX41X1_HVT U136 ( .A1(n273), .A3(n565), .A2(n372), .A4(n562), .S0(n282), 
        .S1(n254), .Y(n459) );
  MUX41X1_HVT U139 ( .A1(n457), .A3(n460), .A2(n459), .A4(n461), .S0(n296), 
        .S1(n286), .Y(n456) );
  AND2X1_HVT U140 ( .A1(n298), .A2(n312), .Y(n455) );
  MUX41X1_HVT U142 ( .A1(n342), .A3(n292), .A2(n359), .A4(n298), .S0(n282), 
        .S1(n320), .Y(n453) );
  OA21X1_HVT U144 ( .A1(n327), .A2(n321), .A3(n567), .Y(n451) );
  NAND2X0_HVT U146 ( .A1(n307), .A2(n306), .Y(n525) );
  MUX41X1_HVT U147 ( .A1(n372), .A3(n525), .A2(n361), .A4(n552), .S0(n283), 
        .S1(n320), .Y(n449) );
  MUX41X1_HVT U148 ( .A1(n449), .A3(n453), .A2(n450), .A4(n454), .S0(in[0]), 
        .S1(n286), .Y(n448) );
  OA21X1_HVT U151 ( .A1(n558), .A2(n321), .A3(n445), .Y(n446) );
  AND2X1_HVT U154 ( .A1(n290), .A2(n297), .Y(n442) );
  NAND2X0_HVT U158 ( .A1(n249), .A2(n378), .Y(n438) );
  MUX41X1_HVT U159 ( .A1(n585), .A3(n292), .A2(n438), .A4(n331), .S0(n314), 
        .S1(n255), .Y(n437) );
  MUX41X1_HVT U160 ( .A1(n437), .A3(n443), .A2(n439), .A4(n444), .S0(n296), 
        .S1(n287), .Y(n436) );
  MUX41X1_HVT U165 ( .A1(n576), .A3(n347), .A2(n552), .A4(n433), .S0(n254), 
        .S1(n315), .Y(n432) );
  NAND2X0_HVT U166 ( .A1(n306), .A2(n542), .Y(n431) );
  NAND2X0_HVT U167 ( .A1(n379), .A2(n313), .Y(n430) );
  MUX41X1_HVT U168 ( .A1(n364), .A3(n298), .A2(n430), .A4(n431), .S0(n315), 
        .S1(n319), .Y(n429) );
  OA21X1_HVT U170 ( .A1(n278), .A2(n321), .A3(n567), .Y(n427) );
  MUX41X1_HVT U172 ( .A1(n426), .A3(n432), .A2(n429), .A4(n434), .S0(in[0]), 
        .S1(n286), .Y(n425) );
  MUX21X2_HVT U173 ( .A1(n425), .A2(n436), .S0(in[6]), .Y(out[5]) );
  NAND2X0_HVT U174 ( .A1(n250), .A2(n591), .Y(n584) );
  MUX41X1_HVT U176 ( .A1(n295), .A3(n424), .A2(n369), .A4(n584), .S0(n255), 
        .S1(n314), .Y(n423) );
  NAND2X0_HVT U177 ( .A1(n307), .A2(n294), .Y(n422) );
  MUX41X1_HVT U178 ( .A1(n580), .A3(n422), .A2(n373), .A4(n560), .S0(n283), 
        .S1(n320), .Y(n421) );
  MUX41X1_HVT U179 ( .A1(n570), .A3(n374), .A2(n328), .A4(n373), .S0(n314), 
        .S1(n254), .Y(n420) );
  MUX41X1_HVT U180 ( .A1(n330), .A3(n589), .A2(n585), .A4(n272), .S0(n288), 
        .S1(n314), .Y(n419) );
  MUX41X1_HVT U181 ( .A1(n419), .A3(n421), .A2(n420), .A4(n423), .S0(n296), 
        .S1(n287), .Y(n418) );
  OA21X1_HVT U184 ( .A1(n564), .A2(n321), .A3(n342), .Y(n415) );
  MUX41X1_HVT U186 ( .A1(n275), .A3(n559), .A2(n525), .A4(n552), .S0(n315), 
        .S1(n319), .Y(n413) );
  MUX41X1_HVT U189 ( .A1(n411), .A3(n584), .A2(n412), .A4(n360), .S0(n288), 
        .S1(n314), .Y(n410) );
  MUX41X1_HVT U190 ( .A1(n410), .A3(n413), .A2(n414), .A4(n417), .S0(n287), 
        .S1(in[0]), .Y(n409) );
  MUX41X1_HVT U193 ( .A1(n556), .A3(n563), .A2(n550), .A4(n408), .S0(n315), 
        .S1(n319), .Y(n407) );
  MUX41X1_HVT U195 ( .A1(n591), .A3(n365), .A2(n597), .A4(n561), .S0(n315), 
        .S1(n254), .Y(n405) );
  AO21X1_HVT U197 ( .A1(n277), .A2(n289), .A3(n362), .Y(n403) );
  MUX41X1_HVT U199 ( .A1(n402), .A3(n406), .A2(n405), .A4(n407), .S0(in[0]), 
        .S1(n287), .Y(n401) );
  NAND2X0_HVT U208 ( .A1(n48), .A2(n302), .Y(n485) );
  NAND2X0_HVT U212 ( .A1(n248), .A2(n299), .Y(n542) );
  NAND2X0_HVT U214 ( .A1(n591), .A2(n313), .Y(n393) );
  NAND2X0_HVT U215 ( .A1(n485), .A2(n300), .Y(n392) );
  AO21X1_HVT U216 ( .A1(n312), .A2(n376), .A3(n321), .Y(n495) );
  NAND2X0_HVT U218 ( .A1(n376), .A2(n48), .Y(n445) );
  NAND2X0_HVT U220 ( .A1(n289), .A2(n393), .Y(n517) );
  MUX41X1_HVT U1 ( .A1(n264), .A3(n336), .A2(n536), .A4(n329), .S0(n320), .S1(
        n23), .Y(n535) );
  IBUFFX16_HVT U2 ( .A(n317), .Y(n23) );
  MUX21X1_HVT U3 ( .A1(n539), .A2(n541), .S0(n284), .Y(n538) );
  XOR2X2_HVT U6 ( .A1(n591), .A2(n309), .Y(n552) );
  IBUFFX2_HVT U7 ( .A(n312), .Y(n48) );
  IBUFFX2_HVT U8 ( .A(n312), .Y(n50) );
  INVX1_HVT U9 ( .A(in[1]), .Y(n312) );
  IBUFFX2_HVT U10 ( .A(n312), .Y(n307) );
  MUX41X1_HVT U11 ( .A1(n571), .A3(n557), .A2(n298), .A4(n371), .S0(n121), 
        .S1(n314), .Y(n406) );
  IBUFFX16_HVT U12 ( .A(n288), .Y(n121) );
  NAND2X0_HVT U14 ( .A1(n345), .A2(n168), .Y(n210) );
  NAND2X0_HVT U16 ( .A1(n213), .A2(n283), .Y(n211) );
  NAND2X0_HVT U17 ( .A1(n210), .A2(n211), .Y(n467) );
  IBUFFX2_HVT U18 ( .A(n283), .Y(n168) );
  MUX21X2_HVT U19 ( .A1(n379), .A2(n378), .S0(n310), .Y(n571) );
  INVX0_HVT U20 ( .A(n568), .Y(n347) );
  INVX2_HVT U22 ( .A(n216), .Y(n591) );
  MUX21X2_HVT U23 ( .A1(n305), .A2(n507), .S0(n279), .Y(n506) );
  INVX1_HVT U25 ( .A(n312), .Y(n309) );
  MUX21X1_HVT U26 ( .A1(n462), .A2(n348), .S0(n212), .Y(n461) );
  IBUFFX16_HVT U27 ( .A(n285), .Y(n212) );
  MUX21X2_HVT U28 ( .A1(n505), .A2(n506), .S0(n315), .Y(n503) );
  INVX1_HVT U29 ( .A(n386), .Y(n348) );
  INVX0_HVT U30 ( .A(n347), .Y(n213) );
  MUX21X1_HVT U31 ( .A1(n291), .A2(n262), .S0(n307), .Y(n568) );
  IBUFFX2_HVT U32 ( .A(n312), .Y(n308) );
  MUX41X1_HVT U34 ( .A1(n355), .A3(n562), .A2(n566), .A4(n586), .S0(n316), 
        .S1(n319), .Y(n397) );
  IBUFFX2_HVT U36 ( .A(n316), .Y(n314) );
  IBUFFX2_HVT U37 ( .A(n566), .Y(n349) );
  XNOR2X2_HVT U38 ( .A1(n380), .A2(in[3]), .Y(n216) );
  NAND2X0_HVT U39 ( .A1(n520), .A2(n217), .Y(n218) );
  NAND2X0_HVT U40 ( .A1(n510), .A2(n231), .Y(n219) );
  NAND2X2_HVT U41 ( .A1(n218), .A2(n219), .Y(out[1]) );
  INVX1_HVT U43 ( .A(n231), .Y(n217) );
  IBUFFX2_HVT U44 ( .A(in[6]), .Y(n231) );
  MUX21X2_HVT U45 ( .A1(n272), .A2(n581), .S0(n242), .Y(n400) );
  MUX21X2_HVT U46 ( .A1(n274), .A2(n337), .S0(n282), .Y(n465) );
  NAND2X0_HVT U47 ( .A1(n594), .A2(n232), .Y(n233) );
  NAND2X0_HVT U48 ( .A1(n458), .A2(n241), .Y(n234) );
  NAND2X0_HVT U49 ( .A1(n233), .A2(n234), .Y(n457) );
  INVX0_HVT U50 ( .A(n241), .Y(n232) );
  MUX21X1_HVT U52 ( .A1(n293), .A2(n297), .S0(in[1]), .Y(n575) );
  MUX21X1_HVT U54 ( .A1(n575), .A2(n354), .S0(n289), .Y(n458) );
  IBUFFX2_HVT U55 ( .A(n285), .Y(n241) );
  MUX41X1_HVT U60 ( .A1(n398), .A3(n397), .A2(n396), .A4(n395), .S0(n269), 
        .S1(n256), .Y(n394) );
  NAND2X0_HVT U63 ( .A1(n399), .A2(n235), .Y(n236) );
  NAND2X0_HVT U64 ( .A1(n400), .A2(n284), .Y(n237) );
  NAND2X0_HVT U65 ( .A1(n236), .A2(n237), .Y(n398) );
  IBUFFX2_HVT U67 ( .A(n284), .Y(n235) );
  MUX21X1_HVT U70 ( .A1(n292), .A2(n291), .S0(in[1]), .Y(n581) );
  NAND2X0_HVT U71 ( .A1(n401), .A2(n238), .Y(n239) );
  NAND2X0_HVT U72 ( .A1(n394), .A2(n243), .Y(n240) );
  NAND2X0_HVT U76 ( .A1(n239), .A2(n240), .Y(out[7]) );
  INVX1_HVT U79 ( .A(n243), .Y(n238) );
  MUX41X2_HVT U81 ( .A1(n262), .A3(n595), .A2(n374), .A4(n266), .S0(n315), 
        .S1(n319), .Y(n395) );
  INVX0_HVT U88 ( .A(n296), .Y(n256) );
  OA21X2_HVT U89 ( .A1(n590), .A2(n321), .A3(n353), .Y(n399) );
  IBUFFX2_HVT U91 ( .A(in[6]), .Y(n243) );
  MUX41X1_HVT U92 ( .A1(n585), .A3(n543), .A2(n575), .A4(n350), .S0(n316), 
        .S1(n319), .Y(n396) );
  INVX0_HVT U94 ( .A(n581), .Y(n337) );
  IBUFFX2_HVT U95 ( .A(n312), .Y(n311) );
  INVX1_HVT U99 ( .A(n590), .Y(n332) );
  IBUFFX16_HVT U100 ( .A(n288), .Y(n242) );
  MUX21X2_HVT U102 ( .A1(n404), .A2(n403), .S0(n284), .Y(n402) );
  AND2X1_HVT U104 ( .A1(n309), .A2(n304), .Y(n244) );
  INVX8_HVT U106 ( .A(n244), .Y(n595) );
  NAND2X0_HVT U107 ( .A1(n480), .A2(n245), .Y(n246) );
  NAND2X0_HVT U108 ( .A1(n477), .A2(n269), .Y(n247) );
  NAND2X0_HVT U109 ( .A1(n246), .A2(n247), .Y(n476) );
  IBUFFX2_HVT U111 ( .A(n269), .Y(n245) );
  NBUFFX2_HVT U112 ( .A(n309), .Y(n248) );
  NBUFFX2_HVT U113 ( .A(n309), .Y(n249) );
  NBUFFX2_HVT U114 ( .A(n309), .Y(n250) );
  INVX0_HVT U115 ( .A(in[7]), .Y(n322) );
  INVX1_HVT U116 ( .A(n312), .Y(n310) );
  INVX1_HVT U117 ( .A(n286), .Y(n269) );
  INVX1_HVT U119 ( .A(n322), .Y(n320) );
  INVX0_HVT U120 ( .A(n282), .Y(n251) );
  INVX2_HVT U121 ( .A(in[7]), .Y(n321) );
  MUX41X1_HVT U122 ( .A1(n326), .A3(n303), .A2(n276), .A4(n486), .S0(n251), 
        .S1(n321), .Y(n443) );
  NAND2X0_HVT U124 ( .A1(n325), .A2(n251), .Y(n252) );
  NAND2X0_HVT U126 ( .A1(n475), .A2(n283), .Y(n253) );
  NAND2X0_HVT U127 ( .A1(n252), .A2(n253), .Y(n474) );
  MUX21X2_HVT U129 ( .A1(n470), .A2(n469), .S0(n269), .Y(n468) );
  MUX21X1_HVT U130 ( .A1(n474), .A2(n473), .S0(n290), .Y(n470) );
  MUX21X2_HVT U133 ( .A1(n554), .A2(n529), .S0(n284), .Y(n528) );
  MUX21X2_HVT U134 ( .A1(n409), .A2(n418), .S0(in[6]), .Y(out[6]) );
  INVX1_HVT U137 ( .A(n322), .Y(n254) );
  INVX1_HVT U138 ( .A(n322), .Y(n255) );
  INVX1_HVT U141 ( .A(n322), .Y(n319) );
  INVX1_HVT U143 ( .A(in[2]), .Y(n316) );
  INVX1_HVT U145 ( .A(n274), .Y(n259) );
  INVX0_HVT U149 ( .A(n338), .Y(n258) );
  INVX0_HVT U150 ( .A(n263), .Y(n480) );
  INVX0_HVT U152 ( .A(n343), .Y(n265) );
  OA21X1_HVT U153 ( .A1(n352), .A2(n316), .A3(n339), .Y(n487) );
  XNOR2X1_HVT U155 ( .A1(n308), .A2(in[2]), .Y(n271) );
  INVX0_HVT U156 ( .A(in[6]), .Y(n268) );
  INVX0_HVT U157 ( .A(n567), .Y(n266) );
  INVX0_HVT U161 ( .A(n585), .Y(n264) );
  INVX1_HVT U162 ( .A(n435), .Y(n260) );
  INVX1_HVT U163 ( .A(n257), .Y(n434) );
  MUX41X1_HVT U164 ( .A1(n260), .A3(n259), .A2(n261), .A4(n258), .S0(n316), 
        .S1(n321), .Y(n257) );
  NAND2X0_HVT U169 ( .A1(n591), .A2(n525), .Y(n261) );
  MUX41X1_HVT U171 ( .A1(n349), .A3(n455), .A2(n353), .A4(n573), .S0(n251), 
        .S1(n322), .Y(n454) );
  MUX21X2_HVT U175 ( .A1(n448), .A2(n456), .S0(in[6]), .Y(out[4]) );
  IBUFFX2_HVT U182 ( .A(n380), .Y(n262) );
  INVX1_HVT U183 ( .A(in[4]), .Y(n380) );
  MUX41X1_HVT U185 ( .A1(n344), .A3(n356), .A2(n301), .A4(n354), .S0(n322), 
        .S1(n251), .Y(n417) );
  MUX41X1_HVT U187 ( .A1(n266), .A3(n265), .A2(n267), .A4(n264), .S0(n251), 
        .S1(n321), .Y(n263) );
  NAND2X0_HVT U188 ( .A1(n310), .A2(n293), .Y(n267) );
  MUX21X2_HVT U191 ( .A1(n499), .A2(n489), .S0(n268), .Y(out[2]) );
  MUX41X1_HVT U192 ( .A1(n497), .A3(n492), .A2(n493), .A4(n490), .S0(n256), 
        .S1(n269), .Y(n489) );
  MUX21X2_HVT U194 ( .A1(n498), .A2(n276), .S0(n270), .Y(n497) );
  MUX41X1_HVT U196 ( .A1(n482), .A3(n488), .A2(n484), .A4(n487), .S0(in[5]), 
        .S1(n289), .Y(n481) );
  NBUFFX2_HVT U198 ( .A(in[2]), .Y(n284) );
  NBUFFX2_HVT U200 ( .A(in[2]), .Y(n282) );
  IBUFFX2_HVT U201 ( .A(n316), .Y(n315) );
  MUX21X2_HVT U202 ( .A1(n305), .A2(n483), .S0(n271), .Y(n482) );
  MUX21X2_HVT U203 ( .A1(n535), .A2(n537), .S0(n284), .Y(n534) );
  INVX0_HVT U204 ( .A(in[3]), .Y(n377) );
  MUX21X2_HVT U205 ( .A1(n545), .A2(n549), .S0(n285), .Y(n544) );
  XNOR2X1_HVT U206 ( .A1(n314), .A2(n255), .Y(n270) );
  INVX1_HVT U207 ( .A(n301), .Y(n375) );
  NBUFFX2_HVT U209 ( .A(n216), .Y(n293) );
  NBUFFX2_HVT U210 ( .A(n216), .Y(n292) );
  AND2X1_HVT U211 ( .A1(n216), .A2(n542), .Y(n272) );
  NBUFFX2_HVT U213 ( .A(n593), .Y(n301) );
  INVX1_HVT U217 ( .A(n303), .Y(n379) );
  MUX21X1_HVT U219 ( .A1(n375), .A2(n378), .S0(n318), .Y(n546) );
  MUX21X1_HVT U221 ( .A1(n567), .A2(n486), .S0(n282), .Y(n484) );
  NBUFFX2_HVT U222 ( .A(n593), .Y(n302) );
  MUX21X1_HVT U223 ( .A1(n333), .A2(n376), .S0(n318), .Y(n531) );
  AND2X1_HVT U224 ( .A1(n304), .A2(n525), .Y(n273) );
  MUX21X1_HVT U225 ( .A1(n216), .A2(n378), .S0(n307), .Y(n590) );
  MUX21X1_HVT U226 ( .A1(n304), .A2(n292), .S0(n311), .Y(n557) );
  MUX21X1_HVT U227 ( .A1(n292), .A2(n295), .S0(n48), .Y(n494) );
  MUX21X1_HVT U228 ( .A1(n378), .A2(n293), .S0(n311), .Y(n435) );
  MUX21X1_HVT U229 ( .A1(n302), .A2(n591), .S0(n310), .Y(n561) );
  MUX21X1_HVT U230 ( .A1(n375), .A2(n379), .S0(n250), .Y(n424) );
  MUX21X1_HVT U231 ( .A1(n293), .A2(n375), .S0(n308), .Y(n502) );
  MUX21X1_HVT U232 ( .A1(n591), .A2(n376), .S0(n249), .Y(n384) );
  MUX21X1_HVT U233 ( .A1(n591), .A2(n379), .S0(n249), .Y(n573) );
  MUX21X1_HVT U234 ( .A1(n591), .A2(n295), .S0(n311), .Y(n522) );
  MUX21X1_HVT U235 ( .A1(n302), .A2(n300), .S0(n250), .Y(n509) );
  MUX21X1_HVT U236 ( .A1(n291), .A2(n591), .S0(n307), .Y(n387) );
  MUX21X1_HVT U237 ( .A1(n378), .A2(n375), .S0(n309), .Y(n560) );
  MUX21X1_HVT U238 ( .A1(n291), .A2(n379), .S0(n48), .Y(n558) );
  MUX21X1_HVT U239 ( .A1(n295), .A2(n375), .S0(n48), .Y(n569) );
  MUX21X1_HVT U240 ( .A1(n370), .A2(n300), .S0(n289), .Y(n462) );
  MUX21X1_HVT U241 ( .A1(n478), .A2(n479), .S0(n289), .Y(n477) );
  MUX21X1_HVT U242 ( .A1(n326), .A2(n350), .S0(n282), .Y(n479) );
  NAND2X0_HVT U243 ( .A1(n294), .A2(n377), .Y(n593) );
  MUX21X1_HVT U244 ( .A1(n375), .A2(n294), .S0(n249), .Y(n385) );
  NBUFFX2_HVT U245 ( .A(n596), .Y(n303) );
  MUX21X1_HVT U246 ( .A1(n378), .A2(n291), .S0(n48), .Y(n564) );
  MUX21X1_HVT U247 ( .A1(n376), .A2(n375), .S0(n50), .Y(n579) );
  MUX21X1_HVT U248 ( .A1(n294), .A2(n291), .S0(n249), .Y(n475) );
  NBUFFX2_HVT U249 ( .A(n596), .Y(n304) );
  MUX21X1_HVT U250 ( .A1(n291), .A2(n306), .S0(n308), .Y(n411) );
  MUX21X1_HVT U251 ( .A1(n597), .A2(n304), .S0(n310), .Y(n412) );
  INVX1_HVT U252 ( .A(n298), .Y(n376) );
  INVX1_HVT U253 ( .A(n597), .Y(n378) );
  MUX21X1_HVT U254 ( .A1(n305), .A2(n299), .S0(n50), .Y(n583) );
  MUX21X1_HVT U255 ( .A1(n301), .A2(n306), .S0(n50), .Y(n504) );
  MUX21X1_HVT U256 ( .A1(n291), .A2(n378), .S0(n48), .Y(n587) );
  MUX21X1_HVT U257 ( .A1(n266), .A2(n583), .S0(n315), .Y(n498) );
  NBUFFX2_HVT U258 ( .A(n596), .Y(n305) );
  XOR2X1_HVT U259 ( .A1(n308), .A2(n376), .Y(n553) );
  MUX21X1_HVT U260 ( .A1(n291), .A2(n295), .S0(n248), .Y(n408) );
  XOR2X1_HVT U261 ( .A1(n303), .A2(n248), .Y(n550) );
  XNOR2X1_HVT U262 ( .A1(n301), .A2(n308), .Y(n274) );
  AND2X1_HVT U263 ( .A1(n250), .A2(n379), .Y(n275) );
  MUX21X1_HVT U264 ( .A1(n597), .A2(n299), .S0(n309), .Y(n567) );
  MUX21X1_HVT U265 ( .A1(n302), .A2(n291), .S0(n250), .Y(n586) );
  AND2X1_HVT U266 ( .A1(n306), .A2(n485), .Y(n276) );
  MUX21X1_HVT U267 ( .A1(n303), .A2(n294), .S0(n249), .Y(n391) );
  MUX21X1_HVT U268 ( .A1(n303), .A2(n302), .S0(n308), .Y(n383) );
  XNOR2X1_HVT U269 ( .A1(n306), .A2(n307), .Y(n277) );
  MUX21X1_HVT U270 ( .A1(n299), .A2(n291), .S0(n311), .Y(n389) );
  MUX21X1_HVT U271 ( .A1(n300), .A2(n294), .S0(n310), .Y(n527) );
  MUX21X1_HVT U272 ( .A1(n300), .A2(n306), .S0(n285), .Y(n472) );
  XOR2X1_HVT U273 ( .A1(n294), .A2(n308), .Y(n572) );
  NBUFFX2_HVT U274 ( .A(n289), .Y(n290) );
  NBUFFX2_HVT U275 ( .A(n289), .Y(n288) );
  NBUFFX2_HVT U276 ( .A(in[7]), .Y(n289) );
  NBUFFX2_HVT U277 ( .A(n377), .Y(n291) );
  NBUFFX2_HVT U278 ( .A(in[2]), .Y(n283) );
  NBUFFX2_HVT U279 ( .A(in[2]), .Y(n285) );
  NBUFFX2_HVT U280 ( .A(n318), .Y(n287) );
  NBUFFX2_HVT U281 ( .A(in[2]), .Y(n281) );
  NBUFFX2_HVT U282 ( .A(n317), .Y(n286) );
  MUX21X1_HVT U283 ( .A1(n496), .A2(n348), .S0(n285), .Y(n493) );
  MUX21X1_HVT U284 ( .A1(n415), .A2(n416), .S0(n284), .Y(n414) );
  MUX21X1_HVT U285 ( .A1(n512), .A2(n297), .S0(n289), .Y(n416) );
  XOR2X1_HVT U286 ( .A1(n311), .A2(n297), .Y(n551) );
  MUX21X1_HVT U287 ( .A1(n299), .A2(n292), .S0(n50), .Y(n491) );
  MUX21X1_HVT U288 ( .A1(n519), .A2(n518), .S0(n284), .Y(n516) );
  MUX21X1_HVT U289 ( .A1(n577), .A2(n300), .S0(n290), .Y(n519) );
  MUX21X1_HVT U290 ( .A1(n428), .A2(n427), .S0(n285), .Y(n426) );
  MUX21X1_HVT U291 ( .A1(n300), .A2(n365), .S0(n290), .Y(n428) );
  MUX21X1_HVT U292 ( .A1(n446), .A2(n447), .S0(n281), .Y(n444) );
  MUX21X1_HVT U293 ( .A1(n367), .A2(n376), .S0(n289), .Y(n447) );
  MUX21X1_HVT U294 ( .A1(n376), .A2(n379), .S0(n50), .Y(n433) );
  AND2X1_HVT U295 ( .A1(n216), .A2(n313), .Y(n278) );
  MUX21X1_HVT U296 ( .A1(n297), .A2(n375), .S0(n307), .Y(n559) );
  MUX21X1_HVT U297 ( .A1(n378), .A2(n365), .S0(n290), .Y(n529) );
  XOR2X1_HVT U298 ( .A1(n321), .A2(n571), .Y(n554) );
  MUX21X1_HVT U299 ( .A1(n452), .A2(n451), .S0(n285), .Y(n450) );
  MUX21X1_HVT U300 ( .A1(n569), .A2(n244), .S0(n290), .Y(n452) );
  NAND2X0_HVT U301 ( .A1(in[3]), .A2(n295), .Y(n596) );
  NBUFFX2_HVT U302 ( .A(n380), .Y(n295) );
  MUX21X1_HVT U303 ( .A1(n379), .A2(n297), .S0(n307), .Y(n578) );
  MUX21X1_HVT U304 ( .A1(n351), .A2(n595), .S0(n283), .Y(n488) );
  MUX21X1_HVT U305 ( .A1(n440), .A2(n441), .S0(n283), .Y(n439) );
  MUX21X1_HVT U306 ( .A1(n442), .A2(n305), .S0(n279), .Y(n441) );
  MUX21X1_HVT U307 ( .A1(n560), .A2(n368), .S0(n288), .Y(n440) );
  MUX21X1_HVT U308 ( .A1(n580), .A2(n349), .S0(n283), .Y(n464) );
  MUX21X1_HVT U309 ( .A1(n595), .A2(n312), .S0(n284), .Y(n471) );
  NBUFFX2_HVT U310 ( .A(n588), .Y(n298) );
  MUX21X1_HVT U311 ( .A1(n547), .A2(n548), .S0(n288), .Y(n545) );
  MUX21X1_HVT U312 ( .A1(n297), .A2(n563), .S0(n318), .Y(n548) );
  XOR2X1_HVT U313 ( .A1(n310), .A2(n287), .Y(n555) );
  MUX21X1_HVT U314 ( .A1(n297), .A2(n376), .S0(n310), .Y(n388) );
  NBUFFX2_HVT U315 ( .A(n588), .Y(n299) );
  MUX21X1_HVT U316 ( .A1(n213), .A2(n392), .S0(n288), .Y(n386) );
  MUX21X1_HVT U317 ( .A1(n302), .A2(n297), .S0(n308), .Y(n589) );
  MUX21X1_HVT U318 ( .A1(n335), .A2(n313), .S0(n318), .Y(n533) );
  MUX21X1_HVT U319 ( .A1(n357), .A2(n373), .S0(n289), .Y(n404) );
  MUX21X1_HVT U320 ( .A1(n297), .A2(n294), .S0(n290), .Y(n507) );
  NBUFFX2_HVT U321 ( .A(n597), .Y(n306) );
  NBUFFX2_HVT U322 ( .A(n380), .Y(n294) );
  NBUFFX2_HVT U323 ( .A(n588), .Y(n300) );
  XNOR2X1_HVT U324 ( .A1(n321), .A2(n250), .Y(n279) );
  AND2X1_HVT U325 ( .A1(n291), .A2(n313), .Y(n280) );
  NBUFFX2_HVT U326 ( .A(in[5]), .Y(n318) );
  NBUFFX2_HVT U327 ( .A(in[5]), .Y(n317) );
  MUX21X1_HVT U328 ( .A1(n375), .A2(n262), .S0(n310), .Y(n566) );
  MUX21X1_HVT U329 ( .A1(n262), .A2(n591), .S0(n311), .Y(n390) );
  MUX21X1_HVT U330 ( .A1(n262), .A2(n378), .S0(n48), .Y(n562) );
  MUX21X1_HVT U331 ( .A1(n262), .A2(n376), .S0(n50), .Y(n580) );
  NAND2X0_HVT U332 ( .A1(in[4]), .A2(n377), .Y(n588) );
  NAND2X0_HVT U333 ( .A1(in[3]), .A2(in[4]), .Y(n597) );
  MUX21X1_HVT U334 ( .A1(n262), .A2(n305), .S0(n311), .Y(n577) );
  MUX21X1_HVT U335 ( .A1(n306), .A2(n262), .S0(n311), .Y(n570) );
  MUX21X1_HVT U336 ( .A1(n297), .A2(n262), .S0(n282), .Y(n483) );
  MUX21X1_HVT U337 ( .A1(n262), .A2(n299), .S0(n50), .Y(n382) );
  MUX21X1_HVT U338 ( .A1(n262), .A2(n306), .S0(n307), .Y(n381) );
  INVX0_HVT U339 ( .A(in[1]), .Y(n313) );
  NBUFFX2_HVT U340 ( .A(in[3]), .Y(n297) );
  NBUFFX2_HVT U341 ( .A(in[0]), .Y(n296) );
  INVX0_HVT U342 ( .A(n576), .Y(n323) );
  INVX0_HVT U343 ( .A(n574), .Y(n324) );
  INVX0_HVT U344 ( .A(n565), .Y(n325) );
  INVX0_HVT U345 ( .A(n563), .Y(n326) );
  INVX0_HVT U346 ( .A(n430), .Y(n327) );
  INVX0_HVT U347 ( .A(n393), .Y(n328) );
  INVX0_HVT U348 ( .A(n582), .Y(n329) );
  INVX0_HVT U349 ( .A(n594), .Y(n330) );
  INVX0_HVT U350 ( .A(n592), .Y(n331) );
  INVX0_HVT U351 ( .A(n589), .Y(n333) );
  INVX0_HVT U352 ( .A(n587), .Y(n334) );
  INVX0_HVT U353 ( .A(n586), .Y(n335) );
  INVX0_HVT U354 ( .A(n583), .Y(n336) );
  INVX0_HVT U355 ( .A(n580), .Y(n338) );
  INVX0_HVT U356 ( .A(n579), .Y(n339) );
  INVX0_HVT U357 ( .A(n578), .Y(n340) );
  INVX0_HVT U358 ( .A(n577), .Y(n341) );
  INVX0_HVT U359 ( .A(n575), .Y(n342) );
  INVX0_HVT U360 ( .A(n573), .Y(n343) );
  INVX0_HVT U361 ( .A(n572), .Y(n344) );
  INVX0_HVT U362 ( .A(n570), .Y(n345) );
  INVX0_HVT U363 ( .A(n569), .Y(n346) );
  INVX0_HVT U364 ( .A(n564), .Y(n350) );
  INVX0_HVT U365 ( .A(n562), .Y(n351) );
  INVX0_HVT U366 ( .A(n561), .Y(n352) );
  INVX0_HVT U367 ( .A(n560), .Y(n353) );
  INVX0_HVT U368 ( .A(n559), .Y(n354) );
  INVX0_HVT U369 ( .A(n558), .Y(n355) );
  INVX0_HVT U370 ( .A(n557), .Y(n356) );
  INVX0_HVT U371 ( .A(n556), .Y(n357) );
  INVX0_HVT U372 ( .A(n525), .Y(n358) );
  INVX0_HVT U373 ( .A(n485), .Y(n359) );
  INVX0_HVT U374 ( .A(n392), .Y(n360) );
  INVX0_HVT U375 ( .A(n542), .Y(n361) );
  INVX0_HVT U376 ( .A(n445), .Y(n362) );
  INVX0_HVT U377 ( .A(n391), .Y(n363) );
  INVX0_HVT U378 ( .A(n390), .Y(n364) );
  INVX0_HVT U379 ( .A(n389), .Y(n365) );
  INVX0_HVT U380 ( .A(n388), .Y(n366) );
  INVX0_HVT U381 ( .A(n387), .Y(n367) );
  INVX0_HVT U382 ( .A(n504), .Y(n368) );
  INVX0_HVT U383 ( .A(n494), .Y(n369) );
  INVX0_HVT U384 ( .A(n385), .Y(n370) );
  INVX0_HVT U385 ( .A(n384), .Y(n371) );
  INVX0_HVT U386 ( .A(n383), .Y(n372) );
  INVX0_HVT U387 ( .A(n382), .Y(n373) );
  INVX0_HVT U388 ( .A(n381), .Y(n374) );
endmodule

