
module inv_add_round_keys ( state, subkey, out );
  input [127:0] state;
  input [127:0] subkey;
  output [127:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121;

  XOR2X2_HVT U1 ( .A1(state[9]), .A2(subkey[9]), .Y(out[9]) );
  XOR2X2_HVT U5 ( .A1(state[96]), .A2(subkey[96]), .Y(out[96]) );
  XOR2X2_HVT U6 ( .A1(state[95]), .A2(subkey[95]), .Y(out[95]) );
  XOR2X2_HVT U8 ( .A1(state[93]), .A2(subkey[93]), .Y(out[93]) );
  XOR2X2_HVT U9 ( .A1(subkey[92]), .A2(state[92]), .Y(out[92]) );
  XOR2X2_HVT U12 ( .A1(subkey[8]), .A2(state[8]), .Y(out[8]) );
  XOR2X2_HVT U17 ( .A1(state[85]), .A2(subkey[85]), .Y(out[85]) );
  XOR2X2_HVT U18 ( .A1(state[84]), .A2(subkey[84]), .Y(out[84]) );
  XOR2X2_HVT U19 ( .A1(state[83]), .A2(subkey[83]), .Y(out[83]) );
  XOR2X2_HVT U22 ( .A1(state[80]), .A2(subkey[80]), .Y(out[80]) );
  XOR2X2_HVT U23 ( .A1(state[7]), .A2(subkey[7]), .Y(out[7]) );
  XOR2X2_HVT U24 ( .A1(state[79]), .A2(subkey[79]), .Y(out[79]) );
  XOR2X2_HVT U25 ( .A1(state[78]), .A2(subkey[78]), .Y(out[78]) );
  XOR2X2_HVT U27 ( .A1(subkey[76]), .A2(state[76]), .Y(out[76]) );
  XOR2X2_HVT U28 ( .A1(state[75]), .A2(subkey[75]), .Y(out[75]) );
  XOR2X2_HVT U30 ( .A1(state[73]), .A2(subkey[73]), .Y(out[73]) );
  XOR2X2_HVT U31 ( .A1(state[72]), .A2(subkey[72]), .Y(out[72]) );
  XOR2X2_HVT U32 ( .A1(state[71]), .A2(subkey[71]), .Y(out[71]) );
  XOR2X2_HVT U33 ( .A1(state[70]), .A2(subkey[70]), .Y(out[70]) );
  XOR2X2_HVT U34 ( .A1(state[6]), .A2(subkey[6]), .Y(out[6]) );
  XOR2X2_HVT U35 ( .A1(subkey[69]), .A2(state[69]), .Y(out[69]) );
  XOR2X2_HVT U36 ( .A1(subkey[68]), .A2(state[68]), .Y(out[68]) );
  XOR2X2_HVT U37 ( .A1(state[67]), .A2(subkey[67]), .Y(out[67]) );
  XOR2X2_HVT U38 ( .A1(state[66]), .A2(subkey[66]), .Y(out[66]) );
  XOR2X2_HVT U39 ( .A1(state[65]), .A2(subkey[65]), .Y(out[65]) );
  XOR2X2_HVT U42 ( .A1(state[62]), .A2(subkey[62]), .Y(out[62]) );
  XOR2X2_HVT U43 ( .A1(state[61]), .A2(subkey[61]), .Y(out[61]) );
  XOR2X2_HVT U44 ( .A1(state[60]), .A2(subkey[60]), .Y(out[60]) );
  XOR2X2_HVT U45 ( .A1(state[5]), .A2(subkey[5]), .Y(out[5]) );
  XOR2X2_HVT U47 ( .A1(state[58]), .A2(subkey[58]), .Y(out[58]) );
  XOR2X2_HVT U48 ( .A1(state[57]), .A2(subkey[57]), .Y(out[57]) );
  XOR2X2_HVT U49 ( .A1(state[56]), .A2(subkey[56]), .Y(out[56]) );
  XOR2X2_HVT U50 ( .A1(state[55]), .A2(subkey[55]), .Y(out[55]) );
  XOR2X2_HVT U51 ( .A1(state[54]), .A2(subkey[54]), .Y(out[54]) );
  XOR2X2_HVT U52 ( .A1(state[53]), .A2(subkey[53]), .Y(out[53]) );
  XOR2X2_HVT U53 ( .A1(state[52]), .A2(subkey[52]), .Y(out[52]) );
  XOR2X2_HVT U54 ( .A1(state[51]), .A2(subkey[51]), .Y(out[51]) );
  XOR2X2_HVT U60 ( .A1(state[46]), .A2(subkey[46]), .Y(out[46]) );
  XOR2X2_HVT U62 ( .A1(subkey[44]), .A2(state[44]), .Y(out[44]) );
  XOR2X2_HVT U63 ( .A1(state[43]), .A2(subkey[43]), .Y(out[43]) );
  XOR2X2_HVT U70 ( .A1(state[37]), .A2(subkey[37]), .Y(out[37]) );
  XOR2X2_HVT U71 ( .A1(subkey[36]), .A2(state[36]), .Y(out[36]) );
  XOR2X2_HVT U72 ( .A1(state[35]), .A2(subkey[35]), .Y(out[35]) );
  XOR2X2_HVT U77 ( .A1(state[30]), .A2(subkey[30]), .Y(out[30]) );
  XOR2X2_HVT U80 ( .A1(subkey[28]), .A2(state[28]), .Y(out[28]) );
  XOR2X2_HVT U83 ( .A1(state[25]), .A2(subkey[25]), .Y(out[25]) );
  XOR2X2_HVT U86 ( .A1(state[22]), .A2(subkey[22]), .Y(out[22]) );
  XOR2X2_HVT U87 ( .A1(state[21]), .A2(subkey[21]), .Y(out[21]) );
  XOR2X2_HVT U88 ( .A1(subkey[20]), .A2(state[20]), .Y(out[20]) );
  XOR2X2_HVT U94 ( .A1(state[15]), .A2(subkey[15]), .Y(out[15]) );
  XOR2X2_HVT U96 ( .A1(state[13]), .A2(subkey[13]), .Y(out[13]) );
  XOR2X2_HVT U97 ( .A1(state[12]), .A2(subkey[12]), .Y(out[12]) );
  XOR2X2_HVT U99 ( .A1(state[126]), .A2(subkey[126]), .Y(out[126]) );
  XOR2X2_HVT U101 ( .A1(subkey[124]), .A2(state[124]), .Y(out[124]) );
  XOR2X2_HVT U103 ( .A1(state[122]), .A2(subkey[122]), .Y(out[122]) );
  XOR2X2_HVT U104 ( .A1(subkey[121]), .A2(state[121]), .Y(out[121]) );
  XOR2X2_HVT U106 ( .A1(state[11]), .A2(subkey[11]), .Y(out[11]) );
  XOR2X2_HVT U108 ( .A1(state[118]), .A2(subkey[118]), .Y(out[118]) );
  XOR2X2_HVT U110 ( .A1(state[116]), .A2(subkey[116]), .Y(out[116]) );
  XOR2X2_HVT U111 ( .A1(state[115]), .A2(subkey[115]), .Y(out[115]) );
  XOR2X2_HVT U114 ( .A1(state[112]), .A2(subkey[112]), .Y(out[112]) );
  XOR2X2_HVT U115 ( .A1(state[111]), .A2(subkey[111]), .Y(out[111]) );
  XOR2X2_HVT U118 ( .A1(state[109]), .A2(subkey[109]), .Y(out[109]) );
  XOR2X2_HVT U119 ( .A1(subkey[108]), .A2(state[108]), .Y(out[108]) );
  XOR2X2_HVT U120 ( .A1(state[107]), .A2(subkey[107]), .Y(out[107]) );
  XOR2X2_HVT U121 ( .A1(state[106]), .A2(subkey[106]), .Y(out[106]) );
  XOR2X2_HVT U125 ( .A1(state[102]), .A2(subkey[102]), .Y(out[102]) );
  XOR2X2_HVT U126 ( .A1(state[101]), .A2(subkey[101]), .Y(out[101]) );
  XOR2X2_HVT U127 ( .A1(subkey[100]), .A2(state[100]), .Y(out[100]) );
  XOR2X2_HVT U128 ( .A1(state[0]), .A2(subkey[0]), .Y(out[0]) );
  XOR2X2_HVT U2 ( .A1(state[10]), .A2(subkey[10]), .Y(out[10]) );
  XOR2X2_HVT U3 ( .A1(state[38]), .A2(subkey[38]), .Y(out[38]) );
  XOR2X2_HVT U4 ( .A1(state[104]), .A2(subkey[104]), .Y(out[104]) );
  NAND2X0_HVT U7 ( .A1(state[117]), .A2(n2), .Y(n3) );
  NAND2X0_HVT U10 ( .A1(n1), .A2(subkey[117]), .Y(n4) );
  NAND2X0_HVT U11 ( .A1(n3), .A2(n4), .Y(out[117]) );
  INVX0_HVT U13 ( .A(state[117]), .Y(n1) );
  INVX0_HVT U14 ( .A(subkey[117]), .Y(n2) );
  NAND2X0_HVT U15 ( .A1(state[42]), .A2(n6), .Y(n7) );
  NAND2X0_HVT U16 ( .A1(n5), .A2(subkey[42]), .Y(n8) );
  NAND2X0_HVT U20 ( .A1(n7), .A2(n8), .Y(out[42]) );
  INVX0_HVT U21 ( .A(state[42]), .Y(n5) );
  INVX0_HVT U26 ( .A(subkey[42]), .Y(n6) );
  INVX0_HVT U29 ( .A(state[77]), .Y(n18) );
  XOR2X2_HVT U40 ( .A1(state[24]), .A2(subkey[24]), .Y(out[24]) );
  INVX1_HVT U41 ( .A(state[47]), .Y(n53) );
  INVX0_HVT U46 ( .A(state[119]), .Y(n117) );
  NAND2X0_HVT U55 ( .A1(state[45]), .A2(n10), .Y(n11) );
  NAND2X0_HVT U56 ( .A1(n9), .A2(subkey[45]), .Y(n12) );
  NAND2X0_HVT U57 ( .A1(n11), .A2(n12), .Y(out[45]) );
  INVX0_HVT U58 ( .A(state[45]), .Y(n9) );
  INVX0_HVT U59 ( .A(subkey[45]), .Y(n10) );
  NAND2X0_HVT U61 ( .A1(subkey[2]), .A2(n14), .Y(n15) );
  NAND2X0_HVT U64 ( .A1(n13), .A2(state[2]), .Y(n16) );
  NAND2X0_HVT U65 ( .A1(n15), .A2(n16), .Y(out[2]) );
  IBUFFX2_HVT U66 ( .A(subkey[2]), .Y(n13) );
  INVX0_HVT U67 ( .A(state[2]), .Y(n14) );
  INVX0_HVT U68 ( .A(state[103]), .Y(n109) );
  XOR2X2_HVT U69 ( .A1(state[19]), .A2(subkey[19]), .Y(out[19]) );
  INVX0_HVT U73 ( .A(state[59]), .Y(n86) );
  XNOR2X2_HVT U74 ( .A1(state[88]), .A2(n17), .Y(out[88]) );
  IBUFFX16_HVT U75 ( .A(subkey[88]), .Y(n17) );
  INVX0_HVT U76 ( .A(state[41]), .Y(n105) );
  INVX0_HVT U78 ( .A(state[64]), .Y(n27) );
  NAND2X0_HVT U79 ( .A1(state[77]), .A2(n19), .Y(n20) );
  NAND2X0_HVT U81 ( .A1(n18), .A2(subkey[77]), .Y(n21) );
  NAND2X0_HVT U82 ( .A1(n20), .A2(n21), .Y(out[77]) );
  INVX0_HVT U84 ( .A(subkey[77]), .Y(n19) );
  XNOR2X2_HVT U85 ( .A1(state[33]), .A2(n22), .Y(out[33]) );
  IBUFFX16_HVT U89 ( .A(subkey[33]), .Y(n22) );
  NAND2X0_HVT U90 ( .A1(state[97]), .A2(n24), .Y(n25) );
  NAND2X0_HVT U91 ( .A1(n23), .A2(subkey[97]), .Y(n26) );
  NAND2X0_HVT U92 ( .A1(n25), .A2(n26), .Y(out[97]) );
  INVX1_HVT U93 ( .A(state[97]), .Y(n23) );
  INVX0_HVT U95 ( .A(subkey[97]), .Y(n24) );
  NAND2X0_HVT U98 ( .A1(state[64]), .A2(n39), .Y(n29) );
  NAND2X0_HVT U100 ( .A1(n27), .A2(n28), .Y(n30) );
  NAND2X0_HVT U102 ( .A1(n29), .A2(n30), .Y(out[64]) );
  INVX0_HVT U105 ( .A(n39), .Y(n28) );
  INVX1_HVT U107 ( .A(subkey[64]), .Y(n39) );
  NAND2X0_HVT U109 ( .A1(state[1]), .A2(n32), .Y(n33) );
  NAND2X0_HVT U112 ( .A1(n31), .A2(subkey[1]), .Y(n34) );
  NAND2X0_HVT U113 ( .A1(n33), .A2(n34), .Y(out[1]) );
  INVX0_HVT U116 ( .A(state[1]), .Y(n31) );
  INVX0_HVT U117 ( .A(subkey[1]), .Y(n32) );
  NAND2X0_HVT U122 ( .A1(n36), .A2(state[89]), .Y(n37) );
  NAND2X0_HVT U123 ( .A1(n35), .A2(subkey[89]), .Y(n38) );
  NAND2X0_HVT U124 ( .A1(n37), .A2(n38), .Y(out[89]) );
  INVX1_HVT U129 ( .A(state[89]), .Y(n35) );
  INVX0_HVT U130 ( .A(subkey[89]), .Y(n36) );
  XNOR2X2_HVT U131 ( .A1(state[99]), .A2(n40), .Y(out[99]) );
  IBUFFX16_HVT U132 ( .A(subkey[99]), .Y(n40) );
  INVX1_HVT U133 ( .A(state[39]), .Y(n112) );
  XOR2X2_HVT U134 ( .A1(state[48]), .A2(n41), .Y(out[48]) );
  IBUFFX16_HVT U135 ( .A(n108), .Y(n41) );
  XNOR2X2_HVT U136 ( .A1(state[114]), .A2(n42), .Y(out[114]) );
  IBUFFX16_HVT U137 ( .A(subkey[114]), .Y(n42) );
  INVX1_HVT U138 ( .A(state[127]), .Y(n100) );
  INVX0_HVT U139 ( .A(state[125]), .Y(n47) );
  NAND2X0_HVT U140 ( .A1(n44), .A2(state[87]), .Y(n45) );
  NAND2X0_HVT U141 ( .A1(n43), .A2(subkey[87]), .Y(n46) );
  NAND2X0_HVT U142 ( .A1(n46), .A2(n45), .Y(out[87]) );
  INVX1_HVT U143 ( .A(state[87]), .Y(n43) );
  INVX0_HVT U144 ( .A(subkey[87]), .Y(n44) );
  NAND2X0_HVT U145 ( .A1(n48), .A2(state[125]), .Y(n49) );
  NAND2X0_HVT U146 ( .A1(n47), .A2(subkey[125]), .Y(n50) );
  NAND2X0_HVT U147 ( .A1(n49), .A2(n50), .Y(out[125]) );
  INVX0_HVT U148 ( .A(subkey[125]), .Y(n48) );
  XNOR2X2_HVT U149 ( .A1(state[17]), .A2(n51), .Y(out[17]) );
  IBUFFX16_HVT U150 ( .A(subkey[17]), .Y(n51) );
  XNOR2X2_HVT U151 ( .A1(state[50]), .A2(n52), .Y(out[50]) );
  IBUFFX16_HVT U152 ( .A(subkey[50]), .Y(n52) );
  NAND2X0_HVT U153 ( .A1(n54), .A2(state[47]), .Y(n55) );
  NAND2X0_HVT U154 ( .A1(n53), .A2(subkey[47]), .Y(n56) );
  NAND2X0_HVT U155 ( .A1(n55), .A2(n56), .Y(out[47]) );
  INVX0_HVT U156 ( .A(subkey[47]), .Y(n54) );
  INVX0_HVT U157 ( .A(state[98]), .Y(n61) );
  NAND2X0_HVT U158 ( .A1(n58), .A2(state[18]), .Y(n59) );
  NAND2X0_HVT U159 ( .A1(n57), .A2(subkey[18]), .Y(n60) );
  NAND2X0_HVT U160 ( .A1(n60), .A2(n59), .Y(out[18]) );
  INVX1_HVT U161 ( .A(state[18]), .Y(n57) );
  INVX0_HVT U162 ( .A(subkey[18]), .Y(n58) );
  NAND2X0_HVT U163 ( .A1(state[98]), .A2(n66), .Y(n63) );
  NAND2X0_HVT U164 ( .A1(n61), .A2(n62), .Y(n64) );
  NAND2X0_HVT U165 ( .A1(n63), .A2(n64), .Y(out[98]) );
  INVX0_HVT U166 ( .A(n66), .Y(n62) );
  INVX1_HVT U167 ( .A(subkey[98]), .Y(n66) );
  XNOR2X2_HVT U168 ( .A1(state[90]), .A2(n65), .Y(out[90]) );
  IBUFFX16_HVT U169 ( .A(subkey[90]), .Y(n65) );
  XOR2X2_HVT U170 ( .A1(state[105]), .A2(subkey[105]), .Y(out[105]) );
  INVX1_HVT U171 ( .A(state[31]), .Y(n67) );
  INVX1_HVT U172 ( .A(state[23]), .Y(n82) );
  INVX0_HVT U173 ( .A(subkey[123]), .Y(n98) );
  INVX0_HVT U174 ( .A(subkey[34]), .Y(n77) );
  INVX0_HVT U175 ( .A(subkey[82]), .Y(n121) );
  INVX0_HVT U176 ( .A(subkey[74]), .Y(n99) );
  INVX0_HVT U177 ( .A(subkey[48]), .Y(n108) );
  INVX0_HVT U178 ( .A(subkey[3]), .Y(n71) );
  INVX0_HVT U179 ( .A(subkey[32]), .Y(n72) );
  INVX0_HVT U180 ( .A(subkey[103]), .Y(n116) );
  NAND2X0_HVT U181 ( .A1(n68), .A2(state[31]), .Y(n69) );
  NAND2X0_HVT U182 ( .A1(n67), .A2(subkey[31]), .Y(n70) );
  NAND2X0_HVT U183 ( .A1(n70), .A2(n69), .Y(out[31]) );
  INVX0_HVT U184 ( .A(subkey[31]), .Y(n68) );
  XNOR2X2_HVT U185 ( .A1(state[3]), .A2(n71), .Y(out[3]) );
  INVX0_HVT U186 ( .A(state[110]), .Y(n90) );
  XNOR2X2_HVT U187 ( .A1(state[32]), .A2(n72), .Y(out[32]) );
  NAND2X0_HVT U188 ( .A1(n74), .A2(subkey[29]), .Y(n75) );
  NAND2X0_HVT U189 ( .A1(state[29]), .A2(n73), .Y(n76) );
  NAND2X0_HVT U190 ( .A1(n75), .A2(n76), .Y(out[29]) );
  IBUFFX2_HVT U191 ( .A(subkey[29]), .Y(n73) );
  INVX1_HVT U192 ( .A(state[29]), .Y(n74) );
  XNOR2X2_HVT U193 ( .A1(state[34]), .A2(n77), .Y(out[34]) );
  NAND2X0_HVT U194 ( .A1(n79), .A2(state[16]), .Y(n80) );
  NAND2X0_HVT U195 ( .A1(n78), .A2(subkey[16]), .Y(n81) );
  NAND2X0_HVT U196 ( .A1(n81), .A2(n80), .Y(out[16]) );
  INVX0_HVT U197 ( .A(state[16]), .Y(n78) );
  INVX0_HVT U198 ( .A(subkey[16]), .Y(n79) );
  NAND2X0_HVT U199 ( .A1(n83), .A2(state[23]), .Y(n84) );
  NAND2X0_HVT U200 ( .A1(n82), .A2(subkey[23]), .Y(n85) );
  NAND2X0_HVT U201 ( .A1(n85), .A2(n84), .Y(out[23]) );
  INVX0_HVT U202 ( .A(subkey[23]), .Y(n83) );
  NAND2X0_HVT U203 ( .A1(n87), .A2(state[59]), .Y(n88) );
  NAND2X0_HVT U204 ( .A1(n86), .A2(subkey[59]), .Y(n89) );
  NAND2X0_HVT U205 ( .A1(n88), .A2(n89), .Y(out[59]) );
  INVX0_HVT U206 ( .A(subkey[59]), .Y(n87) );
  XOR2X2_HVT U207 ( .A1(state[14]), .A2(subkey[14]), .Y(out[14]) );
  NAND2X0_HVT U208 ( .A1(n91), .A2(state[110]), .Y(n92) );
  NAND2X0_HVT U209 ( .A1(n90), .A2(subkey[110]), .Y(n93) );
  NAND2X0_HVT U210 ( .A1(n92), .A2(n93), .Y(out[110]) );
  INVX0_HVT U211 ( .A(subkey[110]), .Y(n91) );
  NAND2X0_HVT U212 ( .A1(n95), .A2(subkey[4]), .Y(n96) );
  NAND2X0_HVT U213 ( .A1(state[4]), .A2(n94), .Y(n97) );
  NAND2X0_HVT U214 ( .A1(n96), .A2(n97), .Y(out[4]) );
  INVX0_HVT U215 ( .A(subkey[4]), .Y(n94) );
  INVX1_HVT U216 ( .A(state[4]), .Y(n95) );
  XNOR2X2_HVT U217 ( .A1(state[123]), .A2(n98), .Y(out[123]) );
  XNOR2X2_HVT U218 ( .A1(state[74]), .A2(n99), .Y(out[74]) );
  NAND2X0_HVT U219 ( .A1(n101), .A2(state[127]), .Y(n102) );
  NAND2X0_HVT U220 ( .A1(n100), .A2(subkey[127]), .Y(n103) );
  NAND2X0_HVT U221 ( .A1(n103), .A2(n102), .Y(out[127]) );
  INVX0_HVT U222 ( .A(subkey[127]), .Y(n101) );
  XOR2X2_HVT U223 ( .A1(state[63]), .A2(subkey[63]), .Y(out[63]) );
  NAND2X0_HVT U224 ( .A1(subkey[41]), .A2(n105), .Y(n106) );
  NAND2X0_HVT U225 ( .A1(state[41]), .A2(n104), .Y(n107) );
  NAND2X0_HVT U226 ( .A1(n106), .A2(n107), .Y(out[41]) );
  INVX0_HVT U227 ( .A(subkey[41]), .Y(n104) );
  XOR2X2_HVT U228 ( .A1(state[94]), .A2(subkey[94]), .Y(out[94]) );
  NAND2X0_HVT U229 ( .A1(n116), .A2(state[103]), .Y(n110) );
  NAND2X0_HVT U230 ( .A1(n109), .A2(subkey[103]), .Y(n111) );
  NAND2X0_HVT U231 ( .A1(n111), .A2(n110), .Y(out[103]) );
  NAND2X0_HVT U232 ( .A1(n113), .A2(state[39]), .Y(n114) );
  NAND2X0_HVT U233 ( .A1(n112), .A2(subkey[39]), .Y(n115) );
  NAND2X0_HVT U234 ( .A1(n114), .A2(n115), .Y(out[39]) );
  INVX0_HVT U235 ( .A(subkey[39]), .Y(n113) );
  XOR2X2_HVT U236 ( .A1(state[40]), .A2(subkey[40]), .Y(out[40]) );
  NAND2X0_HVT U237 ( .A1(n118), .A2(state[119]), .Y(n119) );
  NAND2X0_HVT U238 ( .A1(n117), .A2(subkey[119]), .Y(n120) );
  NAND2X0_HVT U239 ( .A1(n120), .A2(n119), .Y(out[119]) );
  INVX0_HVT U240 ( .A(subkey[119]), .Y(n118) );
  XNOR2X2_HVT U241 ( .A1(state[82]), .A2(n121), .Y(out[82]) );
  XOR2X2_HVT U242 ( .A1(state[120]), .A2(subkey[120]), .Y(out[120]) );
  XOR2X2_HVT U243 ( .A1(state[86]), .A2(subkey[86]), .Y(out[86]) );
  XOR2X2_HVT U244 ( .A1(state[26]), .A2(subkey[26]), .Y(out[26]) );
  XOR2X2_HVT U245 ( .A1(state[113]), .A2(subkey[113]), .Y(out[113]) );
  XOR2X2_HVT U246 ( .A1(state[81]), .A2(subkey[81]), .Y(out[81]) );
  XOR2X2_HVT U247 ( .A1(state[91]), .A2(subkey[91]), .Y(out[91]) );
  XOR2X2_HVT U248 ( .A1(state[27]), .A2(subkey[27]), .Y(out[27]) );
  XOR2X2_HVT U249 ( .A1(state[49]), .A2(subkey[49]), .Y(out[49]) );
endmodule

