
module aes ( plaintext, key, clk, reset, start, cipher_text, ready );
  input [127:0] plaintext;
  input [127:0] key;
  output [127:0] cipher_text;
  input clk, reset, start;
  output ready;
  wire   n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, d, n6,
         n7, n8, n9, n11, n12, n13, n14, n15, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n1, n2, n3, n4, n5,
         n10, n16, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n404, n405, n406, n407, n408, n409, n410, n411, n412, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n437,
         n438, n439, n440, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n468, n469, n470, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n483, n484, n485, n486,
         n487, n488, n490, n491, n492, n494, n495, n496, n497, n499, n500,
         n501, n502, n503, n504, n505, n507, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n525,
         n526, n527, n529, n531, n533, n535, n537, n538, n539, n541, n543,
         n544, n545, n546, n548, n550, n551, n552, n553, n554, n555, n557,
         n559, n561, n563, n565, n567, n569, n570, n571, n572, n574, n576,
         n578, n581, n583, n584, n585, n586, n587, n588, n589, n591, n593,
         n595, n596, n597, n598, n600, n602, n604, n606, n608, n609, n610,
         n611, n612, n613, n615, n623, n624, n625, n627, n629, n631, n632,
         n634, n635, n636, n637, n639, n641, n643, n645, n647, n649, n650,
         n651, n653, n654, n655, n657, n659, n661, n662, n663, n664, n666,
         n668, n670, n672, n674, n676, n677, n678, n679, n681, n683, n684,
         n685, n686, n688, n689, n690, n692, n693, n694, n695, n697, n699,
         n701, n703, n704, n705, n707, n709, n711, n713, n714, n715, n716,
         n718, n720, n722, n724, n726, n727, n728, n729, n731, n733, n735,
         n736, n737, n738, n739, n740, n742, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n756, n757, n758, n759, n760, n761,
         n762, n764, n766, n768, n770, n772, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n795, n797, n799, n801, n802, n803, n804, n806,
         n808, n810, n812, n814, n816, n818, n820, n822, n824, n825, n826,
         n827, n834, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915;
  wire   [127:0] adk_out0;
  wire   [127:0] adk_in;
  wire   [3:0] round_number;
  wire   [127:0] key_round;
  wire   [127:0] keyout;
  tri   clk;
  tri   reset;

  DFFX1_HVT d_reg ( .D(n289), .CLK(clk), .Q(d), .QN(n9) );
  DFFX1_HVT \round_number_reg[3]  ( .D(n288), .CLK(clk), .Q(round_number[3])
         );
  DFFX1_HVT \round_number_reg[0]  ( .D(n287), .CLK(clk), .Q(round_number[0]), 
        .QN(n8) );
  DFFX1_HVT \round_number_reg[1]  ( .D(n286), .CLK(clk), .Q(round_number[1]), 
        .QN(n7) );
  DFFX1_HVT \round_number_reg[2]  ( .D(n285), .CLK(clk), .Q(round_number[2]), 
        .QN(n6) );
  DFFX1_HVT \adk_in_reg[0]  ( .D(n284), .CLK(clk), .Q(adk_in[0]) );
  DFFX1_HVT \adk_in_reg[1]  ( .D(n283), .CLK(clk), .Q(adk_in[1]), .QN(n468) );
  DFFX1_HVT \adk_in_reg[2]  ( .D(n282), .CLK(clk), .Q(adk_in[2]) );
  DFFX1_HVT \adk_in_reg[3]  ( .D(n281), .CLK(clk), .Q(adk_in[3]), .QN(n361) );
  DFFX1_HVT \adk_in_reg[4]  ( .D(n280), .CLK(clk), .Q(adk_in[4]), .QN(n537) );
  DFFX1_HVT \adk_in_reg[5]  ( .D(n279), .CLK(clk), .Q(adk_in[5]) );
  DFFX1_HVT \adk_in_reg[6]  ( .D(n278), .CLK(clk), .Q(adk_in[6]) );
  DFFX1_HVT \adk_in_reg[7]  ( .D(n277), .CLK(clk), .Q(adk_in[7]) );
  DFFX1_HVT \adk_in_reg[8]  ( .D(n276), .CLK(clk), .Q(adk_in[8]) );
  DFFX1_HVT \adk_in_reg[9]  ( .D(n275), .CLK(clk), .Q(adk_in[9]) );
  DFFX1_HVT \adk_in_reg[10]  ( .D(n274), .CLK(clk), .Q(adk_in[10]), .QN(n703)
         );
  DFFX1_HVT \adk_in_reg[11]  ( .D(n273), .CLK(clk), .Q(adk_in[11]) );
  DFFX1_HVT \adk_in_reg[12]  ( .D(n272), .CLK(clk), .Q(adk_in[12]), .QN(n407)
         );
  DFFX1_HVT \adk_in_reg[13]  ( .D(n271), .CLK(clk), .Q(adk_in[13]) );
  DFFX1_HVT \adk_in_reg[14]  ( .D(n270), .CLK(clk), .Q(adk_in[14]) );
  DFFX1_HVT \adk_in_reg[15]  ( .D(n269), .CLK(clk), .Q(adk_in[15]) );
  DFFX1_HVT \adk_in_reg[16]  ( .D(n268), .CLK(clk), .Q(adk_in[16]) );
  DFFX1_HVT \adk_in_reg[17]  ( .D(n267), .CLK(clk), .Q(adk_in[17]) );
  DFFX1_HVT \adk_in_reg[18]  ( .D(n266), .CLK(clk), .Q(adk_in[18]) );
  DFFX1_HVT \adk_in_reg[19]  ( .D(n265), .CLK(clk), .Q(adk_in[19]) );
  DFFX1_HVT \adk_in_reg[20]  ( .D(n264), .CLK(clk), .Q(adk_in[20]), .QN(n611)
         );
  DFFX1_HVT \adk_in_reg[21]  ( .D(n263), .CLK(clk), .Q(adk_in[21]) );
  DFFX1_HVT \adk_in_reg[22]  ( .D(n262), .CLK(clk), .Q(adk_in[22]) );
  DFFX1_HVT \adk_in_reg[23]  ( .D(n261), .CLK(clk), .Q(adk_in[23]) );
  DFFX1_HVT \adk_in_reg[24]  ( .D(n260), .CLK(clk), .Q(adk_in[24]) );
  DFFX1_HVT \adk_in_reg[25]  ( .D(n259), .CLK(clk), .Q(adk_in[25]) );
  DFFX1_HVT \adk_in_reg[26]  ( .D(n258), .CLK(clk), .Q(adk_in[26]) );
  DFFX1_HVT \adk_in_reg[27]  ( .D(n257), .CLK(clk), .Q(adk_in[27]) );
  DFFX1_HVT \adk_in_reg[28]  ( .D(n256), .CLK(clk), .Q(adk_in[28]) );
  DFFX1_HVT \adk_in_reg[29]  ( .D(n255), .CLK(clk), .Q(adk_in[29]) );
  DFFX1_HVT \adk_in_reg[30]  ( .D(n254), .CLK(clk), .Q(adk_in[30]) );
  DFFX1_HVT \adk_in_reg[31]  ( .D(n253), .CLK(clk), .Q(adk_in[31]) );
  DFFX1_HVT \adk_in_reg[32]  ( .D(n252), .CLK(clk), .Q(adk_in[32]) );
  DFFX1_HVT \adk_in_reg[33]  ( .D(n251), .CLK(clk), .Q(adk_in[33]), .QN(n381)
         );
  DFFX1_HVT \adk_in_reg[34]  ( .D(n250), .CLK(clk), .Q(adk_in[34]) );
  DFFX1_HVT \adk_in_reg[35]  ( .D(n249), .CLK(clk), .Q(adk_in[35]) );
  DFFX1_HVT \adk_in_reg[36]  ( .D(n248), .CLK(clk), .Q(adk_in[36]) );
  DFFX1_HVT \adk_in_reg[37]  ( .D(n247), .CLK(clk), .Q(adk_in[37]) );
  DFFX1_HVT \adk_in_reg[38]  ( .D(n246), .CLK(clk), .Q(adk_in[38]) );
  DFFX1_HVT \adk_in_reg[39]  ( .D(n245), .CLK(clk), .Q(adk_in[39]), .QN(n623)
         );
  DFFX1_HVT \adk_in_reg[40]  ( .D(n244), .CLK(clk), .Q(adk_in[40]) );
  DFFX1_HVT \adk_in_reg[41]  ( .D(n243), .CLK(clk), .Q(adk_in[41]) );
  DFFX1_HVT \adk_in_reg[42]  ( .D(n242), .CLK(clk), .Q(adk_in[42]) );
  DFFX1_HVT \adk_in_reg[43]  ( .D(n241), .CLK(clk), .Q(adk_in[43]) );
  DFFX1_HVT \adk_in_reg[44]  ( .D(n240), .CLK(clk), .Q(adk_in[44]) );
  DFFX1_HVT \adk_in_reg[45]  ( .D(n239), .CLK(clk), .Q(adk_in[45]) );
  DFFX1_HVT \adk_in_reg[46]  ( .D(n238), .CLK(clk), .Q(adk_in[46]) );
  DFFX1_HVT \adk_in_reg[47]  ( .D(n237), .CLK(clk), .Q(adk_in[47]) );
  DFFX1_HVT \adk_in_reg[48]  ( .D(n236), .CLK(clk), .Q(adk_in[48]) );
  DFFX1_HVT \adk_in_reg[49]  ( .D(n235), .CLK(clk), .Q(adk_in[49]), .QN(n309)
         );
  DFFX1_HVT \adk_in_reg[50]  ( .D(n234), .CLK(clk), .Q(adk_in[50]) );
  DFFX1_HVT \adk_in_reg[51]  ( .D(n233), .CLK(clk), .Q(adk_in[51]) );
  DFFX1_HVT \adk_in_reg[52]  ( .D(n232), .CLK(clk), .Q(adk_in[52]), .QN(n635)
         );
  DFFX1_HVT \adk_in_reg[53]  ( .D(n231), .CLK(clk), .Q(adk_in[53]) );
  DFFX1_HVT \adk_in_reg[54]  ( .D(n230), .CLK(clk), .Q(adk_in[54]) );
  DFFX1_HVT \adk_in_reg[55]  ( .D(n229), .CLK(clk), .Q(adk_in[55]) );
  DFFX1_HVT \adk_in_reg[56]  ( .D(n228), .CLK(clk), .Q(adk_in[56]) );
  DFFX1_HVT \adk_in_reg[57]  ( .D(n227), .CLK(clk), .Q(adk_in[57]) );
  DFFX1_HVT \adk_in_reg[58]  ( .D(n226), .CLK(clk), .Q(adk_in[58]) );
  DFFX1_HVT \adk_in_reg[59]  ( .D(n225), .CLK(clk), .Q(adk_in[59]) );
  DFFX1_HVT \adk_in_reg[60]  ( .D(n224), .CLK(clk), .Q(adk_in[60]), .QN(n634)
         );
  DFFX1_HVT \adk_in_reg[61]  ( .D(n223), .CLK(clk), .Q(adk_in[61]) );
  DFFX1_HVT \adk_in_reg[62]  ( .D(n222), .CLK(clk), .Q(adk_in[62]) );
  DFFX1_HVT \adk_in_reg[63]  ( .D(n221), .CLK(clk), .Q(adk_in[63]), .QN(n649)
         );
  DFFX1_HVT \adk_in_reg[64]  ( .D(n220), .CLK(clk), .Q(adk_in[64]) );
  DFFX1_HVT \adk_in_reg[65]  ( .D(n219), .CLK(clk), .Q(adk_in[65]) );
  DFFX1_HVT \adk_in_reg[66]  ( .D(n218), .CLK(clk), .Q(adk_in[66]), .QN(n351)
         );
  DFFX1_HVT \adk_in_reg[67]  ( .D(n217), .CLK(clk), .Q(adk_in[67]) );
  DFFX1_HVT \adk_in_reg[68]  ( .D(n216), .CLK(clk), .Q(adk_in[68]) );
  DFFX1_HVT \adk_in_reg[69]  ( .D(n215), .CLK(clk), .Q(adk_in[69]) );
  DFFX1_HVT \adk_in_reg[70]  ( .D(n214), .CLK(clk), .Q(adk_in[70]) );
  DFFX1_HVT \adk_in_reg[71]  ( .D(n213), .CLK(clk), .Q(adk_in[71]) );
  DFFX1_HVT \adk_in_reg[72]  ( .D(n212), .CLK(clk), .Q(adk_in[72]) );
  DFFX1_HVT \adk_in_reg[73]  ( .D(n211), .CLK(clk), .Q(adk_in[73]) );
  DFFX1_HVT \adk_in_reg[74]  ( .D(n210), .CLK(clk), .Q(adk_in[74]) );
  DFFX1_HVT \adk_in_reg[75]  ( .D(n209), .CLK(clk), .Q(adk_in[75]) );
  DFFX1_HVT \adk_in_reg[76]  ( .D(n208), .CLK(clk), .Q(adk_in[76]), .QN(n490)
         );
  DFFX1_HVT \adk_in_reg[78]  ( .D(n206), .CLK(clk), .Q(adk_in[78]) );
  DFFX1_HVT \adk_in_reg[79]  ( .D(n205), .CLK(clk), .Q(adk_in[79]) );
  DFFX1_HVT \adk_in_reg[80]  ( .D(n204), .CLK(clk), .Q(adk_in[80]) );
  DFFX1_HVT \adk_in_reg[81]  ( .D(n203), .CLK(clk), .Q(adk_in[81]), .QN(n483)
         );
  DFFX1_HVT \adk_in_reg[82]  ( .D(n202), .CLK(clk), .Q(adk_in[82]) );
  DFFX1_HVT \adk_in_reg[83]  ( .D(n201), .CLK(clk), .Q(adk_in[83]), .QN(n342)
         );
  DFFX1_HVT \adk_in_reg[84]  ( .D(n200), .CLK(clk), .Q(adk_in[84]), .QN(n365)
         );
  DFFX1_HVT \adk_in_reg[85]  ( .D(n199), .CLK(clk), .Q(adk_in[85]) );
  DFFX1_HVT \adk_in_reg[86]  ( .D(n198), .CLK(clk), .Q(adk_in[86]) );
  DFFX1_HVT \adk_in_reg[87]  ( .D(n197), .CLK(clk), .Q(adk_in[87]) );
  DFFX1_HVT \adk_in_reg[88]  ( .D(n196), .CLK(clk), .Q(adk_in[88]) );
  DFFX1_HVT \adk_in_reg[89]  ( .D(n195), .CLK(clk), .Q(adk_in[89]), .QN(n461)
         );
  DFFX1_HVT \adk_in_reg[90]  ( .D(n194), .CLK(clk), .Q(adk_in[90]) );
  DFFX1_HVT \adk_in_reg[91]  ( .D(n193), .CLK(clk), .Q(adk_in[91]) );
  DFFX1_HVT \adk_in_reg[92]  ( .D(n192), .CLK(clk), .Q(adk_in[92]) );
  DFFX1_HVT \adk_in_reg[93]  ( .D(n191), .CLK(clk), .Q(adk_in[93]) );
  DFFX1_HVT \adk_in_reg[94]  ( .D(n190), .CLK(clk), .Q(adk_in[94]) );
  DFFX1_HVT \adk_in_reg[95]  ( .D(n189), .CLK(clk), .Q(adk_in[95]) );
  DFFX1_HVT \adk_in_reg[96]  ( .D(n188), .CLK(clk), .Q(adk_in[96]) );
  DFFX1_HVT \adk_in_reg[97]  ( .D(n187), .CLK(clk), .Q(adk_in[97]), .QN(n448)
         );
  DFFX1_HVT \adk_in_reg[98]  ( .D(n186), .CLK(clk), .Q(adk_in[98]) );
  DFFX1_HVT \adk_in_reg[99]  ( .D(n185), .CLK(clk), .Q(adk_in[99]) );
  DFFX1_HVT \adk_in_reg[100]  ( .D(n184), .CLK(clk), .Q(adk_in[100]) );
  DFFX1_HVT \adk_in_reg[101]  ( .D(n183), .CLK(clk), .Q(adk_in[101]) );
  DFFX1_HVT \adk_in_reg[102]  ( .D(n182), .CLK(clk), .Q(adk_in[102]) );
  DFFX1_HVT \adk_in_reg[103]  ( .D(n181), .CLK(clk), .Q(adk_in[103]) );
  DFFX1_HVT \adk_in_reg[104]  ( .D(n180), .CLK(clk), .Q(adk_in[104]) );
  DFFX1_HVT \adk_in_reg[105]  ( .D(n179), .CLK(clk), .Q(adk_in[105]) );
  DFFX1_HVT \adk_in_reg[106]  ( .D(n178), .CLK(clk), .Q(adk_in[106]) );
  DFFX1_HVT \adk_in_reg[107]  ( .D(n177), .CLK(clk), .Q(adk_in[107]) );
  DFFX1_HVT \adk_in_reg[108]  ( .D(n176), .CLK(clk), .Q(adk_in[108]) );
  DFFX1_HVT \adk_in_reg[109]  ( .D(n175), .CLK(clk), .Q(adk_in[109]) );
  DFFX1_HVT \adk_in_reg[111]  ( .D(n173), .CLK(clk), .Q(adk_in[111]), .QN(n525) );
  DFFX1_HVT \adk_in_reg[112]  ( .D(n172), .CLK(clk), .Q(adk_in[112]) );
  DFFX1_HVT \adk_in_reg[113]  ( .D(n171), .CLK(clk), .Q(adk_in[113]), .QN(n370) );
  DFFX1_HVT \adk_in_reg[114]  ( .D(n170), .CLK(clk), .Q(adk_in[114]) );
  DFFX1_HVT \adk_in_reg[115]  ( .D(n169), .CLK(clk), .Q(adk_in[115]) );
  DFFX1_HVT \adk_in_reg[116]  ( .D(n168), .CLK(clk), .Q(adk_in[116]) );
  DFFX1_HVT \adk_in_reg[117]  ( .D(n167), .CLK(clk), .Q(adk_in[117]) );
  DFFX1_HVT \adk_in_reg[118]  ( .D(n166), .CLK(clk), .Q(adk_in[118]) );
  DFFX1_HVT \adk_in_reg[119]  ( .D(n165), .CLK(clk), .Q(adk_in[119]) );
  DFFX1_HVT \adk_in_reg[120]  ( .D(n164), .CLK(clk), .Q(adk_in[120]) );
  DFFX1_HVT \adk_in_reg[121]  ( .D(n163), .CLK(clk), .Q(adk_in[121]), .QN(n518) );
  DFFX1_HVT \adk_in_reg[122]  ( .D(n162), .CLK(clk), .Q(adk_in[122]), .QN(n738) );
  DFFX1_HVT \adk_in_reg[123]  ( .D(n161), .CLK(clk), .Q(adk_in[123]) );
  DFFX1_HVT \adk_in_reg[124]  ( .D(n160), .CLK(clk), .Q(adk_in[124]) );
  DFFX1_HVT \adk_in_reg[125]  ( .D(n159), .CLK(clk), .Q(adk_in[125]) );
  DFFX1_HVT \adk_in_reg[126]  ( .D(n158), .CLK(clk), .Q(adk_in[126]) );
  DFFX1_HVT \adk_in_reg[127]  ( .D(n157), .CLK(clk), .Q(adk_in[127]), .QN(n367) );
  DFFX1_HVT \key_round_reg[0]  ( .D(n156), .CLK(clk), .Q(key_round[0]) );
  DFFX1_HVT \key_round_reg[1]  ( .D(n155), .CLK(clk), .Q(key_round[1]), .QN(
        n368) );
  DFFX1_HVT \key_round_reg[2]  ( .D(n154), .CLK(clk), .Q(key_round[2]), .QN(
        n653) );
  DFFX1_HVT \key_round_reg[3]  ( .D(n153), .CLK(clk), .Q(key_round[3]) );
  DFFX1_HVT \key_round_reg[4]  ( .D(n152), .CLK(clk), .Q(key_round[4]) );
  DFFX1_HVT \key_round_reg[5]  ( .D(n151), .CLK(clk), .Q(key_round[5]) );
  DFFX1_HVT \key_round_reg[6]  ( .D(n150), .CLK(clk), .Q(key_round[6]) );
  DFFX1_HVT \key_round_reg[7]  ( .D(n149), .CLK(clk), .Q(key_round[7]), .QN(
        n363) );
  DFFX1_HVT \key_round_reg[8]  ( .D(n148), .CLK(clk), .Q(key_round[8]) );
  DFFX1_HVT \key_round_reg[9]  ( .D(n147), .CLK(clk), .Q(key_round[9]) );
  DFFX1_HVT \key_round_reg[10]  ( .D(n146), .CLK(clk), .Q(key_round[10]), .QN(
        n688) );
  DFFX1_HVT \key_round_reg[11]  ( .D(n145), .CLK(clk), .Q(key_round[11]) );
  DFFX1_HVT \key_round_reg[12]  ( .D(n144), .CLK(clk), .Q(key_round[12]) );
  DFFX1_HVT \key_round_reg[13]  ( .D(n143), .CLK(clk), .Q(key_round[13]) );
  DFFX1_HVT \key_round_reg[14]  ( .D(n142), .CLK(clk), .Q(key_round[14]) );
  DFFX1_HVT \key_round_reg[15]  ( .D(n141), .CLK(clk), .Q(key_round[15]), .QN(
        n550) );
  DFFX1_HVT \key_round_reg[16]  ( .D(n140), .CLK(clk), .Q(key_round[16]) );
  DFFX1_HVT \key_round_reg[17]  ( .D(n139), .CLK(clk), .Q(key_round[17]) );
  DFFX1_HVT \key_round_reg[18]  ( .D(n138), .CLK(clk), .Q(key_round[18]), .QN(
        n387) );
  DFFX1_HVT \key_round_reg[19]  ( .D(n137), .CLK(clk), .Q(key_round[19]) );
  DFFX1_HVT \key_round_reg[20]  ( .D(n136), .CLK(clk), .Q(key_round[20]) );
  DFFX1_HVT \key_round_reg[21]  ( .D(n135), .CLK(clk), .Q(key_round[21]) );
  DFFX1_HVT \key_round_reg[22]  ( .D(n134), .CLK(clk), .Q(key_round[22]) );
  DFFX1_HVT \key_round_reg[23]  ( .D(n133), .CLK(clk), .Q(key_round[23]) );
  DFFX1_HVT \key_round_reg[24]  ( .D(n132), .CLK(clk), .Q(key_round[24]) );
  DFFX1_HVT \key_round_reg[25]  ( .D(n131), .CLK(clk), .Q(key_round[25]) );
  DFFX1_HVT \key_round_reg[26]  ( .D(n130), .CLK(clk), .Q(key_round[26]) );
  DFFX1_HVT \key_round_reg[27]  ( .D(n129), .CLK(clk), .Q(key_round[27]) );
  DFFX1_HVT \key_round_reg[28]  ( .D(n128), .CLK(clk), .Q(key_round[28]) );
  DFFX1_HVT \key_round_reg[29]  ( .D(n127), .CLK(clk), .Q(key_round[29]) );
  DFFX1_HVT \key_round_reg[30]  ( .D(n126), .CLK(clk), .Q(key_round[30]) );
  DFFX1_HVT \key_round_reg[31]  ( .D(n125), .CLK(clk), .Q(key_round[31]) );
  DFFX1_HVT \key_round_reg[32]  ( .D(n124), .CLK(clk), .Q(key_round[32]) );
  DFFX1_HVT \key_round_reg[33]  ( .D(n123), .CLK(clk), .Q(key_round[33]) );
  DFFX1_HVT \key_round_reg[34]  ( .D(n122), .CLK(clk), .Q(key_round[34]) );
  DFFX1_HVT \key_round_reg[35]  ( .D(n121), .CLK(clk), .Q(key_round[35]) );
  DFFX1_HVT \key_round_reg[36]  ( .D(n120), .CLK(clk), .Q(key_round[36]) );
  DFFX1_HVT \key_round_reg[37]  ( .D(n119), .CLK(clk), .Q(key_round[37]) );
  DFFX1_HVT \key_round_reg[38]  ( .D(n118), .CLK(clk), .Q(key_round[38]) );
  DFFX1_HVT \key_round_reg[39]  ( .D(n117), .CLK(clk), .Q(key_round[39]) );
  DFFX1_HVT \key_round_reg[40]  ( .D(n116), .CLK(clk), .Q(key_round[40]) );
  DFFX1_HVT \key_round_reg[41]  ( .D(n115), .CLK(clk), .Q(key_round[41]) );
  DFFX1_HVT \key_round_reg[42]  ( .D(n114), .CLK(clk), .Q(key_round[42]) );
  DFFX1_HVT \key_round_reg[43]  ( .D(n113), .CLK(clk), .Q(key_round[43]) );
  DFFX1_HVT \key_round_reg[44]  ( .D(n112), .CLK(clk), .Q(key_round[44]) );
  DFFX1_HVT \key_round_reg[45]  ( .D(n111), .CLK(clk), .Q(key_round[45]) );
  DFFX1_HVT \key_round_reg[46]  ( .D(n110), .CLK(clk), .Q(key_round[46]) );
  DFFX1_HVT \key_round_reg[47]  ( .D(n109), .CLK(clk), .Q(key_round[47]) );
  DFFX1_HVT \key_round_reg[48]  ( .D(n108), .CLK(clk), .Q(key_round[48]) );
  DFFX1_HVT \key_round_reg[49]  ( .D(n107), .CLK(clk), .Q(key_round[49]) );
  DFFX1_HVT \key_round_reg[50]  ( .D(n106), .CLK(clk), .Q(key_round[50]) );
  DFFX1_HVT \key_round_reg[51]  ( .D(n105), .CLK(clk), .Q(key_round[51]) );
  DFFX1_HVT \key_round_reg[52]  ( .D(n104), .CLK(clk), .Q(key_round[52]) );
  DFFX1_HVT \key_round_reg[53]  ( .D(n103), .CLK(clk), .Q(key_round[53]) );
  DFFX1_HVT \key_round_reg[54]  ( .D(n102), .CLK(clk), .Q(key_round[54]) );
  DFFX1_HVT \key_round_reg[55]  ( .D(n101), .CLK(clk), .Q(key_round[55]) );
  DFFX1_HVT \key_round_reg[56]  ( .D(n100), .CLK(clk), .Q(key_round[56]) );
  DFFX1_HVT \key_round_reg[57]  ( .D(n99), .CLK(clk), .Q(key_round[57]) );
  DFFX1_HVT \key_round_reg[58]  ( .D(n98), .CLK(clk), .Q(key_round[58]) );
  DFFX1_HVT \key_round_reg[59]  ( .D(n97), .CLK(clk), .Q(key_round[59]) );
  DFFX1_HVT \key_round_reg[60]  ( .D(n96), .CLK(clk), .Q(key_round[60]) );
  DFFX1_HVT \key_round_reg[61]  ( .D(n95), .CLK(clk), .Q(key_round[61]) );
  DFFX1_HVT \key_round_reg[62]  ( .D(n94), .CLK(clk), .Q(key_round[62]) );
  DFFX1_HVT \key_round_reg[63]  ( .D(n93), .CLK(clk), .Q(key_round[63]) );
  DFFX1_HVT \key_round_reg[64]  ( .D(n92), .CLK(clk), .Q(key_round[64]) );
  DFFX1_HVT \key_round_reg[65]  ( .D(n91), .CLK(clk), .Q(key_round[65]) );
  DFFX1_HVT \key_round_reg[66]  ( .D(n90), .CLK(clk), .Q(key_round[66]) );
  DFFX1_HVT \key_round_reg[67]  ( .D(n89), .CLK(clk), .Q(key_round[67]) );
  DFFX1_HVT \key_round_reg[68]  ( .D(n88), .CLK(clk), .Q(key_round[68]) );
  DFFX1_HVT \key_round_reg[69]  ( .D(n87), .CLK(clk), .Q(key_round[69]) );
  DFFX1_HVT \key_round_reg[70]  ( .D(n86), .CLK(clk), .Q(key_round[70]) );
  DFFX1_HVT \key_round_reg[71]  ( .D(n85), .CLK(clk), .Q(key_round[71]) );
  DFFX1_HVT \key_round_reg[72]  ( .D(n84), .CLK(clk), .Q(key_round[72]) );
  DFFX1_HVT \key_round_reg[73]  ( .D(n83), .CLK(clk), .Q(key_round[73]) );
  DFFX1_HVT \key_round_reg[74]  ( .D(n82), .CLK(clk), .Q(key_round[74]) );
  DFFX1_HVT \key_round_reg[75]  ( .D(n81), .CLK(clk), .Q(key_round[75]) );
  DFFX1_HVT \key_round_reg[76]  ( .D(n80), .CLK(clk), .Q(key_round[76]) );
  DFFX1_HVT \key_round_reg[77]  ( .D(n79), .CLK(clk), .Q(key_round[77]) );
  DFFX1_HVT \key_round_reg[78]  ( .D(n78), .CLK(clk), .Q(key_round[78]) );
  DFFX1_HVT \key_round_reg[79]  ( .D(n77), .CLK(clk), .Q(key_round[79]) );
  DFFX1_HVT \key_round_reg[80]  ( .D(n76), .CLK(clk), .Q(key_round[80]) );
  DFFX1_HVT \key_round_reg[81]  ( .D(n75), .CLK(clk), .Q(key_round[81]) );
  DFFX1_HVT \key_round_reg[82]  ( .D(n74), .CLK(clk), .Q(key_round[82]) );
  DFFX1_HVT \key_round_reg[83]  ( .D(n73), .CLK(clk), .Q(key_round[83]) );
  DFFX1_HVT \key_round_reg[84]  ( .D(n72), .CLK(clk), .Q(key_round[84]) );
  DFFX1_HVT \key_round_reg[85]  ( .D(n71), .CLK(clk), .Q(key_round[85]) );
  DFFX1_HVT \key_round_reg[86]  ( .D(n70), .CLK(clk), .Q(key_round[86]) );
  DFFX1_HVT \key_round_reg[87]  ( .D(n69), .CLK(clk), .Q(key_round[87]) );
  DFFX1_HVT \key_round_reg[88]  ( .D(n68), .CLK(clk), .Q(key_round[88]) );
  DFFX1_HVT \key_round_reg[89]  ( .D(n67), .CLK(clk), .Q(key_round[89]) );
  DFFX1_HVT \key_round_reg[90]  ( .D(n66), .CLK(clk), .Q(key_round[90]) );
  DFFX1_HVT \key_round_reg[91]  ( .D(n65), .CLK(clk), .Q(key_round[91]) );
  DFFX1_HVT \key_round_reg[92]  ( .D(n64), .CLK(clk), .Q(key_round[92]) );
  DFFX1_HVT \key_round_reg[93]  ( .D(n63), .CLK(clk), .Q(key_round[93]) );
  DFFX1_HVT \key_round_reg[94]  ( .D(n62), .CLK(clk), .Q(key_round[94]) );
  DFFX1_HVT \key_round_reg[95]  ( .D(n61), .CLK(clk), .Q(key_round[95]) );
  DFFX1_HVT \key_round_reg[96]  ( .D(n60), .CLK(clk), .Q(key_round[96]) );
  DFFX1_HVT \key_round_reg[97]  ( .D(n59), .CLK(clk), .Q(key_round[97]) );
  DFFX1_HVT \key_round_reg[98]  ( .D(n58), .CLK(clk), .Q(key_round[98]) );
  DFFX1_HVT \key_round_reg[99]  ( .D(n57), .CLK(clk), .Q(key_round[99]) );
  DFFX1_HVT \key_round_reg[100]  ( .D(n56), .CLK(clk), .Q(key_round[100]) );
  DFFX1_HVT \key_round_reg[101]  ( .D(n55), .CLK(clk), .Q(key_round[101]) );
  DFFX1_HVT \key_round_reg[102]  ( .D(n54), .CLK(clk), .Q(key_round[102]) );
  DFFX1_HVT \key_round_reg[103]  ( .D(n53), .CLK(clk), .Q(key_round[103]) );
  DFFX1_HVT \key_round_reg[104]  ( .D(n52), .CLK(clk), .Q(key_round[104]) );
  DFFX1_HVT \key_round_reg[105]  ( .D(n51), .CLK(clk), .Q(key_round[105]) );
  DFFX1_HVT \key_round_reg[106]  ( .D(n50), .CLK(clk), .Q(key_round[106]) );
  DFFX1_HVT \key_round_reg[107]  ( .D(n49), .CLK(clk), .Q(key_round[107]) );
  DFFX1_HVT \key_round_reg[108]  ( .D(n48), .CLK(clk), .Q(key_round[108]) );
  DFFX1_HVT \key_round_reg[109]  ( .D(n47), .CLK(clk), .Q(key_round[109]) );
  DFFX1_HVT \key_round_reg[110]  ( .D(n46), .CLK(clk), .Q(key_round[110]) );
  DFFX1_HVT \key_round_reg[111]  ( .D(n45), .CLK(clk), .Q(key_round[111]) );
  DFFX1_HVT \key_round_reg[112]  ( .D(n44), .CLK(clk), .Q(key_round[112]) );
  DFFX1_HVT \key_round_reg[113]  ( .D(n43), .CLK(clk), .Q(key_round[113]) );
  DFFX1_HVT \key_round_reg[114]  ( .D(n42), .CLK(clk), .Q(key_round[114]) );
  DFFX1_HVT \key_round_reg[115]  ( .D(n41), .CLK(clk), .Q(key_round[115]) );
  DFFX1_HVT \key_round_reg[116]  ( .D(n40), .CLK(clk), .Q(key_round[116]) );
  DFFX1_HVT \key_round_reg[117]  ( .D(n39), .CLK(clk), .Q(key_round[117]) );
  DFFX1_HVT \key_round_reg[118]  ( .D(n38), .CLK(clk), .Q(key_round[118]) );
  DFFX1_HVT \key_round_reg[119]  ( .D(n37), .CLK(clk), .Q(key_round[119]) );
  DFFX1_HVT \key_round_reg[120]  ( .D(n36), .CLK(clk), .Q(key_round[120]) );
  DFFX1_HVT \key_round_reg[121]  ( .D(n35), .CLK(clk), .Q(key_round[121]) );
  DFFX1_HVT \key_round_reg[122]  ( .D(n34), .CLK(clk), .Q(key_round[122]) );
  DFFX1_HVT \key_round_reg[123]  ( .D(n33), .CLK(clk), .Q(key_round[123]) );
  DFFX1_HVT \key_round_reg[124]  ( .D(n32), .CLK(clk), .Q(key_round[124]) );
  DFFX1_HVT \key_round_reg[125]  ( .D(n31), .CLK(clk), .Q(key_round[125]) );
  DFFX1_HVT \key_round_reg[126]  ( .D(n30), .CLK(clk), .Q(key_round[126]) );
  DFFX1_HVT \key_round_reg[127]  ( .D(n29), .CLK(clk), .Q(key_round[127]) );
  DFFX1_HVT ready_reg ( .D(n28), .CLK(clk), .Q(ready) );
  NOR4X1_HVT U3 ( .A1(round_number[0]), .A2(round_number[1]), .A3(
        round_number[2]), .A4(round_number[3]), .Y(n18) );
  AO22X1_HVT U8 ( .A1(n11), .A2(ready), .A3(n913), .A4(n915), .Y(n28) );
  AND2X1_HVT U9 ( .A1(n13), .A2(n14), .Y(n11) );
  AO222X1_HVT U10 ( .A1(keyout[127]), .A2(n887), .A3(key[127]), .A4(n861), 
        .A5(key_round[127]), .A6(n856), .Y(n29) );
  AO222X1_HVT U11 ( .A1(keyout[126]), .A2(n887), .A3(key[126]), .A4(n861), 
        .A5(key_round[126]), .A6(n856), .Y(n30) );
  AO222X1_HVT U12 ( .A1(keyout[125]), .A2(n887), .A3(key[125]), .A4(n861), 
        .A5(key_round[125]), .A6(n856), .Y(n31) );
  AO222X1_HVT U13 ( .A1(keyout[124]), .A2(n887), .A3(key[124]), .A4(n861), 
        .A5(key_round[124]), .A6(n856), .Y(n32) );
  AO222X1_HVT U14 ( .A1(keyout[123]), .A2(n887), .A3(key[123]), .A4(n861), 
        .A5(key_round[123]), .A6(n856), .Y(n33) );
  AO222X1_HVT U15 ( .A1(keyout[122]), .A2(n887), .A3(key[122]), .A4(n861), 
        .A5(key_round[122]), .A6(n856), .Y(n34) );
  AO222X1_HVT U16 ( .A1(keyout[121]), .A2(n887), .A3(key[121]), .A4(n861), 
        .A5(key_round[121]), .A6(n856), .Y(n35) );
  AO222X1_HVT U17 ( .A1(keyout[120]), .A2(n887), .A3(key[120]), .A4(n861), 
        .A5(key_round[120]), .A6(n856), .Y(n36) );
  AO222X1_HVT U18 ( .A1(keyout[119]), .A2(n887), .A3(key[119]), .A4(n861), 
        .A5(key_round[119]), .A6(n856), .Y(n37) );
  AO222X1_HVT U19 ( .A1(keyout[118]), .A2(n887), .A3(key[118]), .A4(n861), 
        .A5(key_round[118]), .A6(n856), .Y(n38) );
  AO222X1_HVT U20 ( .A1(keyout[117]), .A2(n887), .A3(key[117]), .A4(n861), 
        .A5(key_round[117]), .A6(n855), .Y(n39) );
  AO222X1_HVT U21 ( .A1(keyout[116]), .A2(n887), .A3(key[116]), .A4(n861), 
        .A5(key_round[116]), .A6(n855), .Y(n40) );
  AO222X1_HVT U22 ( .A1(keyout[115]), .A2(n888), .A3(key[115]), .A4(n862), 
        .A5(key_round[115]), .A6(n855), .Y(n41) );
  AO222X1_HVT U23 ( .A1(keyout[114]), .A2(n888), .A3(key[114]), .A4(n862), 
        .A5(key_round[114]), .A6(n855), .Y(n42) );
  AO222X1_HVT U24 ( .A1(keyout[113]), .A2(n888), .A3(key[113]), .A4(n862), 
        .A5(key_round[113]), .A6(n855), .Y(n43) );
  AO222X1_HVT U25 ( .A1(keyout[112]), .A2(n888), .A3(key[112]), .A4(n862), 
        .A5(key_round[112]), .A6(n855), .Y(n44) );
  AO222X1_HVT U26 ( .A1(keyout[111]), .A2(n888), .A3(key[111]), .A4(n862), 
        .A5(key_round[111]), .A6(n855), .Y(n45) );
  AO222X1_HVT U27 ( .A1(keyout[110]), .A2(n888), .A3(key[110]), .A4(n862), 
        .A5(key_round[110]), .A6(n855), .Y(n46) );
  AO222X1_HVT U28 ( .A1(keyout[109]), .A2(n888), .A3(key[109]), .A4(n862), 
        .A5(key_round[109]), .A6(n855), .Y(n47) );
  AO222X1_HVT U29 ( .A1(keyout[108]), .A2(n888), .A3(key[108]), .A4(n862), 
        .A5(key_round[108]), .A6(n855), .Y(n48) );
  AO222X1_HVT U30 ( .A1(keyout[107]), .A2(n888), .A3(key[107]), .A4(n862), 
        .A5(key_round[107]), .A6(n855), .Y(n49) );
  AO222X1_HVT U31 ( .A1(keyout[106]), .A2(n888), .A3(key[106]), .A4(n862), 
        .A5(key_round[106]), .A6(n855), .Y(n50) );
  AO222X1_HVT U32 ( .A1(keyout[105]), .A2(n888), .A3(key[105]), .A4(n862), 
        .A5(key_round[105]), .A6(n855), .Y(n51) );
  AO222X1_HVT U33 ( .A1(keyout[104]), .A2(n888), .A3(key[104]), .A4(n862), 
        .A5(key_round[104]), .A6(n854), .Y(n52) );
  AO222X1_HVT U34 ( .A1(keyout[103]), .A2(n889), .A3(key[103]), .A4(n863), 
        .A5(key_round[103]), .A6(n854), .Y(n53) );
  AO222X1_HVT U35 ( .A1(keyout[102]), .A2(n889), .A3(key[102]), .A4(n863), 
        .A5(key_round[102]), .A6(n854), .Y(n54) );
  AO222X1_HVT U36 ( .A1(keyout[101]), .A2(n889), .A3(key[101]), .A4(n863), 
        .A5(key_round[101]), .A6(n854), .Y(n55) );
  AO222X1_HVT U37 ( .A1(keyout[100]), .A2(n889), .A3(key[100]), .A4(n863), 
        .A5(key_round[100]), .A6(n854), .Y(n56) );
  AO222X1_HVT U38 ( .A1(keyout[99]), .A2(n889), .A3(key[99]), .A4(n863), .A5(
        key_round[99]), .A6(n854), .Y(n57) );
  AO222X1_HVT U39 ( .A1(keyout[98]), .A2(n889), .A3(key[98]), .A4(n863), .A5(
        key_round[98]), .A6(n854), .Y(n58) );
  AO222X1_HVT U40 ( .A1(keyout[97]), .A2(n889), .A3(key[97]), .A4(n863), .A5(
        key_round[97]), .A6(n854), .Y(n59) );
  AO222X1_HVT U41 ( .A1(keyout[96]), .A2(n889), .A3(key[96]), .A4(n863), .A5(
        key_round[96]), .A6(n854), .Y(n60) );
  AO222X1_HVT U42 ( .A1(keyout[95]), .A2(n889), .A3(key[95]), .A4(n863), .A5(
        key_round[95]), .A6(n854), .Y(n61) );
  AO222X1_HVT U43 ( .A1(keyout[94]), .A2(n889), .A3(key[94]), .A4(n863), .A5(
        key_round[94]), .A6(n854), .Y(n62) );
  AO222X1_HVT U44 ( .A1(keyout[93]), .A2(n889), .A3(key[93]), .A4(n863), .A5(
        key_round[93]), .A6(n854), .Y(n63) );
  AO222X1_HVT U45 ( .A1(keyout[92]), .A2(n889), .A3(key[92]), .A4(n863), .A5(
        key_round[92]), .A6(n854), .Y(n64) );
  AO222X1_HVT U46 ( .A1(keyout[91]), .A2(n890), .A3(key[91]), .A4(n864), .A5(
        key_round[91]), .A6(n853), .Y(n65) );
  AO222X1_HVT U47 ( .A1(keyout[90]), .A2(n890), .A3(key[90]), .A4(n864), .A5(
        key_round[90]), .A6(n853), .Y(n66) );
  AO222X1_HVT U48 ( .A1(keyout[89]), .A2(n890), .A3(key[89]), .A4(n864), .A5(
        key_round[89]), .A6(n853), .Y(n67) );
  AO222X1_HVT U49 ( .A1(keyout[88]), .A2(n890), .A3(key[88]), .A4(n864), .A5(
        key_round[88]), .A6(n853), .Y(n68) );
  AO222X1_HVT U50 ( .A1(keyout[87]), .A2(n890), .A3(key[87]), .A4(n864), .A5(
        key_round[87]), .A6(n853), .Y(n69) );
  AO222X1_HVT U51 ( .A1(keyout[86]), .A2(n890), .A3(key[86]), .A4(n864), .A5(
        key_round[86]), .A6(n853), .Y(n70) );
  AO222X1_HVT U52 ( .A1(keyout[85]), .A2(n890), .A3(key[85]), .A4(n864), .A5(
        key_round[85]), .A6(n853), .Y(n71) );
  AO222X1_HVT U53 ( .A1(keyout[84]), .A2(n890), .A3(key[84]), .A4(n864), .A5(
        key_round[84]), .A6(n853), .Y(n72) );
  AO222X1_HVT U54 ( .A1(keyout[83]), .A2(n890), .A3(key[83]), .A4(n864), .A5(
        key_round[83]), .A6(n853), .Y(n73) );
  AO222X1_HVT U55 ( .A1(keyout[82]), .A2(n890), .A3(key[82]), .A4(n864), .A5(
        key_round[82]), .A6(n853), .Y(n74) );
  AO222X1_HVT U56 ( .A1(keyout[81]), .A2(n890), .A3(key[81]), .A4(n864), .A5(
        key_round[81]), .A6(n853), .Y(n75) );
  AO222X1_HVT U57 ( .A1(keyout[80]), .A2(n890), .A3(key[80]), .A4(n864), .A5(
        key_round[80]), .A6(n853), .Y(n76) );
  AO222X1_HVT U58 ( .A1(keyout[79]), .A2(n891), .A3(key[79]), .A4(n865), .A5(
        key_round[79]), .A6(n853), .Y(n77) );
  AO222X1_HVT U59 ( .A1(keyout[78]), .A2(n891), .A3(key[78]), .A4(n865), .A5(
        key_round[78]), .A6(n852), .Y(n78) );
  AO222X1_HVT U60 ( .A1(keyout[77]), .A2(n891), .A3(key[77]), .A4(n865), .A5(
        key_round[77]), .A6(n852), .Y(n79) );
  AO222X1_HVT U61 ( .A1(keyout[76]), .A2(n891), .A3(key[76]), .A4(n865), .A5(
        key_round[76]), .A6(n852), .Y(n80) );
  AO222X1_HVT U62 ( .A1(keyout[75]), .A2(n891), .A3(key[75]), .A4(n865), .A5(
        key_round[75]), .A6(n852), .Y(n81) );
  AO222X1_HVT U63 ( .A1(keyout[74]), .A2(n891), .A3(key[74]), .A4(n865), .A5(
        key_round[74]), .A6(n852), .Y(n82) );
  AO222X1_HVT U64 ( .A1(keyout[73]), .A2(n891), .A3(key[73]), .A4(n865), .A5(
        key_round[73]), .A6(n852), .Y(n83) );
  AO222X1_HVT U65 ( .A1(keyout[72]), .A2(n891), .A3(key[72]), .A4(n865), .A5(
        key_round[72]), .A6(n852), .Y(n84) );
  AO222X1_HVT U66 ( .A1(keyout[71]), .A2(n891), .A3(key[71]), .A4(n865), .A5(
        key_round[71]), .A6(n852), .Y(n85) );
  AO222X1_HVT U67 ( .A1(keyout[70]), .A2(n891), .A3(key[70]), .A4(n865), .A5(
        key_round[70]), .A6(n852), .Y(n86) );
  AO222X1_HVT U68 ( .A1(keyout[69]), .A2(n891), .A3(key[69]), .A4(n865), .A5(
        key_round[69]), .A6(n852), .Y(n87) );
  AO222X1_HVT U69 ( .A1(keyout[68]), .A2(n891), .A3(key[68]), .A4(n865), .A5(
        key_round[68]), .A6(n852), .Y(n88) );
  AO222X1_HVT U70 ( .A1(keyout[67]), .A2(n892), .A3(key[67]), .A4(n866), .A5(
        key_round[67]), .A6(n852), .Y(n89) );
  AO222X1_HVT U71 ( .A1(keyout[66]), .A2(n892), .A3(key[66]), .A4(n866), .A5(
        key_round[66]), .A6(n852), .Y(n90) );
  AO222X1_HVT U72 ( .A1(keyout[65]), .A2(n892), .A3(key[65]), .A4(n866), .A5(
        key_round[65]), .A6(n851), .Y(n91) );
  AO222X1_HVT U73 ( .A1(keyout[64]), .A2(n892), .A3(key[64]), .A4(n866), .A5(
        key_round[64]), .A6(n851), .Y(n92) );
  AO222X1_HVT U74 ( .A1(keyout[63]), .A2(n892), .A3(key[63]), .A4(n866), .A5(
        key_round[63]), .A6(n851), .Y(n93) );
  AO222X1_HVT U75 ( .A1(keyout[62]), .A2(n892), .A3(key[62]), .A4(n866), .A5(
        key_round[62]), .A6(n851), .Y(n94) );
  AO222X1_HVT U76 ( .A1(keyout[61]), .A2(n892), .A3(key[61]), .A4(n866), .A5(
        key_round[61]), .A6(n851), .Y(n95) );
  AO222X1_HVT U77 ( .A1(keyout[60]), .A2(n892), .A3(key[60]), .A4(n866), .A5(
        key_round[60]), .A6(n851), .Y(n96) );
  AO222X1_HVT U78 ( .A1(keyout[59]), .A2(n892), .A3(key[59]), .A4(n866), .A5(
        key_round[59]), .A6(n851), .Y(n97) );
  AO222X1_HVT U79 ( .A1(keyout[58]), .A2(n892), .A3(key[58]), .A4(n866), .A5(
        key_round[58]), .A6(n851), .Y(n98) );
  AO222X1_HVT U80 ( .A1(keyout[57]), .A2(n892), .A3(key[57]), .A4(n866), .A5(
        key_round[57]), .A6(n851), .Y(n99) );
  AO222X1_HVT U81 ( .A1(keyout[56]), .A2(n892), .A3(key[56]), .A4(n866), .A5(
        key_round[56]), .A6(n851), .Y(n100) );
  AO222X1_HVT U82 ( .A1(keyout[55]), .A2(n893), .A3(key[55]), .A4(n867), .A5(
        key_round[55]), .A6(n851), .Y(n101) );
  AO222X1_HVT U83 ( .A1(keyout[54]), .A2(n893), .A3(key[54]), .A4(n867), .A5(
        key_round[54]), .A6(n851), .Y(n102) );
  AO222X1_HVT U84 ( .A1(keyout[53]), .A2(n893), .A3(key[53]), .A4(n867), .A5(
        key_round[53]), .A6(n851), .Y(n103) );
  AO222X1_HVT U85 ( .A1(keyout[52]), .A2(n893), .A3(key[52]), .A4(n867), .A5(
        key_round[52]), .A6(n850), .Y(n104) );
  AO222X1_HVT U86 ( .A1(keyout[51]), .A2(n893), .A3(key[51]), .A4(n867), .A5(
        key_round[51]), .A6(n850), .Y(n105) );
  AO222X1_HVT U87 ( .A1(keyout[50]), .A2(n893), .A3(key[50]), .A4(n867), .A5(
        key_round[50]), .A6(n850), .Y(n106) );
  AO222X1_HVT U88 ( .A1(keyout[49]), .A2(n893), .A3(key[49]), .A4(n867), .A5(
        key_round[49]), .A6(n850), .Y(n107) );
  AO222X1_HVT U89 ( .A1(keyout[48]), .A2(n893), .A3(key[48]), .A4(n867), .A5(
        key_round[48]), .A6(n850), .Y(n108) );
  AO222X1_HVT U90 ( .A1(keyout[47]), .A2(n893), .A3(key[47]), .A4(n867), .A5(
        key_round[47]), .A6(n850), .Y(n109) );
  AO222X1_HVT U91 ( .A1(keyout[46]), .A2(n893), .A3(key[46]), .A4(n867), .A5(
        key_round[46]), .A6(n850), .Y(n110) );
  AO222X1_HVT U92 ( .A1(keyout[45]), .A2(n893), .A3(key[45]), .A4(n867), .A5(
        key_round[45]), .A6(n850), .Y(n111) );
  AO222X1_HVT U93 ( .A1(keyout[44]), .A2(n893), .A3(key[44]), .A4(n867), .A5(
        key_round[44]), .A6(n850), .Y(n112) );
  AO222X1_HVT U94 ( .A1(keyout[43]), .A2(n894), .A3(key[43]), .A4(n868), .A5(
        key_round[43]), .A6(n850), .Y(n113) );
  AO222X1_HVT U95 ( .A1(keyout[42]), .A2(n894), .A3(key[42]), .A4(n868), .A5(
        key_round[42]), .A6(n850), .Y(n114) );
  AO222X1_HVT U96 ( .A1(keyout[41]), .A2(n894), .A3(key[41]), .A4(n868), .A5(
        key_round[41]), .A6(n850), .Y(n115) );
  AO222X1_HVT U97 ( .A1(keyout[40]), .A2(n894), .A3(key[40]), .A4(n868), .A5(
        key_round[40]), .A6(n850), .Y(n116) );
  AO222X1_HVT U98 ( .A1(keyout[39]), .A2(n894), .A3(key[39]), .A4(n868), .A5(
        key_round[39]), .A6(n849), .Y(n117) );
  AO222X1_HVT U99 ( .A1(keyout[38]), .A2(n894), .A3(key[38]), .A4(n868), .A5(
        key_round[38]), .A6(n849), .Y(n118) );
  AO222X1_HVT U100 ( .A1(keyout[37]), .A2(n894), .A3(key[37]), .A4(n868), .A5(
        key_round[37]), .A6(n849), .Y(n119) );
  AO222X1_HVT U101 ( .A1(keyout[36]), .A2(n894), .A3(key[36]), .A4(n868), .A5(
        key_round[36]), .A6(n849), .Y(n120) );
  AO222X1_HVT U102 ( .A1(keyout[35]), .A2(n894), .A3(key[35]), .A4(n868), .A5(
        key_round[35]), .A6(n849), .Y(n121) );
  AO222X1_HVT U103 ( .A1(keyout[34]), .A2(n894), .A3(key[34]), .A4(n868), .A5(
        key_round[34]), .A6(n849), .Y(n122) );
  AO222X1_HVT U104 ( .A1(keyout[33]), .A2(n894), .A3(key[33]), .A4(n868), .A5(
        key_round[33]), .A6(n849), .Y(n123) );
  AO222X1_HVT U105 ( .A1(keyout[32]), .A2(n894), .A3(key[32]), .A4(n868), .A5(
        key_round[32]), .A6(n849), .Y(n124) );
  AO222X1_HVT U106 ( .A1(keyout[31]), .A2(n895), .A3(key[31]), .A4(n869), .A5(
        key_round[31]), .A6(n849), .Y(n125) );
  AO222X1_HVT U107 ( .A1(keyout[30]), .A2(n895), .A3(key[30]), .A4(n869), .A5(
        key_round[30]), .A6(n849), .Y(n126) );
  AO222X1_HVT U108 ( .A1(keyout[29]), .A2(n895), .A3(key[29]), .A4(n869), .A5(
        key_round[29]), .A6(n849), .Y(n127) );
  AO222X1_HVT U109 ( .A1(keyout[28]), .A2(n895), .A3(key[28]), .A4(n869), .A5(
        key_round[28]), .A6(n849), .Y(n128) );
  AO222X1_HVT U110 ( .A1(keyout[27]), .A2(n895), .A3(key[27]), .A4(n869), .A5(
        key_round[27]), .A6(n849), .Y(n129) );
  AO222X1_HVT U111 ( .A1(keyout[26]), .A2(n895), .A3(key[26]), .A4(n869), .A5(
        key_round[26]), .A6(n848), .Y(n130) );
  AO222X1_HVT U112 ( .A1(keyout[25]), .A2(n895), .A3(key[25]), .A4(n869), .A5(
        key_round[25]), .A6(n848), .Y(n131) );
  AO222X1_HVT U113 ( .A1(keyout[24]), .A2(n895), .A3(key[24]), .A4(n869), .A5(
        key_round[24]), .A6(n848), .Y(n132) );
  AO222X1_HVT U114 ( .A1(keyout[23]), .A2(n895), .A3(key[23]), .A4(n869), .A5(
        key_round[23]), .A6(n848), .Y(n133) );
  AO222X1_HVT U115 ( .A1(keyout[22]), .A2(n895), .A3(key[22]), .A4(n869), .A5(
        key_round[22]), .A6(n848), .Y(n134) );
  AO222X1_HVT U116 ( .A1(keyout[21]), .A2(n895), .A3(key[21]), .A4(n869), .A5(
        key_round[21]), .A6(n848), .Y(n135) );
  AO222X1_HVT U117 ( .A1(keyout[20]), .A2(n895), .A3(key[20]), .A4(n869), .A5(
        key_round[20]), .A6(n848), .Y(n136) );
  AO222X1_HVT U118 ( .A1(keyout[19]), .A2(n896), .A3(key[19]), .A4(n870), .A5(
        key_round[19]), .A6(n848), .Y(n137) );
  AO222X1_HVT U119 ( .A1(keyout[18]), .A2(n896), .A3(key[18]), .A4(n870), .A5(
        key_round[18]), .A6(n848), .Y(n138) );
  AO222X1_HVT U120 ( .A1(keyout[17]), .A2(n896), .A3(key[17]), .A4(n870), .A5(
        key_round[17]), .A6(n848), .Y(n139) );
  AO222X1_HVT U121 ( .A1(keyout[16]), .A2(n896), .A3(key[16]), .A4(n870), .A5(
        key_round[16]), .A6(n848), .Y(n140) );
  AO222X1_HVT U122 ( .A1(keyout[15]), .A2(n896), .A3(key[15]), .A4(n870), .A5(
        key_round[15]), .A6(n848), .Y(n141) );
  AO222X1_HVT U123 ( .A1(keyout[14]), .A2(n896), .A3(key[14]), .A4(n870), .A5(
        key_round[14]), .A6(n848), .Y(n142) );
  AO222X1_HVT U124 ( .A1(keyout[13]), .A2(n896), .A3(key[13]), .A4(n870), .A5(
        key_round[13]), .A6(n847), .Y(n143) );
  AO222X1_HVT U125 ( .A1(keyout[12]), .A2(n896), .A3(key[12]), .A4(n870), .A5(
        key_round[12]), .A6(n847), .Y(n144) );
  AO222X1_HVT U126 ( .A1(n896), .A2(keyout[11]), .A3(key[11]), .A4(n870), .A5(
        key_round[11]), .A6(n847), .Y(n145) );
  AO222X1_HVT U127 ( .A1(keyout[10]), .A2(n896), .A3(key[10]), .A4(n870), .A5(
        key_round[10]), .A6(n847), .Y(n146) );
  AO222X1_HVT U128 ( .A1(keyout[9]), .A2(n896), .A3(key[9]), .A4(n870), .A5(
        key_round[9]), .A6(n847), .Y(n147) );
  AO222X1_HVT U129 ( .A1(keyout[8]), .A2(n896), .A3(key[8]), .A4(n870), .A5(
        key_round[8]), .A6(n847), .Y(n148) );
  AO222X1_HVT U130 ( .A1(keyout[7]), .A2(n897), .A3(key[7]), .A4(n871), .A5(
        key_round[7]), .A6(n847), .Y(n149) );
  AO222X1_HVT U131 ( .A1(keyout[6]), .A2(n897), .A3(key[6]), .A4(n871), .A5(
        key_round[6]), .A6(n847), .Y(n150) );
  AO222X1_HVT U132 ( .A1(keyout[5]), .A2(n897), .A3(key[5]), .A4(n871), .A5(
        key_round[5]), .A6(n847), .Y(n151) );
  AO222X1_HVT U133 ( .A1(keyout[4]), .A2(n897), .A3(key[4]), .A4(n871), .A5(
        key_round[4]), .A6(n847), .Y(n152) );
  AO222X1_HVT U134 ( .A1(keyout[3]), .A2(n897), .A3(key[3]), .A4(n871), .A5(
        key_round[3]), .A6(n847), .Y(n153) );
  AO222X1_HVT U135 ( .A1(keyout[2]), .A2(n897), .A3(key[2]), .A4(n871), .A5(
        key_round[2]), .A6(n847), .Y(n154) );
  AO222X1_HVT U136 ( .A1(keyout[1]), .A2(n897), .A3(key[1]), .A4(n871), .A5(
        key_round[1]), .A6(n847), .Y(n155) );
  AO222X1_HVT U137 ( .A1(keyout[0]), .A2(n897), .A3(key[0]), .A4(n871), .A5(
        key_round[0]), .A6(n846), .Y(n156) );
  AO222X1_HVT U139 ( .A1(n897), .A2(n917), .A3(adk_out0[126]), .A4(n871), .A5(
        adk_in[126]), .A6(n846), .Y(n158) );
  AO222X1_HVT U143 ( .A1(n921), .A2(n898), .A3(adk_out0[122]), .A4(n872), .A5(
        adk_in[122]), .A6(n846), .Y(n162) );
  AO222X1_HVT U145 ( .A1(n923), .A2(n898), .A3(adk_out0[120]), .A4(n872), .A5(
        adk_in[120]), .A6(n846), .Y(n164) );
  AO222X1_HVT U146 ( .A1(n924), .A2(n898), .A3(adk_out0[119]), .A4(n872), .A5(
        adk_in[119]), .A6(n846), .Y(n165) );
  AO222X1_HVT U147 ( .A1(n898), .A2(n925), .A3(adk_out0[118]), .A4(n872), .A5(
        adk_in[118]), .A6(n846), .Y(n166) );
  AO222X1_HVT U151 ( .A1(n929), .A2(n898), .A3(adk_out0[114]), .A4(n872), .A5(
        adk_in[114]), .A6(n845), .Y(n170) );
  AO222X1_HVT U153 ( .A1(n931), .A2(n898), .A3(adk_out0[112]), .A4(n872), .A5(
        adk_in[112]), .A6(n845), .Y(n172) );
  AO222X1_HVT U155 ( .A1(n899), .A2(n933), .A3(adk_out0[110]), .A4(n873), .A5(
        adk_in[110]), .A6(n845), .Y(n174) );
  AO222X1_HVT U156 ( .A1(n899), .A2(n934), .A3(adk_out0[109]), .A4(n873), .A5(
        adk_in[109]), .A6(n845), .Y(n175) );
  AO222X1_HVT U157 ( .A1(n899), .A2(n935), .A3(adk_out0[108]), .A4(n873), .A5(
        adk_in[108]), .A6(n845), .Y(n176) );
  AO222X1_HVT U160 ( .A1(n899), .A2(n938), .A3(adk_out0[105]), .A4(n873), .A5(
        adk_in[105]), .A6(n845), .Y(n179) );
  AO222X1_HVT U161 ( .A1(n899), .A2(n939), .A3(adk_out0[104]), .A4(n873), .A5(
        adk_in[104]), .A6(n845), .Y(n180) );
  AO222X1_HVT U163 ( .A1(n940), .A2(n899), .A3(adk_out0[102]), .A4(n873), .A5(
        adk_in[102]), .A6(n844), .Y(n182) );
  AO222X1_HVT U164 ( .A1(n941), .A2(n899), .A3(adk_out0[101]), .A4(n873), .A5(
        adk_in[101]), .A6(n844), .Y(n183) );
  AO222X1_HVT U167 ( .A1(n944), .A2(n900), .A3(adk_out0[98]), .A4(n874), .A5(
        adk_in[98]), .A6(n844), .Y(n186) );
  AO222X1_HVT U168 ( .A1(n900), .A2(n945), .A3(adk_out0[97]), .A4(n874), .A5(
        adk_in[97]), .A6(n844), .Y(n187) );
  AO222X1_HVT U169 ( .A1(n900), .A2(n946), .A3(adk_out0[96]), .A4(n874), .A5(
        adk_in[96]), .A6(n844), .Y(n188) );
  AO222X1_HVT U170 ( .A1(n900), .A2(n947), .A3(adk_out0[95]), .A4(n874), .A5(
        adk_in[95]), .A6(n844), .Y(n189) );
  AO222X1_HVT U175 ( .A1(n900), .A2(n952), .A3(adk_out0[90]), .A4(n874), .A5(
        adk_in[90]), .A6(n844), .Y(n194) );
  AO222X1_HVT U177 ( .A1(n900), .A2(n954), .A3(adk_out0[88]), .A4(n874), .A5(
        adk_in[88]), .A6(n843), .Y(n196) );
  AO222X1_HVT U179 ( .A1(n901), .A2(n956), .A3(adk_out0[86]), .A4(n875), .A5(
        adk_in[86]), .A6(n843), .Y(n198) );
  AO222X1_HVT U180 ( .A1(n901), .A2(n957), .A3(adk_out0[85]), .A4(n875), .A5(
        adk_in[85]), .A6(n843), .Y(n199) );
  AO222X1_HVT U186 ( .A1(n901), .A2(n963), .A3(adk_out0[79]), .A4(n875), .A5(
        adk_in[79]), .A6(n843), .Y(n205) );
  AO222X1_HVT U187 ( .A1(n964), .A2(n901), .A3(adk_out0[78]), .A4(n875), .A5(
        adk_in[78]), .A6(n843), .Y(n206) );
  AO222X1_HVT U191 ( .A1(n902), .A2(n968), .A3(adk_out0[74]), .A4(n876), .A5(
        adk_in[74]), .A6(n842), .Y(n210) );
  AO222X1_HVT U192 ( .A1(n902), .A2(n969), .A3(adk_out0[73]), .A4(n876), .A5(
        adk_in[73]), .A6(n842), .Y(n211) );
  AO222X1_HVT U193 ( .A1(n902), .A2(n970), .A3(adk_out0[72]), .A4(n876), .A5(
        adk_in[72]), .A6(n842), .Y(n212) );
  AO222X1_HVT U194 ( .A1(n902), .A2(n971), .A3(adk_out0[71]), .A4(n876), .A5(
        adk_in[71]), .A6(n842), .Y(n213) );
  AO222X1_HVT U195 ( .A1(n972), .A2(n902), .A3(adk_out0[70]), .A4(n876), .A5(
        adk_in[70]), .A6(n842), .Y(n214) );
  AO222X1_HVT U199 ( .A1(n976), .A2(n902), .A3(adk_out0[66]), .A4(n876), .A5(
        adk_in[66]), .A6(n842), .Y(n218) );
  AO222X1_HVT U201 ( .A1(n902), .A2(n978), .A3(adk_out0[64]), .A4(n876), .A5(
        adk_in[64]), .A6(n842), .Y(n220) );
  AO222X1_HVT U215 ( .A1(n904), .A2(n992), .A3(adk_out0[50]), .A4(n878), .A5(
        adk_in[50]), .A6(n840), .Y(n234) );
  AO222X1_HVT U216 ( .A1(n904), .A2(n993), .A3(adk_out0[49]), .A4(n878), .A5(
        adk_in[49]), .A6(n840), .Y(n235) );
  AO222X1_HVT U217 ( .A1(n994), .A2(n904), .A3(adk_out0[48]), .A4(n878), .A5(
        adk_in[48]), .A6(n840), .Y(n236) );
  AO222X1_HVT U225 ( .A1(n904), .A2(n1002), .A3(adk_out0[40]), .A4(n878), .A5(
        adk_in[40]), .A6(n840), .Y(n244) );
  AO222X1_HVT U228 ( .A1(n1005), .A2(n905), .A3(adk_out0[37]), .A4(n879), .A5(
        adk_in[37]), .A6(n839), .Y(n247) );
  AO222X1_HVT U233 ( .A1(n905), .A2(n1010), .A3(adk_out0[32]), .A4(n879), .A5(
        adk_in[32]), .A6(n839), .Y(n252) );
  AO222X1_HVT U234 ( .A1(n905), .A2(n1011), .A3(adk_out0[31]), .A4(n879), .A5(
        adk_in[31]), .A6(n839), .Y(n253) );
  AO222X1_HVT U239 ( .A1(n906), .A2(n1016), .A3(adk_out0[26]), .A4(n880), .A5(
        adk_in[26]), .A6(n839), .Y(n258) );
  AO222X1_HVT U244 ( .A1(n1021), .A2(n906), .A3(adk_out0[21]), .A4(n880), .A5(
        adk_in[21]), .A6(n838), .Y(n263) );
  AO222X1_HVT U247 ( .A1(n906), .A2(n1024), .A3(adk_out0[18]), .A4(n880), .A5(
        adk_in[18]), .A6(n838), .Y(n266) );
  AO222X1_HVT U248 ( .A1(n1025), .A2(n906), .A3(adk_out0[17]), .A4(n880), .A5(
        adk_in[17]), .A6(n838), .Y(n267) );
  AO222X1_HVT U251 ( .A1(n907), .A2(n1028), .A3(adk_out0[14]), .A4(n881), .A5(
        adk_in[14]), .A6(n838), .Y(n270) );
  AO222X1_HVT U257 ( .A1(n1034), .A2(n907), .A3(adk_out0[8]), .A4(n881), .A5(
        adk_in[8]), .A6(n837), .Y(n276) );
  AO222X1_HVT U258 ( .A1(n907), .A2(n1035), .A3(adk_out0[7]), .A4(n881), .A5(
        adk_in[7]), .A6(n837), .Y(n277) );
  AO222X1_HVT U259 ( .A1(n1036), .A2(n907), .A3(adk_out0[6]), .A4(n881), .A5(
        adk_in[6]), .A6(n837), .Y(n278) );
  AO222X1_HVT U260 ( .A1(n1037), .A2(n907), .A3(adk_out0[5]), .A4(n881), .A5(
        adk_in[5]), .A6(n837), .Y(n279) );
  AO222X1_HVT U265 ( .A1(n908), .A2(n1042), .A3(adk_out0[0]), .A4(n882), .A5(
        adk_in[0]), .A6(n837), .Y(n284) );
  NOR2X0_HVT U267 ( .A1(n837), .A2(n18), .Y(n15) );
  AO22X1_HVT U268 ( .A1(round_number[2]), .A2(n19), .A3(n20), .A4(n21), .Y(
        n285) );
  AND2X1_HVT U269 ( .A1(round_number[1]), .A2(n6), .Y(n20) );
  AO22X1_HVT U270 ( .A1(round_number[1]), .A2(n22), .A3(n21), .A4(n7), .Y(n286) );
  AO22X1_HVT U271 ( .A1(n23), .A2(round_number[0]), .A3(n859), .A4(n8), .Y(
        n287) );
  AO22X1_HVT U272 ( .A1(round_number[3]), .A2(n19), .A3(n24), .A4(
        round_number[2]), .Y(n288) );
  AND2X1_HVT U273 ( .A1(n21), .A2(round_number[1]), .Y(n24) );
  AND2X1_HVT U274 ( .A1(round_number[0]), .A2(n858), .Y(n21) );
  AO21X1_HVT U275 ( .A1(n860), .A2(n7), .A3(n22), .Y(n19) );
  AO21X1_HVT U276 ( .A1(n860), .A2(n8), .A3(n23), .Y(n22) );
  AOI21X1_HVT U277 ( .A1(start), .A2(n914), .A3(n860), .Y(n23) );
  OR2X1_HVT U278 ( .A1(n25), .A2(reset), .Y(n17) );
  NAND2X0_HVT U279 ( .A1(n26), .A2(n13), .Y(n289) );
  AND2X1_HVT U280 ( .A1(n915), .A2(n12), .Y(n13) );
  NAND4X0_HVT U281 ( .A1(n8), .A2(n6), .A3(n9), .A4(n27), .Y(n12) );
  AND2X1_HVT U282 ( .A1(round_number[3]), .A2(round_number[1]), .Y(n27) );
  AO21X1_HVT U283 ( .A1(start), .A2(n914), .A3(n9), .Y(n26) );
  NAND3X0_HVT U284 ( .A1(n25), .A2(n915), .A3(d), .Y(n14) );
  OA21X1_HVT U285 ( .A1(round_number[1]), .A2(round_number[2]), .A3(
        round_number[3]), .Y(n25) );
  add_round_keys_0 adk_0 ( .state(plaintext), .subkey(key), .out(adk_out0) );
  round r1 ( .in({adk_in[127:123], n739, n519, adk_in[120:114], n371, 
        adk_in[112], n526, adk_in[110:98], n449, adk_in[96:90], n462, 
        adk_in[88:85], n366, n343, adk_in[82], n484, adk_in[80:77], n491, 
        adk_in[75:67], n352, adk_in[65:64], n650, adk_in[62:53], n636, 
        adk_in[51:50], n310, adk_in[48:40], n624, adk_in[38:34], n382, 
        adk_in[32:21], n612, adk_in[19:13], n408, adk_in[11], n704, 
        adk_in[9:5], n538, adk_in[3:2], n469, adk_in[0]}), .round_num(
        round_number), .keyin({key_round[127:19], n388, key_round[17:16], n551, 
        key_round[14:11], n689, key_round[9:8], n364, key_round[6:3], n654, 
        n369, key_round[0]}), .keyout(keyout), .out({n916, n917, n918, n919, 
        n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
        n932, n933, n934, n935, n936, n937, n938, n939, cipher_text[103], n940, 
        n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
        n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
        n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
        n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
        n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
        n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
        n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
        n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
        n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
        n1040, n1041, n1042}) );
  DFFX1_HVT \adk_in_reg[110]  ( .D(n174), .CLK(clk), .Q(adk_in[110]) );
  DFFX2_HVT \adk_in_reg[77]  ( .D(n207), .CLK(clk), .Q(adk_in[77]) );
  AO222X1_HVT U4 ( .A1(n1), .A2(n916), .A3(adk_out0[127]), .A4(n886), .A5(n2), 
        .A6(n3), .Y(n157) );
  IBUFFX16_HVT U5 ( .A(n910), .Y(n1) );
  IBUFFX16_HVT U6 ( .A(n367), .Y(n2) );
  IBUFFX16_HVT U7 ( .A(n858), .Y(n3) );
  INVX0_HVT U138 ( .A(n916), .Y(n718) );
  NAND2X0_HVT U140 ( .A1(n937), .A2(n899), .Y(n4) );
  NAND2X0_HVT U141 ( .A1(adk_out0[106]), .A2(n873), .Y(n5) );
  NAND2X0_HVT U142 ( .A1(adk_in[106]), .A2(n845), .Y(n10) );
  NAND3X0_HVT U144 ( .A1(n4), .A2(n5), .A3(n10), .Y(n178) );
  INVX1_HVT U148 ( .A(n666), .Y(cipher_text[1]) );
  INVX1_HVT U149 ( .A(n699), .Y(cipher_text[42]) );
  INVX1_HVT U150 ( .A(n1000), .Y(n699) );
  NBUFFX16_HVT U152 ( .A(n984), .Y(cipher_text[58]) );
  INVX1_HVT U154 ( .A(n1041), .Y(n666) );
  INVX0_HVT U158 ( .A(n931), .Y(n16) );
  INVX0_HVT U159 ( .A(n16), .Y(cipher_text[112]) );
  INVX2_HVT U162 ( .A(n688), .Y(n689) );
  INVX1_HVT U165 ( .A(n600), .Y(cipher_text[56]) );
  INVX0_HVT U166 ( .A(n772), .Y(n291) );
  INVX1_HVT U171 ( .A(n999), .Y(n772) );
  NAND2X0_HVT U172 ( .A1(n1019), .A2(n906), .Y(n292) );
  NAND2X0_HVT U173 ( .A1(adk_out0[23]), .A2(n880), .Y(n293) );
  NAND2X0_HVT U174 ( .A1(adk_in[23]), .A2(n838), .Y(n294) );
  NAND3X0_HVT U176 ( .A1(n292), .A2(n293), .A3(n294), .Y(n261) );
  NAND2X0_HVT U178 ( .A1(n984), .A2(n903), .Y(n295) );
  NAND2X0_HVT U181 ( .A1(adk_out0[58]), .A2(n877), .Y(n296) );
  NAND2X0_HVT U182 ( .A1(adk_in[58]), .A2(n841), .Y(n297) );
  NAND3X0_HVT U183 ( .A1(n295), .A2(n296), .A3(n297), .Y(n226) );
  INVX1_HVT U184 ( .A(n643), .Y(cipher_text[9]) );
  INVX4_HVT U185 ( .A(n351), .Y(n352) );
  INVX1_HVT U188 ( .A(n488), .Y(cipher_text[100]) );
  INVX1_HVT U189 ( .A(n926), .Y(n657) );
  NAND2X0_HVT U190 ( .A1(n927), .A2(n898), .Y(n298) );
  NAND2X0_HVT U196 ( .A1(adk_out0[116]), .A2(n872), .Y(n299) );
  NAND2X0_HVT U197 ( .A1(adk_in[116]), .A2(n846), .Y(n300) );
  NAND3X0_HVT U198 ( .A1(n298), .A2(n299), .A3(n300), .Y(n168) );
  INVX1_HVT U200 ( .A(n986), .Y(n600) );
  INVX1_HVT U202 ( .A(n942), .Y(n488) );
  NAND2X0_HVT U203 ( .A1(n904), .A2(n996), .Y(n301) );
  NAND2X0_HVT U204 ( .A1(adk_out0[46]), .A2(n878), .Y(n302) );
  NAND2X0_HVT U205 ( .A1(adk_in[46]), .A2(n840), .Y(n303) );
  NAND3X0_HVT U206 ( .A1(n301), .A2(n302), .A3(n303), .Y(n238) );
  INVX0_HVT U207 ( .A(n1038), .Y(n808) );
  INVX0_HVT U208 ( .A(n647), .Y(cipher_text[76]) );
  INVX0_HVT U209 ( .A(n966), .Y(n647) );
  NAND2X0_HVT U210 ( .A1(n899), .A2(n942), .Y(n304) );
  NAND2X0_HVT U211 ( .A1(adk_out0[100]), .A2(n873), .Y(n305) );
  NAND2X0_HVT U212 ( .A1(adk_in[100]), .A2(n844), .Y(n306) );
  NAND3X0_HVT U213 ( .A1(n304), .A2(n305), .A3(n306), .Y(n184) );
  INVX0_HVT U214 ( .A(n997), .Y(n523) );
  INVX1_HVT U218 ( .A(n523), .Y(cipher_text[45]) );
  INVX1_HVT U219 ( .A(n943), .Y(n307) );
  INVX1_HVT U220 ( .A(n307), .Y(cipher_text[99]) );
  INVX1_HVT U221 ( .A(n309), .Y(n310) );
  INVX0_HVT U222 ( .A(n810), .Y(n311) );
  INVX1_HVT U223 ( .A(n983), .Y(n810) );
  INVX0_HVT U224 ( .A(n1014), .Y(n729) );
  INVX1_HVT U226 ( .A(n623), .Y(n624) );
  NBUFFX4_HVT U227 ( .A(n1013), .Y(cipher_text[29]) );
  NAND2X0_HVT U229 ( .A1(n571), .A2(n570), .Y(n312) );
  NAND2X0_HVT U230 ( .A1(n313), .A2(n569), .Y(n181) );
  INVX0_HVT U231 ( .A(n312), .Y(n313) );
  NAND2X0_HVT U232 ( .A1(n926), .A2(n898), .Y(n314) );
  NAND2X0_HVT U235 ( .A1(adk_out0[117]), .A2(n872), .Y(n315) );
  NAND2X0_HVT U236 ( .A1(adk_in[117]), .A2(n846), .Y(n316) );
  NAND3X0_HVT U237 ( .A1(n314), .A2(n315), .A3(n316), .Y(n167) );
  INVX1_HVT U238 ( .A(n606), .Y(cipher_text[81]) );
  NAND2X0_HVT U240 ( .A1(n1029), .A2(n907), .Y(n317) );
  NAND2X0_HVT U241 ( .A1(adk_out0[13]), .A2(n881), .Y(n318) );
  NAND2X0_HVT U242 ( .A1(adk_in[13]), .A2(n838), .Y(n319) );
  NAND3X0_HVT U243 ( .A1(n317), .A2(n318), .A3(n319), .Y(n271) );
  INVX1_HVT U245 ( .A(n505), .Y(cipher_text[25]) );
  NAND2X0_HVT U246 ( .A1(n902), .A2(n973), .Y(n320) );
  NAND2X0_HVT U249 ( .A1(adk_out0[69]), .A2(n876), .Y(n321) );
  NAND2X0_HVT U250 ( .A1(adk_in[69]), .A2(n842), .Y(n322) );
  NAND3X0_HVT U252 ( .A1(n320), .A2(n321), .A3(n322), .Y(n215) );
  INVX0_HVT U253 ( .A(n1023), .Y(n812) );
  INVX0_HVT U254 ( .A(n742), .Y(n323) );
  INVX1_HVT U255 ( .A(n967), .Y(n742) );
  INVX0_HVT U256 ( .A(n953), .Y(n701) );
  INVX0_HVT U261 ( .A(n989), .Y(n602) );
  NAND2X0_HVT U262 ( .A1(n1032), .A2(n907), .Y(n324) );
  NAND2X0_HVT U263 ( .A1(adk_out0[10]), .A2(n881), .Y(n325) );
  NAND2X0_HVT U264 ( .A1(adk_in[10]), .A2(n837), .Y(n326) );
  NAND3X0_HVT U266 ( .A1(n324), .A2(n325), .A3(n326), .Y(n274) );
  INVX0_HVT U286 ( .A(n1031), .Y(n481) );
  NAND2X0_HVT U287 ( .A1(n1000), .A2(n904), .Y(n327) );
  NAND2X0_HVT U288 ( .A1(adk_out0[42]), .A2(n878), .Y(n328) );
  NAND2X0_HVT U289 ( .A1(adk_in[42]), .A2(n840), .Y(n329) );
  NAND3X0_HVT U290 ( .A1(n327), .A2(n328), .A3(n329), .Y(n242) );
  INVX1_HVT U291 ( .A(n808), .Y(cipher_text[4]) );
  INVX1_HVT U292 ( .A(n533), .Y(cipher_text[39]) );
  INVX1_HVT U293 ( .A(n574), .Y(cipher_text[15]) );
  INVX1_HVT U294 ( .A(n1027), .Y(n574) );
  NAND2X0_HVT U295 ( .A1(n1033), .A2(n907), .Y(n330) );
  NAND2X0_HVT U296 ( .A1(adk_out0[9]), .A2(n881), .Y(n331) );
  NAND2X0_HVT U297 ( .A1(adk_in[9]), .A2(n837), .Y(n332) );
  NAND3X0_HVT U298 ( .A1(n330), .A2(n331), .A3(n332), .Y(n275) );
  NAND2X0_HVT U299 ( .A1(n1041), .A2(n908), .Y(n333) );
  NAND2X0_HVT U300 ( .A1(adk_out0[1]), .A2(n882), .Y(n334) );
  NAND2X0_HVT U301 ( .A1(adk_in[1]), .A2(n837), .Y(n335) );
  NAND3X0_HVT U302 ( .A1(n333), .A2(n334), .A3(n335), .Y(n283) );
  INVX2_HVT U303 ( .A(n635), .Y(n636) );
  INVX0_HVT U304 ( .A(n647), .Y(n336) );
  INVX0_HVT U305 ( .A(n572), .Y(n337) );
  INVX1_HVT U306 ( .A(n988), .Y(n572) );
  INVX0_HVT U307 ( .A(n548), .Y(cipher_text[57]) );
  INVX0_HVT U308 ( .A(n1022), .Y(n799) );
  INVX0_HVT U309 ( .A(n533), .Y(n338) );
  INVX1_HVT U310 ( .A(n1003), .Y(n533) );
  NAND2X0_HVT U311 ( .A1(n1027), .A2(n907), .Y(n339) );
  NAND2X0_HVT U312 ( .A1(adk_out0[15]), .A2(n881), .Y(n340) );
  NAND2X0_HVT U313 ( .A1(adk_in[15]), .A2(n838), .Y(n341) );
  NAND3X0_HVT U314 ( .A1(n339), .A2(n340), .A3(n341), .Y(n269) );
  INVX2_HVT U315 ( .A(n649), .Y(n650) );
  INVX0_HVT U316 ( .A(n1008), .Y(n686) );
  INVX1_HVT U317 ( .A(n342), .Y(n343) );
  INVX1_HVT U318 ( .A(n818), .Y(cipher_text[124]) );
  INVX1_HVT U319 ( .A(n919), .Y(n818) );
  INVX0_HVT U320 ( .A(n548), .Y(n344) );
  NAND2X0_HVT U321 ( .A1(n903), .A2(n337), .Y(n345) );
  NAND2X0_HVT U322 ( .A1(adk_out0[54]), .A2(n877), .Y(n346) );
  NAND2X0_HVT U323 ( .A1(adk_in[54]), .A2(n841), .Y(n347) );
  NAND3X0_HVT U324 ( .A1(n345), .A2(n346), .A3(n347), .Y(n230) );
  INVX0_HVT U325 ( .A(n1030), .Y(n754) );
  INVX1_HVT U326 ( .A(n1017), .Y(n505) );
  NAND2X0_HVT U327 ( .A1(n902), .A2(n977), .Y(n348) );
  NAND2X0_HVT U328 ( .A1(adk_out0[65]), .A2(n876), .Y(n349) );
  NAND2X0_HVT U329 ( .A1(adk_in[65]), .A2(n842), .Y(n350) );
  NAND3X0_HVT U330 ( .A1(n348), .A2(n349), .A3(n350), .Y(n219) );
  INVX1_HVT U331 ( .A(n766), .Y(cipher_text[36]) );
  INVX0_HVT U332 ( .A(n923), .Y(n353) );
  INVX0_HVT U333 ( .A(n353), .Y(cipher_text[120]) );
  INVX1_HVT U334 ( .A(n602), .Y(cipher_text[53]) );
  INVX1_HVT U335 ( .A(n982), .Y(n797) );
  NAND2X0_HVT U336 ( .A1(n1026), .A2(n906), .Y(n355) );
  NAND2X0_HVT U337 ( .A1(adk_out0[16]), .A2(n880), .Y(n356) );
  NAND2X0_HVT U338 ( .A1(adk_in[16]), .A2(n838), .Y(n357) );
  NAND3X0_HVT U339 ( .A1(n355), .A2(n356), .A3(n357), .Y(n268) );
  INVX1_HVT U340 ( .A(n1026), .Y(n724) );
  NAND2X0_HVT U341 ( .A1(n906), .A2(n1017), .Y(n358) );
  NAND2X0_HVT U342 ( .A1(adk_out0[25]), .A2(n880), .Y(n359) );
  NAND2X0_HVT U343 ( .A1(adk_in[25]), .A2(n839), .Y(n360) );
  NAND3X0_HVT U344 ( .A1(n358), .A2(n359), .A3(n360), .Y(n259) );
  INVX1_HVT U345 ( .A(n490), .Y(n491) );
  INVX0_HVT U346 ( .A(n1001), .Y(n668) );
  INVX1_HVT U347 ( .A(n361), .Y(n362) );
  INVX1_HVT U348 ( .A(n363), .Y(n364) );
  INVX1_HVT U349 ( .A(n365), .Y(n366) );
  INVX1_HVT U350 ( .A(n387), .Y(n388) );
  INVX1_HVT U351 ( .A(n368), .Y(n369) );
  INVX1_HVT U352 ( .A(n370), .Y(n371) );
  NBUFFX2_HVT U353 ( .A(n1018), .Y(cipher_text[24]) );
  NBUFFX4_HVT U354 ( .A(n949), .Y(cipher_text[93]) );
  NAND2X0_HVT U355 ( .A1(n980), .A2(n903), .Y(n372) );
  NAND2X0_HVT U356 ( .A1(adk_out0[62]), .A2(n877), .Y(n373) );
  NAND2X0_HVT U357 ( .A1(adk_in[62]), .A2(n841), .Y(n374) );
  NAND3X0_HVT U358 ( .A1(n372), .A2(n373), .A3(n374), .Y(n222) );
  INVX0_HVT U359 ( .A(n962), .Y(n764) );
  INVX1_HVT U360 ( .A(n764), .Y(cipher_text[80]) );
  INVX0_HVT U361 ( .A(n979), .Y(n655) );
  NAND2X0_HVT U362 ( .A1(n338), .A2(n905), .Y(n375) );
  NAND2X0_HVT U363 ( .A1(adk_out0[39]), .A2(n879), .Y(n376) );
  NAND2X0_HVT U364 ( .A1(adk_in[39]), .A2(n840), .Y(n377) );
  NAND3X0_HVT U365 ( .A1(n375), .A2(n376), .A3(n377), .Y(n245) );
  NAND2X0_HVT U366 ( .A1(n986), .A2(n903), .Y(n378) );
  NAND2X0_HVT U367 ( .A1(adk_out0[56]), .A2(n877), .Y(n379) );
  NAND2X0_HVT U368 ( .A1(adk_in[56]), .A2(n841), .Y(n380) );
  NAND3X0_HVT U369 ( .A1(n378), .A2(n379), .A3(n380), .Y(n228) );
  INVX1_HVT U370 ( .A(n381), .Y(n382) );
  NAND2X0_HVT U371 ( .A1(n1018), .A2(n906), .Y(n383) );
  NAND2X0_HVT U372 ( .A1(adk_out0[24]), .A2(n880), .Y(n384) );
  NAND2X0_HVT U373 ( .A1(adk_in[24]), .A2(n838), .Y(n385) );
  NAND3X0_HVT U374 ( .A1(n383), .A2(n384), .A3(n385), .Y(n260) );
  INVX1_HVT U375 ( .A(n909), .Y(n906) );
  INVX0_HVT U376 ( .A(n668), .Y(n386) );
  INVX0_HVT U377 ( .A(n655), .Y(n389) );
  NAND2X0_HVT U378 ( .A1(n974), .A2(n902), .Y(n390) );
  NAND2X0_HVT U379 ( .A1(adk_out0[68]), .A2(n876), .Y(n391) );
  NAND2X0_HVT U380 ( .A1(adk_in[68]), .A2(n842), .Y(n392) );
  NAND3X0_HVT U381 ( .A1(n390), .A2(n391), .A3(n392), .Y(n216) );
  NAND2X0_HVT U382 ( .A1(n907), .A2(n1038), .Y(n393) );
  NAND2X0_HVT U383 ( .A1(adk_out0[4]), .A2(n881), .Y(n394) );
  NAND2X0_HVT U384 ( .A1(adk_in[4]), .A2(n837), .Y(n395) );
  NAND3X0_HVT U385 ( .A1(n393), .A2(n394), .A3(n395), .Y(n280) );
  INVX1_HVT U386 ( .A(n909), .Y(n907) );
  INVX1_HVT U387 ( .A(n768), .Y(cipher_text[115]) );
  INVX1_HVT U388 ( .A(n928), .Y(n768) );
  NAND2X0_HVT U389 ( .A1(n901), .A2(n336), .Y(n396) );
  NAND2X0_HVT U390 ( .A1(adk_out0[76]), .A2(n875), .Y(n397) );
  NAND2X0_HVT U391 ( .A1(adk_in[76]), .A2(n842), .Y(n398) );
  NAND3X0_HVT U392 ( .A1(n396), .A2(n397), .A3(n398), .Y(n208) );
  INVX1_HVT U393 ( .A(n550), .Y(n551) );
  AND2X1_HVT U394 ( .A1(n585), .A2(n584), .Y(n399) );
  AND2X1_HVT U395 ( .A1(n761), .A2(n760), .Y(n400) );
  AND2X1_HVT U396 ( .A1(n610), .A2(n609), .Y(n401) );
  INVX0_HVT U397 ( .A(n921), .Y(n402) );
  INVX0_HVT U398 ( .A(n402), .Y(cipher_text[122]) );
  NAND2X0_HVT U399 ( .A1(n900), .A2(n951), .Y(n404) );
  NAND2X0_HVT U400 ( .A1(adk_out0[91]), .A2(n874), .Y(n405) );
  NAND2X0_HVT U401 ( .A1(adk_in[91]), .A2(n844), .Y(n406) );
  NAND3X0_HVT U402 ( .A1(n404), .A2(n405), .A3(n406), .Y(n193) );
  INVX2_HVT U403 ( .A(n407), .Y(n408) );
  NAND2X0_HVT U404 ( .A1(n899), .A2(n936), .Y(n409) );
  NAND2X0_HVT U405 ( .A1(adk_out0[107]), .A2(n873), .Y(n410) );
  NAND2X0_HVT U406 ( .A1(adk_in[107]), .A2(n845), .Y(n411) );
  NAND3X0_HVT U407 ( .A1(n409), .A2(n410), .A3(n411), .Y(n177) );
  INVX1_HVT U408 ( .A(n948), .Y(n576) );
  INVX0_HVT U409 ( .A(n941), .Y(n412) );
  INVX0_HVT U410 ( .A(n412), .Y(cipher_text[101]) );
  NAND2X0_HVT U411 ( .A1(n905), .A2(n1006), .Y(n414) );
  NAND2X0_HVT U412 ( .A1(adk_out0[36]), .A2(n879), .Y(n415) );
  NAND2X0_HVT U413 ( .A1(adk_in[36]), .A2(n839), .Y(n416) );
  NAND3X0_HVT U414 ( .A1(n414), .A2(n415), .A3(n416), .Y(n248) );
  NAND2X0_HVT U415 ( .A1(n949), .A2(n900), .Y(n417) );
  NAND2X0_HVT U416 ( .A1(adk_out0[93]), .A2(n874), .Y(n418) );
  NAND2X0_HVT U417 ( .A1(adk_in[93]), .A2(n844), .Y(n419) );
  NAND3X0_HVT U418 ( .A1(n417), .A2(n418), .A3(n419), .Y(n191) );
  NAND2X0_HVT U419 ( .A1(n897), .A2(n918), .Y(n420) );
  NAND2X0_HVT U420 ( .A1(adk_out0[125]), .A2(n871), .Y(n421) );
  NAND2X0_HVT U421 ( .A1(adk_in[125]), .A2(n846), .Y(n422) );
  NAND3X0_HVT U422 ( .A1(n420), .A2(n421), .A3(n422), .Y(n159) );
  NAND2X0_HVT U423 ( .A1(n981), .A2(n903), .Y(n423) );
  NAND2X0_HVT U424 ( .A1(adk_out0[61]), .A2(n877), .Y(n424) );
  NAND2X0_HVT U425 ( .A1(adk_in[61]), .A2(n841), .Y(n425) );
  NAND3X0_HVT U426 ( .A1(n423), .A2(n424), .A3(n425), .Y(n223) );
  INVX0_HVT U427 ( .A(n959), .Y(n770) );
  NAND2X0_HVT U428 ( .A1(n930), .A2(n898), .Y(n426) );
  NAND2X0_HVT U429 ( .A1(adk_out0[113]), .A2(n872), .Y(n427) );
  NAND2X0_HVT U430 ( .A1(adk_in[113]), .A2(n845), .Y(n428) );
  NAND3X0_HVT U431 ( .A1(n426), .A2(n427), .A3(n428), .Y(n171) );
  NAND2X0_HVT U432 ( .A1(n900), .A2(n948), .Y(n429) );
  NAND2X0_HVT U433 ( .A1(adk_out0[94]), .A2(n874), .Y(n430) );
  NAND2X0_HVT U434 ( .A1(adk_in[94]), .A2(n844), .Y(n431) );
  NAND3X0_HVT U435 ( .A1(n429), .A2(n430), .A3(n431), .Y(n190) );
  INVX1_HVT U436 ( .A(n731), .Y(cipher_text[121]) );
  NAND2X0_HVT U437 ( .A1(n898), .A2(n928), .Y(n432) );
  NAND2X0_HVT U438 ( .A1(adk_out0[115]), .A2(n872), .Y(n433) );
  NAND2X0_HVT U439 ( .A1(adk_in[115]), .A2(n845), .Y(n434) );
  NAND3X0_HVT U440 ( .A1(n432), .A2(n433), .A3(n434), .Y(n169) );
  INVX1_HVT U441 ( .A(n922), .Y(n731) );
  INVX0_HVT U442 ( .A(n950), .Y(n814) );
  INVX1_HVT U443 ( .A(n770), .Y(cipher_text[83]) );
  NAND2X0_HVT U444 ( .A1(n400), .A2(n759), .Y(n185) );
  INVX0_HVT U445 ( .A(n940), .Y(n435) );
  INVX0_HVT U446 ( .A(n435), .Y(cipher_text[102]) );
  NAND2X0_HVT U447 ( .A1(n901), .A2(n961), .Y(n437) );
  NAND2X0_HVT U448 ( .A1(adk_out0[81]), .A2(n875), .Y(n438) );
  NAND2X0_HVT U449 ( .A1(adk_in[81]), .A2(n843), .Y(n439) );
  NAND3X0_HVT U450 ( .A1(n437), .A2(n438), .A3(n439), .Y(n203) );
  INVX0_HVT U451 ( .A(n990), .Y(n820) );
  INVX0_HVT U452 ( .A(n998), .Y(n804) );
  INVX0_HVT U453 ( .A(n937), .Y(n440) );
  INVX0_HVT U454 ( .A(n440), .Y(cipher_text[106]) );
  NAND2X0_HVT U455 ( .A1(n955), .A2(n901), .Y(n442) );
  NAND2X0_HVT U456 ( .A1(adk_out0[87]), .A2(n875), .Y(n443) );
  NAND2X0_HVT U457 ( .A1(adk_in[87]), .A2(n843), .Y(n444) );
  NAND3X0_HVT U458 ( .A1(n442), .A2(n443), .A3(n444), .Y(n197) );
  NAND2X0_HVT U459 ( .A1(n997), .A2(n904), .Y(n445) );
  NAND2X0_HVT U460 ( .A1(adk_out0[45]), .A2(n878), .Y(n446) );
  NAND2X0_HVT U461 ( .A1(adk_in[45]), .A2(n840), .Y(n447) );
  NAND3X0_HVT U462 ( .A1(n445), .A2(n446), .A3(n447), .Y(n239) );
  INVX1_HVT U463 ( .A(n448), .Y(n449) );
  INVX1_HVT U464 ( .A(n546), .Y(cipher_text[38]) );
  NAND2X0_HVT U465 ( .A1(n903), .A2(n389), .Y(n450) );
  NAND2X0_HVT U466 ( .A1(adk_out0[63]), .A2(n877), .Y(n451) );
  NAND2X0_HVT U467 ( .A1(adk_in[63]), .A2(n841), .Y(n452) );
  NAND3X0_HVT U468 ( .A1(n450), .A2(n451), .A3(n452), .Y(n221) );
  INVX0_HVT U469 ( .A(n1039), .Y(n792) );
  INVX2_HVT U470 ( .A(n611), .Y(n612) );
  NAND2X0_HVT U471 ( .A1(n1020), .A2(n906), .Y(n453) );
  NAND2X0_HVT U472 ( .A1(adk_out0[22]), .A2(n880), .Y(n454) );
  NAND2X0_HVT U473 ( .A1(adk_in[22]), .A2(n838), .Y(n455) );
  NAND3X0_HVT U474 ( .A1(n453), .A2(n454), .A3(n455), .Y(n262) );
  INVX1_HVT U475 ( .A(n1020), .Y(n456) );
  INVX1_HVT U476 ( .A(n456), .Y(cipher_text[22]) );
  INVX1_HVT U477 ( .A(n814), .Y(cipher_text[92]) );
  NAND2X0_HVT U478 ( .A1(n1012), .A2(n905), .Y(n458) );
  NAND2X0_HVT U479 ( .A1(adk_out0[30]), .A2(n879), .Y(n459) );
  NAND2X0_HVT U480 ( .A1(adk_in[30]), .A2(n839), .Y(n460) );
  NAND3X0_HVT U481 ( .A1(n458), .A2(n459), .A3(n460), .Y(n254) );
  INVX1_HVT U482 ( .A(n668), .Y(cipher_text[41]) );
  INVX1_HVT U483 ( .A(n461), .Y(n462) );
  INVX0_HVT U484 ( .A(n991), .Y(n604) );
  INVX0_HVT U485 ( .A(n958), .Y(n822) );
  NAND2X0_HVT U486 ( .A1(n959), .A2(n901), .Y(n463) );
  NAND2X0_HVT U487 ( .A1(adk_out0[83]), .A2(n875), .Y(n464) );
  NAND2X0_HVT U488 ( .A1(adk_in[83]), .A2(n843), .Y(n465) );
  NAND3X0_HVT U489 ( .A1(n463), .A2(n464), .A3(n465), .Y(n201) );
  INVX0_HVT U490 ( .A(n1035), .Y(n466) );
  INVX0_HVT U491 ( .A(n466), .Y(cipher_text[7]) );
  INVX1_HVT U492 ( .A(n468), .Y(n469) );
  INVX1_HVT U493 ( .A(n686), .Y(cipher_text[34]) );
  INVX0_HVT U494 ( .A(n927), .Y(n470) );
  INVX0_HVT U495 ( .A(n470), .Y(cipher_text[116]) );
  NAND2X0_HVT U496 ( .A1(n962), .A2(n901), .Y(n472) );
  NAND2X0_HVT U497 ( .A1(adk_out0[80]), .A2(n875), .Y(n473) );
  NAND2X0_HVT U498 ( .A1(adk_in[80]), .A2(n843), .Y(n474) );
  NAND3X0_HVT U499 ( .A1(n472), .A2(n473), .A3(n474), .Y(n204) );
  NAND2X0_HVT U500 ( .A1(n386), .A2(n904), .Y(n475) );
  NAND2X0_HVT U501 ( .A1(adk_out0[41]), .A2(n878), .Y(n476) );
  NAND2X0_HVT U502 ( .A1(adk_in[41]), .A2(n840), .Y(n477) );
  NAND3X0_HVT U503 ( .A1(n475), .A2(n476), .A3(n477), .Y(n243) );
  NAND2X0_HVT U504 ( .A1(n898), .A2(n922), .Y(n478) );
  NAND2X0_HVT U505 ( .A1(adk_out0[121]), .A2(n872), .Y(n479) );
  NAND2X0_HVT U506 ( .A1(adk_in[121]), .A2(n846), .Y(n480) );
  NAND3X0_HVT U507 ( .A1(n478), .A2(n479), .A3(n480), .Y(n163) );
  INVX1_HVT U508 ( .A(n910), .Y(n898) );
  INVX1_HVT U509 ( .A(n701), .Y(cipher_text[89]) );
  INVX1_HVT U510 ( .A(n481), .Y(cipher_text[11]) );
  INVX1_HVT U511 ( .A(n483), .Y(n484) );
  NAND2X0_HVT U512 ( .A1(n919), .A2(n897), .Y(n485) );
  NAND2X0_HVT U513 ( .A1(adk_out0[124]), .A2(n871), .Y(n486) );
  NAND2X0_HVT U514 ( .A1(adk_in[124]), .A2(n846), .Y(n487) );
  NAND3X0_HVT U515 ( .A1(n485), .A2(n486), .A3(n487), .Y(n160) );
  INVX0_HVT U516 ( .A(n939), .Y(n492) );
  INVX0_HVT U517 ( .A(n492), .Y(cipher_text[104]) );
  INVX0_HVT U518 ( .A(n985), .Y(n548) );
  NAND2X0_HVT U519 ( .A1(n901), .A2(n960), .Y(n494) );
  NAND2X0_HVT U520 ( .A1(adk_out0[82]), .A2(n875), .Y(n495) );
  NAND2X0_HVT U521 ( .A1(adk_in[82]), .A2(n843), .Y(n496) );
  NAND3X0_HVT U522 ( .A1(n494), .A2(n495), .A3(n496), .Y(n202) );
  INVX1_HVT U523 ( .A(n960), .Y(n707) );
  INVX0_HVT U524 ( .A(n925), .Y(n497) );
  INVX0_HVT U525 ( .A(n497), .Y(cipher_text[118]) );
  NAND2X0_HVT U526 ( .A1(n989), .A2(n903), .Y(n499) );
  NAND2X0_HVT U527 ( .A1(adk_out0[53]), .A2(n877), .Y(n500) );
  NAND2X0_HVT U528 ( .A1(adk_in[53]), .A2(n841), .Y(n501) );
  NAND3X0_HVT U529 ( .A1(n499), .A2(n500), .A3(n501), .Y(n231) );
  INVX1_HVT U530 ( .A(n909), .Y(n903) );
  NAND2X0_HVT U531 ( .A1(n1013), .A2(n905), .Y(n502) );
  NAND2X0_HVT U532 ( .A1(adk_out0[29]), .A2(n879), .Y(n503) );
  NAND2X0_HVT U533 ( .A1(adk_in[29]), .A2(n839), .Y(n504) );
  NAND3X0_HVT U534 ( .A1(n502), .A2(n503), .A3(n504), .Y(n255) );
  INVX0_HVT U535 ( .A(n1028), .Y(n507) );
  INVX0_HVT U536 ( .A(n507), .Y(cipher_text[14]) );
  INVX1_HVT U537 ( .A(n565), .Y(cipher_text[111]) );
  INVX1_HVT U538 ( .A(n932), .Y(n565) );
  NAND2X0_HVT U539 ( .A1(n953), .A2(n900), .Y(n509) );
  NAND2X0_HVT U540 ( .A1(adk_out0[89]), .A2(n874), .Y(n510) );
  NAND2X0_HVT U541 ( .A1(adk_in[89]), .A2(n843), .Y(n511) );
  NAND3X0_HVT U542 ( .A1(n509), .A2(n510), .A3(n511), .Y(n195) );
  INVX0_HVT U543 ( .A(n1007), .Y(n695) );
  NAND2X0_HVT U544 ( .A1(n899), .A2(n932), .Y(n512) );
  NAND2X0_HVT U545 ( .A1(adk_out0[111]), .A2(n873), .Y(n513) );
  NAND2X0_HVT U546 ( .A1(adk_in[111]), .A2(n845), .Y(n514) );
  NAND3X0_HVT U547 ( .A1(n512), .A2(n513), .A3(n514), .Y(n173) );
  NAND2X0_HVT U548 ( .A1(n900), .A2(n950), .Y(n515) );
  NAND2X0_HVT U549 ( .A1(adk_out0[92]), .A2(n874), .Y(n516) );
  NAND2X0_HVT U550 ( .A1(adk_in[92]), .A2(n844), .Y(n517) );
  NAND3X0_HVT U551 ( .A1(n515), .A2(n516), .A3(n517), .Y(n192) );
  INVX1_HVT U552 ( .A(n910), .Y(n900) );
  INVX1_HVT U553 ( .A(n518), .Y(n519) );
  NAND2X0_HVT U554 ( .A1(n1008), .A2(n905), .Y(n520) );
  NAND2X0_HVT U555 ( .A1(adk_out0[34]), .A2(n879), .Y(n521) );
  NAND2X0_HVT U556 ( .A1(adk_in[34]), .A2(n839), .Y(n522) );
  NAND3X0_HVT U557 ( .A1(n520), .A2(n521), .A3(n522), .Y(n250) );
  INVX1_HVT U558 ( .A(n909), .Y(n905) );
  INVX1_HVT U559 ( .A(n525), .Y(n526) );
  INVX0_HVT U560 ( .A(n1019), .Y(n527) );
  INVX0_HVT U561 ( .A(n527), .Y(cipher_text[23]) );
  INVX0_HVT U562 ( .A(n954), .Y(n529) );
  INVX0_HVT U563 ( .A(n529), .Y(cipher_text[88]) );
  INVX0_HVT U564 ( .A(n1037), .Y(n531) );
  INVX0_HVT U565 ( .A(n531), .Y(cipher_text[5]) );
  INVX1_HVT U566 ( .A(n930), .Y(n535) );
  INVX1_HVT U567 ( .A(n535), .Y(cipher_text[113]) );
  INVX2_HVT U568 ( .A(n537), .Y(n538) );
  INVX0_HVT U569 ( .A(n996), .Y(n539) );
  INVX0_HVT U570 ( .A(n539), .Y(cipher_text[46]) );
  INVX0_HVT U571 ( .A(n924), .Y(n541) );
  INVX0_HVT U572 ( .A(n541), .Y(cipher_text[119]) );
  NAND2X0_HVT U573 ( .A1(n1004), .A2(n905), .Y(n543) );
  NAND2X0_HVT U574 ( .A1(adk_out0[38]), .A2(n879), .Y(n544) );
  NAND2X0_HVT U575 ( .A1(adk_in[38]), .A2(n840), .Y(n545) );
  NAND3X0_HVT U576 ( .A1(n543), .A2(n544), .A3(n545), .Y(n246) );
  INVX0_HVT U577 ( .A(n1004), .Y(n546) );
  NAND2X0_HVT U578 ( .A1(n908), .A2(n982), .Y(n552) );
  NAND2X0_HVT U579 ( .A1(adk_out0[60]), .A2(n877), .Y(n553) );
  NAND2X0_HVT U580 ( .A1(n631), .A2(n841), .Y(n554) );
  NAND3X0_HVT U581 ( .A1(n552), .A2(n553), .A3(n554), .Y(n224) );
  INVX0_HVT U582 ( .A(n972), .Y(n555) );
  INVX0_HVT U583 ( .A(n555), .Y(cipher_text[70]) );
  INVX0_HVT U584 ( .A(n993), .Y(n557) );
  INVX0_HVT U585 ( .A(n557), .Y(cipher_text[49]) );
  NAND2X0_HVT U586 ( .A1(n399), .A2(n583), .Y(n251) );
  INVX0_HVT U587 ( .A(n1009), .Y(n559) );
  INVX0_HVT U588 ( .A(n559), .Y(cipher_text[33]) );
  INVX0_HVT U589 ( .A(n1005), .Y(n561) );
  INVX0_HVT U590 ( .A(n561), .Y(cipher_text[37]) );
  INVX0_HVT U591 ( .A(n1021), .Y(n563) );
  INVX0_HVT U592 ( .A(n563), .Y(cipher_text[21]) );
  INVX0_HVT U593 ( .A(n956), .Y(n567) );
  INVX0_HVT U594 ( .A(n567), .Y(cipher_text[86]) );
  INVX2_HVT U595 ( .A(n738), .Y(n739) );
  NAND2X0_HVT U596 ( .A1(cipher_text[103]), .A2(n899), .Y(n569) );
  NAND2X0_HVT U597 ( .A1(adk_out0[103]), .A2(n873), .Y(n570) );
  NAND2X0_HVT U598 ( .A1(adk_in[103]), .A2(n845), .Y(n571) );
  NAND2X0_HVT U599 ( .A1(n401), .A2(n608), .Y(n227) );
  INVX0_HVT U600 ( .A(n572), .Y(cipher_text[54]) );
  INVX0_HVT U601 ( .A(n576), .Y(cipher_text[94]) );
  INVX1_HVT U602 ( .A(n799), .Y(cipher_text[20]) );
  INVX0_HVT U603 ( .A(n947), .Y(n578) );
  INVX0_HVT U604 ( .A(n578), .Y(cipher_text[95]) );
  NBUFFX2_HVT U605 ( .A(n955), .Y(cipher_text[87]) );
  INVX0_HVT U606 ( .A(n1029), .Y(n581) );
  INVX0_HVT U607 ( .A(n581), .Y(cipher_text[13]) );
  NAND2X0_HVT U608 ( .A1(n1009), .A2(n905), .Y(n583) );
  NAND2X0_HVT U609 ( .A1(adk_out0[33]), .A2(n879), .Y(n584) );
  NAND2X0_HVT U610 ( .A1(adk_in[33]), .A2(n839), .Y(n585) );
  NAND2X0_HVT U611 ( .A1(n987), .A2(n903), .Y(n586) );
  NAND2X0_HVT U612 ( .A1(adk_out0[55]), .A2(n877), .Y(n587) );
  NAND2X0_HVT U613 ( .A1(adk_in[55]), .A2(n841), .Y(n588) );
  NAND3X0_HVT U614 ( .A1(n586), .A2(n587), .A3(n588), .Y(n229) );
  INVX1_HVT U615 ( .A(n987), .Y(n589) );
  INVX1_HVT U616 ( .A(n589), .Y(cipher_text[55]) );
  INVX0_HVT U617 ( .A(n1012), .Y(n591) );
  INVX0_HVT U618 ( .A(n591), .Y(cipher_text[30]) );
  INVX0_HVT U619 ( .A(n1002), .Y(n593) );
  INVX0_HVT U620 ( .A(n593), .Y(cipher_text[40]) );
  NAND2X0_HVT U621 ( .A1(n995), .A2(n904), .Y(n595) );
  NAND2X0_HVT U622 ( .A1(adk_out0[47]), .A2(n878), .Y(n596) );
  NAND2X0_HVT U623 ( .A1(adk_in[47]), .A2(n840), .Y(n597) );
  NAND3X0_HVT U624 ( .A1(n595), .A2(n596), .A3(n597), .Y(n237) );
  INVX1_HVT U625 ( .A(n995), .Y(n598) );
  INVX1_HVT U626 ( .A(n598), .Y(cipher_text[47]) );
  INVX1_HVT U627 ( .A(n604), .Y(cipher_text[51]) );
  INVX0_HVT U628 ( .A(n961), .Y(n606) );
  NAND2X0_HVT U629 ( .A1(n344), .A2(n903), .Y(n608) );
  NAND2X0_HVT U630 ( .A1(adk_out0[57]), .A2(n877), .Y(n609) );
  NAND2X0_HVT U631 ( .A1(adk_in[57]), .A2(n841), .Y(n610) );
  INVX0_HVT U632 ( .A(n945), .Y(n613) );
  INVX0_HVT U633 ( .A(n613), .Y(cipher_text[97]) );
  AND2X1_HVT U634 ( .A1(n746), .A2(n747), .Y(n615) );
  INVX1_HVT U635 ( .A(n836), .Y(n886) );
  INVX1_HVT U636 ( .A(n886), .Y(n885) );
  INVX1_HVT U637 ( .A(n886), .Y(n884) );
  NBUFFX2_HVT U638 ( .A(n970), .Y(cipher_text[72]) );
  NBUFFX2_HVT U639 ( .A(n1034), .Y(cipher_text[8]) );
  NBUFFX2_HVT U640 ( .A(n1010), .Y(cipher_text[32]) );
  NBUFFX2_HVT U641 ( .A(n978), .Y(cipher_text[64]) );
  NBUFFX2_HVT U642 ( .A(n944), .Y(cipher_text[98]) );
  NBUFFX2_HVT U643 ( .A(n933), .Y(cipher_text[110]) );
  INVX0_HVT U644 ( .A(n957), .Y(n625) );
  INVX0_HVT U645 ( .A(n625), .Y(cipher_text[85]) );
  INVX0_HVT U646 ( .A(n973), .Y(n627) );
  INVX0_HVT U647 ( .A(n627), .Y(cipher_text[69]) );
  INVX0_HVT U648 ( .A(n917), .Y(n629) );
  INVX0_HVT U649 ( .A(n629), .Y(cipher_text[126]) );
  INVX1_HVT U650 ( .A(n634), .Y(n631) );
  INVX0_HVT U651 ( .A(n964), .Y(n632) );
  INVX0_HVT U652 ( .A(n632), .Y(cipher_text[78]) );
  INVX0_HVT U653 ( .A(n980), .Y(n637) );
  INVX0_HVT U654 ( .A(n637), .Y(cipher_text[62]) );
  INVX0_HVT U655 ( .A(n935), .Y(n639) );
  INVX0_HVT U656 ( .A(n639), .Y(cipher_text[108]) );
  INVX0_HVT U657 ( .A(n946), .Y(n641) );
  INVX0_HVT U658 ( .A(n641), .Y(cipher_text[96]) );
  INVX0_HVT U659 ( .A(n1033), .Y(n643) );
  INVX0_HVT U660 ( .A(n1015), .Y(n645) );
  INVX0_HVT U661 ( .A(n645), .Y(cipher_text[27]) );
  INVX1_HVT U662 ( .A(n820), .Y(cipher_text[52]) );
  INVX0_HVT U663 ( .A(n1036), .Y(n651) );
  INVX0_HVT U664 ( .A(n651), .Y(cipher_text[6]) );
  INVX1_HVT U665 ( .A(n772), .Y(cipher_text[43]) );
  INVX1_HVT U666 ( .A(n653), .Y(n654) );
  NAND2X0_HVT U667 ( .A1(n615), .A2(n745), .Y(n273) );
  INVX0_HVT U668 ( .A(n655), .Y(cipher_text[63]) );
  INVX0_HVT U669 ( .A(n657), .Y(cipher_text[117]) );
  INVX0_HVT U670 ( .A(n934), .Y(n659) );
  INVX0_HVT U671 ( .A(n659), .Y(cipher_text[109]) );
  INVX0_HVT U672 ( .A(n975), .Y(n806) );
  INVX1_HVT U673 ( .A(n806), .Y(cipher_text[67]) );
  NAND2X0_HVT U674 ( .A1(n990), .A2(n903), .Y(n661) );
  NAND2X0_HVT U675 ( .A1(adk_out0[52]), .A2(n877), .Y(n662) );
  NAND2X0_HVT U676 ( .A1(adk_in[52]), .A2(n841), .Y(n663) );
  NAND3X0_HVT U677 ( .A1(n661), .A2(n662), .A3(n663), .Y(n232) );
  INVX0_HVT U678 ( .A(n971), .Y(n664) );
  INVX0_HVT U679 ( .A(n664), .Y(cipher_text[71]) );
  INVX0_HVT U680 ( .A(n992), .Y(n670) );
  INVX0_HVT U681 ( .A(n670), .Y(cipher_text[50]) );
  INVX0_HVT U682 ( .A(n1042), .Y(n672) );
  INVX0_HVT U683 ( .A(n672), .Y(cipher_text[0]) );
  INVX1_HVT U684 ( .A(n810), .Y(cipher_text[59]) );
  INVX0_HVT U685 ( .A(n1024), .Y(n674) );
  INVX0_HVT U686 ( .A(n674), .Y(cipher_text[18]) );
  NAND2X0_HVT U687 ( .A1(n1040), .A2(n908), .Y(n676) );
  NAND2X0_HVT U688 ( .A1(adk_out0[2]), .A2(n882), .Y(n677) );
  NAND2X0_HVT U689 ( .A1(adk_in[2]), .A2(n837), .Y(n678) );
  NAND3X0_HVT U690 ( .A1(n676), .A2(n677), .A3(n678), .Y(n282) );
  INVX1_HVT U691 ( .A(n1040), .Y(n679) );
  INVX1_HVT U692 ( .A(n679), .Y(cipher_text[2]) );
  INVX0_HVT U693 ( .A(n1032), .Y(n681) );
  INVX0_HVT U694 ( .A(n681), .Y(cipher_text[10]) );
  NAND2X0_HVT U695 ( .A1(n903), .A2(n311), .Y(n683) );
  NAND2X0_HVT U696 ( .A1(adk_out0[59]), .A2(n877), .Y(n684) );
  NAND2X0_HVT U697 ( .A1(adk_in[59]), .A2(n841), .Y(n685) );
  NAND3X0_HVT U698 ( .A1(n683), .A2(n684), .A3(n685), .Y(n225) );
  INVX0_HVT U699 ( .A(n929), .Y(n690) );
  INVX0_HVT U700 ( .A(n690), .Y(cipher_text[114]) );
  NAND2X0_HVT U701 ( .A1(n904), .A2(n291), .Y(n692) );
  NAND2X0_HVT U702 ( .A1(adk_out0[43]), .A2(n878), .Y(n693) );
  NAND2X0_HVT U703 ( .A1(adk_in[43]), .A2(n840), .Y(n694) );
  NAND3X0_HVT U704 ( .A1(n692), .A2(n693), .A3(n694), .Y(n241) );
  INVX1_HVT U705 ( .A(n695), .Y(cipher_text[35]) );
  INVX0_HVT U706 ( .A(n994), .Y(n697) );
  INVX0_HVT U707 ( .A(n697), .Y(cipher_text[48]) );
  INVX1_HVT U708 ( .A(n703), .Y(n704) );
  INVX0_HVT U709 ( .A(n938), .Y(n705) );
  INVX0_HVT U710 ( .A(n705), .Y(cipher_text[105]) );
  INVX0_HVT U711 ( .A(n707), .Y(cipher_text[82]) );
  INVX0_HVT U712 ( .A(n977), .Y(n709) );
  INVX0_HVT U713 ( .A(n709), .Y(cipher_text[65]) );
  INVX0_HVT U714 ( .A(n969), .Y(n711) );
  INVX0_HVT U715 ( .A(n711), .Y(cipher_text[73]) );
  NAND2X0_HVT U716 ( .A1(n920), .A2(n898), .Y(n713) );
  NAND2X0_HVT U717 ( .A1(adk_out0[123]), .A2(n872), .Y(n714) );
  NAND2X0_HVT U718 ( .A1(adk_in[123]), .A2(n846), .Y(n715) );
  NAND3X0_HVT U719 ( .A1(n713), .A2(n714), .A3(n715), .Y(n161) );
  INVX0_HVT U720 ( .A(n920), .Y(n716) );
  INVX0_HVT U721 ( .A(n716), .Y(cipher_text[123]) );
  INVX0_HVT U722 ( .A(n718), .Y(cipher_text[127]) );
  INVX0_HVT U723 ( .A(n968), .Y(n720) );
  INVX0_HVT U724 ( .A(n720), .Y(cipher_text[74]) );
  INVX0_HVT U725 ( .A(n976), .Y(n722) );
  INVX0_HVT U726 ( .A(n722), .Y(cipher_text[66]) );
  INVX0_HVT U727 ( .A(n724), .Y(cipher_text[16]) );
  NAND2X0_HVT U728 ( .A1(n1014), .A2(n905), .Y(n726) );
  NAND2X0_HVT U729 ( .A1(adk_out0[28]), .A2(n879), .Y(n727) );
  NAND2X0_HVT U730 ( .A1(adk_in[28]), .A2(n839), .Y(n728) );
  NAND3X0_HVT U731 ( .A1(n726), .A2(n727), .A3(n728), .Y(n256) );
  INVX1_HVT U732 ( .A(n729), .Y(cipher_text[28]) );
  INVX0_HVT U733 ( .A(n1025), .Y(n733) );
  INVX0_HVT U734 ( .A(n733), .Y(cipher_text[17]) );
  NAND2X0_HVT U735 ( .A1(n975), .A2(n902), .Y(n735) );
  NAND2X0_HVT U736 ( .A1(adk_out0[67]), .A2(n876), .Y(n736) );
  NAND2X0_HVT U737 ( .A1(adk_in[67]), .A2(n842), .Y(n737) );
  NAND3X0_HVT U738 ( .A1(n735), .A2(n736), .A3(n737), .Y(n217) );
  INVX1_HVT U739 ( .A(n910), .Y(n902) );
  INVX0_HVT U740 ( .A(n952), .Y(n740) );
  INVX0_HVT U741 ( .A(n740), .Y(cipher_text[90]) );
  INVX1_HVT U742 ( .A(n742), .Y(cipher_text[75]) );
  NBUFFX2_HVT U743 ( .A(n1011), .Y(cipher_text[31]) );
  NAND2X0_HVT U744 ( .A1(n1031), .A2(n15), .Y(n745) );
  NAND2X0_HVT U745 ( .A1(adk_in[11]), .A2(n17), .Y(n746) );
  NAND2X0_HVT U746 ( .A1(adk_out0[11]), .A2(n881), .Y(n747) );
  INVX1_HVT U747 ( .A(n812), .Y(cipher_text[19]) );
  NAND2X0_HVT U748 ( .A1(n1022), .A2(n906), .Y(n748) );
  NAND2X0_HVT U749 ( .A1(adk_out0[20]), .A2(n880), .Y(n749) );
  NAND2X0_HVT U750 ( .A1(adk_in[20]), .A2(n838), .Y(n750) );
  NAND3X0_HVT U751 ( .A1(n748), .A2(n749), .A3(n750), .Y(n264) );
  NAND2X0_HVT U752 ( .A1(n1030), .A2(n907), .Y(n751) );
  NAND2X0_HVT U753 ( .A1(adk_out0[12]), .A2(n881), .Y(n752) );
  NAND2X0_HVT U754 ( .A1(adk_in[12]), .A2(n838), .Y(n753) );
  NAND3X0_HVT U755 ( .A1(n751), .A2(n752), .A3(n753), .Y(n272) );
  INVX1_HVT U756 ( .A(n754), .Y(cipher_text[12]) );
  NAND2X0_HVT U757 ( .A1(n906), .A2(n1023), .Y(n756) );
  NAND2X0_HVT U758 ( .A1(adk_out0[19]), .A2(n880), .Y(n757) );
  NAND2X0_HVT U759 ( .A1(adk_in[19]), .A2(n838), .Y(n758) );
  NAND3X0_HVT U760 ( .A1(n756), .A2(n757), .A3(n758), .Y(n265) );
  INVX1_HVT U761 ( .A(n857), .Y(n838) );
  NAND2X0_HVT U762 ( .A1(n943), .A2(n900), .Y(n759) );
  NAND2X0_HVT U763 ( .A1(adk_out0[99]), .A2(n874), .Y(n760) );
  NAND2X0_HVT U764 ( .A1(adk_in[99]), .A2(n844), .Y(n761) );
  INVX0_HVT U765 ( .A(n963), .Y(n762) );
  INVX0_HVT U766 ( .A(n762), .Y(cipher_text[79]) );
  INVX0_HVT U767 ( .A(n1006), .Y(n766) );
  INVX1_HVT U768 ( .A(n804), .Y(cipher_text[44]) );
  NAND2X0_HVT U769 ( .A1(n998), .A2(n904), .Y(n774) );
  NAND2X0_HVT U770 ( .A1(adk_out0[44]), .A2(n878), .Y(n775) );
  NAND2X0_HVT U771 ( .A1(adk_in[44]), .A2(n840), .Y(n776) );
  NAND3X0_HVT U772 ( .A1(n774), .A2(n775), .A3(n776), .Y(n240) );
  INVX1_HVT U773 ( .A(n909), .Y(n904) );
  INVX1_HVT U774 ( .A(n857), .Y(n840) );
  NAND2X0_HVT U775 ( .A1(n1015), .A2(n906), .Y(n777) );
  NAND2X0_HVT U776 ( .A1(adk_out0[27]), .A2(n880), .Y(n778) );
  NAND2X0_HVT U777 ( .A1(adk_in[27]), .A2(n839), .Y(n779) );
  NAND3X0_HVT U778 ( .A1(n777), .A2(n778), .A3(n779), .Y(n257) );
  NAND2X0_HVT U779 ( .A1(n901), .A2(n958), .Y(n780) );
  NAND2X0_HVT U780 ( .A1(adk_out0[84]), .A2(n875), .Y(n781) );
  NAND2X0_HVT U781 ( .A1(adk_in[84]), .A2(n843), .Y(n782) );
  NAND3X0_HVT U782 ( .A1(n780), .A2(n781), .A3(n782), .Y(n200) );
  INVX1_HVT U783 ( .A(n910), .Y(n901) );
  NAND2X0_HVT U784 ( .A1(n991), .A2(n904), .Y(n783) );
  NAND2X0_HVT U785 ( .A1(adk_out0[51]), .A2(n878), .Y(n784) );
  NAND2X0_HVT U786 ( .A1(adk_in[51]), .A2(n841), .Y(n785) );
  NAND3X0_HVT U787 ( .A1(n783), .A2(n784), .A3(n785), .Y(n233) );
  INVX1_HVT U788 ( .A(n857), .Y(n841) );
  NAND2X0_HVT U789 ( .A1(n1007), .A2(n905), .Y(n786) );
  NAND2X0_HVT U790 ( .A1(adk_out0[35]), .A2(n879), .Y(n787) );
  NAND2X0_HVT U791 ( .A1(adk_in[35]), .A2(n839), .Y(n788) );
  NAND3X0_HVT U792 ( .A1(n786), .A2(n787), .A3(n788), .Y(n249) );
  INVX1_HVT U793 ( .A(n857), .Y(n839) );
  NAND2X0_HVT U794 ( .A1(n1039), .A2(n908), .Y(n789) );
  NAND2X0_HVT U795 ( .A1(adk_out0[3]), .A2(n882), .Y(n790) );
  NAND2X0_HVT U796 ( .A1(n362), .A2(n837), .Y(n791) );
  NAND3X0_HVT U797 ( .A1(n789), .A2(n790), .A3(n791), .Y(n281) );
  INVX1_HVT U798 ( .A(n792), .Y(cipher_text[3]) );
  INVX0_HVT U799 ( .A(n883), .Y(n882) );
  NBUFFX2_HVT U800 ( .A(n974), .Y(cipher_text[68]) );
  INVX0_HVT U801 ( .A(n936), .Y(n795) );
  INVX0_HVT U802 ( .A(n795), .Y(cipher_text[107]) );
  INVX0_HVT U803 ( .A(n797), .Y(cipher_text[60]) );
  NAND2X0_HVT U804 ( .A1(n902), .A2(n323), .Y(n801) );
  NAND2X0_HVT U805 ( .A1(adk_out0[75]), .A2(n876), .Y(n802) );
  NAND2X0_HVT U806 ( .A1(adk_in[75]), .A2(n842), .Y(n803) );
  NAND3X0_HVT U807 ( .A1(n801), .A2(n802), .A3(n803), .Y(n209) );
  INVX1_HVT U808 ( .A(n857), .Y(n842) );
  INVX0_HVT U809 ( .A(n951), .Y(n816) );
  INVX0_HVT U810 ( .A(n816), .Y(cipher_text[91]) );
  INVX0_HVT U811 ( .A(n822), .Y(cipher_text[84]) );
  NAND2X0_HVT U812 ( .A1(n965), .A2(n901), .Y(n824) );
  NAND2X0_HVT U813 ( .A1(adk_out0[77]), .A2(n875), .Y(n825) );
  NAND2X0_HVT U814 ( .A1(adk_in[77]), .A2(n843), .Y(n826) );
  NAND3X0_HVT U815 ( .A1(n824), .A2(n825), .A3(n826), .Y(n207) );
  INVX1_HVT U816 ( .A(n965), .Y(n827) );
  INVX1_HVT U817 ( .A(n827), .Y(cipher_text[77]) );
  NBUFFX2_HVT U818 ( .A(n981), .Y(cipher_text[61]) );
  NBUFFX2_HVT U819 ( .A(n918), .Y(cipher_text[125]) );
  INVX0_HVT U820 ( .A(n1016), .Y(n834) );
  INVX0_HVT U821 ( .A(n834), .Y(cipher_text[26]) );
  INVX0_HVT U822 ( .A(n886), .Y(n883) );
  INVX0_HVT U823 ( .A(n909), .Y(n908) );
  INVX0_HVT U824 ( .A(n15), .Y(n912) );
  INVX0_HVT U825 ( .A(n17), .Y(n858) );
  INVX0_HVT U826 ( .A(n17), .Y(n860) );
  INVX0_HVT U827 ( .A(n17), .Y(n859) );
  INVX1_HVT U828 ( .A(n911), .Y(n891) );
  INVX1_HVT U829 ( .A(n911), .Y(n892) );
  INVX1_HVT U830 ( .A(n911), .Y(n893) );
  INVX1_HVT U831 ( .A(n911), .Y(n894) );
  INVX1_HVT U832 ( .A(n911), .Y(n895) );
  INVX1_HVT U833 ( .A(n910), .Y(n897) );
  INVX1_HVT U834 ( .A(n910), .Y(n899) );
  INVX1_HVT U835 ( .A(n911), .Y(n896) );
  INVX1_HVT U836 ( .A(n912), .Y(n887) );
  INVX1_HVT U837 ( .A(n912), .Y(n888) );
  INVX1_HVT U838 ( .A(n912), .Y(n889) );
  INVX1_HVT U839 ( .A(n912), .Y(n890) );
  INVX1_HVT U840 ( .A(n883), .Y(n877) );
  INVX1_HVT U841 ( .A(n883), .Y(n878) );
  INVX1_HVT U842 ( .A(n883), .Y(n879) );
  INVX1_HVT U843 ( .A(n883), .Y(n880) );
  INVX1_HVT U844 ( .A(n884), .Y(n865) );
  INVX1_HVT U845 ( .A(n884), .Y(n866) );
  INVX1_HVT U846 ( .A(n884), .Y(n867) );
  INVX1_HVT U847 ( .A(n884), .Y(n868) );
  INVX1_HVT U848 ( .A(n884), .Y(n869) );
  INVX1_HVT U849 ( .A(n885), .Y(n871) );
  INVX1_HVT U850 ( .A(n885), .Y(n872) );
  INVX1_HVT U851 ( .A(n885), .Y(n873) );
  INVX1_HVT U852 ( .A(n884), .Y(n874) );
  INVX1_HVT U853 ( .A(n885), .Y(n875) );
  INVX1_HVT U854 ( .A(n883), .Y(n881) );
  INVX1_HVT U855 ( .A(n884), .Y(n870) );
  INVX1_HVT U856 ( .A(n836), .Y(n876) );
  INVX1_HVT U857 ( .A(n885), .Y(n861) );
  INVX1_HVT U858 ( .A(n885), .Y(n862) );
  INVX1_HVT U859 ( .A(n885), .Y(n863) );
  INVX1_HVT U860 ( .A(n885), .Y(n864) );
  INVX1_HVT U861 ( .A(n15), .Y(n909) );
  INVX1_HVT U862 ( .A(n857), .Y(n837) );
  INVX1_HVT U863 ( .A(n15), .Y(n911) );
  INVX1_HVT U864 ( .A(n15), .Y(n910) );
  INVX1_HVT U865 ( .A(n859), .Y(n848) );
  INVX1_HVT U866 ( .A(n859), .Y(n852) );
  INVX1_HVT U867 ( .A(n859), .Y(n851) );
  INVX1_HVT U868 ( .A(n859), .Y(n850) );
  INVX1_HVT U869 ( .A(n859), .Y(n849) );
  INVX1_HVT U870 ( .A(n858), .Y(n847) );
  INVX1_HVT U871 ( .A(n858), .Y(n846) );
  INVX1_HVT U872 ( .A(n858), .Y(n845) );
  INVX1_HVT U873 ( .A(n858), .Y(n844) );
  INVX1_HVT U874 ( .A(n858), .Y(n843) );
  INVX1_HVT U875 ( .A(n859), .Y(n853) );
  INVX1_HVT U876 ( .A(n860), .Y(n854) );
  INVX1_HVT U877 ( .A(n860), .Y(n855) );
  INVX1_HVT U878 ( .A(n858), .Y(n856) );
  INVX1_HVT U879 ( .A(n17), .Y(n857) );
  NAND2X0_HVT U880 ( .A1(n857), .A2(n18), .Y(n836) );
  INVX0_HVT U881 ( .A(n12), .Y(n913) );
  INVX0_HVT U882 ( .A(n14), .Y(n914) );
  INVX0_HVT U883 ( .A(reset), .Y(n915) );
endmodule

