
module sbox_12 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n210, n211, n212, n213, n216, n217, n218, n219, n224, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588;

  NAND2X0_HVT U4 ( .A1(n294), .A2(n586), .Y(n585) );
  NAND2X0_HVT U5 ( .A1(n302), .A2(n284), .Y(n583) );
  NAND2X0_HVT U13 ( .A1(n575), .A2(n298), .Y(n576) );
  NAND2X0_HVT U15 ( .A1(n586), .A2(n285), .Y(n573) );
  NAND2X0_HVT U21 ( .A1(n294), .A2(n305), .Y(n567) );
  NAND2X0_HVT U24 ( .A1(n289), .A2(n305), .Y(n565) );
  NAND2X0_HVT U33 ( .A1(n363), .A2(n305), .Y(n556) );
  NAND2X0_HVT U35 ( .A1(n288), .A2(n305), .Y(n554) );
  NAND2X0_HVT U42 ( .A1(n210), .A2(n289), .Y(n547) );
  MUX41X1_HVT U51 ( .A1(n352), .A3(n312), .A2(n330), .A4(n331), .S0(n256), 
        .S1(n308), .Y(n538) );
  NAND2X0_HVT U53 ( .A1(n535), .A2(n546), .Y(n536) );
  NAND2X0_HVT U56 ( .A1(n294), .A2(n531), .Y(n532) );
  MUX41X1_HVT U57 ( .A1(n353), .A3(n569), .A2(n532), .A4(n578), .S0(n283), 
        .S1(n308), .Y(n530) );
  NAND2X0_HVT U58 ( .A1(n298), .A2(n586), .Y(n529) );
  MUX41X1_HVT U59 ( .A1(n274), .A3(n529), .A2(n272), .A4(n329), .S0(n256), 
        .S1(n308), .Y(n528) );
  MUX41X1_HVT U61 ( .A1(n270), .A3(n328), .A2(n327), .A4(n285), .S0(n256), 
        .S1(n279), .Y(n526) );
  NAND2X0_HVT U62 ( .A1(n305), .A2(n296), .Y(n525) );
  MUX41X1_HVT U63 ( .A1(n525), .A3(n319), .A2(n347), .A4(n326), .S0(n256), 
        .S1(n308), .Y(n524) );
  AO21X1_HVT U66 ( .A1(n324), .A2(n280), .A3(n346), .Y(n521) );
  MUX41X1_HVT U68 ( .A1(n322), .A3(n521), .A2(n520), .A4(n522), .S0(n275), 
        .S1(n310), .Y(n519) );
  MUX41X1_HVT U69 ( .A1(n519), .A3(n527), .A2(n523), .A4(n533), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n291), .A2(n514), .Y(n515) );
  MUX41X1_HVT U74 ( .A1(n516), .A3(n563), .A2(n515), .A4(n565), .S0(n275), 
        .S1(n259), .Y(n513) );
  MUX41X1_HVT U75 ( .A1(n350), .A3(n355), .A2(n367), .A4(n333), .S0(n275), 
        .S1(n259), .Y(n512) );
  MUX41X1_HVT U82 ( .A1(n544), .A3(n331), .A2(n313), .A4(n574), .S0(n275), 
        .S1(n309), .Y(n504) );
  AND2X1_HVT U83 ( .A1(n303), .A2(n216), .Y(n503) );
  NAND2X0_HVT U85 ( .A1(n305), .A2(n366), .Y(n501) );
  MUX41X1_HVT U90 ( .A1(n543), .A3(n547), .A2(n352), .A4(n498), .S0(n276), 
        .S1(n309), .Y(n497) );
  AO21X1_HVT U93 ( .A1(n282), .A2(n493), .A3(n351), .Y(n494) );
  MUX41X1_HVT U96 ( .A1(n313), .A3(n269), .A2(n354), .A4(n491), .S0(n275), 
        .S1(n309), .Y(n490) );
  MUX41X1_HVT U97 ( .A1(n350), .A3(n269), .A2(n300), .A4(n573), .S0(n275), 
        .S1(n309), .Y(n489) );
  MUX41X1_HVT U98 ( .A1(n489), .A3(n492), .A2(n490), .A4(n497), .S0(in[0]), 
        .S1(n308), .Y(n488) );
  NAND2X0_HVT U101 ( .A1(n484), .A2(n483), .Y(n485) );
  MUX41X1_HVT U103 ( .A1(n586), .A3(n323), .A2(n242), .A4(n554), .S0(n275), 
        .S1(n309), .Y(n481) );
  MUX41X1_HVT U105 ( .A1(n335), .A3(n541), .A2(n480), .A4(n349), .S0(n275), 
        .S1(n309), .Y(n479) );
  MUX41X1_HVT U106 ( .A1(n479), .A3(n482), .A2(n481), .A4(n486), .S0(in[0]), 
        .S1(n308), .Y(n478) );
  OA21X1_HVT U109 ( .A1(n252), .A2(n307), .A3(n329), .Y(n476) );
  NAND2X0_HVT U110 ( .A1(n295), .A2(n474), .Y(n475) );
  AND2X1_HVT U115 ( .A1(n301), .A2(n285), .Y(n469) );
  MUX41X1_HVT U116 ( .A1(n576), .A3(n469), .A2(n333), .A4(n558), .S0(n276), 
        .S1(n283), .Y(n468) );
  NAND2X0_HVT U123 ( .A1(n460), .A2(n459), .Y(n461) );
  MUX41X1_HVT U125 ( .A1(n567), .A3(n274), .A2(n322), .A4(n358), .S0(n276), 
        .S1(n259), .Y(n457) );
  MUX41X1_HVT U135 ( .A1(n359), .A3(n364), .A2(n583), .A4(n562), .S0(n247), 
        .S1(n256), .Y(n448) );
  MUX41X1_HVT U136 ( .A1(n267), .A3(n556), .A2(n360), .A4(n553), .S0(n276), 
        .S1(n256), .Y(n447) );
  MUX41X1_HVT U139 ( .A1(n445), .A3(n448), .A2(n447), .A4(n449), .S0(in[0]), 
        .S1(n279), .Y(n444) );
  AND2X1_HVT U140 ( .A1(n290), .A2(n304), .Y(n443) );
  MUX41X1_HVT U141 ( .A1(n564), .A3(n341), .A2(n443), .A4(n338), .S0(n278), 
        .S1(n256), .Y(n442) );
  MUX41X1_HVT U142 ( .A1(n332), .A3(n286), .A2(n348), .A4(n290), .S0(n276), 
        .S1(n256), .Y(n441) );
  NAND2X0_HVT U146 ( .A1(n210), .A2(n298), .Y(n514) );
  OA21X1_HVT U151 ( .A1(n549), .A2(n232), .A3(n433), .Y(n434) );
  MUX41X1_HVT U153 ( .A1(n475), .A3(n270), .A2(n587), .A4(n315), .S0(n276), 
        .S1(n310), .Y(n431) );
  AND2X1_HVT U154 ( .A1(n282), .A2(n289), .Y(n430) );
  NAND2X0_HVT U158 ( .A1(n299), .A2(n366), .Y(n426) );
  MUX41X1_HVT U159 ( .A1(n254), .A3(n286), .A2(n426), .A4(n321), .S0(n244), 
        .S1(n310), .Y(n425) );
  AND2X1_HVT U162 ( .A1(n582), .A2(n514), .Y(n422) );
  MUX41X1_HVT U163 ( .A1(n328), .A3(n422), .A2(n268), .A4(n423), .S0(n306), 
        .S1(n309), .Y(n421) );
  NAND2X0_HVT U166 ( .A1(n298), .A2(n531), .Y(n418) );
  NAND2X0_HVT U167 ( .A1(n367), .A2(n305), .Y(n417) );
  MUX41X1_HVT U168 ( .A1(n353), .A3(n290), .A2(n417), .A4(n418), .S0(n247), 
        .S1(n283), .Y(n416) );
  NAND2X0_HVT U174 ( .A1(n303), .A2(n582), .Y(n575) );
  MUX41X1_HVT U176 ( .A1(n368), .A3(n411), .A2(n357), .A4(n212), .S0(n282), 
        .S1(n306), .Y(n410) );
  NAND2X0_HVT U177 ( .A1(n210), .A2(n287), .Y(n409) );
  MUX41X1_HVT U178 ( .A1(n571), .A3(n409), .A2(n361), .A4(n551), .S0(n244), 
        .S1(n259), .Y(n408) );
  MUX41X1_HVT U179 ( .A1(n561), .A3(n362), .A2(n317), .A4(n361), .S0(n306), 
        .S1(n310), .Y(n407) );
  MUX41X1_HVT U180 ( .A1(n320), .A3(n580), .A2(n254), .A4(n266), .S0(n282), 
        .S1(n247), .Y(n406) );
  MUX41X1_HVT U181 ( .A1(n406), .A3(n408), .A2(n407), .A4(n410), .S0(in[0]), 
        .S1(n279), .Y(n405) );
  OA21X1_HVT U184 ( .A1(n555), .A2(n261), .A3(n332), .Y(n402) );
  MUX41X1_HVT U189 ( .A1(n398), .A3(n212), .A2(n399), .A4(n349), .S0(n282), 
        .S1(n244), .Y(n397) );
  MUX41X1_HVT U193 ( .A1(n547), .A3(n554), .A2(n539), .A4(n395), .S0(n247), 
        .S1(n309), .Y(n394) );
  MUX41X1_HVT U195 ( .A1(n582), .A3(n354), .A2(n297), .A4(n552), .S0(n306), 
        .S1(n310), .Y(n392) );
  AO21X1_HVT U197 ( .A1(n271), .A2(n283), .A3(n351), .Y(n390) );
  OA21X1_HVT U201 ( .A1(n581), .A2(n232), .A3(n341), .Y(n386) );
  MUX41X1_HVT U203 ( .A1(n553), .A3(n343), .A2(n577), .A4(n557), .S0(n306), 
        .S1(n309), .Y(n384) );
  MUX41X1_HVT U205 ( .A1(in[4]), .A3(n586), .A2(n362), .A4(n218), .S0(n244), 
        .S1(n310), .Y(n382) );
  NAND2X0_HVT U208 ( .A1(n302), .A2(n294), .Y(n474) );
  NAND2X0_HVT U212 ( .A1(n301), .A2(n291), .Y(n531) );
  NAND2X0_HVT U214 ( .A1(n582), .A2(n305), .Y(n380) );
  NAND2X0_HVT U215 ( .A1(n474), .A2(n292), .Y(n379) );
  AO21X1_HVT U216 ( .A1(n304), .A2(n364), .A3(n232), .Y(n484) );
  NAND2X0_HVT U218 ( .A1(n364), .A2(n300), .Y(n433) );
  NAND2X0_HVT U220 ( .A1(n281), .A2(n380), .Y(n506) );
  INVX2_HVT U1 ( .A(n311), .Y(n310) );
  INVX4_HVT U2 ( .A(n311), .Y(n309) );
  INVX0_HVT U3 ( .A(n304), .Y(n302) );
  INVX1_HVT U6 ( .A(n304), .Y(n300) );
  INVX0_HVT U7 ( .A(n294), .Y(n253) );
  INVX0_HVT U8 ( .A(n297), .Y(n219) );
  INVX0_HVT U9 ( .A(n291), .Y(n224) );
  XOR2X1_HVT U10 ( .A1(n582), .A2(n299), .Y(n543) );
  XOR2X1_HVT U11 ( .A1(n232), .A2(n562), .Y(n545) );
  INVX0_HVT U12 ( .A(n213), .Y(n511) );
  NAND2X0_HVT U14 ( .A1(n386), .A2(n231), .Y(n250) );
  MUX21X1_HVT U16 ( .A1(n314), .A2(n463), .S0(n278), .Y(n462) );
  INVX0_HVT U17 ( .A(n252), .Y(n552) );
  MUX21X1_HVT U18 ( .A1(n218), .A2(n574), .S0(n278), .Y(n487) );
  INVX1_HVT U19 ( .A(n568), .Y(n331) );
  NBUFFX2_HVT U20 ( .A(in[5]), .Y(n280) );
  NAND2X0_HVT U22 ( .A1(n300), .A2(n295), .Y(n586) );
  OA21X1_HVT U23 ( .A1(n272), .A2(n232), .A3(n558), .Y(n414) );
  INVX1_HVT U25 ( .A(n306), .Y(n231) );
  INVX0_HVT U26 ( .A(in[6]), .Y(n262) );
  INVX1_HVT U27 ( .A(in[4]), .Y(n368) );
  INVX0_HVT U28 ( .A(n261), .Y(n259) );
  INVX0_HVT U29 ( .A(n283), .Y(n261) );
  INVX0_HVT U30 ( .A(n281), .Y(n232) );
  INVX1_HVT U31 ( .A(in[0]), .Y(n257) );
  INVX0_HVT U32 ( .A(n288), .Y(n216) );
  INVX1_HVT U34 ( .A(n279), .Y(n243) );
  INVX1_HVT U36 ( .A(n255), .Y(n244) );
  INVX1_HVT U37 ( .A(n278), .Y(n255) );
  INVX1_HVT U38 ( .A(in[2]), .Y(n307) );
  INVX0_HVT U39 ( .A(n255), .Y(n247) );
  INVX1_HVT U40 ( .A(in[7]), .Y(n311) );
  MUX41X1_HVT U41 ( .A1(n355), .A3(n271), .A2(n501), .A4(n267), .S0(n310), 
        .S1(n275), .Y(n500) );
  MUX41X1_HVT U43 ( .A1(n332), .A3(n572), .A2(n582), .A4(n503), .S0(n309), 
        .S1(n275), .Y(n502) );
  INVX1_HVT U44 ( .A(n566), .Y(n332) );
  INVX1_HVT U45 ( .A(n260), .Y(n582) );
  IBUFFX2_HVT U46 ( .A(n304), .Y(n23) );
  INVX1_HVT U47 ( .A(n304), .Y(n210) );
  NAND2X0_HVT U48 ( .A1(n235), .A2(n236), .Y(out[4]) );
  IBUFFX2_HVT U49 ( .A(n304), .Y(n301) );
  MUX41X1_HVT U50 ( .A1(n394), .A3(n392), .A2(n393), .A4(n389), .S0(n257), 
        .S1(n243), .Y(n388) );
  MUX21X2_HVT U52 ( .A1(n560), .A2(n318), .S0(n281), .Y(n440) );
  AO21X2_HVT U54 ( .A1(n278), .A2(n290), .A3(n582), .Y(n466) );
  INVX0_HVT U55 ( .A(n299), .Y(n217) );
  INVX0_HVT U60 ( .A(n304), .Y(n299) );
  INVX0_HVT U64 ( .A(n575), .Y(n211) );
  INVX1_HVT U65 ( .A(n211), .Y(n212) );
  MUX21X2_HVT U67 ( .A1(n526), .A2(n524), .S0(n231), .Y(n523) );
  MUX41X1_HVT U70 ( .A1(n421), .A3(n416), .A2(n419), .A4(n413), .S0(n257), 
        .S1(n243), .Y(n412) );
  INVX0_HVT U71 ( .A(n576), .Y(n347) );
  INVX0_HVT U72 ( .A(n347), .Y(n254) );
  MUX21X1_HVT U76 ( .A1(n216), .A2(n260), .S0(n217), .Y(n213) );
  MUX21X2_HVT U77 ( .A1(n405), .A2(n396), .S0(n262), .Y(out[6]) );
  IBUFFX2_HVT U78 ( .A(n304), .Y(n303) );
  MUX21X2_HVT U79 ( .A1(n462), .A2(n461), .S0(n282), .Y(n458) );
  OA21X1_HVT U80 ( .A1(n316), .A2(n261), .A3(n558), .Y(n439) );
  IBUFFX2_HVT U81 ( .A(n218), .Y(n558) );
  INVX1_HVT U84 ( .A(n242), .Y(n560) );
  MUX21X2_HVT U86 ( .A1(n270), .A2(n487), .S0(n542), .Y(n486) );
  MUX21X1_HVT U87 ( .A1(n219), .A2(n224), .S0(n303), .Y(n218) );
  MUX21X2_HVT U88 ( .A1(n518), .A2(n545), .S0(n231), .Y(n517) );
  IBUFFX2_HVT U89 ( .A(in[1]), .Y(n305) );
  MUX21X1_HVT U91 ( .A1(n367), .A2(n366), .S0(n210), .Y(n562) );
  IBUFFX2_HVT U92 ( .A(n580), .Y(n323) );
  INVX1_HVT U94 ( .A(n239), .Y(n518) );
  MUX41X1_HVT U95 ( .A1(n258), .A3(n511), .A2(n356), .A4(n580), .S0(n261), 
        .S1(n231), .Y(n510) );
  INVX1_HVT U99 ( .A(n376), .Y(n354) );
  MUX21X1_HVT U100 ( .A1(n364), .A2(n258), .S0(n232), .Y(n435) );
  MUX41X1_HVT U102 ( .A1(n432), .A3(n427), .A2(n431), .A4(n425), .S0(n257), 
        .S1(n243), .Y(n424) );
  NAND2X0_HVT U104 ( .A1(n507), .A2(n247), .Y(n233) );
  NAND2X0_HVT U107 ( .A1(n508), .A2(n231), .Y(n234) );
  NAND2X0_HVT U108 ( .A1(n233), .A2(n234), .Y(n505) );
  AND3X2_HVT U111 ( .A1(n295), .A2(n531), .A3(n506), .Y(n507) );
  MUX21X1_HVT U112 ( .A1(n568), .A2(n292), .S0(n281), .Y(n508) );
  IBUFFX2_HVT U113 ( .A(n311), .Y(n256) );
  MUX41X1_HVT U114 ( .A1(n543), .A3(n514), .A2(n350), .A4(n360), .S0(n261), 
        .S1(n255), .Y(n437) );
  NAND2X0_HVT U117 ( .A1(n444), .A2(in[6]), .Y(n235) );
  NAND2X0_HVT U118 ( .A1(n436), .A2(n262), .Y(n236) );
  NAND2X0_HVT U119 ( .A1(n450), .A2(n244), .Y(n237) );
  NAND2X0_HVT U120 ( .A1(n337), .A2(n255), .Y(n238) );
  NAND2X0_HVT U121 ( .A1(n237), .A2(n238), .Y(n449) );
  MUX21X2_HVT U122 ( .A1(n434), .A2(n435), .S0(n244), .Y(n432) );
  MUX21X2_HVT U124 ( .A1(n457), .A2(n458), .S0(n280), .Y(n456) );
  MUX21X2_HVT U126 ( .A1(n465), .A2(n468), .S0(n280), .Y(n464) );
  MUX21X1_HVT U127 ( .A1(n297), .A2(n376), .S0(n281), .Y(n239) );
  MUX41X1_HVT U128 ( .A1(n517), .A3(n512), .A2(n513), .A4(n510), .S0(n257), 
        .S1(n243), .Y(n509) );
  NAND2X0_HVT U129 ( .A1(n388), .A2(in[6]), .Y(n240) );
  NAND2X0_HVT U130 ( .A1(n381), .A2(n262), .Y(n241) );
  NAND2X0_HVT U131 ( .A1(n240), .A2(n241), .Y(out[7]) );
  MUX21X1_HVT U132 ( .A1(n216), .A2(n293), .S0(n303), .Y(n242) );
  MUX41X1_HVT U133 ( .A1(n505), .A3(n502), .A2(n504), .A4(n500), .S0(n257), 
        .S1(n243), .Y(n499) );
  MUX21X2_HVT U134 ( .A1(n439), .A2(n440), .S0(n255), .Y(n438) );
  INVX1_HVT U137 ( .A(n374), .Y(n337) );
  MUX21X2_HVT U138 ( .A1(n412), .A2(n424), .S0(in[6]), .Y(out[5]) );
  MUX21X2_HVT U143 ( .A1(n494), .A2(n495), .S0(n278), .Y(n492) );
  NAND2X0_HVT U144 ( .A1(n585), .A2(n244), .Y(n245) );
  NAND2X0_HVT U145 ( .A1(n446), .A2(n307), .Y(n246) );
  NAND2X0_HVT U147 ( .A1(n246), .A2(n245), .Y(n445) );
  NAND2X0_HVT U148 ( .A1(n429), .A2(n247), .Y(n248) );
  NAND2X0_HVT U149 ( .A1(n428), .A2(n255), .Y(n249) );
  NAND2X0_HVT U150 ( .A1(n248), .A2(n249), .Y(n427) );
  MUX21X2_HVT U152 ( .A1(n296), .A2(n496), .S0(n273), .Y(n495) );
  NAND2X0_HVT U155 ( .A1(n387), .A2(n277), .Y(n251) );
  NAND2X0_HVT U156 ( .A1(n250), .A2(n251), .Y(n385) );
  INVX2_HVT U157 ( .A(in[1]), .Y(n304) );
  MUX21X1_HVT U160 ( .A1(n253), .A2(n260), .S0(n302), .Y(n252) );
  MUX41X1_HVT U161 ( .A1(n576), .A3(n532), .A2(n566), .A4(n339), .S0(n231), 
        .S1(n310), .Y(n383) );
  MUX41X1_HVT U164 ( .A1(n567), .A3(n336), .A2(n543), .A4(n420), .S0(n256), 
        .S1(in[2]), .Y(n419) );
  MUX41X1_HVT U165 ( .A1(n385), .A3(n383), .A2(n384), .A4(n382), .S0(n257), 
        .S1(n243), .Y(n381) );
  MUX41X1_HVT U169 ( .A1(n550), .A3(n269), .A2(n543), .A4(n514), .S0(n255), 
        .S1(n310), .Y(n400) );
  AND3X2_HVT U170 ( .A1(n278), .A2(n305), .A3(in[4]), .Y(n454) );
  MUX21X1_HVT U171 ( .A1(n285), .A2(n284), .S0(n300), .Y(n572) );
  MUX21X1_HVT U172 ( .A1(n289), .A2(n260), .S0(n300), .Y(n258) );
  MUX21X1_HVT U173 ( .A1(n572), .A2(n266), .S0(n282), .Y(n387) );
  XNOR2X2_HVT U175 ( .A1(n368), .A2(in[3]), .Y(n260) );
  IBUFFX2_HVT U182 ( .A(n572), .Y(n327) );
  MUX41X1_HVT U183 ( .A1(n334), .A3(n344), .A2(n293), .A4(n342), .S0(n261), 
        .S1(n307), .Y(n404) );
  MUX21X2_HVT U185 ( .A1(n499), .A2(n509), .S0(in[6]), .Y(out[1]) );
  MUX41X1_HVT U186 ( .A1(n441), .A3(n437), .A2(n442), .A4(n438), .S0(n257), 
        .S1(n308), .Y(n436) );
  MUX41X1_HVT U187 ( .A1(n452), .A3(n454), .A2(n453), .A4(n455), .S0(n280), 
        .S1(n283), .Y(n451) );
  MUX41X1_HVT U188 ( .A1(n290), .A3(n359), .A2(n562), .A4(n548), .S0(n261), 
        .S1(n307), .Y(n393) );
  MUX41X1_HVT U190 ( .A1(n401), .A3(n404), .A2(n397), .A4(n400), .S0(n279), 
        .S1(n257), .Y(n396) );
  XOR2X1_HVT U191 ( .A1(n305), .A2(n307), .Y(n540) );
  MUX41X1_HVT U192 ( .A1(n456), .A3(n451), .A2(n470), .A4(n464), .S0(n257), 
        .S1(in[6]), .Y(out[3]) );
  XOR2X1_HVT U194 ( .A1(n307), .A2(n232), .Y(n542) );
  MUX21X2_HVT U196 ( .A1(n478), .A2(n488), .S0(in[6]), .Y(out[2]) );
  MUX41X1_HVT U198 ( .A1(n471), .A3(n473), .A2(n477), .A4(n476), .S0(n310), 
        .S1(n280), .Y(n470) );
  NAND2X0_HVT U199 ( .A1(n472), .A2(n263), .Y(n264) );
  NAND2X0_HVT U200 ( .A1(n296), .A2(n540), .Y(n265) );
  NAND2X0_HVT U202 ( .A1(n264), .A2(n265), .Y(n471) );
  INVX0_HVT U204 ( .A(n540), .Y(n263) );
  INVX0_HVT U206 ( .A(in[3]), .Y(n365) );
  INVX1_HVT U207 ( .A(n293), .Y(n363) );
  MUX21X1_HVT U209 ( .A1(n268), .A2(n327), .S0(n276), .Y(n453) );
  NBUFFX2_HVT U210 ( .A(n260), .Y(n285) );
  NBUFFX2_HVT U211 ( .A(n260), .Y(n286) );
  AND2X1_HVT U213 ( .A1(n286), .A2(n531), .Y(n266) );
  NBUFFX2_HVT U217 ( .A(n584), .Y(n293) );
  INVX1_HVT U219 ( .A(n587), .Y(n367) );
  MUX21X1_HVT U221 ( .A1(n363), .A2(n366), .S0(n280), .Y(n535) );
  NBUFFX2_HVT U222 ( .A(n584), .Y(n294) );
  MUX21X1_HVT U223 ( .A1(n558), .A2(n475), .S0(n276), .Y(n473) );
  MUX21X1_HVT U224 ( .A1(n323), .A2(n364), .S0(n280), .Y(n520) );
  AND2X1_HVT U225 ( .A1(n295), .A2(n514), .Y(n267) );
  MUX21X1_HVT U226 ( .A1(n286), .A2(n366), .S0(n301), .Y(n581) );
  MUX21X1_HVT U227 ( .A1(n295), .A2(n285), .S0(n210), .Y(n548) );
  MUX21X1_HVT U228 ( .A1(n285), .A2(n288), .S0(n302), .Y(n483) );
  MUX21X1_HVT U229 ( .A1(n566), .A2(n342), .S0(n282), .Y(n446) );
  MUX21X1_HVT U230 ( .A1(n363), .A2(n367), .S0(n302), .Y(n411) );
  MUX21X1_HVT U231 ( .A1(n366), .A2(n285), .S0(n299), .Y(n423) );
  MUX21X1_HVT U232 ( .A1(n285), .A2(n363), .S0(n303), .Y(n491) );
  MUX21X1_HVT U233 ( .A1(n582), .A2(n364), .S0(n301), .Y(n372) );
  MUX21X1_HVT U234 ( .A1(n582), .A2(n367), .S0(n299), .Y(n564) );
  MUX21X1_HVT U235 ( .A1(n294), .A2(n292), .S0(n23), .Y(n498) );
  MUX21X1_HVT U236 ( .A1(n366), .A2(n363), .S0(n210), .Y(n551) );
  MUX21X1_HVT U237 ( .A1(n366), .A2(n284), .S0(n300), .Y(n555) );
  MUX21X1_HVT U238 ( .A1(n284), .A2(n367), .S0(n23), .Y(n549) );
  MUX21X1_HVT U239 ( .A1(n358), .A2(n292), .S0(n282), .Y(n450) );
  MUX21X1_HVT U240 ( .A1(n466), .A2(n467), .S0(n283), .Y(n465) );
  MUX21X1_HVT U241 ( .A1(n315), .A2(n339), .S0(n276), .Y(n467) );
  NAND2X0_HVT U242 ( .A1(n287), .A2(n365), .Y(n584) );
  MUX21X1_HVT U243 ( .A1(n363), .A2(n287), .S0(n210), .Y(n373) );
  INVX1_HVT U244 ( .A(n297), .Y(n366) );
  MUX21X1_HVT U245 ( .A1(n287), .A2(n284), .S0(n23), .Y(n463) );
  NBUFFX2_HVT U246 ( .A(n587), .Y(n295) );
  XOR2X1_HVT U247 ( .A1(n300), .A2(n364), .Y(n544) );
  MUX21X1_HVT U248 ( .A1(n284), .A2(n298), .S0(n301), .Y(n398) );
  MUX21X1_HVT U249 ( .A1(n297), .A2(n295), .S0(n210), .Y(n399) );
  MUX21X1_HVT U250 ( .A1(n364), .A2(n363), .S0(n303), .Y(n570) );
  INVX1_HVT U251 ( .A(n290), .Y(n364) );
  MUX21X1_HVT U252 ( .A1(n296), .A2(n291), .S0(n301), .Y(n574) );
  MUX21X1_HVT U253 ( .A1(n293), .A2(n298), .S0(n301), .Y(n493) );
  MUX21X1_HVT U254 ( .A1(n284), .A2(n366), .S0(n301), .Y(n578) );
  NBUFFX2_HVT U255 ( .A(n587), .Y(n296) );
  MUX21X1_HVT U256 ( .A1(n284), .A2(n288), .S0(n210), .Y(n395) );
  XOR2X1_HVT U257 ( .A1(n296), .A2(n210), .Y(n539) );
  MUX21X1_HVT U258 ( .A1(n296), .A2(n287), .S0(n301), .Y(n378) );
  XNOR2X1_HVT U259 ( .A1(n293), .A2(n23), .Y(n268) );
  AND2X1_HVT U260 ( .A1(n23), .A2(n367), .Y(n269) );
  MUX21X1_HVT U261 ( .A1(n294), .A2(n284), .S0(n23), .Y(n577) );
  MUX21X1_HVT U262 ( .A1(n296), .A2(n294), .S0(n300), .Y(n371) );
  AND2X1_HVT U263 ( .A1(n298), .A2(n474), .Y(n270) );
  XNOR2X1_HVT U264 ( .A1(n297), .A2(n299), .Y(n271) );
  MUX21X1_HVT U265 ( .A1(n291), .A2(n284), .S0(n302), .Y(n376) );
  MUX21X1_HVT U266 ( .A1(n292), .A2(n287), .S0(n23), .Y(n516) );
  MUX21X1_HVT U267 ( .A1(n292), .A2(n298), .S0(n278), .Y(n460) );
  XOR2X1_HVT U268 ( .A1(n287), .A2(n300), .Y(n563) );
  NBUFFX2_HVT U269 ( .A(in[7]), .Y(n283) );
  NBUFFX2_HVT U270 ( .A(in[7]), .Y(n281) );
  NBUFFX2_HVT U271 ( .A(in[7]), .Y(n282) );
  NBUFFX2_HVT U272 ( .A(n365), .Y(n284) );
  NBUFFX2_HVT U273 ( .A(in[2]), .Y(n276) );
  NBUFFX2_HVT U274 ( .A(in[5]), .Y(n279) );
  NBUFFX2_HVT U275 ( .A(in[2]), .Y(n278) );
  NBUFFX2_HVT U276 ( .A(n306), .Y(n277) );
  NBUFFX2_HVT U277 ( .A(in[2]), .Y(n275) );
  MUX21X1_HVT U278 ( .A1(n286), .A2(n289), .S0(n299), .Y(n566) );
  MUX21X1_HVT U279 ( .A1(n485), .A2(n337), .S0(n244), .Y(n482) );
  MUX21X1_HVT U280 ( .A1(n402), .A2(n403), .S0(n277), .Y(n401) );
  MUX21X1_HVT U281 ( .A1(n501), .A2(n289), .S0(n281), .Y(n403) );
  XOR2X1_HVT U282 ( .A1(n299), .A2(n289), .Y(n541) );
  MUX21X1_HVT U283 ( .A1(n291), .A2(n286), .S0(n299), .Y(n480) );
  MUX21X1_HVT U284 ( .A1(n415), .A2(n414), .S0(n278), .Y(n413) );
  MUX21X1_HVT U285 ( .A1(n292), .A2(n354), .S0(n281), .Y(n415) );
  AND2X1_HVT U286 ( .A1(n286), .A2(n305), .Y(n272) );
  MUX21X1_HVT U287 ( .A1(n289), .A2(n363), .S0(n302), .Y(n550) );
  MUX21X1_HVT U288 ( .A1(n364), .A2(n367), .S0(n303), .Y(n420) );
  NAND2X0_HVT U289 ( .A1(in[3]), .A2(n288), .Y(n587) );
  NBUFFX2_HVT U290 ( .A(n368), .Y(n288) );
  NBUFFX2_HVT U291 ( .A(n588), .Y(n297) );
  MUX21X1_HVT U292 ( .A1(n367), .A2(n289), .S0(n301), .Y(n569) );
  MUX21X1_HVT U293 ( .A1(n340), .A2(n586), .S0(n276), .Y(n477) );
  MUX21X1_HVT U294 ( .A1(n430), .A2(n296), .S0(n273), .Y(n429) );
  MUX21X1_HVT U295 ( .A1(n551), .A2(n356), .S0(n283), .Y(n428) );
  MUX21X1_HVT U296 ( .A1(n571), .A2(n338), .S0(n278), .Y(n452) );
  MUX21X1_HVT U297 ( .A1(n536), .A2(n537), .S0(n283), .Y(n534) );
  MUX21X1_HVT U298 ( .A1(n289), .A2(n554), .S0(n280), .Y(n537) );
  XOR2X1_HVT U299 ( .A1(n23), .A2(n279), .Y(n546) );
  MUX21X1_HVT U300 ( .A1(n586), .A2(n304), .S0(n277), .Y(n459) );
  NBUFFX2_HVT U301 ( .A(n579), .Y(n290) );
  MUX21X1_HVT U302 ( .A1(n289), .A2(n364), .S0(n23), .Y(n375) );
  MUX21X1_HVT U303 ( .A1(n559), .A2(n379), .S0(n282), .Y(n374) );
  MUX21X1_HVT U304 ( .A1(n294), .A2(n289), .S0(n302), .Y(n580) );
  MUX21X1_HVT U305 ( .A1(n325), .A2(n305), .S0(n280), .Y(n522) );
  NBUFFX2_HVT U306 ( .A(n579), .Y(n291) );
  MUX21X1_HVT U307 ( .A1(n335), .A2(n559), .S0(n275), .Y(n455) );
  MUX21X1_HVT U308 ( .A1(n345), .A2(n361), .S0(n281), .Y(n391) );
  MUX21X1_HVT U309 ( .A1(n289), .A2(n287), .S0(n281), .Y(n496) );
  NBUFFX2_HVT U310 ( .A(n588), .Y(n298) );
  NBUFFX2_HVT U311 ( .A(n368), .Y(n287) );
  NBUFFX2_HVT U312 ( .A(n579), .Y(n292) );
  XNOR2X1_HVT U313 ( .A1(n232), .A2(n23), .Y(n273) );
  AND2X1_HVT U314 ( .A1(n284), .A2(n305), .Y(n274) );
  INVX1_HVT U315 ( .A(n307), .Y(n306) );
  NBUFFX2_HVT U316 ( .A(in[5]), .Y(n308) );
  MUX21X1_HVT U317 ( .A1(n391), .A2(n390), .S0(n277), .Y(n389) );
  MUX21X1_HVT U318 ( .A1(n534), .A2(n538), .S0(n247), .Y(n533) );
  MUX21X1_HVT U319 ( .A1(n528), .A2(n530), .S0(n277), .Y(n527) );
  MUX21X1_HVT U320 ( .A1(n363), .A2(n216), .S0(n299), .Y(n557) );
  NAND2X0_HVT U321 ( .A1(in[3]), .A2(in[4]), .Y(n588) );
  MUX21X1_HVT U322 ( .A1(n216), .A2(n582), .S0(n303), .Y(n377) );
  MUX21X1_HVT U323 ( .A1(n216), .A2(n366), .S0(n302), .Y(n553) );
  MUX21X1_HVT U324 ( .A1(n216), .A2(n364), .S0(n302), .Y(n571) );
  NAND2X0_HVT U325 ( .A1(in[4]), .A2(n365), .Y(n579) );
  MUX21X1_HVT U326 ( .A1(n216), .A2(n296), .S0(n303), .Y(n568) );
  MUX21X1_HVT U327 ( .A1(n298), .A2(n216), .S0(n300), .Y(n561) );
  MUX21X1_HVT U328 ( .A1(n289), .A2(n216), .S0(n276), .Y(n472) );
  MUX21X1_HVT U329 ( .A1(n216), .A2(n291), .S0(n300), .Y(n370) );
  MUX21X1_HVT U330 ( .A1(n216), .A2(n298), .S0(n303), .Y(n369) );
  MUX21X1_HVT U331 ( .A1(n284), .A2(n216), .S0(n210), .Y(n559) );
  NBUFFX2_HVT U332 ( .A(in[3]), .Y(n289) );
  INVX0_HVT U333 ( .A(n567), .Y(n312) );
  INVX0_HVT U334 ( .A(n565), .Y(n313) );
  INVX0_HVT U335 ( .A(n556), .Y(n314) );
  INVX0_HVT U336 ( .A(n554), .Y(n315) );
  INVX0_HVT U337 ( .A(n417), .Y(n316) );
  INVX0_HVT U338 ( .A(n380), .Y(n317) );
  INVX0_HVT U339 ( .A(n586), .Y(n318) );
  INVX0_HVT U340 ( .A(n573), .Y(n319) );
  INVX0_HVT U341 ( .A(n585), .Y(n320) );
  INVX0_HVT U342 ( .A(n583), .Y(n321) );
  INVX0_HVT U343 ( .A(n581), .Y(n322) );
  INVX0_HVT U344 ( .A(n578), .Y(n324) );
  INVX0_HVT U345 ( .A(n577), .Y(n325) );
  INVX0_HVT U346 ( .A(n574), .Y(n326) );
  INVX0_HVT U347 ( .A(n571), .Y(n328) );
  INVX0_HVT U348 ( .A(n570), .Y(n329) );
  INVX0_HVT U349 ( .A(n569), .Y(n330) );
  INVX0_HVT U350 ( .A(n564), .Y(n333) );
  INVX0_HVT U351 ( .A(n563), .Y(n334) );
  INVX0_HVT U352 ( .A(n561), .Y(n335) );
  INVX0_HVT U353 ( .A(n559), .Y(n336) );
  INVX0_HVT U354 ( .A(n557), .Y(n338) );
  INVX0_HVT U355 ( .A(n555), .Y(n339) );
  INVX0_HVT U356 ( .A(n553), .Y(n340) );
  INVX0_HVT U357 ( .A(n551), .Y(n341) );
  INVX0_HVT U358 ( .A(n550), .Y(n342) );
  INVX0_HVT U359 ( .A(n549), .Y(n343) );
  INVX0_HVT U360 ( .A(n548), .Y(n344) );
  INVX0_HVT U361 ( .A(n547), .Y(n345) );
  INVX0_HVT U362 ( .A(n514), .Y(n346) );
  INVX0_HVT U363 ( .A(n474), .Y(n348) );
  INVX0_HVT U364 ( .A(n379), .Y(n349) );
  INVX0_HVT U365 ( .A(n531), .Y(n350) );
  INVX0_HVT U366 ( .A(n433), .Y(n351) );
  INVX0_HVT U367 ( .A(n378), .Y(n352) );
  INVX0_HVT U368 ( .A(n377), .Y(n353) );
  INVX0_HVT U369 ( .A(n375), .Y(n355) );
  INVX0_HVT U370 ( .A(n493), .Y(n356) );
  INVX0_HVT U371 ( .A(n483), .Y(n357) );
  INVX0_HVT U372 ( .A(n373), .Y(n358) );
  INVX0_HVT U373 ( .A(n372), .Y(n359) );
  INVX0_HVT U374 ( .A(n371), .Y(n360) );
  INVX0_HVT U375 ( .A(n370), .Y(n361) );
  INVX0_HVT U376 ( .A(n369), .Y(n362) );
endmodule

