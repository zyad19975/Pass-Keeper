
module inv_sbox_9 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n184, n196, n197, n198, n199, n200, n201, n202, n205, n208, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645;

  NAND2X0_HVT U4 ( .A1(n302), .A2(n362), .Y(n642) );
  NAND2X0_HVT U5 ( .A1(n642), .A2(n357), .Y(n641) );
  NAND2X0_HVT U7 ( .A1(n367), .A2(n359), .Y(n638) );
  NAND2X0_HVT U8 ( .A1(n368), .A2(n357), .Y(n637) );
  NAND2X0_HVT U9 ( .A1(n364), .A2(n637), .Y(n636) );
  NAND2X0_HVT U10 ( .A1(n365), .A2(n634), .Y(n635) );
  NAND2X0_HVT U11 ( .A1(n304), .A2(n363), .Y(n633) );
  NAND2X0_HVT U12 ( .A1(n370), .A2(n344), .Y(n632) );
  NAND2X0_HVT U13 ( .A1(n360), .A2(n637), .Y(n631) );
  NAND2X0_HVT U15 ( .A1(n354), .A2(n367), .Y(n629) );
  NAND2X0_HVT U19 ( .A1(n369), .A2(n436), .Y(n624) );
  NAND2X0_HVT U25 ( .A1(n319), .A2(n345), .Y(n640) );
  NAND2X0_HVT U32 ( .A1(n347), .A2(n287), .Y(n612) );
  NAND2X0_HVT U35 ( .A1(n637), .A2(n437), .Y(n609) );
  NAND2X0_HVT U38 ( .A1(n344), .A2(n304), .Y(n606) );
  NAND2X0_HVT U42 ( .A1(n639), .A2(n437), .Y(n602) );
  OA21X1_HVT U53 ( .A1(n378), .A2(n594), .A3(n405), .Y(n592) );
  NAND2X0_HVT U55 ( .A1(n360), .A2(n642), .Y(n590) );
  MUX41X1_HVT U65 ( .A1(n398), .A3(n400), .A2(n399), .A4(n606), .S0(n337), 
        .S1(n376), .Y(n579) );
  NAND2X0_HVT U66 ( .A1(n367), .A2(n331), .Y(n578) );
  MUX41X1_HVT U67 ( .A1(n395), .A3(n419), .A2(n397), .A4(n578), .S0(n341), 
        .S1(n334), .Y(n577) );
  NAND2X0_HVT U72 ( .A1(n355), .A2(n638), .Y(n573) );
  MUX41X1_HVT U73 ( .A1(n617), .A3(n573), .A2(n318), .A4(n344), .S0(n341), 
        .S1(n333), .Y(n572) );
  MUX41X1_HVT U74 ( .A1(n635), .A3(n184), .A2(n409), .A4(n401), .S0(n337), 
        .S1(n376), .Y(n571) );
  MUX41X1_HVT U78 ( .A1(n568), .A3(n572), .A2(n571), .A4(n574), .S0(n352), 
        .S1(n349), .Y(n567) );
  NAND2X0_HVT U81 ( .A1(n363), .A2(n638), .Y(n564) );
  AND2X1_HVT U82 ( .A1(n289), .A2(n358), .Y(n563) );
  MUX41X1_HVT U83 ( .A1(n563), .A3(n407), .A2(n314), .A4(n564), .S0(n336), 
        .S1(n376), .Y(n562) );
  MUX41X1_HVT U84 ( .A1(n329), .A3(n406), .A2(n422), .A4(n619), .S0(n337), 
        .S1(n376), .Y(n561) );
  MUX41X1_HVT U85 ( .A1(n561), .A3(n565), .A2(n562), .A4(n566), .S0(n352), 
        .S1(n349), .Y(n560) );
  MUX41X1_HVT U88 ( .A1(n397), .A3(n382), .A2(n614), .A4(n598), .S0(n336), 
        .S1(n375), .Y(n558) );
  NAND2X0_HVT U89 ( .A1(n286), .A2(n196), .Y(n557) );
  MUX41X1_HVT U90 ( .A1(n435), .A3(n638), .A2(n597), .A4(n557), .S0(n336), 
        .S1(n376), .Y(n556) );
  MUX41X1_HVT U99 ( .A1(n612), .A3(n399), .A2(n596), .A4(n354), .S0(n376), 
        .S1(n334), .Y(n547) );
  NAND2X0_HVT U100 ( .A1(n287), .A2(n432), .Y(n546) );
  MUX41X1_HVT U101 ( .A1(n426), .A3(n632), .A2(n227), .A4(n546), .S0(n376), 
        .S1(n334), .Y(n545) );
  AND2X1_HVT U104 ( .A1(n638), .A2(n356), .Y(n543) );
  MUX41X1_HVT U105 ( .A1(n630), .A3(n427), .A2(n564), .A4(n543), .S0(n337), 
        .S1(n375), .Y(n542) );
  MUX41X1_HVT U107 ( .A1(n426), .A3(n358), .A2(n541), .A4(n388), .S0(n336), 
        .S1(n288), .Y(n540) );
  MUX41X1_HVT U108 ( .A1(n401), .A3(n355), .A2(n269), .A4(n361), .S0(n337), 
        .S1(n312), .Y(n539) );
  MUX41X1_HVT U109 ( .A1(n425), .A3(n382), .A2(n422), .A4(n416), .S0(n336), 
        .S1(n312), .Y(n538) );
  MUX41X1_HVT U110 ( .A1(n538), .A3(n540), .A2(n539), .A4(n542), .S0(in[5]), 
        .S1(n349), .Y(n537) );
  AO21X1_HVT U112 ( .A1(n413), .A2(n341), .A3(n620), .Y(n535) );
  NAND2X0_HVT U114 ( .A1(n365), .A2(n638), .Y(n533) );
  MUX41X1_HVT U115 ( .A1(n533), .A3(n633), .A2(n413), .A4(n358), .S0(n376), 
        .S1(n334), .Y(n532) );
  MUX41X1_HVT U116 ( .A1(n412), .A3(n406), .A2(n382), .A4(n629), .S0(n335), 
        .S1(n288), .Y(n531) );
  NAND2X0_HVT U118 ( .A1(n304), .A2(n313), .Y(n529) );
  MUX41X1_HVT U119 ( .A1(n428), .A3(n530), .A2(n607), .A4(n529), .S0(n335), 
        .S1(n288), .Y(n528) );
  MUX41X1_HVT U120 ( .A1(n528), .A3(n532), .A2(n531), .A4(n534), .S0(n352), 
        .S1(n298), .Y(n527) );
  MUX41X1_HVT U122 ( .A1(n417), .A3(n325), .A2(n598), .A4(n420), .S0(n335), 
        .S1(n312), .Y(n526) );
  MUX41X1_HVT U124 ( .A1(n327), .A3(n525), .A2(n621), .A4(n311), .S0(n343), 
        .S1(n335), .Y(n524) );
  AOI21X1_HVT U127 ( .A1(n340), .A2(n520), .A3(n389), .Y(n521) );
  NAND2X0_HVT U129 ( .A1(n339), .A2(n365), .Y(n518) );
  MUX41X1_HVT U130 ( .A1(n518), .A3(n519), .A2(n522), .A4(n521), .S0(n343), 
        .S1(n298), .Y(n517) );
  AND2X1_HVT U131 ( .A1(n331), .A2(n287), .Y(n516) );
  MUX41X1_HVT U132 ( .A1(n386), .A3(n516), .A2(n430), .A4(n395), .S0(n343), 
        .S1(n333), .Y(n515) );
  MUX41X1_HVT U133 ( .A1(n431), .A3(n388), .A2(n590), .A4(n387), .S0(n341), 
        .S1(n334), .Y(n514) );
  MUX41X1_HVT U136 ( .A1(n595), .A3(n546), .A2(n512), .A4(n393), .S0(n339), 
        .S1(n312), .Y(n511) );
  MUX41X1_HVT U137 ( .A1(n637), .A3(n615), .A2(n619), .A4(n424), .S0(n341), 
        .S1(n338), .Y(n510) );
  MUX41X1_HVT U139 ( .A1(n509), .A3(n513), .A2(n517), .A4(n523), .S0(n352), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n409), .A3(n326), .A2(n403), .A4(n633), .S0(n343), 
        .S1(n334), .Y(n508) );
  NAND2X0_HVT U141 ( .A1(n354), .A2(n286), .Y(n507) );
  MUX41X1_HVT U142 ( .A1(n507), .A3(n605), .A2(n429), .A4(n403), .S0(n340), 
        .S1(n375), .Y(n506) );
  MUX41X1_HVT U145 ( .A1(n613), .A3(n427), .A2(n504), .A4(n564), .S0(n340), 
        .S1(n296), .Y(n503) );
  MUX41X1_HVT U146 ( .A1(n503), .A3(n505), .A2(n506), .A4(n508), .S0(n350), 
        .S1(n352), .Y(n502) );
  AO21X1_HVT U148 ( .A1(n343), .A2(n390), .A3(n432), .Y(n500) );
  MUX41X1_HVT U151 ( .A1(n314), .A3(n411), .A2(n297), .A4(n498), .S0(n343), 
        .S1(n333), .Y(n497) );
  OA21X1_HVT U153 ( .A1(n383), .A2(n283), .A3(n392), .Y(n495) );
  MUX41X1_HVT U155 ( .A1(n403), .A3(n633), .A2(n625), .A4(n404), .S0(n338), 
        .S1(n296), .Y(n493) );
  NAND2X0_HVT U159 ( .A1(n489), .A2(n488), .Y(n490) );
  MUX41X1_HVT U162 ( .A1(n332), .A3(n400), .A2(n609), .A4(n486), .S0(n338), 
        .S1(n295), .Y(n485) );
  NAND2X0_HVT U163 ( .A1(n369), .A2(n196), .Y(n484) );
  NAND2X0_HVT U166 ( .A1(n634), .A2(n480), .Y(n481) );
  MUX41X1_HVT U174 ( .A1(n423), .A3(n590), .A2(n431), .A4(n437), .S0(n338), 
        .S1(n295), .Y(n472) );
  NAND2X0_HVT U177 ( .A1(n370), .A2(n313), .Y(n470) );
  MUX41X1_HVT U178 ( .A1(n328), .A3(n470), .A2(n435), .A4(n600), .S0(n338), 
        .S1(n296), .Y(n469) );
  AND2X1_HVT U179 ( .A1(n289), .A2(n356), .Y(n468) );
  OA21X1_HVT U189 ( .A1(n406), .A2(n379), .A3(n584), .Y(n459) );
  MUX41X1_HVT U190 ( .A1(n460), .A3(n461), .A2(n459), .A4(n462), .S0(n350), 
        .S1(n333), .Y(n458) );
  NAND2X0_HVT U191 ( .A1(n379), .A2(n394), .Y(n457) );
  AND2X1_HVT U192 ( .A1(n410), .A2(n455), .Y(n456) );
  NAND2X0_HVT U194 ( .A1(n602), .A2(n455), .Y(n453) );
  NAND2X0_HVT U198 ( .A1(n367), .A2(n437), .Y(n634) );
  NAND2X0_HVT U200 ( .A1(n357), .A2(n286), .Y(n520) );
  AO21X1_HVT U204 ( .A1(n355), .A2(n642), .A3(n283), .Y(n480) );
  AO21X1_HVT U206 ( .A1(n369), .A2(n432), .A3(n378), .Y(n455) );
  NAND2X0_HVT U207 ( .A1(n286), .A2(n435), .Y(n584) );
  NBUFFX2_HVT U1 ( .A(n438), .Y(n346) );
  NBUFFX2_HVT U2 ( .A(n438), .Y(n347) );
  NBUFFX2_HVT U3 ( .A(n410), .Y(n184) );
  IBUFFX2_HVT U6 ( .A(n640), .Y(n196) );
  INVX0_HVT U14 ( .A(n356), .Y(n433) );
  NBUFFX4_HVT U16 ( .A(n628), .Y(n353) );
  INVX0_HVT U17 ( .A(n318), .Y(n321) );
  MUX21X2_HVT U18 ( .A1(n319), .A2(n363), .S0(n286), .Y(n318) );
  IBUFFX2_HVT U20 ( .A(n371), .Y(n197) );
  INVX1_HVT U21 ( .A(n367), .Y(n229) );
  INVX1_HVT U22 ( .A(n369), .Y(n224) );
  INVX2_HVT U23 ( .A(n246), .Y(n231) );
  INVX1_HVT U24 ( .A(n287), .Y(n271) );
  INVX1_HVT U26 ( .A(n371), .Y(n369) );
  INVX1_HVT U27 ( .A(in[5]), .Y(n198) );
  MUX21X1_HVT U28 ( .A1(n244), .A2(n448), .S0(n342), .Y(n243) );
  IBUFFX2_HVT U29 ( .A(n346), .Y(n228) );
  MUX21X1_HVT U30 ( .A1(n331), .A2(n436), .S0(n285), .Y(n603) );
  INVX2_HVT U31 ( .A(n371), .Y(n302) );
  INVX0_HVT U33 ( .A(n619), .Y(n403) );
  MUX21X1_HVT U34 ( .A1(n435), .A2(n433), .S0(n368), .Y(n616) );
  MUX21X1_HVT U36 ( .A1(n321), .A2(n322), .S0(n342), .Y(n320) );
  INVX1_HVT U37 ( .A(n342), .Y(n323) );
  XNOR2X2_HVT U39 ( .A1(n346), .A2(n434), .Y(n628) );
  MUX21X1_HVT U40 ( .A1(n347), .A2(n433), .S0(n302), .Y(n498) );
  MUX21X1_HVT U41 ( .A1(n347), .A2(n435), .S0(n224), .Y(n475) );
  MUX41X1_HVT U43 ( .A1(n497), .A3(n493), .A2(n499), .A4(n494), .S0(n198), 
        .S1(n199), .Y(n492) );
  IBUFFX16_HVT U44 ( .A(n299), .Y(n199) );
  INVX1_HVT U45 ( .A(n598), .Y(n416) );
  XOR2X2_HVT U46 ( .A1(n355), .A2(n197), .Y(n598) );
  MUX21X2_HVT U47 ( .A1(n524), .A2(n526), .S0(n350), .Y(n523) );
  INVX0_HVT U48 ( .A(n645), .Y(n200) );
  INVX0_HVT U49 ( .A(n200), .Y(n201) );
  NAND2X0_HVT U50 ( .A1(n478), .A2(n202), .Y(n205) );
  NAND2X0_HVT U51 ( .A1(n471), .A2(n284), .Y(n208) );
  NAND2X0_HVT U52 ( .A1(n205), .A2(n208), .Y(out[6]) );
  INVX0_HVT U54 ( .A(n284), .Y(n202) );
  MUX41X1_HVT U56 ( .A1(n602), .A3(n401), .A2(n418), .A4(n414), .S0(n281), 
        .S1(n218), .Y(n464) );
  IBUFFX16_HVT U57 ( .A(n333), .Y(n218) );
  AO21X2_HVT U58 ( .A1(n584), .A2(n341), .A3(n623), .Y(n585) );
  OA21X2_HVT U59 ( .A1(n384), .A2(n379), .A3(n623), .Y(n569) );
  MUX41X1_HVT U60 ( .A1(n456), .A3(n457), .A2(n454), .A4(n453), .S0(n336), 
        .S1(n219), .Y(n452) );
  IBUFFX16_HVT U61 ( .A(n350), .Y(n219) );
  INVX1_HVT U62 ( .A(n623), .Y(n401) );
  MUX41X1_HVT U63 ( .A1(n475), .A3(n557), .A2(n622), .A4(n324), .S0(n316), 
        .S1(n220), .Y(n474) );
  IBUFFX16_HVT U64 ( .A(n225), .Y(n220) );
  NBUFFX4_HVT U68 ( .A(n434), .Y(n345) );
  INVX2_HVT U69 ( .A(n303), .Y(n370) );
  NAND2X0_HVT U70 ( .A1(n567), .A2(n221), .Y(n222) );
  NAND2X0_HVT U71 ( .A1(n560), .A2(n264), .Y(n223) );
  NAND2X0_HVT U75 ( .A1(n222), .A2(n223), .Y(out[1]) );
  INVX0_HVT U76 ( .A(n264), .Y(n221) );
  INVX1_HVT U77 ( .A(n610), .Y(n410) );
  INVX1_HVT U79 ( .A(n269), .Y(n618) );
  MUX21X1_HVT U80 ( .A1(n490), .A2(n491), .S0(n340), .Y(n487) );
  IBUFFX16_HVT U86 ( .A(n295), .Y(n225) );
  MUX21X2_HVT U87 ( .A1(n537), .A2(n527), .S0(n226), .Y(out[3]) );
  IBUFFX16_HVT U91 ( .A(in[7]), .Y(n226) );
  MUX21X1_HVT U92 ( .A1(n353), .A2(n228), .S0(n229), .Y(n227) );
  INVX8_HVT U93 ( .A(n227), .Y(n608) );
  INVX1_HVT U94 ( .A(n353), .Y(n437) );
  MUX41X1_HVT U95 ( .A1(n608), .A3(n361), .A2(n435), .A4(n364), .S0(n268), 
        .S1(n230), .Y(n473) );
  IBUFFX16_HVT U96 ( .A(n295), .Y(n230) );
  NAND2X0_HVT U97 ( .A1(n345), .A2(n231), .Y(n232) );
  NAND2X0_HVT U98 ( .A1(n354), .A2(n246), .Y(n233) );
  NAND2X0_HVT U102 ( .A1(n232), .A2(n233), .Y(n623) );
  IBUFFX2_HVT U103 ( .A(n367), .Y(n246) );
  IBUFFX2_HVT U106 ( .A(in[7]), .Y(n264) );
  NAND2X0_HVT U111 ( .A1(n593), .A2(n234), .Y(n235) );
  NAND2X0_HVT U113 ( .A1(n592), .A2(n339), .Y(n236) );
  NAND2X0_HVT U117 ( .A1(n235), .A2(n236), .Y(n591) );
  IBUFFX2_HVT U121 ( .A(n339), .Y(n234) );
  NAND2X0_HVT U123 ( .A1(n582), .A2(n237), .Y(n238) );
  NAND2X0_HVT U125 ( .A1(n575), .A2(n310), .Y(n239) );
  NAND2X0_HVT U126 ( .A1(n238), .A2(n239), .Y(out[0]) );
  INVX0_HVT U128 ( .A(n310), .Y(n237) );
  MUX21X1_HVT U134 ( .A1(n404), .A2(n396), .S0(n342), .Y(n593) );
  INVX1_HVT U135 ( .A(in[3]), .Y(n434) );
  INVX0_HVT U138 ( .A(n434), .Y(n313) );
  MUX41X1_HVT U143 ( .A1(n641), .A3(n636), .A2(n418), .A4(n421), .S0(n245), 
        .S1(n379), .Y(n565) );
  INVX1_HVT U144 ( .A(n378), .Y(n376) );
  MUX41X1_HVT U147 ( .A1(n418), .A3(n269), .A2(n354), .A4(n590), .S0(n259), 
        .S1(n258), .Y(n589) );
  NAND2X0_HVT U149 ( .A1(n331), .A2(n240), .Y(n241) );
  NAND2X0_HVT U150 ( .A1(n433), .A2(n257), .Y(n242) );
  NAND2X0_HVT U152 ( .A1(n241), .A2(n242), .Y(n451) );
  INVX0_HVT U154 ( .A(n257), .Y(n240) );
  INVX0_HVT U156 ( .A(n316), .Y(n258) );
  IBUFFX2_HVT U157 ( .A(n283), .Y(n259) );
  IBUFFX2_HVT U158 ( .A(n303), .Y(n257) );
  INVX0_HVT U160 ( .A(n451), .Y(n418) );
  INVX1_HVT U161 ( .A(in[4]), .Y(n378) );
  INVX1_HVT U164 ( .A(n243), .Y(n462) );
  NAND2X0_HVT U165 ( .A1(n437), .A2(n304), .Y(n244) );
  IBUFFX2_HVT U167 ( .A(n448), .Y(n421) );
  IBUFFX16_HVT U168 ( .A(n336), .Y(n245) );
  MUX41X1_HVT U169 ( .A1(n401), .A3(n607), .A2(n484), .A4(n636), .S0(n247), 
        .S1(n248), .Y(n483) );
  IBUFFX16_HVT U170 ( .A(n335), .Y(n247) );
  IBUFFX16_HVT U171 ( .A(n296), .Y(n248) );
  MUX21X1_HVT U172 ( .A1(n401), .A2(n581), .S0(n330), .Y(n580) );
  MUX41X1_HVT U173 ( .A1(n545), .A3(n547), .A2(n548), .A4(n550), .S0(n349), 
        .S1(n352), .Y(n544) );
  NAND2X0_HVT U175 ( .A1(n551), .A2(n249), .Y(n250) );
  NAND2X0_HVT U176 ( .A1(n544), .A2(n290), .Y(n251) );
  NAND2X0_HVT U180 ( .A1(n250), .A2(n251), .Y(out[2]) );
  INVX0_HVT U181 ( .A(n290), .Y(n249) );
  MUX41X2_HVT U182 ( .A1(n419), .A3(n631), .A2(n404), .A4(n424), .S0(n337), 
        .S1(n375), .Y(n550) );
  NAND2X0_HVT U183 ( .A1(n641), .A2(n252), .Y(n253) );
  NAND2X0_HVT U184 ( .A1(n403), .A2(n260), .Y(n254) );
  NAND2X0_HVT U185 ( .A1(n253), .A2(n254), .Y(n588) );
  INVX1_HVT U186 ( .A(n260), .Y(n252) );
  IBUFFX2_HVT U187 ( .A(n340), .Y(n260) );
  MUX41X1_HVT U188 ( .A1(n425), .A3(n549), .A2(n616), .A4(n411), .S0(n255), 
        .S1(n375), .Y(n548) );
  IBUFFX16_HVT U193 ( .A(n337), .Y(n255) );
  MUX41X1_HVT U195 ( .A1(n587), .A3(n591), .A2(n583), .A4(n589), .S0(n352), 
        .S1(n256), .Y(n582) );
  IBUFFX16_HVT U196 ( .A(n349), .Y(n256) );
  IBUFFX2_HVT U197 ( .A(n371), .Y(n285) );
  IBUFFX2_HVT U199 ( .A(n601), .Y(n414) );
  MUX41X1_HVT U201 ( .A1(n269), .A3(n423), .A2(n329), .A4(n385), .S0(n291), 
        .S1(n283), .Y(n559) );
  MUX21X1_HVT U202 ( .A1(n315), .A2(n353), .S0(n285), .Y(n314) );
  NAND2X0_HVT U203 ( .A1(n465), .A2(n261), .Y(n262) );
  NAND2X0_HVT U205 ( .A1(n464), .A2(n282), .Y(n263) );
  NAND2X0_HVT U208 ( .A1(n263), .A2(n262), .Y(n463) );
  INVX0_HVT U209 ( .A(n282), .Y(n261) );
  IBUFFX2_HVT U210 ( .A(n350), .Y(n282) );
  INVX1_HVT U211 ( .A(in[6]), .Y(n438) );
  NAND2X0_HVT U212 ( .A1(n347), .A2(n265), .Y(n266) );
  NAND2X0_HVT U213 ( .A1(n355), .A2(n303), .Y(n267) );
  NAND2X0_HVT U214 ( .A1(n266), .A2(n267), .Y(n619) );
  INVX0_HVT U215 ( .A(n303), .Y(n265) );
  IBUFFX16_HVT U216 ( .A(n338), .Y(n268) );
  MUX21X1_HVT U217 ( .A1(n270), .A2(n361), .S0(n271), .Y(n269) );
  IBUFFX16_HVT U218 ( .A(n346), .Y(n270) );
  MUX21X1_HVT U219 ( .A1(n618), .A2(n621), .S0(n343), .Y(n482) );
  INVX1_HVT U220 ( .A(n371), .Y(n366) );
  MUX41X1_HVT U221 ( .A1(n552), .A3(n556), .A2(n558), .A4(n559), .S0(n349), 
        .S1(n352), .Y(n551) );
  NAND2X0_HVT U222 ( .A1(n553), .A2(n272), .Y(n273) );
  NAND2X0_HVT U223 ( .A1(n554), .A2(n339), .Y(n274) );
  NAND2X0_HVT U224 ( .A1(n273), .A2(n274), .Y(n552) );
  IBUFFX2_HVT U225 ( .A(n339), .Y(n272) );
  INVX2_HVT U226 ( .A(n351), .Y(n352) );
  INVX2_HVT U227 ( .A(n348), .Y(n349) );
  NAND2X1_HVT U228 ( .A1(n495), .A2(n275), .Y(n276) );
  NAND2X0_HVT U229 ( .A1(n496), .A2(n340), .Y(n277) );
  NAND2X0_HVT U230 ( .A1(n276), .A2(n277), .Y(n494) );
  IBUFFX2_HVT U231 ( .A(n340), .Y(n275) );
  NAND2X0_HVT U232 ( .A1(n502), .A2(n278), .Y(n279) );
  NAND2X0_HVT U233 ( .A1(n492), .A2(n310), .Y(n280) );
  NAND2X0_HVT U234 ( .A1(n279), .A2(n280), .Y(out[5]) );
  INVX0_HVT U235 ( .A(n310), .Y(n278) );
  MUX21X1_HVT U236 ( .A1(n619), .A2(n329), .S0(n343), .Y(n496) );
  MUX21X2_HVT U237 ( .A1(n601), .A2(n420), .S0(n342), .Y(n491) );
  IBUFFX16_HVT U238 ( .A(n341), .Y(n281) );
  NBUFFX2_HVT U239 ( .A(n379), .Y(n283) );
  IBUFFX2_HVT U240 ( .A(in[7]), .Y(n284) );
  AO21X1_HVT U241 ( .A1(n287), .A2(n365), .A3(n378), .Y(n488) );
  INVX1_HVT U242 ( .A(n366), .Y(n286) );
  INVX1_HVT U243 ( .A(n366), .Y(n287) );
  INVX0_HVT U244 ( .A(n366), .Y(n303) );
  OR2X1_HVT U245 ( .A1(n434), .A2(n438), .Y(n643) );
  INVX1_HVT U246 ( .A(n371), .Y(n368) );
  INVX1_HVT U247 ( .A(n371), .Y(n367) );
  NBUFFX2_HVT U248 ( .A(n375), .Y(n288) );
  INVX1_HVT U249 ( .A(n378), .Y(n375) );
  IBUFFX2_HVT U250 ( .A(in[7]), .Y(n290) );
  INVX1_HVT U251 ( .A(n387), .Y(n289) );
  INVX0_HVT U252 ( .A(n639), .Y(n387) );
  IBUFFX16_HVT U253 ( .A(n335), .Y(n291) );
  NAND2X0_HVT U254 ( .A1(n327), .A2(n292), .Y(n293) );
  NAND2X0_HVT U255 ( .A1(n415), .A2(n305), .Y(n294) );
  NAND2X0_HVT U256 ( .A1(n293), .A2(n294), .Y(n454) );
  INVX0_HVT U257 ( .A(n305), .Y(n292) );
  INVX0_HVT U258 ( .A(n341), .Y(n305) );
  INVX2_HVT U259 ( .A(n323), .Y(n312) );
  NBUFFX4_HVT U260 ( .A(n374), .Y(n295) );
  NBUFFX2_HVT U261 ( .A(n374), .Y(n296) );
  IBUFFX2_HVT U262 ( .A(n378), .Y(n374) );
  NAND2X0_HVT U263 ( .A1(n197), .A2(n365), .Y(n639) );
  INVX1_HVT U264 ( .A(n438), .Y(n331) );
  INVX0_HVT U265 ( .A(n297), .Y(n622) );
  MUX21X1_HVT U266 ( .A1(n590), .A2(n311), .S0(n323), .Y(n586) );
  INVX0_HVT U267 ( .A(in[7]), .Y(n310) );
  INVX0_HVT U268 ( .A(n298), .Y(n299) );
  INVX1_HVT U269 ( .A(n366), .Y(n304) );
  MUX21X1_HVT U270 ( .A1(n363), .A2(n353), .S0(n286), .Y(n297) );
  MUX21X2_HVT U271 ( .A1(n535), .A2(n536), .S0(n340), .Y(n534) );
  MUX21X1_HVT U272 ( .A1(n347), .A2(n345), .S0(n286), .Y(n599) );
  MUX41X1_HVT U273 ( .A1(n385), .A3(n314), .A2(n388), .A4(n642), .S0(n337), 
        .S1(n323), .Y(n465) );
  INVX0_HVT U274 ( .A(n378), .Y(n377) );
  INVX0_HVT U275 ( .A(n602), .Y(n388) );
  INVX0_HVT U276 ( .A(n599), .Y(n415) );
  MUX21X2_HVT U277 ( .A1(n402), .A2(n588), .S0(n330), .Y(n587) );
  MUX41X1_HVT U278 ( .A1(n472), .A3(n474), .A2(n473), .A4(n476), .S0(n352), 
        .S1(n298), .Y(n471) );
  IBUFFX2_HVT U279 ( .A(n348), .Y(n298) );
  MUX41X1_HVT U280 ( .A1(n391), .A3(n633), .A2(n435), .A4(n289), .S0(n316), 
        .S1(n379), .Y(n574) );
  MUX41X1_HVT U281 ( .A1(n328), .A3(n327), .A2(n324), .A4(n477), .S0(n377), 
        .S1(n338), .Y(n476) );
  IBUFFX2_HVT U282 ( .A(in[4]), .Y(n379) );
  NAND2X0_HVT U283 ( .A1(n467), .A2(n299), .Y(n300) );
  NAND2X0_HVT U284 ( .A1(n469), .A2(n349), .Y(n301) );
  NAND2X0_HVT U285 ( .A1(n300), .A2(n301), .Y(n466) );
  MUX41X1_HVT U286 ( .A1(n466), .A3(n458), .A2(n463), .A4(n452), .S0(n310), 
        .S1(n351), .Y(out[7]) );
  INVX1_HVT U287 ( .A(in[5]), .Y(n351) );
  INVX1_HVT U288 ( .A(in[0]), .Y(n371) );
  INVX0_HVT U289 ( .A(n320), .Y(n460) );
  MUX41X1_HVT U290 ( .A1(n599), .A3(n468), .A2(n380), .A4(n612), .S0(n316), 
        .S1(n283), .Y(n467) );
  NAND2X0_HVT U291 ( .A1(n329), .A2(n305), .Y(n306) );
  NAND2X0_HVT U292 ( .A1(n596), .A2(n343), .Y(n307) );
  NAND2X0_HVT U293 ( .A1(n306), .A2(n307), .Y(n461) );
  XOR2X1_HVT U294 ( .A1(n356), .A2(n368), .Y(n596) );
  MUX41X1_HVT U295 ( .A1(n487), .A3(n485), .A2(n483), .A4(n479), .S0(n299), 
        .S1(n351), .Y(n478) );
  NAND2X0_HVT U296 ( .A1(n481), .A2(n316), .Y(n308) );
  NAND2X0_HVT U297 ( .A1(n482), .A2(n339), .Y(n309) );
  NAND2X0_HVT U298 ( .A1(n308), .A2(n309), .Y(n479) );
  MUX41X1_HVT U299 ( .A1(n627), .A3(n408), .A2(n626), .A4(n406), .S0(n316), 
        .S1(n379), .Y(n566) );
  INVX1_HVT U300 ( .A(n317), .Y(n477) );
  INVX1_HVT U301 ( .A(n603), .Y(n322) );
  INVX1_HVT U302 ( .A(n311), .Y(n621) );
  INVX0_HVT U303 ( .A(n344), .Y(n315) );
  INVX0_HVT U304 ( .A(n346), .Y(n319) );
  INVX0_HVT U305 ( .A(n335), .Y(n316) );
  MUX21X1_HVT U306 ( .A1(n345), .A2(n361), .S0(n304), .Y(n311) );
  MUX41X1_HVT U307 ( .A1(n364), .A3(n396), .A2(n313), .A4(n395), .S0(n316), 
        .S1(n283), .Y(n576) );
  NBUFFX2_HVT U308 ( .A(n434), .Y(n344) );
  MUX21X2_HVT U309 ( .A1(n586), .A2(n585), .S0(n339), .Y(n583) );
  MUX41X1_HVT U310 ( .A1(n580), .A3(n577), .A2(n579), .A4(n576), .S0(n351), 
        .S1(n299), .Y(n575) );
  MUX21X1_HVT U311 ( .A1(n358), .A2(n365), .S0(n304), .Y(n317) );
  INVX1_HVT U312 ( .A(n358), .Y(n436) );
  INVX1_HVT U313 ( .A(n361), .Y(n432) );
  MUX41X1_HVT U314 ( .A1(n621), .A3(n624), .A2(n414), .A4(n196), .S0(n316), 
        .S1(n323), .Y(n505) );
  MUX21X2_HVT U315 ( .A1(n297), .A2(n642), .S0(n339), .Y(n581) );
  INVX0_HVT U316 ( .A(in[1]), .Y(n348) );
  NBUFFX2_HVT U317 ( .A(n644), .Y(n361) );
  NBUFFX2_HVT U318 ( .A(n644), .Y(n362) );
  NBUFFX2_HVT U319 ( .A(n644), .Y(n363) );
  AND2X1_HVT U320 ( .A1(n639), .A2(n362), .Y(n324) );
  AND2X1_HVT U321 ( .A1(n362), .A2(n629), .Y(n325) );
  NAND2X0_HVT U322 ( .A1(n344), .A2(n346), .Y(n644) );
  MUX21X1_HVT U323 ( .A1(n432), .A2(n437), .S0(n369), .Y(n611) );
  MUX21X1_HVT U324 ( .A1(n437), .A2(n345), .S0(n368), .Y(n605) );
  MUX21X1_HVT U325 ( .A1(n432), .A2(n436), .S0(n367), .Y(n594) );
  MUX21X1_HVT U326 ( .A1(n501), .A2(n500), .S0(n339), .Y(n499) );
  MUX21X1_HVT U327 ( .A1(n430), .A2(n386), .S0(n341), .Y(n501) );
  MUX21X1_HVT U328 ( .A1(n354), .A2(n433), .S0(n367), .Y(n610) );
  MUX21X1_HVT U329 ( .A1(n437), .A2(n347), .S0(n368), .Y(n441) );
  MUX21X1_HVT U330 ( .A1(n356), .A2(n363), .S0(n368), .Y(n440) );
  MUX21X1_HVT U331 ( .A1(n355), .A2(n435), .S0(n367), .Y(n613) );
  MUX21X1_HVT U332 ( .A1(n345), .A2(n432), .S0(n370), .Y(n614) );
  MUX21X1_HVT U333 ( .A1(n611), .A2(n325), .S0(n340), .Y(n519) );
  MUX21X1_HVT U334 ( .A1(n356), .A2(n359), .S0(n285), .Y(n486) );
  MUX21X1_HVT U335 ( .A1(n361), .A2(n357), .S0(n302), .Y(n504) );
  MUX21X1_HVT U336 ( .A1(n429), .A2(n326), .S0(n339), .Y(n522) );
  XOR2X1_HVT U337 ( .A1(n358), .A2(n285), .Y(n597) );
  XNOR2X1_HVT U338 ( .A1(n361), .A2(n302), .Y(n326) );
  MUX21X1_HVT U339 ( .A1(n331), .A2(n435), .S0(n197), .Y(n620) );
  MUX21X1_HVT U340 ( .A1(n357), .A2(n331), .S0(n369), .Y(n615) );
  MUX21X1_HVT U341 ( .A1(n345), .A2(n436), .S0(n302), .Y(n601) );
  XOR2X1_HVT U342 ( .A1(n370), .A2(n331), .Y(n595) );
  MUX21X1_HVT U343 ( .A1(n432), .A2(n331), .S0(n285), .Y(n512) );
  MUX21X1_HVT U344 ( .A1(n436), .A2(n345), .S0(n370), .Y(n449) );
  MUX21X1_HVT U345 ( .A1(n435), .A2(n355), .S0(n367), .Y(n446) );
  MUX21X1_HVT U346 ( .A1(n345), .A2(n362), .S0(n197), .Y(n448) );
  MUX21X1_HVT U347 ( .A1(n360), .A2(n362), .S0(n197), .Y(n626) );
  MUX21X1_HVT U348 ( .A1(n364), .A2(n363), .S0(n197), .Y(n630) );
  MUX21X1_HVT U349 ( .A1(n359), .A2(n345), .S0(n370), .Y(n625) );
  MUX21X1_HVT U350 ( .A1(n389), .A2(n603), .S0(n342), .Y(n536) );
  MUX21X1_HVT U351 ( .A1(n555), .A2(n359), .S0(n302), .Y(n554) );
  MUX21X1_HVT U352 ( .A1(n391), .A2(n354), .S0(n342), .Y(n553) );
  MUX21X1_HVT U353 ( .A1(n354), .A2(n347), .S0(n342), .Y(n555) );
  XOR2X1_HVT U354 ( .A1(n364), .A2(n370), .Y(n607) );
  MUX21X1_HVT U355 ( .A1(n347), .A2(n363), .S0(n285), .Y(n541) );
  MUX21X1_HVT U356 ( .A1(n331), .A2(n364), .S0(n369), .Y(n627) );
  MUX21X1_HVT U357 ( .A1(n360), .A2(n347), .S0(n368), .Y(n525) );
  MUX21X1_HVT U358 ( .A1(n344), .A2(n331), .S0(n197), .Y(n442) );
  MUX21X1_HVT U359 ( .A1(n331), .A2(n360), .S0(n285), .Y(n450) );
  MUX21X1_HVT U360 ( .A1(n347), .A2(n355), .S0(n370), .Y(n604) );
  MUX21X1_HVT U361 ( .A1(n344), .A2(n359), .S0(n369), .Y(n443) );
  MUX21X1_HVT U362 ( .A1(n359), .A2(n331), .S0(n302), .Y(n447) );
  AND2X1_HVT U363 ( .A1(n368), .A2(n347), .Y(n327) );
  NBUFFX2_HVT U364 ( .A(n377), .Y(n341) );
  NBUFFX2_HVT U365 ( .A(n377), .Y(n343) );
  NBUFFX2_HVT U366 ( .A(n377), .Y(n342) );
  NBUFFX2_HVT U367 ( .A(n640), .Y(n356) );
  NBUFFX2_HVT U368 ( .A(n201), .Y(n364) );
  NBUFFX2_HVT U369 ( .A(n628), .Y(n354) );
  AND2X1_HVT U370 ( .A1(n436), .A2(n287), .Y(n328) );
  NBUFFX2_HVT U371 ( .A(n640), .Y(n357) );
  NBUFFX2_HVT U372 ( .A(n643), .Y(n358) );
  NBUFFX2_HVT U373 ( .A(n628), .Y(n355) );
  AND2X1_HVT U374 ( .A1(n360), .A2(n304), .Y(n329) );
  NBUFFX2_HVT U375 ( .A(n643), .Y(n360) );
  MUX21X1_HVT U376 ( .A1(n570), .A2(n569), .S0(n340), .Y(n568) );
  MUX21X1_HVT U377 ( .A1(n420), .A2(n381), .S0(n341), .Y(n570) );
  NBUFFX2_HVT U378 ( .A(n201), .Y(n365) );
  NBUFFX2_HVT U379 ( .A(n643), .Y(n359) );
  NBUFFX2_HVT U380 ( .A(n373), .Y(n338) );
  NBUFFX2_HVT U381 ( .A(n372), .Y(n340) );
  NBUFFX2_HVT U382 ( .A(n372), .Y(n339) );
  XNOR2X1_HVT U383 ( .A1(n378), .A2(n335), .Y(n330) );
  NBUFFX2_HVT U384 ( .A(n373), .Y(n335) );
  NBUFFX2_HVT U385 ( .A(n372), .Y(n333) );
  NBUFFX2_HVT U386 ( .A(n372), .Y(n334) );
  NBUFFX2_HVT U387 ( .A(n373), .Y(n337) );
  NBUFFX2_HVT U388 ( .A(n373), .Y(n336) );
  INVX1_HVT U389 ( .A(n348), .Y(n350) );
  NAND2X0_HVT U390 ( .A1(n315), .A2(n346), .Y(n645) );
  MUX21X1_HVT U391 ( .A1(n514), .A2(n515), .S0(n298), .Y(n513) );
  MUX21X1_HVT U392 ( .A1(n510), .A2(n511), .S0(n350), .Y(n509) );
  INVX0_HVT U393 ( .A(n332), .Y(n600) );
  MUX21X1_HVT U394 ( .A1(n435), .A2(n313), .S0(n369), .Y(n439) );
  MUX21X1_HVT U395 ( .A1(n357), .A2(n313), .S0(n370), .Y(n549) );
  MUX21X1_HVT U396 ( .A1(n436), .A2(n433), .S0(n197), .Y(n530) );
  MUX21X1_HVT U397 ( .A1(n313), .A2(n357), .S0(n302), .Y(n444) );
  MUX21X1_HVT U398 ( .A1(n364), .A2(n313), .S0(n368), .Y(n489) );
  MUX21X1_HVT U399 ( .A1(n347), .A2(n313), .S0(n302), .Y(n617) );
  MUX21X1_HVT U400 ( .A1(n313), .A2(n365), .S0(n285), .Y(n445) );
  NBUFFX2_HVT U401 ( .A(in[2]), .Y(n373) );
  NBUFFX2_HVT U402 ( .A(in[2]), .Y(n372) );
  MUX21X1_HVT U403 ( .A1(n365), .A2(n356), .S0(n287), .Y(n332) );
  INVX1_HVT U404 ( .A(n645), .Y(n435) );
  INVX0_HVT U405 ( .A(n633), .Y(n380) );
  INVX0_HVT U406 ( .A(n612), .Y(n381) );
  INVX0_HVT U407 ( .A(n606), .Y(n382) );
  INVX0_HVT U408 ( .A(n546), .Y(n383) );
  INVX0_HVT U409 ( .A(n507), .Y(n384) );
  INVX0_HVT U410 ( .A(n642), .Y(n385) );
  INVX0_HVT U411 ( .A(n641), .Y(n386) );
  INVX0_HVT U412 ( .A(n638), .Y(n389) );
  INVX0_HVT U413 ( .A(n637), .Y(n390) );
  INVX0_HVT U414 ( .A(n609), .Y(n391) );
  INVX0_HVT U415 ( .A(n631), .Y(n392) );
  INVX0_HVT U416 ( .A(n636), .Y(n393) );
  INVX0_HVT U417 ( .A(n632), .Y(n394) );
  INVX0_HVT U418 ( .A(n630), .Y(n395) );
  INVX0_HVT U419 ( .A(n629), .Y(n396) );
  INVX0_HVT U420 ( .A(n627), .Y(n397) );
  INVX0_HVT U421 ( .A(n626), .Y(n398) );
  INVX0_HVT U422 ( .A(n625), .Y(n399) );
  INVX0_HVT U423 ( .A(n624), .Y(n400) );
  INVX0_HVT U424 ( .A(n620), .Y(n402) );
  INVX0_HVT U425 ( .A(n617), .Y(n404) );
  INVX0_HVT U426 ( .A(n616), .Y(n405) );
  INVX0_HVT U427 ( .A(n615), .Y(n406) );
  INVX0_HVT U428 ( .A(n614), .Y(n407) );
  INVX0_HVT U429 ( .A(n613), .Y(n408) );
  INVX0_HVT U430 ( .A(n611), .Y(n409) );
  INVX0_HVT U431 ( .A(n607), .Y(n411) );
  INVX0_HVT U432 ( .A(n605), .Y(n412) );
  INVX0_HVT U433 ( .A(n604), .Y(n413) );
  INVX0_HVT U434 ( .A(n635), .Y(n417) );
  INVX0_HVT U435 ( .A(n450), .Y(n419) );
  INVX0_HVT U436 ( .A(n449), .Y(n420) );
  INVX0_HVT U437 ( .A(n447), .Y(n422) );
  INVX0_HVT U438 ( .A(n446), .Y(n423) );
  INVX0_HVT U439 ( .A(n445), .Y(n424) );
  INVX0_HVT U440 ( .A(n444), .Y(n425) );
  INVX0_HVT U441 ( .A(n443), .Y(n426) );
  INVX0_HVT U442 ( .A(n442), .Y(n427) );
  INVX0_HVT U443 ( .A(n489), .Y(n428) );
  INVX0_HVT U444 ( .A(n441), .Y(n429) );
  INVX0_HVT U445 ( .A(n440), .Y(n430) );
  INVX0_HVT U446 ( .A(n439), .Y(n431) );
endmodule

