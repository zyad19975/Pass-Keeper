
module ram_dp_DATA_WIDTH4_ADDR_WIDTH4_6 ( clk, rst, write, a_addr, a_din, 
        b_din, b_dout );
  input [3:0] a_addr;
  input [3:0] a_din;
  input [3:0] b_din;
  output [15:0] b_dout;
  input clk, rst, write;
  wire   N17, N18, N19, N20, \mem[15][15] , \mem[15][14] , \mem[15][13] ,
         \mem[15][12] , \mem[15][11] , \mem[15][10] , \mem[15][9] ,
         \mem[15][8] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][15] ,
         \mem[14][14] , \mem[14][13] , \mem[14][12] , \mem[14][11] ,
         \mem[14][10] , \mem[14][9] , \mem[14][8] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][15] , \mem[13][14] , \mem[13][13] ,
         \mem[13][12] , \mem[13][11] , \mem[13][10] , \mem[13][9] ,
         \mem[13][8] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][15] ,
         \mem[12][14] , \mem[12][13] , \mem[12][12] , \mem[12][11] ,
         \mem[12][10] , \mem[12][9] , \mem[12][8] , \mem[12][7] , \mem[12][6] ,
         \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] , \mem[12][1] ,
         \mem[12][0] , \mem[11][15] , \mem[11][14] , \mem[11][13] ,
         \mem[11][12] , \mem[11][11] , \mem[11][10] , \mem[11][9] ,
         \mem[11][8] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][15] , \mem[9][14] , \mem[9][13] , \mem[9][12] ,
         \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] , \mem[9][7] ,
         \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] ,
         \mem[9][1] , \mem[9][0] , \mem[8][15] , \mem[8][14] , \mem[8][13] ,
         \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] , \mem[8][8] ,
         \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] , \mem[8][3] ,
         \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][15] , \mem[7][14] ,
         \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] ,
         \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][15] ,
         \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] ,
         \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][15] , \mem[3][14] , \mem[3][13] ,
         \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] ,
         \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] ,
         \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][15] ,
         \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310,
         N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453,
         N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464,
         N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519,
         N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530,
         N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177;
  assign N17 = b_din[0];
  assign N18 = b_din[1];
  assign N19 = b_din[2];
  assign N20 = b_din[3];

  DFFNX1_HVT \b_dout_reg[15]  ( .D(n162), .CLK(clk), .Q(b_dout[15]) );
  DFFNX1_HVT \b_dout_reg[14]  ( .D(n163), .CLK(clk), .Q(b_dout[14]) );
  DFFNX1_HVT \b_dout_reg[13]  ( .D(n164), .CLK(clk), .Q(b_dout[13]) );
  DFFNX1_HVT \b_dout_reg[12]  ( .D(n165), .CLK(clk), .Q(b_dout[12]) );
  DFFNX1_HVT \b_dout_reg[11]  ( .D(n166), .CLK(clk), .Q(b_dout[11]) );
  DFFNX1_HVT \b_dout_reg[10]  ( .D(n167), .CLK(clk), .Q(b_dout[10]) );
  DFFNX1_HVT \b_dout_reg[9]  ( .D(n168), .CLK(clk), .Q(b_dout[9]) );
  DFFNX1_HVT \b_dout_reg[8]  ( .D(n169), .CLK(clk), .Q(b_dout[8]) );
  DFFNX1_HVT \b_dout_reg[7]  ( .D(n170), .CLK(clk), .Q(b_dout[7]) );
  DFFNX1_HVT \b_dout_reg[6]  ( .D(n171), .CLK(clk), .Q(b_dout[6]) );
  DFFNX1_HVT \b_dout_reg[5]  ( .D(n172), .CLK(clk), .Q(b_dout[5]) );
  DFFNX1_HVT \b_dout_reg[4]  ( .D(n173), .CLK(clk), .Q(b_dout[4]) );
  DFFNX1_HVT \b_dout_reg[3]  ( .D(n174), .CLK(clk), .Q(b_dout[3]) );
  DFFNX1_HVT \b_dout_reg[2]  ( .D(n175), .CLK(clk), .Q(b_dout[2]) );
  DFFNX1_HVT \b_dout_reg[1]  ( .D(n176), .CLK(clk), .Q(b_dout[1]) );
  DFFNX1_HVT \b_dout_reg[0]  ( .D(n177), .CLK(clk), .Q(b_dout[0]) );
  LATCHX1_HVT \mem_reg[15][15]  ( .CLK(N552), .D(n6), .Q(\mem[15][15] ) );
  LATCHX1_HVT \mem_reg[15][14]  ( .CLK(N551), .D(n6), .Q(\mem[15][14] ) );
  LATCHX1_HVT \mem_reg[15][13]  ( .CLK(N550), .D(n6), .Q(\mem[15][13] ) );
  LATCHX1_HVT \mem_reg[15][12]  ( .CLK(N549), .D(n11), .Q(\mem[15][12] ) );
  LATCHX1_HVT \mem_reg[15][11]  ( .CLK(N548), .D(n6), .Q(\mem[15][11] ) );
  LATCHX1_HVT \mem_reg[15][10]  ( .CLK(N547), .D(n6), .Q(\mem[15][10] ) );
  LATCHX1_HVT \mem_reg[15][9]  ( .CLK(N546), .D(n6), .Q(\mem[15][9] ) );
  LATCHX1_HVT \mem_reg[15][8]  ( .CLK(N545), .D(n6), .Q(\mem[15][8] ) );
  LATCHX1_HVT \mem_reg[15][7]  ( .CLK(N544), .D(n7), .Q(\mem[15][7] ) );
  LATCHX1_HVT \mem_reg[15][6]  ( .CLK(N543), .D(n7), .Q(\mem[15][6] ) );
  LATCHX1_HVT \mem_reg[15][5]  ( .CLK(N542), .D(n7), .Q(\mem[15][5] ) );
  LATCHX1_HVT \mem_reg[15][4]  ( .CLK(N541), .D(n7), .Q(\mem[15][4] ) );
  LATCHX1_HVT \mem_reg[15][3]  ( .CLK(N540), .D(n7), .Q(\mem[15][3] ) );
  LATCHX1_HVT \mem_reg[15][2]  ( .CLK(N539), .D(n7), .Q(\mem[15][2] ) );
  LATCHX1_HVT \mem_reg[15][1]  ( .CLK(N538), .D(n7), .Q(\mem[15][1] ) );
  LATCHX1_HVT \mem_reg[15][0]  ( .CLK(N537), .D(n7), .Q(\mem[15][0] ) );
  LATCHX1_HVT \mem_reg[14][15]  ( .CLK(N536), .D(n1), .Q(\mem[14][15] ) );
  LATCHX1_HVT \mem_reg[14][14]  ( .CLK(N535), .D(n17), .Q(\mem[14][14] ) );
  LATCHX1_HVT \mem_reg[14][13]  ( .CLK(N534), .D(n11), .Q(\mem[14][13] ) );
  LATCHX1_HVT \mem_reg[14][12]  ( .CLK(N533), .D(n11), .Q(\mem[14][12] ) );
  LATCHX1_HVT \mem_reg[14][11]  ( .CLK(N532), .D(n11), .Q(\mem[14][11] ) );
  LATCHX1_HVT \mem_reg[14][10]  ( .CLK(N531), .D(n12), .Q(\mem[14][10] ) );
  LATCHX1_HVT \mem_reg[14][9]  ( .CLK(N530), .D(n12), .Q(\mem[14][9] ) );
  LATCHX1_HVT \mem_reg[14][8]  ( .CLK(N529), .D(n12), .Q(\mem[14][8] ) );
  LATCHX1_HVT \mem_reg[14][7]  ( .CLK(N528), .D(n12), .Q(\mem[14][7] ) );
  LATCHX1_HVT \mem_reg[14][6]  ( .CLK(N527), .D(n12), .Q(\mem[14][6] ) );
  LATCHX1_HVT \mem_reg[14][5]  ( .CLK(N526), .D(n12), .Q(\mem[14][5] ) );
  LATCHX1_HVT \mem_reg[14][4]  ( .CLK(N525), .D(n12), .Q(\mem[14][4] ) );
  LATCHX1_HVT \mem_reg[14][3]  ( .CLK(N524), .D(n12), .Q(\mem[14][3] ) );
  LATCHX1_HVT \mem_reg[14][2]  ( .CLK(N523), .D(n12), .Q(\mem[14][2] ) );
  LATCHX1_HVT \mem_reg[14][1]  ( .CLK(N522), .D(n12), .Q(\mem[14][1] ) );
  LATCHX1_HVT \mem_reg[14][0]  ( .CLK(N521), .D(n12), .Q(\mem[14][0] ) );
  LATCHX1_HVT \mem_reg[13][15]  ( .CLK(N520), .D(n7), .Q(\mem[13][15] ) );
  LATCHX1_HVT \mem_reg[13][14]  ( .CLK(N519), .D(n7), .Q(\mem[13][14] ) );
  LATCHX1_HVT \mem_reg[13][13]  ( .CLK(N518), .D(n7), .Q(\mem[13][13] ) );
  LATCHX1_HVT \mem_reg[13][12]  ( .CLK(N517), .D(n7), .Q(\mem[13][12] ) );
  LATCHX1_HVT \mem_reg[13][11]  ( .CLK(N516), .D(n8), .Q(\mem[13][11] ) );
  LATCHX1_HVT \mem_reg[13][10]  ( .CLK(N515), .D(n8), .Q(\mem[13][10] ) );
  LATCHX1_HVT \mem_reg[13][9]  ( .CLK(N514), .D(n8), .Q(\mem[13][9] ) );
  LATCHX1_HVT \mem_reg[13][8]  ( .CLK(N513), .D(n8), .Q(\mem[13][8] ) );
  LATCHX1_HVT \mem_reg[13][7]  ( .CLK(N512), .D(n8), .Q(\mem[13][7] ) );
  LATCHX1_HVT \mem_reg[13][6]  ( .CLK(N511), .D(n8), .Q(\mem[13][6] ) );
  LATCHX1_HVT \mem_reg[13][5]  ( .CLK(N510), .D(n8), .Q(\mem[13][5] ) );
  LATCHX1_HVT \mem_reg[13][4]  ( .CLK(N509), .D(n8), .Q(\mem[13][4] ) );
  LATCHX1_HVT \mem_reg[13][3]  ( .CLK(N508), .D(n8), .Q(\mem[13][3] ) );
  LATCHX1_HVT \mem_reg[13][2]  ( .CLK(N507), .D(n8), .Q(\mem[13][2] ) );
  LATCHX1_HVT \mem_reg[13][1]  ( .CLK(N506), .D(n8), .Q(\mem[13][1] ) );
  LATCHX1_HVT \mem_reg[13][0]  ( .CLK(N505), .D(n8), .Q(\mem[13][0] ) );
  LATCHX1_HVT \mem_reg[12][15]  ( .CLK(N504), .D(n12), .Q(\mem[12][15] ) );
  LATCHX1_HVT \mem_reg[12][14]  ( .CLK(N503), .D(n13), .Q(\mem[12][14] ) );
  LATCHX1_HVT \mem_reg[12][13]  ( .CLK(N502), .D(n13), .Q(\mem[12][13] ) );
  LATCHX1_HVT \mem_reg[12][12]  ( .CLK(N501), .D(n13), .Q(\mem[12][12] ) );
  LATCHX1_HVT \mem_reg[12][11]  ( .CLK(N500), .D(n13), .Q(\mem[12][11] ) );
  LATCHX1_HVT \mem_reg[12][10]  ( .CLK(N499), .D(n13), .Q(\mem[12][10] ) );
  LATCHX1_HVT \mem_reg[12][9]  ( .CLK(N498), .D(n13), .Q(\mem[12][9] ) );
  LATCHX1_HVT \mem_reg[12][8]  ( .CLK(N497), .D(n13), .Q(\mem[12][8] ) );
  LATCHX1_HVT \mem_reg[12][7]  ( .CLK(N496), .D(n13), .Q(\mem[12][7] ) );
  LATCHX1_HVT \mem_reg[12][6]  ( .CLK(N494), .D(n13), .Q(\mem[12][6] ) );
  LATCHX1_HVT \mem_reg[12][5]  ( .CLK(N493), .D(n13), .Q(\mem[12][5] ) );
  LATCHX1_HVT \mem_reg[12][4]  ( .CLK(N492), .D(n13), .Q(\mem[12][4] ) );
  LATCHX1_HVT \mem_reg[12][3]  ( .CLK(N491), .D(n13), .Q(\mem[12][3] ) );
  LATCHX1_HVT \mem_reg[12][2]  ( .CLK(N490), .D(n14), .Q(\mem[12][2] ) );
  LATCHX1_HVT \mem_reg[12][1]  ( .CLK(N489), .D(n14), .Q(\mem[12][1] ) );
  LATCHX1_HVT \mem_reg[12][0]  ( .CLK(N488), .D(n14), .Q(\mem[12][0] ) );
  LATCHX1_HVT \mem_reg[11][15]  ( .CLK(N487), .D(n9), .Q(\mem[11][15] ) );
  LATCHX1_HVT \mem_reg[11][14]  ( .CLK(N486), .D(n9), .Q(\mem[11][14] ) );
  LATCHX1_HVT \mem_reg[11][13]  ( .CLK(N485), .D(n9), .Q(\mem[11][13] ) );
  LATCHX1_HVT \mem_reg[11][12]  ( .CLK(N484), .D(n9), .Q(\mem[11][12] ) );
  LATCHX1_HVT \mem_reg[11][11]  ( .CLK(N483), .D(n9), .Q(\mem[11][11] ) );
  LATCHX1_HVT \mem_reg[11][10]  ( .CLK(N482), .D(n9), .Q(\mem[11][10] ) );
  LATCHX1_HVT \mem_reg[11][9]  ( .CLK(N481), .D(n9), .Q(\mem[11][9] ) );
  LATCHX1_HVT \mem_reg[11][8]  ( .CLK(N480), .D(n9), .Q(\mem[11][8] ) );
  LATCHX1_HVT \mem_reg[11][7]  ( .CLK(N479), .D(n9), .Q(\mem[11][7] ) );
  LATCHX1_HVT \mem_reg[11][6]  ( .CLK(N478), .D(n9), .Q(\mem[11][6] ) );
  LATCHX1_HVT \mem_reg[11][5]  ( .CLK(N477), .D(n9), .Q(\mem[11][5] ) );
  LATCHX1_HVT \mem_reg[11][4]  ( .CLK(N476), .D(n9), .Q(\mem[11][4] ) );
  LATCHX1_HVT \mem_reg[11][3]  ( .CLK(N475), .D(n10), .Q(\mem[11][3] ) );
  LATCHX1_HVT \mem_reg[11][2]  ( .CLK(N474), .D(n10), .Q(\mem[11][2] ) );
  LATCHX1_HVT \mem_reg[11][1]  ( .CLK(N473), .D(n10), .Q(\mem[11][1] ) );
  LATCHX1_HVT \mem_reg[11][0]  ( .CLK(N472), .D(n10), .Q(\mem[11][0] ) );
  LATCHX1_HVT \mem_reg[10][15]  ( .CLK(N471), .D(n14), .Q(\mem[10][15] ) );
  LATCHX1_HVT \mem_reg[10][14]  ( .CLK(N470), .D(n14), .Q(\mem[10][14] ) );
  LATCHX1_HVT \mem_reg[10][13]  ( .CLK(N469), .D(n14), .Q(\mem[10][13] ) );
  LATCHX1_HVT \mem_reg[10][12]  ( .CLK(N468), .D(n14), .Q(\mem[10][12] ) );
  LATCHX1_HVT \mem_reg[10][11]  ( .CLK(N467), .D(n14), .Q(\mem[10][11] ) );
  LATCHX1_HVT \mem_reg[10][10]  ( .CLK(N466), .D(n14), .Q(\mem[10][10] ) );
  LATCHX1_HVT \mem_reg[10][9]  ( .CLK(N465), .D(n14), .Q(\mem[10][9] ) );
  LATCHX1_HVT \mem_reg[10][8]  ( .CLK(N464), .D(n14), .Q(\mem[10][8] ) );
  LATCHX1_HVT \mem_reg[10][7]  ( .CLK(N463), .D(n14), .Q(\mem[10][7] ) );
  LATCHX1_HVT \mem_reg[10][6]  ( .CLK(N462), .D(n15), .Q(\mem[10][6] ) );
  LATCHX1_HVT \mem_reg[10][5]  ( .CLK(N461), .D(n15), .Q(\mem[10][5] ) );
  LATCHX1_HVT \mem_reg[10][4]  ( .CLK(N460), .D(n15), .Q(\mem[10][4] ) );
  LATCHX1_HVT \mem_reg[10][3]  ( .CLK(N459), .D(n15), .Q(\mem[10][3] ) );
  LATCHX1_HVT \mem_reg[10][2]  ( .CLK(N458), .D(n15), .Q(\mem[10][2] ) );
  LATCHX1_HVT \mem_reg[10][1]  ( .CLK(N457), .D(n15), .Q(\mem[10][1] ) );
  LATCHX1_HVT \mem_reg[10][0]  ( .CLK(N456), .D(n15), .Q(\mem[10][0] ) );
  LATCHX1_HVT \mem_reg[9][15]  ( .CLK(N455), .D(n10), .Q(\mem[9][15] ) );
  LATCHX1_HVT \mem_reg[9][14]  ( .CLK(N454), .D(n10), .Q(\mem[9][14] ) );
  LATCHX1_HVT \mem_reg[9][13]  ( .CLK(N453), .D(n10), .Q(\mem[9][13] ) );
  LATCHX1_HVT \mem_reg[9][12]  ( .CLK(N452), .D(n10), .Q(\mem[9][12] ) );
  LATCHX1_HVT \mem_reg[9][11]  ( .CLK(N451), .D(n10), .Q(\mem[9][11] ) );
  LATCHX1_HVT \mem_reg[9][10]  ( .CLK(N450), .D(n10), .Q(\mem[9][10] ) );
  LATCHX1_HVT \mem_reg[9][9]  ( .CLK(N449), .D(n10), .Q(\mem[9][9] ) );
  LATCHX1_HVT \mem_reg[9][8]  ( .CLK(N448), .D(n10), .Q(\mem[9][8] ) );
  LATCHX1_HVT \mem_reg[9][7]  ( .CLK(N447), .D(n11), .Q(\mem[9][7] ) );
  LATCHX1_HVT \mem_reg[9][6]  ( .CLK(N446), .D(n11), .Q(\mem[9][6] ) );
  LATCHX1_HVT \mem_reg[9][5]  ( .CLK(N445), .D(n11), .Q(\mem[9][5] ) );
  LATCHX1_HVT \mem_reg[9][4]  ( .CLK(N444), .D(n11), .Q(\mem[9][4] ) );
  LATCHX1_HVT \mem_reg[9][3]  ( .CLK(N443), .D(n11), .Q(\mem[9][3] ) );
  LATCHX1_HVT \mem_reg[9][2]  ( .CLK(N442), .D(n11), .Q(\mem[9][2] ) );
  LATCHX1_HVT \mem_reg[9][1]  ( .CLK(N441), .D(n11), .Q(\mem[9][1] ) );
  LATCHX1_HVT \mem_reg[9][0]  ( .CLK(N440), .D(n11), .Q(\mem[9][0] ) );
  LATCHX1_HVT \mem_reg[8][15]  ( .CLK(N439), .D(n15), .Q(\mem[8][15] ) );
  LATCHX1_HVT \mem_reg[8][14]  ( .CLK(N438), .D(n15), .Q(\mem[8][14] ) );
  LATCHX1_HVT \mem_reg[8][13]  ( .CLK(N437), .D(n15), .Q(\mem[8][13] ) );
  LATCHX1_HVT \mem_reg[8][12]  ( .CLK(N436), .D(n15), .Q(\mem[8][12] ) );
  LATCHX1_HVT \mem_reg[8][11]  ( .CLK(N435), .D(n15), .Q(\mem[8][11] ) );
  LATCHX1_HVT \mem_reg[8][10]  ( .CLK(N434), .D(n16), .Q(\mem[8][10] ) );
  LATCHX1_HVT \mem_reg[8][9]  ( .CLK(N433), .D(n16), .Q(\mem[8][9] ) );
  LATCHX1_HVT \mem_reg[8][8]  ( .CLK(N432), .D(n16), .Q(\mem[8][8] ) );
  LATCHX1_HVT \mem_reg[8][7]  ( .CLK(N431), .D(n16), .Q(\mem[8][7] ) );
  LATCHX1_HVT \mem_reg[8][6]  ( .CLK(N430), .D(n16), .Q(\mem[8][6] ) );
  LATCHX1_HVT \mem_reg[8][5]  ( .CLK(N429), .D(n16), .Q(\mem[8][5] ) );
  LATCHX1_HVT \mem_reg[8][4]  ( .CLK(N428), .D(n16), .Q(\mem[8][4] ) );
  LATCHX1_HVT \mem_reg[8][3]  ( .CLK(N427), .D(n16), .Q(\mem[8][3] ) );
  LATCHX1_HVT \mem_reg[8][2]  ( .CLK(N426), .D(n16), .Q(\mem[8][2] ) );
  LATCHX1_HVT \mem_reg[8][1]  ( .CLK(N425), .D(n16), .Q(\mem[8][1] ) );
  LATCHX1_HVT \mem_reg[8][0]  ( .CLK(N424), .D(n16), .Q(\mem[8][0] ) );
  LATCHX1_HVT \mem_reg[7][15]  ( .CLK(N423), .D(n6), .Q(\mem[7][15] ) );
  LATCHX1_HVT \mem_reg[7][14]  ( .CLK(N422), .D(n1), .Q(\mem[7][14] ) );
  LATCHX1_HVT \mem_reg[7][13]  ( .CLK(N421), .D(n1), .Q(\mem[7][13] ) );
  LATCHX1_HVT \mem_reg[7][12]  ( .CLK(N420), .D(n1), .Q(\mem[7][12] ) );
  LATCHX1_HVT \mem_reg[7][11]  ( .CLK(N419), .D(n1), .Q(\mem[7][11] ) );
  LATCHX1_HVT \mem_reg[7][10]  ( .CLK(N418), .D(n1), .Q(\mem[7][10] ) );
  LATCHX1_HVT \mem_reg[7][9]  ( .CLK(N417), .D(n1), .Q(\mem[7][9] ) );
  LATCHX1_HVT \mem_reg[7][8]  ( .CLK(N416), .D(n1), .Q(\mem[7][8] ) );
  LATCHX1_HVT \mem_reg[7][7]  ( .CLK(N415), .D(n1), .Q(\mem[7][7] ) );
  LATCHX1_HVT \mem_reg[7][6]  ( .CLK(N414), .D(n1), .Q(\mem[7][6] ) );
  LATCHX1_HVT \mem_reg[7][5]  ( .CLK(N413), .D(n1), .Q(\mem[7][5] ) );
  LATCHX1_HVT \mem_reg[7][4]  ( .CLK(N412), .D(n1), .Q(\mem[7][4] ) );
  LATCHX1_HVT \mem_reg[7][3]  ( .CLK(N411), .D(n2), .Q(\mem[7][3] ) );
  LATCHX1_HVT \mem_reg[7][2]  ( .CLK(N410), .D(n2), .Q(\mem[7][2] ) );
  LATCHX1_HVT \mem_reg[7][1]  ( .CLK(N409), .D(n2), .Q(\mem[7][1] ) );
  LATCHX1_HVT \mem_reg[7][0]  ( .CLK(N408), .D(n2), .Q(\mem[7][0] ) );
  LATCHX1_HVT \mem_reg[6][15]  ( .CLK(N407), .D(n16), .Q(\mem[6][15] ) );
  LATCHX1_HVT \mem_reg[6][14]  ( .CLK(N406), .D(n17), .Q(\mem[6][14] ) );
  LATCHX1_HVT \mem_reg[6][13]  ( .CLK(N405), .D(n17), .Q(\mem[6][13] ) );
  LATCHX1_HVT \mem_reg[6][12]  ( .CLK(N404), .D(n17), .Q(\mem[6][12] ) );
  LATCHX1_HVT \mem_reg[6][11]  ( .CLK(N403), .D(n17), .Q(\mem[6][11] ) );
  LATCHX1_HVT \mem_reg[6][10]  ( .CLK(N402), .D(n17), .Q(\mem[6][10] ) );
  LATCHX1_HVT \mem_reg[6][9]  ( .CLK(N401), .D(n17), .Q(\mem[6][9] ) );
  LATCHX1_HVT \mem_reg[6][8]  ( .CLK(N400), .D(n17), .Q(\mem[6][8] ) );
  LATCHX1_HVT \mem_reg[6][7]  ( .CLK(N399), .D(n17), .Q(\mem[6][7] ) );
  LATCHX1_HVT \mem_reg[6][6]  ( .CLK(N398), .D(n17), .Q(\mem[6][6] ) );
  LATCHX1_HVT \mem_reg[6][5]  ( .CLK(N397), .D(n17), .Q(\mem[6][5] ) );
  LATCHX1_HVT \mem_reg[6][4]  ( .CLK(N396), .D(n18), .Q(\mem[6][4] ) );
  LATCHX1_HVT \mem_reg[6][3]  ( .CLK(N395), .D(n17), .Q(\mem[6][3] ) );
  LATCHX1_HVT \mem_reg[6][2]  ( .CLK(N394), .D(n18), .Q(\mem[6][2] ) );
  LATCHX1_HVT \mem_reg[6][1]  ( .CLK(N393), .D(n18), .Q(\mem[6][1] ) );
  LATCHX1_HVT \mem_reg[6][0]  ( .CLK(N392), .D(n18), .Q(\mem[6][0] ) );
  LATCHX1_HVT \mem_reg[5][15]  ( .CLK(N391), .D(n2), .Q(\mem[5][15] ) );
  LATCHX1_HVT \mem_reg[5][14]  ( .CLK(N390), .D(n2), .Q(\mem[5][14] ) );
  LATCHX1_HVT \mem_reg[5][13]  ( .CLK(N389), .D(n2), .Q(\mem[5][13] ) );
  LATCHX1_HVT \mem_reg[5][12]  ( .CLK(N388), .D(n2), .Q(\mem[5][12] ) );
  LATCHX1_HVT \mem_reg[5][11]  ( .CLK(N387), .D(n2), .Q(\mem[5][11] ) );
  LATCHX1_HVT \mem_reg[5][10]  ( .CLK(N386), .D(n2), .Q(\mem[5][10] ) );
  LATCHX1_HVT \mem_reg[5][9]  ( .CLK(N385), .D(n2), .Q(\mem[5][9] ) );
  LATCHX1_HVT \mem_reg[5][8]  ( .CLK(N384), .D(n2), .Q(\mem[5][8] ) );
  LATCHX1_HVT \mem_reg[5][7]  ( .CLK(N383), .D(n3), .Q(\mem[5][7] ) );
  LATCHX1_HVT \mem_reg[5][6]  ( .CLK(N382), .D(n3), .Q(\mem[5][6] ) );
  LATCHX1_HVT \mem_reg[5][5]  ( .CLK(N381), .D(n3), .Q(\mem[5][5] ) );
  LATCHX1_HVT \mem_reg[5][4]  ( .CLK(N380), .D(n3), .Q(\mem[5][4] ) );
  LATCHX1_HVT \mem_reg[5][3]  ( .CLK(N379), .D(n3), .Q(\mem[5][3] ) );
  LATCHX1_HVT \mem_reg[5][2]  ( .CLK(N378), .D(n3), .Q(\mem[5][2] ) );
  LATCHX1_HVT \mem_reg[5][1]  ( .CLK(N377), .D(n3), .Q(\mem[5][1] ) );
  LATCHX1_HVT \mem_reg[5][0]  ( .CLK(N376), .D(n3), .Q(\mem[5][0] ) );
  LATCHX1_HVT \mem_reg[4][15]  ( .CLK(N375), .D(n18), .Q(\mem[4][15] ) );
  LATCHX1_HVT \mem_reg[4][14]  ( .CLK(N374), .D(n18), .Q(\mem[4][14] ) );
  LATCHX1_HVT \mem_reg[4][13]  ( .CLK(N373), .D(n18), .Q(\mem[4][13] ) );
  LATCHX1_HVT \mem_reg[4][12]  ( .CLK(N372), .D(n18), .Q(\mem[4][12] ) );
  LATCHX1_HVT \mem_reg[4][11]  ( .CLK(N371), .D(n18), .Q(\mem[4][11] ) );
  LATCHX1_HVT \mem_reg[4][10]  ( .CLK(N370), .D(n18), .Q(\mem[4][10] ) );
  LATCHX1_HVT \mem_reg[4][9]  ( .CLK(N369), .D(n18), .Q(\mem[4][9] ) );
  LATCHX1_HVT \mem_reg[4][8]  ( .CLK(N368), .D(n19), .Q(\mem[4][8] ) );
  LATCHX1_HVT \mem_reg[4][7]  ( .CLK(N367), .D(n18), .Q(\mem[4][7] ) );
  LATCHX1_HVT \mem_reg[4][6]  ( .CLK(N366), .D(n19), .Q(\mem[4][6] ) );
  LATCHX1_HVT \mem_reg[4][5]  ( .CLK(N365), .D(n19), .Q(\mem[4][5] ) );
  LATCHX1_HVT \mem_reg[4][4]  ( .CLK(N364), .D(n19), .Q(\mem[4][4] ) );
  LATCHX1_HVT \mem_reg[4][3]  ( .CLK(N363), .D(n19), .Q(\mem[4][3] ) );
  LATCHX1_HVT \mem_reg[4][2]  ( .CLK(N362), .D(n19), .Q(\mem[4][2] ) );
  LATCHX1_HVT \mem_reg[4][1]  ( .CLK(N361), .D(n19), .Q(\mem[4][1] ) );
  LATCHX1_HVT \mem_reg[4][0]  ( .CLK(N360), .D(n19), .Q(\mem[4][0] ) );
  LATCHX1_HVT \mem_reg[3][15]  ( .CLK(N359), .D(n3), .Q(\mem[3][15] ) );
  LATCHX1_HVT \mem_reg[3][14]  ( .CLK(N358), .D(n3), .Q(\mem[3][14] ) );
  LATCHX1_HVT \mem_reg[3][13]  ( .CLK(N357), .D(n3), .Q(\mem[3][13] ) );
  LATCHX1_HVT \mem_reg[3][12]  ( .CLK(N356), .D(n3), .Q(\mem[3][12] ) );
  LATCHX1_HVT \mem_reg[3][11]  ( .CLK(N355), .D(n4), .Q(\mem[3][11] ) );
  LATCHX1_HVT \mem_reg[3][10]  ( .CLK(N354), .D(n4), .Q(\mem[3][10] ) );
  LATCHX1_HVT \mem_reg[3][9]  ( .CLK(N353), .D(n4), .Q(\mem[3][9] ) );
  LATCHX1_HVT \mem_reg[3][8]  ( .CLK(N352), .D(n4), .Q(\mem[3][8] ) );
  LATCHX1_HVT \mem_reg[3][7]  ( .CLK(N351), .D(n4), .Q(\mem[3][7] ) );
  LATCHX1_HVT \mem_reg[3][6]  ( .CLK(N350), .D(n4), .Q(\mem[3][6] ) );
  LATCHX1_HVT \mem_reg[3][5]  ( .CLK(N349), .D(n4), .Q(\mem[3][5] ) );
  LATCHX1_HVT \mem_reg[3][4]  ( .CLK(N348), .D(n4), .Q(\mem[3][4] ) );
  LATCHX1_HVT \mem_reg[3][3]  ( .CLK(N347), .D(n4), .Q(\mem[3][3] ) );
  LATCHX1_HVT \mem_reg[3][2]  ( .CLK(N346), .D(n4), .Q(\mem[3][2] ) );
  LATCHX1_HVT \mem_reg[3][1]  ( .CLK(N345), .D(n4), .Q(\mem[3][1] ) );
  LATCHX1_HVT \mem_reg[3][0]  ( .CLK(N344), .D(n4), .Q(\mem[3][0] ) );
  LATCHX1_HVT \mem_reg[2][15]  ( .CLK(N343), .D(n19), .Q(\mem[2][15] ) );
  LATCHX1_HVT \mem_reg[2][14]  ( .CLK(N342), .D(n19), .Q(\mem[2][14] ) );
  LATCHX1_HVT \mem_reg[2][13]  ( .CLK(N341), .D(n19), .Q(\mem[2][13] ) );
  LATCHX1_HVT \mem_reg[2][12]  ( .CLK(N340), .D(n20), .Q(\mem[2][12] ) );
  LATCHX1_HVT \mem_reg[2][11]  ( .CLK(N339), .D(n19), .Q(\mem[2][11] ) );
  LATCHX1_HVT \mem_reg[2][10]  ( .CLK(N338), .D(n20), .Q(\mem[2][10] ) );
  LATCHX1_HVT \mem_reg[2][9]  ( .CLK(N337), .D(n20), .Q(\mem[2][9] ) );
  LATCHX1_HVT \mem_reg[2][8]  ( .CLK(N336), .D(n20), .Q(\mem[2][8] ) );
  LATCHX1_HVT \mem_reg[2][7]  ( .CLK(N335), .D(n20), .Q(\mem[2][7] ) );
  LATCHX1_HVT \mem_reg[2][6]  ( .CLK(N334), .D(n20), .Q(\mem[2][6] ) );
  LATCHX1_HVT \mem_reg[2][5]  ( .CLK(N333), .D(n20), .Q(\mem[2][5] ) );
  LATCHX1_HVT \mem_reg[2][4]  ( .CLK(N332), .D(n20), .Q(\mem[2][4] ) );
  LATCHX1_HVT \mem_reg[2][3]  ( .CLK(N331), .D(n20), .Q(\mem[2][3] ) );
  LATCHX1_HVT \mem_reg[2][2]  ( .CLK(N330), .D(n20), .Q(\mem[2][2] ) );
  LATCHX1_HVT \mem_reg[2][1]  ( .CLK(N329), .D(n20), .Q(\mem[2][1] ) );
  LATCHX1_HVT \mem_reg[2][0]  ( .CLK(N328), .D(n21), .Q(\mem[2][0] ) );
  LATCHX1_HVT \mem_reg[1][15]  ( .CLK(N327), .D(n5), .Q(\mem[1][15] ) );
  LATCHX1_HVT \mem_reg[1][14]  ( .CLK(N326), .D(n5), .Q(\mem[1][14] ) );
  LATCHX1_HVT \mem_reg[1][13]  ( .CLK(N325), .D(n5), .Q(\mem[1][13] ) );
  LATCHX1_HVT \mem_reg[1][12]  ( .CLK(N324), .D(n5), .Q(\mem[1][12] ) );
  LATCHX1_HVT \mem_reg[1][11]  ( .CLK(N323), .D(n5), .Q(\mem[1][11] ) );
  LATCHX1_HVT \mem_reg[1][10]  ( .CLK(N322), .D(n5), .Q(\mem[1][10] ) );
  LATCHX1_HVT \mem_reg[1][9]  ( .CLK(N321), .D(n5), .Q(\mem[1][9] ) );
  LATCHX1_HVT \mem_reg[1][8]  ( .CLK(N320), .D(n5), .Q(\mem[1][8] ) );
  LATCHX1_HVT \mem_reg[1][7]  ( .CLK(N319), .D(n5), .Q(\mem[1][7] ) );
  LATCHX1_HVT \mem_reg[1][6]  ( .CLK(N318), .D(n5), .Q(\mem[1][6] ) );
  LATCHX1_HVT \mem_reg[1][5]  ( .CLK(N317), .D(n5), .Q(\mem[1][5] ) );
  LATCHX1_HVT \mem_reg[1][4]  ( .CLK(N316), .D(n5), .Q(\mem[1][4] ) );
  LATCHX1_HVT \mem_reg[1][3]  ( .CLK(N315), .D(n6), .Q(\mem[1][3] ) );
  LATCHX1_HVT \mem_reg[1][2]  ( .CLK(N314), .D(n6), .Q(\mem[1][2] ) );
  LATCHX1_HVT \mem_reg[1][1]  ( .CLK(N313), .D(n6), .Q(\mem[1][1] ) );
  LATCHX1_HVT \mem_reg[1][0]  ( .CLK(N312), .D(n6), .Q(\mem[1][0] ) );
  LATCHX1_HVT \mem_reg[0][15]  ( .CLK(N311), .D(n20), .Q(\mem[0][15] ) );
  LATCHX1_HVT \mem_reg[0][14]  ( .CLK(N310), .D(n21), .Q(\mem[0][14] ) );
  LATCHX1_HVT \mem_reg[0][13]  ( .CLK(N309), .D(n21), .Q(\mem[0][13] ) );
  LATCHX1_HVT \mem_reg[0][12]  ( .CLK(N308), .D(n21), .Q(\mem[0][12] ) );
  LATCHX1_HVT \mem_reg[0][11]  ( .CLK(N307), .D(n21), .Q(\mem[0][11] ) );
  LATCHX1_HVT \mem_reg[0][10]  ( .CLK(N306), .D(n21), .Q(\mem[0][10] ) );
  LATCHX1_HVT \mem_reg[0][9]  ( .CLK(N305), .D(n21), .Q(\mem[0][9] ) );
  LATCHX1_HVT \mem_reg[0][8]  ( .CLK(N304), .D(n21), .Q(\mem[0][8] ) );
  LATCHX1_HVT \mem_reg[0][7]  ( .CLK(N303), .D(n21), .Q(\mem[0][7] ) );
  LATCHX1_HVT \mem_reg[0][6]  ( .CLK(N302), .D(n21), .Q(\mem[0][6] ) );
  LATCHX1_HVT \mem_reg[0][5]  ( .CLK(N301), .D(n21), .Q(\mem[0][5] ) );
  LATCHX1_HVT \mem_reg[0][4]  ( .CLK(N300), .D(N495), .Q(\mem[0][4] ) );
  LATCHX1_HVT \mem_reg[0][3]  ( .CLK(N299), .D(n21), .Q(\mem[0][3] ) );
  LATCHX1_HVT \mem_reg[0][2]  ( .CLK(N298), .D(N495), .Q(\mem[0][2] ) );
  LATCHX1_HVT \mem_reg[0][1]  ( .CLK(N297), .D(N495), .Q(\mem[0][1] ) );
  LATCHX1_HVT \mem_reg[0][0]  ( .CLK(N296), .D(N495), .Q(\mem[0][0] ) );
  INVX1_HVT U3 ( .A(n23), .Y(n5) );
  INVX1_HVT U4 ( .A(n22), .Y(n21) );
  INVX1_HVT U5 ( .A(n22), .Y(n20) );
  INVX1_HVT U6 ( .A(n22), .Y(n4) );
  INVX1_HVT U7 ( .A(n22), .Y(n19) );
  INVX1_HVT U8 ( .A(n23), .Y(n3) );
  INVX1_HVT U9 ( .A(n22), .Y(n18) );
  INVX1_HVT U10 ( .A(n22), .Y(n2) );
  INVX1_HVT U11 ( .A(n23), .Y(n16) );
  INVX1_HVT U12 ( .A(n23), .Y(n15) );
  INVX1_HVT U13 ( .A(n22), .Y(n10) );
  INVX1_HVT U14 ( .A(n23), .Y(n9) );
  INVX1_HVT U15 ( .A(n23), .Y(n14) );
  INVX1_HVT U16 ( .A(n23), .Y(n13) );
  INVX1_HVT U17 ( .A(n22), .Y(n8) );
  INVX1_HVT U18 ( .A(n23), .Y(n12) );
  INVX1_HVT U19 ( .A(n22), .Y(n17) );
  INVX1_HVT U20 ( .A(n22), .Y(n1) );
  INVX1_HVT U21 ( .A(n23), .Y(n7) );
  INVX1_HVT U22 ( .A(n23), .Y(n11) );
  INVX1_HVT U23 ( .A(n22), .Y(n6) );
  INVX1_HVT U24 ( .A(N495), .Y(n22) );
  INVX1_HVT U25 ( .A(N495), .Y(n23) );
  MUX41X1_HVT U26 ( .A1(\mem[12][0] ), .A3(\mem[14][0] ), .A2(\mem[13][0] ), 
        .A4(\mem[15][0] ), .S0(N18), .S1(N17), .Y(n24) );
  MUX41X1_HVT U27 ( .A1(\mem[8][0] ), .A3(\mem[10][0] ), .A2(\mem[9][0] ), 
        .A4(\mem[11][0] ), .S0(N18), .S1(N17), .Y(n25) );
  MUX41X1_HVT U28 ( .A1(\mem[4][0] ), .A3(\mem[6][0] ), .A2(\mem[5][0] ), .A4(
        \mem[7][0] ), .S0(N18), .S1(N17), .Y(n26) );
  MUX41X1_HVT U29 ( .A1(\mem[0][0] ), .A3(\mem[2][0] ), .A2(\mem[1][0] ), .A4(
        \mem[3][0] ), .S0(N18), .S1(N17), .Y(n27) );
  MUX41X1_HVT U30 ( .A1(n27), .A3(n25), .A2(n26), .A4(n24), .S0(N20), .S1(N19), 
        .Y(N295) );
  MUX41X1_HVT U31 ( .A1(\mem[12][1] ), .A3(\mem[14][1] ), .A2(\mem[13][1] ), 
        .A4(\mem[15][1] ), .S0(N18), .S1(N17), .Y(n28) );
  MUX41X1_HVT U32 ( .A1(\mem[8][1] ), .A3(\mem[10][1] ), .A2(\mem[9][1] ), 
        .A4(\mem[11][1] ), .S0(N18), .S1(N17), .Y(n29) );
  MUX41X1_HVT U33 ( .A1(\mem[4][1] ), .A3(\mem[6][1] ), .A2(\mem[5][1] ), .A4(
        \mem[7][1] ), .S0(N18), .S1(N17), .Y(n30) );
  MUX41X1_HVT U34 ( .A1(\mem[0][1] ), .A3(\mem[2][1] ), .A2(\mem[1][1] ), .A4(
        \mem[3][1] ), .S0(N18), .S1(N17), .Y(n31) );
  MUX41X1_HVT U35 ( .A1(n31), .A3(n29), .A2(n30), .A4(n28), .S0(N20), .S1(N19), 
        .Y(N294) );
  MUX41X1_HVT U36 ( .A1(\mem[12][2] ), .A3(\mem[14][2] ), .A2(\mem[13][2] ), 
        .A4(\mem[15][2] ), .S0(N18), .S1(N17), .Y(n32) );
  MUX41X1_HVT U37 ( .A1(\mem[8][2] ), .A3(\mem[10][2] ), .A2(\mem[9][2] ), 
        .A4(\mem[11][2] ), .S0(N18), .S1(N17), .Y(n33) );
  MUX41X1_HVT U38 ( .A1(\mem[4][2] ), .A3(\mem[6][2] ), .A2(\mem[5][2] ), .A4(
        \mem[7][2] ), .S0(N18), .S1(N17), .Y(n34) );
  MUX41X1_HVT U39 ( .A1(\mem[0][2] ), .A3(\mem[2][2] ), .A2(\mem[1][2] ), .A4(
        \mem[3][2] ), .S0(N18), .S1(N17), .Y(n35) );
  MUX41X1_HVT U40 ( .A1(n35), .A3(n33), .A2(n34), .A4(n32), .S0(N20), .S1(N19), 
        .Y(N293) );
  MUX41X1_HVT U41 ( .A1(\mem[12][3] ), .A3(\mem[14][3] ), .A2(\mem[13][3] ), 
        .A4(\mem[15][3] ), .S0(N18), .S1(N17), .Y(n36) );
  MUX41X1_HVT U42 ( .A1(\mem[8][3] ), .A3(\mem[10][3] ), .A2(\mem[9][3] ), 
        .A4(\mem[11][3] ), .S0(N18), .S1(N17), .Y(n37) );
  MUX41X1_HVT U43 ( .A1(\mem[4][3] ), .A3(\mem[6][3] ), .A2(\mem[5][3] ), .A4(
        \mem[7][3] ), .S0(N18), .S1(N17), .Y(n38) );
  MUX41X1_HVT U44 ( .A1(\mem[0][3] ), .A3(\mem[2][3] ), .A2(\mem[1][3] ), .A4(
        \mem[3][3] ), .S0(N18), .S1(N17), .Y(n39) );
  MUX41X1_HVT U45 ( .A1(n39), .A3(n37), .A2(n38), .A4(n36), .S0(N20), .S1(N19), 
        .Y(N292) );
  MUX41X1_HVT U46 ( .A1(\mem[12][4] ), .A3(\mem[14][4] ), .A2(\mem[13][4] ), 
        .A4(\mem[15][4] ), .S0(N18), .S1(N17), .Y(n40) );
  MUX41X1_HVT U47 ( .A1(\mem[8][4] ), .A3(\mem[10][4] ), .A2(\mem[9][4] ), 
        .A4(\mem[11][4] ), .S0(N18), .S1(N17), .Y(n41) );
  MUX41X1_HVT U48 ( .A1(\mem[4][4] ), .A3(\mem[6][4] ), .A2(\mem[5][4] ), .A4(
        \mem[7][4] ), .S0(N18), .S1(N17), .Y(n42) );
  MUX41X1_HVT U49 ( .A1(\mem[0][4] ), .A3(\mem[2][4] ), .A2(\mem[1][4] ), .A4(
        \mem[3][4] ), .S0(N18), .S1(N17), .Y(n43) );
  MUX41X1_HVT U50 ( .A1(n43), .A3(n41), .A2(n42), .A4(n40), .S0(N20), .S1(N19), 
        .Y(N291) );
  MUX41X1_HVT U51 ( .A1(\mem[12][5] ), .A3(\mem[14][5] ), .A2(\mem[13][5] ), 
        .A4(\mem[15][5] ), .S0(N18), .S1(N17), .Y(n44) );
  MUX41X1_HVT U52 ( .A1(\mem[8][5] ), .A3(\mem[10][5] ), .A2(\mem[9][5] ), 
        .A4(\mem[11][5] ), .S0(N18), .S1(N17), .Y(n45) );
  MUX41X1_HVT U53 ( .A1(\mem[4][5] ), .A3(\mem[6][5] ), .A2(\mem[5][5] ), .A4(
        \mem[7][5] ), .S0(N18), .S1(N17), .Y(n46) );
  MUX41X1_HVT U54 ( .A1(\mem[0][5] ), .A3(\mem[2][5] ), .A2(\mem[1][5] ), .A4(
        \mem[3][5] ), .S0(N18), .S1(N17), .Y(n47) );
  MUX41X1_HVT U55 ( .A1(n47), .A3(n45), .A2(n46), .A4(n44), .S0(N20), .S1(N19), 
        .Y(N290) );
  MUX41X1_HVT U56 ( .A1(\mem[12][6] ), .A3(\mem[14][6] ), .A2(\mem[13][6] ), 
        .A4(\mem[15][6] ), .S0(N18), .S1(N17), .Y(n48) );
  MUX41X1_HVT U57 ( .A1(\mem[8][6] ), .A3(\mem[10][6] ), .A2(\mem[9][6] ), 
        .A4(\mem[11][6] ), .S0(N18), .S1(N17), .Y(n49) );
  MUX41X1_HVT U58 ( .A1(\mem[4][6] ), .A3(\mem[6][6] ), .A2(\mem[5][6] ), .A4(
        \mem[7][6] ), .S0(N18), .S1(N17), .Y(n50) );
  MUX41X1_HVT U59 ( .A1(\mem[0][6] ), .A3(\mem[2][6] ), .A2(\mem[1][6] ), .A4(
        \mem[3][6] ), .S0(N18), .S1(N17), .Y(n51) );
  MUX41X1_HVT U60 ( .A1(n51), .A3(n49), .A2(n50), .A4(n48), .S0(N20), .S1(N19), 
        .Y(N289) );
  MUX41X1_HVT U61 ( .A1(\mem[12][7] ), .A3(\mem[14][7] ), .A2(\mem[13][7] ), 
        .A4(\mem[15][7] ), .S0(N18), .S1(N17), .Y(n52) );
  MUX41X1_HVT U62 ( .A1(\mem[8][7] ), .A3(\mem[10][7] ), .A2(\mem[9][7] ), 
        .A4(\mem[11][7] ), .S0(N18), .S1(N17), .Y(n53) );
  MUX41X1_HVT U63 ( .A1(\mem[4][7] ), .A3(\mem[6][7] ), .A2(\mem[5][7] ), .A4(
        \mem[7][7] ), .S0(N18), .S1(N17), .Y(n54) );
  MUX41X1_HVT U64 ( .A1(\mem[0][7] ), .A3(\mem[2][7] ), .A2(\mem[1][7] ), .A4(
        \mem[3][7] ), .S0(N18), .S1(N17), .Y(n55) );
  MUX41X1_HVT U65 ( .A1(n55), .A3(n53), .A2(n54), .A4(n52), .S0(N20), .S1(N19), 
        .Y(N288) );
  MUX41X1_HVT U66 ( .A1(\mem[12][8] ), .A3(\mem[14][8] ), .A2(\mem[13][8] ), 
        .A4(\mem[15][8] ), .S0(N18), .S1(N17), .Y(n56) );
  MUX41X1_HVT U67 ( .A1(\mem[8][8] ), .A3(\mem[10][8] ), .A2(\mem[9][8] ), 
        .A4(\mem[11][8] ), .S0(N18), .S1(N17), .Y(n57) );
  MUX41X1_HVT U68 ( .A1(\mem[4][8] ), .A3(\mem[6][8] ), .A2(\mem[5][8] ), .A4(
        \mem[7][8] ), .S0(N18), .S1(N17), .Y(n58) );
  MUX41X1_HVT U69 ( .A1(\mem[0][8] ), .A3(\mem[2][8] ), .A2(\mem[1][8] ), .A4(
        \mem[3][8] ), .S0(N18), .S1(N17), .Y(n59) );
  MUX41X1_HVT U70 ( .A1(n59), .A3(n57), .A2(n58), .A4(n56), .S0(N20), .S1(N19), 
        .Y(N287) );
  MUX41X1_HVT U71 ( .A1(\mem[12][9] ), .A3(\mem[14][9] ), .A2(\mem[13][9] ), 
        .A4(\mem[15][9] ), .S0(N18), .S1(N17), .Y(n60) );
  MUX41X1_HVT U72 ( .A1(\mem[8][9] ), .A3(\mem[10][9] ), .A2(\mem[9][9] ), 
        .A4(\mem[11][9] ), .S0(N18), .S1(N17), .Y(n61) );
  MUX41X1_HVT U73 ( .A1(\mem[4][9] ), .A3(\mem[6][9] ), .A2(\mem[5][9] ), .A4(
        \mem[7][9] ), .S0(N18), .S1(N17), .Y(n78) );
  MUX41X1_HVT U74 ( .A1(\mem[0][9] ), .A3(\mem[2][9] ), .A2(\mem[1][9] ), .A4(
        \mem[3][9] ), .S0(N18), .S1(N17), .Y(n79) );
  MUX41X1_HVT U75 ( .A1(n79), .A3(n61), .A2(n78), .A4(n60), .S0(N20), .S1(N19), 
        .Y(N286) );
  MUX41X1_HVT U76 ( .A1(\mem[12][10] ), .A3(\mem[14][10] ), .A2(\mem[13][10] ), 
        .A4(\mem[15][10] ), .S0(N18), .S1(N17), .Y(n80) );
  MUX41X1_HVT U77 ( .A1(\mem[8][10] ), .A3(\mem[10][10] ), .A2(\mem[9][10] ), 
        .A4(\mem[11][10] ), .S0(N18), .S1(N17), .Y(n81) );
  MUX41X1_HVT U78 ( .A1(\mem[4][10] ), .A3(\mem[6][10] ), .A2(\mem[5][10] ), 
        .A4(\mem[7][10] ), .S0(N18), .S1(N17), .Y(n82) );
  MUX41X1_HVT U79 ( .A1(\mem[0][10] ), .A3(\mem[2][10] ), .A2(\mem[1][10] ), 
        .A4(\mem[3][10] ), .S0(N18), .S1(N17), .Y(n83) );
  MUX41X1_HVT U80 ( .A1(n83), .A3(n81), .A2(n82), .A4(n80), .S0(N20), .S1(N19), 
        .Y(N285) );
  MUX41X1_HVT U81 ( .A1(\mem[12][11] ), .A3(\mem[14][11] ), .A2(\mem[13][11] ), 
        .A4(\mem[15][11] ), .S0(N18), .S1(N17), .Y(n84) );
  MUX41X1_HVT U82 ( .A1(\mem[8][11] ), .A3(\mem[10][11] ), .A2(\mem[9][11] ), 
        .A4(\mem[11][11] ), .S0(N18), .S1(N17), .Y(n85) );
  MUX41X1_HVT U83 ( .A1(\mem[4][11] ), .A3(\mem[6][11] ), .A2(\mem[5][11] ), 
        .A4(\mem[7][11] ), .S0(N18), .S1(N17), .Y(n86) );
  MUX41X1_HVT U84 ( .A1(\mem[0][11] ), .A3(\mem[2][11] ), .A2(\mem[1][11] ), 
        .A4(\mem[3][11] ), .S0(N18), .S1(N17), .Y(n87) );
  MUX41X1_HVT U85 ( .A1(n87), .A3(n85), .A2(n86), .A4(n84), .S0(N20), .S1(N19), 
        .Y(N284) );
  MUX41X1_HVT U86 ( .A1(\mem[12][12] ), .A3(\mem[14][12] ), .A2(\mem[13][12] ), 
        .A4(\mem[15][12] ), .S0(N18), .S1(N17), .Y(n88) );
  MUX41X1_HVT U87 ( .A1(\mem[8][12] ), .A3(\mem[10][12] ), .A2(\mem[9][12] ), 
        .A4(\mem[11][12] ), .S0(N18), .S1(N17), .Y(n89) );
  MUX41X1_HVT U88 ( .A1(\mem[4][12] ), .A3(\mem[6][12] ), .A2(\mem[5][12] ), 
        .A4(\mem[7][12] ), .S0(N18), .S1(N17), .Y(n90) );
  MUX41X1_HVT U89 ( .A1(\mem[0][12] ), .A3(\mem[2][12] ), .A2(\mem[1][12] ), 
        .A4(\mem[3][12] ), .S0(N18), .S1(N17), .Y(n91) );
  MUX41X1_HVT U90 ( .A1(n91), .A3(n89), .A2(n90), .A4(n88), .S0(N20), .S1(N19), 
        .Y(N283) );
  MUX41X1_HVT U91 ( .A1(\mem[12][13] ), .A3(\mem[14][13] ), .A2(\mem[13][13] ), 
        .A4(\mem[15][13] ), .S0(N18), .S1(N17), .Y(n92) );
  MUX41X1_HVT U92 ( .A1(\mem[8][13] ), .A3(\mem[10][13] ), .A2(\mem[9][13] ), 
        .A4(\mem[11][13] ), .S0(N18), .S1(N17), .Y(n93) );
  MUX41X1_HVT U93 ( .A1(\mem[4][13] ), .A3(\mem[6][13] ), .A2(\mem[5][13] ), 
        .A4(\mem[7][13] ), .S0(N18), .S1(N17), .Y(n94) );
  MUX41X1_HVT U94 ( .A1(\mem[0][13] ), .A3(\mem[2][13] ), .A2(\mem[1][13] ), 
        .A4(\mem[3][13] ), .S0(N18), .S1(N17), .Y(n95) );
  MUX41X1_HVT U95 ( .A1(n95), .A3(n93), .A2(n94), .A4(n92), .S0(N20), .S1(N19), 
        .Y(N282) );
  MUX41X1_HVT U96 ( .A1(\mem[12][14] ), .A3(\mem[14][14] ), .A2(\mem[13][14] ), 
        .A4(\mem[15][14] ), .S0(N18), .S1(N17), .Y(n96) );
  MUX41X1_HVT U97 ( .A1(\mem[8][14] ), .A3(\mem[10][14] ), .A2(\mem[9][14] ), 
        .A4(\mem[11][14] ), .S0(N18), .S1(N17), .Y(n97) );
  MUX41X1_HVT U98 ( .A1(\mem[4][14] ), .A3(\mem[6][14] ), .A2(\mem[5][14] ), 
        .A4(\mem[7][14] ), .S0(N18), .S1(N17), .Y(n98) );
  MUX41X1_HVT U99 ( .A1(\mem[0][14] ), .A3(\mem[2][14] ), .A2(\mem[1][14] ), 
        .A4(\mem[3][14] ), .S0(N18), .S1(N17), .Y(n99) );
  MUX41X1_HVT U100 ( .A1(n99), .A3(n97), .A2(n98), .A4(n96), .S0(N20), .S1(N19), .Y(N281) );
  MUX41X1_HVT U101 ( .A1(\mem[12][15] ), .A3(\mem[14][15] ), .A2(\mem[13][15] ), .A4(\mem[15][15] ), .S0(N18), .S1(N17), .Y(n100) );
  MUX41X1_HVT U102 ( .A1(\mem[8][15] ), .A3(\mem[10][15] ), .A2(\mem[9][15] ), 
        .A4(\mem[11][15] ), .S0(N18), .S1(N17), .Y(n101) );
  MUX41X1_HVT U103 ( .A1(\mem[4][15] ), .A3(\mem[6][15] ), .A2(\mem[5][15] ), 
        .A4(\mem[7][15] ), .S0(N18), .S1(N17), .Y(n102) );
  MUX41X1_HVT U104 ( .A1(\mem[0][15] ), .A3(\mem[2][15] ), .A2(\mem[1][15] ), 
        .A4(\mem[3][15] ), .S0(N18), .S1(N17), .Y(n103) );
  MUX41X1_HVT U105 ( .A1(n103), .A3(n101), .A2(n102), .A4(n100), .S0(N20), 
        .S1(N19), .Y(N280) );
  MUX21X1_HVT U106 ( .A1(b_dout[15]), .A2(N280), .S0(n104), .Y(n162) );
  MUX21X1_HVT U107 ( .A1(b_dout[14]), .A2(N281), .S0(n104), .Y(n163) );
  MUX21X1_HVT U108 ( .A1(b_dout[13]), .A2(N282), .S0(n104), .Y(n164) );
  MUX21X1_HVT U109 ( .A1(b_dout[12]), .A2(N283), .S0(n104), .Y(n165) );
  MUX21X1_HVT U110 ( .A1(b_dout[11]), .A2(N284), .S0(n104), .Y(n166) );
  MUX21X1_HVT U111 ( .A1(b_dout[10]), .A2(N285), .S0(n104), .Y(n167) );
  MUX21X1_HVT U112 ( .A1(b_dout[9]), .A2(N286), .S0(n104), .Y(n168) );
  MUX21X1_HVT U113 ( .A1(b_dout[8]), .A2(N287), .S0(n104), .Y(n169) );
  MUX21X1_HVT U114 ( .A1(b_dout[7]), .A2(N288), .S0(n104), .Y(n170) );
  MUX21X1_HVT U115 ( .A1(b_dout[6]), .A2(N289), .S0(n104), .Y(n171) );
  MUX21X1_HVT U116 ( .A1(b_dout[5]), .A2(N290), .S0(n104), .Y(n172) );
  MUX21X1_HVT U117 ( .A1(b_dout[4]), .A2(N291), .S0(n104), .Y(n173) );
  MUX21X1_HVT U118 ( .A1(b_dout[3]), .A2(N292), .S0(n104), .Y(n174) );
  MUX21X1_HVT U119 ( .A1(b_dout[2]), .A2(N293), .S0(n104), .Y(n175) );
  MUX21X1_HVT U120 ( .A1(b_dout[1]), .A2(N294), .S0(n104), .Y(n176) );
  MUX21X1_HVT U121 ( .A1(b_dout[0]), .A2(N295), .S0(n104), .Y(n177) );
  NOR2X0_HVT U122 ( .A1(write), .A2(rst), .Y(n104) );
  AO21X1_HVT U123 ( .A1(n105), .A2(n106), .A3(rst), .Y(N552) );
  AO21X1_HVT U124 ( .A1(n107), .A2(n106), .A3(rst), .Y(N551) );
  AO21X1_HVT U125 ( .A1(n108), .A2(n106), .A3(rst), .Y(N550) );
  AO21X1_HVT U126 ( .A1(n109), .A2(n106), .A3(rst), .Y(N549) );
  AO21X1_HVT U127 ( .A1(n110), .A2(n106), .A3(rst), .Y(N548) );
  AO21X1_HVT U128 ( .A1(n111), .A2(n106), .A3(rst), .Y(N547) );
  AO21X1_HVT U129 ( .A1(n112), .A2(n106), .A3(rst), .Y(N546) );
  AO21X1_HVT U130 ( .A1(n113), .A2(n106), .A3(rst), .Y(N545) );
  AO21X1_HVT U131 ( .A1(n114), .A2(n106), .A3(rst), .Y(N544) );
  AO21X1_HVT U132 ( .A1(n115), .A2(n106), .A3(rst), .Y(N543) );
  AO21X1_HVT U133 ( .A1(n116), .A2(n106), .A3(rst), .Y(N542) );
  AO21X1_HVT U134 ( .A1(n117), .A2(n106), .A3(rst), .Y(N541) );
  AO21X1_HVT U135 ( .A1(n118), .A2(n106), .A3(rst), .Y(N540) );
  AO21X1_HVT U136 ( .A1(n119), .A2(n106), .A3(rst), .Y(N539) );
  AO21X1_HVT U137 ( .A1(n120), .A2(n106), .A3(rst), .Y(N538) );
  AO21X1_HVT U138 ( .A1(n121), .A2(n106), .A3(rst), .Y(N537) );
  AND2X1_HVT U139 ( .A1(n122), .A2(n123), .Y(n106) );
  AO21X1_HVT U140 ( .A1(n124), .A2(n105), .A3(rst), .Y(N536) );
  AO21X1_HVT U141 ( .A1(n124), .A2(n107), .A3(rst), .Y(N535) );
  AO21X1_HVT U142 ( .A1(n124), .A2(n108), .A3(rst), .Y(N534) );
  AO21X1_HVT U143 ( .A1(n124), .A2(n109), .A3(rst), .Y(N533) );
  AO21X1_HVT U144 ( .A1(n124), .A2(n110), .A3(rst), .Y(N532) );
  AO21X1_HVT U145 ( .A1(n124), .A2(n111), .A3(rst), .Y(N531) );
  AO21X1_HVT U146 ( .A1(n124), .A2(n112), .A3(rst), .Y(N530) );
  AO21X1_HVT U147 ( .A1(n124), .A2(n113), .A3(rst), .Y(N529) );
  AO21X1_HVT U148 ( .A1(n124), .A2(n114), .A3(rst), .Y(N528) );
  AO21X1_HVT U149 ( .A1(n124), .A2(n115), .A3(rst), .Y(N527) );
  AO21X1_HVT U150 ( .A1(n124), .A2(n116), .A3(rst), .Y(N526) );
  AO21X1_HVT U151 ( .A1(n124), .A2(n117), .A3(rst), .Y(N525) );
  AO21X1_HVT U152 ( .A1(n124), .A2(n118), .A3(rst), .Y(N524) );
  AO21X1_HVT U153 ( .A1(n124), .A2(n119), .A3(rst), .Y(N523) );
  AO21X1_HVT U154 ( .A1(n124), .A2(n120), .A3(rst), .Y(N522) );
  AO21X1_HVT U155 ( .A1(n124), .A2(n121), .A3(rst), .Y(N521) );
  AND2X1_HVT U156 ( .A1(n125), .A2(n123), .Y(n124) );
  AO21X1_HVT U157 ( .A1(n126), .A2(n105), .A3(rst), .Y(N520) );
  AO21X1_HVT U158 ( .A1(n126), .A2(n107), .A3(rst), .Y(N519) );
  AO21X1_HVT U159 ( .A1(n126), .A2(n108), .A3(rst), .Y(N518) );
  AO21X1_HVT U160 ( .A1(n126), .A2(n109), .A3(rst), .Y(N517) );
  AO21X1_HVT U161 ( .A1(n126), .A2(n110), .A3(rst), .Y(N516) );
  AO21X1_HVT U162 ( .A1(n126), .A2(n111), .A3(rst), .Y(N515) );
  AO21X1_HVT U163 ( .A1(n126), .A2(n112), .A3(rst), .Y(N514) );
  AO21X1_HVT U164 ( .A1(n126), .A2(n113), .A3(rst), .Y(N513) );
  AO21X1_HVT U165 ( .A1(n126), .A2(n114), .A3(rst), .Y(N512) );
  AO21X1_HVT U166 ( .A1(n126), .A2(n115), .A3(rst), .Y(N511) );
  AO21X1_HVT U167 ( .A1(n126), .A2(n116), .A3(rst), .Y(N510) );
  AO21X1_HVT U168 ( .A1(n126), .A2(n117), .A3(rst), .Y(N509) );
  AO21X1_HVT U169 ( .A1(n126), .A2(n118), .A3(rst), .Y(N508) );
  AO21X1_HVT U170 ( .A1(n126), .A2(n119), .A3(rst), .Y(N507) );
  AO21X1_HVT U171 ( .A1(n126), .A2(n120), .A3(rst), .Y(N506) );
  AO21X1_HVT U172 ( .A1(n126), .A2(n121), .A3(rst), .Y(N505) );
  AND2X1_HVT U173 ( .A1(n127), .A2(n122), .Y(n126) );
  AO21X1_HVT U174 ( .A1(n128), .A2(n105), .A3(rst), .Y(N504) );
  AO21X1_HVT U175 ( .A1(n128), .A2(n107), .A3(rst), .Y(N503) );
  AO21X1_HVT U176 ( .A1(n128), .A2(n108), .A3(rst), .Y(N502) );
  AO21X1_HVT U177 ( .A1(n128), .A2(n109), .A3(rst), .Y(N501) );
  AO21X1_HVT U178 ( .A1(n128), .A2(n110), .A3(rst), .Y(N500) );
  AO21X1_HVT U179 ( .A1(n128), .A2(n111), .A3(rst), .Y(N499) );
  AO21X1_HVT U180 ( .A1(n128), .A2(n112), .A3(rst), .Y(N498) );
  AO21X1_HVT U181 ( .A1(n128), .A2(n113), .A3(rst), .Y(N497) );
  AO21X1_HVT U182 ( .A1(n128), .A2(n114), .A3(rst), .Y(N496) );
  AO21X1_HVT U183 ( .A1(n128), .A2(n115), .A3(rst), .Y(N494) );
  AO21X1_HVT U184 ( .A1(n128), .A2(n116), .A3(rst), .Y(N493) );
  AO21X1_HVT U185 ( .A1(n128), .A2(n117), .A3(rst), .Y(N492) );
  AO21X1_HVT U186 ( .A1(n128), .A2(n118), .A3(rst), .Y(N491) );
  AO21X1_HVT U187 ( .A1(n128), .A2(n119), .A3(rst), .Y(N490) );
  AO21X1_HVT U188 ( .A1(n128), .A2(n120), .A3(rst), .Y(N489) );
  AO21X1_HVT U189 ( .A1(n128), .A2(n121), .A3(rst), .Y(N488) );
  AND2X1_HVT U190 ( .A1(n127), .A2(n125), .Y(n128) );
  AO21X1_HVT U191 ( .A1(n129), .A2(n105), .A3(rst), .Y(N487) );
  AO21X1_HVT U192 ( .A1(n129), .A2(n107), .A3(rst), .Y(N486) );
  AO21X1_HVT U193 ( .A1(n129), .A2(n108), .A3(rst), .Y(N485) );
  AO21X1_HVT U194 ( .A1(n129), .A2(n109), .A3(rst), .Y(N484) );
  AO21X1_HVT U195 ( .A1(n129), .A2(n110), .A3(rst), .Y(N483) );
  AO21X1_HVT U196 ( .A1(n129), .A2(n111), .A3(rst), .Y(N482) );
  AO21X1_HVT U197 ( .A1(n129), .A2(n112), .A3(rst), .Y(N481) );
  AO21X1_HVT U198 ( .A1(n129), .A2(n113), .A3(rst), .Y(N480) );
  AO21X1_HVT U199 ( .A1(n129), .A2(n114), .A3(rst), .Y(N479) );
  AO21X1_HVT U200 ( .A1(n129), .A2(n115), .A3(rst), .Y(N478) );
  AO21X1_HVT U201 ( .A1(n129), .A2(n116), .A3(rst), .Y(N477) );
  AO21X1_HVT U202 ( .A1(n129), .A2(n117), .A3(rst), .Y(N476) );
  AO21X1_HVT U203 ( .A1(n129), .A2(n118), .A3(rst), .Y(N475) );
  AO21X1_HVT U204 ( .A1(n129), .A2(n119), .A3(rst), .Y(N474) );
  AO21X1_HVT U205 ( .A1(n129), .A2(n120), .A3(rst), .Y(N473) );
  AO21X1_HVT U206 ( .A1(n129), .A2(n121), .A3(rst), .Y(N472) );
  AND2X1_HVT U207 ( .A1(n130), .A2(n122), .Y(n129) );
  AO21X1_HVT U208 ( .A1(n131), .A2(n105), .A3(rst), .Y(N471) );
  AO21X1_HVT U209 ( .A1(n131), .A2(n107), .A3(rst), .Y(N470) );
  AO21X1_HVT U210 ( .A1(n131), .A2(n108), .A3(rst), .Y(N469) );
  AO21X1_HVT U211 ( .A1(n131), .A2(n109), .A3(rst), .Y(N468) );
  AO21X1_HVT U212 ( .A1(n131), .A2(n110), .A3(rst), .Y(N467) );
  AO21X1_HVT U213 ( .A1(n131), .A2(n111), .A3(rst), .Y(N466) );
  AO21X1_HVT U214 ( .A1(n131), .A2(n112), .A3(rst), .Y(N465) );
  AO21X1_HVT U215 ( .A1(n131), .A2(n113), .A3(rst), .Y(N464) );
  AO21X1_HVT U216 ( .A1(n131), .A2(n114), .A3(rst), .Y(N463) );
  AO21X1_HVT U217 ( .A1(n131), .A2(n115), .A3(rst), .Y(N462) );
  AO21X1_HVT U218 ( .A1(n131), .A2(n116), .A3(rst), .Y(N461) );
  AO21X1_HVT U219 ( .A1(n131), .A2(n117), .A3(rst), .Y(N460) );
  AO21X1_HVT U220 ( .A1(n131), .A2(n118), .A3(rst), .Y(N459) );
  AO21X1_HVT U221 ( .A1(n131), .A2(n119), .A3(rst), .Y(N458) );
  AO21X1_HVT U222 ( .A1(n131), .A2(n120), .A3(rst), .Y(N457) );
  AO21X1_HVT U223 ( .A1(n131), .A2(n121), .A3(rst), .Y(N456) );
  AND2X1_HVT U224 ( .A1(n130), .A2(n125), .Y(n131) );
  AO21X1_HVT U225 ( .A1(n132), .A2(n105), .A3(rst), .Y(N455) );
  AO21X1_HVT U226 ( .A1(n132), .A2(n107), .A3(rst), .Y(N454) );
  AO21X1_HVT U227 ( .A1(n132), .A2(n108), .A3(rst), .Y(N453) );
  AO21X1_HVT U228 ( .A1(n132), .A2(n109), .A3(rst), .Y(N452) );
  AO21X1_HVT U229 ( .A1(n132), .A2(n110), .A3(rst), .Y(N451) );
  AO21X1_HVT U230 ( .A1(n132), .A2(n111), .A3(rst), .Y(N450) );
  AO21X1_HVT U231 ( .A1(n132), .A2(n112), .A3(rst), .Y(N449) );
  AO21X1_HVT U232 ( .A1(n132), .A2(n113), .A3(rst), .Y(N448) );
  AO21X1_HVT U233 ( .A1(n132), .A2(n114), .A3(rst), .Y(N447) );
  AO21X1_HVT U234 ( .A1(n132), .A2(n115), .A3(rst), .Y(N446) );
  AO21X1_HVT U235 ( .A1(n132), .A2(n116), .A3(rst), .Y(N445) );
  AO21X1_HVT U236 ( .A1(n132), .A2(n117), .A3(rst), .Y(N444) );
  AO21X1_HVT U237 ( .A1(n132), .A2(n118), .A3(rst), .Y(N443) );
  AO21X1_HVT U238 ( .A1(n132), .A2(n119), .A3(rst), .Y(N442) );
  AO21X1_HVT U239 ( .A1(n132), .A2(n120), .A3(rst), .Y(N441) );
  AO21X1_HVT U240 ( .A1(n132), .A2(n121), .A3(rst), .Y(N440) );
  AND2X1_HVT U241 ( .A1(n133), .A2(n122), .Y(n132) );
  AND3X1_HVT U242 ( .A1(a_din[0]), .A2(N495), .A3(a_din[3]), .Y(n122) );
  AO21X1_HVT U243 ( .A1(n134), .A2(n105), .A3(rst), .Y(N439) );
  AO21X1_HVT U244 ( .A1(n134), .A2(n107), .A3(rst), .Y(N438) );
  AO21X1_HVT U245 ( .A1(n134), .A2(n108), .A3(rst), .Y(N437) );
  AO21X1_HVT U246 ( .A1(n134), .A2(n109), .A3(rst), .Y(N436) );
  AO21X1_HVT U247 ( .A1(n134), .A2(n110), .A3(rst), .Y(N435) );
  AO21X1_HVT U248 ( .A1(n134), .A2(n111), .A3(rst), .Y(N434) );
  AO21X1_HVT U249 ( .A1(n134), .A2(n112), .A3(rst), .Y(N433) );
  AO21X1_HVT U250 ( .A1(n134), .A2(n113), .A3(rst), .Y(N432) );
  AO21X1_HVT U251 ( .A1(n134), .A2(n114), .A3(rst), .Y(N431) );
  AO21X1_HVT U252 ( .A1(n134), .A2(n115), .A3(rst), .Y(N430) );
  AO21X1_HVT U253 ( .A1(n134), .A2(n116), .A3(rst), .Y(N429) );
  AO21X1_HVT U254 ( .A1(n134), .A2(n117), .A3(rst), .Y(N428) );
  AO21X1_HVT U255 ( .A1(n134), .A2(n118), .A3(rst), .Y(N427) );
  AO21X1_HVT U256 ( .A1(n134), .A2(n119), .A3(rst), .Y(N426) );
  AO21X1_HVT U257 ( .A1(n134), .A2(n120), .A3(rst), .Y(N425) );
  AO21X1_HVT U258 ( .A1(n134), .A2(n121), .A3(rst), .Y(N424) );
  AND2X1_HVT U259 ( .A1(n133), .A2(n125), .Y(n134) );
  AND3X1_HVT U260 ( .A1(N495), .A2(n135), .A3(a_din[3]), .Y(n125) );
  AO21X1_HVT U261 ( .A1(n136), .A2(n105), .A3(rst), .Y(N423) );
  AO21X1_HVT U262 ( .A1(n136), .A2(n107), .A3(rst), .Y(N422) );
  AO21X1_HVT U263 ( .A1(n136), .A2(n108), .A3(rst), .Y(N421) );
  AO21X1_HVT U264 ( .A1(n136), .A2(n109), .A3(rst), .Y(N420) );
  AO21X1_HVT U265 ( .A1(n136), .A2(n110), .A3(rst), .Y(N419) );
  AO21X1_HVT U266 ( .A1(n136), .A2(n111), .A3(rst), .Y(N418) );
  AO21X1_HVT U267 ( .A1(n136), .A2(n112), .A3(rst), .Y(N417) );
  AO21X1_HVT U268 ( .A1(n136), .A2(n113), .A3(rst), .Y(N416) );
  AO21X1_HVT U269 ( .A1(n136), .A2(n114), .A3(rst), .Y(N415) );
  AO21X1_HVT U270 ( .A1(n136), .A2(n115), .A3(rst), .Y(N414) );
  AO21X1_HVT U271 ( .A1(n136), .A2(n116), .A3(rst), .Y(N413) );
  AO21X1_HVT U272 ( .A1(n136), .A2(n117), .A3(rst), .Y(N412) );
  AO21X1_HVT U273 ( .A1(n136), .A2(n118), .A3(rst), .Y(N411) );
  AO21X1_HVT U274 ( .A1(n136), .A2(n119), .A3(rst), .Y(N410) );
  AO21X1_HVT U275 ( .A1(n136), .A2(n120), .A3(rst), .Y(N409) );
  AO21X1_HVT U276 ( .A1(n136), .A2(n121), .A3(rst), .Y(N408) );
  AND2X1_HVT U277 ( .A1(n137), .A2(n123), .Y(n136) );
  AO21X1_HVT U278 ( .A1(n138), .A2(n105), .A3(rst), .Y(N407) );
  AO21X1_HVT U279 ( .A1(n138), .A2(n107), .A3(rst), .Y(N406) );
  AO21X1_HVT U280 ( .A1(n138), .A2(n108), .A3(rst), .Y(N405) );
  AO21X1_HVT U281 ( .A1(n138), .A2(n109), .A3(rst), .Y(N404) );
  AO21X1_HVT U282 ( .A1(n138), .A2(n110), .A3(rst), .Y(N403) );
  AO21X1_HVT U283 ( .A1(n138), .A2(n111), .A3(rst), .Y(N402) );
  AO21X1_HVT U284 ( .A1(n138), .A2(n112), .A3(rst), .Y(N401) );
  AO21X1_HVT U285 ( .A1(n138), .A2(n113), .A3(rst), .Y(N400) );
  AO21X1_HVT U286 ( .A1(n138), .A2(n114), .A3(rst), .Y(N399) );
  AO21X1_HVT U287 ( .A1(n138), .A2(n115), .A3(rst), .Y(N398) );
  AO21X1_HVT U288 ( .A1(n138), .A2(n116), .A3(rst), .Y(N397) );
  AO21X1_HVT U289 ( .A1(n138), .A2(n117), .A3(rst), .Y(N396) );
  AO21X1_HVT U290 ( .A1(n138), .A2(n118), .A3(rst), .Y(N395) );
  AO21X1_HVT U291 ( .A1(n138), .A2(n119), .A3(rst), .Y(N394) );
  AO21X1_HVT U292 ( .A1(n138), .A2(n120), .A3(rst), .Y(N393) );
  AO21X1_HVT U293 ( .A1(n138), .A2(n121), .A3(rst), .Y(N392) );
  AND2X1_HVT U294 ( .A1(n139), .A2(n123), .Y(n138) );
  AND2X1_HVT U295 ( .A1(a_din[2]), .A2(a_din[1]), .Y(n123) );
  AO21X1_HVT U296 ( .A1(n140), .A2(n105), .A3(rst), .Y(N391) );
  AO21X1_HVT U297 ( .A1(n140), .A2(n107), .A3(rst), .Y(N390) );
  AO21X1_HVT U298 ( .A1(n140), .A2(n108), .A3(rst), .Y(N389) );
  AO21X1_HVT U299 ( .A1(n140), .A2(n109), .A3(rst), .Y(N388) );
  AO21X1_HVT U300 ( .A1(n140), .A2(n110), .A3(rst), .Y(N387) );
  AO21X1_HVT U301 ( .A1(n140), .A2(n111), .A3(rst), .Y(N386) );
  AO21X1_HVT U302 ( .A1(n140), .A2(n112), .A3(rst), .Y(N385) );
  AO21X1_HVT U303 ( .A1(n140), .A2(n113), .A3(rst), .Y(N384) );
  AO21X1_HVT U304 ( .A1(n140), .A2(n114), .A3(rst), .Y(N383) );
  AO21X1_HVT U305 ( .A1(n140), .A2(n115), .A3(rst), .Y(N382) );
  AO21X1_HVT U306 ( .A1(n140), .A2(n116), .A3(rst), .Y(N381) );
  AO21X1_HVT U307 ( .A1(n140), .A2(n117), .A3(rst), .Y(N380) );
  AO21X1_HVT U308 ( .A1(n140), .A2(n118), .A3(rst), .Y(N379) );
  AO21X1_HVT U309 ( .A1(n140), .A2(n119), .A3(rst), .Y(N378) );
  AO21X1_HVT U310 ( .A1(n140), .A2(n120), .A3(rst), .Y(N377) );
  AO21X1_HVT U311 ( .A1(n140), .A2(n121), .A3(rst), .Y(N376) );
  AND2X1_HVT U312 ( .A1(n137), .A2(n127), .Y(n140) );
  AO21X1_HVT U313 ( .A1(n141), .A2(n105), .A3(rst), .Y(N375) );
  AO21X1_HVT U314 ( .A1(n141), .A2(n107), .A3(rst), .Y(N374) );
  AO21X1_HVT U315 ( .A1(n141), .A2(n108), .A3(rst), .Y(N373) );
  AO21X1_HVT U316 ( .A1(n141), .A2(n109), .A3(rst), .Y(N372) );
  AO21X1_HVT U317 ( .A1(n141), .A2(n110), .A3(rst), .Y(N371) );
  AO21X1_HVT U318 ( .A1(n141), .A2(n111), .A3(rst), .Y(N370) );
  AO21X1_HVT U319 ( .A1(n141), .A2(n112), .A3(rst), .Y(N369) );
  AO21X1_HVT U320 ( .A1(n141), .A2(n113), .A3(rst), .Y(N368) );
  AO21X1_HVT U321 ( .A1(n141), .A2(n114), .A3(rst), .Y(N367) );
  AO21X1_HVT U322 ( .A1(n141), .A2(n115), .A3(rst), .Y(N366) );
  AO21X1_HVT U323 ( .A1(n141), .A2(n116), .A3(rst), .Y(N365) );
  AO21X1_HVT U324 ( .A1(n141), .A2(n117), .A3(rst), .Y(N364) );
  AO21X1_HVT U325 ( .A1(n141), .A2(n118), .A3(rst), .Y(N363) );
  AO21X1_HVT U326 ( .A1(n141), .A2(n119), .A3(rst), .Y(N362) );
  AO21X1_HVT U327 ( .A1(n141), .A2(n120), .A3(rst), .Y(N361) );
  AO21X1_HVT U328 ( .A1(n141), .A2(n121), .A3(rst), .Y(N360) );
  AND2X1_HVT U329 ( .A1(n139), .A2(n127), .Y(n141) );
  AND2X1_HVT U330 ( .A1(a_din[2]), .A2(n142), .Y(n127) );
  AO21X1_HVT U331 ( .A1(n143), .A2(n105), .A3(rst), .Y(N359) );
  AO21X1_HVT U332 ( .A1(n143), .A2(n107), .A3(rst), .Y(N358) );
  AO21X1_HVT U333 ( .A1(n143), .A2(n108), .A3(rst), .Y(N357) );
  AO21X1_HVT U334 ( .A1(n143), .A2(n109), .A3(rst), .Y(N356) );
  AO21X1_HVT U335 ( .A1(n143), .A2(n110), .A3(rst), .Y(N355) );
  AO21X1_HVT U336 ( .A1(n143), .A2(n111), .A3(rst), .Y(N354) );
  AO21X1_HVT U337 ( .A1(n143), .A2(n112), .A3(rst), .Y(N353) );
  AO21X1_HVT U338 ( .A1(n143), .A2(n113), .A3(rst), .Y(N352) );
  AO21X1_HVT U339 ( .A1(n143), .A2(n114), .A3(rst), .Y(N351) );
  AO21X1_HVT U340 ( .A1(n143), .A2(n115), .A3(rst), .Y(N350) );
  AO21X1_HVT U341 ( .A1(n143), .A2(n116), .A3(rst), .Y(N349) );
  AO21X1_HVT U342 ( .A1(n143), .A2(n117), .A3(rst), .Y(N348) );
  AO21X1_HVT U343 ( .A1(n143), .A2(n118), .A3(rst), .Y(N347) );
  AO21X1_HVT U344 ( .A1(n143), .A2(n119), .A3(rst), .Y(N346) );
  AO21X1_HVT U345 ( .A1(n143), .A2(n120), .A3(rst), .Y(N345) );
  AO21X1_HVT U346 ( .A1(n143), .A2(n121), .A3(rst), .Y(N344) );
  AND2X1_HVT U347 ( .A1(n137), .A2(n130), .Y(n143) );
  AO21X1_HVT U348 ( .A1(n144), .A2(n105), .A3(rst), .Y(N343) );
  AO21X1_HVT U349 ( .A1(n144), .A2(n107), .A3(rst), .Y(N342) );
  AO21X1_HVT U350 ( .A1(n144), .A2(n108), .A3(rst), .Y(N341) );
  AO21X1_HVT U351 ( .A1(n144), .A2(n109), .A3(rst), .Y(N340) );
  AO21X1_HVT U352 ( .A1(n144), .A2(n110), .A3(rst), .Y(N339) );
  AO21X1_HVT U353 ( .A1(n144), .A2(n111), .A3(rst), .Y(N338) );
  AO21X1_HVT U354 ( .A1(n144), .A2(n112), .A3(rst), .Y(N337) );
  AO21X1_HVT U355 ( .A1(n144), .A2(n113), .A3(rst), .Y(N336) );
  AO21X1_HVT U356 ( .A1(n144), .A2(n114), .A3(rst), .Y(N335) );
  AO21X1_HVT U357 ( .A1(n144), .A2(n115), .A3(rst), .Y(N334) );
  AO21X1_HVT U358 ( .A1(n144), .A2(n116), .A3(rst), .Y(N333) );
  AO21X1_HVT U359 ( .A1(n144), .A2(n117), .A3(rst), .Y(N332) );
  AO21X1_HVT U360 ( .A1(n144), .A2(n118), .A3(rst), .Y(N331) );
  AO21X1_HVT U361 ( .A1(n144), .A2(n119), .A3(rst), .Y(N330) );
  AO21X1_HVT U362 ( .A1(n144), .A2(n120), .A3(rst), .Y(N329) );
  AO21X1_HVT U363 ( .A1(n144), .A2(n121), .A3(rst), .Y(N328) );
  AND2X1_HVT U364 ( .A1(n139), .A2(n130), .Y(n144) );
  AND2X1_HVT U365 ( .A1(a_din[1]), .A2(n145), .Y(n130) );
  AO21X1_HVT U366 ( .A1(n146), .A2(n105), .A3(rst), .Y(N327) );
  AO21X1_HVT U367 ( .A1(n146), .A2(n107), .A3(rst), .Y(N326) );
  AO21X1_HVT U368 ( .A1(n146), .A2(n108), .A3(rst), .Y(N325) );
  AO21X1_HVT U369 ( .A1(n146), .A2(n109), .A3(rst), .Y(N324) );
  AO21X1_HVT U370 ( .A1(n146), .A2(n110), .A3(rst), .Y(N323) );
  AO21X1_HVT U371 ( .A1(n146), .A2(n111), .A3(rst), .Y(N322) );
  AO21X1_HVT U372 ( .A1(n146), .A2(n112), .A3(rst), .Y(N321) );
  AO21X1_HVT U373 ( .A1(n146), .A2(n113), .A3(rst), .Y(N320) );
  AO21X1_HVT U374 ( .A1(n146), .A2(n114), .A3(rst), .Y(N319) );
  AO21X1_HVT U375 ( .A1(n146), .A2(n115), .A3(rst), .Y(N318) );
  AO21X1_HVT U376 ( .A1(n146), .A2(n116), .A3(rst), .Y(N317) );
  AO21X1_HVT U377 ( .A1(n146), .A2(n117), .A3(rst), .Y(N316) );
  AO21X1_HVT U378 ( .A1(n146), .A2(n118), .A3(rst), .Y(N315) );
  AO21X1_HVT U379 ( .A1(n146), .A2(n119), .A3(rst), .Y(N314) );
  AO21X1_HVT U380 ( .A1(n146), .A2(n120), .A3(rst), .Y(N313) );
  AO21X1_HVT U381 ( .A1(n146), .A2(n121), .A3(rst), .Y(N312) );
  AND2X1_HVT U382 ( .A1(n137), .A2(n133), .Y(n146) );
  AND3X1_HVT U383 ( .A1(N495), .A2(n147), .A3(a_din[0]), .Y(n137) );
  AO21X1_HVT U384 ( .A1(n148), .A2(n105), .A3(rst), .Y(N311) );
  AND2X1_HVT U385 ( .A1(n149), .A2(n150), .Y(n105) );
  AO21X1_HVT U386 ( .A1(n148), .A2(n107), .A3(rst), .Y(N310) );
  AND2X1_HVT U387 ( .A1(n151), .A2(n149), .Y(n107) );
  AO21X1_HVT U388 ( .A1(n148), .A2(n108), .A3(rst), .Y(N309) );
  AND2X1_HVT U389 ( .A1(n152), .A2(n149), .Y(n108) );
  AO21X1_HVT U390 ( .A1(n148), .A2(n109), .A3(rst), .Y(N308) );
  AND2X1_HVT U391 ( .A1(n153), .A2(n149), .Y(n109) );
  AND2X1_HVT U392 ( .A1(a_addr[3]), .A2(a_addr[2]), .Y(n149) );
  AO21X1_HVT U393 ( .A1(n148), .A2(n110), .A3(rst), .Y(N307) );
  AND2X1_HVT U394 ( .A1(n154), .A2(n150), .Y(n110) );
  AO21X1_HVT U395 ( .A1(n148), .A2(n111), .A3(rst), .Y(N306) );
  AND2X1_HVT U396 ( .A1(n154), .A2(n151), .Y(n111) );
  AO21X1_HVT U397 ( .A1(n148), .A2(n112), .A3(rst), .Y(N305) );
  AND2X1_HVT U398 ( .A1(n154), .A2(n152), .Y(n112) );
  AO21X1_HVT U399 ( .A1(n148), .A2(n113), .A3(rst), .Y(N304) );
  AND2X1_HVT U400 ( .A1(n154), .A2(n153), .Y(n113) );
  AND2X1_HVT U401 ( .A1(a_addr[3]), .A2(n155), .Y(n154) );
  AO21X1_HVT U402 ( .A1(n148), .A2(n114), .A3(rst), .Y(N303) );
  AND2X1_HVT U403 ( .A1(n156), .A2(n150), .Y(n114) );
  AO21X1_HVT U404 ( .A1(n148), .A2(n115), .A3(rst), .Y(N302) );
  AND2X1_HVT U405 ( .A1(n156), .A2(n151), .Y(n115) );
  AO21X1_HVT U406 ( .A1(n148), .A2(n116), .A3(rst), .Y(N301) );
  AND2X1_HVT U407 ( .A1(n156), .A2(n152), .Y(n116) );
  AO21X1_HVT U408 ( .A1(n148), .A2(n117), .A3(rst), .Y(N300) );
  AND2X1_HVT U409 ( .A1(n156), .A2(n153), .Y(n117) );
  AND2X1_HVT U410 ( .A1(a_addr[2]), .A2(n157), .Y(n156) );
  AO21X1_HVT U411 ( .A1(n148), .A2(n118), .A3(rst), .Y(N299) );
  AND2X1_HVT U412 ( .A1(n158), .A2(n150), .Y(n118) );
  AND2X1_HVT U413 ( .A1(a_addr[1]), .A2(a_addr[0]), .Y(n150) );
  AO21X1_HVT U414 ( .A1(n148), .A2(n119), .A3(rst), .Y(N298) );
  AND2X1_HVT U415 ( .A1(n158), .A2(n151), .Y(n119) );
  AND2X1_HVT U416 ( .A1(a_addr[1]), .A2(n159), .Y(n151) );
  AO21X1_HVT U417 ( .A1(n148), .A2(n120), .A3(rst), .Y(N297) );
  AND2X1_HVT U418 ( .A1(n158), .A2(n152), .Y(n120) );
  AND2X1_HVT U419 ( .A1(a_addr[0]), .A2(n160), .Y(n152) );
  AO21X1_HVT U420 ( .A1(n148), .A2(n121), .A3(rst), .Y(N296) );
  AND2X1_HVT U421 ( .A1(n158), .A2(n153), .Y(n121) );
  AND2X1_HVT U422 ( .A1(n159), .A2(n160), .Y(n153) );
  INVX0_HVT U423 ( .A(a_addr[1]), .Y(n160) );
  INVX0_HVT U424 ( .A(a_addr[0]), .Y(n159) );
  AND2X1_HVT U425 ( .A1(n155), .A2(n157), .Y(n158) );
  INVX0_HVT U426 ( .A(a_addr[3]), .Y(n157) );
  INVX0_HVT U427 ( .A(a_addr[2]), .Y(n155) );
  AND2X1_HVT U428 ( .A1(n139), .A2(n133), .Y(n148) );
  AND2X1_HVT U429 ( .A1(n142), .A2(n145), .Y(n133) );
  INVX0_HVT U430 ( .A(a_din[2]), .Y(n145) );
  INVX0_HVT U431 ( .A(a_din[1]), .Y(n142) );
  AND3X1_HVT U432 ( .A1(n135), .A2(n147), .A3(N495), .Y(n139) );
  AND2X1_HVT U433 ( .A1(write), .A2(n161), .Y(N495) );
  INVX0_HVT U434 ( .A(rst), .Y(n161) );
  INVX0_HVT U435 ( .A(a_din[3]), .Y(n147) );
  INVX0_HVT U436 ( .A(a_din[0]), .Y(n135) );
endmodule

