
module sbox_14 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n10, n19, n23, n32, n50, n118, n119, n132, n140, n160, n210, n211,
         n212, n213, n216, n217, n218, n219, n221, n231, n232, n236, n238,
         n242, n243, n245, n255, n261, n264, n268, n271, n273, n274, n277,
         n282, n283, n285, n289, n290, n293, n296, n297, n300, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796;

  NAND2X0_HVT U4 ( .A1(n340), .A2(n794), .Y(n793) );
  NAND2X0_HVT U5 ( .A1(n330), .A2(n523), .Y(n791) );
  NAND2X0_HVT U13 ( .A1(n784), .A2(n245), .Y(n785) );
  NAND2X0_HVT U15 ( .A1(n794), .A2(n474), .Y(n782) );
  NAND2X0_HVT U21 ( .A1(n340), .A2(n343), .Y(n777) );
  NAND2X0_HVT U24 ( .A1(n433), .A2(n419), .Y(n775) );
  NAND2X0_HVT U33 ( .A1(n560), .A2(n343), .Y(n767) );
  NAND2X0_HVT U35 ( .A1(n273), .A2(n411), .Y(n765) );
  NAND2X0_HVT U42 ( .A1(n361), .A2(n433), .Y(n758) );
  NAND2X0_HVT U53 ( .A1(n747), .A2(n757), .Y(n748) );
  NAND2X0_HVT U56 ( .A1(n316), .A2(n743), .Y(n744) );
  MUX41X1_HVT U57 ( .A1(n119), .A3(n779), .A2(n744), .A4(n787), .S0(n483), 
        .S1(n532), .Y(n742) );
  NAND2X0_HVT U62 ( .A1(n419), .A2(n525), .Y(n737) );
  AO21X1_HVT U66 ( .A1(n432), .A2(n532), .A3(n581), .Y(n733) );
  MUX41X1_HVT U68 ( .A1(n548), .A3(n733), .A2(n732), .A4(n734), .S0(n392), 
        .S1(n535), .Y(n731) );
  NAND2X0_HVT U73 ( .A1(n465), .A2(n726), .Y(n727) );
  MUX41X1_HVT U77 ( .A1(n788), .A3(n561), .A2(n723), .A4(n553), .S0(n479), 
        .S1(n216), .Y(n722) );
  AND2X1_HVT U83 ( .A1(n314), .A2(n437), .Y(n715) );
  NAND2X0_HVT U85 ( .A1(n19), .A2(n486), .Y(n713) );
  NAND2X0_HVT U101 ( .A1(n696), .A2(n695), .Y(n697) );
  MUX41X1_HVT U103 ( .A1(n794), .A3(n566), .A2(n556), .A4(n765), .S0(n283), 
        .S1(n398), .Y(n693) );
  MUX41X1_HVT U105 ( .A1(n573), .A3(n752), .A2(n692), .A4(n563), .S0(n515), 
        .S1(n398), .Y(n691) );
  NAND2X0_HVT U110 ( .A1(n308), .A2(n686), .Y(n687) );
  AND2X1_HVT U115 ( .A1(n218), .A2(n319), .Y(n683) );
  NAND2X0_HVT U123 ( .A1(n673), .A2(n674), .Y(n675) );
  MUX41X1_HVT U125 ( .A1(n777), .A3(n512), .A2(n548), .A4(n559), .S0(n515), 
        .S1(n446), .Y(n672) );
  MUX41X1_HVT U135 ( .A1(n552), .A3(n462), .A2(n791), .A4(n772), .S0(n515), 
        .S1(n535), .Y(n664) );
  AND2X1_HVT U140 ( .A1(n372), .A2(n436), .Y(n659) );
  NAND2X0_HVT U158 ( .A1(n314), .A2(n486), .Y(n643) );
  MUX41X1_HVT U159 ( .A1(n785), .A3(n474), .A2(n643), .A4(n582), .S0(n283), 
        .S1(n398), .Y(n642) );
  AND2X1_HVT U162 ( .A1(n359), .A2(n726), .Y(n639) );
  MUX41X1_HVT U163 ( .A1(n574), .A3(n639), .A2(n507), .A4(n640), .S0(n392), 
        .S1(n536), .Y(n638) );
  MUX41X1_HVT U165 ( .A1(n777), .A3(n572), .A2(n754), .A4(n637), .S0(n446), 
        .S1(n140), .Y(n636) );
  NAND2X0_HVT U166 ( .A1(n245), .A2(n743), .Y(n635) );
  NAND2X0_HVT U167 ( .A1(n491), .A2(n411), .Y(n634) );
  MUX41X1_HVT U168 ( .A1(n119), .A3(n372), .A2(n634), .A4(n635), .S0(n516), 
        .S1(n535), .Y(n633) );
  NAND2X0_HVT U174 ( .A1(n456), .A2(n469), .Y(n784) );
  NAND2X0_HVT U177 ( .A1(n327), .A2(n421), .Y(n626) );
  MUX41X1_HVT U180 ( .A1(n547), .A3(n243), .A2(n785), .A4(n504), .S0(n353), 
        .S1(n381), .Y(n623) );
  MUX41X1_HVT U189 ( .A1(n615), .A3(n213), .A2(n616), .A4(n563), .S0(n353), 
        .S1(n517), .Y(n614) );
  MUX41X1_HVT U195 ( .A1(n359), .A3(n407), .A2(n245), .A4(n763), .S0(n283), 
        .S1(n478), .Y(n609) );
  MUX41X1_HVT U203 ( .A1(n764), .A3(n540), .A2(n786), .A4(n768), .S0(n517), 
        .S1(n446), .Y(n601) );
  NAND2X0_HVT U208 ( .A1(n217), .A2(n361), .Y(n686) );
  NAND2X0_HVT U214 ( .A1(n359), .A2(n19), .Y(n597) );
  NAND2X0_HVT U215 ( .A1(n686), .A2(n465), .Y(n596) );
  NAND2X0_HVT U218 ( .A1(n460), .A2(n218), .Y(n649) );
  NAND2X0_HVT U220 ( .A1(n364), .A2(n597), .Y(n718) );
  INVX0_HVT U241 ( .A(n775), .Y(n585) );
  INVX0_HVT U242 ( .A(n758), .Y(n584) );
  INVX0_HVT U245 ( .A(n791), .Y(n582) );
  INVX0_HVT U256 ( .A(n649), .Y(n575) );
  INVX0_HVT U268 ( .A(n777), .Y(n564) );
  INVX0_HVT U270 ( .A(n596), .Y(n563) );
  INVX0_HVT U278 ( .A(n767), .Y(n557) );
  INVX0_HVT U280 ( .A(n770), .Y(n556) );
  INVX0_HVT U283 ( .A(n387), .Y(n555) );
  INVX0_HVT U284 ( .A(n597), .Y(n554) );
  INVX0_HVT U289 ( .A(n695), .Y(n550) );
  INVX0_HVT U294 ( .A(n789), .Y(n548) );
  INVX0_HVT U295 ( .A(n793), .Y(n547) );
  INVX0_HVT U306 ( .A(n634), .Y(n541) );
  INVX1_HVT U1 ( .A(n537), .Y(n497) );
  INVX1_HVT U2 ( .A(n306), .Y(n364) );
  INVX1_HVT U3 ( .A(n336), .Y(n337) );
  OA21X1_HVT U6 ( .A1(n416), .A2(n766), .A3(n282), .Y(n619) );
  NBUFFX2_HVT U7 ( .A(n456), .Y(n264) );
  INVX1_HVT U8 ( .A(n726), .Y(n581) );
  AO21X1_HVT U9 ( .A1(n436), .A2(n460), .A3(n320), .Y(n696) );
  XNOR2X1_HVT U10 ( .A1(n264), .A2(n530), .Y(n514) );
  AO21X1_HVT U11 ( .A1(n140), .A2(n372), .A3(n470), .Y(n680) );
  INVX1_HVT U12 ( .A(n485), .Y(n409) );
  MUX21X1_HVT U14 ( .A1(n793), .A2(n662), .S0(n368), .Y(n661) );
  INVX1_HVT U16 ( .A(n459), .Y(n462) );
  XOR2X1_HVT U17 ( .A1(n217), .A2(n242), .Y(n507) );
  INVX1_HVT U18 ( .A(n759), .Y(n544) );
  INVX1_HVT U19 ( .A(n773), .Y(n567) );
  INVX1_HVT U20 ( .A(n586), .Y(n569) );
  INVX1_HVT U22 ( .A(n496), .Y(n446) );
  MUX21X1_HVT U23 ( .A1(n748), .A2(n749), .S0(n536), .Y(n746) );
  AND3X1_HVT U25 ( .A1(n308), .A2(n743), .A3(n718), .Y(n719) );
  MUX21X1_HVT U26 ( .A1(n316), .A2(n464), .S0(n393), .Y(n710) );
  MUX21X1_HVT U27 ( .A1(n560), .A2(n319), .S0(n318), .Y(n703) );
  INVX1_HVT U28 ( .A(n313), .Y(n774) );
  INVX1_HVT U29 ( .A(n686), .Y(n562) );
  INVX1_HVT U30 ( .A(n318), .Y(n314) );
  INVX1_HVT U31 ( .A(n594), .Y(n407) );
  INVX1_HVT U32 ( .A(n376), .Y(n343) );
  INVX1_HVT U34 ( .A(n436), .Y(n456) );
  NBUFFX2_HVT U36 ( .A(n529), .Y(n436) );
  INVX1_HVT U37 ( .A(n529), .Y(n457) );
  INVX0_HVT U38 ( .A(n515), .Y(n440) );
  INVX1_HVT U39 ( .A(n489), .Y(n140) );
  INVX1_HVT U40 ( .A(n530), .Y(n50) );
  INVX1_HVT U41 ( .A(n381), .Y(n368) );
  AND2X1_HVT U43 ( .A1(n354), .A2(n355), .Y(n10) );
  INVX0_HVT U44 ( .A(n551), .Y(n472) );
  INVX1_HVT U45 ( .A(n306), .Y(n535) );
  INVX1_HVT U46 ( .A(n519), .Y(n477) );
  INVX0_HVT U47 ( .A(n583), .Y(n433) );
  INVX1_HVT U48 ( .A(n315), .Y(n316) );
  NAND2X0_HVT U49 ( .A1(n342), .A2(n19), .Y(n23) );
  NAND2X0_HVT U50 ( .A1(n580), .A2(n393), .Y(n32) );
  NAND2X0_HVT U51 ( .A1(n23), .A2(n32), .Y(n764) );
  INVX0_HVT U52 ( .A(n393), .Y(n19) );
  INVX1_HVT U54 ( .A(n764), .Y(n571) );
  MUX21X1_HVT U55 ( .A1(n783), .A2(n485), .S0(n50), .Y(n699) );
  MUX21X1_HVT U58 ( .A1(n315), .A2(n468), .S0(n456), .Y(n391) );
  INVX1_HVT U59 ( .A(n788), .Y(n566) );
  INVX0_HVT U60 ( .A(in[3]), .Y(n336) );
  INVX1_HVT U61 ( .A(n391), .Y(n763) );
  MUX21X2_HVT U63 ( .A1(n573), .A2(n769), .S0(n283), .Y(n670) );
  INVX1_HVT U64 ( .A(n792), .Y(n560) );
  INVX1_HVT U65 ( .A(n427), .Y(n217) );
  MUX21X1_HVT U67 ( .A1(n345), .A2(n507), .S0(n50), .Y(n668) );
  INVX1_HVT U69 ( .A(n455), .Y(n768) );
  MUX21X1_HVT U70 ( .A1(n273), .A2(n526), .S0(n329), .Y(n595) );
  INVX1_HVT U71 ( .A(n471), .Y(n118) );
  INVX1_HVT U72 ( .A(n551), .Y(n471) );
  INVX1_HVT U74 ( .A(n531), .Y(n530) );
  MUX21X2_HVT U75 ( .A1(n792), .A2(n461), .S0(n318), .Y(n312) );
  INVX1_HVT U76 ( .A(n454), .Y(n315) );
  INVX1_HVT U78 ( .A(n337), .Y(n583) );
  INVX1_HVT U79 ( .A(n427), .Y(n454) );
  MUX21X2_HVT U80 ( .A1(n503), .A2(n523), .S0(n411), .Y(n769) );
  INVX1_HVT U81 ( .A(n528), .Y(n318) );
  INVX0_HVT U82 ( .A(n577), .Y(n461) );
  MUX41X1_HVT U84 ( .A1(n666), .A3(n671), .A2(n678), .A4(n684), .S0(n520), 
        .S1(in[6]), .Y(out[3]) );
  INVX0_HVT U86 ( .A(n743), .Y(n578) );
  INVX1_HVT U87 ( .A(n522), .Y(n503) );
  NBUFFX2_HVT U88 ( .A(n390), .Y(n526) );
  INVX1_HVT U89 ( .A(n517), .Y(n369) );
  NAND2X0_HVT U90 ( .A1(n706), .A2(n400), .Y(n481) );
  MUX21X1_HVT U91 ( .A1(n311), .A2(n493), .S0(n492), .Y(n490) );
  OA21X1_HVT U92 ( .A1(n510), .A2(n320), .A3(n415), .Y(n631) );
  MUX21X1_HVT U93 ( .A1(n463), .A2(n513), .S0(n338), .Y(n637) );
  INVX1_HVT U94 ( .A(n410), .Y(n338) );
  AO21X1_HVT U95 ( .A1(n508), .A2(n364), .A3(n575), .Y(n607) );
  INVX1_HVT U96 ( .A(n211), .Y(n753) );
  AND3X1_HVT U97 ( .A1(n381), .A2(n19), .A3(n437), .Y(n669) );
  OA21X1_HVT U98 ( .A1(n541), .A2(n416), .A3(n409), .Y(n655) );
  MUX21X1_HVT U99 ( .A1(n651), .A2(n650), .S0(n400), .Y(n648) );
  INVX1_HVT U100 ( .A(n341), .Y(n761) );
  INVX1_HVT U102 ( .A(n488), .Y(n353) );
  INVX0_HVT U104 ( .A(n306), .Y(n478) );
  INVX0_HVT U106 ( .A(n497), .Y(n398) );
  INVX1_HVT U107 ( .A(n518), .Y(n367) );
  INVX1_HVT U108 ( .A(n519), .Y(n488) );
  INVX0_HVT U109 ( .A(n533), .Y(n467) );
  INVX1_HVT U111 ( .A(n496), .Y(n537) );
  INVX0_HVT U112 ( .A(n497), .Y(n479) );
  INVX0_HVT U113 ( .A(n529), .Y(n443) );
  INVX1_HVT U114 ( .A(n533), .Y(n424) );
  INVX0_HVT U116 ( .A(n411), .Y(n218) );
  INVX1_HVT U117 ( .A(in[1]), .Y(n529) );
  NBUFFX2_HVT U118 ( .A(n537), .Y(n519) );
  NBUFFX2_HVT U119 ( .A(n503), .Y(n342) );
  AND2X1_HVT U120 ( .A1(n303), .A2(n304), .Y(n119) );
  AND2X1_HVT U121 ( .A1(n385), .A2(n386), .Y(n132) );
  INVX0_HVT U122 ( .A(n242), .Y(n361) );
  INVX0_HVT U124 ( .A(n277), .Y(n282) );
  INVX0_HVT U126 ( .A(n549), .Y(n277) );
  INVX1_HVT U127 ( .A(n373), .Y(n325) );
  MUX41X1_HVT U128 ( .A1(n617), .A3(n614), .A2(n621), .A4(n618), .S0(n367), 
        .S1(n520), .Y(n613) );
  MUX21X2_HVT U129 ( .A1(n274), .A2(n217), .S0(n318), .Y(n788) );
  MUX41X1_HVT U130 ( .A1(n554), .A3(n570), .A2(n771), .A4(n569), .S0(n516), 
        .S1(n488), .Y(n624) );
  MUX41X1_HVT U131 ( .A1(n668), .A3(n670), .A2(n667), .A4(n669), .S0(n518), 
        .S1(n477), .Y(n666) );
  NBUFFX2_HVT U132 ( .A(n337), .Y(n521) );
  INVX1_HVT U133 ( .A(n771), .Y(n573) );
  NAND2X0_HVT U134 ( .A1(n794), .A2(n140), .Y(n160) );
  NAND2X0_HVT U136 ( .A1(n571), .A2(n489), .Y(n210) );
  NAND2X0_HVT U137 ( .A1(n160), .A2(n210), .Y(n689) );
  XNOR2X1_HVT U138 ( .A1(n531), .A2(n306), .Y(n211) );
  MUX41X1_HVT U139 ( .A1(n691), .A3(n693), .A2(n694), .A4(n698), .S0(n458), 
        .S1(n520), .Y(n690) );
  INVX1_HVT U141 ( .A(n531), .Y(n305) );
  NBUFFX2_HVT U142 ( .A(n443), .Y(n212) );
  INVX1_HVT U143 ( .A(n468), .Y(n470) );
  NOR2X0_HVT U144 ( .A1(n337), .A2(n395), .Y(n427) );
  INVX1_HVT U145 ( .A(n705), .Y(n561) );
  MUX41X1_HVT U146 ( .A1(n716), .A3(n717), .A2(n712), .A4(n714), .S0(n458), 
        .S1(n331), .Y(n711) );
  INVX1_HVT U147 ( .A(in[0]), .Y(n331) );
  INVX1_HVT U148 ( .A(n373), .Y(n480) );
  MUX21X1_HVT U149 ( .A1(n631), .A2(n632), .S0(n400), .Y(n630) );
  NBUFFX2_HVT U150 ( .A(n784), .Y(n213) );
  NBUFFX2_HVT U151 ( .A(n530), .Y(n216) );
  INVX0_HVT U152 ( .A(n427), .Y(n792) );
  XNOR2X1_HVT U153 ( .A1(n525), .A2(n343), .Y(n751) );
  INVX1_HVT U154 ( .A(n357), .Y(n358) );
  INVX1_HVT U155 ( .A(n357), .Y(n245) );
  XNOR2X2_HVT U156 ( .A1(n330), .A2(n459), .Y(n755) );
  NAND2X0_HVT U157 ( .A1(n221), .A2(n218), .Y(n219) );
  NAND2X0_HVT U160 ( .A1(n219), .A2(n767), .Y(n590) );
  INVX1_HVT U161 ( .A(n528), .Y(n411) );
  INVX0_HVT U164 ( .A(n497), .Y(n483) );
  NBUFFX2_HVT U169 ( .A(n522), .Y(n221) );
  NBUFFX2_HVT U170 ( .A(n373), .Y(n522) );
  INVX0_HVT U171 ( .A(n472), .Y(n474) );
  INVX0_HVT U172 ( .A(n528), .Y(n348) );
  INVX0_HVT U173 ( .A(n528), .Y(n419) );
  AO21X1_HVT U175 ( .A1(n705), .A2(n446), .A3(n575), .Y(n706) );
  INVX0_HVT U176 ( .A(n432), .Y(n787) );
  MUX21X2_HVT U178 ( .A1(n486), .A2(n407), .S0(n519), .Y(n730) );
  MUX41X1_HVT U179 ( .A1(n689), .A3(n688), .A2(n132), .A4(n685), .S0(n483), 
        .S1(n467), .Y(n684) );
  MUX41X1_HVT U181 ( .A1(n773), .A3(n728), .A2(n775), .A4(n727), .S0(n356), 
        .S1(n479), .Y(n725) );
  MUX21X1_HVT U182 ( .A1(n697), .A2(n538), .S0(n516), .Y(n694) );
  NAND2X0_HVT U183 ( .A1(n462), .A2(n532), .Y(n231) );
  NAND2X0_HVT U184 ( .A1(n566), .A2(n367), .Y(n232) );
  NAND2X0_HVT U185 ( .A1(n231), .A2(n232), .Y(n732) );
  INVX1_HVT U186 ( .A(n516), .Y(n489) );
  NAND2X0_HVT U187 ( .A1(n795), .A2(n212), .Y(n236) );
  NAND2X0_HVT U188 ( .A1(n342), .A2(n419), .Y(n238) );
  NAND2X0_HVT U190 ( .A1(n236), .A2(n238), .Y(n778) );
  MUX21X1_HVT U191 ( .A1(n778), .A2(n372), .S0(n519), .Y(n720) );
  INVX1_HVT U192 ( .A(n457), .Y(n242) );
  INVX0_HVT U193 ( .A(n337), .Y(n332) );
  MUX21X1_HVT U194 ( .A1(n561), .A2(n762), .S0(n488), .Y(n645) );
  MUX21X1_HVT U196 ( .A1(n580), .A2(n319), .S0(n264), .Y(n640) );
  INVX0_HVT U197 ( .A(n468), .Y(n359) );
  INVX0_HVT U198 ( .A(n566), .Y(n243) );
  INVX1_HVT U199 ( .A(n332), .Y(n326) );
  MUX41X1_HVT U200 ( .A1(n509), .A3(n578), .A2(n782), .A4(n218), .S0(n356), 
        .S1(n536), .Y(n701) );
  MUX21X1_HVT U201 ( .A1(n217), .A2(n524), .S0(n348), .Y(n341) );
  MUX41X1_HVT U202 ( .A1(n544), .A3(n567), .A2(n341), .A4(n316), .S0(n353), 
        .S1(n50), .Y(n621) );
  INVX0_HVT U204 ( .A(n348), .Y(n327) );
  MUX41X1_HVT U205 ( .A1(n709), .A3(n702), .A2(n704), .A4(n701), .S0(n331), 
        .S1(n424), .Y(n700) );
  MUX41X1_HVT U206 ( .A1(n506), .A3(n345), .A2(n574), .A4(n474), .S0(n533), 
        .S1(n478), .Y(n738) );
  INVX1_HVT U207 ( .A(n463), .Y(n372) );
  NAND2X0_HVT U209 ( .A1(n679), .A2(n424), .Y(n255) );
  NAND2X0_HVT U210 ( .A1(n682), .A2(n458), .Y(n261) );
  NAND2X0_HVT U211 ( .A1(n255), .A2(n261), .Y(n678) );
  INVX1_HVT U212 ( .A(n436), .Y(n393) );
  INVX0_HVT U213 ( .A(n529), .Y(n528) );
  MUX41X1_HVT U216 ( .A1(n576), .A3(n578), .A2(n313), .A4(n311), .S0(n356), 
        .S1(n479), .Y(n724) );
  INVX1_HVT U217 ( .A(in[7]), .Y(n496) );
  MUX41X1_HVT U219 ( .A1(n758), .A3(n710), .A2(n754), .A4(n543), .S0(n483), 
        .S1(n440), .Y(n709) );
  NAND2X0_HVT U221 ( .A1(n524), .A2(n329), .Y(n268) );
  NAND2X0_HVT U222 ( .A1(n469), .A2(n393), .Y(n271) );
  NAND2X0_HVT U223 ( .A1(n271), .A2(n268), .Y(n592) );
  INVX0_HVT U224 ( .A(n592), .Y(n553) );
  INVX0_HVT U225 ( .A(n461), .Y(n463) );
  INVX0_HVT U226 ( .A(n480), .Y(n394) );
  INVX1_HVT U227 ( .A(n307), .Y(n468) );
  INVX1_HVT U228 ( .A(n325), .Y(n273) );
  NBUFFX2_HVT U229 ( .A(n521), .Y(n274) );
  INVX1_HVT U230 ( .A(n795), .Y(n491) );
  NAND2X0_HVT U231 ( .A1(n687), .A2(n283), .Y(n285) );
  NAND2X0_HVT U232 ( .A1(n415), .A2(n489), .Y(n289) );
  NAND2X0_HVT U233 ( .A1(n285), .A2(n289), .Y(n685) );
  INVX0_HVT U234 ( .A(n531), .Y(n283) );
  MUX41X1_HVT U235 ( .A1(n585), .A3(n783), .A2(n755), .A4(n545), .S0(n283), 
        .S1(n497), .Y(n716) );
  NAND2X0_HVT U236 ( .A1(n433), .A2(n361), .Y(n290) );
  NAND2X0_HVT U237 ( .A1(n473), .A2(n348), .Y(n293) );
  NAND2X0_HVT U238 ( .A1(n290), .A2(n293), .Y(n776) );
  INVX0_HVT U239 ( .A(n471), .Y(n473) );
  INVX0_HVT U240 ( .A(n776), .Y(n549) );
  INVX1_HVT U243 ( .A(n329), .Y(n330) );
  INVX0_HVT U244 ( .A(n782), .Y(n546) );
  NAND2X0_HVT U246 ( .A1(n524), .A2(n212), .Y(n296) );
  NAND2X0_HVT U247 ( .A1(n340), .A2(n419), .Y(n297) );
  NAND2X0_HVT U248 ( .A1(n296), .A2(n297), .Y(n786) );
  INVX0_HVT U249 ( .A(n786), .Y(n565) );
  OR2X1_HVT U250 ( .A1(n580), .A2(n484), .Y(n741) );
  INVX1_HVT U251 ( .A(n484), .Y(n794) );
  MUX21X1_HVT U252 ( .A1(n523), .A2(n513), .S0(n212), .Y(n760) );
  NAND2X0_HVT U253 ( .A1(n326), .A2(n480), .Y(n300) );
  NAND2X0_HVT U254 ( .A1(n437), .A2(n343), .Y(n303) );
  NAND2X0_HVT U255 ( .A1(n470), .A2(n327), .Y(n304) );
  MUX41X1_HVT U257 ( .A1(n317), .A3(n542), .A2(n754), .A4(n578), .S0(n400), 
        .S1(n446), .Y(n653) );
  INVX1_HVT U258 ( .A(n328), .Y(n728) );
  MUX41X1_HVT U259 ( .A1(n648), .A3(n644), .A2(n647), .A4(n642), .S0(n331), 
        .S1(n467), .Y(n641) );
  MUX21X1_HVT U260 ( .A1(n553), .A2(n462), .S0(n364), .Y(n651) );
  MUX41X1_HVT U261 ( .A1(n633), .A3(n630), .A2(n638), .A4(n636), .S0(n424), 
        .S1(n520), .Y(n629) );
  INVX1_HVT U262 ( .A(n515), .Y(n400) );
  INVX1_HVT U263 ( .A(n515), .Y(n356) );
  INVX1_HVT U264 ( .A(n537), .Y(n306) );
  NAND2X0_HVT U265 ( .A1(n334), .A2(n333), .Y(n307) );
  NBUFFX2_HVT U266 ( .A(n305), .Y(n516) );
  INVX1_HVT U267 ( .A(n242), .Y(n321) );
  MUX21X1_HVT U269 ( .A1(n780), .A2(n455), .S0(n216), .Y(n667) );
  NBUFFX2_HVT U271 ( .A(n526), .Y(n308) );
  NAND2X0_HVT U272 ( .A1(n358), .A2(n218), .Y(n309) );
  NAND2X0_HVT U273 ( .A1(n526), .A2(n348), .Y(n310) );
  NAND2X0_HVT U274 ( .A1(n309), .A2(n310), .Y(n449) );
  INVX0_HVT U275 ( .A(n449), .Y(n772) );
  MUX41X1_HVT U276 ( .A1(n552), .A3(n372), .A2(n759), .A4(n772), .S0(n353), 
        .S1(n368), .Y(n610) );
  INVX1_HVT U277 ( .A(n50), .Y(n381) );
  NBUFFX2_HVT U279 ( .A(n491), .Y(n311) );
  INVX0_HVT U281 ( .A(n390), .Y(n513) );
  MUX21X1_HVT U282 ( .A1(n340), .A2(n526), .S0(n318), .Y(n588) );
  INVX1_HVT U285 ( .A(n471), .Y(n319) );
  AND2X1_HVT U286 ( .A1(n408), .A2(n379), .Y(n313) );
  NBUFFX2_HVT U287 ( .A(n583), .Y(n523) );
  INVX0_HVT U288 ( .A(n581), .Y(n317) );
  NAND2X0_HVT U290 ( .A1(n457), .A2(n334), .Y(n726) );
  MUX21X2_HVT U291 ( .A1(n473), .A2(n324), .S0(n348), .Y(n759) );
  MUX21X1_HVT U292 ( .A1(n580), .A2(n560), .S0(n314), .Y(n762) );
  MUX21X1_HVT U293 ( .A1(n273), .A2(n454), .S0(n410), .Y(n455) );
  NBUFFX2_HVT U296 ( .A(n497), .Y(n320) );
  INVX0_HVT U297 ( .A(n778), .Y(n545) );
  NAND2X0_HVT U298 ( .A1(n245), .A2(n321), .Y(n322) );
  NAND2X0_HVT U299 ( .A1(n433), .A2(n419), .Y(n323) );
  NAND2X0_HVT U300 ( .A1(n322), .A2(n323), .Y(n432) );
  INVX0_HVT U301 ( .A(n513), .Y(n324) );
  INVX1_HVT U302 ( .A(n527), .Y(n486) );
  INVX1_HVT U303 ( .A(n527), .Y(n580) );
  XOR2X2_HVT U304 ( .A1(n221), .A2(n456), .Y(n773) );
  MUX41X1_HVT U305 ( .A1(n724), .A3(n729), .A2(n722), .A4(n725), .S0(n520), 
        .S1(n424), .Y(n721) );
  INVX1_HVT U307 ( .A(in[2]), .Y(n531) );
  INVX1_HVT U308 ( .A(n511), .Y(n492) );
  MUX21X1_HVT U309 ( .A1(n503), .A2(n360), .S0(n329), .Y(n328) );
  INVX0_HVT U310 ( .A(n360), .Y(n464) );
  INVX1_HVT U311 ( .A(n443), .Y(n329) );
  MUX41X1_HVT U312 ( .A1(n508), .A3(n505), .A2(n576), .A4(n713), .S0(n515), 
        .S1(n320), .Y(n712) );
  INVX1_HVT U313 ( .A(n514), .Y(n384) );
  MUX21X1_HVT U314 ( .A1(n358), .A2(n525), .S0(n314), .Y(n616) );
  INVX0_HVT U315 ( .A(in[4]), .Y(n373) );
  MUX41X1_HVT U316 ( .A1(n611), .A3(n609), .A2(n610), .A4(n606), .S0(n331), 
        .S1(n424), .Y(n605) );
  NAND2X0_HVT U317 ( .A1(n373), .A2(n332), .Y(n333) );
  NAND2X0_HVT U318 ( .A1(n326), .A2(n395), .Y(n334) );
  NAND2X0_HVT U319 ( .A1(n300), .A2(n333), .Y(n790) );
  INVX0_HVT U320 ( .A(n790), .Y(n551) );
  AND2X1_HVT U321 ( .A1(n350), .A2(n349), .Y(n335) );
  INVX1_HVT U322 ( .A(n364), .Y(n416) );
  INVX1_HVT U323 ( .A(n769), .Y(n572) );
  INVX1_HVT U324 ( .A(n528), .Y(n410) );
  INVX1_HVT U325 ( .A(n498), .Y(n339) );
  INVX1_HVT U326 ( .A(in[6]), .Y(n498) );
  INVX0_HVT U327 ( .A(n315), .Y(n340) );
  INVX1_HVT U328 ( .A(n410), .Y(n376) );
  OA21X1_HVT U329 ( .A1(n368), .A2(n391), .A3(n312), .Y(n688) );
  MUX41X1_HVT U330 ( .A1(n282), .A3(n474), .A2(n562), .A4(n465), .S0(n515), 
        .S1(n478), .Y(n657) );
  INVX0_HVT U331 ( .A(n360), .Y(n465) );
  NBUFFX2_HVT U332 ( .A(n305), .Y(n515) );
  MUX41X1_HVT U333 ( .A1(n654), .A3(n653), .A2(n658), .A4(n657), .S0(n424), 
        .S1(n520), .Y(n652) );
  MUX21X1_HVT U334 ( .A1(n433), .A2(n765), .S0(n532), .Y(n749) );
  NAND2X0_HVT U335 ( .A1(n487), .A2(n338), .Y(n344) );
  NAND2X0_HVT U336 ( .A1(n238), .A2(n344), .Y(n780) );
  INVX1_HVT U337 ( .A(n765), .Y(n568) );
  AND2X1_HVT U338 ( .A1(n362), .A2(n363), .Y(n345) );
  NAND2X0_HVT U339 ( .A1(n584), .A2(n488), .Y(n346) );
  NAND2X0_HVT U340 ( .A1(n446), .A2(n570), .Y(n347) );
  NAND2X0_HVT U341 ( .A1(n346), .A2(n347), .Y(n608) );
  INVX1_HVT U342 ( .A(n468), .Y(n469) );
  MUX21X1_HVT U343 ( .A1(n504), .A2(n781), .S0(n477), .Y(n604) );
  NAND2X0_HVT U344 ( .A1(n525), .A2(n348), .Y(n349) );
  NAND2X0_HVT U345 ( .A1(n464), .A2(n361), .Y(n350) );
  NAND2X0_HVT U346 ( .A1(n349), .A2(n350), .Y(n783) );
  NAND2X0_HVT U347 ( .A1(n538), .A2(n369), .Y(n351) );
  NAND2X0_HVT U348 ( .A1(n10), .A2(n516), .Y(n352) );
  NAND2X0_HVT U349 ( .A1(n351), .A2(n352), .Y(n665) );
  NAND2X0_HVT U350 ( .A1(n462), .A2(n353), .Y(n354) );
  NAND2X0_HVT U351 ( .A1(n590), .A2(n477), .Y(n355) );
  MUX41X1_HVT U352 ( .A1(n509), .A3(n585), .A2(n703), .A4(n407), .S0(n356), 
        .S1(n536), .Y(n702) );
  MUX21X1_HVT U353 ( .A1(n491), .A2(n560), .S0(n419), .Y(n628) );
  INVX0_HVT U354 ( .A(n796), .Y(n357) );
  MUX21X1_HVT U355 ( .A1(n464), .A2(n319), .S0(n376), .Y(n692) );
  AND2X1_HVT U356 ( .A1(n583), .A2(n325), .Y(n360) );
  MUX41X1_HVT U357 ( .A1(n762), .A3(n570), .A2(n626), .A4(n780), .S0(n356), 
        .S1(n416), .Y(n625) );
  NAND2X0_HVT U358 ( .A1(n524), .A2(n212), .Y(n362) );
  NAND2X0_HVT U359 ( .A1(n118), .A2(n419), .Y(n363) );
  NAND2X0_HVT U360 ( .A1(n362), .A2(n363), .Y(n781) );
  INVX0_HVT U361 ( .A(n437), .Y(n421) );
  INVX0_HVT U362 ( .A(n762), .Y(n558) );
  INVX0_HVT U363 ( .A(n366), .Y(n577) );
  INVX0_HVT U364 ( .A(n366), .Y(n487) );
  MUX41X1_HVT U365 ( .A1(n421), .A3(n628), .A2(n550), .A4(n213), .S0(n364), 
        .S1(n530), .Y(n627) );
  NAND2X0_HVT U366 ( .A1(n463), .A2(n264), .Y(n365) );
  NAND2X0_HVT U367 ( .A1(n325), .A2(n583), .Y(n366) );
  MUX41X1_HVT U368 ( .A1(n785), .A3(n744), .A2(n277), .A4(n579), .S0(n369), 
        .S1(n535), .Y(n600) );
  INVX0_HVT U369 ( .A(n766), .Y(n579) );
  INVX0_HVT U370 ( .A(n780), .Y(n574) );
  MUX41X1_HVT U371 ( .A1(n625), .A3(n627), .A2(n623), .A4(n624), .S0(n518), 
        .S1(n331), .Y(n622) );
  OA21X1_HVT U372 ( .A1(n789), .A2(n320), .A3(n558), .Y(n603) );
  NAND2X0_HVT U373 ( .A1(n756), .A2(n369), .Y(n370) );
  NAND2X0_HVT U374 ( .A1(n730), .A2(n516), .Y(n371) );
  NAND2X0_HVT U375 ( .A1(n371), .A2(n370), .Y(n729) );
  MUX41X1_HVT U376 ( .A1(n664), .A3(n661), .A2(n665), .A4(n663), .S0(n331), 
        .S1(n518), .Y(n660) );
  NAND2X0_HVT U377 ( .A1(n565), .A2(n467), .Y(n374) );
  NAND2X0_HVT U378 ( .A1(n19), .A2(n533), .Y(n375) );
  NAND2X0_HVT U379 ( .A1(n374), .A2(n375), .Y(n734) );
  MUX21X1_HVT U380 ( .A1(n523), .A2(n273), .S0(n457), .Y(n612) );
  NAND2X0_HVT U381 ( .A1(n274), .A2(n376), .Y(n377) );
  NAND2X0_HVT U382 ( .A1(n491), .A2(n410), .Y(n378) );
  NAND2X0_HVT U383 ( .A1(n377), .A2(n378), .Y(n779) );
  INVX1_HVT U384 ( .A(n593), .Y(n576) );
  NAND2X0_HVT U385 ( .A1(n470), .A2(n411), .Y(n379) );
  NAND2X0_HVT U386 ( .A1(n421), .A2(n218), .Y(n380) );
  NAND2X0_HVT U387 ( .A1(n379), .A2(n380), .Y(n723) );
  MUX41X1_HVT U388 ( .A1(n602), .A3(n601), .A2(n600), .A4(n599), .S0(n424), 
        .S1(n331), .Y(n598) );
  NAND2X0_HVT U389 ( .A1(n719), .A2(n381), .Y(n382) );
  NAND2X0_HVT U390 ( .A1(n720), .A2(n369), .Y(n383) );
  NAND2X0_HVT U391 ( .A1(n383), .A2(n382), .Y(n717) );
  NAND2X0_HVT U392 ( .A1(n311), .A2(n384), .Y(n385) );
  NAND2X0_HVT U393 ( .A1(n420), .A2(n514), .Y(n386) );
  INVX1_HVT U394 ( .A(n440), .Y(n392) );
  NAND2X0_HVT U395 ( .A1(n784), .A2(n245), .Y(n387) );
  MUX41X1_HVT U396 ( .A1(n687), .A3(n506), .A2(n308), .A4(n568), .S0(n216), 
        .S1(n536), .Y(n647) );
  NAND2X0_HVT U397 ( .A1(n619), .A2(n369), .Y(n388) );
  NAND2X0_HVT U398 ( .A1(n620), .A2(n517), .Y(n389) );
  NAND2X0_HVT U399 ( .A1(n388), .A2(n389), .Y(n618) );
  MUX21X1_HVT U400 ( .A1(n580), .A2(n523), .S0(n264), .Y(n766) );
  NAND2X0_HVT U401 ( .A1(n521), .A2(n394), .Y(n390) );
  MUX41X1_HVT U402 ( .A1(n774), .A3(n558), .A2(n659), .A4(n455), .S0(n392), 
        .S1(n535), .Y(n658) );
  MUX41X1_HVT U403 ( .A1(n313), .A3(n415), .A2(n387), .A4(n683), .S0(n140), 
        .S1(n416), .Y(n682) );
  INVX1_HVT U404 ( .A(n760), .Y(n540) );
  NBUFFX2_HVT U405 ( .A(in[4]), .Y(n395) );
  NAND2X0_HVT U406 ( .A1(n646), .A2(n392), .Y(n396) );
  NAND2X0_HVT U407 ( .A1(n645), .A2(n440), .Y(n397) );
  NAND2X0_HVT U408 ( .A1(n396), .A2(n397), .Y(n644) );
  NAND2X0_HVT U409 ( .A1(n540), .A2(n398), .Y(n399) );
  AND2X1_HVT U410 ( .A1(n399), .A2(n649), .Y(n650) );
  MUX41X1_HVT U411 ( .A1(n767), .A3(n505), .A2(n764), .A4(n542), .S0(n400), 
        .S1(n483), .Y(n663) );
  INVX1_HVT U412 ( .A(n595), .Y(n543) );
  NAND2X0_HVT U413 ( .A1(n746), .A2(n369), .Y(n401) );
  NAND2X0_HVT U414 ( .A1(n750), .A2(n516), .Y(n402) );
  NAND2X0_HVT U415 ( .A1(n402), .A2(n401), .Y(n745) );
  INVX1_HVT U416 ( .A(n588), .Y(n542) );
  NAND2X0_HVT U417 ( .A1(n738), .A2(n140), .Y(n403) );
  NAND2X0_HVT U418 ( .A1(n736), .A2(n440), .Y(n404) );
  NAND2X0_HVT U419 ( .A1(n404), .A2(n403), .Y(n735) );
  MUX41X1_HVT U420 ( .A1(n539), .A3(n545), .A2(n543), .A4(n564), .S0(n478), 
        .S1(n367), .Y(n750) );
  MUX41X1_HVT U421 ( .A1(n737), .A3(n546), .A2(n555), .A4(n335), .S0(n353), 
        .S1(n458), .Y(n736) );
  NAND2X0_HVT U422 ( .A1(n450), .A2(n451), .Y(out[1]) );
  INVX1_HVT U423 ( .A(n589), .Y(n552) );
  NAND2X0_HVT U424 ( .A1(n652), .A2(n498), .Y(n405) );
  NAND2X0_HVT U425 ( .A1(n660), .A2(n339), .Y(n406) );
  NAND2X0_HVT U426 ( .A1(n405), .A2(n406), .Y(out[4]) );
  INVX1_HVT U427 ( .A(n591), .Y(n538) );
  NAND2X0_HVT U428 ( .A1(n491), .A2(n327), .Y(n408) );
  INVX0_HVT U429 ( .A(n590), .Y(n559) );
  OR2X1_HVT U430 ( .A1(n242), .A2(n360), .Y(n743) );
  MUX41X1_HVT U431 ( .A1(n735), .A3(n745), .A2(n731), .A4(n739), .S0(n339), 
        .S1(n331), .Y(out[0]) );
  NAND2X0_HVT U432 ( .A1(n442), .A2(n441), .Y(out[6]) );
  NAND2X0_HVT U433 ( .A1(n675), .A2(n414), .Y(n412) );
  AND2X1_HVT U434 ( .A1(n412), .A2(n413), .Y(n429) );
  OR2X1_HVT U435 ( .A1(n424), .A2(n466), .Y(n413) );
  AND2X1_HVT U436 ( .A1(n519), .A2(n458), .Y(n414) );
  AND2X1_HVT U437 ( .A1(n422), .A2(n423), .Y(n415) );
  MUX41X1_HVT U438 ( .A1(n758), .A3(n765), .A2(n751), .A4(n612), .S0(n517), 
        .S1(n478), .Y(n611) );
  NAND2X0_HVT U439 ( .A1(n416), .A2(n776), .Y(n417) );
  NAND2X0_HVT U440 ( .A1(n341), .A2(n364), .Y(n418) );
  NAND2X0_HVT U441 ( .A1(n417), .A2(n418), .Y(n662) );
  MUX21X1_HVT U442 ( .A1(n523), .A2(n421), .S0(n216), .Y(n420) );
  NAND2X0_HVT U443 ( .A1(n486), .A2(n19), .Y(n422) );
  NAND2X0_HVT U444 ( .A1(n460), .A2(n212), .Y(n423) );
  NAND2X0_HVT U445 ( .A1(n365), .A2(n422), .Y(n485) );
  INVX0_HVT U446 ( .A(n779), .Y(n539) );
  NAND2X0_HVT U447 ( .A1(n681), .A2(n398), .Y(n475) );
  NAND2X0_HVT U448 ( .A1(n740), .A2(n369), .Y(n425) );
  NAND2X0_HVT U449 ( .A1(n742), .A2(n517), .Y(n426) );
  NAND2X0_HVT U450 ( .A1(n425), .A2(n426), .Y(n739) );
  NAND2X0_HVT U451 ( .A1(n672), .A2(n424), .Y(n428) );
  NAND2X0_HVT U452 ( .A1(n429), .A2(n428), .Y(n671) );
  INVX1_HVT U453 ( .A(n467), .Y(n458) );
  NAND2X0_HVT U454 ( .A1(n506), .A2(n211), .Y(n430) );
  NAND2X0_HVT U455 ( .A1(n699), .A2(n753), .Y(n431) );
  NAND2X0_HVT U456 ( .A1(n430), .A2(n431), .Y(n698) );
  NAND2X0_HVT U457 ( .A1(n655), .A2(n392), .Y(n434) );
  NAND2X0_HVT U458 ( .A1(n656), .A2(n400), .Y(n435) );
  NAND2X0_HVT U459 ( .A1(n434), .A2(n435), .Y(n654) );
  NBUFFX2_HVT U460 ( .A(n503), .Y(n437) );
  NAND2X0_HVT U461 ( .A1(n607), .A2(n283), .Y(n438) );
  NAND2X0_HVT U462 ( .A1(n608), .A2(n400), .Y(n439) );
  NAND2X0_HVT U463 ( .A1(n438), .A2(n439), .Y(n606) );
  NAND2X0_HVT U464 ( .A1(n613), .A2(n498), .Y(n441) );
  NAND2X0_HVT U465 ( .A1(n622), .A2(n339), .Y(n442) );
  NAND2X0_HVT U466 ( .A1(n500), .A2(n499), .Y(out[5]) );
  MUX41X1_HVT U467 ( .A1(n761), .A3(n509), .A2(n754), .A4(n317), .S0(n440), 
        .S1(n535), .Y(n617) );
  NAND2X0_HVT U468 ( .A1(n598), .A2(n498), .Y(n444) );
  NAND2X0_HVT U469 ( .A1(n605), .A2(in[6]), .Y(n445) );
  NAND2X0_HVT U470 ( .A1(n445), .A2(n444), .Y(out[7]) );
  XOR2X2_HVT U471 ( .A1(n469), .A2(n321), .Y(n754) );
  NAND2X0_HVT U472 ( .A1(n488), .A2(n449), .Y(n447) );
  NAND2X0_HVT U473 ( .A1(n478), .A2(n772), .Y(n448) );
  NAND2X0_HVT U474 ( .A1(n447), .A2(n448), .Y(n756) );
  NAND2X0_HVT U475 ( .A1(n711), .A2(n498), .Y(n450) );
  NAND2X0_HVT U476 ( .A1(n721), .A2(n339), .Y(n451) );
  MUX21X1_HVT U477 ( .A1(n118), .A2(n486), .S0(n361), .Y(n789) );
  NAND2X0_HVT U478 ( .A1(n603), .A2(n369), .Y(n452) );
  NAND2X0_HVT U479 ( .A1(n604), .A2(n517), .Y(n453) );
  NAND2X0_HVT U480 ( .A1(n452), .A2(n453), .Y(n602) );
  INVX1_HVT U481 ( .A(n587), .Y(n570) );
  INVX1_HVT U482 ( .A(n487), .Y(n459) );
  INVX1_HVT U483 ( .A(n459), .Y(n460) );
  MUX41X1_HVT U484 ( .A1(n312), .A3(n510), .A2(n741), .A4(n512), .S0(n477), 
        .S1(n367), .Y(n740) );
  NAND2X0_HVT U485 ( .A1(n676), .A2(n488), .Y(n466) );
  MUX21X1_HVT U486 ( .A1(n557), .A2(n677), .S0(n381), .Y(n676) );
  MUX41X1_HVT U487 ( .A1(n794), .A3(n437), .A2(n485), .A4(n569), .S0(n369), 
        .S1(n479), .Y(n599) );
  NAND2X0_HVT U488 ( .A1(n680), .A2(n477), .Y(n476) );
  NAND2X0_HVT U489 ( .A1(n475), .A2(n476), .Y(n679) );
  NAND2X0_HVT U490 ( .A1(n707), .A2(n516), .Y(n482) );
  NAND2X0_HVT U491 ( .A1(n481), .A2(n482), .Y(n704) );
  INVX1_HVT U492 ( .A(n490), .Y(n646) );
  INVX1_HVT U493 ( .A(n497), .Y(n536) );
  AND2X1_HVT U494 ( .A1(n390), .A2(n443), .Y(n484) );
  NAND2X0_HVT U495 ( .A1(n446), .A2(n274), .Y(n493) );
  NAND2X0_HVT U496 ( .A1(n308), .A2(n492), .Y(n494) );
  NAND2X0_HVT U497 ( .A1(n708), .A2(n511), .Y(n495) );
  NAND2X0_HVT U498 ( .A1(n495), .A2(n494), .Y(n707) );
  NAND2X0_HVT U499 ( .A1(n502), .A2(n501), .Y(out[2]) );
  MUX41X1_HVT U500 ( .A1(n781), .A3(n715), .A2(n549), .A4(n470), .S0(n283), 
        .S1(n320), .Y(n714) );
  NAND2X0_HVT U501 ( .A1(n629), .A2(n498), .Y(n499) );
  NAND2X0_HVT U502 ( .A1(n641), .A2(n339), .Y(n500) );
  NAND2X0_HVT U503 ( .A1(n690), .A2(n498), .Y(n501) );
  NAND2X0_HVT U504 ( .A1(n700), .A2(n339), .Y(n502) );
  AND2X1_HVT U505 ( .A1(n474), .A2(n743), .Y(n504) );
  MUX21X1_HVT U506 ( .A1(n560), .A2(n486), .S0(n532), .Y(n747) );
  AND2X1_HVT U507 ( .A1(n526), .A2(n726), .Y(n505) );
  MUX21X1_HVT U508 ( .A1(n474), .A2(n221), .S0(n338), .Y(n695) );
  MUX21X1_HVT U509 ( .A1(n359), .A2(n460), .S0(n330), .Y(n589) );
  MUX21X1_HVT U510 ( .A1(n394), .A2(n560), .S0(n330), .Y(n770) );
  NBUFFX2_HVT U511 ( .A(n795), .Y(n525) );
  MUX21X1_HVT U512 ( .A1(n568), .A2(n579), .S0(n140), .Y(n681) );
  MUX21X1_HVT U513 ( .A1(n273), .A2(n524), .S0(n393), .Y(n677) );
  MUX21X1_HVT U514 ( .A1(n524), .A2(n358), .S0(n327), .Y(n615) );
  MUX21X1_HVT U515 ( .A1(n454), .A2(n358), .S0(n212), .Y(n705) );
  AND2X1_HVT U516 ( .A1(n245), .A2(n686), .Y(n506) );
  XNOR2X1_HVT U517 ( .A1(n358), .A2(n457), .Y(n508) );
  AND2X1_HVT U518 ( .A1(n376), .A2(n513), .Y(n509) );
  MUX21X1_HVT U519 ( .A1(n461), .A2(n524), .S0(n212), .Y(n594) );
  MUX21X1_HVT U520 ( .A1(n372), .A2(n358), .S0(n216), .Y(n674) );
  NBUFFX2_HVT U521 ( .A(n583), .Y(n524) );
  NBUFFX2_HVT U522 ( .A(n533), .Y(n518) );
  MUX21X1_HVT U523 ( .A1(n713), .A2(n433), .S0(n364), .Y(n620) );
  XOR2X1_HVT U524 ( .A1(n338), .A2(n274), .Y(n752) );
  MUX21X1_HVT U525 ( .A1(n465), .A2(n407), .S0(n519), .Y(n632) );
  MUX21X1_HVT U526 ( .A1(n770), .A2(n484), .S0(n446), .Y(n656) );
  NAND2X0_HVT U527 ( .A1(n521), .A2(n394), .Y(n795) );
  AND2X1_HVT U528 ( .A1(n118), .A2(n329), .Y(n510) );
  NBUFFX2_HVT U529 ( .A(n796), .Y(n527) );
  XOR2X1_HVT U530 ( .A1(n338), .A2(n518), .Y(n757) );
  MUX21X1_HVT U531 ( .A1(n769), .A2(n596), .S0(n483), .Y(n591) );
  MUX21X1_HVT U532 ( .A1(n794), .A2(n436), .S0(n216), .Y(n673) );
  MUX21X1_HVT U533 ( .A1(n433), .A2(n487), .S0(n321), .Y(n593) );
  MUX21X1_HVT U534 ( .A1(n274), .A2(n273), .S0(n519), .Y(n708) );
  XNOR2X1_HVT U535 ( .A1(n497), .A2(n361), .Y(n511) );
  AND2X1_HVT U536 ( .A1(n523), .A2(n411), .Y(n512) );
  NBUFFX2_HVT U537 ( .A(n533), .Y(n532) );
  NAND2X0_HVT U538 ( .A1(n395), .A2(n337), .Y(n796) );
  MUX21X1_HVT U539 ( .A1(n437), .A2(n464), .S0(n376), .Y(n587) );
  MUX21X1_HVT U540 ( .A1(n527), .A2(n503), .S0(n321), .Y(n771) );
  MUX21X1_HVT U541 ( .A1(n342), .A2(n527), .S0(n321), .Y(n586) );
  INVX1_HVT U542 ( .A(n534), .Y(n533) );
  INVX0_HVT U543 ( .A(in[5]), .Y(n534) );
  NBUFFX2_HVT U544 ( .A(in[0]), .Y(n520) );
  NBUFFX2_HVT U545 ( .A(n305), .Y(n517) );
endmodule

