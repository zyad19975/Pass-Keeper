
module aes ( plaintext, key, clk, reset, start, cipher_text, ready );
  input [127:0] plaintext;
  input [127:0] key;
  output [127:0] cipher_text;
  input clk, reset, start;
  output ready;
  wire   n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, d, n6, n7, n8, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n1,
         n2, n3, n4, n5, n10, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n479, n481, n482, n483, n484, n485, n486, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n498, n499, n500, n501, n502,
         n503, n504, n506, n507, n508, n509, n511, n512, n513, n514, n516,
         n518, n520, n522, n524, n525, n526, n527, n528, n529, n530, n532,
         n534, n536, n538, n540, n541, n542, n543, n544, n545, n546, n548,
         n550, n553, n554, n555, n556, n558, n559, n560, n561, n562, n563,
         n564, n565, n567, n568, n569, n570, n571, n572, n574, n576, n577,
         n578, n579, n581, n582, n583, n584, n586, n587, n588, n593, n594,
         n600, n601, n602, n603, n604, n616, n617, n619, n620, n622, n628,
         n629, n630, n631, n632, n633, n634, n635, n637, n638, n639, n640,
         n642, n644, n645, n646, n647, n648, n649, n651, n653, n654, n655,
         n656, n658, n660, n661, n662, n663, n665, n667, n668, n669, n671,
         n672, n673, n674, n676, n679, n681, n682, n683, n684, n686, n687,
         n688, n689, n690, n692, n694, n695, n696, n697, n699, n701, n702,
         n704, n706, n707, n708, n709, n711, n712, n713, n714, n715, n716,
         n717, n719, n721, n723, n725, n728, n730, n732, n734, n736, n737,
         n738, n739, n741, n742, n743, n745, n747, n748, n749, n750, n751,
         n752, n753, n755, n756, n757, n758, n760, n762, n763, n764, n765,
         n767, n772, n774, n776, n780, n782, n783, n784, n785, n787, n789,
         n791, n794, n795, n796, n797, n799, n801, n802, n803, n804, n805,
         n806, n807, n809, n811, n812, n813, n814, n816, n818, n820, n822,
         n824, n825, n826, n827, n829, n831, n833, n837, n839, n840, n841,
         n842, n844, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923;
  wire   [127:0] adk_out0;
  wire   [127:0] adk_in;
  wire   [3:0] round_number;
  wire   [127:0] key_round;
  wire   [127:0] keyout;

  DFFX1_HVT d_reg ( .D(n289), .CLK(clk), .Q(d), .QN(n9) );
  DFFX1_HVT \round_number_reg[3]  ( .D(n288), .CLK(clk), .Q(round_number[3])
         );
  DFFX1_HVT \round_number_reg[0]  ( .D(n287), .CLK(clk), .Q(round_number[0]), 
        .QN(n8) );
  DFFX1_HVT \round_number_reg[1]  ( .D(n286), .CLK(clk), .Q(round_number[1]), 
        .QN(n7) );
  DFFX1_HVT \round_number_reg[2]  ( .D(n285), .CLK(clk), .Q(round_number[2]), 
        .QN(n6) );
  DFFX1_HVT \adk_in_reg[0]  ( .D(n284), .CLK(clk), .Q(adk_in[0]) );
  DFFX1_HVT \adk_in_reg[1]  ( .D(n283), .CLK(clk), .Q(adk_in[1]), .QN(n300) );
  DFFX1_HVT \adk_in_reg[2]  ( .D(n282), .CLK(clk), .Q(adk_in[2]) );
  DFFX1_HVT \adk_in_reg[3]  ( .D(n281), .CLK(clk), .Q(adk_in[3]) );
  DFFX1_HVT \adk_in_reg[4]  ( .D(n280), .CLK(clk), .Q(adk_in[4]) );
  DFFX1_HVT \adk_in_reg[5]  ( .D(n279), .CLK(clk), .Q(adk_in[5]) );
  DFFX1_HVT \adk_in_reg[6]  ( .D(n278), .CLK(clk), .Q(adk_in[6]) );
  DFFX1_HVT \adk_in_reg[7]  ( .D(n277), .CLK(clk), .Q(adk_in[7]) );
  DFFX1_HVT \adk_in_reg[8]  ( .D(n276), .CLK(clk), .Q(adk_in[8]) );
  DFFX1_HVT \adk_in_reg[9]  ( .D(n275), .CLK(clk), .Q(adk_in[9]), .QN(n296) );
  DFFX1_HVT \adk_in_reg[10]  ( .D(n274), .CLK(clk), .Q(adk_in[10]) );
  DFFX1_HVT \adk_in_reg[11]  ( .D(n273), .CLK(clk), .Q(adk_in[11]) );
  DFFX1_HVT \adk_in_reg[12]  ( .D(n272), .CLK(clk), .Q(adk_in[12]), .QN(n619)
         );
  DFFX1_HVT \adk_in_reg[13]  ( .D(n271), .CLK(clk), .Q(adk_in[13]) );
  DFFX1_HVT \adk_in_reg[14]  ( .D(n270), .CLK(clk), .Q(adk_in[14]) );
  DFFX1_HVT \adk_in_reg[15]  ( .D(n269), .CLK(clk), .Q(adk_in[15]), .QN(n604)
         );
  DFFX1_HVT \adk_in_reg[16]  ( .D(n268), .CLK(clk), .Q(adk_in[16]) );
  DFFX1_HVT \adk_in_reg[17]  ( .D(n267), .CLK(clk), .Q(adk_in[17]), .QN(n369)
         );
  DFFX1_HVT \adk_in_reg[18]  ( .D(n266), .CLK(clk), .Q(adk_in[18]) );
  DFFX1_HVT \adk_in_reg[19]  ( .D(n265), .CLK(clk), .Q(adk_in[19]) );
  DFFX1_HVT \adk_in_reg[20]  ( .D(n264), .CLK(clk), .Q(adk_in[20]) );
  DFFX1_HVT \adk_in_reg[21]  ( .D(n263), .CLK(clk), .Q(adk_in[21]) );
  DFFX1_HVT \adk_in_reg[22]  ( .D(n262), .CLK(clk), .Q(adk_in[22]) );
  DFFX1_HVT \adk_in_reg[23]  ( .D(n261), .CLK(clk), .Q(adk_in[23]) );
  DFFX1_HVT \adk_in_reg[24]  ( .D(n260), .CLK(clk), .Q(adk_in[24]) );
  DFFX1_HVT \adk_in_reg[25]  ( .D(n259), .CLK(clk), .Q(adk_in[25]) );
  DFFX1_HVT \adk_in_reg[26]  ( .D(n258), .CLK(clk), .Q(adk_in[26]) );
  DFFX1_HVT \adk_in_reg[27]  ( .D(n257), .CLK(clk), .Q(adk_in[27]) );
  DFFX1_HVT \adk_in_reg[28]  ( .D(n256), .CLK(clk), .Q(adk_in[28]), .QN(n630)
         );
  DFFX1_HVT \adk_in_reg[29]  ( .D(n255), .CLK(clk), .Q(adk_in[29]) );
  DFFX1_HVT \adk_in_reg[30]  ( .D(n254), .CLK(clk), .Q(adk_in[30]) );
  DFFX1_HVT \adk_in_reg[31]  ( .D(n253), .CLK(clk), .Q(adk_in[31]), .QN(n434)
         );
  DFFX1_HVT \adk_in_reg[32]  ( .D(n252), .CLK(clk), .Q(adk_in[32]) );
  DFFX1_HVT \adk_in_reg[33]  ( .D(n251), .CLK(clk), .Q(adk_in[33]), .QN(n4) );
  DFFX1_HVT \adk_in_reg[34]  ( .D(n250), .CLK(clk), .Q(adk_in[34]) );
  DFFX1_HVT \adk_in_reg[35]  ( .D(n249), .CLK(clk), .Q(adk_in[35]) );
  DFFX1_HVT \adk_in_reg[36]  ( .D(n248), .CLK(clk), .Q(adk_in[36]) );
  DFFX1_HVT \adk_in_reg[37]  ( .D(n247), .CLK(clk), .Q(adk_in[37]) );
  DFFX1_HVT \adk_in_reg[38]  ( .D(n246), .CLK(clk), .Q(adk_in[38]) );
  DFFX1_HVT \adk_in_reg[39]  ( .D(n245), .CLK(clk), .Q(adk_in[39]) );
  DFFX1_HVT \adk_in_reg[40]  ( .D(n244), .CLK(clk), .Q(adk_in[40]) );
  DFFX1_HVT \adk_in_reg[41]  ( .D(n243), .CLK(clk), .Q(adk_in[41]), .QN(n380)
         );
  DFFX1_HVT \adk_in_reg[42]  ( .D(n242), .CLK(clk), .Q(adk_in[42]) );
  DFFX1_HVT \adk_in_reg[43]  ( .D(n241), .CLK(clk), .Q(adk_in[43]) );
  DFFX1_HVT \adk_in_reg[44]  ( .D(n240), .CLK(clk), .Q(adk_in[44]) );
  DFFX1_HVT \adk_in_reg[45]  ( .D(n239), .CLK(clk), .Q(adk_in[45]) );
  DFFX1_HVT \adk_in_reg[46]  ( .D(n238), .CLK(clk), .Q(adk_in[46]) );
  DFFX1_HVT \adk_in_reg[47]  ( .D(n237), .CLK(clk), .Q(adk_in[47]) );
  DFFX1_HVT \adk_in_reg[48]  ( .D(n236), .CLK(clk), .Q(adk_in[48]) );
  DFFX1_HVT \adk_in_reg[49]  ( .D(n235), .CLK(clk), .Q(adk_in[49]), .QN(n436)
         );
  DFFX1_HVT \adk_in_reg[50]  ( .D(n234), .CLK(clk), .Q(adk_in[50]) );
  DFFX1_HVT \adk_in_reg[51]  ( .D(n233), .CLK(clk), .Q(adk_in[51]) );
  DFFX1_HVT \adk_in_reg[52]  ( .D(n232), .CLK(clk), .Q(adk_in[52]), .QN(n298)
         );
  DFFX1_HVT \adk_in_reg[53]  ( .D(n231), .CLK(clk), .Q(adk_in[53]) );
  DFFX1_HVT \adk_in_reg[54]  ( .D(n230), .CLK(clk), .Q(adk_in[54]) );
  DFFX1_HVT \adk_in_reg[55]  ( .D(n229), .CLK(clk), .Q(adk_in[55]), .QN(n689)
         );
  DFFX1_HVT \adk_in_reg[56]  ( .D(n228), .CLK(clk), .Q(adk_in[56]) );
  DFFX1_HVT \adk_in_reg[57]  ( .D(n227), .CLK(clk), .Q(adk_in[57]) );
  DFFX1_HVT \adk_in_reg[58]  ( .D(n226), .CLK(clk), .Q(adk_in[58]) );
  DFFX1_HVT \adk_in_reg[59]  ( .D(n225), .CLK(clk), .Q(adk_in[59]) );
  DFFX1_HVT \adk_in_reg[60]  ( .D(n224), .CLK(clk), .Q(adk_in[60]), .QN(n667)
         );
  DFFX1_HVT \adk_in_reg[61]  ( .D(n223), .CLK(clk), .Q(adk_in[61]) );
  DFFX1_HVT \adk_in_reg[62]  ( .D(n222), .CLK(clk), .Q(adk_in[62]) );
  DFFX1_HVT \adk_in_reg[63]  ( .D(n221), .CLK(clk), .Q(adk_in[63]) );
  DFFX1_HVT \adk_in_reg[64]  ( .D(n220), .CLK(clk), .Q(adk_in[64]) );
  DFFX1_HVT \adk_in_reg[65]  ( .D(n219), .CLK(clk), .Q(adk_in[65]) );
  DFFX1_HVT \adk_in_reg[66]  ( .D(n218), .CLK(clk), .Q(adk_in[66]) );
  DFFX1_HVT \adk_in_reg[67]  ( .D(n217), .CLK(clk), .Q(adk_in[67]) );
  DFFX1_HVT \adk_in_reg[68]  ( .D(n216), .CLK(clk), .Q(adk_in[68]) );
  DFFX1_HVT \adk_in_reg[69]  ( .D(n215), .CLK(clk), .Q(adk_in[69]) );
  DFFX1_HVT \adk_in_reg[70]  ( .D(n214), .CLK(clk), .Q(adk_in[70]) );
  DFFX1_HVT \adk_in_reg[71]  ( .D(n213), .CLK(clk), .Q(adk_in[71]), .QN(n558)
         );
  DFFX1_HVT \adk_in_reg[72]  ( .D(n212), .CLK(clk), .Q(adk_in[72]) );
  DFFX1_HVT \adk_in_reg[73]  ( .D(n211), .CLK(clk), .Q(adk_in[73]) );
  DFFX1_HVT \adk_in_reg[74]  ( .D(n210), .CLK(clk), .Q(adk_in[74]) );
  DFFX1_HVT \adk_in_reg[75]  ( .D(n209), .CLK(clk), .Q(adk_in[75]) );
  DFFX1_HVT \adk_in_reg[76]  ( .D(n208), .CLK(clk), .Q(adk_in[76]) );
  DFFX1_HVT \adk_in_reg[77]  ( .D(n207), .CLK(clk), .Q(adk_in[77]) );
  DFFX1_HVT \adk_in_reg[78]  ( .D(n206), .CLK(clk), .Q(adk_in[78]) );
  DFFX1_HVT \adk_in_reg[79]  ( .D(n205), .CLK(clk), .Q(adk_in[79]) );
  DFFX1_HVT \adk_in_reg[80]  ( .D(n204), .CLK(clk), .Q(adk_in[80]) );
  DFFX1_HVT \adk_in_reg[81]  ( .D(n203), .CLK(clk), .Q(adk_in[81]) );
  DFFX1_HVT \adk_in_reg[82]  ( .D(n202), .CLK(clk), .Q(adk_in[82]) );
  DFFX1_HVT \adk_in_reg[83]  ( .D(n201), .CLK(clk), .Q(adk_in[83]) );
  DFFX1_HVT \adk_in_reg[84]  ( .D(n200), .CLK(clk), .Q(adk_in[84]) );
  DFFX1_HVT \adk_in_reg[85]  ( .D(n199), .CLK(clk), .Q(adk_in[85]) );
  DFFX1_HVT \adk_in_reg[87]  ( .D(n197), .CLK(clk), .Q(adk_in[87]), .QN(n511)
         );
  DFFX1_HVT \adk_in_reg[88]  ( .D(n196), .CLK(clk), .Q(adk_in[88]) );
  DFFX1_HVT \adk_in_reg[89]  ( .D(n195), .CLK(clk), .Q(adk_in[89]) );
  DFFX1_HVT \adk_in_reg[90]  ( .D(n194), .CLK(clk), .Q(adk_in[90]) );
  DFFX1_HVT \adk_in_reg[91]  ( .D(n193), .CLK(clk), .Q(adk_in[91]) );
  DFFX1_HVT \adk_in_reg[92]  ( .D(n192), .CLK(clk), .Q(adk_in[92]), .QN(n484)
         );
  DFFX1_HVT \adk_in_reg[93]  ( .D(n191), .CLK(clk), .Q(adk_in[93]) );
  DFFX1_HVT \adk_in_reg[94]  ( .D(n190), .CLK(clk), .Q(adk_in[94]) );
  DFFX1_HVT \adk_in_reg[95]  ( .D(n189), .CLK(clk), .Q(adk_in[95]) );
  DFFX1_HVT \adk_in_reg[96]  ( .D(n188), .CLK(clk), .Q(adk_in[96]) );
  DFFX1_HVT \adk_in_reg[97]  ( .D(n187), .CLK(clk), .Q(adk_in[97]) );
  DFFX1_HVT \adk_in_reg[98]  ( .D(n186), .CLK(clk), .Q(adk_in[98]) );
  DFFX1_HVT \adk_in_reg[99]  ( .D(n185), .CLK(clk), .Q(adk_in[99]) );
  DFFX1_HVT \adk_in_reg[100]  ( .D(n184), .CLK(clk), .Q(adk_in[100]), .QN(n466) );
  DFFX1_HVT \adk_in_reg[101]  ( .D(n183), .CLK(clk), .Q(adk_in[101]) );
  DFFX1_HVT \adk_in_reg[102]  ( .D(n182), .CLK(clk), .Q(adk_in[102]) );
  DFFX1_HVT \adk_in_reg[103]  ( .D(n181), .CLK(clk), .Q(adk_in[103]) );
  DFFX1_HVT \adk_in_reg[104]  ( .D(n180), .CLK(clk), .Q(adk_in[104]) );
  DFFX1_HVT \adk_in_reg[105]  ( .D(n179), .CLK(clk), .Q(adk_in[105]), .QN(n409) );
  DFFX1_HVT \adk_in_reg[106]  ( .D(n178), .CLK(clk), .Q(adk_in[106]) );
  DFFX1_HVT \adk_in_reg[107]  ( .D(n177), .CLK(clk), .Q(adk_in[107]) );
  DFFX1_HVT \adk_in_reg[108]  ( .D(n176), .CLK(clk), .Q(adk_in[108]), .QN(n644) );
  DFFX1_HVT \adk_in_reg[109]  ( .D(n175), .CLK(clk), .Q(adk_in[109]) );
  DFFX1_HVT \adk_in_reg[110]  ( .D(n174), .CLK(clk), .Q(adk_in[110]) );
  DFFX1_HVT \adk_in_reg[111]  ( .D(n173), .CLK(clk), .Q(adk_in[111]), .QN(n594) );
  DFFX1_HVT \adk_in_reg[112]  ( .D(n172), .CLK(clk), .Q(adk_in[112]) );
  DFFX1_HVT \adk_in_reg[113]  ( .D(n171), .CLK(clk), .Q(adk_in[113]), .QN(n317) );
  DFFX1_HVT \adk_in_reg[114]  ( .D(n170), .CLK(clk), .Q(adk_in[114]), .QN(n741) );
  DFFX1_HVT \adk_in_reg[115]  ( .D(n169), .CLK(clk), .Q(adk_in[115]) );
  DFFX1_HVT \adk_in_reg[116]  ( .D(n168), .CLK(clk), .Q(adk_in[116]), .QN(n441) );
  DFFX1_HVT \adk_in_reg[117]  ( .D(n167), .CLK(clk), .Q(adk_in[117]) );
  DFFX1_HVT \adk_in_reg[118]  ( .D(n166), .CLK(clk), .Q(adk_in[118]) );
  DFFX1_HVT \adk_in_reg[119]  ( .D(n165), .CLK(clk), .Q(adk_in[119]) );
  DFFX1_HVT \adk_in_reg[120]  ( .D(n164), .CLK(clk), .Q(adk_in[120]) );
  DFFX1_HVT \adk_in_reg[121]  ( .D(n163), .CLK(clk), .Q(adk_in[121]), .QN(n513) );
  DFFX1_HVT \adk_in_reg[122]  ( .D(n162), .CLK(clk), .Q(adk_in[122]) );
  DFFX1_HVT \adk_in_reg[123]  ( .D(n161), .CLK(clk), .Q(adk_in[123]) );
  DFFX1_HVT \adk_in_reg[124]  ( .D(n160), .CLK(clk), .Q(adk_in[124]), .QN(n617) );
  DFFX1_HVT \adk_in_reg[125]  ( .D(n159), .CLK(clk), .Q(adk_in[125]) );
  DFFX1_HVT \adk_in_reg[126]  ( .D(n158), .CLK(clk), .Q(adk_in[126]) );
  DFFX1_HVT \adk_in_reg[127]  ( .D(n157), .CLK(clk), .Q(adk_in[127]), .QN(n488) );
  DFFX1_HVT \key_round_reg[0]  ( .D(n156), .CLK(clk), .Q(key_round[0]) );
  DFFX1_HVT \key_round_reg[1]  ( .D(n155), .CLK(clk), .Q(key_round[1]) );
  DFFX1_HVT \key_round_reg[2]  ( .D(n154), .CLK(clk), .Q(key_round[2]) );
  DFFX1_HVT \key_round_reg[3]  ( .D(n153), .CLK(clk), .Q(key_round[3]) );
  DFFX1_HVT \key_round_reg[4]  ( .D(n152), .CLK(clk), .Q(key_round[4]) );
  DFFX1_HVT \key_round_reg[5]  ( .D(n151), .CLK(clk), .Q(key_round[5]) );
  DFFX1_HVT \key_round_reg[6]  ( .D(n150), .CLK(clk), .Q(key_round[6]) );
  DFFX1_HVT \key_round_reg[7]  ( .D(n149), .CLK(clk), .Q(key_round[7]), .QN(
        n628) );
  DFFX1_HVT \key_round_reg[8]  ( .D(n148), .CLK(clk), .Q(key_round[8]) );
  DFFX1_HVT \key_round_reg[9]  ( .D(n147), .CLK(clk), .Q(key_round[9]), .QN(
        n310) );
  DFFX1_HVT \key_round_reg[10]  ( .D(n146), .CLK(clk), .Q(key_round[10]) );
  DFFX1_HVT \key_round_reg[11]  ( .D(n145), .CLK(clk), .Q(key_round[11]) );
  DFFX1_HVT \key_round_reg[12]  ( .D(n144), .CLK(clk), .Q(key_round[12]) );
  DFFX1_HVT \key_round_reg[13]  ( .D(n143), .CLK(clk), .Q(key_round[13]) );
  DFFX1_HVT \key_round_reg[14]  ( .D(n142), .CLK(clk), .Q(key_round[14]) );
  DFFX1_HVT \key_round_reg[15]  ( .D(n141), .CLK(clk), .Q(key_round[15]) );
  DFFX1_HVT \key_round_reg[16]  ( .D(n140), .CLK(clk), .Q(key_round[16]) );
  DFFX1_HVT \key_round_reg[17]  ( .D(n139), .CLK(clk), .Q(key_round[17]), .QN(
        n346) );
  DFFX1_HVT \key_round_reg[18]  ( .D(n138), .CLK(clk), .Q(key_round[18]), .QN(
        n587) );
  DFFX1_HVT \key_round_reg[19]  ( .D(n137), .CLK(clk), .Q(key_round[19]) );
  DFFX1_HVT \key_round_reg[20]  ( .D(n136), .CLK(clk), .Q(key_round[20]) );
  DFFX1_HVT \key_round_reg[21]  ( .D(n135), .CLK(clk), .Q(key_round[21]) );
  DFFX1_HVT \key_round_reg[22]  ( .D(n134), .CLK(clk), .Q(key_round[22]) );
  DFFX1_HVT \key_round_reg[23]  ( .D(n133), .CLK(clk), .Q(key_round[23]), .QN(
        n292) );
  DFFX1_HVT \key_round_reg[24]  ( .D(n132), .CLK(clk), .Q(key_round[24]) );
  DFFX1_HVT \key_round_reg[25]  ( .D(n131), .CLK(clk), .Q(key_round[25]) );
  DFFX1_HVT \key_round_reg[26]  ( .D(n130), .CLK(clk), .Q(key_round[26]) );
  DFFX1_HVT \key_round_reg[27]  ( .D(n129), .CLK(clk), .Q(key_round[27]) );
  DFFX1_HVT \key_round_reg[28]  ( .D(n128), .CLK(clk), .Q(key_round[28]) );
  DFFX1_HVT \key_round_reg[29]  ( .D(n127), .CLK(clk), .Q(key_round[29]) );
  DFFX1_HVT \key_round_reg[30]  ( .D(n126), .CLK(clk), .Q(key_round[30]) );
  DFFX1_HVT \key_round_reg[31]  ( .D(n125), .CLK(clk), .Q(key_round[31]), .QN(
        n701) );
  DFFX1_HVT \key_round_reg[32]  ( .D(n124), .CLK(clk), .Q(key_round[32]) );
  DFFX1_HVT \key_round_reg[33]  ( .D(n123), .CLK(clk), .Q(key_round[33]) );
  DFFX1_HVT \key_round_reg[34]  ( .D(n122), .CLK(clk), .Q(key_round[34]) );
  DFFX1_HVT \key_round_reg[35]  ( .D(n121), .CLK(clk), .Q(key_round[35]) );
  DFFX1_HVT \key_round_reg[36]  ( .D(n120), .CLK(clk), .Q(key_round[36]) );
  DFFX1_HVT \key_round_reg[37]  ( .D(n119), .CLK(clk), .Q(key_round[37]) );
  DFFX1_HVT \key_round_reg[38]  ( .D(n118), .CLK(clk), .Q(key_round[38]) );
  DFFX1_HVT \key_round_reg[39]  ( .D(n117), .CLK(clk), .Q(key_round[39]) );
  DFFX1_HVT \key_round_reg[40]  ( .D(n116), .CLK(clk), .Q(key_round[40]) );
  DFFX1_HVT \key_round_reg[41]  ( .D(n115), .CLK(clk), .Q(key_round[41]) );
  DFFX1_HVT \key_round_reg[42]  ( .D(n114), .CLK(clk), .Q(key_round[42]) );
  DFFX1_HVT \key_round_reg[43]  ( .D(n113), .CLK(clk), .Q(key_round[43]) );
  DFFX1_HVT \key_round_reg[44]  ( .D(n112), .CLK(clk), .Q(key_round[44]) );
  DFFX1_HVT \key_round_reg[45]  ( .D(n111), .CLK(clk), .Q(key_round[45]) );
  DFFX1_HVT \key_round_reg[46]  ( .D(n110), .CLK(clk), .Q(key_round[46]) );
  DFFX1_HVT \key_round_reg[47]  ( .D(n109), .CLK(clk), .Q(key_round[47]) );
  DFFX1_HVT \key_round_reg[48]  ( .D(n108), .CLK(clk), .Q(key_round[48]) );
  DFFX1_HVT \key_round_reg[49]  ( .D(n107), .CLK(clk), .Q(key_round[49]) );
  DFFX1_HVT \key_round_reg[50]  ( .D(n106), .CLK(clk), .Q(key_round[50]) );
  DFFX1_HVT \key_round_reg[51]  ( .D(n105), .CLK(clk), .Q(key_round[51]) );
  DFFX1_HVT \key_round_reg[52]  ( .D(n104), .CLK(clk), .Q(key_round[52]) );
  DFFX1_HVT \key_round_reg[53]  ( .D(n103), .CLK(clk), .Q(key_round[53]) );
  DFFX1_HVT \key_round_reg[54]  ( .D(n102), .CLK(clk), .Q(key_round[54]) );
  DFFX1_HVT \key_round_reg[55]  ( .D(n101), .CLK(clk), .Q(key_round[55]) );
  DFFX1_HVT \key_round_reg[56]  ( .D(n100), .CLK(clk), .Q(key_round[56]) );
  DFFX1_HVT \key_round_reg[57]  ( .D(n99), .CLK(clk), .Q(key_round[57]) );
  DFFX1_HVT \key_round_reg[58]  ( .D(n98), .CLK(clk), .Q(key_round[58]) );
  DFFX1_HVT \key_round_reg[59]  ( .D(n97), .CLK(clk), .Q(key_round[59]) );
  DFFX1_HVT \key_round_reg[60]  ( .D(n96), .CLK(clk), .Q(key_round[60]) );
  DFFX1_HVT \key_round_reg[61]  ( .D(n95), .CLK(clk), .Q(key_round[61]) );
  DFFX1_HVT \key_round_reg[62]  ( .D(n94), .CLK(clk), .Q(key_round[62]) );
  DFFX1_HVT \key_round_reg[63]  ( .D(n93), .CLK(clk), .Q(key_round[63]) );
  DFFX1_HVT \key_round_reg[64]  ( .D(n92), .CLK(clk), .Q(key_round[64]) );
  DFFX1_HVT \key_round_reg[65]  ( .D(n91), .CLK(clk), .Q(key_round[65]) );
  DFFX1_HVT \key_round_reg[66]  ( .D(n90), .CLK(clk), .Q(key_round[66]) );
  DFFX1_HVT \key_round_reg[67]  ( .D(n89), .CLK(clk), .Q(key_round[67]) );
  DFFX1_HVT \key_round_reg[68]  ( .D(n88), .CLK(clk), .Q(key_round[68]) );
  DFFX1_HVT \key_round_reg[69]  ( .D(n87), .CLK(clk), .Q(key_round[69]) );
  DFFX1_HVT \key_round_reg[70]  ( .D(n86), .CLK(clk), .Q(key_round[70]) );
  DFFX1_HVT \key_round_reg[71]  ( .D(n85), .CLK(clk), .Q(key_round[71]) );
  DFFX1_HVT \key_round_reg[72]  ( .D(n84), .CLK(clk), .Q(key_round[72]) );
  DFFX1_HVT \key_round_reg[73]  ( .D(n83), .CLK(clk), .Q(key_round[73]) );
  DFFX1_HVT \key_round_reg[74]  ( .D(n82), .CLK(clk), .Q(key_round[74]) );
  DFFX1_HVT \key_round_reg[75]  ( .D(n81), .CLK(clk), .Q(key_round[75]) );
  DFFX1_HVT \key_round_reg[76]  ( .D(n80), .CLK(clk), .Q(key_round[76]) );
  DFFX1_HVT \key_round_reg[77]  ( .D(n79), .CLK(clk), .Q(key_round[77]) );
  DFFX1_HVT \key_round_reg[78]  ( .D(n78), .CLK(clk), .Q(key_round[78]) );
  DFFX1_HVT \key_round_reg[79]  ( .D(n77), .CLK(clk), .Q(key_round[79]) );
  DFFX1_HVT \key_round_reg[80]  ( .D(n76), .CLK(clk), .Q(key_round[80]) );
  DFFX1_HVT \key_round_reg[81]  ( .D(n75), .CLK(clk), .Q(key_round[81]) );
  DFFX1_HVT \key_round_reg[82]  ( .D(n74), .CLK(clk), .Q(key_round[82]) );
  DFFX1_HVT \key_round_reg[83]  ( .D(n73), .CLK(clk), .Q(key_round[83]) );
  DFFX1_HVT \key_round_reg[84]  ( .D(n72), .CLK(clk), .Q(key_round[84]) );
  DFFX1_HVT \key_round_reg[85]  ( .D(n71), .CLK(clk), .Q(key_round[85]) );
  DFFX1_HVT \key_round_reg[86]  ( .D(n70), .CLK(clk), .Q(key_round[86]) );
  DFFX1_HVT \key_round_reg[87]  ( .D(n69), .CLK(clk), .Q(key_round[87]) );
  DFFX1_HVT \key_round_reg[88]  ( .D(n68), .CLK(clk), .Q(key_round[88]) );
  DFFX1_HVT \key_round_reg[89]  ( .D(n67), .CLK(clk), .Q(key_round[89]) );
  DFFX1_HVT \key_round_reg[90]  ( .D(n66), .CLK(clk), .Q(key_round[90]) );
  DFFX1_HVT \key_round_reg[91]  ( .D(n65), .CLK(clk), .Q(key_round[91]) );
  DFFX1_HVT \key_round_reg[92]  ( .D(n64), .CLK(clk), .Q(key_round[92]) );
  DFFX1_HVT \key_round_reg[93]  ( .D(n63), .CLK(clk), .Q(key_round[93]) );
  DFFX1_HVT \key_round_reg[94]  ( .D(n62), .CLK(clk), .Q(key_round[94]) );
  DFFX1_HVT \key_round_reg[95]  ( .D(n61), .CLK(clk), .Q(key_round[95]) );
  DFFX1_HVT \key_round_reg[96]  ( .D(n60), .CLK(clk), .Q(key_round[96]) );
  DFFX1_HVT \key_round_reg[97]  ( .D(n59), .CLK(clk), .Q(key_round[97]) );
  DFFX1_HVT \key_round_reg[98]  ( .D(n58), .CLK(clk), .Q(key_round[98]) );
  DFFX1_HVT \key_round_reg[99]  ( .D(n57), .CLK(clk), .Q(key_round[99]) );
  DFFX1_HVT \key_round_reg[100]  ( .D(n56), .CLK(clk), .Q(key_round[100]) );
  DFFX1_HVT \key_round_reg[101]  ( .D(n55), .CLK(clk), .Q(key_round[101]) );
  DFFX1_HVT \key_round_reg[102]  ( .D(n54), .CLK(clk), .Q(key_round[102]) );
  DFFX1_HVT \key_round_reg[103]  ( .D(n53), .CLK(clk), .Q(key_round[103]) );
  DFFX1_HVT \key_round_reg[104]  ( .D(n52), .CLK(clk), .Q(key_round[104]) );
  DFFX1_HVT \key_round_reg[105]  ( .D(n51), .CLK(clk), .Q(key_round[105]) );
  DFFX1_HVT \key_round_reg[106]  ( .D(n50), .CLK(clk), .Q(key_round[106]) );
  DFFX1_HVT \key_round_reg[107]  ( .D(n49), .CLK(clk), .Q(key_round[107]) );
  DFFX1_HVT \key_round_reg[108]  ( .D(n48), .CLK(clk), .Q(key_round[108]) );
  DFFX1_HVT \key_round_reg[109]  ( .D(n47), .CLK(clk), .Q(key_round[109]) );
  DFFX1_HVT \key_round_reg[110]  ( .D(n46), .CLK(clk), .Q(key_round[110]) );
  DFFX1_HVT \key_round_reg[111]  ( .D(n45), .CLK(clk), .Q(key_round[111]) );
  DFFX1_HVT \key_round_reg[112]  ( .D(n44), .CLK(clk), .Q(key_round[112]) );
  DFFX1_HVT \key_round_reg[113]  ( .D(n43), .CLK(clk), .Q(key_round[113]) );
  DFFX1_HVT \key_round_reg[114]  ( .D(n42), .CLK(clk), .Q(key_round[114]) );
  DFFX1_HVT \key_round_reg[115]  ( .D(n41), .CLK(clk), .Q(key_round[115]) );
  DFFX1_HVT \key_round_reg[116]  ( .D(n40), .CLK(clk), .Q(key_round[116]) );
  DFFX1_HVT \key_round_reg[117]  ( .D(n39), .CLK(clk), .Q(key_round[117]) );
  DFFX1_HVT \key_round_reg[118]  ( .D(n38), .CLK(clk), .Q(key_round[118]) );
  DFFX1_HVT \key_round_reg[119]  ( .D(n37), .CLK(clk), .Q(key_round[119]) );
  DFFX1_HVT \key_round_reg[120]  ( .D(n36), .CLK(clk), .Q(key_round[120]) );
  DFFX1_HVT \key_round_reg[121]  ( .D(n35), .CLK(clk), .Q(key_round[121]) );
  DFFX1_HVT \key_round_reg[122]  ( .D(n34), .CLK(clk), .Q(key_round[122]) );
  DFFX1_HVT \key_round_reg[123]  ( .D(n33), .CLK(clk), .Q(key_round[123]) );
  DFFX1_HVT \key_round_reg[124]  ( .D(n32), .CLK(clk), .Q(key_round[124]) );
  DFFX1_HVT \key_round_reg[125]  ( .D(n31), .CLK(clk), .Q(key_round[125]) );
  DFFX1_HVT \key_round_reg[126]  ( .D(n30), .CLK(clk), .Q(key_round[126]) );
  DFFX1_HVT \key_round_reg[127]  ( .D(n29), .CLK(clk), .Q(key_round[127]) );
  DFFX1_HVT ready_reg ( .D(n28), .CLK(clk), .Q(ready) );
  NOR4X1_HVT U3 ( .A1(round_number[0]), .A2(round_number[1]), .A3(
        round_number[2]), .A4(round_number[3]), .Y(n18) );
  AO22X1_HVT U8 ( .A1(n11), .A2(ready), .A3(n922), .A4(n921), .Y(n28) );
  AND2X1_HVT U9 ( .A1(n13), .A2(n14), .Y(n11) );
  AO222X1_HVT U10 ( .A1(keyout[127]), .A2(n895), .A3(key[127]), .A4(n869), 
        .A5(key_round[127]), .A6(n864), .Y(n29) );
  AO222X1_HVT U11 ( .A1(keyout[126]), .A2(n895), .A3(key[126]), .A4(n869), 
        .A5(key_round[126]), .A6(n864), .Y(n30) );
  AO222X1_HVT U12 ( .A1(keyout[125]), .A2(n895), .A3(key[125]), .A4(n869), 
        .A5(key_round[125]), .A6(n864), .Y(n31) );
  AO222X1_HVT U13 ( .A1(keyout[124]), .A2(n895), .A3(key[124]), .A4(n869), 
        .A5(key_round[124]), .A6(n864), .Y(n32) );
  AO222X1_HVT U14 ( .A1(keyout[123]), .A2(n895), .A3(key[123]), .A4(n869), 
        .A5(key_round[123]), .A6(n864), .Y(n33) );
  AO222X1_HVT U15 ( .A1(keyout[122]), .A2(n895), .A3(key[122]), .A4(n869), 
        .A5(key_round[122]), .A6(n864), .Y(n34) );
  AO222X1_HVT U16 ( .A1(keyout[121]), .A2(n895), .A3(key[121]), .A4(n869), 
        .A5(key_round[121]), .A6(n864), .Y(n35) );
  AO222X1_HVT U17 ( .A1(keyout[120]), .A2(n895), .A3(key[120]), .A4(n869), 
        .A5(key_round[120]), .A6(n864), .Y(n36) );
  AO222X1_HVT U18 ( .A1(keyout[119]), .A2(n895), .A3(key[119]), .A4(n869), 
        .A5(key_round[119]), .A6(n864), .Y(n37) );
  AO222X1_HVT U19 ( .A1(keyout[118]), .A2(n895), .A3(key[118]), .A4(n869), 
        .A5(key_round[118]), .A6(n864), .Y(n38) );
  AO222X1_HVT U20 ( .A1(keyout[117]), .A2(n895), .A3(key[117]), .A4(n869), 
        .A5(key_round[117]), .A6(n863), .Y(n39) );
  AO222X1_HVT U21 ( .A1(keyout[116]), .A2(n895), .A3(key[116]), .A4(n869), 
        .A5(key_round[116]), .A6(n863), .Y(n40) );
  AO222X1_HVT U22 ( .A1(keyout[115]), .A2(n896), .A3(key[115]), .A4(n870), 
        .A5(key_round[115]), .A6(n863), .Y(n41) );
  AO222X1_HVT U23 ( .A1(keyout[114]), .A2(n896), .A3(key[114]), .A4(n870), 
        .A5(key_round[114]), .A6(n863), .Y(n42) );
  AO222X1_HVT U24 ( .A1(keyout[113]), .A2(n896), .A3(key[113]), .A4(n870), 
        .A5(key_round[113]), .A6(n863), .Y(n43) );
  AO222X1_HVT U25 ( .A1(keyout[112]), .A2(n896), .A3(key[112]), .A4(n870), 
        .A5(key_round[112]), .A6(n863), .Y(n44) );
  AO222X1_HVT U26 ( .A1(keyout[111]), .A2(n896), .A3(key[111]), .A4(n870), 
        .A5(key_round[111]), .A6(n863), .Y(n45) );
  AO222X1_HVT U27 ( .A1(keyout[110]), .A2(n896), .A3(key[110]), .A4(n870), 
        .A5(key_round[110]), .A6(n863), .Y(n46) );
  AO222X1_HVT U28 ( .A1(keyout[109]), .A2(n896), .A3(key[109]), .A4(n870), 
        .A5(key_round[109]), .A6(n863), .Y(n47) );
  AO222X1_HVT U29 ( .A1(keyout[108]), .A2(n896), .A3(key[108]), .A4(n870), 
        .A5(key_round[108]), .A6(n863), .Y(n48) );
  AO222X1_HVT U30 ( .A1(keyout[107]), .A2(n896), .A3(key[107]), .A4(n870), 
        .A5(key_round[107]), .A6(n863), .Y(n49) );
  AO222X1_HVT U31 ( .A1(keyout[106]), .A2(n896), .A3(key[106]), .A4(n870), 
        .A5(key_round[106]), .A6(n863), .Y(n50) );
  AO222X1_HVT U32 ( .A1(keyout[105]), .A2(n896), .A3(key[105]), .A4(n870), 
        .A5(key_round[105]), .A6(n863), .Y(n51) );
  AO222X1_HVT U33 ( .A1(keyout[104]), .A2(n896), .A3(key[104]), .A4(n870), 
        .A5(key_round[104]), .A6(n862), .Y(n52) );
  AO222X1_HVT U34 ( .A1(keyout[103]), .A2(n897), .A3(key[103]), .A4(n871), 
        .A5(key_round[103]), .A6(n862), .Y(n53) );
  AO222X1_HVT U35 ( .A1(keyout[102]), .A2(n897), .A3(key[102]), .A4(n871), 
        .A5(key_round[102]), .A6(n862), .Y(n54) );
  AO222X1_HVT U36 ( .A1(keyout[101]), .A2(n897), .A3(key[101]), .A4(n871), 
        .A5(key_round[101]), .A6(n862), .Y(n55) );
  AO222X1_HVT U37 ( .A1(keyout[100]), .A2(n897), .A3(key[100]), .A4(n871), 
        .A5(key_round[100]), .A6(n862), .Y(n56) );
  AO222X1_HVT U38 ( .A1(keyout[99]), .A2(n897), .A3(key[99]), .A4(n871), .A5(
        key_round[99]), .A6(n862), .Y(n57) );
  AO222X1_HVT U39 ( .A1(keyout[98]), .A2(n897), .A3(key[98]), .A4(n871), .A5(
        key_round[98]), .A6(n862), .Y(n58) );
  AO222X1_HVT U40 ( .A1(keyout[97]), .A2(n897), .A3(key[97]), .A4(n871), .A5(
        key_round[97]), .A6(n862), .Y(n59) );
  AO222X1_HVT U41 ( .A1(keyout[96]), .A2(n897), .A3(key[96]), .A4(n871), .A5(
        key_round[96]), .A6(n862), .Y(n60) );
  AO222X1_HVT U42 ( .A1(keyout[95]), .A2(n897), .A3(key[95]), .A4(n871), .A5(
        key_round[95]), .A6(n862), .Y(n61) );
  AO222X1_HVT U43 ( .A1(keyout[94]), .A2(n897), .A3(key[94]), .A4(n871), .A5(
        key_round[94]), .A6(n862), .Y(n62) );
  AO222X1_HVT U44 ( .A1(keyout[93]), .A2(n897), .A3(key[93]), .A4(n871), .A5(
        key_round[93]), .A6(n862), .Y(n63) );
  AO222X1_HVT U45 ( .A1(keyout[92]), .A2(n897), .A3(key[92]), .A4(n871), .A5(
        key_round[92]), .A6(n862), .Y(n64) );
  AO222X1_HVT U46 ( .A1(keyout[91]), .A2(n898), .A3(key[91]), .A4(n872), .A5(
        key_round[91]), .A6(n861), .Y(n65) );
  AO222X1_HVT U47 ( .A1(keyout[90]), .A2(n898), .A3(key[90]), .A4(n872), .A5(
        key_round[90]), .A6(n861), .Y(n66) );
  AO222X1_HVT U48 ( .A1(keyout[89]), .A2(n898), .A3(key[89]), .A4(n872), .A5(
        key_round[89]), .A6(n861), .Y(n67) );
  AO222X1_HVT U49 ( .A1(keyout[88]), .A2(n898), .A3(key[88]), .A4(n872), .A5(
        key_round[88]), .A6(n861), .Y(n68) );
  AO222X1_HVT U50 ( .A1(keyout[87]), .A2(n898), .A3(key[87]), .A4(n872), .A5(
        key_round[87]), .A6(n861), .Y(n69) );
  AO222X1_HVT U51 ( .A1(keyout[86]), .A2(n898), .A3(key[86]), .A4(n872), .A5(
        key_round[86]), .A6(n861), .Y(n70) );
  AO222X1_HVT U52 ( .A1(keyout[85]), .A2(n898), .A3(key[85]), .A4(n872), .A5(
        key_round[85]), .A6(n861), .Y(n71) );
  AO222X1_HVT U53 ( .A1(keyout[84]), .A2(n898), .A3(key[84]), .A4(n872), .A5(
        key_round[84]), .A6(n861), .Y(n72) );
  AO222X1_HVT U54 ( .A1(keyout[83]), .A2(n898), .A3(key[83]), .A4(n872), .A5(
        key_round[83]), .A6(n861), .Y(n73) );
  AO222X1_HVT U55 ( .A1(keyout[82]), .A2(n898), .A3(key[82]), .A4(n872), .A5(
        key_round[82]), .A6(n861), .Y(n74) );
  AO222X1_HVT U56 ( .A1(keyout[81]), .A2(n898), .A3(key[81]), .A4(n872), .A5(
        key_round[81]), .A6(n861), .Y(n75) );
  AO222X1_HVT U57 ( .A1(keyout[80]), .A2(n898), .A3(key[80]), .A4(n872), .A5(
        key_round[80]), .A6(n861), .Y(n76) );
  AO222X1_HVT U58 ( .A1(n899), .A2(keyout[79]), .A3(key[79]), .A4(n873), .A5(
        key_round[79]), .A6(n861), .Y(n77) );
  AO222X1_HVT U59 ( .A1(keyout[78]), .A2(n899), .A3(key[78]), .A4(n873), .A5(
        key_round[78]), .A6(n860), .Y(n78) );
  AO222X1_HVT U60 ( .A1(keyout[77]), .A2(n899), .A3(key[77]), .A4(n873), .A5(
        key_round[77]), .A6(n860), .Y(n79) );
  AO222X1_HVT U61 ( .A1(keyout[76]), .A2(n899), .A3(key[76]), .A4(n873), .A5(
        key_round[76]), .A6(n860), .Y(n80) );
  AO222X1_HVT U62 ( .A1(keyout[75]), .A2(n899), .A3(key[75]), .A4(n873), .A5(
        key_round[75]), .A6(n860), .Y(n81) );
  AO222X1_HVT U63 ( .A1(keyout[74]), .A2(n899), .A3(key[74]), .A4(n873), .A5(
        key_round[74]), .A6(n860), .Y(n82) );
  AO222X1_HVT U64 ( .A1(keyout[73]), .A2(n899), .A3(key[73]), .A4(n873), .A5(
        key_round[73]), .A6(n860), .Y(n83) );
  AO222X1_HVT U65 ( .A1(keyout[72]), .A2(n899), .A3(key[72]), .A4(n873), .A5(
        key_round[72]), .A6(n860), .Y(n84) );
  AO222X1_HVT U66 ( .A1(keyout[71]), .A2(n899), .A3(key[71]), .A4(n873), .A5(
        key_round[71]), .A6(n860), .Y(n85) );
  AO222X1_HVT U67 ( .A1(keyout[70]), .A2(n899), .A3(key[70]), .A4(n873), .A5(
        key_round[70]), .A6(n860), .Y(n86) );
  AO222X1_HVT U68 ( .A1(keyout[69]), .A2(n899), .A3(key[69]), .A4(n873), .A5(
        key_round[69]), .A6(n860), .Y(n87) );
  AO222X1_HVT U69 ( .A1(keyout[68]), .A2(n899), .A3(key[68]), .A4(n873), .A5(
        key_round[68]), .A6(n860), .Y(n88) );
  AO222X1_HVT U70 ( .A1(keyout[67]), .A2(n900), .A3(key[67]), .A4(n874), .A5(
        key_round[67]), .A6(n860), .Y(n89) );
  AO222X1_HVT U71 ( .A1(keyout[66]), .A2(n900), .A3(key[66]), .A4(n874), .A5(
        key_round[66]), .A6(n860), .Y(n90) );
  AO222X1_HVT U72 ( .A1(keyout[65]), .A2(n900), .A3(key[65]), .A4(n874), .A5(
        key_round[65]), .A6(n859), .Y(n91) );
  AO222X1_HVT U73 ( .A1(keyout[64]), .A2(n900), .A3(key[64]), .A4(n874), .A5(
        key_round[64]), .A6(n859), .Y(n92) );
  AO222X1_HVT U74 ( .A1(keyout[63]), .A2(n900), .A3(key[63]), .A4(n874), .A5(
        key_round[63]), .A6(n859), .Y(n93) );
  AO222X1_HVT U75 ( .A1(keyout[62]), .A2(n900), .A3(key[62]), .A4(n874), .A5(
        key_round[62]), .A6(n859), .Y(n94) );
  AO222X1_HVT U76 ( .A1(keyout[61]), .A2(n900), .A3(key[61]), .A4(n874), .A5(
        key_round[61]), .A6(n859), .Y(n95) );
  AO222X1_HVT U77 ( .A1(keyout[60]), .A2(n900), .A3(key[60]), .A4(n874), .A5(
        key_round[60]), .A6(n859), .Y(n96) );
  AO222X1_HVT U78 ( .A1(keyout[59]), .A2(n900), .A3(key[59]), .A4(n874), .A5(
        key_round[59]), .A6(n859), .Y(n97) );
  AO222X1_HVT U79 ( .A1(keyout[58]), .A2(n900), .A3(key[58]), .A4(n874), .A5(
        key_round[58]), .A6(n859), .Y(n98) );
  AO222X1_HVT U80 ( .A1(keyout[57]), .A2(n900), .A3(key[57]), .A4(n874), .A5(
        key_round[57]), .A6(n859), .Y(n99) );
  AO222X1_HVT U81 ( .A1(keyout[56]), .A2(n900), .A3(key[56]), .A4(n874), .A5(
        key_round[56]), .A6(n859), .Y(n100) );
  AO222X1_HVT U82 ( .A1(keyout[55]), .A2(n901), .A3(key[55]), .A4(n875), .A5(
        key_round[55]), .A6(n859), .Y(n101) );
  AO222X1_HVT U83 ( .A1(keyout[54]), .A2(n901), .A3(key[54]), .A4(n875), .A5(
        key_round[54]), .A6(n859), .Y(n102) );
  AO222X1_HVT U84 ( .A1(keyout[53]), .A2(n901), .A3(key[53]), .A4(n875), .A5(
        key_round[53]), .A6(n859), .Y(n103) );
  AO222X1_HVT U85 ( .A1(keyout[52]), .A2(n901), .A3(key[52]), .A4(n875), .A5(
        key_round[52]), .A6(n858), .Y(n104) );
  AO222X1_HVT U86 ( .A1(n901), .A2(keyout[51]), .A3(key[51]), .A4(n875), .A5(
        key_round[51]), .A6(n858), .Y(n105) );
  AO222X1_HVT U87 ( .A1(keyout[50]), .A2(n901), .A3(key[50]), .A4(n875), .A5(
        key_round[50]), .A6(n858), .Y(n106) );
  AO222X1_HVT U88 ( .A1(keyout[49]), .A2(n901), .A3(key[49]), .A4(n875), .A5(
        key_round[49]), .A6(n858), .Y(n107) );
  AO222X1_HVT U89 ( .A1(keyout[48]), .A2(n901), .A3(key[48]), .A4(n875), .A5(
        key_round[48]), .A6(n858), .Y(n108) );
  AO222X1_HVT U90 ( .A1(keyout[47]), .A2(n901), .A3(key[47]), .A4(n875), .A5(
        key_round[47]), .A6(n858), .Y(n109) );
  AO222X1_HVT U91 ( .A1(keyout[46]), .A2(n901), .A3(key[46]), .A4(n875), .A5(
        key_round[46]), .A6(n858), .Y(n110) );
  AO222X1_HVT U92 ( .A1(keyout[45]), .A2(n901), .A3(key[45]), .A4(n875), .A5(
        key_round[45]), .A6(n858), .Y(n111) );
  AO222X1_HVT U93 ( .A1(keyout[44]), .A2(n901), .A3(key[44]), .A4(n875), .A5(
        key_round[44]), .A6(n858), .Y(n112) );
  AO222X1_HVT U94 ( .A1(keyout[43]), .A2(n902), .A3(key[43]), .A4(n876), .A5(
        key_round[43]), .A6(n858), .Y(n113) );
  AO222X1_HVT U95 ( .A1(keyout[42]), .A2(n902), .A3(key[42]), .A4(n876), .A5(
        key_round[42]), .A6(n858), .Y(n114) );
  AO222X1_HVT U96 ( .A1(keyout[41]), .A2(n902), .A3(key[41]), .A4(n876), .A5(
        key_round[41]), .A6(n858), .Y(n115) );
  AO222X1_HVT U97 ( .A1(keyout[40]), .A2(n902), .A3(key[40]), .A4(n876), .A5(
        key_round[40]), .A6(n858), .Y(n116) );
  AO222X1_HVT U98 ( .A1(keyout[39]), .A2(n902), .A3(key[39]), .A4(n876), .A5(
        key_round[39]), .A6(n857), .Y(n117) );
  AO222X1_HVT U99 ( .A1(keyout[38]), .A2(n902), .A3(key[38]), .A4(n876), .A5(
        key_round[38]), .A6(n857), .Y(n118) );
  AO222X1_HVT U100 ( .A1(keyout[37]), .A2(n902), .A3(key[37]), .A4(n876), .A5(
        key_round[37]), .A6(n857), .Y(n119) );
  AO222X1_HVT U101 ( .A1(keyout[36]), .A2(n902), .A3(key[36]), .A4(n876), .A5(
        key_round[36]), .A6(n857), .Y(n120) );
  AO222X1_HVT U102 ( .A1(keyout[35]), .A2(n902), .A3(key[35]), .A4(n876), .A5(
        key_round[35]), .A6(n857), .Y(n121) );
  AO222X1_HVT U103 ( .A1(keyout[34]), .A2(n902), .A3(key[34]), .A4(n876), .A5(
        key_round[34]), .A6(n857), .Y(n122) );
  AO222X1_HVT U104 ( .A1(keyout[33]), .A2(n902), .A3(key[33]), .A4(n876), .A5(
        key_round[33]), .A6(n857), .Y(n123) );
  AO222X1_HVT U105 ( .A1(keyout[32]), .A2(n902), .A3(key[32]), .A4(n876), .A5(
        key_round[32]), .A6(n857), .Y(n124) );
  AO222X1_HVT U106 ( .A1(keyout[31]), .A2(n903), .A3(key[31]), .A4(n877), .A5(
        key_round[31]), .A6(n857), .Y(n125) );
  AO222X1_HVT U107 ( .A1(keyout[30]), .A2(n903), .A3(key[30]), .A4(n877), .A5(
        key_round[30]), .A6(n857), .Y(n126) );
  AO222X1_HVT U108 ( .A1(keyout[29]), .A2(n903), .A3(key[29]), .A4(n877), .A5(
        key_round[29]), .A6(n857), .Y(n127) );
  AO222X1_HVT U109 ( .A1(keyout[28]), .A2(n903), .A3(key[28]), .A4(n877), .A5(
        key_round[28]), .A6(n857), .Y(n128) );
  AO222X1_HVT U110 ( .A1(keyout[27]), .A2(n903), .A3(key[27]), .A4(n877), .A5(
        key_round[27]), .A6(n857), .Y(n129) );
  AO222X1_HVT U111 ( .A1(keyout[26]), .A2(n903), .A3(key[26]), .A4(n877), .A5(
        key_round[26]), .A6(n856), .Y(n130) );
  AO222X1_HVT U112 ( .A1(keyout[25]), .A2(n903), .A3(key[25]), .A4(n877), .A5(
        key_round[25]), .A6(n856), .Y(n131) );
  AO222X1_HVT U113 ( .A1(keyout[24]), .A2(n903), .A3(key[24]), .A4(n877), .A5(
        key_round[24]), .A6(n856), .Y(n132) );
  AO222X1_HVT U114 ( .A1(keyout[23]), .A2(n903), .A3(key[23]), .A4(n877), .A5(
        key_round[23]), .A6(n856), .Y(n133) );
  AO222X1_HVT U115 ( .A1(keyout[22]), .A2(n903), .A3(key[22]), .A4(n877), .A5(
        key_round[22]), .A6(n856), .Y(n134) );
  AO222X1_HVT U116 ( .A1(keyout[21]), .A2(n903), .A3(key[21]), .A4(n877), .A5(
        key_round[21]), .A6(n856), .Y(n135) );
  AO222X1_HVT U117 ( .A1(keyout[20]), .A2(n903), .A3(key[20]), .A4(n877), .A5(
        key_round[20]), .A6(n856), .Y(n136) );
  AO222X1_HVT U118 ( .A1(keyout[19]), .A2(n904), .A3(key[19]), .A4(n878), .A5(
        key_round[19]), .A6(n856), .Y(n137) );
  AO222X1_HVT U119 ( .A1(keyout[18]), .A2(n904), .A3(key[18]), .A4(n878), .A5(
        key_round[18]), .A6(n856), .Y(n138) );
  AO222X1_HVT U120 ( .A1(keyout[17]), .A2(n904), .A3(key[17]), .A4(n878), .A5(
        key_round[17]), .A6(n856), .Y(n139) );
  AO222X1_HVT U121 ( .A1(keyout[16]), .A2(n904), .A3(key[16]), .A4(n878), .A5(
        key_round[16]), .A6(n856), .Y(n140) );
  AO222X1_HVT U122 ( .A1(keyout[15]), .A2(n904), .A3(key[15]), .A4(n878), .A5(
        key_round[15]), .A6(n856), .Y(n141) );
  AO222X1_HVT U123 ( .A1(keyout[14]), .A2(n904), .A3(key[14]), .A4(n878), .A5(
        key_round[14]), .A6(n856), .Y(n142) );
  AO222X1_HVT U124 ( .A1(keyout[13]), .A2(n904), .A3(key[13]), .A4(n878), .A5(
        key_round[13]), .A6(n855), .Y(n143) );
  AO222X1_HVT U125 ( .A1(keyout[12]), .A2(n904), .A3(key[12]), .A4(n878), .A5(
        key_round[12]), .A6(n855), .Y(n144) );
  AO222X1_HVT U126 ( .A1(keyout[11]), .A2(n904), .A3(key[11]), .A4(n878), .A5(
        key_round[11]), .A6(n855), .Y(n145) );
  AO222X1_HVT U127 ( .A1(keyout[10]), .A2(n904), .A3(key[10]), .A4(n878), .A5(
        key_round[10]), .A6(n855), .Y(n146) );
  AO222X1_HVT U128 ( .A1(keyout[9]), .A2(n904), .A3(key[9]), .A4(n878), .A5(
        key_round[9]), .A6(n855), .Y(n147) );
  AO222X1_HVT U129 ( .A1(keyout[8]), .A2(n904), .A3(key[8]), .A4(n878), .A5(
        key_round[8]), .A6(n855), .Y(n148) );
  AO222X1_HVT U130 ( .A1(keyout[7]), .A2(n905), .A3(key[7]), .A4(n879), .A5(
        key_round[7]), .A6(n855), .Y(n149) );
  AO222X1_HVT U131 ( .A1(keyout[6]), .A2(n905), .A3(key[6]), .A4(n879), .A5(
        key_round[6]), .A6(n855), .Y(n150) );
  AO222X1_HVT U132 ( .A1(keyout[5]), .A2(n905), .A3(key[5]), .A4(n879), .A5(
        key_round[5]), .A6(n855), .Y(n151) );
  AO222X1_HVT U133 ( .A1(keyout[4]), .A2(n905), .A3(key[4]), .A4(n879), .A5(
        key_round[4]), .A6(n855), .Y(n152) );
  AO222X1_HVT U134 ( .A1(keyout[3]), .A2(n905), .A3(key[3]), .A4(n879), .A5(
        key_round[3]), .A6(n855), .Y(n153) );
  AO222X1_HVT U135 ( .A1(keyout[2]), .A2(n905), .A3(key[2]), .A4(n879), .A5(
        key_round[2]), .A6(n855), .Y(n154) );
  AO222X1_HVT U136 ( .A1(keyout[1]), .A2(n905), .A3(key[1]), .A4(n879), .A5(
        key_round[1]), .A6(n855), .Y(n155) );
  AO222X1_HVT U137 ( .A1(keyout[0]), .A2(n905), .A3(key[0]), .A4(n879), .A5(
        key_round[0]), .A6(n854), .Y(n156) );
  AO222X1_HVT U145 ( .A1(n906), .A2(n931), .A3(adk_out0[120]), .A4(n880), .A5(
        adk_in[120]), .A6(n854), .Y(n164) );
  AO222X1_HVT U146 ( .A1(n906), .A2(n932), .A3(adk_out0[119]), .A4(n880), .A5(
        adk_in[119]), .A6(n854), .Y(n165) );
  AO222X1_HVT U147 ( .A1(n906), .A2(n933), .A3(adk_out0[118]), .A4(n880), .A5(
        adk_in[118]), .A6(n854), .Y(n166) );
  AO222X1_HVT U151 ( .A1(n906), .A2(n937), .A3(adk_out0[114]), .A4(n880), .A5(
        adk_in[114]), .A6(n853), .Y(n170) );
  AO222X1_HVT U153 ( .A1(n906), .A2(n939), .A3(adk_out0[112]), .A4(n880), .A5(
        adk_in[112]), .A6(n853), .Y(n172) );
  AO222X1_HVT U155 ( .A1(n907), .A2(n941), .A3(adk_out0[110]), .A4(n881), .A5(
        adk_in[110]), .A6(n853), .Y(n174) );
  AO222X1_HVT U163 ( .A1(n907), .A2(n949), .A3(adk_out0[102]), .A4(n881), .A5(
        adk_in[102]), .A6(n852), .Y(n182) );
  AO222X1_HVT U165 ( .A1(n907), .A2(n951), .A3(adk_out0[100]), .A4(n881), .A5(
        adk_in[100]), .A6(n852), .Y(n184) );
  AO222X1_HVT U167 ( .A1(n908), .A2(n953), .A3(adk_out0[98]), .A4(n882), .A5(
        adk_in[98]), .A6(n852), .Y(n186) );
  AO222X1_HVT U172 ( .A1(n908), .A2(n958), .A3(adk_out0[93]), .A4(n882), .A5(
        adk_in[93]), .A6(n852), .Y(n191) );
  AO222X1_HVT U177 ( .A1(n908), .A2(n963), .A3(adk_out0[88]), .A4(n882), .A5(
        adk_in[88]), .A6(n851), .Y(n196) );
  AO222X1_HVT U179 ( .A1(n909), .A2(n965), .A3(adk_out0[86]), .A4(n883), .A5(
        adk_in[86]), .A6(n851), .Y(n198) );
  AO222X1_HVT U183 ( .A1(n909), .A2(n969), .A3(adk_out0[82]), .A4(n883), .A5(
        adk_in[82]), .A6(n851), .Y(n202) );
  AO222X1_HVT U184 ( .A1(n909), .A2(n970), .A3(adk_out0[81]), .A4(n883), .A5(
        adk_in[81]), .A6(n851), .Y(n203) );
  AO222X1_HVT U193 ( .A1(n979), .A2(n910), .A3(adk_out0[72]), .A4(n884), .A5(
        adk_in[72]), .A6(n850), .Y(n212) );
  AO222X1_HVT U195 ( .A1(n910), .A2(n981), .A3(adk_out0[70]), .A4(n884), .A5(
        adk_in[70]), .A6(n850), .Y(n214) );
  AO222X1_HVT U211 ( .A1(n911), .A2(n997), .A3(adk_out0[54]), .A4(n885), .A5(
        adk_in[54]), .A6(n849), .Y(n230) );
  AO222X1_HVT U212 ( .A1(n998), .A2(n911), .A3(adk_out0[53]), .A4(n885), .A5(
        adk_in[53]), .A6(n849), .Y(n231) );
  AO222X1_HVT U223 ( .A1(n912), .A2(n1009), .A3(adk_out0[42]), .A4(n886), .A5(
        adk_in[42]), .A6(n362), .Y(n242) );
  AO222X1_HVT U225 ( .A1(n912), .A2(n1011), .A3(adk_out0[40]), .A4(n886), .A5(
        adk_in[40]), .A6(n850), .Y(n244) );
  AO222X1_HVT U227 ( .A1(n913), .A2(n1013), .A3(adk_out0[38]), .A4(n887), .A5(
        adk_in[38]), .A6(n864), .Y(n246) );
  AO222X1_HVT U231 ( .A1(n913), .A2(n1017), .A3(adk_out0[34]), .A4(n887), .A5(
        adk_in[34]), .A6(n848), .Y(n250) );
  AO222X1_HVT U233 ( .A1(n913), .A2(n1019), .A3(adk_out0[32]), .A4(n887), .A5(
        adk_in[32]), .A6(n848), .Y(n252) );
  AO222X1_HVT U236 ( .A1(n913), .A2(n1022), .A3(adk_out0[29]), .A4(n887), .A5(
        adk_in[29]), .A6(n848), .Y(n255) );
  AO222X1_HVT U239 ( .A1(n914), .A2(n1025), .A3(adk_out0[26]), .A4(n888), .A5(
        adk_in[26]), .A6(n848), .Y(n258) );
  AO222X1_HVT U241 ( .A1(n1027), .A2(n914), .A3(adk_out0[24]), .A4(n888), .A5(
        adk_in[24]), .A6(n847), .Y(n260) );
  AO222X1_HVT U243 ( .A1(n914), .A2(n1029), .A3(adk_out0[22]), .A4(n888), .A5(
        adk_in[22]), .A6(n847), .Y(n262) );
  AO222X1_HVT U244 ( .A1(n914), .A2(n1030), .A3(adk_out0[21]), .A4(n888), .A5(
        adk_in[21]), .A6(n847), .Y(n263) );
  AO222X1_HVT U248 ( .A1(n914), .A2(n1034), .A3(adk_out0[17]), .A4(n888), .A5(
        adk_in[17]), .A6(n847), .Y(n267) );
  AO222X1_HVT U249 ( .A1(n914), .A2(n1035), .A3(adk_out0[16]), .A4(n888), .A5(
        adk_in[16]), .A6(n847), .Y(n268) );
  AO222X1_HVT U251 ( .A1(n1037), .A2(n915), .A3(adk_out0[14]), .A4(n889), .A5(
        adk_in[14]), .A6(n847), .Y(n270) );
  AO222X1_HVT U255 ( .A1(n1041), .A2(n915), .A3(adk_out0[10]), .A4(n889), .A5(
        adk_in[10]), .A6(n846), .Y(n274) );
  AO222X1_HVT U258 ( .A1(n915), .A2(n1044), .A3(adk_out0[7]), .A4(n889), .A5(
        adk_in[7]), .A6(n846), .Y(n277) );
  AO222X1_HVT U263 ( .A1(n916), .A2(n1049), .A3(adk_out0[2]), .A4(n890), .A5(
        adk_in[2]), .A6(n846), .Y(n282) );
  AO222X1_HVT U265 ( .A1(n1051), .A2(n916), .A3(adk_out0[0]), .A4(n890), .A5(
        adk_in[0]), .A6(n846), .Y(n284) );
  AND2X1_HVT U266 ( .A1(n865), .A2(n18), .Y(n16) );
  NOR2X0_HVT U267 ( .A1(n846), .A2(n18), .Y(n15) );
  AO22X1_HVT U268 ( .A1(round_number[2]), .A2(n19), .A3(n20), .A4(n21), .Y(
        n285) );
  AND2X1_HVT U269 ( .A1(round_number[1]), .A2(n6), .Y(n20) );
  AO22X1_HVT U270 ( .A1(round_number[1]), .A2(n22), .A3(n21), .A4(n7), .Y(n286) );
  AO22X1_HVT U271 ( .A1(n23), .A2(round_number[0]), .A3(n867), .A4(n8), .Y(
        n287) );
  AO22X1_HVT U272 ( .A1(round_number[3]), .A2(n19), .A3(n24), .A4(
        round_number[2]), .Y(n288) );
  AND2X1_HVT U273 ( .A1(n21), .A2(round_number[1]), .Y(n24) );
  AND2X1_HVT U274 ( .A1(round_number[0]), .A2(n866), .Y(n21) );
  AO21X1_HVT U275 ( .A1(n868), .A2(n7), .A3(n22), .Y(n19) );
  AO21X1_HVT U276 ( .A1(n868), .A2(n8), .A3(n23), .Y(n22) );
  AOI21X1_HVT U277 ( .A1(start), .A2(n923), .A3(n868), .Y(n23) );
  OR2X1_HVT U278 ( .A1(n25), .A2(reset), .Y(n17) );
  NAND2X0_HVT U279 ( .A1(n26), .A2(n13), .Y(n289) );
  AND2X1_HVT U280 ( .A1(n921), .A2(n12), .Y(n13) );
  NAND4X0_HVT U281 ( .A1(n8), .A2(n6), .A3(n9), .A4(n27), .Y(n12) );
  AND2X1_HVT U282 ( .A1(round_number[3]), .A2(round_number[1]), .Y(n27) );
  AO21X1_HVT U283 ( .A1(start), .A2(n923), .A3(n9), .Y(n26) );
  NAND3X0_HVT U284 ( .A1(n25), .A2(n921), .A3(d), .Y(n14) );
  OA21X1_HVT U285 ( .A1(round_number[1]), .A2(round_number[2]), .A3(
        round_number[3]), .Y(n25) );
  add_round_keys_0 adk_0 ( .state(plaintext), .subkey(key), .out(adk_out0) );
  round r1 ( .in({n489, adk_in[126:122], n514, adk_in[120:117], n442, 
        adk_in[115], n742, n318, adk_in[112:109], n645, adk_in[107:106], n410, 
        adk_in[104:101], n467, adk_in[99:93], n485, adk_in[91:88], n512, 
        adk_in[86:72], n559, adk_in[70:61], n668, adk_in[59:56], n690, 
        adk_in[54:53], n299, adk_in[51:50], n437, adk_in[48:42], n381, 
        adk_in[40:34], n5, adk_in[32], n435, adk_in[30:29], n631, 
        adk_in[27:18], n370, adk_in[16:13], n620, adk_in[11:10], n297, 
        adk_in[8:2], n301, adk_in[0]}), .round_num(round_number), .keyin({
        key_round[127:32], n702, key_round[30:24], n293, key_round[22:19], 
        n588, n347, key_round[16:10], n311, key_round[8], n629, key_round[6:0]}), .keyout(keyout), .out({n924, n925, n926, n927, n928, n929, n930, n931, n932, 
        n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, 
        n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, 
        n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
        n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
        n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
        n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
        n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
        n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
        n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
        n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
        n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051}) );
  DFFX1_HVT \adk_in_reg[86]  ( .D(n198), .CLK(clk), .Q(adk_in[86]) );
  NBUFFX16_HVT U4 ( .A(n987), .Y(cipher_text[64]) );
  OAI222X2_HVT U5 ( .A1(n669), .A2(n600), .A3(n601), .A4(n602), .A5(n604), 
        .A6(n603), .Y(n269) );
  NBUFFX4_HVT U6 ( .A(n973), .Y(cipher_text[78]) );
  NAND2X0_HVT U7 ( .A1(n294), .A2(n927), .Y(n1) );
  NAND2X0_HVT U138 ( .A1(adk_out0[124]), .A2(n890), .Y(n2) );
  NAND2X0_HVT U139 ( .A1(n295), .A2(n362), .Y(n3) );
  NAND3X0_HVT U140 ( .A1(n1), .A2(n2), .A3(n3), .Y(n160) );
  INVX1_HVT U141 ( .A(n616), .Y(n294) );
  INVX1_HVT U142 ( .A(n891), .Y(n890) );
  INVX1_HVT U143 ( .A(n4), .Y(n5) );
  NBUFFX4_HVT U144 ( .A(n1002), .Y(cipher_text[49]) );
  NBUFFX4_HVT U148 ( .A(n964), .Y(cipher_text[87]) );
  INVX0_HVT U149 ( .A(n975), .Y(n739) );
  NBUFFX16_HVT U150 ( .A(n984), .Y(cipher_text[67]) );
  NAND2X0_HVT U152 ( .A1(n964), .A2(n909), .Y(n10) );
  NAND2X0_HVT U154 ( .A1(adk_out0[87]), .A2(n883), .Y(n290) );
  NAND2X0_HVT U156 ( .A1(adk_in[87]), .A2(n851), .Y(n291) );
  NAND3X0_HVT U157 ( .A1(n10), .A2(n290), .A3(n291), .Y(n197) );
  INVX1_HVT U158 ( .A(n674), .Y(cipher_text[8]) );
  INVX1_HVT U159 ( .A(n1043), .Y(n674) );
  NBUFFX4_HVT U160 ( .A(n1007), .Y(cipher_text[44]) );
  INVX2_HVT U161 ( .A(n346), .Y(n347) );
  INVX1_HVT U162 ( .A(n663), .Y(cipher_text[95]) );
  INVX1_HVT U164 ( .A(n441), .Y(n442) );
  INVX2_HVT U166 ( .A(n434), .Y(n435) );
  NBUFFX2_HVT U168 ( .A(n1023), .Y(cipher_text[28]) );
  NBUFFX16_HVT U169 ( .A(n1032), .Y(cipher_text[19]) );
  NBUFFX2_HVT U170 ( .A(n1003), .Y(cipher_text[48]) );
  NBUFFX2_HVT U171 ( .A(n982), .Y(cipher_text[69]) );
  NBUFFX16_HVT U173 ( .A(n937), .Y(cipher_text[114]) );
  INVX1_HVT U174 ( .A(n617), .Y(n295) );
  INVX1_HVT U175 ( .A(n292), .Y(n293) );
  INVX2_HVT U176 ( .A(n689), .Y(n690) );
  INVX1_HVT U178 ( .A(n296), .Y(n297) );
  INVX1_HVT U180 ( .A(n298), .Y(n299) );
  INVX1_HVT U181 ( .A(n300), .Y(n301) );
  INVX0_HVT U182 ( .A(n944), .Y(n807) );
  NBUFFX2_HVT U185 ( .A(n946), .Y(cipher_text[105]) );
  INVX0_HVT U186 ( .A(n829), .Y(n302) );
  NAND2X0_HVT U187 ( .A1(n906), .A2(n928), .Y(n303) );
  NAND2X0_HVT U188 ( .A1(adk_out0[123]), .A2(n880), .Y(n304) );
  NAND2X0_HVT U189 ( .A1(adk_in[123]), .A2(n854), .Y(n305) );
  NAND3X0_HVT U190 ( .A1(n303), .A2(n304), .A3(n305), .Y(n161) );
  INVX1_HVT U191 ( .A(n667), .Y(n668) );
  INVX1_HVT U192 ( .A(n466), .Y(n467) );
  INVX1_HVT U194 ( .A(n484), .Y(n485) );
  INVX1_HVT U196 ( .A(n630), .Y(n631) );
  NBUFFX2_HVT U197 ( .A(n935), .Y(cipher_text[116]) );
  NBUFFX2_HVT U198 ( .A(n1004), .Y(cipher_text[47]) );
  NBUFFX2_HVT U199 ( .A(n996), .Y(cipher_text[55]) );
  INVX0_HVT U200 ( .A(n967), .Y(n837) );
  INVX1_HVT U201 ( .A(n488), .Y(n489) );
  AND2X1_HVT U202 ( .A1(n673), .A2(n672), .Y(n306) );
  INVX0_HVT U203 ( .A(n1008), .Y(n816) );
  INVX1_HVT U204 ( .A(n868), .Y(n362) );
  INVX0_HVT U205 ( .A(n966), .Y(n842) );
  INVX1_HVT U206 ( .A(n496), .Y(cipher_text[13]) );
  INVX1_HVT U207 ( .A(n1038), .Y(n496) );
  INVX0_HVT U208 ( .A(n1033), .Y(n509) );
  NAND2X0_HVT U209 ( .A1(n926), .A2(n905), .Y(n307) );
  NAND2X0_HVT U210 ( .A1(adk_out0[125]), .A2(n879), .Y(n308) );
  NAND2X0_HVT U213 ( .A1(adk_in[125]), .A2(n854), .Y(n309) );
  NAND3X0_HVT U214 ( .A1(n307), .A2(n308), .A3(n309), .Y(n159) );
  INVX1_HVT U215 ( .A(n918), .Y(n905) );
  INVX1_HVT U216 ( .A(n310), .Y(n311) );
  NAND2X0_HVT U217 ( .A1(n995), .A2(n911), .Y(n312) );
  NAND2X0_HVT U218 ( .A1(adk_out0[56]), .A2(n885), .Y(n313) );
  NAND2X0_HVT U219 ( .A1(adk_in[56]), .A2(n849), .Y(n314) );
  NAND3X0_HVT U220 ( .A1(n312), .A2(n313), .A3(n314), .Y(n228) );
  INVX0_HVT U221 ( .A(n925), .Y(n432) );
  INVX0_HVT U222 ( .A(n980), .Y(n315) );
  INVX0_HVT U224 ( .A(n315), .Y(cipher_text[71]) );
  INVX0_HVT U226 ( .A(n948), .Y(n649) );
  INVX1_HVT U228 ( .A(n317), .Y(n318) );
  NAND2X0_HVT U229 ( .A1(n911), .A2(n993), .Y(n319) );
  NAND2X0_HVT U230 ( .A1(adk_out0[58]), .A2(n885), .Y(n320) );
  NAND2X0_HVT U232 ( .A1(adk_in[58]), .A2(n849), .Y(n321) );
  NAND3X0_HVT U234 ( .A1(n319), .A2(n320), .A3(n321), .Y(n226) );
  INVX0_HVT U235 ( .A(n1018), .Y(n774) );
  NAND2X0_HVT U237 ( .A1(n913), .A2(n1012), .Y(n322) );
  NAND2X0_HVT U238 ( .A1(adk_out0[39]), .A2(n887), .Y(n323) );
  NAND2X0_HVT U240 ( .A1(adk_in[39]), .A2(n362), .Y(n324) );
  NAND3X0_HVT U242 ( .A1(n322), .A2(n323), .A3(n324), .Y(n245) );
  INVX1_HVT U245 ( .A(n787), .Y(cipher_text[4]) );
  NAND2X0_HVT U246 ( .A1(n996), .A2(n911), .Y(n325) );
  NAND2X0_HVT U247 ( .A1(adk_out0[55]), .A2(n885), .Y(n326) );
  NAND2X0_HVT U250 ( .A1(adk_in[55]), .A2(n849), .Y(n327) );
  NAND3X0_HVT U252 ( .A1(n325), .A2(n326), .A3(n327), .Y(n229) );
  NAND2X0_HVT U253 ( .A1(n1038), .A2(n915), .Y(n328) );
  NAND2X0_HVT U254 ( .A1(adk_out0[13]), .A2(n889), .Y(n329) );
  NAND2X0_HVT U256 ( .A1(adk_in[13]), .A2(n847), .Y(n330) );
  NAND3X0_HVT U257 ( .A1(n328), .A2(n329), .A3(n330), .Y(n271) );
  INVX0_HVT U259 ( .A(n1042), .Y(n656) );
  INVX1_HVT U260 ( .A(n955), .Y(n520) );
  INVX0_HVT U261 ( .A(n1028), .Y(n767) );
  INVX0_HVT U262 ( .A(n934), .Y(n504) );
  NBUFFX2_HVT U264 ( .A(n1001), .Y(cipher_text[50]) );
  NBUFFX2_HVT U286 ( .A(n1026), .Y(cipher_text[25]) );
  INVX1_HVT U287 ( .A(n656), .Y(cipher_text[9]) );
  INVX0_HVT U288 ( .A(n930), .Y(n760) );
  INVX0_HVT U289 ( .A(n961), .Y(n743) );
  INVX1_HVT U290 ( .A(n760), .Y(cipher_text[121]) );
  INVX0_HVT U291 ( .A(n991), .Y(n822) );
  NAND2X0_HVT U292 ( .A1(n907), .A2(n946), .Y(n331) );
  NAND2X0_HVT U293 ( .A1(adk_out0[105]), .A2(n881), .Y(n332) );
  NAND2X0_HVT U294 ( .A1(adk_in[105]), .A2(n853), .Y(n333) );
  NAND3X0_HVT U295 ( .A1(n331), .A2(n332), .A3(n333), .Y(n179) );
  NAND2X0_HVT U296 ( .A1(n908), .A2(n962), .Y(n334) );
  NAND2X0_HVT U297 ( .A1(adk_out0[89]), .A2(n882), .Y(n335) );
  NAND2X0_HVT U298 ( .A1(adk_in[89]), .A2(n851), .Y(n336) );
  NAND3X0_HVT U299 ( .A1(n334), .A2(n335), .A3(n336), .Y(n195) );
  NAND2X0_HVT U300 ( .A1(n915), .A2(n1047), .Y(n337) );
  NAND2X0_HVT U301 ( .A1(adk_out0[4]), .A2(n889), .Y(n338) );
  NAND2X0_HVT U302 ( .A1(adk_in[4]), .A2(n846), .Y(n339) );
  NAND3X0_HVT U303 ( .A1(n337), .A2(n338), .A3(n339), .Y(n280) );
  NAND2X0_HVT U304 ( .A1(n945), .A2(n907), .Y(n340) );
  NAND2X0_HVT U305 ( .A1(adk_out0[106]), .A2(n881), .Y(n341) );
  NAND2X0_HVT U306 ( .A1(adk_in[106]), .A2(n853), .Y(n342) );
  NAND3X0_HVT U307 ( .A1(n340), .A2(n341), .A3(n342), .Y(n178) );
  NAND2X0_HVT U308 ( .A1(n955), .A2(n908), .Y(n343) );
  NAND2X0_HVT U309 ( .A1(adk_out0[96]), .A2(n882), .Y(n344) );
  NAND2X0_HVT U310 ( .A1(adk_in[96]), .A2(n852), .Y(n345) );
  NAND3X0_HVT U311 ( .A1(n343), .A2(n344), .A3(n345), .Y(n188) );
  INVX0_HVT U312 ( .A(n927), .Y(n833) );
  NAND2X0_HVT U313 ( .A1(n908), .A2(n952), .Y(n348) );
  NAND2X0_HVT U314 ( .A1(adk_out0[99]), .A2(n882), .Y(n349) );
  NAND2X0_HVT U315 ( .A1(adk_in[99]), .A2(n852), .Y(n350) );
  NAND3X0_HVT U316 ( .A1(n348), .A2(n349), .A3(n350), .Y(n185) );
  NBUFFX2_HVT U317 ( .A(n1031), .Y(cipher_text[20]) );
  INVX0_HVT U318 ( .A(n816), .Y(cipher_text[43]) );
  NAND2X0_HVT U319 ( .A1(n930), .A2(n906), .Y(n351) );
  NAND2X0_HVT U320 ( .A1(adk_out0[121]), .A2(n880), .Y(n352) );
  NAND2X0_HVT U321 ( .A1(adk_in[121]), .A2(n854), .Y(n353) );
  NAND3X0_HVT U322 ( .A1(n351), .A2(n352), .A3(n353), .Y(n163) );
  INVX1_HVT U323 ( .A(n743), .Y(cipher_text[90]) );
  INVX1_HVT U324 ( .A(n509), .Y(cipher_text[18]) );
  NAND2X0_HVT U325 ( .A1(n1018), .A2(n913), .Y(n354) );
  NAND2X0_HVT U326 ( .A1(adk_out0[33]), .A2(n887), .Y(n355) );
  NAND2X0_HVT U327 ( .A1(adk_in[33]), .A2(n848), .Y(n356) );
  NAND3X0_HVT U328 ( .A1(n354), .A2(n355), .A3(n356), .Y(n251) );
  INVX0_HVT U329 ( .A(n1015), .Y(n831) );
  INVX0_HVT U330 ( .A(n986), .Y(n753) );
  INVX0_HVT U331 ( .A(n1050), .Y(n721) );
  INVX1_HVT U332 ( .A(n628), .Y(n629) );
  NAND2X0_HVT U333 ( .A1(n1042), .A2(n915), .Y(n357) );
  NAND2X0_HVT U334 ( .A1(adk_out0[9]), .A2(n889), .Y(n358) );
  NAND2X0_HVT U335 ( .A1(adk_in[9]), .A2(n846), .Y(n359) );
  NAND3X0_HVT U336 ( .A1(n357), .A2(n358), .A3(n359), .Y(n275) );
  NBUFFX2_HVT U337 ( .A(n942), .Y(cipher_text[109]) );
  AO222X1_HVT U338 ( .A1(n360), .A2(n940), .A3(adk_out0[111]), .A4(n890), .A5(
        n361), .A6(n362), .Y(n173) );
  IBUFFX16_HVT U339 ( .A(n593), .Y(n360) );
  IBUFFX16_HVT U340 ( .A(n594), .Y(n361) );
  INVX0_HVT U341 ( .A(n940), .Y(n809) );
  INVX1_HVT U342 ( .A(n619), .Y(n620) );
  NAND2X0_HVT U343 ( .A1(n913), .A2(n1023), .Y(n363) );
  NAND2X0_HVT U344 ( .A1(adk_out0[28]), .A2(n887), .Y(n364) );
  NAND2X0_HVT U345 ( .A1(adk_in[28]), .A2(n848), .Y(n365) );
  NAND3X0_HVT U346 ( .A1(n363), .A2(n364), .A3(n365), .Y(n256) );
  NAND2X0_HVT U347 ( .A1(n910), .A2(n982), .Y(n366) );
  NAND2X0_HVT U348 ( .A1(adk_out0[69]), .A2(n884), .Y(n367) );
  NAND2X0_HVT U349 ( .A1(adk_in[69]), .A2(n850), .Y(n368) );
  NAND3X0_HVT U350 ( .A1(n366), .A2(n367), .A3(n368), .Y(n215) );
  INVX1_HVT U351 ( .A(n369), .Y(n370) );
  NAND2X0_HVT U352 ( .A1(n1002), .A2(n912), .Y(n371) );
  NAND2X0_HVT U353 ( .A1(adk_out0[49]), .A2(n886), .Y(n372) );
  NAND2X0_HVT U354 ( .A1(adk_in[49]), .A2(n362), .Y(n373) );
  NAND3X0_HVT U355 ( .A1(n371), .A2(n372), .A3(n373), .Y(n235) );
  NAND2X0_HVT U356 ( .A1(n942), .A2(n907), .Y(n374) );
  NAND2X0_HVT U357 ( .A1(adk_out0[109]), .A2(n881), .Y(n375) );
  NAND2X0_HVT U358 ( .A1(adk_in[109]), .A2(n853), .Y(n376) );
  NAND3X0_HVT U359 ( .A1(n374), .A2(n375), .A3(n376), .Y(n175) );
  INVX1_HVT U360 ( .A(n692), .Y(cipher_text[108]) );
  INVX0_HVT U361 ( .A(n943), .Y(n692) );
  NAND2X0_HVT U362 ( .A1(n1001), .A2(n912), .Y(n377) );
  NAND2X0_HVT U363 ( .A1(adk_out0[50]), .A2(n886), .Y(n378) );
  NAND2X0_HVT U364 ( .A1(adk_in[50]), .A2(n362), .Y(n379) );
  NAND3X0_HVT U365 ( .A1(n377), .A2(n378), .A3(n379), .Y(n234) );
  INVX1_HVT U366 ( .A(n704), .Y(cipher_text[41]) );
  INVX1_HVT U367 ( .A(n380), .Y(n381) );
  NAND2X0_HVT U368 ( .A1(n909), .A2(n973), .Y(n382) );
  NAND2X0_HVT U369 ( .A1(adk_out0[78]), .A2(n883), .Y(n383) );
  NAND2X0_HVT U370 ( .A1(adk_in[78]), .A2(n851), .Y(n384) );
  NAND3X0_HVT U371 ( .A1(n382), .A2(n383), .A3(n384), .Y(n206) );
  INVX1_HVT U372 ( .A(n918), .Y(n909) );
  NAND2X0_HVT U373 ( .A1(n306), .A2(n671), .Y(n213) );
  NAND2X0_HVT U374 ( .A1(n1033), .A2(n914), .Y(n385) );
  NAND2X0_HVT U375 ( .A1(adk_out0[18]), .A2(n888), .Y(n386) );
  NAND2X0_HVT U376 ( .A1(adk_in[18]), .A2(n847), .Y(n387) );
  NAND3X0_HVT U377 ( .A1(n385), .A2(n386), .A3(n387), .Y(n266) );
  INVX1_HVT U378 ( .A(n534), .Y(cipher_text[6]) );
  INVX1_HVT U379 ( .A(n1045), .Y(n534) );
  NAND2X0_HVT U380 ( .A1(n1045), .A2(n915), .Y(n388) );
  NAND2X0_HVT U381 ( .A1(adk_out0[6]), .A2(n889), .Y(n389) );
  NAND2X0_HVT U382 ( .A1(adk_in[6]), .A2(n846), .Y(n390) );
  NAND3X0_HVT U383 ( .A1(n388), .A2(n389), .A3(n390), .Y(n278) );
  INVX1_HVT U384 ( .A(n753), .Y(cipher_text[65]) );
  INVX0_HVT U385 ( .A(n1016), .Y(n791) );
  INVX0_HVT U386 ( .A(n989), .Y(n635) );
  INVX1_HVT U387 ( .A(n725), .Y(cipher_text[5]) );
  INVX1_HVT U388 ( .A(n635), .Y(cipher_text[62]) );
  INVX0_HVT U389 ( .A(n1005), .Y(n584) );
  INVX1_HVT U390 ( .A(n1046), .Y(n725) );
  NAND2X0_HVT U391 ( .A1(n961), .A2(n908), .Y(n391) );
  NAND2X0_HVT U392 ( .A1(adk_out0[90]), .A2(n882), .Y(n392) );
  NAND2X0_HVT U393 ( .A1(adk_in[90]), .A2(n852), .Y(n393) );
  NAND3X0_HVT U394 ( .A1(n391), .A2(n392), .A3(n393), .Y(n194) );
  INVX0_HVT U395 ( .A(n968), .Y(n734) );
  NAND2X0_HVT U396 ( .A1(n986), .A2(n910), .Y(n394) );
  NAND2X0_HVT U397 ( .A1(adk_out0[65]), .A2(n884), .Y(n395) );
  NAND2X0_HVT U398 ( .A1(adk_in[65]), .A2(n850), .Y(n396) );
  NAND3X0_HVT U399 ( .A1(n394), .A2(n395), .A3(n396), .Y(n219) );
  INVX1_HVT U400 ( .A(n721), .Y(cipher_text[1]) );
  NAND2X0_HVT U401 ( .A1(n1043), .A2(n915), .Y(n397) );
  NAND2X0_HVT U402 ( .A1(adk_out0[8]), .A2(n889), .Y(n398) );
  NAND2X0_HVT U403 ( .A1(adk_in[8]), .A2(n846), .Y(n399) );
  NAND3X0_HVT U404 ( .A1(n397), .A2(n398), .A3(n399), .Y(n276) );
  NAND2X0_HVT U405 ( .A1(n912), .A2(n1006), .Y(n400) );
  NAND2X0_HVT U406 ( .A1(adk_out0[45]), .A2(n886), .Y(n401) );
  NAND2X0_HVT U407 ( .A1(adk_in[45]), .A2(n362), .Y(n402) );
  NAND3X0_HVT U408 ( .A1(n400), .A2(n401), .A3(n402), .Y(n239) );
  INVX0_HVT U409 ( .A(n976), .Y(n814) );
  NAND2X0_HVT U410 ( .A1(n912), .A2(n1010), .Y(n403) );
  NAND2X0_HVT U411 ( .A1(adk_out0[41]), .A2(n886), .Y(n404) );
  NAND2X0_HVT U412 ( .A1(adk_in[41]), .A2(n362), .Y(n405) );
  NAND3X0_HVT U413 ( .A1(n403), .A2(n404), .A3(n405), .Y(n243) );
  NAND2X0_HVT U414 ( .A1(n1046), .A2(n915), .Y(n406) );
  NAND2X0_HVT U415 ( .A1(adk_out0[5]), .A2(n889), .Y(n407) );
  NAND2X0_HVT U416 ( .A1(adk_in[5]), .A2(n846), .Y(n408) );
  NAND3X0_HVT U417 ( .A1(n406), .A2(n407), .A3(n408), .Y(n279) );
  INVX1_HVT U418 ( .A(n409), .Y(n410) );
  INVX0_HVT U419 ( .A(n990), .Y(n844) );
  NAND2X0_HVT U420 ( .A1(n989), .A2(n911), .Y(n411) );
  NAND2X0_HVT U421 ( .A1(adk_out0[62]), .A2(n885), .Y(n412) );
  NAND2X0_HVT U422 ( .A1(adk_in[62]), .A2(n849), .Y(n413) );
  NAND3X0_HVT U423 ( .A1(n411), .A2(n412), .A3(n413), .Y(n222) );
  NAND2X0_HVT U424 ( .A1(n1003), .A2(n912), .Y(n414) );
  NAND2X0_HVT U425 ( .A1(adk_out0[48]), .A2(n886), .Y(n415) );
  NAND2X0_HVT U426 ( .A1(adk_in[48]), .A2(n362), .Y(n416) );
  NAND3X0_HVT U427 ( .A1(n414), .A2(n415), .A3(n416), .Y(n236) );
  INVX0_HVT U428 ( .A(n972), .Y(n684) );
  NAND2X0_HVT U429 ( .A1(n943), .A2(n907), .Y(n417) );
  NAND2X0_HVT U430 ( .A1(adk_out0[108]), .A2(n881), .Y(n418) );
  NAND2X0_HVT U431 ( .A1(adk_in[108]), .A2(n853), .Y(n419) );
  NAND3X0_HVT U432 ( .A1(n417), .A2(n418), .A3(n419), .Y(n176) );
  INVX1_HVT U433 ( .A(n918), .Y(n907) );
  NAND2X0_HVT U434 ( .A1(n1021), .A2(n913), .Y(n420) );
  NAND2X0_HVT U435 ( .A1(adk_out0[30]), .A2(n887), .Y(n421) );
  NAND2X0_HVT U436 ( .A1(adk_in[30]), .A2(n848), .Y(n422) );
  NAND3X0_HVT U437 ( .A1(n420), .A2(n421), .A3(n422), .Y(n254) );
  NAND2X0_HVT U438 ( .A1(n914), .A2(n1031), .Y(n423) );
  NAND2X0_HVT U439 ( .A1(adk_out0[20]), .A2(n888), .Y(n424) );
  NAND2X0_HVT U440 ( .A1(adk_in[20]), .A2(n847), .Y(n425) );
  NAND3X0_HVT U441 ( .A1(n423), .A2(n424), .A3(n425), .Y(n264) );
  NAND2X0_HVT U442 ( .A1(n908), .A2(n954), .Y(n426) );
  NAND2X0_HVT U443 ( .A1(adk_out0[97]), .A2(n882), .Y(n427) );
  NAND2X0_HVT U444 ( .A1(adk_in[97]), .A2(n852), .Y(n428) );
  NAND3X0_HVT U445 ( .A1(n426), .A2(n427), .A3(n428), .Y(n187) );
  NBUFFX2_HVT U446 ( .A(n1039), .Y(cipher_text[12]) );
  NAND2X0_HVT U447 ( .A1(n925), .A2(n905), .Y(n429) );
  NAND2X0_HVT U448 ( .A1(adk_out0[126]), .A2(n879), .Y(n430) );
  NAND2X0_HVT U449 ( .A1(adk_in[126]), .A2(n854), .Y(n431) );
  NAND3X0_HVT U450 ( .A1(n429), .A2(n430), .A3(n431), .Y(n158) );
  INVX1_HVT U451 ( .A(n432), .Y(cipher_text[126]) );
  INVX1_HVT U452 ( .A(n765), .Y(cipher_text[66]) );
  INVX1_HVT U453 ( .A(n436), .Y(n437) );
  NAND2X0_HVT U454 ( .A1(n984), .A2(n15), .Y(n438) );
  NAND2X0_HVT U455 ( .A1(adk_out0[67]), .A2(n16), .Y(n439) );
  NAND2X0_HVT U456 ( .A1(adk_in[67]), .A2(n17), .Y(n440) );
  NAND3X0_HVT U457 ( .A1(n438), .A2(n439), .A3(n440), .Y(n217) );
  NBUFFX2_HVT U458 ( .A(n938), .Y(cipher_text[113]) );
  NAND2X0_HVT U459 ( .A1(n990), .A2(n911), .Y(n443) );
  NAND2X0_HVT U460 ( .A1(adk_out0[61]), .A2(n885), .Y(n444) );
  NAND2X0_HVT U461 ( .A1(adk_in[61]), .A2(n849), .Y(n445) );
  NAND3X0_HVT U462 ( .A1(n443), .A2(n444), .A3(n445), .Y(n223) );
  NAND2X0_HVT U463 ( .A1(n987), .A2(n910), .Y(n446) );
  NAND2X0_HVT U464 ( .A1(adk_out0[64]), .A2(n884), .Y(n447) );
  NAND2X0_HVT U465 ( .A1(adk_in[64]), .A2(n850), .Y(n448) );
  NAND3X0_HVT U466 ( .A1(n446), .A2(n447), .A3(n448), .Y(n220) );
  NAND2X0_HVT U467 ( .A1(n974), .A2(n909), .Y(n449) );
  NAND2X0_HVT U468 ( .A1(adk_out0[77]), .A2(n883), .Y(n450) );
  NAND2X0_HVT U469 ( .A1(adk_in[77]), .A2(n851), .Y(n451) );
  NAND3X0_HVT U470 ( .A1(n449), .A2(n450), .A3(n451), .Y(n207) );
  INVX0_HVT U471 ( .A(n974), .Y(n452) );
  INVX0_HVT U472 ( .A(n452), .Y(cipher_text[77]) );
  NAND2X0_HVT U473 ( .A1(n914), .A2(n1026), .Y(n454) );
  NAND2X0_HVT U474 ( .A1(adk_out0[25]), .A2(n888), .Y(n455) );
  NAND2X0_HVT U475 ( .A1(adk_in[25]), .A2(n848), .Y(n456) );
  NAND3X0_HVT U476 ( .A1(n454), .A2(n455), .A3(n456), .Y(n259) );
  INVX0_HVT U477 ( .A(n957), .Y(n658) );
  NAND2X0_HVT U478 ( .A1(n971), .A2(n909), .Y(n457) );
  NAND2X0_HVT U479 ( .A1(adk_out0[80]), .A2(n883), .Y(n458) );
  NAND2X0_HVT U480 ( .A1(adk_in[80]), .A2(n851), .Y(n459) );
  NAND3X0_HVT U481 ( .A1(n457), .A2(n458), .A3(n459), .Y(n204) );
  INVX1_HVT U482 ( .A(n985), .Y(n765) );
  NAND2X0_HVT U483 ( .A1(n914), .A2(n1032), .Y(n460) );
  NAND2X0_HVT U484 ( .A1(adk_out0[19]), .A2(n888), .Y(n461) );
  NAND2X0_HVT U485 ( .A1(adk_in[19]), .A2(n847), .Y(n462) );
  NAND3X0_HVT U486 ( .A1(n460), .A2(n461), .A3(n462), .Y(n265) );
  NAND2X0_HVT U487 ( .A1(n1004), .A2(n912), .Y(n463) );
  NAND2X0_HVT U488 ( .A1(adk_out0[47]), .A2(n886), .Y(n464) );
  NAND2X0_HVT U489 ( .A1(adk_in[47]), .A2(n362), .Y(n465) );
  NAND3X0_HVT U490 ( .A1(n463), .A2(n464), .A3(n465), .Y(n237) );
  INVX1_HVT U491 ( .A(n758), .Y(cipher_text[68]) );
  INVX0_HVT U492 ( .A(n776), .Y(cipher_text[57]) );
  NAND2X0_HVT U493 ( .A1(n916), .A2(n1050), .Y(n468) );
  NAND2X0_HVT U494 ( .A1(adk_out0[1]), .A2(n890), .Y(n469) );
  NAND2X0_HVT U495 ( .A1(adk_in[1]), .A2(n846), .Y(n470) );
  NAND3X0_HVT U496 ( .A1(n468), .A2(n469), .A3(n470), .Y(n283) );
  NAND2X0_HVT U497 ( .A1(n915), .A2(n1039), .Y(n471) );
  NAND2X0_HVT U498 ( .A1(adk_out0[12]), .A2(n889), .Y(n472) );
  NAND2X0_HVT U499 ( .A1(adk_in[12]), .A2(n847), .Y(n473) );
  NAND3X0_HVT U500 ( .A1(n471), .A2(n472), .A3(n473), .Y(n272) );
  NAND2X0_HVT U501 ( .A1(n947), .A2(n907), .Y(n474) );
  NAND2X0_HVT U502 ( .A1(adk_out0[104]), .A2(n881), .Y(n475) );
  NAND2X0_HVT U503 ( .A1(adk_in[104]), .A2(n853), .Y(n476) );
  NAND3X0_HVT U504 ( .A1(n474), .A2(n475), .A3(n476), .Y(n180) );
  INVX1_HVT U505 ( .A(n947), .Y(n477) );
  INVX1_HVT U506 ( .A(n477), .Y(cipher_text[104]) );
  INVX0_HVT U507 ( .A(n949), .Y(n479) );
  INVX0_HVT U508 ( .A(n479), .Y(cipher_text[102]) );
  NAND2X0_HVT U509 ( .A1(n908), .A2(n960), .Y(n481) );
  NAND2X0_HVT U510 ( .A1(adk_out0[91]), .A2(n882), .Y(n482) );
  NAND2X0_HVT U511 ( .A1(adk_in[91]), .A2(n852), .Y(n483) );
  NAND3X0_HVT U512 ( .A1(n481), .A2(n482), .A3(n483), .Y(n193) );
  INVX1_HVT U513 ( .A(n772), .Y(cipher_text[127]) );
  INVX1_HVT U514 ( .A(n924), .Y(n772) );
  INVX0_HVT U515 ( .A(n941), .Y(n486) );
  INVX0_HVT U516 ( .A(n486), .Y(cipher_text[110]) );
  NAND2X0_HVT U517 ( .A1(n905), .A2(n924), .Y(n490) );
  NAND2X0_HVT U518 ( .A1(adk_out0[127]), .A2(n879), .Y(n491) );
  NAND2X0_HVT U519 ( .A1(adk_in[127]), .A2(n854), .Y(n492) );
  NAND3X0_HVT U520 ( .A1(n490), .A2(n491), .A3(n492), .Y(n157) );
  NAND2X0_HVT U521 ( .A1(n910), .A2(n985), .Y(n493) );
  NAND2X0_HVT U522 ( .A1(adk_out0[66]), .A2(n884), .Y(n494) );
  NAND2X0_HVT U523 ( .A1(adk_in[66]), .A2(n850), .Y(n495) );
  NAND3X0_HVT U524 ( .A1(n493), .A2(n494), .A3(n495), .Y(n218) );
  INVX1_HVT U525 ( .A(n918), .Y(n910) );
  INVX0_HVT U526 ( .A(n994), .Y(n776) );
  NAND2X0_HVT U527 ( .A1(n906), .A2(n938), .Y(n498) );
  NAND2X0_HVT U528 ( .A1(adk_out0[113]), .A2(n880), .Y(n499) );
  NAND2X0_HVT U529 ( .A1(adk_in[113]), .A2(n853), .Y(n500) );
  NAND3X0_HVT U530 ( .A1(n498), .A2(n499), .A3(n500), .Y(n171) );
  INVX1_HVT U531 ( .A(n918), .Y(n906) );
  NAND2X0_HVT U532 ( .A1(n934), .A2(n906), .Y(n501) );
  NAND2X0_HVT U533 ( .A1(adk_out0[117]), .A2(n880), .Y(n502) );
  NAND2X0_HVT U534 ( .A1(adk_in[117]), .A2(n854), .Y(n503) );
  NAND3X0_HVT U535 ( .A1(n501), .A2(n502), .A3(n503), .Y(n167) );
  INVX1_HVT U536 ( .A(n504), .Y(cipher_text[117]) );
  NAND2X0_HVT U537 ( .A1(n913), .A2(n1020), .Y(n506) );
  NAND2X0_HVT U538 ( .A1(adk_out0[31]), .A2(n887), .Y(n507) );
  NAND2X0_HVT U539 ( .A1(adk_in[31]), .A2(n848), .Y(n508) );
  NAND3X0_HVT U540 ( .A1(n506), .A2(n507), .A3(n508), .Y(n253) );
  INVX1_HVT U541 ( .A(n917), .Y(n913) );
  INVX1_HVT U542 ( .A(n511), .Y(n512) );
  INVX0_HVT U543 ( .A(n1024), .Y(n785) );
  INVX1_HVT U544 ( .A(n513), .Y(n514) );
  NBUFFX2_HVT U545 ( .A(n1025), .Y(cipher_text[26]) );
  INVX0_HVT U546 ( .A(n933), .Y(n516) );
  INVX0_HVT U547 ( .A(n516), .Y(cipher_text[118]) );
  INVX1_HVT U548 ( .A(n734), .Y(cipher_text[83]) );
  INVX0_HVT U549 ( .A(n926), .Y(n518) );
  INVX0_HVT U550 ( .A(n518), .Y(cipher_text[125]) );
  INVX0_HVT U551 ( .A(n520), .Y(cipher_text[96]) );
  NBUFFX2_HVT U552 ( .A(n978), .Y(cipher_text[73]) );
  INVX0_HVT U553 ( .A(n965), .Y(n522) );
  INVX0_HVT U554 ( .A(n522), .Y(cipher_text[86]) );
  NAND2X0_HVT U555 ( .A1(n909), .A2(n968), .Y(n524) );
  NAND2X0_HVT U556 ( .A1(adk_out0[83]), .A2(n883), .Y(n525) );
  NAND2X0_HVT U557 ( .A1(adk_in[83]), .A2(n851), .Y(n526) );
  NAND3X0_HVT U558 ( .A1(n524), .A2(n525), .A3(n526), .Y(n201) );
  NAND2X0_HVT U559 ( .A1(n910), .A2(n977), .Y(n527) );
  NAND2X0_HVT U560 ( .A1(adk_out0[74]), .A2(n884), .Y(n528) );
  NAND2X0_HVT U561 ( .A1(adk_in[74]), .A2(n850), .Y(n529) );
  NAND3X0_HVT U562 ( .A1(n527), .A2(n528), .A3(n529), .Y(n210) );
  INVX1_HVT U563 ( .A(n977), .Y(n530) );
  INVX1_HVT U564 ( .A(n530), .Y(cipher_text[74]) );
  INVX0_HVT U565 ( .A(n999), .Y(n829) );
  INVX1_HVT U566 ( .A(n822), .Y(cipher_text[60]) );
  INVX0_HVT U567 ( .A(n1022), .Y(n532) );
  INVX0_HVT U568 ( .A(n532), .Y(cipher_text[29]) );
  INVX1_HVT U569 ( .A(n837), .Y(cipher_text[84]) );
  INVX0_HVT U570 ( .A(n1006), .Y(n536) );
  INVX0_HVT U571 ( .A(n536), .Y(cipher_text[45]) );
  INVX0_HVT U572 ( .A(n1037), .Y(n538) );
  INVX0_HVT U573 ( .A(n538), .Y(cipher_text[14]) );
  NAND2X0_HVT U574 ( .A1(n911), .A2(n302), .Y(n540) );
  NAND2X0_HVT U575 ( .A1(adk_out0[52]), .A2(n885), .Y(n541) );
  NAND2X0_HVT U576 ( .A1(adk_in[52]), .A2(n849), .Y(n542) );
  NAND3X0_HVT U577 ( .A1(n540), .A2(n541), .A3(n542), .Y(n232) );
  NAND2X0_HVT U578 ( .A1(n910), .A2(n978), .Y(n543) );
  NAND2X0_HVT U579 ( .A1(adk_out0[73]), .A2(n884), .Y(n544) );
  NAND2X0_HVT U580 ( .A1(adk_in[73]), .A2(n850), .Y(n545) );
  NAND3X0_HVT U581 ( .A1(n543), .A2(n544), .A3(n545), .Y(n211) );
  INVX0_HVT U582 ( .A(n1030), .Y(n546) );
  INVX0_HVT U583 ( .A(n546), .Y(cipher_text[21]) );
  INVX0_HVT U584 ( .A(n997), .Y(n548) );
  INVX0_HVT U585 ( .A(n548), .Y(cipher_text[54]) );
  INVX0_HVT U586 ( .A(n1011), .Y(n550) );
  INVX0_HVT U587 ( .A(n550), .Y(cipher_text[40]) );
  NBUFFX2_HVT U588 ( .A(n979), .Y(cipher_text[72]) );
  NAND2X0_HVT U589 ( .A1(n991), .A2(n911), .Y(n553) );
  NAND2X0_HVT U590 ( .A1(adk_out0[60]), .A2(n885), .Y(n554) );
  NAND2X0_HVT U591 ( .A1(adk_in[60]), .A2(n849), .Y(n555) );
  NAND3X0_HVT U592 ( .A1(n553), .A2(n554), .A3(n555), .Y(n224) );
  INVX1_HVT U593 ( .A(n917), .Y(n911) );
  INVX1_HVT U594 ( .A(n767), .Y(cipher_text[23]) );
  INVX0_HVT U595 ( .A(n963), .Y(n556) );
  INVX0_HVT U596 ( .A(n556), .Y(cipher_text[88]) );
  INVX1_HVT U597 ( .A(n558), .Y(n559) );
  NAND2X0_HVT U598 ( .A1(n908), .A2(n957), .Y(n560) );
  NAND2X0_HVT U599 ( .A1(adk_out0[94]), .A2(n882), .Y(n561) );
  NAND2X0_HVT U600 ( .A1(adk_in[94]), .A2(n852), .Y(n562) );
  NAND3X0_HVT U601 ( .A1(n560), .A2(n561), .A3(n562), .Y(n190) );
  NAND2X0_HVT U602 ( .A1(n1028), .A2(n914), .Y(n563) );
  NAND2X0_HVT U603 ( .A1(adk_out0[23]), .A2(n888), .Y(n564) );
  NAND2X0_HVT U604 ( .A1(adk_in[23]), .A2(n847), .Y(n565) );
  NAND3X0_HVT U605 ( .A1(n563), .A2(n564), .A3(n565), .Y(n261) );
  INVX1_HVT U606 ( .A(n917), .Y(n914) );
  INVX0_HVT U607 ( .A(n827), .Y(cipher_text[11]) );
  NBUFFX2_HVT U608 ( .A(n1044), .Y(cipher_text[7]) );
  NAND2X0_HVT U609 ( .A1(n906), .A2(n935), .Y(n567) );
  NAND2X0_HVT U610 ( .A1(adk_out0[116]), .A2(n880), .Y(n568) );
  NAND2X0_HVT U611 ( .A1(adk_in[116]), .A2(n854), .Y(n569) );
  NAND3X0_HVT U612 ( .A1(n567), .A2(n568), .A3(n569), .Y(n168) );
  NAND2X0_HVT U613 ( .A1(n1007), .A2(n912), .Y(n570) );
  NAND2X0_HVT U614 ( .A1(adk_out0[44]), .A2(n886), .Y(n571) );
  NAND2X0_HVT U615 ( .A1(adk_in[44]), .A2(n362), .Y(n572) );
  NAND3X0_HVT U616 ( .A1(n570), .A2(n571), .A3(n572), .Y(n240) );
  INVX1_HVT U617 ( .A(n917), .Y(n912) );
  NBUFFX2_HVT U618 ( .A(n1029), .Y(cipher_text[22]) );
  INVX1_HVT U619 ( .A(n1021), .Y(n574) );
  INVX1_HVT U620 ( .A(n574), .Y(cipher_text[30]) );
  NAND2X0_HVT U621 ( .A1(n988), .A2(n911), .Y(n576) );
  NAND2X0_HVT U622 ( .A1(adk_out0[63]), .A2(n885), .Y(n577) );
  NAND2X0_HVT U623 ( .A1(adk_in[63]), .A2(n849), .Y(n578) );
  NAND3X0_HVT U624 ( .A1(n576), .A2(n577), .A3(n578), .Y(n221) );
  INVX1_HVT U625 ( .A(n988), .Y(n579) );
  INVX1_HVT U626 ( .A(n579), .Y(cipher_text[63]) );
  NAND2X0_HVT U627 ( .A1(n1005), .A2(n912), .Y(n581) );
  NAND2X0_HVT U628 ( .A1(adk_out0[46]), .A2(n886), .Y(n582) );
  NAND2X0_HVT U629 ( .A1(adk_in[46]), .A2(n362), .Y(n583) );
  NAND3X0_HVT U630 ( .A1(n581), .A2(n582), .A3(n583), .Y(n238) );
  INVX1_HVT U631 ( .A(n584), .Y(cipher_text[46]) );
  INVX0_HVT U632 ( .A(n915), .Y(n600) );
  INVX1_HVT U633 ( .A(n644), .Y(n645) );
  INVX0_HVT U634 ( .A(n907), .Y(n593) );
  INVX1_HVT U635 ( .A(adk_out0[15]), .Y(n601) );
  INVX0_HVT U636 ( .A(n847), .Y(n603) );
  INVX0_HVT U637 ( .A(n889), .Y(n602) );
  AND2X1_HVT U638 ( .A1(n803), .A2(n802), .Y(n586) );
  INVX1_HVT U639 ( .A(n587), .Y(n588) );
  NBUFFX2_HVT U640 ( .A(n945), .Y(cipher_text[106]) );
  NBUFFX2_HVT U641 ( .A(n1041), .Y(cipher_text[10]) );
  NBUFFX2_HVT U642 ( .A(n951), .Y(cipher_text[100]) );
  NBUFFX2_HVT U643 ( .A(n995), .Y(cipher_text[56]) );
  NBUFFX2_HVT U644 ( .A(n1019), .Y(cipher_text[32]) );
  INVX1_HVT U645 ( .A(n1036), .Y(n669) );
  NBUFFX2_HVT U646 ( .A(n993), .Y(cipher_text[58]) );
  NBUFFX2_HVT U647 ( .A(n981), .Y(cipher_text[70]) );
  NBUFFX2_HVT U648 ( .A(n962), .Y(cipher_text[89]) );
  IBUFFX16_HVT U649 ( .A(n905), .Y(n616) );
  NBUFFX2_HVT U650 ( .A(n1012), .Y(cipher_text[39]) );
  NBUFFX2_HVT U651 ( .A(n1035), .Y(cipher_text[16]) );
  INVX0_HVT U652 ( .A(n998), .Y(n622) );
  INVX0_HVT U653 ( .A(n622), .Y(cipher_text[53]) );
  NAND2X0_HVT U654 ( .A1(n911), .A2(n994), .Y(n632) );
  NAND2X0_HVT U655 ( .A1(adk_out0[57]), .A2(n885), .Y(n633) );
  NAND2X0_HVT U656 ( .A1(adk_in[57]), .A2(n849), .Y(n634) );
  NAND3X0_HVT U657 ( .A1(n632), .A2(n633), .A3(n634), .Y(n227) );
  NAND2X0_HVT U658 ( .A1(n967), .A2(n909), .Y(n637) );
  NAND2X0_HVT U659 ( .A1(adk_out0[84]), .A2(n883), .Y(n638) );
  NAND2X0_HVT U660 ( .A1(adk_in[84]), .A2(n851), .Y(n639) );
  NAND3X0_HVT U661 ( .A1(n637), .A2(n638), .A3(n639), .Y(n200) );
  INVX0_HVT U662 ( .A(n936), .Y(n640) );
  INVX0_HVT U663 ( .A(n640), .Y(cipher_text[115]) );
  INVX0_HVT U664 ( .A(n958), .Y(n642) );
  INVX0_HVT U665 ( .A(n642), .Y(cipher_text[93]) );
  INVX1_HVT U666 ( .A(n950), .Y(n709) );
  NAND2X0_HVT U667 ( .A1(n948), .A2(n907), .Y(n646) );
  NAND2X0_HVT U668 ( .A1(adk_out0[103]), .A2(n881), .Y(n647) );
  NAND2X0_HVT U669 ( .A1(adk_in[103]), .A2(n853), .Y(n648) );
  NAND3X0_HVT U670 ( .A1(n646), .A2(n647), .A3(n648), .Y(n181) );
  INVX1_HVT U671 ( .A(n649), .Y(cipher_text[103]) );
  INVX0_HVT U672 ( .A(n953), .Y(n651) );
  INVX0_HVT U673 ( .A(n651), .Y(cipher_text[98]) );
  NAND2X0_HVT U674 ( .A1(n950), .A2(n907), .Y(n653) );
  NAND2X0_HVT U675 ( .A1(adk_out0[101]), .A2(n881), .Y(n654) );
  NAND2X0_HVT U676 ( .A1(adk_in[101]), .A2(n852), .Y(n655) );
  NAND3X0_HVT U677 ( .A1(n653), .A2(n654), .A3(n655), .Y(n183) );
  INVX1_HVT U678 ( .A(n658), .Y(cipher_text[94]) );
  INVX0_HVT U679 ( .A(n1040), .Y(n827) );
  NAND2X0_HVT U680 ( .A1(n956), .A2(n908), .Y(n660) );
  NAND2X0_HVT U681 ( .A1(adk_out0[95]), .A2(n882), .Y(n661) );
  NAND2X0_HVT U682 ( .A1(adk_in[95]), .A2(n852), .Y(n662) );
  NAND3X0_HVT U683 ( .A1(n660), .A2(n661), .A3(n662), .Y(n189) );
  INVX0_HVT U684 ( .A(n956), .Y(n663) );
  INVX1_HVT U685 ( .A(n918), .Y(n908) );
  INVX0_HVT U686 ( .A(n939), .Y(n665) );
  INVX0_HVT U687 ( .A(n665), .Y(cipher_text[112]) );
  INVX0_HVT U688 ( .A(n669), .Y(cipher_text[15]) );
  NAND2X0_HVT U689 ( .A1(n980), .A2(n910), .Y(n671) );
  NAND2X0_HVT U690 ( .A1(adk_out0[71]), .A2(n884), .Y(n672) );
  NAND2X0_HVT U691 ( .A1(adk_in[71]), .A2(n850), .Y(n673) );
  INVX0_HVT U692 ( .A(n954), .Y(n676) );
  INVX0_HVT U693 ( .A(n676), .Y(cipher_text[97]) );
  NBUFFX2_HVT U694 ( .A(n969), .Y(cipher_text[82]) );
  NAND2X0_HVT U695 ( .A1(n586), .A2(n801), .Y(n192) );
  INVX0_HVT U696 ( .A(n959), .Y(n679) );
  INVX0_HVT U697 ( .A(n679), .Y(cipher_text[92]) );
  NAND2X0_HVT U698 ( .A1(n972), .A2(n909), .Y(n681) );
  NAND2X0_HVT U699 ( .A1(adk_out0[79]), .A2(n883), .Y(n682) );
  NAND2X0_HVT U700 ( .A1(adk_in[79]), .A2(n851), .Y(n683) );
  NAND3X0_HVT U701 ( .A1(n681), .A2(n682), .A3(n683), .Y(n205) );
  INVX1_HVT U702 ( .A(n684), .Y(cipher_text[79]) );
  INVX0_HVT U703 ( .A(n983), .Y(n758) );
  INVX1_HVT U704 ( .A(n818), .Y(cipher_text[59]) );
  NAND2X0_HVT U705 ( .A1(n992), .A2(n911), .Y(n686) );
  NAND2X0_HVT U706 ( .A1(adk_out0[59]), .A2(n885), .Y(n687) );
  NAND2X0_HVT U707 ( .A1(adk_in[59]), .A2(n849), .Y(n688) );
  NAND3X0_HVT U708 ( .A1(n686), .A2(n687), .A3(n688), .Y(n225) );
  NAND2X0_HVT U709 ( .A1(n913), .A2(n1014), .Y(n694) );
  NAND2X0_HVT U710 ( .A1(adk_out0[37]), .A2(n887), .Y(n695) );
  NAND2X0_HVT U711 ( .A1(adk_in[37]), .A2(n848), .Y(n696) );
  NAND3X0_HVT U712 ( .A1(n694), .A2(n695), .A3(n696), .Y(n247) );
  INVX1_HVT U713 ( .A(n1014), .Y(n697) );
  INVX1_HVT U714 ( .A(n697), .Y(cipher_text[37]) );
  INVX0_HVT U715 ( .A(n1013), .Y(n699) );
  INVX0_HVT U716 ( .A(n699), .Y(cipher_text[38]) );
  INVX1_HVT U717 ( .A(n701), .Y(n702) );
  INVX0_HVT U718 ( .A(n1010), .Y(n704) );
  INVX1_HVT U719 ( .A(n831), .Y(cipher_text[36]) );
  NAND2X0_HVT U720 ( .A1(n913), .A2(n1015), .Y(n706) );
  NAND2X0_HVT U721 ( .A1(adk_out0[36]), .A2(n887), .Y(n707) );
  NAND2X0_HVT U722 ( .A1(adk_in[36]), .A2(n848), .Y(n708) );
  NAND3X0_HVT U723 ( .A1(n706), .A2(n707), .A3(n708), .Y(n248) );
  INVX1_HVT U724 ( .A(n709), .Y(cipher_text[101]) );
  NAND2X0_HVT U725 ( .A1(n915), .A2(n1040), .Y(n711) );
  NAND2X0_HVT U726 ( .A1(adk_out0[11]), .A2(n889), .Y(n712) );
  NAND2X0_HVT U727 ( .A1(adk_in[11]), .A2(n846), .Y(n713) );
  NAND3X0_HVT U728 ( .A1(n711), .A2(n712), .A3(n713), .Y(n273) );
  NAND2X0_HVT U729 ( .A1(n929), .A2(n906), .Y(n714) );
  NAND2X0_HVT U730 ( .A1(adk_out0[122]), .A2(n880), .Y(n715) );
  NAND2X0_HVT U731 ( .A1(adk_in[122]), .A2(n854), .Y(n716) );
  NAND3X0_HVT U732 ( .A1(n714), .A2(n715), .A3(n716), .Y(n162) );
  INVX1_HVT U733 ( .A(n929), .Y(n717) );
  INVX1_HVT U734 ( .A(n717), .Y(cipher_text[122]) );
  INVX0_HVT U735 ( .A(n1051), .Y(n719) );
  INVX0_HVT U736 ( .A(n719), .Y(cipher_text[0]) );
  INVX0_HVT U737 ( .A(n1020), .Y(n723) );
  INVX0_HVT U738 ( .A(n723), .Y(cipher_text[31]) );
  NBUFFX2_HVT U739 ( .A(n1000), .Y(cipher_text[51]) );
  INVX0_HVT U740 ( .A(n932), .Y(n728) );
  INVX0_HVT U741 ( .A(n728), .Y(cipher_text[119]) );
  INVX0_HVT U742 ( .A(n952), .Y(n730) );
  INVX0_HVT U743 ( .A(n730), .Y(cipher_text[99]) );
  INVX0_HVT U744 ( .A(n1034), .Y(n732) );
  INVX0_HVT U745 ( .A(n732), .Y(cipher_text[17]) );
  INVX1_HVT U746 ( .A(n791), .Y(cipher_text[35]) );
  NAND2X0_HVT U747 ( .A1(n909), .A2(n975), .Y(n736) );
  NAND2X0_HVT U748 ( .A1(adk_out0[76]), .A2(n883), .Y(n737) );
  NAND2X0_HVT U749 ( .A1(adk_in[76]), .A2(n850), .Y(n738) );
  NAND3X0_HVT U750 ( .A1(n736), .A2(n737), .A3(n738), .Y(n208) );
  INVX1_HVT U751 ( .A(n739), .Y(cipher_text[76]) );
  INVX1_HVT U752 ( .A(n741), .Y(n742) );
  INVX0_HVT U753 ( .A(n931), .Y(n745) );
  INVX0_HVT U754 ( .A(n745), .Y(cipher_text[120]) );
  NAND2X0_HVT U755 ( .A1(n913), .A2(n1016), .Y(n747) );
  NAND2X0_HVT U756 ( .A1(adk_out0[35]), .A2(n887), .Y(n748) );
  NAND2X0_HVT U757 ( .A1(adk_in[35]), .A2(n848), .Y(n749) );
  NAND3X0_HVT U758 ( .A1(n747), .A2(n748), .A3(n749), .Y(n249) );
  NAND2X0_HVT U759 ( .A1(n1008), .A2(n912), .Y(n750) );
  NAND2X0_HVT U760 ( .A1(adk_out0[43]), .A2(n886), .Y(n751) );
  NAND2X0_HVT U761 ( .A1(adk_in[43]), .A2(n864), .Y(n752) );
  NAND3X0_HVT U762 ( .A1(n750), .A2(n751), .A3(n752), .Y(n241) );
  NAND2X0_HVT U763 ( .A1(n983), .A2(n910), .Y(n755) );
  NAND2X0_HVT U764 ( .A1(adk_out0[68]), .A2(n884), .Y(n756) );
  NAND2X0_HVT U765 ( .A1(adk_in[68]), .A2(n850), .Y(n757) );
  NAND3X0_HVT U766 ( .A1(n755), .A2(n756), .A3(n757), .Y(n216) );
  INVX1_HVT U767 ( .A(n814), .Y(cipher_text[75]) );
  NAND2X0_HVT U768 ( .A1(n912), .A2(n1000), .Y(n762) );
  NAND2X0_HVT U769 ( .A1(adk_out0[51]), .A2(n886), .Y(n763) );
  NAND2X0_HVT U770 ( .A1(adk_in[51]), .A2(n849), .Y(n764) );
  NAND3X0_HVT U771 ( .A1(n762), .A2(n763), .A3(n764), .Y(n233) );
  NBUFFX2_HVT U772 ( .A(n1027), .Y(cipher_text[24]) );
  NBUFFX2_HVT U773 ( .A(n1049), .Y(cipher_text[2]) );
  INVX0_HVT U774 ( .A(n774), .Y(cipher_text[33]) );
  INVX1_HVT U775 ( .A(n797), .Y(cipher_text[3]) );
  NBUFFX2_HVT U776 ( .A(n1009), .Y(cipher_text[42]) );
  NBUFFX2_HVT U777 ( .A(n1017), .Y(cipher_text[34]) );
  INVX0_HVT U778 ( .A(n971), .Y(n780) );
  INVX0_HVT U779 ( .A(n780), .Y(cipher_text[80]) );
  NAND2X0_HVT U780 ( .A1(n914), .A2(n1024), .Y(n782) );
  NAND2X0_HVT U781 ( .A1(adk_out0[27]), .A2(n888), .Y(n783) );
  NAND2X0_HVT U782 ( .A1(adk_in[27]), .A2(n848), .Y(n784) );
  NAND3X0_HVT U783 ( .A1(n782), .A2(n783), .A3(n784), .Y(n257) );
  INVX1_HVT U784 ( .A(n785), .Y(cipher_text[27]) );
  INVX0_HVT U785 ( .A(n1047), .Y(n787) );
  INVX0_HVT U786 ( .A(n970), .Y(n789) );
  INVX0_HVT U787 ( .A(n789), .Y(cipher_text[81]) );
  NAND2X0_HVT U788 ( .A1(n1048), .A2(n916), .Y(n794) );
  NAND2X0_HVT U789 ( .A1(adk_out0[3]), .A2(n890), .Y(n795) );
  NAND2X0_HVT U790 ( .A1(adk_in[3]), .A2(n846), .Y(n796) );
  NAND3X0_HVT U791 ( .A1(n794), .A2(n795), .A3(n796), .Y(n281) );
  INVX0_HVT U792 ( .A(n1048), .Y(n797) );
  INVX0_HVT U793 ( .A(n917), .Y(n916) );
  INVX1_HVT U794 ( .A(n865), .Y(n846) );
  INVX0_HVT U795 ( .A(n960), .Y(n799) );
  INVX0_HVT U796 ( .A(n799), .Y(cipher_text[91]) );
  NAND2X0_HVT U797 ( .A1(n959), .A2(n908), .Y(n801) );
  NAND2X0_HVT U798 ( .A1(adk_out0[92]), .A2(n882), .Y(n802) );
  NAND2X0_HVT U799 ( .A1(adk_in[92]), .A2(n852), .Y(n803) );
  NAND2X0_HVT U800 ( .A1(n976), .A2(n910), .Y(n804) );
  NAND2X0_HVT U801 ( .A1(adk_out0[75]), .A2(n884), .Y(n805) );
  NAND2X0_HVT U802 ( .A1(adk_in[75]), .A2(n850), .Y(n806) );
  NAND3X0_HVT U803 ( .A1(n804), .A2(n805), .A3(n806), .Y(n209) );
  INVX1_HVT U804 ( .A(n807), .Y(cipher_text[107]) );
  INVX0_HVT U805 ( .A(n809), .Y(cipher_text[111]) );
  NAND2X0_HVT U806 ( .A1(n936), .A2(n906), .Y(n811) );
  NAND2X0_HVT U807 ( .A1(adk_out0[115]), .A2(n880), .Y(n812) );
  NAND2X0_HVT U808 ( .A1(adk_in[115]), .A2(n853), .Y(n813) );
  NAND3X0_HVT U809 ( .A1(n811), .A2(n812), .A3(n813), .Y(n169) );
  INVX0_HVT U810 ( .A(n992), .Y(n818) );
  INVX0_HVT U811 ( .A(n928), .Y(n820) );
  INVX0_HVT U812 ( .A(n820), .Y(cipher_text[123]) );
  NAND2X0_HVT U813 ( .A1(n907), .A2(n944), .Y(n824) );
  NAND2X0_HVT U814 ( .A1(adk_out0[107]), .A2(n881), .Y(n825) );
  NAND2X0_HVT U815 ( .A1(adk_in[107]), .A2(n853), .Y(n826) );
  NAND3X0_HVT U816 ( .A1(n824), .A2(n825), .A3(n826), .Y(n177) );
  INVX0_HVT U817 ( .A(n829), .Y(cipher_text[52]) );
  INVX0_HVT U818 ( .A(n833), .Y(cipher_text[124]) );
  NAND2X0_HVT U819 ( .A1(n966), .A2(n909), .Y(n839) );
  NAND2X0_HVT U820 ( .A1(adk_out0[85]), .A2(n883), .Y(n840) );
  NAND2X0_HVT U821 ( .A1(adk_in[85]), .A2(n851), .Y(n841) );
  NAND3X0_HVT U822 ( .A1(n839), .A2(n840), .A3(n841), .Y(n199) );
  INVX1_HVT U823 ( .A(n842), .Y(cipher_text[85]) );
  INVX0_HVT U824 ( .A(n844), .Y(cipher_text[61]) );
  IBUFFX2_HVT U825 ( .A(n17), .Y(n867) );
  INVX0_HVT U826 ( .A(n17), .Y(n868) );
  INVX0_HVT U827 ( .A(n866), .Y(n864) );
  INVX0_HVT U828 ( .A(n15), .Y(n920) );
  INVX0_HVT U829 ( .A(n16), .Y(n894) );
  INVX1_HVT U830 ( .A(n919), .Y(n899) );
  INVX1_HVT U831 ( .A(n919), .Y(n900) );
  INVX1_HVT U832 ( .A(n919), .Y(n901) );
  INVX1_HVT U833 ( .A(n919), .Y(n902) );
  INVX1_HVT U834 ( .A(n919), .Y(n903) );
  INVX1_HVT U835 ( .A(n917), .Y(n915) );
  INVX1_HVT U836 ( .A(n919), .Y(n904) );
  INVX1_HVT U837 ( .A(n920), .Y(n895) );
  INVX1_HVT U838 ( .A(n920), .Y(n896) );
  INVX1_HVT U839 ( .A(n920), .Y(n897) );
  INVX1_HVT U840 ( .A(n920), .Y(n898) );
  INVX1_HVT U841 ( .A(n891), .Y(n885) );
  INVX1_HVT U842 ( .A(n891), .Y(n886) );
  INVX1_HVT U843 ( .A(n891), .Y(n887) );
  INVX1_HVT U844 ( .A(n891), .Y(n888) );
  INVX1_HVT U845 ( .A(n893), .Y(n873) );
  INVX1_HVT U846 ( .A(n893), .Y(n874) );
  INVX1_HVT U847 ( .A(n893), .Y(n875) );
  INVX1_HVT U848 ( .A(n893), .Y(n876) );
  INVX1_HVT U849 ( .A(n893), .Y(n877) );
  INVX1_HVT U850 ( .A(n892), .Y(n879) );
  INVX1_HVT U851 ( .A(n892), .Y(n880) );
  INVX1_HVT U852 ( .A(n892), .Y(n881) );
  INVX1_HVT U853 ( .A(n892), .Y(n882) );
  INVX1_HVT U854 ( .A(n892), .Y(n883) );
  INVX1_HVT U855 ( .A(n891), .Y(n889) );
  INVX1_HVT U856 ( .A(n893), .Y(n878) );
  INVX1_HVT U857 ( .A(n892), .Y(n884) );
  INVX1_HVT U858 ( .A(n894), .Y(n869) );
  INVX1_HVT U859 ( .A(n894), .Y(n870) );
  INVX1_HVT U860 ( .A(n894), .Y(n871) );
  INVX1_HVT U861 ( .A(n867), .Y(n856) );
  INVX1_HVT U862 ( .A(n867), .Y(n860) );
  INVX1_HVT U863 ( .A(n867), .Y(n859) );
  INVX1_HVT U864 ( .A(n867), .Y(n858) );
  INVX1_HVT U865 ( .A(n867), .Y(n857) );
  INVX1_HVT U866 ( .A(n866), .Y(n855) );
  INVX1_HVT U867 ( .A(n866), .Y(n854) );
  INVX1_HVT U868 ( .A(n866), .Y(n853) );
  INVX1_HVT U869 ( .A(n866), .Y(n852) );
  INVX1_HVT U870 ( .A(n866), .Y(n851) );
  INVX1_HVT U871 ( .A(n865), .Y(n847) );
  INVX1_HVT U872 ( .A(n865), .Y(n849) );
  INVX1_HVT U873 ( .A(n865), .Y(n848) );
  INVX1_HVT U874 ( .A(n894), .Y(n872) );
  INVX1_HVT U875 ( .A(n865), .Y(n850) );
  INVX1_HVT U876 ( .A(n867), .Y(n861) );
  INVX1_HVT U877 ( .A(n868), .Y(n862) );
  INVX1_HVT U878 ( .A(n868), .Y(n863) );
  INVX1_HVT U879 ( .A(n15), .Y(n917) );
  INVX1_HVT U880 ( .A(n17), .Y(n865) );
  INVX1_HVT U881 ( .A(n15), .Y(n919) );
  INVX1_HVT U882 ( .A(n15), .Y(n918) );
  INVX1_HVT U883 ( .A(n16), .Y(n891) );
  INVX1_HVT U884 ( .A(n16), .Y(n893) );
  INVX1_HVT U885 ( .A(n16), .Y(n892) );
  INVX1_HVT U886 ( .A(n17), .Y(n866) );
  INVX1_HVT U887 ( .A(reset), .Y(n921) );
  INVX0_HVT U888 ( .A(n12), .Y(n922) );
  INVX0_HVT U889 ( .A(n14), .Y(n923) );
endmodule

