
module RAM_memory ( data, addr, we, clk, rst, q );
  input [255:0] data;
  input [3:0] addr;
  output [255:0] q;
  input we, clk, rst;
  wire   N9, N10, N11, N12, \ram[15][255] , \ram[15][254] , \ram[15][253] ,
         \ram[15][252] , \ram[15][251] , \ram[15][250] , \ram[15][249] ,
         \ram[15][248] , \ram[15][247] , \ram[15][246] , \ram[15][245] ,
         \ram[15][244] , \ram[15][243] , \ram[15][242] , \ram[15][241] ,
         \ram[15][240] , \ram[15][239] , \ram[15][238] , \ram[15][237] ,
         \ram[15][236] , \ram[15][235] , \ram[15][234] , \ram[15][233] ,
         \ram[15][232] , \ram[15][231] , \ram[15][230] , \ram[15][229] ,
         \ram[15][228] , \ram[15][227] , \ram[15][226] , \ram[15][225] ,
         \ram[15][224] , \ram[15][223] , \ram[15][222] , \ram[15][221] ,
         \ram[15][220] , \ram[15][219] , \ram[15][218] , \ram[15][217] ,
         \ram[15][216] , \ram[15][215] , \ram[15][214] , \ram[15][213] ,
         \ram[15][212] , \ram[15][211] , \ram[15][210] , \ram[15][209] ,
         \ram[15][208] , \ram[15][207] , \ram[15][206] , \ram[15][205] ,
         \ram[15][204] , \ram[15][203] , \ram[15][202] , \ram[15][201] ,
         \ram[15][200] , \ram[15][199] , \ram[15][198] , \ram[15][197] ,
         \ram[15][196] , \ram[15][195] , \ram[15][194] , \ram[15][193] ,
         \ram[15][192] , \ram[15][191] , \ram[15][190] , \ram[15][189] ,
         \ram[15][188] , \ram[15][187] , \ram[15][186] , \ram[15][185] ,
         \ram[15][184] , \ram[15][183] , \ram[15][182] , \ram[15][181] ,
         \ram[15][180] , \ram[15][179] , \ram[15][178] , \ram[15][177] ,
         \ram[15][176] , \ram[15][175] , \ram[15][174] , \ram[15][173] ,
         \ram[15][172] , \ram[15][171] , \ram[15][170] , \ram[15][169] ,
         \ram[15][168] , \ram[15][167] , \ram[15][166] , \ram[15][165] ,
         \ram[15][164] , \ram[15][163] , \ram[15][162] , \ram[15][161] ,
         \ram[15][160] , \ram[15][159] , \ram[15][158] , \ram[15][157] ,
         \ram[15][156] , \ram[15][155] , \ram[15][154] , \ram[15][153] ,
         \ram[15][152] , \ram[15][151] , \ram[15][150] , \ram[15][149] ,
         \ram[15][148] , \ram[15][147] , \ram[15][146] , \ram[15][145] ,
         \ram[15][144] , \ram[15][143] , \ram[15][142] , \ram[15][141] ,
         \ram[15][140] , \ram[15][139] , \ram[15][138] , \ram[15][137] ,
         \ram[15][136] , \ram[15][135] , \ram[15][134] , \ram[15][133] ,
         \ram[15][132] , \ram[15][131] , \ram[15][130] , \ram[15][129] ,
         \ram[15][128] , \ram[15][127] , \ram[15][126] , \ram[15][125] ,
         \ram[15][124] , \ram[15][123] , \ram[15][122] , \ram[15][121] ,
         \ram[15][120] , \ram[15][119] , \ram[15][118] , \ram[15][117] ,
         \ram[15][116] , \ram[15][115] , \ram[15][114] , \ram[15][113] ,
         \ram[15][112] , \ram[15][111] , \ram[15][110] , \ram[15][109] ,
         \ram[15][108] , \ram[15][107] , \ram[15][106] , \ram[15][105] ,
         \ram[15][104] , \ram[15][103] , \ram[15][102] , \ram[15][101] ,
         \ram[15][100] , \ram[15][99] , \ram[15][98] , \ram[15][97] ,
         \ram[15][96] , \ram[15][95] , \ram[15][94] , \ram[15][93] ,
         \ram[15][92] , \ram[15][91] , \ram[15][90] , \ram[15][89] ,
         \ram[15][88] , \ram[15][87] , \ram[15][86] , \ram[15][85] ,
         \ram[15][84] , \ram[15][83] , \ram[15][82] , \ram[15][81] ,
         \ram[15][80] , \ram[15][79] , \ram[15][78] , \ram[15][77] ,
         \ram[15][76] , \ram[15][75] , \ram[15][74] , \ram[15][73] ,
         \ram[15][72] , \ram[15][71] , \ram[15][70] , \ram[15][69] ,
         \ram[15][68] , \ram[15][67] , \ram[15][66] , \ram[15][65] ,
         \ram[15][64] , \ram[15][63] , \ram[15][62] , \ram[15][61] ,
         \ram[15][60] , \ram[15][59] , \ram[15][58] , \ram[15][57] ,
         \ram[15][56] , \ram[15][55] , \ram[15][54] , \ram[15][53] ,
         \ram[15][52] , \ram[15][51] , \ram[15][50] , \ram[15][49] ,
         \ram[15][48] , \ram[15][47] , \ram[15][46] , \ram[15][45] ,
         \ram[15][44] , \ram[15][43] , \ram[15][42] , \ram[15][41] ,
         \ram[15][40] , \ram[15][39] , \ram[15][38] , \ram[15][37] ,
         \ram[15][36] , \ram[15][35] , \ram[15][34] , \ram[15][33] ,
         \ram[15][32] , \ram[15][31] , \ram[15][30] , \ram[15][29] ,
         \ram[15][28] , \ram[15][27] , \ram[15][26] , \ram[15][25] ,
         \ram[15][24] , \ram[15][23] , \ram[15][22] , \ram[15][21] ,
         \ram[15][20] , \ram[15][19] , \ram[15][18] , \ram[15][17] ,
         \ram[15][16] , \ram[15][15] , \ram[15][14] , \ram[15][13] ,
         \ram[15][12] , \ram[15][11] , \ram[15][10] , \ram[15][9] ,
         \ram[15][8] , \ram[15][7] , \ram[15][6] , \ram[15][5] , \ram[15][4] ,
         \ram[15][3] , \ram[15][2] , \ram[15][1] , \ram[15][0] ,
         \ram[14][255] , \ram[14][254] , \ram[14][253] , \ram[14][252] ,
         \ram[14][251] , \ram[14][250] , \ram[14][249] , \ram[14][248] ,
         \ram[14][247] , \ram[14][246] , \ram[14][245] , \ram[14][244] ,
         \ram[14][243] , \ram[14][242] , \ram[14][241] , \ram[14][240] ,
         \ram[14][239] , \ram[14][238] , \ram[14][237] , \ram[14][236] ,
         \ram[14][235] , \ram[14][234] , \ram[14][233] , \ram[14][232] ,
         \ram[14][231] , \ram[14][230] , \ram[14][229] , \ram[14][228] ,
         \ram[14][227] , \ram[14][226] , \ram[14][225] , \ram[14][224] ,
         \ram[14][223] , \ram[14][222] , \ram[14][221] , \ram[14][220] ,
         \ram[14][219] , \ram[14][218] , \ram[14][217] , \ram[14][216] ,
         \ram[14][215] , \ram[14][214] , \ram[14][213] , \ram[14][212] ,
         \ram[14][211] , \ram[14][210] , \ram[14][209] , \ram[14][208] ,
         \ram[14][207] , \ram[14][206] , \ram[14][205] , \ram[14][204] ,
         \ram[14][203] , \ram[14][202] , \ram[14][201] , \ram[14][200] ,
         \ram[14][199] , \ram[14][198] , \ram[14][197] , \ram[14][196] ,
         \ram[14][195] , \ram[14][194] , \ram[14][193] , \ram[14][192] ,
         \ram[14][191] , \ram[14][190] , \ram[14][189] , \ram[14][188] ,
         \ram[14][187] , \ram[14][186] , \ram[14][185] , \ram[14][184] ,
         \ram[14][183] , \ram[14][182] , \ram[14][181] , \ram[14][180] ,
         \ram[14][179] , \ram[14][178] , \ram[14][177] , \ram[14][176] ,
         \ram[14][175] , \ram[14][174] , \ram[14][173] , \ram[14][172] ,
         \ram[14][171] , \ram[14][170] , \ram[14][169] , \ram[14][168] ,
         \ram[14][167] , \ram[14][166] , \ram[14][165] , \ram[14][164] ,
         \ram[14][163] , \ram[14][162] , \ram[14][161] , \ram[14][160] ,
         \ram[14][159] , \ram[14][158] , \ram[14][157] , \ram[14][156] ,
         \ram[14][155] , \ram[14][154] , \ram[14][153] , \ram[14][152] ,
         \ram[14][151] , \ram[14][150] , \ram[14][149] , \ram[14][148] ,
         \ram[14][147] , \ram[14][146] , \ram[14][145] , \ram[14][144] ,
         \ram[14][143] , \ram[14][142] , \ram[14][141] , \ram[14][140] ,
         \ram[14][139] , \ram[14][138] , \ram[14][137] , \ram[14][136] ,
         \ram[14][135] , \ram[14][134] , \ram[14][133] , \ram[14][132] ,
         \ram[14][131] , \ram[14][130] , \ram[14][129] , \ram[14][128] ,
         \ram[14][127] , \ram[14][126] , \ram[14][125] , \ram[14][124] ,
         \ram[14][123] , \ram[14][122] , \ram[14][121] , \ram[14][120] ,
         \ram[14][119] , \ram[14][118] , \ram[14][117] , \ram[14][116] ,
         \ram[14][115] , \ram[14][114] , \ram[14][113] , \ram[14][112] ,
         \ram[14][111] , \ram[14][110] , \ram[14][109] , \ram[14][108] ,
         \ram[14][107] , \ram[14][106] , \ram[14][105] , \ram[14][104] ,
         \ram[14][103] , \ram[14][102] , \ram[14][101] , \ram[14][100] ,
         \ram[14][99] , \ram[14][98] , \ram[14][97] , \ram[14][96] ,
         \ram[14][95] , \ram[14][94] , \ram[14][93] , \ram[14][92] ,
         \ram[14][91] , \ram[14][90] , \ram[14][89] , \ram[14][88] ,
         \ram[14][87] , \ram[14][86] , \ram[14][85] , \ram[14][84] ,
         \ram[14][83] , \ram[14][82] , \ram[14][81] , \ram[14][80] ,
         \ram[14][79] , \ram[14][78] , \ram[14][77] , \ram[14][76] ,
         \ram[14][75] , \ram[14][74] , \ram[14][73] , \ram[14][72] ,
         \ram[14][71] , \ram[14][70] , \ram[14][69] , \ram[14][68] ,
         \ram[14][67] , \ram[14][66] , \ram[14][65] , \ram[14][64] ,
         \ram[14][63] , \ram[14][62] , \ram[14][61] , \ram[14][60] ,
         \ram[14][59] , \ram[14][58] , \ram[14][57] , \ram[14][56] ,
         \ram[14][55] , \ram[14][54] , \ram[14][53] , \ram[14][52] ,
         \ram[14][51] , \ram[14][50] , \ram[14][49] , \ram[14][48] ,
         \ram[14][47] , \ram[14][46] , \ram[14][45] , \ram[14][44] ,
         \ram[14][43] , \ram[14][42] , \ram[14][41] , \ram[14][40] ,
         \ram[14][39] , \ram[14][38] , \ram[14][37] , \ram[14][36] ,
         \ram[14][35] , \ram[14][34] , \ram[14][33] , \ram[14][32] ,
         \ram[14][31] , \ram[14][30] , \ram[14][29] , \ram[14][28] ,
         \ram[14][27] , \ram[14][26] , \ram[14][25] , \ram[14][24] ,
         \ram[14][23] , \ram[14][22] , \ram[14][21] , \ram[14][20] ,
         \ram[14][19] , \ram[14][18] , \ram[14][17] , \ram[14][16] ,
         \ram[14][15] , \ram[14][14] , \ram[14][13] , \ram[14][12] ,
         \ram[14][11] , \ram[14][10] , \ram[14][9] , \ram[14][8] ,
         \ram[14][7] , \ram[14][6] , \ram[14][5] , \ram[14][4] , \ram[14][3] ,
         \ram[14][2] , \ram[14][1] , \ram[14][0] , \ram[13][255] ,
         \ram[13][254] , \ram[13][253] , \ram[13][252] , \ram[13][251] ,
         \ram[13][250] , \ram[13][249] , \ram[13][248] , \ram[13][247] ,
         \ram[13][246] , \ram[13][245] , \ram[13][244] , \ram[13][243] ,
         \ram[13][242] , \ram[13][241] , \ram[13][240] , \ram[13][239] ,
         \ram[13][238] , \ram[13][237] , \ram[13][236] , \ram[13][235] ,
         \ram[13][234] , \ram[13][233] , \ram[13][232] , \ram[13][231] ,
         \ram[13][230] , \ram[13][229] , \ram[13][228] , \ram[13][227] ,
         \ram[13][226] , \ram[13][225] , \ram[13][224] , \ram[13][223] ,
         \ram[13][222] , \ram[13][221] , \ram[13][220] , \ram[13][219] ,
         \ram[13][218] , \ram[13][217] , \ram[13][216] , \ram[13][215] ,
         \ram[13][214] , \ram[13][213] , \ram[13][212] , \ram[13][211] ,
         \ram[13][210] , \ram[13][209] , \ram[13][208] , \ram[13][207] ,
         \ram[13][206] , \ram[13][205] , \ram[13][204] , \ram[13][203] ,
         \ram[13][202] , \ram[13][201] , \ram[13][200] , \ram[13][199] ,
         \ram[13][198] , \ram[13][197] , \ram[13][196] , \ram[13][195] ,
         \ram[13][194] , \ram[13][193] , \ram[13][192] , \ram[13][191] ,
         \ram[13][190] , \ram[13][189] , \ram[13][188] , \ram[13][187] ,
         \ram[13][186] , \ram[13][185] , \ram[13][184] , \ram[13][183] ,
         \ram[13][182] , \ram[13][181] , \ram[13][180] , \ram[13][179] ,
         \ram[13][178] , \ram[13][177] , \ram[13][176] , \ram[13][175] ,
         \ram[13][174] , \ram[13][173] , \ram[13][172] , \ram[13][171] ,
         \ram[13][170] , \ram[13][169] , \ram[13][168] , \ram[13][167] ,
         \ram[13][166] , \ram[13][165] , \ram[13][164] , \ram[13][163] ,
         \ram[13][162] , \ram[13][161] , \ram[13][160] , \ram[13][159] ,
         \ram[13][158] , \ram[13][157] , \ram[13][156] , \ram[13][155] ,
         \ram[13][154] , \ram[13][153] , \ram[13][152] , \ram[13][151] ,
         \ram[13][150] , \ram[13][149] , \ram[13][148] , \ram[13][147] ,
         \ram[13][146] , \ram[13][145] , \ram[13][144] , \ram[13][143] ,
         \ram[13][142] , \ram[13][141] , \ram[13][140] , \ram[13][139] ,
         \ram[13][138] , \ram[13][137] , \ram[13][136] , \ram[13][135] ,
         \ram[13][134] , \ram[13][133] , \ram[13][132] , \ram[13][131] ,
         \ram[13][130] , \ram[13][129] , \ram[13][128] , \ram[13][127] ,
         \ram[13][126] , \ram[13][125] , \ram[13][124] , \ram[13][123] ,
         \ram[13][122] , \ram[13][121] , \ram[13][120] , \ram[13][119] ,
         \ram[13][118] , \ram[13][117] , \ram[13][116] , \ram[13][115] ,
         \ram[13][114] , \ram[13][113] , \ram[13][112] , \ram[13][111] ,
         \ram[13][110] , \ram[13][109] , \ram[13][108] , \ram[13][107] ,
         \ram[13][106] , \ram[13][105] , \ram[13][104] , \ram[13][103] ,
         \ram[13][102] , \ram[13][101] , \ram[13][100] , \ram[13][99] ,
         \ram[13][98] , \ram[13][97] , \ram[13][96] , \ram[13][95] ,
         \ram[13][94] , \ram[13][93] , \ram[13][92] , \ram[13][91] ,
         \ram[13][90] , \ram[13][89] , \ram[13][88] , \ram[13][87] ,
         \ram[13][86] , \ram[13][85] , \ram[13][84] , \ram[13][83] ,
         \ram[13][82] , \ram[13][81] , \ram[13][80] , \ram[13][79] ,
         \ram[13][78] , \ram[13][77] , \ram[13][76] , \ram[13][75] ,
         \ram[13][74] , \ram[13][73] , \ram[13][72] , \ram[13][71] ,
         \ram[13][70] , \ram[13][69] , \ram[13][68] , \ram[13][67] ,
         \ram[13][66] , \ram[13][65] , \ram[13][64] , \ram[13][63] ,
         \ram[13][62] , \ram[13][61] , \ram[13][60] , \ram[13][59] ,
         \ram[13][58] , \ram[13][57] , \ram[13][56] , \ram[13][55] ,
         \ram[13][54] , \ram[13][53] , \ram[13][52] , \ram[13][51] ,
         \ram[13][50] , \ram[13][49] , \ram[13][48] , \ram[13][47] ,
         \ram[13][46] , \ram[13][45] , \ram[13][44] , \ram[13][43] ,
         \ram[13][42] , \ram[13][41] , \ram[13][40] , \ram[13][39] ,
         \ram[13][38] , \ram[13][37] , \ram[13][36] , \ram[13][35] ,
         \ram[13][34] , \ram[13][33] , \ram[13][32] , \ram[13][31] ,
         \ram[13][30] , \ram[13][29] , \ram[13][28] , \ram[13][27] ,
         \ram[13][26] , \ram[13][25] , \ram[13][24] , \ram[13][23] ,
         \ram[13][22] , \ram[13][21] , \ram[13][20] , \ram[13][19] ,
         \ram[13][18] , \ram[13][17] , \ram[13][16] , \ram[13][15] ,
         \ram[13][14] , \ram[13][13] , \ram[13][12] , \ram[13][11] ,
         \ram[13][10] , \ram[13][9] , \ram[13][8] , \ram[13][7] , \ram[13][6] ,
         \ram[13][5] , \ram[13][4] , \ram[13][3] , \ram[13][2] , \ram[13][1] ,
         \ram[13][0] , \ram[12][255] , \ram[12][254] , \ram[12][253] ,
         \ram[12][252] , \ram[12][251] , \ram[12][250] , \ram[12][249] ,
         \ram[12][248] , \ram[12][247] , \ram[12][246] , \ram[12][245] ,
         \ram[12][244] , \ram[12][243] , \ram[12][242] , \ram[12][241] ,
         \ram[12][240] , \ram[12][239] , \ram[12][238] , \ram[12][237] ,
         \ram[12][236] , \ram[12][235] , \ram[12][234] , \ram[12][233] ,
         \ram[12][232] , \ram[12][231] , \ram[12][230] , \ram[12][229] ,
         \ram[12][228] , \ram[12][227] , \ram[12][226] , \ram[12][225] ,
         \ram[12][224] , \ram[12][223] , \ram[12][222] , \ram[12][221] ,
         \ram[12][220] , \ram[12][219] , \ram[12][218] , \ram[12][217] ,
         \ram[12][216] , \ram[12][215] , \ram[12][214] , \ram[12][213] ,
         \ram[12][212] , \ram[12][211] , \ram[12][210] , \ram[12][209] ,
         \ram[12][208] , \ram[12][207] , \ram[12][206] , \ram[12][205] ,
         \ram[12][204] , \ram[12][203] , \ram[12][202] , \ram[12][201] ,
         \ram[12][200] , \ram[12][199] , \ram[12][198] , \ram[12][197] ,
         \ram[12][196] , \ram[12][195] , \ram[12][194] , \ram[12][193] ,
         \ram[12][192] , \ram[12][191] , \ram[12][190] , \ram[12][189] ,
         \ram[12][188] , \ram[12][187] , \ram[12][186] , \ram[12][185] ,
         \ram[12][184] , \ram[12][183] , \ram[12][182] , \ram[12][181] ,
         \ram[12][180] , \ram[12][179] , \ram[12][178] , \ram[12][177] ,
         \ram[12][176] , \ram[12][175] , \ram[12][174] , \ram[12][173] ,
         \ram[12][172] , \ram[12][171] , \ram[12][170] , \ram[12][169] ,
         \ram[12][168] , \ram[12][167] , \ram[12][166] , \ram[12][165] ,
         \ram[12][164] , \ram[12][163] , \ram[12][162] , \ram[12][161] ,
         \ram[12][160] , \ram[12][159] , \ram[12][158] , \ram[12][157] ,
         \ram[12][156] , \ram[12][155] , \ram[12][154] , \ram[12][153] ,
         \ram[12][152] , \ram[12][151] , \ram[12][150] , \ram[12][149] ,
         \ram[12][148] , \ram[12][147] , \ram[12][146] , \ram[12][145] ,
         \ram[12][144] , \ram[12][143] , \ram[12][142] , \ram[12][141] ,
         \ram[12][140] , \ram[12][139] , \ram[12][138] , \ram[12][137] ,
         \ram[12][136] , \ram[12][135] , \ram[12][134] , \ram[12][133] ,
         \ram[12][132] , \ram[12][131] , \ram[12][130] , \ram[12][129] ,
         \ram[12][128] , \ram[12][127] , \ram[12][126] , \ram[12][125] ,
         \ram[12][124] , \ram[12][123] , \ram[12][122] , \ram[12][121] ,
         \ram[12][120] , \ram[12][119] , \ram[12][118] , \ram[12][117] ,
         \ram[12][116] , \ram[12][115] , \ram[12][114] , \ram[12][113] ,
         \ram[12][112] , \ram[12][111] , \ram[12][110] , \ram[12][109] ,
         \ram[12][108] , \ram[12][107] , \ram[12][106] , \ram[12][105] ,
         \ram[12][104] , \ram[12][103] , \ram[12][102] , \ram[12][101] ,
         \ram[12][100] , \ram[12][99] , \ram[12][98] , \ram[12][97] ,
         \ram[12][96] , \ram[12][95] , \ram[12][94] , \ram[12][93] ,
         \ram[12][92] , \ram[12][91] , \ram[12][90] , \ram[12][89] ,
         \ram[12][88] , \ram[12][87] , \ram[12][86] , \ram[12][85] ,
         \ram[12][84] , \ram[12][83] , \ram[12][82] , \ram[12][81] ,
         \ram[12][80] , \ram[12][79] , \ram[12][78] , \ram[12][77] ,
         \ram[12][76] , \ram[12][75] , \ram[12][74] , \ram[12][73] ,
         \ram[12][72] , \ram[12][71] , \ram[12][70] , \ram[12][69] ,
         \ram[12][68] , \ram[12][67] , \ram[12][66] , \ram[12][65] ,
         \ram[12][64] , \ram[12][63] , \ram[12][62] , \ram[12][61] ,
         \ram[12][60] , \ram[12][59] , \ram[12][58] , \ram[12][57] ,
         \ram[12][56] , \ram[12][55] , \ram[12][54] , \ram[12][53] ,
         \ram[12][52] , \ram[12][51] , \ram[12][50] , \ram[12][49] ,
         \ram[12][48] , \ram[12][47] , \ram[12][46] , \ram[12][45] ,
         \ram[12][44] , \ram[12][43] , \ram[12][42] , \ram[12][41] ,
         \ram[12][40] , \ram[12][39] , \ram[12][38] , \ram[12][37] ,
         \ram[12][36] , \ram[12][35] , \ram[12][34] , \ram[12][33] ,
         \ram[12][32] , \ram[12][31] , \ram[12][30] , \ram[12][29] ,
         \ram[12][28] , \ram[12][27] , \ram[12][26] , \ram[12][25] ,
         \ram[12][24] , \ram[12][23] , \ram[12][22] , \ram[12][21] ,
         \ram[12][20] , \ram[12][19] , \ram[12][18] , \ram[12][17] ,
         \ram[12][16] , \ram[12][15] , \ram[12][14] , \ram[12][13] ,
         \ram[12][12] , \ram[12][11] , \ram[12][10] , \ram[12][9] ,
         \ram[12][8] , \ram[12][7] , \ram[12][6] , \ram[12][5] , \ram[12][4] ,
         \ram[12][3] , \ram[12][2] , \ram[12][1] , \ram[12][0] ,
         \ram[11][255] , \ram[11][254] , \ram[11][253] , \ram[11][252] ,
         \ram[11][251] , \ram[11][250] , \ram[11][249] , \ram[11][248] ,
         \ram[11][247] , \ram[11][246] , \ram[11][245] , \ram[11][244] ,
         \ram[11][243] , \ram[11][242] , \ram[11][241] , \ram[11][240] ,
         \ram[11][239] , \ram[11][238] , \ram[11][237] , \ram[11][236] ,
         \ram[11][235] , \ram[11][234] , \ram[11][233] , \ram[11][232] ,
         \ram[11][231] , \ram[11][230] , \ram[11][229] , \ram[11][228] ,
         \ram[11][227] , \ram[11][226] , \ram[11][225] , \ram[11][224] ,
         \ram[11][223] , \ram[11][222] , \ram[11][221] , \ram[11][220] ,
         \ram[11][219] , \ram[11][218] , \ram[11][217] , \ram[11][216] ,
         \ram[11][215] , \ram[11][214] , \ram[11][213] , \ram[11][212] ,
         \ram[11][211] , \ram[11][210] , \ram[11][209] , \ram[11][208] ,
         \ram[11][207] , \ram[11][206] , \ram[11][205] , \ram[11][204] ,
         \ram[11][203] , \ram[11][202] , \ram[11][201] , \ram[11][200] ,
         \ram[11][199] , \ram[11][198] , \ram[11][197] , \ram[11][196] ,
         \ram[11][195] , \ram[11][194] , \ram[11][193] , \ram[11][192] ,
         \ram[11][191] , \ram[11][190] , \ram[11][189] , \ram[11][188] ,
         \ram[11][187] , \ram[11][186] , \ram[11][185] , \ram[11][184] ,
         \ram[11][183] , \ram[11][182] , \ram[11][181] , \ram[11][180] ,
         \ram[11][179] , \ram[11][178] , \ram[11][177] , \ram[11][176] ,
         \ram[11][175] , \ram[11][174] , \ram[11][173] , \ram[11][172] ,
         \ram[11][171] , \ram[11][170] , \ram[11][169] , \ram[11][168] ,
         \ram[11][167] , \ram[11][166] , \ram[11][165] , \ram[11][164] ,
         \ram[11][163] , \ram[11][162] , \ram[11][161] , \ram[11][160] ,
         \ram[11][159] , \ram[11][158] , \ram[11][157] , \ram[11][156] ,
         \ram[11][155] , \ram[11][154] , \ram[11][153] , \ram[11][152] ,
         \ram[11][151] , \ram[11][150] , \ram[11][149] , \ram[11][148] ,
         \ram[11][147] , \ram[11][146] , \ram[11][145] , \ram[11][144] ,
         \ram[11][143] , \ram[11][142] , \ram[11][141] , \ram[11][140] ,
         \ram[11][139] , \ram[11][138] , \ram[11][137] , \ram[11][136] ,
         \ram[11][135] , \ram[11][134] , \ram[11][133] , \ram[11][132] ,
         \ram[11][131] , \ram[11][130] , \ram[11][129] , \ram[11][128] ,
         \ram[11][127] , \ram[11][126] , \ram[11][125] , \ram[11][124] ,
         \ram[11][123] , \ram[11][122] , \ram[11][121] , \ram[11][120] ,
         \ram[11][119] , \ram[11][118] , \ram[11][117] , \ram[11][116] ,
         \ram[11][115] , \ram[11][114] , \ram[11][113] , \ram[11][112] ,
         \ram[11][111] , \ram[11][110] , \ram[11][109] , \ram[11][108] ,
         \ram[11][107] , \ram[11][106] , \ram[11][105] , \ram[11][104] ,
         \ram[11][103] , \ram[11][102] , \ram[11][101] , \ram[11][100] ,
         \ram[11][99] , \ram[11][98] , \ram[11][97] , \ram[11][96] ,
         \ram[11][95] , \ram[11][94] , \ram[11][93] , \ram[11][92] ,
         \ram[11][91] , \ram[11][90] , \ram[11][89] , \ram[11][88] ,
         \ram[11][87] , \ram[11][86] , \ram[11][85] , \ram[11][84] ,
         \ram[11][83] , \ram[11][82] , \ram[11][81] , \ram[11][80] ,
         \ram[11][79] , \ram[11][78] , \ram[11][77] , \ram[11][76] ,
         \ram[11][75] , \ram[11][74] , \ram[11][73] , \ram[11][72] ,
         \ram[11][71] , \ram[11][70] , \ram[11][69] , \ram[11][68] ,
         \ram[11][67] , \ram[11][66] , \ram[11][65] , \ram[11][64] ,
         \ram[11][63] , \ram[11][62] , \ram[11][61] , \ram[11][60] ,
         \ram[11][59] , \ram[11][58] , \ram[11][57] , \ram[11][56] ,
         \ram[11][55] , \ram[11][54] , \ram[11][53] , \ram[11][52] ,
         \ram[11][51] , \ram[11][50] , \ram[11][49] , \ram[11][48] ,
         \ram[11][47] , \ram[11][46] , \ram[11][45] , \ram[11][44] ,
         \ram[11][43] , \ram[11][42] , \ram[11][41] , \ram[11][40] ,
         \ram[11][39] , \ram[11][38] , \ram[11][37] , \ram[11][36] ,
         \ram[11][35] , \ram[11][34] , \ram[11][33] , \ram[11][32] ,
         \ram[11][31] , \ram[11][30] , \ram[11][29] , \ram[11][28] ,
         \ram[11][27] , \ram[11][26] , \ram[11][25] , \ram[11][24] ,
         \ram[11][23] , \ram[11][22] , \ram[11][21] , \ram[11][20] ,
         \ram[11][19] , \ram[11][18] , \ram[11][17] , \ram[11][16] ,
         \ram[11][15] , \ram[11][14] , \ram[11][13] , \ram[11][12] ,
         \ram[11][11] , \ram[11][10] , \ram[11][9] , \ram[11][8] ,
         \ram[11][7] , \ram[11][6] , \ram[11][5] , \ram[11][4] , \ram[11][3] ,
         \ram[11][2] , \ram[11][1] , \ram[11][0] , \ram[10][255] ,
         \ram[10][254] , \ram[10][253] , \ram[10][252] , \ram[10][251] ,
         \ram[10][250] , \ram[10][249] , \ram[10][248] , \ram[10][247] ,
         \ram[10][246] , \ram[10][245] , \ram[10][244] , \ram[10][243] ,
         \ram[10][242] , \ram[10][241] , \ram[10][240] , \ram[10][239] ,
         \ram[10][238] , \ram[10][237] , \ram[10][236] , \ram[10][235] ,
         \ram[10][234] , \ram[10][233] , \ram[10][232] , \ram[10][231] ,
         \ram[10][230] , \ram[10][229] , \ram[10][228] , \ram[10][227] ,
         \ram[10][226] , \ram[10][225] , \ram[10][224] , \ram[10][223] ,
         \ram[10][222] , \ram[10][221] , \ram[10][220] , \ram[10][219] ,
         \ram[10][218] , \ram[10][217] , \ram[10][216] , \ram[10][215] ,
         \ram[10][214] , \ram[10][213] , \ram[10][212] , \ram[10][211] ,
         \ram[10][210] , \ram[10][209] , \ram[10][208] , \ram[10][207] ,
         \ram[10][206] , \ram[10][205] , \ram[10][204] , \ram[10][203] ,
         \ram[10][202] , \ram[10][201] , \ram[10][200] , \ram[10][199] ,
         \ram[10][198] , \ram[10][197] , \ram[10][196] , \ram[10][195] ,
         \ram[10][194] , \ram[10][193] , \ram[10][192] , \ram[10][191] ,
         \ram[10][190] , \ram[10][189] , \ram[10][188] , \ram[10][187] ,
         \ram[10][186] , \ram[10][185] , \ram[10][184] , \ram[10][183] ,
         \ram[10][182] , \ram[10][181] , \ram[10][180] , \ram[10][179] ,
         \ram[10][178] , \ram[10][177] , \ram[10][176] , \ram[10][175] ,
         \ram[10][174] , \ram[10][173] , \ram[10][172] , \ram[10][171] ,
         \ram[10][170] , \ram[10][169] , \ram[10][168] , \ram[10][167] ,
         \ram[10][166] , \ram[10][165] , \ram[10][164] , \ram[10][163] ,
         \ram[10][162] , \ram[10][161] , \ram[10][160] , \ram[10][159] ,
         \ram[10][158] , \ram[10][157] , \ram[10][156] , \ram[10][155] ,
         \ram[10][154] , \ram[10][153] , \ram[10][152] , \ram[10][151] ,
         \ram[10][150] , \ram[10][149] , \ram[10][148] , \ram[10][147] ,
         \ram[10][146] , \ram[10][145] , \ram[10][144] , \ram[10][143] ,
         \ram[10][142] , \ram[10][141] , \ram[10][140] , \ram[10][139] ,
         \ram[10][138] , \ram[10][137] , \ram[10][136] , \ram[10][135] ,
         \ram[10][134] , \ram[10][133] , \ram[10][132] , \ram[10][131] ,
         \ram[10][130] , \ram[10][129] , \ram[10][128] , \ram[10][127] ,
         \ram[10][126] , \ram[10][125] , \ram[10][124] , \ram[10][123] ,
         \ram[10][122] , \ram[10][121] , \ram[10][120] , \ram[10][119] ,
         \ram[10][118] , \ram[10][117] , \ram[10][116] , \ram[10][115] ,
         \ram[10][114] , \ram[10][113] , \ram[10][112] , \ram[10][111] ,
         \ram[10][110] , \ram[10][109] , \ram[10][108] , \ram[10][107] ,
         \ram[10][106] , \ram[10][105] , \ram[10][104] , \ram[10][103] ,
         \ram[10][102] , \ram[10][101] , \ram[10][100] , \ram[10][99] ,
         \ram[10][98] , \ram[10][97] , \ram[10][96] , \ram[10][95] ,
         \ram[10][94] , \ram[10][93] , \ram[10][92] , \ram[10][91] ,
         \ram[10][90] , \ram[10][89] , \ram[10][88] , \ram[10][87] ,
         \ram[10][86] , \ram[10][85] , \ram[10][84] , \ram[10][83] ,
         \ram[10][82] , \ram[10][81] , \ram[10][80] , \ram[10][79] ,
         \ram[10][78] , \ram[10][77] , \ram[10][76] , \ram[10][75] ,
         \ram[10][74] , \ram[10][73] , \ram[10][72] , \ram[10][71] ,
         \ram[10][70] , \ram[10][69] , \ram[10][68] , \ram[10][67] ,
         \ram[10][66] , \ram[10][65] , \ram[10][64] , \ram[10][63] ,
         \ram[10][62] , \ram[10][61] , \ram[10][60] , \ram[10][59] ,
         \ram[10][58] , \ram[10][57] , \ram[10][56] , \ram[10][55] ,
         \ram[10][54] , \ram[10][53] , \ram[10][52] , \ram[10][51] ,
         \ram[10][50] , \ram[10][49] , \ram[10][48] , \ram[10][47] ,
         \ram[10][46] , \ram[10][45] , \ram[10][44] , \ram[10][43] ,
         \ram[10][42] , \ram[10][41] , \ram[10][40] , \ram[10][39] ,
         \ram[10][38] , \ram[10][37] , \ram[10][36] , \ram[10][35] ,
         \ram[10][34] , \ram[10][33] , \ram[10][32] , \ram[10][31] ,
         \ram[10][30] , \ram[10][29] , \ram[10][28] , \ram[10][27] ,
         \ram[10][26] , \ram[10][25] , \ram[10][24] , \ram[10][23] ,
         \ram[10][22] , \ram[10][21] , \ram[10][20] , \ram[10][19] ,
         \ram[10][18] , \ram[10][17] , \ram[10][16] , \ram[10][15] ,
         \ram[10][14] , \ram[10][13] , \ram[10][12] , \ram[10][11] ,
         \ram[10][10] , \ram[10][9] , \ram[10][8] , \ram[10][7] , \ram[10][6] ,
         \ram[10][5] , \ram[10][4] , \ram[10][3] , \ram[10][2] , \ram[10][1] ,
         \ram[10][0] , \ram[9][255] , \ram[9][254] , \ram[9][253] ,
         \ram[9][252] , \ram[9][251] , \ram[9][250] , \ram[9][249] ,
         \ram[9][248] , \ram[9][247] , \ram[9][246] , \ram[9][245] ,
         \ram[9][244] , \ram[9][243] , \ram[9][242] , \ram[9][241] ,
         \ram[9][240] , \ram[9][239] , \ram[9][238] , \ram[9][237] ,
         \ram[9][236] , \ram[9][235] , \ram[9][234] , \ram[9][233] ,
         \ram[9][232] , \ram[9][231] , \ram[9][230] , \ram[9][229] ,
         \ram[9][228] , \ram[9][227] , \ram[9][226] , \ram[9][225] ,
         \ram[9][224] , \ram[9][223] , \ram[9][222] , \ram[9][221] ,
         \ram[9][220] , \ram[9][219] , \ram[9][218] , \ram[9][217] ,
         \ram[9][216] , \ram[9][215] , \ram[9][214] , \ram[9][213] ,
         \ram[9][212] , \ram[9][211] , \ram[9][210] , \ram[9][209] ,
         \ram[9][208] , \ram[9][207] , \ram[9][206] , \ram[9][205] ,
         \ram[9][204] , \ram[9][203] , \ram[9][202] , \ram[9][201] ,
         \ram[9][200] , \ram[9][199] , \ram[9][198] , \ram[9][197] ,
         \ram[9][196] , \ram[9][195] , \ram[9][194] , \ram[9][193] ,
         \ram[9][192] , \ram[9][191] , \ram[9][190] , \ram[9][189] ,
         \ram[9][188] , \ram[9][187] , \ram[9][186] , \ram[9][185] ,
         \ram[9][184] , \ram[9][183] , \ram[9][182] , \ram[9][181] ,
         \ram[9][180] , \ram[9][179] , \ram[9][178] , \ram[9][177] ,
         \ram[9][176] , \ram[9][175] , \ram[9][174] , \ram[9][173] ,
         \ram[9][172] , \ram[9][171] , \ram[9][170] , \ram[9][169] ,
         \ram[9][168] , \ram[9][167] , \ram[9][166] , \ram[9][165] ,
         \ram[9][164] , \ram[9][163] , \ram[9][162] , \ram[9][161] ,
         \ram[9][160] , \ram[9][159] , \ram[9][158] , \ram[9][157] ,
         \ram[9][156] , \ram[9][155] , \ram[9][154] , \ram[9][153] ,
         \ram[9][152] , \ram[9][151] , \ram[9][150] , \ram[9][149] ,
         \ram[9][148] , \ram[9][147] , \ram[9][146] , \ram[9][145] ,
         \ram[9][144] , \ram[9][143] , \ram[9][142] , \ram[9][141] ,
         \ram[9][140] , \ram[9][139] , \ram[9][138] , \ram[9][137] ,
         \ram[9][136] , \ram[9][135] , \ram[9][134] , \ram[9][133] ,
         \ram[9][132] , \ram[9][131] , \ram[9][130] , \ram[9][129] ,
         \ram[9][128] , \ram[9][127] , \ram[9][126] , \ram[9][125] ,
         \ram[9][124] , \ram[9][123] , \ram[9][122] , \ram[9][121] ,
         \ram[9][120] , \ram[9][119] , \ram[9][118] , \ram[9][117] ,
         \ram[9][116] , \ram[9][115] , \ram[9][114] , \ram[9][113] ,
         \ram[9][112] , \ram[9][111] , \ram[9][110] , \ram[9][109] ,
         \ram[9][108] , \ram[9][107] , \ram[9][106] , \ram[9][105] ,
         \ram[9][104] , \ram[9][103] , \ram[9][102] , \ram[9][101] ,
         \ram[9][100] , \ram[9][99] , \ram[9][98] , \ram[9][97] , \ram[9][96] ,
         \ram[9][95] , \ram[9][94] , \ram[9][93] , \ram[9][92] , \ram[9][91] ,
         \ram[9][90] , \ram[9][89] , \ram[9][88] , \ram[9][87] , \ram[9][86] ,
         \ram[9][85] , \ram[9][84] , \ram[9][83] , \ram[9][82] , \ram[9][81] ,
         \ram[9][80] , \ram[9][79] , \ram[9][78] , \ram[9][77] , \ram[9][76] ,
         \ram[9][75] , \ram[9][74] , \ram[9][73] , \ram[9][72] , \ram[9][71] ,
         \ram[9][70] , \ram[9][69] , \ram[9][68] , \ram[9][67] , \ram[9][66] ,
         \ram[9][65] , \ram[9][64] , \ram[9][63] , \ram[9][62] , \ram[9][61] ,
         \ram[9][60] , \ram[9][59] , \ram[9][58] , \ram[9][57] , \ram[9][56] ,
         \ram[9][55] , \ram[9][54] , \ram[9][53] , \ram[9][52] , \ram[9][51] ,
         \ram[9][50] , \ram[9][49] , \ram[9][48] , \ram[9][47] , \ram[9][46] ,
         \ram[9][45] , \ram[9][44] , \ram[9][43] , \ram[9][42] , \ram[9][41] ,
         \ram[9][40] , \ram[9][39] , \ram[9][38] , \ram[9][37] , \ram[9][36] ,
         \ram[9][35] , \ram[9][34] , \ram[9][33] , \ram[9][32] , \ram[9][31] ,
         \ram[9][30] , \ram[9][29] , \ram[9][28] , \ram[9][27] , \ram[9][26] ,
         \ram[9][25] , \ram[9][24] , \ram[9][23] , \ram[9][22] , \ram[9][21] ,
         \ram[9][20] , \ram[9][19] , \ram[9][18] , \ram[9][17] , \ram[9][16] ,
         \ram[9][15] , \ram[9][14] , \ram[9][13] , \ram[9][12] , \ram[9][11] ,
         \ram[9][10] , \ram[9][9] , \ram[9][8] , \ram[9][7] , \ram[9][6] ,
         \ram[9][5] , \ram[9][4] , \ram[9][3] , \ram[9][2] , \ram[9][1] ,
         \ram[9][0] , \ram[8][255] , \ram[8][254] , \ram[8][253] ,
         \ram[8][252] , \ram[8][251] , \ram[8][250] , \ram[8][249] ,
         \ram[8][248] , \ram[8][247] , \ram[8][246] , \ram[8][245] ,
         \ram[8][244] , \ram[8][243] , \ram[8][242] , \ram[8][241] ,
         \ram[8][240] , \ram[8][239] , \ram[8][238] , \ram[8][237] ,
         \ram[8][236] , \ram[8][235] , \ram[8][234] , \ram[8][233] ,
         \ram[8][232] , \ram[8][231] , \ram[8][230] , \ram[8][229] ,
         \ram[8][228] , \ram[8][227] , \ram[8][226] , \ram[8][225] ,
         \ram[8][224] , \ram[8][223] , \ram[8][222] , \ram[8][221] ,
         \ram[8][220] , \ram[8][219] , \ram[8][218] , \ram[8][217] ,
         \ram[8][216] , \ram[8][215] , \ram[8][214] , \ram[8][213] ,
         \ram[8][212] , \ram[8][211] , \ram[8][210] , \ram[8][209] ,
         \ram[8][208] , \ram[8][207] , \ram[8][206] , \ram[8][205] ,
         \ram[8][204] , \ram[8][203] , \ram[8][202] , \ram[8][201] ,
         \ram[8][200] , \ram[8][199] , \ram[8][198] , \ram[8][197] ,
         \ram[8][196] , \ram[8][195] , \ram[8][194] , \ram[8][193] ,
         \ram[8][192] , \ram[8][191] , \ram[8][190] , \ram[8][189] ,
         \ram[8][188] , \ram[8][187] , \ram[8][186] , \ram[8][185] ,
         \ram[8][184] , \ram[8][183] , \ram[8][182] , \ram[8][181] ,
         \ram[8][180] , \ram[8][179] , \ram[8][178] , \ram[8][177] ,
         \ram[8][176] , \ram[8][175] , \ram[8][174] , \ram[8][173] ,
         \ram[8][172] , \ram[8][171] , \ram[8][170] , \ram[8][169] ,
         \ram[8][168] , \ram[8][167] , \ram[8][166] , \ram[8][165] ,
         \ram[8][164] , \ram[8][163] , \ram[8][162] , \ram[8][161] ,
         \ram[8][160] , \ram[8][159] , \ram[8][158] , \ram[8][157] ,
         \ram[8][156] , \ram[8][155] , \ram[8][154] , \ram[8][153] ,
         \ram[8][152] , \ram[8][151] , \ram[8][150] , \ram[8][149] ,
         \ram[8][148] , \ram[8][147] , \ram[8][146] , \ram[8][145] ,
         \ram[8][144] , \ram[8][143] , \ram[8][142] , \ram[8][141] ,
         \ram[8][140] , \ram[8][139] , \ram[8][138] , \ram[8][137] ,
         \ram[8][136] , \ram[8][135] , \ram[8][134] , \ram[8][133] ,
         \ram[8][132] , \ram[8][131] , \ram[8][130] , \ram[8][129] ,
         \ram[8][128] , \ram[8][127] , \ram[8][126] , \ram[8][125] ,
         \ram[8][124] , \ram[8][123] , \ram[8][122] , \ram[8][121] ,
         \ram[8][120] , \ram[8][119] , \ram[8][118] , \ram[8][117] ,
         \ram[8][116] , \ram[8][115] , \ram[8][114] , \ram[8][113] ,
         \ram[8][112] , \ram[8][111] , \ram[8][110] , \ram[8][109] ,
         \ram[8][108] , \ram[8][107] , \ram[8][106] , \ram[8][105] ,
         \ram[8][104] , \ram[8][103] , \ram[8][102] , \ram[8][101] ,
         \ram[8][100] , \ram[8][99] , \ram[8][98] , \ram[8][97] , \ram[8][96] ,
         \ram[8][95] , \ram[8][94] , \ram[8][93] , \ram[8][92] , \ram[8][91] ,
         \ram[8][90] , \ram[8][89] , \ram[8][88] , \ram[8][87] , \ram[8][86] ,
         \ram[8][85] , \ram[8][84] , \ram[8][83] , \ram[8][82] , \ram[8][81] ,
         \ram[8][80] , \ram[8][79] , \ram[8][78] , \ram[8][77] , \ram[8][76] ,
         \ram[8][75] , \ram[8][74] , \ram[8][73] , \ram[8][72] , \ram[8][71] ,
         \ram[8][70] , \ram[8][69] , \ram[8][68] , \ram[8][67] , \ram[8][66] ,
         \ram[8][65] , \ram[8][64] , \ram[8][63] , \ram[8][62] , \ram[8][61] ,
         \ram[8][60] , \ram[8][59] , \ram[8][58] , \ram[8][57] , \ram[8][56] ,
         \ram[8][55] , \ram[8][54] , \ram[8][53] , \ram[8][52] , \ram[8][51] ,
         \ram[8][50] , \ram[8][49] , \ram[8][48] , \ram[8][47] , \ram[8][46] ,
         \ram[8][45] , \ram[8][44] , \ram[8][43] , \ram[8][42] , \ram[8][41] ,
         \ram[8][40] , \ram[8][39] , \ram[8][38] , \ram[8][37] , \ram[8][36] ,
         \ram[8][35] , \ram[8][34] , \ram[8][33] , \ram[8][32] , \ram[8][31] ,
         \ram[8][30] , \ram[8][29] , \ram[8][28] , \ram[8][27] , \ram[8][26] ,
         \ram[8][25] , \ram[8][24] , \ram[8][23] , \ram[8][22] , \ram[8][21] ,
         \ram[8][20] , \ram[8][19] , \ram[8][18] , \ram[8][17] , \ram[8][16] ,
         \ram[8][15] , \ram[8][14] , \ram[8][13] , \ram[8][12] , \ram[8][11] ,
         \ram[8][10] , \ram[8][9] , \ram[8][8] , \ram[8][7] , \ram[8][6] ,
         \ram[8][5] , \ram[8][4] , \ram[8][3] , \ram[8][2] , \ram[8][1] ,
         \ram[8][0] , \ram[7][255] , \ram[7][254] , \ram[7][253] ,
         \ram[7][252] , \ram[7][251] , \ram[7][250] , \ram[7][249] ,
         \ram[7][248] , \ram[7][247] , \ram[7][246] , \ram[7][245] ,
         \ram[7][244] , \ram[7][243] , \ram[7][242] , \ram[7][241] ,
         \ram[7][240] , \ram[7][239] , \ram[7][238] , \ram[7][237] ,
         \ram[7][236] , \ram[7][235] , \ram[7][234] , \ram[7][233] ,
         \ram[7][232] , \ram[7][231] , \ram[7][230] , \ram[7][229] ,
         \ram[7][228] , \ram[7][227] , \ram[7][226] , \ram[7][225] ,
         \ram[7][224] , \ram[7][223] , \ram[7][222] , \ram[7][221] ,
         \ram[7][220] , \ram[7][219] , \ram[7][218] , \ram[7][217] ,
         \ram[7][216] , \ram[7][215] , \ram[7][214] , \ram[7][213] ,
         \ram[7][212] , \ram[7][211] , \ram[7][210] , \ram[7][209] ,
         \ram[7][208] , \ram[7][207] , \ram[7][206] , \ram[7][205] ,
         \ram[7][204] , \ram[7][203] , \ram[7][202] , \ram[7][201] ,
         \ram[7][200] , \ram[7][199] , \ram[7][198] , \ram[7][197] ,
         \ram[7][196] , \ram[7][195] , \ram[7][194] , \ram[7][193] ,
         \ram[7][192] , \ram[7][191] , \ram[7][190] , \ram[7][189] ,
         \ram[7][188] , \ram[7][187] , \ram[7][186] , \ram[7][185] ,
         \ram[7][184] , \ram[7][183] , \ram[7][182] , \ram[7][181] ,
         \ram[7][180] , \ram[7][179] , \ram[7][178] , \ram[7][177] ,
         \ram[7][176] , \ram[7][175] , \ram[7][174] , \ram[7][173] ,
         \ram[7][172] , \ram[7][171] , \ram[7][170] , \ram[7][169] ,
         \ram[7][168] , \ram[7][167] , \ram[7][166] , \ram[7][165] ,
         \ram[7][164] , \ram[7][163] , \ram[7][162] , \ram[7][161] ,
         \ram[7][160] , \ram[7][159] , \ram[7][158] , \ram[7][157] ,
         \ram[7][156] , \ram[7][155] , \ram[7][154] , \ram[7][153] ,
         \ram[7][152] , \ram[7][151] , \ram[7][150] , \ram[7][149] ,
         \ram[7][148] , \ram[7][147] , \ram[7][146] , \ram[7][145] ,
         \ram[7][144] , \ram[7][143] , \ram[7][142] , \ram[7][141] ,
         \ram[7][140] , \ram[7][139] , \ram[7][138] , \ram[7][137] ,
         \ram[7][136] , \ram[7][135] , \ram[7][134] , \ram[7][133] ,
         \ram[7][132] , \ram[7][131] , \ram[7][130] , \ram[7][129] ,
         \ram[7][128] , \ram[7][127] , \ram[7][126] , \ram[7][125] ,
         \ram[7][124] , \ram[7][123] , \ram[7][122] , \ram[7][121] ,
         \ram[7][120] , \ram[7][119] , \ram[7][118] , \ram[7][117] ,
         \ram[7][116] , \ram[7][115] , \ram[7][114] , \ram[7][113] ,
         \ram[7][112] , \ram[7][111] , \ram[7][110] , \ram[7][109] ,
         \ram[7][108] , \ram[7][107] , \ram[7][106] , \ram[7][105] ,
         \ram[7][104] , \ram[7][103] , \ram[7][102] , \ram[7][101] ,
         \ram[7][100] , \ram[7][99] , \ram[7][98] , \ram[7][97] , \ram[7][96] ,
         \ram[7][95] , \ram[7][94] , \ram[7][93] , \ram[7][92] , \ram[7][91] ,
         \ram[7][90] , \ram[7][89] , \ram[7][88] , \ram[7][87] , \ram[7][86] ,
         \ram[7][85] , \ram[7][84] , \ram[7][83] , \ram[7][82] , \ram[7][81] ,
         \ram[7][80] , \ram[7][79] , \ram[7][78] , \ram[7][77] , \ram[7][76] ,
         \ram[7][75] , \ram[7][74] , \ram[7][73] , \ram[7][72] , \ram[7][71] ,
         \ram[7][70] , \ram[7][69] , \ram[7][68] , \ram[7][67] , \ram[7][66] ,
         \ram[7][65] , \ram[7][64] , \ram[7][63] , \ram[7][62] , \ram[7][61] ,
         \ram[7][60] , \ram[7][59] , \ram[7][58] , \ram[7][57] , \ram[7][56] ,
         \ram[7][55] , \ram[7][54] , \ram[7][53] , \ram[7][52] , \ram[7][51] ,
         \ram[7][50] , \ram[7][49] , \ram[7][48] , \ram[7][47] , \ram[7][46] ,
         \ram[7][45] , \ram[7][44] , \ram[7][43] , \ram[7][42] , \ram[7][41] ,
         \ram[7][40] , \ram[7][39] , \ram[7][38] , \ram[7][37] , \ram[7][36] ,
         \ram[7][35] , \ram[7][34] , \ram[7][33] , \ram[7][32] , \ram[7][31] ,
         \ram[7][30] , \ram[7][29] , \ram[7][28] , \ram[7][27] , \ram[7][26] ,
         \ram[7][25] , \ram[7][24] , \ram[7][23] , \ram[7][22] , \ram[7][21] ,
         \ram[7][20] , \ram[7][19] , \ram[7][18] , \ram[7][17] , \ram[7][16] ,
         \ram[7][15] , \ram[7][14] , \ram[7][13] , \ram[7][12] , \ram[7][11] ,
         \ram[7][10] , \ram[7][9] , \ram[7][8] , \ram[7][7] , \ram[7][6] ,
         \ram[7][5] , \ram[7][4] , \ram[7][3] , \ram[7][2] , \ram[7][1] ,
         \ram[7][0] , \ram[6][255] , \ram[6][254] , \ram[6][253] ,
         \ram[6][252] , \ram[6][251] , \ram[6][250] , \ram[6][249] ,
         \ram[6][248] , \ram[6][247] , \ram[6][246] , \ram[6][245] ,
         \ram[6][244] , \ram[6][243] , \ram[6][242] , \ram[6][241] ,
         \ram[6][240] , \ram[6][239] , \ram[6][238] , \ram[6][237] ,
         \ram[6][236] , \ram[6][235] , \ram[6][234] , \ram[6][233] ,
         \ram[6][232] , \ram[6][231] , \ram[6][230] , \ram[6][229] ,
         \ram[6][228] , \ram[6][227] , \ram[6][226] , \ram[6][225] ,
         \ram[6][224] , \ram[6][223] , \ram[6][222] , \ram[6][221] ,
         \ram[6][220] , \ram[6][219] , \ram[6][218] , \ram[6][217] ,
         \ram[6][216] , \ram[6][215] , \ram[6][214] , \ram[6][213] ,
         \ram[6][212] , \ram[6][211] , \ram[6][210] , \ram[6][209] ,
         \ram[6][208] , \ram[6][207] , \ram[6][206] , \ram[6][205] ,
         \ram[6][204] , \ram[6][203] , \ram[6][202] , \ram[6][201] ,
         \ram[6][200] , \ram[6][199] , \ram[6][198] , \ram[6][197] ,
         \ram[6][196] , \ram[6][195] , \ram[6][194] , \ram[6][193] ,
         \ram[6][192] , \ram[6][191] , \ram[6][190] , \ram[6][189] ,
         \ram[6][188] , \ram[6][187] , \ram[6][186] , \ram[6][185] ,
         \ram[6][184] , \ram[6][183] , \ram[6][182] , \ram[6][181] ,
         \ram[6][180] , \ram[6][179] , \ram[6][178] , \ram[6][177] ,
         \ram[6][176] , \ram[6][175] , \ram[6][174] , \ram[6][173] ,
         \ram[6][172] , \ram[6][171] , \ram[6][170] , \ram[6][169] ,
         \ram[6][168] , \ram[6][167] , \ram[6][166] , \ram[6][165] ,
         \ram[6][164] , \ram[6][163] , \ram[6][162] , \ram[6][161] ,
         \ram[6][160] , \ram[6][159] , \ram[6][158] , \ram[6][157] ,
         \ram[6][156] , \ram[6][155] , \ram[6][154] , \ram[6][153] ,
         \ram[6][152] , \ram[6][151] , \ram[6][150] , \ram[6][149] ,
         \ram[6][148] , \ram[6][147] , \ram[6][146] , \ram[6][145] ,
         \ram[6][144] , \ram[6][143] , \ram[6][142] , \ram[6][141] ,
         \ram[6][140] , \ram[6][139] , \ram[6][138] , \ram[6][137] ,
         \ram[6][136] , \ram[6][135] , \ram[6][134] , \ram[6][133] ,
         \ram[6][132] , \ram[6][131] , \ram[6][130] , \ram[6][129] ,
         \ram[6][128] , \ram[6][127] , \ram[6][126] , \ram[6][125] ,
         \ram[6][124] , \ram[6][123] , \ram[6][122] , \ram[6][121] ,
         \ram[6][120] , \ram[6][119] , \ram[6][118] , \ram[6][117] ,
         \ram[6][116] , \ram[6][115] , \ram[6][114] , \ram[6][113] ,
         \ram[6][112] , \ram[6][111] , \ram[6][110] , \ram[6][109] ,
         \ram[6][108] , \ram[6][107] , \ram[6][106] , \ram[6][105] ,
         \ram[6][104] , \ram[6][103] , \ram[6][102] , \ram[6][101] ,
         \ram[6][100] , \ram[6][99] , \ram[6][98] , \ram[6][97] , \ram[6][96] ,
         \ram[6][95] , \ram[6][94] , \ram[6][93] , \ram[6][92] , \ram[6][91] ,
         \ram[6][90] , \ram[6][89] , \ram[6][88] , \ram[6][87] , \ram[6][86] ,
         \ram[6][85] , \ram[6][84] , \ram[6][83] , \ram[6][82] , \ram[6][81] ,
         \ram[6][80] , \ram[6][79] , \ram[6][78] , \ram[6][77] , \ram[6][76] ,
         \ram[6][75] , \ram[6][74] , \ram[6][73] , \ram[6][72] , \ram[6][71] ,
         \ram[6][70] , \ram[6][69] , \ram[6][68] , \ram[6][67] , \ram[6][66] ,
         \ram[6][65] , \ram[6][64] , \ram[6][63] , \ram[6][62] , \ram[6][61] ,
         \ram[6][60] , \ram[6][59] , \ram[6][58] , \ram[6][57] , \ram[6][56] ,
         \ram[6][55] , \ram[6][54] , \ram[6][53] , \ram[6][52] , \ram[6][51] ,
         \ram[6][50] , \ram[6][49] , \ram[6][48] , \ram[6][47] , \ram[6][46] ,
         \ram[6][45] , \ram[6][44] , \ram[6][43] , \ram[6][42] , \ram[6][41] ,
         \ram[6][40] , \ram[6][39] , \ram[6][38] , \ram[6][37] , \ram[6][36] ,
         \ram[6][35] , \ram[6][34] , \ram[6][33] , \ram[6][32] , \ram[6][31] ,
         \ram[6][30] , \ram[6][29] , \ram[6][28] , \ram[6][27] , \ram[6][26] ,
         \ram[6][25] , \ram[6][24] , \ram[6][23] , \ram[6][22] , \ram[6][21] ,
         \ram[6][20] , \ram[6][19] , \ram[6][18] , \ram[6][17] , \ram[6][16] ,
         \ram[6][15] , \ram[6][14] , \ram[6][13] , \ram[6][12] , \ram[6][11] ,
         \ram[6][10] , \ram[6][9] , \ram[6][8] , \ram[6][7] , \ram[6][6] ,
         \ram[6][5] , \ram[6][4] , \ram[6][3] , \ram[6][2] , \ram[6][1] ,
         \ram[6][0] , \ram[5][255] , \ram[5][254] , \ram[5][253] ,
         \ram[5][252] , \ram[5][251] , \ram[5][250] , \ram[5][249] ,
         \ram[5][248] , \ram[5][247] , \ram[5][246] , \ram[5][245] ,
         \ram[5][244] , \ram[5][243] , \ram[5][242] , \ram[5][241] ,
         \ram[5][240] , \ram[5][239] , \ram[5][238] , \ram[5][237] ,
         \ram[5][236] , \ram[5][235] , \ram[5][234] , \ram[5][233] ,
         \ram[5][232] , \ram[5][231] , \ram[5][230] , \ram[5][229] ,
         \ram[5][228] , \ram[5][227] , \ram[5][226] , \ram[5][225] ,
         \ram[5][224] , \ram[5][223] , \ram[5][222] , \ram[5][221] ,
         \ram[5][220] , \ram[5][219] , \ram[5][218] , \ram[5][217] ,
         \ram[5][216] , \ram[5][215] , \ram[5][214] , \ram[5][213] ,
         \ram[5][212] , \ram[5][211] , \ram[5][210] , \ram[5][209] ,
         \ram[5][208] , \ram[5][207] , \ram[5][206] , \ram[5][205] ,
         \ram[5][204] , \ram[5][203] , \ram[5][202] , \ram[5][201] ,
         \ram[5][200] , \ram[5][199] , \ram[5][198] , \ram[5][197] ,
         \ram[5][196] , \ram[5][195] , \ram[5][194] , \ram[5][193] ,
         \ram[5][192] , \ram[5][191] , \ram[5][190] , \ram[5][189] ,
         \ram[5][188] , \ram[5][187] , \ram[5][186] , \ram[5][185] ,
         \ram[5][184] , \ram[5][183] , \ram[5][182] , \ram[5][181] ,
         \ram[5][180] , \ram[5][179] , \ram[5][178] , \ram[5][177] ,
         \ram[5][176] , \ram[5][175] , \ram[5][174] , \ram[5][173] ,
         \ram[5][172] , \ram[5][171] , \ram[5][170] , \ram[5][169] ,
         \ram[5][168] , \ram[5][167] , \ram[5][166] , \ram[5][165] ,
         \ram[5][164] , \ram[5][163] , \ram[5][162] , \ram[5][161] ,
         \ram[5][160] , \ram[5][159] , \ram[5][158] , \ram[5][157] ,
         \ram[5][156] , \ram[5][155] , \ram[5][154] , \ram[5][153] ,
         \ram[5][152] , \ram[5][151] , \ram[5][150] , \ram[5][149] ,
         \ram[5][148] , \ram[5][147] , \ram[5][146] , \ram[5][145] ,
         \ram[5][144] , \ram[5][143] , \ram[5][142] , \ram[5][141] ,
         \ram[5][140] , \ram[5][139] , \ram[5][138] , \ram[5][137] ,
         \ram[5][136] , \ram[5][135] , \ram[5][134] , \ram[5][133] ,
         \ram[5][132] , \ram[5][131] , \ram[5][130] , \ram[5][129] ,
         \ram[5][128] , \ram[5][127] , \ram[5][126] , \ram[5][125] ,
         \ram[5][124] , \ram[5][123] , \ram[5][122] , \ram[5][121] ,
         \ram[5][120] , \ram[5][119] , \ram[5][118] , \ram[5][117] ,
         \ram[5][116] , \ram[5][115] , \ram[5][114] , \ram[5][113] ,
         \ram[5][112] , \ram[5][111] , \ram[5][110] , \ram[5][109] ,
         \ram[5][108] , \ram[5][107] , \ram[5][106] , \ram[5][105] ,
         \ram[5][104] , \ram[5][103] , \ram[5][102] , \ram[5][101] ,
         \ram[5][100] , \ram[5][99] , \ram[5][98] , \ram[5][97] , \ram[5][96] ,
         \ram[5][95] , \ram[5][94] , \ram[5][93] , \ram[5][92] , \ram[5][91] ,
         \ram[5][90] , \ram[5][89] , \ram[5][88] , \ram[5][87] , \ram[5][86] ,
         \ram[5][85] , \ram[5][84] , \ram[5][83] , \ram[5][82] , \ram[5][81] ,
         \ram[5][80] , \ram[5][79] , \ram[5][78] , \ram[5][77] , \ram[5][76] ,
         \ram[5][75] , \ram[5][74] , \ram[5][73] , \ram[5][72] , \ram[5][71] ,
         \ram[5][70] , \ram[5][69] , \ram[5][68] , \ram[5][67] , \ram[5][66] ,
         \ram[5][65] , \ram[5][64] , \ram[5][63] , \ram[5][62] , \ram[5][61] ,
         \ram[5][60] , \ram[5][59] , \ram[5][58] , \ram[5][57] , \ram[5][56] ,
         \ram[5][55] , \ram[5][54] , \ram[5][53] , \ram[5][52] , \ram[5][51] ,
         \ram[5][50] , \ram[5][49] , \ram[5][48] , \ram[5][47] , \ram[5][46] ,
         \ram[5][45] , \ram[5][44] , \ram[5][43] , \ram[5][42] , \ram[5][41] ,
         \ram[5][40] , \ram[5][39] , \ram[5][38] , \ram[5][37] , \ram[5][36] ,
         \ram[5][35] , \ram[5][34] , \ram[5][33] , \ram[5][32] , \ram[5][31] ,
         \ram[5][30] , \ram[5][29] , \ram[5][28] , \ram[5][27] , \ram[5][26] ,
         \ram[5][25] , \ram[5][24] , \ram[5][23] , \ram[5][22] , \ram[5][21] ,
         \ram[5][20] , \ram[5][19] , \ram[5][18] , \ram[5][17] , \ram[5][16] ,
         \ram[5][15] , \ram[5][14] , \ram[5][13] , \ram[5][12] , \ram[5][11] ,
         \ram[5][10] , \ram[5][9] , \ram[5][8] , \ram[5][7] , \ram[5][6] ,
         \ram[5][5] , \ram[5][4] , \ram[5][3] , \ram[5][2] , \ram[5][1] ,
         \ram[5][0] , \ram[4][255] , \ram[4][254] , \ram[4][253] ,
         \ram[4][252] , \ram[4][251] , \ram[4][250] , \ram[4][249] ,
         \ram[4][248] , \ram[4][247] , \ram[4][246] , \ram[4][245] ,
         \ram[4][244] , \ram[4][243] , \ram[4][242] , \ram[4][241] ,
         \ram[4][240] , \ram[4][239] , \ram[4][238] , \ram[4][237] ,
         \ram[4][236] , \ram[4][235] , \ram[4][234] , \ram[4][233] ,
         \ram[4][232] , \ram[4][231] , \ram[4][230] , \ram[4][229] ,
         \ram[4][228] , \ram[4][227] , \ram[4][226] , \ram[4][225] ,
         \ram[4][224] , \ram[4][223] , \ram[4][222] , \ram[4][221] ,
         \ram[4][220] , \ram[4][219] , \ram[4][218] , \ram[4][217] ,
         \ram[4][216] , \ram[4][215] , \ram[4][214] , \ram[4][213] ,
         \ram[4][212] , \ram[4][211] , \ram[4][210] , \ram[4][209] ,
         \ram[4][208] , \ram[4][207] , \ram[4][206] , \ram[4][205] ,
         \ram[4][204] , \ram[4][203] , \ram[4][202] , \ram[4][201] ,
         \ram[4][200] , \ram[4][199] , \ram[4][198] , \ram[4][197] ,
         \ram[4][196] , \ram[4][195] , \ram[4][194] , \ram[4][193] ,
         \ram[4][192] , \ram[4][191] , \ram[4][190] , \ram[4][189] ,
         \ram[4][188] , \ram[4][187] , \ram[4][186] , \ram[4][185] ,
         \ram[4][184] , \ram[4][183] , \ram[4][182] , \ram[4][181] ,
         \ram[4][180] , \ram[4][179] , \ram[4][178] , \ram[4][177] ,
         \ram[4][176] , \ram[4][175] , \ram[4][174] , \ram[4][173] ,
         \ram[4][172] , \ram[4][171] , \ram[4][170] , \ram[4][169] ,
         \ram[4][168] , \ram[4][167] , \ram[4][166] , \ram[4][165] ,
         \ram[4][164] , \ram[4][163] , \ram[4][162] , \ram[4][161] ,
         \ram[4][160] , \ram[4][159] , \ram[4][158] , \ram[4][157] ,
         \ram[4][156] , \ram[4][155] , \ram[4][154] , \ram[4][153] ,
         \ram[4][152] , \ram[4][151] , \ram[4][150] , \ram[4][149] ,
         \ram[4][148] , \ram[4][147] , \ram[4][146] , \ram[4][145] ,
         \ram[4][144] , \ram[4][143] , \ram[4][142] , \ram[4][141] ,
         \ram[4][140] , \ram[4][139] , \ram[4][138] , \ram[4][137] ,
         \ram[4][136] , \ram[4][135] , \ram[4][134] , \ram[4][133] ,
         \ram[4][132] , \ram[4][131] , \ram[4][130] , \ram[4][129] ,
         \ram[4][128] , \ram[4][127] , \ram[4][126] , \ram[4][125] ,
         \ram[4][124] , \ram[4][123] , \ram[4][122] , \ram[4][121] ,
         \ram[4][120] , \ram[4][119] , \ram[4][118] , \ram[4][117] ,
         \ram[4][116] , \ram[4][115] , \ram[4][114] , \ram[4][113] ,
         \ram[4][112] , \ram[4][111] , \ram[4][110] , \ram[4][109] ,
         \ram[4][108] , \ram[4][107] , \ram[4][106] , \ram[4][105] ,
         \ram[4][104] , \ram[4][103] , \ram[4][102] , \ram[4][101] ,
         \ram[4][100] , \ram[4][99] , \ram[4][98] , \ram[4][97] , \ram[4][96] ,
         \ram[4][95] , \ram[4][94] , \ram[4][93] , \ram[4][92] , \ram[4][91] ,
         \ram[4][90] , \ram[4][89] , \ram[4][88] , \ram[4][87] , \ram[4][86] ,
         \ram[4][85] , \ram[4][84] , \ram[4][83] , \ram[4][82] , \ram[4][81] ,
         \ram[4][80] , \ram[4][79] , \ram[4][78] , \ram[4][77] , \ram[4][76] ,
         \ram[4][75] , \ram[4][74] , \ram[4][73] , \ram[4][72] , \ram[4][71] ,
         \ram[4][70] , \ram[4][69] , \ram[4][68] , \ram[4][67] , \ram[4][66] ,
         \ram[4][65] , \ram[4][64] , \ram[4][63] , \ram[4][62] , \ram[4][61] ,
         \ram[4][60] , \ram[4][59] , \ram[4][58] , \ram[4][57] , \ram[4][56] ,
         \ram[4][55] , \ram[4][54] , \ram[4][53] , \ram[4][52] , \ram[4][51] ,
         \ram[4][50] , \ram[4][49] , \ram[4][48] , \ram[4][47] , \ram[4][46] ,
         \ram[4][45] , \ram[4][44] , \ram[4][43] , \ram[4][42] , \ram[4][41] ,
         \ram[4][40] , \ram[4][39] , \ram[4][38] , \ram[4][37] , \ram[4][36] ,
         \ram[4][35] , \ram[4][34] , \ram[4][33] , \ram[4][32] , \ram[4][31] ,
         \ram[4][30] , \ram[4][29] , \ram[4][28] , \ram[4][27] , \ram[4][26] ,
         \ram[4][25] , \ram[4][24] , \ram[4][23] , \ram[4][22] , \ram[4][21] ,
         \ram[4][20] , \ram[4][19] , \ram[4][18] , \ram[4][17] , \ram[4][16] ,
         \ram[4][15] , \ram[4][14] , \ram[4][13] , \ram[4][12] , \ram[4][11] ,
         \ram[4][10] , \ram[4][9] , \ram[4][8] , \ram[4][7] , \ram[4][6] ,
         \ram[4][5] , \ram[4][4] , \ram[4][3] , \ram[4][2] , \ram[4][1] ,
         \ram[4][0] , \ram[3][255] , \ram[3][254] , \ram[3][253] ,
         \ram[3][252] , \ram[3][251] , \ram[3][250] , \ram[3][249] ,
         \ram[3][248] , \ram[3][247] , \ram[3][246] , \ram[3][245] ,
         \ram[3][244] , \ram[3][243] , \ram[3][242] , \ram[3][241] ,
         \ram[3][240] , \ram[3][239] , \ram[3][238] , \ram[3][237] ,
         \ram[3][236] , \ram[3][235] , \ram[3][234] , \ram[3][233] ,
         \ram[3][232] , \ram[3][231] , \ram[3][230] , \ram[3][229] ,
         \ram[3][228] , \ram[3][227] , \ram[3][226] , \ram[3][225] ,
         \ram[3][224] , \ram[3][223] , \ram[3][222] , \ram[3][221] ,
         \ram[3][220] , \ram[3][219] , \ram[3][218] , \ram[3][217] ,
         \ram[3][216] , \ram[3][215] , \ram[3][214] , \ram[3][213] ,
         \ram[3][212] , \ram[3][211] , \ram[3][210] , \ram[3][209] ,
         \ram[3][208] , \ram[3][207] , \ram[3][206] , \ram[3][205] ,
         \ram[3][204] , \ram[3][203] , \ram[3][202] , \ram[3][201] ,
         \ram[3][200] , \ram[3][199] , \ram[3][198] , \ram[3][197] ,
         \ram[3][196] , \ram[3][195] , \ram[3][194] , \ram[3][193] ,
         \ram[3][192] , \ram[3][191] , \ram[3][190] , \ram[3][189] ,
         \ram[3][188] , \ram[3][187] , \ram[3][186] , \ram[3][185] ,
         \ram[3][184] , \ram[3][183] , \ram[3][182] , \ram[3][181] ,
         \ram[3][180] , \ram[3][179] , \ram[3][178] , \ram[3][177] ,
         \ram[3][176] , \ram[3][175] , \ram[3][174] , \ram[3][173] ,
         \ram[3][172] , \ram[3][171] , \ram[3][170] , \ram[3][169] ,
         \ram[3][168] , \ram[3][167] , \ram[3][166] , \ram[3][165] ,
         \ram[3][164] , \ram[3][163] , \ram[3][162] , \ram[3][161] ,
         \ram[3][160] , \ram[3][159] , \ram[3][158] , \ram[3][157] ,
         \ram[3][156] , \ram[3][155] , \ram[3][154] , \ram[3][153] ,
         \ram[3][152] , \ram[3][151] , \ram[3][150] , \ram[3][149] ,
         \ram[3][148] , \ram[3][147] , \ram[3][146] , \ram[3][145] ,
         \ram[3][144] , \ram[3][143] , \ram[3][142] , \ram[3][141] ,
         \ram[3][140] , \ram[3][139] , \ram[3][138] , \ram[3][137] ,
         \ram[3][136] , \ram[3][135] , \ram[3][134] , \ram[3][133] ,
         \ram[3][132] , \ram[3][131] , \ram[3][130] , \ram[3][129] ,
         \ram[3][128] , \ram[3][127] , \ram[3][126] , \ram[3][125] ,
         \ram[3][124] , \ram[3][123] , \ram[3][122] , \ram[3][121] ,
         \ram[3][120] , \ram[3][119] , \ram[3][118] , \ram[3][117] ,
         \ram[3][116] , \ram[3][115] , \ram[3][114] , \ram[3][113] ,
         \ram[3][112] , \ram[3][111] , \ram[3][110] , \ram[3][109] ,
         \ram[3][108] , \ram[3][107] , \ram[3][106] , \ram[3][105] ,
         \ram[3][104] , \ram[3][103] , \ram[3][102] , \ram[3][101] ,
         \ram[3][100] , \ram[3][99] , \ram[3][98] , \ram[3][97] , \ram[3][96] ,
         \ram[3][95] , \ram[3][94] , \ram[3][93] , \ram[3][92] , \ram[3][91] ,
         \ram[3][90] , \ram[3][89] , \ram[3][88] , \ram[3][87] , \ram[3][86] ,
         \ram[3][85] , \ram[3][84] , \ram[3][83] , \ram[3][82] , \ram[3][81] ,
         \ram[3][80] , \ram[3][79] , \ram[3][78] , \ram[3][77] , \ram[3][76] ,
         \ram[3][75] , \ram[3][74] , \ram[3][73] , \ram[3][72] , \ram[3][71] ,
         \ram[3][70] , \ram[3][69] , \ram[3][68] , \ram[3][67] , \ram[3][66] ,
         \ram[3][65] , \ram[3][64] , \ram[3][63] , \ram[3][62] , \ram[3][61] ,
         \ram[3][60] , \ram[3][59] , \ram[3][58] , \ram[3][57] , \ram[3][56] ,
         \ram[3][55] , \ram[3][54] , \ram[3][53] , \ram[3][52] , \ram[3][51] ,
         \ram[3][50] , \ram[3][49] , \ram[3][48] , \ram[3][47] , \ram[3][46] ,
         \ram[3][45] , \ram[3][44] , \ram[3][43] , \ram[3][42] , \ram[3][41] ,
         \ram[3][40] , \ram[3][39] , \ram[3][38] , \ram[3][37] , \ram[3][36] ,
         \ram[3][35] , \ram[3][34] , \ram[3][33] , \ram[3][32] , \ram[3][31] ,
         \ram[3][30] , \ram[3][29] , \ram[3][28] , \ram[3][27] , \ram[3][26] ,
         \ram[3][25] , \ram[3][24] , \ram[3][23] , \ram[3][22] , \ram[3][21] ,
         \ram[3][20] , \ram[3][19] , \ram[3][18] , \ram[3][17] , \ram[3][16] ,
         \ram[3][15] , \ram[3][14] , \ram[3][13] , \ram[3][12] , \ram[3][11] ,
         \ram[3][10] , \ram[3][9] , \ram[3][8] , \ram[3][7] , \ram[3][6] ,
         \ram[3][5] , \ram[3][4] , \ram[3][3] , \ram[3][2] , \ram[3][1] ,
         \ram[3][0] , \ram[2][255] , \ram[2][254] , \ram[2][253] ,
         \ram[2][252] , \ram[2][251] , \ram[2][250] , \ram[2][249] ,
         \ram[2][248] , \ram[2][247] , \ram[2][246] , \ram[2][245] ,
         \ram[2][244] , \ram[2][243] , \ram[2][242] , \ram[2][241] ,
         \ram[2][240] , \ram[2][239] , \ram[2][238] , \ram[2][237] ,
         \ram[2][236] , \ram[2][235] , \ram[2][234] , \ram[2][233] ,
         \ram[2][232] , \ram[2][231] , \ram[2][230] , \ram[2][229] ,
         \ram[2][228] , \ram[2][227] , \ram[2][226] , \ram[2][225] ,
         \ram[2][224] , \ram[2][223] , \ram[2][222] , \ram[2][221] ,
         \ram[2][220] , \ram[2][219] , \ram[2][218] , \ram[2][217] ,
         \ram[2][216] , \ram[2][215] , \ram[2][214] , \ram[2][213] ,
         \ram[2][212] , \ram[2][211] , \ram[2][210] , \ram[2][209] ,
         \ram[2][208] , \ram[2][207] , \ram[2][206] , \ram[2][205] ,
         \ram[2][204] , \ram[2][203] , \ram[2][202] , \ram[2][201] ,
         \ram[2][200] , \ram[2][199] , \ram[2][198] , \ram[2][197] ,
         \ram[2][196] , \ram[2][195] , \ram[2][194] , \ram[2][193] ,
         \ram[2][192] , \ram[2][191] , \ram[2][190] , \ram[2][189] ,
         \ram[2][188] , \ram[2][187] , \ram[2][186] , \ram[2][185] ,
         \ram[2][184] , \ram[2][183] , \ram[2][182] , \ram[2][181] ,
         \ram[2][180] , \ram[2][179] , \ram[2][178] , \ram[2][177] ,
         \ram[2][176] , \ram[2][175] , \ram[2][174] , \ram[2][173] ,
         \ram[2][172] , \ram[2][171] , \ram[2][170] , \ram[2][169] ,
         \ram[2][168] , \ram[2][167] , \ram[2][166] , \ram[2][165] ,
         \ram[2][164] , \ram[2][163] , \ram[2][162] , \ram[2][161] ,
         \ram[2][160] , \ram[2][159] , \ram[2][158] , \ram[2][157] ,
         \ram[2][156] , \ram[2][155] , \ram[2][154] , \ram[2][153] ,
         \ram[2][152] , \ram[2][151] , \ram[2][150] , \ram[2][149] ,
         \ram[2][148] , \ram[2][147] , \ram[2][146] , \ram[2][145] ,
         \ram[2][144] , \ram[2][143] , \ram[2][142] , \ram[2][141] ,
         \ram[2][140] , \ram[2][139] , \ram[2][138] , \ram[2][137] ,
         \ram[2][136] , \ram[2][135] , \ram[2][134] , \ram[2][133] ,
         \ram[2][132] , \ram[2][131] , \ram[2][130] , \ram[2][129] ,
         \ram[2][128] , \ram[2][127] , \ram[2][126] , \ram[2][125] ,
         \ram[2][124] , \ram[2][123] , \ram[2][122] , \ram[2][121] ,
         \ram[2][120] , \ram[2][119] , \ram[2][118] , \ram[2][117] ,
         \ram[2][116] , \ram[2][115] , \ram[2][114] , \ram[2][113] ,
         \ram[2][112] , \ram[2][111] , \ram[2][110] , \ram[2][109] ,
         \ram[2][108] , \ram[2][107] , \ram[2][106] , \ram[2][105] ,
         \ram[2][104] , \ram[2][103] , \ram[2][102] , \ram[2][101] ,
         \ram[2][100] , \ram[2][99] , \ram[2][98] , \ram[2][97] , \ram[2][96] ,
         \ram[2][95] , \ram[2][94] , \ram[2][93] , \ram[2][92] , \ram[2][91] ,
         \ram[2][90] , \ram[2][89] , \ram[2][88] , \ram[2][87] , \ram[2][86] ,
         \ram[2][85] , \ram[2][84] , \ram[2][83] , \ram[2][82] , \ram[2][81] ,
         \ram[2][80] , \ram[2][79] , \ram[2][78] , \ram[2][77] , \ram[2][76] ,
         \ram[2][75] , \ram[2][74] , \ram[2][73] , \ram[2][72] , \ram[2][71] ,
         \ram[2][70] , \ram[2][69] , \ram[2][68] , \ram[2][67] , \ram[2][66] ,
         \ram[2][65] , \ram[2][64] , \ram[2][63] , \ram[2][62] , \ram[2][61] ,
         \ram[2][60] , \ram[2][59] , \ram[2][58] , \ram[2][57] , \ram[2][56] ,
         \ram[2][55] , \ram[2][54] , \ram[2][53] , \ram[2][52] , \ram[2][51] ,
         \ram[2][50] , \ram[2][49] , \ram[2][48] , \ram[2][47] , \ram[2][46] ,
         \ram[2][45] , \ram[2][44] , \ram[2][43] , \ram[2][42] , \ram[2][41] ,
         \ram[2][40] , \ram[2][39] , \ram[2][38] , \ram[2][37] , \ram[2][36] ,
         \ram[2][35] , \ram[2][34] , \ram[2][33] , \ram[2][32] , \ram[2][31] ,
         \ram[2][30] , \ram[2][29] , \ram[2][28] , \ram[2][27] , \ram[2][26] ,
         \ram[2][25] , \ram[2][24] , \ram[2][23] , \ram[2][22] , \ram[2][21] ,
         \ram[2][20] , \ram[2][19] , \ram[2][18] , \ram[2][17] , \ram[2][16] ,
         \ram[2][15] , \ram[2][14] , \ram[2][13] , \ram[2][12] , \ram[2][11] ,
         \ram[2][10] , \ram[2][9] , \ram[2][8] , \ram[2][7] , \ram[2][6] ,
         \ram[2][5] , \ram[2][4] , \ram[2][3] , \ram[2][2] , \ram[2][1] ,
         \ram[2][0] , \ram[1][255] , \ram[1][254] , \ram[1][253] ,
         \ram[1][252] , \ram[1][251] , \ram[1][250] , \ram[1][249] ,
         \ram[1][248] , \ram[1][247] , \ram[1][246] , \ram[1][245] ,
         \ram[1][244] , \ram[1][243] , \ram[1][242] , \ram[1][241] ,
         \ram[1][240] , \ram[1][239] , \ram[1][238] , \ram[1][237] ,
         \ram[1][236] , \ram[1][235] , \ram[1][234] , \ram[1][233] ,
         \ram[1][232] , \ram[1][231] , \ram[1][230] , \ram[1][229] ,
         \ram[1][228] , \ram[1][227] , \ram[1][226] , \ram[1][225] ,
         \ram[1][224] , \ram[1][223] , \ram[1][222] , \ram[1][221] ,
         \ram[1][220] , \ram[1][219] , \ram[1][218] , \ram[1][217] ,
         \ram[1][216] , \ram[1][215] , \ram[1][214] , \ram[1][213] ,
         \ram[1][212] , \ram[1][211] , \ram[1][210] , \ram[1][209] ,
         \ram[1][208] , \ram[1][207] , \ram[1][206] , \ram[1][205] ,
         \ram[1][204] , \ram[1][203] , \ram[1][202] , \ram[1][201] ,
         \ram[1][200] , \ram[1][199] , \ram[1][198] , \ram[1][197] ,
         \ram[1][196] , \ram[1][195] , \ram[1][194] , \ram[1][193] ,
         \ram[1][192] , \ram[1][191] , \ram[1][190] , \ram[1][189] ,
         \ram[1][188] , \ram[1][187] , \ram[1][186] , \ram[1][185] ,
         \ram[1][184] , \ram[1][183] , \ram[1][182] , \ram[1][181] ,
         \ram[1][180] , \ram[1][179] , \ram[1][178] , \ram[1][177] ,
         \ram[1][176] , \ram[1][175] , \ram[1][174] , \ram[1][173] ,
         \ram[1][172] , \ram[1][171] , \ram[1][170] , \ram[1][169] ,
         \ram[1][168] , \ram[1][167] , \ram[1][166] , \ram[1][165] ,
         \ram[1][164] , \ram[1][163] , \ram[1][162] , \ram[1][161] ,
         \ram[1][160] , \ram[1][159] , \ram[1][158] , \ram[1][157] ,
         \ram[1][156] , \ram[1][155] , \ram[1][154] , \ram[1][153] ,
         \ram[1][152] , \ram[1][151] , \ram[1][150] , \ram[1][149] ,
         \ram[1][148] , \ram[1][147] , \ram[1][146] , \ram[1][145] ,
         \ram[1][144] , \ram[1][143] , \ram[1][142] , \ram[1][141] ,
         \ram[1][140] , \ram[1][139] , \ram[1][138] , \ram[1][137] ,
         \ram[1][136] , \ram[1][135] , \ram[1][134] , \ram[1][133] ,
         \ram[1][132] , \ram[1][131] , \ram[1][130] , \ram[1][129] ,
         \ram[1][128] , \ram[1][127] , \ram[1][126] , \ram[1][125] ,
         \ram[1][124] , \ram[1][123] , \ram[1][122] , \ram[1][121] ,
         \ram[1][120] , \ram[1][119] , \ram[1][118] , \ram[1][117] ,
         \ram[1][116] , \ram[1][115] , \ram[1][114] , \ram[1][113] ,
         \ram[1][112] , \ram[1][111] , \ram[1][110] , \ram[1][109] ,
         \ram[1][108] , \ram[1][107] , \ram[1][106] , \ram[1][105] ,
         \ram[1][104] , \ram[1][103] , \ram[1][102] , \ram[1][101] ,
         \ram[1][100] , \ram[1][99] , \ram[1][98] , \ram[1][97] , \ram[1][96] ,
         \ram[1][95] , \ram[1][94] , \ram[1][93] , \ram[1][92] , \ram[1][91] ,
         \ram[1][90] , \ram[1][89] , \ram[1][88] , \ram[1][87] , \ram[1][86] ,
         \ram[1][85] , \ram[1][84] , \ram[1][83] , \ram[1][82] , \ram[1][81] ,
         \ram[1][80] , \ram[1][79] , \ram[1][78] , \ram[1][77] , \ram[1][76] ,
         \ram[1][75] , \ram[1][74] , \ram[1][73] , \ram[1][72] , \ram[1][71] ,
         \ram[1][70] , \ram[1][69] , \ram[1][68] , \ram[1][67] , \ram[1][66] ,
         \ram[1][65] , \ram[1][64] , \ram[1][63] , \ram[1][62] , \ram[1][61] ,
         \ram[1][60] , \ram[1][59] , \ram[1][58] , \ram[1][57] , \ram[1][56] ,
         \ram[1][55] , \ram[1][54] , \ram[1][53] , \ram[1][52] , \ram[1][51] ,
         \ram[1][50] , \ram[1][49] , \ram[1][48] , \ram[1][47] , \ram[1][46] ,
         \ram[1][45] , \ram[1][44] , \ram[1][43] , \ram[1][42] , \ram[1][41] ,
         \ram[1][40] , \ram[1][39] , \ram[1][38] , \ram[1][37] , \ram[1][36] ,
         \ram[1][35] , \ram[1][34] , \ram[1][33] , \ram[1][32] , \ram[1][31] ,
         \ram[1][30] , \ram[1][29] , \ram[1][28] , \ram[1][27] , \ram[1][26] ,
         \ram[1][25] , \ram[1][24] , \ram[1][23] , \ram[1][22] , \ram[1][21] ,
         \ram[1][20] , \ram[1][19] , \ram[1][18] , \ram[1][17] , \ram[1][16] ,
         \ram[1][15] , \ram[1][14] , \ram[1][13] , \ram[1][12] , \ram[1][11] ,
         \ram[1][10] , \ram[1][9] , \ram[1][8] , \ram[1][7] , \ram[1][6] ,
         \ram[1][5] , \ram[1][4] , \ram[1][3] , \ram[1][2] , \ram[1][1] ,
         \ram[1][0] , \ram[0][255] , \ram[0][254] , \ram[0][253] ,
         \ram[0][252] , \ram[0][251] , \ram[0][250] , \ram[0][249] ,
         \ram[0][248] , \ram[0][247] , \ram[0][246] , \ram[0][245] ,
         \ram[0][244] , \ram[0][243] , \ram[0][242] , \ram[0][241] ,
         \ram[0][240] , \ram[0][239] , \ram[0][238] , \ram[0][237] ,
         \ram[0][236] , \ram[0][235] , \ram[0][234] , \ram[0][233] ,
         \ram[0][232] , \ram[0][231] , \ram[0][230] , \ram[0][229] ,
         \ram[0][228] , \ram[0][227] , \ram[0][226] , \ram[0][225] ,
         \ram[0][224] , \ram[0][223] , \ram[0][222] , \ram[0][221] ,
         \ram[0][220] , \ram[0][219] , \ram[0][218] , \ram[0][217] ,
         \ram[0][216] , \ram[0][215] , \ram[0][214] , \ram[0][213] ,
         \ram[0][212] , \ram[0][211] , \ram[0][210] , \ram[0][209] ,
         \ram[0][208] , \ram[0][207] , \ram[0][206] , \ram[0][205] ,
         \ram[0][204] , \ram[0][203] , \ram[0][202] , \ram[0][201] ,
         \ram[0][200] , \ram[0][199] , \ram[0][198] , \ram[0][197] ,
         \ram[0][196] , \ram[0][195] , \ram[0][194] , \ram[0][193] ,
         \ram[0][192] , \ram[0][191] , \ram[0][190] , \ram[0][189] ,
         \ram[0][188] , \ram[0][187] , \ram[0][186] , \ram[0][185] ,
         \ram[0][184] , \ram[0][183] , \ram[0][182] , \ram[0][181] ,
         \ram[0][180] , \ram[0][179] , \ram[0][178] , \ram[0][177] ,
         \ram[0][176] , \ram[0][175] , \ram[0][174] , \ram[0][173] ,
         \ram[0][172] , \ram[0][171] , \ram[0][170] , \ram[0][169] ,
         \ram[0][168] , \ram[0][167] , \ram[0][166] , \ram[0][165] ,
         \ram[0][164] , \ram[0][163] , \ram[0][162] , \ram[0][161] ,
         \ram[0][160] , \ram[0][159] , \ram[0][158] , \ram[0][157] ,
         \ram[0][156] , \ram[0][155] , \ram[0][154] , \ram[0][153] ,
         \ram[0][152] , \ram[0][151] , \ram[0][150] , \ram[0][149] ,
         \ram[0][148] , \ram[0][147] , \ram[0][146] , \ram[0][145] ,
         \ram[0][144] , \ram[0][143] , \ram[0][142] , \ram[0][141] ,
         \ram[0][140] , \ram[0][139] , \ram[0][138] , \ram[0][137] ,
         \ram[0][136] , \ram[0][135] , \ram[0][134] , \ram[0][133] ,
         \ram[0][132] , \ram[0][131] , \ram[0][130] , \ram[0][129] ,
         \ram[0][128] , \ram[0][127] , \ram[0][126] , \ram[0][125] ,
         \ram[0][124] , \ram[0][123] , \ram[0][122] , \ram[0][121] ,
         \ram[0][120] , \ram[0][119] , \ram[0][118] , \ram[0][117] ,
         \ram[0][116] , \ram[0][115] , \ram[0][114] , \ram[0][113] ,
         \ram[0][112] , \ram[0][111] , \ram[0][110] , \ram[0][109] ,
         \ram[0][108] , \ram[0][107] , \ram[0][106] , \ram[0][105] ,
         \ram[0][104] , \ram[0][103] , \ram[0][102] , \ram[0][101] ,
         \ram[0][100] , \ram[0][99] , \ram[0][98] , \ram[0][97] , \ram[0][96] ,
         \ram[0][95] , \ram[0][94] , \ram[0][93] , \ram[0][92] , \ram[0][91] ,
         \ram[0][90] , \ram[0][89] , \ram[0][88] , \ram[0][87] , \ram[0][86] ,
         \ram[0][85] , \ram[0][84] , \ram[0][83] , \ram[0][82] , \ram[0][81] ,
         \ram[0][80] , \ram[0][79] , \ram[0][78] , \ram[0][77] , \ram[0][76] ,
         \ram[0][75] , \ram[0][74] , \ram[0][73] , \ram[0][72] , \ram[0][71] ,
         \ram[0][70] , \ram[0][69] , \ram[0][68] , \ram[0][67] , \ram[0][66] ,
         \ram[0][65] , \ram[0][64] , \ram[0][63] , \ram[0][62] , \ram[0][61] ,
         \ram[0][60] , \ram[0][59] , \ram[0][58] , \ram[0][57] , \ram[0][56] ,
         \ram[0][55] , \ram[0][54] , \ram[0][53] , \ram[0][52] , \ram[0][51] ,
         \ram[0][50] , \ram[0][49] , \ram[0][48] , \ram[0][47] , \ram[0][46] ,
         \ram[0][45] , \ram[0][44] , \ram[0][43] , \ram[0][42] , \ram[0][41] ,
         \ram[0][40] , \ram[0][39] , \ram[0][38] , \ram[0][37] , \ram[0][36] ,
         \ram[0][35] , \ram[0][34] , \ram[0][33] , \ram[0][32] , \ram[0][31] ,
         \ram[0][30] , \ram[0][29] , \ram[0][28] , \ram[0][27] , \ram[0][26] ,
         \ram[0][25] , \ram[0][24] , \ram[0][23] , \ram[0][22] , \ram[0][21] ,
         \ram[0][20] , \ram[0][19] , \ram[0][18] , \ram[0][17] , \ram[0][16] ,
         \ram[0][15] , \ram[0][14] , \ram[0][13] , \ram[0][12] , \ram[0][11] ,
         \ram[0][10] , \ram[0][9] , \ram[0][8] , \ram[0][7] , \ram[0][6] ,
         \ram[0][5] , \ram[0][4] , \ram[0][3] , \ram[0][2] , \ram[0][1] ,
         \ram[0][0] , N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96,
         N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108,
         N109, N110, N111, N112, N113, N114, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175,
         N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N276,
         N279, N282, N285, N288, N291, N294, N297, N300, N303, N306, N309,
         N312, N315, N318, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640;
  assign N9 = addr[0];
  assign N10 = addr[1];
  assign N11 = addr[2];
  assign N12 = addr[3];

  LATCHX1_HVT \ram_reg[15][255]  ( .CLK(N318), .D(N273), .Q(\ram[15][255] ) );
  LATCHX1_HVT \ram_reg[15][254]  ( .CLK(N318), .D(N272), .Q(\ram[15][254] ) );
  LATCHX1_HVT \ram_reg[15][253]  ( .CLK(N318), .D(N271), .Q(\ram[15][253] ) );
  LATCHX1_HVT \ram_reg[15][252]  ( .CLK(N318), .D(N270), .Q(\ram[15][252] ) );
  LATCHX1_HVT \ram_reg[15][251]  ( .CLK(n21), .D(N269), .Q(\ram[15][251] ) );
  LATCHX1_HVT \ram_reg[15][250]  ( .CLK(n13), .D(N268), .Q(\ram[15][250] ) );
  LATCHX1_HVT \ram_reg[15][249]  ( .CLK(n13), .D(N267), .Q(\ram[15][249] ) );
  LATCHX1_HVT \ram_reg[15][248]  ( .CLK(n13), .D(N266), .Q(\ram[15][248] ) );
  LATCHX1_HVT \ram_reg[15][247]  ( .CLK(n13), .D(N265), .Q(\ram[15][247] ) );
  LATCHX1_HVT \ram_reg[15][246]  ( .CLK(n13), .D(N264), .Q(\ram[15][246] ) );
  LATCHX1_HVT \ram_reg[15][245]  ( .CLK(n13), .D(N263), .Q(\ram[15][245] ) );
  LATCHX1_HVT \ram_reg[15][244]  ( .CLK(n13), .D(N262), .Q(\ram[15][244] ) );
  LATCHX1_HVT \ram_reg[15][243]  ( .CLK(n13), .D(N261), .Q(\ram[15][243] ) );
  LATCHX1_HVT \ram_reg[15][242]  ( .CLK(n13), .D(N260), .Q(\ram[15][242] ) );
  LATCHX1_HVT \ram_reg[15][241]  ( .CLK(n12), .D(N259), .Q(\ram[15][241] ) );
  LATCHX1_HVT \ram_reg[15][240]  ( .CLK(n12), .D(N258), .Q(\ram[15][240] ) );
  LATCHX1_HVT \ram_reg[15][239]  ( .CLK(n12), .D(N257), .Q(\ram[15][239] ) );
  LATCHX1_HVT \ram_reg[15][238]  ( .CLK(n12), .D(N256), .Q(\ram[15][238] ) );
  LATCHX1_HVT \ram_reg[15][237]  ( .CLK(n12), .D(N255), .Q(\ram[15][237] ) );
  LATCHX1_HVT \ram_reg[15][236]  ( .CLK(n12), .D(N254), .Q(\ram[15][236] ) );
  LATCHX1_HVT \ram_reg[15][235]  ( .CLK(n12), .D(N253), .Q(\ram[15][235] ) );
  LATCHX1_HVT \ram_reg[15][234]  ( .CLK(n12), .D(N252), .Q(\ram[15][234] ) );
  LATCHX1_HVT \ram_reg[15][233]  ( .CLK(n12), .D(N251), .Q(\ram[15][233] ) );
  LATCHX1_HVT \ram_reg[15][232]  ( .CLK(n12), .D(N250), .Q(\ram[15][232] ) );
  LATCHX1_HVT \ram_reg[15][231]  ( .CLK(n12), .D(N249), .Q(\ram[15][231] ) );
  LATCHX1_HVT \ram_reg[15][230]  ( .CLK(n11), .D(N248), .Q(\ram[15][230] ) );
  LATCHX1_HVT \ram_reg[15][229]  ( .CLK(n11), .D(N247), .Q(\ram[15][229] ) );
  LATCHX1_HVT \ram_reg[15][228]  ( .CLK(n11), .D(N246), .Q(\ram[15][228] ) );
  LATCHX1_HVT \ram_reg[15][227]  ( .CLK(n21), .D(N245), .Q(\ram[15][227] ) );
  LATCHX1_HVT \ram_reg[15][226]  ( .CLK(n21), .D(N244), .Q(\ram[15][226] ) );
  LATCHX1_HVT \ram_reg[15][225]  ( .CLK(n21), .D(N243), .Q(\ram[15][225] ) );
  LATCHX1_HVT \ram_reg[15][224]  ( .CLK(n21), .D(N242), .Q(\ram[15][224] ) );
  LATCHX1_HVT \ram_reg[15][223]  ( .CLK(n21), .D(N241), .Q(\ram[15][223] ) );
  LATCHX1_HVT \ram_reg[15][222]  ( .CLK(n21), .D(N240), .Q(\ram[15][222] ) );
  LATCHX1_HVT \ram_reg[15][221]  ( .CLK(n21), .D(N239), .Q(\ram[15][221] ) );
  LATCHX1_HVT \ram_reg[15][220]  ( .CLK(n21), .D(N238), .Q(\ram[15][220] ) );
  LATCHX1_HVT \ram_reg[15][219]  ( .CLK(n21), .D(N237), .Q(\ram[15][219] ) );
  LATCHX1_HVT \ram_reg[15][218]  ( .CLK(n21), .D(N236), .Q(\ram[15][218] ) );
  LATCHX1_HVT \ram_reg[15][217]  ( .CLK(n20), .D(N235), .Q(\ram[15][217] ) );
  LATCHX1_HVT \ram_reg[15][216]  ( .CLK(n20), .D(N234), .Q(\ram[15][216] ) );
  LATCHX1_HVT \ram_reg[15][215]  ( .CLK(n20), .D(N233), .Q(\ram[15][215] ) );
  LATCHX1_HVT \ram_reg[15][214]  ( .CLK(n20), .D(N232), .Q(\ram[15][214] ) );
  LATCHX1_HVT \ram_reg[15][213]  ( .CLK(n20), .D(N231), .Q(\ram[15][213] ) );
  LATCHX1_HVT \ram_reg[15][212]  ( .CLK(n20), .D(N230), .Q(\ram[15][212] ) );
  LATCHX1_HVT \ram_reg[15][211]  ( .CLK(n20), .D(N229), .Q(\ram[15][211] ) );
  LATCHX1_HVT \ram_reg[15][210]  ( .CLK(n20), .D(N228), .Q(\ram[15][210] ) );
  LATCHX1_HVT \ram_reg[15][209]  ( .CLK(n20), .D(N227), .Q(\ram[15][209] ) );
  LATCHX1_HVT \ram_reg[15][208]  ( .CLK(n20), .D(N226), .Q(\ram[15][208] ) );
  LATCHX1_HVT \ram_reg[15][207]  ( .CLK(n19), .D(N225), .Q(\ram[15][207] ) );
  LATCHX1_HVT \ram_reg[15][206]  ( .CLK(n19), .D(N224), .Q(\ram[15][206] ) );
  LATCHX1_HVT \ram_reg[15][205]  ( .CLK(n19), .D(N223), .Q(\ram[15][205] ) );
  LATCHX1_HVT \ram_reg[15][204]  ( .CLK(n19), .D(N222), .Q(\ram[15][204] ) );
  LATCHX1_HVT \ram_reg[15][203]  ( .CLK(n19), .D(N221), .Q(\ram[15][203] ) );
  LATCHX1_HVT \ram_reg[15][202]  ( .CLK(n19), .D(N220), .Q(\ram[15][202] ) );
  LATCHX1_HVT \ram_reg[15][201]  ( .CLK(n19), .D(N219), .Q(\ram[15][201] ) );
  LATCHX1_HVT \ram_reg[15][200]  ( .CLK(n19), .D(N218), .Q(\ram[15][200] ) );
  LATCHX1_HVT \ram_reg[15][199]  ( .CLK(n19), .D(N217), .Q(\ram[15][199] ) );
  LATCHX1_HVT \ram_reg[15][198]  ( .CLK(n19), .D(N216), .Q(\ram[15][198] ) );
  LATCHX1_HVT \ram_reg[15][197]  ( .CLK(n19), .D(N214), .Q(\ram[15][197] ) );
  LATCHX1_HVT \ram_reg[15][196]  ( .CLK(n18), .D(N213), .Q(\ram[15][196] ) );
  LATCHX1_HVT \ram_reg[15][195]  ( .CLK(n18), .D(N212), .Q(\ram[15][195] ) );
  LATCHX1_HVT \ram_reg[15][194]  ( .CLK(n18), .D(N211), .Q(\ram[15][194] ) );
  LATCHX1_HVT \ram_reg[15][193]  ( .CLK(n18), .D(N210), .Q(\ram[15][193] ) );
  LATCHX1_HVT \ram_reg[15][192]  ( .CLK(n18), .D(N209), .Q(\ram[15][192] ) );
  LATCHX1_HVT \ram_reg[15][191]  ( .CLK(n18), .D(N208), .Q(\ram[15][191] ) );
  LATCHX1_HVT \ram_reg[15][190]  ( .CLK(n18), .D(N207), .Q(\ram[15][190] ) );
  LATCHX1_HVT \ram_reg[15][189]  ( .CLK(n18), .D(N206), .Q(\ram[15][189] ) );
  LATCHX1_HVT \ram_reg[15][188]  ( .CLK(n18), .D(N205), .Q(\ram[15][188] ) );
  LATCHX1_HVT \ram_reg[15][187]  ( .CLK(n18), .D(N204), .Q(\ram[15][187] ) );
  LATCHX1_HVT \ram_reg[15][186]  ( .CLK(n18), .D(N203), .Q(\ram[15][186] ) );
  LATCHX1_HVT \ram_reg[15][185]  ( .CLK(n17), .D(N202), .Q(\ram[15][185] ) );
  LATCHX1_HVT \ram_reg[15][184]  ( .CLK(n17), .D(N201), .Q(\ram[15][184] ) );
  LATCHX1_HVT \ram_reg[15][183]  ( .CLK(n17), .D(N200), .Q(\ram[15][183] ) );
  LATCHX1_HVT \ram_reg[15][182]  ( .CLK(n17), .D(N199), .Q(\ram[15][182] ) );
  LATCHX1_HVT \ram_reg[15][181]  ( .CLK(n17), .D(N198), .Q(\ram[15][181] ) );
  LATCHX1_HVT \ram_reg[15][180]  ( .CLK(n17), .D(N197), .Q(\ram[15][180] ) );
  LATCHX1_HVT \ram_reg[15][179]  ( .CLK(n17), .D(N196), .Q(\ram[15][179] ) );
  LATCHX1_HVT \ram_reg[15][178]  ( .CLK(n17), .D(N195), .Q(\ram[15][178] ) );
  LATCHX1_HVT \ram_reg[15][177]  ( .CLK(n17), .D(N194), .Q(\ram[15][177] ) );
  LATCHX1_HVT \ram_reg[15][176]  ( .CLK(n17), .D(N193), .Q(\ram[15][176] ) );
  LATCHX1_HVT \ram_reg[15][175]  ( .CLK(n17), .D(N192), .Q(\ram[15][175] ) );
  LATCHX1_HVT \ram_reg[15][174]  ( .CLK(n16), .D(N191), .Q(\ram[15][174] ) );
  LATCHX1_HVT \ram_reg[15][173]  ( .CLK(n16), .D(N190), .Q(\ram[15][173] ) );
  LATCHX1_HVT \ram_reg[15][172]  ( .CLK(n16), .D(N189), .Q(\ram[15][172] ) );
  LATCHX1_HVT \ram_reg[15][171]  ( .CLK(n16), .D(N188), .Q(\ram[15][171] ) );
  LATCHX1_HVT \ram_reg[15][170]  ( .CLK(n16), .D(N187), .Q(\ram[15][170] ) );
  LATCHX1_HVT \ram_reg[15][169]  ( .CLK(n16), .D(N186), .Q(\ram[15][169] ) );
  LATCHX1_HVT \ram_reg[15][168]  ( .CLK(n16), .D(N185), .Q(\ram[15][168] ) );
  LATCHX1_HVT \ram_reg[15][167]  ( .CLK(n16), .D(N184), .Q(\ram[15][167] ) );
  LATCHX1_HVT \ram_reg[15][166]  ( .CLK(n16), .D(N183), .Q(\ram[15][166] ) );
  LATCHX1_HVT \ram_reg[15][165]  ( .CLK(n16), .D(N182), .Q(\ram[15][165] ) );
  LATCHX1_HVT \ram_reg[15][164]  ( .CLK(n16), .D(N181), .Q(\ram[15][164] ) );
  LATCHX1_HVT \ram_reg[15][163]  ( .CLK(n15), .D(N180), .Q(\ram[15][163] ) );
  LATCHX1_HVT \ram_reg[15][162]  ( .CLK(n15), .D(N179), .Q(\ram[15][162] ) );
  LATCHX1_HVT \ram_reg[15][161]  ( .CLK(n15), .D(N178), .Q(\ram[15][161] ) );
  LATCHX1_HVT \ram_reg[15][160]  ( .CLK(n15), .D(N177), .Q(\ram[15][160] ) );
  LATCHX1_HVT \ram_reg[15][159]  ( .CLK(n15), .D(N176), .Q(\ram[15][159] ) );
  LATCHX1_HVT \ram_reg[15][158]  ( .CLK(n15), .D(N175), .Q(\ram[15][158] ) );
  LATCHX1_HVT \ram_reg[15][157]  ( .CLK(n15), .D(N174), .Q(\ram[15][157] ) );
  LATCHX1_HVT \ram_reg[15][156]  ( .CLK(n15), .D(N173), .Q(\ram[15][156] ) );
  LATCHX1_HVT \ram_reg[15][155]  ( .CLK(n15), .D(N172), .Q(\ram[15][155] ) );
  LATCHX1_HVT \ram_reg[15][154]  ( .CLK(n15), .D(N171), .Q(\ram[15][154] ) );
  LATCHX1_HVT \ram_reg[15][153]  ( .CLK(n15), .D(N170), .Q(\ram[15][153] ) );
  LATCHX1_HVT \ram_reg[15][152]  ( .CLK(n14), .D(N169), .Q(\ram[15][152] ) );
  LATCHX1_HVT \ram_reg[15][151]  ( .CLK(n14), .D(N168), .Q(\ram[15][151] ) );
  LATCHX1_HVT \ram_reg[15][150]  ( .CLK(n14), .D(N167), .Q(\ram[15][150] ) );
  LATCHX1_HVT \ram_reg[15][149]  ( .CLK(n14), .D(N166), .Q(\ram[15][149] ) );
  LATCHX1_HVT \ram_reg[15][148]  ( .CLK(n14), .D(N165), .Q(\ram[15][148] ) );
  LATCHX1_HVT \ram_reg[15][147]  ( .CLK(n14), .D(N164), .Q(\ram[15][147] ) );
  LATCHX1_HVT \ram_reg[15][146]  ( .CLK(n14), .D(N163), .Q(\ram[15][146] ) );
  LATCHX1_HVT \ram_reg[15][145]  ( .CLK(n14), .D(N162), .Q(\ram[15][145] ) );
  LATCHX1_HVT \ram_reg[15][144]  ( .CLK(n14), .D(N161), .Q(\ram[15][144] ) );
  LATCHX1_HVT \ram_reg[15][143]  ( .CLK(n14), .D(N160), .Q(\ram[15][143] ) );
  LATCHX1_HVT \ram_reg[15][142]  ( .CLK(n14), .D(N159), .Q(\ram[15][142] ) );
  LATCHX1_HVT \ram_reg[15][141]  ( .CLK(n13), .D(N158), .Q(\ram[15][141] ) );
  LATCHX1_HVT \ram_reg[15][140]  ( .CLK(n13), .D(N157), .Q(\ram[15][140] ) );
  LATCHX1_HVT \ram_reg[15][139]  ( .CLK(n13), .D(N156), .Q(\ram[15][139] ) );
  LATCHX1_HVT \ram_reg[15][138]  ( .CLK(n12), .D(N155), .Q(\ram[15][138] ) );
  LATCHX1_HVT \ram_reg[15][137]  ( .CLK(n21), .D(N154), .Q(\ram[15][137] ) );
  LATCHX1_HVT \ram_reg[15][136]  ( .CLK(n20), .D(N153), .Q(\ram[15][136] ) );
  LATCHX1_HVT \ram_reg[15][135]  ( .CLK(n20), .D(N152), .Q(\ram[15][135] ) );
  LATCHX1_HVT \ram_reg[15][134]  ( .CLK(n19), .D(N151), .Q(\ram[15][134] ) );
  LATCHX1_HVT \ram_reg[15][133]  ( .CLK(n18), .D(N150), .Q(\ram[15][133] ) );
  LATCHX1_HVT \ram_reg[15][132]  ( .CLK(n17), .D(N149), .Q(\ram[15][132] ) );
  LATCHX1_HVT \ram_reg[15][131]  ( .CLK(n16), .D(N148), .Q(\ram[15][131] ) );
  LATCHX1_HVT \ram_reg[15][130]  ( .CLK(n15), .D(N147), .Q(\ram[15][130] ) );
  LATCHX1_HVT \ram_reg[15][129]  ( .CLK(n14), .D(N146), .Q(\ram[15][129] ) );
  LATCHX1_HVT \ram_reg[15][128]  ( .CLK(n11), .D(N145), .Q(\ram[15][128] ) );
  LATCHX1_HVT \ram_reg[15][127]  ( .CLK(n2), .D(N144), .Q(\ram[15][127] ) );
  LATCHX1_HVT \ram_reg[15][126]  ( .CLK(n2), .D(N143), .Q(\ram[15][126] ) );
  LATCHX1_HVT \ram_reg[15][125]  ( .CLK(n2), .D(N142), .Q(\ram[15][125] ) );
  LATCHX1_HVT \ram_reg[15][124]  ( .CLK(n2), .D(N141), .Q(\ram[15][124] ) );
  LATCHX1_HVT \ram_reg[15][123]  ( .CLK(n2), .D(N140), .Q(\ram[15][123] ) );
  LATCHX1_HVT \ram_reg[15][122]  ( .CLK(n1), .D(N139), .Q(\ram[15][122] ) );
  LATCHX1_HVT \ram_reg[15][121]  ( .CLK(n2), .D(N138), .Q(\ram[15][121] ) );
  LATCHX1_HVT \ram_reg[15][120]  ( .CLK(n2), .D(N137), .Q(\ram[15][120] ) );
  LATCHX1_HVT \ram_reg[15][119]  ( .CLK(n11), .D(N136), .Q(\ram[15][119] ) );
  LATCHX1_HVT \ram_reg[15][118]  ( .CLK(n10), .D(N135), .Q(\ram[15][118] ) );
  LATCHX1_HVT \ram_reg[15][117]  ( .CLK(n10), .D(N134), .Q(\ram[15][117] ) );
  LATCHX1_HVT \ram_reg[15][116]  ( .CLK(n9), .D(N133), .Q(\ram[15][116] ) );
  LATCHX1_HVT \ram_reg[15][115]  ( .CLK(n4), .D(N132), .Q(\ram[15][115] ) );
  LATCHX1_HVT \ram_reg[15][114]  ( .CLK(n9), .D(N131), .Q(\ram[15][114] ) );
  LATCHX1_HVT \ram_reg[15][113]  ( .CLK(n9), .D(N130), .Q(\ram[15][113] ) );
  LATCHX1_HVT \ram_reg[15][112]  ( .CLK(n10), .D(N129), .Q(\ram[15][112] ) );
  LATCHX1_HVT \ram_reg[15][111]  ( .CLK(n8), .D(N128), .Q(\ram[15][111] ) );
  LATCHX1_HVT \ram_reg[15][110]  ( .CLK(n8), .D(N127), .Q(\ram[15][110] ) );
  LATCHX1_HVT \ram_reg[15][109]  ( .CLK(n8), .D(N126), .Q(\ram[15][109] ) );
  LATCHX1_HVT \ram_reg[15][108]  ( .CLK(n5), .D(N125), .Q(\ram[15][108] ) );
  LATCHX1_HVT \ram_reg[15][107]  ( .CLK(n2), .D(N124), .Q(\ram[15][107] ) );
  LATCHX1_HVT \ram_reg[15][106]  ( .CLK(n8), .D(N123), .Q(\ram[15][106] ) );
  LATCHX1_HVT \ram_reg[15][105]  ( .CLK(n8), .D(N122), .Q(\ram[15][105] ) );
  LATCHX1_HVT \ram_reg[15][104]  ( .CLK(n8), .D(N121), .Q(\ram[15][104] ) );
  LATCHX1_HVT \ram_reg[15][103]  ( .CLK(n7), .D(N120), .Q(\ram[15][103] ) );
  LATCHX1_HVT \ram_reg[15][102]  ( .CLK(n6), .D(N119), .Q(\ram[15][102] ) );
  LATCHX1_HVT \ram_reg[15][101]  ( .CLK(n6), .D(N118), .Q(\ram[15][101] ) );
  LATCHX1_HVT \ram_reg[15][100]  ( .CLK(n7), .D(N117), .Q(\ram[15][100] ) );
  LATCHX1_HVT \ram_reg[15][99]  ( .CLK(n5), .D(N116), .Q(\ram[15][99] ) );
  LATCHX1_HVT \ram_reg[15][98]  ( .CLK(n6), .D(N114), .Q(\ram[15][98] ) );
  LATCHX1_HVT \ram_reg[15][97]  ( .CLK(n7), .D(N113), .Q(\ram[15][97] ) );
  LATCHX1_HVT \ram_reg[15][96]  ( .CLK(n11), .D(N112), .Q(\ram[15][96] ) );
  LATCHX1_HVT \ram_reg[15][95]  ( .CLK(n3), .D(N111), .Q(\ram[15][95] ) );
  LATCHX1_HVT \ram_reg[15][94]  ( .CLK(n3), .D(N110), .Q(\ram[15][94] ) );
  LATCHX1_HVT \ram_reg[15][93]  ( .CLK(n3), .D(N109), .Q(\ram[15][93] ) );
  LATCHX1_HVT \ram_reg[15][92]  ( .CLK(n2), .D(N108), .Q(\ram[15][92] ) );
  LATCHX1_HVT \ram_reg[15][91]  ( .CLK(n2), .D(N107), .Q(\ram[15][91] ) );
  LATCHX1_HVT \ram_reg[15][90]  ( .CLK(n3), .D(N106), .Q(\ram[15][90] ) );
  LATCHX1_HVT \ram_reg[15][89]  ( .CLK(n2), .D(N105), .Q(\ram[15][89] ) );
  LATCHX1_HVT \ram_reg[15][88]  ( .CLK(n3), .D(N104), .Q(\ram[15][88] ) );
  LATCHX1_HVT \ram_reg[15][87]  ( .CLK(n11), .D(N103), .Q(\ram[15][87] ) );
  LATCHX1_HVT \ram_reg[15][86]  ( .CLK(n10), .D(N102), .Q(\ram[15][86] ) );
  LATCHX1_HVT \ram_reg[15][85]  ( .CLK(n9), .D(N101), .Q(\ram[15][85] ) );
  LATCHX1_HVT \ram_reg[15][84]  ( .CLK(n9), .D(N100), .Q(\ram[15][84] ) );
  LATCHX1_HVT \ram_reg[15][83]  ( .CLK(n4), .D(N99), .Q(\ram[15][83] ) );
  LATCHX1_HVT \ram_reg[15][82]  ( .CLK(n10), .D(N98), .Q(\ram[15][82] ) );
  LATCHX1_HVT \ram_reg[15][81]  ( .CLK(n9), .D(N97), .Q(\ram[15][81] ) );
  LATCHX1_HVT \ram_reg[15][80]  ( .CLK(n10), .D(N96), .Q(\ram[15][80] ) );
  LATCHX1_HVT \ram_reg[15][79]  ( .CLK(n4), .D(N95), .Q(\ram[15][79] ) );
  LATCHX1_HVT \ram_reg[15][78]  ( .CLK(n3), .D(N94), .Q(\ram[15][78] ) );
  LATCHX1_HVT \ram_reg[15][77]  ( .CLK(n4), .D(N93), .Q(\ram[15][77] ) );
  LATCHX1_HVT \ram_reg[15][76]  ( .CLK(n3), .D(N92), .Q(\ram[15][76] ) );
  LATCHX1_HVT \ram_reg[15][75]  ( .CLK(n3), .D(N91), .Q(\ram[15][75] ) );
  LATCHX1_HVT \ram_reg[15][74]  ( .CLK(n1), .D(N90), .Q(\ram[15][74] ) );
  LATCHX1_HVT \ram_reg[15][73]  ( .CLK(n4), .D(N89), .Q(\ram[15][73] ) );
  LATCHX1_HVT \ram_reg[15][72]  ( .CLK(n4), .D(N88), .Q(\ram[15][72] ) );
  LATCHX1_HVT \ram_reg[15][71]  ( .CLK(n7), .D(N87), .Q(\ram[15][71] ) );
  LATCHX1_HVT \ram_reg[15][70]  ( .CLK(n7), .D(N86), .Q(\ram[15][70] ) );
  LATCHX1_HVT \ram_reg[15][69]  ( .CLK(n6), .D(N85), .Q(\ram[15][69] ) );
  LATCHX1_HVT \ram_reg[15][68]  ( .CLK(n7), .D(N84), .Q(\ram[15][68] ) );
  LATCHX1_HVT \ram_reg[15][67]  ( .CLK(n6), .D(N83), .Q(\ram[15][67] ) );
  LATCHX1_HVT \ram_reg[15][66]  ( .CLK(n5), .D(N82), .Q(\ram[15][66] ) );
  LATCHX1_HVT \ram_reg[15][65]  ( .CLK(n6), .D(N81), .Q(\ram[15][65] ) );
  LATCHX1_HVT \ram_reg[15][64]  ( .CLK(n11), .D(N80), .Q(\ram[15][64] ) );
  LATCHX1_HVT \ram_reg[15][63]  ( .CLK(n5), .D(N79), .Q(\ram[15][63] ) );
  LATCHX1_HVT \ram_reg[15][62]  ( .CLK(n5), .D(N78), .Q(\ram[15][62] ) );
  LATCHX1_HVT \ram_reg[15][61]  ( .CLK(n5), .D(N77), .Q(\ram[15][61] ) );
  LATCHX1_HVT \ram_reg[15][60]  ( .CLK(n5), .D(N76), .Q(\ram[15][60] ) );
  LATCHX1_HVT \ram_reg[15][59]  ( .CLK(n5), .D(N75), .Q(\ram[15][59] ) );
  LATCHX1_HVT \ram_reg[15][58]  ( .CLK(n4), .D(N74), .Q(\ram[15][58] ) );
  LATCHX1_HVT \ram_reg[15][57]  ( .CLK(n5), .D(N73), .Q(\ram[15][57] ) );
  LATCHX1_HVT \ram_reg[15][56]  ( .CLK(n5), .D(N72), .Q(\ram[15][56] ) );
  LATCHX1_HVT \ram_reg[15][55]  ( .CLK(n11), .D(N71), .Q(\ram[15][55] ) );
  LATCHX1_HVT \ram_reg[15][54]  ( .CLK(n9), .D(N70), .Q(\ram[15][54] ) );
  LATCHX1_HVT \ram_reg[15][53]  ( .CLK(n9), .D(N69), .Q(\ram[15][53] ) );
  LATCHX1_HVT \ram_reg[15][52]  ( .CLK(n10), .D(N68), .Q(\ram[15][52] ) );
  LATCHX1_HVT \ram_reg[15][51]  ( .CLK(n4), .D(N67), .Q(\ram[15][51] ) );
  LATCHX1_HVT \ram_reg[15][50]  ( .CLK(n1), .D(N66), .Q(\ram[15][50] ) );
  LATCHX1_HVT \ram_reg[15][49]  ( .CLK(n10), .D(N65), .Q(\ram[15][49] ) );
  LATCHX1_HVT \ram_reg[15][48]  ( .CLK(n10), .D(N64), .Q(\ram[15][48] ) );
  LATCHX1_HVT \ram_reg[15][47]  ( .CLK(n8), .D(N63), .Q(\ram[15][47] ) );
  LATCHX1_HVT \ram_reg[15][46]  ( .CLK(n8), .D(N62), .Q(\ram[15][46] ) );
  LATCHX1_HVT \ram_reg[15][45]  ( .CLK(n8), .D(N61), .Q(\ram[15][45] ) );
  LATCHX1_HVT \ram_reg[15][44]  ( .CLK(n8), .D(N60), .Q(\ram[15][44] ) );
  LATCHX1_HVT \ram_reg[15][43]  ( .CLK(n5), .D(N59), .Q(\ram[15][43] ) );
  LATCHX1_HVT \ram_reg[15][42]  ( .CLK(n9), .D(N58), .Q(\ram[15][42] ) );
  LATCHX1_HVT \ram_reg[15][41]  ( .CLK(n2), .D(N57), .Q(\ram[15][41] ) );
  LATCHX1_HVT \ram_reg[15][40]  ( .CLK(n8), .D(N56), .Q(\ram[15][40] ) );
  LATCHX1_HVT \ram_reg[15][39]  ( .CLK(n7), .D(N55), .Q(\ram[15][39] ) );
  LATCHX1_HVT \ram_reg[15][38]  ( .CLK(n7), .D(N54), .Q(\ram[15][38] ) );
  LATCHX1_HVT \ram_reg[15][37]  ( .CLK(n6), .D(N53), .Q(\ram[15][37] ) );
  LATCHX1_HVT \ram_reg[15][36]  ( .CLK(n6), .D(N52), .Q(\ram[15][36] ) );
  LATCHX1_HVT \ram_reg[15][35]  ( .CLK(n6), .D(N51), .Q(\ram[15][35] ) );
  LATCHX1_HVT \ram_reg[15][34]  ( .CLK(n8), .D(N50), .Q(\ram[15][34] ) );
  LATCHX1_HVT \ram_reg[15][33]  ( .CLK(n7), .D(N49), .Q(\ram[15][33] ) );
  LATCHX1_HVT \ram_reg[15][32]  ( .CLK(n11), .D(N48), .Q(\ram[15][32] ) );
  LATCHX1_HVT \ram_reg[15][31]  ( .CLK(n1), .D(N47), .Q(\ram[15][31] ) );
  LATCHX1_HVT \ram_reg[15][30]  ( .CLK(n1), .D(N46), .Q(\ram[15][30] ) );
  LATCHX1_HVT \ram_reg[15][29]  ( .CLK(n1), .D(N45), .Q(\ram[15][29] ) );
  LATCHX1_HVT \ram_reg[15][28]  ( .CLK(n1), .D(N44), .Q(\ram[15][28] ) );
  LATCHX1_HVT \ram_reg[15][27]  ( .CLK(n1), .D(N43), .Q(\ram[15][27] ) );
  LATCHX1_HVT \ram_reg[15][26]  ( .CLK(n1), .D(N42), .Q(\ram[15][26] ) );
  LATCHX1_HVT \ram_reg[15][25]  ( .CLK(n1), .D(N41), .Q(\ram[15][25] ) );
  LATCHX1_HVT \ram_reg[15][24]  ( .CLK(n1), .D(N40), .Q(\ram[15][24] ) );
  LATCHX1_HVT \ram_reg[15][23]  ( .CLK(n11), .D(N39), .Q(\ram[15][23] ) );
  LATCHX1_HVT \ram_reg[15][22]  ( .CLK(n10), .D(N38), .Q(\ram[15][22] ) );
  LATCHX1_HVT \ram_reg[15][21]  ( .CLK(n9), .D(N37), .Q(\ram[15][21] ) );
  LATCHX1_HVT \ram_reg[15][20]  ( .CLK(n9), .D(N36), .Q(\ram[15][20] ) );
  LATCHX1_HVT \ram_reg[15][19]  ( .CLK(n1), .D(N35), .Q(\ram[15][19] ) );
  LATCHX1_HVT \ram_reg[15][18]  ( .CLK(n9), .D(N34), .Q(\ram[15][18] ) );
  LATCHX1_HVT \ram_reg[15][17]  ( .CLK(n10), .D(N33), .Q(\ram[15][17] ) );
  LATCHX1_HVT \ram_reg[15][16]  ( .CLK(n10), .D(N32), .Q(\ram[15][16] ) );
  LATCHX1_HVT \ram_reg[15][15]  ( .CLK(n4), .D(N31), .Q(\ram[15][15] ) );
  LATCHX1_HVT \ram_reg[15][14]  ( .CLK(n4), .D(N30), .Q(\ram[15][14] ) );
  LATCHX1_HVT \ram_reg[15][13]  ( .CLK(n3), .D(N29), .Q(\ram[15][13] ) );
  LATCHX1_HVT \ram_reg[15][12]  ( .CLK(n3), .D(N28), .Q(\ram[15][12] ) );
  LATCHX1_HVT \ram_reg[15][11]  ( .CLK(n4), .D(N27), .Q(\ram[15][11] ) );
  LATCHX1_HVT \ram_reg[15][10]  ( .CLK(n3), .D(N26), .Q(\ram[15][10] ) );
  LATCHX1_HVT \ram_reg[15][9]  ( .CLK(n3), .D(N25), .Q(\ram[15][9] ) );
  LATCHX1_HVT \ram_reg[15][8]  ( .CLK(n4), .D(N24), .Q(\ram[15][8] ) );
  LATCHX1_HVT \ram_reg[15][7]  ( .CLK(n7), .D(N23), .Q(\ram[15][7] ) );
  LATCHX1_HVT \ram_reg[15][6]  ( .CLK(n7), .D(N22), .Q(\ram[15][6] ) );
  LATCHX1_HVT \ram_reg[15][5]  ( .CLK(n6), .D(N21), .Q(\ram[15][5] ) );
  LATCHX1_HVT \ram_reg[15][4]  ( .CLK(n6), .D(N20), .Q(\ram[15][4] ) );
  LATCHX1_HVT \ram_reg[15][3]  ( .CLK(n5), .D(N19), .Q(\ram[15][3] ) );
  LATCHX1_HVT \ram_reg[15][2]  ( .CLK(n6), .D(N18), .Q(\ram[15][2] ) );
  LATCHX1_HVT \ram_reg[15][1]  ( .CLK(n7), .D(N17), .Q(\ram[15][1] ) );
  LATCHX1_HVT \ram_reg[15][0]  ( .CLK(n11), .D(N16), .Q(\ram[15][0] ) );
  LATCHX1_HVT \ram_reg[14][255]  ( .CLK(n24), .D(N273), .Q(\ram[14][255] ) );
  LATCHX1_HVT \ram_reg[14][254]  ( .CLK(n24), .D(N272), .Q(\ram[14][254] ) );
  LATCHX1_HVT \ram_reg[14][253]  ( .CLK(n24), .D(N271), .Q(\ram[14][253] ) );
  LATCHX1_HVT \ram_reg[14][252]  ( .CLK(n24), .D(N270), .Q(\ram[14][252] ) );
  LATCHX1_HVT \ram_reg[14][251]  ( .CLK(N315), .D(N269), .Q(\ram[14][251] ) );
  LATCHX1_HVT \ram_reg[14][250]  ( .CLK(n37), .D(N268), .Q(\ram[14][250] ) );
  LATCHX1_HVT \ram_reg[14][249]  ( .CLK(n37), .D(N267), .Q(\ram[14][249] ) );
  LATCHX1_HVT \ram_reg[14][248]  ( .CLK(n36), .D(N266), .Q(\ram[14][248] ) );
  LATCHX1_HVT \ram_reg[14][247]  ( .CLK(n36), .D(N265), .Q(\ram[14][247] ) );
  LATCHX1_HVT \ram_reg[14][246]  ( .CLK(n36), .D(N264), .Q(\ram[14][246] ) );
  LATCHX1_HVT \ram_reg[14][245]  ( .CLK(n36), .D(N263), .Q(\ram[14][245] ) );
  LATCHX1_HVT \ram_reg[14][244]  ( .CLK(n36), .D(N262), .Q(\ram[14][244] ) );
  LATCHX1_HVT \ram_reg[14][243]  ( .CLK(n36), .D(N261), .Q(\ram[14][243] ) );
  LATCHX1_HVT \ram_reg[14][242]  ( .CLK(n36), .D(N260), .Q(\ram[14][242] ) );
  LATCHX1_HVT \ram_reg[14][241]  ( .CLK(n36), .D(N259), .Q(\ram[14][241] ) );
  LATCHX1_HVT \ram_reg[14][240]  ( .CLK(n36), .D(N258), .Q(\ram[14][240] ) );
  LATCHX1_HVT \ram_reg[14][239]  ( .CLK(n36), .D(N257), .Q(\ram[14][239] ) );
  LATCHX1_HVT \ram_reg[14][238]  ( .CLK(n36), .D(N256), .Q(\ram[14][238] ) );
  LATCHX1_HVT \ram_reg[14][237]  ( .CLK(n35), .D(N255), .Q(\ram[14][237] ) );
  LATCHX1_HVT \ram_reg[14][236]  ( .CLK(n35), .D(N254), .Q(\ram[14][236] ) );
  LATCHX1_HVT \ram_reg[14][235]  ( .CLK(n35), .D(N253), .Q(\ram[14][235] ) );
  LATCHX1_HVT \ram_reg[14][234]  ( .CLK(n35), .D(N252), .Q(\ram[14][234] ) );
  LATCHX1_HVT \ram_reg[14][233]  ( .CLK(n35), .D(N251), .Q(\ram[14][233] ) );
  LATCHX1_HVT \ram_reg[14][232]  ( .CLK(n35), .D(N250), .Q(\ram[14][232] ) );
  LATCHX1_HVT \ram_reg[14][231]  ( .CLK(n35), .D(N249), .Q(\ram[14][231] ) );
  LATCHX1_HVT \ram_reg[14][230]  ( .CLK(n35), .D(N248), .Q(\ram[14][230] ) );
  LATCHX1_HVT \ram_reg[14][229]  ( .CLK(n35), .D(N247), .Q(\ram[14][229] ) );
  LATCHX1_HVT \ram_reg[14][228]  ( .CLK(n35), .D(N246), .Q(\ram[14][228] ) );
  LATCHX1_HVT \ram_reg[14][227]  ( .CLK(N315), .D(N245), .Q(\ram[14][227] ) );
  LATCHX1_HVT \ram_reg[14][226]  ( .CLK(N315), .D(N244), .Q(\ram[14][226] ) );
  LATCHX1_HVT \ram_reg[14][225]  ( .CLK(n44), .D(N243), .Q(\ram[14][225] ) );
  LATCHX1_HVT \ram_reg[14][224]  ( .CLK(n44), .D(N242), .Q(\ram[14][224] ) );
  LATCHX1_HVT \ram_reg[14][223]  ( .CLK(n44), .D(N241), .Q(\ram[14][223] ) );
  LATCHX1_HVT \ram_reg[14][222]  ( .CLK(n44), .D(N240), .Q(\ram[14][222] ) );
  LATCHX1_HVT \ram_reg[14][221]  ( .CLK(n44), .D(N239), .Q(\ram[14][221] ) );
  LATCHX1_HVT \ram_reg[14][220]  ( .CLK(n44), .D(N238), .Q(\ram[14][220] ) );
  LATCHX1_HVT \ram_reg[14][219]  ( .CLK(n44), .D(N237), .Q(\ram[14][219] ) );
  LATCHX1_HVT \ram_reg[14][218]  ( .CLK(n44), .D(N236), .Q(\ram[14][218] ) );
  LATCHX1_HVT \ram_reg[14][217]  ( .CLK(n44), .D(N235), .Q(\ram[14][217] ) );
  LATCHX1_HVT \ram_reg[14][216]  ( .CLK(n44), .D(N234), .Q(\ram[14][216] ) );
  LATCHX1_HVT \ram_reg[14][215]  ( .CLK(n44), .D(N233), .Q(\ram[14][215] ) );
  LATCHX1_HVT \ram_reg[14][214]  ( .CLK(n43), .D(N232), .Q(\ram[14][214] ) );
  LATCHX1_HVT \ram_reg[14][213]  ( .CLK(n43), .D(N231), .Q(\ram[14][213] ) );
  LATCHX1_HVT \ram_reg[14][212]  ( .CLK(n43), .D(N230), .Q(\ram[14][212] ) );
  LATCHX1_HVT \ram_reg[14][211]  ( .CLK(n43), .D(N229), .Q(\ram[14][211] ) );
  LATCHX1_HVT \ram_reg[14][210]  ( .CLK(n43), .D(N228), .Q(\ram[14][210] ) );
  LATCHX1_HVT \ram_reg[14][209]  ( .CLK(n43), .D(N227), .Q(\ram[14][209] ) );
  LATCHX1_HVT \ram_reg[14][208]  ( .CLK(n43), .D(N226), .Q(\ram[14][208] ) );
  LATCHX1_HVT \ram_reg[14][207]  ( .CLK(n43), .D(N225), .Q(\ram[14][207] ) );
  LATCHX1_HVT \ram_reg[14][206]  ( .CLK(n43), .D(N224), .Q(\ram[14][206] ) );
  LATCHX1_HVT \ram_reg[14][205]  ( .CLK(n43), .D(N223), .Q(\ram[14][205] ) );
  LATCHX1_HVT \ram_reg[14][204]  ( .CLK(n43), .D(N222), .Q(\ram[14][204] ) );
  LATCHX1_HVT \ram_reg[14][203]  ( .CLK(n42), .D(N221), .Q(\ram[14][203] ) );
  LATCHX1_HVT \ram_reg[14][202]  ( .CLK(n42), .D(N220), .Q(\ram[14][202] ) );
  LATCHX1_HVT \ram_reg[14][201]  ( .CLK(n42), .D(N219), .Q(\ram[14][201] ) );
  LATCHX1_HVT \ram_reg[14][200]  ( .CLK(n42), .D(N218), .Q(\ram[14][200] ) );
  LATCHX1_HVT \ram_reg[14][199]  ( .CLK(n42), .D(N217), .Q(\ram[14][199] ) );
  LATCHX1_HVT \ram_reg[14][198]  ( .CLK(n42), .D(N216), .Q(\ram[14][198] ) );
  LATCHX1_HVT \ram_reg[14][197]  ( .CLK(n42), .D(N214), .Q(\ram[14][197] ) );
  LATCHX1_HVT \ram_reg[14][196]  ( .CLK(n42), .D(N213), .Q(\ram[14][196] ) );
  LATCHX1_HVT \ram_reg[14][195]  ( .CLK(n42), .D(N212), .Q(\ram[14][195] ) );
  LATCHX1_HVT \ram_reg[14][194]  ( .CLK(n42), .D(N211), .Q(\ram[14][194] ) );
  LATCHX1_HVT \ram_reg[14][193]  ( .CLK(n42), .D(N210), .Q(\ram[14][193] ) );
  LATCHX1_HVT \ram_reg[14][192]  ( .CLK(n41), .D(N209), .Q(\ram[14][192] ) );
  LATCHX1_HVT \ram_reg[14][191]  ( .CLK(n41), .D(N208), .Q(\ram[14][191] ) );
  LATCHX1_HVT \ram_reg[14][190]  ( .CLK(n41), .D(N207), .Q(\ram[14][190] ) );
  LATCHX1_HVT \ram_reg[14][189]  ( .CLK(n41), .D(N206), .Q(\ram[14][189] ) );
  LATCHX1_HVT \ram_reg[14][188]  ( .CLK(n41), .D(N205), .Q(\ram[14][188] ) );
  LATCHX1_HVT \ram_reg[14][187]  ( .CLK(n41), .D(N204), .Q(\ram[14][187] ) );
  LATCHX1_HVT \ram_reg[14][186]  ( .CLK(n41), .D(N203), .Q(\ram[14][186] ) );
  LATCHX1_HVT \ram_reg[14][185]  ( .CLK(n41), .D(N202), .Q(\ram[14][185] ) );
  LATCHX1_HVT \ram_reg[14][184]  ( .CLK(n41), .D(N201), .Q(\ram[14][184] ) );
  LATCHX1_HVT \ram_reg[14][183]  ( .CLK(n41), .D(N200), .Q(\ram[14][183] ) );
  LATCHX1_HVT \ram_reg[14][182]  ( .CLK(n41), .D(N199), .Q(\ram[14][182] ) );
  LATCHX1_HVT \ram_reg[14][181]  ( .CLK(n40), .D(N198), .Q(\ram[14][181] ) );
  LATCHX1_HVT \ram_reg[14][180]  ( .CLK(n40), .D(N197), .Q(\ram[14][180] ) );
  LATCHX1_HVT \ram_reg[14][179]  ( .CLK(n40), .D(N196), .Q(\ram[14][179] ) );
  LATCHX1_HVT \ram_reg[14][178]  ( .CLK(n40), .D(N195), .Q(\ram[14][178] ) );
  LATCHX1_HVT \ram_reg[14][177]  ( .CLK(n40), .D(N194), .Q(\ram[14][177] ) );
  LATCHX1_HVT \ram_reg[14][176]  ( .CLK(n40), .D(N193), .Q(\ram[14][176] ) );
  LATCHX1_HVT \ram_reg[14][175]  ( .CLK(n40), .D(N192), .Q(\ram[14][175] ) );
  LATCHX1_HVT \ram_reg[14][174]  ( .CLK(n40), .D(N191), .Q(\ram[14][174] ) );
  LATCHX1_HVT \ram_reg[14][173]  ( .CLK(n40), .D(N190), .Q(\ram[14][173] ) );
  LATCHX1_HVT \ram_reg[14][172]  ( .CLK(n40), .D(N189), .Q(\ram[14][172] ) );
  LATCHX1_HVT \ram_reg[14][171]  ( .CLK(n40), .D(N188), .Q(\ram[14][171] ) );
  LATCHX1_HVT \ram_reg[14][170]  ( .CLK(n39), .D(N187), .Q(\ram[14][170] ) );
  LATCHX1_HVT \ram_reg[14][169]  ( .CLK(n39), .D(N186), .Q(\ram[14][169] ) );
  LATCHX1_HVT \ram_reg[14][168]  ( .CLK(n39), .D(N185), .Q(\ram[14][168] ) );
  LATCHX1_HVT \ram_reg[14][167]  ( .CLK(n39), .D(N184), .Q(\ram[14][167] ) );
  LATCHX1_HVT \ram_reg[14][166]  ( .CLK(n39), .D(N183), .Q(\ram[14][166] ) );
  LATCHX1_HVT \ram_reg[14][165]  ( .CLK(n39), .D(N182), .Q(\ram[14][165] ) );
  LATCHX1_HVT \ram_reg[14][164]  ( .CLK(n39), .D(N181), .Q(\ram[14][164] ) );
  LATCHX1_HVT \ram_reg[14][163]  ( .CLK(n39), .D(N180), .Q(\ram[14][163] ) );
  LATCHX1_HVT \ram_reg[14][162]  ( .CLK(n39), .D(N179), .Q(\ram[14][162] ) );
  LATCHX1_HVT \ram_reg[14][161]  ( .CLK(n39), .D(N178), .Q(\ram[14][161] ) );
  LATCHX1_HVT \ram_reg[14][160]  ( .CLK(n39), .D(N177), .Q(\ram[14][160] ) );
  LATCHX1_HVT \ram_reg[14][159]  ( .CLK(n38), .D(N176), .Q(\ram[14][159] ) );
  LATCHX1_HVT \ram_reg[14][158]  ( .CLK(n38), .D(N175), .Q(\ram[14][158] ) );
  LATCHX1_HVT \ram_reg[14][157]  ( .CLK(n38), .D(N174), .Q(\ram[14][157] ) );
  LATCHX1_HVT \ram_reg[14][156]  ( .CLK(n38), .D(N173), .Q(\ram[14][156] ) );
  LATCHX1_HVT \ram_reg[14][155]  ( .CLK(n38), .D(N172), .Q(\ram[14][155] ) );
  LATCHX1_HVT \ram_reg[14][154]  ( .CLK(n38), .D(N171), .Q(\ram[14][154] ) );
  LATCHX1_HVT \ram_reg[14][153]  ( .CLK(n38), .D(N170), .Q(\ram[14][153] ) );
  LATCHX1_HVT \ram_reg[14][152]  ( .CLK(n38), .D(N169), .Q(\ram[14][152] ) );
  LATCHX1_HVT \ram_reg[14][151]  ( .CLK(n38), .D(N168), .Q(\ram[14][151] ) );
  LATCHX1_HVT \ram_reg[14][150]  ( .CLK(n38), .D(N167), .Q(\ram[14][150] ) );
  LATCHX1_HVT \ram_reg[14][149]  ( .CLK(n38), .D(N166), .Q(\ram[14][149] ) );
  LATCHX1_HVT \ram_reg[14][148]  ( .CLK(n37), .D(N165), .Q(\ram[14][148] ) );
  LATCHX1_HVT \ram_reg[14][147]  ( .CLK(n37), .D(N164), .Q(\ram[14][147] ) );
  LATCHX1_HVT \ram_reg[14][146]  ( .CLK(n37), .D(N163), .Q(\ram[14][146] ) );
  LATCHX1_HVT \ram_reg[14][145]  ( .CLK(n37), .D(N162), .Q(\ram[14][145] ) );
  LATCHX1_HVT \ram_reg[14][144]  ( .CLK(n37), .D(N161), .Q(\ram[14][144] ) );
  LATCHX1_HVT \ram_reg[14][143]  ( .CLK(n37), .D(N160), .Q(\ram[14][143] ) );
  LATCHX1_HVT \ram_reg[14][142]  ( .CLK(n37), .D(N159), .Q(\ram[14][142] ) );
  LATCHX1_HVT \ram_reg[14][141]  ( .CLK(n37), .D(N158), .Q(\ram[14][141] ) );
  LATCHX1_HVT \ram_reg[14][140]  ( .CLK(n37), .D(N157), .Q(\ram[14][140] ) );
  LATCHX1_HVT \ram_reg[14][139]  ( .CLK(n36), .D(N156), .Q(\ram[14][139] ) );
  LATCHX1_HVT \ram_reg[14][138]  ( .CLK(n35), .D(N155), .Q(\ram[14][138] ) );
  LATCHX1_HVT \ram_reg[14][137]  ( .CLK(N315), .D(N154), .Q(\ram[14][137] ) );
  LATCHX1_HVT \ram_reg[14][136]  ( .CLK(n44), .D(N153), .Q(\ram[14][136] ) );
  LATCHX1_HVT \ram_reg[14][135]  ( .CLK(n43), .D(N152), .Q(\ram[14][135] ) );
  LATCHX1_HVT \ram_reg[14][134]  ( .CLK(n42), .D(N151), .Q(\ram[14][134] ) );
  LATCHX1_HVT \ram_reg[14][133]  ( .CLK(n41), .D(N150), .Q(\ram[14][133] ) );
  LATCHX1_HVT \ram_reg[14][132]  ( .CLK(n40), .D(N149), .Q(\ram[14][132] ) );
  LATCHX1_HVT \ram_reg[14][131]  ( .CLK(n39), .D(N148), .Q(\ram[14][131] ) );
  LATCHX1_HVT \ram_reg[14][130]  ( .CLK(n38), .D(N147), .Q(\ram[14][130] ) );
  LATCHX1_HVT \ram_reg[14][129]  ( .CLK(n37), .D(N146), .Q(\ram[14][129] ) );
  LATCHX1_HVT \ram_reg[14][128]  ( .CLK(n35), .D(N145), .Q(\ram[14][128] ) );
  LATCHX1_HVT \ram_reg[14][127]  ( .CLK(n26), .D(N144), .Q(\ram[14][127] ) );
  LATCHX1_HVT \ram_reg[14][126]  ( .CLK(n25), .D(N143), .Q(\ram[14][126] ) );
  LATCHX1_HVT \ram_reg[14][125]  ( .CLK(n25), .D(N142), .Q(\ram[14][125] ) );
  LATCHX1_HVT \ram_reg[14][124]  ( .CLK(n25), .D(N141), .Q(\ram[14][124] ) );
  LATCHX1_HVT \ram_reg[14][123]  ( .CLK(n25), .D(N140), .Q(\ram[14][123] ) );
  LATCHX1_HVT \ram_reg[14][122]  ( .CLK(n25), .D(N139), .Q(\ram[14][122] ) );
  LATCHX1_HVT \ram_reg[14][121]  ( .CLK(n25), .D(N138), .Q(\ram[14][121] ) );
  LATCHX1_HVT \ram_reg[14][120]  ( .CLK(n25), .D(N137), .Q(\ram[14][120] ) );
  LATCHX1_HVT \ram_reg[14][119]  ( .CLK(n34), .D(N136), .Q(\ram[14][119] ) );
  LATCHX1_HVT \ram_reg[14][118]  ( .CLK(n33), .D(N135), .Q(\ram[14][118] ) );
  LATCHX1_HVT \ram_reg[14][117]  ( .CLK(n33), .D(N134), .Q(\ram[14][117] ) );
  LATCHX1_HVT \ram_reg[14][116]  ( .CLK(n32), .D(N133), .Q(\ram[14][116] ) );
  LATCHX1_HVT \ram_reg[14][115]  ( .CLK(n28), .D(N132), .Q(\ram[14][115] ) );
  LATCHX1_HVT \ram_reg[14][114]  ( .CLK(n33), .D(N131), .Q(\ram[14][114] ) );
  LATCHX1_HVT \ram_reg[14][113]  ( .CLK(n32), .D(N130), .Q(\ram[14][113] ) );
  LATCHX1_HVT \ram_reg[14][112]  ( .CLK(n34), .D(N129), .Q(\ram[14][112] ) );
  LATCHX1_HVT \ram_reg[14][111]  ( .CLK(n32), .D(N128), .Q(\ram[14][111] ) );
  LATCHX1_HVT \ram_reg[14][110]  ( .CLK(n32), .D(N127), .Q(\ram[14][110] ) );
  LATCHX1_HVT \ram_reg[14][109]  ( .CLK(n31), .D(N126), .Q(\ram[14][109] ) );
  LATCHX1_HVT \ram_reg[14][108]  ( .CLK(n28), .D(N125), .Q(\ram[14][108] ) );
  LATCHX1_HVT \ram_reg[14][107]  ( .CLK(n25), .D(N124), .Q(\ram[14][107] ) );
  LATCHX1_HVT \ram_reg[14][106]  ( .CLK(n31), .D(N123), .Q(\ram[14][106] ) );
  LATCHX1_HVT \ram_reg[14][105]  ( .CLK(n31), .D(N122), .Q(\ram[14][105] ) );
  LATCHX1_HVT \ram_reg[14][104]  ( .CLK(n31), .D(N121), .Q(\ram[14][104] ) );
  LATCHX1_HVT \ram_reg[14][103]  ( .CLK(n31), .D(N120), .Q(\ram[14][103] ) );
  LATCHX1_HVT \ram_reg[14][102]  ( .CLK(n30), .D(N119), .Q(\ram[14][102] ) );
  LATCHX1_HVT \ram_reg[14][101]  ( .CLK(n29), .D(N118), .Q(\ram[14][101] ) );
  LATCHX1_HVT \ram_reg[14][100]  ( .CLK(n30), .D(N117), .Q(\ram[14][100] ) );
  LATCHX1_HVT \ram_reg[14][99]  ( .CLK(n29), .D(N116), .Q(\ram[14][99] ) );
  LATCHX1_HVT \ram_reg[14][98]  ( .CLK(n29), .D(N114), .Q(\ram[14][98] ) );
  LATCHX1_HVT \ram_reg[14][97]  ( .CLK(n30), .D(N113), .Q(\ram[14][97] ) );
  LATCHX1_HVT \ram_reg[14][96]  ( .CLK(n34), .D(N112), .Q(\ram[14][96] ) );
  LATCHX1_HVT \ram_reg[14][95]  ( .CLK(n26), .D(N111), .Q(\ram[14][95] ) );
  LATCHX1_HVT \ram_reg[14][94]  ( .CLK(n26), .D(N110), .Q(\ram[14][94] ) );
  LATCHX1_HVT \ram_reg[14][93]  ( .CLK(n26), .D(N109), .Q(\ram[14][93] ) );
  LATCHX1_HVT \ram_reg[14][92]  ( .CLK(n26), .D(N108), .Q(\ram[14][92] ) );
  LATCHX1_HVT \ram_reg[14][91]  ( .CLK(n26), .D(N107), .Q(\ram[14][91] ) );
  LATCHX1_HVT \ram_reg[14][90]  ( .CLK(n26), .D(N106), .Q(\ram[14][90] ) );
  LATCHX1_HVT \ram_reg[14][89]  ( .CLK(n26), .D(N105), .Q(\ram[14][89] ) );
  LATCHX1_HVT \ram_reg[14][88]  ( .CLK(n26), .D(N104), .Q(\ram[14][88] ) );
  LATCHX1_HVT \ram_reg[14][87]  ( .CLK(n34), .D(N103), .Q(\ram[14][87] ) );
  LATCHX1_HVT \ram_reg[14][86]  ( .CLK(n34), .D(N102), .Q(\ram[14][86] ) );
  LATCHX1_HVT \ram_reg[14][85]  ( .CLK(n32), .D(N101), .Q(\ram[14][85] ) );
  LATCHX1_HVT \ram_reg[14][84]  ( .CLK(n33), .D(N100), .Q(\ram[14][84] ) );
  LATCHX1_HVT \ram_reg[14][83]  ( .CLK(n28), .D(N99), .Q(\ram[14][83] ) );
  LATCHX1_HVT \ram_reg[14][82]  ( .CLK(n33), .D(N98), .Q(\ram[14][82] ) );
  LATCHX1_HVT \ram_reg[14][81]  ( .CLK(n32), .D(N97), .Q(\ram[14][81] ) );
  LATCHX1_HVT \ram_reg[14][80]  ( .CLK(n33), .D(N96), .Q(\ram[14][80] ) );
  LATCHX1_HVT \ram_reg[14][79]  ( .CLK(n27), .D(N95), .Q(\ram[14][79] ) );
  LATCHX1_HVT \ram_reg[14][78]  ( .CLK(n27), .D(N94), .Q(\ram[14][78] ) );
  LATCHX1_HVT \ram_reg[14][77]  ( .CLK(n27), .D(N93), .Q(\ram[14][77] ) );
  LATCHX1_HVT \ram_reg[14][76]  ( .CLK(n27), .D(N92), .Q(\ram[14][76] ) );
  LATCHX1_HVT \ram_reg[14][75]  ( .CLK(n26), .D(N91), .Q(\ram[14][75] ) );
  LATCHX1_HVT \ram_reg[14][74]  ( .CLK(n25), .D(N90), .Q(\ram[14][74] ) );
  LATCHX1_HVT \ram_reg[14][73]  ( .CLK(n27), .D(N89), .Q(\ram[14][73] ) );
  LATCHX1_HVT \ram_reg[14][72]  ( .CLK(n27), .D(N88), .Q(\ram[14][72] ) );
  LATCHX1_HVT \ram_reg[14][71]  ( .CLK(n31), .D(N87), .Q(\ram[14][71] ) );
  LATCHX1_HVT \ram_reg[14][70]  ( .CLK(n30), .D(N86), .Q(\ram[14][70] ) );
  LATCHX1_HVT \ram_reg[14][69]  ( .CLK(n29), .D(N85), .Q(\ram[14][69] ) );
  LATCHX1_HVT \ram_reg[14][68]  ( .CLK(n30), .D(N84), .Q(\ram[14][68] ) );
  LATCHX1_HVT \ram_reg[14][67]  ( .CLK(n29), .D(N83), .Q(\ram[14][67] ) );
  LATCHX1_HVT \ram_reg[14][66]  ( .CLK(n29), .D(N82), .Q(\ram[14][66] ) );
  LATCHX1_HVT \ram_reg[14][65]  ( .CLK(n30), .D(N81), .Q(\ram[14][65] ) );
  LATCHX1_HVT \ram_reg[14][64]  ( .CLK(n34), .D(N80), .Q(\ram[14][64] ) );
  LATCHX1_HVT \ram_reg[14][63]  ( .CLK(n28), .D(N79), .Q(\ram[14][63] ) );
  LATCHX1_HVT \ram_reg[14][62]  ( .CLK(n28), .D(N78), .Q(\ram[14][62] ) );
  LATCHX1_HVT \ram_reg[14][61]  ( .CLK(n28), .D(N77), .Q(\ram[14][61] ) );
  LATCHX1_HVT \ram_reg[14][60]  ( .CLK(n28), .D(N76), .Q(\ram[14][60] ) );
  LATCHX1_HVT \ram_reg[14][59]  ( .CLK(n28), .D(N75), .Q(\ram[14][59] ) );
  LATCHX1_HVT \ram_reg[14][58]  ( .CLK(n28), .D(N74), .Q(\ram[14][58] ) );
  LATCHX1_HVT \ram_reg[14][57]  ( .CLK(n28), .D(N73), .Q(\ram[14][57] ) );
  LATCHX1_HVT \ram_reg[14][56]  ( .CLK(n28), .D(N72), .Q(\ram[14][56] ) );
  LATCHX1_HVT \ram_reg[14][55]  ( .CLK(n34), .D(N71), .Q(\ram[14][55] ) );
  LATCHX1_HVT \ram_reg[14][54]  ( .CLK(n33), .D(N70), .Q(\ram[14][54] ) );
  LATCHX1_HVT \ram_reg[14][53]  ( .CLK(n32), .D(N69), .Q(\ram[14][53] ) );
  LATCHX1_HVT \ram_reg[14][52]  ( .CLK(n33), .D(N68), .Q(\ram[14][52] ) );
  LATCHX1_HVT \ram_reg[14][51]  ( .CLK(n28), .D(N67), .Q(\ram[14][51] ) );
  LATCHX1_HVT \ram_reg[14][50]  ( .CLK(n24), .D(N66), .Q(\ram[14][50] ) );
  LATCHX1_HVT \ram_reg[14][49]  ( .CLK(n33), .D(N65), .Q(\ram[14][49] ) );
  LATCHX1_HVT \ram_reg[14][48]  ( .CLK(n34), .D(N64), .Q(\ram[14][48] ) );
  LATCHX1_HVT \ram_reg[14][47]  ( .CLK(n32), .D(N63), .Q(\ram[14][47] ) );
  LATCHX1_HVT \ram_reg[14][46]  ( .CLK(n31), .D(N62), .Q(\ram[14][46] ) );
  LATCHX1_HVT \ram_reg[14][45]  ( .CLK(n31), .D(N61), .Q(\ram[14][45] ) );
  LATCHX1_HVT \ram_reg[14][44]  ( .CLK(n31), .D(N60), .Q(\ram[14][44] ) );
  LATCHX1_HVT \ram_reg[14][43]  ( .CLK(n29), .D(N59), .Q(\ram[14][43] ) );
  LATCHX1_HVT \ram_reg[14][42]  ( .CLK(n32), .D(N58), .Q(\ram[14][42] ) );
  LATCHX1_HVT \ram_reg[14][41]  ( .CLK(n25), .D(N57), .Q(\ram[14][41] ) );
  LATCHX1_HVT \ram_reg[14][40]  ( .CLK(n32), .D(N56), .Q(\ram[14][40] ) );
  LATCHX1_HVT \ram_reg[14][39]  ( .CLK(n31), .D(N55), .Q(\ram[14][39] ) );
  LATCHX1_HVT \ram_reg[14][38]  ( .CLK(n30), .D(N54), .Q(\ram[14][38] ) );
  LATCHX1_HVT \ram_reg[14][37]  ( .CLK(n29), .D(N53), .Q(\ram[14][37] ) );
  LATCHX1_HVT \ram_reg[14][36]  ( .CLK(n30), .D(N52), .Q(\ram[14][36] ) );
  LATCHX1_HVT \ram_reg[14][35]  ( .CLK(n29), .D(N51), .Q(\ram[14][35] ) );
  LATCHX1_HVT \ram_reg[14][34]  ( .CLK(n31), .D(N50), .Q(\ram[14][34] ) );
  LATCHX1_HVT \ram_reg[14][33]  ( .CLK(n30), .D(N49), .Q(\ram[14][33] ) );
  LATCHX1_HVT \ram_reg[14][32]  ( .CLK(n34), .D(N48), .Q(\ram[14][32] ) );
  LATCHX1_HVT \ram_reg[14][31]  ( .CLK(n25), .D(N47), .Q(\ram[14][31] ) );
  LATCHX1_HVT \ram_reg[14][30]  ( .CLK(n24), .D(N46), .Q(\ram[14][30] ) );
  LATCHX1_HVT \ram_reg[14][29]  ( .CLK(n24), .D(N45), .Q(\ram[14][29] ) );
  LATCHX1_HVT \ram_reg[14][28]  ( .CLK(n24), .D(N44), .Q(\ram[14][28] ) );
  LATCHX1_HVT \ram_reg[14][27]  ( .CLK(n25), .D(N43), .Q(\ram[14][27] ) );
  LATCHX1_HVT \ram_reg[14][26]  ( .CLK(n24), .D(N42), .Q(\ram[14][26] ) );
  LATCHX1_HVT \ram_reg[14][25]  ( .CLK(n24), .D(N41), .Q(\ram[14][25] ) );
  LATCHX1_HVT \ram_reg[14][24]  ( .CLK(n24), .D(N40), .Q(\ram[14][24] ) );
  LATCHX1_HVT \ram_reg[14][23]  ( .CLK(n34), .D(N39), .Q(\ram[14][23] ) );
  LATCHX1_HVT \ram_reg[14][22]  ( .CLK(n33), .D(N38), .Q(\ram[14][22] ) );
  LATCHX1_HVT \ram_reg[14][21]  ( .CLK(n33), .D(N37), .Q(\ram[14][21] ) );
  LATCHX1_HVT \ram_reg[14][20]  ( .CLK(n32), .D(N36), .Q(\ram[14][20] ) );
  LATCHX1_HVT \ram_reg[14][19]  ( .CLK(n24), .D(N35), .Q(\ram[14][19] ) );
  LATCHX1_HVT \ram_reg[14][18]  ( .CLK(n32), .D(N34), .Q(\ram[14][18] ) );
  LATCHX1_HVT \ram_reg[14][17]  ( .CLK(n33), .D(N33), .Q(\ram[14][17] ) );
  LATCHX1_HVT \ram_reg[14][16]  ( .CLK(n34), .D(N32), .Q(\ram[14][16] ) );
  LATCHX1_HVT \ram_reg[14][15]  ( .CLK(n27), .D(N31), .Q(\ram[14][15] ) );
  LATCHX1_HVT \ram_reg[14][14]  ( .CLK(n27), .D(N30), .Q(\ram[14][14] ) );
  LATCHX1_HVT \ram_reg[14][13]  ( .CLK(n26), .D(N29), .Q(\ram[14][13] ) );
  LATCHX1_HVT \ram_reg[14][12]  ( .CLK(n27), .D(N28), .Q(\ram[14][12] ) );
  LATCHX1_HVT \ram_reg[14][11]  ( .CLK(n27), .D(N27), .Q(\ram[14][11] ) );
  LATCHX1_HVT \ram_reg[14][10]  ( .CLK(n26), .D(N26), .Q(\ram[14][10] ) );
  LATCHX1_HVT \ram_reg[14][9]  ( .CLK(n27), .D(N25), .Q(\ram[14][9] ) );
  LATCHX1_HVT \ram_reg[14][8]  ( .CLK(n27), .D(N24), .Q(\ram[14][8] ) );
  LATCHX1_HVT \ram_reg[14][7]  ( .CLK(n31), .D(N23), .Q(\ram[14][7] ) );
  LATCHX1_HVT \ram_reg[14][6]  ( .CLK(n30), .D(N22), .Q(\ram[14][6] ) );
  LATCHX1_HVT \ram_reg[14][5]  ( .CLK(n29), .D(N21), .Q(\ram[14][5] ) );
  LATCHX1_HVT \ram_reg[14][4]  ( .CLK(n30), .D(N20), .Q(\ram[14][4] ) );
  LATCHX1_HVT \ram_reg[14][3]  ( .CLK(n29), .D(N19), .Q(\ram[14][3] ) );
  LATCHX1_HVT \ram_reg[14][2]  ( .CLK(n29), .D(N18), .Q(\ram[14][2] ) );
  LATCHX1_HVT \ram_reg[14][1]  ( .CLK(n30), .D(N17), .Q(\ram[14][1] ) );
  LATCHX1_HVT \ram_reg[14][0]  ( .CLK(n34), .D(N16), .Q(\ram[14][0] ) );
  LATCHX1_HVT \ram_reg[13][255]  ( .CLK(n47), .D(N273), .Q(\ram[13][255] ) );
  LATCHX1_HVT \ram_reg[13][254]  ( .CLK(n47), .D(N272), .Q(\ram[13][254] ) );
  LATCHX1_HVT \ram_reg[13][253]  ( .CLK(N312), .D(N271), .Q(\ram[13][253] ) );
  LATCHX1_HVT \ram_reg[13][252]  ( .CLK(N312), .D(N270), .Q(\ram[13][252] ) );
  LATCHX1_HVT \ram_reg[13][251]  ( .CLK(N312), .D(N269), .Q(\ram[13][251] ) );
  LATCHX1_HVT \ram_reg[13][250]  ( .CLK(n59), .D(N268), .Q(\ram[13][250] ) );
  LATCHX1_HVT \ram_reg[13][249]  ( .CLK(n59), .D(N267), .Q(\ram[13][249] ) );
  LATCHX1_HVT \ram_reg[13][248]  ( .CLK(n59), .D(N266), .Q(\ram[13][248] ) );
  LATCHX1_HVT \ram_reg[13][247]  ( .CLK(n59), .D(N265), .Q(\ram[13][247] ) );
  LATCHX1_HVT \ram_reg[13][246]  ( .CLK(n59), .D(N264), .Q(\ram[13][246] ) );
  LATCHX1_HVT \ram_reg[13][245]  ( .CLK(n59), .D(N263), .Q(\ram[13][245] ) );
  LATCHX1_HVT \ram_reg[13][244]  ( .CLK(n59), .D(N262), .Q(\ram[13][244] ) );
  LATCHX1_HVT \ram_reg[13][243]  ( .CLK(n59), .D(N261), .Q(\ram[13][243] ) );
  LATCHX1_HVT \ram_reg[13][242]  ( .CLK(n59), .D(N260), .Q(\ram[13][242] ) );
  LATCHX1_HVT \ram_reg[13][241]  ( .CLK(n59), .D(N259), .Q(\ram[13][241] ) );
  LATCHX1_HVT \ram_reg[13][240]  ( .CLK(n59), .D(N258), .Q(\ram[13][240] ) );
  LATCHX1_HVT \ram_reg[13][239]  ( .CLK(n58), .D(N257), .Q(\ram[13][239] ) );
  LATCHX1_HVT \ram_reg[13][238]  ( .CLK(n58), .D(N256), .Q(\ram[13][238] ) );
  LATCHX1_HVT \ram_reg[13][237]  ( .CLK(n58), .D(N255), .Q(\ram[13][237] ) );
  LATCHX1_HVT \ram_reg[13][236]  ( .CLK(n58), .D(N254), .Q(\ram[13][236] ) );
  LATCHX1_HVT \ram_reg[13][235]  ( .CLK(n58), .D(N253), .Q(\ram[13][235] ) );
  LATCHX1_HVT \ram_reg[13][234]  ( .CLK(n58), .D(N252), .Q(\ram[13][234] ) );
  LATCHX1_HVT \ram_reg[13][233]  ( .CLK(n58), .D(N251), .Q(\ram[13][233] ) );
  LATCHX1_HVT \ram_reg[13][232]  ( .CLK(n58), .D(N250), .Q(\ram[13][232] ) );
  LATCHX1_HVT \ram_reg[13][231]  ( .CLK(n58), .D(N249), .Q(\ram[13][231] ) );
  LATCHX1_HVT \ram_reg[13][230]  ( .CLK(n58), .D(N248), .Q(\ram[13][230] ) );
  LATCHX1_HVT \ram_reg[13][229]  ( .CLK(n58), .D(N247), .Q(\ram[13][229] ) );
  LATCHX1_HVT \ram_reg[13][228]  ( .CLK(n57), .D(N246), .Q(\ram[13][228] ) );
  LATCHX1_HVT \ram_reg[13][227]  ( .CLK(n67), .D(N245), .Q(\ram[13][227] ) );
  LATCHX1_HVT \ram_reg[13][226]  ( .CLK(n67), .D(N244), .Q(\ram[13][226] ) );
  LATCHX1_HVT \ram_reg[13][225]  ( .CLK(n67), .D(N243), .Q(\ram[13][225] ) );
  LATCHX1_HVT \ram_reg[13][224]  ( .CLK(n67), .D(N242), .Q(\ram[13][224] ) );
  LATCHX1_HVT \ram_reg[13][223]  ( .CLK(n67), .D(N241), .Q(\ram[13][223] ) );
  LATCHX1_HVT \ram_reg[13][222]  ( .CLK(n67), .D(N240), .Q(\ram[13][222] ) );
  LATCHX1_HVT \ram_reg[13][221]  ( .CLK(n67), .D(N239), .Q(\ram[13][221] ) );
  LATCHX1_HVT \ram_reg[13][220]  ( .CLK(n67), .D(N238), .Q(\ram[13][220] ) );
  LATCHX1_HVT \ram_reg[13][219]  ( .CLK(n67), .D(N237), .Q(\ram[13][219] ) );
  LATCHX1_HVT \ram_reg[13][218]  ( .CLK(n67), .D(N236), .Q(\ram[13][218] ) );
  LATCHX1_HVT \ram_reg[13][217]  ( .CLK(n67), .D(N235), .Q(\ram[13][217] ) );
  LATCHX1_HVT \ram_reg[13][216]  ( .CLK(n66), .D(N234), .Q(\ram[13][216] ) );
  LATCHX1_HVT \ram_reg[13][215]  ( .CLK(n66), .D(N233), .Q(\ram[13][215] ) );
  LATCHX1_HVT \ram_reg[13][214]  ( .CLK(n66), .D(N232), .Q(\ram[13][214] ) );
  LATCHX1_HVT \ram_reg[13][213]  ( .CLK(n66), .D(N231), .Q(\ram[13][213] ) );
  LATCHX1_HVT \ram_reg[13][212]  ( .CLK(n66), .D(N230), .Q(\ram[13][212] ) );
  LATCHX1_HVT \ram_reg[13][211]  ( .CLK(n66), .D(N229), .Q(\ram[13][211] ) );
  LATCHX1_HVT \ram_reg[13][210]  ( .CLK(n66), .D(N228), .Q(\ram[13][210] ) );
  LATCHX1_HVT \ram_reg[13][209]  ( .CLK(n66), .D(N227), .Q(\ram[13][209] ) );
  LATCHX1_HVT \ram_reg[13][208]  ( .CLK(n66), .D(N226), .Q(\ram[13][208] ) );
  LATCHX1_HVT \ram_reg[13][207]  ( .CLK(n66), .D(N225), .Q(\ram[13][207] ) );
  LATCHX1_HVT \ram_reg[13][206]  ( .CLK(n66), .D(N224), .Q(\ram[13][206] ) );
  LATCHX1_HVT \ram_reg[13][205]  ( .CLK(n65), .D(N223), .Q(\ram[13][205] ) );
  LATCHX1_HVT \ram_reg[13][204]  ( .CLK(n65), .D(N222), .Q(\ram[13][204] ) );
  LATCHX1_HVT \ram_reg[13][203]  ( .CLK(n65), .D(N221), .Q(\ram[13][203] ) );
  LATCHX1_HVT \ram_reg[13][202]  ( .CLK(n65), .D(N220), .Q(\ram[13][202] ) );
  LATCHX1_HVT \ram_reg[13][201]  ( .CLK(n65), .D(N219), .Q(\ram[13][201] ) );
  LATCHX1_HVT \ram_reg[13][200]  ( .CLK(n65), .D(N218), .Q(\ram[13][200] ) );
  LATCHX1_HVT \ram_reg[13][199]  ( .CLK(n65), .D(N217), .Q(\ram[13][199] ) );
  LATCHX1_HVT \ram_reg[13][198]  ( .CLK(n65), .D(N216), .Q(\ram[13][198] ) );
  LATCHX1_HVT \ram_reg[13][197]  ( .CLK(n65), .D(N214), .Q(\ram[13][197] ) );
  LATCHX1_HVT \ram_reg[13][196]  ( .CLK(n65), .D(N213), .Q(\ram[13][196] ) );
  LATCHX1_HVT \ram_reg[13][195]  ( .CLK(n65), .D(N212), .Q(\ram[13][195] ) );
  LATCHX1_HVT \ram_reg[13][194]  ( .CLK(n64), .D(N211), .Q(\ram[13][194] ) );
  LATCHX1_HVT \ram_reg[13][193]  ( .CLK(n64), .D(N210), .Q(\ram[13][193] ) );
  LATCHX1_HVT \ram_reg[13][192]  ( .CLK(n64), .D(N209), .Q(\ram[13][192] ) );
  LATCHX1_HVT \ram_reg[13][191]  ( .CLK(n64), .D(N208), .Q(\ram[13][191] ) );
  LATCHX1_HVT \ram_reg[13][190]  ( .CLK(n64), .D(N207), .Q(\ram[13][190] ) );
  LATCHX1_HVT \ram_reg[13][189]  ( .CLK(n64), .D(N206), .Q(\ram[13][189] ) );
  LATCHX1_HVT \ram_reg[13][188]  ( .CLK(n64), .D(N205), .Q(\ram[13][188] ) );
  LATCHX1_HVT \ram_reg[13][187]  ( .CLK(n64), .D(N204), .Q(\ram[13][187] ) );
  LATCHX1_HVT \ram_reg[13][186]  ( .CLK(n64), .D(N203), .Q(\ram[13][186] ) );
  LATCHX1_HVT \ram_reg[13][185]  ( .CLK(n64), .D(N202), .Q(\ram[13][185] ) );
  LATCHX1_HVT \ram_reg[13][184]  ( .CLK(n64), .D(N201), .Q(\ram[13][184] ) );
  LATCHX1_HVT \ram_reg[13][183]  ( .CLK(n63), .D(N200), .Q(\ram[13][183] ) );
  LATCHX1_HVT \ram_reg[13][182]  ( .CLK(n63), .D(N199), .Q(\ram[13][182] ) );
  LATCHX1_HVT \ram_reg[13][181]  ( .CLK(n63), .D(N198), .Q(\ram[13][181] ) );
  LATCHX1_HVT \ram_reg[13][180]  ( .CLK(n63), .D(N197), .Q(\ram[13][180] ) );
  LATCHX1_HVT \ram_reg[13][179]  ( .CLK(n63), .D(N196), .Q(\ram[13][179] ) );
  LATCHX1_HVT \ram_reg[13][178]  ( .CLK(n63), .D(N195), .Q(\ram[13][178] ) );
  LATCHX1_HVT \ram_reg[13][177]  ( .CLK(n63), .D(N194), .Q(\ram[13][177] ) );
  LATCHX1_HVT \ram_reg[13][176]  ( .CLK(n63), .D(N193), .Q(\ram[13][176] ) );
  LATCHX1_HVT \ram_reg[13][175]  ( .CLK(n63), .D(N192), .Q(\ram[13][175] ) );
  LATCHX1_HVT \ram_reg[13][174]  ( .CLK(n63), .D(N191), .Q(\ram[13][174] ) );
  LATCHX1_HVT \ram_reg[13][173]  ( .CLK(n63), .D(N190), .Q(\ram[13][173] ) );
  LATCHX1_HVT \ram_reg[13][172]  ( .CLK(n62), .D(N189), .Q(\ram[13][172] ) );
  LATCHX1_HVT \ram_reg[13][171]  ( .CLK(n62), .D(N188), .Q(\ram[13][171] ) );
  LATCHX1_HVT \ram_reg[13][170]  ( .CLK(n62), .D(N187), .Q(\ram[13][170] ) );
  LATCHX1_HVT \ram_reg[13][169]  ( .CLK(n62), .D(N186), .Q(\ram[13][169] ) );
  LATCHX1_HVT \ram_reg[13][168]  ( .CLK(n62), .D(N185), .Q(\ram[13][168] ) );
  LATCHX1_HVT \ram_reg[13][167]  ( .CLK(n62), .D(N184), .Q(\ram[13][167] ) );
  LATCHX1_HVT \ram_reg[13][166]  ( .CLK(n62), .D(N183), .Q(\ram[13][166] ) );
  LATCHX1_HVT \ram_reg[13][165]  ( .CLK(n62), .D(N182), .Q(\ram[13][165] ) );
  LATCHX1_HVT \ram_reg[13][164]  ( .CLK(n62), .D(N181), .Q(\ram[13][164] ) );
  LATCHX1_HVT \ram_reg[13][163]  ( .CLK(n62), .D(N180), .Q(\ram[13][163] ) );
  LATCHX1_HVT \ram_reg[13][162]  ( .CLK(n62), .D(N179), .Q(\ram[13][162] ) );
  LATCHX1_HVT \ram_reg[13][161]  ( .CLK(n61), .D(N178), .Q(\ram[13][161] ) );
  LATCHX1_HVT \ram_reg[13][160]  ( .CLK(n61), .D(N177), .Q(\ram[13][160] ) );
  LATCHX1_HVT \ram_reg[13][159]  ( .CLK(n61), .D(N176), .Q(\ram[13][159] ) );
  LATCHX1_HVT \ram_reg[13][158]  ( .CLK(n61), .D(N175), .Q(\ram[13][158] ) );
  LATCHX1_HVT \ram_reg[13][157]  ( .CLK(n61), .D(N174), .Q(\ram[13][157] ) );
  LATCHX1_HVT \ram_reg[13][156]  ( .CLK(n61), .D(N173), .Q(\ram[13][156] ) );
  LATCHX1_HVT \ram_reg[13][155]  ( .CLK(n61), .D(N172), .Q(\ram[13][155] ) );
  LATCHX1_HVT \ram_reg[13][154]  ( .CLK(n61), .D(N171), .Q(\ram[13][154] ) );
  LATCHX1_HVT \ram_reg[13][153]  ( .CLK(n61), .D(N170), .Q(\ram[13][153] ) );
  LATCHX1_HVT \ram_reg[13][152]  ( .CLK(n61), .D(N169), .Q(\ram[13][152] ) );
  LATCHX1_HVT \ram_reg[13][151]  ( .CLK(n61), .D(N168), .Q(\ram[13][151] ) );
  LATCHX1_HVT \ram_reg[13][150]  ( .CLK(n60), .D(N167), .Q(\ram[13][150] ) );
  LATCHX1_HVT \ram_reg[13][149]  ( .CLK(n60), .D(N166), .Q(\ram[13][149] ) );
  LATCHX1_HVT \ram_reg[13][148]  ( .CLK(n60), .D(N165), .Q(\ram[13][148] ) );
  LATCHX1_HVT \ram_reg[13][147]  ( .CLK(n60), .D(N164), .Q(\ram[13][147] ) );
  LATCHX1_HVT \ram_reg[13][146]  ( .CLK(n60), .D(N163), .Q(\ram[13][146] ) );
  LATCHX1_HVT \ram_reg[13][145]  ( .CLK(n60), .D(N162), .Q(\ram[13][145] ) );
  LATCHX1_HVT \ram_reg[13][144]  ( .CLK(n60), .D(N161), .Q(\ram[13][144] ) );
  LATCHX1_HVT \ram_reg[13][143]  ( .CLK(n60), .D(N160), .Q(\ram[13][143] ) );
  LATCHX1_HVT \ram_reg[13][142]  ( .CLK(n60), .D(N159), .Q(\ram[13][142] ) );
  LATCHX1_HVT \ram_reg[13][141]  ( .CLK(n60), .D(N158), .Q(\ram[13][141] ) );
  LATCHX1_HVT \ram_reg[13][140]  ( .CLK(n60), .D(N157), .Q(\ram[13][140] ) );
  LATCHX1_HVT \ram_reg[13][139]  ( .CLK(n59), .D(N156), .Q(\ram[13][139] ) );
  LATCHX1_HVT \ram_reg[13][138]  ( .CLK(n58), .D(N155), .Q(\ram[13][138] ) );
  LATCHX1_HVT \ram_reg[13][137]  ( .CLK(N312), .D(N154), .Q(\ram[13][137] ) );
  LATCHX1_HVT \ram_reg[13][136]  ( .CLK(n67), .D(N153), .Q(\ram[13][136] ) );
  LATCHX1_HVT \ram_reg[13][135]  ( .CLK(n66), .D(N152), .Q(\ram[13][135] ) );
  LATCHX1_HVT \ram_reg[13][134]  ( .CLK(n65), .D(N151), .Q(\ram[13][134] ) );
  LATCHX1_HVT \ram_reg[13][133]  ( .CLK(n64), .D(N150), .Q(\ram[13][133] ) );
  LATCHX1_HVT \ram_reg[13][132]  ( .CLK(n63), .D(N149), .Q(\ram[13][132] ) );
  LATCHX1_HVT \ram_reg[13][131]  ( .CLK(n62), .D(N148), .Q(\ram[13][131] ) );
  LATCHX1_HVT \ram_reg[13][130]  ( .CLK(n61), .D(N147), .Q(\ram[13][130] ) );
  LATCHX1_HVT \ram_reg[13][129]  ( .CLK(n60), .D(N146), .Q(\ram[13][129] ) );
  LATCHX1_HVT \ram_reg[13][128]  ( .CLK(n57), .D(N145), .Q(\ram[13][128] ) );
  LATCHX1_HVT \ram_reg[13][127]  ( .CLK(n48), .D(N144), .Q(\ram[13][127] ) );
  LATCHX1_HVT \ram_reg[13][126]  ( .CLK(n48), .D(N143), .Q(\ram[13][126] ) );
  LATCHX1_HVT \ram_reg[13][125]  ( .CLK(n48), .D(N142), .Q(\ram[13][125] ) );
  LATCHX1_HVT \ram_reg[13][124]  ( .CLK(n48), .D(N141), .Q(\ram[13][124] ) );
  LATCHX1_HVT \ram_reg[13][123]  ( .CLK(n48), .D(N140), .Q(\ram[13][123] ) );
  LATCHX1_HVT \ram_reg[13][122]  ( .CLK(n48), .D(N139), .Q(\ram[13][122] ) );
  LATCHX1_HVT \ram_reg[13][121]  ( .CLK(n48), .D(N138), .Q(\ram[13][121] ) );
  LATCHX1_HVT \ram_reg[13][120]  ( .CLK(n48), .D(N137), .Q(\ram[13][120] ) );
  LATCHX1_HVT \ram_reg[13][119]  ( .CLK(n57), .D(N136), .Q(\ram[13][119] ) );
  LATCHX1_HVT \ram_reg[13][118]  ( .CLK(n56), .D(N135), .Q(\ram[13][118] ) );
  LATCHX1_HVT \ram_reg[13][117]  ( .CLK(n56), .D(N134), .Q(\ram[13][117] ) );
  LATCHX1_HVT \ram_reg[13][116]  ( .CLK(n55), .D(N133), .Q(\ram[13][116] ) );
  LATCHX1_HVT \ram_reg[13][115]  ( .CLK(n50), .D(N132), .Q(\ram[13][115] ) );
  LATCHX1_HVT \ram_reg[13][114]  ( .CLK(n56), .D(N131), .Q(\ram[13][114] ) );
  LATCHX1_HVT \ram_reg[13][113]  ( .CLK(n55), .D(N130), .Q(\ram[13][113] ) );
  LATCHX1_HVT \ram_reg[13][112]  ( .CLK(n57), .D(N129), .Q(\ram[13][112] ) );
  LATCHX1_HVT \ram_reg[13][111]  ( .CLK(n55), .D(N128), .Q(\ram[13][111] ) );
  LATCHX1_HVT \ram_reg[13][110]  ( .CLK(n54), .D(N127), .Q(\ram[13][110] ) );
  LATCHX1_HVT \ram_reg[13][109]  ( .CLK(n54), .D(N126), .Q(\ram[13][109] ) );
  LATCHX1_HVT \ram_reg[13][108]  ( .CLK(n51), .D(N125), .Q(\ram[13][108] ) );
  LATCHX1_HVT \ram_reg[13][107]  ( .CLK(n48), .D(N124), .Q(\ram[13][107] ) );
  LATCHX1_HVT \ram_reg[13][106]  ( .CLK(n54), .D(N123), .Q(\ram[13][106] ) );
  LATCHX1_HVT \ram_reg[13][105]  ( .CLK(n54), .D(N122), .Q(\ram[13][105] ) );
  LATCHX1_HVT \ram_reg[13][104]  ( .CLK(n54), .D(N121), .Q(\ram[13][104] ) );
  LATCHX1_HVT \ram_reg[13][103]  ( .CLK(n54), .D(N120), .Q(\ram[13][103] ) );
  LATCHX1_HVT \ram_reg[13][102]  ( .CLK(n53), .D(N119), .Q(\ram[13][102] ) );
  LATCHX1_HVT \ram_reg[13][101]  ( .CLK(n52), .D(N118), .Q(\ram[13][101] ) );
  LATCHX1_HVT \ram_reg[13][100]  ( .CLK(n53), .D(N117), .Q(\ram[13][100] ) );
  LATCHX1_HVT \ram_reg[13][99]  ( .CLK(n52), .D(N116), .Q(\ram[13][99] ) );
  LATCHX1_HVT \ram_reg[13][98]  ( .CLK(n52), .D(N114), .Q(\ram[13][98] ) );
  LATCHX1_HVT \ram_reg[13][97]  ( .CLK(n53), .D(N113), .Q(\ram[13][97] ) );
  LATCHX1_HVT \ram_reg[13][96]  ( .CLK(n57), .D(N112), .Q(\ram[13][96] ) );
  LATCHX1_HVT \ram_reg[13][95]  ( .CLK(n49), .D(N111), .Q(\ram[13][95] ) );
  LATCHX1_HVT \ram_reg[13][94]  ( .CLK(n49), .D(N110), .Q(\ram[13][94] ) );
  LATCHX1_HVT \ram_reg[13][93]  ( .CLK(n49), .D(N109), .Q(\ram[13][93] ) );
  LATCHX1_HVT \ram_reg[13][92]  ( .CLK(n49), .D(N108), .Q(\ram[13][92] ) );
  LATCHX1_HVT \ram_reg[13][91]  ( .CLK(n49), .D(N107), .Q(\ram[13][91] ) );
  LATCHX1_HVT \ram_reg[13][90]  ( .CLK(n49), .D(N106), .Q(\ram[13][90] ) );
  LATCHX1_HVT \ram_reg[13][89]  ( .CLK(n48), .D(N105), .Q(\ram[13][89] ) );
  LATCHX1_HVT \ram_reg[13][88]  ( .CLK(n49), .D(N104), .Q(\ram[13][88] ) );
  LATCHX1_HVT \ram_reg[13][87]  ( .CLK(n57), .D(N103), .Q(\ram[13][87] ) );
  LATCHX1_HVT \ram_reg[13][86]  ( .CLK(n57), .D(N102), .Q(\ram[13][86] ) );
  LATCHX1_HVT \ram_reg[13][85]  ( .CLK(n55), .D(N101), .Q(\ram[13][85] ) );
  LATCHX1_HVT \ram_reg[13][84]  ( .CLK(n56), .D(N100), .Q(\ram[13][84] ) );
  LATCHX1_HVT \ram_reg[13][83]  ( .CLK(n50), .D(N99), .Q(\ram[13][83] ) );
  LATCHX1_HVT \ram_reg[13][82]  ( .CLK(n56), .D(N98), .Q(\ram[13][82] ) );
  LATCHX1_HVT \ram_reg[13][81]  ( .CLK(n55), .D(N97), .Q(\ram[13][81] ) );
  LATCHX1_HVT \ram_reg[13][80]  ( .CLK(n56), .D(N96), .Q(\ram[13][80] ) );
  LATCHX1_HVT \ram_reg[13][79]  ( .CLK(n50), .D(N95), .Q(\ram[13][79] ) );
  LATCHX1_HVT \ram_reg[13][78]  ( .CLK(n50), .D(N94), .Q(\ram[13][78] ) );
  LATCHX1_HVT \ram_reg[13][77]  ( .CLK(n50), .D(N93), .Q(\ram[13][77] ) );
  LATCHX1_HVT \ram_reg[13][76]  ( .CLK(n49), .D(N92), .Q(\ram[13][76] ) );
  LATCHX1_HVT \ram_reg[13][75]  ( .CLK(n49), .D(N91), .Q(\ram[13][75] ) );
  LATCHX1_HVT \ram_reg[13][74]  ( .CLK(n48), .D(N90), .Q(\ram[13][74] ) );
  LATCHX1_HVT \ram_reg[13][73]  ( .CLK(n50), .D(N89), .Q(\ram[13][73] ) );
  LATCHX1_HVT \ram_reg[13][72]  ( .CLK(n50), .D(N88), .Q(\ram[13][72] ) );
  LATCHX1_HVT \ram_reg[13][71]  ( .CLK(n53), .D(N87), .Q(\ram[13][71] ) );
  LATCHX1_HVT \ram_reg[13][70]  ( .CLK(n53), .D(N86), .Q(\ram[13][70] ) );
  LATCHX1_HVT \ram_reg[13][69]  ( .CLK(n52), .D(N85), .Q(\ram[13][69] ) );
  LATCHX1_HVT \ram_reg[13][68]  ( .CLK(n53), .D(N84), .Q(\ram[13][68] ) );
  LATCHX1_HVT \ram_reg[13][67]  ( .CLK(n52), .D(N83), .Q(\ram[13][67] ) );
  LATCHX1_HVT \ram_reg[13][66]  ( .CLK(n51), .D(N82), .Q(\ram[13][66] ) );
  LATCHX1_HVT \ram_reg[13][65]  ( .CLK(n52), .D(N81), .Q(\ram[13][65] ) );
  LATCHX1_HVT \ram_reg[13][64]  ( .CLK(n57), .D(N80), .Q(\ram[13][64] ) );
  LATCHX1_HVT \ram_reg[13][63]  ( .CLK(n51), .D(N79), .Q(\ram[13][63] ) );
  LATCHX1_HVT \ram_reg[13][62]  ( .CLK(n51), .D(N78), .Q(\ram[13][62] ) );
  LATCHX1_HVT \ram_reg[13][61]  ( .CLK(n51), .D(N77), .Q(\ram[13][61] ) );
  LATCHX1_HVT \ram_reg[13][60]  ( .CLK(n51), .D(N76), .Q(\ram[13][60] ) );
  LATCHX1_HVT \ram_reg[13][59]  ( .CLK(n51), .D(N75), .Q(\ram[13][59] ) );
  LATCHX1_HVT \ram_reg[13][58]  ( .CLK(n51), .D(N74), .Q(\ram[13][58] ) );
  LATCHX1_HVT \ram_reg[13][57]  ( .CLK(n51), .D(N73), .Q(\ram[13][57] ) );
  LATCHX1_HVT \ram_reg[13][56]  ( .CLK(n51), .D(N72), .Q(\ram[13][56] ) );
  LATCHX1_HVT \ram_reg[13][55]  ( .CLK(n57), .D(N71), .Q(\ram[13][55] ) );
  LATCHX1_HVT \ram_reg[13][54]  ( .CLK(n55), .D(N70), .Q(\ram[13][54] ) );
  LATCHX1_HVT \ram_reg[13][53]  ( .CLK(n55), .D(N69), .Q(\ram[13][53] ) );
  LATCHX1_HVT \ram_reg[13][52]  ( .CLK(n56), .D(N68), .Q(\ram[13][52] ) );
  LATCHX1_HVT \ram_reg[13][51]  ( .CLK(n51), .D(N67), .Q(\ram[13][51] ) );
  LATCHX1_HVT \ram_reg[13][50]  ( .CLK(n47), .D(N66), .Q(\ram[13][50] ) );
  LATCHX1_HVT \ram_reg[13][49]  ( .CLK(n56), .D(N65), .Q(\ram[13][49] ) );
  LATCHX1_HVT \ram_reg[13][48]  ( .CLK(n56), .D(N64), .Q(\ram[13][48] ) );
  LATCHX1_HVT \ram_reg[13][47]  ( .CLK(n55), .D(N63), .Q(\ram[13][47] ) );
  LATCHX1_HVT \ram_reg[13][46]  ( .CLK(n54), .D(N62), .Q(\ram[13][46] ) );
  LATCHX1_HVT \ram_reg[13][45]  ( .CLK(n54), .D(N61), .Q(\ram[13][45] ) );
  LATCHX1_HVT \ram_reg[13][44]  ( .CLK(n54), .D(N60), .Q(\ram[13][44] ) );
  LATCHX1_HVT \ram_reg[13][43]  ( .CLK(n51), .D(N59), .Q(\ram[13][43] ) );
  LATCHX1_HVT \ram_reg[13][42]  ( .CLK(n55), .D(N58), .Q(\ram[13][42] ) );
  LATCHX1_HVT \ram_reg[13][41]  ( .CLK(n48), .D(N57), .Q(\ram[13][41] ) );
  LATCHX1_HVT \ram_reg[13][40]  ( .CLK(n54), .D(N56), .Q(\ram[13][40] ) );
  LATCHX1_HVT \ram_reg[13][39]  ( .CLK(n53), .D(N55), .Q(\ram[13][39] ) );
  LATCHX1_HVT \ram_reg[13][38]  ( .CLK(n53), .D(N54), .Q(\ram[13][38] ) );
  LATCHX1_HVT \ram_reg[13][37]  ( .CLK(n52), .D(N53), .Q(\ram[13][37] ) );
  LATCHX1_HVT \ram_reg[13][36]  ( .CLK(n52), .D(N52), .Q(\ram[13][36] ) );
  LATCHX1_HVT \ram_reg[13][35]  ( .CLK(n52), .D(N51), .Q(\ram[13][35] ) );
  LATCHX1_HVT \ram_reg[13][34]  ( .CLK(n54), .D(N50), .Q(\ram[13][34] ) );
  LATCHX1_HVT \ram_reg[13][33]  ( .CLK(n53), .D(N49), .Q(\ram[13][33] ) );
  LATCHX1_HVT \ram_reg[13][32]  ( .CLK(n57), .D(N48), .Q(\ram[13][32] ) );
  LATCHX1_HVT \ram_reg[13][31]  ( .CLK(n47), .D(N47), .Q(\ram[13][31] ) );
  LATCHX1_HVT \ram_reg[13][30]  ( .CLK(n47), .D(N46), .Q(\ram[13][30] ) );
  LATCHX1_HVT \ram_reg[13][29]  ( .CLK(n47), .D(N45), .Q(\ram[13][29] ) );
  LATCHX1_HVT \ram_reg[13][28]  ( .CLK(n47), .D(N44), .Q(\ram[13][28] ) );
  LATCHX1_HVT \ram_reg[13][27]  ( .CLK(n47), .D(N43), .Q(\ram[13][27] ) );
  LATCHX1_HVT \ram_reg[13][26]  ( .CLK(n47), .D(N42), .Q(\ram[13][26] ) );
  LATCHX1_HVT \ram_reg[13][25]  ( .CLK(n47), .D(N41), .Q(\ram[13][25] ) );
  LATCHX1_HVT \ram_reg[13][24]  ( .CLK(n47), .D(N40), .Q(\ram[13][24] ) );
  LATCHX1_HVT \ram_reg[13][23]  ( .CLK(n57), .D(N39), .Q(\ram[13][23] ) );
  LATCHX1_HVT \ram_reg[13][22]  ( .CLK(n56), .D(N38), .Q(\ram[13][22] ) );
  LATCHX1_HVT \ram_reg[13][21]  ( .CLK(n55), .D(N37), .Q(\ram[13][21] ) );
  LATCHX1_HVT \ram_reg[13][20]  ( .CLK(n55), .D(N36), .Q(\ram[13][20] ) );
  LATCHX1_HVT \ram_reg[13][19]  ( .CLK(n47), .D(N35), .Q(\ram[13][19] ) );
  LATCHX1_HVT \ram_reg[13][18]  ( .CLK(n55), .D(N34), .Q(\ram[13][18] ) );
  LATCHX1_HVT \ram_reg[13][17]  ( .CLK(n56), .D(N33), .Q(\ram[13][17] ) );
  LATCHX1_HVT \ram_reg[13][16]  ( .CLK(n56), .D(N32), .Q(\ram[13][16] ) );
  LATCHX1_HVT \ram_reg[13][15]  ( .CLK(n50), .D(N31), .Q(\ram[13][15] ) );
  LATCHX1_HVT \ram_reg[13][14]  ( .CLK(n50), .D(N30), .Q(\ram[13][14] ) );
  LATCHX1_HVT \ram_reg[13][13]  ( .CLK(n49), .D(N29), .Q(\ram[13][13] ) );
  LATCHX1_HVT \ram_reg[13][12]  ( .CLK(n50), .D(N28), .Q(\ram[13][12] ) );
  LATCHX1_HVT \ram_reg[13][11]  ( .CLK(n50), .D(N27), .Q(\ram[13][11] ) );
  LATCHX1_HVT \ram_reg[13][10]  ( .CLK(n49), .D(N26), .Q(\ram[13][10] ) );
  LATCHX1_HVT \ram_reg[13][9]  ( .CLK(n49), .D(N25), .Q(\ram[13][9] ) );
  LATCHX1_HVT \ram_reg[13][8]  ( .CLK(n50), .D(N24), .Q(\ram[13][8] ) );
  LATCHX1_HVT \ram_reg[13][7]  ( .CLK(n54), .D(N23), .Q(\ram[13][7] ) );
  LATCHX1_HVT \ram_reg[13][6]  ( .CLK(n53), .D(N22), .Q(\ram[13][6] ) );
  LATCHX1_HVT \ram_reg[13][5]  ( .CLK(n52), .D(N21), .Q(\ram[13][5] ) );
  LATCHX1_HVT \ram_reg[13][4]  ( .CLK(n53), .D(N20), .Q(\ram[13][4] ) );
  LATCHX1_HVT \ram_reg[13][3]  ( .CLK(n52), .D(N19), .Q(\ram[13][3] ) );
  LATCHX1_HVT \ram_reg[13][2]  ( .CLK(n52), .D(N18), .Q(\ram[13][2] ) );
  LATCHX1_HVT \ram_reg[13][1]  ( .CLK(n53), .D(N17), .Q(\ram[13][1] ) );
  LATCHX1_HVT \ram_reg[13][0]  ( .CLK(n57), .D(N16), .Q(\ram[13][0] ) );
  LATCHX1_HVT \ram_reg[12][255]  ( .CLK(N309), .D(N273), .Q(\ram[12][255] ) );
  LATCHX1_HVT \ram_reg[12][254]  ( .CLK(N309), .D(N272), .Q(\ram[12][254] ) );
  LATCHX1_HVT \ram_reg[12][253]  ( .CLK(N309), .D(N271), .Q(\ram[12][253] ) );
  LATCHX1_HVT \ram_reg[12][252]  ( .CLK(N309), .D(N270), .Q(\ram[12][252] ) );
  LATCHX1_HVT \ram_reg[12][251]  ( .CLK(n90), .D(N269), .Q(\ram[12][251] ) );
  LATCHX1_HVT \ram_reg[12][250]  ( .CLK(n82), .D(N268), .Q(\ram[12][250] ) );
  LATCHX1_HVT \ram_reg[12][249]  ( .CLK(n82), .D(N267), .Q(\ram[12][249] ) );
  LATCHX1_HVT \ram_reg[12][248]  ( .CLK(n82), .D(N266), .Q(\ram[12][248] ) );
  LATCHX1_HVT \ram_reg[12][247]  ( .CLK(n82), .D(N265), .Q(\ram[12][247] ) );
  LATCHX1_HVT \ram_reg[12][246]  ( .CLK(n82), .D(N264), .Q(\ram[12][246] ) );
  LATCHX1_HVT \ram_reg[12][245]  ( .CLK(n82), .D(N263), .Q(\ram[12][245] ) );
  LATCHX1_HVT \ram_reg[12][244]  ( .CLK(n82), .D(N262), .Q(\ram[12][244] ) );
  LATCHX1_HVT \ram_reg[12][243]  ( .CLK(n82), .D(N261), .Q(\ram[12][243] ) );
  LATCHX1_HVT \ram_reg[12][242]  ( .CLK(n82), .D(N260), .Q(\ram[12][242] ) );
  LATCHX1_HVT \ram_reg[12][241]  ( .CLK(n81), .D(N259), .Q(\ram[12][241] ) );
  LATCHX1_HVT \ram_reg[12][240]  ( .CLK(n81), .D(N258), .Q(\ram[12][240] ) );
  LATCHX1_HVT \ram_reg[12][239]  ( .CLK(n81), .D(N257), .Q(\ram[12][239] ) );
  LATCHX1_HVT \ram_reg[12][238]  ( .CLK(n81), .D(N256), .Q(\ram[12][238] ) );
  LATCHX1_HVT \ram_reg[12][237]  ( .CLK(n81), .D(N255), .Q(\ram[12][237] ) );
  LATCHX1_HVT \ram_reg[12][236]  ( .CLK(n81), .D(N254), .Q(\ram[12][236] ) );
  LATCHX1_HVT \ram_reg[12][235]  ( .CLK(n81), .D(N253), .Q(\ram[12][235] ) );
  LATCHX1_HVT \ram_reg[12][234]  ( .CLK(n81), .D(N252), .Q(\ram[12][234] ) );
  LATCHX1_HVT \ram_reg[12][233]  ( .CLK(n81), .D(N251), .Q(\ram[12][233] ) );
  LATCHX1_HVT \ram_reg[12][232]  ( .CLK(n81), .D(N250), .Q(\ram[12][232] ) );
  LATCHX1_HVT \ram_reg[12][231]  ( .CLK(n81), .D(N249), .Q(\ram[12][231] ) );
  LATCHX1_HVT \ram_reg[12][230]  ( .CLK(n80), .D(N248), .Q(\ram[12][230] ) );
  LATCHX1_HVT \ram_reg[12][229]  ( .CLK(n80), .D(N247), .Q(\ram[12][229] ) );
  LATCHX1_HVT \ram_reg[12][228]  ( .CLK(n80), .D(N246), .Q(\ram[12][228] ) );
  LATCHX1_HVT \ram_reg[12][227]  ( .CLK(n90), .D(N245), .Q(\ram[12][227] ) );
  LATCHX1_HVT \ram_reg[12][226]  ( .CLK(n90), .D(N244), .Q(\ram[12][226] ) );
  LATCHX1_HVT \ram_reg[12][225]  ( .CLK(n90), .D(N243), .Q(\ram[12][225] ) );
  LATCHX1_HVT \ram_reg[12][224]  ( .CLK(n90), .D(N242), .Q(\ram[12][224] ) );
  LATCHX1_HVT \ram_reg[12][223]  ( .CLK(n90), .D(N241), .Q(\ram[12][223] ) );
  LATCHX1_HVT \ram_reg[12][222]  ( .CLK(n90), .D(N240), .Q(\ram[12][222] ) );
  LATCHX1_HVT \ram_reg[12][221]  ( .CLK(n90), .D(N239), .Q(\ram[12][221] ) );
  LATCHX1_HVT \ram_reg[12][220]  ( .CLK(n90), .D(N238), .Q(\ram[12][220] ) );
  LATCHX1_HVT \ram_reg[12][219]  ( .CLK(n90), .D(N237), .Q(\ram[12][219] ) );
  LATCHX1_HVT \ram_reg[12][218]  ( .CLK(n90), .D(N236), .Q(\ram[12][218] ) );
  LATCHX1_HVT \ram_reg[12][217]  ( .CLK(n89), .D(N235), .Q(\ram[12][217] ) );
  LATCHX1_HVT \ram_reg[12][216]  ( .CLK(n89), .D(N234), .Q(\ram[12][216] ) );
  LATCHX1_HVT \ram_reg[12][215]  ( .CLK(n89), .D(N233), .Q(\ram[12][215] ) );
  LATCHX1_HVT \ram_reg[12][214]  ( .CLK(n89), .D(N232), .Q(\ram[12][214] ) );
  LATCHX1_HVT \ram_reg[12][213]  ( .CLK(n89), .D(N231), .Q(\ram[12][213] ) );
  LATCHX1_HVT \ram_reg[12][212]  ( .CLK(n89), .D(N230), .Q(\ram[12][212] ) );
  LATCHX1_HVT \ram_reg[12][211]  ( .CLK(n89), .D(N229), .Q(\ram[12][211] ) );
  LATCHX1_HVT \ram_reg[12][210]  ( .CLK(n89), .D(N228), .Q(\ram[12][210] ) );
  LATCHX1_HVT \ram_reg[12][209]  ( .CLK(n89), .D(N227), .Q(\ram[12][209] ) );
  LATCHX1_HVT \ram_reg[12][208]  ( .CLK(n89), .D(N226), .Q(\ram[12][208] ) );
  LATCHX1_HVT \ram_reg[12][207]  ( .CLK(n88), .D(N225), .Q(\ram[12][207] ) );
  LATCHX1_HVT \ram_reg[12][206]  ( .CLK(n88), .D(N224), .Q(\ram[12][206] ) );
  LATCHX1_HVT \ram_reg[12][205]  ( .CLK(n88), .D(N223), .Q(\ram[12][205] ) );
  LATCHX1_HVT \ram_reg[12][204]  ( .CLK(n88), .D(N222), .Q(\ram[12][204] ) );
  LATCHX1_HVT \ram_reg[12][203]  ( .CLK(n88), .D(N221), .Q(\ram[12][203] ) );
  LATCHX1_HVT \ram_reg[12][202]  ( .CLK(n88), .D(N220), .Q(\ram[12][202] ) );
  LATCHX1_HVT \ram_reg[12][201]  ( .CLK(n88), .D(N219), .Q(\ram[12][201] ) );
  LATCHX1_HVT \ram_reg[12][200]  ( .CLK(n88), .D(N218), .Q(\ram[12][200] ) );
  LATCHX1_HVT \ram_reg[12][199]  ( .CLK(n88), .D(N217), .Q(\ram[12][199] ) );
  LATCHX1_HVT \ram_reg[12][198]  ( .CLK(n88), .D(N216), .Q(\ram[12][198] ) );
  LATCHX1_HVT \ram_reg[12][197]  ( .CLK(n88), .D(N214), .Q(\ram[12][197] ) );
  LATCHX1_HVT \ram_reg[12][196]  ( .CLK(n87), .D(N213), .Q(\ram[12][196] ) );
  LATCHX1_HVT \ram_reg[12][195]  ( .CLK(n87), .D(N212), .Q(\ram[12][195] ) );
  LATCHX1_HVT \ram_reg[12][194]  ( .CLK(n87), .D(N211), .Q(\ram[12][194] ) );
  LATCHX1_HVT \ram_reg[12][193]  ( .CLK(n87), .D(N210), .Q(\ram[12][193] ) );
  LATCHX1_HVT \ram_reg[12][192]  ( .CLK(n87), .D(N209), .Q(\ram[12][192] ) );
  LATCHX1_HVT \ram_reg[12][191]  ( .CLK(n87), .D(N208), .Q(\ram[12][191] ) );
  LATCHX1_HVT \ram_reg[12][190]  ( .CLK(n87), .D(N207), .Q(\ram[12][190] ) );
  LATCHX1_HVT \ram_reg[12][189]  ( .CLK(n87), .D(N206), .Q(\ram[12][189] ) );
  LATCHX1_HVT \ram_reg[12][188]  ( .CLK(n87), .D(N205), .Q(\ram[12][188] ) );
  LATCHX1_HVT \ram_reg[12][187]  ( .CLK(n87), .D(N204), .Q(\ram[12][187] ) );
  LATCHX1_HVT \ram_reg[12][186]  ( .CLK(n87), .D(N203), .Q(\ram[12][186] ) );
  LATCHX1_HVT \ram_reg[12][185]  ( .CLK(n86), .D(N202), .Q(\ram[12][185] ) );
  LATCHX1_HVT \ram_reg[12][184]  ( .CLK(n86), .D(N201), .Q(\ram[12][184] ) );
  LATCHX1_HVT \ram_reg[12][183]  ( .CLK(n86), .D(N200), .Q(\ram[12][183] ) );
  LATCHX1_HVT \ram_reg[12][182]  ( .CLK(n86), .D(N199), .Q(\ram[12][182] ) );
  LATCHX1_HVT \ram_reg[12][181]  ( .CLK(n86), .D(N198), .Q(\ram[12][181] ) );
  LATCHX1_HVT \ram_reg[12][180]  ( .CLK(n86), .D(N197), .Q(\ram[12][180] ) );
  LATCHX1_HVT \ram_reg[12][179]  ( .CLK(n86), .D(N196), .Q(\ram[12][179] ) );
  LATCHX1_HVT \ram_reg[12][178]  ( .CLK(n86), .D(N195), .Q(\ram[12][178] ) );
  LATCHX1_HVT \ram_reg[12][177]  ( .CLK(n86), .D(N194), .Q(\ram[12][177] ) );
  LATCHX1_HVT \ram_reg[12][176]  ( .CLK(n86), .D(N193), .Q(\ram[12][176] ) );
  LATCHX1_HVT \ram_reg[12][175]  ( .CLK(n86), .D(N192), .Q(\ram[12][175] ) );
  LATCHX1_HVT \ram_reg[12][174]  ( .CLK(n85), .D(N191), .Q(\ram[12][174] ) );
  LATCHX1_HVT \ram_reg[12][173]  ( .CLK(n85), .D(N190), .Q(\ram[12][173] ) );
  LATCHX1_HVT \ram_reg[12][172]  ( .CLK(n85), .D(N189), .Q(\ram[12][172] ) );
  LATCHX1_HVT \ram_reg[12][171]  ( .CLK(n85), .D(N188), .Q(\ram[12][171] ) );
  LATCHX1_HVT \ram_reg[12][170]  ( .CLK(n85), .D(N187), .Q(\ram[12][170] ) );
  LATCHX1_HVT \ram_reg[12][169]  ( .CLK(n85), .D(N186), .Q(\ram[12][169] ) );
  LATCHX1_HVT \ram_reg[12][168]  ( .CLK(n85), .D(N185), .Q(\ram[12][168] ) );
  LATCHX1_HVT \ram_reg[12][167]  ( .CLK(n85), .D(N184), .Q(\ram[12][167] ) );
  LATCHX1_HVT \ram_reg[12][166]  ( .CLK(n85), .D(N183), .Q(\ram[12][166] ) );
  LATCHX1_HVT \ram_reg[12][165]  ( .CLK(n85), .D(N182), .Q(\ram[12][165] ) );
  LATCHX1_HVT \ram_reg[12][164]  ( .CLK(n85), .D(N181), .Q(\ram[12][164] ) );
  LATCHX1_HVT \ram_reg[12][163]  ( .CLK(n84), .D(N180), .Q(\ram[12][163] ) );
  LATCHX1_HVT \ram_reg[12][162]  ( .CLK(n84), .D(N179), .Q(\ram[12][162] ) );
  LATCHX1_HVT \ram_reg[12][161]  ( .CLK(n84), .D(N178), .Q(\ram[12][161] ) );
  LATCHX1_HVT \ram_reg[12][160]  ( .CLK(n84), .D(N177), .Q(\ram[12][160] ) );
  LATCHX1_HVT \ram_reg[12][159]  ( .CLK(n84), .D(N176), .Q(\ram[12][159] ) );
  LATCHX1_HVT \ram_reg[12][158]  ( .CLK(n84), .D(N175), .Q(\ram[12][158] ) );
  LATCHX1_HVT \ram_reg[12][157]  ( .CLK(n84), .D(N174), .Q(\ram[12][157] ) );
  LATCHX1_HVT \ram_reg[12][156]  ( .CLK(n84), .D(N173), .Q(\ram[12][156] ) );
  LATCHX1_HVT \ram_reg[12][155]  ( .CLK(n84), .D(N172), .Q(\ram[12][155] ) );
  LATCHX1_HVT \ram_reg[12][154]  ( .CLK(n84), .D(N171), .Q(\ram[12][154] ) );
  LATCHX1_HVT \ram_reg[12][153]  ( .CLK(n84), .D(N170), .Q(\ram[12][153] ) );
  LATCHX1_HVT \ram_reg[12][152]  ( .CLK(n83), .D(N169), .Q(\ram[12][152] ) );
  LATCHX1_HVT \ram_reg[12][151]  ( .CLK(n83), .D(N168), .Q(\ram[12][151] ) );
  LATCHX1_HVT \ram_reg[12][150]  ( .CLK(n83), .D(N167), .Q(\ram[12][150] ) );
  LATCHX1_HVT \ram_reg[12][149]  ( .CLK(n83), .D(N166), .Q(\ram[12][149] ) );
  LATCHX1_HVT \ram_reg[12][148]  ( .CLK(n83), .D(N165), .Q(\ram[12][148] ) );
  LATCHX1_HVT \ram_reg[12][147]  ( .CLK(n83), .D(N164), .Q(\ram[12][147] ) );
  LATCHX1_HVT \ram_reg[12][146]  ( .CLK(n83), .D(N163), .Q(\ram[12][146] ) );
  LATCHX1_HVT \ram_reg[12][145]  ( .CLK(n83), .D(N162), .Q(\ram[12][145] ) );
  LATCHX1_HVT \ram_reg[12][144]  ( .CLK(n83), .D(N161), .Q(\ram[12][144] ) );
  LATCHX1_HVT \ram_reg[12][143]  ( .CLK(n83), .D(N160), .Q(\ram[12][143] ) );
  LATCHX1_HVT \ram_reg[12][142]  ( .CLK(n83), .D(N159), .Q(\ram[12][142] ) );
  LATCHX1_HVT \ram_reg[12][141]  ( .CLK(n82), .D(N158), .Q(\ram[12][141] ) );
  LATCHX1_HVT \ram_reg[12][140]  ( .CLK(n82), .D(N157), .Q(\ram[12][140] ) );
  LATCHX1_HVT \ram_reg[12][139]  ( .CLK(n82), .D(N156), .Q(\ram[12][139] ) );
  LATCHX1_HVT \ram_reg[12][138]  ( .CLK(n81), .D(N155), .Q(\ram[12][138] ) );
  LATCHX1_HVT \ram_reg[12][137]  ( .CLK(n90), .D(N154), .Q(\ram[12][137] ) );
  LATCHX1_HVT \ram_reg[12][136]  ( .CLK(n89), .D(N153), .Q(\ram[12][136] ) );
  LATCHX1_HVT \ram_reg[12][135]  ( .CLK(n89), .D(N152), .Q(\ram[12][135] ) );
  LATCHX1_HVT \ram_reg[12][134]  ( .CLK(n88), .D(N151), .Q(\ram[12][134] ) );
  LATCHX1_HVT \ram_reg[12][133]  ( .CLK(n87), .D(N150), .Q(\ram[12][133] ) );
  LATCHX1_HVT \ram_reg[12][132]  ( .CLK(n86), .D(N149), .Q(\ram[12][132] ) );
  LATCHX1_HVT \ram_reg[12][131]  ( .CLK(n85), .D(N148), .Q(\ram[12][131] ) );
  LATCHX1_HVT \ram_reg[12][130]  ( .CLK(n84), .D(N147), .Q(\ram[12][130] ) );
  LATCHX1_HVT \ram_reg[12][129]  ( .CLK(n83), .D(N146), .Q(\ram[12][129] ) );
  LATCHX1_HVT \ram_reg[12][128]  ( .CLK(n80), .D(N145), .Q(\ram[12][128] ) );
  LATCHX1_HVT \ram_reg[12][127]  ( .CLK(n71), .D(N144), .Q(\ram[12][127] ) );
  LATCHX1_HVT \ram_reg[12][126]  ( .CLK(n71), .D(N143), .Q(\ram[12][126] ) );
  LATCHX1_HVT \ram_reg[12][125]  ( .CLK(n71), .D(N142), .Q(\ram[12][125] ) );
  LATCHX1_HVT \ram_reg[12][124]  ( .CLK(n71), .D(N141), .Q(\ram[12][124] ) );
  LATCHX1_HVT \ram_reg[12][123]  ( .CLK(n71), .D(N140), .Q(\ram[12][123] ) );
  LATCHX1_HVT \ram_reg[12][122]  ( .CLK(n70), .D(N139), .Q(\ram[12][122] ) );
  LATCHX1_HVT \ram_reg[12][121]  ( .CLK(n71), .D(N138), .Q(\ram[12][121] ) );
  LATCHX1_HVT \ram_reg[12][120]  ( .CLK(n71), .D(N137), .Q(\ram[12][120] ) );
  LATCHX1_HVT \ram_reg[12][119]  ( .CLK(n80), .D(N136), .Q(\ram[12][119] ) );
  LATCHX1_HVT \ram_reg[12][118]  ( .CLK(n79), .D(N135), .Q(\ram[12][118] ) );
  LATCHX1_HVT \ram_reg[12][117]  ( .CLK(n79), .D(N134), .Q(\ram[12][117] ) );
  LATCHX1_HVT \ram_reg[12][116]  ( .CLK(n78), .D(N133), .Q(\ram[12][116] ) );
  LATCHX1_HVT \ram_reg[12][115]  ( .CLK(n73), .D(N132), .Q(\ram[12][115] ) );
  LATCHX1_HVT \ram_reg[12][114]  ( .CLK(n78), .D(N131), .Q(\ram[12][114] ) );
  LATCHX1_HVT \ram_reg[12][113]  ( .CLK(n78), .D(N130), .Q(\ram[12][113] ) );
  LATCHX1_HVT \ram_reg[12][112]  ( .CLK(n79), .D(N129), .Q(\ram[12][112] ) );
  LATCHX1_HVT \ram_reg[12][111]  ( .CLK(n77), .D(N128), .Q(\ram[12][111] ) );
  LATCHX1_HVT \ram_reg[12][110]  ( .CLK(n77), .D(N127), .Q(\ram[12][110] ) );
  LATCHX1_HVT \ram_reg[12][109]  ( .CLK(n77), .D(N126), .Q(\ram[12][109] ) );
  LATCHX1_HVT \ram_reg[12][108]  ( .CLK(n74), .D(N125), .Q(\ram[12][108] ) );
  LATCHX1_HVT \ram_reg[12][107]  ( .CLK(n71), .D(N124), .Q(\ram[12][107] ) );
  LATCHX1_HVT \ram_reg[12][106]  ( .CLK(n77), .D(N123), .Q(\ram[12][106] ) );
  LATCHX1_HVT \ram_reg[12][105]  ( .CLK(n77), .D(N122), .Q(\ram[12][105] ) );
  LATCHX1_HVT \ram_reg[12][104]  ( .CLK(n77), .D(N121), .Q(\ram[12][104] ) );
  LATCHX1_HVT \ram_reg[12][103]  ( .CLK(n76), .D(N120), .Q(\ram[12][103] ) );
  LATCHX1_HVT \ram_reg[12][102]  ( .CLK(n75), .D(N119), .Q(\ram[12][102] ) );
  LATCHX1_HVT \ram_reg[12][101]  ( .CLK(n75), .D(N118), .Q(\ram[12][101] ) );
  LATCHX1_HVT \ram_reg[12][100]  ( .CLK(n76), .D(N117), .Q(\ram[12][100] ) );
  LATCHX1_HVT \ram_reg[12][99]  ( .CLK(n74), .D(N116), .Q(\ram[12][99] ) );
  LATCHX1_HVT \ram_reg[12][98]  ( .CLK(n75), .D(N114), .Q(\ram[12][98] ) );
  LATCHX1_HVT \ram_reg[12][97]  ( .CLK(n76), .D(N113), .Q(\ram[12][97] ) );
  LATCHX1_HVT \ram_reg[12][96]  ( .CLK(n80), .D(N112), .Q(\ram[12][96] ) );
  LATCHX1_HVT \ram_reg[12][95]  ( .CLK(n72), .D(N111), .Q(\ram[12][95] ) );
  LATCHX1_HVT \ram_reg[12][94]  ( .CLK(n72), .D(N110), .Q(\ram[12][94] ) );
  LATCHX1_HVT \ram_reg[12][93]  ( .CLK(n72), .D(N109), .Q(\ram[12][93] ) );
  LATCHX1_HVT \ram_reg[12][92]  ( .CLK(n71), .D(N108), .Q(\ram[12][92] ) );
  LATCHX1_HVT \ram_reg[12][91]  ( .CLK(n71), .D(N107), .Q(\ram[12][91] ) );
  LATCHX1_HVT \ram_reg[12][90]  ( .CLK(n72), .D(N106), .Q(\ram[12][90] ) );
  LATCHX1_HVT \ram_reg[12][89]  ( .CLK(n71), .D(N105), .Q(\ram[12][89] ) );
  LATCHX1_HVT \ram_reg[12][88]  ( .CLK(n72), .D(N104), .Q(\ram[12][88] ) );
  LATCHX1_HVT \ram_reg[12][87]  ( .CLK(n80), .D(N103), .Q(\ram[12][87] ) );
  LATCHX1_HVT \ram_reg[12][86]  ( .CLK(n79), .D(N102), .Q(\ram[12][86] ) );
  LATCHX1_HVT \ram_reg[12][85]  ( .CLK(n78), .D(N101), .Q(\ram[12][85] ) );
  LATCHX1_HVT \ram_reg[12][84]  ( .CLK(n78), .D(N100), .Q(\ram[12][84] ) );
  LATCHX1_HVT \ram_reg[12][83]  ( .CLK(n73), .D(N99), .Q(\ram[12][83] ) );
  LATCHX1_HVT \ram_reg[12][82]  ( .CLK(n79), .D(N98), .Q(\ram[12][82] ) );
  LATCHX1_HVT \ram_reg[12][81]  ( .CLK(n78), .D(N97), .Q(\ram[12][81] ) );
  LATCHX1_HVT \ram_reg[12][80]  ( .CLK(n79), .D(N96), .Q(\ram[12][80] ) );
  LATCHX1_HVT \ram_reg[12][79]  ( .CLK(n73), .D(N95), .Q(\ram[12][79] ) );
  LATCHX1_HVT \ram_reg[12][78]  ( .CLK(n72), .D(N94), .Q(\ram[12][78] ) );
  LATCHX1_HVT \ram_reg[12][77]  ( .CLK(n73), .D(N93), .Q(\ram[12][77] ) );
  LATCHX1_HVT \ram_reg[12][76]  ( .CLK(n72), .D(N92), .Q(\ram[12][76] ) );
  LATCHX1_HVT \ram_reg[12][75]  ( .CLK(n72), .D(N91), .Q(\ram[12][75] ) );
  LATCHX1_HVT \ram_reg[12][74]  ( .CLK(n70), .D(N90), .Q(\ram[12][74] ) );
  LATCHX1_HVT \ram_reg[12][73]  ( .CLK(n73), .D(N89), .Q(\ram[12][73] ) );
  LATCHX1_HVT \ram_reg[12][72]  ( .CLK(n73), .D(N88), .Q(\ram[12][72] ) );
  LATCHX1_HVT \ram_reg[12][71]  ( .CLK(n76), .D(N87), .Q(\ram[12][71] ) );
  LATCHX1_HVT \ram_reg[12][70]  ( .CLK(n76), .D(N86), .Q(\ram[12][70] ) );
  LATCHX1_HVT \ram_reg[12][69]  ( .CLK(n75), .D(N85), .Q(\ram[12][69] ) );
  LATCHX1_HVT \ram_reg[12][68]  ( .CLK(n76), .D(N84), .Q(\ram[12][68] ) );
  LATCHX1_HVT \ram_reg[12][67]  ( .CLK(n75), .D(N83), .Q(\ram[12][67] ) );
  LATCHX1_HVT \ram_reg[12][66]  ( .CLK(n74), .D(N82), .Q(\ram[12][66] ) );
  LATCHX1_HVT \ram_reg[12][65]  ( .CLK(n75), .D(N81), .Q(\ram[12][65] ) );
  LATCHX1_HVT \ram_reg[12][64]  ( .CLK(n80), .D(N80), .Q(\ram[12][64] ) );
  LATCHX1_HVT \ram_reg[12][63]  ( .CLK(n74), .D(N79), .Q(\ram[12][63] ) );
  LATCHX1_HVT \ram_reg[12][62]  ( .CLK(n74), .D(N78), .Q(\ram[12][62] ) );
  LATCHX1_HVT \ram_reg[12][61]  ( .CLK(n74), .D(N77), .Q(\ram[12][61] ) );
  LATCHX1_HVT \ram_reg[12][60]  ( .CLK(n74), .D(N76), .Q(\ram[12][60] ) );
  LATCHX1_HVT \ram_reg[12][59]  ( .CLK(n74), .D(N75), .Q(\ram[12][59] ) );
  LATCHX1_HVT \ram_reg[12][58]  ( .CLK(n73), .D(N74), .Q(\ram[12][58] ) );
  LATCHX1_HVT \ram_reg[12][57]  ( .CLK(n74), .D(N73), .Q(\ram[12][57] ) );
  LATCHX1_HVT \ram_reg[12][56]  ( .CLK(n74), .D(N72), .Q(\ram[12][56] ) );
  LATCHX1_HVT \ram_reg[12][55]  ( .CLK(n80), .D(N71), .Q(\ram[12][55] ) );
  LATCHX1_HVT \ram_reg[12][54]  ( .CLK(n78), .D(N70), .Q(\ram[12][54] ) );
  LATCHX1_HVT \ram_reg[12][53]  ( .CLK(n78), .D(N69), .Q(\ram[12][53] ) );
  LATCHX1_HVT \ram_reg[12][52]  ( .CLK(n79), .D(N68), .Q(\ram[12][52] ) );
  LATCHX1_HVT \ram_reg[12][51]  ( .CLK(n73), .D(N67), .Q(\ram[12][51] ) );
  LATCHX1_HVT \ram_reg[12][50]  ( .CLK(n70), .D(N66), .Q(\ram[12][50] ) );
  LATCHX1_HVT \ram_reg[12][49]  ( .CLK(n79), .D(N65), .Q(\ram[12][49] ) );
  LATCHX1_HVT \ram_reg[12][48]  ( .CLK(n79), .D(N64), .Q(\ram[12][48] ) );
  LATCHX1_HVT \ram_reg[12][47]  ( .CLK(n77), .D(N63), .Q(\ram[12][47] ) );
  LATCHX1_HVT \ram_reg[12][46]  ( .CLK(n77), .D(N62), .Q(\ram[12][46] ) );
  LATCHX1_HVT \ram_reg[12][45]  ( .CLK(n77), .D(N61), .Q(\ram[12][45] ) );
  LATCHX1_HVT \ram_reg[12][44]  ( .CLK(n77), .D(N60), .Q(\ram[12][44] ) );
  LATCHX1_HVT \ram_reg[12][43]  ( .CLK(n74), .D(N59), .Q(\ram[12][43] ) );
  LATCHX1_HVT \ram_reg[12][42]  ( .CLK(n78), .D(N58), .Q(\ram[12][42] ) );
  LATCHX1_HVT \ram_reg[12][41]  ( .CLK(n71), .D(N57), .Q(\ram[12][41] ) );
  LATCHX1_HVT \ram_reg[12][40]  ( .CLK(n77), .D(N56), .Q(\ram[12][40] ) );
  LATCHX1_HVT \ram_reg[12][39]  ( .CLK(n76), .D(N55), .Q(\ram[12][39] ) );
  LATCHX1_HVT \ram_reg[12][38]  ( .CLK(n76), .D(N54), .Q(\ram[12][38] ) );
  LATCHX1_HVT \ram_reg[12][37]  ( .CLK(n75), .D(N53), .Q(\ram[12][37] ) );
  LATCHX1_HVT \ram_reg[12][36]  ( .CLK(n75), .D(N52), .Q(\ram[12][36] ) );
  LATCHX1_HVT \ram_reg[12][35]  ( .CLK(n75), .D(N51), .Q(\ram[12][35] ) );
  LATCHX1_HVT \ram_reg[12][34]  ( .CLK(n77), .D(N50), .Q(\ram[12][34] ) );
  LATCHX1_HVT \ram_reg[12][33]  ( .CLK(n76), .D(N49), .Q(\ram[12][33] ) );
  LATCHX1_HVT \ram_reg[12][32]  ( .CLK(n80), .D(N48), .Q(\ram[12][32] ) );
  LATCHX1_HVT \ram_reg[12][31]  ( .CLK(n70), .D(N47), .Q(\ram[12][31] ) );
  LATCHX1_HVT \ram_reg[12][30]  ( .CLK(n70), .D(N46), .Q(\ram[12][30] ) );
  LATCHX1_HVT \ram_reg[12][29]  ( .CLK(n70), .D(N45), .Q(\ram[12][29] ) );
  LATCHX1_HVT \ram_reg[12][28]  ( .CLK(n70), .D(N44), .Q(\ram[12][28] ) );
  LATCHX1_HVT \ram_reg[12][27]  ( .CLK(n70), .D(N43), .Q(\ram[12][27] ) );
  LATCHX1_HVT \ram_reg[12][26]  ( .CLK(n70), .D(N42), .Q(\ram[12][26] ) );
  LATCHX1_HVT \ram_reg[12][25]  ( .CLK(n70), .D(N41), .Q(\ram[12][25] ) );
  LATCHX1_HVT \ram_reg[12][24]  ( .CLK(n70), .D(N40), .Q(\ram[12][24] ) );
  LATCHX1_HVT \ram_reg[12][23]  ( .CLK(n80), .D(N39), .Q(\ram[12][23] ) );
  LATCHX1_HVT \ram_reg[12][22]  ( .CLK(n79), .D(N38), .Q(\ram[12][22] ) );
  LATCHX1_HVT \ram_reg[12][21]  ( .CLK(n78), .D(N37), .Q(\ram[12][21] ) );
  LATCHX1_HVT \ram_reg[12][20]  ( .CLK(n78), .D(N36), .Q(\ram[12][20] ) );
  LATCHX1_HVT \ram_reg[12][19]  ( .CLK(n70), .D(N35), .Q(\ram[12][19] ) );
  LATCHX1_HVT \ram_reg[12][18]  ( .CLK(n78), .D(N34), .Q(\ram[12][18] ) );
  LATCHX1_HVT \ram_reg[12][17]  ( .CLK(n79), .D(N33), .Q(\ram[12][17] ) );
  LATCHX1_HVT \ram_reg[12][16]  ( .CLK(n79), .D(N32), .Q(\ram[12][16] ) );
  LATCHX1_HVT \ram_reg[12][15]  ( .CLK(n73), .D(N31), .Q(\ram[12][15] ) );
  LATCHX1_HVT \ram_reg[12][14]  ( .CLK(n73), .D(N30), .Q(\ram[12][14] ) );
  LATCHX1_HVT \ram_reg[12][13]  ( .CLK(n72), .D(N29), .Q(\ram[12][13] ) );
  LATCHX1_HVT \ram_reg[12][12]  ( .CLK(n72), .D(N28), .Q(\ram[12][12] ) );
  LATCHX1_HVT \ram_reg[12][11]  ( .CLK(n73), .D(N27), .Q(\ram[12][11] ) );
  LATCHX1_HVT \ram_reg[12][10]  ( .CLK(n72), .D(N26), .Q(\ram[12][10] ) );
  LATCHX1_HVT \ram_reg[12][9]  ( .CLK(n72), .D(N25), .Q(\ram[12][9] ) );
  LATCHX1_HVT \ram_reg[12][8]  ( .CLK(n73), .D(N24), .Q(\ram[12][8] ) );
  LATCHX1_HVT \ram_reg[12][7]  ( .CLK(n76), .D(N23), .Q(\ram[12][7] ) );
  LATCHX1_HVT \ram_reg[12][6]  ( .CLK(n76), .D(N22), .Q(\ram[12][6] ) );
  LATCHX1_HVT \ram_reg[12][5]  ( .CLK(n75), .D(N21), .Q(\ram[12][5] ) );
  LATCHX1_HVT \ram_reg[12][4]  ( .CLK(n75), .D(N20), .Q(\ram[12][4] ) );
  LATCHX1_HVT \ram_reg[12][3]  ( .CLK(n74), .D(N19), .Q(\ram[12][3] ) );
  LATCHX1_HVT \ram_reg[12][2]  ( .CLK(n75), .D(N18), .Q(\ram[12][2] ) );
  LATCHX1_HVT \ram_reg[12][1]  ( .CLK(n76), .D(N17), .Q(\ram[12][1] ) );
  LATCHX1_HVT \ram_reg[12][0]  ( .CLK(n80), .D(N16), .Q(\ram[12][0] ) );
  LATCHX1_HVT \ram_reg[11][255]  ( .CLK(n93), .D(N273), .Q(\ram[11][255] ) );
  LATCHX1_HVT \ram_reg[11][254]  ( .CLK(N306), .D(N272), .Q(\ram[11][254] ) );
  LATCHX1_HVT \ram_reg[11][253]  ( .CLK(N306), .D(N271), .Q(\ram[11][253] ) );
  LATCHX1_HVT \ram_reg[11][252]  ( .CLK(N306), .D(N270), .Q(\ram[11][252] ) );
  LATCHX1_HVT \ram_reg[11][251]  ( .CLK(N306), .D(N269), .Q(\ram[11][251] ) );
  LATCHX1_HVT \ram_reg[11][250]  ( .CLK(n105), .D(N268), .Q(\ram[11][250] ) );
  LATCHX1_HVT \ram_reg[11][249]  ( .CLK(n105), .D(N267), .Q(\ram[11][249] ) );
  LATCHX1_HVT \ram_reg[11][248]  ( .CLK(n105), .D(N266), .Q(\ram[11][248] ) );
  LATCHX1_HVT \ram_reg[11][247]  ( .CLK(n105), .D(N265), .Q(\ram[11][247] ) );
  LATCHX1_HVT \ram_reg[11][246]  ( .CLK(n105), .D(N264), .Q(\ram[11][246] ) );
  LATCHX1_HVT \ram_reg[11][245]  ( .CLK(n105), .D(N263), .Q(\ram[11][245] ) );
  LATCHX1_HVT \ram_reg[11][244]  ( .CLK(n105), .D(N262), .Q(\ram[11][244] ) );
  LATCHX1_HVT \ram_reg[11][243]  ( .CLK(n105), .D(N261), .Q(\ram[11][243] ) );
  LATCHX1_HVT \ram_reg[11][242]  ( .CLK(n105), .D(N260), .Q(\ram[11][242] ) );
  LATCHX1_HVT \ram_reg[11][241]  ( .CLK(n105), .D(N259), .Q(\ram[11][241] ) );
  LATCHX1_HVT \ram_reg[11][240]  ( .CLK(n104), .D(N258), .Q(\ram[11][240] ) );
  LATCHX1_HVT \ram_reg[11][239]  ( .CLK(n104), .D(N257), .Q(\ram[11][239] ) );
  LATCHX1_HVT \ram_reg[11][238]  ( .CLK(n104), .D(N256), .Q(\ram[11][238] ) );
  LATCHX1_HVT \ram_reg[11][237]  ( .CLK(n104), .D(N255), .Q(\ram[11][237] ) );
  LATCHX1_HVT \ram_reg[11][236]  ( .CLK(n104), .D(N254), .Q(\ram[11][236] ) );
  LATCHX1_HVT \ram_reg[11][235]  ( .CLK(n104), .D(N253), .Q(\ram[11][235] ) );
  LATCHX1_HVT \ram_reg[11][234]  ( .CLK(n104), .D(N252), .Q(\ram[11][234] ) );
  LATCHX1_HVT \ram_reg[11][233]  ( .CLK(n104), .D(N251), .Q(\ram[11][233] ) );
  LATCHX1_HVT \ram_reg[11][232]  ( .CLK(n104), .D(N250), .Q(\ram[11][232] ) );
  LATCHX1_HVT \ram_reg[11][231]  ( .CLK(n104), .D(N249), .Q(\ram[11][231] ) );
  LATCHX1_HVT \ram_reg[11][230]  ( .CLK(n104), .D(N248), .Q(\ram[11][230] ) );
  LATCHX1_HVT \ram_reg[11][229]  ( .CLK(n103), .D(N247), .Q(\ram[11][229] ) );
  LATCHX1_HVT \ram_reg[11][228]  ( .CLK(n103), .D(N246), .Q(\ram[11][228] ) );
  LATCHX1_HVT \ram_reg[11][227]  ( .CLK(n113), .D(N245), .Q(\ram[11][227] ) );
  LATCHX1_HVT \ram_reg[11][226]  ( .CLK(n113), .D(N244), .Q(\ram[11][226] ) );
  LATCHX1_HVT \ram_reg[11][225]  ( .CLK(n113), .D(N243), .Q(\ram[11][225] ) );
  LATCHX1_HVT \ram_reg[11][224]  ( .CLK(n113), .D(N242), .Q(\ram[11][224] ) );
  LATCHX1_HVT \ram_reg[11][223]  ( .CLK(n113), .D(N241), .Q(\ram[11][223] ) );
  LATCHX1_HVT \ram_reg[11][222]  ( .CLK(n113), .D(N240), .Q(\ram[11][222] ) );
  LATCHX1_HVT \ram_reg[11][221]  ( .CLK(n113), .D(N239), .Q(\ram[11][221] ) );
  LATCHX1_HVT \ram_reg[11][220]  ( .CLK(n113), .D(N238), .Q(\ram[11][220] ) );
  LATCHX1_HVT \ram_reg[11][219]  ( .CLK(n113), .D(N237), .Q(\ram[11][219] ) );
  LATCHX1_HVT \ram_reg[11][218]  ( .CLK(n113), .D(N236), .Q(\ram[11][218] ) );
  LATCHX1_HVT \ram_reg[11][217]  ( .CLK(n112), .D(N235), .Q(\ram[11][217] ) );
  LATCHX1_HVT \ram_reg[11][216]  ( .CLK(n112), .D(N234), .Q(\ram[11][216] ) );
  LATCHX1_HVT \ram_reg[11][215]  ( .CLK(n112), .D(N233), .Q(\ram[11][215] ) );
  LATCHX1_HVT \ram_reg[11][214]  ( .CLK(n112), .D(N232), .Q(\ram[11][214] ) );
  LATCHX1_HVT \ram_reg[11][213]  ( .CLK(n112), .D(N231), .Q(\ram[11][213] ) );
  LATCHX1_HVT \ram_reg[11][212]  ( .CLK(n112), .D(N230), .Q(\ram[11][212] ) );
  LATCHX1_HVT \ram_reg[11][211]  ( .CLK(n112), .D(N229), .Q(\ram[11][211] ) );
  LATCHX1_HVT \ram_reg[11][210]  ( .CLK(n112), .D(N228), .Q(\ram[11][210] ) );
  LATCHX1_HVT \ram_reg[11][209]  ( .CLK(n112), .D(N227), .Q(\ram[11][209] ) );
  LATCHX1_HVT \ram_reg[11][208]  ( .CLK(n112), .D(N226), .Q(\ram[11][208] ) );
  LATCHX1_HVT \ram_reg[11][207]  ( .CLK(n112), .D(N225), .Q(\ram[11][207] ) );
  LATCHX1_HVT \ram_reg[11][206]  ( .CLK(n111), .D(N224), .Q(\ram[11][206] ) );
  LATCHX1_HVT \ram_reg[11][205]  ( .CLK(n111), .D(N223), .Q(\ram[11][205] ) );
  LATCHX1_HVT \ram_reg[11][204]  ( .CLK(n111), .D(N222), .Q(\ram[11][204] ) );
  LATCHX1_HVT \ram_reg[11][203]  ( .CLK(n111), .D(N221), .Q(\ram[11][203] ) );
  LATCHX1_HVT \ram_reg[11][202]  ( .CLK(n111), .D(N220), .Q(\ram[11][202] ) );
  LATCHX1_HVT \ram_reg[11][201]  ( .CLK(n111), .D(N219), .Q(\ram[11][201] ) );
  LATCHX1_HVT \ram_reg[11][200]  ( .CLK(n111), .D(N218), .Q(\ram[11][200] ) );
  LATCHX1_HVT \ram_reg[11][199]  ( .CLK(n111), .D(N217), .Q(\ram[11][199] ) );
  LATCHX1_HVT \ram_reg[11][198]  ( .CLK(n111), .D(N216), .Q(\ram[11][198] ) );
  LATCHX1_HVT \ram_reg[11][197]  ( .CLK(n111), .D(N214), .Q(\ram[11][197] ) );
  LATCHX1_HVT \ram_reg[11][196]  ( .CLK(n111), .D(N213), .Q(\ram[11][196] ) );
  LATCHX1_HVT \ram_reg[11][195]  ( .CLK(n110), .D(N212), .Q(\ram[11][195] ) );
  LATCHX1_HVT \ram_reg[11][194]  ( .CLK(n110), .D(N211), .Q(\ram[11][194] ) );
  LATCHX1_HVT \ram_reg[11][193]  ( .CLK(n110), .D(N210), .Q(\ram[11][193] ) );
  LATCHX1_HVT \ram_reg[11][192]  ( .CLK(n110), .D(N209), .Q(\ram[11][192] ) );
  LATCHX1_HVT \ram_reg[11][191]  ( .CLK(n110), .D(N208), .Q(\ram[11][191] ) );
  LATCHX1_HVT \ram_reg[11][190]  ( .CLK(n110), .D(N207), .Q(\ram[11][190] ) );
  LATCHX1_HVT \ram_reg[11][189]  ( .CLK(n110), .D(N206), .Q(\ram[11][189] ) );
  LATCHX1_HVT \ram_reg[11][188]  ( .CLK(n110), .D(N205), .Q(\ram[11][188] ) );
  LATCHX1_HVT \ram_reg[11][187]  ( .CLK(n110), .D(N204), .Q(\ram[11][187] ) );
  LATCHX1_HVT \ram_reg[11][186]  ( .CLK(n110), .D(N203), .Q(\ram[11][186] ) );
  LATCHX1_HVT \ram_reg[11][185]  ( .CLK(n110), .D(N202), .Q(\ram[11][185] ) );
  LATCHX1_HVT \ram_reg[11][184]  ( .CLK(n109), .D(N201), .Q(\ram[11][184] ) );
  LATCHX1_HVT \ram_reg[11][183]  ( .CLK(n109), .D(N200), .Q(\ram[11][183] ) );
  LATCHX1_HVT \ram_reg[11][182]  ( .CLK(n109), .D(N199), .Q(\ram[11][182] ) );
  LATCHX1_HVT \ram_reg[11][181]  ( .CLK(n109), .D(N198), .Q(\ram[11][181] ) );
  LATCHX1_HVT \ram_reg[11][180]  ( .CLK(n109), .D(N197), .Q(\ram[11][180] ) );
  LATCHX1_HVT \ram_reg[11][179]  ( .CLK(n109), .D(N196), .Q(\ram[11][179] ) );
  LATCHX1_HVT \ram_reg[11][178]  ( .CLK(n109), .D(N195), .Q(\ram[11][178] ) );
  LATCHX1_HVT \ram_reg[11][177]  ( .CLK(n109), .D(N194), .Q(\ram[11][177] ) );
  LATCHX1_HVT \ram_reg[11][176]  ( .CLK(n109), .D(N193), .Q(\ram[11][176] ) );
  LATCHX1_HVT \ram_reg[11][175]  ( .CLK(n109), .D(N192), .Q(\ram[11][175] ) );
  LATCHX1_HVT \ram_reg[11][174]  ( .CLK(n109), .D(N191), .Q(\ram[11][174] ) );
  LATCHX1_HVT \ram_reg[11][173]  ( .CLK(n108), .D(N190), .Q(\ram[11][173] ) );
  LATCHX1_HVT \ram_reg[11][172]  ( .CLK(n108), .D(N189), .Q(\ram[11][172] ) );
  LATCHX1_HVT \ram_reg[11][171]  ( .CLK(n108), .D(N188), .Q(\ram[11][171] ) );
  LATCHX1_HVT \ram_reg[11][170]  ( .CLK(n108), .D(N187), .Q(\ram[11][170] ) );
  LATCHX1_HVT \ram_reg[11][169]  ( .CLK(n108), .D(N186), .Q(\ram[11][169] ) );
  LATCHX1_HVT \ram_reg[11][168]  ( .CLK(n108), .D(N185), .Q(\ram[11][168] ) );
  LATCHX1_HVT \ram_reg[11][167]  ( .CLK(n108), .D(N184), .Q(\ram[11][167] ) );
  LATCHX1_HVT \ram_reg[11][166]  ( .CLK(n108), .D(N183), .Q(\ram[11][166] ) );
  LATCHX1_HVT \ram_reg[11][165]  ( .CLK(n108), .D(N182), .Q(\ram[11][165] ) );
  LATCHX1_HVT \ram_reg[11][164]  ( .CLK(n108), .D(N181), .Q(\ram[11][164] ) );
  LATCHX1_HVT \ram_reg[11][163]  ( .CLK(n108), .D(N180), .Q(\ram[11][163] ) );
  LATCHX1_HVT \ram_reg[11][162]  ( .CLK(n107), .D(N179), .Q(\ram[11][162] ) );
  LATCHX1_HVT \ram_reg[11][161]  ( .CLK(n107), .D(N178), .Q(\ram[11][161] ) );
  LATCHX1_HVT \ram_reg[11][160]  ( .CLK(n107), .D(N177), .Q(\ram[11][160] ) );
  LATCHX1_HVT \ram_reg[11][159]  ( .CLK(n107), .D(N176), .Q(\ram[11][159] ) );
  LATCHX1_HVT \ram_reg[11][158]  ( .CLK(n107), .D(N175), .Q(\ram[11][158] ) );
  LATCHX1_HVT \ram_reg[11][157]  ( .CLK(n107), .D(N174), .Q(\ram[11][157] ) );
  LATCHX1_HVT \ram_reg[11][156]  ( .CLK(n107), .D(N173), .Q(\ram[11][156] ) );
  LATCHX1_HVT \ram_reg[11][155]  ( .CLK(n107), .D(N172), .Q(\ram[11][155] ) );
  LATCHX1_HVT \ram_reg[11][154]  ( .CLK(n107), .D(N171), .Q(\ram[11][154] ) );
  LATCHX1_HVT \ram_reg[11][153]  ( .CLK(n107), .D(N170), .Q(\ram[11][153] ) );
  LATCHX1_HVT \ram_reg[11][152]  ( .CLK(n107), .D(N169), .Q(\ram[11][152] ) );
  LATCHX1_HVT \ram_reg[11][151]  ( .CLK(n106), .D(N168), .Q(\ram[11][151] ) );
  LATCHX1_HVT \ram_reg[11][150]  ( .CLK(n106), .D(N167), .Q(\ram[11][150] ) );
  LATCHX1_HVT \ram_reg[11][149]  ( .CLK(n106), .D(N166), .Q(\ram[11][149] ) );
  LATCHX1_HVT \ram_reg[11][148]  ( .CLK(n106), .D(N165), .Q(\ram[11][148] ) );
  LATCHX1_HVT \ram_reg[11][147]  ( .CLK(n106), .D(N164), .Q(\ram[11][147] ) );
  LATCHX1_HVT \ram_reg[11][146]  ( .CLK(n106), .D(N163), .Q(\ram[11][146] ) );
  LATCHX1_HVT \ram_reg[11][145]  ( .CLK(n106), .D(N162), .Q(\ram[11][145] ) );
  LATCHX1_HVT \ram_reg[11][144]  ( .CLK(n106), .D(N161), .Q(\ram[11][144] ) );
  LATCHX1_HVT \ram_reg[11][143]  ( .CLK(n106), .D(N160), .Q(\ram[11][143] ) );
  LATCHX1_HVT \ram_reg[11][142]  ( .CLK(n106), .D(N159), .Q(\ram[11][142] ) );
  LATCHX1_HVT \ram_reg[11][141]  ( .CLK(n106), .D(N158), .Q(\ram[11][141] ) );
  LATCHX1_HVT \ram_reg[11][140]  ( .CLK(n105), .D(N157), .Q(\ram[11][140] ) );
  LATCHX1_HVT \ram_reg[11][139]  ( .CLK(n105), .D(N156), .Q(\ram[11][139] ) );
  LATCHX1_HVT \ram_reg[11][138]  ( .CLK(n104), .D(N155), .Q(\ram[11][138] ) );
  LATCHX1_HVT \ram_reg[11][137]  ( .CLK(n113), .D(N154), .Q(\ram[11][137] ) );
  LATCHX1_HVT \ram_reg[11][136]  ( .CLK(n113), .D(N153), .Q(\ram[11][136] ) );
  LATCHX1_HVT \ram_reg[11][135]  ( .CLK(n112), .D(N152), .Q(\ram[11][135] ) );
  LATCHX1_HVT \ram_reg[11][134]  ( .CLK(n111), .D(N151), .Q(\ram[11][134] ) );
  LATCHX1_HVT \ram_reg[11][133]  ( .CLK(n110), .D(N150), .Q(\ram[11][133] ) );
  LATCHX1_HVT \ram_reg[11][132]  ( .CLK(n109), .D(N149), .Q(\ram[11][132] ) );
  LATCHX1_HVT \ram_reg[11][131]  ( .CLK(n108), .D(N148), .Q(\ram[11][131] ) );
  LATCHX1_HVT \ram_reg[11][130]  ( .CLK(n107), .D(N147), .Q(\ram[11][130] ) );
  LATCHX1_HVT \ram_reg[11][129]  ( .CLK(n106), .D(N146), .Q(\ram[11][129] ) );
  LATCHX1_HVT \ram_reg[11][128]  ( .CLK(n103), .D(N145), .Q(\ram[11][128] ) );
  LATCHX1_HVT \ram_reg[11][127]  ( .CLK(n94), .D(N144), .Q(\ram[11][127] ) );
  LATCHX1_HVT \ram_reg[11][126]  ( .CLK(n94), .D(N143), .Q(\ram[11][126] ) );
  LATCHX1_HVT \ram_reg[11][125]  ( .CLK(n94), .D(N142), .Q(\ram[11][125] ) );
  LATCHX1_HVT \ram_reg[11][124]  ( .CLK(n94), .D(N141), .Q(\ram[11][124] ) );
  LATCHX1_HVT \ram_reg[11][123]  ( .CLK(n94), .D(N140), .Q(\ram[11][123] ) );
  LATCHX1_HVT \ram_reg[11][122]  ( .CLK(n94), .D(N139), .Q(\ram[11][122] ) );
  LATCHX1_HVT \ram_reg[11][121]  ( .CLK(n94), .D(N138), .Q(\ram[11][121] ) );
  LATCHX1_HVT \ram_reg[11][120]  ( .CLK(n94), .D(N137), .Q(\ram[11][120] ) );
  LATCHX1_HVT \ram_reg[11][119]  ( .CLK(n103), .D(N136), .Q(\ram[11][119] ) );
  LATCHX1_HVT \ram_reg[11][118]  ( .CLK(n102), .D(N135), .Q(\ram[11][118] ) );
  LATCHX1_HVT \ram_reg[11][117]  ( .CLK(n102), .D(N134), .Q(\ram[11][117] ) );
  LATCHX1_HVT \ram_reg[11][116]  ( .CLK(n101), .D(N133), .Q(\ram[11][116] ) );
  LATCHX1_HVT \ram_reg[11][115]  ( .CLK(n96), .D(N132), .Q(\ram[11][115] ) );
  LATCHX1_HVT \ram_reg[11][114]  ( .CLK(n101), .D(N131), .Q(\ram[11][114] ) );
  LATCHX1_HVT \ram_reg[11][113]  ( .CLK(n101), .D(N130), .Q(\ram[11][113] ) );
  LATCHX1_HVT \ram_reg[11][112]  ( .CLK(n102), .D(N129), .Q(\ram[11][112] ) );
  LATCHX1_HVT \ram_reg[11][111]  ( .CLK(n101), .D(N128), .Q(\ram[11][111] ) );
  LATCHX1_HVT \ram_reg[11][110]  ( .CLK(n100), .D(N127), .Q(\ram[11][110] ) );
  LATCHX1_HVT \ram_reg[11][109]  ( .CLK(n100), .D(N126), .Q(\ram[11][109] ) );
  LATCHX1_HVT \ram_reg[11][108]  ( .CLK(n97), .D(N125), .Q(\ram[11][108] ) );
  LATCHX1_HVT \ram_reg[11][107]  ( .CLK(n94), .D(N124), .Q(\ram[11][107] ) );
  LATCHX1_HVT \ram_reg[11][106]  ( .CLK(n100), .D(N123), .Q(\ram[11][106] ) );
  LATCHX1_HVT \ram_reg[11][105]  ( .CLK(n100), .D(N122), .Q(\ram[11][105] ) );
  LATCHX1_HVT \ram_reg[11][104]  ( .CLK(n100), .D(N121), .Q(\ram[11][104] ) );
  LATCHX1_HVT \ram_reg[11][103]  ( .CLK(n99), .D(N120), .Q(\ram[11][103] ) );
  LATCHX1_HVT \ram_reg[11][102]  ( .CLK(n98), .D(N119), .Q(\ram[11][102] ) );
  LATCHX1_HVT \ram_reg[11][101]  ( .CLK(n98), .D(N118), .Q(\ram[11][101] ) );
  LATCHX1_HVT \ram_reg[11][100]  ( .CLK(n99), .D(N117), .Q(\ram[11][100] ) );
  LATCHX1_HVT \ram_reg[11][99]  ( .CLK(n97), .D(N116), .Q(\ram[11][99] ) );
  LATCHX1_HVT \ram_reg[11][98]  ( .CLK(n98), .D(N114), .Q(\ram[11][98] ) );
  LATCHX1_HVT \ram_reg[11][97]  ( .CLK(n99), .D(N113), .Q(\ram[11][97] ) );
  LATCHX1_HVT \ram_reg[11][96]  ( .CLK(n103), .D(N112), .Q(\ram[11][96] ) );
  LATCHX1_HVT \ram_reg[11][95]  ( .CLK(n95), .D(N111), .Q(\ram[11][95] ) );
  LATCHX1_HVT \ram_reg[11][94]  ( .CLK(n95), .D(N110), .Q(\ram[11][94] ) );
  LATCHX1_HVT \ram_reg[11][93]  ( .CLK(n95), .D(N109), .Q(\ram[11][93] ) );
  LATCHX1_HVT \ram_reg[11][92]  ( .CLK(n95), .D(N108), .Q(\ram[11][92] ) );
  LATCHX1_HVT \ram_reg[11][91]  ( .CLK(n94), .D(N107), .Q(\ram[11][91] ) );
  LATCHX1_HVT \ram_reg[11][90]  ( .CLK(n95), .D(N106), .Q(\ram[11][90] ) );
  LATCHX1_HVT \ram_reg[11][89]  ( .CLK(n94), .D(N105), .Q(\ram[11][89] ) );
  LATCHX1_HVT \ram_reg[11][88]  ( .CLK(n95), .D(N104), .Q(\ram[11][88] ) );
  LATCHX1_HVT \ram_reg[11][87]  ( .CLK(n103), .D(N103), .Q(\ram[11][87] ) );
  LATCHX1_HVT \ram_reg[11][86]  ( .CLK(n103), .D(N102), .Q(\ram[11][86] ) );
  LATCHX1_HVT \ram_reg[11][85]  ( .CLK(n101), .D(N101), .Q(\ram[11][85] ) );
  LATCHX1_HVT \ram_reg[11][84]  ( .CLK(n102), .D(N100), .Q(\ram[11][84] ) );
  LATCHX1_HVT \ram_reg[11][83]  ( .CLK(n96), .D(N99), .Q(\ram[11][83] ) );
  LATCHX1_HVT \ram_reg[11][82]  ( .CLK(n102), .D(N98), .Q(\ram[11][82] ) );
  LATCHX1_HVT \ram_reg[11][81]  ( .CLK(n101), .D(N97), .Q(\ram[11][81] ) );
  LATCHX1_HVT \ram_reg[11][80]  ( .CLK(n102), .D(N96), .Q(\ram[11][80] ) );
  LATCHX1_HVT \ram_reg[11][79]  ( .CLK(n96), .D(N95), .Q(\ram[11][79] ) );
  LATCHX1_HVT \ram_reg[11][78]  ( .CLK(n95), .D(N94), .Q(\ram[11][78] ) );
  LATCHX1_HVT \ram_reg[11][77]  ( .CLK(n96), .D(N93), .Q(\ram[11][77] ) );
  LATCHX1_HVT \ram_reg[11][76]  ( .CLK(n95), .D(N92), .Q(\ram[11][76] ) );
  LATCHX1_HVT \ram_reg[11][75]  ( .CLK(n95), .D(N91), .Q(\ram[11][75] ) );
  LATCHX1_HVT \ram_reg[11][74]  ( .CLK(n93), .D(N90), .Q(\ram[11][74] ) );
  LATCHX1_HVT \ram_reg[11][73]  ( .CLK(n96), .D(N89), .Q(\ram[11][73] ) );
  LATCHX1_HVT \ram_reg[11][72]  ( .CLK(n96), .D(N88), .Q(\ram[11][72] ) );
  LATCHX1_HVT \ram_reg[11][71]  ( .CLK(n99), .D(N87), .Q(\ram[11][71] ) );
  LATCHX1_HVT \ram_reg[11][70]  ( .CLK(n99), .D(N86), .Q(\ram[11][70] ) );
  LATCHX1_HVT \ram_reg[11][69]  ( .CLK(n98), .D(N85), .Q(\ram[11][69] ) );
  LATCHX1_HVT \ram_reg[11][68]  ( .CLK(n99), .D(N84), .Q(\ram[11][68] ) );
  LATCHX1_HVT \ram_reg[11][67]  ( .CLK(n98), .D(N83), .Q(\ram[11][67] ) );
  LATCHX1_HVT \ram_reg[11][66]  ( .CLK(n97), .D(N82), .Q(\ram[11][66] ) );
  LATCHX1_HVT \ram_reg[11][65]  ( .CLK(n98), .D(N81), .Q(\ram[11][65] ) );
  LATCHX1_HVT \ram_reg[11][64]  ( .CLK(n103), .D(N80), .Q(\ram[11][64] ) );
  LATCHX1_HVT \ram_reg[11][63]  ( .CLK(n97), .D(N79), .Q(\ram[11][63] ) );
  LATCHX1_HVT \ram_reg[11][62]  ( .CLK(n97), .D(N78), .Q(\ram[11][62] ) );
  LATCHX1_HVT \ram_reg[11][61]  ( .CLK(n97), .D(N77), .Q(\ram[11][61] ) );
  LATCHX1_HVT \ram_reg[11][60]  ( .CLK(n97), .D(N76), .Q(\ram[11][60] ) );
  LATCHX1_HVT \ram_reg[11][59]  ( .CLK(n97), .D(N75), .Q(\ram[11][59] ) );
  LATCHX1_HVT \ram_reg[11][58]  ( .CLK(n97), .D(N74), .Q(\ram[11][58] ) );
  LATCHX1_HVT \ram_reg[11][57]  ( .CLK(n97), .D(N73), .Q(\ram[11][57] ) );
  LATCHX1_HVT \ram_reg[11][56]  ( .CLK(n97), .D(N72), .Q(\ram[11][56] ) );
  LATCHX1_HVT \ram_reg[11][55]  ( .CLK(n103), .D(N71), .Q(\ram[11][55] ) );
  LATCHX1_HVT \ram_reg[11][54]  ( .CLK(n101), .D(N70), .Q(\ram[11][54] ) );
  LATCHX1_HVT \ram_reg[11][53]  ( .CLK(n101), .D(N69), .Q(\ram[11][53] ) );
  LATCHX1_HVT \ram_reg[11][52]  ( .CLK(n102), .D(N68), .Q(\ram[11][52] ) );
  LATCHX1_HVT \ram_reg[11][51]  ( .CLK(n96), .D(N67), .Q(\ram[11][51] ) );
  LATCHX1_HVT \ram_reg[11][50]  ( .CLK(n93), .D(N66), .Q(\ram[11][50] ) );
  LATCHX1_HVT \ram_reg[11][49]  ( .CLK(n102), .D(N65), .Q(\ram[11][49] ) );
  LATCHX1_HVT \ram_reg[11][48]  ( .CLK(n102), .D(N64), .Q(\ram[11][48] ) );
  LATCHX1_HVT \ram_reg[11][47]  ( .CLK(n100), .D(N63), .Q(\ram[11][47] ) );
  LATCHX1_HVT \ram_reg[11][46]  ( .CLK(n100), .D(N62), .Q(\ram[11][46] ) );
  LATCHX1_HVT \ram_reg[11][45]  ( .CLK(n100), .D(N61), .Q(\ram[11][45] ) );
  LATCHX1_HVT \ram_reg[11][44]  ( .CLK(n100), .D(N60), .Q(\ram[11][44] ) );
  LATCHX1_HVT \ram_reg[11][43]  ( .CLK(n97), .D(N59), .Q(\ram[11][43] ) );
  LATCHX1_HVT \ram_reg[11][42]  ( .CLK(n101), .D(N58), .Q(\ram[11][42] ) );
  LATCHX1_HVT \ram_reg[11][41]  ( .CLK(n94), .D(N57), .Q(\ram[11][41] ) );
  LATCHX1_HVT \ram_reg[11][40]  ( .CLK(n100), .D(N56), .Q(\ram[11][40] ) );
  LATCHX1_HVT \ram_reg[11][39]  ( .CLK(n99), .D(N55), .Q(\ram[11][39] ) );
  LATCHX1_HVT \ram_reg[11][38]  ( .CLK(n99), .D(N54), .Q(\ram[11][38] ) );
  LATCHX1_HVT \ram_reg[11][37]  ( .CLK(n98), .D(N53), .Q(\ram[11][37] ) );
  LATCHX1_HVT \ram_reg[11][36]  ( .CLK(n98), .D(N52), .Q(\ram[11][36] ) );
  LATCHX1_HVT \ram_reg[11][35]  ( .CLK(n98), .D(N51), .Q(\ram[11][35] ) );
  LATCHX1_HVT \ram_reg[11][34]  ( .CLK(n100), .D(N50), .Q(\ram[11][34] ) );
  LATCHX1_HVT \ram_reg[11][33]  ( .CLK(n99), .D(N49), .Q(\ram[11][33] ) );
  LATCHX1_HVT \ram_reg[11][32]  ( .CLK(n103), .D(N48), .Q(\ram[11][32] ) );
  LATCHX1_HVT \ram_reg[11][31]  ( .CLK(n93), .D(N47), .Q(\ram[11][31] ) );
  LATCHX1_HVT \ram_reg[11][30]  ( .CLK(n93), .D(N46), .Q(\ram[11][30] ) );
  LATCHX1_HVT \ram_reg[11][29]  ( .CLK(n93), .D(N45), .Q(\ram[11][29] ) );
  LATCHX1_HVT \ram_reg[11][28]  ( .CLK(n93), .D(N44), .Q(\ram[11][28] ) );
  LATCHX1_HVT \ram_reg[11][27]  ( .CLK(n93), .D(N43), .Q(\ram[11][27] ) );
  LATCHX1_HVT \ram_reg[11][26]  ( .CLK(n93), .D(N42), .Q(\ram[11][26] ) );
  LATCHX1_HVT \ram_reg[11][25]  ( .CLK(n93), .D(N41), .Q(\ram[11][25] ) );
  LATCHX1_HVT \ram_reg[11][24]  ( .CLK(n93), .D(N40), .Q(\ram[11][24] ) );
  LATCHX1_HVT \ram_reg[11][23]  ( .CLK(n103), .D(N39), .Q(\ram[11][23] ) );
  LATCHX1_HVT \ram_reg[11][22]  ( .CLK(n102), .D(N38), .Q(\ram[11][22] ) );
  LATCHX1_HVT \ram_reg[11][21]  ( .CLK(n101), .D(N37), .Q(\ram[11][21] ) );
  LATCHX1_HVT \ram_reg[11][20]  ( .CLK(n101), .D(N36), .Q(\ram[11][20] ) );
  LATCHX1_HVT \ram_reg[11][19]  ( .CLK(n93), .D(N35), .Q(\ram[11][19] ) );
  LATCHX1_HVT \ram_reg[11][18]  ( .CLK(n101), .D(N34), .Q(\ram[11][18] ) );
  LATCHX1_HVT \ram_reg[11][17]  ( .CLK(n102), .D(N33), .Q(\ram[11][17] ) );
  LATCHX1_HVT \ram_reg[11][16]  ( .CLK(n102), .D(N32), .Q(\ram[11][16] ) );
  LATCHX1_HVT \ram_reg[11][15]  ( .CLK(n96), .D(N31), .Q(\ram[11][15] ) );
  LATCHX1_HVT \ram_reg[11][14]  ( .CLK(n96), .D(N30), .Q(\ram[11][14] ) );
  LATCHX1_HVT \ram_reg[11][13]  ( .CLK(n95), .D(N29), .Q(\ram[11][13] ) );
  LATCHX1_HVT \ram_reg[11][12]  ( .CLK(n96), .D(N28), .Q(\ram[11][12] ) );
  LATCHX1_HVT \ram_reg[11][11]  ( .CLK(n96), .D(N27), .Q(\ram[11][11] ) );
  LATCHX1_HVT \ram_reg[11][10]  ( .CLK(n95), .D(N26), .Q(\ram[11][10] ) );
  LATCHX1_HVT \ram_reg[11][9]  ( .CLK(n95), .D(N25), .Q(\ram[11][9] ) );
  LATCHX1_HVT \ram_reg[11][8]  ( .CLK(n96), .D(N24), .Q(\ram[11][8] ) );
  LATCHX1_HVT \ram_reg[11][7]  ( .CLK(n100), .D(N23), .Q(\ram[11][7] ) );
  LATCHX1_HVT \ram_reg[11][6]  ( .CLK(n99), .D(N22), .Q(\ram[11][6] ) );
  LATCHX1_HVT \ram_reg[11][5]  ( .CLK(n98), .D(N21), .Q(\ram[11][5] ) );
  LATCHX1_HVT \ram_reg[11][4]  ( .CLK(n99), .D(N20), .Q(\ram[11][4] ) );
  LATCHX1_HVT \ram_reg[11][3]  ( .CLK(n98), .D(N19), .Q(\ram[11][3] ) );
  LATCHX1_HVT \ram_reg[11][2]  ( .CLK(n98), .D(N18), .Q(\ram[11][2] ) );
  LATCHX1_HVT \ram_reg[11][1]  ( .CLK(n99), .D(N17), .Q(\ram[11][1] ) );
  LATCHX1_HVT \ram_reg[11][0]  ( .CLK(n103), .D(N16), .Q(\ram[11][0] ) );
  LATCHX1_HVT \ram_reg[10][255]  ( .CLK(N303), .D(N273), .Q(\ram[10][255] ) );
  LATCHX1_HVT \ram_reg[10][254]  ( .CLK(N303), .D(N272), .Q(\ram[10][254] ) );
  LATCHX1_HVT \ram_reg[10][253]  ( .CLK(N303), .D(N271), .Q(\ram[10][253] ) );
  LATCHX1_HVT \ram_reg[10][252]  ( .CLK(N303), .D(N270), .Q(\ram[10][252] ) );
  LATCHX1_HVT \ram_reg[10][251]  ( .CLK(n136), .D(N269), .Q(\ram[10][251] ) );
  LATCHX1_HVT \ram_reg[10][250]  ( .CLK(n128), .D(N268), .Q(\ram[10][250] ) );
  LATCHX1_HVT \ram_reg[10][249]  ( .CLK(n128), .D(N267), .Q(\ram[10][249] ) );
  LATCHX1_HVT \ram_reg[10][248]  ( .CLK(n128), .D(N266), .Q(\ram[10][248] ) );
  LATCHX1_HVT \ram_reg[10][247]  ( .CLK(n128), .D(N265), .Q(\ram[10][247] ) );
  LATCHX1_HVT \ram_reg[10][246]  ( .CLK(n128), .D(N264), .Q(\ram[10][246] ) );
  LATCHX1_HVT \ram_reg[10][245]  ( .CLK(n128), .D(N263), .Q(\ram[10][245] ) );
  LATCHX1_HVT \ram_reg[10][244]  ( .CLK(n128), .D(N262), .Q(\ram[10][244] ) );
  LATCHX1_HVT \ram_reg[10][243]  ( .CLK(n128), .D(N261), .Q(\ram[10][243] ) );
  LATCHX1_HVT \ram_reg[10][242]  ( .CLK(n128), .D(N260), .Q(\ram[10][242] ) );
  LATCHX1_HVT \ram_reg[10][241]  ( .CLK(n127), .D(N259), .Q(\ram[10][241] ) );
  LATCHX1_HVT \ram_reg[10][240]  ( .CLK(n127), .D(N258), .Q(\ram[10][240] ) );
  LATCHX1_HVT \ram_reg[10][239]  ( .CLK(n127), .D(N257), .Q(\ram[10][239] ) );
  LATCHX1_HVT \ram_reg[10][238]  ( .CLK(n127), .D(N256), .Q(\ram[10][238] ) );
  LATCHX1_HVT \ram_reg[10][237]  ( .CLK(n127), .D(N255), .Q(\ram[10][237] ) );
  LATCHX1_HVT \ram_reg[10][236]  ( .CLK(n127), .D(N254), .Q(\ram[10][236] ) );
  LATCHX1_HVT \ram_reg[10][235]  ( .CLK(n127), .D(N253), .Q(\ram[10][235] ) );
  LATCHX1_HVT \ram_reg[10][234]  ( .CLK(n127), .D(N252), .Q(\ram[10][234] ) );
  LATCHX1_HVT \ram_reg[10][233]  ( .CLK(n127), .D(N251), .Q(\ram[10][233] ) );
  LATCHX1_HVT \ram_reg[10][232]  ( .CLK(n127), .D(N250), .Q(\ram[10][232] ) );
  LATCHX1_HVT \ram_reg[10][231]  ( .CLK(n127), .D(N249), .Q(\ram[10][231] ) );
  LATCHX1_HVT \ram_reg[10][230]  ( .CLK(n126), .D(N248), .Q(\ram[10][230] ) );
  LATCHX1_HVT \ram_reg[10][229]  ( .CLK(n126), .D(N247), .Q(\ram[10][229] ) );
  LATCHX1_HVT \ram_reg[10][228]  ( .CLK(n126), .D(N246), .Q(\ram[10][228] ) );
  LATCHX1_HVT \ram_reg[10][227]  ( .CLK(n136), .D(N245), .Q(\ram[10][227] ) );
  LATCHX1_HVT \ram_reg[10][226]  ( .CLK(n136), .D(N244), .Q(\ram[10][226] ) );
  LATCHX1_HVT \ram_reg[10][225]  ( .CLK(n136), .D(N243), .Q(\ram[10][225] ) );
  LATCHX1_HVT \ram_reg[10][224]  ( .CLK(n136), .D(N242), .Q(\ram[10][224] ) );
  LATCHX1_HVT \ram_reg[10][223]  ( .CLK(n136), .D(N241), .Q(\ram[10][223] ) );
  LATCHX1_HVT \ram_reg[10][222]  ( .CLK(n136), .D(N240), .Q(\ram[10][222] ) );
  LATCHX1_HVT \ram_reg[10][221]  ( .CLK(n136), .D(N239), .Q(\ram[10][221] ) );
  LATCHX1_HVT \ram_reg[10][220]  ( .CLK(n136), .D(N238), .Q(\ram[10][220] ) );
  LATCHX1_HVT \ram_reg[10][219]  ( .CLK(n136), .D(N237), .Q(\ram[10][219] ) );
  LATCHX1_HVT \ram_reg[10][218]  ( .CLK(n136), .D(N236), .Q(\ram[10][218] ) );
  LATCHX1_HVT \ram_reg[10][217]  ( .CLK(n135), .D(N235), .Q(\ram[10][217] ) );
  LATCHX1_HVT \ram_reg[10][216]  ( .CLK(n135), .D(N234), .Q(\ram[10][216] ) );
  LATCHX1_HVT \ram_reg[10][215]  ( .CLK(n135), .D(N233), .Q(\ram[10][215] ) );
  LATCHX1_HVT \ram_reg[10][214]  ( .CLK(n135), .D(N232), .Q(\ram[10][214] ) );
  LATCHX1_HVT \ram_reg[10][213]  ( .CLK(n135), .D(N231), .Q(\ram[10][213] ) );
  LATCHX1_HVT \ram_reg[10][212]  ( .CLK(n135), .D(N230), .Q(\ram[10][212] ) );
  LATCHX1_HVT \ram_reg[10][211]  ( .CLK(n135), .D(N229), .Q(\ram[10][211] ) );
  LATCHX1_HVT \ram_reg[10][210]  ( .CLK(n135), .D(N228), .Q(\ram[10][210] ) );
  LATCHX1_HVT \ram_reg[10][209]  ( .CLK(n135), .D(N227), .Q(\ram[10][209] ) );
  LATCHX1_HVT \ram_reg[10][208]  ( .CLK(n135), .D(N226), .Q(\ram[10][208] ) );
  LATCHX1_HVT \ram_reg[10][207]  ( .CLK(n134), .D(N225), .Q(\ram[10][207] ) );
  LATCHX1_HVT \ram_reg[10][206]  ( .CLK(n134), .D(N224), .Q(\ram[10][206] ) );
  LATCHX1_HVT \ram_reg[10][205]  ( .CLK(n134), .D(N223), .Q(\ram[10][205] ) );
  LATCHX1_HVT \ram_reg[10][204]  ( .CLK(n134), .D(N222), .Q(\ram[10][204] ) );
  LATCHX1_HVT \ram_reg[10][203]  ( .CLK(n134), .D(N221), .Q(\ram[10][203] ) );
  LATCHX1_HVT \ram_reg[10][202]  ( .CLK(n134), .D(N220), .Q(\ram[10][202] ) );
  LATCHX1_HVT \ram_reg[10][201]  ( .CLK(n134), .D(N219), .Q(\ram[10][201] ) );
  LATCHX1_HVT \ram_reg[10][200]  ( .CLK(n134), .D(N218), .Q(\ram[10][200] ) );
  LATCHX1_HVT \ram_reg[10][199]  ( .CLK(n134), .D(N217), .Q(\ram[10][199] ) );
  LATCHX1_HVT \ram_reg[10][198]  ( .CLK(n134), .D(N216), .Q(\ram[10][198] ) );
  LATCHX1_HVT \ram_reg[10][197]  ( .CLK(n134), .D(N214), .Q(\ram[10][197] ) );
  LATCHX1_HVT \ram_reg[10][196]  ( .CLK(n133), .D(N213), .Q(\ram[10][196] ) );
  LATCHX1_HVT \ram_reg[10][195]  ( .CLK(n133), .D(N212), .Q(\ram[10][195] ) );
  LATCHX1_HVT \ram_reg[10][194]  ( .CLK(n133), .D(N211), .Q(\ram[10][194] ) );
  LATCHX1_HVT \ram_reg[10][193]  ( .CLK(n133), .D(N210), .Q(\ram[10][193] ) );
  LATCHX1_HVT \ram_reg[10][192]  ( .CLK(n133), .D(N209), .Q(\ram[10][192] ) );
  LATCHX1_HVT \ram_reg[10][191]  ( .CLK(n133), .D(N208), .Q(\ram[10][191] ) );
  LATCHX1_HVT \ram_reg[10][190]  ( .CLK(n133), .D(N207), .Q(\ram[10][190] ) );
  LATCHX1_HVT \ram_reg[10][189]  ( .CLK(n133), .D(N206), .Q(\ram[10][189] ) );
  LATCHX1_HVT \ram_reg[10][188]  ( .CLK(n133), .D(N205), .Q(\ram[10][188] ) );
  LATCHX1_HVT \ram_reg[10][187]  ( .CLK(n133), .D(N204), .Q(\ram[10][187] ) );
  LATCHX1_HVT \ram_reg[10][186]  ( .CLK(n133), .D(N203), .Q(\ram[10][186] ) );
  LATCHX1_HVT \ram_reg[10][185]  ( .CLK(n132), .D(N202), .Q(\ram[10][185] ) );
  LATCHX1_HVT \ram_reg[10][184]  ( .CLK(n132), .D(N201), .Q(\ram[10][184] ) );
  LATCHX1_HVT \ram_reg[10][183]  ( .CLK(n132), .D(N200), .Q(\ram[10][183] ) );
  LATCHX1_HVT \ram_reg[10][182]  ( .CLK(n132), .D(N199), .Q(\ram[10][182] ) );
  LATCHX1_HVT \ram_reg[10][181]  ( .CLK(n132), .D(N198), .Q(\ram[10][181] ) );
  LATCHX1_HVT \ram_reg[10][180]  ( .CLK(n132), .D(N197), .Q(\ram[10][180] ) );
  LATCHX1_HVT \ram_reg[10][179]  ( .CLK(n132), .D(N196), .Q(\ram[10][179] ) );
  LATCHX1_HVT \ram_reg[10][178]  ( .CLK(n132), .D(N195), .Q(\ram[10][178] ) );
  LATCHX1_HVT \ram_reg[10][177]  ( .CLK(n132), .D(N194), .Q(\ram[10][177] ) );
  LATCHX1_HVT \ram_reg[10][176]  ( .CLK(n132), .D(N193), .Q(\ram[10][176] ) );
  LATCHX1_HVT \ram_reg[10][175]  ( .CLK(n132), .D(N192), .Q(\ram[10][175] ) );
  LATCHX1_HVT \ram_reg[10][174]  ( .CLK(n131), .D(N191), .Q(\ram[10][174] ) );
  LATCHX1_HVT \ram_reg[10][173]  ( .CLK(n131), .D(N190), .Q(\ram[10][173] ) );
  LATCHX1_HVT \ram_reg[10][172]  ( .CLK(n131), .D(N189), .Q(\ram[10][172] ) );
  LATCHX1_HVT \ram_reg[10][171]  ( .CLK(n131), .D(N188), .Q(\ram[10][171] ) );
  LATCHX1_HVT \ram_reg[10][170]  ( .CLK(n131), .D(N187), .Q(\ram[10][170] ) );
  LATCHX1_HVT \ram_reg[10][169]  ( .CLK(n131), .D(N186), .Q(\ram[10][169] ) );
  LATCHX1_HVT \ram_reg[10][168]  ( .CLK(n131), .D(N185), .Q(\ram[10][168] ) );
  LATCHX1_HVT \ram_reg[10][167]  ( .CLK(n131), .D(N184), .Q(\ram[10][167] ) );
  LATCHX1_HVT \ram_reg[10][166]  ( .CLK(n131), .D(N183), .Q(\ram[10][166] ) );
  LATCHX1_HVT \ram_reg[10][165]  ( .CLK(n131), .D(N182), .Q(\ram[10][165] ) );
  LATCHX1_HVT \ram_reg[10][164]  ( .CLK(n131), .D(N181), .Q(\ram[10][164] ) );
  LATCHX1_HVT \ram_reg[10][163]  ( .CLK(n130), .D(N180), .Q(\ram[10][163] ) );
  LATCHX1_HVT \ram_reg[10][162]  ( .CLK(n130), .D(N179), .Q(\ram[10][162] ) );
  LATCHX1_HVT \ram_reg[10][161]  ( .CLK(n130), .D(N178), .Q(\ram[10][161] ) );
  LATCHX1_HVT \ram_reg[10][160]  ( .CLK(n130), .D(N177), .Q(\ram[10][160] ) );
  LATCHX1_HVT \ram_reg[10][159]  ( .CLK(n130), .D(N176), .Q(\ram[10][159] ) );
  LATCHX1_HVT \ram_reg[10][158]  ( .CLK(n130), .D(N175), .Q(\ram[10][158] ) );
  LATCHX1_HVT \ram_reg[10][157]  ( .CLK(n130), .D(N174), .Q(\ram[10][157] ) );
  LATCHX1_HVT \ram_reg[10][156]  ( .CLK(n130), .D(N173), .Q(\ram[10][156] ) );
  LATCHX1_HVT \ram_reg[10][155]  ( .CLK(n130), .D(N172), .Q(\ram[10][155] ) );
  LATCHX1_HVT \ram_reg[10][154]  ( .CLK(n130), .D(N171), .Q(\ram[10][154] ) );
  LATCHX1_HVT \ram_reg[10][153]  ( .CLK(n130), .D(N170), .Q(\ram[10][153] ) );
  LATCHX1_HVT \ram_reg[10][152]  ( .CLK(n129), .D(N169), .Q(\ram[10][152] ) );
  LATCHX1_HVT \ram_reg[10][151]  ( .CLK(n129), .D(N168), .Q(\ram[10][151] ) );
  LATCHX1_HVT \ram_reg[10][150]  ( .CLK(n129), .D(N167), .Q(\ram[10][150] ) );
  LATCHX1_HVT \ram_reg[10][149]  ( .CLK(n129), .D(N166), .Q(\ram[10][149] ) );
  LATCHX1_HVT \ram_reg[10][148]  ( .CLK(n129), .D(N165), .Q(\ram[10][148] ) );
  LATCHX1_HVT \ram_reg[10][147]  ( .CLK(n129), .D(N164), .Q(\ram[10][147] ) );
  LATCHX1_HVT \ram_reg[10][146]  ( .CLK(n129), .D(N163), .Q(\ram[10][146] ) );
  LATCHX1_HVT \ram_reg[10][145]  ( .CLK(n129), .D(N162), .Q(\ram[10][145] ) );
  LATCHX1_HVT \ram_reg[10][144]  ( .CLK(n129), .D(N161), .Q(\ram[10][144] ) );
  LATCHX1_HVT \ram_reg[10][143]  ( .CLK(n129), .D(N160), .Q(\ram[10][143] ) );
  LATCHX1_HVT \ram_reg[10][142]  ( .CLK(n129), .D(N159), .Q(\ram[10][142] ) );
  LATCHX1_HVT \ram_reg[10][141]  ( .CLK(n128), .D(N158), .Q(\ram[10][141] ) );
  LATCHX1_HVT \ram_reg[10][140]  ( .CLK(n128), .D(N157), .Q(\ram[10][140] ) );
  LATCHX1_HVT \ram_reg[10][139]  ( .CLK(n128), .D(N156), .Q(\ram[10][139] ) );
  LATCHX1_HVT \ram_reg[10][138]  ( .CLK(n127), .D(N155), .Q(\ram[10][138] ) );
  LATCHX1_HVT \ram_reg[10][137]  ( .CLK(n136), .D(N154), .Q(\ram[10][137] ) );
  LATCHX1_HVT \ram_reg[10][136]  ( .CLK(n135), .D(N153), .Q(\ram[10][136] ) );
  LATCHX1_HVT \ram_reg[10][135]  ( .CLK(n135), .D(N152), .Q(\ram[10][135] ) );
  LATCHX1_HVT \ram_reg[10][134]  ( .CLK(n134), .D(N151), .Q(\ram[10][134] ) );
  LATCHX1_HVT \ram_reg[10][133]  ( .CLK(n133), .D(N150), .Q(\ram[10][133] ) );
  LATCHX1_HVT \ram_reg[10][132]  ( .CLK(n132), .D(N149), .Q(\ram[10][132] ) );
  LATCHX1_HVT \ram_reg[10][131]  ( .CLK(n131), .D(N148), .Q(\ram[10][131] ) );
  LATCHX1_HVT \ram_reg[10][130]  ( .CLK(n130), .D(N147), .Q(\ram[10][130] ) );
  LATCHX1_HVT \ram_reg[10][129]  ( .CLK(n129), .D(N146), .Q(\ram[10][129] ) );
  LATCHX1_HVT \ram_reg[10][128]  ( .CLK(n126), .D(N145), .Q(\ram[10][128] ) );
  LATCHX1_HVT \ram_reg[10][127]  ( .CLK(n117), .D(N144), .Q(\ram[10][127] ) );
  LATCHX1_HVT \ram_reg[10][126]  ( .CLK(n117), .D(N143), .Q(\ram[10][126] ) );
  LATCHX1_HVT \ram_reg[10][125]  ( .CLK(n117), .D(N142), .Q(\ram[10][125] ) );
  LATCHX1_HVT \ram_reg[10][124]  ( .CLK(n117), .D(N141), .Q(\ram[10][124] ) );
  LATCHX1_HVT \ram_reg[10][123]  ( .CLK(n117), .D(N140), .Q(\ram[10][123] ) );
  LATCHX1_HVT \ram_reg[10][122]  ( .CLK(n116), .D(N139), .Q(\ram[10][122] ) );
  LATCHX1_HVT \ram_reg[10][121]  ( .CLK(n117), .D(N138), .Q(\ram[10][121] ) );
  LATCHX1_HVT \ram_reg[10][120]  ( .CLK(n117), .D(N137), .Q(\ram[10][120] ) );
  LATCHX1_HVT \ram_reg[10][119]  ( .CLK(n126), .D(N136), .Q(\ram[10][119] ) );
  LATCHX1_HVT \ram_reg[10][118]  ( .CLK(n125), .D(N135), .Q(\ram[10][118] ) );
  LATCHX1_HVT \ram_reg[10][117]  ( .CLK(n125), .D(N134), .Q(\ram[10][117] ) );
  LATCHX1_HVT \ram_reg[10][116]  ( .CLK(n124), .D(N133), .Q(\ram[10][116] ) );
  LATCHX1_HVT \ram_reg[10][115]  ( .CLK(n119), .D(N132), .Q(\ram[10][115] ) );
  LATCHX1_HVT \ram_reg[10][114]  ( .CLK(n124), .D(N131), .Q(\ram[10][114] ) );
  LATCHX1_HVT \ram_reg[10][113]  ( .CLK(n124), .D(N130), .Q(\ram[10][113] ) );
  LATCHX1_HVT \ram_reg[10][112]  ( .CLK(n125), .D(N129), .Q(\ram[10][112] ) );
  LATCHX1_HVT \ram_reg[10][111]  ( .CLK(n123), .D(N128), .Q(\ram[10][111] ) );
  LATCHX1_HVT \ram_reg[10][110]  ( .CLK(n123), .D(N127), .Q(\ram[10][110] ) );
  LATCHX1_HVT \ram_reg[10][109]  ( .CLK(n123), .D(N126), .Q(\ram[10][109] ) );
  LATCHX1_HVT \ram_reg[10][108]  ( .CLK(n120), .D(N125), .Q(\ram[10][108] ) );
  LATCHX1_HVT \ram_reg[10][107]  ( .CLK(n117), .D(N124), .Q(\ram[10][107] ) );
  LATCHX1_HVT \ram_reg[10][106]  ( .CLK(n123), .D(N123), .Q(\ram[10][106] ) );
  LATCHX1_HVT \ram_reg[10][105]  ( .CLK(n123), .D(N122), .Q(\ram[10][105] ) );
  LATCHX1_HVT \ram_reg[10][104]  ( .CLK(n123), .D(N121), .Q(\ram[10][104] ) );
  LATCHX1_HVT \ram_reg[10][103]  ( .CLK(n122), .D(N120), .Q(\ram[10][103] ) );
  LATCHX1_HVT \ram_reg[10][102]  ( .CLK(n121), .D(N119), .Q(\ram[10][102] ) );
  LATCHX1_HVT \ram_reg[10][101]  ( .CLK(n121), .D(N118), .Q(\ram[10][101] ) );
  LATCHX1_HVT \ram_reg[10][100]  ( .CLK(n122), .D(N117), .Q(\ram[10][100] ) );
  LATCHX1_HVT \ram_reg[10][99]  ( .CLK(n120), .D(N116), .Q(\ram[10][99] ) );
  LATCHX1_HVT \ram_reg[10][98]  ( .CLK(n121), .D(N114), .Q(\ram[10][98] ) );
  LATCHX1_HVT \ram_reg[10][97]  ( .CLK(n122), .D(N113), .Q(\ram[10][97] ) );
  LATCHX1_HVT \ram_reg[10][96]  ( .CLK(n126), .D(N112), .Q(\ram[10][96] ) );
  LATCHX1_HVT \ram_reg[10][95]  ( .CLK(n118), .D(N111), .Q(\ram[10][95] ) );
  LATCHX1_HVT \ram_reg[10][94]  ( .CLK(n118), .D(N110), .Q(\ram[10][94] ) );
  LATCHX1_HVT \ram_reg[10][93]  ( .CLK(n118), .D(N109), .Q(\ram[10][93] ) );
  LATCHX1_HVT \ram_reg[10][92]  ( .CLK(n117), .D(N108), .Q(\ram[10][92] ) );
  LATCHX1_HVT \ram_reg[10][91]  ( .CLK(n117), .D(N107), .Q(\ram[10][91] ) );
  LATCHX1_HVT \ram_reg[10][90]  ( .CLK(n118), .D(N106), .Q(\ram[10][90] ) );
  LATCHX1_HVT \ram_reg[10][89]  ( .CLK(n117), .D(N105), .Q(\ram[10][89] ) );
  LATCHX1_HVT \ram_reg[10][88]  ( .CLK(n118), .D(N104), .Q(\ram[10][88] ) );
  LATCHX1_HVT \ram_reg[10][87]  ( .CLK(n126), .D(N103), .Q(\ram[10][87] ) );
  LATCHX1_HVT \ram_reg[10][86]  ( .CLK(n125), .D(N102), .Q(\ram[10][86] ) );
  LATCHX1_HVT \ram_reg[10][85]  ( .CLK(n124), .D(N101), .Q(\ram[10][85] ) );
  LATCHX1_HVT \ram_reg[10][84]  ( .CLK(n124), .D(N100), .Q(\ram[10][84] ) );
  LATCHX1_HVT \ram_reg[10][83]  ( .CLK(n119), .D(N99), .Q(\ram[10][83] ) );
  LATCHX1_HVT \ram_reg[10][82]  ( .CLK(n125), .D(N98), .Q(\ram[10][82] ) );
  LATCHX1_HVT \ram_reg[10][81]  ( .CLK(n124), .D(N97), .Q(\ram[10][81] ) );
  LATCHX1_HVT \ram_reg[10][80]  ( .CLK(n125), .D(N96), .Q(\ram[10][80] ) );
  LATCHX1_HVT \ram_reg[10][79]  ( .CLK(n119), .D(N95), .Q(\ram[10][79] ) );
  LATCHX1_HVT \ram_reg[10][78]  ( .CLK(n118), .D(N94), .Q(\ram[10][78] ) );
  LATCHX1_HVT \ram_reg[10][77]  ( .CLK(n119), .D(N93), .Q(\ram[10][77] ) );
  LATCHX1_HVT \ram_reg[10][76]  ( .CLK(n118), .D(N92), .Q(\ram[10][76] ) );
  LATCHX1_HVT \ram_reg[10][75]  ( .CLK(n118), .D(N91), .Q(\ram[10][75] ) );
  LATCHX1_HVT \ram_reg[10][74]  ( .CLK(n116), .D(N90), .Q(\ram[10][74] ) );
  LATCHX1_HVT \ram_reg[10][73]  ( .CLK(n119), .D(N89), .Q(\ram[10][73] ) );
  LATCHX1_HVT \ram_reg[10][72]  ( .CLK(n119), .D(N88), .Q(\ram[10][72] ) );
  LATCHX1_HVT \ram_reg[10][71]  ( .CLK(n122), .D(N87), .Q(\ram[10][71] ) );
  LATCHX1_HVT \ram_reg[10][70]  ( .CLK(n122), .D(N86), .Q(\ram[10][70] ) );
  LATCHX1_HVT \ram_reg[10][69]  ( .CLK(n121), .D(N85), .Q(\ram[10][69] ) );
  LATCHX1_HVT \ram_reg[10][68]  ( .CLK(n122), .D(N84), .Q(\ram[10][68] ) );
  LATCHX1_HVT \ram_reg[10][67]  ( .CLK(n121), .D(N83), .Q(\ram[10][67] ) );
  LATCHX1_HVT \ram_reg[10][66]  ( .CLK(n120), .D(N82), .Q(\ram[10][66] ) );
  LATCHX1_HVT \ram_reg[10][65]  ( .CLK(n121), .D(N81), .Q(\ram[10][65] ) );
  LATCHX1_HVT \ram_reg[10][64]  ( .CLK(n126), .D(N80), .Q(\ram[10][64] ) );
  LATCHX1_HVT \ram_reg[10][63]  ( .CLK(n120), .D(N79), .Q(\ram[10][63] ) );
  LATCHX1_HVT \ram_reg[10][62]  ( .CLK(n120), .D(N78), .Q(\ram[10][62] ) );
  LATCHX1_HVT \ram_reg[10][61]  ( .CLK(n120), .D(N77), .Q(\ram[10][61] ) );
  LATCHX1_HVT \ram_reg[10][60]  ( .CLK(n120), .D(N76), .Q(\ram[10][60] ) );
  LATCHX1_HVT \ram_reg[10][59]  ( .CLK(n120), .D(N75), .Q(\ram[10][59] ) );
  LATCHX1_HVT \ram_reg[10][58]  ( .CLK(n119), .D(N74), .Q(\ram[10][58] ) );
  LATCHX1_HVT \ram_reg[10][57]  ( .CLK(n120), .D(N73), .Q(\ram[10][57] ) );
  LATCHX1_HVT \ram_reg[10][56]  ( .CLK(n120), .D(N72), .Q(\ram[10][56] ) );
  LATCHX1_HVT \ram_reg[10][55]  ( .CLK(n126), .D(N71), .Q(\ram[10][55] ) );
  LATCHX1_HVT \ram_reg[10][54]  ( .CLK(n124), .D(N70), .Q(\ram[10][54] ) );
  LATCHX1_HVT \ram_reg[10][53]  ( .CLK(n124), .D(N69), .Q(\ram[10][53] ) );
  LATCHX1_HVT \ram_reg[10][52]  ( .CLK(n125), .D(N68), .Q(\ram[10][52] ) );
  LATCHX1_HVT \ram_reg[10][51]  ( .CLK(n119), .D(N67), .Q(\ram[10][51] ) );
  LATCHX1_HVT \ram_reg[10][50]  ( .CLK(n116), .D(N66), .Q(\ram[10][50] ) );
  LATCHX1_HVT \ram_reg[10][49]  ( .CLK(n125), .D(N65), .Q(\ram[10][49] ) );
  LATCHX1_HVT \ram_reg[10][48]  ( .CLK(n125), .D(N64), .Q(\ram[10][48] ) );
  LATCHX1_HVT \ram_reg[10][47]  ( .CLK(n123), .D(N63), .Q(\ram[10][47] ) );
  LATCHX1_HVT \ram_reg[10][46]  ( .CLK(n123), .D(N62), .Q(\ram[10][46] ) );
  LATCHX1_HVT \ram_reg[10][45]  ( .CLK(n123), .D(N61), .Q(\ram[10][45] ) );
  LATCHX1_HVT \ram_reg[10][44]  ( .CLK(n123), .D(N60), .Q(\ram[10][44] ) );
  LATCHX1_HVT \ram_reg[10][43]  ( .CLK(n120), .D(N59), .Q(\ram[10][43] ) );
  LATCHX1_HVT \ram_reg[10][42]  ( .CLK(n124), .D(N58), .Q(\ram[10][42] ) );
  LATCHX1_HVT \ram_reg[10][41]  ( .CLK(n117), .D(N57), .Q(\ram[10][41] ) );
  LATCHX1_HVT \ram_reg[10][40]  ( .CLK(n123), .D(N56), .Q(\ram[10][40] ) );
  LATCHX1_HVT \ram_reg[10][39]  ( .CLK(n122), .D(N55), .Q(\ram[10][39] ) );
  LATCHX1_HVT \ram_reg[10][38]  ( .CLK(n122), .D(N54), .Q(\ram[10][38] ) );
  LATCHX1_HVT \ram_reg[10][37]  ( .CLK(n121), .D(N53), .Q(\ram[10][37] ) );
  LATCHX1_HVT \ram_reg[10][36]  ( .CLK(n121), .D(N52), .Q(\ram[10][36] ) );
  LATCHX1_HVT \ram_reg[10][35]  ( .CLK(n121), .D(N51), .Q(\ram[10][35] ) );
  LATCHX1_HVT \ram_reg[10][34]  ( .CLK(n123), .D(N50), .Q(\ram[10][34] ) );
  LATCHX1_HVT \ram_reg[10][33]  ( .CLK(n122), .D(N49), .Q(\ram[10][33] ) );
  LATCHX1_HVT \ram_reg[10][32]  ( .CLK(n126), .D(N48), .Q(\ram[10][32] ) );
  LATCHX1_HVT \ram_reg[10][31]  ( .CLK(n116), .D(N47), .Q(\ram[10][31] ) );
  LATCHX1_HVT \ram_reg[10][30]  ( .CLK(n116), .D(N46), .Q(\ram[10][30] ) );
  LATCHX1_HVT \ram_reg[10][29]  ( .CLK(n116), .D(N45), .Q(\ram[10][29] ) );
  LATCHX1_HVT \ram_reg[10][28]  ( .CLK(n116), .D(N44), .Q(\ram[10][28] ) );
  LATCHX1_HVT \ram_reg[10][27]  ( .CLK(n116), .D(N43), .Q(\ram[10][27] ) );
  LATCHX1_HVT \ram_reg[10][26]  ( .CLK(n116), .D(N42), .Q(\ram[10][26] ) );
  LATCHX1_HVT \ram_reg[10][25]  ( .CLK(n116), .D(N41), .Q(\ram[10][25] ) );
  LATCHX1_HVT \ram_reg[10][24]  ( .CLK(n116), .D(N40), .Q(\ram[10][24] ) );
  LATCHX1_HVT \ram_reg[10][23]  ( .CLK(n126), .D(N39), .Q(\ram[10][23] ) );
  LATCHX1_HVT \ram_reg[10][22]  ( .CLK(n125), .D(N38), .Q(\ram[10][22] ) );
  LATCHX1_HVT \ram_reg[10][21]  ( .CLK(n124), .D(N37), .Q(\ram[10][21] ) );
  LATCHX1_HVT \ram_reg[10][20]  ( .CLK(n124), .D(N36), .Q(\ram[10][20] ) );
  LATCHX1_HVT \ram_reg[10][19]  ( .CLK(n116), .D(N35), .Q(\ram[10][19] ) );
  LATCHX1_HVT \ram_reg[10][18]  ( .CLK(n124), .D(N34), .Q(\ram[10][18] ) );
  LATCHX1_HVT \ram_reg[10][17]  ( .CLK(n125), .D(N33), .Q(\ram[10][17] ) );
  LATCHX1_HVT \ram_reg[10][16]  ( .CLK(n125), .D(N32), .Q(\ram[10][16] ) );
  LATCHX1_HVT \ram_reg[10][15]  ( .CLK(n119), .D(N31), .Q(\ram[10][15] ) );
  LATCHX1_HVT \ram_reg[10][14]  ( .CLK(n119), .D(N30), .Q(\ram[10][14] ) );
  LATCHX1_HVT \ram_reg[10][13]  ( .CLK(n118), .D(N29), .Q(\ram[10][13] ) );
  LATCHX1_HVT \ram_reg[10][12]  ( .CLK(n118), .D(N28), .Q(\ram[10][12] ) );
  LATCHX1_HVT \ram_reg[10][11]  ( .CLK(n119), .D(N27), .Q(\ram[10][11] ) );
  LATCHX1_HVT \ram_reg[10][10]  ( .CLK(n118), .D(N26), .Q(\ram[10][10] ) );
  LATCHX1_HVT \ram_reg[10][9]  ( .CLK(n118), .D(N25), .Q(\ram[10][9] ) );
  LATCHX1_HVT \ram_reg[10][8]  ( .CLK(n119), .D(N24), .Q(\ram[10][8] ) );
  LATCHX1_HVT \ram_reg[10][7]  ( .CLK(n122), .D(N23), .Q(\ram[10][7] ) );
  LATCHX1_HVT \ram_reg[10][6]  ( .CLK(n122), .D(N22), .Q(\ram[10][6] ) );
  LATCHX1_HVT \ram_reg[10][5]  ( .CLK(n121), .D(N21), .Q(\ram[10][5] ) );
  LATCHX1_HVT \ram_reg[10][4]  ( .CLK(n121), .D(N20), .Q(\ram[10][4] ) );
  LATCHX1_HVT \ram_reg[10][3]  ( .CLK(n120), .D(N19), .Q(\ram[10][3] ) );
  LATCHX1_HVT \ram_reg[10][2]  ( .CLK(n121), .D(N18), .Q(\ram[10][2] ) );
  LATCHX1_HVT \ram_reg[10][1]  ( .CLK(n122), .D(N17), .Q(\ram[10][1] ) );
  LATCHX1_HVT \ram_reg[10][0]  ( .CLK(n126), .D(N16), .Q(\ram[10][0] ) );
  LATCHX1_HVT \ram_reg[9][255]  ( .CLK(N300), .D(N273), .Q(\ram[9][255] ) );
  LATCHX1_HVT \ram_reg[9][254]  ( .CLK(N300), .D(N272), .Q(\ram[9][254] ) );
  LATCHX1_HVT \ram_reg[9][253]  ( .CLK(N300), .D(N271), .Q(\ram[9][253] ) );
  LATCHX1_HVT \ram_reg[9][252]  ( .CLK(N300), .D(N270), .Q(\ram[9][252] ) );
  LATCHX1_HVT \ram_reg[9][251]  ( .CLK(n159), .D(N269), .Q(\ram[9][251] ) );
  LATCHX1_HVT \ram_reg[9][250]  ( .CLK(n151), .D(N268), .Q(\ram[9][250] ) );
  LATCHX1_HVT \ram_reg[9][249]  ( .CLK(n151), .D(N267), .Q(\ram[9][249] ) );
  LATCHX1_HVT \ram_reg[9][248]  ( .CLK(n151), .D(N266), .Q(\ram[9][248] ) );
  LATCHX1_HVT \ram_reg[9][247]  ( .CLK(n151), .D(N265), .Q(\ram[9][247] ) );
  LATCHX1_HVT \ram_reg[9][246]  ( .CLK(n151), .D(N264), .Q(\ram[9][246] ) );
  LATCHX1_HVT \ram_reg[9][245]  ( .CLK(n151), .D(N263), .Q(\ram[9][245] ) );
  LATCHX1_HVT \ram_reg[9][244]  ( .CLK(n151), .D(N262), .Q(\ram[9][244] ) );
  LATCHX1_HVT \ram_reg[9][243]  ( .CLK(n151), .D(N261), .Q(\ram[9][243] ) );
  LATCHX1_HVT \ram_reg[9][242]  ( .CLK(n151), .D(N260), .Q(\ram[9][242] ) );
  LATCHX1_HVT \ram_reg[9][241]  ( .CLK(n150), .D(N259), .Q(\ram[9][241] ) );
  LATCHX1_HVT \ram_reg[9][240]  ( .CLK(n150), .D(N258), .Q(\ram[9][240] ) );
  LATCHX1_HVT \ram_reg[9][239]  ( .CLK(n150), .D(N257), .Q(\ram[9][239] ) );
  LATCHX1_HVT \ram_reg[9][238]  ( .CLK(n150), .D(N256), .Q(\ram[9][238] ) );
  LATCHX1_HVT \ram_reg[9][237]  ( .CLK(n150), .D(N255), .Q(\ram[9][237] ) );
  LATCHX1_HVT \ram_reg[9][236]  ( .CLK(n150), .D(N254), .Q(\ram[9][236] ) );
  LATCHX1_HVT \ram_reg[9][235]  ( .CLK(n150), .D(N253), .Q(\ram[9][235] ) );
  LATCHX1_HVT \ram_reg[9][234]  ( .CLK(n150), .D(N252), .Q(\ram[9][234] ) );
  LATCHX1_HVT \ram_reg[9][233]  ( .CLK(n150), .D(N251), .Q(\ram[9][233] ) );
  LATCHX1_HVT \ram_reg[9][232]  ( .CLK(n150), .D(N250), .Q(\ram[9][232] ) );
  LATCHX1_HVT \ram_reg[9][231]  ( .CLK(n150), .D(N249), .Q(\ram[9][231] ) );
  LATCHX1_HVT \ram_reg[9][230]  ( .CLK(n149), .D(N248), .Q(\ram[9][230] ) );
  LATCHX1_HVT \ram_reg[9][229]  ( .CLK(n149), .D(N247), .Q(\ram[9][229] ) );
  LATCHX1_HVT \ram_reg[9][228]  ( .CLK(n149), .D(N246), .Q(\ram[9][228] ) );
  LATCHX1_HVT \ram_reg[9][227]  ( .CLK(n159), .D(N245), .Q(\ram[9][227] ) );
  LATCHX1_HVT \ram_reg[9][226]  ( .CLK(n159), .D(N244), .Q(\ram[9][226] ) );
  LATCHX1_HVT \ram_reg[9][225]  ( .CLK(n159), .D(N243), .Q(\ram[9][225] ) );
  LATCHX1_HVT \ram_reg[9][224]  ( .CLK(n159), .D(N242), .Q(\ram[9][224] ) );
  LATCHX1_HVT \ram_reg[9][223]  ( .CLK(n159), .D(N241), .Q(\ram[9][223] ) );
  LATCHX1_HVT \ram_reg[9][222]  ( .CLK(n159), .D(N240), .Q(\ram[9][222] ) );
  LATCHX1_HVT \ram_reg[9][221]  ( .CLK(n159), .D(N239), .Q(\ram[9][221] ) );
  LATCHX1_HVT \ram_reg[9][220]  ( .CLK(n159), .D(N238), .Q(\ram[9][220] ) );
  LATCHX1_HVT \ram_reg[9][219]  ( .CLK(n159), .D(N237), .Q(\ram[9][219] ) );
  LATCHX1_HVT \ram_reg[9][218]  ( .CLK(n159), .D(N236), .Q(\ram[9][218] ) );
  LATCHX1_HVT \ram_reg[9][217]  ( .CLK(n158), .D(N235), .Q(\ram[9][217] ) );
  LATCHX1_HVT \ram_reg[9][216]  ( .CLK(n158), .D(N234), .Q(\ram[9][216] ) );
  LATCHX1_HVT \ram_reg[9][215]  ( .CLK(n158), .D(N233), .Q(\ram[9][215] ) );
  LATCHX1_HVT \ram_reg[9][214]  ( .CLK(n158), .D(N232), .Q(\ram[9][214] ) );
  LATCHX1_HVT \ram_reg[9][213]  ( .CLK(n158), .D(N231), .Q(\ram[9][213] ) );
  LATCHX1_HVT \ram_reg[9][212]  ( .CLK(n158), .D(N230), .Q(\ram[9][212] ) );
  LATCHX1_HVT \ram_reg[9][211]  ( .CLK(n158), .D(N229), .Q(\ram[9][211] ) );
  LATCHX1_HVT \ram_reg[9][210]  ( .CLK(n158), .D(N228), .Q(\ram[9][210] ) );
  LATCHX1_HVT \ram_reg[9][209]  ( .CLK(n158), .D(N227), .Q(\ram[9][209] ) );
  LATCHX1_HVT \ram_reg[9][208]  ( .CLK(n158), .D(N226), .Q(\ram[9][208] ) );
  LATCHX1_HVT \ram_reg[9][207]  ( .CLK(n157), .D(N225), .Q(\ram[9][207] ) );
  LATCHX1_HVT \ram_reg[9][206]  ( .CLK(n157), .D(N224), .Q(\ram[9][206] ) );
  LATCHX1_HVT \ram_reg[9][205]  ( .CLK(n157), .D(N223), .Q(\ram[9][205] ) );
  LATCHX1_HVT \ram_reg[9][204]  ( .CLK(n157), .D(N222), .Q(\ram[9][204] ) );
  LATCHX1_HVT \ram_reg[9][203]  ( .CLK(n157), .D(N221), .Q(\ram[9][203] ) );
  LATCHX1_HVT \ram_reg[9][202]  ( .CLK(n157), .D(N220), .Q(\ram[9][202] ) );
  LATCHX1_HVT \ram_reg[9][201]  ( .CLK(n157), .D(N219), .Q(\ram[9][201] ) );
  LATCHX1_HVT \ram_reg[9][200]  ( .CLK(n157), .D(N218), .Q(\ram[9][200] ) );
  LATCHX1_HVT \ram_reg[9][199]  ( .CLK(n157), .D(N217), .Q(\ram[9][199] ) );
  LATCHX1_HVT \ram_reg[9][198]  ( .CLK(n157), .D(N216), .Q(\ram[9][198] ) );
  LATCHX1_HVT \ram_reg[9][197]  ( .CLK(n157), .D(N214), .Q(\ram[9][197] ) );
  LATCHX1_HVT \ram_reg[9][196]  ( .CLK(n156), .D(N213), .Q(\ram[9][196] ) );
  LATCHX1_HVT \ram_reg[9][195]  ( .CLK(n156), .D(N212), .Q(\ram[9][195] ) );
  LATCHX1_HVT \ram_reg[9][194]  ( .CLK(n156), .D(N211), .Q(\ram[9][194] ) );
  LATCHX1_HVT \ram_reg[9][193]  ( .CLK(n156), .D(N210), .Q(\ram[9][193] ) );
  LATCHX1_HVT \ram_reg[9][192]  ( .CLK(n156), .D(N209), .Q(\ram[9][192] ) );
  LATCHX1_HVT \ram_reg[9][191]  ( .CLK(n156), .D(N208), .Q(\ram[9][191] ) );
  LATCHX1_HVT \ram_reg[9][190]  ( .CLK(n156), .D(N207), .Q(\ram[9][190] ) );
  LATCHX1_HVT \ram_reg[9][189]  ( .CLK(n156), .D(N206), .Q(\ram[9][189] ) );
  LATCHX1_HVT \ram_reg[9][188]  ( .CLK(n156), .D(N205), .Q(\ram[9][188] ) );
  LATCHX1_HVT \ram_reg[9][187]  ( .CLK(n156), .D(N204), .Q(\ram[9][187] ) );
  LATCHX1_HVT \ram_reg[9][186]  ( .CLK(n156), .D(N203), .Q(\ram[9][186] ) );
  LATCHX1_HVT \ram_reg[9][185]  ( .CLK(n155), .D(N202), .Q(\ram[9][185] ) );
  LATCHX1_HVT \ram_reg[9][184]  ( .CLK(n155), .D(N201), .Q(\ram[9][184] ) );
  LATCHX1_HVT \ram_reg[9][183]  ( .CLK(n155), .D(N200), .Q(\ram[9][183] ) );
  LATCHX1_HVT \ram_reg[9][182]  ( .CLK(n155), .D(N199), .Q(\ram[9][182] ) );
  LATCHX1_HVT \ram_reg[9][181]  ( .CLK(n155), .D(N198), .Q(\ram[9][181] ) );
  LATCHX1_HVT \ram_reg[9][180]  ( .CLK(n155), .D(N197), .Q(\ram[9][180] ) );
  LATCHX1_HVT \ram_reg[9][179]  ( .CLK(n155), .D(N196), .Q(\ram[9][179] ) );
  LATCHX1_HVT \ram_reg[9][178]  ( .CLK(n155), .D(N195), .Q(\ram[9][178] ) );
  LATCHX1_HVT \ram_reg[9][177]  ( .CLK(n155), .D(N194), .Q(\ram[9][177] ) );
  LATCHX1_HVT \ram_reg[9][176]  ( .CLK(n155), .D(N193), .Q(\ram[9][176] ) );
  LATCHX1_HVT \ram_reg[9][175]  ( .CLK(n155), .D(N192), .Q(\ram[9][175] ) );
  LATCHX1_HVT \ram_reg[9][174]  ( .CLK(n154), .D(N191), .Q(\ram[9][174] ) );
  LATCHX1_HVT \ram_reg[9][173]  ( .CLK(n154), .D(N190), .Q(\ram[9][173] ) );
  LATCHX1_HVT \ram_reg[9][172]  ( .CLK(n154), .D(N189), .Q(\ram[9][172] ) );
  LATCHX1_HVT \ram_reg[9][171]  ( .CLK(n154), .D(N188), .Q(\ram[9][171] ) );
  LATCHX1_HVT \ram_reg[9][170]  ( .CLK(n154), .D(N187), .Q(\ram[9][170] ) );
  LATCHX1_HVT \ram_reg[9][169]  ( .CLK(n154), .D(N186), .Q(\ram[9][169] ) );
  LATCHX1_HVT \ram_reg[9][168]  ( .CLK(n154), .D(N185), .Q(\ram[9][168] ) );
  LATCHX1_HVT \ram_reg[9][167]  ( .CLK(n154), .D(N184), .Q(\ram[9][167] ) );
  LATCHX1_HVT \ram_reg[9][166]  ( .CLK(n154), .D(N183), .Q(\ram[9][166] ) );
  LATCHX1_HVT \ram_reg[9][165]  ( .CLK(n154), .D(N182), .Q(\ram[9][165] ) );
  LATCHX1_HVT \ram_reg[9][164]  ( .CLK(n154), .D(N181), .Q(\ram[9][164] ) );
  LATCHX1_HVT \ram_reg[9][163]  ( .CLK(n153), .D(N180), .Q(\ram[9][163] ) );
  LATCHX1_HVT \ram_reg[9][162]  ( .CLK(n153), .D(N179), .Q(\ram[9][162] ) );
  LATCHX1_HVT \ram_reg[9][161]  ( .CLK(n153), .D(N178), .Q(\ram[9][161] ) );
  LATCHX1_HVT \ram_reg[9][160]  ( .CLK(n153), .D(N177), .Q(\ram[9][160] ) );
  LATCHX1_HVT \ram_reg[9][159]  ( .CLK(n153), .D(N176), .Q(\ram[9][159] ) );
  LATCHX1_HVT \ram_reg[9][158]  ( .CLK(n153), .D(N175), .Q(\ram[9][158] ) );
  LATCHX1_HVT \ram_reg[9][157]  ( .CLK(n153), .D(N174), .Q(\ram[9][157] ) );
  LATCHX1_HVT \ram_reg[9][156]  ( .CLK(n153), .D(N173), .Q(\ram[9][156] ) );
  LATCHX1_HVT \ram_reg[9][155]  ( .CLK(n153), .D(N172), .Q(\ram[9][155] ) );
  LATCHX1_HVT \ram_reg[9][154]  ( .CLK(n153), .D(N171), .Q(\ram[9][154] ) );
  LATCHX1_HVT \ram_reg[9][153]  ( .CLK(n153), .D(N170), .Q(\ram[9][153] ) );
  LATCHX1_HVT \ram_reg[9][152]  ( .CLK(n152), .D(N169), .Q(\ram[9][152] ) );
  LATCHX1_HVT \ram_reg[9][151]  ( .CLK(n152), .D(N168), .Q(\ram[9][151] ) );
  LATCHX1_HVT \ram_reg[9][150]  ( .CLK(n152), .D(N167), .Q(\ram[9][150] ) );
  LATCHX1_HVT \ram_reg[9][149]  ( .CLK(n152), .D(N166), .Q(\ram[9][149] ) );
  LATCHX1_HVT \ram_reg[9][148]  ( .CLK(n152), .D(N165), .Q(\ram[9][148] ) );
  LATCHX1_HVT \ram_reg[9][147]  ( .CLK(n152), .D(N164), .Q(\ram[9][147] ) );
  LATCHX1_HVT \ram_reg[9][146]  ( .CLK(n152), .D(N163), .Q(\ram[9][146] ) );
  LATCHX1_HVT \ram_reg[9][145]  ( .CLK(n152), .D(N162), .Q(\ram[9][145] ) );
  LATCHX1_HVT \ram_reg[9][144]  ( .CLK(n152), .D(N161), .Q(\ram[9][144] ) );
  LATCHX1_HVT \ram_reg[9][143]  ( .CLK(n152), .D(N160), .Q(\ram[9][143] ) );
  LATCHX1_HVT \ram_reg[9][142]  ( .CLK(n152), .D(N159), .Q(\ram[9][142] ) );
  LATCHX1_HVT \ram_reg[9][141]  ( .CLK(n151), .D(N158), .Q(\ram[9][141] ) );
  LATCHX1_HVT \ram_reg[9][140]  ( .CLK(n151), .D(N157), .Q(\ram[9][140] ) );
  LATCHX1_HVT \ram_reg[9][139]  ( .CLK(n151), .D(N156), .Q(\ram[9][139] ) );
  LATCHX1_HVT \ram_reg[9][138]  ( .CLK(n150), .D(N155), .Q(\ram[9][138] ) );
  LATCHX1_HVT \ram_reg[9][137]  ( .CLK(n159), .D(N154), .Q(\ram[9][137] ) );
  LATCHX1_HVT \ram_reg[9][136]  ( .CLK(n158), .D(N153), .Q(\ram[9][136] ) );
  LATCHX1_HVT \ram_reg[9][135]  ( .CLK(n158), .D(N152), .Q(\ram[9][135] ) );
  LATCHX1_HVT \ram_reg[9][134]  ( .CLK(n157), .D(N151), .Q(\ram[9][134] ) );
  LATCHX1_HVT \ram_reg[9][133]  ( .CLK(n156), .D(N150), .Q(\ram[9][133] ) );
  LATCHX1_HVT \ram_reg[9][132]  ( .CLK(n155), .D(N149), .Q(\ram[9][132] ) );
  LATCHX1_HVT \ram_reg[9][131]  ( .CLK(n154), .D(N148), .Q(\ram[9][131] ) );
  LATCHX1_HVT \ram_reg[9][130]  ( .CLK(n153), .D(N147), .Q(\ram[9][130] ) );
  LATCHX1_HVT \ram_reg[9][129]  ( .CLK(n152), .D(N146), .Q(\ram[9][129] ) );
  LATCHX1_HVT \ram_reg[9][128]  ( .CLK(n149), .D(N145), .Q(\ram[9][128] ) );
  LATCHX1_HVT \ram_reg[9][127]  ( .CLK(n140), .D(N144), .Q(\ram[9][127] ) );
  LATCHX1_HVT \ram_reg[9][126]  ( .CLK(n140), .D(N143), .Q(\ram[9][126] ) );
  LATCHX1_HVT \ram_reg[9][125]  ( .CLK(n140), .D(N142), .Q(\ram[9][125] ) );
  LATCHX1_HVT \ram_reg[9][124]  ( .CLK(n140), .D(N141), .Q(\ram[9][124] ) );
  LATCHX1_HVT \ram_reg[9][123]  ( .CLK(n140), .D(N140), .Q(\ram[9][123] ) );
  LATCHX1_HVT \ram_reg[9][122]  ( .CLK(n139), .D(N139), .Q(\ram[9][122] ) );
  LATCHX1_HVT \ram_reg[9][121]  ( .CLK(n140), .D(N138), .Q(\ram[9][121] ) );
  LATCHX1_HVT \ram_reg[9][120]  ( .CLK(n140), .D(N137), .Q(\ram[9][120] ) );
  LATCHX1_HVT \ram_reg[9][119]  ( .CLK(n149), .D(N136), .Q(\ram[9][119] ) );
  LATCHX1_HVT \ram_reg[9][118]  ( .CLK(n148), .D(N135), .Q(\ram[9][118] ) );
  LATCHX1_HVT \ram_reg[9][117]  ( .CLK(n148), .D(N134), .Q(\ram[9][117] ) );
  LATCHX1_HVT \ram_reg[9][116]  ( .CLK(n147), .D(N133), .Q(\ram[9][116] ) );
  LATCHX1_HVT \ram_reg[9][115]  ( .CLK(n142), .D(N132), .Q(\ram[9][115] ) );
  LATCHX1_HVT \ram_reg[9][114]  ( .CLK(n147), .D(N131), .Q(\ram[9][114] ) );
  LATCHX1_HVT \ram_reg[9][113]  ( .CLK(n147), .D(N130), .Q(\ram[9][113] ) );
  LATCHX1_HVT \ram_reg[9][112]  ( .CLK(n148), .D(N129), .Q(\ram[9][112] ) );
  LATCHX1_HVT \ram_reg[9][111]  ( .CLK(n146), .D(N128), .Q(\ram[9][111] ) );
  LATCHX1_HVT \ram_reg[9][110]  ( .CLK(n146), .D(N127), .Q(\ram[9][110] ) );
  LATCHX1_HVT \ram_reg[9][109]  ( .CLK(n146), .D(N126), .Q(\ram[9][109] ) );
  LATCHX1_HVT \ram_reg[9][108]  ( .CLK(n143), .D(N125), .Q(\ram[9][108] ) );
  LATCHX1_HVT \ram_reg[9][107]  ( .CLK(n140), .D(N124), .Q(\ram[9][107] ) );
  LATCHX1_HVT \ram_reg[9][106]  ( .CLK(n146), .D(N123), .Q(\ram[9][106] ) );
  LATCHX1_HVT \ram_reg[9][105]  ( .CLK(n146), .D(N122), .Q(\ram[9][105] ) );
  LATCHX1_HVT \ram_reg[9][104]  ( .CLK(n146), .D(N121), .Q(\ram[9][104] ) );
  LATCHX1_HVT \ram_reg[9][103]  ( .CLK(n145), .D(N120), .Q(\ram[9][103] ) );
  LATCHX1_HVT \ram_reg[9][102]  ( .CLK(n144), .D(N119), .Q(\ram[9][102] ) );
  LATCHX1_HVT \ram_reg[9][101]  ( .CLK(n144), .D(N118), .Q(\ram[9][101] ) );
  LATCHX1_HVT \ram_reg[9][100]  ( .CLK(n145), .D(N117), .Q(\ram[9][100] ) );
  LATCHX1_HVT \ram_reg[9][99]  ( .CLK(n143), .D(N116), .Q(\ram[9][99] ) );
  LATCHX1_HVT \ram_reg[9][98]  ( .CLK(n144), .D(N114), .Q(\ram[9][98] ) );
  LATCHX1_HVT \ram_reg[9][97]  ( .CLK(n145), .D(N113), .Q(\ram[9][97] ) );
  LATCHX1_HVT \ram_reg[9][96]  ( .CLK(n149), .D(N112), .Q(\ram[9][96] ) );
  LATCHX1_HVT \ram_reg[9][95]  ( .CLK(n141), .D(N111), .Q(\ram[9][95] ) );
  LATCHX1_HVT \ram_reg[9][94]  ( .CLK(n141), .D(N110), .Q(\ram[9][94] ) );
  LATCHX1_HVT \ram_reg[9][93]  ( .CLK(n141), .D(N109), .Q(\ram[9][93] ) );
  LATCHX1_HVT \ram_reg[9][92]  ( .CLK(n140), .D(N108), .Q(\ram[9][92] ) );
  LATCHX1_HVT \ram_reg[9][91]  ( .CLK(n140), .D(N107), .Q(\ram[9][91] ) );
  LATCHX1_HVT \ram_reg[9][90]  ( .CLK(n141), .D(N106), .Q(\ram[9][90] ) );
  LATCHX1_HVT \ram_reg[9][89]  ( .CLK(n140), .D(N105), .Q(\ram[9][89] ) );
  LATCHX1_HVT \ram_reg[9][88]  ( .CLK(n141), .D(N104), .Q(\ram[9][88] ) );
  LATCHX1_HVT \ram_reg[9][87]  ( .CLK(n149), .D(N103), .Q(\ram[9][87] ) );
  LATCHX1_HVT \ram_reg[9][86]  ( .CLK(n148), .D(N102), .Q(\ram[9][86] ) );
  LATCHX1_HVT \ram_reg[9][85]  ( .CLK(n147), .D(N101), .Q(\ram[9][85] ) );
  LATCHX1_HVT \ram_reg[9][84]  ( .CLK(n147), .D(N100), .Q(\ram[9][84] ) );
  LATCHX1_HVT \ram_reg[9][83]  ( .CLK(n142), .D(N99), .Q(\ram[9][83] ) );
  LATCHX1_HVT \ram_reg[9][82]  ( .CLK(n148), .D(N98), .Q(\ram[9][82] ) );
  LATCHX1_HVT \ram_reg[9][81]  ( .CLK(n147), .D(N97), .Q(\ram[9][81] ) );
  LATCHX1_HVT \ram_reg[9][80]  ( .CLK(n148), .D(N96), .Q(\ram[9][80] ) );
  LATCHX1_HVT \ram_reg[9][79]  ( .CLK(n142), .D(N95), .Q(\ram[9][79] ) );
  LATCHX1_HVT \ram_reg[9][78]  ( .CLK(n141), .D(N94), .Q(\ram[9][78] ) );
  LATCHX1_HVT \ram_reg[9][77]  ( .CLK(n142), .D(N93), .Q(\ram[9][77] ) );
  LATCHX1_HVT \ram_reg[9][76]  ( .CLK(n141), .D(N92), .Q(\ram[9][76] ) );
  LATCHX1_HVT \ram_reg[9][75]  ( .CLK(n141), .D(N91), .Q(\ram[9][75] ) );
  LATCHX1_HVT \ram_reg[9][74]  ( .CLK(n139), .D(N90), .Q(\ram[9][74] ) );
  LATCHX1_HVT \ram_reg[9][73]  ( .CLK(n142), .D(N89), .Q(\ram[9][73] ) );
  LATCHX1_HVT \ram_reg[9][72]  ( .CLK(n142), .D(N88), .Q(\ram[9][72] ) );
  LATCHX1_HVT \ram_reg[9][71]  ( .CLK(n145), .D(N87), .Q(\ram[9][71] ) );
  LATCHX1_HVT \ram_reg[9][70]  ( .CLK(n145), .D(N86), .Q(\ram[9][70] ) );
  LATCHX1_HVT \ram_reg[9][69]  ( .CLK(n144), .D(N85), .Q(\ram[9][69] ) );
  LATCHX1_HVT \ram_reg[9][68]  ( .CLK(n145), .D(N84), .Q(\ram[9][68] ) );
  LATCHX1_HVT \ram_reg[9][67]  ( .CLK(n144), .D(N83), .Q(\ram[9][67] ) );
  LATCHX1_HVT \ram_reg[9][66]  ( .CLK(n143), .D(N82), .Q(\ram[9][66] ) );
  LATCHX1_HVT \ram_reg[9][65]  ( .CLK(n144), .D(N81), .Q(\ram[9][65] ) );
  LATCHX1_HVT \ram_reg[9][64]  ( .CLK(n149), .D(N80), .Q(\ram[9][64] ) );
  LATCHX1_HVT \ram_reg[9][63]  ( .CLK(n143), .D(N79), .Q(\ram[9][63] ) );
  LATCHX1_HVT \ram_reg[9][62]  ( .CLK(n143), .D(N78), .Q(\ram[9][62] ) );
  LATCHX1_HVT \ram_reg[9][61]  ( .CLK(n143), .D(N77), .Q(\ram[9][61] ) );
  LATCHX1_HVT \ram_reg[9][60]  ( .CLK(n143), .D(N76), .Q(\ram[9][60] ) );
  LATCHX1_HVT \ram_reg[9][59]  ( .CLK(n143), .D(N75), .Q(\ram[9][59] ) );
  LATCHX1_HVT \ram_reg[9][58]  ( .CLK(n142), .D(N74), .Q(\ram[9][58] ) );
  LATCHX1_HVT \ram_reg[9][57]  ( .CLK(n143), .D(N73), .Q(\ram[9][57] ) );
  LATCHX1_HVT \ram_reg[9][56]  ( .CLK(n143), .D(N72), .Q(\ram[9][56] ) );
  LATCHX1_HVT \ram_reg[9][55]  ( .CLK(n149), .D(N71), .Q(\ram[9][55] ) );
  LATCHX1_HVT \ram_reg[9][54]  ( .CLK(n147), .D(N70), .Q(\ram[9][54] ) );
  LATCHX1_HVT \ram_reg[9][53]  ( .CLK(n147), .D(N69), .Q(\ram[9][53] ) );
  LATCHX1_HVT \ram_reg[9][52]  ( .CLK(n148), .D(N68), .Q(\ram[9][52] ) );
  LATCHX1_HVT \ram_reg[9][51]  ( .CLK(n142), .D(N67), .Q(\ram[9][51] ) );
  LATCHX1_HVT \ram_reg[9][50]  ( .CLK(n139), .D(N66), .Q(\ram[9][50] ) );
  LATCHX1_HVT \ram_reg[9][49]  ( .CLK(n148), .D(N65), .Q(\ram[9][49] ) );
  LATCHX1_HVT \ram_reg[9][48]  ( .CLK(n148), .D(N64), .Q(\ram[9][48] ) );
  LATCHX1_HVT \ram_reg[9][47]  ( .CLK(n146), .D(N63), .Q(\ram[9][47] ) );
  LATCHX1_HVT \ram_reg[9][46]  ( .CLK(n146), .D(N62), .Q(\ram[9][46] ) );
  LATCHX1_HVT \ram_reg[9][45]  ( .CLK(n146), .D(N61), .Q(\ram[9][45] ) );
  LATCHX1_HVT \ram_reg[9][44]  ( .CLK(n146), .D(N60), .Q(\ram[9][44] ) );
  LATCHX1_HVT \ram_reg[9][43]  ( .CLK(n143), .D(N59), .Q(\ram[9][43] ) );
  LATCHX1_HVT \ram_reg[9][42]  ( .CLK(n147), .D(N58), .Q(\ram[9][42] ) );
  LATCHX1_HVT \ram_reg[9][41]  ( .CLK(n140), .D(N57), .Q(\ram[9][41] ) );
  LATCHX1_HVT \ram_reg[9][40]  ( .CLK(n146), .D(N56), .Q(\ram[9][40] ) );
  LATCHX1_HVT \ram_reg[9][39]  ( .CLK(n145), .D(N55), .Q(\ram[9][39] ) );
  LATCHX1_HVT \ram_reg[9][38]  ( .CLK(n145), .D(N54), .Q(\ram[9][38] ) );
  LATCHX1_HVT \ram_reg[9][37]  ( .CLK(n144), .D(N53), .Q(\ram[9][37] ) );
  LATCHX1_HVT \ram_reg[9][36]  ( .CLK(n144), .D(N52), .Q(\ram[9][36] ) );
  LATCHX1_HVT \ram_reg[9][35]  ( .CLK(n144), .D(N51), .Q(\ram[9][35] ) );
  LATCHX1_HVT \ram_reg[9][34]  ( .CLK(n146), .D(N50), .Q(\ram[9][34] ) );
  LATCHX1_HVT \ram_reg[9][33]  ( .CLK(n145), .D(N49), .Q(\ram[9][33] ) );
  LATCHX1_HVT \ram_reg[9][32]  ( .CLK(n149), .D(N48), .Q(\ram[9][32] ) );
  LATCHX1_HVT \ram_reg[9][31]  ( .CLK(n139), .D(N47), .Q(\ram[9][31] ) );
  LATCHX1_HVT \ram_reg[9][30]  ( .CLK(n139), .D(N46), .Q(\ram[9][30] ) );
  LATCHX1_HVT \ram_reg[9][29]  ( .CLK(n139), .D(N45), .Q(\ram[9][29] ) );
  LATCHX1_HVT \ram_reg[9][28]  ( .CLK(n139), .D(N44), .Q(\ram[9][28] ) );
  LATCHX1_HVT \ram_reg[9][27]  ( .CLK(n139), .D(N43), .Q(\ram[9][27] ) );
  LATCHX1_HVT \ram_reg[9][26]  ( .CLK(n139), .D(N42), .Q(\ram[9][26] ) );
  LATCHX1_HVT \ram_reg[9][25]  ( .CLK(n139), .D(N41), .Q(\ram[9][25] ) );
  LATCHX1_HVT \ram_reg[9][24]  ( .CLK(n139), .D(N40), .Q(\ram[9][24] ) );
  LATCHX1_HVT \ram_reg[9][23]  ( .CLK(n149), .D(N39), .Q(\ram[9][23] ) );
  LATCHX1_HVT \ram_reg[9][22]  ( .CLK(n148), .D(N38), .Q(\ram[9][22] ) );
  LATCHX1_HVT \ram_reg[9][21]  ( .CLK(n147), .D(N37), .Q(\ram[9][21] ) );
  LATCHX1_HVT \ram_reg[9][20]  ( .CLK(n147), .D(N36), .Q(\ram[9][20] ) );
  LATCHX1_HVT \ram_reg[9][19]  ( .CLK(n139), .D(N35), .Q(\ram[9][19] ) );
  LATCHX1_HVT \ram_reg[9][18]  ( .CLK(n147), .D(N34), .Q(\ram[9][18] ) );
  LATCHX1_HVT \ram_reg[9][17]  ( .CLK(n148), .D(N33), .Q(\ram[9][17] ) );
  LATCHX1_HVT \ram_reg[9][16]  ( .CLK(n148), .D(N32), .Q(\ram[9][16] ) );
  LATCHX1_HVT \ram_reg[9][15]  ( .CLK(n142), .D(N31), .Q(\ram[9][15] ) );
  LATCHX1_HVT \ram_reg[9][14]  ( .CLK(n142), .D(N30), .Q(\ram[9][14] ) );
  LATCHX1_HVT \ram_reg[9][13]  ( .CLK(n141), .D(N29), .Q(\ram[9][13] ) );
  LATCHX1_HVT \ram_reg[9][12]  ( .CLK(n141), .D(N28), .Q(\ram[9][12] ) );
  LATCHX1_HVT \ram_reg[9][11]  ( .CLK(n142), .D(N27), .Q(\ram[9][11] ) );
  LATCHX1_HVT \ram_reg[9][10]  ( .CLK(n141), .D(N26), .Q(\ram[9][10] ) );
  LATCHX1_HVT \ram_reg[9][9]  ( .CLK(n141), .D(N25), .Q(\ram[9][9] ) );
  LATCHX1_HVT \ram_reg[9][8]  ( .CLK(n142), .D(N24), .Q(\ram[9][8] ) );
  LATCHX1_HVT \ram_reg[9][7]  ( .CLK(n145), .D(N23), .Q(\ram[9][7] ) );
  LATCHX1_HVT \ram_reg[9][6]  ( .CLK(n145), .D(N22), .Q(\ram[9][6] ) );
  LATCHX1_HVT \ram_reg[9][5]  ( .CLK(n144), .D(N21), .Q(\ram[9][5] ) );
  LATCHX1_HVT \ram_reg[9][4]  ( .CLK(n144), .D(N20), .Q(\ram[9][4] ) );
  LATCHX1_HVT \ram_reg[9][3]  ( .CLK(n143), .D(N19), .Q(\ram[9][3] ) );
  LATCHX1_HVT \ram_reg[9][2]  ( .CLK(n144), .D(N18), .Q(\ram[9][2] ) );
  LATCHX1_HVT \ram_reg[9][1]  ( .CLK(n145), .D(N17), .Q(\ram[9][1] ) );
  LATCHX1_HVT \ram_reg[9][0]  ( .CLK(n149), .D(N16), .Q(\ram[9][0] ) );
  LATCHX1_HVT \ram_reg[8][255]  ( .CLK(N297), .D(N273), .Q(\ram[8][255] ) );
  LATCHX1_HVT \ram_reg[8][254]  ( .CLK(N297), .D(N272), .Q(\ram[8][254] ) );
  LATCHX1_HVT \ram_reg[8][253]  ( .CLK(N297), .D(N271), .Q(\ram[8][253] ) );
  LATCHX1_HVT \ram_reg[8][252]  ( .CLK(N297), .D(N270), .Q(\ram[8][252] ) );
  LATCHX1_HVT \ram_reg[8][251]  ( .CLK(n182), .D(N269), .Q(\ram[8][251] ) );
  LATCHX1_HVT \ram_reg[8][250]  ( .CLK(n174), .D(N268), .Q(\ram[8][250] ) );
  LATCHX1_HVT \ram_reg[8][249]  ( .CLK(n174), .D(N267), .Q(\ram[8][249] ) );
  LATCHX1_HVT \ram_reg[8][248]  ( .CLK(n174), .D(N266), .Q(\ram[8][248] ) );
  LATCHX1_HVT \ram_reg[8][247]  ( .CLK(n174), .D(N265), .Q(\ram[8][247] ) );
  LATCHX1_HVT \ram_reg[8][246]  ( .CLK(n174), .D(N264), .Q(\ram[8][246] ) );
  LATCHX1_HVT \ram_reg[8][245]  ( .CLK(n174), .D(N263), .Q(\ram[8][245] ) );
  LATCHX1_HVT \ram_reg[8][244]  ( .CLK(n174), .D(N262), .Q(\ram[8][244] ) );
  LATCHX1_HVT \ram_reg[8][243]  ( .CLK(n174), .D(N261), .Q(\ram[8][243] ) );
  LATCHX1_HVT \ram_reg[8][242]  ( .CLK(n174), .D(N260), .Q(\ram[8][242] ) );
  LATCHX1_HVT \ram_reg[8][241]  ( .CLK(n173), .D(N259), .Q(\ram[8][241] ) );
  LATCHX1_HVT \ram_reg[8][240]  ( .CLK(n173), .D(N258), .Q(\ram[8][240] ) );
  LATCHX1_HVT \ram_reg[8][239]  ( .CLK(n173), .D(N257), .Q(\ram[8][239] ) );
  LATCHX1_HVT \ram_reg[8][238]  ( .CLK(n173), .D(N256), .Q(\ram[8][238] ) );
  LATCHX1_HVT \ram_reg[8][237]  ( .CLK(n173), .D(N255), .Q(\ram[8][237] ) );
  LATCHX1_HVT \ram_reg[8][236]  ( .CLK(n173), .D(N254), .Q(\ram[8][236] ) );
  LATCHX1_HVT \ram_reg[8][235]  ( .CLK(n173), .D(N253), .Q(\ram[8][235] ) );
  LATCHX1_HVT \ram_reg[8][234]  ( .CLK(n173), .D(N252), .Q(\ram[8][234] ) );
  LATCHX1_HVT \ram_reg[8][233]  ( .CLK(n173), .D(N251), .Q(\ram[8][233] ) );
  LATCHX1_HVT \ram_reg[8][232]  ( .CLK(n173), .D(N250), .Q(\ram[8][232] ) );
  LATCHX1_HVT \ram_reg[8][231]  ( .CLK(n173), .D(N249), .Q(\ram[8][231] ) );
  LATCHX1_HVT \ram_reg[8][230]  ( .CLK(n172), .D(N248), .Q(\ram[8][230] ) );
  LATCHX1_HVT \ram_reg[8][229]  ( .CLK(n172), .D(N247), .Q(\ram[8][229] ) );
  LATCHX1_HVT \ram_reg[8][228]  ( .CLK(n172), .D(N246), .Q(\ram[8][228] ) );
  LATCHX1_HVT \ram_reg[8][227]  ( .CLK(n182), .D(N245), .Q(\ram[8][227] ) );
  LATCHX1_HVT \ram_reg[8][226]  ( .CLK(n182), .D(N244), .Q(\ram[8][226] ) );
  LATCHX1_HVT \ram_reg[8][225]  ( .CLK(n182), .D(N243), .Q(\ram[8][225] ) );
  LATCHX1_HVT \ram_reg[8][224]  ( .CLK(n182), .D(N242), .Q(\ram[8][224] ) );
  LATCHX1_HVT \ram_reg[8][223]  ( .CLK(n182), .D(N241), .Q(\ram[8][223] ) );
  LATCHX1_HVT \ram_reg[8][222]  ( .CLK(n182), .D(N240), .Q(\ram[8][222] ) );
  LATCHX1_HVT \ram_reg[8][221]  ( .CLK(n182), .D(N239), .Q(\ram[8][221] ) );
  LATCHX1_HVT \ram_reg[8][220]  ( .CLK(n182), .D(N238), .Q(\ram[8][220] ) );
  LATCHX1_HVT \ram_reg[8][219]  ( .CLK(n182), .D(N237), .Q(\ram[8][219] ) );
  LATCHX1_HVT \ram_reg[8][218]  ( .CLK(n182), .D(N236), .Q(\ram[8][218] ) );
  LATCHX1_HVT \ram_reg[8][217]  ( .CLK(n181), .D(N235), .Q(\ram[8][217] ) );
  LATCHX1_HVT \ram_reg[8][216]  ( .CLK(n181), .D(N234), .Q(\ram[8][216] ) );
  LATCHX1_HVT \ram_reg[8][215]  ( .CLK(n181), .D(N233), .Q(\ram[8][215] ) );
  LATCHX1_HVT \ram_reg[8][214]  ( .CLK(n181), .D(N232), .Q(\ram[8][214] ) );
  LATCHX1_HVT \ram_reg[8][213]  ( .CLK(n181), .D(N231), .Q(\ram[8][213] ) );
  LATCHX1_HVT \ram_reg[8][212]  ( .CLK(n181), .D(N230), .Q(\ram[8][212] ) );
  LATCHX1_HVT \ram_reg[8][211]  ( .CLK(n181), .D(N229), .Q(\ram[8][211] ) );
  LATCHX1_HVT \ram_reg[8][210]  ( .CLK(n181), .D(N228), .Q(\ram[8][210] ) );
  LATCHX1_HVT \ram_reg[8][209]  ( .CLK(n181), .D(N227), .Q(\ram[8][209] ) );
  LATCHX1_HVT \ram_reg[8][208]  ( .CLK(n181), .D(N226), .Q(\ram[8][208] ) );
  LATCHX1_HVT \ram_reg[8][207]  ( .CLK(n180), .D(N225), .Q(\ram[8][207] ) );
  LATCHX1_HVT \ram_reg[8][206]  ( .CLK(n180), .D(N224), .Q(\ram[8][206] ) );
  LATCHX1_HVT \ram_reg[8][205]  ( .CLK(n180), .D(N223), .Q(\ram[8][205] ) );
  LATCHX1_HVT \ram_reg[8][204]  ( .CLK(n180), .D(N222), .Q(\ram[8][204] ) );
  LATCHX1_HVT \ram_reg[8][203]  ( .CLK(n180), .D(N221), .Q(\ram[8][203] ) );
  LATCHX1_HVT \ram_reg[8][202]  ( .CLK(n180), .D(N220), .Q(\ram[8][202] ) );
  LATCHX1_HVT \ram_reg[8][201]  ( .CLK(n180), .D(N219), .Q(\ram[8][201] ) );
  LATCHX1_HVT \ram_reg[8][200]  ( .CLK(n180), .D(N218), .Q(\ram[8][200] ) );
  LATCHX1_HVT \ram_reg[8][199]  ( .CLK(n180), .D(N217), .Q(\ram[8][199] ) );
  LATCHX1_HVT \ram_reg[8][198]  ( .CLK(n180), .D(N216), .Q(\ram[8][198] ) );
  LATCHX1_HVT \ram_reg[8][197]  ( .CLK(n180), .D(N214), .Q(\ram[8][197] ) );
  LATCHX1_HVT \ram_reg[8][196]  ( .CLK(n179), .D(N213), .Q(\ram[8][196] ) );
  LATCHX1_HVT \ram_reg[8][195]  ( .CLK(n179), .D(N212), .Q(\ram[8][195] ) );
  LATCHX1_HVT \ram_reg[8][194]  ( .CLK(n179), .D(N211), .Q(\ram[8][194] ) );
  LATCHX1_HVT \ram_reg[8][193]  ( .CLK(n179), .D(N210), .Q(\ram[8][193] ) );
  LATCHX1_HVT \ram_reg[8][192]  ( .CLK(n179), .D(N209), .Q(\ram[8][192] ) );
  LATCHX1_HVT \ram_reg[8][191]  ( .CLK(n179), .D(N208), .Q(\ram[8][191] ) );
  LATCHX1_HVT \ram_reg[8][190]  ( .CLK(n179), .D(N207), .Q(\ram[8][190] ) );
  LATCHX1_HVT \ram_reg[8][189]  ( .CLK(n179), .D(N206), .Q(\ram[8][189] ) );
  LATCHX1_HVT \ram_reg[8][188]  ( .CLK(n179), .D(N205), .Q(\ram[8][188] ) );
  LATCHX1_HVT \ram_reg[8][187]  ( .CLK(n179), .D(N204), .Q(\ram[8][187] ) );
  LATCHX1_HVT \ram_reg[8][186]  ( .CLK(n179), .D(N203), .Q(\ram[8][186] ) );
  LATCHX1_HVT \ram_reg[8][185]  ( .CLK(n178), .D(N202), .Q(\ram[8][185] ) );
  LATCHX1_HVT \ram_reg[8][184]  ( .CLK(n178), .D(N201), .Q(\ram[8][184] ) );
  LATCHX1_HVT \ram_reg[8][183]  ( .CLK(n178), .D(N200), .Q(\ram[8][183] ) );
  LATCHX1_HVT \ram_reg[8][182]  ( .CLK(n178), .D(N199), .Q(\ram[8][182] ) );
  LATCHX1_HVT \ram_reg[8][181]  ( .CLK(n178), .D(N198), .Q(\ram[8][181] ) );
  LATCHX1_HVT \ram_reg[8][180]  ( .CLK(n178), .D(N197), .Q(\ram[8][180] ) );
  LATCHX1_HVT \ram_reg[8][179]  ( .CLK(n178), .D(N196), .Q(\ram[8][179] ) );
  LATCHX1_HVT \ram_reg[8][178]  ( .CLK(n178), .D(N195), .Q(\ram[8][178] ) );
  LATCHX1_HVT \ram_reg[8][177]  ( .CLK(n178), .D(N194), .Q(\ram[8][177] ) );
  LATCHX1_HVT \ram_reg[8][176]  ( .CLK(n178), .D(N193), .Q(\ram[8][176] ) );
  LATCHX1_HVT \ram_reg[8][175]  ( .CLK(n178), .D(N192), .Q(\ram[8][175] ) );
  LATCHX1_HVT \ram_reg[8][174]  ( .CLK(n177), .D(N191), .Q(\ram[8][174] ) );
  LATCHX1_HVT \ram_reg[8][173]  ( .CLK(n177), .D(N190), .Q(\ram[8][173] ) );
  LATCHX1_HVT \ram_reg[8][172]  ( .CLK(n177), .D(N189), .Q(\ram[8][172] ) );
  LATCHX1_HVT \ram_reg[8][171]  ( .CLK(n177), .D(N188), .Q(\ram[8][171] ) );
  LATCHX1_HVT \ram_reg[8][170]  ( .CLK(n177), .D(N187), .Q(\ram[8][170] ) );
  LATCHX1_HVT \ram_reg[8][169]  ( .CLK(n177), .D(N186), .Q(\ram[8][169] ) );
  LATCHX1_HVT \ram_reg[8][168]  ( .CLK(n177), .D(N185), .Q(\ram[8][168] ) );
  LATCHX1_HVT \ram_reg[8][167]  ( .CLK(n177), .D(N184), .Q(\ram[8][167] ) );
  LATCHX1_HVT \ram_reg[8][166]  ( .CLK(n177), .D(N183), .Q(\ram[8][166] ) );
  LATCHX1_HVT \ram_reg[8][165]  ( .CLK(n177), .D(N182), .Q(\ram[8][165] ) );
  LATCHX1_HVT \ram_reg[8][164]  ( .CLK(n177), .D(N181), .Q(\ram[8][164] ) );
  LATCHX1_HVT \ram_reg[8][163]  ( .CLK(n176), .D(N180), .Q(\ram[8][163] ) );
  LATCHX1_HVT \ram_reg[8][162]  ( .CLK(n176), .D(N179), .Q(\ram[8][162] ) );
  LATCHX1_HVT \ram_reg[8][161]  ( .CLK(n176), .D(N178), .Q(\ram[8][161] ) );
  LATCHX1_HVT \ram_reg[8][160]  ( .CLK(n176), .D(N177), .Q(\ram[8][160] ) );
  LATCHX1_HVT \ram_reg[8][159]  ( .CLK(n176), .D(N176), .Q(\ram[8][159] ) );
  LATCHX1_HVT \ram_reg[8][158]  ( .CLK(n176), .D(N175), .Q(\ram[8][158] ) );
  LATCHX1_HVT \ram_reg[8][157]  ( .CLK(n176), .D(N174), .Q(\ram[8][157] ) );
  LATCHX1_HVT \ram_reg[8][156]  ( .CLK(n176), .D(N173), .Q(\ram[8][156] ) );
  LATCHX1_HVT \ram_reg[8][155]  ( .CLK(n176), .D(N172), .Q(\ram[8][155] ) );
  LATCHX1_HVT \ram_reg[8][154]  ( .CLK(n176), .D(N171), .Q(\ram[8][154] ) );
  LATCHX1_HVT \ram_reg[8][153]  ( .CLK(n176), .D(N170), .Q(\ram[8][153] ) );
  LATCHX1_HVT \ram_reg[8][152]  ( .CLK(n175), .D(N169), .Q(\ram[8][152] ) );
  LATCHX1_HVT \ram_reg[8][151]  ( .CLK(n175), .D(N168), .Q(\ram[8][151] ) );
  LATCHX1_HVT \ram_reg[8][150]  ( .CLK(n175), .D(N167), .Q(\ram[8][150] ) );
  LATCHX1_HVT \ram_reg[8][149]  ( .CLK(n175), .D(N166), .Q(\ram[8][149] ) );
  LATCHX1_HVT \ram_reg[8][148]  ( .CLK(n175), .D(N165), .Q(\ram[8][148] ) );
  LATCHX1_HVT \ram_reg[8][147]  ( .CLK(n175), .D(N164), .Q(\ram[8][147] ) );
  LATCHX1_HVT \ram_reg[8][146]  ( .CLK(n175), .D(N163), .Q(\ram[8][146] ) );
  LATCHX1_HVT \ram_reg[8][145]  ( .CLK(n175), .D(N162), .Q(\ram[8][145] ) );
  LATCHX1_HVT \ram_reg[8][144]  ( .CLK(n175), .D(N161), .Q(\ram[8][144] ) );
  LATCHX1_HVT \ram_reg[8][143]  ( .CLK(n175), .D(N160), .Q(\ram[8][143] ) );
  LATCHX1_HVT \ram_reg[8][142]  ( .CLK(n175), .D(N159), .Q(\ram[8][142] ) );
  LATCHX1_HVT \ram_reg[8][141]  ( .CLK(n174), .D(N158), .Q(\ram[8][141] ) );
  LATCHX1_HVT \ram_reg[8][140]  ( .CLK(n174), .D(N157), .Q(\ram[8][140] ) );
  LATCHX1_HVT \ram_reg[8][139]  ( .CLK(n174), .D(N156), .Q(\ram[8][139] ) );
  LATCHX1_HVT \ram_reg[8][138]  ( .CLK(n173), .D(N155), .Q(\ram[8][138] ) );
  LATCHX1_HVT \ram_reg[8][137]  ( .CLK(n182), .D(N154), .Q(\ram[8][137] ) );
  LATCHX1_HVT \ram_reg[8][136]  ( .CLK(n181), .D(N153), .Q(\ram[8][136] ) );
  LATCHX1_HVT \ram_reg[8][135]  ( .CLK(n181), .D(N152), .Q(\ram[8][135] ) );
  LATCHX1_HVT \ram_reg[8][134]  ( .CLK(n180), .D(N151), .Q(\ram[8][134] ) );
  LATCHX1_HVT \ram_reg[8][133]  ( .CLK(n179), .D(N150), .Q(\ram[8][133] ) );
  LATCHX1_HVT \ram_reg[8][132]  ( .CLK(n178), .D(N149), .Q(\ram[8][132] ) );
  LATCHX1_HVT \ram_reg[8][131]  ( .CLK(n177), .D(N148), .Q(\ram[8][131] ) );
  LATCHX1_HVT \ram_reg[8][130]  ( .CLK(n176), .D(N147), .Q(\ram[8][130] ) );
  LATCHX1_HVT \ram_reg[8][129]  ( .CLK(n175), .D(N146), .Q(\ram[8][129] ) );
  LATCHX1_HVT \ram_reg[8][128]  ( .CLK(n172), .D(N145), .Q(\ram[8][128] ) );
  LATCHX1_HVT \ram_reg[8][127]  ( .CLK(n163), .D(N144), .Q(\ram[8][127] ) );
  LATCHX1_HVT \ram_reg[8][126]  ( .CLK(n163), .D(N143), .Q(\ram[8][126] ) );
  LATCHX1_HVT \ram_reg[8][125]  ( .CLK(n163), .D(N142), .Q(\ram[8][125] ) );
  LATCHX1_HVT \ram_reg[8][124]  ( .CLK(n163), .D(N141), .Q(\ram[8][124] ) );
  LATCHX1_HVT \ram_reg[8][123]  ( .CLK(n163), .D(N140), .Q(\ram[8][123] ) );
  LATCHX1_HVT \ram_reg[8][122]  ( .CLK(n162), .D(N139), .Q(\ram[8][122] ) );
  LATCHX1_HVT \ram_reg[8][121]  ( .CLK(n163), .D(N138), .Q(\ram[8][121] ) );
  LATCHX1_HVT \ram_reg[8][120]  ( .CLK(n163), .D(N137), .Q(\ram[8][120] ) );
  LATCHX1_HVT \ram_reg[8][119]  ( .CLK(n172), .D(N136), .Q(\ram[8][119] ) );
  LATCHX1_HVT \ram_reg[8][118]  ( .CLK(n171), .D(N135), .Q(\ram[8][118] ) );
  LATCHX1_HVT \ram_reg[8][117]  ( .CLK(n171), .D(N134), .Q(\ram[8][117] ) );
  LATCHX1_HVT \ram_reg[8][116]  ( .CLK(n170), .D(N133), .Q(\ram[8][116] ) );
  LATCHX1_HVT \ram_reg[8][115]  ( .CLK(n165), .D(N132), .Q(\ram[8][115] ) );
  LATCHX1_HVT \ram_reg[8][114]  ( .CLK(n170), .D(N131), .Q(\ram[8][114] ) );
  LATCHX1_HVT \ram_reg[8][113]  ( .CLK(n170), .D(N130), .Q(\ram[8][113] ) );
  LATCHX1_HVT \ram_reg[8][112]  ( .CLK(n171), .D(N129), .Q(\ram[8][112] ) );
  LATCHX1_HVT \ram_reg[8][111]  ( .CLK(n169), .D(N128), .Q(\ram[8][111] ) );
  LATCHX1_HVT \ram_reg[8][110]  ( .CLK(n169), .D(N127), .Q(\ram[8][110] ) );
  LATCHX1_HVT \ram_reg[8][109]  ( .CLK(n169), .D(N126), .Q(\ram[8][109] ) );
  LATCHX1_HVT \ram_reg[8][108]  ( .CLK(n166), .D(N125), .Q(\ram[8][108] ) );
  LATCHX1_HVT \ram_reg[8][107]  ( .CLK(n163), .D(N124), .Q(\ram[8][107] ) );
  LATCHX1_HVT \ram_reg[8][106]  ( .CLK(n169), .D(N123), .Q(\ram[8][106] ) );
  LATCHX1_HVT \ram_reg[8][105]  ( .CLK(n169), .D(N122), .Q(\ram[8][105] ) );
  LATCHX1_HVT \ram_reg[8][104]  ( .CLK(n169), .D(N121), .Q(\ram[8][104] ) );
  LATCHX1_HVT \ram_reg[8][103]  ( .CLK(n168), .D(N120), .Q(\ram[8][103] ) );
  LATCHX1_HVT \ram_reg[8][102]  ( .CLK(n167), .D(N119), .Q(\ram[8][102] ) );
  LATCHX1_HVT \ram_reg[8][101]  ( .CLK(n167), .D(N118), .Q(\ram[8][101] ) );
  LATCHX1_HVT \ram_reg[8][100]  ( .CLK(n168), .D(N117), .Q(\ram[8][100] ) );
  LATCHX1_HVT \ram_reg[8][99]  ( .CLK(n166), .D(N116), .Q(\ram[8][99] ) );
  LATCHX1_HVT \ram_reg[8][98]  ( .CLK(n167), .D(N114), .Q(\ram[8][98] ) );
  LATCHX1_HVT \ram_reg[8][97]  ( .CLK(n168), .D(N113), .Q(\ram[8][97] ) );
  LATCHX1_HVT \ram_reg[8][96]  ( .CLK(n172), .D(N112), .Q(\ram[8][96] ) );
  LATCHX1_HVT \ram_reg[8][95]  ( .CLK(n164), .D(N111), .Q(\ram[8][95] ) );
  LATCHX1_HVT \ram_reg[8][94]  ( .CLK(n164), .D(N110), .Q(\ram[8][94] ) );
  LATCHX1_HVT \ram_reg[8][93]  ( .CLK(n164), .D(N109), .Q(\ram[8][93] ) );
  LATCHX1_HVT \ram_reg[8][92]  ( .CLK(n163), .D(N108), .Q(\ram[8][92] ) );
  LATCHX1_HVT \ram_reg[8][91]  ( .CLK(n163), .D(N107), .Q(\ram[8][91] ) );
  LATCHX1_HVT \ram_reg[8][90]  ( .CLK(n164), .D(N106), .Q(\ram[8][90] ) );
  LATCHX1_HVT \ram_reg[8][89]  ( .CLK(n163), .D(N105), .Q(\ram[8][89] ) );
  LATCHX1_HVT \ram_reg[8][88]  ( .CLK(n164), .D(N104), .Q(\ram[8][88] ) );
  LATCHX1_HVT \ram_reg[8][87]  ( .CLK(n172), .D(N103), .Q(\ram[8][87] ) );
  LATCHX1_HVT \ram_reg[8][86]  ( .CLK(n171), .D(N102), .Q(\ram[8][86] ) );
  LATCHX1_HVT \ram_reg[8][85]  ( .CLK(n170), .D(N101), .Q(\ram[8][85] ) );
  LATCHX1_HVT \ram_reg[8][84]  ( .CLK(n170), .D(N100), .Q(\ram[8][84] ) );
  LATCHX1_HVT \ram_reg[8][83]  ( .CLK(n165), .D(N99), .Q(\ram[8][83] ) );
  LATCHX1_HVT \ram_reg[8][82]  ( .CLK(n171), .D(N98), .Q(\ram[8][82] ) );
  LATCHX1_HVT \ram_reg[8][81]  ( .CLK(n170), .D(N97), .Q(\ram[8][81] ) );
  LATCHX1_HVT \ram_reg[8][80]  ( .CLK(n171), .D(N96), .Q(\ram[8][80] ) );
  LATCHX1_HVT \ram_reg[8][79]  ( .CLK(n165), .D(N95), .Q(\ram[8][79] ) );
  LATCHX1_HVT \ram_reg[8][78]  ( .CLK(n164), .D(N94), .Q(\ram[8][78] ) );
  LATCHX1_HVT \ram_reg[8][77]  ( .CLK(n165), .D(N93), .Q(\ram[8][77] ) );
  LATCHX1_HVT \ram_reg[8][76]  ( .CLK(n164), .D(N92), .Q(\ram[8][76] ) );
  LATCHX1_HVT \ram_reg[8][75]  ( .CLK(n164), .D(N91), .Q(\ram[8][75] ) );
  LATCHX1_HVT \ram_reg[8][74]  ( .CLK(n162), .D(N90), .Q(\ram[8][74] ) );
  LATCHX1_HVT \ram_reg[8][73]  ( .CLK(n165), .D(N89), .Q(\ram[8][73] ) );
  LATCHX1_HVT \ram_reg[8][72]  ( .CLK(n165), .D(N88), .Q(\ram[8][72] ) );
  LATCHX1_HVT \ram_reg[8][71]  ( .CLK(n168), .D(N87), .Q(\ram[8][71] ) );
  LATCHX1_HVT \ram_reg[8][70]  ( .CLK(n168), .D(N86), .Q(\ram[8][70] ) );
  LATCHX1_HVT \ram_reg[8][69]  ( .CLK(n167), .D(N85), .Q(\ram[8][69] ) );
  LATCHX1_HVT \ram_reg[8][68]  ( .CLK(n168), .D(N84), .Q(\ram[8][68] ) );
  LATCHX1_HVT \ram_reg[8][67]  ( .CLK(n167), .D(N83), .Q(\ram[8][67] ) );
  LATCHX1_HVT \ram_reg[8][66]  ( .CLK(n166), .D(N82), .Q(\ram[8][66] ) );
  LATCHX1_HVT \ram_reg[8][65]  ( .CLK(n167), .D(N81), .Q(\ram[8][65] ) );
  LATCHX1_HVT \ram_reg[8][64]  ( .CLK(n172), .D(N80), .Q(\ram[8][64] ) );
  LATCHX1_HVT \ram_reg[8][63]  ( .CLK(n166), .D(N79), .Q(\ram[8][63] ) );
  LATCHX1_HVT \ram_reg[8][62]  ( .CLK(n166), .D(N78), .Q(\ram[8][62] ) );
  LATCHX1_HVT \ram_reg[8][61]  ( .CLK(n166), .D(N77), .Q(\ram[8][61] ) );
  LATCHX1_HVT \ram_reg[8][60]  ( .CLK(n166), .D(N76), .Q(\ram[8][60] ) );
  LATCHX1_HVT \ram_reg[8][59]  ( .CLK(n166), .D(N75), .Q(\ram[8][59] ) );
  LATCHX1_HVT \ram_reg[8][58]  ( .CLK(n165), .D(N74), .Q(\ram[8][58] ) );
  LATCHX1_HVT \ram_reg[8][57]  ( .CLK(n166), .D(N73), .Q(\ram[8][57] ) );
  LATCHX1_HVT \ram_reg[8][56]  ( .CLK(n166), .D(N72), .Q(\ram[8][56] ) );
  LATCHX1_HVT \ram_reg[8][55]  ( .CLK(n172), .D(N71), .Q(\ram[8][55] ) );
  LATCHX1_HVT \ram_reg[8][54]  ( .CLK(n170), .D(N70), .Q(\ram[8][54] ) );
  LATCHX1_HVT \ram_reg[8][53]  ( .CLK(n170), .D(N69), .Q(\ram[8][53] ) );
  LATCHX1_HVT \ram_reg[8][52]  ( .CLK(n171), .D(N68), .Q(\ram[8][52] ) );
  LATCHX1_HVT \ram_reg[8][51]  ( .CLK(n165), .D(N67), .Q(\ram[8][51] ) );
  LATCHX1_HVT \ram_reg[8][50]  ( .CLK(n162), .D(N66), .Q(\ram[8][50] ) );
  LATCHX1_HVT \ram_reg[8][49]  ( .CLK(n171), .D(N65), .Q(\ram[8][49] ) );
  LATCHX1_HVT \ram_reg[8][48]  ( .CLK(n171), .D(N64), .Q(\ram[8][48] ) );
  LATCHX1_HVT \ram_reg[8][47]  ( .CLK(n169), .D(N63), .Q(\ram[8][47] ) );
  LATCHX1_HVT \ram_reg[8][46]  ( .CLK(n169), .D(N62), .Q(\ram[8][46] ) );
  LATCHX1_HVT \ram_reg[8][45]  ( .CLK(n169), .D(N61), .Q(\ram[8][45] ) );
  LATCHX1_HVT \ram_reg[8][44]  ( .CLK(n169), .D(N60), .Q(\ram[8][44] ) );
  LATCHX1_HVT \ram_reg[8][43]  ( .CLK(n166), .D(N59), .Q(\ram[8][43] ) );
  LATCHX1_HVT \ram_reg[8][42]  ( .CLK(n170), .D(N58), .Q(\ram[8][42] ) );
  LATCHX1_HVT \ram_reg[8][41]  ( .CLK(n163), .D(N57), .Q(\ram[8][41] ) );
  LATCHX1_HVT \ram_reg[8][40]  ( .CLK(n169), .D(N56), .Q(\ram[8][40] ) );
  LATCHX1_HVT \ram_reg[8][39]  ( .CLK(n168), .D(N55), .Q(\ram[8][39] ) );
  LATCHX1_HVT \ram_reg[8][38]  ( .CLK(n168), .D(N54), .Q(\ram[8][38] ) );
  LATCHX1_HVT \ram_reg[8][37]  ( .CLK(n167), .D(N53), .Q(\ram[8][37] ) );
  LATCHX1_HVT \ram_reg[8][36]  ( .CLK(n167), .D(N52), .Q(\ram[8][36] ) );
  LATCHX1_HVT \ram_reg[8][35]  ( .CLK(n167), .D(N51), .Q(\ram[8][35] ) );
  LATCHX1_HVT \ram_reg[8][34]  ( .CLK(n169), .D(N50), .Q(\ram[8][34] ) );
  LATCHX1_HVT \ram_reg[8][33]  ( .CLK(n168), .D(N49), .Q(\ram[8][33] ) );
  LATCHX1_HVT \ram_reg[8][32]  ( .CLK(n172), .D(N48), .Q(\ram[8][32] ) );
  LATCHX1_HVT \ram_reg[8][31]  ( .CLK(n162), .D(N47), .Q(\ram[8][31] ) );
  LATCHX1_HVT \ram_reg[8][30]  ( .CLK(n162), .D(N46), .Q(\ram[8][30] ) );
  LATCHX1_HVT \ram_reg[8][29]  ( .CLK(n162), .D(N45), .Q(\ram[8][29] ) );
  LATCHX1_HVT \ram_reg[8][28]  ( .CLK(n162), .D(N44), .Q(\ram[8][28] ) );
  LATCHX1_HVT \ram_reg[8][27]  ( .CLK(n162), .D(N43), .Q(\ram[8][27] ) );
  LATCHX1_HVT \ram_reg[8][26]  ( .CLK(n162), .D(N42), .Q(\ram[8][26] ) );
  LATCHX1_HVT \ram_reg[8][25]  ( .CLK(n162), .D(N41), .Q(\ram[8][25] ) );
  LATCHX1_HVT \ram_reg[8][24]  ( .CLK(n162), .D(N40), .Q(\ram[8][24] ) );
  LATCHX1_HVT \ram_reg[8][23]  ( .CLK(n172), .D(N39), .Q(\ram[8][23] ) );
  LATCHX1_HVT \ram_reg[8][22]  ( .CLK(n171), .D(N38), .Q(\ram[8][22] ) );
  LATCHX1_HVT \ram_reg[8][21]  ( .CLK(n170), .D(N37), .Q(\ram[8][21] ) );
  LATCHX1_HVT \ram_reg[8][20]  ( .CLK(n170), .D(N36), .Q(\ram[8][20] ) );
  LATCHX1_HVT \ram_reg[8][19]  ( .CLK(n162), .D(N35), .Q(\ram[8][19] ) );
  LATCHX1_HVT \ram_reg[8][18]  ( .CLK(n170), .D(N34), .Q(\ram[8][18] ) );
  LATCHX1_HVT \ram_reg[8][17]  ( .CLK(n171), .D(N33), .Q(\ram[8][17] ) );
  LATCHX1_HVT \ram_reg[8][16]  ( .CLK(n171), .D(N32), .Q(\ram[8][16] ) );
  LATCHX1_HVT \ram_reg[8][15]  ( .CLK(n165), .D(N31), .Q(\ram[8][15] ) );
  LATCHX1_HVT \ram_reg[8][14]  ( .CLK(n165), .D(N30), .Q(\ram[8][14] ) );
  LATCHX1_HVT \ram_reg[8][13]  ( .CLK(n164), .D(N29), .Q(\ram[8][13] ) );
  LATCHX1_HVT \ram_reg[8][12]  ( .CLK(n164), .D(N28), .Q(\ram[8][12] ) );
  LATCHX1_HVT \ram_reg[8][11]  ( .CLK(n165), .D(N27), .Q(\ram[8][11] ) );
  LATCHX1_HVT \ram_reg[8][10]  ( .CLK(n164), .D(N26), .Q(\ram[8][10] ) );
  LATCHX1_HVT \ram_reg[8][9]  ( .CLK(n164), .D(N25), .Q(\ram[8][9] ) );
  LATCHX1_HVT \ram_reg[8][8]  ( .CLK(n165), .D(N24), .Q(\ram[8][8] ) );
  LATCHX1_HVT \ram_reg[8][7]  ( .CLK(n168), .D(N23), .Q(\ram[8][7] ) );
  LATCHX1_HVT \ram_reg[8][6]  ( .CLK(n168), .D(N22), .Q(\ram[8][6] ) );
  LATCHX1_HVT \ram_reg[8][5]  ( .CLK(n167), .D(N21), .Q(\ram[8][5] ) );
  LATCHX1_HVT \ram_reg[8][4]  ( .CLK(n167), .D(N20), .Q(\ram[8][4] ) );
  LATCHX1_HVT \ram_reg[8][3]  ( .CLK(n166), .D(N19), .Q(\ram[8][3] ) );
  LATCHX1_HVT \ram_reg[8][2]  ( .CLK(n167), .D(N18), .Q(\ram[8][2] ) );
  LATCHX1_HVT \ram_reg[8][1]  ( .CLK(n168), .D(N17), .Q(\ram[8][1] ) );
  LATCHX1_HVT \ram_reg[8][0]  ( .CLK(n172), .D(N16), .Q(\ram[8][0] ) );
  LATCHX1_HVT \ram_reg[7][255]  ( .CLK(n185), .D(N273), .Q(\ram[7][255] ) );
  LATCHX1_HVT \ram_reg[7][254]  ( .CLK(n185), .D(N272), .Q(\ram[7][254] ) );
  LATCHX1_HVT \ram_reg[7][253]  ( .CLK(n185), .D(N271), .Q(\ram[7][253] ) );
  LATCHX1_HVT \ram_reg[7][252]  ( .CLK(N294), .D(N270), .Q(\ram[7][252] ) );
  LATCHX1_HVT \ram_reg[7][251]  ( .CLK(N294), .D(N269), .Q(\ram[7][251] ) );
  LATCHX1_HVT \ram_reg[7][250]  ( .CLK(n198), .D(N268), .Q(\ram[7][250] ) );
  LATCHX1_HVT \ram_reg[7][249]  ( .CLK(n197), .D(N267), .Q(\ram[7][249] ) );
  LATCHX1_HVT \ram_reg[7][248]  ( .CLK(n197), .D(N266), .Q(\ram[7][248] ) );
  LATCHX1_HVT \ram_reg[7][247]  ( .CLK(n197), .D(N265), .Q(\ram[7][247] ) );
  LATCHX1_HVT \ram_reg[7][246]  ( .CLK(n197), .D(N264), .Q(\ram[7][246] ) );
  LATCHX1_HVT \ram_reg[7][245]  ( .CLK(n197), .D(N263), .Q(\ram[7][245] ) );
  LATCHX1_HVT \ram_reg[7][244]  ( .CLK(n197), .D(N262), .Q(\ram[7][244] ) );
  LATCHX1_HVT \ram_reg[7][243]  ( .CLK(n197), .D(N261), .Q(\ram[7][243] ) );
  LATCHX1_HVT \ram_reg[7][242]  ( .CLK(n197), .D(N260), .Q(\ram[7][242] ) );
  LATCHX1_HVT \ram_reg[7][241]  ( .CLK(n197), .D(N259), .Q(\ram[7][241] ) );
  LATCHX1_HVT \ram_reg[7][240]  ( .CLK(n197), .D(N258), .Q(\ram[7][240] ) );
  LATCHX1_HVT \ram_reg[7][239]  ( .CLK(n197), .D(N257), .Q(\ram[7][239] ) );
  LATCHX1_HVT \ram_reg[7][238]  ( .CLK(n196), .D(N256), .Q(\ram[7][238] ) );
  LATCHX1_HVT \ram_reg[7][237]  ( .CLK(n196), .D(N255), .Q(\ram[7][237] ) );
  LATCHX1_HVT \ram_reg[7][236]  ( .CLK(n196), .D(N254), .Q(\ram[7][236] ) );
  LATCHX1_HVT \ram_reg[7][235]  ( .CLK(n196), .D(N253), .Q(\ram[7][235] ) );
  LATCHX1_HVT \ram_reg[7][234]  ( .CLK(n196), .D(N252), .Q(\ram[7][234] ) );
  LATCHX1_HVT \ram_reg[7][233]  ( .CLK(n196), .D(N251), .Q(\ram[7][233] ) );
  LATCHX1_HVT \ram_reg[7][232]  ( .CLK(n196), .D(N250), .Q(\ram[7][232] ) );
  LATCHX1_HVT \ram_reg[7][231]  ( .CLK(n196), .D(N249), .Q(\ram[7][231] ) );
  LATCHX1_HVT \ram_reg[7][230]  ( .CLK(n196), .D(N248), .Q(\ram[7][230] ) );
  LATCHX1_HVT \ram_reg[7][229]  ( .CLK(n196), .D(N247), .Q(\ram[7][229] ) );
  LATCHX1_HVT \ram_reg[7][228]  ( .CLK(n196), .D(N246), .Q(\ram[7][228] ) );
  LATCHX1_HVT \ram_reg[7][227]  ( .CLK(N294), .D(N245), .Q(\ram[7][227] ) );
  LATCHX1_HVT \ram_reg[7][226]  ( .CLK(n205), .D(N244), .Q(\ram[7][226] ) );
  LATCHX1_HVT \ram_reg[7][225]  ( .CLK(n205), .D(N243), .Q(\ram[7][225] ) );
  LATCHX1_HVT \ram_reg[7][224]  ( .CLK(n205), .D(N242), .Q(\ram[7][224] ) );
  LATCHX1_HVT \ram_reg[7][223]  ( .CLK(n205), .D(N241), .Q(\ram[7][223] ) );
  LATCHX1_HVT \ram_reg[7][222]  ( .CLK(n205), .D(N240), .Q(\ram[7][222] ) );
  LATCHX1_HVT \ram_reg[7][221]  ( .CLK(n205), .D(N239), .Q(\ram[7][221] ) );
  LATCHX1_HVT \ram_reg[7][220]  ( .CLK(n205), .D(N238), .Q(\ram[7][220] ) );
  LATCHX1_HVT \ram_reg[7][219]  ( .CLK(n205), .D(N237), .Q(\ram[7][219] ) );
  LATCHX1_HVT \ram_reg[7][218]  ( .CLK(n205), .D(N236), .Q(\ram[7][218] ) );
  LATCHX1_HVT \ram_reg[7][217]  ( .CLK(n205), .D(N235), .Q(\ram[7][217] ) );
  LATCHX1_HVT \ram_reg[7][216]  ( .CLK(n205), .D(N234), .Q(\ram[7][216] ) );
  LATCHX1_HVT \ram_reg[7][215]  ( .CLK(n204), .D(N233), .Q(\ram[7][215] ) );
  LATCHX1_HVT \ram_reg[7][214]  ( .CLK(n204), .D(N232), .Q(\ram[7][214] ) );
  LATCHX1_HVT \ram_reg[7][213]  ( .CLK(n204), .D(N231), .Q(\ram[7][213] ) );
  LATCHX1_HVT \ram_reg[7][212]  ( .CLK(n204), .D(N230), .Q(\ram[7][212] ) );
  LATCHX1_HVT \ram_reg[7][211]  ( .CLK(n204), .D(N229), .Q(\ram[7][211] ) );
  LATCHX1_HVT \ram_reg[7][210]  ( .CLK(n204), .D(N228), .Q(\ram[7][210] ) );
  LATCHX1_HVT \ram_reg[7][209]  ( .CLK(n204), .D(N227), .Q(\ram[7][209] ) );
  LATCHX1_HVT \ram_reg[7][208]  ( .CLK(n204), .D(N226), .Q(\ram[7][208] ) );
  LATCHX1_HVT \ram_reg[7][207]  ( .CLK(n204), .D(N225), .Q(\ram[7][207] ) );
  LATCHX1_HVT \ram_reg[7][206]  ( .CLK(n204), .D(N224), .Q(\ram[7][206] ) );
  LATCHX1_HVT \ram_reg[7][205]  ( .CLK(n204), .D(N223), .Q(\ram[7][205] ) );
  LATCHX1_HVT \ram_reg[7][204]  ( .CLK(n203), .D(N222), .Q(\ram[7][204] ) );
  LATCHX1_HVT \ram_reg[7][203]  ( .CLK(n203), .D(N221), .Q(\ram[7][203] ) );
  LATCHX1_HVT \ram_reg[7][202]  ( .CLK(n203), .D(N220), .Q(\ram[7][202] ) );
  LATCHX1_HVT \ram_reg[7][201]  ( .CLK(n203), .D(N219), .Q(\ram[7][201] ) );
  LATCHX1_HVT \ram_reg[7][200]  ( .CLK(n203), .D(N218), .Q(\ram[7][200] ) );
  LATCHX1_HVT \ram_reg[7][199]  ( .CLK(n203), .D(N217), .Q(\ram[7][199] ) );
  LATCHX1_HVT \ram_reg[7][198]  ( .CLK(n203), .D(N216), .Q(\ram[7][198] ) );
  LATCHX1_HVT \ram_reg[7][197]  ( .CLK(n203), .D(N214), .Q(\ram[7][197] ) );
  LATCHX1_HVT \ram_reg[7][196]  ( .CLK(n203), .D(N213), .Q(\ram[7][196] ) );
  LATCHX1_HVT \ram_reg[7][195]  ( .CLK(n203), .D(N212), .Q(\ram[7][195] ) );
  LATCHX1_HVT \ram_reg[7][194]  ( .CLK(n203), .D(N211), .Q(\ram[7][194] ) );
  LATCHX1_HVT \ram_reg[7][193]  ( .CLK(n202), .D(N210), .Q(\ram[7][193] ) );
  LATCHX1_HVT \ram_reg[7][192]  ( .CLK(n202), .D(N209), .Q(\ram[7][192] ) );
  LATCHX1_HVT \ram_reg[7][191]  ( .CLK(n202), .D(N208), .Q(\ram[7][191] ) );
  LATCHX1_HVT \ram_reg[7][190]  ( .CLK(n202), .D(N207), .Q(\ram[7][190] ) );
  LATCHX1_HVT \ram_reg[7][189]  ( .CLK(n202), .D(N206), .Q(\ram[7][189] ) );
  LATCHX1_HVT \ram_reg[7][188]  ( .CLK(n202), .D(N205), .Q(\ram[7][188] ) );
  LATCHX1_HVT \ram_reg[7][187]  ( .CLK(n202), .D(N204), .Q(\ram[7][187] ) );
  LATCHX1_HVT \ram_reg[7][186]  ( .CLK(n202), .D(N203), .Q(\ram[7][186] ) );
  LATCHX1_HVT \ram_reg[7][185]  ( .CLK(n202), .D(N202), .Q(\ram[7][185] ) );
  LATCHX1_HVT \ram_reg[7][184]  ( .CLK(n202), .D(N201), .Q(\ram[7][184] ) );
  LATCHX1_HVT \ram_reg[7][183]  ( .CLK(n202), .D(N200), .Q(\ram[7][183] ) );
  LATCHX1_HVT \ram_reg[7][182]  ( .CLK(n201), .D(N199), .Q(\ram[7][182] ) );
  LATCHX1_HVT \ram_reg[7][181]  ( .CLK(n201), .D(N198), .Q(\ram[7][181] ) );
  LATCHX1_HVT \ram_reg[7][180]  ( .CLK(n201), .D(N197), .Q(\ram[7][180] ) );
  LATCHX1_HVT \ram_reg[7][179]  ( .CLK(n201), .D(N196), .Q(\ram[7][179] ) );
  LATCHX1_HVT \ram_reg[7][178]  ( .CLK(n201), .D(N195), .Q(\ram[7][178] ) );
  LATCHX1_HVT \ram_reg[7][177]  ( .CLK(n201), .D(N194), .Q(\ram[7][177] ) );
  LATCHX1_HVT \ram_reg[7][176]  ( .CLK(n201), .D(N193), .Q(\ram[7][176] ) );
  LATCHX1_HVT \ram_reg[7][175]  ( .CLK(n201), .D(N192), .Q(\ram[7][175] ) );
  LATCHX1_HVT \ram_reg[7][174]  ( .CLK(n201), .D(N191), .Q(\ram[7][174] ) );
  LATCHX1_HVT \ram_reg[7][173]  ( .CLK(n201), .D(N190), .Q(\ram[7][173] ) );
  LATCHX1_HVT \ram_reg[7][172]  ( .CLK(n201), .D(N189), .Q(\ram[7][172] ) );
  LATCHX1_HVT \ram_reg[7][171]  ( .CLK(n200), .D(N188), .Q(\ram[7][171] ) );
  LATCHX1_HVT \ram_reg[7][170]  ( .CLK(n200), .D(N187), .Q(\ram[7][170] ) );
  LATCHX1_HVT \ram_reg[7][169]  ( .CLK(n200), .D(N186), .Q(\ram[7][169] ) );
  LATCHX1_HVT \ram_reg[7][168]  ( .CLK(n200), .D(N185), .Q(\ram[7][168] ) );
  LATCHX1_HVT \ram_reg[7][167]  ( .CLK(n200), .D(N184), .Q(\ram[7][167] ) );
  LATCHX1_HVT \ram_reg[7][166]  ( .CLK(n200), .D(N183), .Q(\ram[7][166] ) );
  LATCHX1_HVT \ram_reg[7][165]  ( .CLK(n200), .D(N182), .Q(\ram[7][165] ) );
  LATCHX1_HVT \ram_reg[7][164]  ( .CLK(n200), .D(N181), .Q(\ram[7][164] ) );
  LATCHX1_HVT \ram_reg[7][163]  ( .CLK(n200), .D(N180), .Q(\ram[7][163] ) );
  LATCHX1_HVT \ram_reg[7][162]  ( .CLK(n200), .D(N179), .Q(\ram[7][162] ) );
  LATCHX1_HVT \ram_reg[7][161]  ( .CLK(n200), .D(N178), .Q(\ram[7][161] ) );
  LATCHX1_HVT \ram_reg[7][160]  ( .CLK(n199), .D(N177), .Q(\ram[7][160] ) );
  LATCHX1_HVT \ram_reg[7][159]  ( .CLK(n199), .D(N176), .Q(\ram[7][159] ) );
  LATCHX1_HVT \ram_reg[7][158]  ( .CLK(n199), .D(N175), .Q(\ram[7][158] ) );
  LATCHX1_HVT \ram_reg[7][157]  ( .CLK(n199), .D(N174), .Q(\ram[7][157] ) );
  LATCHX1_HVT \ram_reg[7][156]  ( .CLK(n199), .D(N173), .Q(\ram[7][156] ) );
  LATCHX1_HVT \ram_reg[7][155]  ( .CLK(n199), .D(N172), .Q(\ram[7][155] ) );
  LATCHX1_HVT \ram_reg[7][154]  ( .CLK(n199), .D(N171), .Q(\ram[7][154] ) );
  LATCHX1_HVT \ram_reg[7][153]  ( .CLK(n199), .D(N170), .Q(\ram[7][153] ) );
  LATCHX1_HVT \ram_reg[7][152]  ( .CLK(n199), .D(N169), .Q(\ram[7][152] ) );
  LATCHX1_HVT \ram_reg[7][151]  ( .CLK(n199), .D(N168), .Q(\ram[7][151] ) );
  LATCHX1_HVT \ram_reg[7][150]  ( .CLK(n199), .D(N167), .Q(\ram[7][150] ) );
  LATCHX1_HVT \ram_reg[7][149]  ( .CLK(n198), .D(N166), .Q(\ram[7][149] ) );
  LATCHX1_HVT \ram_reg[7][148]  ( .CLK(n198), .D(N165), .Q(\ram[7][148] ) );
  LATCHX1_HVT \ram_reg[7][147]  ( .CLK(n198), .D(N164), .Q(\ram[7][147] ) );
  LATCHX1_HVT \ram_reg[7][146]  ( .CLK(n198), .D(N163), .Q(\ram[7][146] ) );
  LATCHX1_HVT \ram_reg[7][145]  ( .CLK(n198), .D(N162), .Q(\ram[7][145] ) );
  LATCHX1_HVT \ram_reg[7][144]  ( .CLK(n198), .D(N161), .Q(\ram[7][144] ) );
  LATCHX1_HVT \ram_reg[7][143]  ( .CLK(n198), .D(N160), .Q(\ram[7][143] ) );
  LATCHX1_HVT \ram_reg[7][142]  ( .CLK(n198), .D(N159), .Q(\ram[7][142] ) );
  LATCHX1_HVT \ram_reg[7][141]  ( .CLK(n198), .D(N158), .Q(\ram[7][141] ) );
  LATCHX1_HVT \ram_reg[7][140]  ( .CLK(n198), .D(N157), .Q(\ram[7][140] ) );
  LATCHX1_HVT \ram_reg[7][139]  ( .CLK(n197), .D(N156), .Q(\ram[7][139] ) );
  LATCHX1_HVT \ram_reg[7][138]  ( .CLK(n196), .D(N155), .Q(\ram[7][138] ) );
  LATCHX1_HVT \ram_reg[7][137]  ( .CLK(N294), .D(N154), .Q(\ram[7][137] ) );
  LATCHX1_HVT \ram_reg[7][136]  ( .CLK(n205), .D(N153), .Q(\ram[7][136] ) );
  LATCHX1_HVT \ram_reg[7][135]  ( .CLK(n204), .D(N152), .Q(\ram[7][135] ) );
  LATCHX1_HVT \ram_reg[7][134]  ( .CLK(n203), .D(N151), .Q(\ram[7][134] ) );
  LATCHX1_HVT \ram_reg[7][133]  ( .CLK(n202), .D(N150), .Q(\ram[7][133] ) );
  LATCHX1_HVT \ram_reg[7][132]  ( .CLK(n201), .D(N149), .Q(\ram[7][132] ) );
  LATCHX1_HVT \ram_reg[7][131]  ( .CLK(n200), .D(N148), .Q(\ram[7][131] ) );
  LATCHX1_HVT \ram_reg[7][130]  ( .CLK(n199), .D(N147), .Q(\ram[7][130] ) );
  LATCHX1_HVT \ram_reg[7][129]  ( .CLK(n198), .D(N146), .Q(\ram[7][129] ) );
  LATCHX1_HVT \ram_reg[7][128]  ( .CLK(n195), .D(N145), .Q(\ram[7][128] ) );
  LATCHX1_HVT \ram_reg[7][127]  ( .CLK(n186), .D(N144), .Q(\ram[7][127] ) );
  LATCHX1_HVT \ram_reg[7][126]  ( .CLK(n186), .D(N143), .Q(\ram[7][126] ) );
  LATCHX1_HVT \ram_reg[7][125]  ( .CLK(n186), .D(N142), .Q(\ram[7][125] ) );
  LATCHX1_HVT \ram_reg[7][124]  ( .CLK(n186), .D(N141), .Q(\ram[7][124] ) );
  LATCHX1_HVT \ram_reg[7][123]  ( .CLK(n186), .D(N140), .Q(\ram[7][123] ) );
  LATCHX1_HVT \ram_reg[7][122]  ( .CLK(n186), .D(N139), .Q(\ram[7][122] ) );
  LATCHX1_HVT \ram_reg[7][121]  ( .CLK(n186), .D(N138), .Q(\ram[7][121] ) );
  LATCHX1_HVT \ram_reg[7][120]  ( .CLK(n186), .D(N137), .Q(\ram[7][120] ) );
  LATCHX1_HVT \ram_reg[7][119]  ( .CLK(n195), .D(N136), .Q(\ram[7][119] ) );
  LATCHX1_HVT \ram_reg[7][118]  ( .CLK(n194), .D(N135), .Q(\ram[7][118] ) );
  LATCHX1_HVT \ram_reg[7][117]  ( .CLK(n194), .D(N134), .Q(\ram[7][117] ) );
  LATCHX1_HVT \ram_reg[7][116]  ( .CLK(n193), .D(N133), .Q(\ram[7][116] ) );
  LATCHX1_HVT \ram_reg[7][115]  ( .CLK(n188), .D(N132), .Q(\ram[7][115] ) );
  LATCHX1_HVT \ram_reg[7][114]  ( .CLK(n194), .D(N131), .Q(\ram[7][114] ) );
  LATCHX1_HVT \ram_reg[7][113]  ( .CLK(n193), .D(N130), .Q(\ram[7][113] ) );
  LATCHX1_HVT \ram_reg[7][112]  ( .CLK(n195), .D(N129), .Q(\ram[7][112] ) );
  LATCHX1_HVT \ram_reg[7][111]  ( .CLK(n193), .D(N128), .Q(\ram[7][111] ) );
  LATCHX1_HVT \ram_reg[7][110]  ( .CLK(n193), .D(N127), .Q(\ram[7][110] ) );
  LATCHX1_HVT \ram_reg[7][109]  ( .CLK(n192), .D(N126), .Q(\ram[7][109] ) );
  LATCHX1_HVT \ram_reg[7][108]  ( .CLK(n189), .D(N125), .Q(\ram[7][108] ) );
  LATCHX1_HVT \ram_reg[7][107]  ( .CLK(n186), .D(N124), .Q(\ram[7][107] ) );
  LATCHX1_HVT \ram_reg[7][106]  ( .CLK(n192), .D(N123), .Q(\ram[7][106] ) );
  LATCHX1_HVT \ram_reg[7][105]  ( .CLK(n192), .D(N122), .Q(\ram[7][105] ) );
  LATCHX1_HVT \ram_reg[7][104]  ( .CLK(n192), .D(N121), .Q(\ram[7][104] ) );
  LATCHX1_HVT \ram_reg[7][103]  ( .CLK(n192), .D(N120), .Q(\ram[7][103] ) );
  LATCHX1_HVT \ram_reg[7][102]  ( .CLK(n191), .D(N119), .Q(\ram[7][102] ) );
  LATCHX1_HVT \ram_reg[7][101]  ( .CLK(n190), .D(N118), .Q(\ram[7][101] ) );
  LATCHX1_HVT \ram_reg[7][100]  ( .CLK(n191), .D(N117), .Q(\ram[7][100] ) );
  LATCHX1_HVT \ram_reg[7][99]  ( .CLK(n190), .D(N116), .Q(\ram[7][99] ) );
  LATCHX1_HVT \ram_reg[7][98]  ( .CLK(n190), .D(N114), .Q(\ram[7][98] ) );
  LATCHX1_HVT \ram_reg[7][97]  ( .CLK(n191), .D(N113), .Q(\ram[7][97] ) );
  LATCHX1_HVT \ram_reg[7][96]  ( .CLK(n195), .D(N112), .Q(\ram[7][96] ) );
  LATCHX1_HVT \ram_reg[7][95]  ( .CLK(n187), .D(N111), .Q(\ram[7][95] ) );
  LATCHX1_HVT \ram_reg[7][94]  ( .CLK(n187), .D(N110), .Q(\ram[7][94] ) );
  LATCHX1_HVT \ram_reg[7][93]  ( .CLK(n187), .D(N109), .Q(\ram[7][93] ) );
  LATCHX1_HVT \ram_reg[7][92]  ( .CLK(n187), .D(N108), .Q(\ram[7][92] ) );
  LATCHX1_HVT \ram_reg[7][91]  ( .CLK(n187), .D(N107), .Q(\ram[7][91] ) );
  LATCHX1_HVT \ram_reg[7][90]  ( .CLK(n187), .D(N106), .Q(\ram[7][90] ) );
  LATCHX1_HVT \ram_reg[7][89]  ( .CLK(n187), .D(N105), .Q(\ram[7][89] ) );
  LATCHX1_HVT \ram_reg[7][88]  ( .CLK(n187), .D(N104), .Q(\ram[7][88] ) );
  LATCHX1_HVT \ram_reg[7][87]  ( .CLK(n195), .D(N103), .Q(\ram[7][87] ) );
  LATCHX1_HVT \ram_reg[7][86]  ( .CLK(n195), .D(N102), .Q(\ram[7][86] ) );
  LATCHX1_HVT \ram_reg[7][85]  ( .CLK(n193), .D(N101), .Q(\ram[7][85] ) );
  LATCHX1_HVT \ram_reg[7][84]  ( .CLK(n194), .D(N100), .Q(\ram[7][84] ) );
  LATCHX1_HVT \ram_reg[7][83]  ( .CLK(n189), .D(N99), .Q(\ram[7][83] ) );
  LATCHX1_HVT \ram_reg[7][82]  ( .CLK(n194), .D(N98), .Q(\ram[7][82] ) );
  LATCHX1_HVT \ram_reg[7][81]  ( .CLK(n193), .D(N97), .Q(\ram[7][81] ) );
  LATCHX1_HVT \ram_reg[7][80]  ( .CLK(n194), .D(N96), .Q(\ram[7][80] ) );
  LATCHX1_HVT \ram_reg[7][79]  ( .CLK(n188), .D(N95), .Q(\ram[7][79] ) );
  LATCHX1_HVT \ram_reg[7][78]  ( .CLK(n188), .D(N94), .Q(\ram[7][78] ) );
  LATCHX1_HVT \ram_reg[7][77]  ( .CLK(n188), .D(N93), .Q(\ram[7][77] ) );
  LATCHX1_HVT \ram_reg[7][76]  ( .CLK(n187), .D(N92), .Q(\ram[7][76] ) );
  LATCHX1_HVT \ram_reg[7][75]  ( .CLK(n187), .D(N91), .Q(\ram[7][75] ) );
  LATCHX1_HVT \ram_reg[7][74]  ( .CLK(n186), .D(N90), .Q(\ram[7][74] ) );
  LATCHX1_HVT \ram_reg[7][73]  ( .CLK(n188), .D(N89), .Q(\ram[7][73] ) );
  LATCHX1_HVT \ram_reg[7][72]  ( .CLK(n188), .D(N88), .Q(\ram[7][72] ) );
  LATCHX1_HVT \ram_reg[7][71]  ( .CLK(n192), .D(N87), .Q(\ram[7][71] ) );
  LATCHX1_HVT \ram_reg[7][70]  ( .CLK(n191), .D(N86), .Q(\ram[7][70] ) );
  LATCHX1_HVT \ram_reg[7][69]  ( .CLK(n190), .D(N85), .Q(\ram[7][69] ) );
  LATCHX1_HVT \ram_reg[7][68]  ( .CLK(n191), .D(N84), .Q(\ram[7][68] ) );
  LATCHX1_HVT \ram_reg[7][67]  ( .CLK(n190), .D(N83), .Q(\ram[7][67] ) );
  LATCHX1_HVT \ram_reg[7][66]  ( .CLK(n190), .D(N82), .Q(\ram[7][66] ) );
  LATCHX1_HVT \ram_reg[7][65]  ( .CLK(n191), .D(N81), .Q(\ram[7][65] ) );
  LATCHX1_HVT \ram_reg[7][64]  ( .CLK(n195), .D(N80), .Q(\ram[7][64] ) );
  LATCHX1_HVT \ram_reg[7][63]  ( .CLK(n189), .D(N79), .Q(\ram[7][63] ) );
  LATCHX1_HVT \ram_reg[7][62]  ( .CLK(n189), .D(N78), .Q(\ram[7][62] ) );
  LATCHX1_HVT \ram_reg[7][61]  ( .CLK(n189), .D(N77), .Q(\ram[7][61] ) );
  LATCHX1_HVT \ram_reg[7][60]  ( .CLK(n189), .D(N76), .Q(\ram[7][60] ) );
  LATCHX1_HVT \ram_reg[7][59]  ( .CLK(n189), .D(N75), .Q(\ram[7][59] ) );
  LATCHX1_HVT \ram_reg[7][58]  ( .CLK(n189), .D(N74), .Q(\ram[7][58] ) );
  LATCHX1_HVT \ram_reg[7][57]  ( .CLK(n189), .D(N73), .Q(\ram[7][57] ) );
  LATCHX1_HVT \ram_reg[7][56]  ( .CLK(n189), .D(N72), .Q(\ram[7][56] ) );
  LATCHX1_HVT \ram_reg[7][55]  ( .CLK(n195), .D(N71), .Q(\ram[7][55] ) );
  LATCHX1_HVT \ram_reg[7][54]  ( .CLK(n193), .D(N70), .Q(\ram[7][54] ) );
  LATCHX1_HVT \ram_reg[7][53]  ( .CLK(n193), .D(N69), .Q(\ram[7][53] ) );
  LATCHX1_HVT \ram_reg[7][52]  ( .CLK(n194), .D(N68), .Q(\ram[7][52] ) );
  LATCHX1_HVT \ram_reg[7][51]  ( .CLK(n189), .D(N67), .Q(\ram[7][51] ) );
  LATCHX1_HVT \ram_reg[7][50]  ( .CLK(n185), .D(N66), .Q(\ram[7][50] ) );
  LATCHX1_HVT \ram_reg[7][49]  ( .CLK(n194), .D(N65), .Q(\ram[7][49] ) );
  LATCHX1_HVT \ram_reg[7][48]  ( .CLK(n194), .D(N64), .Q(\ram[7][48] ) );
  LATCHX1_HVT \ram_reg[7][47]  ( .CLK(n193), .D(N63), .Q(\ram[7][47] ) );
  LATCHX1_HVT \ram_reg[7][46]  ( .CLK(n192), .D(N62), .Q(\ram[7][46] ) );
  LATCHX1_HVT \ram_reg[7][45]  ( .CLK(n192), .D(N61), .Q(\ram[7][45] ) );
  LATCHX1_HVT \ram_reg[7][44]  ( .CLK(n192), .D(N60), .Q(\ram[7][44] ) );
  LATCHX1_HVT \ram_reg[7][43]  ( .CLK(n189), .D(N59), .Q(\ram[7][43] ) );
  LATCHX1_HVT \ram_reg[7][42]  ( .CLK(n193), .D(N58), .Q(\ram[7][42] ) );
  LATCHX1_HVT \ram_reg[7][41]  ( .CLK(n186), .D(N57), .Q(\ram[7][41] ) );
  LATCHX1_HVT \ram_reg[7][40]  ( .CLK(n192), .D(N56), .Q(\ram[7][40] ) );
  LATCHX1_HVT \ram_reg[7][39]  ( .CLK(n191), .D(N55), .Q(\ram[7][39] ) );
  LATCHX1_HVT \ram_reg[7][38]  ( .CLK(n191), .D(N54), .Q(\ram[7][38] ) );
  LATCHX1_HVT \ram_reg[7][37]  ( .CLK(n190), .D(N53), .Q(\ram[7][37] ) );
  LATCHX1_HVT \ram_reg[7][36]  ( .CLK(n190), .D(N52), .Q(\ram[7][36] ) );
  LATCHX1_HVT \ram_reg[7][35]  ( .CLK(n190), .D(N51), .Q(\ram[7][35] ) );
  LATCHX1_HVT \ram_reg[7][34]  ( .CLK(n192), .D(N50), .Q(\ram[7][34] ) );
  LATCHX1_HVT \ram_reg[7][33]  ( .CLK(n191), .D(N49), .Q(\ram[7][33] ) );
  LATCHX1_HVT \ram_reg[7][32]  ( .CLK(n195), .D(N48), .Q(\ram[7][32] ) );
  LATCHX1_HVT \ram_reg[7][31]  ( .CLK(n185), .D(N47), .Q(\ram[7][31] ) );
  LATCHX1_HVT \ram_reg[7][30]  ( .CLK(n185), .D(N46), .Q(\ram[7][30] ) );
  LATCHX1_HVT \ram_reg[7][29]  ( .CLK(n185), .D(N45), .Q(\ram[7][29] ) );
  LATCHX1_HVT \ram_reg[7][28]  ( .CLK(n185), .D(N44), .Q(\ram[7][28] ) );
  LATCHX1_HVT \ram_reg[7][27]  ( .CLK(n186), .D(N43), .Q(\ram[7][27] ) );
  LATCHX1_HVT \ram_reg[7][26]  ( .CLK(n185), .D(N42), .Q(\ram[7][26] ) );
  LATCHX1_HVT \ram_reg[7][25]  ( .CLK(n185), .D(N41), .Q(\ram[7][25] ) );
  LATCHX1_HVT \ram_reg[7][24]  ( .CLK(n185), .D(N40), .Q(\ram[7][24] ) );
  LATCHX1_HVT \ram_reg[7][23]  ( .CLK(n195), .D(N39), .Q(\ram[7][23] ) );
  LATCHX1_HVT \ram_reg[7][22]  ( .CLK(n194), .D(N38), .Q(\ram[7][22] ) );
  LATCHX1_HVT \ram_reg[7][21]  ( .CLK(n194), .D(N37), .Q(\ram[7][21] ) );
  LATCHX1_HVT \ram_reg[7][20]  ( .CLK(n193), .D(N36), .Q(\ram[7][20] ) );
  LATCHX1_HVT \ram_reg[7][19]  ( .CLK(n185), .D(N35), .Q(\ram[7][19] ) );
  LATCHX1_HVT \ram_reg[7][18]  ( .CLK(n193), .D(N34), .Q(\ram[7][18] ) );
  LATCHX1_HVT \ram_reg[7][17]  ( .CLK(n194), .D(N33), .Q(\ram[7][17] ) );
  LATCHX1_HVT \ram_reg[7][16]  ( .CLK(n195), .D(N32), .Q(\ram[7][16] ) );
  LATCHX1_HVT \ram_reg[7][15]  ( .CLK(n188), .D(N31), .Q(\ram[7][15] ) );
  LATCHX1_HVT \ram_reg[7][14]  ( .CLK(n188), .D(N30), .Q(\ram[7][14] ) );
  LATCHX1_HVT \ram_reg[7][13]  ( .CLK(n187), .D(N29), .Q(\ram[7][13] ) );
  LATCHX1_HVT \ram_reg[7][12]  ( .CLK(n188), .D(N28), .Q(\ram[7][12] ) );
  LATCHX1_HVT \ram_reg[7][11]  ( .CLK(n188), .D(N27), .Q(\ram[7][11] ) );
  LATCHX1_HVT \ram_reg[7][10]  ( .CLK(n187), .D(N26), .Q(\ram[7][10] ) );
  LATCHX1_HVT \ram_reg[7][9]  ( .CLK(n188), .D(N25), .Q(\ram[7][9] ) );
  LATCHX1_HVT \ram_reg[7][8]  ( .CLK(n188), .D(N24), .Q(\ram[7][8] ) );
  LATCHX1_HVT \ram_reg[7][7]  ( .CLK(n192), .D(N23), .Q(\ram[7][7] ) );
  LATCHX1_HVT \ram_reg[7][6]  ( .CLK(n191), .D(N22), .Q(\ram[7][6] ) );
  LATCHX1_HVT \ram_reg[7][5]  ( .CLK(n190), .D(N21), .Q(\ram[7][5] ) );
  LATCHX1_HVT \ram_reg[7][4]  ( .CLK(n191), .D(N20), .Q(\ram[7][4] ) );
  LATCHX1_HVT \ram_reg[7][3]  ( .CLK(n190), .D(N19), .Q(\ram[7][3] ) );
  LATCHX1_HVT \ram_reg[7][2]  ( .CLK(n190), .D(N18), .Q(\ram[7][2] ) );
  LATCHX1_HVT \ram_reg[7][1]  ( .CLK(n191), .D(N17), .Q(\ram[7][1] ) );
  LATCHX1_HVT \ram_reg[7][0]  ( .CLK(n195), .D(N16), .Q(\ram[7][0] ) );
  LATCHX1_HVT \ram_reg[6][255]  ( .CLK(N291), .D(N273), .Q(\ram[6][255] ) );
  LATCHX1_HVT \ram_reg[6][254]  ( .CLK(N291), .D(N272), .Q(\ram[6][254] ) );
  LATCHX1_HVT \ram_reg[6][253]  ( .CLK(N291), .D(N271), .Q(\ram[6][253] ) );
  LATCHX1_HVT \ram_reg[6][252]  ( .CLK(N291), .D(N270), .Q(\ram[6][252] ) );
  LATCHX1_HVT \ram_reg[6][251]  ( .CLK(n228), .D(N269), .Q(\ram[6][251] ) );
  LATCHX1_HVT \ram_reg[6][250]  ( .CLK(n220), .D(N268), .Q(\ram[6][250] ) );
  LATCHX1_HVT \ram_reg[6][249]  ( .CLK(n220), .D(N267), .Q(\ram[6][249] ) );
  LATCHX1_HVT \ram_reg[6][248]  ( .CLK(n220), .D(N266), .Q(\ram[6][248] ) );
  LATCHX1_HVT \ram_reg[6][247]  ( .CLK(n220), .D(N265), .Q(\ram[6][247] ) );
  LATCHX1_HVT \ram_reg[6][246]  ( .CLK(n220), .D(N264), .Q(\ram[6][246] ) );
  LATCHX1_HVT \ram_reg[6][245]  ( .CLK(n220), .D(N263), .Q(\ram[6][245] ) );
  LATCHX1_HVT \ram_reg[6][244]  ( .CLK(n220), .D(N262), .Q(\ram[6][244] ) );
  LATCHX1_HVT \ram_reg[6][243]  ( .CLK(n220), .D(N261), .Q(\ram[6][243] ) );
  LATCHX1_HVT \ram_reg[6][242]  ( .CLK(n220), .D(N260), .Q(\ram[6][242] ) );
  LATCHX1_HVT \ram_reg[6][241]  ( .CLK(n219), .D(N259), .Q(\ram[6][241] ) );
  LATCHX1_HVT \ram_reg[6][240]  ( .CLK(n219), .D(N258), .Q(\ram[6][240] ) );
  LATCHX1_HVT \ram_reg[6][239]  ( .CLK(n219), .D(N257), .Q(\ram[6][239] ) );
  LATCHX1_HVT \ram_reg[6][238]  ( .CLK(n219), .D(N256), .Q(\ram[6][238] ) );
  LATCHX1_HVT \ram_reg[6][237]  ( .CLK(n219), .D(N255), .Q(\ram[6][237] ) );
  LATCHX1_HVT \ram_reg[6][236]  ( .CLK(n219), .D(N254), .Q(\ram[6][236] ) );
  LATCHX1_HVT \ram_reg[6][235]  ( .CLK(n219), .D(N253), .Q(\ram[6][235] ) );
  LATCHX1_HVT \ram_reg[6][234]  ( .CLK(n219), .D(N252), .Q(\ram[6][234] ) );
  LATCHX1_HVT \ram_reg[6][233]  ( .CLK(n219), .D(N251), .Q(\ram[6][233] ) );
  LATCHX1_HVT \ram_reg[6][232]  ( .CLK(n219), .D(N250), .Q(\ram[6][232] ) );
  LATCHX1_HVT \ram_reg[6][231]  ( .CLK(n219), .D(N249), .Q(\ram[6][231] ) );
  LATCHX1_HVT \ram_reg[6][230]  ( .CLK(n218), .D(N248), .Q(\ram[6][230] ) );
  LATCHX1_HVT \ram_reg[6][229]  ( .CLK(n218), .D(N247), .Q(\ram[6][229] ) );
  LATCHX1_HVT \ram_reg[6][228]  ( .CLK(n218), .D(N246), .Q(\ram[6][228] ) );
  LATCHX1_HVT \ram_reg[6][227]  ( .CLK(n228), .D(N245), .Q(\ram[6][227] ) );
  LATCHX1_HVT \ram_reg[6][226]  ( .CLK(n228), .D(N244), .Q(\ram[6][226] ) );
  LATCHX1_HVT \ram_reg[6][225]  ( .CLK(n228), .D(N243), .Q(\ram[6][225] ) );
  LATCHX1_HVT \ram_reg[6][224]  ( .CLK(n228), .D(N242), .Q(\ram[6][224] ) );
  LATCHX1_HVT \ram_reg[6][223]  ( .CLK(n228), .D(N241), .Q(\ram[6][223] ) );
  LATCHX1_HVT \ram_reg[6][222]  ( .CLK(n228), .D(N240), .Q(\ram[6][222] ) );
  LATCHX1_HVT \ram_reg[6][221]  ( .CLK(n228), .D(N239), .Q(\ram[6][221] ) );
  LATCHX1_HVT \ram_reg[6][220]  ( .CLK(n228), .D(N238), .Q(\ram[6][220] ) );
  LATCHX1_HVT \ram_reg[6][219]  ( .CLK(n228), .D(N237), .Q(\ram[6][219] ) );
  LATCHX1_HVT \ram_reg[6][218]  ( .CLK(n228), .D(N236), .Q(\ram[6][218] ) );
  LATCHX1_HVT \ram_reg[6][217]  ( .CLK(n227), .D(N235), .Q(\ram[6][217] ) );
  LATCHX1_HVT \ram_reg[6][216]  ( .CLK(n227), .D(N234), .Q(\ram[6][216] ) );
  LATCHX1_HVT \ram_reg[6][215]  ( .CLK(n227), .D(N233), .Q(\ram[6][215] ) );
  LATCHX1_HVT \ram_reg[6][214]  ( .CLK(n227), .D(N232), .Q(\ram[6][214] ) );
  LATCHX1_HVT \ram_reg[6][213]  ( .CLK(n227), .D(N231), .Q(\ram[6][213] ) );
  LATCHX1_HVT \ram_reg[6][212]  ( .CLK(n227), .D(N230), .Q(\ram[6][212] ) );
  LATCHX1_HVT \ram_reg[6][211]  ( .CLK(n227), .D(N229), .Q(\ram[6][211] ) );
  LATCHX1_HVT \ram_reg[6][210]  ( .CLK(n227), .D(N228), .Q(\ram[6][210] ) );
  LATCHX1_HVT \ram_reg[6][209]  ( .CLK(n227), .D(N227), .Q(\ram[6][209] ) );
  LATCHX1_HVT \ram_reg[6][208]  ( .CLK(n227), .D(N226), .Q(\ram[6][208] ) );
  LATCHX1_HVT \ram_reg[6][207]  ( .CLK(n226), .D(N225), .Q(\ram[6][207] ) );
  LATCHX1_HVT \ram_reg[6][206]  ( .CLK(n226), .D(N224), .Q(\ram[6][206] ) );
  LATCHX1_HVT \ram_reg[6][205]  ( .CLK(n226), .D(N223), .Q(\ram[6][205] ) );
  LATCHX1_HVT \ram_reg[6][204]  ( .CLK(n226), .D(N222), .Q(\ram[6][204] ) );
  LATCHX1_HVT \ram_reg[6][203]  ( .CLK(n226), .D(N221), .Q(\ram[6][203] ) );
  LATCHX1_HVT \ram_reg[6][202]  ( .CLK(n226), .D(N220), .Q(\ram[6][202] ) );
  LATCHX1_HVT \ram_reg[6][201]  ( .CLK(n226), .D(N219), .Q(\ram[6][201] ) );
  LATCHX1_HVT \ram_reg[6][200]  ( .CLK(n226), .D(N218), .Q(\ram[6][200] ) );
  LATCHX1_HVT \ram_reg[6][199]  ( .CLK(n226), .D(N217), .Q(\ram[6][199] ) );
  LATCHX1_HVT \ram_reg[6][198]  ( .CLK(n226), .D(N216), .Q(\ram[6][198] ) );
  LATCHX1_HVT \ram_reg[6][197]  ( .CLK(n226), .D(N214), .Q(\ram[6][197] ) );
  LATCHX1_HVT \ram_reg[6][196]  ( .CLK(n225), .D(N213), .Q(\ram[6][196] ) );
  LATCHX1_HVT \ram_reg[6][195]  ( .CLK(n225), .D(N212), .Q(\ram[6][195] ) );
  LATCHX1_HVT \ram_reg[6][194]  ( .CLK(n225), .D(N211), .Q(\ram[6][194] ) );
  LATCHX1_HVT \ram_reg[6][193]  ( .CLK(n225), .D(N210), .Q(\ram[6][193] ) );
  LATCHX1_HVT \ram_reg[6][192]  ( .CLK(n225), .D(N209), .Q(\ram[6][192] ) );
  LATCHX1_HVT \ram_reg[6][191]  ( .CLK(n225), .D(N208), .Q(\ram[6][191] ) );
  LATCHX1_HVT \ram_reg[6][190]  ( .CLK(n225), .D(N207), .Q(\ram[6][190] ) );
  LATCHX1_HVT \ram_reg[6][189]  ( .CLK(n225), .D(N206), .Q(\ram[6][189] ) );
  LATCHX1_HVT \ram_reg[6][188]  ( .CLK(n225), .D(N205), .Q(\ram[6][188] ) );
  LATCHX1_HVT \ram_reg[6][187]  ( .CLK(n225), .D(N204), .Q(\ram[6][187] ) );
  LATCHX1_HVT \ram_reg[6][186]  ( .CLK(n225), .D(N203), .Q(\ram[6][186] ) );
  LATCHX1_HVT \ram_reg[6][185]  ( .CLK(n224), .D(N202), .Q(\ram[6][185] ) );
  LATCHX1_HVT \ram_reg[6][184]  ( .CLK(n224), .D(N201), .Q(\ram[6][184] ) );
  LATCHX1_HVT \ram_reg[6][183]  ( .CLK(n224), .D(N200), .Q(\ram[6][183] ) );
  LATCHX1_HVT \ram_reg[6][182]  ( .CLK(n224), .D(N199), .Q(\ram[6][182] ) );
  LATCHX1_HVT \ram_reg[6][181]  ( .CLK(n224), .D(N198), .Q(\ram[6][181] ) );
  LATCHX1_HVT \ram_reg[6][180]  ( .CLK(n224), .D(N197), .Q(\ram[6][180] ) );
  LATCHX1_HVT \ram_reg[6][179]  ( .CLK(n224), .D(N196), .Q(\ram[6][179] ) );
  LATCHX1_HVT \ram_reg[6][178]  ( .CLK(n224), .D(N195), .Q(\ram[6][178] ) );
  LATCHX1_HVT \ram_reg[6][177]  ( .CLK(n224), .D(N194), .Q(\ram[6][177] ) );
  LATCHX1_HVT \ram_reg[6][176]  ( .CLK(n224), .D(N193), .Q(\ram[6][176] ) );
  LATCHX1_HVT \ram_reg[6][175]  ( .CLK(n224), .D(N192), .Q(\ram[6][175] ) );
  LATCHX1_HVT \ram_reg[6][174]  ( .CLK(n223), .D(N191), .Q(\ram[6][174] ) );
  LATCHX1_HVT \ram_reg[6][173]  ( .CLK(n223), .D(N190), .Q(\ram[6][173] ) );
  LATCHX1_HVT \ram_reg[6][172]  ( .CLK(n223), .D(N189), .Q(\ram[6][172] ) );
  LATCHX1_HVT \ram_reg[6][171]  ( .CLK(n223), .D(N188), .Q(\ram[6][171] ) );
  LATCHX1_HVT \ram_reg[6][170]  ( .CLK(n223), .D(N187), .Q(\ram[6][170] ) );
  LATCHX1_HVT \ram_reg[6][169]  ( .CLK(n223), .D(N186), .Q(\ram[6][169] ) );
  LATCHX1_HVT \ram_reg[6][168]  ( .CLK(n223), .D(N185), .Q(\ram[6][168] ) );
  LATCHX1_HVT \ram_reg[6][167]  ( .CLK(n223), .D(N184), .Q(\ram[6][167] ) );
  LATCHX1_HVT \ram_reg[6][166]  ( .CLK(n223), .D(N183), .Q(\ram[6][166] ) );
  LATCHX1_HVT \ram_reg[6][165]  ( .CLK(n223), .D(N182), .Q(\ram[6][165] ) );
  LATCHX1_HVT \ram_reg[6][164]  ( .CLK(n223), .D(N181), .Q(\ram[6][164] ) );
  LATCHX1_HVT \ram_reg[6][163]  ( .CLK(n222), .D(N180), .Q(\ram[6][163] ) );
  LATCHX1_HVT \ram_reg[6][162]  ( .CLK(n222), .D(N179), .Q(\ram[6][162] ) );
  LATCHX1_HVT \ram_reg[6][161]  ( .CLK(n222), .D(N178), .Q(\ram[6][161] ) );
  LATCHX1_HVT \ram_reg[6][160]  ( .CLK(n222), .D(N177), .Q(\ram[6][160] ) );
  LATCHX1_HVT \ram_reg[6][159]  ( .CLK(n222), .D(N176), .Q(\ram[6][159] ) );
  LATCHX1_HVT \ram_reg[6][158]  ( .CLK(n222), .D(N175), .Q(\ram[6][158] ) );
  LATCHX1_HVT \ram_reg[6][157]  ( .CLK(n222), .D(N174), .Q(\ram[6][157] ) );
  LATCHX1_HVT \ram_reg[6][156]  ( .CLK(n222), .D(N173), .Q(\ram[6][156] ) );
  LATCHX1_HVT \ram_reg[6][155]  ( .CLK(n222), .D(N172), .Q(\ram[6][155] ) );
  LATCHX1_HVT \ram_reg[6][154]  ( .CLK(n222), .D(N171), .Q(\ram[6][154] ) );
  LATCHX1_HVT \ram_reg[6][153]  ( .CLK(n222), .D(N170), .Q(\ram[6][153] ) );
  LATCHX1_HVT \ram_reg[6][152]  ( .CLK(n221), .D(N169), .Q(\ram[6][152] ) );
  LATCHX1_HVT \ram_reg[6][151]  ( .CLK(n221), .D(N168), .Q(\ram[6][151] ) );
  LATCHX1_HVT \ram_reg[6][150]  ( .CLK(n221), .D(N167), .Q(\ram[6][150] ) );
  LATCHX1_HVT \ram_reg[6][149]  ( .CLK(n221), .D(N166), .Q(\ram[6][149] ) );
  LATCHX1_HVT \ram_reg[6][148]  ( .CLK(n221), .D(N165), .Q(\ram[6][148] ) );
  LATCHX1_HVT \ram_reg[6][147]  ( .CLK(n221), .D(N164), .Q(\ram[6][147] ) );
  LATCHX1_HVT \ram_reg[6][146]  ( .CLK(n221), .D(N163), .Q(\ram[6][146] ) );
  LATCHX1_HVT \ram_reg[6][145]  ( .CLK(n221), .D(N162), .Q(\ram[6][145] ) );
  LATCHX1_HVT \ram_reg[6][144]  ( .CLK(n221), .D(N161), .Q(\ram[6][144] ) );
  LATCHX1_HVT \ram_reg[6][143]  ( .CLK(n221), .D(N160), .Q(\ram[6][143] ) );
  LATCHX1_HVT \ram_reg[6][142]  ( .CLK(n221), .D(N159), .Q(\ram[6][142] ) );
  LATCHX1_HVT \ram_reg[6][141]  ( .CLK(n220), .D(N158), .Q(\ram[6][141] ) );
  LATCHX1_HVT \ram_reg[6][140]  ( .CLK(n220), .D(N157), .Q(\ram[6][140] ) );
  LATCHX1_HVT \ram_reg[6][139]  ( .CLK(n220), .D(N156), .Q(\ram[6][139] ) );
  LATCHX1_HVT \ram_reg[6][138]  ( .CLK(n219), .D(N155), .Q(\ram[6][138] ) );
  LATCHX1_HVT \ram_reg[6][137]  ( .CLK(n228), .D(N154), .Q(\ram[6][137] ) );
  LATCHX1_HVT \ram_reg[6][136]  ( .CLK(n227), .D(N153), .Q(\ram[6][136] ) );
  LATCHX1_HVT \ram_reg[6][135]  ( .CLK(n227), .D(N152), .Q(\ram[6][135] ) );
  LATCHX1_HVT \ram_reg[6][134]  ( .CLK(n226), .D(N151), .Q(\ram[6][134] ) );
  LATCHX1_HVT \ram_reg[6][133]  ( .CLK(n225), .D(N150), .Q(\ram[6][133] ) );
  LATCHX1_HVT \ram_reg[6][132]  ( .CLK(n224), .D(N149), .Q(\ram[6][132] ) );
  LATCHX1_HVT \ram_reg[6][131]  ( .CLK(n223), .D(N148), .Q(\ram[6][131] ) );
  LATCHX1_HVT \ram_reg[6][130]  ( .CLK(n222), .D(N147), .Q(\ram[6][130] ) );
  LATCHX1_HVT \ram_reg[6][129]  ( .CLK(n221), .D(N146), .Q(\ram[6][129] ) );
  LATCHX1_HVT \ram_reg[6][128]  ( .CLK(n218), .D(N145), .Q(\ram[6][128] ) );
  LATCHX1_HVT \ram_reg[6][127]  ( .CLK(n209), .D(N144), .Q(\ram[6][127] ) );
  LATCHX1_HVT \ram_reg[6][126]  ( .CLK(n209), .D(N143), .Q(\ram[6][126] ) );
  LATCHX1_HVT \ram_reg[6][125]  ( .CLK(n209), .D(N142), .Q(\ram[6][125] ) );
  LATCHX1_HVT \ram_reg[6][124]  ( .CLK(n209), .D(N141), .Q(\ram[6][124] ) );
  LATCHX1_HVT \ram_reg[6][123]  ( .CLK(n209), .D(N140), .Q(\ram[6][123] ) );
  LATCHX1_HVT \ram_reg[6][122]  ( .CLK(n208), .D(N139), .Q(\ram[6][122] ) );
  LATCHX1_HVT \ram_reg[6][121]  ( .CLK(n209), .D(N138), .Q(\ram[6][121] ) );
  LATCHX1_HVT \ram_reg[6][120]  ( .CLK(n209), .D(N137), .Q(\ram[6][120] ) );
  LATCHX1_HVT \ram_reg[6][119]  ( .CLK(n218), .D(N136), .Q(\ram[6][119] ) );
  LATCHX1_HVT \ram_reg[6][118]  ( .CLK(n217), .D(N135), .Q(\ram[6][118] ) );
  LATCHX1_HVT \ram_reg[6][117]  ( .CLK(n217), .D(N134), .Q(\ram[6][117] ) );
  LATCHX1_HVT \ram_reg[6][116]  ( .CLK(n216), .D(N133), .Q(\ram[6][116] ) );
  LATCHX1_HVT \ram_reg[6][115]  ( .CLK(n211), .D(N132), .Q(\ram[6][115] ) );
  LATCHX1_HVT \ram_reg[6][114]  ( .CLK(n216), .D(N131), .Q(\ram[6][114] ) );
  LATCHX1_HVT \ram_reg[6][113]  ( .CLK(n216), .D(N130), .Q(\ram[6][113] ) );
  LATCHX1_HVT \ram_reg[6][112]  ( .CLK(n217), .D(N129), .Q(\ram[6][112] ) );
  LATCHX1_HVT \ram_reg[6][111]  ( .CLK(n215), .D(N128), .Q(\ram[6][111] ) );
  LATCHX1_HVT \ram_reg[6][110]  ( .CLK(n215), .D(N127), .Q(\ram[6][110] ) );
  LATCHX1_HVT \ram_reg[6][109]  ( .CLK(n215), .D(N126), .Q(\ram[6][109] ) );
  LATCHX1_HVT \ram_reg[6][108]  ( .CLK(n212), .D(N125), .Q(\ram[6][108] ) );
  LATCHX1_HVT \ram_reg[6][107]  ( .CLK(n209), .D(N124), .Q(\ram[6][107] ) );
  LATCHX1_HVT \ram_reg[6][106]  ( .CLK(n215), .D(N123), .Q(\ram[6][106] ) );
  LATCHX1_HVT \ram_reg[6][105]  ( .CLK(n215), .D(N122), .Q(\ram[6][105] ) );
  LATCHX1_HVT \ram_reg[6][104]  ( .CLK(n215), .D(N121), .Q(\ram[6][104] ) );
  LATCHX1_HVT \ram_reg[6][103]  ( .CLK(n214), .D(N120), .Q(\ram[6][103] ) );
  LATCHX1_HVT \ram_reg[6][102]  ( .CLK(n213), .D(N119), .Q(\ram[6][102] ) );
  LATCHX1_HVT \ram_reg[6][101]  ( .CLK(n213), .D(N118), .Q(\ram[6][101] ) );
  LATCHX1_HVT \ram_reg[6][100]  ( .CLK(n214), .D(N117), .Q(\ram[6][100] ) );
  LATCHX1_HVT \ram_reg[6][99]  ( .CLK(n212), .D(N116), .Q(\ram[6][99] ) );
  LATCHX1_HVT \ram_reg[6][98]  ( .CLK(n213), .D(N114), .Q(\ram[6][98] ) );
  LATCHX1_HVT \ram_reg[6][97]  ( .CLK(n214), .D(N113), .Q(\ram[6][97] ) );
  LATCHX1_HVT \ram_reg[6][96]  ( .CLK(n218), .D(N112), .Q(\ram[6][96] ) );
  LATCHX1_HVT \ram_reg[6][95]  ( .CLK(n210), .D(N111), .Q(\ram[6][95] ) );
  LATCHX1_HVT \ram_reg[6][94]  ( .CLK(n210), .D(N110), .Q(\ram[6][94] ) );
  LATCHX1_HVT \ram_reg[6][93]  ( .CLK(n210), .D(N109), .Q(\ram[6][93] ) );
  LATCHX1_HVT \ram_reg[6][92]  ( .CLK(n209), .D(N108), .Q(\ram[6][92] ) );
  LATCHX1_HVT \ram_reg[6][91]  ( .CLK(n209), .D(N107), .Q(\ram[6][91] ) );
  LATCHX1_HVT \ram_reg[6][90]  ( .CLK(n210), .D(N106), .Q(\ram[6][90] ) );
  LATCHX1_HVT \ram_reg[6][89]  ( .CLK(n209), .D(N105), .Q(\ram[6][89] ) );
  LATCHX1_HVT \ram_reg[6][88]  ( .CLK(n210), .D(N104), .Q(\ram[6][88] ) );
  LATCHX1_HVT \ram_reg[6][87]  ( .CLK(n218), .D(N103), .Q(\ram[6][87] ) );
  LATCHX1_HVT \ram_reg[6][86]  ( .CLK(n217), .D(N102), .Q(\ram[6][86] ) );
  LATCHX1_HVT \ram_reg[6][85]  ( .CLK(n216), .D(N101), .Q(\ram[6][85] ) );
  LATCHX1_HVT \ram_reg[6][84]  ( .CLK(n216), .D(N100), .Q(\ram[6][84] ) );
  LATCHX1_HVT \ram_reg[6][83]  ( .CLK(n211), .D(N99), .Q(\ram[6][83] ) );
  LATCHX1_HVT \ram_reg[6][82]  ( .CLK(n217), .D(N98), .Q(\ram[6][82] ) );
  LATCHX1_HVT \ram_reg[6][81]  ( .CLK(n216), .D(N97), .Q(\ram[6][81] ) );
  LATCHX1_HVT \ram_reg[6][80]  ( .CLK(n217), .D(N96), .Q(\ram[6][80] ) );
  LATCHX1_HVT \ram_reg[6][79]  ( .CLK(n211), .D(N95), .Q(\ram[6][79] ) );
  LATCHX1_HVT \ram_reg[6][78]  ( .CLK(n210), .D(N94), .Q(\ram[6][78] ) );
  LATCHX1_HVT \ram_reg[6][77]  ( .CLK(n211), .D(N93), .Q(\ram[6][77] ) );
  LATCHX1_HVT \ram_reg[6][76]  ( .CLK(n210), .D(N92), .Q(\ram[6][76] ) );
  LATCHX1_HVT \ram_reg[6][75]  ( .CLK(n210), .D(N91), .Q(\ram[6][75] ) );
  LATCHX1_HVT \ram_reg[6][74]  ( .CLK(n208), .D(N90), .Q(\ram[6][74] ) );
  LATCHX1_HVT \ram_reg[6][73]  ( .CLK(n211), .D(N89), .Q(\ram[6][73] ) );
  LATCHX1_HVT \ram_reg[6][72]  ( .CLK(n211), .D(N88), .Q(\ram[6][72] ) );
  LATCHX1_HVT \ram_reg[6][71]  ( .CLK(n214), .D(N87), .Q(\ram[6][71] ) );
  LATCHX1_HVT \ram_reg[6][70]  ( .CLK(n214), .D(N86), .Q(\ram[6][70] ) );
  LATCHX1_HVT \ram_reg[6][69]  ( .CLK(n213), .D(N85), .Q(\ram[6][69] ) );
  LATCHX1_HVT \ram_reg[6][68]  ( .CLK(n214), .D(N84), .Q(\ram[6][68] ) );
  LATCHX1_HVT \ram_reg[6][67]  ( .CLK(n213), .D(N83), .Q(\ram[6][67] ) );
  LATCHX1_HVT \ram_reg[6][66]  ( .CLK(n212), .D(N82), .Q(\ram[6][66] ) );
  LATCHX1_HVT \ram_reg[6][65]  ( .CLK(n213), .D(N81), .Q(\ram[6][65] ) );
  LATCHX1_HVT \ram_reg[6][64]  ( .CLK(n218), .D(N80), .Q(\ram[6][64] ) );
  LATCHX1_HVT \ram_reg[6][63]  ( .CLK(n212), .D(N79), .Q(\ram[6][63] ) );
  LATCHX1_HVT \ram_reg[6][62]  ( .CLK(n212), .D(N78), .Q(\ram[6][62] ) );
  LATCHX1_HVT \ram_reg[6][61]  ( .CLK(n212), .D(N77), .Q(\ram[6][61] ) );
  LATCHX1_HVT \ram_reg[6][60]  ( .CLK(n212), .D(N76), .Q(\ram[6][60] ) );
  LATCHX1_HVT \ram_reg[6][59]  ( .CLK(n212), .D(N75), .Q(\ram[6][59] ) );
  LATCHX1_HVT \ram_reg[6][58]  ( .CLK(n211), .D(N74), .Q(\ram[6][58] ) );
  LATCHX1_HVT \ram_reg[6][57]  ( .CLK(n212), .D(N73), .Q(\ram[6][57] ) );
  LATCHX1_HVT \ram_reg[6][56]  ( .CLK(n212), .D(N72), .Q(\ram[6][56] ) );
  LATCHX1_HVT \ram_reg[6][55]  ( .CLK(n218), .D(N71), .Q(\ram[6][55] ) );
  LATCHX1_HVT \ram_reg[6][54]  ( .CLK(n216), .D(N70), .Q(\ram[6][54] ) );
  LATCHX1_HVT \ram_reg[6][53]  ( .CLK(n216), .D(N69), .Q(\ram[6][53] ) );
  LATCHX1_HVT \ram_reg[6][52]  ( .CLK(n217), .D(N68), .Q(\ram[6][52] ) );
  LATCHX1_HVT \ram_reg[6][51]  ( .CLK(n211), .D(N67), .Q(\ram[6][51] ) );
  LATCHX1_HVT \ram_reg[6][50]  ( .CLK(n208), .D(N66), .Q(\ram[6][50] ) );
  LATCHX1_HVT \ram_reg[6][49]  ( .CLK(n217), .D(N65), .Q(\ram[6][49] ) );
  LATCHX1_HVT \ram_reg[6][48]  ( .CLK(n217), .D(N64), .Q(\ram[6][48] ) );
  LATCHX1_HVT \ram_reg[6][47]  ( .CLK(n215), .D(N63), .Q(\ram[6][47] ) );
  LATCHX1_HVT \ram_reg[6][46]  ( .CLK(n215), .D(N62), .Q(\ram[6][46] ) );
  LATCHX1_HVT \ram_reg[6][45]  ( .CLK(n215), .D(N61), .Q(\ram[6][45] ) );
  LATCHX1_HVT \ram_reg[6][44]  ( .CLK(n215), .D(N60), .Q(\ram[6][44] ) );
  LATCHX1_HVT \ram_reg[6][43]  ( .CLK(n212), .D(N59), .Q(\ram[6][43] ) );
  LATCHX1_HVT \ram_reg[6][42]  ( .CLK(n216), .D(N58), .Q(\ram[6][42] ) );
  LATCHX1_HVT \ram_reg[6][41]  ( .CLK(n209), .D(N57), .Q(\ram[6][41] ) );
  LATCHX1_HVT \ram_reg[6][40]  ( .CLK(n215), .D(N56), .Q(\ram[6][40] ) );
  LATCHX1_HVT \ram_reg[6][39]  ( .CLK(n214), .D(N55), .Q(\ram[6][39] ) );
  LATCHX1_HVT \ram_reg[6][38]  ( .CLK(n214), .D(N54), .Q(\ram[6][38] ) );
  LATCHX1_HVT \ram_reg[6][37]  ( .CLK(n213), .D(N53), .Q(\ram[6][37] ) );
  LATCHX1_HVT \ram_reg[6][36]  ( .CLK(n213), .D(N52), .Q(\ram[6][36] ) );
  LATCHX1_HVT \ram_reg[6][35]  ( .CLK(n213), .D(N51), .Q(\ram[6][35] ) );
  LATCHX1_HVT \ram_reg[6][34]  ( .CLK(n215), .D(N50), .Q(\ram[6][34] ) );
  LATCHX1_HVT \ram_reg[6][33]  ( .CLK(n214), .D(N49), .Q(\ram[6][33] ) );
  LATCHX1_HVT \ram_reg[6][32]  ( .CLK(n218), .D(N48), .Q(\ram[6][32] ) );
  LATCHX1_HVT \ram_reg[6][31]  ( .CLK(n208), .D(N47), .Q(\ram[6][31] ) );
  LATCHX1_HVT \ram_reg[6][30]  ( .CLK(n208), .D(N46), .Q(\ram[6][30] ) );
  LATCHX1_HVT \ram_reg[6][29]  ( .CLK(n208), .D(N45), .Q(\ram[6][29] ) );
  LATCHX1_HVT \ram_reg[6][28]  ( .CLK(n208), .D(N44), .Q(\ram[6][28] ) );
  LATCHX1_HVT \ram_reg[6][27]  ( .CLK(n208), .D(N43), .Q(\ram[6][27] ) );
  LATCHX1_HVT \ram_reg[6][26]  ( .CLK(n208), .D(N42), .Q(\ram[6][26] ) );
  LATCHX1_HVT \ram_reg[6][25]  ( .CLK(n208), .D(N41), .Q(\ram[6][25] ) );
  LATCHX1_HVT \ram_reg[6][24]  ( .CLK(n208), .D(N40), .Q(\ram[6][24] ) );
  LATCHX1_HVT \ram_reg[6][23]  ( .CLK(n218), .D(N39), .Q(\ram[6][23] ) );
  LATCHX1_HVT \ram_reg[6][22]  ( .CLK(n217), .D(N38), .Q(\ram[6][22] ) );
  LATCHX1_HVT \ram_reg[6][21]  ( .CLK(n216), .D(N37), .Q(\ram[6][21] ) );
  LATCHX1_HVT \ram_reg[6][20]  ( .CLK(n216), .D(N36), .Q(\ram[6][20] ) );
  LATCHX1_HVT \ram_reg[6][19]  ( .CLK(n208), .D(N35), .Q(\ram[6][19] ) );
  LATCHX1_HVT \ram_reg[6][18]  ( .CLK(n216), .D(N34), .Q(\ram[6][18] ) );
  LATCHX1_HVT \ram_reg[6][17]  ( .CLK(n217), .D(N33), .Q(\ram[6][17] ) );
  LATCHX1_HVT \ram_reg[6][16]  ( .CLK(n217), .D(N32), .Q(\ram[6][16] ) );
  LATCHX1_HVT \ram_reg[6][15]  ( .CLK(n211), .D(N31), .Q(\ram[6][15] ) );
  LATCHX1_HVT \ram_reg[6][14]  ( .CLK(n211), .D(N30), .Q(\ram[6][14] ) );
  LATCHX1_HVT \ram_reg[6][13]  ( .CLK(n210), .D(N29), .Q(\ram[6][13] ) );
  LATCHX1_HVT \ram_reg[6][12]  ( .CLK(n210), .D(N28), .Q(\ram[6][12] ) );
  LATCHX1_HVT \ram_reg[6][11]  ( .CLK(n211), .D(N27), .Q(\ram[6][11] ) );
  LATCHX1_HVT \ram_reg[6][10]  ( .CLK(n210), .D(N26), .Q(\ram[6][10] ) );
  LATCHX1_HVT \ram_reg[6][9]  ( .CLK(n210), .D(N25), .Q(\ram[6][9] ) );
  LATCHX1_HVT \ram_reg[6][8]  ( .CLK(n211), .D(N24), .Q(\ram[6][8] ) );
  LATCHX1_HVT \ram_reg[6][7]  ( .CLK(n214), .D(N23), .Q(\ram[6][7] ) );
  LATCHX1_HVT \ram_reg[6][6]  ( .CLK(n214), .D(N22), .Q(\ram[6][6] ) );
  LATCHX1_HVT \ram_reg[6][5]  ( .CLK(n213), .D(N21), .Q(\ram[6][5] ) );
  LATCHX1_HVT \ram_reg[6][4]  ( .CLK(n213), .D(N20), .Q(\ram[6][4] ) );
  LATCHX1_HVT \ram_reg[6][3]  ( .CLK(n212), .D(N19), .Q(\ram[6][3] ) );
  LATCHX1_HVT \ram_reg[6][2]  ( .CLK(n213), .D(N18), .Q(\ram[6][2] ) );
  LATCHX1_HVT \ram_reg[6][1]  ( .CLK(n214), .D(N17), .Q(\ram[6][1] ) );
  LATCHX1_HVT \ram_reg[6][0]  ( .CLK(n218), .D(N16), .Q(\ram[6][0] ) );
  LATCHX1_HVT \ram_reg[5][255]  ( .CLK(N288), .D(N273), .Q(\ram[5][255] ) );
  LATCHX1_HVT \ram_reg[5][254]  ( .CLK(N288), .D(N272), .Q(\ram[5][254] ) );
  LATCHX1_HVT \ram_reg[5][253]  ( .CLK(N288), .D(N271), .Q(\ram[5][253] ) );
  LATCHX1_HVT \ram_reg[5][252]  ( .CLK(N288), .D(N270), .Q(\ram[5][252] ) );
  LATCHX1_HVT \ram_reg[5][251]  ( .CLK(n251), .D(N269), .Q(\ram[5][251] ) );
  LATCHX1_HVT \ram_reg[5][250]  ( .CLK(n243), .D(N268), .Q(\ram[5][250] ) );
  LATCHX1_HVT \ram_reg[5][249]  ( .CLK(n243), .D(N267), .Q(\ram[5][249] ) );
  LATCHX1_HVT \ram_reg[5][248]  ( .CLK(n243), .D(N266), .Q(\ram[5][248] ) );
  LATCHX1_HVT \ram_reg[5][247]  ( .CLK(n243), .D(N265), .Q(\ram[5][247] ) );
  LATCHX1_HVT \ram_reg[5][246]  ( .CLK(n243), .D(N264), .Q(\ram[5][246] ) );
  LATCHX1_HVT \ram_reg[5][245]  ( .CLK(n243), .D(N263), .Q(\ram[5][245] ) );
  LATCHX1_HVT \ram_reg[5][244]  ( .CLK(n243), .D(N262), .Q(\ram[5][244] ) );
  LATCHX1_HVT \ram_reg[5][243]  ( .CLK(n243), .D(N261), .Q(\ram[5][243] ) );
  LATCHX1_HVT \ram_reg[5][242]  ( .CLK(n243), .D(N260), .Q(\ram[5][242] ) );
  LATCHX1_HVT \ram_reg[5][241]  ( .CLK(n242), .D(N259), .Q(\ram[5][241] ) );
  LATCHX1_HVT \ram_reg[5][240]  ( .CLK(n242), .D(N258), .Q(\ram[5][240] ) );
  LATCHX1_HVT \ram_reg[5][239]  ( .CLK(n242), .D(N257), .Q(\ram[5][239] ) );
  LATCHX1_HVT \ram_reg[5][238]  ( .CLK(n242), .D(N256), .Q(\ram[5][238] ) );
  LATCHX1_HVT \ram_reg[5][237]  ( .CLK(n242), .D(N255), .Q(\ram[5][237] ) );
  LATCHX1_HVT \ram_reg[5][236]  ( .CLK(n242), .D(N254), .Q(\ram[5][236] ) );
  LATCHX1_HVT \ram_reg[5][235]  ( .CLK(n242), .D(N253), .Q(\ram[5][235] ) );
  LATCHX1_HVT \ram_reg[5][234]  ( .CLK(n242), .D(N252), .Q(\ram[5][234] ) );
  LATCHX1_HVT \ram_reg[5][233]  ( .CLK(n242), .D(N251), .Q(\ram[5][233] ) );
  LATCHX1_HVT \ram_reg[5][232]  ( .CLK(n242), .D(N250), .Q(\ram[5][232] ) );
  LATCHX1_HVT \ram_reg[5][231]  ( .CLK(n242), .D(N249), .Q(\ram[5][231] ) );
  LATCHX1_HVT \ram_reg[5][230]  ( .CLK(n241), .D(N248), .Q(\ram[5][230] ) );
  LATCHX1_HVT \ram_reg[5][229]  ( .CLK(n241), .D(N247), .Q(\ram[5][229] ) );
  LATCHX1_HVT \ram_reg[5][228]  ( .CLK(n241), .D(N246), .Q(\ram[5][228] ) );
  LATCHX1_HVT \ram_reg[5][227]  ( .CLK(n251), .D(N245), .Q(\ram[5][227] ) );
  LATCHX1_HVT \ram_reg[5][226]  ( .CLK(n251), .D(N244), .Q(\ram[5][226] ) );
  LATCHX1_HVT \ram_reg[5][225]  ( .CLK(n251), .D(N243), .Q(\ram[5][225] ) );
  LATCHX1_HVT \ram_reg[5][224]  ( .CLK(n251), .D(N242), .Q(\ram[5][224] ) );
  LATCHX1_HVT \ram_reg[5][223]  ( .CLK(n251), .D(N241), .Q(\ram[5][223] ) );
  LATCHX1_HVT \ram_reg[5][222]  ( .CLK(n251), .D(N240), .Q(\ram[5][222] ) );
  LATCHX1_HVT \ram_reg[5][221]  ( .CLK(n251), .D(N239), .Q(\ram[5][221] ) );
  LATCHX1_HVT \ram_reg[5][220]  ( .CLK(n251), .D(N238), .Q(\ram[5][220] ) );
  LATCHX1_HVT \ram_reg[5][219]  ( .CLK(n251), .D(N237), .Q(\ram[5][219] ) );
  LATCHX1_HVT \ram_reg[5][218]  ( .CLK(n251), .D(N236), .Q(\ram[5][218] ) );
  LATCHX1_HVT \ram_reg[5][217]  ( .CLK(n250), .D(N235), .Q(\ram[5][217] ) );
  LATCHX1_HVT \ram_reg[5][216]  ( .CLK(n250), .D(N234), .Q(\ram[5][216] ) );
  LATCHX1_HVT \ram_reg[5][215]  ( .CLK(n250), .D(N233), .Q(\ram[5][215] ) );
  LATCHX1_HVT \ram_reg[5][214]  ( .CLK(n250), .D(N232), .Q(\ram[5][214] ) );
  LATCHX1_HVT \ram_reg[5][213]  ( .CLK(n250), .D(N231), .Q(\ram[5][213] ) );
  LATCHX1_HVT \ram_reg[5][212]  ( .CLK(n250), .D(N230), .Q(\ram[5][212] ) );
  LATCHX1_HVT \ram_reg[5][211]  ( .CLK(n250), .D(N229), .Q(\ram[5][211] ) );
  LATCHX1_HVT \ram_reg[5][210]  ( .CLK(n250), .D(N228), .Q(\ram[5][210] ) );
  LATCHX1_HVT \ram_reg[5][209]  ( .CLK(n250), .D(N227), .Q(\ram[5][209] ) );
  LATCHX1_HVT \ram_reg[5][208]  ( .CLK(n250), .D(N226), .Q(\ram[5][208] ) );
  LATCHX1_HVT \ram_reg[5][207]  ( .CLK(n249), .D(N225), .Q(\ram[5][207] ) );
  LATCHX1_HVT \ram_reg[5][206]  ( .CLK(n249), .D(N224), .Q(\ram[5][206] ) );
  LATCHX1_HVT \ram_reg[5][205]  ( .CLK(n249), .D(N223), .Q(\ram[5][205] ) );
  LATCHX1_HVT \ram_reg[5][204]  ( .CLK(n249), .D(N222), .Q(\ram[5][204] ) );
  LATCHX1_HVT \ram_reg[5][203]  ( .CLK(n249), .D(N221), .Q(\ram[5][203] ) );
  LATCHX1_HVT \ram_reg[5][202]  ( .CLK(n249), .D(N220), .Q(\ram[5][202] ) );
  LATCHX1_HVT \ram_reg[5][201]  ( .CLK(n249), .D(N219), .Q(\ram[5][201] ) );
  LATCHX1_HVT \ram_reg[5][200]  ( .CLK(n249), .D(N218), .Q(\ram[5][200] ) );
  LATCHX1_HVT \ram_reg[5][199]  ( .CLK(n249), .D(N217), .Q(\ram[5][199] ) );
  LATCHX1_HVT \ram_reg[5][198]  ( .CLK(n249), .D(N216), .Q(\ram[5][198] ) );
  LATCHX1_HVT \ram_reg[5][197]  ( .CLK(n249), .D(N214), .Q(\ram[5][197] ) );
  LATCHX1_HVT \ram_reg[5][196]  ( .CLK(n248), .D(N213), .Q(\ram[5][196] ) );
  LATCHX1_HVT \ram_reg[5][195]  ( .CLK(n248), .D(N212), .Q(\ram[5][195] ) );
  LATCHX1_HVT \ram_reg[5][194]  ( .CLK(n248), .D(N211), .Q(\ram[5][194] ) );
  LATCHX1_HVT \ram_reg[5][193]  ( .CLK(n248), .D(N210), .Q(\ram[5][193] ) );
  LATCHX1_HVT \ram_reg[5][192]  ( .CLK(n248), .D(N209), .Q(\ram[5][192] ) );
  LATCHX1_HVT \ram_reg[5][191]  ( .CLK(n248), .D(N208), .Q(\ram[5][191] ) );
  LATCHX1_HVT \ram_reg[5][190]  ( .CLK(n248), .D(N207), .Q(\ram[5][190] ) );
  LATCHX1_HVT \ram_reg[5][189]  ( .CLK(n248), .D(N206), .Q(\ram[5][189] ) );
  LATCHX1_HVT \ram_reg[5][188]  ( .CLK(n248), .D(N205), .Q(\ram[5][188] ) );
  LATCHX1_HVT \ram_reg[5][187]  ( .CLK(n248), .D(N204), .Q(\ram[5][187] ) );
  LATCHX1_HVT \ram_reg[5][186]  ( .CLK(n248), .D(N203), .Q(\ram[5][186] ) );
  LATCHX1_HVT \ram_reg[5][185]  ( .CLK(n247), .D(N202), .Q(\ram[5][185] ) );
  LATCHX1_HVT \ram_reg[5][184]  ( .CLK(n247), .D(N201), .Q(\ram[5][184] ) );
  LATCHX1_HVT \ram_reg[5][183]  ( .CLK(n247), .D(N200), .Q(\ram[5][183] ) );
  LATCHX1_HVT \ram_reg[5][182]  ( .CLK(n247), .D(N199), .Q(\ram[5][182] ) );
  LATCHX1_HVT \ram_reg[5][181]  ( .CLK(n247), .D(N198), .Q(\ram[5][181] ) );
  LATCHX1_HVT \ram_reg[5][180]  ( .CLK(n247), .D(N197), .Q(\ram[5][180] ) );
  LATCHX1_HVT \ram_reg[5][179]  ( .CLK(n247), .D(N196), .Q(\ram[5][179] ) );
  LATCHX1_HVT \ram_reg[5][178]  ( .CLK(n247), .D(N195), .Q(\ram[5][178] ) );
  LATCHX1_HVT \ram_reg[5][177]  ( .CLK(n247), .D(N194), .Q(\ram[5][177] ) );
  LATCHX1_HVT \ram_reg[5][176]  ( .CLK(n247), .D(N193), .Q(\ram[5][176] ) );
  LATCHX1_HVT \ram_reg[5][175]  ( .CLK(n247), .D(N192), .Q(\ram[5][175] ) );
  LATCHX1_HVT \ram_reg[5][174]  ( .CLK(n246), .D(N191), .Q(\ram[5][174] ) );
  LATCHX1_HVT \ram_reg[5][173]  ( .CLK(n246), .D(N190), .Q(\ram[5][173] ) );
  LATCHX1_HVT \ram_reg[5][172]  ( .CLK(n246), .D(N189), .Q(\ram[5][172] ) );
  LATCHX1_HVT \ram_reg[5][171]  ( .CLK(n246), .D(N188), .Q(\ram[5][171] ) );
  LATCHX1_HVT \ram_reg[5][170]  ( .CLK(n246), .D(N187), .Q(\ram[5][170] ) );
  LATCHX1_HVT \ram_reg[5][169]  ( .CLK(n246), .D(N186), .Q(\ram[5][169] ) );
  LATCHX1_HVT \ram_reg[5][168]  ( .CLK(n246), .D(N185), .Q(\ram[5][168] ) );
  LATCHX1_HVT \ram_reg[5][167]  ( .CLK(n246), .D(N184), .Q(\ram[5][167] ) );
  LATCHX1_HVT \ram_reg[5][166]  ( .CLK(n246), .D(N183), .Q(\ram[5][166] ) );
  LATCHX1_HVT \ram_reg[5][165]  ( .CLK(n246), .D(N182), .Q(\ram[5][165] ) );
  LATCHX1_HVT \ram_reg[5][164]  ( .CLK(n246), .D(N181), .Q(\ram[5][164] ) );
  LATCHX1_HVT \ram_reg[5][163]  ( .CLK(n245), .D(N180), .Q(\ram[5][163] ) );
  LATCHX1_HVT \ram_reg[5][162]  ( .CLK(n245), .D(N179), .Q(\ram[5][162] ) );
  LATCHX1_HVT \ram_reg[5][161]  ( .CLK(n245), .D(N178), .Q(\ram[5][161] ) );
  LATCHX1_HVT \ram_reg[5][160]  ( .CLK(n245), .D(N177), .Q(\ram[5][160] ) );
  LATCHX1_HVT \ram_reg[5][159]  ( .CLK(n245), .D(N176), .Q(\ram[5][159] ) );
  LATCHX1_HVT \ram_reg[5][158]  ( .CLK(n245), .D(N175), .Q(\ram[5][158] ) );
  LATCHX1_HVT \ram_reg[5][157]  ( .CLK(n245), .D(N174), .Q(\ram[5][157] ) );
  LATCHX1_HVT \ram_reg[5][156]  ( .CLK(n245), .D(N173), .Q(\ram[5][156] ) );
  LATCHX1_HVT \ram_reg[5][155]  ( .CLK(n245), .D(N172), .Q(\ram[5][155] ) );
  LATCHX1_HVT \ram_reg[5][154]  ( .CLK(n245), .D(N171), .Q(\ram[5][154] ) );
  LATCHX1_HVT \ram_reg[5][153]  ( .CLK(n245), .D(N170), .Q(\ram[5][153] ) );
  LATCHX1_HVT \ram_reg[5][152]  ( .CLK(n244), .D(N169), .Q(\ram[5][152] ) );
  LATCHX1_HVT \ram_reg[5][151]  ( .CLK(n244), .D(N168), .Q(\ram[5][151] ) );
  LATCHX1_HVT \ram_reg[5][150]  ( .CLK(n244), .D(N167), .Q(\ram[5][150] ) );
  LATCHX1_HVT \ram_reg[5][149]  ( .CLK(n244), .D(N166), .Q(\ram[5][149] ) );
  LATCHX1_HVT \ram_reg[5][148]  ( .CLK(n244), .D(N165), .Q(\ram[5][148] ) );
  LATCHX1_HVT \ram_reg[5][147]  ( .CLK(n244), .D(N164), .Q(\ram[5][147] ) );
  LATCHX1_HVT \ram_reg[5][146]  ( .CLK(n244), .D(N163), .Q(\ram[5][146] ) );
  LATCHX1_HVT \ram_reg[5][145]  ( .CLK(n244), .D(N162), .Q(\ram[5][145] ) );
  LATCHX1_HVT \ram_reg[5][144]  ( .CLK(n244), .D(N161), .Q(\ram[5][144] ) );
  LATCHX1_HVT \ram_reg[5][143]  ( .CLK(n244), .D(N160), .Q(\ram[5][143] ) );
  LATCHX1_HVT \ram_reg[5][142]  ( .CLK(n244), .D(N159), .Q(\ram[5][142] ) );
  LATCHX1_HVT \ram_reg[5][141]  ( .CLK(n243), .D(N158), .Q(\ram[5][141] ) );
  LATCHX1_HVT \ram_reg[5][140]  ( .CLK(n243), .D(N157), .Q(\ram[5][140] ) );
  LATCHX1_HVT \ram_reg[5][139]  ( .CLK(n243), .D(N156), .Q(\ram[5][139] ) );
  LATCHX1_HVT \ram_reg[5][138]  ( .CLK(n242), .D(N155), .Q(\ram[5][138] ) );
  LATCHX1_HVT \ram_reg[5][137]  ( .CLK(n251), .D(N154), .Q(\ram[5][137] ) );
  LATCHX1_HVT \ram_reg[5][136]  ( .CLK(n250), .D(N153), .Q(\ram[5][136] ) );
  LATCHX1_HVT \ram_reg[5][135]  ( .CLK(n250), .D(N152), .Q(\ram[5][135] ) );
  LATCHX1_HVT \ram_reg[5][134]  ( .CLK(n249), .D(N151), .Q(\ram[5][134] ) );
  LATCHX1_HVT \ram_reg[5][133]  ( .CLK(n248), .D(N150), .Q(\ram[5][133] ) );
  LATCHX1_HVT \ram_reg[5][132]  ( .CLK(n247), .D(N149), .Q(\ram[5][132] ) );
  LATCHX1_HVT \ram_reg[5][131]  ( .CLK(n246), .D(N148), .Q(\ram[5][131] ) );
  LATCHX1_HVT \ram_reg[5][130]  ( .CLK(n245), .D(N147), .Q(\ram[5][130] ) );
  LATCHX1_HVT \ram_reg[5][129]  ( .CLK(n244), .D(N146), .Q(\ram[5][129] ) );
  LATCHX1_HVT \ram_reg[5][128]  ( .CLK(n241), .D(N145), .Q(\ram[5][128] ) );
  LATCHX1_HVT \ram_reg[5][127]  ( .CLK(n232), .D(N144), .Q(\ram[5][127] ) );
  LATCHX1_HVT \ram_reg[5][126]  ( .CLK(n232), .D(N143), .Q(\ram[5][126] ) );
  LATCHX1_HVT \ram_reg[5][125]  ( .CLK(n232), .D(N142), .Q(\ram[5][125] ) );
  LATCHX1_HVT \ram_reg[5][124]  ( .CLK(n232), .D(N141), .Q(\ram[5][124] ) );
  LATCHX1_HVT \ram_reg[5][123]  ( .CLK(n232), .D(N140), .Q(\ram[5][123] ) );
  LATCHX1_HVT \ram_reg[5][122]  ( .CLK(n231), .D(N139), .Q(\ram[5][122] ) );
  LATCHX1_HVT \ram_reg[5][121]  ( .CLK(n232), .D(N138), .Q(\ram[5][121] ) );
  LATCHX1_HVT \ram_reg[5][120]  ( .CLK(n232), .D(N137), .Q(\ram[5][120] ) );
  LATCHX1_HVT \ram_reg[5][119]  ( .CLK(n241), .D(N136), .Q(\ram[5][119] ) );
  LATCHX1_HVT \ram_reg[5][118]  ( .CLK(n240), .D(N135), .Q(\ram[5][118] ) );
  LATCHX1_HVT \ram_reg[5][117]  ( .CLK(n240), .D(N134), .Q(\ram[5][117] ) );
  LATCHX1_HVT \ram_reg[5][116]  ( .CLK(n239), .D(N133), .Q(\ram[5][116] ) );
  LATCHX1_HVT \ram_reg[5][115]  ( .CLK(n234), .D(N132), .Q(\ram[5][115] ) );
  LATCHX1_HVT \ram_reg[5][114]  ( .CLK(n239), .D(N131), .Q(\ram[5][114] ) );
  LATCHX1_HVT \ram_reg[5][113]  ( .CLK(n239), .D(N130), .Q(\ram[5][113] ) );
  LATCHX1_HVT \ram_reg[5][112]  ( .CLK(n240), .D(N129), .Q(\ram[5][112] ) );
  LATCHX1_HVT \ram_reg[5][111]  ( .CLK(n238), .D(N128), .Q(\ram[5][111] ) );
  LATCHX1_HVT \ram_reg[5][110]  ( .CLK(n238), .D(N127), .Q(\ram[5][110] ) );
  LATCHX1_HVT \ram_reg[5][109]  ( .CLK(n238), .D(N126), .Q(\ram[5][109] ) );
  LATCHX1_HVT \ram_reg[5][108]  ( .CLK(n235), .D(N125), .Q(\ram[5][108] ) );
  LATCHX1_HVT \ram_reg[5][107]  ( .CLK(n232), .D(N124), .Q(\ram[5][107] ) );
  LATCHX1_HVT \ram_reg[5][106]  ( .CLK(n238), .D(N123), .Q(\ram[5][106] ) );
  LATCHX1_HVT \ram_reg[5][105]  ( .CLK(n238), .D(N122), .Q(\ram[5][105] ) );
  LATCHX1_HVT \ram_reg[5][104]  ( .CLK(n238), .D(N121), .Q(\ram[5][104] ) );
  LATCHX1_HVT \ram_reg[5][103]  ( .CLK(n237), .D(N120), .Q(\ram[5][103] ) );
  LATCHX1_HVT \ram_reg[5][102]  ( .CLK(n236), .D(N119), .Q(\ram[5][102] ) );
  LATCHX1_HVT \ram_reg[5][101]  ( .CLK(n236), .D(N118), .Q(\ram[5][101] ) );
  LATCHX1_HVT \ram_reg[5][100]  ( .CLK(n237), .D(N117), .Q(\ram[5][100] ) );
  LATCHX1_HVT \ram_reg[5][99]  ( .CLK(n235), .D(N116), .Q(\ram[5][99] ) );
  LATCHX1_HVT \ram_reg[5][98]  ( .CLK(n236), .D(N114), .Q(\ram[5][98] ) );
  LATCHX1_HVT \ram_reg[5][97]  ( .CLK(n237), .D(N113), .Q(\ram[5][97] ) );
  LATCHX1_HVT \ram_reg[5][96]  ( .CLK(n241), .D(N112), .Q(\ram[5][96] ) );
  LATCHX1_HVT \ram_reg[5][95]  ( .CLK(n233), .D(N111), .Q(\ram[5][95] ) );
  LATCHX1_HVT \ram_reg[5][94]  ( .CLK(n233), .D(N110), .Q(\ram[5][94] ) );
  LATCHX1_HVT \ram_reg[5][93]  ( .CLK(n233), .D(N109), .Q(\ram[5][93] ) );
  LATCHX1_HVT \ram_reg[5][92]  ( .CLK(n232), .D(N108), .Q(\ram[5][92] ) );
  LATCHX1_HVT \ram_reg[5][91]  ( .CLK(n232), .D(N107), .Q(\ram[5][91] ) );
  LATCHX1_HVT \ram_reg[5][90]  ( .CLK(n233), .D(N106), .Q(\ram[5][90] ) );
  LATCHX1_HVT \ram_reg[5][89]  ( .CLK(n232), .D(N105), .Q(\ram[5][89] ) );
  LATCHX1_HVT \ram_reg[5][88]  ( .CLK(n233), .D(N104), .Q(\ram[5][88] ) );
  LATCHX1_HVT \ram_reg[5][87]  ( .CLK(n241), .D(N103), .Q(\ram[5][87] ) );
  LATCHX1_HVT \ram_reg[5][86]  ( .CLK(n240), .D(N102), .Q(\ram[5][86] ) );
  LATCHX1_HVT \ram_reg[5][85]  ( .CLK(n239), .D(N101), .Q(\ram[5][85] ) );
  LATCHX1_HVT \ram_reg[5][84]  ( .CLK(n239), .D(N100), .Q(\ram[5][84] ) );
  LATCHX1_HVT \ram_reg[5][83]  ( .CLK(n234), .D(N99), .Q(\ram[5][83] ) );
  LATCHX1_HVT \ram_reg[5][82]  ( .CLK(n240), .D(N98), .Q(\ram[5][82] ) );
  LATCHX1_HVT \ram_reg[5][81]  ( .CLK(n239), .D(N97), .Q(\ram[5][81] ) );
  LATCHX1_HVT \ram_reg[5][80]  ( .CLK(n240), .D(N96), .Q(\ram[5][80] ) );
  LATCHX1_HVT \ram_reg[5][79]  ( .CLK(n234), .D(N95), .Q(\ram[5][79] ) );
  LATCHX1_HVT \ram_reg[5][78]  ( .CLK(n233), .D(N94), .Q(\ram[5][78] ) );
  LATCHX1_HVT \ram_reg[5][77]  ( .CLK(n234), .D(N93), .Q(\ram[5][77] ) );
  LATCHX1_HVT \ram_reg[5][76]  ( .CLK(n233), .D(N92), .Q(\ram[5][76] ) );
  LATCHX1_HVT \ram_reg[5][75]  ( .CLK(n233), .D(N91), .Q(\ram[5][75] ) );
  LATCHX1_HVT \ram_reg[5][74]  ( .CLK(n231), .D(N90), .Q(\ram[5][74] ) );
  LATCHX1_HVT \ram_reg[5][73]  ( .CLK(n234), .D(N89), .Q(\ram[5][73] ) );
  LATCHX1_HVT \ram_reg[5][72]  ( .CLK(n234), .D(N88), .Q(\ram[5][72] ) );
  LATCHX1_HVT \ram_reg[5][71]  ( .CLK(n237), .D(N87), .Q(\ram[5][71] ) );
  LATCHX1_HVT \ram_reg[5][70]  ( .CLK(n237), .D(N86), .Q(\ram[5][70] ) );
  LATCHX1_HVT \ram_reg[5][69]  ( .CLK(n236), .D(N85), .Q(\ram[5][69] ) );
  LATCHX1_HVT \ram_reg[5][68]  ( .CLK(n237), .D(N84), .Q(\ram[5][68] ) );
  LATCHX1_HVT \ram_reg[5][67]  ( .CLK(n236), .D(N83), .Q(\ram[5][67] ) );
  LATCHX1_HVT \ram_reg[5][66]  ( .CLK(n235), .D(N82), .Q(\ram[5][66] ) );
  LATCHX1_HVT \ram_reg[5][65]  ( .CLK(n236), .D(N81), .Q(\ram[5][65] ) );
  LATCHX1_HVT \ram_reg[5][64]  ( .CLK(n241), .D(N80), .Q(\ram[5][64] ) );
  LATCHX1_HVT \ram_reg[5][63]  ( .CLK(n235), .D(N79), .Q(\ram[5][63] ) );
  LATCHX1_HVT \ram_reg[5][62]  ( .CLK(n235), .D(N78), .Q(\ram[5][62] ) );
  LATCHX1_HVT \ram_reg[5][61]  ( .CLK(n235), .D(N77), .Q(\ram[5][61] ) );
  LATCHX1_HVT \ram_reg[5][60]  ( .CLK(n235), .D(N76), .Q(\ram[5][60] ) );
  LATCHX1_HVT \ram_reg[5][59]  ( .CLK(n235), .D(N75), .Q(\ram[5][59] ) );
  LATCHX1_HVT \ram_reg[5][58]  ( .CLK(n234), .D(N74), .Q(\ram[5][58] ) );
  LATCHX1_HVT \ram_reg[5][57]  ( .CLK(n235), .D(N73), .Q(\ram[5][57] ) );
  LATCHX1_HVT \ram_reg[5][56]  ( .CLK(n235), .D(N72), .Q(\ram[5][56] ) );
  LATCHX1_HVT \ram_reg[5][55]  ( .CLK(n241), .D(N71), .Q(\ram[5][55] ) );
  LATCHX1_HVT \ram_reg[5][54]  ( .CLK(n239), .D(N70), .Q(\ram[5][54] ) );
  LATCHX1_HVT \ram_reg[5][53]  ( .CLK(n239), .D(N69), .Q(\ram[5][53] ) );
  LATCHX1_HVT \ram_reg[5][52]  ( .CLK(n240), .D(N68), .Q(\ram[5][52] ) );
  LATCHX1_HVT \ram_reg[5][51]  ( .CLK(n234), .D(N67), .Q(\ram[5][51] ) );
  LATCHX1_HVT \ram_reg[5][50]  ( .CLK(n231), .D(N66), .Q(\ram[5][50] ) );
  LATCHX1_HVT \ram_reg[5][49]  ( .CLK(n240), .D(N65), .Q(\ram[5][49] ) );
  LATCHX1_HVT \ram_reg[5][48]  ( .CLK(n240), .D(N64), .Q(\ram[5][48] ) );
  LATCHX1_HVT \ram_reg[5][47]  ( .CLK(n238), .D(N63), .Q(\ram[5][47] ) );
  LATCHX1_HVT \ram_reg[5][46]  ( .CLK(n238), .D(N62), .Q(\ram[5][46] ) );
  LATCHX1_HVT \ram_reg[5][45]  ( .CLK(n238), .D(N61), .Q(\ram[5][45] ) );
  LATCHX1_HVT \ram_reg[5][44]  ( .CLK(n238), .D(N60), .Q(\ram[5][44] ) );
  LATCHX1_HVT \ram_reg[5][43]  ( .CLK(n235), .D(N59), .Q(\ram[5][43] ) );
  LATCHX1_HVT \ram_reg[5][42]  ( .CLK(n239), .D(N58), .Q(\ram[5][42] ) );
  LATCHX1_HVT \ram_reg[5][41]  ( .CLK(n232), .D(N57), .Q(\ram[5][41] ) );
  LATCHX1_HVT \ram_reg[5][40]  ( .CLK(n238), .D(N56), .Q(\ram[5][40] ) );
  LATCHX1_HVT \ram_reg[5][39]  ( .CLK(n237), .D(N55), .Q(\ram[5][39] ) );
  LATCHX1_HVT \ram_reg[5][38]  ( .CLK(n237), .D(N54), .Q(\ram[5][38] ) );
  LATCHX1_HVT \ram_reg[5][37]  ( .CLK(n236), .D(N53), .Q(\ram[5][37] ) );
  LATCHX1_HVT \ram_reg[5][36]  ( .CLK(n236), .D(N52), .Q(\ram[5][36] ) );
  LATCHX1_HVT \ram_reg[5][35]  ( .CLK(n236), .D(N51), .Q(\ram[5][35] ) );
  LATCHX1_HVT \ram_reg[5][34]  ( .CLK(n238), .D(N50), .Q(\ram[5][34] ) );
  LATCHX1_HVT \ram_reg[5][33]  ( .CLK(n237), .D(N49), .Q(\ram[5][33] ) );
  LATCHX1_HVT \ram_reg[5][32]  ( .CLK(n241), .D(N48), .Q(\ram[5][32] ) );
  LATCHX1_HVT \ram_reg[5][31]  ( .CLK(n231), .D(N47), .Q(\ram[5][31] ) );
  LATCHX1_HVT \ram_reg[5][30]  ( .CLK(n231), .D(N46), .Q(\ram[5][30] ) );
  LATCHX1_HVT \ram_reg[5][29]  ( .CLK(n231), .D(N45), .Q(\ram[5][29] ) );
  LATCHX1_HVT \ram_reg[5][28]  ( .CLK(n231), .D(N44), .Q(\ram[5][28] ) );
  LATCHX1_HVT \ram_reg[5][27]  ( .CLK(n231), .D(N43), .Q(\ram[5][27] ) );
  LATCHX1_HVT \ram_reg[5][26]  ( .CLK(n231), .D(N42), .Q(\ram[5][26] ) );
  LATCHX1_HVT \ram_reg[5][25]  ( .CLK(n231), .D(N41), .Q(\ram[5][25] ) );
  LATCHX1_HVT \ram_reg[5][24]  ( .CLK(n231), .D(N40), .Q(\ram[5][24] ) );
  LATCHX1_HVT \ram_reg[5][23]  ( .CLK(n241), .D(N39), .Q(\ram[5][23] ) );
  LATCHX1_HVT \ram_reg[5][22]  ( .CLK(n240), .D(N38), .Q(\ram[5][22] ) );
  LATCHX1_HVT \ram_reg[5][21]  ( .CLK(n239), .D(N37), .Q(\ram[5][21] ) );
  LATCHX1_HVT \ram_reg[5][20]  ( .CLK(n239), .D(N36), .Q(\ram[5][20] ) );
  LATCHX1_HVT \ram_reg[5][19]  ( .CLK(n231), .D(N35), .Q(\ram[5][19] ) );
  LATCHX1_HVT \ram_reg[5][18]  ( .CLK(n239), .D(N34), .Q(\ram[5][18] ) );
  LATCHX1_HVT \ram_reg[5][17]  ( .CLK(n240), .D(N33), .Q(\ram[5][17] ) );
  LATCHX1_HVT \ram_reg[5][16]  ( .CLK(n240), .D(N32), .Q(\ram[5][16] ) );
  LATCHX1_HVT \ram_reg[5][15]  ( .CLK(n234), .D(N31), .Q(\ram[5][15] ) );
  LATCHX1_HVT \ram_reg[5][14]  ( .CLK(n234), .D(N30), .Q(\ram[5][14] ) );
  LATCHX1_HVT \ram_reg[5][13]  ( .CLK(n233), .D(N29), .Q(\ram[5][13] ) );
  LATCHX1_HVT \ram_reg[5][12]  ( .CLK(n233), .D(N28), .Q(\ram[5][12] ) );
  LATCHX1_HVT \ram_reg[5][11]  ( .CLK(n234), .D(N27), .Q(\ram[5][11] ) );
  LATCHX1_HVT \ram_reg[5][10]  ( .CLK(n233), .D(N26), .Q(\ram[5][10] ) );
  LATCHX1_HVT \ram_reg[5][9]  ( .CLK(n233), .D(N25), .Q(\ram[5][9] ) );
  LATCHX1_HVT \ram_reg[5][8]  ( .CLK(n234), .D(N24), .Q(\ram[5][8] ) );
  LATCHX1_HVT \ram_reg[5][7]  ( .CLK(n237), .D(N23), .Q(\ram[5][7] ) );
  LATCHX1_HVT \ram_reg[5][6]  ( .CLK(n237), .D(N22), .Q(\ram[5][6] ) );
  LATCHX1_HVT \ram_reg[5][5]  ( .CLK(n236), .D(N21), .Q(\ram[5][5] ) );
  LATCHX1_HVT \ram_reg[5][4]  ( .CLK(n236), .D(N20), .Q(\ram[5][4] ) );
  LATCHX1_HVT \ram_reg[5][3]  ( .CLK(n235), .D(N19), .Q(\ram[5][3] ) );
  LATCHX1_HVT \ram_reg[5][2]  ( .CLK(n236), .D(N18), .Q(\ram[5][2] ) );
  LATCHX1_HVT \ram_reg[5][1]  ( .CLK(n237), .D(N17), .Q(\ram[5][1] ) );
  LATCHX1_HVT \ram_reg[5][0]  ( .CLK(n241), .D(N16), .Q(\ram[5][0] ) );
  LATCHX1_HVT \ram_reg[4][255]  ( .CLK(N285), .D(N273), .Q(\ram[4][255] ) );
  LATCHX1_HVT \ram_reg[4][254]  ( .CLK(N285), .D(N272), .Q(\ram[4][254] ) );
  LATCHX1_HVT \ram_reg[4][253]  ( .CLK(N285), .D(N271), .Q(\ram[4][253] ) );
  LATCHX1_HVT \ram_reg[4][252]  ( .CLK(N285), .D(N270), .Q(\ram[4][252] ) );
  LATCHX1_HVT \ram_reg[4][251]  ( .CLK(n274), .D(N269), .Q(\ram[4][251] ) );
  LATCHX1_HVT \ram_reg[4][250]  ( .CLK(n266), .D(N268), .Q(\ram[4][250] ) );
  LATCHX1_HVT \ram_reg[4][249]  ( .CLK(n266), .D(N267), .Q(\ram[4][249] ) );
  LATCHX1_HVT \ram_reg[4][248]  ( .CLK(n266), .D(N266), .Q(\ram[4][248] ) );
  LATCHX1_HVT \ram_reg[4][247]  ( .CLK(n266), .D(N265), .Q(\ram[4][247] ) );
  LATCHX1_HVT \ram_reg[4][246]  ( .CLK(n266), .D(N264), .Q(\ram[4][246] ) );
  LATCHX1_HVT \ram_reg[4][245]  ( .CLK(n266), .D(N263), .Q(\ram[4][245] ) );
  LATCHX1_HVT \ram_reg[4][244]  ( .CLK(n266), .D(N262), .Q(\ram[4][244] ) );
  LATCHX1_HVT \ram_reg[4][243]  ( .CLK(n266), .D(N261), .Q(\ram[4][243] ) );
  LATCHX1_HVT \ram_reg[4][242]  ( .CLK(n266), .D(N260), .Q(\ram[4][242] ) );
  LATCHX1_HVT \ram_reg[4][241]  ( .CLK(n265), .D(N259), .Q(\ram[4][241] ) );
  LATCHX1_HVT \ram_reg[4][240]  ( .CLK(n265), .D(N258), .Q(\ram[4][240] ) );
  LATCHX1_HVT \ram_reg[4][239]  ( .CLK(n265), .D(N257), .Q(\ram[4][239] ) );
  LATCHX1_HVT \ram_reg[4][238]  ( .CLK(n265), .D(N256), .Q(\ram[4][238] ) );
  LATCHX1_HVT \ram_reg[4][237]  ( .CLK(n265), .D(N255), .Q(\ram[4][237] ) );
  LATCHX1_HVT \ram_reg[4][236]  ( .CLK(n265), .D(N254), .Q(\ram[4][236] ) );
  LATCHX1_HVT \ram_reg[4][235]  ( .CLK(n265), .D(N253), .Q(\ram[4][235] ) );
  LATCHX1_HVT \ram_reg[4][234]  ( .CLK(n265), .D(N252), .Q(\ram[4][234] ) );
  LATCHX1_HVT \ram_reg[4][233]  ( .CLK(n265), .D(N251), .Q(\ram[4][233] ) );
  LATCHX1_HVT \ram_reg[4][232]  ( .CLK(n265), .D(N250), .Q(\ram[4][232] ) );
  LATCHX1_HVT \ram_reg[4][231]  ( .CLK(n265), .D(N249), .Q(\ram[4][231] ) );
  LATCHX1_HVT \ram_reg[4][230]  ( .CLK(n264), .D(N248), .Q(\ram[4][230] ) );
  LATCHX1_HVT \ram_reg[4][229]  ( .CLK(n264), .D(N247), .Q(\ram[4][229] ) );
  LATCHX1_HVT \ram_reg[4][228]  ( .CLK(n264), .D(N246), .Q(\ram[4][228] ) );
  LATCHX1_HVT \ram_reg[4][227]  ( .CLK(n274), .D(N245), .Q(\ram[4][227] ) );
  LATCHX1_HVT \ram_reg[4][226]  ( .CLK(n274), .D(N244), .Q(\ram[4][226] ) );
  LATCHX1_HVT \ram_reg[4][225]  ( .CLK(n274), .D(N243), .Q(\ram[4][225] ) );
  LATCHX1_HVT \ram_reg[4][224]  ( .CLK(n274), .D(N242), .Q(\ram[4][224] ) );
  LATCHX1_HVT \ram_reg[4][223]  ( .CLK(n274), .D(N241), .Q(\ram[4][223] ) );
  LATCHX1_HVT \ram_reg[4][222]  ( .CLK(n274), .D(N240), .Q(\ram[4][222] ) );
  LATCHX1_HVT \ram_reg[4][221]  ( .CLK(n274), .D(N239), .Q(\ram[4][221] ) );
  LATCHX1_HVT \ram_reg[4][220]  ( .CLK(n274), .D(N238), .Q(\ram[4][220] ) );
  LATCHX1_HVT \ram_reg[4][219]  ( .CLK(n274), .D(N237), .Q(\ram[4][219] ) );
  LATCHX1_HVT \ram_reg[4][218]  ( .CLK(n274), .D(N236), .Q(\ram[4][218] ) );
  LATCHX1_HVT \ram_reg[4][217]  ( .CLK(n273), .D(N235), .Q(\ram[4][217] ) );
  LATCHX1_HVT \ram_reg[4][216]  ( .CLK(n273), .D(N234), .Q(\ram[4][216] ) );
  LATCHX1_HVT \ram_reg[4][215]  ( .CLK(n273), .D(N233), .Q(\ram[4][215] ) );
  LATCHX1_HVT \ram_reg[4][214]  ( .CLK(n273), .D(N232), .Q(\ram[4][214] ) );
  LATCHX1_HVT \ram_reg[4][213]  ( .CLK(n273), .D(N231), .Q(\ram[4][213] ) );
  LATCHX1_HVT \ram_reg[4][212]  ( .CLK(n273), .D(N230), .Q(\ram[4][212] ) );
  LATCHX1_HVT \ram_reg[4][211]  ( .CLK(n273), .D(N229), .Q(\ram[4][211] ) );
  LATCHX1_HVT \ram_reg[4][210]  ( .CLK(n273), .D(N228), .Q(\ram[4][210] ) );
  LATCHX1_HVT \ram_reg[4][209]  ( .CLK(n273), .D(N227), .Q(\ram[4][209] ) );
  LATCHX1_HVT \ram_reg[4][208]  ( .CLK(n273), .D(N226), .Q(\ram[4][208] ) );
  LATCHX1_HVT \ram_reg[4][207]  ( .CLK(n272), .D(N225), .Q(\ram[4][207] ) );
  LATCHX1_HVT \ram_reg[4][206]  ( .CLK(n272), .D(N224), .Q(\ram[4][206] ) );
  LATCHX1_HVT \ram_reg[4][205]  ( .CLK(n272), .D(N223), .Q(\ram[4][205] ) );
  LATCHX1_HVT \ram_reg[4][204]  ( .CLK(n272), .D(N222), .Q(\ram[4][204] ) );
  LATCHX1_HVT \ram_reg[4][203]  ( .CLK(n272), .D(N221), .Q(\ram[4][203] ) );
  LATCHX1_HVT \ram_reg[4][202]  ( .CLK(n272), .D(N220), .Q(\ram[4][202] ) );
  LATCHX1_HVT \ram_reg[4][201]  ( .CLK(n272), .D(N219), .Q(\ram[4][201] ) );
  LATCHX1_HVT \ram_reg[4][200]  ( .CLK(n272), .D(N218), .Q(\ram[4][200] ) );
  LATCHX1_HVT \ram_reg[4][199]  ( .CLK(n272), .D(N217), .Q(\ram[4][199] ) );
  LATCHX1_HVT \ram_reg[4][198]  ( .CLK(n272), .D(N216), .Q(\ram[4][198] ) );
  LATCHX1_HVT \ram_reg[4][197]  ( .CLK(n272), .D(N214), .Q(\ram[4][197] ) );
  LATCHX1_HVT \ram_reg[4][196]  ( .CLK(n271), .D(N213), .Q(\ram[4][196] ) );
  LATCHX1_HVT \ram_reg[4][195]  ( .CLK(n271), .D(N212), .Q(\ram[4][195] ) );
  LATCHX1_HVT \ram_reg[4][194]  ( .CLK(n271), .D(N211), .Q(\ram[4][194] ) );
  LATCHX1_HVT \ram_reg[4][193]  ( .CLK(n271), .D(N210), .Q(\ram[4][193] ) );
  LATCHX1_HVT \ram_reg[4][192]  ( .CLK(n271), .D(N209), .Q(\ram[4][192] ) );
  LATCHX1_HVT \ram_reg[4][191]  ( .CLK(n271), .D(N208), .Q(\ram[4][191] ) );
  LATCHX1_HVT \ram_reg[4][190]  ( .CLK(n271), .D(N207), .Q(\ram[4][190] ) );
  LATCHX1_HVT \ram_reg[4][189]  ( .CLK(n271), .D(N206), .Q(\ram[4][189] ) );
  LATCHX1_HVT \ram_reg[4][188]  ( .CLK(n271), .D(N205), .Q(\ram[4][188] ) );
  LATCHX1_HVT \ram_reg[4][187]  ( .CLK(n271), .D(N204), .Q(\ram[4][187] ) );
  LATCHX1_HVT \ram_reg[4][186]  ( .CLK(n271), .D(N203), .Q(\ram[4][186] ) );
  LATCHX1_HVT \ram_reg[4][185]  ( .CLK(n270), .D(N202), .Q(\ram[4][185] ) );
  LATCHX1_HVT \ram_reg[4][184]  ( .CLK(n270), .D(N201), .Q(\ram[4][184] ) );
  LATCHX1_HVT \ram_reg[4][183]  ( .CLK(n270), .D(N200), .Q(\ram[4][183] ) );
  LATCHX1_HVT \ram_reg[4][182]  ( .CLK(n270), .D(N199), .Q(\ram[4][182] ) );
  LATCHX1_HVT \ram_reg[4][181]  ( .CLK(n270), .D(N198), .Q(\ram[4][181] ) );
  LATCHX1_HVT \ram_reg[4][180]  ( .CLK(n270), .D(N197), .Q(\ram[4][180] ) );
  LATCHX1_HVT \ram_reg[4][179]  ( .CLK(n270), .D(N196), .Q(\ram[4][179] ) );
  LATCHX1_HVT \ram_reg[4][178]  ( .CLK(n270), .D(N195), .Q(\ram[4][178] ) );
  LATCHX1_HVT \ram_reg[4][177]  ( .CLK(n270), .D(N194), .Q(\ram[4][177] ) );
  LATCHX1_HVT \ram_reg[4][176]  ( .CLK(n270), .D(N193), .Q(\ram[4][176] ) );
  LATCHX1_HVT \ram_reg[4][175]  ( .CLK(n270), .D(N192), .Q(\ram[4][175] ) );
  LATCHX1_HVT \ram_reg[4][174]  ( .CLK(n269), .D(N191), .Q(\ram[4][174] ) );
  LATCHX1_HVT \ram_reg[4][173]  ( .CLK(n269), .D(N190), .Q(\ram[4][173] ) );
  LATCHX1_HVT \ram_reg[4][172]  ( .CLK(n269), .D(N189), .Q(\ram[4][172] ) );
  LATCHX1_HVT \ram_reg[4][171]  ( .CLK(n269), .D(N188), .Q(\ram[4][171] ) );
  LATCHX1_HVT \ram_reg[4][170]  ( .CLK(n269), .D(N187), .Q(\ram[4][170] ) );
  LATCHX1_HVT \ram_reg[4][169]  ( .CLK(n269), .D(N186), .Q(\ram[4][169] ) );
  LATCHX1_HVT \ram_reg[4][168]  ( .CLK(n269), .D(N185), .Q(\ram[4][168] ) );
  LATCHX1_HVT \ram_reg[4][167]  ( .CLK(n269), .D(N184), .Q(\ram[4][167] ) );
  LATCHX1_HVT \ram_reg[4][166]  ( .CLK(n269), .D(N183), .Q(\ram[4][166] ) );
  LATCHX1_HVT \ram_reg[4][165]  ( .CLK(n269), .D(N182), .Q(\ram[4][165] ) );
  LATCHX1_HVT \ram_reg[4][164]  ( .CLK(n269), .D(N181), .Q(\ram[4][164] ) );
  LATCHX1_HVT \ram_reg[4][163]  ( .CLK(n268), .D(N180), .Q(\ram[4][163] ) );
  LATCHX1_HVT \ram_reg[4][162]  ( .CLK(n268), .D(N179), .Q(\ram[4][162] ) );
  LATCHX1_HVT \ram_reg[4][161]  ( .CLK(n268), .D(N178), .Q(\ram[4][161] ) );
  LATCHX1_HVT \ram_reg[4][160]  ( .CLK(n268), .D(N177), .Q(\ram[4][160] ) );
  LATCHX1_HVT \ram_reg[4][159]  ( .CLK(n268), .D(N176), .Q(\ram[4][159] ) );
  LATCHX1_HVT \ram_reg[4][158]  ( .CLK(n268), .D(N175), .Q(\ram[4][158] ) );
  LATCHX1_HVT \ram_reg[4][157]  ( .CLK(n268), .D(N174), .Q(\ram[4][157] ) );
  LATCHX1_HVT \ram_reg[4][156]  ( .CLK(n268), .D(N173), .Q(\ram[4][156] ) );
  LATCHX1_HVT \ram_reg[4][155]  ( .CLK(n268), .D(N172), .Q(\ram[4][155] ) );
  LATCHX1_HVT \ram_reg[4][154]  ( .CLK(n268), .D(N171), .Q(\ram[4][154] ) );
  LATCHX1_HVT \ram_reg[4][153]  ( .CLK(n268), .D(N170), .Q(\ram[4][153] ) );
  LATCHX1_HVT \ram_reg[4][152]  ( .CLK(n267), .D(N169), .Q(\ram[4][152] ) );
  LATCHX1_HVT \ram_reg[4][151]  ( .CLK(n267), .D(N168), .Q(\ram[4][151] ) );
  LATCHX1_HVT \ram_reg[4][150]  ( .CLK(n267), .D(N167), .Q(\ram[4][150] ) );
  LATCHX1_HVT \ram_reg[4][149]  ( .CLK(n267), .D(N166), .Q(\ram[4][149] ) );
  LATCHX1_HVT \ram_reg[4][148]  ( .CLK(n267), .D(N165), .Q(\ram[4][148] ) );
  LATCHX1_HVT \ram_reg[4][147]  ( .CLK(n267), .D(N164), .Q(\ram[4][147] ) );
  LATCHX1_HVT \ram_reg[4][146]  ( .CLK(n267), .D(N163), .Q(\ram[4][146] ) );
  LATCHX1_HVT \ram_reg[4][145]  ( .CLK(n267), .D(N162), .Q(\ram[4][145] ) );
  LATCHX1_HVT \ram_reg[4][144]  ( .CLK(n267), .D(N161), .Q(\ram[4][144] ) );
  LATCHX1_HVT \ram_reg[4][143]  ( .CLK(n267), .D(N160), .Q(\ram[4][143] ) );
  LATCHX1_HVT \ram_reg[4][142]  ( .CLK(n267), .D(N159), .Q(\ram[4][142] ) );
  LATCHX1_HVT \ram_reg[4][141]  ( .CLK(n266), .D(N158), .Q(\ram[4][141] ) );
  LATCHX1_HVT \ram_reg[4][140]  ( .CLK(n266), .D(N157), .Q(\ram[4][140] ) );
  LATCHX1_HVT \ram_reg[4][139]  ( .CLK(n266), .D(N156), .Q(\ram[4][139] ) );
  LATCHX1_HVT \ram_reg[4][138]  ( .CLK(n265), .D(N155), .Q(\ram[4][138] ) );
  LATCHX1_HVT \ram_reg[4][137]  ( .CLK(n274), .D(N154), .Q(\ram[4][137] ) );
  LATCHX1_HVT \ram_reg[4][136]  ( .CLK(n273), .D(N153), .Q(\ram[4][136] ) );
  LATCHX1_HVT \ram_reg[4][135]  ( .CLK(n273), .D(N152), .Q(\ram[4][135] ) );
  LATCHX1_HVT \ram_reg[4][134]  ( .CLK(n272), .D(N151), .Q(\ram[4][134] ) );
  LATCHX1_HVT \ram_reg[4][133]  ( .CLK(n271), .D(N150), .Q(\ram[4][133] ) );
  LATCHX1_HVT \ram_reg[4][132]  ( .CLK(n270), .D(N149), .Q(\ram[4][132] ) );
  LATCHX1_HVT \ram_reg[4][131]  ( .CLK(n269), .D(N148), .Q(\ram[4][131] ) );
  LATCHX1_HVT \ram_reg[4][130]  ( .CLK(n268), .D(N147), .Q(\ram[4][130] ) );
  LATCHX1_HVT \ram_reg[4][129]  ( .CLK(n267), .D(N146), .Q(\ram[4][129] ) );
  LATCHX1_HVT \ram_reg[4][128]  ( .CLK(n264), .D(N145), .Q(\ram[4][128] ) );
  LATCHX1_HVT \ram_reg[4][127]  ( .CLK(n255), .D(N144), .Q(\ram[4][127] ) );
  LATCHX1_HVT \ram_reg[4][126]  ( .CLK(n255), .D(N143), .Q(\ram[4][126] ) );
  LATCHX1_HVT \ram_reg[4][125]  ( .CLK(n255), .D(N142), .Q(\ram[4][125] ) );
  LATCHX1_HVT \ram_reg[4][124]  ( .CLK(n255), .D(N141), .Q(\ram[4][124] ) );
  LATCHX1_HVT \ram_reg[4][123]  ( .CLK(n255), .D(N140), .Q(\ram[4][123] ) );
  LATCHX1_HVT \ram_reg[4][122]  ( .CLK(n254), .D(N139), .Q(\ram[4][122] ) );
  LATCHX1_HVT \ram_reg[4][121]  ( .CLK(n255), .D(N138), .Q(\ram[4][121] ) );
  LATCHX1_HVT \ram_reg[4][120]  ( .CLK(n255), .D(N137), .Q(\ram[4][120] ) );
  LATCHX1_HVT \ram_reg[4][119]  ( .CLK(n264), .D(N136), .Q(\ram[4][119] ) );
  LATCHX1_HVT \ram_reg[4][118]  ( .CLK(n263), .D(N135), .Q(\ram[4][118] ) );
  LATCHX1_HVT \ram_reg[4][117]  ( .CLK(n263), .D(N134), .Q(\ram[4][117] ) );
  LATCHX1_HVT \ram_reg[4][116]  ( .CLK(n262), .D(N133), .Q(\ram[4][116] ) );
  LATCHX1_HVT \ram_reg[4][115]  ( .CLK(n257), .D(N132), .Q(\ram[4][115] ) );
  LATCHX1_HVT \ram_reg[4][114]  ( .CLK(n262), .D(N131), .Q(\ram[4][114] ) );
  LATCHX1_HVT \ram_reg[4][113]  ( .CLK(n262), .D(N130), .Q(\ram[4][113] ) );
  LATCHX1_HVT \ram_reg[4][112]  ( .CLK(n263), .D(N129), .Q(\ram[4][112] ) );
  LATCHX1_HVT \ram_reg[4][111]  ( .CLK(n261), .D(N128), .Q(\ram[4][111] ) );
  LATCHX1_HVT \ram_reg[4][110]  ( .CLK(n261), .D(N127), .Q(\ram[4][110] ) );
  LATCHX1_HVT \ram_reg[4][109]  ( .CLK(n261), .D(N126), .Q(\ram[4][109] ) );
  LATCHX1_HVT \ram_reg[4][108]  ( .CLK(n258), .D(N125), .Q(\ram[4][108] ) );
  LATCHX1_HVT \ram_reg[4][107]  ( .CLK(n255), .D(N124), .Q(\ram[4][107] ) );
  LATCHX1_HVT \ram_reg[4][106]  ( .CLK(n261), .D(N123), .Q(\ram[4][106] ) );
  LATCHX1_HVT \ram_reg[4][105]  ( .CLK(n261), .D(N122), .Q(\ram[4][105] ) );
  LATCHX1_HVT \ram_reg[4][104]  ( .CLK(n261), .D(N121), .Q(\ram[4][104] ) );
  LATCHX1_HVT \ram_reg[4][103]  ( .CLK(n260), .D(N120), .Q(\ram[4][103] ) );
  LATCHX1_HVT \ram_reg[4][102]  ( .CLK(n259), .D(N119), .Q(\ram[4][102] ) );
  LATCHX1_HVT \ram_reg[4][101]  ( .CLK(n259), .D(N118), .Q(\ram[4][101] ) );
  LATCHX1_HVT \ram_reg[4][100]  ( .CLK(n260), .D(N117), .Q(\ram[4][100] ) );
  LATCHX1_HVT \ram_reg[4][99]  ( .CLK(n258), .D(N116), .Q(\ram[4][99] ) );
  LATCHX1_HVT \ram_reg[4][98]  ( .CLK(n259), .D(N114), .Q(\ram[4][98] ) );
  LATCHX1_HVT \ram_reg[4][97]  ( .CLK(n260), .D(N113), .Q(\ram[4][97] ) );
  LATCHX1_HVT \ram_reg[4][96]  ( .CLK(n264), .D(N112), .Q(\ram[4][96] ) );
  LATCHX1_HVT \ram_reg[4][95]  ( .CLK(n256), .D(N111), .Q(\ram[4][95] ) );
  LATCHX1_HVT \ram_reg[4][94]  ( .CLK(n256), .D(N110), .Q(\ram[4][94] ) );
  LATCHX1_HVT \ram_reg[4][93]  ( .CLK(n256), .D(N109), .Q(\ram[4][93] ) );
  LATCHX1_HVT \ram_reg[4][92]  ( .CLK(n255), .D(N108), .Q(\ram[4][92] ) );
  LATCHX1_HVT \ram_reg[4][91]  ( .CLK(n255), .D(N107), .Q(\ram[4][91] ) );
  LATCHX1_HVT \ram_reg[4][90]  ( .CLK(n256), .D(N106), .Q(\ram[4][90] ) );
  LATCHX1_HVT \ram_reg[4][89]  ( .CLK(n255), .D(N105), .Q(\ram[4][89] ) );
  LATCHX1_HVT \ram_reg[4][88]  ( .CLK(n256), .D(N104), .Q(\ram[4][88] ) );
  LATCHX1_HVT \ram_reg[4][87]  ( .CLK(n264), .D(N103), .Q(\ram[4][87] ) );
  LATCHX1_HVT \ram_reg[4][86]  ( .CLK(n263), .D(N102), .Q(\ram[4][86] ) );
  LATCHX1_HVT \ram_reg[4][85]  ( .CLK(n262), .D(N101), .Q(\ram[4][85] ) );
  LATCHX1_HVT \ram_reg[4][84]  ( .CLK(n262), .D(N100), .Q(\ram[4][84] ) );
  LATCHX1_HVT \ram_reg[4][83]  ( .CLK(n257), .D(N99), .Q(\ram[4][83] ) );
  LATCHX1_HVT \ram_reg[4][82]  ( .CLK(n263), .D(N98), .Q(\ram[4][82] ) );
  LATCHX1_HVT \ram_reg[4][81]  ( .CLK(n262), .D(N97), .Q(\ram[4][81] ) );
  LATCHX1_HVT \ram_reg[4][80]  ( .CLK(n263), .D(N96), .Q(\ram[4][80] ) );
  LATCHX1_HVT \ram_reg[4][79]  ( .CLK(n257), .D(N95), .Q(\ram[4][79] ) );
  LATCHX1_HVT \ram_reg[4][78]  ( .CLK(n256), .D(N94), .Q(\ram[4][78] ) );
  LATCHX1_HVT \ram_reg[4][77]  ( .CLK(n257), .D(N93), .Q(\ram[4][77] ) );
  LATCHX1_HVT \ram_reg[4][76]  ( .CLK(n256), .D(N92), .Q(\ram[4][76] ) );
  LATCHX1_HVT \ram_reg[4][75]  ( .CLK(n256), .D(N91), .Q(\ram[4][75] ) );
  LATCHX1_HVT \ram_reg[4][74]  ( .CLK(n254), .D(N90), .Q(\ram[4][74] ) );
  LATCHX1_HVT \ram_reg[4][73]  ( .CLK(n257), .D(N89), .Q(\ram[4][73] ) );
  LATCHX1_HVT \ram_reg[4][72]  ( .CLK(n257), .D(N88), .Q(\ram[4][72] ) );
  LATCHX1_HVT \ram_reg[4][71]  ( .CLK(n260), .D(N87), .Q(\ram[4][71] ) );
  LATCHX1_HVT \ram_reg[4][70]  ( .CLK(n260), .D(N86), .Q(\ram[4][70] ) );
  LATCHX1_HVT \ram_reg[4][69]  ( .CLK(n259), .D(N85), .Q(\ram[4][69] ) );
  LATCHX1_HVT \ram_reg[4][68]  ( .CLK(n260), .D(N84), .Q(\ram[4][68] ) );
  LATCHX1_HVT \ram_reg[4][67]  ( .CLK(n259), .D(N83), .Q(\ram[4][67] ) );
  LATCHX1_HVT \ram_reg[4][66]  ( .CLK(n258), .D(N82), .Q(\ram[4][66] ) );
  LATCHX1_HVT \ram_reg[4][65]  ( .CLK(n259), .D(N81), .Q(\ram[4][65] ) );
  LATCHX1_HVT \ram_reg[4][64]  ( .CLK(n264), .D(N80), .Q(\ram[4][64] ) );
  LATCHX1_HVT \ram_reg[4][63]  ( .CLK(n258), .D(N79), .Q(\ram[4][63] ) );
  LATCHX1_HVT \ram_reg[4][62]  ( .CLK(n258), .D(N78), .Q(\ram[4][62] ) );
  LATCHX1_HVT \ram_reg[4][61]  ( .CLK(n258), .D(N77), .Q(\ram[4][61] ) );
  LATCHX1_HVT \ram_reg[4][60]  ( .CLK(n258), .D(N76), .Q(\ram[4][60] ) );
  LATCHX1_HVT \ram_reg[4][59]  ( .CLK(n258), .D(N75), .Q(\ram[4][59] ) );
  LATCHX1_HVT \ram_reg[4][58]  ( .CLK(n257), .D(N74), .Q(\ram[4][58] ) );
  LATCHX1_HVT \ram_reg[4][57]  ( .CLK(n258), .D(N73), .Q(\ram[4][57] ) );
  LATCHX1_HVT \ram_reg[4][56]  ( .CLK(n258), .D(N72), .Q(\ram[4][56] ) );
  LATCHX1_HVT \ram_reg[4][55]  ( .CLK(n264), .D(N71), .Q(\ram[4][55] ) );
  LATCHX1_HVT \ram_reg[4][54]  ( .CLK(n262), .D(N70), .Q(\ram[4][54] ) );
  LATCHX1_HVT \ram_reg[4][53]  ( .CLK(n262), .D(N69), .Q(\ram[4][53] ) );
  LATCHX1_HVT \ram_reg[4][52]  ( .CLK(n263), .D(N68), .Q(\ram[4][52] ) );
  LATCHX1_HVT \ram_reg[4][51]  ( .CLK(n257), .D(N67), .Q(\ram[4][51] ) );
  LATCHX1_HVT \ram_reg[4][50]  ( .CLK(n254), .D(N66), .Q(\ram[4][50] ) );
  LATCHX1_HVT \ram_reg[4][49]  ( .CLK(n263), .D(N65), .Q(\ram[4][49] ) );
  LATCHX1_HVT \ram_reg[4][48]  ( .CLK(n263), .D(N64), .Q(\ram[4][48] ) );
  LATCHX1_HVT \ram_reg[4][47]  ( .CLK(n261), .D(N63), .Q(\ram[4][47] ) );
  LATCHX1_HVT \ram_reg[4][46]  ( .CLK(n261), .D(N62), .Q(\ram[4][46] ) );
  LATCHX1_HVT \ram_reg[4][45]  ( .CLK(n261), .D(N61), .Q(\ram[4][45] ) );
  LATCHX1_HVT \ram_reg[4][44]  ( .CLK(n261), .D(N60), .Q(\ram[4][44] ) );
  LATCHX1_HVT \ram_reg[4][43]  ( .CLK(n258), .D(N59), .Q(\ram[4][43] ) );
  LATCHX1_HVT \ram_reg[4][42]  ( .CLK(n262), .D(N58), .Q(\ram[4][42] ) );
  LATCHX1_HVT \ram_reg[4][41]  ( .CLK(n255), .D(N57), .Q(\ram[4][41] ) );
  LATCHX1_HVT \ram_reg[4][40]  ( .CLK(n261), .D(N56), .Q(\ram[4][40] ) );
  LATCHX1_HVT \ram_reg[4][39]  ( .CLK(n260), .D(N55), .Q(\ram[4][39] ) );
  LATCHX1_HVT \ram_reg[4][38]  ( .CLK(n260), .D(N54), .Q(\ram[4][38] ) );
  LATCHX1_HVT \ram_reg[4][37]  ( .CLK(n259), .D(N53), .Q(\ram[4][37] ) );
  LATCHX1_HVT \ram_reg[4][36]  ( .CLK(n259), .D(N52), .Q(\ram[4][36] ) );
  LATCHX1_HVT \ram_reg[4][35]  ( .CLK(n259), .D(N51), .Q(\ram[4][35] ) );
  LATCHX1_HVT \ram_reg[4][34]  ( .CLK(n261), .D(N50), .Q(\ram[4][34] ) );
  LATCHX1_HVT \ram_reg[4][33]  ( .CLK(n260), .D(N49), .Q(\ram[4][33] ) );
  LATCHX1_HVT \ram_reg[4][32]  ( .CLK(n264), .D(N48), .Q(\ram[4][32] ) );
  LATCHX1_HVT \ram_reg[4][31]  ( .CLK(n254), .D(N47), .Q(\ram[4][31] ) );
  LATCHX1_HVT \ram_reg[4][30]  ( .CLK(n254), .D(N46), .Q(\ram[4][30] ) );
  LATCHX1_HVT \ram_reg[4][29]  ( .CLK(n254), .D(N45), .Q(\ram[4][29] ) );
  LATCHX1_HVT \ram_reg[4][28]  ( .CLK(n254), .D(N44), .Q(\ram[4][28] ) );
  LATCHX1_HVT \ram_reg[4][27]  ( .CLK(n254), .D(N43), .Q(\ram[4][27] ) );
  LATCHX1_HVT \ram_reg[4][26]  ( .CLK(n254), .D(N42), .Q(\ram[4][26] ) );
  LATCHX1_HVT \ram_reg[4][25]  ( .CLK(n254), .D(N41), .Q(\ram[4][25] ) );
  LATCHX1_HVT \ram_reg[4][24]  ( .CLK(n254), .D(N40), .Q(\ram[4][24] ) );
  LATCHX1_HVT \ram_reg[4][23]  ( .CLK(n264), .D(N39), .Q(\ram[4][23] ) );
  LATCHX1_HVT \ram_reg[4][22]  ( .CLK(n263), .D(N38), .Q(\ram[4][22] ) );
  LATCHX1_HVT \ram_reg[4][21]  ( .CLK(n262), .D(N37), .Q(\ram[4][21] ) );
  LATCHX1_HVT \ram_reg[4][20]  ( .CLK(n262), .D(N36), .Q(\ram[4][20] ) );
  LATCHX1_HVT \ram_reg[4][19]  ( .CLK(n254), .D(N35), .Q(\ram[4][19] ) );
  LATCHX1_HVT \ram_reg[4][18]  ( .CLK(n262), .D(N34), .Q(\ram[4][18] ) );
  LATCHX1_HVT \ram_reg[4][17]  ( .CLK(n263), .D(N33), .Q(\ram[4][17] ) );
  LATCHX1_HVT \ram_reg[4][16]  ( .CLK(n263), .D(N32), .Q(\ram[4][16] ) );
  LATCHX1_HVT \ram_reg[4][15]  ( .CLK(n257), .D(N31), .Q(\ram[4][15] ) );
  LATCHX1_HVT \ram_reg[4][14]  ( .CLK(n257), .D(N30), .Q(\ram[4][14] ) );
  LATCHX1_HVT \ram_reg[4][13]  ( .CLK(n256), .D(N29), .Q(\ram[4][13] ) );
  LATCHX1_HVT \ram_reg[4][12]  ( .CLK(n256), .D(N28), .Q(\ram[4][12] ) );
  LATCHX1_HVT \ram_reg[4][11]  ( .CLK(n257), .D(N27), .Q(\ram[4][11] ) );
  LATCHX1_HVT \ram_reg[4][10]  ( .CLK(n256), .D(N26), .Q(\ram[4][10] ) );
  LATCHX1_HVT \ram_reg[4][9]  ( .CLK(n256), .D(N25), .Q(\ram[4][9] ) );
  LATCHX1_HVT \ram_reg[4][8]  ( .CLK(n257), .D(N24), .Q(\ram[4][8] ) );
  LATCHX1_HVT \ram_reg[4][7]  ( .CLK(n260), .D(N23), .Q(\ram[4][7] ) );
  LATCHX1_HVT \ram_reg[4][6]  ( .CLK(n260), .D(N22), .Q(\ram[4][6] ) );
  LATCHX1_HVT \ram_reg[4][5]  ( .CLK(n259), .D(N21), .Q(\ram[4][5] ) );
  LATCHX1_HVT \ram_reg[4][4]  ( .CLK(n259), .D(N20), .Q(\ram[4][4] ) );
  LATCHX1_HVT \ram_reg[4][3]  ( .CLK(n258), .D(N19), .Q(\ram[4][3] ) );
  LATCHX1_HVT \ram_reg[4][2]  ( .CLK(n259), .D(N18), .Q(\ram[4][2] ) );
  LATCHX1_HVT \ram_reg[4][1]  ( .CLK(n260), .D(N17), .Q(\ram[4][1] ) );
  LATCHX1_HVT \ram_reg[4][0]  ( .CLK(n264), .D(N16), .Q(\ram[4][0] ) );
  LATCHX1_HVT \ram_reg[3][255]  ( .CLK(N282), .D(N273), .Q(\ram[3][255] ) );
  LATCHX1_HVT \ram_reg[3][254]  ( .CLK(N282), .D(N272), .Q(\ram[3][254] ) );
  LATCHX1_HVT \ram_reg[3][253]  ( .CLK(N282), .D(N271), .Q(\ram[3][253] ) );
  LATCHX1_HVT \ram_reg[3][252]  ( .CLK(N282), .D(N270), .Q(\ram[3][252] ) );
  LATCHX1_HVT \ram_reg[3][251]  ( .CLK(n297), .D(N269), .Q(\ram[3][251] ) );
  LATCHX1_HVT \ram_reg[3][250]  ( .CLK(n289), .D(N268), .Q(\ram[3][250] ) );
  LATCHX1_HVT \ram_reg[3][249]  ( .CLK(n289), .D(N267), .Q(\ram[3][249] ) );
  LATCHX1_HVT \ram_reg[3][248]  ( .CLK(n289), .D(N266), .Q(\ram[3][248] ) );
  LATCHX1_HVT \ram_reg[3][247]  ( .CLK(n289), .D(N265), .Q(\ram[3][247] ) );
  LATCHX1_HVT \ram_reg[3][246]  ( .CLK(n289), .D(N264), .Q(\ram[3][246] ) );
  LATCHX1_HVT \ram_reg[3][245]  ( .CLK(n289), .D(N263), .Q(\ram[3][245] ) );
  LATCHX1_HVT \ram_reg[3][244]  ( .CLK(n289), .D(N262), .Q(\ram[3][244] ) );
  LATCHX1_HVT \ram_reg[3][243]  ( .CLK(n289), .D(N261), .Q(\ram[3][243] ) );
  LATCHX1_HVT \ram_reg[3][242]  ( .CLK(n289), .D(N260), .Q(\ram[3][242] ) );
  LATCHX1_HVT \ram_reg[3][241]  ( .CLK(n288), .D(N259), .Q(\ram[3][241] ) );
  LATCHX1_HVT \ram_reg[3][240]  ( .CLK(n288), .D(N258), .Q(\ram[3][240] ) );
  LATCHX1_HVT \ram_reg[3][239]  ( .CLK(n288), .D(N257), .Q(\ram[3][239] ) );
  LATCHX1_HVT \ram_reg[3][238]  ( .CLK(n288), .D(N256), .Q(\ram[3][238] ) );
  LATCHX1_HVT \ram_reg[3][237]  ( .CLK(n288), .D(N255), .Q(\ram[3][237] ) );
  LATCHX1_HVT \ram_reg[3][236]  ( .CLK(n288), .D(N254), .Q(\ram[3][236] ) );
  LATCHX1_HVT \ram_reg[3][235]  ( .CLK(n288), .D(N253), .Q(\ram[3][235] ) );
  LATCHX1_HVT \ram_reg[3][234]  ( .CLK(n288), .D(N252), .Q(\ram[3][234] ) );
  LATCHX1_HVT \ram_reg[3][233]  ( .CLK(n288), .D(N251), .Q(\ram[3][233] ) );
  LATCHX1_HVT \ram_reg[3][232]  ( .CLK(n288), .D(N250), .Q(\ram[3][232] ) );
  LATCHX1_HVT \ram_reg[3][231]  ( .CLK(n288), .D(N249), .Q(\ram[3][231] ) );
  LATCHX1_HVT \ram_reg[3][230]  ( .CLK(n287), .D(N248), .Q(\ram[3][230] ) );
  LATCHX1_HVT \ram_reg[3][229]  ( .CLK(n287), .D(N247), .Q(\ram[3][229] ) );
  LATCHX1_HVT \ram_reg[3][228]  ( .CLK(n287), .D(N246), .Q(\ram[3][228] ) );
  LATCHX1_HVT \ram_reg[3][227]  ( .CLK(n297), .D(N245), .Q(\ram[3][227] ) );
  LATCHX1_HVT \ram_reg[3][226]  ( .CLK(n297), .D(N244), .Q(\ram[3][226] ) );
  LATCHX1_HVT \ram_reg[3][225]  ( .CLK(n297), .D(N243), .Q(\ram[3][225] ) );
  LATCHX1_HVT \ram_reg[3][224]  ( .CLK(n297), .D(N242), .Q(\ram[3][224] ) );
  LATCHX1_HVT \ram_reg[3][223]  ( .CLK(n297), .D(N241), .Q(\ram[3][223] ) );
  LATCHX1_HVT \ram_reg[3][222]  ( .CLK(n297), .D(N240), .Q(\ram[3][222] ) );
  LATCHX1_HVT \ram_reg[3][221]  ( .CLK(n297), .D(N239), .Q(\ram[3][221] ) );
  LATCHX1_HVT \ram_reg[3][220]  ( .CLK(n297), .D(N238), .Q(\ram[3][220] ) );
  LATCHX1_HVT \ram_reg[3][219]  ( .CLK(n297), .D(N237), .Q(\ram[3][219] ) );
  LATCHX1_HVT \ram_reg[3][218]  ( .CLK(n297), .D(N236), .Q(\ram[3][218] ) );
  LATCHX1_HVT \ram_reg[3][217]  ( .CLK(n296), .D(N235), .Q(\ram[3][217] ) );
  LATCHX1_HVT \ram_reg[3][216]  ( .CLK(n296), .D(N234), .Q(\ram[3][216] ) );
  LATCHX1_HVT \ram_reg[3][215]  ( .CLK(n296), .D(N233), .Q(\ram[3][215] ) );
  LATCHX1_HVT \ram_reg[3][214]  ( .CLK(n296), .D(N232), .Q(\ram[3][214] ) );
  LATCHX1_HVT \ram_reg[3][213]  ( .CLK(n296), .D(N231), .Q(\ram[3][213] ) );
  LATCHX1_HVT \ram_reg[3][212]  ( .CLK(n296), .D(N230), .Q(\ram[3][212] ) );
  LATCHX1_HVT \ram_reg[3][211]  ( .CLK(n296), .D(N229), .Q(\ram[3][211] ) );
  LATCHX1_HVT \ram_reg[3][210]  ( .CLK(n296), .D(N228), .Q(\ram[3][210] ) );
  LATCHX1_HVT \ram_reg[3][209]  ( .CLK(n296), .D(N227), .Q(\ram[3][209] ) );
  LATCHX1_HVT \ram_reg[3][208]  ( .CLK(n296), .D(N226), .Q(\ram[3][208] ) );
  LATCHX1_HVT \ram_reg[3][207]  ( .CLK(n295), .D(N225), .Q(\ram[3][207] ) );
  LATCHX1_HVT \ram_reg[3][206]  ( .CLK(n295), .D(N224), .Q(\ram[3][206] ) );
  LATCHX1_HVT \ram_reg[3][205]  ( .CLK(n295), .D(N223), .Q(\ram[3][205] ) );
  LATCHX1_HVT \ram_reg[3][204]  ( .CLK(n295), .D(N222), .Q(\ram[3][204] ) );
  LATCHX1_HVT \ram_reg[3][203]  ( .CLK(n295), .D(N221), .Q(\ram[3][203] ) );
  LATCHX1_HVT \ram_reg[3][202]  ( .CLK(n295), .D(N220), .Q(\ram[3][202] ) );
  LATCHX1_HVT \ram_reg[3][201]  ( .CLK(n295), .D(N219), .Q(\ram[3][201] ) );
  LATCHX1_HVT \ram_reg[3][200]  ( .CLK(n295), .D(N218), .Q(\ram[3][200] ) );
  LATCHX1_HVT \ram_reg[3][199]  ( .CLK(n295), .D(N217), .Q(\ram[3][199] ) );
  LATCHX1_HVT \ram_reg[3][198]  ( .CLK(n295), .D(N216), .Q(\ram[3][198] ) );
  LATCHX1_HVT \ram_reg[3][197]  ( .CLK(n295), .D(N214), .Q(\ram[3][197] ) );
  LATCHX1_HVT \ram_reg[3][196]  ( .CLK(n294), .D(N213), .Q(\ram[3][196] ) );
  LATCHX1_HVT \ram_reg[3][195]  ( .CLK(n294), .D(N212), .Q(\ram[3][195] ) );
  LATCHX1_HVT \ram_reg[3][194]  ( .CLK(n294), .D(N211), .Q(\ram[3][194] ) );
  LATCHX1_HVT \ram_reg[3][193]  ( .CLK(n294), .D(N210), .Q(\ram[3][193] ) );
  LATCHX1_HVT \ram_reg[3][192]  ( .CLK(n294), .D(N209), .Q(\ram[3][192] ) );
  LATCHX1_HVT \ram_reg[3][191]  ( .CLK(n294), .D(N208), .Q(\ram[3][191] ) );
  LATCHX1_HVT \ram_reg[3][190]  ( .CLK(n294), .D(N207), .Q(\ram[3][190] ) );
  LATCHX1_HVT \ram_reg[3][189]  ( .CLK(n294), .D(N206), .Q(\ram[3][189] ) );
  LATCHX1_HVT \ram_reg[3][188]  ( .CLK(n294), .D(N205), .Q(\ram[3][188] ) );
  LATCHX1_HVT \ram_reg[3][187]  ( .CLK(n294), .D(N204), .Q(\ram[3][187] ) );
  LATCHX1_HVT \ram_reg[3][186]  ( .CLK(n294), .D(N203), .Q(\ram[3][186] ) );
  LATCHX1_HVT \ram_reg[3][185]  ( .CLK(n293), .D(N202), .Q(\ram[3][185] ) );
  LATCHX1_HVT \ram_reg[3][184]  ( .CLK(n293), .D(N201), .Q(\ram[3][184] ) );
  LATCHX1_HVT \ram_reg[3][183]  ( .CLK(n293), .D(N200), .Q(\ram[3][183] ) );
  LATCHX1_HVT \ram_reg[3][182]  ( .CLK(n293), .D(N199), .Q(\ram[3][182] ) );
  LATCHX1_HVT \ram_reg[3][181]  ( .CLK(n293), .D(N198), .Q(\ram[3][181] ) );
  LATCHX1_HVT \ram_reg[3][180]  ( .CLK(n293), .D(N197), .Q(\ram[3][180] ) );
  LATCHX1_HVT \ram_reg[3][179]  ( .CLK(n293), .D(N196), .Q(\ram[3][179] ) );
  LATCHX1_HVT \ram_reg[3][178]  ( .CLK(n293), .D(N195), .Q(\ram[3][178] ) );
  LATCHX1_HVT \ram_reg[3][177]  ( .CLK(n293), .D(N194), .Q(\ram[3][177] ) );
  LATCHX1_HVT \ram_reg[3][176]  ( .CLK(n293), .D(N193), .Q(\ram[3][176] ) );
  LATCHX1_HVT \ram_reg[3][175]  ( .CLK(n293), .D(N192), .Q(\ram[3][175] ) );
  LATCHX1_HVT \ram_reg[3][174]  ( .CLK(n292), .D(N191), .Q(\ram[3][174] ) );
  LATCHX1_HVT \ram_reg[3][173]  ( .CLK(n292), .D(N190), .Q(\ram[3][173] ) );
  LATCHX1_HVT \ram_reg[3][172]  ( .CLK(n292), .D(N189), .Q(\ram[3][172] ) );
  LATCHX1_HVT \ram_reg[3][171]  ( .CLK(n292), .D(N188), .Q(\ram[3][171] ) );
  LATCHX1_HVT \ram_reg[3][170]  ( .CLK(n292), .D(N187), .Q(\ram[3][170] ) );
  LATCHX1_HVT \ram_reg[3][169]  ( .CLK(n292), .D(N186), .Q(\ram[3][169] ) );
  LATCHX1_HVT \ram_reg[3][168]  ( .CLK(n292), .D(N185), .Q(\ram[3][168] ) );
  LATCHX1_HVT \ram_reg[3][167]  ( .CLK(n292), .D(N184), .Q(\ram[3][167] ) );
  LATCHX1_HVT \ram_reg[3][166]  ( .CLK(n292), .D(N183), .Q(\ram[3][166] ) );
  LATCHX1_HVT \ram_reg[3][165]  ( .CLK(n292), .D(N182), .Q(\ram[3][165] ) );
  LATCHX1_HVT \ram_reg[3][164]  ( .CLK(n292), .D(N181), .Q(\ram[3][164] ) );
  LATCHX1_HVT \ram_reg[3][163]  ( .CLK(n291), .D(N180), .Q(\ram[3][163] ) );
  LATCHX1_HVT \ram_reg[3][162]  ( .CLK(n291), .D(N179), .Q(\ram[3][162] ) );
  LATCHX1_HVT \ram_reg[3][161]  ( .CLK(n291), .D(N178), .Q(\ram[3][161] ) );
  LATCHX1_HVT \ram_reg[3][160]  ( .CLK(n291), .D(N177), .Q(\ram[3][160] ) );
  LATCHX1_HVT \ram_reg[3][159]  ( .CLK(n291), .D(N176), .Q(\ram[3][159] ) );
  LATCHX1_HVT \ram_reg[3][158]  ( .CLK(n291), .D(N175), .Q(\ram[3][158] ) );
  LATCHX1_HVT \ram_reg[3][157]  ( .CLK(n291), .D(N174), .Q(\ram[3][157] ) );
  LATCHX1_HVT \ram_reg[3][156]  ( .CLK(n291), .D(N173), .Q(\ram[3][156] ) );
  LATCHX1_HVT \ram_reg[3][155]  ( .CLK(n291), .D(N172), .Q(\ram[3][155] ) );
  LATCHX1_HVT \ram_reg[3][154]  ( .CLK(n291), .D(N171), .Q(\ram[3][154] ) );
  LATCHX1_HVT \ram_reg[3][153]  ( .CLK(n291), .D(N170), .Q(\ram[3][153] ) );
  LATCHX1_HVT \ram_reg[3][152]  ( .CLK(n290), .D(N169), .Q(\ram[3][152] ) );
  LATCHX1_HVT \ram_reg[3][151]  ( .CLK(n290), .D(N168), .Q(\ram[3][151] ) );
  LATCHX1_HVT \ram_reg[3][150]  ( .CLK(n290), .D(N167), .Q(\ram[3][150] ) );
  LATCHX1_HVT \ram_reg[3][149]  ( .CLK(n290), .D(N166), .Q(\ram[3][149] ) );
  LATCHX1_HVT \ram_reg[3][148]  ( .CLK(n290), .D(N165), .Q(\ram[3][148] ) );
  LATCHX1_HVT \ram_reg[3][147]  ( .CLK(n290), .D(N164), .Q(\ram[3][147] ) );
  LATCHX1_HVT \ram_reg[3][146]  ( .CLK(n290), .D(N163), .Q(\ram[3][146] ) );
  LATCHX1_HVT \ram_reg[3][145]  ( .CLK(n290), .D(N162), .Q(\ram[3][145] ) );
  LATCHX1_HVT \ram_reg[3][144]  ( .CLK(n290), .D(N161), .Q(\ram[3][144] ) );
  LATCHX1_HVT \ram_reg[3][143]  ( .CLK(n290), .D(N160), .Q(\ram[3][143] ) );
  LATCHX1_HVT \ram_reg[3][142]  ( .CLK(n290), .D(N159), .Q(\ram[3][142] ) );
  LATCHX1_HVT \ram_reg[3][141]  ( .CLK(n289), .D(N158), .Q(\ram[3][141] ) );
  LATCHX1_HVT \ram_reg[3][140]  ( .CLK(n289), .D(N157), .Q(\ram[3][140] ) );
  LATCHX1_HVT \ram_reg[3][139]  ( .CLK(n289), .D(N156), .Q(\ram[3][139] ) );
  LATCHX1_HVT \ram_reg[3][138]  ( .CLK(n288), .D(N155), .Q(\ram[3][138] ) );
  LATCHX1_HVT \ram_reg[3][137]  ( .CLK(n297), .D(N154), .Q(\ram[3][137] ) );
  LATCHX1_HVT \ram_reg[3][136]  ( .CLK(n296), .D(N153), .Q(\ram[3][136] ) );
  LATCHX1_HVT \ram_reg[3][135]  ( .CLK(n296), .D(N152), .Q(\ram[3][135] ) );
  LATCHX1_HVT \ram_reg[3][134]  ( .CLK(n295), .D(N151), .Q(\ram[3][134] ) );
  LATCHX1_HVT \ram_reg[3][133]  ( .CLK(n294), .D(N150), .Q(\ram[3][133] ) );
  LATCHX1_HVT \ram_reg[3][132]  ( .CLK(n293), .D(N149), .Q(\ram[3][132] ) );
  LATCHX1_HVT \ram_reg[3][131]  ( .CLK(n292), .D(N148), .Q(\ram[3][131] ) );
  LATCHX1_HVT \ram_reg[3][130]  ( .CLK(n291), .D(N147), .Q(\ram[3][130] ) );
  LATCHX1_HVT \ram_reg[3][129]  ( .CLK(n290), .D(N146), .Q(\ram[3][129] ) );
  LATCHX1_HVT \ram_reg[3][128]  ( .CLK(n287), .D(N145), .Q(\ram[3][128] ) );
  LATCHX1_HVT \ram_reg[3][127]  ( .CLK(n278), .D(N144), .Q(\ram[3][127] ) );
  LATCHX1_HVT \ram_reg[3][126]  ( .CLK(n278), .D(N143), .Q(\ram[3][126] ) );
  LATCHX1_HVT \ram_reg[3][125]  ( .CLK(n278), .D(N142), .Q(\ram[3][125] ) );
  LATCHX1_HVT \ram_reg[3][124]  ( .CLK(n278), .D(N141), .Q(\ram[3][124] ) );
  LATCHX1_HVT \ram_reg[3][123]  ( .CLK(n278), .D(N140), .Q(\ram[3][123] ) );
  LATCHX1_HVT \ram_reg[3][122]  ( .CLK(n277), .D(N139), .Q(\ram[3][122] ) );
  LATCHX1_HVT \ram_reg[3][121]  ( .CLK(n278), .D(N138), .Q(\ram[3][121] ) );
  LATCHX1_HVT \ram_reg[3][120]  ( .CLK(n278), .D(N137), .Q(\ram[3][120] ) );
  LATCHX1_HVT \ram_reg[3][119]  ( .CLK(n287), .D(N136), .Q(\ram[3][119] ) );
  LATCHX1_HVT \ram_reg[3][118]  ( .CLK(n286), .D(N135), .Q(\ram[3][118] ) );
  LATCHX1_HVT \ram_reg[3][117]  ( .CLK(n286), .D(N134), .Q(\ram[3][117] ) );
  LATCHX1_HVT \ram_reg[3][116]  ( .CLK(n285), .D(N133), .Q(\ram[3][116] ) );
  LATCHX1_HVT \ram_reg[3][115]  ( .CLK(n280), .D(N132), .Q(\ram[3][115] ) );
  LATCHX1_HVT \ram_reg[3][114]  ( .CLK(n285), .D(N131), .Q(\ram[3][114] ) );
  LATCHX1_HVT \ram_reg[3][113]  ( .CLK(n285), .D(N130), .Q(\ram[3][113] ) );
  LATCHX1_HVT \ram_reg[3][112]  ( .CLK(n286), .D(N129), .Q(\ram[3][112] ) );
  LATCHX1_HVT \ram_reg[3][111]  ( .CLK(n284), .D(N128), .Q(\ram[3][111] ) );
  LATCHX1_HVT \ram_reg[3][110]  ( .CLK(n284), .D(N127), .Q(\ram[3][110] ) );
  LATCHX1_HVT \ram_reg[3][109]  ( .CLK(n284), .D(N126), .Q(\ram[3][109] ) );
  LATCHX1_HVT \ram_reg[3][108]  ( .CLK(n281), .D(N125), .Q(\ram[3][108] ) );
  LATCHX1_HVT \ram_reg[3][107]  ( .CLK(n278), .D(N124), .Q(\ram[3][107] ) );
  LATCHX1_HVT \ram_reg[3][106]  ( .CLK(n284), .D(N123), .Q(\ram[3][106] ) );
  LATCHX1_HVT \ram_reg[3][105]  ( .CLK(n284), .D(N122), .Q(\ram[3][105] ) );
  LATCHX1_HVT \ram_reg[3][104]  ( .CLK(n284), .D(N121), .Q(\ram[3][104] ) );
  LATCHX1_HVT \ram_reg[3][103]  ( .CLK(n283), .D(N120), .Q(\ram[3][103] ) );
  LATCHX1_HVT \ram_reg[3][102]  ( .CLK(n282), .D(N119), .Q(\ram[3][102] ) );
  LATCHX1_HVT \ram_reg[3][101]  ( .CLK(n282), .D(N118), .Q(\ram[3][101] ) );
  LATCHX1_HVT \ram_reg[3][100]  ( .CLK(n283), .D(N117), .Q(\ram[3][100] ) );
  LATCHX1_HVT \ram_reg[3][99]  ( .CLK(n281), .D(N116), .Q(\ram[3][99] ) );
  LATCHX1_HVT \ram_reg[3][98]  ( .CLK(n282), .D(N114), .Q(\ram[3][98] ) );
  LATCHX1_HVT \ram_reg[3][97]  ( .CLK(n283), .D(N113), .Q(\ram[3][97] ) );
  LATCHX1_HVT \ram_reg[3][96]  ( .CLK(n287), .D(N112), .Q(\ram[3][96] ) );
  LATCHX1_HVT \ram_reg[3][95]  ( .CLK(n279), .D(N111), .Q(\ram[3][95] ) );
  LATCHX1_HVT \ram_reg[3][94]  ( .CLK(n279), .D(N110), .Q(\ram[3][94] ) );
  LATCHX1_HVT \ram_reg[3][93]  ( .CLK(n279), .D(N109), .Q(\ram[3][93] ) );
  LATCHX1_HVT \ram_reg[3][92]  ( .CLK(n278), .D(N108), .Q(\ram[3][92] ) );
  LATCHX1_HVT \ram_reg[3][91]  ( .CLK(n278), .D(N107), .Q(\ram[3][91] ) );
  LATCHX1_HVT \ram_reg[3][90]  ( .CLK(n279), .D(N106), .Q(\ram[3][90] ) );
  LATCHX1_HVT \ram_reg[3][89]  ( .CLK(n278), .D(N105), .Q(\ram[3][89] ) );
  LATCHX1_HVT \ram_reg[3][88]  ( .CLK(n279), .D(N104), .Q(\ram[3][88] ) );
  LATCHX1_HVT \ram_reg[3][87]  ( .CLK(n287), .D(N103), .Q(\ram[3][87] ) );
  LATCHX1_HVT \ram_reg[3][86]  ( .CLK(n286), .D(N102), .Q(\ram[3][86] ) );
  LATCHX1_HVT \ram_reg[3][85]  ( .CLK(n285), .D(N101), .Q(\ram[3][85] ) );
  LATCHX1_HVT \ram_reg[3][84]  ( .CLK(n285), .D(N100), .Q(\ram[3][84] ) );
  LATCHX1_HVT \ram_reg[3][83]  ( .CLK(n280), .D(N99), .Q(\ram[3][83] ) );
  LATCHX1_HVT \ram_reg[3][82]  ( .CLK(n286), .D(N98), .Q(\ram[3][82] ) );
  LATCHX1_HVT \ram_reg[3][81]  ( .CLK(n285), .D(N97), .Q(\ram[3][81] ) );
  LATCHX1_HVT \ram_reg[3][80]  ( .CLK(n286), .D(N96), .Q(\ram[3][80] ) );
  LATCHX1_HVT \ram_reg[3][79]  ( .CLK(n280), .D(N95), .Q(\ram[3][79] ) );
  LATCHX1_HVT \ram_reg[3][78]  ( .CLK(n279), .D(N94), .Q(\ram[3][78] ) );
  LATCHX1_HVT \ram_reg[3][77]  ( .CLK(n280), .D(N93), .Q(\ram[3][77] ) );
  LATCHX1_HVT \ram_reg[3][76]  ( .CLK(n279), .D(N92), .Q(\ram[3][76] ) );
  LATCHX1_HVT \ram_reg[3][75]  ( .CLK(n279), .D(N91), .Q(\ram[3][75] ) );
  LATCHX1_HVT \ram_reg[3][74]  ( .CLK(n277), .D(N90), .Q(\ram[3][74] ) );
  LATCHX1_HVT \ram_reg[3][73]  ( .CLK(n280), .D(N89), .Q(\ram[3][73] ) );
  LATCHX1_HVT \ram_reg[3][72]  ( .CLK(n280), .D(N88), .Q(\ram[3][72] ) );
  LATCHX1_HVT \ram_reg[3][71]  ( .CLK(n283), .D(N87), .Q(\ram[3][71] ) );
  LATCHX1_HVT \ram_reg[3][70]  ( .CLK(n283), .D(N86), .Q(\ram[3][70] ) );
  LATCHX1_HVT \ram_reg[3][69]  ( .CLK(n282), .D(N85), .Q(\ram[3][69] ) );
  LATCHX1_HVT \ram_reg[3][68]  ( .CLK(n283), .D(N84), .Q(\ram[3][68] ) );
  LATCHX1_HVT \ram_reg[3][67]  ( .CLK(n282), .D(N83), .Q(\ram[3][67] ) );
  LATCHX1_HVT \ram_reg[3][66]  ( .CLK(n281), .D(N82), .Q(\ram[3][66] ) );
  LATCHX1_HVT \ram_reg[3][65]  ( .CLK(n282), .D(N81), .Q(\ram[3][65] ) );
  LATCHX1_HVT \ram_reg[3][64]  ( .CLK(n287), .D(N80), .Q(\ram[3][64] ) );
  LATCHX1_HVT \ram_reg[3][63]  ( .CLK(n281), .D(N79), .Q(\ram[3][63] ) );
  LATCHX1_HVT \ram_reg[3][62]  ( .CLK(n281), .D(N78), .Q(\ram[3][62] ) );
  LATCHX1_HVT \ram_reg[3][61]  ( .CLK(n281), .D(N77), .Q(\ram[3][61] ) );
  LATCHX1_HVT \ram_reg[3][60]  ( .CLK(n281), .D(N76), .Q(\ram[3][60] ) );
  LATCHX1_HVT \ram_reg[3][59]  ( .CLK(n281), .D(N75), .Q(\ram[3][59] ) );
  LATCHX1_HVT \ram_reg[3][58]  ( .CLK(n280), .D(N74), .Q(\ram[3][58] ) );
  LATCHX1_HVT \ram_reg[3][57]  ( .CLK(n281), .D(N73), .Q(\ram[3][57] ) );
  LATCHX1_HVT \ram_reg[3][56]  ( .CLK(n281), .D(N72), .Q(\ram[3][56] ) );
  LATCHX1_HVT \ram_reg[3][55]  ( .CLK(n287), .D(N71), .Q(\ram[3][55] ) );
  LATCHX1_HVT \ram_reg[3][54]  ( .CLK(n285), .D(N70), .Q(\ram[3][54] ) );
  LATCHX1_HVT \ram_reg[3][53]  ( .CLK(n285), .D(N69), .Q(\ram[3][53] ) );
  LATCHX1_HVT \ram_reg[3][52]  ( .CLK(n286), .D(N68), .Q(\ram[3][52] ) );
  LATCHX1_HVT \ram_reg[3][51]  ( .CLK(n280), .D(N67), .Q(\ram[3][51] ) );
  LATCHX1_HVT \ram_reg[3][50]  ( .CLK(n277), .D(N66), .Q(\ram[3][50] ) );
  LATCHX1_HVT \ram_reg[3][49]  ( .CLK(n286), .D(N65), .Q(\ram[3][49] ) );
  LATCHX1_HVT \ram_reg[3][48]  ( .CLK(n286), .D(N64), .Q(\ram[3][48] ) );
  LATCHX1_HVT \ram_reg[3][47]  ( .CLK(n284), .D(N63), .Q(\ram[3][47] ) );
  LATCHX1_HVT \ram_reg[3][46]  ( .CLK(n284), .D(N62), .Q(\ram[3][46] ) );
  LATCHX1_HVT \ram_reg[3][45]  ( .CLK(n284), .D(N61), .Q(\ram[3][45] ) );
  LATCHX1_HVT \ram_reg[3][44]  ( .CLK(n284), .D(N60), .Q(\ram[3][44] ) );
  LATCHX1_HVT \ram_reg[3][43]  ( .CLK(n281), .D(N59), .Q(\ram[3][43] ) );
  LATCHX1_HVT \ram_reg[3][42]  ( .CLK(n285), .D(N58), .Q(\ram[3][42] ) );
  LATCHX1_HVT \ram_reg[3][41]  ( .CLK(n278), .D(N57), .Q(\ram[3][41] ) );
  LATCHX1_HVT \ram_reg[3][40]  ( .CLK(n284), .D(N56), .Q(\ram[3][40] ) );
  LATCHX1_HVT \ram_reg[3][39]  ( .CLK(n283), .D(N55), .Q(\ram[3][39] ) );
  LATCHX1_HVT \ram_reg[3][38]  ( .CLK(n283), .D(N54), .Q(\ram[3][38] ) );
  LATCHX1_HVT \ram_reg[3][37]  ( .CLK(n282), .D(N53), .Q(\ram[3][37] ) );
  LATCHX1_HVT \ram_reg[3][36]  ( .CLK(n282), .D(N52), .Q(\ram[3][36] ) );
  LATCHX1_HVT \ram_reg[3][35]  ( .CLK(n282), .D(N51), .Q(\ram[3][35] ) );
  LATCHX1_HVT \ram_reg[3][34]  ( .CLK(n284), .D(N50), .Q(\ram[3][34] ) );
  LATCHX1_HVT \ram_reg[3][33]  ( .CLK(n283), .D(N49), .Q(\ram[3][33] ) );
  LATCHX1_HVT \ram_reg[3][32]  ( .CLK(n287), .D(N48), .Q(\ram[3][32] ) );
  LATCHX1_HVT \ram_reg[3][31]  ( .CLK(n277), .D(N47), .Q(\ram[3][31] ) );
  LATCHX1_HVT \ram_reg[3][30]  ( .CLK(n277), .D(N46), .Q(\ram[3][30] ) );
  LATCHX1_HVT \ram_reg[3][29]  ( .CLK(n277), .D(N45), .Q(\ram[3][29] ) );
  LATCHX1_HVT \ram_reg[3][28]  ( .CLK(n277), .D(N44), .Q(\ram[3][28] ) );
  LATCHX1_HVT \ram_reg[3][27]  ( .CLK(n277), .D(N43), .Q(\ram[3][27] ) );
  LATCHX1_HVT \ram_reg[3][26]  ( .CLK(n277), .D(N42), .Q(\ram[3][26] ) );
  LATCHX1_HVT \ram_reg[3][25]  ( .CLK(n277), .D(N41), .Q(\ram[3][25] ) );
  LATCHX1_HVT \ram_reg[3][24]  ( .CLK(n277), .D(N40), .Q(\ram[3][24] ) );
  LATCHX1_HVT \ram_reg[3][23]  ( .CLK(n287), .D(N39), .Q(\ram[3][23] ) );
  LATCHX1_HVT \ram_reg[3][22]  ( .CLK(n286), .D(N38), .Q(\ram[3][22] ) );
  LATCHX1_HVT \ram_reg[3][21]  ( .CLK(n285), .D(N37), .Q(\ram[3][21] ) );
  LATCHX1_HVT \ram_reg[3][20]  ( .CLK(n285), .D(N36), .Q(\ram[3][20] ) );
  LATCHX1_HVT \ram_reg[3][19]  ( .CLK(n277), .D(N35), .Q(\ram[3][19] ) );
  LATCHX1_HVT \ram_reg[3][18]  ( .CLK(n285), .D(N34), .Q(\ram[3][18] ) );
  LATCHX1_HVT \ram_reg[3][17]  ( .CLK(n286), .D(N33), .Q(\ram[3][17] ) );
  LATCHX1_HVT \ram_reg[3][16]  ( .CLK(n286), .D(N32), .Q(\ram[3][16] ) );
  LATCHX1_HVT \ram_reg[3][15]  ( .CLK(n280), .D(N31), .Q(\ram[3][15] ) );
  LATCHX1_HVT \ram_reg[3][14]  ( .CLK(n280), .D(N30), .Q(\ram[3][14] ) );
  LATCHX1_HVT \ram_reg[3][13]  ( .CLK(n279), .D(N29), .Q(\ram[3][13] ) );
  LATCHX1_HVT \ram_reg[3][12]  ( .CLK(n279), .D(N28), .Q(\ram[3][12] ) );
  LATCHX1_HVT \ram_reg[3][11]  ( .CLK(n280), .D(N27), .Q(\ram[3][11] ) );
  LATCHX1_HVT \ram_reg[3][10]  ( .CLK(n279), .D(N26), .Q(\ram[3][10] ) );
  LATCHX1_HVT \ram_reg[3][9]  ( .CLK(n279), .D(N25), .Q(\ram[3][9] ) );
  LATCHX1_HVT \ram_reg[3][8]  ( .CLK(n280), .D(N24), .Q(\ram[3][8] ) );
  LATCHX1_HVT \ram_reg[3][7]  ( .CLK(n283), .D(N23), .Q(\ram[3][7] ) );
  LATCHX1_HVT \ram_reg[3][6]  ( .CLK(n283), .D(N22), .Q(\ram[3][6] ) );
  LATCHX1_HVT \ram_reg[3][5]  ( .CLK(n282), .D(N21), .Q(\ram[3][5] ) );
  LATCHX1_HVT \ram_reg[3][4]  ( .CLK(n282), .D(N20), .Q(\ram[3][4] ) );
  LATCHX1_HVT \ram_reg[3][3]  ( .CLK(n281), .D(N19), .Q(\ram[3][3] ) );
  LATCHX1_HVT \ram_reg[3][2]  ( .CLK(n282), .D(N18), .Q(\ram[3][2] ) );
  LATCHX1_HVT \ram_reg[3][1]  ( .CLK(n283), .D(N17), .Q(\ram[3][1] ) );
  LATCHX1_HVT \ram_reg[3][0]  ( .CLK(n287), .D(N16), .Q(\ram[3][0] ) );
  LATCHX1_HVT \ram_reg[2][255]  ( .CLK(N279), .D(N273), .Q(\ram[2][255] ) );
  LATCHX1_HVT \ram_reg[2][254]  ( .CLK(N279), .D(N272), .Q(\ram[2][254] ) );
  LATCHX1_HVT \ram_reg[2][253]  ( .CLK(N279), .D(N271), .Q(\ram[2][253] ) );
  LATCHX1_HVT \ram_reg[2][252]  ( .CLK(N279), .D(N270), .Q(\ram[2][252] ) );
  LATCHX1_HVT \ram_reg[2][251]  ( .CLK(n320), .D(N269), .Q(\ram[2][251] ) );
  LATCHX1_HVT \ram_reg[2][250]  ( .CLK(n312), .D(N268), .Q(\ram[2][250] ) );
  LATCHX1_HVT \ram_reg[2][249]  ( .CLK(n312), .D(N267), .Q(\ram[2][249] ) );
  LATCHX1_HVT \ram_reg[2][248]  ( .CLK(n312), .D(N266), .Q(\ram[2][248] ) );
  LATCHX1_HVT \ram_reg[2][247]  ( .CLK(n312), .D(N265), .Q(\ram[2][247] ) );
  LATCHX1_HVT \ram_reg[2][246]  ( .CLK(n312), .D(N264), .Q(\ram[2][246] ) );
  LATCHX1_HVT \ram_reg[2][245]  ( .CLK(n312), .D(N263), .Q(\ram[2][245] ) );
  LATCHX1_HVT \ram_reg[2][244]  ( .CLK(n312), .D(N262), .Q(\ram[2][244] ) );
  LATCHX1_HVT \ram_reg[2][243]  ( .CLK(n312), .D(N261), .Q(\ram[2][243] ) );
  LATCHX1_HVT \ram_reg[2][242]  ( .CLK(n312), .D(N260), .Q(\ram[2][242] ) );
  LATCHX1_HVT \ram_reg[2][241]  ( .CLK(n311), .D(N259), .Q(\ram[2][241] ) );
  LATCHX1_HVT \ram_reg[2][240]  ( .CLK(n311), .D(N258), .Q(\ram[2][240] ) );
  LATCHX1_HVT \ram_reg[2][239]  ( .CLK(n311), .D(N257), .Q(\ram[2][239] ) );
  LATCHX1_HVT \ram_reg[2][238]  ( .CLK(n311), .D(N256), .Q(\ram[2][238] ) );
  LATCHX1_HVT \ram_reg[2][237]  ( .CLK(n311), .D(N255), .Q(\ram[2][237] ) );
  LATCHX1_HVT \ram_reg[2][236]  ( .CLK(n311), .D(N254), .Q(\ram[2][236] ) );
  LATCHX1_HVT \ram_reg[2][235]  ( .CLK(n311), .D(N253), .Q(\ram[2][235] ) );
  LATCHX1_HVT \ram_reg[2][234]  ( .CLK(n311), .D(N252), .Q(\ram[2][234] ) );
  LATCHX1_HVT \ram_reg[2][233]  ( .CLK(n311), .D(N251), .Q(\ram[2][233] ) );
  LATCHX1_HVT \ram_reg[2][232]  ( .CLK(n311), .D(N250), .Q(\ram[2][232] ) );
  LATCHX1_HVT \ram_reg[2][231]  ( .CLK(n311), .D(N249), .Q(\ram[2][231] ) );
  LATCHX1_HVT \ram_reg[2][230]  ( .CLK(n310), .D(N248), .Q(\ram[2][230] ) );
  LATCHX1_HVT \ram_reg[2][229]  ( .CLK(n310), .D(N247), .Q(\ram[2][229] ) );
  LATCHX1_HVT \ram_reg[2][228]  ( .CLK(n310), .D(N246), .Q(\ram[2][228] ) );
  LATCHX1_HVT \ram_reg[2][227]  ( .CLK(n320), .D(N245), .Q(\ram[2][227] ) );
  LATCHX1_HVT \ram_reg[2][226]  ( .CLK(n320), .D(N244), .Q(\ram[2][226] ) );
  LATCHX1_HVT \ram_reg[2][225]  ( .CLK(n320), .D(N243), .Q(\ram[2][225] ) );
  LATCHX1_HVT \ram_reg[2][224]  ( .CLK(n320), .D(N242), .Q(\ram[2][224] ) );
  LATCHX1_HVT \ram_reg[2][223]  ( .CLK(n320), .D(N241), .Q(\ram[2][223] ) );
  LATCHX1_HVT \ram_reg[2][222]  ( .CLK(n320), .D(N240), .Q(\ram[2][222] ) );
  LATCHX1_HVT \ram_reg[2][221]  ( .CLK(n320), .D(N239), .Q(\ram[2][221] ) );
  LATCHX1_HVT \ram_reg[2][220]  ( .CLK(n320), .D(N238), .Q(\ram[2][220] ) );
  LATCHX1_HVT \ram_reg[2][219]  ( .CLK(n320), .D(N237), .Q(\ram[2][219] ) );
  LATCHX1_HVT \ram_reg[2][218]  ( .CLK(n320), .D(N236), .Q(\ram[2][218] ) );
  LATCHX1_HVT \ram_reg[2][217]  ( .CLK(n319), .D(N235), .Q(\ram[2][217] ) );
  LATCHX1_HVT \ram_reg[2][216]  ( .CLK(n319), .D(N234), .Q(\ram[2][216] ) );
  LATCHX1_HVT \ram_reg[2][215]  ( .CLK(n319), .D(N233), .Q(\ram[2][215] ) );
  LATCHX1_HVT \ram_reg[2][214]  ( .CLK(n319), .D(N232), .Q(\ram[2][214] ) );
  LATCHX1_HVT \ram_reg[2][213]  ( .CLK(n319), .D(N231), .Q(\ram[2][213] ) );
  LATCHX1_HVT \ram_reg[2][212]  ( .CLK(n319), .D(N230), .Q(\ram[2][212] ) );
  LATCHX1_HVT \ram_reg[2][211]  ( .CLK(n319), .D(N229), .Q(\ram[2][211] ) );
  LATCHX1_HVT \ram_reg[2][210]  ( .CLK(n319), .D(N228), .Q(\ram[2][210] ) );
  LATCHX1_HVT \ram_reg[2][209]  ( .CLK(n319), .D(N227), .Q(\ram[2][209] ) );
  LATCHX1_HVT \ram_reg[2][208]  ( .CLK(n319), .D(N226), .Q(\ram[2][208] ) );
  LATCHX1_HVT \ram_reg[2][207]  ( .CLK(n318), .D(N225), .Q(\ram[2][207] ) );
  LATCHX1_HVT \ram_reg[2][206]  ( .CLK(n318), .D(N224), .Q(\ram[2][206] ) );
  LATCHX1_HVT \ram_reg[2][205]  ( .CLK(n318), .D(N223), .Q(\ram[2][205] ) );
  LATCHX1_HVT \ram_reg[2][204]  ( .CLK(n318), .D(N222), .Q(\ram[2][204] ) );
  LATCHX1_HVT \ram_reg[2][203]  ( .CLK(n318), .D(N221), .Q(\ram[2][203] ) );
  LATCHX1_HVT \ram_reg[2][202]  ( .CLK(n318), .D(N220), .Q(\ram[2][202] ) );
  LATCHX1_HVT \ram_reg[2][201]  ( .CLK(n318), .D(N219), .Q(\ram[2][201] ) );
  LATCHX1_HVT \ram_reg[2][200]  ( .CLK(n318), .D(N218), .Q(\ram[2][200] ) );
  LATCHX1_HVT \ram_reg[2][199]  ( .CLK(n318), .D(N217), .Q(\ram[2][199] ) );
  LATCHX1_HVT \ram_reg[2][198]  ( .CLK(n318), .D(N216), .Q(\ram[2][198] ) );
  LATCHX1_HVT \ram_reg[2][197]  ( .CLK(n318), .D(N214), .Q(\ram[2][197] ) );
  LATCHX1_HVT \ram_reg[2][196]  ( .CLK(n317), .D(N213), .Q(\ram[2][196] ) );
  LATCHX1_HVT \ram_reg[2][195]  ( .CLK(n317), .D(N212), .Q(\ram[2][195] ) );
  LATCHX1_HVT \ram_reg[2][194]  ( .CLK(n317), .D(N211), .Q(\ram[2][194] ) );
  LATCHX1_HVT \ram_reg[2][193]  ( .CLK(n317), .D(N210), .Q(\ram[2][193] ) );
  LATCHX1_HVT \ram_reg[2][192]  ( .CLK(n317), .D(N209), .Q(\ram[2][192] ) );
  LATCHX1_HVT \ram_reg[2][191]  ( .CLK(n317), .D(N208), .Q(\ram[2][191] ) );
  LATCHX1_HVT \ram_reg[2][190]  ( .CLK(n317), .D(N207), .Q(\ram[2][190] ) );
  LATCHX1_HVT \ram_reg[2][189]  ( .CLK(n317), .D(N206), .Q(\ram[2][189] ) );
  LATCHX1_HVT \ram_reg[2][188]  ( .CLK(n317), .D(N205), .Q(\ram[2][188] ) );
  LATCHX1_HVT \ram_reg[2][187]  ( .CLK(n317), .D(N204), .Q(\ram[2][187] ) );
  LATCHX1_HVT \ram_reg[2][186]  ( .CLK(n317), .D(N203), .Q(\ram[2][186] ) );
  LATCHX1_HVT \ram_reg[2][185]  ( .CLK(n316), .D(N202), .Q(\ram[2][185] ) );
  LATCHX1_HVT \ram_reg[2][184]  ( .CLK(n316), .D(N201), .Q(\ram[2][184] ) );
  LATCHX1_HVT \ram_reg[2][183]  ( .CLK(n316), .D(N200), .Q(\ram[2][183] ) );
  LATCHX1_HVT \ram_reg[2][182]  ( .CLK(n316), .D(N199), .Q(\ram[2][182] ) );
  LATCHX1_HVT \ram_reg[2][181]  ( .CLK(n316), .D(N198), .Q(\ram[2][181] ) );
  LATCHX1_HVT \ram_reg[2][180]  ( .CLK(n316), .D(N197), .Q(\ram[2][180] ) );
  LATCHX1_HVT \ram_reg[2][179]  ( .CLK(n316), .D(N196), .Q(\ram[2][179] ) );
  LATCHX1_HVT \ram_reg[2][178]  ( .CLK(n316), .D(N195), .Q(\ram[2][178] ) );
  LATCHX1_HVT \ram_reg[2][177]  ( .CLK(n316), .D(N194), .Q(\ram[2][177] ) );
  LATCHX1_HVT \ram_reg[2][176]  ( .CLK(n316), .D(N193), .Q(\ram[2][176] ) );
  LATCHX1_HVT \ram_reg[2][175]  ( .CLK(n316), .D(N192), .Q(\ram[2][175] ) );
  LATCHX1_HVT \ram_reg[2][174]  ( .CLK(n315), .D(N191), .Q(\ram[2][174] ) );
  LATCHX1_HVT \ram_reg[2][173]  ( .CLK(n315), .D(N190), .Q(\ram[2][173] ) );
  LATCHX1_HVT \ram_reg[2][172]  ( .CLK(n315), .D(N189), .Q(\ram[2][172] ) );
  LATCHX1_HVT \ram_reg[2][171]  ( .CLK(n315), .D(N188), .Q(\ram[2][171] ) );
  LATCHX1_HVT \ram_reg[2][170]  ( .CLK(n315), .D(N187), .Q(\ram[2][170] ) );
  LATCHX1_HVT \ram_reg[2][169]  ( .CLK(n315), .D(N186), .Q(\ram[2][169] ) );
  LATCHX1_HVT \ram_reg[2][168]  ( .CLK(n315), .D(N185), .Q(\ram[2][168] ) );
  LATCHX1_HVT \ram_reg[2][167]  ( .CLK(n315), .D(N184), .Q(\ram[2][167] ) );
  LATCHX1_HVT \ram_reg[2][166]  ( .CLK(n315), .D(N183), .Q(\ram[2][166] ) );
  LATCHX1_HVT \ram_reg[2][165]  ( .CLK(n315), .D(N182), .Q(\ram[2][165] ) );
  LATCHX1_HVT \ram_reg[2][164]  ( .CLK(n315), .D(N181), .Q(\ram[2][164] ) );
  LATCHX1_HVT \ram_reg[2][163]  ( .CLK(n314), .D(N180), .Q(\ram[2][163] ) );
  LATCHX1_HVT \ram_reg[2][162]  ( .CLK(n314), .D(N179), .Q(\ram[2][162] ) );
  LATCHX1_HVT \ram_reg[2][161]  ( .CLK(n314), .D(N178), .Q(\ram[2][161] ) );
  LATCHX1_HVT \ram_reg[2][160]  ( .CLK(n314), .D(N177), .Q(\ram[2][160] ) );
  LATCHX1_HVT \ram_reg[2][159]  ( .CLK(n314), .D(N176), .Q(\ram[2][159] ) );
  LATCHX1_HVT \ram_reg[2][158]  ( .CLK(n314), .D(N175), .Q(\ram[2][158] ) );
  LATCHX1_HVT \ram_reg[2][157]  ( .CLK(n314), .D(N174), .Q(\ram[2][157] ) );
  LATCHX1_HVT \ram_reg[2][156]  ( .CLK(n314), .D(N173), .Q(\ram[2][156] ) );
  LATCHX1_HVT \ram_reg[2][155]  ( .CLK(n314), .D(N172), .Q(\ram[2][155] ) );
  LATCHX1_HVT \ram_reg[2][154]  ( .CLK(n314), .D(N171), .Q(\ram[2][154] ) );
  LATCHX1_HVT \ram_reg[2][153]  ( .CLK(n314), .D(N170), .Q(\ram[2][153] ) );
  LATCHX1_HVT \ram_reg[2][152]  ( .CLK(n313), .D(N169), .Q(\ram[2][152] ) );
  LATCHX1_HVT \ram_reg[2][151]  ( .CLK(n313), .D(N168), .Q(\ram[2][151] ) );
  LATCHX1_HVT \ram_reg[2][150]  ( .CLK(n313), .D(N167), .Q(\ram[2][150] ) );
  LATCHX1_HVT \ram_reg[2][149]  ( .CLK(n313), .D(N166), .Q(\ram[2][149] ) );
  LATCHX1_HVT \ram_reg[2][148]  ( .CLK(n313), .D(N165), .Q(\ram[2][148] ) );
  LATCHX1_HVT \ram_reg[2][147]  ( .CLK(n313), .D(N164), .Q(\ram[2][147] ) );
  LATCHX1_HVT \ram_reg[2][146]  ( .CLK(n313), .D(N163), .Q(\ram[2][146] ) );
  LATCHX1_HVT \ram_reg[2][145]  ( .CLK(n313), .D(N162), .Q(\ram[2][145] ) );
  LATCHX1_HVT \ram_reg[2][144]  ( .CLK(n313), .D(N161), .Q(\ram[2][144] ) );
  LATCHX1_HVT \ram_reg[2][143]  ( .CLK(n313), .D(N160), .Q(\ram[2][143] ) );
  LATCHX1_HVT \ram_reg[2][142]  ( .CLK(n313), .D(N159), .Q(\ram[2][142] ) );
  LATCHX1_HVT \ram_reg[2][141]  ( .CLK(n312), .D(N158), .Q(\ram[2][141] ) );
  LATCHX1_HVT \ram_reg[2][140]  ( .CLK(n312), .D(N157), .Q(\ram[2][140] ) );
  LATCHX1_HVT \ram_reg[2][139]  ( .CLK(n312), .D(N156), .Q(\ram[2][139] ) );
  LATCHX1_HVT \ram_reg[2][138]  ( .CLK(n311), .D(N155), .Q(\ram[2][138] ) );
  LATCHX1_HVT \ram_reg[2][137]  ( .CLK(n320), .D(N154), .Q(\ram[2][137] ) );
  LATCHX1_HVT \ram_reg[2][136]  ( .CLK(n319), .D(N153), .Q(\ram[2][136] ) );
  LATCHX1_HVT \ram_reg[2][135]  ( .CLK(n319), .D(N152), .Q(\ram[2][135] ) );
  LATCHX1_HVT \ram_reg[2][134]  ( .CLK(n318), .D(N151), .Q(\ram[2][134] ) );
  LATCHX1_HVT \ram_reg[2][133]  ( .CLK(n317), .D(N150), .Q(\ram[2][133] ) );
  LATCHX1_HVT \ram_reg[2][132]  ( .CLK(n316), .D(N149), .Q(\ram[2][132] ) );
  LATCHX1_HVT \ram_reg[2][131]  ( .CLK(n315), .D(N148), .Q(\ram[2][131] ) );
  LATCHX1_HVT \ram_reg[2][130]  ( .CLK(n314), .D(N147), .Q(\ram[2][130] ) );
  LATCHX1_HVT \ram_reg[2][129]  ( .CLK(n313), .D(N146), .Q(\ram[2][129] ) );
  LATCHX1_HVT \ram_reg[2][128]  ( .CLK(n310), .D(N145), .Q(\ram[2][128] ) );
  LATCHX1_HVT \ram_reg[2][127]  ( .CLK(n301), .D(N144), .Q(\ram[2][127] ) );
  LATCHX1_HVT \ram_reg[2][126]  ( .CLK(n301), .D(N143), .Q(\ram[2][126] ) );
  LATCHX1_HVT \ram_reg[2][125]  ( .CLK(n301), .D(N142), .Q(\ram[2][125] ) );
  LATCHX1_HVT \ram_reg[2][124]  ( .CLK(n301), .D(N141), .Q(\ram[2][124] ) );
  LATCHX1_HVT \ram_reg[2][123]  ( .CLK(n301), .D(N140), .Q(\ram[2][123] ) );
  LATCHX1_HVT \ram_reg[2][122]  ( .CLK(n300), .D(N139), .Q(\ram[2][122] ) );
  LATCHX1_HVT \ram_reg[2][121]  ( .CLK(n301), .D(N138), .Q(\ram[2][121] ) );
  LATCHX1_HVT \ram_reg[2][120]  ( .CLK(n301), .D(N137), .Q(\ram[2][120] ) );
  LATCHX1_HVT \ram_reg[2][119]  ( .CLK(n310), .D(N136), .Q(\ram[2][119] ) );
  LATCHX1_HVT \ram_reg[2][118]  ( .CLK(n309), .D(N135), .Q(\ram[2][118] ) );
  LATCHX1_HVT \ram_reg[2][117]  ( .CLK(n309), .D(N134), .Q(\ram[2][117] ) );
  LATCHX1_HVT \ram_reg[2][116]  ( .CLK(n308), .D(N133), .Q(\ram[2][116] ) );
  LATCHX1_HVT \ram_reg[2][115]  ( .CLK(n303), .D(N132), .Q(\ram[2][115] ) );
  LATCHX1_HVT \ram_reg[2][114]  ( .CLK(n308), .D(N131), .Q(\ram[2][114] ) );
  LATCHX1_HVT \ram_reg[2][113]  ( .CLK(n308), .D(N130), .Q(\ram[2][113] ) );
  LATCHX1_HVT \ram_reg[2][112]  ( .CLK(n309), .D(N129), .Q(\ram[2][112] ) );
  LATCHX1_HVT \ram_reg[2][111]  ( .CLK(n307), .D(N128), .Q(\ram[2][111] ) );
  LATCHX1_HVT \ram_reg[2][110]  ( .CLK(n307), .D(N127), .Q(\ram[2][110] ) );
  LATCHX1_HVT \ram_reg[2][109]  ( .CLK(n307), .D(N126), .Q(\ram[2][109] ) );
  LATCHX1_HVT \ram_reg[2][108]  ( .CLK(n304), .D(N125), .Q(\ram[2][108] ) );
  LATCHX1_HVT \ram_reg[2][107]  ( .CLK(n301), .D(N124), .Q(\ram[2][107] ) );
  LATCHX1_HVT \ram_reg[2][106]  ( .CLK(n307), .D(N123), .Q(\ram[2][106] ) );
  LATCHX1_HVT \ram_reg[2][105]  ( .CLK(n307), .D(N122), .Q(\ram[2][105] ) );
  LATCHX1_HVT \ram_reg[2][104]  ( .CLK(n307), .D(N121), .Q(\ram[2][104] ) );
  LATCHX1_HVT \ram_reg[2][103]  ( .CLK(n306), .D(N120), .Q(\ram[2][103] ) );
  LATCHX1_HVT \ram_reg[2][102]  ( .CLK(n305), .D(N119), .Q(\ram[2][102] ) );
  LATCHX1_HVT \ram_reg[2][101]  ( .CLK(n305), .D(N118), .Q(\ram[2][101] ) );
  LATCHX1_HVT \ram_reg[2][100]  ( .CLK(n306), .D(N117), .Q(\ram[2][100] ) );
  LATCHX1_HVT \ram_reg[2][99]  ( .CLK(n304), .D(N116), .Q(\ram[2][99] ) );
  LATCHX1_HVT \ram_reg[2][98]  ( .CLK(n305), .D(N114), .Q(\ram[2][98] ) );
  LATCHX1_HVT \ram_reg[2][97]  ( .CLK(n306), .D(N113), .Q(\ram[2][97] ) );
  LATCHX1_HVT \ram_reg[2][96]  ( .CLK(n310), .D(N112), .Q(\ram[2][96] ) );
  LATCHX1_HVT \ram_reg[2][95]  ( .CLK(n302), .D(N111), .Q(\ram[2][95] ) );
  LATCHX1_HVT \ram_reg[2][94]  ( .CLK(n302), .D(N110), .Q(\ram[2][94] ) );
  LATCHX1_HVT \ram_reg[2][93]  ( .CLK(n302), .D(N109), .Q(\ram[2][93] ) );
  LATCHX1_HVT \ram_reg[2][92]  ( .CLK(n301), .D(N108), .Q(\ram[2][92] ) );
  LATCHX1_HVT \ram_reg[2][91]  ( .CLK(n301), .D(N107), .Q(\ram[2][91] ) );
  LATCHX1_HVT \ram_reg[2][90]  ( .CLK(n302), .D(N106), .Q(\ram[2][90] ) );
  LATCHX1_HVT \ram_reg[2][89]  ( .CLK(n301), .D(N105), .Q(\ram[2][89] ) );
  LATCHX1_HVT \ram_reg[2][88]  ( .CLK(n302), .D(N104), .Q(\ram[2][88] ) );
  LATCHX1_HVT \ram_reg[2][87]  ( .CLK(n310), .D(N103), .Q(\ram[2][87] ) );
  LATCHX1_HVT \ram_reg[2][86]  ( .CLK(n309), .D(N102), .Q(\ram[2][86] ) );
  LATCHX1_HVT \ram_reg[2][85]  ( .CLK(n308), .D(N101), .Q(\ram[2][85] ) );
  LATCHX1_HVT \ram_reg[2][84]  ( .CLK(n308), .D(N100), .Q(\ram[2][84] ) );
  LATCHX1_HVT \ram_reg[2][83]  ( .CLK(n303), .D(N99), .Q(\ram[2][83] ) );
  LATCHX1_HVT \ram_reg[2][82]  ( .CLK(n309), .D(N98), .Q(\ram[2][82] ) );
  LATCHX1_HVT \ram_reg[2][81]  ( .CLK(n308), .D(N97), .Q(\ram[2][81] ) );
  LATCHX1_HVT \ram_reg[2][80]  ( .CLK(n309), .D(N96), .Q(\ram[2][80] ) );
  LATCHX1_HVT \ram_reg[2][79]  ( .CLK(n303), .D(N95), .Q(\ram[2][79] ) );
  LATCHX1_HVT \ram_reg[2][78]  ( .CLK(n302), .D(N94), .Q(\ram[2][78] ) );
  LATCHX1_HVT \ram_reg[2][77]  ( .CLK(n303), .D(N93), .Q(\ram[2][77] ) );
  LATCHX1_HVT \ram_reg[2][76]  ( .CLK(n302), .D(N92), .Q(\ram[2][76] ) );
  LATCHX1_HVT \ram_reg[2][75]  ( .CLK(n302), .D(N91), .Q(\ram[2][75] ) );
  LATCHX1_HVT \ram_reg[2][74]  ( .CLK(n300), .D(N90), .Q(\ram[2][74] ) );
  LATCHX1_HVT \ram_reg[2][73]  ( .CLK(n303), .D(N89), .Q(\ram[2][73] ) );
  LATCHX1_HVT \ram_reg[2][72]  ( .CLK(n303), .D(N88), .Q(\ram[2][72] ) );
  LATCHX1_HVT \ram_reg[2][71]  ( .CLK(n306), .D(N87), .Q(\ram[2][71] ) );
  LATCHX1_HVT \ram_reg[2][70]  ( .CLK(n306), .D(N86), .Q(\ram[2][70] ) );
  LATCHX1_HVT \ram_reg[2][69]  ( .CLK(n305), .D(N85), .Q(\ram[2][69] ) );
  LATCHX1_HVT \ram_reg[2][68]  ( .CLK(n306), .D(N84), .Q(\ram[2][68] ) );
  LATCHX1_HVT \ram_reg[2][67]  ( .CLK(n305), .D(N83), .Q(\ram[2][67] ) );
  LATCHX1_HVT \ram_reg[2][66]  ( .CLK(n304), .D(N82), .Q(\ram[2][66] ) );
  LATCHX1_HVT \ram_reg[2][65]  ( .CLK(n305), .D(N81), .Q(\ram[2][65] ) );
  LATCHX1_HVT \ram_reg[2][64]  ( .CLK(n310), .D(N80), .Q(\ram[2][64] ) );
  LATCHX1_HVT \ram_reg[2][63]  ( .CLK(n304), .D(N79), .Q(\ram[2][63] ) );
  LATCHX1_HVT \ram_reg[2][62]  ( .CLK(n304), .D(N78), .Q(\ram[2][62] ) );
  LATCHX1_HVT \ram_reg[2][61]  ( .CLK(n304), .D(N77), .Q(\ram[2][61] ) );
  LATCHX1_HVT \ram_reg[2][60]  ( .CLK(n304), .D(N76), .Q(\ram[2][60] ) );
  LATCHX1_HVT \ram_reg[2][59]  ( .CLK(n304), .D(N75), .Q(\ram[2][59] ) );
  LATCHX1_HVT \ram_reg[2][58]  ( .CLK(n303), .D(N74), .Q(\ram[2][58] ) );
  LATCHX1_HVT \ram_reg[2][57]  ( .CLK(n304), .D(N73), .Q(\ram[2][57] ) );
  LATCHX1_HVT \ram_reg[2][56]  ( .CLK(n304), .D(N72), .Q(\ram[2][56] ) );
  LATCHX1_HVT \ram_reg[2][55]  ( .CLK(n310), .D(N71), .Q(\ram[2][55] ) );
  LATCHX1_HVT \ram_reg[2][54]  ( .CLK(n308), .D(N70), .Q(\ram[2][54] ) );
  LATCHX1_HVT \ram_reg[2][53]  ( .CLK(n308), .D(N69), .Q(\ram[2][53] ) );
  LATCHX1_HVT \ram_reg[2][52]  ( .CLK(n309), .D(N68), .Q(\ram[2][52] ) );
  LATCHX1_HVT \ram_reg[2][51]  ( .CLK(n303), .D(N67), .Q(\ram[2][51] ) );
  LATCHX1_HVT \ram_reg[2][50]  ( .CLK(n300), .D(N66), .Q(\ram[2][50] ) );
  LATCHX1_HVT \ram_reg[2][49]  ( .CLK(n309), .D(N65), .Q(\ram[2][49] ) );
  LATCHX1_HVT \ram_reg[2][48]  ( .CLK(n309), .D(N64), .Q(\ram[2][48] ) );
  LATCHX1_HVT \ram_reg[2][47]  ( .CLK(n307), .D(N63), .Q(\ram[2][47] ) );
  LATCHX1_HVT \ram_reg[2][46]  ( .CLK(n307), .D(N62), .Q(\ram[2][46] ) );
  LATCHX1_HVT \ram_reg[2][45]  ( .CLK(n307), .D(N61), .Q(\ram[2][45] ) );
  LATCHX1_HVT \ram_reg[2][44]  ( .CLK(n307), .D(N60), .Q(\ram[2][44] ) );
  LATCHX1_HVT \ram_reg[2][43]  ( .CLK(n304), .D(N59), .Q(\ram[2][43] ) );
  LATCHX1_HVT \ram_reg[2][42]  ( .CLK(n308), .D(N58), .Q(\ram[2][42] ) );
  LATCHX1_HVT \ram_reg[2][41]  ( .CLK(n301), .D(N57), .Q(\ram[2][41] ) );
  LATCHX1_HVT \ram_reg[2][40]  ( .CLK(n307), .D(N56), .Q(\ram[2][40] ) );
  LATCHX1_HVT \ram_reg[2][39]  ( .CLK(n306), .D(N55), .Q(\ram[2][39] ) );
  LATCHX1_HVT \ram_reg[2][38]  ( .CLK(n306), .D(N54), .Q(\ram[2][38] ) );
  LATCHX1_HVT \ram_reg[2][37]  ( .CLK(n305), .D(N53), .Q(\ram[2][37] ) );
  LATCHX1_HVT \ram_reg[2][36]  ( .CLK(n305), .D(N52), .Q(\ram[2][36] ) );
  LATCHX1_HVT \ram_reg[2][35]  ( .CLK(n305), .D(N51), .Q(\ram[2][35] ) );
  LATCHX1_HVT \ram_reg[2][34]  ( .CLK(n307), .D(N50), .Q(\ram[2][34] ) );
  LATCHX1_HVT \ram_reg[2][33]  ( .CLK(n306), .D(N49), .Q(\ram[2][33] ) );
  LATCHX1_HVT \ram_reg[2][32]  ( .CLK(n310), .D(N48), .Q(\ram[2][32] ) );
  LATCHX1_HVT \ram_reg[2][31]  ( .CLK(n300), .D(N47), .Q(\ram[2][31] ) );
  LATCHX1_HVT \ram_reg[2][30]  ( .CLK(n300), .D(N46), .Q(\ram[2][30] ) );
  LATCHX1_HVT \ram_reg[2][29]  ( .CLK(n300), .D(N45), .Q(\ram[2][29] ) );
  LATCHX1_HVT \ram_reg[2][28]  ( .CLK(n300), .D(N44), .Q(\ram[2][28] ) );
  LATCHX1_HVT \ram_reg[2][27]  ( .CLK(n300), .D(N43), .Q(\ram[2][27] ) );
  LATCHX1_HVT \ram_reg[2][26]  ( .CLK(n300), .D(N42), .Q(\ram[2][26] ) );
  LATCHX1_HVT \ram_reg[2][25]  ( .CLK(n300), .D(N41), .Q(\ram[2][25] ) );
  LATCHX1_HVT \ram_reg[2][24]  ( .CLK(n300), .D(N40), .Q(\ram[2][24] ) );
  LATCHX1_HVT \ram_reg[2][23]  ( .CLK(n310), .D(N39), .Q(\ram[2][23] ) );
  LATCHX1_HVT \ram_reg[2][22]  ( .CLK(n309), .D(N38), .Q(\ram[2][22] ) );
  LATCHX1_HVT \ram_reg[2][21]  ( .CLK(n308), .D(N37), .Q(\ram[2][21] ) );
  LATCHX1_HVT \ram_reg[2][20]  ( .CLK(n308), .D(N36), .Q(\ram[2][20] ) );
  LATCHX1_HVT \ram_reg[2][19]  ( .CLK(n300), .D(N35), .Q(\ram[2][19] ) );
  LATCHX1_HVT \ram_reg[2][18]  ( .CLK(n308), .D(N34), .Q(\ram[2][18] ) );
  LATCHX1_HVT \ram_reg[2][17]  ( .CLK(n309), .D(N33), .Q(\ram[2][17] ) );
  LATCHX1_HVT \ram_reg[2][16]  ( .CLK(n309), .D(N32), .Q(\ram[2][16] ) );
  LATCHX1_HVT \ram_reg[2][15]  ( .CLK(n303), .D(N31), .Q(\ram[2][15] ) );
  LATCHX1_HVT \ram_reg[2][14]  ( .CLK(n303), .D(N30), .Q(\ram[2][14] ) );
  LATCHX1_HVT \ram_reg[2][13]  ( .CLK(n302), .D(N29), .Q(\ram[2][13] ) );
  LATCHX1_HVT \ram_reg[2][12]  ( .CLK(n302), .D(N28), .Q(\ram[2][12] ) );
  LATCHX1_HVT \ram_reg[2][11]  ( .CLK(n303), .D(N27), .Q(\ram[2][11] ) );
  LATCHX1_HVT \ram_reg[2][10]  ( .CLK(n302), .D(N26), .Q(\ram[2][10] ) );
  LATCHX1_HVT \ram_reg[2][9]  ( .CLK(n302), .D(N25), .Q(\ram[2][9] ) );
  LATCHX1_HVT \ram_reg[2][8]  ( .CLK(n303), .D(N24), .Q(\ram[2][8] ) );
  LATCHX1_HVT \ram_reg[2][7]  ( .CLK(n306), .D(N23), .Q(\ram[2][7] ) );
  LATCHX1_HVT \ram_reg[2][6]  ( .CLK(n306), .D(N22), .Q(\ram[2][6] ) );
  LATCHX1_HVT \ram_reg[2][5]  ( .CLK(n305), .D(N21), .Q(\ram[2][5] ) );
  LATCHX1_HVT \ram_reg[2][4]  ( .CLK(n305), .D(N20), .Q(\ram[2][4] ) );
  LATCHX1_HVT \ram_reg[2][3]  ( .CLK(n304), .D(N19), .Q(\ram[2][3] ) );
  LATCHX1_HVT \ram_reg[2][2]  ( .CLK(n305), .D(N18), .Q(\ram[2][2] ) );
  LATCHX1_HVT \ram_reg[2][1]  ( .CLK(n306), .D(N17), .Q(\ram[2][1] ) );
  LATCHX1_HVT \ram_reg[2][0]  ( .CLK(n310), .D(N16), .Q(\ram[2][0] ) );
  LATCHX1_HVT \ram_reg[1][255]  ( .CLK(N276), .D(N273), .Q(\ram[1][255] ) );
  LATCHX1_HVT \ram_reg[1][254]  ( .CLK(N276), .D(N272), .Q(\ram[1][254] ) );
  LATCHX1_HVT \ram_reg[1][253]  ( .CLK(N276), .D(N271), .Q(\ram[1][253] ) );
  LATCHX1_HVT \ram_reg[1][252]  ( .CLK(N276), .D(N270), .Q(\ram[1][252] ) );
  LATCHX1_HVT \ram_reg[1][251]  ( .CLK(n343), .D(N269), .Q(\ram[1][251] ) );
  LATCHX1_HVT \ram_reg[1][250]  ( .CLK(n335), .D(N268), .Q(\ram[1][250] ) );
  LATCHX1_HVT \ram_reg[1][249]  ( .CLK(n335), .D(N267), .Q(\ram[1][249] ) );
  LATCHX1_HVT \ram_reg[1][248]  ( .CLK(n335), .D(N266), .Q(\ram[1][248] ) );
  LATCHX1_HVT \ram_reg[1][247]  ( .CLK(n335), .D(N265), .Q(\ram[1][247] ) );
  LATCHX1_HVT \ram_reg[1][246]  ( .CLK(n335), .D(N264), .Q(\ram[1][246] ) );
  LATCHX1_HVT \ram_reg[1][245]  ( .CLK(n335), .D(N263), .Q(\ram[1][245] ) );
  LATCHX1_HVT \ram_reg[1][244]  ( .CLK(n335), .D(N262), .Q(\ram[1][244] ) );
  LATCHX1_HVT \ram_reg[1][243]  ( .CLK(n335), .D(N261), .Q(\ram[1][243] ) );
  LATCHX1_HVT \ram_reg[1][242]  ( .CLK(n335), .D(N260), .Q(\ram[1][242] ) );
  LATCHX1_HVT \ram_reg[1][241]  ( .CLK(n334), .D(N259), .Q(\ram[1][241] ) );
  LATCHX1_HVT \ram_reg[1][240]  ( .CLK(n334), .D(N258), .Q(\ram[1][240] ) );
  LATCHX1_HVT \ram_reg[1][239]  ( .CLK(n334), .D(N257), .Q(\ram[1][239] ) );
  LATCHX1_HVT \ram_reg[1][238]  ( .CLK(n334), .D(N256), .Q(\ram[1][238] ) );
  LATCHX1_HVT \ram_reg[1][237]  ( .CLK(n334), .D(N255), .Q(\ram[1][237] ) );
  LATCHX1_HVT \ram_reg[1][236]  ( .CLK(n334), .D(N254), .Q(\ram[1][236] ) );
  LATCHX1_HVT \ram_reg[1][235]  ( .CLK(n334), .D(N253), .Q(\ram[1][235] ) );
  LATCHX1_HVT \ram_reg[1][234]  ( .CLK(n334), .D(N252), .Q(\ram[1][234] ) );
  LATCHX1_HVT \ram_reg[1][233]  ( .CLK(n334), .D(N251), .Q(\ram[1][233] ) );
  LATCHX1_HVT \ram_reg[1][232]  ( .CLK(n334), .D(N250), .Q(\ram[1][232] ) );
  LATCHX1_HVT \ram_reg[1][231]  ( .CLK(n334), .D(N249), .Q(\ram[1][231] ) );
  LATCHX1_HVT \ram_reg[1][230]  ( .CLK(n333), .D(N248), .Q(\ram[1][230] ) );
  LATCHX1_HVT \ram_reg[1][229]  ( .CLK(n333), .D(N247), .Q(\ram[1][229] ) );
  LATCHX1_HVT \ram_reg[1][228]  ( .CLK(n333), .D(N246), .Q(\ram[1][228] ) );
  LATCHX1_HVT \ram_reg[1][227]  ( .CLK(n343), .D(N245), .Q(\ram[1][227] ) );
  LATCHX1_HVT \ram_reg[1][226]  ( .CLK(n343), .D(N244), .Q(\ram[1][226] ) );
  LATCHX1_HVT \ram_reg[1][225]  ( .CLK(n343), .D(N243), .Q(\ram[1][225] ) );
  LATCHX1_HVT \ram_reg[1][224]  ( .CLK(n343), .D(N242), .Q(\ram[1][224] ) );
  LATCHX1_HVT \ram_reg[1][223]  ( .CLK(n343), .D(N241), .Q(\ram[1][223] ) );
  LATCHX1_HVT \ram_reg[1][222]  ( .CLK(n343), .D(N240), .Q(\ram[1][222] ) );
  LATCHX1_HVT \ram_reg[1][221]  ( .CLK(n343), .D(N239), .Q(\ram[1][221] ) );
  LATCHX1_HVT \ram_reg[1][220]  ( .CLK(n343), .D(N238), .Q(\ram[1][220] ) );
  LATCHX1_HVT \ram_reg[1][219]  ( .CLK(n343), .D(N237), .Q(\ram[1][219] ) );
  LATCHX1_HVT \ram_reg[1][218]  ( .CLK(n343), .D(N236), .Q(\ram[1][218] ) );
  LATCHX1_HVT \ram_reg[1][217]  ( .CLK(n342), .D(N235), .Q(\ram[1][217] ) );
  LATCHX1_HVT \ram_reg[1][216]  ( .CLK(n342), .D(N234), .Q(\ram[1][216] ) );
  LATCHX1_HVT \ram_reg[1][215]  ( .CLK(n342), .D(N233), .Q(\ram[1][215] ) );
  LATCHX1_HVT \ram_reg[1][214]  ( .CLK(n342), .D(N232), .Q(\ram[1][214] ) );
  LATCHX1_HVT \ram_reg[1][213]  ( .CLK(n342), .D(N231), .Q(\ram[1][213] ) );
  LATCHX1_HVT \ram_reg[1][212]  ( .CLK(n342), .D(N230), .Q(\ram[1][212] ) );
  LATCHX1_HVT \ram_reg[1][211]  ( .CLK(n342), .D(N229), .Q(\ram[1][211] ) );
  LATCHX1_HVT \ram_reg[1][210]  ( .CLK(n342), .D(N228), .Q(\ram[1][210] ) );
  LATCHX1_HVT \ram_reg[1][209]  ( .CLK(n342), .D(N227), .Q(\ram[1][209] ) );
  LATCHX1_HVT \ram_reg[1][208]  ( .CLK(n342), .D(N226), .Q(\ram[1][208] ) );
  LATCHX1_HVT \ram_reg[1][207]  ( .CLK(n341), .D(N225), .Q(\ram[1][207] ) );
  LATCHX1_HVT \ram_reg[1][206]  ( .CLK(n341), .D(N224), .Q(\ram[1][206] ) );
  LATCHX1_HVT \ram_reg[1][205]  ( .CLK(n341), .D(N223), .Q(\ram[1][205] ) );
  LATCHX1_HVT \ram_reg[1][204]  ( .CLK(n341), .D(N222), .Q(\ram[1][204] ) );
  LATCHX1_HVT \ram_reg[1][203]  ( .CLK(n341), .D(N221), .Q(\ram[1][203] ) );
  LATCHX1_HVT \ram_reg[1][202]  ( .CLK(n341), .D(N220), .Q(\ram[1][202] ) );
  LATCHX1_HVT \ram_reg[1][201]  ( .CLK(n341), .D(N219), .Q(\ram[1][201] ) );
  LATCHX1_HVT \ram_reg[1][200]  ( .CLK(n341), .D(N218), .Q(\ram[1][200] ) );
  LATCHX1_HVT \ram_reg[1][199]  ( .CLK(n341), .D(N217), .Q(\ram[1][199] ) );
  LATCHX1_HVT \ram_reg[1][198]  ( .CLK(n341), .D(N216), .Q(\ram[1][198] ) );
  LATCHX1_HVT \ram_reg[1][197]  ( .CLK(n341), .D(N214), .Q(\ram[1][197] ) );
  LATCHX1_HVT \ram_reg[1][196]  ( .CLK(n340), .D(N213), .Q(\ram[1][196] ) );
  LATCHX1_HVT \ram_reg[1][195]  ( .CLK(n340), .D(N212), .Q(\ram[1][195] ) );
  LATCHX1_HVT \ram_reg[1][194]  ( .CLK(n340), .D(N211), .Q(\ram[1][194] ) );
  LATCHX1_HVT \ram_reg[1][193]  ( .CLK(n340), .D(N210), .Q(\ram[1][193] ) );
  LATCHX1_HVT \ram_reg[1][192]  ( .CLK(n340), .D(N209), .Q(\ram[1][192] ) );
  LATCHX1_HVT \ram_reg[1][191]  ( .CLK(n340), .D(N208), .Q(\ram[1][191] ) );
  LATCHX1_HVT \ram_reg[1][190]  ( .CLK(n340), .D(N207), .Q(\ram[1][190] ) );
  LATCHX1_HVT \ram_reg[1][189]  ( .CLK(n340), .D(N206), .Q(\ram[1][189] ) );
  LATCHX1_HVT \ram_reg[1][188]  ( .CLK(n340), .D(N205), .Q(\ram[1][188] ) );
  LATCHX1_HVT \ram_reg[1][187]  ( .CLK(n340), .D(N204), .Q(\ram[1][187] ) );
  LATCHX1_HVT \ram_reg[1][186]  ( .CLK(n340), .D(N203), .Q(\ram[1][186] ) );
  LATCHX1_HVT \ram_reg[1][185]  ( .CLK(n339), .D(N202), .Q(\ram[1][185] ) );
  LATCHX1_HVT \ram_reg[1][184]  ( .CLK(n339), .D(N201), .Q(\ram[1][184] ) );
  LATCHX1_HVT \ram_reg[1][183]  ( .CLK(n339), .D(N200), .Q(\ram[1][183] ) );
  LATCHX1_HVT \ram_reg[1][182]  ( .CLK(n339), .D(N199), .Q(\ram[1][182] ) );
  LATCHX1_HVT \ram_reg[1][181]  ( .CLK(n339), .D(N198), .Q(\ram[1][181] ) );
  LATCHX1_HVT \ram_reg[1][180]  ( .CLK(n339), .D(N197), .Q(\ram[1][180] ) );
  LATCHX1_HVT \ram_reg[1][179]  ( .CLK(n339), .D(N196), .Q(\ram[1][179] ) );
  LATCHX1_HVT \ram_reg[1][178]  ( .CLK(n339), .D(N195), .Q(\ram[1][178] ) );
  LATCHX1_HVT \ram_reg[1][177]  ( .CLK(n339), .D(N194), .Q(\ram[1][177] ) );
  LATCHX1_HVT \ram_reg[1][176]  ( .CLK(n339), .D(N193), .Q(\ram[1][176] ) );
  LATCHX1_HVT \ram_reg[1][175]  ( .CLK(n339), .D(N192), .Q(\ram[1][175] ) );
  LATCHX1_HVT \ram_reg[1][174]  ( .CLK(n338), .D(N191), .Q(\ram[1][174] ) );
  LATCHX1_HVT \ram_reg[1][173]  ( .CLK(n338), .D(N190), .Q(\ram[1][173] ) );
  LATCHX1_HVT \ram_reg[1][172]  ( .CLK(n338), .D(N189), .Q(\ram[1][172] ) );
  LATCHX1_HVT \ram_reg[1][171]  ( .CLK(n338), .D(N188), .Q(\ram[1][171] ) );
  LATCHX1_HVT \ram_reg[1][170]  ( .CLK(n338), .D(N187), .Q(\ram[1][170] ) );
  LATCHX1_HVT \ram_reg[1][169]  ( .CLK(n338), .D(N186), .Q(\ram[1][169] ) );
  LATCHX1_HVT \ram_reg[1][168]  ( .CLK(n338), .D(N185), .Q(\ram[1][168] ) );
  LATCHX1_HVT \ram_reg[1][167]  ( .CLK(n338), .D(N184), .Q(\ram[1][167] ) );
  LATCHX1_HVT \ram_reg[1][166]  ( .CLK(n338), .D(N183), .Q(\ram[1][166] ) );
  LATCHX1_HVT \ram_reg[1][165]  ( .CLK(n338), .D(N182), .Q(\ram[1][165] ) );
  LATCHX1_HVT \ram_reg[1][164]  ( .CLK(n338), .D(N181), .Q(\ram[1][164] ) );
  LATCHX1_HVT \ram_reg[1][163]  ( .CLK(n337), .D(N180), .Q(\ram[1][163] ) );
  LATCHX1_HVT \ram_reg[1][162]  ( .CLK(n337), .D(N179), .Q(\ram[1][162] ) );
  LATCHX1_HVT \ram_reg[1][161]  ( .CLK(n337), .D(N178), .Q(\ram[1][161] ) );
  LATCHX1_HVT \ram_reg[1][160]  ( .CLK(n337), .D(N177), .Q(\ram[1][160] ) );
  LATCHX1_HVT \ram_reg[1][159]  ( .CLK(n337), .D(N176), .Q(\ram[1][159] ) );
  LATCHX1_HVT \ram_reg[1][158]  ( .CLK(n337), .D(N175), .Q(\ram[1][158] ) );
  LATCHX1_HVT \ram_reg[1][157]  ( .CLK(n337), .D(N174), .Q(\ram[1][157] ) );
  LATCHX1_HVT \ram_reg[1][156]  ( .CLK(n337), .D(N173), .Q(\ram[1][156] ) );
  LATCHX1_HVT \ram_reg[1][155]  ( .CLK(n337), .D(N172), .Q(\ram[1][155] ) );
  LATCHX1_HVT \ram_reg[1][154]  ( .CLK(n337), .D(N171), .Q(\ram[1][154] ) );
  LATCHX1_HVT \ram_reg[1][153]  ( .CLK(n337), .D(N170), .Q(\ram[1][153] ) );
  LATCHX1_HVT \ram_reg[1][152]  ( .CLK(n336), .D(N169), .Q(\ram[1][152] ) );
  LATCHX1_HVT \ram_reg[1][151]  ( .CLK(n336), .D(N168), .Q(\ram[1][151] ) );
  LATCHX1_HVT \ram_reg[1][150]  ( .CLK(n336), .D(N167), .Q(\ram[1][150] ) );
  LATCHX1_HVT \ram_reg[1][149]  ( .CLK(n336), .D(N166), .Q(\ram[1][149] ) );
  LATCHX1_HVT \ram_reg[1][148]  ( .CLK(n336), .D(N165), .Q(\ram[1][148] ) );
  LATCHX1_HVT \ram_reg[1][147]  ( .CLK(n336), .D(N164), .Q(\ram[1][147] ) );
  LATCHX1_HVT \ram_reg[1][146]  ( .CLK(n336), .D(N163), .Q(\ram[1][146] ) );
  LATCHX1_HVT \ram_reg[1][145]  ( .CLK(n336), .D(N162), .Q(\ram[1][145] ) );
  LATCHX1_HVT \ram_reg[1][144]  ( .CLK(n336), .D(N161), .Q(\ram[1][144] ) );
  LATCHX1_HVT \ram_reg[1][143]  ( .CLK(n336), .D(N160), .Q(\ram[1][143] ) );
  LATCHX1_HVT \ram_reg[1][142]  ( .CLK(n336), .D(N159), .Q(\ram[1][142] ) );
  LATCHX1_HVT \ram_reg[1][141]  ( .CLK(n335), .D(N158), .Q(\ram[1][141] ) );
  LATCHX1_HVT \ram_reg[1][140]  ( .CLK(n335), .D(N157), .Q(\ram[1][140] ) );
  LATCHX1_HVT \ram_reg[1][139]  ( .CLK(n335), .D(N156), .Q(\ram[1][139] ) );
  LATCHX1_HVT \ram_reg[1][138]  ( .CLK(n334), .D(N155), .Q(\ram[1][138] ) );
  LATCHX1_HVT \ram_reg[1][137]  ( .CLK(n343), .D(N154), .Q(\ram[1][137] ) );
  LATCHX1_HVT \ram_reg[1][136]  ( .CLK(n342), .D(N153), .Q(\ram[1][136] ) );
  LATCHX1_HVT \ram_reg[1][135]  ( .CLK(n342), .D(N152), .Q(\ram[1][135] ) );
  LATCHX1_HVT \ram_reg[1][134]  ( .CLK(n341), .D(N151), .Q(\ram[1][134] ) );
  LATCHX1_HVT \ram_reg[1][133]  ( .CLK(n340), .D(N150), .Q(\ram[1][133] ) );
  LATCHX1_HVT \ram_reg[1][132]  ( .CLK(n339), .D(N149), .Q(\ram[1][132] ) );
  LATCHX1_HVT \ram_reg[1][131]  ( .CLK(n338), .D(N148), .Q(\ram[1][131] ) );
  LATCHX1_HVT \ram_reg[1][130]  ( .CLK(n337), .D(N147), .Q(\ram[1][130] ) );
  LATCHX1_HVT \ram_reg[1][129]  ( .CLK(n336), .D(N146), .Q(\ram[1][129] ) );
  LATCHX1_HVT \ram_reg[1][128]  ( .CLK(n333), .D(N145), .Q(\ram[1][128] ) );
  LATCHX1_HVT \ram_reg[1][127]  ( .CLK(n324), .D(N144), .Q(\ram[1][127] ) );
  LATCHX1_HVT \ram_reg[1][126]  ( .CLK(n324), .D(N143), .Q(\ram[1][126] ) );
  LATCHX1_HVT \ram_reg[1][125]  ( .CLK(n324), .D(N142), .Q(\ram[1][125] ) );
  LATCHX1_HVT \ram_reg[1][124]  ( .CLK(n324), .D(N141), .Q(\ram[1][124] ) );
  LATCHX1_HVT \ram_reg[1][123]  ( .CLK(n324), .D(N140), .Q(\ram[1][123] ) );
  LATCHX1_HVT \ram_reg[1][122]  ( .CLK(n323), .D(N139), .Q(\ram[1][122] ) );
  LATCHX1_HVT \ram_reg[1][121]  ( .CLK(n324), .D(N138), .Q(\ram[1][121] ) );
  LATCHX1_HVT \ram_reg[1][120]  ( .CLK(n324), .D(N137), .Q(\ram[1][120] ) );
  LATCHX1_HVT \ram_reg[1][119]  ( .CLK(n333), .D(N136), .Q(\ram[1][119] ) );
  LATCHX1_HVT \ram_reg[1][118]  ( .CLK(n332), .D(N135), .Q(\ram[1][118] ) );
  LATCHX1_HVT \ram_reg[1][117]  ( .CLK(n332), .D(N134), .Q(\ram[1][117] ) );
  LATCHX1_HVT \ram_reg[1][116]  ( .CLK(n331), .D(N133), .Q(\ram[1][116] ) );
  LATCHX1_HVT \ram_reg[1][115]  ( .CLK(n326), .D(N132), .Q(\ram[1][115] ) );
  LATCHX1_HVT \ram_reg[1][114]  ( .CLK(n331), .D(N131), .Q(\ram[1][114] ) );
  LATCHX1_HVT \ram_reg[1][113]  ( .CLK(n331), .D(N130), .Q(\ram[1][113] ) );
  LATCHX1_HVT \ram_reg[1][112]  ( .CLK(n332), .D(N129), .Q(\ram[1][112] ) );
  LATCHX1_HVT \ram_reg[1][111]  ( .CLK(n330), .D(N128), .Q(\ram[1][111] ) );
  LATCHX1_HVT \ram_reg[1][110]  ( .CLK(n330), .D(N127), .Q(\ram[1][110] ) );
  LATCHX1_HVT \ram_reg[1][109]  ( .CLK(n330), .D(N126), .Q(\ram[1][109] ) );
  LATCHX1_HVT \ram_reg[1][108]  ( .CLK(n327), .D(N125), .Q(\ram[1][108] ) );
  LATCHX1_HVT \ram_reg[1][107]  ( .CLK(n324), .D(N124), .Q(\ram[1][107] ) );
  LATCHX1_HVT \ram_reg[1][106]  ( .CLK(n330), .D(N123), .Q(\ram[1][106] ) );
  LATCHX1_HVT \ram_reg[1][105]  ( .CLK(n330), .D(N122), .Q(\ram[1][105] ) );
  LATCHX1_HVT \ram_reg[1][104]  ( .CLK(n330), .D(N121), .Q(\ram[1][104] ) );
  LATCHX1_HVT \ram_reg[1][103]  ( .CLK(n329), .D(N120), .Q(\ram[1][103] ) );
  LATCHX1_HVT \ram_reg[1][102]  ( .CLK(n328), .D(N119), .Q(\ram[1][102] ) );
  LATCHX1_HVT \ram_reg[1][101]  ( .CLK(n328), .D(N118), .Q(\ram[1][101] ) );
  LATCHX1_HVT \ram_reg[1][100]  ( .CLK(n329), .D(N117), .Q(\ram[1][100] ) );
  LATCHX1_HVT \ram_reg[1][99]  ( .CLK(n327), .D(N116), .Q(\ram[1][99] ) );
  LATCHX1_HVT \ram_reg[1][98]  ( .CLK(n328), .D(N114), .Q(\ram[1][98] ) );
  LATCHX1_HVT \ram_reg[1][97]  ( .CLK(n329), .D(N113), .Q(\ram[1][97] ) );
  LATCHX1_HVT \ram_reg[1][96]  ( .CLK(n333), .D(N112), .Q(\ram[1][96] ) );
  LATCHX1_HVT \ram_reg[1][95]  ( .CLK(n325), .D(N111), .Q(\ram[1][95] ) );
  LATCHX1_HVT \ram_reg[1][94]  ( .CLK(n325), .D(N110), .Q(\ram[1][94] ) );
  LATCHX1_HVT \ram_reg[1][93]  ( .CLK(n325), .D(N109), .Q(\ram[1][93] ) );
  LATCHX1_HVT \ram_reg[1][92]  ( .CLK(n324), .D(N108), .Q(\ram[1][92] ) );
  LATCHX1_HVT \ram_reg[1][91]  ( .CLK(n324), .D(N107), .Q(\ram[1][91] ) );
  LATCHX1_HVT \ram_reg[1][90]  ( .CLK(n325), .D(N106), .Q(\ram[1][90] ) );
  LATCHX1_HVT \ram_reg[1][89]  ( .CLK(n324), .D(N105), .Q(\ram[1][89] ) );
  LATCHX1_HVT \ram_reg[1][88]  ( .CLK(n325), .D(N104), .Q(\ram[1][88] ) );
  LATCHX1_HVT \ram_reg[1][87]  ( .CLK(n333), .D(N103), .Q(\ram[1][87] ) );
  LATCHX1_HVT \ram_reg[1][86]  ( .CLK(n332), .D(N102), .Q(\ram[1][86] ) );
  LATCHX1_HVT \ram_reg[1][85]  ( .CLK(n331), .D(N101), .Q(\ram[1][85] ) );
  LATCHX1_HVT \ram_reg[1][84]  ( .CLK(n331), .D(N100), .Q(\ram[1][84] ) );
  LATCHX1_HVT \ram_reg[1][83]  ( .CLK(n326), .D(N99), .Q(\ram[1][83] ) );
  LATCHX1_HVT \ram_reg[1][82]  ( .CLK(n332), .D(N98), .Q(\ram[1][82] ) );
  LATCHX1_HVT \ram_reg[1][81]  ( .CLK(n331), .D(N97), .Q(\ram[1][81] ) );
  LATCHX1_HVT \ram_reg[1][80]  ( .CLK(n332), .D(N96), .Q(\ram[1][80] ) );
  LATCHX1_HVT \ram_reg[1][79]  ( .CLK(n326), .D(N95), .Q(\ram[1][79] ) );
  LATCHX1_HVT \ram_reg[1][78]  ( .CLK(n325), .D(N94), .Q(\ram[1][78] ) );
  LATCHX1_HVT \ram_reg[1][77]  ( .CLK(n326), .D(N93), .Q(\ram[1][77] ) );
  LATCHX1_HVT \ram_reg[1][76]  ( .CLK(n325), .D(N92), .Q(\ram[1][76] ) );
  LATCHX1_HVT \ram_reg[1][75]  ( .CLK(n325), .D(N91), .Q(\ram[1][75] ) );
  LATCHX1_HVT \ram_reg[1][74]  ( .CLK(n323), .D(N90), .Q(\ram[1][74] ) );
  LATCHX1_HVT \ram_reg[1][73]  ( .CLK(n326), .D(N89), .Q(\ram[1][73] ) );
  LATCHX1_HVT \ram_reg[1][72]  ( .CLK(n326), .D(N88), .Q(\ram[1][72] ) );
  LATCHX1_HVT \ram_reg[1][71]  ( .CLK(n329), .D(N87), .Q(\ram[1][71] ) );
  LATCHX1_HVT \ram_reg[1][70]  ( .CLK(n329), .D(N86), .Q(\ram[1][70] ) );
  LATCHX1_HVT \ram_reg[1][69]  ( .CLK(n328), .D(N85), .Q(\ram[1][69] ) );
  LATCHX1_HVT \ram_reg[1][68]  ( .CLK(n329), .D(N84), .Q(\ram[1][68] ) );
  LATCHX1_HVT \ram_reg[1][67]  ( .CLK(n328), .D(N83), .Q(\ram[1][67] ) );
  LATCHX1_HVT \ram_reg[1][66]  ( .CLK(n327), .D(N82), .Q(\ram[1][66] ) );
  LATCHX1_HVT \ram_reg[1][65]  ( .CLK(n328), .D(N81), .Q(\ram[1][65] ) );
  LATCHX1_HVT \ram_reg[1][64]  ( .CLK(n333), .D(N80), .Q(\ram[1][64] ) );
  LATCHX1_HVT \ram_reg[1][63]  ( .CLK(n327), .D(N79), .Q(\ram[1][63] ) );
  LATCHX1_HVT \ram_reg[1][62]  ( .CLK(n327), .D(N78), .Q(\ram[1][62] ) );
  LATCHX1_HVT \ram_reg[1][61]  ( .CLK(n327), .D(N77), .Q(\ram[1][61] ) );
  LATCHX1_HVT \ram_reg[1][60]  ( .CLK(n327), .D(N76), .Q(\ram[1][60] ) );
  LATCHX1_HVT \ram_reg[1][59]  ( .CLK(n327), .D(N75), .Q(\ram[1][59] ) );
  LATCHX1_HVT \ram_reg[1][58]  ( .CLK(n326), .D(N74), .Q(\ram[1][58] ) );
  LATCHX1_HVT \ram_reg[1][57]  ( .CLK(n327), .D(N73), .Q(\ram[1][57] ) );
  LATCHX1_HVT \ram_reg[1][56]  ( .CLK(n327), .D(N72), .Q(\ram[1][56] ) );
  LATCHX1_HVT \ram_reg[1][55]  ( .CLK(n333), .D(N71), .Q(\ram[1][55] ) );
  LATCHX1_HVT \ram_reg[1][54]  ( .CLK(n331), .D(N70), .Q(\ram[1][54] ) );
  LATCHX1_HVT \ram_reg[1][53]  ( .CLK(n331), .D(N69), .Q(\ram[1][53] ) );
  LATCHX1_HVT \ram_reg[1][52]  ( .CLK(n332), .D(N68), .Q(\ram[1][52] ) );
  LATCHX1_HVT \ram_reg[1][51]  ( .CLK(n326), .D(N67), .Q(\ram[1][51] ) );
  LATCHX1_HVT \ram_reg[1][50]  ( .CLK(n323), .D(N66), .Q(\ram[1][50] ) );
  LATCHX1_HVT \ram_reg[1][49]  ( .CLK(n332), .D(N65), .Q(\ram[1][49] ) );
  LATCHX1_HVT \ram_reg[1][48]  ( .CLK(n332), .D(N64), .Q(\ram[1][48] ) );
  LATCHX1_HVT \ram_reg[1][47]  ( .CLK(n330), .D(N63), .Q(\ram[1][47] ) );
  LATCHX1_HVT \ram_reg[1][46]  ( .CLK(n330), .D(N62), .Q(\ram[1][46] ) );
  LATCHX1_HVT \ram_reg[1][45]  ( .CLK(n330), .D(N61), .Q(\ram[1][45] ) );
  LATCHX1_HVT \ram_reg[1][44]  ( .CLK(n330), .D(N60), .Q(\ram[1][44] ) );
  LATCHX1_HVT \ram_reg[1][43]  ( .CLK(n327), .D(N59), .Q(\ram[1][43] ) );
  LATCHX1_HVT \ram_reg[1][42]  ( .CLK(n331), .D(N58), .Q(\ram[1][42] ) );
  LATCHX1_HVT \ram_reg[1][41]  ( .CLK(n324), .D(N57), .Q(\ram[1][41] ) );
  LATCHX1_HVT \ram_reg[1][40]  ( .CLK(n330), .D(N56), .Q(\ram[1][40] ) );
  LATCHX1_HVT \ram_reg[1][39]  ( .CLK(n329), .D(N55), .Q(\ram[1][39] ) );
  LATCHX1_HVT \ram_reg[1][38]  ( .CLK(n329), .D(N54), .Q(\ram[1][38] ) );
  LATCHX1_HVT \ram_reg[1][37]  ( .CLK(n328), .D(N53), .Q(\ram[1][37] ) );
  LATCHX1_HVT \ram_reg[1][36]  ( .CLK(n328), .D(N52), .Q(\ram[1][36] ) );
  LATCHX1_HVT \ram_reg[1][35]  ( .CLK(n328), .D(N51), .Q(\ram[1][35] ) );
  LATCHX1_HVT \ram_reg[1][34]  ( .CLK(n330), .D(N50), .Q(\ram[1][34] ) );
  LATCHX1_HVT \ram_reg[1][33]  ( .CLK(n329), .D(N49), .Q(\ram[1][33] ) );
  LATCHX1_HVT \ram_reg[1][32]  ( .CLK(n333), .D(N48), .Q(\ram[1][32] ) );
  LATCHX1_HVT \ram_reg[1][31]  ( .CLK(n323), .D(N47), .Q(\ram[1][31] ) );
  LATCHX1_HVT \ram_reg[1][30]  ( .CLK(n323), .D(N46), .Q(\ram[1][30] ) );
  LATCHX1_HVT \ram_reg[1][29]  ( .CLK(n323), .D(N45), .Q(\ram[1][29] ) );
  LATCHX1_HVT \ram_reg[1][28]  ( .CLK(n323), .D(N44), .Q(\ram[1][28] ) );
  LATCHX1_HVT \ram_reg[1][27]  ( .CLK(n323), .D(N43), .Q(\ram[1][27] ) );
  LATCHX1_HVT \ram_reg[1][26]  ( .CLK(n323), .D(N42), .Q(\ram[1][26] ) );
  LATCHX1_HVT \ram_reg[1][25]  ( .CLK(n323), .D(N41), .Q(\ram[1][25] ) );
  LATCHX1_HVT \ram_reg[1][24]  ( .CLK(n323), .D(N40), .Q(\ram[1][24] ) );
  LATCHX1_HVT \ram_reg[1][23]  ( .CLK(n333), .D(N39), .Q(\ram[1][23] ) );
  LATCHX1_HVT \ram_reg[1][22]  ( .CLK(n332), .D(N38), .Q(\ram[1][22] ) );
  LATCHX1_HVT \ram_reg[1][21]  ( .CLK(n331), .D(N37), .Q(\ram[1][21] ) );
  LATCHX1_HVT \ram_reg[1][20]  ( .CLK(n331), .D(N36), .Q(\ram[1][20] ) );
  LATCHX1_HVT \ram_reg[1][19]  ( .CLK(n323), .D(N35), .Q(\ram[1][19] ) );
  LATCHX1_HVT \ram_reg[1][18]  ( .CLK(n331), .D(N34), .Q(\ram[1][18] ) );
  LATCHX1_HVT \ram_reg[1][17]  ( .CLK(n332), .D(N33), .Q(\ram[1][17] ) );
  LATCHX1_HVT \ram_reg[1][16]  ( .CLK(n332), .D(N32), .Q(\ram[1][16] ) );
  LATCHX1_HVT \ram_reg[1][15]  ( .CLK(n326), .D(N31), .Q(\ram[1][15] ) );
  LATCHX1_HVT \ram_reg[1][14]  ( .CLK(n326), .D(N30), .Q(\ram[1][14] ) );
  LATCHX1_HVT \ram_reg[1][13]  ( .CLK(n325), .D(N29), .Q(\ram[1][13] ) );
  LATCHX1_HVT \ram_reg[1][12]  ( .CLK(n325), .D(N28), .Q(\ram[1][12] ) );
  LATCHX1_HVT \ram_reg[1][11]  ( .CLK(n326), .D(N27), .Q(\ram[1][11] ) );
  LATCHX1_HVT \ram_reg[1][10]  ( .CLK(n325), .D(N26), .Q(\ram[1][10] ) );
  LATCHX1_HVT \ram_reg[1][9]  ( .CLK(n325), .D(N25), .Q(\ram[1][9] ) );
  LATCHX1_HVT \ram_reg[1][8]  ( .CLK(n326), .D(N24), .Q(\ram[1][8] ) );
  LATCHX1_HVT \ram_reg[1][7]  ( .CLK(n329), .D(N23), .Q(\ram[1][7] ) );
  LATCHX1_HVT \ram_reg[1][6]  ( .CLK(n329), .D(N22), .Q(\ram[1][6] ) );
  LATCHX1_HVT \ram_reg[1][5]  ( .CLK(n328), .D(N21), .Q(\ram[1][5] ) );
  LATCHX1_HVT \ram_reg[1][4]  ( .CLK(n328), .D(N20), .Q(\ram[1][4] ) );
  LATCHX1_HVT \ram_reg[1][3]  ( .CLK(n327), .D(N19), .Q(\ram[1][3] ) );
  LATCHX1_HVT \ram_reg[1][2]  ( .CLK(n328), .D(N18), .Q(\ram[1][2] ) );
  LATCHX1_HVT \ram_reg[1][1]  ( .CLK(n329), .D(N17), .Q(\ram[1][1] ) );
  LATCHX1_HVT \ram_reg[1][0]  ( .CLK(n333), .D(N16), .Q(\ram[1][0] ) );
  LATCHX1_HVT \ram_reg[0][255]  ( .CLK(N215), .D(N273), .Q(\ram[0][255] ) );
  LATCHX1_HVT \ram_reg[0][254]  ( .CLK(N215), .D(N272), .Q(\ram[0][254] ) );
  LATCHX1_HVT \ram_reg[0][253]  ( .CLK(N215), .D(N271), .Q(\ram[0][253] ) );
  LATCHX1_HVT \ram_reg[0][252]  ( .CLK(N215), .D(N270), .Q(\ram[0][252] ) );
  LATCHX1_HVT \ram_reg[0][251]  ( .CLK(n366), .D(N269), .Q(\ram[0][251] ) );
  LATCHX1_HVT \ram_reg[0][250]  ( .CLK(n358), .D(N268), .Q(\ram[0][250] ) );
  LATCHX1_HVT \ram_reg[0][249]  ( .CLK(n358), .D(N267), .Q(\ram[0][249] ) );
  LATCHX1_HVT \ram_reg[0][248]  ( .CLK(n358), .D(N266), .Q(\ram[0][248] ) );
  LATCHX1_HVT \ram_reg[0][247]  ( .CLK(n358), .D(N265), .Q(\ram[0][247] ) );
  LATCHX1_HVT \ram_reg[0][246]  ( .CLK(n358), .D(N264), .Q(\ram[0][246] ) );
  LATCHX1_HVT \ram_reg[0][245]  ( .CLK(n358), .D(N263), .Q(\ram[0][245] ) );
  LATCHX1_HVT \ram_reg[0][244]  ( .CLK(n358), .D(N262), .Q(\ram[0][244] ) );
  LATCHX1_HVT \ram_reg[0][243]  ( .CLK(n358), .D(N261), .Q(\ram[0][243] ) );
  LATCHX1_HVT \ram_reg[0][242]  ( .CLK(n358), .D(N260), .Q(\ram[0][242] ) );
  LATCHX1_HVT \ram_reg[0][241]  ( .CLK(n357), .D(N259), .Q(\ram[0][241] ) );
  LATCHX1_HVT \ram_reg[0][240]  ( .CLK(n357), .D(N258), .Q(\ram[0][240] ) );
  LATCHX1_HVT \ram_reg[0][239]  ( .CLK(n357), .D(N257), .Q(\ram[0][239] ) );
  LATCHX1_HVT \ram_reg[0][238]  ( .CLK(n357), .D(N256), .Q(\ram[0][238] ) );
  LATCHX1_HVT \ram_reg[0][237]  ( .CLK(n357), .D(N255), .Q(\ram[0][237] ) );
  LATCHX1_HVT \ram_reg[0][236]  ( .CLK(n357), .D(N254), .Q(\ram[0][236] ) );
  LATCHX1_HVT \ram_reg[0][235]  ( .CLK(n357), .D(N253), .Q(\ram[0][235] ) );
  LATCHX1_HVT \ram_reg[0][234]  ( .CLK(n357), .D(N252), .Q(\ram[0][234] ) );
  LATCHX1_HVT \ram_reg[0][233]  ( .CLK(n357), .D(N251), .Q(\ram[0][233] ) );
  LATCHX1_HVT \ram_reg[0][232]  ( .CLK(n357), .D(N250), .Q(\ram[0][232] ) );
  LATCHX1_HVT \ram_reg[0][231]  ( .CLK(n357), .D(N249), .Q(\ram[0][231] ) );
  LATCHX1_HVT \ram_reg[0][230]  ( .CLK(n356), .D(N248), .Q(\ram[0][230] ) );
  LATCHX1_HVT \ram_reg[0][229]  ( .CLK(n356), .D(N247), .Q(\ram[0][229] ) );
  LATCHX1_HVT \ram_reg[0][228]  ( .CLK(n356), .D(N246), .Q(\ram[0][228] ) );
  LATCHX1_HVT \ram_reg[0][227]  ( .CLK(n366), .D(N245), .Q(\ram[0][227] ) );
  LATCHX1_HVT \ram_reg[0][226]  ( .CLK(n366), .D(N244), .Q(\ram[0][226] ) );
  LATCHX1_HVT \ram_reg[0][225]  ( .CLK(n366), .D(N243), .Q(\ram[0][225] ) );
  LATCHX1_HVT \ram_reg[0][224]  ( .CLK(n366), .D(N242), .Q(\ram[0][224] ) );
  LATCHX1_HVT \ram_reg[0][223]  ( .CLK(n366), .D(N241), .Q(\ram[0][223] ) );
  LATCHX1_HVT \ram_reg[0][222]  ( .CLK(n366), .D(N240), .Q(\ram[0][222] ) );
  LATCHX1_HVT \ram_reg[0][221]  ( .CLK(n366), .D(N239), .Q(\ram[0][221] ) );
  LATCHX1_HVT \ram_reg[0][220]  ( .CLK(n366), .D(N238), .Q(\ram[0][220] ) );
  LATCHX1_HVT \ram_reg[0][219]  ( .CLK(n366), .D(N237), .Q(\ram[0][219] ) );
  LATCHX1_HVT \ram_reg[0][218]  ( .CLK(n366), .D(N236), .Q(\ram[0][218] ) );
  LATCHX1_HVT \ram_reg[0][217]  ( .CLK(n365), .D(N235), .Q(\ram[0][217] ) );
  LATCHX1_HVT \ram_reg[0][216]  ( .CLK(n365), .D(N234), .Q(\ram[0][216] ) );
  LATCHX1_HVT \ram_reg[0][215]  ( .CLK(n365), .D(N233), .Q(\ram[0][215] ) );
  LATCHX1_HVT \ram_reg[0][214]  ( .CLK(n365), .D(N232), .Q(\ram[0][214] ) );
  LATCHX1_HVT \ram_reg[0][213]  ( .CLK(n365), .D(N231), .Q(\ram[0][213] ) );
  LATCHX1_HVT \ram_reg[0][212]  ( .CLK(n365), .D(N230), .Q(\ram[0][212] ) );
  LATCHX1_HVT \ram_reg[0][211]  ( .CLK(n365), .D(N229), .Q(\ram[0][211] ) );
  LATCHX1_HVT \ram_reg[0][210]  ( .CLK(n365), .D(N228), .Q(\ram[0][210] ) );
  LATCHX1_HVT \ram_reg[0][209]  ( .CLK(n365), .D(N227), .Q(\ram[0][209] ) );
  LATCHX1_HVT \ram_reg[0][208]  ( .CLK(n365), .D(N226), .Q(\ram[0][208] ) );
  LATCHX1_HVT \ram_reg[0][207]  ( .CLK(n364), .D(N225), .Q(\ram[0][207] ) );
  LATCHX1_HVT \ram_reg[0][206]  ( .CLK(n364), .D(N224), .Q(\ram[0][206] ) );
  LATCHX1_HVT \ram_reg[0][205]  ( .CLK(n364), .D(N223), .Q(\ram[0][205] ) );
  LATCHX1_HVT \ram_reg[0][204]  ( .CLK(n364), .D(N222), .Q(\ram[0][204] ) );
  LATCHX1_HVT \ram_reg[0][203]  ( .CLK(n364), .D(N221), .Q(\ram[0][203] ) );
  LATCHX1_HVT \ram_reg[0][202]  ( .CLK(n364), .D(N220), .Q(\ram[0][202] ) );
  LATCHX1_HVT \ram_reg[0][201]  ( .CLK(n364), .D(N219), .Q(\ram[0][201] ) );
  LATCHX1_HVT \ram_reg[0][200]  ( .CLK(n364), .D(N218), .Q(\ram[0][200] ) );
  LATCHX1_HVT \ram_reg[0][199]  ( .CLK(n364), .D(N217), .Q(\ram[0][199] ) );
  LATCHX1_HVT \ram_reg[0][198]  ( .CLK(n364), .D(N216), .Q(\ram[0][198] ) );
  LATCHX1_HVT \ram_reg[0][197]  ( .CLK(n364), .D(N214), .Q(\ram[0][197] ) );
  LATCHX1_HVT \ram_reg[0][196]  ( .CLK(n363), .D(N213), .Q(\ram[0][196] ) );
  LATCHX1_HVT \ram_reg[0][195]  ( .CLK(n363), .D(N212), .Q(\ram[0][195] ) );
  LATCHX1_HVT \ram_reg[0][194]  ( .CLK(n363), .D(N211), .Q(\ram[0][194] ) );
  LATCHX1_HVT \ram_reg[0][193]  ( .CLK(n363), .D(N210), .Q(\ram[0][193] ) );
  LATCHX1_HVT \ram_reg[0][192]  ( .CLK(n363), .D(N209), .Q(\ram[0][192] ) );
  LATCHX1_HVT \ram_reg[0][191]  ( .CLK(n363), .D(N208), .Q(\ram[0][191] ) );
  LATCHX1_HVT \ram_reg[0][190]  ( .CLK(n363), .D(N207), .Q(\ram[0][190] ) );
  LATCHX1_HVT \ram_reg[0][189]  ( .CLK(n363), .D(N206), .Q(\ram[0][189] ) );
  LATCHX1_HVT \ram_reg[0][188]  ( .CLK(n363), .D(N205), .Q(\ram[0][188] ) );
  LATCHX1_HVT \ram_reg[0][187]  ( .CLK(n363), .D(N204), .Q(\ram[0][187] ) );
  LATCHX1_HVT \ram_reg[0][186]  ( .CLK(n363), .D(N203), .Q(\ram[0][186] ) );
  LATCHX1_HVT \ram_reg[0][185]  ( .CLK(n362), .D(N202), .Q(\ram[0][185] ) );
  LATCHX1_HVT \ram_reg[0][184]  ( .CLK(n362), .D(N201), .Q(\ram[0][184] ) );
  LATCHX1_HVT \ram_reg[0][183]  ( .CLK(n362), .D(N200), .Q(\ram[0][183] ) );
  LATCHX1_HVT \ram_reg[0][182]  ( .CLK(n362), .D(N199), .Q(\ram[0][182] ) );
  LATCHX1_HVT \ram_reg[0][181]  ( .CLK(n362), .D(N198), .Q(\ram[0][181] ) );
  LATCHX1_HVT \ram_reg[0][180]  ( .CLK(n362), .D(N197), .Q(\ram[0][180] ) );
  LATCHX1_HVT \ram_reg[0][179]  ( .CLK(n362), .D(N196), .Q(\ram[0][179] ) );
  LATCHX1_HVT \ram_reg[0][178]  ( .CLK(n362), .D(N195), .Q(\ram[0][178] ) );
  LATCHX1_HVT \ram_reg[0][177]  ( .CLK(n362), .D(N194), .Q(\ram[0][177] ) );
  LATCHX1_HVT \ram_reg[0][176]  ( .CLK(n362), .D(N193), .Q(\ram[0][176] ) );
  LATCHX1_HVT \ram_reg[0][175]  ( .CLK(n362), .D(N192), .Q(\ram[0][175] ) );
  LATCHX1_HVT \ram_reg[0][174]  ( .CLK(n361), .D(N191), .Q(\ram[0][174] ) );
  LATCHX1_HVT \ram_reg[0][173]  ( .CLK(n361), .D(N190), .Q(\ram[0][173] ) );
  LATCHX1_HVT \ram_reg[0][172]  ( .CLK(n361), .D(N189), .Q(\ram[0][172] ) );
  LATCHX1_HVT \ram_reg[0][171]  ( .CLK(n361), .D(N188), .Q(\ram[0][171] ) );
  LATCHX1_HVT \ram_reg[0][170]  ( .CLK(n361), .D(N187), .Q(\ram[0][170] ) );
  LATCHX1_HVT \ram_reg[0][169]  ( .CLK(n361), .D(N186), .Q(\ram[0][169] ) );
  LATCHX1_HVT \ram_reg[0][168]  ( .CLK(n361), .D(N185), .Q(\ram[0][168] ) );
  LATCHX1_HVT \ram_reg[0][167]  ( .CLK(n361), .D(N184), .Q(\ram[0][167] ) );
  LATCHX1_HVT \ram_reg[0][166]  ( .CLK(n361), .D(N183), .Q(\ram[0][166] ) );
  LATCHX1_HVT \ram_reg[0][165]  ( .CLK(n361), .D(N182), .Q(\ram[0][165] ) );
  LATCHX1_HVT \ram_reg[0][164]  ( .CLK(n361), .D(N181), .Q(\ram[0][164] ) );
  LATCHX1_HVT \ram_reg[0][163]  ( .CLK(n360), .D(N180), .Q(\ram[0][163] ) );
  LATCHX1_HVT \ram_reg[0][162]  ( .CLK(n360), .D(N179), .Q(\ram[0][162] ) );
  LATCHX1_HVT \ram_reg[0][161]  ( .CLK(n360), .D(N178), .Q(\ram[0][161] ) );
  LATCHX1_HVT \ram_reg[0][160]  ( .CLK(n360), .D(N177), .Q(\ram[0][160] ) );
  LATCHX1_HVT \ram_reg[0][159]  ( .CLK(n360), .D(N176), .Q(\ram[0][159] ) );
  LATCHX1_HVT \ram_reg[0][158]  ( .CLK(n360), .D(N175), .Q(\ram[0][158] ) );
  LATCHX1_HVT \ram_reg[0][157]  ( .CLK(n360), .D(N174), .Q(\ram[0][157] ) );
  LATCHX1_HVT \ram_reg[0][156]  ( .CLK(n360), .D(N173), .Q(\ram[0][156] ) );
  LATCHX1_HVT \ram_reg[0][155]  ( .CLK(n360), .D(N172), .Q(\ram[0][155] ) );
  LATCHX1_HVT \ram_reg[0][154]  ( .CLK(n360), .D(N171), .Q(\ram[0][154] ) );
  LATCHX1_HVT \ram_reg[0][153]  ( .CLK(n360), .D(N170), .Q(\ram[0][153] ) );
  LATCHX1_HVT \ram_reg[0][152]  ( .CLK(n359), .D(N169), .Q(\ram[0][152] ) );
  LATCHX1_HVT \ram_reg[0][151]  ( .CLK(n359), .D(N168), .Q(\ram[0][151] ) );
  LATCHX1_HVT \ram_reg[0][150]  ( .CLK(n359), .D(N167), .Q(\ram[0][150] ) );
  LATCHX1_HVT \ram_reg[0][149]  ( .CLK(n359), .D(N166), .Q(\ram[0][149] ) );
  LATCHX1_HVT \ram_reg[0][148]  ( .CLK(n359), .D(N165), .Q(\ram[0][148] ) );
  LATCHX1_HVT \ram_reg[0][147]  ( .CLK(n359), .D(N164), .Q(\ram[0][147] ) );
  LATCHX1_HVT \ram_reg[0][146]  ( .CLK(n359), .D(N163), .Q(\ram[0][146] ) );
  LATCHX1_HVT \ram_reg[0][145]  ( .CLK(n359), .D(N162), .Q(\ram[0][145] ) );
  LATCHX1_HVT \ram_reg[0][144]  ( .CLK(n359), .D(N161), .Q(\ram[0][144] ) );
  LATCHX1_HVT \ram_reg[0][143]  ( .CLK(n359), .D(N160), .Q(\ram[0][143] ) );
  LATCHX1_HVT \ram_reg[0][142]  ( .CLK(n359), .D(N159), .Q(\ram[0][142] ) );
  LATCHX1_HVT \ram_reg[0][141]  ( .CLK(n358), .D(N158), .Q(\ram[0][141] ) );
  LATCHX1_HVT \ram_reg[0][140]  ( .CLK(n358), .D(N157), .Q(\ram[0][140] ) );
  LATCHX1_HVT \ram_reg[0][139]  ( .CLK(n358), .D(N156), .Q(\ram[0][139] ) );
  LATCHX1_HVT \ram_reg[0][138]  ( .CLK(n357), .D(N155), .Q(\ram[0][138] ) );
  LATCHX1_HVT \ram_reg[0][137]  ( .CLK(n366), .D(N154), .Q(\ram[0][137] ) );
  LATCHX1_HVT \ram_reg[0][136]  ( .CLK(n365), .D(N153), .Q(\ram[0][136] ) );
  LATCHX1_HVT \ram_reg[0][135]  ( .CLK(n365), .D(N152), .Q(\ram[0][135] ) );
  LATCHX1_HVT \ram_reg[0][134]  ( .CLK(n364), .D(N151), .Q(\ram[0][134] ) );
  LATCHX1_HVT \ram_reg[0][133]  ( .CLK(n363), .D(N150), .Q(\ram[0][133] ) );
  LATCHX1_HVT \ram_reg[0][132]  ( .CLK(n362), .D(N149), .Q(\ram[0][132] ) );
  LATCHX1_HVT \ram_reg[0][131]  ( .CLK(n361), .D(N148), .Q(\ram[0][131] ) );
  LATCHX1_HVT \ram_reg[0][130]  ( .CLK(n360), .D(N147), .Q(\ram[0][130] ) );
  LATCHX1_HVT \ram_reg[0][129]  ( .CLK(n359), .D(N146), .Q(\ram[0][129] ) );
  LATCHX1_HVT \ram_reg[0][128]  ( .CLK(n356), .D(N145), .Q(\ram[0][128] ) );
  LATCHX1_HVT \ram_reg[0][127]  ( .CLK(n347), .D(N144), .Q(\ram[0][127] ) );
  LATCHX1_HVT \ram_reg[0][126]  ( .CLK(n347), .D(N143), .Q(\ram[0][126] ) );
  LATCHX1_HVT \ram_reg[0][125]  ( .CLK(n347), .D(N142), .Q(\ram[0][125] ) );
  LATCHX1_HVT \ram_reg[0][124]  ( .CLK(n347), .D(N141), .Q(\ram[0][124] ) );
  LATCHX1_HVT \ram_reg[0][123]  ( .CLK(n347), .D(N140), .Q(\ram[0][123] ) );
  LATCHX1_HVT \ram_reg[0][122]  ( .CLK(n346), .D(N139), .Q(\ram[0][122] ) );
  LATCHX1_HVT \ram_reg[0][121]  ( .CLK(n347), .D(N138), .Q(\ram[0][121] ) );
  LATCHX1_HVT \ram_reg[0][120]  ( .CLK(n347), .D(N137), .Q(\ram[0][120] ) );
  LATCHX1_HVT \ram_reg[0][119]  ( .CLK(n356), .D(N136), .Q(\ram[0][119] ) );
  LATCHX1_HVT \ram_reg[0][118]  ( .CLK(n355), .D(N135), .Q(\ram[0][118] ) );
  LATCHX1_HVT \ram_reg[0][117]  ( .CLK(n355), .D(N134), .Q(\ram[0][117] ) );
  LATCHX1_HVT \ram_reg[0][116]  ( .CLK(n354), .D(N133), .Q(\ram[0][116] ) );
  LATCHX1_HVT \ram_reg[0][115]  ( .CLK(n349), .D(N132), .Q(\ram[0][115] ) );
  LATCHX1_HVT \ram_reg[0][114]  ( .CLK(n354), .D(N131), .Q(\ram[0][114] ) );
  LATCHX1_HVT \ram_reg[0][113]  ( .CLK(n354), .D(N130), .Q(\ram[0][113] ) );
  LATCHX1_HVT \ram_reg[0][112]  ( .CLK(n355), .D(N129), .Q(\ram[0][112] ) );
  LATCHX1_HVT \ram_reg[0][111]  ( .CLK(n353), .D(N128), .Q(\ram[0][111] ) );
  LATCHX1_HVT \ram_reg[0][110]  ( .CLK(n353), .D(N127), .Q(\ram[0][110] ) );
  LATCHX1_HVT \ram_reg[0][109]  ( .CLK(n353), .D(N126), .Q(\ram[0][109] ) );
  LATCHX1_HVT \ram_reg[0][108]  ( .CLK(n350), .D(N125), .Q(\ram[0][108] ) );
  LATCHX1_HVT \ram_reg[0][107]  ( .CLK(n347), .D(N124), .Q(\ram[0][107] ) );
  LATCHX1_HVT \ram_reg[0][106]  ( .CLK(n353), .D(N123), .Q(\ram[0][106] ) );
  LATCHX1_HVT \ram_reg[0][105]  ( .CLK(n353), .D(N122), .Q(\ram[0][105] ) );
  LATCHX1_HVT \ram_reg[0][104]  ( .CLK(n353), .D(N121), .Q(\ram[0][104] ) );
  LATCHX1_HVT \ram_reg[0][103]  ( .CLK(n352), .D(N120), .Q(\ram[0][103] ) );
  LATCHX1_HVT \ram_reg[0][102]  ( .CLK(n351), .D(N119), .Q(\ram[0][102] ) );
  LATCHX1_HVT \ram_reg[0][101]  ( .CLK(n351), .D(N118), .Q(\ram[0][101] ) );
  LATCHX1_HVT \ram_reg[0][100]  ( .CLK(n352), .D(N117), .Q(\ram[0][100] ) );
  LATCHX1_HVT \ram_reg[0][99]  ( .CLK(n350), .D(N116), .Q(\ram[0][99] ) );
  LATCHX1_HVT \ram_reg[0][98]  ( .CLK(n351), .D(N114), .Q(\ram[0][98] ) );
  LATCHX1_HVT \ram_reg[0][97]  ( .CLK(n352), .D(N113), .Q(\ram[0][97] ) );
  LATCHX1_HVT \ram_reg[0][96]  ( .CLK(n356), .D(N112), .Q(\ram[0][96] ) );
  LATCHX1_HVT \ram_reg[0][95]  ( .CLK(n348), .D(N111), .Q(\ram[0][95] ) );
  LATCHX1_HVT \ram_reg[0][94]  ( .CLK(n348), .D(N110), .Q(\ram[0][94] ) );
  LATCHX1_HVT \ram_reg[0][93]  ( .CLK(n348), .D(N109), .Q(\ram[0][93] ) );
  LATCHX1_HVT \ram_reg[0][92]  ( .CLK(n347), .D(N108), .Q(\ram[0][92] ) );
  LATCHX1_HVT \ram_reg[0][91]  ( .CLK(n347), .D(N107), .Q(\ram[0][91] ) );
  LATCHX1_HVT \ram_reg[0][90]  ( .CLK(n348), .D(N106), .Q(\ram[0][90] ) );
  LATCHX1_HVT \ram_reg[0][89]  ( .CLK(n347), .D(N105), .Q(\ram[0][89] ) );
  LATCHX1_HVT \ram_reg[0][88]  ( .CLK(n348), .D(N104), .Q(\ram[0][88] ) );
  LATCHX1_HVT \ram_reg[0][87]  ( .CLK(n356), .D(N103), .Q(\ram[0][87] ) );
  LATCHX1_HVT \ram_reg[0][86]  ( .CLK(n355), .D(N102), .Q(\ram[0][86] ) );
  LATCHX1_HVT \ram_reg[0][85]  ( .CLK(n354), .D(N101), .Q(\ram[0][85] ) );
  LATCHX1_HVT \ram_reg[0][84]  ( .CLK(n354), .D(N100), .Q(\ram[0][84] ) );
  LATCHX1_HVT \ram_reg[0][83]  ( .CLK(n349), .D(N99), .Q(\ram[0][83] ) );
  LATCHX1_HVT \ram_reg[0][82]  ( .CLK(n355), .D(N98), .Q(\ram[0][82] ) );
  LATCHX1_HVT \ram_reg[0][81]  ( .CLK(n354), .D(N97), .Q(\ram[0][81] ) );
  LATCHX1_HVT \ram_reg[0][80]  ( .CLK(n355), .D(N96), .Q(\ram[0][80] ) );
  LATCHX1_HVT \ram_reg[0][79]  ( .CLK(n349), .D(N95), .Q(\ram[0][79] ) );
  LATCHX1_HVT \ram_reg[0][78]  ( .CLK(n348), .D(N94), .Q(\ram[0][78] ) );
  LATCHX1_HVT \ram_reg[0][77]  ( .CLK(n349), .D(N93), .Q(\ram[0][77] ) );
  LATCHX1_HVT \ram_reg[0][76]  ( .CLK(n348), .D(N92), .Q(\ram[0][76] ) );
  LATCHX1_HVT \ram_reg[0][75]  ( .CLK(n348), .D(N91), .Q(\ram[0][75] ) );
  LATCHX1_HVT \ram_reg[0][74]  ( .CLK(n346), .D(N90), .Q(\ram[0][74] ) );
  LATCHX1_HVT \ram_reg[0][73]  ( .CLK(n349), .D(N89), .Q(\ram[0][73] ) );
  LATCHX1_HVT \ram_reg[0][72]  ( .CLK(n349), .D(N88), .Q(\ram[0][72] ) );
  LATCHX1_HVT \ram_reg[0][71]  ( .CLK(n352), .D(N87), .Q(\ram[0][71] ) );
  LATCHX1_HVT \ram_reg[0][70]  ( .CLK(n352), .D(N86), .Q(\ram[0][70] ) );
  LATCHX1_HVT \ram_reg[0][69]  ( .CLK(n351), .D(N85), .Q(\ram[0][69] ) );
  LATCHX1_HVT \ram_reg[0][68]  ( .CLK(n352), .D(N84), .Q(\ram[0][68] ) );
  LATCHX1_HVT \ram_reg[0][67]  ( .CLK(n351), .D(N83), .Q(\ram[0][67] ) );
  LATCHX1_HVT \ram_reg[0][66]  ( .CLK(n350), .D(N82), .Q(\ram[0][66] ) );
  LATCHX1_HVT \ram_reg[0][65]  ( .CLK(n351), .D(N81), .Q(\ram[0][65] ) );
  LATCHX1_HVT \ram_reg[0][64]  ( .CLK(n356), .D(N80), .Q(\ram[0][64] ) );
  LATCHX1_HVT \ram_reg[0][63]  ( .CLK(n350), .D(N79), .Q(\ram[0][63] ) );
  LATCHX1_HVT \ram_reg[0][62]  ( .CLK(n350), .D(N78), .Q(\ram[0][62] ) );
  LATCHX1_HVT \ram_reg[0][61]  ( .CLK(n350), .D(N77), .Q(\ram[0][61] ) );
  LATCHX1_HVT \ram_reg[0][60]  ( .CLK(n350), .D(N76), .Q(\ram[0][60] ) );
  LATCHX1_HVT \ram_reg[0][59]  ( .CLK(n350), .D(N75), .Q(\ram[0][59] ) );
  LATCHX1_HVT \ram_reg[0][58]  ( .CLK(n349), .D(N74), .Q(\ram[0][58] ) );
  LATCHX1_HVT \ram_reg[0][57]  ( .CLK(n350), .D(N73), .Q(\ram[0][57] ) );
  LATCHX1_HVT \ram_reg[0][56]  ( .CLK(n350), .D(N72), .Q(\ram[0][56] ) );
  LATCHX1_HVT \ram_reg[0][55]  ( .CLK(n356), .D(N71), .Q(\ram[0][55] ) );
  LATCHX1_HVT \ram_reg[0][54]  ( .CLK(n354), .D(N70), .Q(\ram[0][54] ) );
  LATCHX1_HVT \ram_reg[0][53]  ( .CLK(n354), .D(N69), .Q(\ram[0][53] ) );
  LATCHX1_HVT \ram_reg[0][52]  ( .CLK(n355), .D(N68), .Q(\ram[0][52] ) );
  LATCHX1_HVT \ram_reg[0][51]  ( .CLK(n349), .D(N67), .Q(\ram[0][51] ) );
  LATCHX1_HVT \ram_reg[0][50]  ( .CLK(n346), .D(N66), .Q(\ram[0][50] ) );
  LATCHX1_HVT \ram_reg[0][49]  ( .CLK(n355), .D(N65), .Q(\ram[0][49] ) );
  LATCHX1_HVT \ram_reg[0][48]  ( .CLK(n355), .D(N64), .Q(\ram[0][48] ) );
  LATCHX1_HVT \ram_reg[0][47]  ( .CLK(n353), .D(N63), .Q(\ram[0][47] ) );
  LATCHX1_HVT \ram_reg[0][46]  ( .CLK(n353), .D(N62), .Q(\ram[0][46] ) );
  LATCHX1_HVT \ram_reg[0][45]  ( .CLK(n353), .D(N61), .Q(\ram[0][45] ) );
  LATCHX1_HVT \ram_reg[0][44]  ( .CLK(n353), .D(N60), .Q(\ram[0][44] ) );
  LATCHX1_HVT \ram_reg[0][43]  ( .CLK(n350), .D(N59), .Q(\ram[0][43] ) );
  LATCHX1_HVT \ram_reg[0][42]  ( .CLK(n354), .D(N58), .Q(\ram[0][42] ) );
  LATCHX1_HVT \ram_reg[0][41]  ( .CLK(n347), .D(N57), .Q(\ram[0][41] ) );
  LATCHX1_HVT \ram_reg[0][40]  ( .CLK(n353), .D(N56), .Q(\ram[0][40] ) );
  LATCHX1_HVT \ram_reg[0][39]  ( .CLK(n352), .D(N55), .Q(\ram[0][39] ) );
  LATCHX1_HVT \ram_reg[0][38]  ( .CLK(n352), .D(N54), .Q(\ram[0][38] ) );
  LATCHX1_HVT \ram_reg[0][37]  ( .CLK(n351), .D(N53), .Q(\ram[0][37] ) );
  LATCHX1_HVT \ram_reg[0][36]  ( .CLK(n351), .D(N52), .Q(\ram[0][36] ) );
  LATCHX1_HVT \ram_reg[0][35]  ( .CLK(n351), .D(N51), .Q(\ram[0][35] ) );
  LATCHX1_HVT \ram_reg[0][34]  ( .CLK(n353), .D(N50), .Q(\ram[0][34] ) );
  LATCHX1_HVT \ram_reg[0][33]  ( .CLK(n352), .D(N49), .Q(\ram[0][33] ) );
  LATCHX1_HVT \ram_reg[0][32]  ( .CLK(n356), .D(N48), .Q(\ram[0][32] ) );
  LATCHX1_HVT \ram_reg[0][31]  ( .CLK(n346), .D(N47), .Q(\ram[0][31] ) );
  LATCHX1_HVT \ram_reg[0][30]  ( .CLK(n346), .D(N46), .Q(\ram[0][30] ) );
  LATCHX1_HVT \ram_reg[0][29]  ( .CLK(n346), .D(N45), .Q(\ram[0][29] ) );
  LATCHX1_HVT \ram_reg[0][28]  ( .CLK(n346), .D(N44), .Q(\ram[0][28] ) );
  LATCHX1_HVT \ram_reg[0][27]  ( .CLK(n346), .D(N43), .Q(\ram[0][27] ) );
  LATCHX1_HVT \ram_reg[0][26]  ( .CLK(n346), .D(N42), .Q(\ram[0][26] ) );
  LATCHX1_HVT \ram_reg[0][25]  ( .CLK(n346), .D(N41), .Q(\ram[0][25] ) );
  LATCHX1_HVT \ram_reg[0][24]  ( .CLK(n346), .D(N40), .Q(\ram[0][24] ) );
  LATCHX1_HVT \ram_reg[0][23]  ( .CLK(n356), .D(N39), .Q(\ram[0][23] ) );
  LATCHX1_HVT \ram_reg[0][22]  ( .CLK(n355), .D(N38), .Q(\ram[0][22] ) );
  LATCHX1_HVT \ram_reg[0][21]  ( .CLK(n354), .D(N37), .Q(\ram[0][21] ) );
  LATCHX1_HVT \ram_reg[0][20]  ( .CLK(n354), .D(N36), .Q(\ram[0][20] ) );
  LATCHX1_HVT \ram_reg[0][19]  ( .CLK(n346), .D(N35), .Q(\ram[0][19] ) );
  LATCHX1_HVT \ram_reg[0][18]  ( .CLK(n354), .D(N34), .Q(\ram[0][18] ) );
  LATCHX1_HVT \ram_reg[0][17]  ( .CLK(n355), .D(N33), .Q(\ram[0][17] ) );
  LATCHX1_HVT \ram_reg[0][16]  ( .CLK(n355), .D(N32), .Q(\ram[0][16] ) );
  LATCHX1_HVT \ram_reg[0][15]  ( .CLK(n349), .D(N31), .Q(\ram[0][15] ) );
  LATCHX1_HVT \ram_reg[0][14]  ( .CLK(n349), .D(N30), .Q(\ram[0][14] ) );
  LATCHX1_HVT \ram_reg[0][13]  ( .CLK(n348), .D(N29), .Q(\ram[0][13] ) );
  LATCHX1_HVT \ram_reg[0][12]  ( .CLK(n348), .D(N28), .Q(\ram[0][12] ) );
  LATCHX1_HVT \ram_reg[0][11]  ( .CLK(n349), .D(N27), .Q(\ram[0][11] ) );
  LATCHX1_HVT \ram_reg[0][10]  ( .CLK(n348), .D(N26), .Q(\ram[0][10] ) );
  LATCHX1_HVT \ram_reg[0][9]  ( .CLK(n348), .D(N25), .Q(\ram[0][9] ) );
  LATCHX1_HVT \ram_reg[0][8]  ( .CLK(n349), .D(N24), .Q(\ram[0][8] ) );
  LATCHX1_HVT \ram_reg[0][7]  ( .CLK(n352), .D(N23), .Q(\ram[0][7] ) );
  LATCHX1_HVT \ram_reg[0][6]  ( .CLK(n352), .D(N22), .Q(\ram[0][6] ) );
  LATCHX1_HVT \ram_reg[0][5]  ( .CLK(n351), .D(N21), .Q(\ram[0][5] ) );
  LATCHX1_HVT \ram_reg[0][4]  ( .CLK(n351), .D(N20), .Q(\ram[0][4] ) );
  LATCHX1_HVT \ram_reg[0][3]  ( .CLK(n350), .D(N19), .Q(\ram[0][3] ) );
  LATCHX1_HVT \ram_reg[0][2]  ( .CLK(n351), .D(N18), .Q(\ram[0][2] ) );
  LATCHX1_HVT \ram_reg[0][1]  ( .CLK(n352), .D(N17), .Q(\ram[0][1] ) );
  LATCHX1_HVT \ram_reg[0][0]  ( .CLK(n356), .D(N16), .Q(\ram[0][0] ) );
  INVX1_HVT U3 ( .A(n550), .Y(n547) );
  INVX1_HVT U4 ( .A(n604), .Y(n580) );
  INVX1_HVT U5 ( .A(n602), .Y(n581) );
  INVX1_HVT U6 ( .A(n603), .Y(n582) );
  INVX1_HVT U7 ( .A(n604), .Y(n583) );
  INVX1_HVT U8 ( .A(n550), .Y(n462) );
  INVX1_HVT U9 ( .A(n549), .Y(n463) );
  INVX1_HVT U10 ( .A(n604), .Y(n584) );
  INVX1_HVT U11 ( .A(n604), .Y(n585) );
  INVX1_HVT U12 ( .A(n604), .Y(n586) );
  INVX1_HVT U13 ( .A(n604), .Y(n587) );
  INVX1_HVT U14 ( .A(n604), .Y(n588) );
  INVX1_HVT U15 ( .A(n604), .Y(n589) );
  INVX1_HVT U16 ( .A(n603), .Y(n591) );
  INVX1_HVT U17 ( .A(n603), .Y(n592) );
  INVX1_HVT U18 ( .A(n603), .Y(n593) );
  INVX1_HVT U19 ( .A(n603), .Y(n594) );
  INVX1_HVT U20 ( .A(n603), .Y(n595) );
  INVX1_HVT U21 ( .A(n602), .Y(n596) );
  INVX1_HVT U22 ( .A(n602), .Y(n597) );
  INVX1_HVT U23 ( .A(n602), .Y(n598) );
  INVX1_HVT U24 ( .A(n602), .Y(n599) );
  INVX1_HVT U25 ( .A(n602), .Y(n600) );
  INVX1_HVT U26 ( .A(n603), .Y(n590) );
  INVX1_HVT U27 ( .A(n461), .Y(n446) );
  INVX1_HVT U28 ( .A(n461), .Y(n447) );
  INVX1_HVT U29 ( .A(n461), .Y(n448) );
  INVX1_HVT U30 ( .A(n461), .Y(n449) );
  INVX1_HVT U31 ( .A(n461), .Y(n450) );
  INVX1_HVT U32 ( .A(n461), .Y(n451) );
  INVX1_HVT U33 ( .A(n461), .Y(n452) );
  INVX1_HVT U34 ( .A(n461), .Y(n453) );
  INVX1_HVT U35 ( .A(n579), .Y(n567) );
  INVX1_HVT U36 ( .A(n579), .Y(n568) );
  INVX1_HVT U37 ( .A(n579), .Y(n569) );
  INVX1_HVT U38 ( .A(n579), .Y(n570) );
  INVX1_HVT U39 ( .A(n579), .Y(n571) );
  INVX1_HVT U40 ( .A(n579), .Y(n572) );
  INVX1_HVT U41 ( .A(n579), .Y(n573) );
  INVX1_HVT U42 ( .A(n579), .Y(n574) );
  INVX1_HVT U43 ( .A(n579), .Y(n575) );
  INVX1_HVT U44 ( .A(n579), .Y(n576) );
  INVX1_HVT U45 ( .A(n579), .Y(n577) );
  INVX1_HVT U46 ( .A(n455), .Y(n369) );
  INVX1_HVT U47 ( .A(n455), .Y(n370) );
  INVX1_HVT U48 ( .A(n455), .Y(n371) );
  INVX1_HVT U49 ( .A(n455), .Y(n372) );
  INVX1_HVT U50 ( .A(n455), .Y(n373) );
  INVX1_HVT U51 ( .A(n455), .Y(n374) );
  INVX1_HVT U52 ( .A(n455), .Y(n375) );
  INVX1_HVT U53 ( .A(n455), .Y(n376) );
  INVX1_HVT U54 ( .A(n455), .Y(n377) );
  INVX1_HVT U55 ( .A(n455), .Y(n378) );
  INVX1_HVT U56 ( .A(n455), .Y(n379) );
  INVX1_HVT U57 ( .A(n455), .Y(n380) );
  INVX1_HVT U58 ( .A(n458), .Y(n412) );
  INVX1_HVT U59 ( .A(n458), .Y(n413) );
  INVX1_HVT U60 ( .A(n458), .Y(n414) );
  INVX1_HVT U61 ( .A(n458), .Y(n415) );
  INVX1_HVT U62 ( .A(n458), .Y(n416) );
  INVX1_HVT U63 ( .A(n458), .Y(n417) );
  INVX1_HVT U64 ( .A(n458), .Y(n418) );
  INVX1_HVT U65 ( .A(n458), .Y(n419) );
  INVX1_HVT U66 ( .A(n459), .Y(n420) );
  INVX1_HVT U67 ( .A(n459), .Y(n421) );
  INVX1_HVT U68 ( .A(n459), .Y(n422) );
  INVX1_HVT U69 ( .A(n459), .Y(n423) );
  INVX1_HVT U70 ( .A(n459), .Y(n424) );
  INVX1_HVT U71 ( .A(n459), .Y(n425) );
  INVX1_HVT U72 ( .A(n459), .Y(n426) );
  INVX1_HVT U73 ( .A(n459), .Y(n427) );
  INVX1_HVT U74 ( .A(n459), .Y(n428) );
  INVX1_HVT U75 ( .A(n459), .Y(n429) );
  INVX1_HVT U76 ( .A(n459), .Y(n430) );
  INVX1_HVT U77 ( .A(n459), .Y(n431) );
  INVX1_HVT U78 ( .A(n459), .Y(n432) );
  INVX1_HVT U79 ( .A(n460), .Y(n433) );
  INVX1_HVT U80 ( .A(n460), .Y(n434) );
  INVX1_HVT U81 ( .A(n460), .Y(n435) );
  INVX1_HVT U82 ( .A(n460), .Y(n436) );
  INVX1_HVT U83 ( .A(n460), .Y(n437) );
  INVX1_HVT U84 ( .A(n460), .Y(n438) );
  INVX1_HVT U85 ( .A(n460), .Y(n439) );
  INVX1_HVT U86 ( .A(n460), .Y(n440) );
  INVX1_HVT U87 ( .A(n460), .Y(n441) );
  INVX1_HVT U88 ( .A(n460), .Y(n442) );
  INVX1_HVT U89 ( .A(n460), .Y(n443) );
  INVX1_HVT U90 ( .A(n460), .Y(n444) );
  INVX1_HVT U91 ( .A(n460), .Y(n445) );
  INVX1_HVT U92 ( .A(n456), .Y(n381) );
  INVX1_HVT U93 ( .A(n456), .Y(n382) );
  INVX1_HVT U94 ( .A(n456), .Y(n383) );
  INVX1_HVT U95 ( .A(n456), .Y(n384) );
  INVX1_HVT U96 ( .A(n456), .Y(n385) );
  INVX1_HVT U97 ( .A(n456), .Y(n386) );
  INVX1_HVT U98 ( .A(n456), .Y(n387) );
  INVX1_HVT U99 ( .A(n456), .Y(n388) );
  INVX1_HVT U100 ( .A(n456), .Y(n389) );
  INVX1_HVT U101 ( .A(n456), .Y(n390) );
  INVX1_HVT U102 ( .A(n456), .Y(n391) );
  INVX1_HVT U103 ( .A(n456), .Y(n392) );
  INVX1_HVT U104 ( .A(n456), .Y(n393) );
  INVX1_HVT U105 ( .A(n457), .Y(n394) );
  INVX1_HVT U106 ( .A(n457), .Y(n395) );
  INVX1_HVT U107 ( .A(n457), .Y(n396) );
  INVX1_HVT U108 ( .A(n457), .Y(n397) );
  INVX1_HVT U109 ( .A(n457), .Y(n398) );
  INVX1_HVT U110 ( .A(n457), .Y(n399) );
  INVX1_HVT U111 ( .A(n457), .Y(n400) );
  INVX1_HVT U112 ( .A(n457), .Y(n401) );
  INVX1_HVT U113 ( .A(n457), .Y(n402) );
  INVX1_HVT U114 ( .A(n457), .Y(n403) );
  INVX1_HVT U115 ( .A(n457), .Y(n404) );
  INVX1_HVT U116 ( .A(n457), .Y(n405) );
  INVX1_HVT U117 ( .A(n457), .Y(n406) );
  INVX1_HVT U118 ( .A(n458), .Y(n407) );
  INVX1_HVT U119 ( .A(n458), .Y(n408) );
  INVX1_HVT U120 ( .A(n458), .Y(n409) );
  INVX1_HVT U121 ( .A(n458), .Y(n410) );
  INVX1_HVT U122 ( .A(n458), .Y(n411) );
  INVX1_HVT U123 ( .A(n578), .Y(n558) );
  INVX1_HVT U124 ( .A(n578), .Y(n559) );
  INVX1_HVT U125 ( .A(n578), .Y(n560) );
  INVX1_HVT U126 ( .A(n578), .Y(n561) );
  INVX1_HVT U127 ( .A(n578), .Y(n562) );
  INVX1_HVT U128 ( .A(n578), .Y(n563) );
  INVX1_HVT U129 ( .A(n578), .Y(n564) );
  INVX1_HVT U130 ( .A(n578), .Y(n565) );
  INVX1_HVT U131 ( .A(n578), .Y(n566) );
  INVX1_HVT U132 ( .A(n578), .Y(n557) );
  INVX1_HVT U133 ( .A(n553), .Y(n536) );
  INVX1_HVT U134 ( .A(n550), .Y(n537) );
  INVX1_HVT U135 ( .A(n549), .Y(n538) );
  INVX1_HVT U136 ( .A(n548), .Y(n539) );
  INVX1_HVT U137 ( .A(n556), .Y(n540) );
  INVX1_HVT U138 ( .A(n555), .Y(n541) );
  INVX1_HVT U139 ( .A(n549), .Y(n542) );
  INVX1_HVT U140 ( .A(n548), .Y(n543) );
  INVX1_HVT U141 ( .A(n556), .Y(n544) );
  INVX1_HVT U142 ( .A(n555), .Y(n545) );
  INVX1_HVT U143 ( .A(n554), .Y(n546) );
  INVX1_HVT U144 ( .A(n461), .Y(n454) );
  INVX1_HVT U145 ( .A(n552), .Y(n505) );
  INVX1_HVT U146 ( .A(n550), .Y(n506) );
  INVX1_HVT U147 ( .A(n550), .Y(n507) );
  INVX1_HVT U148 ( .A(n550), .Y(n508) );
  INVX1_HVT U149 ( .A(n550), .Y(n509) );
  INVX1_HVT U150 ( .A(n550), .Y(n510) );
  INVX1_HVT U151 ( .A(n550), .Y(n511) );
  INVX1_HVT U152 ( .A(n549), .Y(n512) );
  INVX1_HVT U153 ( .A(n549), .Y(n513) );
  INVX1_HVT U154 ( .A(n549), .Y(n514) );
  INVX1_HVT U155 ( .A(n549), .Y(n515) );
  INVX1_HVT U156 ( .A(n549), .Y(n516) );
  INVX1_HVT U157 ( .A(n549), .Y(n517) );
  INVX1_HVT U158 ( .A(n548), .Y(n518) );
  INVX1_HVT U159 ( .A(n548), .Y(n519) );
  INVX1_HVT U160 ( .A(n548), .Y(n520) );
  INVX1_HVT U161 ( .A(n548), .Y(n521) );
  INVX1_HVT U162 ( .A(n548), .Y(n522) );
  INVX1_HVT U163 ( .A(n548), .Y(n523) );
  INVX1_HVT U164 ( .A(n556), .Y(n524) );
  INVX1_HVT U165 ( .A(n555), .Y(n525) );
  INVX1_HVT U166 ( .A(n554), .Y(n526) );
  INVX1_HVT U167 ( .A(n553), .Y(n527) );
  INVX1_HVT U168 ( .A(n552), .Y(n528) );
  INVX1_HVT U169 ( .A(n551), .Y(n529) );
  INVX1_HVT U170 ( .A(n548), .Y(n530) );
  INVX1_HVT U171 ( .A(n548), .Y(n531) );
  INVX1_HVT U172 ( .A(n556), .Y(n532) );
  INVX1_HVT U173 ( .A(n555), .Y(n533) );
  INVX1_HVT U174 ( .A(n554), .Y(n534) );
  INVX1_HVT U175 ( .A(n553), .Y(n535) );
  INVX1_HVT U176 ( .A(n556), .Y(n464) );
  INVX1_HVT U177 ( .A(n556), .Y(n465) );
  INVX1_HVT U178 ( .A(n556), .Y(n466) );
  INVX1_HVT U179 ( .A(n556), .Y(n467) );
  INVX1_HVT U180 ( .A(n556), .Y(n468) );
  INVX1_HVT U181 ( .A(n556), .Y(n469) );
  INVX1_HVT U182 ( .A(n555), .Y(n470) );
  INVX1_HVT U183 ( .A(n555), .Y(n471) );
  INVX1_HVT U184 ( .A(n555), .Y(n472) );
  INVX1_HVT U185 ( .A(n555), .Y(n473) );
  INVX1_HVT U186 ( .A(n555), .Y(n474) );
  INVX1_HVT U187 ( .A(n555), .Y(n475) );
  INVX1_HVT U188 ( .A(n554), .Y(n476) );
  INVX1_HVT U189 ( .A(n554), .Y(n477) );
  INVX1_HVT U190 ( .A(n554), .Y(n478) );
  INVX1_HVT U191 ( .A(n554), .Y(n479) );
  INVX1_HVT U192 ( .A(n554), .Y(n480) );
  INVX1_HVT U193 ( .A(n554), .Y(n481) );
  INVX1_HVT U194 ( .A(n553), .Y(n482) );
  INVX1_HVT U195 ( .A(n553), .Y(n483) );
  INVX1_HVT U196 ( .A(n553), .Y(n484) );
  INVX1_HVT U197 ( .A(n553), .Y(n485) );
  INVX1_HVT U198 ( .A(n553), .Y(n486) );
  INVX1_HVT U199 ( .A(n553), .Y(n487) );
  INVX1_HVT U200 ( .A(n552), .Y(n488) );
  INVX1_HVT U201 ( .A(n552), .Y(n489) );
  INVX1_HVT U202 ( .A(n552), .Y(n490) );
  INVX1_HVT U203 ( .A(n552), .Y(n491) );
  INVX1_HVT U204 ( .A(n552), .Y(n492) );
  INVX1_HVT U205 ( .A(n552), .Y(n493) );
  INVX1_HVT U206 ( .A(n551), .Y(n494) );
  INVX1_HVT U207 ( .A(n551), .Y(n495) );
  INVX1_HVT U208 ( .A(n551), .Y(n496) );
  INVX1_HVT U209 ( .A(n551), .Y(n497) );
  INVX1_HVT U210 ( .A(n551), .Y(n498) );
  INVX1_HVT U211 ( .A(n551), .Y(n499) );
  INVX1_HVT U212 ( .A(n551), .Y(n500) );
  INVX1_HVT U213 ( .A(n551), .Y(n501) );
  INVX1_HVT U214 ( .A(n552), .Y(n502) );
  INVX1_HVT U215 ( .A(n550), .Y(n503) );
  INVX1_HVT U216 ( .A(n549), .Y(n504) );
  INVX1_HVT U217 ( .A(n368), .Y(n348) );
  INVX1_HVT U218 ( .A(n367), .Y(n351) );
  INVX1_HVT U219 ( .A(n367), .Y(n352) );
  INVX1_HVT U220 ( .A(n367), .Y(n350) );
  INVX1_HVT U221 ( .A(n367), .Y(n353) );
  INVX1_HVT U222 ( .A(n368), .Y(n349) );
  INVX1_HVT U223 ( .A(n367), .Y(n354) );
  INVX1_HVT U224 ( .A(n367), .Y(n355) );
  INVX1_HVT U225 ( .A(n368), .Y(n346) );
  INVX1_HVT U226 ( .A(n368), .Y(n347) );
  INVX1_HVT U227 ( .A(n368), .Y(n359) );
  INVX1_HVT U228 ( .A(n368), .Y(n360) );
  INVX1_HVT U229 ( .A(n368), .Y(n361) );
  INVX1_HVT U230 ( .A(n368), .Y(n362) );
  INVX1_HVT U231 ( .A(n367), .Y(n363) );
  INVX1_HVT U232 ( .A(n368), .Y(n364) );
  INVX1_HVT U233 ( .A(n367), .Y(n365) );
  INVX1_HVT U234 ( .A(n367), .Y(n356) );
  INVX1_HVT U235 ( .A(n368), .Y(n357) );
  INVX1_HVT U236 ( .A(n367), .Y(n358) );
  INVX1_HVT U237 ( .A(n368), .Y(n366) );
  INVX1_HVT U238 ( .A(n345), .Y(n325) );
  INVX1_HVT U239 ( .A(n345), .Y(n328) );
  INVX1_HVT U240 ( .A(n345), .Y(n329) );
  INVX1_HVT U241 ( .A(n345), .Y(n327) );
  INVX1_HVT U242 ( .A(n345), .Y(n330) );
  INVX1_HVT U243 ( .A(n345), .Y(n326) );
  INVX1_HVT U244 ( .A(n345), .Y(n331) );
  INVX1_HVT U245 ( .A(n345), .Y(n332) );
  INVX1_HVT U246 ( .A(n345), .Y(n323) );
  INVX1_HVT U247 ( .A(n345), .Y(n324) );
  INVX1_HVT U248 ( .A(n344), .Y(n336) );
  INVX1_HVT U249 ( .A(n344), .Y(n337) );
  INVX1_HVT U250 ( .A(n344), .Y(n338) );
  INVX1_HVT U251 ( .A(n344), .Y(n339) );
  INVX1_HVT U252 ( .A(n344), .Y(n340) );
  INVX1_HVT U253 ( .A(n344), .Y(n341) );
  INVX1_HVT U254 ( .A(n344), .Y(n342) );
  INVX1_HVT U255 ( .A(n344), .Y(n333) );
  INVX1_HVT U256 ( .A(n344), .Y(n334) );
  INVX1_HVT U257 ( .A(n344), .Y(n335) );
  INVX1_HVT U258 ( .A(n344), .Y(n343) );
  INVX1_HVT U259 ( .A(n322), .Y(n302) );
  INVX1_HVT U260 ( .A(n321), .Y(n305) );
  INVX1_HVT U261 ( .A(n321), .Y(n306) );
  INVX1_HVT U262 ( .A(n321), .Y(n304) );
  INVX1_HVT U263 ( .A(n321), .Y(n307) );
  INVX1_HVT U264 ( .A(n322), .Y(n303) );
  INVX1_HVT U265 ( .A(n321), .Y(n308) );
  INVX1_HVT U266 ( .A(n321), .Y(n309) );
  INVX1_HVT U267 ( .A(n322), .Y(n300) );
  INVX1_HVT U268 ( .A(n322), .Y(n301) );
  INVX1_HVT U269 ( .A(n322), .Y(n313) );
  INVX1_HVT U270 ( .A(n322), .Y(n314) );
  INVX1_HVT U271 ( .A(n322), .Y(n315) );
  INVX1_HVT U272 ( .A(n322), .Y(n316) );
  INVX1_HVT U273 ( .A(n321), .Y(n317) );
  INVX1_HVT U274 ( .A(n322), .Y(n318) );
  INVX1_HVT U275 ( .A(n321), .Y(n319) );
  INVX1_HVT U276 ( .A(n321), .Y(n310) );
  INVX1_HVT U277 ( .A(n322), .Y(n311) );
  INVX1_HVT U278 ( .A(n321), .Y(n312) );
  INVX1_HVT U279 ( .A(n322), .Y(n320) );
  INVX1_HVT U280 ( .A(n299), .Y(n279) );
  INVX1_HVT U281 ( .A(n299), .Y(n282) );
  INVX1_HVT U282 ( .A(n299), .Y(n283) );
  INVX1_HVT U283 ( .A(n299), .Y(n281) );
  INVX1_HVT U284 ( .A(n299), .Y(n284) );
  INVX1_HVT U285 ( .A(n299), .Y(n280) );
  INVX1_HVT U286 ( .A(n299), .Y(n285) );
  INVX1_HVT U287 ( .A(n299), .Y(n286) );
  INVX1_HVT U288 ( .A(n299), .Y(n277) );
  INVX1_HVT U289 ( .A(n299), .Y(n278) );
  INVX1_HVT U290 ( .A(n298), .Y(n290) );
  INVX1_HVT U291 ( .A(n298), .Y(n291) );
  INVX1_HVT U292 ( .A(n298), .Y(n292) );
  INVX1_HVT U293 ( .A(n298), .Y(n293) );
  INVX1_HVT U294 ( .A(n298), .Y(n294) );
  INVX1_HVT U295 ( .A(n298), .Y(n295) );
  INVX1_HVT U296 ( .A(n298), .Y(n296) );
  INVX1_HVT U297 ( .A(n298), .Y(n287) );
  INVX1_HVT U298 ( .A(n298), .Y(n288) );
  INVX1_HVT U299 ( .A(n298), .Y(n289) );
  INVX1_HVT U300 ( .A(n298), .Y(n297) );
  INVX1_HVT U301 ( .A(n276), .Y(n256) );
  INVX1_HVT U302 ( .A(n275), .Y(n259) );
  INVX1_HVT U303 ( .A(n275), .Y(n260) );
  INVX1_HVT U304 ( .A(n275), .Y(n258) );
  INVX1_HVT U305 ( .A(n275), .Y(n261) );
  INVX1_HVT U306 ( .A(n276), .Y(n257) );
  INVX1_HVT U307 ( .A(n275), .Y(n262) );
  INVX1_HVT U308 ( .A(n275), .Y(n263) );
  INVX1_HVT U309 ( .A(n276), .Y(n254) );
  INVX1_HVT U310 ( .A(n276), .Y(n255) );
  INVX1_HVT U311 ( .A(n276), .Y(n267) );
  INVX1_HVT U312 ( .A(n276), .Y(n268) );
  INVX1_HVT U313 ( .A(n276), .Y(n269) );
  INVX1_HVT U314 ( .A(n276), .Y(n270) );
  INVX1_HVT U315 ( .A(n275), .Y(n271) );
  INVX1_HVT U316 ( .A(n276), .Y(n272) );
  INVX1_HVT U317 ( .A(n275), .Y(n273) );
  INVX1_HVT U318 ( .A(n275), .Y(n264) );
  INVX1_HVT U319 ( .A(n276), .Y(n265) );
  INVX1_HVT U320 ( .A(n275), .Y(n266) );
  INVX1_HVT U321 ( .A(n276), .Y(n274) );
  INVX1_HVT U322 ( .A(n253), .Y(n233) );
  INVX1_HVT U323 ( .A(n253), .Y(n236) );
  INVX1_HVT U324 ( .A(n253), .Y(n237) );
  INVX1_HVT U325 ( .A(n253), .Y(n235) );
  INVX1_HVT U326 ( .A(n253), .Y(n238) );
  INVX1_HVT U327 ( .A(n253), .Y(n234) );
  INVX1_HVT U328 ( .A(n253), .Y(n239) );
  INVX1_HVT U329 ( .A(n253), .Y(n240) );
  INVX1_HVT U330 ( .A(n253), .Y(n231) );
  INVX1_HVT U331 ( .A(n253), .Y(n232) );
  INVX1_HVT U332 ( .A(n252), .Y(n244) );
  INVX1_HVT U333 ( .A(n252), .Y(n245) );
  INVX1_HVT U334 ( .A(n252), .Y(n246) );
  INVX1_HVT U335 ( .A(n252), .Y(n247) );
  INVX1_HVT U336 ( .A(n252), .Y(n248) );
  INVX1_HVT U337 ( .A(n252), .Y(n249) );
  INVX1_HVT U338 ( .A(n252), .Y(n250) );
  INVX1_HVT U339 ( .A(n252), .Y(n241) );
  INVX1_HVT U340 ( .A(n252), .Y(n242) );
  INVX1_HVT U341 ( .A(n252), .Y(n243) );
  INVX1_HVT U342 ( .A(n252), .Y(n251) );
  INVX1_HVT U343 ( .A(n230), .Y(n210) );
  INVX1_HVT U344 ( .A(n229), .Y(n213) );
  INVX1_HVT U345 ( .A(n229), .Y(n214) );
  INVX1_HVT U346 ( .A(n229), .Y(n212) );
  INVX1_HVT U347 ( .A(n229), .Y(n215) );
  INVX1_HVT U348 ( .A(n230), .Y(n211) );
  INVX1_HVT U349 ( .A(n229), .Y(n216) );
  INVX1_HVT U350 ( .A(n229), .Y(n217) );
  INVX1_HVT U351 ( .A(n230), .Y(n208) );
  INVX1_HVT U352 ( .A(n230), .Y(n209) );
  INVX1_HVT U353 ( .A(n230), .Y(n221) );
  INVX1_HVT U354 ( .A(n230), .Y(n222) );
  INVX1_HVT U355 ( .A(n230), .Y(n223) );
  INVX1_HVT U356 ( .A(n230), .Y(n224) );
  INVX1_HVT U357 ( .A(n229), .Y(n225) );
  INVX1_HVT U358 ( .A(n230), .Y(n226) );
  INVX1_HVT U359 ( .A(n229), .Y(n227) );
  INVX1_HVT U360 ( .A(n229), .Y(n218) );
  INVX1_HVT U361 ( .A(n230), .Y(n219) );
  INVX1_HVT U362 ( .A(n229), .Y(n220) );
  INVX1_HVT U363 ( .A(n230), .Y(n228) );
  INVX1_HVT U364 ( .A(n207), .Y(n187) );
  INVX1_HVT U365 ( .A(n207), .Y(n190) );
  INVX1_HVT U366 ( .A(n207), .Y(n191) );
  INVX1_HVT U367 ( .A(n207), .Y(n189) );
  INVX1_HVT U368 ( .A(n207), .Y(n192) );
  INVX1_HVT U369 ( .A(n207), .Y(n188) );
  INVX1_HVT U370 ( .A(n207), .Y(n193) );
  INVX1_HVT U371 ( .A(n207), .Y(n194) );
  INVX1_HVT U372 ( .A(n207), .Y(n186) );
  INVX1_HVT U373 ( .A(n206), .Y(n195) );
  INVX1_HVT U374 ( .A(n206), .Y(n199) );
  INVX1_HVT U375 ( .A(n206), .Y(n200) );
  INVX1_HVT U376 ( .A(n206), .Y(n201) );
  INVX1_HVT U377 ( .A(n206), .Y(n202) );
  INVX1_HVT U378 ( .A(n206), .Y(n203) );
  INVX1_HVT U379 ( .A(n206), .Y(n204) );
  INVX1_HVT U380 ( .A(n206), .Y(n205) );
  INVX1_HVT U381 ( .A(n206), .Y(n196) );
  INVX1_HVT U382 ( .A(n206), .Y(n197) );
  INVX1_HVT U383 ( .A(n206), .Y(n198) );
  INVX1_HVT U384 ( .A(n207), .Y(n185) );
  INVX1_HVT U385 ( .A(n184), .Y(n164) );
  INVX1_HVT U386 ( .A(n183), .Y(n167) );
  INVX1_HVT U387 ( .A(n183), .Y(n168) );
  INVX1_HVT U388 ( .A(n183), .Y(n166) );
  INVX1_HVT U389 ( .A(n183), .Y(n169) );
  INVX1_HVT U390 ( .A(n184), .Y(n165) );
  INVX1_HVT U391 ( .A(n183), .Y(n170) );
  INVX1_HVT U392 ( .A(n183), .Y(n171) );
  INVX1_HVT U393 ( .A(n184), .Y(n162) );
  INVX1_HVT U394 ( .A(n184), .Y(n163) );
  INVX1_HVT U395 ( .A(n184), .Y(n175) );
  INVX1_HVT U396 ( .A(n184), .Y(n176) );
  INVX1_HVT U397 ( .A(n184), .Y(n177) );
  INVX1_HVT U398 ( .A(n184), .Y(n178) );
  INVX1_HVT U399 ( .A(n183), .Y(n179) );
  INVX1_HVT U400 ( .A(n184), .Y(n180) );
  INVX1_HVT U401 ( .A(n183), .Y(n181) );
  INVX1_HVT U402 ( .A(n183), .Y(n172) );
  INVX1_HVT U403 ( .A(n184), .Y(n173) );
  INVX1_HVT U404 ( .A(n183), .Y(n174) );
  INVX1_HVT U405 ( .A(n184), .Y(n182) );
  INVX1_HVT U406 ( .A(n161), .Y(n141) );
  INVX1_HVT U407 ( .A(n161), .Y(n144) );
  INVX1_HVT U408 ( .A(n161), .Y(n145) );
  INVX1_HVT U409 ( .A(n161), .Y(n143) );
  INVX1_HVT U410 ( .A(n161), .Y(n146) );
  INVX1_HVT U411 ( .A(n161), .Y(n142) );
  INVX1_HVT U412 ( .A(n161), .Y(n147) );
  INVX1_HVT U413 ( .A(n161), .Y(n148) );
  INVX1_HVT U414 ( .A(n161), .Y(n139) );
  INVX1_HVT U415 ( .A(n161), .Y(n140) );
  INVX1_HVT U416 ( .A(n160), .Y(n152) );
  INVX1_HVT U417 ( .A(n160), .Y(n153) );
  INVX1_HVT U418 ( .A(n160), .Y(n154) );
  INVX1_HVT U419 ( .A(n160), .Y(n155) );
  INVX1_HVT U420 ( .A(n160), .Y(n156) );
  INVX1_HVT U421 ( .A(n160), .Y(n157) );
  INVX1_HVT U422 ( .A(n160), .Y(n158) );
  INVX1_HVT U423 ( .A(n160), .Y(n149) );
  INVX1_HVT U424 ( .A(n160), .Y(n150) );
  INVX1_HVT U425 ( .A(n160), .Y(n151) );
  INVX1_HVT U426 ( .A(n160), .Y(n159) );
  INVX1_HVT U427 ( .A(n138), .Y(n118) );
  INVX1_HVT U428 ( .A(n137), .Y(n121) );
  INVX1_HVT U429 ( .A(n137), .Y(n122) );
  INVX1_HVT U430 ( .A(n137), .Y(n120) );
  INVX1_HVT U431 ( .A(n137), .Y(n123) );
  INVX1_HVT U432 ( .A(n138), .Y(n119) );
  INVX1_HVT U433 ( .A(n137), .Y(n124) );
  INVX1_HVT U434 ( .A(n137), .Y(n125) );
  INVX1_HVT U435 ( .A(n138), .Y(n116) );
  INVX1_HVT U436 ( .A(n138), .Y(n117) );
  INVX1_HVT U437 ( .A(n138), .Y(n129) );
  INVX1_HVT U438 ( .A(n138), .Y(n130) );
  INVX1_HVT U439 ( .A(n138), .Y(n131) );
  INVX1_HVT U440 ( .A(n138), .Y(n132) );
  INVX1_HVT U441 ( .A(n137), .Y(n133) );
  INVX1_HVT U442 ( .A(n138), .Y(n134) );
  INVX1_HVT U443 ( .A(n137), .Y(n135) );
  INVX1_HVT U444 ( .A(n137), .Y(n126) );
  INVX1_HVT U445 ( .A(n138), .Y(n127) );
  INVX1_HVT U446 ( .A(n137), .Y(n128) );
  INVX1_HVT U447 ( .A(n138), .Y(n136) );
  INVX1_HVT U448 ( .A(n115), .Y(n95) );
  INVX1_HVT U449 ( .A(n115), .Y(n98) );
  INVX1_HVT U450 ( .A(n115), .Y(n99) );
  INVX1_HVT U451 ( .A(n115), .Y(n97) );
  INVX1_HVT U452 ( .A(n115), .Y(n100) );
  INVX1_HVT U453 ( .A(n115), .Y(n96) );
  INVX1_HVT U454 ( .A(n115), .Y(n101) );
  INVX1_HVT U455 ( .A(n115), .Y(n102) );
  INVX1_HVT U456 ( .A(n115), .Y(n94) );
  INVX1_HVT U457 ( .A(n114), .Y(n106) );
  INVX1_HVT U458 ( .A(n114), .Y(n107) );
  INVX1_HVT U459 ( .A(n114), .Y(n108) );
  INVX1_HVT U460 ( .A(n114), .Y(n109) );
  INVX1_HVT U461 ( .A(n114), .Y(n110) );
  INVX1_HVT U462 ( .A(n114), .Y(n111) );
  INVX1_HVT U463 ( .A(n114), .Y(n112) );
  INVX1_HVT U464 ( .A(n114), .Y(n113) );
  INVX1_HVT U465 ( .A(n114), .Y(n103) );
  INVX1_HVT U466 ( .A(n114), .Y(n104) );
  INVX1_HVT U467 ( .A(n114), .Y(n105) );
  INVX1_HVT U468 ( .A(n115), .Y(n93) );
  INVX1_HVT U469 ( .A(n92), .Y(n72) );
  INVX1_HVT U470 ( .A(n91), .Y(n75) );
  INVX1_HVT U471 ( .A(n91), .Y(n76) );
  INVX1_HVT U472 ( .A(n91), .Y(n74) );
  INVX1_HVT U473 ( .A(n91), .Y(n77) );
  INVX1_HVT U474 ( .A(n92), .Y(n73) );
  INVX1_HVT U475 ( .A(n91), .Y(n78) );
  INVX1_HVT U476 ( .A(n91), .Y(n79) );
  INVX1_HVT U477 ( .A(n92), .Y(n70) );
  INVX1_HVT U478 ( .A(n92), .Y(n71) );
  INVX1_HVT U479 ( .A(n92), .Y(n83) );
  INVX1_HVT U480 ( .A(n92), .Y(n84) );
  INVX1_HVT U481 ( .A(n92), .Y(n85) );
  INVX1_HVT U482 ( .A(n92), .Y(n86) );
  INVX1_HVT U483 ( .A(n91), .Y(n87) );
  INVX1_HVT U484 ( .A(n92), .Y(n88) );
  INVX1_HVT U485 ( .A(n91), .Y(n89) );
  INVX1_HVT U486 ( .A(n91), .Y(n80) );
  INVX1_HVT U487 ( .A(n92), .Y(n81) );
  INVX1_HVT U488 ( .A(n91), .Y(n82) );
  INVX1_HVT U489 ( .A(n92), .Y(n90) );
  INVX1_HVT U490 ( .A(n69), .Y(n49) );
  INVX1_HVT U491 ( .A(n69), .Y(n52) );
  INVX1_HVT U492 ( .A(n69), .Y(n53) );
  INVX1_HVT U493 ( .A(n69), .Y(n51) );
  INVX1_HVT U494 ( .A(n69), .Y(n54) );
  INVX1_HVT U495 ( .A(n69), .Y(n50) );
  INVX1_HVT U496 ( .A(n69), .Y(n55) );
  INVX1_HVT U497 ( .A(n69), .Y(n56) );
  INVX1_HVT U498 ( .A(n69), .Y(n48) );
  INVX1_HVT U499 ( .A(n68), .Y(n60) );
  INVX1_HVT U500 ( .A(n68), .Y(n61) );
  INVX1_HVT U501 ( .A(n68), .Y(n62) );
  INVX1_HVT U502 ( .A(n68), .Y(n63) );
  INVX1_HVT U503 ( .A(n68), .Y(n64) );
  INVX1_HVT U504 ( .A(n68), .Y(n65) );
  INVX1_HVT U505 ( .A(n68), .Y(n66) );
  INVX1_HVT U506 ( .A(n68), .Y(n67) );
  INVX1_HVT U507 ( .A(n68), .Y(n57) );
  INVX1_HVT U508 ( .A(n68), .Y(n58) );
  INVX1_HVT U509 ( .A(n68), .Y(n59) );
  INVX1_HVT U510 ( .A(n69), .Y(n47) );
  INVX1_HVT U511 ( .A(n46), .Y(n27) );
  INVX1_HVT U512 ( .A(n45), .Y(n29) );
  INVX1_HVT U513 ( .A(n45), .Y(n30) );
  INVX1_HVT U514 ( .A(n45), .Y(n31) );
  INVX1_HVT U515 ( .A(n45), .Y(n28) );
  INVX1_HVT U516 ( .A(n45), .Y(n32) );
  INVX1_HVT U517 ( .A(n45), .Y(n33) );
  INVX1_HVT U518 ( .A(n46), .Y(n34) );
  INVX1_HVT U519 ( .A(n46), .Y(n25) );
  INVX1_HVT U520 ( .A(n46), .Y(n26) );
  INVX1_HVT U521 ( .A(n46), .Y(n38) );
  INVX1_HVT U522 ( .A(n46), .Y(n39) );
  INVX1_HVT U523 ( .A(n46), .Y(n40) );
  INVX1_HVT U524 ( .A(n45), .Y(n41) );
  INVX1_HVT U525 ( .A(n46), .Y(n42) );
  INVX1_HVT U526 ( .A(n45), .Y(n43) );
  INVX1_HVT U527 ( .A(n46), .Y(n44) );
  INVX1_HVT U528 ( .A(n45), .Y(n35) );
  INVX1_HVT U529 ( .A(n46), .Y(n36) );
  INVX1_HVT U530 ( .A(n45), .Y(n37) );
  INVX1_HVT U531 ( .A(n46), .Y(n24) );
  INVX1_HVT U532 ( .A(n23), .Y(n3) );
  INVX1_HVT U533 ( .A(n23), .Y(n6) );
  INVX1_HVT U534 ( .A(n23), .Y(n7) );
  INVX1_HVT U535 ( .A(n23), .Y(n5) );
  INVX1_HVT U536 ( .A(n23), .Y(n8) );
  INVX1_HVT U537 ( .A(n23), .Y(n4) );
  INVX1_HVT U538 ( .A(n23), .Y(n9) );
  INVX1_HVT U539 ( .A(n23), .Y(n10) );
  INVX1_HVT U540 ( .A(n23), .Y(n1) );
  INVX1_HVT U541 ( .A(n23), .Y(n2) );
  INVX1_HVT U542 ( .A(n22), .Y(n14) );
  INVX1_HVT U543 ( .A(n22), .Y(n15) );
  INVX1_HVT U544 ( .A(n22), .Y(n16) );
  INVX1_HVT U545 ( .A(n22), .Y(n17) );
  INVX1_HVT U546 ( .A(n22), .Y(n18) );
  INVX1_HVT U547 ( .A(n22), .Y(n19) );
  INVX1_HVT U548 ( .A(n22), .Y(n20) );
  INVX1_HVT U549 ( .A(n22), .Y(n11) );
  INVX1_HVT U550 ( .A(n22), .Y(n12) );
  INVX1_HVT U551 ( .A(n22), .Y(n13) );
  INVX1_HVT U552 ( .A(n22), .Y(n21) );
  INVX1_HVT U553 ( .A(n602), .Y(n601) );
  INVX1_HVT U554 ( .A(N309), .Y(n92) );
  INVX1_HVT U555 ( .A(N312), .Y(n69) );
  INVX1_HVT U556 ( .A(N315), .Y(n46) );
  INVX1_HVT U557 ( .A(N282), .Y(n299) );
  INVX1_HVT U558 ( .A(N294), .Y(n207) );
  INVX1_HVT U559 ( .A(N306), .Y(n115) );
  INVX1_HVT U560 ( .A(N318), .Y(n23) );
  INVX1_HVT U561 ( .A(N215), .Y(n368) );
  INVX1_HVT U562 ( .A(N276), .Y(n345) );
  INVX1_HVT U563 ( .A(N279), .Y(n322) );
  INVX1_HVT U564 ( .A(N285), .Y(n276) );
  INVX1_HVT U565 ( .A(N288), .Y(n253) );
  INVX1_HVT U566 ( .A(N291), .Y(n230) );
  INVX1_HVT U567 ( .A(N297), .Y(n184) );
  INVX1_HVT U568 ( .A(N300), .Y(n161) );
  INVX1_HVT U569 ( .A(N303), .Y(n138) );
  INVX1_HVT U570 ( .A(N309), .Y(n91) );
  INVX1_HVT U571 ( .A(N312), .Y(n68) );
  INVX1_HVT U572 ( .A(N315), .Y(n45) );
  INVX1_HVT U573 ( .A(N282), .Y(n298) );
  INVX1_HVT U574 ( .A(N294), .Y(n206) );
  INVX1_HVT U575 ( .A(N306), .Y(n114) );
  INVX1_HVT U576 ( .A(N318), .Y(n22) );
  INVX1_HVT U577 ( .A(N215), .Y(n367) );
  INVX1_HVT U578 ( .A(N276), .Y(n344) );
  INVX1_HVT U579 ( .A(N279), .Y(n321) );
  INVX1_HVT U580 ( .A(N285), .Y(n275) );
  INVX1_HVT U581 ( .A(N288), .Y(n252) );
  INVX1_HVT U582 ( .A(N291), .Y(n229) );
  INVX1_HVT U583 ( .A(N297), .Y(n183) );
  INVX1_HVT U584 ( .A(N300), .Y(n160) );
  INVX1_HVT U585 ( .A(N303), .Y(n137) );
  INVX1_HVT U586 ( .A(N11), .Y(n579) );
  INVX1_HVT U587 ( .A(N11), .Y(n578) );
  INVX1_HVT U588 ( .A(N12), .Y(n604) );
  INVX1_HVT U589 ( .A(N12), .Y(n602) );
  INVX1_HVT U590 ( .A(N12), .Y(n603) );
  INVX1_HVT U591 ( .A(N9), .Y(n458) );
  INVX1_HVT U592 ( .A(N9), .Y(n459) );
  INVX1_HVT U593 ( .A(N9), .Y(n460) );
  INVX1_HVT U594 ( .A(N9), .Y(n456) );
  INVX1_HVT U595 ( .A(N9), .Y(n457) );
  INVX1_HVT U596 ( .A(N9), .Y(n455) );
  INVX1_HVT U597 ( .A(N9), .Y(n461) );
  INVX1_HVT U598 ( .A(N10), .Y(n550) );
  INVX1_HVT U599 ( .A(N10), .Y(n549) );
  INVX1_HVT U600 ( .A(N10), .Y(n548) );
  INVX1_HVT U601 ( .A(N10), .Y(n556) );
  INVX1_HVT U602 ( .A(N10), .Y(n555) );
  INVX1_HVT U603 ( .A(N10), .Y(n554) );
  INVX1_HVT U604 ( .A(N10), .Y(n553) );
  INVX1_HVT U605 ( .A(N10), .Y(n552) );
  INVX1_HVT U606 ( .A(N10), .Y(n551) );
  MUX41X1_HVT U607 ( .A1(\ram[12][0] ), .A3(\ram[14][0] ), .A2(\ram[13][0] ), 
        .A4(\ram[15][0] ), .S0(n462), .S1(n369), .Y(n605) );
  MUX41X1_HVT U608 ( .A1(\ram[8][0] ), .A3(\ram[10][0] ), .A2(\ram[9][0] ), 
        .A4(\ram[11][0] ), .S0(n462), .S1(n369), .Y(n606) );
  MUX41X1_HVT U609 ( .A1(\ram[4][0] ), .A3(\ram[6][0] ), .A2(\ram[5][0] ), 
        .A4(\ram[7][0] ), .S0(n462), .S1(n369), .Y(n607) );
  MUX41X1_HVT U610 ( .A1(\ram[0][0] ), .A3(\ram[2][0] ), .A2(\ram[1][0] ), 
        .A4(\ram[3][0] ), .S0(n462), .S1(n369), .Y(n608) );
  MUX41X1_HVT U611 ( .A1(n608), .A3(n606), .A2(n607), .A4(n605), .S0(n580), 
        .S1(n557), .Y(q[0]) );
  MUX41X1_HVT U612 ( .A1(\ram[12][1] ), .A3(\ram[14][1] ), .A2(\ram[13][1] ), 
        .A4(\ram[15][1] ), .S0(n462), .S1(n369), .Y(n609) );
  MUX41X1_HVT U613 ( .A1(\ram[8][1] ), .A3(\ram[10][1] ), .A2(\ram[9][1] ), 
        .A4(\ram[11][1] ), .S0(n462), .S1(n369), .Y(n610) );
  MUX41X1_HVT U614 ( .A1(\ram[4][1] ), .A3(\ram[6][1] ), .A2(\ram[5][1] ), 
        .A4(\ram[7][1] ), .S0(n462), .S1(n369), .Y(n611) );
  MUX41X1_HVT U615 ( .A1(\ram[0][1] ), .A3(\ram[2][1] ), .A2(\ram[1][1] ), 
        .A4(\ram[3][1] ), .S0(n462), .S1(n369), .Y(n612) );
  MUX41X1_HVT U616 ( .A1(n612), .A3(n610), .A2(n611), .A4(n609), .S0(n580), 
        .S1(n573), .Y(q[1]) );
  MUX41X1_HVT U617 ( .A1(\ram[12][2] ), .A3(\ram[14][2] ), .A2(\ram[13][2] ), 
        .A4(\ram[15][2] ), .S0(n462), .S1(n369), .Y(n613) );
  MUX41X1_HVT U618 ( .A1(\ram[8][2] ), .A3(\ram[10][2] ), .A2(\ram[9][2] ), 
        .A4(\ram[11][2] ), .S0(n462), .S1(n369), .Y(n614) );
  MUX41X1_HVT U619 ( .A1(\ram[4][2] ), .A3(\ram[6][2] ), .A2(\ram[5][2] ), 
        .A4(\ram[7][2] ), .S0(n462), .S1(n369), .Y(n615) );
  MUX41X1_HVT U620 ( .A1(\ram[0][2] ), .A3(\ram[2][2] ), .A2(\ram[1][2] ), 
        .A4(\ram[3][2] ), .S0(n462), .S1(n369), .Y(n616) );
  MUX41X1_HVT U621 ( .A1(n616), .A3(n614), .A2(n615), .A4(n613), .S0(n580), 
        .S1(n567), .Y(q[2]) );
  MUX41X1_HVT U622 ( .A1(\ram[12][3] ), .A3(\ram[14][3] ), .A2(\ram[13][3] ), 
        .A4(\ram[15][3] ), .S0(n463), .S1(n370), .Y(n617) );
  MUX41X1_HVT U623 ( .A1(\ram[8][3] ), .A3(\ram[10][3] ), .A2(\ram[9][3] ), 
        .A4(\ram[11][3] ), .S0(n463), .S1(n370), .Y(n618) );
  MUX41X1_HVT U624 ( .A1(\ram[4][3] ), .A3(\ram[6][3] ), .A2(\ram[5][3] ), 
        .A4(\ram[7][3] ), .S0(n463), .S1(n370), .Y(n619) );
  MUX41X1_HVT U625 ( .A1(\ram[0][3] ), .A3(\ram[2][3] ), .A2(\ram[1][3] ), 
        .A4(\ram[3][3] ), .S0(n463), .S1(n370), .Y(n620) );
  MUX41X1_HVT U626 ( .A1(n620), .A3(n618), .A2(n619), .A4(n617), .S0(n580), 
        .S1(n567), .Y(q[3]) );
  MUX41X1_HVT U627 ( .A1(\ram[12][4] ), .A3(\ram[14][4] ), .A2(\ram[13][4] ), 
        .A4(\ram[15][4] ), .S0(n463), .S1(n370), .Y(n621) );
  MUX41X1_HVT U628 ( .A1(\ram[8][4] ), .A3(\ram[10][4] ), .A2(\ram[9][4] ), 
        .A4(\ram[11][4] ), .S0(n463), .S1(n370), .Y(n622) );
  MUX41X1_HVT U629 ( .A1(\ram[4][4] ), .A3(\ram[6][4] ), .A2(\ram[5][4] ), 
        .A4(\ram[7][4] ), .S0(n463), .S1(n370), .Y(n623) );
  MUX41X1_HVT U630 ( .A1(\ram[0][4] ), .A3(\ram[2][4] ), .A2(\ram[1][4] ), 
        .A4(\ram[3][4] ), .S0(n463), .S1(n370), .Y(n624) );
  MUX41X1_HVT U631 ( .A1(n624), .A3(n622), .A2(n623), .A4(n621), .S0(n580), 
        .S1(n567), .Y(q[4]) );
  MUX41X1_HVT U632 ( .A1(\ram[12][5] ), .A3(\ram[14][5] ), .A2(\ram[13][5] ), 
        .A4(\ram[15][5] ), .S0(n463), .S1(n370), .Y(n625) );
  MUX41X1_HVT U633 ( .A1(\ram[8][5] ), .A3(\ram[10][5] ), .A2(\ram[9][5] ), 
        .A4(\ram[11][5] ), .S0(n463), .S1(n370), .Y(n626) );
  MUX41X1_HVT U634 ( .A1(\ram[4][5] ), .A3(\ram[6][5] ), .A2(\ram[5][5] ), 
        .A4(\ram[7][5] ), .S0(n463), .S1(n370), .Y(n627) );
  MUX41X1_HVT U635 ( .A1(\ram[0][5] ), .A3(\ram[2][5] ), .A2(\ram[1][5] ), 
        .A4(\ram[3][5] ), .S0(n463), .S1(n370), .Y(n628) );
  MUX41X1_HVT U636 ( .A1(n628), .A3(n626), .A2(n627), .A4(n625), .S0(n580), 
        .S1(n568), .Y(q[5]) );
  MUX41X1_HVT U637 ( .A1(\ram[12][6] ), .A3(\ram[14][6] ), .A2(\ram[13][6] ), 
        .A4(\ram[15][6] ), .S0(n464), .S1(n371), .Y(n629) );
  MUX41X1_HVT U638 ( .A1(\ram[8][6] ), .A3(\ram[10][6] ), .A2(\ram[9][6] ), 
        .A4(\ram[11][6] ), .S0(n464), .S1(n371), .Y(n630) );
  MUX41X1_HVT U639 ( .A1(\ram[4][6] ), .A3(\ram[6][6] ), .A2(\ram[5][6] ), 
        .A4(\ram[7][6] ), .S0(n464), .S1(n371), .Y(n631) );
  MUX41X1_HVT U640 ( .A1(\ram[0][6] ), .A3(\ram[2][6] ), .A2(\ram[1][6] ), 
        .A4(\ram[3][6] ), .S0(n464), .S1(n371), .Y(n632) );
  MUX41X1_HVT U641 ( .A1(n632), .A3(n630), .A2(n631), .A4(n629), .S0(n580), 
        .S1(n568), .Y(q[6]) );
  MUX41X1_HVT U642 ( .A1(\ram[12][7] ), .A3(\ram[14][7] ), .A2(\ram[13][7] ), 
        .A4(\ram[15][7] ), .S0(n464), .S1(n371), .Y(n633) );
  MUX41X1_HVT U643 ( .A1(\ram[8][7] ), .A3(\ram[10][7] ), .A2(\ram[9][7] ), 
        .A4(\ram[11][7] ), .S0(n464), .S1(n371), .Y(n634) );
  MUX41X1_HVT U644 ( .A1(\ram[4][7] ), .A3(\ram[6][7] ), .A2(\ram[5][7] ), 
        .A4(\ram[7][7] ), .S0(n464), .S1(n371), .Y(n635) );
  MUX41X1_HVT U645 ( .A1(\ram[0][7] ), .A3(\ram[2][7] ), .A2(\ram[1][7] ), 
        .A4(\ram[3][7] ), .S0(n464), .S1(n371), .Y(n636) );
  MUX41X1_HVT U646 ( .A1(n636), .A3(n634), .A2(n635), .A4(n633), .S0(n580), 
        .S1(n568), .Y(q[7]) );
  MUX41X1_HVT U647 ( .A1(\ram[12][8] ), .A3(\ram[14][8] ), .A2(\ram[13][8] ), 
        .A4(\ram[15][8] ), .S0(n464), .S1(n371), .Y(n637) );
  MUX41X1_HVT U648 ( .A1(\ram[8][8] ), .A3(\ram[10][8] ), .A2(\ram[9][8] ), 
        .A4(\ram[11][8] ), .S0(n464), .S1(n371), .Y(n638) );
  MUX41X1_HVT U649 ( .A1(\ram[4][8] ), .A3(\ram[6][8] ), .A2(\ram[5][8] ), 
        .A4(\ram[7][8] ), .S0(n464), .S1(n371), .Y(n639) );
  MUX41X1_HVT U650 ( .A1(\ram[0][8] ), .A3(\ram[2][8] ), .A2(\ram[1][8] ), 
        .A4(\ram[3][8] ), .S0(n464), .S1(n371), .Y(n640) );
  MUX41X1_HVT U651 ( .A1(n640), .A3(n638), .A2(n639), .A4(n637), .S0(n580), 
        .S1(n568), .Y(q[8]) );
  MUX41X1_HVT U652 ( .A1(\ram[12][9] ), .A3(\ram[14][9] ), .A2(\ram[13][9] ), 
        .A4(\ram[15][9] ), .S0(n465), .S1(n372), .Y(n641) );
  MUX41X1_HVT U653 ( .A1(\ram[8][9] ), .A3(\ram[10][9] ), .A2(\ram[9][9] ), 
        .A4(\ram[11][9] ), .S0(n465), .S1(n372), .Y(n642) );
  MUX41X1_HVT U654 ( .A1(\ram[4][9] ), .A3(\ram[6][9] ), .A2(\ram[5][9] ), 
        .A4(\ram[7][9] ), .S0(n465), .S1(n372), .Y(n643) );
  MUX41X1_HVT U655 ( .A1(\ram[0][9] ), .A3(\ram[2][9] ), .A2(\ram[1][9] ), 
        .A4(\ram[3][9] ), .S0(n465), .S1(n372), .Y(n644) );
  MUX41X1_HVT U656 ( .A1(n644), .A3(n642), .A2(n643), .A4(n641), .S0(n580), 
        .S1(n568), .Y(q[9]) );
  MUX41X1_HVT U657 ( .A1(\ram[12][10] ), .A3(\ram[14][10] ), .A2(\ram[13][10] ), .A4(\ram[15][10] ), .S0(n465), .S1(n372), .Y(n645) );
  MUX41X1_HVT U658 ( .A1(\ram[8][10] ), .A3(\ram[10][10] ), .A2(\ram[9][10] ), 
        .A4(\ram[11][10] ), .S0(n465), .S1(n372), .Y(n646) );
  MUX41X1_HVT U659 ( .A1(\ram[4][10] ), .A3(\ram[6][10] ), .A2(\ram[5][10] ), 
        .A4(\ram[7][10] ), .S0(n465), .S1(n372), .Y(n647) );
  MUX41X1_HVT U660 ( .A1(\ram[0][10] ), .A3(\ram[2][10] ), .A2(\ram[1][10] ), 
        .A4(\ram[3][10] ), .S0(n465), .S1(n372), .Y(n648) );
  MUX41X1_HVT U661 ( .A1(n648), .A3(n646), .A2(n647), .A4(n645), .S0(n580), 
        .S1(n568), .Y(q[10]) );
  MUX41X1_HVT U662 ( .A1(\ram[12][11] ), .A3(\ram[14][11] ), .A2(\ram[13][11] ), .A4(\ram[15][11] ), .S0(n465), .S1(n372), .Y(n649) );
  MUX41X1_HVT U663 ( .A1(\ram[8][11] ), .A3(\ram[10][11] ), .A2(\ram[9][11] ), 
        .A4(\ram[11][11] ), .S0(n465), .S1(n372), .Y(n650) );
  MUX41X1_HVT U664 ( .A1(\ram[4][11] ), .A3(\ram[6][11] ), .A2(\ram[5][11] ), 
        .A4(\ram[7][11] ), .S0(n465), .S1(n372), .Y(n651) );
  MUX41X1_HVT U665 ( .A1(\ram[0][11] ), .A3(\ram[2][11] ), .A2(\ram[1][11] ), 
        .A4(\ram[3][11] ), .S0(n465), .S1(n372), .Y(n652) );
  MUX41X1_HVT U666 ( .A1(n652), .A3(n650), .A2(n651), .A4(n649), .S0(n580), 
        .S1(n568), .Y(q[11]) );
  MUX41X1_HVT U667 ( .A1(\ram[12][12] ), .A3(\ram[14][12] ), .A2(\ram[13][12] ), .A4(\ram[15][12] ), .S0(n466), .S1(n373), .Y(n653) );
  MUX41X1_HVT U668 ( .A1(\ram[8][12] ), .A3(\ram[10][12] ), .A2(\ram[9][12] ), 
        .A4(\ram[11][12] ), .S0(n466), .S1(n373), .Y(n654) );
  MUX41X1_HVT U669 ( .A1(\ram[4][12] ), .A3(\ram[6][12] ), .A2(\ram[5][12] ), 
        .A4(\ram[7][12] ), .S0(n466), .S1(n373), .Y(n655) );
  MUX41X1_HVT U670 ( .A1(\ram[0][12] ), .A3(\ram[2][12] ), .A2(\ram[1][12] ), 
        .A4(\ram[3][12] ), .S0(n466), .S1(n373), .Y(n656) );
  MUX41X1_HVT U671 ( .A1(n656), .A3(n654), .A2(n655), .A4(n653), .S0(n581), 
        .S1(n568), .Y(q[12]) );
  MUX41X1_HVT U672 ( .A1(\ram[12][13] ), .A3(\ram[14][13] ), .A2(\ram[13][13] ), .A4(\ram[15][13] ), .S0(n466), .S1(n373), .Y(n657) );
  MUX41X1_HVT U673 ( .A1(\ram[8][13] ), .A3(\ram[10][13] ), .A2(\ram[9][13] ), 
        .A4(\ram[11][13] ), .S0(n466), .S1(n373), .Y(n658) );
  MUX41X1_HVT U674 ( .A1(\ram[4][13] ), .A3(\ram[6][13] ), .A2(\ram[5][13] ), 
        .A4(\ram[7][13] ), .S0(n466), .S1(n373), .Y(n659) );
  MUX41X1_HVT U675 ( .A1(\ram[0][13] ), .A3(\ram[2][13] ), .A2(\ram[1][13] ), 
        .A4(\ram[3][13] ), .S0(n466), .S1(n373), .Y(n660) );
  MUX41X1_HVT U676 ( .A1(n660), .A3(n658), .A2(n659), .A4(n657), .S0(n581), 
        .S1(n568), .Y(q[13]) );
  MUX41X1_HVT U677 ( .A1(\ram[12][14] ), .A3(\ram[14][14] ), .A2(\ram[13][14] ), .A4(\ram[15][14] ), .S0(n466), .S1(n373), .Y(n661) );
  MUX41X1_HVT U678 ( .A1(\ram[8][14] ), .A3(\ram[10][14] ), .A2(\ram[9][14] ), 
        .A4(\ram[11][14] ), .S0(n466), .S1(n373), .Y(n662) );
  MUX41X1_HVT U679 ( .A1(\ram[4][14] ), .A3(\ram[6][14] ), .A2(\ram[5][14] ), 
        .A4(\ram[7][14] ), .S0(n466), .S1(n373), .Y(n663) );
  MUX41X1_HVT U680 ( .A1(\ram[0][14] ), .A3(\ram[2][14] ), .A2(\ram[1][14] ), 
        .A4(\ram[3][14] ), .S0(n466), .S1(n373), .Y(n664) );
  MUX41X1_HVT U681 ( .A1(n664), .A3(n662), .A2(n663), .A4(n661), .S0(n581), 
        .S1(n568), .Y(q[14]) );
  MUX41X1_HVT U682 ( .A1(\ram[12][15] ), .A3(\ram[14][15] ), .A2(\ram[13][15] ), .A4(\ram[15][15] ), .S0(n467), .S1(n374), .Y(n665) );
  MUX41X1_HVT U683 ( .A1(\ram[8][15] ), .A3(\ram[10][15] ), .A2(\ram[9][15] ), 
        .A4(\ram[11][15] ), .S0(n467), .S1(n374), .Y(n666) );
  MUX41X1_HVT U684 ( .A1(\ram[4][15] ), .A3(\ram[6][15] ), .A2(\ram[5][15] ), 
        .A4(\ram[7][15] ), .S0(n467), .S1(n374), .Y(n667) );
  MUX41X1_HVT U685 ( .A1(\ram[0][15] ), .A3(\ram[2][15] ), .A2(\ram[1][15] ), 
        .A4(\ram[3][15] ), .S0(n467), .S1(n374), .Y(n668) );
  MUX41X1_HVT U686 ( .A1(n668), .A3(n666), .A2(n667), .A4(n665), .S0(n581), 
        .S1(n568), .Y(q[15]) );
  MUX41X1_HVT U687 ( .A1(\ram[12][16] ), .A3(\ram[14][16] ), .A2(\ram[13][16] ), .A4(\ram[15][16] ), .S0(n467), .S1(n374), .Y(n669) );
  MUX41X1_HVT U688 ( .A1(\ram[8][16] ), .A3(\ram[10][16] ), .A2(\ram[9][16] ), 
        .A4(\ram[11][16] ), .S0(n467), .S1(n374), .Y(n670) );
  MUX41X1_HVT U689 ( .A1(\ram[4][16] ), .A3(\ram[6][16] ), .A2(\ram[5][16] ), 
        .A4(\ram[7][16] ), .S0(n467), .S1(n374), .Y(n671) );
  MUX41X1_HVT U690 ( .A1(\ram[0][16] ), .A3(\ram[2][16] ), .A2(\ram[1][16] ), 
        .A4(\ram[3][16] ), .S0(n467), .S1(n374), .Y(n672) );
  MUX41X1_HVT U691 ( .A1(n672), .A3(n670), .A2(n671), .A4(n669), .S0(n581), 
        .S1(n568), .Y(q[16]) );
  MUX41X1_HVT U692 ( .A1(\ram[12][17] ), .A3(\ram[14][17] ), .A2(\ram[13][17] ), .A4(\ram[15][17] ), .S0(n467), .S1(n374), .Y(n673) );
  MUX41X1_HVT U693 ( .A1(\ram[8][17] ), .A3(\ram[10][17] ), .A2(\ram[9][17] ), 
        .A4(\ram[11][17] ), .S0(n467), .S1(n374), .Y(n674) );
  MUX41X1_HVT U694 ( .A1(\ram[4][17] ), .A3(\ram[6][17] ), .A2(\ram[5][17] ), 
        .A4(\ram[7][17] ), .S0(n467), .S1(n374), .Y(n675) );
  MUX41X1_HVT U695 ( .A1(\ram[0][17] ), .A3(\ram[2][17] ), .A2(\ram[1][17] ), 
        .A4(\ram[3][17] ), .S0(n467), .S1(n374), .Y(n676) );
  MUX41X1_HVT U696 ( .A1(n676), .A3(n674), .A2(n675), .A4(n673), .S0(n581), 
        .S1(n569), .Y(q[17]) );
  MUX41X1_HVT U697 ( .A1(\ram[12][18] ), .A3(\ram[14][18] ), .A2(\ram[13][18] ), .A4(\ram[15][18] ), .S0(n468), .S1(n375), .Y(n677) );
  MUX41X1_HVT U698 ( .A1(\ram[8][18] ), .A3(\ram[10][18] ), .A2(\ram[9][18] ), 
        .A4(\ram[11][18] ), .S0(n468), .S1(n375), .Y(n678) );
  MUX41X1_HVT U699 ( .A1(\ram[4][18] ), .A3(\ram[6][18] ), .A2(\ram[5][18] ), 
        .A4(\ram[7][18] ), .S0(n468), .S1(n375), .Y(n679) );
  MUX41X1_HVT U700 ( .A1(\ram[0][18] ), .A3(\ram[2][18] ), .A2(\ram[1][18] ), 
        .A4(\ram[3][18] ), .S0(n468), .S1(n375), .Y(n680) );
  MUX41X1_HVT U701 ( .A1(n680), .A3(n678), .A2(n679), .A4(n677), .S0(n581), 
        .S1(n569), .Y(q[18]) );
  MUX41X1_HVT U702 ( .A1(\ram[12][19] ), .A3(\ram[14][19] ), .A2(\ram[13][19] ), .A4(\ram[15][19] ), .S0(n468), .S1(n375), .Y(n681) );
  MUX41X1_HVT U703 ( .A1(\ram[8][19] ), .A3(\ram[10][19] ), .A2(\ram[9][19] ), 
        .A4(\ram[11][19] ), .S0(n468), .S1(n375), .Y(n682) );
  MUX41X1_HVT U704 ( .A1(\ram[4][19] ), .A3(\ram[6][19] ), .A2(\ram[5][19] ), 
        .A4(\ram[7][19] ), .S0(n468), .S1(n375), .Y(n683) );
  MUX41X1_HVT U705 ( .A1(\ram[0][19] ), .A3(\ram[2][19] ), .A2(\ram[1][19] ), 
        .A4(\ram[3][19] ), .S0(n468), .S1(n375), .Y(n684) );
  MUX41X1_HVT U706 ( .A1(n684), .A3(n682), .A2(n683), .A4(n681), .S0(n581), 
        .S1(n569), .Y(q[19]) );
  MUX41X1_HVT U707 ( .A1(\ram[12][20] ), .A3(\ram[14][20] ), .A2(\ram[13][20] ), .A4(\ram[15][20] ), .S0(n468), .S1(n375), .Y(n685) );
  MUX41X1_HVT U708 ( .A1(\ram[8][20] ), .A3(\ram[10][20] ), .A2(\ram[9][20] ), 
        .A4(\ram[11][20] ), .S0(n468), .S1(n375), .Y(n686) );
  MUX41X1_HVT U709 ( .A1(\ram[4][20] ), .A3(\ram[6][20] ), .A2(\ram[5][20] ), 
        .A4(\ram[7][20] ), .S0(n468), .S1(n375), .Y(n687) );
  MUX41X1_HVT U710 ( .A1(\ram[0][20] ), .A3(\ram[2][20] ), .A2(\ram[1][20] ), 
        .A4(\ram[3][20] ), .S0(n468), .S1(n375), .Y(n688) );
  MUX41X1_HVT U711 ( .A1(n688), .A3(n686), .A2(n687), .A4(n685), .S0(n581), 
        .S1(n569), .Y(q[20]) );
  MUX41X1_HVT U712 ( .A1(\ram[12][21] ), .A3(\ram[14][21] ), .A2(\ram[13][21] ), .A4(\ram[15][21] ), .S0(n469), .S1(n376), .Y(n689) );
  MUX41X1_HVT U713 ( .A1(\ram[8][21] ), .A3(\ram[10][21] ), .A2(\ram[9][21] ), 
        .A4(\ram[11][21] ), .S0(n469), .S1(n376), .Y(n690) );
  MUX41X1_HVT U714 ( .A1(\ram[4][21] ), .A3(\ram[6][21] ), .A2(\ram[5][21] ), 
        .A4(\ram[7][21] ), .S0(n469), .S1(n376), .Y(n691) );
  MUX41X1_HVT U715 ( .A1(\ram[0][21] ), .A3(\ram[2][21] ), .A2(\ram[1][21] ), 
        .A4(\ram[3][21] ), .S0(n469), .S1(n376), .Y(n692) );
  MUX41X1_HVT U716 ( .A1(n692), .A3(n690), .A2(n691), .A4(n689), .S0(n581), 
        .S1(n569), .Y(q[21]) );
  MUX41X1_HVT U717 ( .A1(\ram[12][22] ), .A3(\ram[14][22] ), .A2(\ram[13][22] ), .A4(\ram[15][22] ), .S0(n469), .S1(n376), .Y(n693) );
  MUX41X1_HVT U718 ( .A1(\ram[8][22] ), .A3(\ram[10][22] ), .A2(\ram[9][22] ), 
        .A4(\ram[11][22] ), .S0(n469), .S1(n376), .Y(n694) );
  MUX41X1_HVT U719 ( .A1(\ram[4][22] ), .A3(\ram[6][22] ), .A2(\ram[5][22] ), 
        .A4(\ram[7][22] ), .S0(n469), .S1(n376), .Y(n695) );
  MUX41X1_HVT U720 ( .A1(\ram[0][22] ), .A3(\ram[2][22] ), .A2(\ram[1][22] ), 
        .A4(\ram[3][22] ), .S0(n469), .S1(n376), .Y(n696) );
  MUX41X1_HVT U721 ( .A1(n696), .A3(n694), .A2(n695), .A4(n693), .S0(n581), 
        .S1(n569), .Y(q[22]) );
  MUX41X1_HVT U722 ( .A1(\ram[12][23] ), .A3(\ram[14][23] ), .A2(\ram[13][23] ), .A4(\ram[15][23] ), .S0(n469), .S1(n376), .Y(n697) );
  MUX41X1_HVT U723 ( .A1(\ram[8][23] ), .A3(\ram[10][23] ), .A2(\ram[9][23] ), 
        .A4(\ram[11][23] ), .S0(n469), .S1(n376), .Y(n698) );
  MUX41X1_HVT U724 ( .A1(\ram[4][23] ), .A3(\ram[6][23] ), .A2(\ram[5][23] ), 
        .A4(\ram[7][23] ), .S0(n469), .S1(n376), .Y(n699) );
  MUX41X1_HVT U725 ( .A1(\ram[0][23] ), .A3(\ram[2][23] ), .A2(\ram[1][23] ), 
        .A4(\ram[3][23] ), .S0(n469), .S1(n376), .Y(n700) );
  MUX41X1_HVT U726 ( .A1(n700), .A3(n698), .A2(n699), .A4(n697), .S0(n581), 
        .S1(n569), .Y(q[23]) );
  MUX41X1_HVT U727 ( .A1(\ram[12][24] ), .A3(\ram[14][24] ), .A2(\ram[13][24] ), .A4(\ram[15][24] ), .S0(n470), .S1(n377), .Y(n701) );
  MUX41X1_HVT U728 ( .A1(\ram[8][24] ), .A3(\ram[10][24] ), .A2(\ram[9][24] ), 
        .A4(\ram[11][24] ), .S0(n470), .S1(n377), .Y(n702) );
  MUX41X1_HVT U729 ( .A1(\ram[4][24] ), .A3(\ram[6][24] ), .A2(\ram[5][24] ), 
        .A4(\ram[7][24] ), .S0(n470), .S1(n377), .Y(n703) );
  MUX41X1_HVT U730 ( .A1(\ram[0][24] ), .A3(\ram[2][24] ), .A2(\ram[1][24] ), 
        .A4(\ram[3][24] ), .S0(n470), .S1(n377), .Y(n704) );
  MUX41X1_HVT U731 ( .A1(n704), .A3(n702), .A2(n703), .A4(n701), .S0(n582), 
        .S1(n569), .Y(q[24]) );
  MUX41X1_HVT U732 ( .A1(\ram[12][25] ), .A3(\ram[14][25] ), .A2(\ram[13][25] ), .A4(\ram[15][25] ), .S0(n470), .S1(n377), .Y(n705) );
  MUX41X1_HVT U733 ( .A1(\ram[8][25] ), .A3(\ram[10][25] ), .A2(\ram[9][25] ), 
        .A4(\ram[11][25] ), .S0(n470), .S1(n377), .Y(n706) );
  MUX41X1_HVT U734 ( .A1(\ram[4][25] ), .A3(\ram[6][25] ), .A2(\ram[5][25] ), 
        .A4(\ram[7][25] ), .S0(n470), .S1(n377), .Y(n707) );
  MUX41X1_HVT U735 ( .A1(\ram[0][25] ), .A3(\ram[2][25] ), .A2(\ram[1][25] ), 
        .A4(\ram[3][25] ), .S0(n470), .S1(n377), .Y(n708) );
  MUX41X1_HVT U736 ( .A1(n708), .A3(n706), .A2(n707), .A4(n705), .S0(n582), 
        .S1(n569), .Y(q[25]) );
  MUX41X1_HVT U737 ( .A1(\ram[12][26] ), .A3(\ram[14][26] ), .A2(\ram[13][26] ), .A4(\ram[15][26] ), .S0(n470), .S1(n377), .Y(n709) );
  MUX41X1_HVT U738 ( .A1(\ram[8][26] ), .A3(\ram[10][26] ), .A2(\ram[9][26] ), 
        .A4(\ram[11][26] ), .S0(n470), .S1(n377), .Y(n710) );
  MUX41X1_HVT U739 ( .A1(\ram[4][26] ), .A3(\ram[6][26] ), .A2(\ram[5][26] ), 
        .A4(\ram[7][26] ), .S0(n470), .S1(n377), .Y(n711) );
  MUX41X1_HVT U740 ( .A1(\ram[0][26] ), .A3(\ram[2][26] ), .A2(\ram[1][26] ), 
        .A4(\ram[3][26] ), .S0(n470), .S1(n377), .Y(n712) );
  MUX41X1_HVT U741 ( .A1(n712), .A3(n710), .A2(n711), .A4(n709), .S0(n582), 
        .S1(n569), .Y(q[26]) );
  MUX41X1_HVT U742 ( .A1(\ram[12][27] ), .A3(\ram[14][27] ), .A2(\ram[13][27] ), .A4(\ram[15][27] ), .S0(n471), .S1(n378), .Y(n713) );
  MUX41X1_HVT U743 ( .A1(\ram[8][27] ), .A3(\ram[10][27] ), .A2(\ram[9][27] ), 
        .A4(\ram[11][27] ), .S0(n471), .S1(n378), .Y(n714) );
  MUX41X1_HVT U744 ( .A1(\ram[4][27] ), .A3(\ram[6][27] ), .A2(\ram[5][27] ), 
        .A4(\ram[7][27] ), .S0(n471), .S1(n378), .Y(n715) );
  MUX41X1_HVT U745 ( .A1(\ram[0][27] ), .A3(\ram[2][27] ), .A2(\ram[1][27] ), 
        .A4(\ram[3][27] ), .S0(n471), .S1(n378), .Y(n716) );
  MUX41X1_HVT U746 ( .A1(n716), .A3(n714), .A2(n715), .A4(n713), .S0(n582), 
        .S1(n569), .Y(q[27]) );
  MUX41X1_HVT U747 ( .A1(\ram[12][28] ), .A3(\ram[14][28] ), .A2(\ram[13][28] ), .A4(\ram[15][28] ), .S0(n471), .S1(n378), .Y(n717) );
  MUX41X1_HVT U748 ( .A1(\ram[8][28] ), .A3(\ram[10][28] ), .A2(\ram[9][28] ), 
        .A4(\ram[11][28] ), .S0(n471), .S1(n378), .Y(n718) );
  MUX41X1_HVT U749 ( .A1(\ram[4][28] ), .A3(\ram[6][28] ), .A2(\ram[5][28] ), 
        .A4(\ram[7][28] ), .S0(n471), .S1(n378), .Y(n719) );
  MUX41X1_HVT U750 ( .A1(\ram[0][28] ), .A3(\ram[2][28] ), .A2(\ram[1][28] ), 
        .A4(\ram[3][28] ), .S0(n471), .S1(n378), .Y(n720) );
  MUX41X1_HVT U751 ( .A1(n720), .A3(n718), .A2(n719), .A4(n717), .S0(n582), 
        .S1(n569), .Y(q[28]) );
  MUX41X1_HVT U752 ( .A1(\ram[12][29] ), .A3(\ram[14][29] ), .A2(\ram[13][29] ), .A4(\ram[15][29] ), .S0(n471), .S1(n378), .Y(n721) );
  MUX41X1_HVT U753 ( .A1(\ram[8][29] ), .A3(\ram[10][29] ), .A2(\ram[9][29] ), 
        .A4(\ram[11][29] ), .S0(n471), .S1(n378), .Y(n722) );
  MUX41X1_HVT U754 ( .A1(\ram[4][29] ), .A3(\ram[6][29] ), .A2(\ram[5][29] ), 
        .A4(\ram[7][29] ), .S0(n471), .S1(n378), .Y(n723) );
  MUX41X1_HVT U755 ( .A1(\ram[0][29] ), .A3(\ram[2][29] ), .A2(\ram[1][29] ), 
        .A4(\ram[3][29] ), .S0(n471), .S1(n378), .Y(n724) );
  MUX41X1_HVT U756 ( .A1(n724), .A3(n722), .A2(n723), .A4(n721), .S0(n582), 
        .S1(n570), .Y(q[29]) );
  MUX41X1_HVT U757 ( .A1(\ram[12][30] ), .A3(\ram[14][30] ), .A2(\ram[13][30] ), .A4(\ram[15][30] ), .S0(n472), .S1(n379), .Y(n725) );
  MUX41X1_HVT U758 ( .A1(\ram[8][30] ), .A3(\ram[10][30] ), .A2(\ram[9][30] ), 
        .A4(\ram[11][30] ), .S0(n472), .S1(n379), .Y(n726) );
  MUX41X1_HVT U759 ( .A1(\ram[4][30] ), .A3(\ram[6][30] ), .A2(\ram[5][30] ), 
        .A4(\ram[7][30] ), .S0(n472), .S1(n379), .Y(n727) );
  MUX41X1_HVT U760 ( .A1(\ram[0][30] ), .A3(\ram[2][30] ), .A2(\ram[1][30] ), 
        .A4(\ram[3][30] ), .S0(n472), .S1(n379), .Y(n728) );
  MUX41X1_HVT U761 ( .A1(n728), .A3(n726), .A2(n727), .A4(n725), .S0(n582), 
        .S1(n570), .Y(q[30]) );
  MUX41X1_HVT U762 ( .A1(\ram[12][31] ), .A3(\ram[14][31] ), .A2(\ram[13][31] ), .A4(\ram[15][31] ), .S0(n472), .S1(n379), .Y(n729) );
  MUX41X1_HVT U763 ( .A1(\ram[8][31] ), .A3(\ram[10][31] ), .A2(\ram[9][31] ), 
        .A4(\ram[11][31] ), .S0(n472), .S1(n379), .Y(n730) );
  MUX41X1_HVT U764 ( .A1(\ram[4][31] ), .A3(\ram[6][31] ), .A2(\ram[5][31] ), 
        .A4(\ram[7][31] ), .S0(n472), .S1(n379), .Y(n731) );
  MUX41X1_HVT U765 ( .A1(\ram[0][31] ), .A3(\ram[2][31] ), .A2(\ram[1][31] ), 
        .A4(\ram[3][31] ), .S0(n472), .S1(n379), .Y(n732) );
  MUX41X1_HVT U766 ( .A1(n732), .A3(n730), .A2(n731), .A4(n729), .S0(n582), 
        .S1(n570), .Y(q[31]) );
  MUX41X1_HVT U767 ( .A1(\ram[12][32] ), .A3(\ram[14][32] ), .A2(\ram[13][32] ), .A4(\ram[15][32] ), .S0(n472), .S1(n379), .Y(n733) );
  MUX41X1_HVT U768 ( .A1(\ram[8][32] ), .A3(\ram[10][32] ), .A2(\ram[9][32] ), 
        .A4(\ram[11][32] ), .S0(n472), .S1(n379), .Y(n734) );
  MUX41X1_HVT U769 ( .A1(\ram[4][32] ), .A3(\ram[6][32] ), .A2(\ram[5][32] ), 
        .A4(\ram[7][32] ), .S0(n472), .S1(n379), .Y(n735) );
  MUX41X1_HVT U770 ( .A1(\ram[0][32] ), .A3(\ram[2][32] ), .A2(\ram[1][32] ), 
        .A4(\ram[3][32] ), .S0(n472), .S1(n379), .Y(n736) );
  MUX41X1_HVT U771 ( .A1(n736), .A3(n734), .A2(n735), .A4(n733), .S0(n582), 
        .S1(n570), .Y(q[32]) );
  MUX41X1_HVT U772 ( .A1(\ram[12][33] ), .A3(\ram[14][33] ), .A2(\ram[13][33] ), .A4(\ram[15][33] ), .S0(n473), .S1(n380), .Y(n737) );
  MUX41X1_HVT U773 ( .A1(\ram[8][33] ), .A3(\ram[10][33] ), .A2(\ram[9][33] ), 
        .A4(\ram[11][33] ), .S0(n473), .S1(n380), .Y(n738) );
  MUX41X1_HVT U774 ( .A1(\ram[4][33] ), .A3(\ram[6][33] ), .A2(\ram[5][33] ), 
        .A4(\ram[7][33] ), .S0(n473), .S1(n380), .Y(n739) );
  MUX41X1_HVT U775 ( .A1(\ram[0][33] ), .A3(\ram[2][33] ), .A2(\ram[1][33] ), 
        .A4(\ram[3][33] ), .S0(n473), .S1(n380), .Y(n740) );
  MUX41X1_HVT U776 ( .A1(n740), .A3(n738), .A2(n739), .A4(n737), .S0(n582), 
        .S1(n570), .Y(q[33]) );
  MUX41X1_HVT U777 ( .A1(\ram[12][34] ), .A3(\ram[14][34] ), .A2(\ram[13][34] ), .A4(\ram[15][34] ), .S0(n473), .S1(n380), .Y(n741) );
  MUX41X1_HVT U778 ( .A1(\ram[8][34] ), .A3(\ram[10][34] ), .A2(\ram[9][34] ), 
        .A4(\ram[11][34] ), .S0(n473), .S1(n380), .Y(n742) );
  MUX41X1_HVT U779 ( .A1(\ram[4][34] ), .A3(\ram[6][34] ), .A2(\ram[5][34] ), 
        .A4(\ram[7][34] ), .S0(n473), .S1(n380), .Y(n743) );
  MUX41X1_HVT U780 ( .A1(\ram[0][34] ), .A3(\ram[2][34] ), .A2(\ram[1][34] ), 
        .A4(\ram[3][34] ), .S0(n473), .S1(n380), .Y(n744) );
  MUX41X1_HVT U781 ( .A1(n744), .A3(n742), .A2(n743), .A4(n741), .S0(n582), 
        .S1(n570), .Y(q[34]) );
  MUX41X1_HVT U782 ( .A1(\ram[12][35] ), .A3(\ram[14][35] ), .A2(\ram[13][35] ), .A4(\ram[15][35] ), .S0(n473), .S1(n380), .Y(n745) );
  MUX41X1_HVT U783 ( .A1(\ram[8][35] ), .A3(\ram[10][35] ), .A2(\ram[9][35] ), 
        .A4(\ram[11][35] ), .S0(n473), .S1(n380), .Y(n746) );
  MUX41X1_HVT U784 ( .A1(\ram[4][35] ), .A3(\ram[6][35] ), .A2(\ram[5][35] ), 
        .A4(\ram[7][35] ), .S0(n473), .S1(n380), .Y(n747) );
  MUX41X1_HVT U785 ( .A1(\ram[0][35] ), .A3(\ram[2][35] ), .A2(\ram[1][35] ), 
        .A4(\ram[3][35] ), .S0(n473), .S1(n380), .Y(n748) );
  MUX41X1_HVT U786 ( .A1(n748), .A3(n746), .A2(n747), .A4(n745), .S0(n582), 
        .S1(n570), .Y(q[35]) );
  MUX41X1_HVT U787 ( .A1(\ram[12][36] ), .A3(\ram[14][36] ), .A2(\ram[13][36] ), .A4(\ram[15][36] ), .S0(n474), .S1(n381), .Y(n749) );
  MUX41X1_HVT U788 ( .A1(\ram[8][36] ), .A3(\ram[10][36] ), .A2(\ram[9][36] ), 
        .A4(\ram[11][36] ), .S0(n474), .S1(n381), .Y(n750) );
  MUX41X1_HVT U789 ( .A1(\ram[4][36] ), .A3(\ram[6][36] ), .A2(\ram[5][36] ), 
        .A4(\ram[7][36] ), .S0(n474), .S1(n381), .Y(n751) );
  MUX41X1_HVT U790 ( .A1(\ram[0][36] ), .A3(\ram[2][36] ), .A2(\ram[1][36] ), 
        .A4(\ram[3][36] ), .S0(n474), .S1(n381), .Y(n752) );
  MUX41X1_HVT U791 ( .A1(n752), .A3(n750), .A2(n751), .A4(n749), .S0(n583), 
        .S1(n570), .Y(q[36]) );
  MUX41X1_HVT U792 ( .A1(\ram[12][37] ), .A3(\ram[14][37] ), .A2(\ram[13][37] ), .A4(\ram[15][37] ), .S0(n474), .S1(n381), .Y(n753) );
  MUX41X1_HVT U793 ( .A1(\ram[8][37] ), .A3(\ram[10][37] ), .A2(\ram[9][37] ), 
        .A4(\ram[11][37] ), .S0(n474), .S1(n381), .Y(n754) );
  MUX41X1_HVT U794 ( .A1(\ram[4][37] ), .A3(\ram[6][37] ), .A2(\ram[5][37] ), 
        .A4(\ram[7][37] ), .S0(n474), .S1(n381), .Y(n755) );
  MUX41X1_HVT U795 ( .A1(\ram[0][37] ), .A3(\ram[2][37] ), .A2(\ram[1][37] ), 
        .A4(\ram[3][37] ), .S0(n474), .S1(n381), .Y(n756) );
  MUX41X1_HVT U796 ( .A1(n756), .A3(n754), .A2(n755), .A4(n753), .S0(n583), 
        .S1(n570), .Y(q[37]) );
  MUX41X1_HVT U797 ( .A1(\ram[12][38] ), .A3(\ram[14][38] ), .A2(\ram[13][38] ), .A4(\ram[15][38] ), .S0(n474), .S1(n381), .Y(n757) );
  MUX41X1_HVT U798 ( .A1(\ram[8][38] ), .A3(\ram[10][38] ), .A2(\ram[9][38] ), 
        .A4(\ram[11][38] ), .S0(n474), .S1(n381), .Y(n758) );
  MUX41X1_HVT U799 ( .A1(\ram[4][38] ), .A3(\ram[6][38] ), .A2(\ram[5][38] ), 
        .A4(\ram[7][38] ), .S0(n474), .S1(n381), .Y(n759) );
  MUX41X1_HVT U800 ( .A1(\ram[0][38] ), .A3(\ram[2][38] ), .A2(\ram[1][38] ), 
        .A4(\ram[3][38] ), .S0(n474), .S1(n381), .Y(n760) );
  MUX41X1_HVT U801 ( .A1(n760), .A3(n758), .A2(n759), .A4(n757), .S0(n583), 
        .S1(n570), .Y(q[38]) );
  MUX41X1_HVT U802 ( .A1(\ram[12][39] ), .A3(\ram[14][39] ), .A2(\ram[13][39] ), .A4(\ram[15][39] ), .S0(n475), .S1(n382), .Y(n761) );
  MUX41X1_HVT U803 ( .A1(\ram[8][39] ), .A3(\ram[10][39] ), .A2(\ram[9][39] ), 
        .A4(\ram[11][39] ), .S0(n475), .S1(n382), .Y(n762) );
  MUX41X1_HVT U804 ( .A1(\ram[4][39] ), .A3(\ram[6][39] ), .A2(\ram[5][39] ), 
        .A4(\ram[7][39] ), .S0(n475), .S1(n382), .Y(n763) );
  MUX41X1_HVT U805 ( .A1(\ram[0][39] ), .A3(\ram[2][39] ), .A2(\ram[1][39] ), 
        .A4(\ram[3][39] ), .S0(n475), .S1(n382), .Y(n764) );
  MUX41X1_HVT U806 ( .A1(n764), .A3(n762), .A2(n763), .A4(n761), .S0(n583), 
        .S1(n570), .Y(q[39]) );
  MUX41X1_HVT U807 ( .A1(\ram[12][40] ), .A3(\ram[14][40] ), .A2(\ram[13][40] ), .A4(\ram[15][40] ), .S0(n475), .S1(n382), .Y(n765) );
  MUX41X1_HVT U808 ( .A1(\ram[8][40] ), .A3(\ram[10][40] ), .A2(\ram[9][40] ), 
        .A4(\ram[11][40] ), .S0(n475), .S1(n382), .Y(n766) );
  MUX41X1_HVT U809 ( .A1(\ram[4][40] ), .A3(\ram[6][40] ), .A2(\ram[5][40] ), 
        .A4(\ram[7][40] ), .S0(n475), .S1(n382), .Y(n767) );
  MUX41X1_HVT U810 ( .A1(\ram[0][40] ), .A3(\ram[2][40] ), .A2(\ram[1][40] ), 
        .A4(\ram[3][40] ), .S0(n475), .S1(n382), .Y(n768) );
  MUX41X1_HVT U811 ( .A1(n768), .A3(n766), .A2(n767), .A4(n765), .S0(n583), 
        .S1(n570), .Y(q[40]) );
  MUX41X1_HVT U812 ( .A1(\ram[12][41] ), .A3(\ram[14][41] ), .A2(\ram[13][41] ), .A4(\ram[15][41] ), .S0(n475), .S1(n382), .Y(n769) );
  MUX41X1_HVT U813 ( .A1(\ram[8][41] ), .A3(\ram[10][41] ), .A2(\ram[9][41] ), 
        .A4(\ram[11][41] ), .S0(n475), .S1(n382), .Y(n770) );
  MUX41X1_HVT U814 ( .A1(\ram[4][41] ), .A3(\ram[6][41] ), .A2(\ram[5][41] ), 
        .A4(\ram[7][41] ), .S0(n475), .S1(n382), .Y(n771) );
  MUX41X1_HVT U815 ( .A1(\ram[0][41] ), .A3(\ram[2][41] ), .A2(\ram[1][41] ), 
        .A4(\ram[3][41] ), .S0(n475), .S1(n382), .Y(n772) );
  MUX41X1_HVT U816 ( .A1(n772), .A3(n770), .A2(n771), .A4(n769), .S0(n583), 
        .S1(n571), .Y(q[41]) );
  MUX41X1_HVT U817 ( .A1(\ram[12][42] ), .A3(\ram[14][42] ), .A2(\ram[13][42] ), .A4(\ram[15][42] ), .S0(n476), .S1(n383), .Y(n773) );
  MUX41X1_HVT U818 ( .A1(\ram[8][42] ), .A3(\ram[10][42] ), .A2(\ram[9][42] ), 
        .A4(\ram[11][42] ), .S0(n476), .S1(n383), .Y(n774) );
  MUX41X1_HVT U819 ( .A1(\ram[4][42] ), .A3(\ram[6][42] ), .A2(\ram[5][42] ), 
        .A4(\ram[7][42] ), .S0(n476), .S1(n383), .Y(n775) );
  MUX41X1_HVT U820 ( .A1(\ram[0][42] ), .A3(\ram[2][42] ), .A2(\ram[1][42] ), 
        .A4(\ram[3][42] ), .S0(n476), .S1(n383), .Y(n776) );
  MUX41X1_HVT U821 ( .A1(n776), .A3(n774), .A2(n775), .A4(n773), .S0(n583), 
        .S1(n571), .Y(q[42]) );
  MUX41X1_HVT U822 ( .A1(\ram[12][43] ), .A3(\ram[14][43] ), .A2(\ram[13][43] ), .A4(\ram[15][43] ), .S0(n476), .S1(n383), .Y(n777) );
  MUX41X1_HVT U823 ( .A1(\ram[8][43] ), .A3(\ram[10][43] ), .A2(\ram[9][43] ), 
        .A4(\ram[11][43] ), .S0(n476), .S1(n383), .Y(n778) );
  MUX41X1_HVT U824 ( .A1(\ram[4][43] ), .A3(\ram[6][43] ), .A2(\ram[5][43] ), 
        .A4(\ram[7][43] ), .S0(n476), .S1(n383), .Y(n779) );
  MUX41X1_HVT U825 ( .A1(\ram[0][43] ), .A3(\ram[2][43] ), .A2(\ram[1][43] ), 
        .A4(\ram[3][43] ), .S0(n476), .S1(n383), .Y(n780) );
  MUX41X1_HVT U826 ( .A1(n780), .A3(n778), .A2(n779), .A4(n777), .S0(n583), 
        .S1(n571), .Y(q[43]) );
  MUX41X1_HVT U827 ( .A1(\ram[12][44] ), .A3(\ram[14][44] ), .A2(\ram[13][44] ), .A4(\ram[15][44] ), .S0(n476), .S1(n383), .Y(n781) );
  MUX41X1_HVT U828 ( .A1(\ram[8][44] ), .A3(\ram[10][44] ), .A2(\ram[9][44] ), 
        .A4(\ram[11][44] ), .S0(n476), .S1(n383), .Y(n782) );
  MUX41X1_HVT U829 ( .A1(\ram[4][44] ), .A3(\ram[6][44] ), .A2(\ram[5][44] ), 
        .A4(\ram[7][44] ), .S0(n476), .S1(n383), .Y(n783) );
  MUX41X1_HVT U830 ( .A1(\ram[0][44] ), .A3(\ram[2][44] ), .A2(\ram[1][44] ), 
        .A4(\ram[3][44] ), .S0(n476), .S1(n383), .Y(n784) );
  MUX41X1_HVT U831 ( .A1(n784), .A3(n782), .A2(n783), .A4(n781), .S0(n583), 
        .S1(n571), .Y(q[44]) );
  MUX41X1_HVT U832 ( .A1(\ram[12][45] ), .A3(\ram[14][45] ), .A2(\ram[13][45] ), .A4(\ram[15][45] ), .S0(n477), .S1(n384), .Y(n785) );
  MUX41X1_HVT U833 ( .A1(\ram[8][45] ), .A3(\ram[10][45] ), .A2(\ram[9][45] ), 
        .A4(\ram[11][45] ), .S0(n477), .S1(n384), .Y(n786) );
  MUX41X1_HVT U834 ( .A1(\ram[4][45] ), .A3(\ram[6][45] ), .A2(\ram[5][45] ), 
        .A4(\ram[7][45] ), .S0(n477), .S1(n384), .Y(n787) );
  MUX41X1_HVT U835 ( .A1(\ram[0][45] ), .A3(\ram[2][45] ), .A2(\ram[1][45] ), 
        .A4(\ram[3][45] ), .S0(n477), .S1(n384), .Y(n788) );
  MUX41X1_HVT U836 ( .A1(n788), .A3(n786), .A2(n787), .A4(n785), .S0(n583), 
        .S1(n571), .Y(q[45]) );
  MUX41X1_HVT U837 ( .A1(\ram[12][46] ), .A3(\ram[14][46] ), .A2(\ram[13][46] ), .A4(\ram[15][46] ), .S0(n477), .S1(n384), .Y(n789) );
  MUX41X1_HVT U838 ( .A1(\ram[8][46] ), .A3(\ram[10][46] ), .A2(\ram[9][46] ), 
        .A4(\ram[11][46] ), .S0(n477), .S1(n384), .Y(n790) );
  MUX41X1_HVT U839 ( .A1(\ram[4][46] ), .A3(\ram[6][46] ), .A2(\ram[5][46] ), 
        .A4(\ram[7][46] ), .S0(n477), .S1(n384), .Y(n791) );
  MUX41X1_HVT U840 ( .A1(\ram[0][46] ), .A3(\ram[2][46] ), .A2(\ram[1][46] ), 
        .A4(\ram[3][46] ), .S0(n477), .S1(n384), .Y(n792) );
  MUX41X1_HVT U841 ( .A1(n792), .A3(n790), .A2(n791), .A4(n789), .S0(n583), 
        .S1(n571), .Y(q[46]) );
  MUX41X1_HVT U842 ( .A1(\ram[12][47] ), .A3(\ram[14][47] ), .A2(\ram[13][47] ), .A4(\ram[15][47] ), .S0(n477), .S1(n384), .Y(n793) );
  MUX41X1_HVT U843 ( .A1(\ram[8][47] ), .A3(\ram[10][47] ), .A2(\ram[9][47] ), 
        .A4(\ram[11][47] ), .S0(n477), .S1(n384), .Y(n794) );
  MUX41X1_HVT U844 ( .A1(\ram[4][47] ), .A3(\ram[6][47] ), .A2(\ram[5][47] ), 
        .A4(\ram[7][47] ), .S0(n477), .S1(n384), .Y(n795) );
  MUX41X1_HVT U845 ( .A1(\ram[0][47] ), .A3(\ram[2][47] ), .A2(\ram[1][47] ), 
        .A4(\ram[3][47] ), .S0(n477), .S1(n384), .Y(n796) );
  MUX41X1_HVT U846 ( .A1(n796), .A3(n794), .A2(n795), .A4(n793), .S0(n583), 
        .S1(n571), .Y(q[47]) );
  MUX41X1_HVT U847 ( .A1(\ram[12][48] ), .A3(\ram[14][48] ), .A2(\ram[13][48] ), .A4(\ram[15][48] ), .S0(n478), .S1(n385), .Y(n797) );
  MUX41X1_HVT U848 ( .A1(\ram[8][48] ), .A3(\ram[10][48] ), .A2(\ram[9][48] ), 
        .A4(\ram[11][48] ), .S0(n478), .S1(n385), .Y(n798) );
  MUX41X1_HVT U849 ( .A1(\ram[4][48] ), .A3(\ram[6][48] ), .A2(\ram[5][48] ), 
        .A4(\ram[7][48] ), .S0(n478), .S1(n385), .Y(n799) );
  MUX41X1_HVT U850 ( .A1(\ram[0][48] ), .A3(\ram[2][48] ), .A2(\ram[1][48] ), 
        .A4(\ram[3][48] ), .S0(n478), .S1(n385), .Y(n800) );
  MUX41X1_HVT U851 ( .A1(n800), .A3(n798), .A2(n799), .A4(n797), .S0(n584), 
        .S1(n571), .Y(q[48]) );
  MUX41X1_HVT U852 ( .A1(\ram[12][49] ), .A3(\ram[14][49] ), .A2(\ram[13][49] ), .A4(\ram[15][49] ), .S0(n478), .S1(n385), .Y(n801) );
  MUX41X1_HVT U853 ( .A1(\ram[8][49] ), .A3(\ram[10][49] ), .A2(\ram[9][49] ), 
        .A4(\ram[11][49] ), .S0(n478), .S1(n385), .Y(n802) );
  MUX41X1_HVT U854 ( .A1(\ram[4][49] ), .A3(\ram[6][49] ), .A2(\ram[5][49] ), 
        .A4(\ram[7][49] ), .S0(n478), .S1(n385), .Y(n803) );
  MUX41X1_HVT U855 ( .A1(\ram[0][49] ), .A3(\ram[2][49] ), .A2(\ram[1][49] ), 
        .A4(\ram[3][49] ), .S0(n478), .S1(n385), .Y(n804) );
  MUX41X1_HVT U856 ( .A1(n804), .A3(n802), .A2(n803), .A4(n801), .S0(n584), 
        .S1(n571), .Y(q[49]) );
  MUX41X1_HVT U857 ( .A1(\ram[12][50] ), .A3(\ram[14][50] ), .A2(\ram[13][50] ), .A4(\ram[15][50] ), .S0(n478), .S1(n385), .Y(n805) );
  MUX41X1_HVT U858 ( .A1(\ram[8][50] ), .A3(\ram[10][50] ), .A2(\ram[9][50] ), 
        .A4(\ram[11][50] ), .S0(n478), .S1(n385), .Y(n806) );
  MUX41X1_HVT U859 ( .A1(\ram[4][50] ), .A3(\ram[6][50] ), .A2(\ram[5][50] ), 
        .A4(\ram[7][50] ), .S0(n478), .S1(n385), .Y(n807) );
  MUX41X1_HVT U860 ( .A1(\ram[0][50] ), .A3(\ram[2][50] ), .A2(\ram[1][50] ), 
        .A4(\ram[3][50] ), .S0(n478), .S1(n385), .Y(n808) );
  MUX41X1_HVT U861 ( .A1(n808), .A3(n806), .A2(n807), .A4(n805), .S0(n584), 
        .S1(n571), .Y(q[50]) );
  MUX41X1_HVT U862 ( .A1(\ram[12][51] ), .A3(\ram[14][51] ), .A2(\ram[13][51] ), .A4(\ram[15][51] ), .S0(n479), .S1(n386), .Y(n809) );
  MUX41X1_HVT U863 ( .A1(\ram[8][51] ), .A3(\ram[10][51] ), .A2(\ram[9][51] ), 
        .A4(\ram[11][51] ), .S0(n479), .S1(n386), .Y(n810) );
  MUX41X1_HVT U864 ( .A1(\ram[4][51] ), .A3(\ram[6][51] ), .A2(\ram[5][51] ), 
        .A4(\ram[7][51] ), .S0(n479), .S1(n386), .Y(n811) );
  MUX41X1_HVT U865 ( .A1(\ram[0][51] ), .A3(\ram[2][51] ), .A2(\ram[1][51] ), 
        .A4(\ram[3][51] ), .S0(n479), .S1(n386), .Y(n812) );
  MUX41X1_HVT U866 ( .A1(n812), .A3(n810), .A2(n811), .A4(n809), .S0(n584), 
        .S1(n571), .Y(q[51]) );
  MUX41X1_HVT U867 ( .A1(\ram[12][52] ), .A3(\ram[14][52] ), .A2(\ram[13][52] ), .A4(\ram[15][52] ), .S0(n479), .S1(n386), .Y(n813) );
  MUX41X1_HVT U868 ( .A1(\ram[8][52] ), .A3(\ram[10][52] ), .A2(\ram[9][52] ), 
        .A4(\ram[11][52] ), .S0(n479), .S1(n386), .Y(n814) );
  MUX41X1_HVT U869 ( .A1(\ram[4][52] ), .A3(\ram[6][52] ), .A2(\ram[5][52] ), 
        .A4(\ram[7][52] ), .S0(n479), .S1(n386), .Y(n815) );
  MUX41X1_HVT U870 ( .A1(\ram[0][52] ), .A3(\ram[2][52] ), .A2(\ram[1][52] ), 
        .A4(\ram[3][52] ), .S0(n479), .S1(n386), .Y(n816) );
  MUX41X1_HVT U871 ( .A1(n816), .A3(n814), .A2(n815), .A4(n813), .S0(n584), 
        .S1(n571), .Y(q[52]) );
  MUX41X1_HVT U872 ( .A1(\ram[12][53] ), .A3(\ram[14][53] ), .A2(\ram[13][53] ), .A4(\ram[15][53] ), .S0(n479), .S1(n386), .Y(n817) );
  MUX41X1_HVT U873 ( .A1(\ram[8][53] ), .A3(\ram[10][53] ), .A2(\ram[9][53] ), 
        .A4(\ram[11][53] ), .S0(n479), .S1(n386), .Y(n818) );
  MUX41X1_HVT U874 ( .A1(\ram[4][53] ), .A3(\ram[6][53] ), .A2(\ram[5][53] ), 
        .A4(\ram[7][53] ), .S0(n479), .S1(n386), .Y(n819) );
  MUX41X1_HVT U875 ( .A1(\ram[0][53] ), .A3(\ram[2][53] ), .A2(\ram[1][53] ), 
        .A4(\ram[3][53] ), .S0(n479), .S1(n386), .Y(n820) );
  MUX41X1_HVT U876 ( .A1(n820), .A3(n818), .A2(n819), .A4(n817), .S0(n584), 
        .S1(n572), .Y(q[53]) );
  MUX41X1_HVT U877 ( .A1(\ram[12][54] ), .A3(\ram[14][54] ), .A2(\ram[13][54] ), .A4(\ram[15][54] ), .S0(n480), .S1(n387), .Y(n821) );
  MUX41X1_HVT U878 ( .A1(\ram[8][54] ), .A3(\ram[10][54] ), .A2(\ram[9][54] ), 
        .A4(\ram[11][54] ), .S0(n480), .S1(n387), .Y(n822) );
  MUX41X1_HVT U879 ( .A1(\ram[4][54] ), .A3(\ram[6][54] ), .A2(\ram[5][54] ), 
        .A4(\ram[7][54] ), .S0(n480), .S1(n387), .Y(n823) );
  MUX41X1_HVT U880 ( .A1(\ram[0][54] ), .A3(\ram[2][54] ), .A2(\ram[1][54] ), 
        .A4(\ram[3][54] ), .S0(n480), .S1(n387), .Y(n824) );
  MUX41X1_HVT U881 ( .A1(n824), .A3(n822), .A2(n823), .A4(n821), .S0(n584), 
        .S1(n572), .Y(q[54]) );
  MUX41X1_HVT U882 ( .A1(\ram[12][55] ), .A3(\ram[14][55] ), .A2(\ram[13][55] ), .A4(\ram[15][55] ), .S0(n480), .S1(n387), .Y(n825) );
  MUX41X1_HVT U883 ( .A1(\ram[8][55] ), .A3(\ram[10][55] ), .A2(\ram[9][55] ), 
        .A4(\ram[11][55] ), .S0(n480), .S1(n387), .Y(n826) );
  MUX41X1_HVT U884 ( .A1(\ram[4][55] ), .A3(\ram[6][55] ), .A2(\ram[5][55] ), 
        .A4(\ram[7][55] ), .S0(n480), .S1(n387), .Y(n827) );
  MUX41X1_HVT U885 ( .A1(\ram[0][55] ), .A3(\ram[2][55] ), .A2(\ram[1][55] ), 
        .A4(\ram[3][55] ), .S0(n480), .S1(n387), .Y(n828) );
  MUX41X1_HVT U886 ( .A1(n828), .A3(n826), .A2(n827), .A4(n825), .S0(n584), 
        .S1(n572), .Y(q[55]) );
  MUX41X1_HVT U887 ( .A1(\ram[12][56] ), .A3(\ram[14][56] ), .A2(\ram[13][56] ), .A4(\ram[15][56] ), .S0(n480), .S1(n387), .Y(n829) );
  MUX41X1_HVT U888 ( .A1(\ram[8][56] ), .A3(\ram[10][56] ), .A2(\ram[9][56] ), 
        .A4(\ram[11][56] ), .S0(n480), .S1(n387), .Y(n830) );
  MUX41X1_HVT U889 ( .A1(\ram[4][56] ), .A3(\ram[6][56] ), .A2(\ram[5][56] ), 
        .A4(\ram[7][56] ), .S0(n480), .S1(n387), .Y(n831) );
  MUX41X1_HVT U890 ( .A1(\ram[0][56] ), .A3(\ram[2][56] ), .A2(\ram[1][56] ), 
        .A4(\ram[3][56] ), .S0(n480), .S1(n387), .Y(n832) );
  MUX41X1_HVT U891 ( .A1(n832), .A3(n830), .A2(n831), .A4(n829), .S0(n584), 
        .S1(n572), .Y(q[56]) );
  MUX41X1_HVT U892 ( .A1(\ram[12][57] ), .A3(\ram[14][57] ), .A2(\ram[13][57] ), .A4(\ram[15][57] ), .S0(n481), .S1(n388), .Y(n833) );
  MUX41X1_HVT U893 ( .A1(\ram[8][57] ), .A3(\ram[10][57] ), .A2(\ram[9][57] ), 
        .A4(\ram[11][57] ), .S0(n481), .S1(n388), .Y(n834) );
  MUX41X1_HVT U894 ( .A1(\ram[4][57] ), .A3(\ram[6][57] ), .A2(\ram[5][57] ), 
        .A4(\ram[7][57] ), .S0(n481), .S1(n388), .Y(n835) );
  MUX41X1_HVT U895 ( .A1(\ram[0][57] ), .A3(\ram[2][57] ), .A2(\ram[1][57] ), 
        .A4(\ram[3][57] ), .S0(n481), .S1(n388), .Y(n836) );
  MUX41X1_HVT U896 ( .A1(n836), .A3(n834), .A2(n835), .A4(n833), .S0(n584), 
        .S1(n572), .Y(q[57]) );
  MUX41X1_HVT U897 ( .A1(\ram[12][58] ), .A3(\ram[14][58] ), .A2(\ram[13][58] ), .A4(\ram[15][58] ), .S0(n481), .S1(n388), .Y(n837) );
  MUX41X1_HVT U898 ( .A1(\ram[8][58] ), .A3(\ram[10][58] ), .A2(\ram[9][58] ), 
        .A4(\ram[11][58] ), .S0(n481), .S1(n388), .Y(n838) );
  MUX41X1_HVT U899 ( .A1(\ram[4][58] ), .A3(\ram[6][58] ), .A2(\ram[5][58] ), 
        .A4(\ram[7][58] ), .S0(n481), .S1(n388), .Y(n839) );
  MUX41X1_HVT U900 ( .A1(\ram[0][58] ), .A3(\ram[2][58] ), .A2(\ram[1][58] ), 
        .A4(\ram[3][58] ), .S0(n481), .S1(n388), .Y(n840) );
  MUX41X1_HVT U901 ( .A1(n840), .A3(n838), .A2(n839), .A4(n837), .S0(n584), 
        .S1(n572), .Y(q[58]) );
  MUX41X1_HVT U902 ( .A1(\ram[12][59] ), .A3(\ram[14][59] ), .A2(\ram[13][59] ), .A4(\ram[15][59] ), .S0(n481), .S1(n388), .Y(n841) );
  MUX41X1_HVT U903 ( .A1(\ram[8][59] ), .A3(\ram[10][59] ), .A2(\ram[9][59] ), 
        .A4(\ram[11][59] ), .S0(n481), .S1(n388), .Y(n842) );
  MUX41X1_HVT U904 ( .A1(\ram[4][59] ), .A3(\ram[6][59] ), .A2(\ram[5][59] ), 
        .A4(\ram[7][59] ), .S0(n481), .S1(n388), .Y(n843) );
  MUX41X1_HVT U905 ( .A1(\ram[0][59] ), .A3(\ram[2][59] ), .A2(\ram[1][59] ), 
        .A4(\ram[3][59] ), .S0(n481), .S1(n388), .Y(n844) );
  MUX41X1_HVT U906 ( .A1(n844), .A3(n842), .A2(n843), .A4(n841), .S0(n584), 
        .S1(n572), .Y(q[59]) );
  MUX41X1_HVT U907 ( .A1(\ram[12][60] ), .A3(\ram[14][60] ), .A2(\ram[13][60] ), .A4(\ram[15][60] ), .S0(n482), .S1(n389), .Y(n845) );
  MUX41X1_HVT U908 ( .A1(\ram[8][60] ), .A3(\ram[10][60] ), .A2(\ram[9][60] ), 
        .A4(\ram[11][60] ), .S0(n482), .S1(n389), .Y(n846) );
  MUX41X1_HVT U909 ( .A1(\ram[4][60] ), .A3(\ram[6][60] ), .A2(\ram[5][60] ), 
        .A4(\ram[7][60] ), .S0(n482), .S1(n389), .Y(n847) );
  MUX41X1_HVT U910 ( .A1(\ram[0][60] ), .A3(\ram[2][60] ), .A2(\ram[1][60] ), 
        .A4(\ram[3][60] ), .S0(n482), .S1(n389), .Y(n848) );
  MUX41X1_HVT U911 ( .A1(n848), .A3(n846), .A2(n847), .A4(n845), .S0(n585), 
        .S1(n572), .Y(q[60]) );
  MUX41X1_HVT U912 ( .A1(\ram[12][61] ), .A3(\ram[14][61] ), .A2(\ram[13][61] ), .A4(\ram[15][61] ), .S0(n482), .S1(n389), .Y(n849) );
  MUX41X1_HVT U913 ( .A1(\ram[8][61] ), .A3(\ram[10][61] ), .A2(\ram[9][61] ), 
        .A4(\ram[11][61] ), .S0(n482), .S1(n389), .Y(n850) );
  MUX41X1_HVT U914 ( .A1(\ram[4][61] ), .A3(\ram[6][61] ), .A2(\ram[5][61] ), 
        .A4(\ram[7][61] ), .S0(n482), .S1(n389), .Y(n851) );
  MUX41X1_HVT U915 ( .A1(\ram[0][61] ), .A3(\ram[2][61] ), .A2(\ram[1][61] ), 
        .A4(\ram[3][61] ), .S0(n482), .S1(n389), .Y(n852) );
  MUX41X1_HVT U916 ( .A1(n852), .A3(n850), .A2(n851), .A4(n849), .S0(n585), 
        .S1(n572), .Y(q[61]) );
  MUX41X1_HVT U917 ( .A1(\ram[12][62] ), .A3(\ram[14][62] ), .A2(\ram[13][62] ), .A4(\ram[15][62] ), .S0(n482), .S1(n389), .Y(n853) );
  MUX41X1_HVT U918 ( .A1(\ram[8][62] ), .A3(\ram[10][62] ), .A2(\ram[9][62] ), 
        .A4(\ram[11][62] ), .S0(n482), .S1(n389), .Y(n854) );
  MUX41X1_HVT U919 ( .A1(\ram[4][62] ), .A3(\ram[6][62] ), .A2(\ram[5][62] ), 
        .A4(\ram[7][62] ), .S0(n482), .S1(n389), .Y(n855) );
  MUX41X1_HVT U920 ( .A1(\ram[0][62] ), .A3(\ram[2][62] ), .A2(\ram[1][62] ), 
        .A4(\ram[3][62] ), .S0(n482), .S1(n389), .Y(n856) );
  MUX41X1_HVT U921 ( .A1(n856), .A3(n854), .A2(n855), .A4(n853), .S0(n585), 
        .S1(n572), .Y(q[62]) );
  MUX41X1_HVT U922 ( .A1(\ram[12][63] ), .A3(\ram[14][63] ), .A2(\ram[13][63] ), .A4(\ram[15][63] ), .S0(n483), .S1(n390), .Y(n857) );
  MUX41X1_HVT U923 ( .A1(\ram[8][63] ), .A3(\ram[10][63] ), .A2(\ram[9][63] ), 
        .A4(\ram[11][63] ), .S0(n483), .S1(n390), .Y(n858) );
  MUX41X1_HVT U924 ( .A1(\ram[4][63] ), .A3(\ram[6][63] ), .A2(\ram[5][63] ), 
        .A4(\ram[7][63] ), .S0(n483), .S1(n390), .Y(n859) );
  MUX41X1_HVT U925 ( .A1(\ram[0][63] ), .A3(\ram[2][63] ), .A2(\ram[1][63] ), 
        .A4(\ram[3][63] ), .S0(n483), .S1(n390), .Y(n860) );
  MUX41X1_HVT U926 ( .A1(n860), .A3(n858), .A2(n859), .A4(n857), .S0(n585), 
        .S1(n572), .Y(q[63]) );
  MUX41X1_HVT U927 ( .A1(\ram[12][64] ), .A3(\ram[14][64] ), .A2(\ram[13][64] ), .A4(\ram[15][64] ), .S0(n483), .S1(n390), .Y(n861) );
  MUX41X1_HVT U928 ( .A1(\ram[8][64] ), .A3(\ram[10][64] ), .A2(\ram[9][64] ), 
        .A4(\ram[11][64] ), .S0(n483), .S1(n390), .Y(n862) );
  MUX41X1_HVT U929 ( .A1(\ram[4][64] ), .A3(\ram[6][64] ), .A2(\ram[5][64] ), 
        .A4(\ram[7][64] ), .S0(n483), .S1(n390), .Y(n863) );
  MUX41X1_HVT U930 ( .A1(\ram[0][64] ), .A3(\ram[2][64] ), .A2(\ram[1][64] ), 
        .A4(\ram[3][64] ), .S0(n483), .S1(n390), .Y(n864) );
  MUX41X1_HVT U931 ( .A1(n864), .A3(n862), .A2(n863), .A4(n861), .S0(n585), 
        .S1(n572), .Y(q[64]) );
  MUX41X1_HVT U932 ( .A1(\ram[12][65] ), .A3(\ram[14][65] ), .A2(\ram[13][65] ), .A4(\ram[15][65] ), .S0(n483), .S1(n390), .Y(n865) );
  MUX41X1_HVT U933 ( .A1(\ram[8][65] ), .A3(\ram[10][65] ), .A2(\ram[9][65] ), 
        .A4(\ram[11][65] ), .S0(n483), .S1(n390), .Y(n866) );
  MUX41X1_HVT U934 ( .A1(\ram[4][65] ), .A3(\ram[6][65] ), .A2(\ram[5][65] ), 
        .A4(\ram[7][65] ), .S0(n483), .S1(n390), .Y(n867) );
  MUX41X1_HVT U935 ( .A1(\ram[0][65] ), .A3(\ram[2][65] ), .A2(\ram[1][65] ), 
        .A4(\ram[3][65] ), .S0(n483), .S1(n390), .Y(n868) );
  MUX41X1_HVT U936 ( .A1(n868), .A3(n866), .A2(n867), .A4(n865), .S0(n585), 
        .S1(n573), .Y(q[65]) );
  MUX41X1_HVT U937 ( .A1(\ram[12][66] ), .A3(\ram[14][66] ), .A2(\ram[13][66] ), .A4(\ram[15][66] ), .S0(n484), .S1(n391), .Y(n869) );
  MUX41X1_HVT U938 ( .A1(\ram[8][66] ), .A3(\ram[10][66] ), .A2(\ram[9][66] ), 
        .A4(\ram[11][66] ), .S0(n484), .S1(n391), .Y(n870) );
  MUX41X1_HVT U939 ( .A1(\ram[4][66] ), .A3(\ram[6][66] ), .A2(\ram[5][66] ), 
        .A4(\ram[7][66] ), .S0(n484), .S1(n391), .Y(n871) );
  MUX41X1_HVT U940 ( .A1(\ram[0][66] ), .A3(\ram[2][66] ), .A2(\ram[1][66] ), 
        .A4(\ram[3][66] ), .S0(n484), .S1(n391), .Y(n872) );
  MUX41X1_HVT U941 ( .A1(n872), .A3(n870), .A2(n871), .A4(n869), .S0(n585), 
        .S1(n573), .Y(q[66]) );
  MUX41X1_HVT U942 ( .A1(\ram[12][67] ), .A3(\ram[14][67] ), .A2(\ram[13][67] ), .A4(\ram[15][67] ), .S0(n484), .S1(n391), .Y(n873) );
  MUX41X1_HVT U943 ( .A1(\ram[8][67] ), .A3(\ram[10][67] ), .A2(\ram[9][67] ), 
        .A4(\ram[11][67] ), .S0(n484), .S1(n391), .Y(n874) );
  MUX41X1_HVT U944 ( .A1(\ram[4][67] ), .A3(\ram[6][67] ), .A2(\ram[5][67] ), 
        .A4(\ram[7][67] ), .S0(n484), .S1(n391), .Y(n875) );
  MUX41X1_HVT U945 ( .A1(\ram[0][67] ), .A3(\ram[2][67] ), .A2(\ram[1][67] ), 
        .A4(\ram[3][67] ), .S0(n484), .S1(n391), .Y(n876) );
  MUX41X1_HVT U946 ( .A1(n876), .A3(n874), .A2(n875), .A4(n873), .S0(n585), 
        .S1(n573), .Y(q[67]) );
  MUX41X1_HVT U947 ( .A1(\ram[12][68] ), .A3(\ram[14][68] ), .A2(\ram[13][68] ), .A4(\ram[15][68] ), .S0(n484), .S1(n391), .Y(n877) );
  MUX41X1_HVT U948 ( .A1(\ram[8][68] ), .A3(\ram[10][68] ), .A2(\ram[9][68] ), 
        .A4(\ram[11][68] ), .S0(n484), .S1(n391), .Y(n878) );
  MUX41X1_HVT U949 ( .A1(\ram[4][68] ), .A3(\ram[6][68] ), .A2(\ram[5][68] ), 
        .A4(\ram[7][68] ), .S0(n484), .S1(n391), .Y(n879) );
  MUX41X1_HVT U950 ( .A1(\ram[0][68] ), .A3(\ram[2][68] ), .A2(\ram[1][68] ), 
        .A4(\ram[3][68] ), .S0(n484), .S1(n391), .Y(n880) );
  MUX41X1_HVT U951 ( .A1(n880), .A3(n878), .A2(n879), .A4(n877), .S0(n585), 
        .S1(n573), .Y(q[68]) );
  MUX41X1_HVT U952 ( .A1(\ram[12][69] ), .A3(\ram[14][69] ), .A2(\ram[13][69] ), .A4(\ram[15][69] ), .S0(n485), .S1(n392), .Y(n881) );
  MUX41X1_HVT U953 ( .A1(\ram[8][69] ), .A3(\ram[10][69] ), .A2(\ram[9][69] ), 
        .A4(\ram[11][69] ), .S0(n485), .S1(n392), .Y(n882) );
  MUX41X1_HVT U954 ( .A1(\ram[4][69] ), .A3(\ram[6][69] ), .A2(\ram[5][69] ), 
        .A4(\ram[7][69] ), .S0(n485), .S1(n392), .Y(n883) );
  MUX41X1_HVT U955 ( .A1(\ram[0][69] ), .A3(\ram[2][69] ), .A2(\ram[1][69] ), 
        .A4(\ram[3][69] ), .S0(n485), .S1(n392), .Y(n884) );
  MUX41X1_HVT U956 ( .A1(n884), .A3(n882), .A2(n883), .A4(n881), .S0(n585), 
        .S1(n573), .Y(q[69]) );
  MUX41X1_HVT U957 ( .A1(\ram[12][70] ), .A3(\ram[14][70] ), .A2(\ram[13][70] ), .A4(\ram[15][70] ), .S0(n485), .S1(n392), .Y(n885) );
  MUX41X1_HVT U958 ( .A1(\ram[8][70] ), .A3(\ram[10][70] ), .A2(\ram[9][70] ), 
        .A4(\ram[11][70] ), .S0(n485), .S1(n392), .Y(n886) );
  MUX41X1_HVT U959 ( .A1(\ram[4][70] ), .A3(\ram[6][70] ), .A2(\ram[5][70] ), 
        .A4(\ram[7][70] ), .S0(n485), .S1(n392), .Y(n887) );
  MUX41X1_HVT U960 ( .A1(\ram[0][70] ), .A3(\ram[2][70] ), .A2(\ram[1][70] ), 
        .A4(\ram[3][70] ), .S0(n485), .S1(n392), .Y(n888) );
  MUX41X1_HVT U961 ( .A1(n888), .A3(n886), .A2(n887), .A4(n885), .S0(n585), 
        .S1(n573), .Y(q[70]) );
  MUX41X1_HVT U962 ( .A1(\ram[12][71] ), .A3(\ram[14][71] ), .A2(\ram[13][71] ), .A4(\ram[15][71] ), .S0(n485), .S1(n392), .Y(n889) );
  MUX41X1_HVT U963 ( .A1(\ram[8][71] ), .A3(\ram[10][71] ), .A2(\ram[9][71] ), 
        .A4(\ram[11][71] ), .S0(n485), .S1(n392), .Y(n890) );
  MUX41X1_HVT U964 ( .A1(\ram[4][71] ), .A3(\ram[6][71] ), .A2(\ram[5][71] ), 
        .A4(\ram[7][71] ), .S0(n485), .S1(n392), .Y(n891) );
  MUX41X1_HVT U965 ( .A1(\ram[0][71] ), .A3(\ram[2][71] ), .A2(\ram[1][71] ), 
        .A4(\ram[3][71] ), .S0(n485), .S1(n392), .Y(n892) );
  MUX41X1_HVT U966 ( .A1(n892), .A3(n890), .A2(n891), .A4(n889), .S0(n585), 
        .S1(n573), .Y(q[71]) );
  MUX41X1_HVT U967 ( .A1(\ram[12][72] ), .A3(\ram[14][72] ), .A2(\ram[13][72] ), .A4(\ram[15][72] ), .S0(n486), .S1(n393), .Y(n893) );
  MUX41X1_HVT U968 ( .A1(\ram[8][72] ), .A3(\ram[10][72] ), .A2(\ram[9][72] ), 
        .A4(\ram[11][72] ), .S0(n486), .S1(n393), .Y(n894) );
  MUX41X1_HVT U969 ( .A1(\ram[4][72] ), .A3(\ram[6][72] ), .A2(\ram[5][72] ), 
        .A4(\ram[7][72] ), .S0(n486), .S1(n393), .Y(n895) );
  MUX41X1_HVT U970 ( .A1(\ram[0][72] ), .A3(\ram[2][72] ), .A2(\ram[1][72] ), 
        .A4(\ram[3][72] ), .S0(n486), .S1(n393), .Y(n896) );
  MUX41X1_HVT U971 ( .A1(n896), .A3(n894), .A2(n895), .A4(n893), .S0(n586), 
        .S1(n573), .Y(q[72]) );
  MUX41X1_HVT U972 ( .A1(\ram[12][73] ), .A3(\ram[14][73] ), .A2(\ram[13][73] ), .A4(\ram[15][73] ), .S0(n486), .S1(n393), .Y(n897) );
  MUX41X1_HVT U973 ( .A1(\ram[8][73] ), .A3(\ram[10][73] ), .A2(\ram[9][73] ), 
        .A4(\ram[11][73] ), .S0(n486), .S1(n393), .Y(n898) );
  MUX41X1_HVT U974 ( .A1(\ram[4][73] ), .A3(\ram[6][73] ), .A2(\ram[5][73] ), 
        .A4(\ram[7][73] ), .S0(n486), .S1(n393), .Y(n899) );
  MUX41X1_HVT U975 ( .A1(\ram[0][73] ), .A3(\ram[2][73] ), .A2(\ram[1][73] ), 
        .A4(\ram[3][73] ), .S0(n486), .S1(n393), .Y(n900) );
  MUX41X1_HVT U976 ( .A1(n900), .A3(n898), .A2(n899), .A4(n897), .S0(n586), 
        .S1(n573), .Y(q[73]) );
  MUX41X1_HVT U977 ( .A1(\ram[12][74] ), .A3(\ram[14][74] ), .A2(\ram[13][74] ), .A4(\ram[15][74] ), .S0(n486), .S1(n393), .Y(n901) );
  MUX41X1_HVT U978 ( .A1(\ram[8][74] ), .A3(\ram[10][74] ), .A2(\ram[9][74] ), 
        .A4(\ram[11][74] ), .S0(n486), .S1(n393), .Y(n902) );
  MUX41X1_HVT U979 ( .A1(\ram[4][74] ), .A3(\ram[6][74] ), .A2(\ram[5][74] ), 
        .A4(\ram[7][74] ), .S0(n486), .S1(n393), .Y(n903) );
  MUX41X1_HVT U980 ( .A1(\ram[0][74] ), .A3(\ram[2][74] ), .A2(\ram[1][74] ), 
        .A4(\ram[3][74] ), .S0(n486), .S1(n393), .Y(n904) );
  MUX41X1_HVT U981 ( .A1(n904), .A3(n902), .A2(n903), .A4(n901), .S0(n586), 
        .S1(n573), .Y(q[74]) );
  MUX41X1_HVT U982 ( .A1(\ram[12][75] ), .A3(\ram[14][75] ), .A2(\ram[13][75] ), .A4(\ram[15][75] ), .S0(n487), .S1(n394), .Y(n905) );
  MUX41X1_HVT U983 ( .A1(\ram[8][75] ), .A3(\ram[10][75] ), .A2(\ram[9][75] ), 
        .A4(\ram[11][75] ), .S0(n487), .S1(n394), .Y(n906) );
  MUX41X1_HVT U984 ( .A1(\ram[4][75] ), .A3(\ram[6][75] ), .A2(\ram[5][75] ), 
        .A4(\ram[7][75] ), .S0(n487), .S1(n394), .Y(n907) );
  MUX41X1_HVT U985 ( .A1(\ram[0][75] ), .A3(\ram[2][75] ), .A2(\ram[1][75] ), 
        .A4(\ram[3][75] ), .S0(n487), .S1(n394), .Y(n908) );
  MUX41X1_HVT U986 ( .A1(n908), .A3(n906), .A2(n907), .A4(n905), .S0(n586), 
        .S1(n574), .Y(q[75]) );
  MUX41X1_HVT U987 ( .A1(\ram[12][76] ), .A3(\ram[14][76] ), .A2(\ram[13][76] ), .A4(\ram[15][76] ), .S0(n487), .S1(n394), .Y(n909) );
  MUX41X1_HVT U988 ( .A1(\ram[8][76] ), .A3(\ram[10][76] ), .A2(\ram[9][76] ), 
        .A4(\ram[11][76] ), .S0(n487), .S1(n394), .Y(n910) );
  MUX41X1_HVT U989 ( .A1(\ram[4][76] ), .A3(\ram[6][76] ), .A2(\ram[5][76] ), 
        .A4(\ram[7][76] ), .S0(n487), .S1(n394), .Y(n911) );
  MUX41X1_HVT U990 ( .A1(\ram[0][76] ), .A3(\ram[2][76] ), .A2(\ram[1][76] ), 
        .A4(\ram[3][76] ), .S0(n487), .S1(n394), .Y(n912) );
  MUX41X1_HVT U991 ( .A1(n912), .A3(n910), .A2(n911), .A4(n909), .S0(n586), 
        .S1(n573), .Y(q[76]) );
  MUX41X1_HVT U992 ( .A1(\ram[12][77] ), .A3(\ram[14][77] ), .A2(\ram[13][77] ), .A4(\ram[15][77] ), .S0(n487), .S1(n394), .Y(n913) );
  MUX41X1_HVT U993 ( .A1(\ram[8][77] ), .A3(\ram[10][77] ), .A2(\ram[9][77] ), 
        .A4(\ram[11][77] ), .S0(n487), .S1(n394), .Y(n914) );
  MUX41X1_HVT U994 ( .A1(\ram[4][77] ), .A3(\ram[6][77] ), .A2(\ram[5][77] ), 
        .A4(\ram[7][77] ), .S0(n487), .S1(n394), .Y(n915) );
  MUX41X1_HVT U995 ( .A1(\ram[0][77] ), .A3(\ram[2][77] ), .A2(\ram[1][77] ), 
        .A4(\ram[3][77] ), .S0(n487), .S1(n394), .Y(n916) );
  MUX41X1_HVT U996 ( .A1(n916), .A3(n914), .A2(n915), .A4(n913), .S0(n586), 
        .S1(n574), .Y(q[77]) );
  MUX41X1_HVT U997 ( .A1(\ram[12][78] ), .A3(\ram[14][78] ), .A2(\ram[13][78] ), .A4(\ram[15][78] ), .S0(n488), .S1(n395), .Y(n917) );
  MUX41X1_HVT U998 ( .A1(\ram[8][78] ), .A3(\ram[10][78] ), .A2(\ram[9][78] ), 
        .A4(\ram[11][78] ), .S0(n488), .S1(n395), .Y(n918) );
  MUX41X1_HVT U999 ( .A1(\ram[4][78] ), .A3(\ram[6][78] ), .A2(\ram[5][78] ), 
        .A4(\ram[7][78] ), .S0(n488), .S1(n395), .Y(n919) );
  MUX41X1_HVT U1000 ( .A1(\ram[0][78] ), .A3(\ram[2][78] ), .A2(\ram[1][78] ), 
        .A4(\ram[3][78] ), .S0(n488), .S1(n395), .Y(n920) );
  MUX41X1_HVT U1001 ( .A1(n920), .A3(n918), .A2(n919), .A4(n917), .S0(n586), 
        .S1(n574), .Y(q[78]) );
  MUX41X1_HVT U1002 ( .A1(\ram[12][79] ), .A3(\ram[14][79] ), .A2(
        \ram[13][79] ), .A4(\ram[15][79] ), .S0(n488), .S1(n395), .Y(n921) );
  MUX41X1_HVT U1003 ( .A1(\ram[8][79] ), .A3(\ram[10][79] ), .A2(\ram[9][79] ), 
        .A4(\ram[11][79] ), .S0(n488), .S1(n395), .Y(n922) );
  MUX41X1_HVT U1004 ( .A1(\ram[4][79] ), .A3(\ram[6][79] ), .A2(\ram[5][79] ), 
        .A4(\ram[7][79] ), .S0(n488), .S1(n395), .Y(n923) );
  MUX41X1_HVT U1005 ( .A1(\ram[0][79] ), .A3(\ram[2][79] ), .A2(\ram[1][79] ), 
        .A4(\ram[3][79] ), .S0(n488), .S1(n395), .Y(n924) );
  MUX41X1_HVT U1006 ( .A1(n924), .A3(n922), .A2(n923), .A4(n921), .S0(n586), 
        .S1(n574), .Y(q[79]) );
  MUX41X1_HVT U1007 ( .A1(\ram[12][80] ), .A3(\ram[14][80] ), .A2(
        \ram[13][80] ), .A4(\ram[15][80] ), .S0(n488), .S1(n395), .Y(n925) );
  MUX41X1_HVT U1008 ( .A1(\ram[8][80] ), .A3(\ram[10][80] ), .A2(\ram[9][80] ), 
        .A4(\ram[11][80] ), .S0(n488), .S1(n395), .Y(n926) );
  MUX41X1_HVT U1009 ( .A1(\ram[4][80] ), .A3(\ram[6][80] ), .A2(\ram[5][80] ), 
        .A4(\ram[7][80] ), .S0(n488), .S1(n395), .Y(n927) );
  MUX41X1_HVT U1010 ( .A1(\ram[0][80] ), .A3(\ram[2][80] ), .A2(\ram[1][80] ), 
        .A4(\ram[3][80] ), .S0(n488), .S1(n395), .Y(n928) );
  MUX41X1_HVT U1011 ( .A1(n928), .A3(n926), .A2(n927), .A4(n925), .S0(n586), 
        .S1(n574), .Y(q[80]) );
  MUX41X1_HVT U1012 ( .A1(\ram[12][81] ), .A3(\ram[14][81] ), .A2(
        \ram[13][81] ), .A4(\ram[15][81] ), .S0(n489), .S1(n396), .Y(n929) );
  MUX41X1_HVT U1013 ( .A1(\ram[8][81] ), .A3(\ram[10][81] ), .A2(\ram[9][81] ), 
        .A4(\ram[11][81] ), .S0(n489), .S1(n396), .Y(n930) );
  MUX41X1_HVT U1014 ( .A1(\ram[4][81] ), .A3(\ram[6][81] ), .A2(\ram[5][81] ), 
        .A4(\ram[7][81] ), .S0(n489), .S1(n396), .Y(n931) );
  MUX41X1_HVT U1015 ( .A1(\ram[0][81] ), .A3(\ram[2][81] ), .A2(\ram[1][81] ), 
        .A4(\ram[3][81] ), .S0(n489), .S1(n396), .Y(n932) );
  MUX41X1_HVT U1016 ( .A1(n932), .A3(n930), .A2(n931), .A4(n929), .S0(n586), 
        .S1(n574), .Y(q[81]) );
  MUX41X1_HVT U1017 ( .A1(\ram[12][82] ), .A3(\ram[14][82] ), .A2(
        \ram[13][82] ), .A4(\ram[15][82] ), .S0(n489), .S1(n396), .Y(n933) );
  MUX41X1_HVT U1018 ( .A1(\ram[8][82] ), .A3(\ram[10][82] ), .A2(\ram[9][82] ), 
        .A4(\ram[11][82] ), .S0(n489), .S1(n396), .Y(n934) );
  MUX41X1_HVT U1019 ( .A1(\ram[4][82] ), .A3(\ram[6][82] ), .A2(\ram[5][82] ), 
        .A4(\ram[7][82] ), .S0(n489), .S1(n396), .Y(n935) );
  MUX41X1_HVT U1020 ( .A1(\ram[0][82] ), .A3(\ram[2][82] ), .A2(\ram[1][82] ), 
        .A4(\ram[3][82] ), .S0(n489), .S1(n396), .Y(n936) );
  MUX41X1_HVT U1021 ( .A1(n936), .A3(n934), .A2(n935), .A4(n933), .S0(n586), 
        .S1(n574), .Y(q[82]) );
  MUX41X1_HVT U1022 ( .A1(\ram[12][83] ), .A3(\ram[14][83] ), .A2(
        \ram[13][83] ), .A4(\ram[15][83] ), .S0(n489), .S1(n396), .Y(n937) );
  MUX41X1_HVT U1023 ( .A1(\ram[8][83] ), .A3(\ram[10][83] ), .A2(\ram[9][83] ), 
        .A4(\ram[11][83] ), .S0(n489), .S1(n396), .Y(n938) );
  MUX41X1_HVT U1024 ( .A1(\ram[4][83] ), .A3(\ram[6][83] ), .A2(\ram[5][83] ), 
        .A4(\ram[7][83] ), .S0(n489), .S1(n396), .Y(n939) );
  MUX41X1_HVT U1025 ( .A1(\ram[0][83] ), .A3(\ram[2][83] ), .A2(\ram[1][83] ), 
        .A4(\ram[3][83] ), .S0(n489), .S1(n396), .Y(n940) );
  MUX41X1_HVT U1026 ( .A1(n940), .A3(n938), .A2(n939), .A4(n937), .S0(n586), 
        .S1(n574), .Y(q[83]) );
  MUX41X1_HVT U1027 ( .A1(\ram[12][84] ), .A3(\ram[14][84] ), .A2(
        \ram[13][84] ), .A4(\ram[15][84] ), .S0(n490), .S1(n397), .Y(n941) );
  MUX41X1_HVT U1028 ( .A1(\ram[8][84] ), .A3(\ram[10][84] ), .A2(\ram[9][84] ), 
        .A4(\ram[11][84] ), .S0(n490), .S1(n397), .Y(n942) );
  MUX41X1_HVT U1029 ( .A1(\ram[4][84] ), .A3(\ram[6][84] ), .A2(\ram[5][84] ), 
        .A4(\ram[7][84] ), .S0(n490), .S1(n397), .Y(n943) );
  MUX41X1_HVT U1030 ( .A1(\ram[0][84] ), .A3(\ram[2][84] ), .A2(\ram[1][84] ), 
        .A4(\ram[3][84] ), .S0(n490), .S1(n397), .Y(n944) );
  MUX41X1_HVT U1031 ( .A1(n944), .A3(n942), .A2(n943), .A4(n941), .S0(n587), 
        .S1(n574), .Y(q[84]) );
  MUX41X1_HVT U1032 ( .A1(\ram[12][85] ), .A3(\ram[14][85] ), .A2(
        \ram[13][85] ), .A4(\ram[15][85] ), .S0(n490), .S1(n397), .Y(n945) );
  MUX41X1_HVT U1033 ( .A1(\ram[8][85] ), .A3(\ram[10][85] ), .A2(\ram[9][85] ), 
        .A4(\ram[11][85] ), .S0(n490), .S1(n397), .Y(n946) );
  MUX41X1_HVT U1034 ( .A1(\ram[4][85] ), .A3(\ram[6][85] ), .A2(\ram[5][85] ), 
        .A4(\ram[7][85] ), .S0(n490), .S1(n397), .Y(n947) );
  MUX41X1_HVT U1035 ( .A1(\ram[0][85] ), .A3(\ram[2][85] ), .A2(\ram[1][85] ), 
        .A4(\ram[3][85] ), .S0(n490), .S1(n397), .Y(n948) );
  MUX41X1_HVT U1036 ( .A1(n948), .A3(n946), .A2(n947), .A4(n945), .S0(n587), 
        .S1(n574), .Y(q[85]) );
  MUX41X1_HVT U1037 ( .A1(\ram[12][86] ), .A3(\ram[14][86] ), .A2(
        \ram[13][86] ), .A4(\ram[15][86] ), .S0(n490), .S1(n397), .Y(n949) );
  MUX41X1_HVT U1038 ( .A1(\ram[8][86] ), .A3(\ram[10][86] ), .A2(\ram[9][86] ), 
        .A4(\ram[11][86] ), .S0(n490), .S1(n397), .Y(n950) );
  MUX41X1_HVT U1039 ( .A1(\ram[4][86] ), .A3(\ram[6][86] ), .A2(\ram[5][86] ), 
        .A4(\ram[7][86] ), .S0(n490), .S1(n397), .Y(n951) );
  MUX41X1_HVT U1040 ( .A1(\ram[0][86] ), .A3(\ram[2][86] ), .A2(\ram[1][86] ), 
        .A4(\ram[3][86] ), .S0(n490), .S1(n397), .Y(n952) );
  MUX41X1_HVT U1041 ( .A1(n952), .A3(n950), .A2(n951), .A4(n949), .S0(n587), 
        .S1(n574), .Y(q[86]) );
  MUX41X1_HVT U1042 ( .A1(\ram[12][87] ), .A3(\ram[14][87] ), .A2(
        \ram[13][87] ), .A4(\ram[15][87] ), .S0(n491), .S1(n398), .Y(n953) );
  MUX41X1_HVT U1043 ( .A1(\ram[8][87] ), .A3(\ram[10][87] ), .A2(\ram[9][87] ), 
        .A4(\ram[11][87] ), .S0(n491), .S1(n398), .Y(n954) );
  MUX41X1_HVT U1044 ( .A1(\ram[4][87] ), .A3(\ram[6][87] ), .A2(\ram[5][87] ), 
        .A4(\ram[7][87] ), .S0(n491), .S1(n398), .Y(n955) );
  MUX41X1_HVT U1045 ( .A1(\ram[0][87] ), .A3(\ram[2][87] ), .A2(\ram[1][87] ), 
        .A4(\ram[3][87] ), .S0(n491), .S1(n398), .Y(n956) );
  MUX41X1_HVT U1046 ( .A1(n956), .A3(n954), .A2(n955), .A4(n953), .S0(n587), 
        .S1(n575), .Y(q[87]) );
  MUX41X1_HVT U1047 ( .A1(\ram[12][88] ), .A3(\ram[14][88] ), .A2(
        \ram[13][88] ), .A4(\ram[15][88] ), .S0(n491), .S1(n398), .Y(n957) );
  MUX41X1_HVT U1048 ( .A1(\ram[8][88] ), .A3(\ram[10][88] ), .A2(\ram[9][88] ), 
        .A4(\ram[11][88] ), .S0(n491), .S1(n398), .Y(n958) );
  MUX41X1_HVT U1049 ( .A1(\ram[4][88] ), .A3(\ram[6][88] ), .A2(\ram[5][88] ), 
        .A4(\ram[7][88] ), .S0(n491), .S1(n398), .Y(n959) );
  MUX41X1_HVT U1050 ( .A1(\ram[0][88] ), .A3(\ram[2][88] ), .A2(\ram[1][88] ), 
        .A4(\ram[3][88] ), .S0(n491), .S1(n398), .Y(n960) );
  MUX41X1_HVT U1051 ( .A1(n960), .A3(n958), .A2(n959), .A4(n957), .S0(n587), 
        .S1(n574), .Y(q[88]) );
  MUX41X1_HVT U1052 ( .A1(\ram[12][89] ), .A3(\ram[14][89] ), .A2(
        \ram[13][89] ), .A4(\ram[15][89] ), .S0(n491), .S1(n398), .Y(n961) );
  MUX41X1_HVT U1053 ( .A1(\ram[8][89] ), .A3(\ram[10][89] ), .A2(\ram[9][89] ), 
        .A4(\ram[11][89] ), .S0(n491), .S1(n398), .Y(n962) );
  MUX41X1_HVT U1054 ( .A1(\ram[4][89] ), .A3(\ram[6][89] ), .A2(\ram[5][89] ), 
        .A4(\ram[7][89] ), .S0(n491), .S1(n398), .Y(n963) );
  MUX41X1_HVT U1055 ( .A1(\ram[0][89] ), .A3(\ram[2][89] ), .A2(\ram[1][89] ), 
        .A4(\ram[3][89] ), .S0(n491), .S1(n398), .Y(n964) );
  MUX41X1_HVT U1056 ( .A1(n964), .A3(n962), .A2(n963), .A4(n961), .S0(n587), 
        .S1(n575), .Y(q[89]) );
  MUX41X1_HVT U1057 ( .A1(\ram[12][90] ), .A3(\ram[14][90] ), .A2(
        \ram[13][90] ), .A4(\ram[15][90] ), .S0(n492), .S1(n399), .Y(n965) );
  MUX41X1_HVT U1058 ( .A1(\ram[8][90] ), .A3(\ram[10][90] ), .A2(\ram[9][90] ), 
        .A4(\ram[11][90] ), .S0(n492), .S1(n399), .Y(n966) );
  MUX41X1_HVT U1059 ( .A1(\ram[4][90] ), .A3(\ram[6][90] ), .A2(\ram[5][90] ), 
        .A4(\ram[7][90] ), .S0(n492), .S1(n399), .Y(n967) );
  MUX41X1_HVT U1060 ( .A1(\ram[0][90] ), .A3(\ram[2][90] ), .A2(\ram[1][90] ), 
        .A4(\ram[3][90] ), .S0(n492), .S1(n399), .Y(n968) );
  MUX41X1_HVT U1061 ( .A1(n968), .A3(n966), .A2(n967), .A4(n965), .S0(n587), 
        .S1(n575), .Y(q[90]) );
  MUX41X1_HVT U1062 ( .A1(\ram[12][91] ), .A3(\ram[14][91] ), .A2(
        \ram[13][91] ), .A4(\ram[15][91] ), .S0(n492), .S1(n399), .Y(n969) );
  MUX41X1_HVT U1063 ( .A1(\ram[8][91] ), .A3(\ram[10][91] ), .A2(\ram[9][91] ), 
        .A4(\ram[11][91] ), .S0(n492), .S1(n399), .Y(n970) );
  MUX41X1_HVT U1064 ( .A1(\ram[4][91] ), .A3(\ram[6][91] ), .A2(\ram[5][91] ), 
        .A4(\ram[7][91] ), .S0(n492), .S1(n399), .Y(n971) );
  MUX41X1_HVT U1065 ( .A1(\ram[0][91] ), .A3(\ram[2][91] ), .A2(\ram[1][91] ), 
        .A4(\ram[3][91] ), .S0(n492), .S1(n399), .Y(n972) );
  MUX41X1_HVT U1066 ( .A1(n972), .A3(n970), .A2(n971), .A4(n969), .S0(n587), 
        .S1(n575), .Y(q[91]) );
  MUX41X1_HVT U1067 ( .A1(\ram[12][92] ), .A3(\ram[14][92] ), .A2(
        \ram[13][92] ), .A4(\ram[15][92] ), .S0(n492), .S1(n399), .Y(n973) );
  MUX41X1_HVT U1068 ( .A1(\ram[8][92] ), .A3(\ram[10][92] ), .A2(\ram[9][92] ), 
        .A4(\ram[11][92] ), .S0(n492), .S1(n399), .Y(n974) );
  MUX41X1_HVT U1069 ( .A1(\ram[4][92] ), .A3(\ram[6][92] ), .A2(\ram[5][92] ), 
        .A4(\ram[7][92] ), .S0(n492), .S1(n399), .Y(n975) );
  MUX41X1_HVT U1070 ( .A1(\ram[0][92] ), .A3(\ram[2][92] ), .A2(\ram[1][92] ), 
        .A4(\ram[3][92] ), .S0(n492), .S1(n399), .Y(n976) );
  MUX41X1_HVT U1071 ( .A1(n976), .A3(n974), .A2(n975), .A4(n973), .S0(n587), 
        .S1(n575), .Y(q[92]) );
  MUX41X1_HVT U1072 ( .A1(\ram[12][93] ), .A3(\ram[14][93] ), .A2(
        \ram[13][93] ), .A4(\ram[15][93] ), .S0(n493), .S1(n400), .Y(n977) );
  MUX41X1_HVT U1073 ( .A1(\ram[8][93] ), .A3(\ram[10][93] ), .A2(\ram[9][93] ), 
        .A4(\ram[11][93] ), .S0(n493), .S1(n400), .Y(n978) );
  MUX41X1_HVT U1074 ( .A1(\ram[4][93] ), .A3(\ram[6][93] ), .A2(\ram[5][93] ), 
        .A4(\ram[7][93] ), .S0(n493), .S1(n400), .Y(n979) );
  MUX41X1_HVT U1075 ( .A1(\ram[0][93] ), .A3(\ram[2][93] ), .A2(\ram[1][93] ), 
        .A4(\ram[3][93] ), .S0(n493), .S1(n400), .Y(n980) );
  MUX41X1_HVT U1076 ( .A1(n980), .A3(n978), .A2(n979), .A4(n977), .S0(n587), 
        .S1(n575), .Y(q[93]) );
  MUX41X1_HVT U1077 ( .A1(\ram[12][94] ), .A3(\ram[14][94] ), .A2(
        \ram[13][94] ), .A4(\ram[15][94] ), .S0(n493), .S1(n400), .Y(n981) );
  MUX41X1_HVT U1078 ( .A1(\ram[8][94] ), .A3(\ram[10][94] ), .A2(\ram[9][94] ), 
        .A4(\ram[11][94] ), .S0(n493), .S1(n400), .Y(n982) );
  MUX41X1_HVT U1079 ( .A1(\ram[4][94] ), .A3(\ram[6][94] ), .A2(\ram[5][94] ), 
        .A4(\ram[7][94] ), .S0(n493), .S1(n400), .Y(n983) );
  MUX41X1_HVT U1080 ( .A1(\ram[0][94] ), .A3(\ram[2][94] ), .A2(\ram[1][94] ), 
        .A4(\ram[3][94] ), .S0(n493), .S1(n400), .Y(n984) );
  MUX41X1_HVT U1081 ( .A1(n984), .A3(n982), .A2(n983), .A4(n981), .S0(n587), 
        .S1(n575), .Y(q[94]) );
  MUX41X1_HVT U1082 ( .A1(\ram[12][95] ), .A3(\ram[14][95] ), .A2(
        \ram[13][95] ), .A4(\ram[15][95] ), .S0(n493), .S1(n400), .Y(n985) );
  MUX41X1_HVT U1083 ( .A1(\ram[8][95] ), .A3(\ram[10][95] ), .A2(\ram[9][95] ), 
        .A4(\ram[11][95] ), .S0(n493), .S1(n400), .Y(n986) );
  MUX41X1_HVT U1084 ( .A1(\ram[4][95] ), .A3(\ram[6][95] ), .A2(\ram[5][95] ), 
        .A4(\ram[7][95] ), .S0(n493), .S1(n400), .Y(n987) );
  MUX41X1_HVT U1085 ( .A1(\ram[0][95] ), .A3(\ram[2][95] ), .A2(\ram[1][95] ), 
        .A4(\ram[3][95] ), .S0(n493), .S1(n400), .Y(n988) );
  MUX41X1_HVT U1086 ( .A1(n988), .A3(n986), .A2(n987), .A4(n985), .S0(n587), 
        .S1(n575), .Y(q[95]) );
  MUX41X1_HVT U1087 ( .A1(\ram[12][96] ), .A3(\ram[14][96] ), .A2(
        \ram[13][96] ), .A4(\ram[15][96] ), .S0(n494), .S1(n401), .Y(n989) );
  MUX41X1_HVT U1088 ( .A1(\ram[8][96] ), .A3(\ram[10][96] ), .A2(\ram[9][96] ), 
        .A4(\ram[11][96] ), .S0(n494), .S1(n401), .Y(n990) );
  MUX41X1_HVT U1089 ( .A1(\ram[4][96] ), .A3(\ram[6][96] ), .A2(\ram[5][96] ), 
        .A4(\ram[7][96] ), .S0(n494), .S1(n401), .Y(n991) );
  MUX41X1_HVT U1090 ( .A1(\ram[0][96] ), .A3(\ram[2][96] ), .A2(\ram[1][96] ), 
        .A4(\ram[3][96] ), .S0(n494), .S1(n401), .Y(n992) );
  MUX41X1_HVT U1091 ( .A1(n992), .A3(n990), .A2(n991), .A4(n989), .S0(n588), 
        .S1(n575), .Y(q[96]) );
  MUX41X1_HVT U1092 ( .A1(\ram[12][97] ), .A3(\ram[14][97] ), .A2(
        \ram[13][97] ), .A4(\ram[15][97] ), .S0(n494), .S1(n401), .Y(n993) );
  MUX41X1_HVT U1093 ( .A1(\ram[8][97] ), .A3(\ram[10][97] ), .A2(\ram[9][97] ), 
        .A4(\ram[11][97] ), .S0(n494), .S1(n401), .Y(n994) );
  MUX41X1_HVT U1094 ( .A1(\ram[4][97] ), .A3(\ram[6][97] ), .A2(\ram[5][97] ), 
        .A4(\ram[7][97] ), .S0(n494), .S1(n401), .Y(n995) );
  MUX41X1_HVT U1095 ( .A1(\ram[0][97] ), .A3(\ram[2][97] ), .A2(\ram[1][97] ), 
        .A4(\ram[3][97] ), .S0(n494), .S1(n401), .Y(n996) );
  MUX41X1_HVT U1096 ( .A1(n996), .A3(n994), .A2(n995), .A4(n993), .S0(n588), 
        .S1(n575), .Y(q[97]) );
  MUX41X1_HVT U1097 ( .A1(\ram[12][98] ), .A3(\ram[14][98] ), .A2(
        \ram[13][98] ), .A4(\ram[15][98] ), .S0(n494), .S1(n401), .Y(n997) );
  MUX41X1_HVT U1098 ( .A1(\ram[8][98] ), .A3(\ram[10][98] ), .A2(\ram[9][98] ), 
        .A4(\ram[11][98] ), .S0(n494), .S1(n401), .Y(n998) );
  MUX41X1_HVT U1099 ( .A1(\ram[4][98] ), .A3(\ram[6][98] ), .A2(\ram[5][98] ), 
        .A4(\ram[7][98] ), .S0(n494), .S1(n401), .Y(n999) );
  MUX41X1_HVT U1100 ( .A1(\ram[0][98] ), .A3(\ram[2][98] ), .A2(\ram[1][98] ), 
        .A4(\ram[3][98] ), .S0(n494), .S1(n401), .Y(n1000) );
  MUX41X1_HVT U1101 ( .A1(n1000), .A3(n998), .A2(n999), .A4(n997), .S0(n588), 
        .S1(n575), .Y(q[98]) );
  MUX41X1_HVT U1102 ( .A1(\ram[12][99] ), .A3(\ram[14][99] ), .A2(
        \ram[13][99] ), .A4(\ram[15][99] ), .S0(n495), .S1(n402), .Y(n1001) );
  MUX41X1_HVT U1103 ( .A1(\ram[8][99] ), .A3(\ram[10][99] ), .A2(\ram[9][99] ), 
        .A4(\ram[11][99] ), .S0(n495), .S1(n402), .Y(n1002) );
  MUX41X1_HVT U1104 ( .A1(\ram[4][99] ), .A3(\ram[6][99] ), .A2(\ram[5][99] ), 
        .A4(\ram[7][99] ), .S0(n495), .S1(n402), .Y(n1003) );
  MUX41X1_HVT U1105 ( .A1(\ram[0][99] ), .A3(\ram[2][99] ), .A2(\ram[1][99] ), 
        .A4(\ram[3][99] ), .S0(n495), .S1(n402), .Y(n1004) );
  MUX41X1_HVT U1106 ( .A1(n1004), .A3(n1002), .A2(n1003), .A4(n1001), .S0(n588), .S1(n576), .Y(q[99]) );
  MUX41X1_HVT U1107 ( .A1(\ram[12][100] ), .A3(\ram[14][100] ), .A2(
        \ram[13][100] ), .A4(\ram[15][100] ), .S0(n495), .S1(n402), .Y(n1005)
         );
  MUX41X1_HVT U1108 ( .A1(\ram[8][100] ), .A3(\ram[10][100] ), .A2(
        \ram[9][100] ), .A4(\ram[11][100] ), .S0(n495), .S1(n402), .Y(n1006)
         );
  MUX41X1_HVT U1109 ( .A1(\ram[4][100] ), .A3(\ram[6][100] ), .A2(
        \ram[5][100] ), .A4(\ram[7][100] ), .S0(n495), .S1(n402), .Y(n1007) );
  MUX41X1_HVT U1110 ( .A1(\ram[0][100] ), .A3(\ram[2][100] ), .A2(
        \ram[1][100] ), .A4(\ram[3][100] ), .S0(n495), .S1(n402), .Y(n1008) );
  MUX41X1_HVT U1111 ( .A1(n1008), .A3(n1006), .A2(n1007), .A4(n1005), .S0(n588), .S1(n575), .Y(q[100]) );
  MUX41X1_HVT U1112 ( .A1(\ram[12][101] ), .A3(\ram[14][101] ), .A2(
        \ram[13][101] ), .A4(\ram[15][101] ), .S0(n495), .S1(n402), .Y(n1009)
         );
  MUX41X1_HVT U1113 ( .A1(\ram[8][101] ), .A3(\ram[10][101] ), .A2(
        \ram[9][101] ), .A4(\ram[11][101] ), .S0(n495), .S1(n402), .Y(n1010)
         );
  MUX41X1_HVT U1114 ( .A1(\ram[4][101] ), .A3(\ram[6][101] ), .A2(
        \ram[5][101] ), .A4(\ram[7][101] ), .S0(n495), .S1(n402), .Y(n1011) );
  MUX41X1_HVT U1115 ( .A1(\ram[0][101] ), .A3(\ram[2][101] ), .A2(
        \ram[1][101] ), .A4(\ram[3][101] ), .S0(n495), .S1(n402), .Y(n1012) );
  MUX41X1_HVT U1116 ( .A1(n1012), .A3(n1010), .A2(n1011), .A4(n1009), .S0(n588), .S1(n576), .Y(q[101]) );
  MUX41X1_HVT U1117 ( .A1(\ram[12][102] ), .A3(\ram[14][102] ), .A2(
        \ram[13][102] ), .A4(\ram[15][102] ), .S0(n496), .S1(n403), .Y(n1013)
         );
  MUX41X1_HVT U1118 ( .A1(\ram[8][102] ), .A3(\ram[10][102] ), .A2(
        \ram[9][102] ), .A4(\ram[11][102] ), .S0(n496), .S1(n403), .Y(n1014)
         );
  MUX41X1_HVT U1119 ( .A1(\ram[4][102] ), .A3(\ram[6][102] ), .A2(
        \ram[5][102] ), .A4(\ram[7][102] ), .S0(n496), .S1(n403), .Y(n1015) );
  MUX41X1_HVT U1120 ( .A1(\ram[0][102] ), .A3(\ram[2][102] ), .A2(
        \ram[1][102] ), .A4(\ram[3][102] ), .S0(n496), .S1(n403), .Y(n1016) );
  MUX41X1_HVT U1121 ( .A1(n1016), .A3(n1014), .A2(n1015), .A4(n1013), .S0(n588), .S1(n576), .Y(q[102]) );
  MUX41X1_HVT U1122 ( .A1(\ram[12][103] ), .A3(\ram[14][103] ), .A2(
        \ram[13][103] ), .A4(\ram[15][103] ), .S0(n496), .S1(n403), .Y(n1017)
         );
  MUX41X1_HVT U1123 ( .A1(\ram[8][103] ), .A3(\ram[10][103] ), .A2(
        \ram[9][103] ), .A4(\ram[11][103] ), .S0(n496), .S1(n403), .Y(n1018)
         );
  MUX41X1_HVT U1124 ( .A1(\ram[4][103] ), .A3(\ram[6][103] ), .A2(
        \ram[5][103] ), .A4(\ram[7][103] ), .S0(n496), .S1(n403), .Y(n1019) );
  MUX41X1_HVT U1125 ( .A1(\ram[0][103] ), .A3(\ram[2][103] ), .A2(
        \ram[1][103] ), .A4(\ram[3][103] ), .S0(n496), .S1(n403), .Y(n1020) );
  MUX41X1_HVT U1126 ( .A1(n1020), .A3(n1018), .A2(n1019), .A4(n1017), .S0(n588), .S1(n576), .Y(q[103]) );
  MUX41X1_HVT U1127 ( .A1(\ram[12][104] ), .A3(\ram[14][104] ), .A2(
        \ram[13][104] ), .A4(\ram[15][104] ), .S0(n496), .S1(n403), .Y(n1021)
         );
  MUX41X1_HVT U1128 ( .A1(\ram[8][104] ), .A3(\ram[10][104] ), .A2(
        \ram[9][104] ), .A4(\ram[11][104] ), .S0(n496), .S1(n403), .Y(n1022)
         );
  MUX41X1_HVT U1129 ( .A1(\ram[4][104] ), .A3(\ram[6][104] ), .A2(
        \ram[5][104] ), .A4(\ram[7][104] ), .S0(n496), .S1(n403), .Y(n1023) );
  MUX41X1_HVT U1130 ( .A1(\ram[0][104] ), .A3(\ram[2][104] ), .A2(
        \ram[1][104] ), .A4(\ram[3][104] ), .S0(n496), .S1(n403), .Y(n1024) );
  MUX41X1_HVT U1131 ( .A1(n1024), .A3(n1022), .A2(n1023), .A4(n1021), .S0(n588), .S1(n576), .Y(q[104]) );
  MUX41X1_HVT U1132 ( .A1(\ram[12][105] ), .A3(\ram[14][105] ), .A2(
        \ram[13][105] ), .A4(\ram[15][105] ), .S0(n497), .S1(n404), .Y(n1025)
         );
  MUX41X1_HVT U1133 ( .A1(\ram[8][105] ), .A3(\ram[10][105] ), .A2(
        \ram[9][105] ), .A4(\ram[11][105] ), .S0(n497), .S1(n404), .Y(n1026)
         );
  MUX41X1_HVT U1134 ( .A1(\ram[4][105] ), .A3(\ram[6][105] ), .A2(
        \ram[5][105] ), .A4(\ram[7][105] ), .S0(n497), .S1(n404), .Y(n1027) );
  MUX41X1_HVT U1135 ( .A1(\ram[0][105] ), .A3(\ram[2][105] ), .A2(
        \ram[1][105] ), .A4(\ram[3][105] ), .S0(n497), .S1(n404), .Y(n1028) );
  MUX41X1_HVT U1136 ( .A1(n1028), .A3(n1026), .A2(n1027), .A4(n1025), .S0(n588), .S1(n576), .Y(q[105]) );
  MUX41X1_HVT U1137 ( .A1(\ram[12][106] ), .A3(\ram[14][106] ), .A2(
        \ram[13][106] ), .A4(\ram[15][106] ), .S0(n497), .S1(n404), .Y(n1029)
         );
  MUX41X1_HVT U1138 ( .A1(\ram[8][106] ), .A3(\ram[10][106] ), .A2(
        \ram[9][106] ), .A4(\ram[11][106] ), .S0(n497), .S1(n404), .Y(n1030)
         );
  MUX41X1_HVT U1139 ( .A1(\ram[4][106] ), .A3(\ram[6][106] ), .A2(
        \ram[5][106] ), .A4(\ram[7][106] ), .S0(n497), .S1(n404), .Y(n1031) );
  MUX41X1_HVT U1140 ( .A1(\ram[0][106] ), .A3(\ram[2][106] ), .A2(
        \ram[1][106] ), .A4(\ram[3][106] ), .S0(n497), .S1(n404), .Y(n1032) );
  MUX41X1_HVT U1141 ( .A1(n1032), .A3(n1030), .A2(n1031), .A4(n1029), .S0(n588), .S1(n576), .Y(q[106]) );
  MUX41X1_HVT U1142 ( .A1(\ram[12][107] ), .A3(\ram[14][107] ), .A2(
        \ram[13][107] ), .A4(\ram[15][107] ), .S0(n497), .S1(n404), .Y(n1033)
         );
  MUX41X1_HVT U1143 ( .A1(\ram[8][107] ), .A3(\ram[10][107] ), .A2(
        \ram[9][107] ), .A4(\ram[11][107] ), .S0(n497), .S1(n404), .Y(n1034)
         );
  MUX41X1_HVT U1144 ( .A1(\ram[4][107] ), .A3(\ram[6][107] ), .A2(
        \ram[5][107] ), .A4(\ram[7][107] ), .S0(n497), .S1(n404), .Y(n1035) );
  MUX41X1_HVT U1145 ( .A1(\ram[0][107] ), .A3(\ram[2][107] ), .A2(
        \ram[1][107] ), .A4(\ram[3][107] ), .S0(n497), .S1(n404), .Y(n1036) );
  MUX41X1_HVT U1146 ( .A1(n1036), .A3(n1034), .A2(n1035), .A4(n1033), .S0(n588), .S1(n576), .Y(q[107]) );
  MUX41X1_HVT U1147 ( .A1(\ram[12][108] ), .A3(\ram[14][108] ), .A2(
        \ram[13][108] ), .A4(\ram[15][108] ), .S0(n498), .S1(n405), .Y(n1037)
         );
  MUX41X1_HVT U1148 ( .A1(\ram[8][108] ), .A3(\ram[10][108] ), .A2(
        \ram[9][108] ), .A4(\ram[11][108] ), .S0(n498), .S1(n405), .Y(n1038)
         );
  MUX41X1_HVT U1149 ( .A1(\ram[4][108] ), .A3(\ram[6][108] ), .A2(
        \ram[5][108] ), .A4(\ram[7][108] ), .S0(n498), .S1(n405), .Y(n1039) );
  MUX41X1_HVT U1150 ( .A1(\ram[0][108] ), .A3(\ram[2][108] ), .A2(
        \ram[1][108] ), .A4(\ram[3][108] ), .S0(n498), .S1(n405), .Y(n1040) );
  MUX41X1_HVT U1151 ( .A1(n1040), .A3(n1038), .A2(n1039), .A4(n1037), .S0(n589), .S1(n576), .Y(q[108]) );
  MUX41X1_HVT U1152 ( .A1(\ram[12][109] ), .A3(\ram[14][109] ), .A2(
        \ram[13][109] ), .A4(\ram[15][109] ), .S0(n498), .S1(n405), .Y(n1041)
         );
  MUX41X1_HVT U1153 ( .A1(\ram[8][109] ), .A3(\ram[10][109] ), .A2(
        \ram[9][109] ), .A4(\ram[11][109] ), .S0(n498), .S1(n405), .Y(n1042)
         );
  MUX41X1_HVT U1154 ( .A1(\ram[4][109] ), .A3(\ram[6][109] ), .A2(
        \ram[5][109] ), .A4(\ram[7][109] ), .S0(n498), .S1(n405), .Y(n1043) );
  MUX41X1_HVT U1155 ( .A1(\ram[0][109] ), .A3(\ram[2][109] ), .A2(
        \ram[1][109] ), .A4(\ram[3][109] ), .S0(n498), .S1(n405), .Y(n1044) );
  MUX41X1_HVT U1156 ( .A1(n1044), .A3(n1042), .A2(n1043), .A4(n1041), .S0(n589), .S1(n576), .Y(q[109]) );
  MUX41X1_HVT U1157 ( .A1(\ram[12][110] ), .A3(\ram[14][110] ), .A2(
        \ram[13][110] ), .A4(\ram[15][110] ), .S0(n498), .S1(n405), .Y(n1045)
         );
  MUX41X1_HVT U1158 ( .A1(\ram[8][110] ), .A3(\ram[10][110] ), .A2(
        \ram[9][110] ), .A4(\ram[11][110] ), .S0(n498), .S1(n405), .Y(n1046)
         );
  MUX41X1_HVT U1159 ( .A1(\ram[4][110] ), .A3(\ram[6][110] ), .A2(
        \ram[5][110] ), .A4(\ram[7][110] ), .S0(n498), .S1(n405), .Y(n1047) );
  MUX41X1_HVT U1160 ( .A1(\ram[0][110] ), .A3(\ram[2][110] ), .A2(
        \ram[1][110] ), .A4(\ram[3][110] ), .S0(n498), .S1(n405), .Y(n1048) );
  MUX41X1_HVT U1161 ( .A1(n1048), .A3(n1046), .A2(n1047), .A4(n1045), .S0(n589), .S1(n576), .Y(q[110]) );
  MUX41X1_HVT U1162 ( .A1(\ram[12][111] ), .A3(\ram[14][111] ), .A2(
        \ram[13][111] ), .A4(\ram[15][111] ), .S0(n499), .S1(n406), .Y(n1049)
         );
  MUX41X1_HVT U1163 ( .A1(\ram[8][111] ), .A3(\ram[10][111] ), .A2(
        \ram[9][111] ), .A4(\ram[11][111] ), .S0(n499), .S1(n406), .Y(n1050)
         );
  MUX41X1_HVT U1164 ( .A1(\ram[4][111] ), .A3(\ram[6][111] ), .A2(
        \ram[5][111] ), .A4(\ram[7][111] ), .S0(n499), .S1(n406), .Y(n1051) );
  MUX41X1_HVT U1165 ( .A1(\ram[0][111] ), .A3(\ram[2][111] ), .A2(
        \ram[1][111] ), .A4(\ram[3][111] ), .S0(n499), .S1(n406), .Y(n1052) );
  MUX41X1_HVT U1166 ( .A1(n1052), .A3(n1050), .A2(n1051), .A4(n1049), .S0(n589), .S1(n577), .Y(q[111]) );
  MUX41X1_HVT U1167 ( .A1(\ram[12][112] ), .A3(\ram[14][112] ), .A2(
        \ram[13][112] ), .A4(\ram[15][112] ), .S0(n499), .S1(n406), .Y(n1053)
         );
  MUX41X1_HVT U1168 ( .A1(\ram[8][112] ), .A3(\ram[10][112] ), .A2(
        \ram[9][112] ), .A4(\ram[11][112] ), .S0(n499), .S1(n406), .Y(n1054)
         );
  MUX41X1_HVT U1169 ( .A1(\ram[4][112] ), .A3(\ram[6][112] ), .A2(
        \ram[5][112] ), .A4(\ram[7][112] ), .S0(n499), .S1(n406), .Y(n1055) );
  MUX41X1_HVT U1170 ( .A1(\ram[0][112] ), .A3(\ram[2][112] ), .A2(
        \ram[1][112] ), .A4(\ram[3][112] ), .S0(n499), .S1(n406), .Y(n1056) );
  MUX41X1_HVT U1171 ( .A1(n1056), .A3(n1054), .A2(n1055), .A4(n1053), .S0(n589), .S1(n576), .Y(q[112]) );
  MUX41X1_HVT U1172 ( .A1(\ram[12][113] ), .A3(\ram[14][113] ), .A2(
        \ram[13][113] ), .A4(\ram[15][113] ), .S0(n499), .S1(n406), .Y(n1057)
         );
  MUX41X1_HVT U1173 ( .A1(\ram[8][113] ), .A3(\ram[10][113] ), .A2(
        \ram[9][113] ), .A4(\ram[11][113] ), .S0(n499), .S1(n406), .Y(n1058)
         );
  MUX41X1_HVT U1174 ( .A1(\ram[4][113] ), .A3(\ram[6][113] ), .A2(
        \ram[5][113] ), .A4(\ram[7][113] ), .S0(n499), .S1(n406), .Y(n1059) );
  MUX41X1_HVT U1175 ( .A1(\ram[0][113] ), .A3(\ram[2][113] ), .A2(
        \ram[1][113] ), .A4(\ram[3][113] ), .S0(n499), .S1(n406), .Y(n1060) );
  MUX41X1_HVT U1176 ( .A1(n1060), .A3(n1058), .A2(n1059), .A4(n1057), .S0(n589), .S1(n577), .Y(q[113]) );
  MUX41X1_HVT U1177 ( .A1(\ram[12][114] ), .A3(\ram[14][114] ), .A2(
        \ram[13][114] ), .A4(\ram[15][114] ), .S0(n500), .S1(n407), .Y(n1061)
         );
  MUX41X1_HVT U1178 ( .A1(\ram[8][114] ), .A3(\ram[10][114] ), .A2(
        \ram[9][114] ), .A4(\ram[11][114] ), .S0(n500), .S1(n407), .Y(n1062)
         );
  MUX41X1_HVT U1179 ( .A1(\ram[4][114] ), .A3(\ram[6][114] ), .A2(
        \ram[5][114] ), .A4(\ram[7][114] ), .S0(n500), .S1(n407), .Y(n1063) );
  MUX41X1_HVT U1180 ( .A1(\ram[0][114] ), .A3(\ram[2][114] ), .A2(
        \ram[1][114] ), .A4(\ram[3][114] ), .S0(n500), .S1(n407), .Y(n1064) );
  MUX41X1_HVT U1181 ( .A1(n1064), .A3(n1062), .A2(n1063), .A4(n1061), .S0(n589), .S1(n577), .Y(q[114]) );
  MUX41X1_HVT U1182 ( .A1(\ram[12][115] ), .A3(\ram[14][115] ), .A2(
        \ram[13][115] ), .A4(\ram[15][115] ), .S0(n500), .S1(n407), .Y(n1065)
         );
  MUX41X1_HVT U1183 ( .A1(\ram[8][115] ), .A3(\ram[10][115] ), .A2(
        \ram[9][115] ), .A4(\ram[11][115] ), .S0(n500), .S1(n407), .Y(n1066)
         );
  MUX41X1_HVT U1184 ( .A1(\ram[4][115] ), .A3(\ram[6][115] ), .A2(
        \ram[5][115] ), .A4(\ram[7][115] ), .S0(n500), .S1(n407), .Y(n1067) );
  MUX41X1_HVT U1185 ( .A1(\ram[0][115] ), .A3(\ram[2][115] ), .A2(
        \ram[1][115] ), .A4(\ram[3][115] ), .S0(n500), .S1(n407), .Y(n1068) );
  MUX41X1_HVT U1186 ( .A1(n1068), .A3(n1066), .A2(n1067), .A4(n1065), .S0(n589), .S1(n577), .Y(q[115]) );
  MUX41X1_HVT U1187 ( .A1(\ram[12][116] ), .A3(\ram[14][116] ), .A2(
        \ram[13][116] ), .A4(\ram[15][116] ), .S0(n500), .S1(n407), .Y(n1069)
         );
  MUX41X1_HVT U1188 ( .A1(\ram[8][116] ), .A3(\ram[10][116] ), .A2(
        \ram[9][116] ), .A4(\ram[11][116] ), .S0(n500), .S1(n407), .Y(n1070)
         );
  MUX41X1_HVT U1189 ( .A1(\ram[4][116] ), .A3(\ram[6][116] ), .A2(
        \ram[5][116] ), .A4(\ram[7][116] ), .S0(n500), .S1(n407), .Y(n1071) );
  MUX41X1_HVT U1190 ( .A1(\ram[0][116] ), .A3(\ram[2][116] ), .A2(
        \ram[1][116] ), .A4(\ram[3][116] ), .S0(n500), .S1(n407), .Y(n1072) );
  MUX41X1_HVT U1191 ( .A1(n1072), .A3(n1070), .A2(n1071), .A4(n1069), .S0(n589), .S1(n577), .Y(q[116]) );
  MUX41X1_HVT U1192 ( .A1(\ram[12][117] ), .A3(\ram[14][117] ), .A2(
        \ram[13][117] ), .A4(\ram[15][117] ), .S0(n501), .S1(n408), .Y(n1073)
         );
  MUX41X1_HVT U1193 ( .A1(\ram[8][117] ), .A3(\ram[10][117] ), .A2(
        \ram[9][117] ), .A4(\ram[11][117] ), .S0(n501), .S1(n408), .Y(n1074)
         );
  MUX41X1_HVT U1194 ( .A1(\ram[4][117] ), .A3(\ram[6][117] ), .A2(
        \ram[5][117] ), .A4(\ram[7][117] ), .S0(n501), .S1(n408), .Y(n1075) );
  MUX41X1_HVT U1195 ( .A1(\ram[0][117] ), .A3(\ram[2][117] ), .A2(
        \ram[1][117] ), .A4(\ram[3][117] ), .S0(n501), .S1(n408), .Y(n1076) );
  MUX41X1_HVT U1196 ( .A1(n1076), .A3(n1074), .A2(n1075), .A4(n1073), .S0(n589), .S1(n577), .Y(q[117]) );
  MUX41X1_HVT U1197 ( .A1(\ram[12][118] ), .A3(\ram[14][118] ), .A2(
        \ram[13][118] ), .A4(\ram[15][118] ), .S0(n501), .S1(n408), .Y(n1077)
         );
  MUX41X1_HVT U1198 ( .A1(\ram[8][118] ), .A3(\ram[10][118] ), .A2(
        \ram[9][118] ), .A4(\ram[11][118] ), .S0(n501), .S1(n408), .Y(n1078)
         );
  MUX41X1_HVT U1199 ( .A1(\ram[4][118] ), .A3(\ram[6][118] ), .A2(
        \ram[5][118] ), .A4(\ram[7][118] ), .S0(n501), .S1(n408), .Y(n1079) );
  MUX41X1_HVT U1200 ( .A1(\ram[0][118] ), .A3(\ram[2][118] ), .A2(
        \ram[1][118] ), .A4(\ram[3][118] ), .S0(n501), .S1(n408), .Y(n1080) );
  MUX41X1_HVT U1201 ( .A1(n1080), .A3(n1078), .A2(n1079), .A4(n1077), .S0(n589), .S1(n577), .Y(q[118]) );
  MUX41X1_HVT U1202 ( .A1(\ram[12][119] ), .A3(\ram[14][119] ), .A2(
        \ram[13][119] ), .A4(\ram[15][119] ), .S0(n501), .S1(n408), .Y(n1081)
         );
  MUX41X1_HVT U1203 ( .A1(\ram[8][119] ), .A3(\ram[10][119] ), .A2(
        \ram[9][119] ), .A4(\ram[11][119] ), .S0(n501), .S1(n408), .Y(n1082)
         );
  MUX41X1_HVT U1204 ( .A1(\ram[4][119] ), .A3(\ram[6][119] ), .A2(
        \ram[5][119] ), .A4(\ram[7][119] ), .S0(n501), .S1(n408), .Y(n1083) );
  MUX41X1_HVT U1205 ( .A1(\ram[0][119] ), .A3(\ram[2][119] ), .A2(
        \ram[1][119] ), .A4(\ram[3][119] ), .S0(n501), .S1(n408), .Y(n1084) );
  MUX41X1_HVT U1206 ( .A1(n1084), .A3(n1082), .A2(n1083), .A4(n1081), .S0(n589), .S1(n577), .Y(q[119]) );
  MUX41X1_HVT U1207 ( .A1(\ram[12][120] ), .A3(\ram[14][120] ), .A2(
        \ram[13][120] ), .A4(\ram[15][120] ), .S0(n502), .S1(n409), .Y(n1085)
         );
  MUX41X1_HVT U1208 ( .A1(\ram[8][120] ), .A3(\ram[10][120] ), .A2(
        \ram[9][120] ), .A4(\ram[11][120] ), .S0(n502), .S1(n409), .Y(n1086)
         );
  MUX41X1_HVT U1209 ( .A1(\ram[4][120] ), .A3(\ram[6][120] ), .A2(
        \ram[5][120] ), .A4(\ram[7][120] ), .S0(n502), .S1(n409), .Y(n1087) );
  MUX41X1_HVT U1210 ( .A1(\ram[0][120] ), .A3(\ram[2][120] ), .A2(
        \ram[1][120] ), .A4(\ram[3][120] ), .S0(n502), .S1(n409), .Y(n1088) );
  MUX41X1_HVT U1211 ( .A1(n1088), .A3(n1086), .A2(n1087), .A4(n1085), .S0(n590), .S1(n577), .Y(q[120]) );
  MUX41X1_HVT U1212 ( .A1(\ram[12][121] ), .A3(\ram[14][121] ), .A2(
        \ram[13][121] ), .A4(\ram[15][121] ), .S0(n502), .S1(n409), .Y(n1089)
         );
  MUX41X1_HVT U1213 ( .A1(\ram[8][121] ), .A3(\ram[10][121] ), .A2(
        \ram[9][121] ), .A4(\ram[11][121] ), .S0(n502), .S1(n409), .Y(n1090)
         );
  MUX41X1_HVT U1214 ( .A1(\ram[4][121] ), .A3(\ram[6][121] ), .A2(
        \ram[5][121] ), .A4(\ram[7][121] ), .S0(n502), .S1(n409), .Y(n1091) );
  MUX41X1_HVT U1215 ( .A1(\ram[0][121] ), .A3(\ram[2][121] ), .A2(
        \ram[1][121] ), .A4(\ram[3][121] ), .S0(n502), .S1(n409), .Y(n1092) );
  MUX41X1_HVT U1216 ( .A1(n1092), .A3(n1090), .A2(n1091), .A4(n1089), .S0(n590), .S1(n577), .Y(q[121]) );
  MUX41X1_HVT U1217 ( .A1(\ram[12][122] ), .A3(\ram[14][122] ), .A2(
        \ram[13][122] ), .A4(\ram[15][122] ), .S0(n502), .S1(n409), .Y(n1093)
         );
  MUX41X1_HVT U1218 ( .A1(\ram[8][122] ), .A3(\ram[10][122] ), .A2(
        \ram[9][122] ), .A4(\ram[11][122] ), .S0(n502), .S1(n409), .Y(n1094)
         );
  MUX41X1_HVT U1219 ( .A1(\ram[4][122] ), .A3(\ram[6][122] ), .A2(
        \ram[5][122] ), .A4(\ram[7][122] ), .S0(n502), .S1(n409), .Y(n1095) );
  MUX41X1_HVT U1220 ( .A1(\ram[0][122] ), .A3(\ram[2][122] ), .A2(
        \ram[1][122] ), .A4(\ram[3][122] ), .S0(n502), .S1(n409), .Y(n1096) );
  MUX41X1_HVT U1221 ( .A1(n1096), .A3(n1094), .A2(n1095), .A4(n1093), .S0(n590), .S1(n577), .Y(q[122]) );
  MUX41X1_HVT U1222 ( .A1(\ram[12][123] ), .A3(\ram[14][123] ), .A2(
        \ram[13][123] ), .A4(\ram[15][123] ), .S0(n503), .S1(n410), .Y(n1097)
         );
  MUX41X1_HVT U1223 ( .A1(\ram[8][123] ), .A3(\ram[10][123] ), .A2(
        \ram[9][123] ), .A4(\ram[11][123] ), .S0(n503), .S1(n410), .Y(n1098)
         );
  MUX41X1_HVT U1224 ( .A1(\ram[4][123] ), .A3(\ram[6][123] ), .A2(
        \ram[5][123] ), .A4(\ram[7][123] ), .S0(n503), .S1(n410), .Y(n1099) );
  MUX41X1_HVT U1225 ( .A1(\ram[0][123] ), .A3(\ram[2][123] ), .A2(
        \ram[1][123] ), .A4(\ram[3][123] ), .S0(n503), .S1(n410), .Y(n1100) );
  MUX41X1_HVT U1226 ( .A1(n1100), .A3(n1098), .A2(n1099), .A4(n1097), .S0(n590), .S1(N11), .Y(q[123]) );
  MUX41X1_HVT U1227 ( .A1(\ram[12][124] ), .A3(\ram[14][124] ), .A2(
        \ram[13][124] ), .A4(\ram[15][124] ), .S0(n503), .S1(n410), .Y(n1101)
         );
  MUX41X1_HVT U1228 ( .A1(\ram[8][124] ), .A3(\ram[10][124] ), .A2(
        \ram[9][124] ), .A4(\ram[11][124] ), .S0(n503), .S1(n410), .Y(n1102)
         );
  MUX41X1_HVT U1229 ( .A1(\ram[4][124] ), .A3(\ram[6][124] ), .A2(
        \ram[5][124] ), .A4(\ram[7][124] ), .S0(n503), .S1(n410), .Y(n1103) );
  MUX41X1_HVT U1230 ( .A1(\ram[0][124] ), .A3(\ram[2][124] ), .A2(
        \ram[1][124] ), .A4(\ram[3][124] ), .S0(n503), .S1(n410), .Y(n1104) );
  MUX41X1_HVT U1231 ( .A1(n1104), .A3(n1102), .A2(n1103), .A4(n1101), .S0(n590), .S1(n577), .Y(q[124]) );
  MUX41X1_HVT U1232 ( .A1(\ram[12][125] ), .A3(\ram[14][125] ), .A2(
        \ram[13][125] ), .A4(\ram[15][125] ), .S0(n503), .S1(n410), .Y(n1105)
         );
  MUX41X1_HVT U1233 ( .A1(\ram[8][125] ), .A3(\ram[10][125] ), .A2(
        \ram[9][125] ), .A4(\ram[11][125] ), .S0(n503), .S1(n410), .Y(n1106)
         );
  MUX41X1_HVT U1234 ( .A1(\ram[4][125] ), .A3(\ram[6][125] ), .A2(
        \ram[5][125] ), .A4(\ram[7][125] ), .S0(n503), .S1(n410), .Y(n1107) );
  MUX41X1_HVT U1235 ( .A1(\ram[0][125] ), .A3(\ram[2][125] ), .A2(
        \ram[1][125] ), .A4(\ram[3][125] ), .S0(n503), .S1(n410), .Y(n1108) );
  MUX41X1_HVT U1236 ( .A1(n1108), .A3(n1106), .A2(n1107), .A4(n1105), .S0(n590), .S1(N11), .Y(q[125]) );
  MUX41X1_HVT U1237 ( .A1(\ram[12][126] ), .A3(\ram[14][126] ), .A2(
        \ram[13][126] ), .A4(\ram[15][126] ), .S0(n504), .S1(n411), .Y(n1109)
         );
  MUX41X1_HVT U1238 ( .A1(\ram[8][126] ), .A3(\ram[10][126] ), .A2(
        \ram[9][126] ), .A4(\ram[11][126] ), .S0(n504), .S1(n411), .Y(n1110)
         );
  MUX41X1_HVT U1239 ( .A1(\ram[4][126] ), .A3(\ram[6][126] ), .A2(
        \ram[5][126] ), .A4(\ram[7][126] ), .S0(n504), .S1(n411), .Y(n1111) );
  MUX41X1_HVT U1240 ( .A1(\ram[0][126] ), .A3(\ram[2][126] ), .A2(
        \ram[1][126] ), .A4(\ram[3][126] ), .S0(n504), .S1(n411), .Y(n1112) );
  MUX41X1_HVT U1241 ( .A1(n1112), .A3(n1110), .A2(n1111), .A4(n1109), .S0(n590), .S1(N11), .Y(q[126]) );
  MUX41X1_HVT U1242 ( .A1(\ram[12][127] ), .A3(\ram[14][127] ), .A2(
        \ram[13][127] ), .A4(\ram[15][127] ), .S0(n504), .S1(n411), .Y(n1113)
         );
  MUX41X1_HVT U1243 ( .A1(\ram[8][127] ), .A3(\ram[10][127] ), .A2(
        \ram[9][127] ), .A4(\ram[11][127] ), .S0(n504), .S1(n411), .Y(n1114)
         );
  MUX41X1_HVT U1244 ( .A1(\ram[4][127] ), .A3(\ram[6][127] ), .A2(
        \ram[5][127] ), .A4(\ram[7][127] ), .S0(n504), .S1(n411), .Y(n1115) );
  MUX41X1_HVT U1245 ( .A1(\ram[0][127] ), .A3(\ram[2][127] ), .A2(
        \ram[1][127] ), .A4(\ram[3][127] ), .S0(n504), .S1(n411), .Y(n1116) );
  MUX41X1_HVT U1246 ( .A1(n1116), .A3(n1114), .A2(n1115), .A4(n1113), .S0(n590), .S1(N11), .Y(q[127]) );
  MUX41X1_HVT U1247 ( .A1(\ram[12][128] ), .A3(\ram[14][128] ), .A2(
        \ram[13][128] ), .A4(\ram[15][128] ), .S0(n504), .S1(n411), .Y(n1117)
         );
  MUX41X1_HVT U1248 ( .A1(\ram[8][128] ), .A3(\ram[10][128] ), .A2(
        \ram[9][128] ), .A4(\ram[11][128] ), .S0(n504), .S1(n411), .Y(n1118)
         );
  MUX41X1_HVT U1249 ( .A1(\ram[4][128] ), .A3(\ram[6][128] ), .A2(
        \ram[5][128] ), .A4(\ram[7][128] ), .S0(n504), .S1(n411), .Y(n1119) );
  MUX41X1_HVT U1250 ( .A1(\ram[0][128] ), .A3(\ram[2][128] ), .A2(
        \ram[1][128] ), .A4(\ram[3][128] ), .S0(n504), .S1(n411), .Y(n1120) );
  MUX41X1_HVT U1251 ( .A1(n1120), .A3(n1118), .A2(n1119), .A4(n1117), .S0(n590), .S1(n562), .Y(q[128]) );
  MUX41X1_HVT U1252 ( .A1(\ram[12][129] ), .A3(\ram[14][129] ), .A2(
        \ram[13][129] ), .A4(\ram[15][129] ), .S0(n505), .S1(n412), .Y(n1121)
         );
  MUX41X1_HVT U1253 ( .A1(\ram[8][129] ), .A3(\ram[10][129] ), .A2(
        \ram[9][129] ), .A4(\ram[11][129] ), .S0(n505), .S1(n412), .Y(n1122)
         );
  MUX41X1_HVT U1254 ( .A1(\ram[4][129] ), .A3(\ram[6][129] ), .A2(
        \ram[5][129] ), .A4(\ram[7][129] ), .S0(n505), .S1(n412), .Y(n1123) );
  MUX41X1_HVT U1255 ( .A1(\ram[0][129] ), .A3(\ram[2][129] ), .A2(
        \ram[1][129] ), .A4(\ram[3][129] ), .S0(n505), .S1(n412), .Y(n1124) );
  MUX41X1_HVT U1256 ( .A1(n1124), .A3(n1122), .A2(n1123), .A4(n1121), .S0(n590), .S1(n557), .Y(q[129]) );
  MUX41X1_HVT U1257 ( .A1(\ram[12][130] ), .A3(\ram[14][130] ), .A2(
        \ram[13][130] ), .A4(\ram[15][130] ), .S0(n505), .S1(n412), .Y(n1125)
         );
  MUX41X1_HVT U1258 ( .A1(\ram[8][130] ), .A3(\ram[10][130] ), .A2(
        \ram[9][130] ), .A4(\ram[11][130] ), .S0(n505), .S1(n412), .Y(n1126)
         );
  MUX41X1_HVT U1259 ( .A1(\ram[4][130] ), .A3(\ram[6][130] ), .A2(
        \ram[5][130] ), .A4(\ram[7][130] ), .S0(n505), .S1(n412), .Y(n1127) );
  MUX41X1_HVT U1260 ( .A1(\ram[0][130] ), .A3(\ram[2][130] ), .A2(
        \ram[1][130] ), .A4(\ram[3][130] ), .S0(n505), .S1(n412), .Y(n1128) );
  MUX41X1_HVT U1261 ( .A1(n1128), .A3(n1126), .A2(n1127), .A4(n1125), .S0(n590), .S1(n557), .Y(q[130]) );
  MUX41X1_HVT U1262 ( .A1(\ram[12][131] ), .A3(\ram[14][131] ), .A2(
        \ram[13][131] ), .A4(\ram[15][131] ), .S0(n505), .S1(n412), .Y(n1129)
         );
  MUX41X1_HVT U1263 ( .A1(\ram[8][131] ), .A3(\ram[10][131] ), .A2(
        \ram[9][131] ), .A4(\ram[11][131] ), .S0(n505), .S1(n412), .Y(n1130)
         );
  MUX41X1_HVT U1264 ( .A1(\ram[4][131] ), .A3(\ram[6][131] ), .A2(
        \ram[5][131] ), .A4(\ram[7][131] ), .S0(n505), .S1(n412), .Y(n1131) );
  MUX41X1_HVT U1265 ( .A1(\ram[0][131] ), .A3(\ram[2][131] ), .A2(
        \ram[1][131] ), .A4(\ram[3][131] ), .S0(n505), .S1(n412), .Y(n1132) );
  MUX41X1_HVT U1266 ( .A1(n1132), .A3(n1130), .A2(n1131), .A4(n1129), .S0(n590), .S1(n557), .Y(q[131]) );
  MUX41X1_HVT U1267 ( .A1(\ram[12][132] ), .A3(\ram[14][132] ), .A2(
        \ram[13][132] ), .A4(\ram[15][132] ), .S0(n506), .S1(n413), .Y(n1133)
         );
  MUX41X1_HVT U1268 ( .A1(\ram[8][132] ), .A3(\ram[10][132] ), .A2(
        \ram[9][132] ), .A4(\ram[11][132] ), .S0(n506), .S1(n413), .Y(n1134)
         );
  MUX41X1_HVT U1269 ( .A1(\ram[4][132] ), .A3(\ram[6][132] ), .A2(
        \ram[5][132] ), .A4(\ram[7][132] ), .S0(n506), .S1(n413), .Y(n1135) );
  MUX41X1_HVT U1270 ( .A1(\ram[0][132] ), .A3(\ram[2][132] ), .A2(
        \ram[1][132] ), .A4(\ram[3][132] ), .S0(n506), .S1(n413), .Y(n1136) );
  MUX41X1_HVT U1271 ( .A1(n1136), .A3(n1134), .A2(n1135), .A4(n1133), .S0(n591), .S1(n557), .Y(q[132]) );
  MUX41X1_HVT U1272 ( .A1(\ram[12][133] ), .A3(\ram[14][133] ), .A2(
        \ram[13][133] ), .A4(\ram[15][133] ), .S0(n506), .S1(n413), .Y(n1137)
         );
  MUX41X1_HVT U1273 ( .A1(\ram[8][133] ), .A3(\ram[10][133] ), .A2(
        \ram[9][133] ), .A4(\ram[11][133] ), .S0(n506), .S1(n413), .Y(n1138)
         );
  MUX41X1_HVT U1274 ( .A1(\ram[4][133] ), .A3(\ram[6][133] ), .A2(
        \ram[5][133] ), .A4(\ram[7][133] ), .S0(n506), .S1(n413), .Y(n1139) );
  MUX41X1_HVT U1275 ( .A1(\ram[0][133] ), .A3(\ram[2][133] ), .A2(
        \ram[1][133] ), .A4(\ram[3][133] ), .S0(n506), .S1(n413), .Y(n1140) );
  MUX41X1_HVT U1276 ( .A1(n1140), .A3(n1138), .A2(n1139), .A4(n1137), .S0(n591), .S1(n557), .Y(q[133]) );
  MUX41X1_HVT U1277 ( .A1(\ram[12][134] ), .A3(\ram[14][134] ), .A2(
        \ram[13][134] ), .A4(\ram[15][134] ), .S0(n506), .S1(n413), .Y(n1141)
         );
  MUX41X1_HVT U1278 ( .A1(\ram[8][134] ), .A3(\ram[10][134] ), .A2(
        \ram[9][134] ), .A4(\ram[11][134] ), .S0(n506), .S1(n413), .Y(n1142)
         );
  MUX41X1_HVT U1279 ( .A1(\ram[4][134] ), .A3(\ram[6][134] ), .A2(
        \ram[5][134] ), .A4(\ram[7][134] ), .S0(n506), .S1(n413), .Y(n1143) );
  MUX41X1_HVT U1280 ( .A1(\ram[0][134] ), .A3(\ram[2][134] ), .A2(
        \ram[1][134] ), .A4(\ram[3][134] ), .S0(n506), .S1(n413), .Y(n1144) );
  MUX41X1_HVT U1281 ( .A1(n1144), .A3(n1142), .A2(n1143), .A4(n1141), .S0(n591), .S1(n557), .Y(q[134]) );
  MUX41X1_HVT U1282 ( .A1(\ram[12][135] ), .A3(\ram[14][135] ), .A2(
        \ram[13][135] ), .A4(\ram[15][135] ), .S0(n507), .S1(n414), .Y(n1145)
         );
  MUX41X1_HVT U1283 ( .A1(\ram[8][135] ), .A3(\ram[10][135] ), .A2(
        \ram[9][135] ), .A4(\ram[11][135] ), .S0(n507), .S1(n414), .Y(n1146)
         );
  MUX41X1_HVT U1284 ( .A1(\ram[4][135] ), .A3(\ram[6][135] ), .A2(
        \ram[5][135] ), .A4(\ram[7][135] ), .S0(n507), .S1(n414), .Y(n1147) );
  MUX41X1_HVT U1285 ( .A1(\ram[0][135] ), .A3(\ram[2][135] ), .A2(
        \ram[1][135] ), .A4(\ram[3][135] ), .S0(n507), .S1(n414), .Y(n1148) );
  MUX41X1_HVT U1286 ( .A1(n1148), .A3(n1146), .A2(n1147), .A4(n1145), .S0(n591), .S1(n557), .Y(q[135]) );
  MUX41X1_HVT U1287 ( .A1(\ram[12][136] ), .A3(\ram[14][136] ), .A2(
        \ram[13][136] ), .A4(\ram[15][136] ), .S0(n507), .S1(n414), .Y(n1149)
         );
  MUX41X1_HVT U1288 ( .A1(\ram[8][136] ), .A3(\ram[10][136] ), .A2(
        \ram[9][136] ), .A4(\ram[11][136] ), .S0(n507), .S1(n414), .Y(n1150)
         );
  MUX41X1_HVT U1289 ( .A1(\ram[4][136] ), .A3(\ram[6][136] ), .A2(
        \ram[5][136] ), .A4(\ram[7][136] ), .S0(n507), .S1(n414), .Y(n1151) );
  MUX41X1_HVT U1290 ( .A1(\ram[0][136] ), .A3(\ram[2][136] ), .A2(
        \ram[1][136] ), .A4(\ram[3][136] ), .S0(n507), .S1(n414), .Y(n1152) );
  MUX41X1_HVT U1291 ( .A1(n1152), .A3(n1150), .A2(n1151), .A4(n1149), .S0(n591), .S1(n557), .Y(q[136]) );
  MUX41X1_HVT U1292 ( .A1(\ram[12][137] ), .A3(\ram[14][137] ), .A2(
        \ram[13][137] ), .A4(\ram[15][137] ), .S0(n507), .S1(n414), .Y(n1153)
         );
  MUX41X1_HVT U1293 ( .A1(\ram[8][137] ), .A3(\ram[10][137] ), .A2(
        \ram[9][137] ), .A4(\ram[11][137] ), .S0(n507), .S1(n414), .Y(n1154)
         );
  MUX41X1_HVT U1294 ( .A1(\ram[4][137] ), .A3(\ram[6][137] ), .A2(
        \ram[5][137] ), .A4(\ram[7][137] ), .S0(n507), .S1(n414), .Y(n1155) );
  MUX41X1_HVT U1295 ( .A1(\ram[0][137] ), .A3(\ram[2][137] ), .A2(
        \ram[1][137] ), .A4(\ram[3][137] ), .S0(n507), .S1(n414), .Y(n1156) );
  MUX41X1_HVT U1296 ( .A1(n1156), .A3(n1154), .A2(n1155), .A4(n1153), .S0(n591), .S1(n557), .Y(q[137]) );
  MUX41X1_HVT U1297 ( .A1(\ram[12][138] ), .A3(\ram[14][138] ), .A2(
        \ram[13][138] ), .A4(\ram[15][138] ), .S0(n508), .S1(n415), .Y(n1157)
         );
  MUX41X1_HVT U1298 ( .A1(\ram[8][138] ), .A3(\ram[10][138] ), .A2(
        \ram[9][138] ), .A4(\ram[11][138] ), .S0(n508), .S1(n415), .Y(n1158)
         );
  MUX41X1_HVT U1299 ( .A1(\ram[4][138] ), .A3(\ram[6][138] ), .A2(
        \ram[5][138] ), .A4(\ram[7][138] ), .S0(n508), .S1(n415), .Y(n1159) );
  MUX41X1_HVT U1300 ( .A1(\ram[0][138] ), .A3(\ram[2][138] ), .A2(
        \ram[1][138] ), .A4(\ram[3][138] ), .S0(n508), .S1(n415), .Y(n1160) );
  MUX41X1_HVT U1301 ( .A1(n1160), .A3(n1158), .A2(n1159), .A4(n1157), .S0(n591), .S1(n557), .Y(q[138]) );
  MUX41X1_HVT U1302 ( .A1(\ram[12][139] ), .A3(\ram[14][139] ), .A2(
        \ram[13][139] ), .A4(\ram[15][139] ), .S0(n508), .S1(n415), .Y(n1161)
         );
  MUX41X1_HVT U1303 ( .A1(\ram[8][139] ), .A3(\ram[10][139] ), .A2(
        \ram[9][139] ), .A4(\ram[11][139] ), .S0(n508), .S1(n415), .Y(n1162)
         );
  MUX41X1_HVT U1304 ( .A1(\ram[4][139] ), .A3(\ram[6][139] ), .A2(
        \ram[5][139] ), .A4(\ram[7][139] ), .S0(n508), .S1(n415), .Y(n1163) );
  MUX41X1_HVT U1305 ( .A1(\ram[0][139] ), .A3(\ram[2][139] ), .A2(
        \ram[1][139] ), .A4(\ram[3][139] ), .S0(n508), .S1(n415), .Y(n1164) );
  MUX41X1_HVT U1306 ( .A1(n1164), .A3(n1162), .A2(n1163), .A4(n1161), .S0(n591), .S1(n557), .Y(q[139]) );
  MUX41X1_HVT U1307 ( .A1(\ram[12][140] ), .A3(\ram[14][140] ), .A2(
        \ram[13][140] ), .A4(\ram[15][140] ), .S0(n508), .S1(n415), .Y(n1165)
         );
  MUX41X1_HVT U1308 ( .A1(\ram[8][140] ), .A3(\ram[10][140] ), .A2(
        \ram[9][140] ), .A4(\ram[11][140] ), .S0(n508), .S1(n415), .Y(n1166)
         );
  MUX41X1_HVT U1309 ( .A1(\ram[4][140] ), .A3(\ram[6][140] ), .A2(
        \ram[5][140] ), .A4(\ram[7][140] ), .S0(n508), .S1(n415), .Y(n1167) );
  MUX41X1_HVT U1310 ( .A1(\ram[0][140] ), .A3(\ram[2][140] ), .A2(
        \ram[1][140] ), .A4(\ram[3][140] ), .S0(n508), .S1(n415), .Y(n1168) );
  MUX41X1_HVT U1311 ( .A1(n1168), .A3(n1166), .A2(n1167), .A4(n1165), .S0(n591), .S1(n558), .Y(q[140]) );
  MUX41X1_HVT U1312 ( .A1(\ram[12][141] ), .A3(\ram[14][141] ), .A2(
        \ram[13][141] ), .A4(\ram[15][141] ), .S0(n509), .S1(n416), .Y(n1169)
         );
  MUX41X1_HVT U1313 ( .A1(\ram[8][141] ), .A3(\ram[10][141] ), .A2(
        \ram[9][141] ), .A4(\ram[11][141] ), .S0(n509), .S1(n416), .Y(n1170)
         );
  MUX41X1_HVT U1314 ( .A1(\ram[4][141] ), .A3(\ram[6][141] ), .A2(
        \ram[5][141] ), .A4(\ram[7][141] ), .S0(n509), .S1(n416), .Y(n1171) );
  MUX41X1_HVT U1315 ( .A1(\ram[0][141] ), .A3(\ram[2][141] ), .A2(
        \ram[1][141] ), .A4(\ram[3][141] ), .S0(n509), .S1(n416), .Y(n1172) );
  MUX41X1_HVT U1316 ( .A1(n1172), .A3(n1170), .A2(n1171), .A4(n1169), .S0(n591), .S1(n558), .Y(q[141]) );
  MUX41X1_HVT U1317 ( .A1(\ram[12][142] ), .A3(\ram[14][142] ), .A2(
        \ram[13][142] ), .A4(\ram[15][142] ), .S0(n509), .S1(n416), .Y(n1173)
         );
  MUX41X1_HVT U1318 ( .A1(\ram[8][142] ), .A3(\ram[10][142] ), .A2(
        \ram[9][142] ), .A4(\ram[11][142] ), .S0(n509), .S1(n416), .Y(n1174)
         );
  MUX41X1_HVT U1319 ( .A1(\ram[4][142] ), .A3(\ram[6][142] ), .A2(
        \ram[5][142] ), .A4(\ram[7][142] ), .S0(n509), .S1(n416), .Y(n1175) );
  MUX41X1_HVT U1320 ( .A1(\ram[0][142] ), .A3(\ram[2][142] ), .A2(
        \ram[1][142] ), .A4(\ram[3][142] ), .S0(n509), .S1(n416), .Y(n1176) );
  MUX41X1_HVT U1321 ( .A1(n1176), .A3(n1174), .A2(n1175), .A4(n1173), .S0(n591), .S1(n558), .Y(q[142]) );
  MUX41X1_HVT U1322 ( .A1(\ram[12][143] ), .A3(\ram[14][143] ), .A2(
        \ram[13][143] ), .A4(\ram[15][143] ), .S0(n509), .S1(n416), .Y(n1177)
         );
  MUX41X1_HVT U1323 ( .A1(\ram[8][143] ), .A3(\ram[10][143] ), .A2(
        \ram[9][143] ), .A4(\ram[11][143] ), .S0(n509), .S1(n416), .Y(n1178)
         );
  MUX41X1_HVT U1324 ( .A1(\ram[4][143] ), .A3(\ram[6][143] ), .A2(
        \ram[5][143] ), .A4(\ram[7][143] ), .S0(n509), .S1(n416), .Y(n1179) );
  MUX41X1_HVT U1325 ( .A1(\ram[0][143] ), .A3(\ram[2][143] ), .A2(
        \ram[1][143] ), .A4(\ram[3][143] ), .S0(n509), .S1(n416), .Y(n1180) );
  MUX41X1_HVT U1326 ( .A1(n1180), .A3(n1178), .A2(n1179), .A4(n1177), .S0(n591), .S1(n558), .Y(q[143]) );
  MUX41X1_HVT U1327 ( .A1(\ram[12][144] ), .A3(\ram[14][144] ), .A2(
        \ram[13][144] ), .A4(\ram[15][144] ), .S0(n510), .S1(n417), .Y(n1181)
         );
  MUX41X1_HVT U1328 ( .A1(\ram[8][144] ), .A3(\ram[10][144] ), .A2(
        \ram[9][144] ), .A4(\ram[11][144] ), .S0(n510), .S1(n417), .Y(n1182)
         );
  MUX41X1_HVT U1329 ( .A1(\ram[4][144] ), .A3(\ram[6][144] ), .A2(
        \ram[5][144] ), .A4(\ram[7][144] ), .S0(n510), .S1(n417), .Y(n1183) );
  MUX41X1_HVT U1330 ( .A1(\ram[0][144] ), .A3(\ram[2][144] ), .A2(
        \ram[1][144] ), .A4(\ram[3][144] ), .S0(n510), .S1(n417), .Y(n1184) );
  MUX41X1_HVT U1331 ( .A1(n1184), .A3(n1182), .A2(n1183), .A4(n1181), .S0(n592), .S1(n558), .Y(q[144]) );
  MUX41X1_HVT U1332 ( .A1(\ram[12][145] ), .A3(\ram[14][145] ), .A2(
        \ram[13][145] ), .A4(\ram[15][145] ), .S0(n510), .S1(n417), .Y(n1185)
         );
  MUX41X1_HVT U1333 ( .A1(\ram[8][145] ), .A3(\ram[10][145] ), .A2(
        \ram[9][145] ), .A4(\ram[11][145] ), .S0(n510), .S1(n417), .Y(n1186)
         );
  MUX41X1_HVT U1334 ( .A1(\ram[4][145] ), .A3(\ram[6][145] ), .A2(
        \ram[5][145] ), .A4(\ram[7][145] ), .S0(n510), .S1(n417), .Y(n1187) );
  MUX41X1_HVT U1335 ( .A1(\ram[0][145] ), .A3(\ram[2][145] ), .A2(
        \ram[1][145] ), .A4(\ram[3][145] ), .S0(n510), .S1(n417), .Y(n1188) );
  MUX41X1_HVT U1336 ( .A1(n1188), .A3(n1186), .A2(n1187), .A4(n1185), .S0(n592), .S1(n558), .Y(q[145]) );
  MUX41X1_HVT U1337 ( .A1(\ram[12][146] ), .A3(\ram[14][146] ), .A2(
        \ram[13][146] ), .A4(\ram[15][146] ), .S0(n510), .S1(n417), .Y(n1189)
         );
  MUX41X1_HVT U1338 ( .A1(\ram[8][146] ), .A3(\ram[10][146] ), .A2(
        \ram[9][146] ), .A4(\ram[11][146] ), .S0(n510), .S1(n417), .Y(n1190)
         );
  MUX41X1_HVT U1339 ( .A1(\ram[4][146] ), .A3(\ram[6][146] ), .A2(
        \ram[5][146] ), .A4(\ram[7][146] ), .S0(n510), .S1(n417), .Y(n1191) );
  MUX41X1_HVT U1340 ( .A1(\ram[0][146] ), .A3(\ram[2][146] ), .A2(
        \ram[1][146] ), .A4(\ram[3][146] ), .S0(n510), .S1(n417), .Y(n1192) );
  MUX41X1_HVT U1341 ( .A1(n1192), .A3(n1190), .A2(n1191), .A4(n1189), .S0(n592), .S1(n558), .Y(q[146]) );
  MUX41X1_HVT U1342 ( .A1(\ram[12][147] ), .A3(\ram[14][147] ), .A2(
        \ram[13][147] ), .A4(\ram[15][147] ), .S0(n511), .S1(n418), .Y(n1193)
         );
  MUX41X1_HVT U1343 ( .A1(\ram[8][147] ), .A3(\ram[10][147] ), .A2(
        \ram[9][147] ), .A4(\ram[11][147] ), .S0(n511), .S1(n418), .Y(n1194)
         );
  MUX41X1_HVT U1344 ( .A1(\ram[4][147] ), .A3(\ram[6][147] ), .A2(
        \ram[5][147] ), .A4(\ram[7][147] ), .S0(n511), .S1(n418), .Y(n1195) );
  MUX41X1_HVT U1345 ( .A1(\ram[0][147] ), .A3(\ram[2][147] ), .A2(
        \ram[1][147] ), .A4(\ram[3][147] ), .S0(n511), .S1(n418), .Y(n1196) );
  MUX41X1_HVT U1346 ( .A1(n1196), .A3(n1194), .A2(n1195), .A4(n1193), .S0(n592), .S1(n558), .Y(q[147]) );
  MUX41X1_HVT U1347 ( .A1(\ram[12][148] ), .A3(\ram[14][148] ), .A2(
        \ram[13][148] ), .A4(\ram[15][148] ), .S0(n511), .S1(n418), .Y(n1197)
         );
  MUX41X1_HVT U1348 ( .A1(\ram[8][148] ), .A3(\ram[10][148] ), .A2(
        \ram[9][148] ), .A4(\ram[11][148] ), .S0(n511), .S1(n418), .Y(n1198)
         );
  MUX41X1_HVT U1349 ( .A1(\ram[4][148] ), .A3(\ram[6][148] ), .A2(
        \ram[5][148] ), .A4(\ram[7][148] ), .S0(n511), .S1(n418), .Y(n1199) );
  MUX41X1_HVT U1350 ( .A1(\ram[0][148] ), .A3(\ram[2][148] ), .A2(
        \ram[1][148] ), .A4(\ram[3][148] ), .S0(n511), .S1(n418), .Y(n1200) );
  MUX41X1_HVT U1351 ( .A1(n1200), .A3(n1198), .A2(n1199), .A4(n1197), .S0(n592), .S1(n558), .Y(q[148]) );
  MUX41X1_HVT U1352 ( .A1(\ram[12][149] ), .A3(\ram[14][149] ), .A2(
        \ram[13][149] ), .A4(\ram[15][149] ), .S0(n511), .S1(n418), .Y(n1201)
         );
  MUX41X1_HVT U1353 ( .A1(\ram[8][149] ), .A3(\ram[10][149] ), .A2(
        \ram[9][149] ), .A4(\ram[11][149] ), .S0(n511), .S1(n418), .Y(n1202)
         );
  MUX41X1_HVT U1354 ( .A1(\ram[4][149] ), .A3(\ram[6][149] ), .A2(
        \ram[5][149] ), .A4(\ram[7][149] ), .S0(n511), .S1(n418), .Y(n1203) );
  MUX41X1_HVT U1355 ( .A1(\ram[0][149] ), .A3(\ram[2][149] ), .A2(
        \ram[1][149] ), .A4(\ram[3][149] ), .S0(n511), .S1(n418), .Y(n1204) );
  MUX41X1_HVT U1356 ( .A1(n1204), .A3(n1202), .A2(n1203), .A4(n1201), .S0(n592), .S1(n558), .Y(q[149]) );
  MUX41X1_HVT U1357 ( .A1(\ram[12][150] ), .A3(\ram[14][150] ), .A2(
        \ram[13][150] ), .A4(\ram[15][150] ), .S0(n512), .S1(n419), .Y(n1205)
         );
  MUX41X1_HVT U1358 ( .A1(\ram[8][150] ), .A3(\ram[10][150] ), .A2(
        \ram[9][150] ), .A4(\ram[11][150] ), .S0(n512), .S1(n419), .Y(n1206)
         );
  MUX41X1_HVT U1359 ( .A1(\ram[4][150] ), .A3(\ram[6][150] ), .A2(
        \ram[5][150] ), .A4(\ram[7][150] ), .S0(n512), .S1(n419), .Y(n1207) );
  MUX41X1_HVT U1360 ( .A1(\ram[0][150] ), .A3(\ram[2][150] ), .A2(
        \ram[1][150] ), .A4(\ram[3][150] ), .S0(n512), .S1(n419), .Y(n1208) );
  MUX41X1_HVT U1361 ( .A1(n1208), .A3(n1206), .A2(n1207), .A4(n1205), .S0(n592), .S1(n558), .Y(q[150]) );
  MUX41X1_HVT U1362 ( .A1(\ram[12][151] ), .A3(\ram[14][151] ), .A2(
        \ram[13][151] ), .A4(\ram[15][151] ), .S0(n512), .S1(n419), .Y(n1209)
         );
  MUX41X1_HVT U1363 ( .A1(\ram[8][151] ), .A3(\ram[10][151] ), .A2(
        \ram[9][151] ), .A4(\ram[11][151] ), .S0(n512), .S1(n419), .Y(n1210)
         );
  MUX41X1_HVT U1364 ( .A1(\ram[4][151] ), .A3(\ram[6][151] ), .A2(
        \ram[5][151] ), .A4(\ram[7][151] ), .S0(n512), .S1(n419), .Y(n1211) );
  MUX41X1_HVT U1365 ( .A1(\ram[0][151] ), .A3(\ram[2][151] ), .A2(
        \ram[1][151] ), .A4(\ram[3][151] ), .S0(n512), .S1(n419), .Y(n1212) );
  MUX41X1_HVT U1366 ( .A1(n1212), .A3(n1210), .A2(n1211), .A4(n1209), .S0(n592), .S1(n558), .Y(q[151]) );
  MUX41X1_HVT U1367 ( .A1(\ram[12][152] ), .A3(\ram[14][152] ), .A2(
        \ram[13][152] ), .A4(\ram[15][152] ), .S0(n512), .S1(n419), .Y(n1213)
         );
  MUX41X1_HVT U1368 ( .A1(\ram[8][152] ), .A3(\ram[10][152] ), .A2(
        \ram[9][152] ), .A4(\ram[11][152] ), .S0(n512), .S1(n419), .Y(n1214)
         );
  MUX41X1_HVT U1369 ( .A1(\ram[4][152] ), .A3(\ram[6][152] ), .A2(
        \ram[5][152] ), .A4(\ram[7][152] ), .S0(n512), .S1(n419), .Y(n1215) );
  MUX41X1_HVT U1370 ( .A1(\ram[0][152] ), .A3(\ram[2][152] ), .A2(
        \ram[1][152] ), .A4(\ram[3][152] ), .S0(n512), .S1(n419), .Y(n1216) );
  MUX41X1_HVT U1371 ( .A1(n1216), .A3(n1214), .A2(n1215), .A4(n1213), .S0(n592), .S1(n559), .Y(q[152]) );
  MUX41X1_HVT U1372 ( .A1(\ram[12][153] ), .A3(\ram[14][153] ), .A2(
        \ram[13][153] ), .A4(\ram[15][153] ), .S0(n513), .S1(n420), .Y(n1217)
         );
  MUX41X1_HVT U1373 ( .A1(\ram[8][153] ), .A3(\ram[10][153] ), .A2(
        \ram[9][153] ), .A4(\ram[11][153] ), .S0(n513), .S1(n420), .Y(n1218)
         );
  MUX41X1_HVT U1374 ( .A1(\ram[4][153] ), .A3(\ram[6][153] ), .A2(
        \ram[5][153] ), .A4(\ram[7][153] ), .S0(n513), .S1(n420), .Y(n1219) );
  MUX41X1_HVT U1375 ( .A1(\ram[0][153] ), .A3(\ram[2][153] ), .A2(
        \ram[1][153] ), .A4(\ram[3][153] ), .S0(n513), .S1(n420), .Y(n1220) );
  MUX41X1_HVT U1376 ( .A1(n1220), .A3(n1218), .A2(n1219), .A4(n1217), .S0(n592), .S1(n559), .Y(q[153]) );
  MUX41X1_HVT U1377 ( .A1(\ram[12][154] ), .A3(\ram[14][154] ), .A2(
        \ram[13][154] ), .A4(\ram[15][154] ), .S0(n513), .S1(n420), .Y(n1221)
         );
  MUX41X1_HVT U1378 ( .A1(\ram[8][154] ), .A3(\ram[10][154] ), .A2(
        \ram[9][154] ), .A4(\ram[11][154] ), .S0(n513), .S1(n420), .Y(n1222)
         );
  MUX41X1_HVT U1379 ( .A1(\ram[4][154] ), .A3(\ram[6][154] ), .A2(
        \ram[5][154] ), .A4(\ram[7][154] ), .S0(n513), .S1(n420), .Y(n1223) );
  MUX41X1_HVT U1380 ( .A1(\ram[0][154] ), .A3(\ram[2][154] ), .A2(
        \ram[1][154] ), .A4(\ram[3][154] ), .S0(n513), .S1(n420), .Y(n1224) );
  MUX41X1_HVT U1381 ( .A1(n1224), .A3(n1222), .A2(n1223), .A4(n1221), .S0(n592), .S1(n559), .Y(q[154]) );
  MUX41X1_HVT U1382 ( .A1(\ram[12][155] ), .A3(\ram[14][155] ), .A2(
        \ram[13][155] ), .A4(\ram[15][155] ), .S0(n513), .S1(n420), .Y(n1225)
         );
  MUX41X1_HVT U1383 ( .A1(\ram[8][155] ), .A3(\ram[10][155] ), .A2(
        \ram[9][155] ), .A4(\ram[11][155] ), .S0(n513), .S1(n420), .Y(n1226)
         );
  MUX41X1_HVT U1384 ( .A1(\ram[4][155] ), .A3(\ram[6][155] ), .A2(
        \ram[5][155] ), .A4(\ram[7][155] ), .S0(n513), .S1(n420), .Y(n1227) );
  MUX41X1_HVT U1385 ( .A1(\ram[0][155] ), .A3(\ram[2][155] ), .A2(
        \ram[1][155] ), .A4(\ram[3][155] ), .S0(n513), .S1(n420), .Y(n1228) );
  MUX41X1_HVT U1386 ( .A1(n1228), .A3(n1226), .A2(n1227), .A4(n1225), .S0(n592), .S1(n559), .Y(q[155]) );
  MUX41X1_HVT U1387 ( .A1(\ram[12][156] ), .A3(\ram[14][156] ), .A2(
        \ram[13][156] ), .A4(\ram[15][156] ), .S0(n514), .S1(n421), .Y(n1229)
         );
  MUX41X1_HVT U1388 ( .A1(\ram[8][156] ), .A3(\ram[10][156] ), .A2(
        \ram[9][156] ), .A4(\ram[11][156] ), .S0(n514), .S1(n421), .Y(n1230)
         );
  MUX41X1_HVT U1389 ( .A1(\ram[4][156] ), .A3(\ram[6][156] ), .A2(
        \ram[5][156] ), .A4(\ram[7][156] ), .S0(n514), .S1(n421), .Y(n1231) );
  MUX41X1_HVT U1390 ( .A1(\ram[0][156] ), .A3(\ram[2][156] ), .A2(
        \ram[1][156] ), .A4(\ram[3][156] ), .S0(n514), .S1(n421), .Y(n1232) );
  MUX41X1_HVT U1391 ( .A1(n1232), .A3(n1230), .A2(n1231), .A4(n1229), .S0(n593), .S1(n559), .Y(q[156]) );
  MUX41X1_HVT U1392 ( .A1(\ram[12][157] ), .A3(\ram[14][157] ), .A2(
        \ram[13][157] ), .A4(\ram[15][157] ), .S0(n514), .S1(n421), .Y(n1233)
         );
  MUX41X1_HVT U1393 ( .A1(\ram[8][157] ), .A3(\ram[10][157] ), .A2(
        \ram[9][157] ), .A4(\ram[11][157] ), .S0(n514), .S1(n421), .Y(n1234)
         );
  MUX41X1_HVT U1394 ( .A1(\ram[4][157] ), .A3(\ram[6][157] ), .A2(
        \ram[5][157] ), .A4(\ram[7][157] ), .S0(n514), .S1(n421), .Y(n1235) );
  MUX41X1_HVT U1395 ( .A1(\ram[0][157] ), .A3(\ram[2][157] ), .A2(
        \ram[1][157] ), .A4(\ram[3][157] ), .S0(n514), .S1(n421), .Y(n1236) );
  MUX41X1_HVT U1396 ( .A1(n1236), .A3(n1234), .A2(n1235), .A4(n1233), .S0(n593), .S1(n559), .Y(q[157]) );
  MUX41X1_HVT U1397 ( .A1(\ram[12][158] ), .A3(\ram[14][158] ), .A2(
        \ram[13][158] ), .A4(\ram[15][158] ), .S0(n514), .S1(n421), .Y(n1237)
         );
  MUX41X1_HVT U1398 ( .A1(\ram[8][158] ), .A3(\ram[10][158] ), .A2(
        \ram[9][158] ), .A4(\ram[11][158] ), .S0(n514), .S1(n421), .Y(n1238)
         );
  MUX41X1_HVT U1399 ( .A1(\ram[4][158] ), .A3(\ram[6][158] ), .A2(
        \ram[5][158] ), .A4(\ram[7][158] ), .S0(n514), .S1(n421), .Y(n1239) );
  MUX41X1_HVT U1400 ( .A1(\ram[0][158] ), .A3(\ram[2][158] ), .A2(
        \ram[1][158] ), .A4(\ram[3][158] ), .S0(n514), .S1(n421), .Y(n1240) );
  MUX41X1_HVT U1401 ( .A1(n1240), .A3(n1238), .A2(n1239), .A4(n1237), .S0(n593), .S1(n559), .Y(q[158]) );
  MUX41X1_HVT U1402 ( .A1(\ram[12][159] ), .A3(\ram[14][159] ), .A2(
        \ram[13][159] ), .A4(\ram[15][159] ), .S0(n515), .S1(n422), .Y(n1241)
         );
  MUX41X1_HVT U1403 ( .A1(\ram[8][159] ), .A3(\ram[10][159] ), .A2(
        \ram[9][159] ), .A4(\ram[11][159] ), .S0(n515), .S1(n422), .Y(n1242)
         );
  MUX41X1_HVT U1404 ( .A1(\ram[4][159] ), .A3(\ram[6][159] ), .A2(
        \ram[5][159] ), .A4(\ram[7][159] ), .S0(n515), .S1(n422), .Y(n1243) );
  MUX41X1_HVT U1405 ( .A1(\ram[0][159] ), .A3(\ram[2][159] ), .A2(
        \ram[1][159] ), .A4(\ram[3][159] ), .S0(n515), .S1(n422), .Y(n1244) );
  MUX41X1_HVT U1406 ( .A1(n1244), .A3(n1242), .A2(n1243), .A4(n1241), .S0(n593), .S1(n559), .Y(q[159]) );
  MUX41X1_HVT U1407 ( .A1(\ram[12][160] ), .A3(\ram[14][160] ), .A2(
        \ram[13][160] ), .A4(\ram[15][160] ), .S0(n515), .S1(n422), .Y(n1245)
         );
  MUX41X1_HVT U1408 ( .A1(\ram[8][160] ), .A3(\ram[10][160] ), .A2(
        \ram[9][160] ), .A4(\ram[11][160] ), .S0(n515), .S1(n422), .Y(n1246)
         );
  MUX41X1_HVT U1409 ( .A1(\ram[4][160] ), .A3(\ram[6][160] ), .A2(
        \ram[5][160] ), .A4(\ram[7][160] ), .S0(n515), .S1(n422), .Y(n1247) );
  MUX41X1_HVT U1410 ( .A1(\ram[0][160] ), .A3(\ram[2][160] ), .A2(
        \ram[1][160] ), .A4(\ram[3][160] ), .S0(n515), .S1(n422), .Y(n1248) );
  MUX41X1_HVT U1411 ( .A1(n1248), .A3(n1246), .A2(n1247), .A4(n1245), .S0(n593), .S1(n559), .Y(q[160]) );
  MUX41X1_HVT U1412 ( .A1(\ram[12][161] ), .A3(\ram[14][161] ), .A2(
        \ram[13][161] ), .A4(\ram[15][161] ), .S0(n515), .S1(n422), .Y(n1249)
         );
  MUX41X1_HVT U1413 ( .A1(\ram[8][161] ), .A3(\ram[10][161] ), .A2(
        \ram[9][161] ), .A4(\ram[11][161] ), .S0(n515), .S1(n422), .Y(n1250)
         );
  MUX41X1_HVT U1414 ( .A1(\ram[4][161] ), .A3(\ram[6][161] ), .A2(
        \ram[5][161] ), .A4(\ram[7][161] ), .S0(n515), .S1(n422), .Y(n1251) );
  MUX41X1_HVT U1415 ( .A1(\ram[0][161] ), .A3(\ram[2][161] ), .A2(
        \ram[1][161] ), .A4(\ram[3][161] ), .S0(n515), .S1(n422), .Y(n1252) );
  MUX41X1_HVT U1416 ( .A1(n1252), .A3(n1250), .A2(n1251), .A4(n1249), .S0(n593), .S1(n559), .Y(q[161]) );
  MUX41X1_HVT U1417 ( .A1(\ram[12][162] ), .A3(\ram[14][162] ), .A2(
        \ram[13][162] ), .A4(\ram[15][162] ), .S0(n516), .S1(n423), .Y(n1253)
         );
  MUX41X1_HVT U1418 ( .A1(\ram[8][162] ), .A3(\ram[10][162] ), .A2(
        \ram[9][162] ), .A4(\ram[11][162] ), .S0(n516), .S1(n423), .Y(n1254)
         );
  MUX41X1_HVT U1419 ( .A1(\ram[4][162] ), .A3(\ram[6][162] ), .A2(
        \ram[5][162] ), .A4(\ram[7][162] ), .S0(n516), .S1(n423), .Y(n1255) );
  MUX41X1_HVT U1420 ( .A1(\ram[0][162] ), .A3(\ram[2][162] ), .A2(
        \ram[1][162] ), .A4(\ram[3][162] ), .S0(n516), .S1(n423), .Y(n1256) );
  MUX41X1_HVT U1421 ( .A1(n1256), .A3(n1254), .A2(n1255), .A4(n1253), .S0(n593), .S1(n559), .Y(q[162]) );
  MUX41X1_HVT U1422 ( .A1(\ram[12][163] ), .A3(\ram[14][163] ), .A2(
        \ram[13][163] ), .A4(\ram[15][163] ), .S0(n516), .S1(n423), .Y(n1257)
         );
  MUX41X1_HVT U1423 ( .A1(\ram[8][163] ), .A3(\ram[10][163] ), .A2(
        \ram[9][163] ), .A4(\ram[11][163] ), .S0(n516), .S1(n423), .Y(n1258)
         );
  MUX41X1_HVT U1424 ( .A1(\ram[4][163] ), .A3(\ram[6][163] ), .A2(
        \ram[5][163] ), .A4(\ram[7][163] ), .S0(n516), .S1(n423), .Y(n1259) );
  MUX41X1_HVT U1425 ( .A1(\ram[0][163] ), .A3(\ram[2][163] ), .A2(
        \ram[1][163] ), .A4(\ram[3][163] ), .S0(n516), .S1(n423), .Y(n1260) );
  MUX41X1_HVT U1426 ( .A1(n1260), .A3(n1258), .A2(n1259), .A4(n1257), .S0(n593), .S1(n559), .Y(q[163]) );
  MUX41X1_HVT U1427 ( .A1(\ram[12][164] ), .A3(\ram[14][164] ), .A2(
        \ram[13][164] ), .A4(\ram[15][164] ), .S0(n516), .S1(n423), .Y(n1261)
         );
  MUX41X1_HVT U1428 ( .A1(\ram[8][164] ), .A3(\ram[10][164] ), .A2(
        \ram[9][164] ), .A4(\ram[11][164] ), .S0(n516), .S1(n423), .Y(n1262)
         );
  MUX41X1_HVT U1429 ( .A1(\ram[4][164] ), .A3(\ram[6][164] ), .A2(
        \ram[5][164] ), .A4(\ram[7][164] ), .S0(n516), .S1(n423), .Y(n1263) );
  MUX41X1_HVT U1430 ( .A1(\ram[0][164] ), .A3(\ram[2][164] ), .A2(
        \ram[1][164] ), .A4(\ram[3][164] ), .S0(n516), .S1(n423), .Y(n1264) );
  MUX41X1_HVT U1431 ( .A1(n1264), .A3(n1262), .A2(n1263), .A4(n1261), .S0(n593), .S1(n560), .Y(q[164]) );
  MUX41X1_HVT U1432 ( .A1(\ram[12][165] ), .A3(\ram[14][165] ), .A2(
        \ram[13][165] ), .A4(\ram[15][165] ), .S0(n517), .S1(n424), .Y(n1265)
         );
  MUX41X1_HVT U1433 ( .A1(\ram[8][165] ), .A3(\ram[10][165] ), .A2(
        \ram[9][165] ), .A4(\ram[11][165] ), .S0(n517), .S1(n424), .Y(n1266)
         );
  MUX41X1_HVT U1434 ( .A1(\ram[4][165] ), .A3(\ram[6][165] ), .A2(
        \ram[5][165] ), .A4(\ram[7][165] ), .S0(n517), .S1(n424), .Y(n1267) );
  MUX41X1_HVT U1435 ( .A1(\ram[0][165] ), .A3(\ram[2][165] ), .A2(
        \ram[1][165] ), .A4(\ram[3][165] ), .S0(n517), .S1(n424), .Y(n1268) );
  MUX41X1_HVT U1436 ( .A1(n1268), .A3(n1266), .A2(n1267), .A4(n1265), .S0(n593), .S1(n560), .Y(q[165]) );
  MUX41X1_HVT U1437 ( .A1(\ram[12][166] ), .A3(\ram[14][166] ), .A2(
        \ram[13][166] ), .A4(\ram[15][166] ), .S0(n517), .S1(n424), .Y(n1269)
         );
  MUX41X1_HVT U1438 ( .A1(\ram[8][166] ), .A3(\ram[10][166] ), .A2(
        \ram[9][166] ), .A4(\ram[11][166] ), .S0(n517), .S1(n424), .Y(n1270)
         );
  MUX41X1_HVT U1439 ( .A1(\ram[4][166] ), .A3(\ram[6][166] ), .A2(
        \ram[5][166] ), .A4(\ram[7][166] ), .S0(n517), .S1(n424), .Y(n1271) );
  MUX41X1_HVT U1440 ( .A1(\ram[0][166] ), .A3(\ram[2][166] ), .A2(
        \ram[1][166] ), .A4(\ram[3][166] ), .S0(n517), .S1(n424), .Y(n1272) );
  MUX41X1_HVT U1441 ( .A1(n1272), .A3(n1270), .A2(n1271), .A4(n1269), .S0(n593), .S1(n560), .Y(q[166]) );
  MUX41X1_HVT U1442 ( .A1(\ram[12][167] ), .A3(\ram[14][167] ), .A2(
        \ram[13][167] ), .A4(\ram[15][167] ), .S0(n517), .S1(n424), .Y(n1273)
         );
  MUX41X1_HVT U1443 ( .A1(\ram[8][167] ), .A3(\ram[10][167] ), .A2(
        \ram[9][167] ), .A4(\ram[11][167] ), .S0(n517), .S1(n424), .Y(n1274)
         );
  MUX41X1_HVT U1444 ( .A1(\ram[4][167] ), .A3(\ram[6][167] ), .A2(
        \ram[5][167] ), .A4(\ram[7][167] ), .S0(n517), .S1(n424), .Y(n1275) );
  MUX41X1_HVT U1445 ( .A1(\ram[0][167] ), .A3(\ram[2][167] ), .A2(
        \ram[1][167] ), .A4(\ram[3][167] ), .S0(n517), .S1(n424), .Y(n1276) );
  MUX41X1_HVT U1446 ( .A1(n1276), .A3(n1274), .A2(n1275), .A4(n1273), .S0(n593), .S1(n560), .Y(q[167]) );
  MUX41X1_HVT U1447 ( .A1(\ram[12][168] ), .A3(\ram[14][168] ), .A2(
        \ram[13][168] ), .A4(\ram[15][168] ), .S0(n518), .S1(n425), .Y(n1277)
         );
  MUX41X1_HVT U1448 ( .A1(\ram[8][168] ), .A3(\ram[10][168] ), .A2(
        \ram[9][168] ), .A4(\ram[11][168] ), .S0(n518), .S1(n425), .Y(n1278)
         );
  MUX41X1_HVT U1449 ( .A1(\ram[4][168] ), .A3(\ram[6][168] ), .A2(
        \ram[5][168] ), .A4(\ram[7][168] ), .S0(n518), .S1(n425), .Y(n1279) );
  MUX41X1_HVT U1450 ( .A1(\ram[0][168] ), .A3(\ram[2][168] ), .A2(
        \ram[1][168] ), .A4(\ram[3][168] ), .S0(n518), .S1(n425), .Y(n1280) );
  MUX41X1_HVT U1451 ( .A1(n1280), .A3(n1278), .A2(n1279), .A4(n1277), .S0(n594), .S1(n560), .Y(q[168]) );
  MUX41X1_HVT U1452 ( .A1(\ram[12][169] ), .A3(\ram[14][169] ), .A2(
        \ram[13][169] ), .A4(\ram[15][169] ), .S0(n518), .S1(n425), .Y(n1281)
         );
  MUX41X1_HVT U1453 ( .A1(\ram[8][169] ), .A3(\ram[10][169] ), .A2(
        \ram[9][169] ), .A4(\ram[11][169] ), .S0(n518), .S1(n425), .Y(n1282)
         );
  MUX41X1_HVT U1454 ( .A1(\ram[4][169] ), .A3(\ram[6][169] ), .A2(
        \ram[5][169] ), .A4(\ram[7][169] ), .S0(n518), .S1(n425), .Y(n1283) );
  MUX41X1_HVT U1455 ( .A1(\ram[0][169] ), .A3(\ram[2][169] ), .A2(
        \ram[1][169] ), .A4(\ram[3][169] ), .S0(n518), .S1(n425), .Y(n1284) );
  MUX41X1_HVT U1456 ( .A1(n1284), .A3(n1282), .A2(n1283), .A4(n1281), .S0(n594), .S1(n560), .Y(q[169]) );
  MUX41X1_HVT U1457 ( .A1(\ram[12][170] ), .A3(\ram[14][170] ), .A2(
        \ram[13][170] ), .A4(\ram[15][170] ), .S0(n518), .S1(n425), .Y(n1285)
         );
  MUX41X1_HVT U1458 ( .A1(\ram[8][170] ), .A3(\ram[10][170] ), .A2(
        \ram[9][170] ), .A4(\ram[11][170] ), .S0(n518), .S1(n425), .Y(n1286)
         );
  MUX41X1_HVT U1459 ( .A1(\ram[4][170] ), .A3(\ram[6][170] ), .A2(
        \ram[5][170] ), .A4(\ram[7][170] ), .S0(n518), .S1(n425), .Y(n1287) );
  MUX41X1_HVT U1460 ( .A1(\ram[0][170] ), .A3(\ram[2][170] ), .A2(
        \ram[1][170] ), .A4(\ram[3][170] ), .S0(n518), .S1(n425), .Y(n1288) );
  MUX41X1_HVT U1461 ( .A1(n1288), .A3(n1286), .A2(n1287), .A4(n1285), .S0(n594), .S1(n560), .Y(q[170]) );
  MUX41X1_HVT U1462 ( .A1(\ram[12][171] ), .A3(\ram[14][171] ), .A2(
        \ram[13][171] ), .A4(\ram[15][171] ), .S0(n519), .S1(n426), .Y(n1289)
         );
  MUX41X1_HVT U1463 ( .A1(\ram[8][171] ), .A3(\ram[10][171] ), .A2(
        \ram[9][171] ), .A4(\ram[11][171] ), .S0(n519), .S1(n426), .Y(n1290)
         );
  MUX41X1_HVT U1464 ( .A1(\ram[4][171] ), .A3(\ram[6][171] ), .A2(
        \ram[5][171] ), .A4(\ram[7][171] ), .S0(n519), .S1(n426), .Y(n1291) );
  MUX41X1_HVT U1465 ( .A1(\ram[0][171] ), .A3(\ram[2][171] ), .A2(
        \ram[1][171] ), .A4(\ram[3][171] ), .S0(n519), .S1(n426), .Y(n1292) );
  MUX41X1_HVT U1466 ( .A1(n1292), .A3(n1290), .A2(n1291), .A4(n1289), .S0(n594), .S1(n560), .Y(q[171]) );
  MUX41X1_HVT U1467 ( .A1(\ram[12][172] ), .A3(\ram[14][172] ), .A2(
        \ram[13][172] ), .A4(\ram[15][172] ), .S0(n519), .S1(n426), .Y(n1293)
         );
  MUX41X1_HVT U1468 ( .A1(\ram[8][172] ), .A3(\ram[10][172] ), .A2(
        \ram[9][172] ), .A4(\ram[11][172] ), .S0(n519), .S1(n426), .Y(n1294)
         );
  MUX41X1_HVT U1469 ( .A1(\ram[4][172] ), .A3(\ram[6][172] ), .A2(
        \ram[5][172] ), .A4(\ram[7][172] ), .S0(n519), .S1(n426), .Y(n1295) );
  MUX41X1_HVT U1470 ( .A1(\ram[0][172] ), .A3(\ram[2][172] ), .A2(
        \ram[1][172] ), .A4(\ram[3][172] ), .S0(n519), .S1(n426), .Y(n1296) );
  MUX41X1_HVT U1471 ( .A1(n1296), .A3(n1294), .A2(n1295), .A4(n1293), .S0(n594), .S1(n560), .Y(q[172]) );
  MUX41X1_HVT U1472 ( .A1(\ram[12][173] ), .A3(\ram[14][173] ), .A2(
        \ram[13][173] ), .A4(\ram[15][173] ), .S0(n519), .S1(n426), .Y(n1297)
         );
  MUX41X1_HVT U1473 ( .A1(\ram[8][173] ), .A3(\ram[10][173] ), .A2(
        \ram[9][173] ), .A4(\ram[11][173] ), .S0(n519), .S1(n426), .Y(n1298)
         );
  MUX41X1_HVT U1474 ( .A1(\ram[4][173] ), .A3(\ram[6][173] ), .A2(
        \ram[5][173] ), .A4(\ram[7][173] ), .S0(n519), .S1(n426), .Y(n1299) );
  MUX41X1_HVT U1475 ( .A1(\ram[0][173] ), .A3(\ram[2][173] ), .A2(
        \ram[1][173] ), .A4(\ram[3][173] ), .S0(n519), .S1(n426), .Y(n1300) );
  MUX41X1_HVT U1476 ( .A1(n1300), .A3(n1298), .A2(n1299), .A4(n1297), .S0(n594), .S1(n560), .Y(q[173]) );
  MUX41X1_HVT U1477 ( .A1(\ram[12][174] ), .A3(\ram[14][174] ), .A2(
        \ram[13][174] ), .A4(\ram[15][174] ), .S0(n520), .S1(n427), .Y(n1301)
         );
  MUX41X1_HVT U1478 ( .A1(\ram[8][174] ), .A3(\ram[10][174] ), .A2(
        \ram[9][174] ), .A4(\ram[11][174] ), .S0(n520), .S1(n427), .Y(n1302)
         );
  MUX41X1_HVT U1479 ( .A1(\ram[4][174] ), .A3(\ram[6][174] ), .A2(
        \ram[5][174] ), .A4(\ram[7][174] ), .S0(n520), .S1(n427), .Y(n1303) );
  MUX41X1_HVT U1480 ( .A1(\ram[0][174] ), .A3(\ram[2][174] ), .A2(
        \ram[1][174] ), .A4(\ram[3][174] ), .S0(n520), .S1(n427), .Y(n1304) );
  MUX41X1_HVT U1481 ( .A1(n1304), .A3(n1302), .A2(n1303), .A4(n1301), .S0(n594), .S1(n560), .Y(q[174]) );
  MUX41X1_HVT U1482 ( .A1(\ram[12][175] ), .A3(\ram[14][175] ), .A2(
        \ram[13][175] ), .A4(\ram[15][175] ), .S0(n520), .S1(n427), .Y(n1305)
         );
  MUX41X1_HVT U1483 ( .A1(\ram[8][175] ), .A3(\ram[10][175] ), .A2(
        \ram[9][175] ), .A4(\ram[11][175] ), .S0(n520), .S1(n427), .Y(n1306)
         );
  MUX41X1_HVT U1484 ( .A1(\ram[4][175] ), .A3(\ram[6][175] ), .A2(
        \ram[5][175] ), .A4(\ram[7][175] ), .S0(n520), .S1(n427), .Y(n1307) );
  MUX41X1_HVT U1485 ( .A1(\ram[0][175] ), .A3(\ram[2][175] ), .A2(
        \ram[1][175] ), .A4(\ram[3][175] ), .S0(n520), .S1(n427), .Y(n1308) );
  MUX41X1_HVT U1486 ( .A1(n1308), .A3(n1306), .A2(n1307), .A4(n1305), .S0(n594), .S1(n560), .Y(q[175]) );
  MUX41X1_HVT U1487 ( .A1(\ram[12][176] ), .A3(\ram[14][176] ), .A2(
        \ram[13][176] ), .A4(\ram[15][176] ), .S0(n520), .S1(n427), .Y(n1309)
         );
  MUX41X1_HVT U1488 ( .A1(\ram[8][176] ), .A3(\ram[10][176] ), .A2(
        \ram[9][176] ), .A4(\ram[11][176] ), .S0(n520), .S1(n427), .Y(n1310)
         );
  MUX41X1_HVT U1489 ( .A1(\ram[4][176] ), .A3(\ram[6][176] ), .A2(
        \ram[5][176] ), .A4(\ram[7][176] ), .S0(n520), .S1(n427), .Y(n1311) );
  MUX41X1_HVT U1490 ( .A1(\ram[0][176] ), .A3(\ram[2][176] ), .A2(
        \ram[1][176] ), .A4(\ram[3][176] ), .S0(n520), .S1(n427), .Y(n1312) );
  MUX41X1_HVT U1491 ( .A1(n1312), .A3(n1310), .A2(n1311), .A4(n1309), .S0(n594), .S1(n561), .Y(q[176]) );
  MUX41X1_HVT U1492 ( .A1(\ram[12][177] ), .A3(\ram[14][177] ), .A2(
        \ram[13][177] ), .A4(\ram[15][177] ), .S0(n521), .S1(n428), .Y(n1313)
         );
  MUX41X1_HVT U1493 ( .A1(\ram[8][177] ), .A3(\ram[10][177] ), .A2(
        \ram[9][177] ), .A4(\ram[11][177] ), .S0(n521), .S1(n428), .Y(n1314)
         );
  MUX41X1_HVT U1494 ( .A1(\ram[4][177] ), .A3(\ram[6][177] ), .A2(
        \ram[5][177] ), .A4(\ram[7][177] ), .S0(n521), .S1(n428), .Y(n1315) );
  MUX41X1_HVT U1495 ( .A1(\ram[0][177] ), .A3(\ram[2][177] ), .A2(
        \ram[1][177] ), .A4(\ram[3][177] ), .S0(n521), .S1(n428), .Y(n1316) );
  MUX41X1_HVT U1496 ( .A1(n1316), .A3(n1314), .A2(n1315), .A4(n1313), .S0(n594), .S1(n561), .Y(q[177]) );
  MUX41X1_HVT U1497 ( .A1(\ram[12][178] ), .A3(\ram[14][178] ), .A2(
        \ram[13][178] ), .A4(\ram[15][178] ), .S0(n521), .S1(n428), .Y(n1317)
         );
  MUX41X1_HVT U1498 ( .A1(\ram[8][178] ), .A3(\ram[10][178] ), .A2(
        \ram[9][178] ), .A4(\ram[11][178] ), .S0(n521), .S1(n428), .Y(n1318)
         );
  MUX41X1_HVT U1499 ( .A1(\ram[4][178] ), .A3(\ram[6][178] ), .A2(
        \ram[5][178] ), .A4(\ram[7][178] ), .S0(n521), .S1(n428), .Y(n1319) );
  MUX41X1_HVT U1500 ( .A1(\ram[0][178] ), .A3(\ram[2][178] ), .A2(
        \ram[1][178] ), .A4(\ram[3][178] ), .S0(n521), .S1(n428), .Y(n1320) );
  MUX41X1_HVT U1501 ( .A1(n1320), .A3(n1318), .A2(n1319), .A4(n1317), .S0(n594), .S1(n561), .Y(q[178]) );
  MUX41X1_HVT U1502 ( .A1(\ram[12][179] ), .A3(\ram[14][179] ), .A2(
        \ram[13][179] ), .A4(\ram[15][179] ), .S0(n521), .S1(n428), .Y(n1321)
         );
  MUX41X1_HVT U1503 ( .A1(\ram[8][179] ), .A3(\ram[10][179] ), .A2(
        \ram[9][179] ), .A4(\ram[11][179] ), .S0(n521), .S1(n428), .Y(n1322)
         );
  MUX41X1_HVT U1504 ( .A1(\ram[4][179] ), .A3(\ram[6][179] ), .A2(
        \ram[5][179] ), .A4(\ram[7][179] ), .S0(n521), .S1(n428), .Y(n1323) );
  MUX41X1_HVT U1505 ( .A1(\ram[0][179] ), .A3(\ram[2][179] ), .A2(
        \ram[1][179] ), .A4(\ram[3][179] ), .S0(n521), .S1(n428), .Y(n1324) );
  MUX41X1_HVT U1506 ( .A1(n1324), .A3(n1322), .A2(n1323), .A4(n1321), .S0(n594), .S1(n561), .Y(q[179]) );
  MUX41X1_HVT U1507 ( .A1(\ram[12][180] ), .A3(\ram[14][180] ), .A2(
        \ram[13][180] ), .A4(\ram[15][180] ), .S0(n522), .S1(n429), .Y(n1325)
         );
  MUX41X1_HVT U1508 ( .A1(\ram[8][180] ), .A3(\ram[10][180] ), .A2(
        \ram[9][180] ), .A4(\ram[11][180] ), .S0(n522), .S1(n429), .Y(n1326)
         );
  MUX41X1_HVT U1509 ( .A1(\ram[4][180] ), .A3(\ram[6][180] ), .A2(
        \ram[5][180] ), .A4(\ram[7][180] ), .S0(n522), .S1(n429), .Y(n1327) );
  MUX41X1_HVT U1510 ( .A1(\ram[0][180] ), .A3(\ram[2][180] ), .A2(
        \ram[1][180] ), .A4(\ram[3][180] ), .S0(n522), .S1(n429), .Y(n1328) );
  MUX41X1_HVT U1511 ( .A1(n1328), .A3(n1326), .A2(n1327), .A4(n1325), .S0(n595), .S1(n561), .Y(q[180]) );
  MUX41X1_HVT U1512 ( .A1(\ram[12][181] ), .A3(\ram[14][181] ), .A2(
        \ram[13][181] ), .A4(\ram[15][181] ), .S0(n522), .S1(n429), .Y(n1329)
         );
  MUX41X1_HVT U1513 ( .A1(\ram[8][181] ), .A3(\ram[10][181] ), .A2(
        \ram[9][181] ), .A4(\ram[11][181] ), .S0(n522), .S1(n429), .Y(n1330)
         );
  MUX41X1_HVT U1514 ( .A1(\ram[4][181] ), .A3(\ram[6][181] ), .A2(
        \ram[5][181] ), .A4(\ram[7][181] ), .S0(n522), .S1(n429), .Y(n1331) );
  MUX41X1_HVT U1515 ( .A1(\ram[0][181] ), .A3(\ram[2][181] ), .A2(
        \ram[1][181] ), .A4(\ram[3][181] ), .S0(n522), .S1(n429), .Y(n1332) );
  MUX41X1_HVT U1516 ( .A1(n1332), .A3(n1330), .A2(n1331), .A4(n1329), .S0(n595), .S1(n561), .Y(q[181]) );
  MUX41X1_HVT U1517 ( .A1(\ram[12][182] ), .A3(\ram[14][182] ), .A2(
        \ram[13][182] ), .A4(\ram[15][182] ), .S0(n522), .S1(n429), .Y(n1333)
         );
  MUX41X1_HVT U1518 ( .A1(\ram[8][182] ), .A3(\ram[10][182] ), .A2(
        \ram[9][182] ), .A4(\ram[11][182] ), .S0(n522), .S1(n429), .Y(n1334)
         );
  MUX41X1_HVT U1519 ( .A1(\ram[4][182] ), .A3(\ram[6][182] ), .A2(
        \ram[5][182] ), .A4(\ram[7][182] ), .S0(n522), .S1(n429), .Y(n1335) );
  MUX41X1_HVT U1520 ( .A1(\ram[0][182] ), .A3(\ram[2][182] ), .A2(
        \ram[1][182] ), .A4(\ram[3][182] ), .S0(n522), .S1(n429), .Y(n1336) );
  MUX41X1_HVT U1521 ( .A1(n1336), .A3(n1334), .A2(n1335), .A4(n1333), .S0(n595), .S1(n561), .Y(q[182]) );
  MUX41X1_HVT U1522 ( .A1(\ram[12][183] ), .A3(\ram[14][183] ), .A2(
        \ram[13][183] ), .A4(\ram[15][183] ), .S0(n523), .S1(n430), .Y(n1337)
         );
  MUX41X1_HVT U1523 ( .A1(\ram[8][183] ), .A3(\ram[10][183] ), .A2(
        \ram[9][183] ), .A4(\ram[11][183] ), .S0(n523), .S1(n430), .Y(n1338)
         );
  MUX41X1_HVT U1524 ( .A1(\ram[4][183] ), .A3(\ram[6][183] ), .A2(
        \ram[5][183] ), .A4(\ram[7][183] ), .S0(n523), .S1(n430), .Y(n1339) );
  MUX41X1_HVT U1525 ( .A1(\ram[0][183] ), .A3(\ram[2][183] ), .A2(
        \ram[1][183] ), .A4(\ram[3][183] ), .S0(n523), .S1(n430), .Y(n1340) );
  MUX41X1_HVT U1526 ( .A1(n1340), .A3(n1338), .A2(n1339), .A4(n1337), .S0(n595), .S1(n561), .Y(q[183]) );
  MUX41X1_HVT U1527 ( .A1(\ram[12][184] ), .A3(\ram[14][184] ), .A2(
        \ram[13][184] ), .A4(\ram[15][184] ), .S0(n523), .S1(n430), .Y(n1341)
         );
  MUX41X1_HVT U1528 ( .A1(\ram[8][184] ), .A3(\ram[10][184] ), .A2(
        \ram[9][184] ), .A4(\ram[11][184] ), .S0(n523), .S1(n430), .Y(n1342)
         );
  MUX41X1_HVT U1529 ( .A1(\ram[4][184] ), .A3(\ram[6][184] ), .A2(
        \ram[5][184] ), .A4(\ram[7][184] ), .S0(n523), .S1(n430), .Y(n1343) );
  MUX41X1_HVT U1530 ( .A1(\ram[0][184] ), .A3(\ram[2][184] ), .A2(
        \ram[1][184] ), .A4(\ram[3][184] ), .S0(n523), .S1(n430), .Y(n1344) );
  MUX41X1_HVT U1531 ( .A1(n1344), .A3(n1342), .A2(n1343), .A4(n1341), .S0(n595), .S1(n561), .Y(q[184]) );
  MUX41X1_HVT U1532 ( .A1(\ram[12][185] ), .A3(\ram[14][185] ), .A2(
        \ram[13][185] ), .A4(\ram[15][185] ), .S0(n523), .S1(n430), .Y(n1345)
         );
  MUX41X1_HVT U1533 ( .A1(\ram[8][185] ), .A3(\ram[10][185] ), .A2(
        \ram[9][185] ), .A4(\ram[11][185] ), .S0(n523), .S1(n430), .Y(n1346)
         );
  MUX41X1_HVT U1534 ( .A1(\ram[4][185] ), .A3(\ram[6][185] ), .A2(
        \ram[5][185] ), .A4(\ram[7][185] ), .S0(n523), .S1(n430), .Y(n1347) );
  MUX41X1_HVT U1535 ( .A1(\ram[0][185] ), .A3(\ram[2][185] ), .A2(
        \ram[1][185] ), .A4(\ram[3][185] ), .S0(n523), .S1(n430), .Y(n1348) );
  MUX41X1_HVT U1536 ( .A1(n1348), .A3(n1346), .A2(n1347), .A4(n1345), .S0(n595), .S1(n561), .Y(q[185]) );
  MUX41X1_HVT U1537 ( .A1(\ram[12][186] ), .A3(\ram[14][186] ), .A2(
        \ram[13][186] ), .A4(\ram[15][186] ), .S0(n524), .S1(n431), .Y(n1349)
         );
  MUX41X1_HVT U1538 ( .A1(\ram[8][186] ), .A3(\ram[10][186] ), .A2(
        \ram[9][186] ), .A4(\ram[11][186] ), .S0(n524), .S1(n431), .Y(n1350)
         );
  MUX41X1_HVT U1539 ( .A1(\ram[4][186] ), .A3(\ram[6][186] ), .A2(
        \ram[5][186] ), .A4(\ram[7][186] ), .S0(n524), .S1(n431), .Y(n1351) );
  MUX41X1_HVT U1540 ( .A1(\ram[0][186] ), .A3(\ram[2][186] ), .A2(
        \ram[1][186] ), .A4(\ram[3][186] ), .S0(n524), .S1(n431), .Y(n1352) );
  MUX41X1_HVT U1541 ( .A1(n1352), .A3(n1350), .A2(n1351), .A4(n1349), .S0(n595), .S1(n561), .Y(q[186]) );
  MUX41X1_HVT U1542 ( .A1(\ram[12][187] ), .A3(\ram[14][187] ), .A2(
        \ram[13][187] ), .A4(\ram[15][187] ), .S0(n524), .S1(n431), .Y(n1353)
         );
  MUX41X1_HVT U1543 ( .A1(\ram[8][187] ), .A3(\ram[10][187] ), .A2(
        \ram[9][187] ), .A4(\ram[11][187] ), .S0(n524), .S1(n431), .Y(n1354)
         );
  MUX41X1_HVT U1544 ( .A1(\ram[4][187] ), .A3(\ram[6][187] ), .A2(
        \ram[5][187] ), .A4(\ram[7][187] ), .S0(n524), .S1(n431), .Y(n1355) );
  MUX41X1_HVT U1545 ( .A1(\ram[0][187] ), .A3(\ram[2][187] ), .A2(
        \ram[1][187] ), .A4(\ram[3][187] ), .S0(n524), .S1(n431), .Y(n1356) );
  MUX41X1_HVT U1546 ( .A1(n1356), .A3(n1354), .A2(n1355), .A4(n1353), .S0(n595), .S1(n561), .Y(q[187]) );
  MUX41X1_HVT U1547 ( .A1(\ram[12][188] ), .A3(\ram[14][188] ), .A2(
        \ram[13][188] ), .A4(\ram[15][188] ), .S0(n524), .S1(n431), .Y(n1357)
         );
  MUX41X1_HVT U1548 ( .A1(\ram[8][188] ), .A3(\ram[10][188] ), .A2(
        \ram[9][188] ), .A4(\ram[11][188] ), .S0(n524), .S1(n431), .Y(n1358)
         );
  MUX41X1_HVT U1549 ( .A1(\ram[4][188] ), .A3(\ram[6][188] ), .A2(
        \ram[5][188] ), .A4(\ram[7][188] ), .S0(n524), .S1(n431), .Y(n1359) );
  MUX41X1_HVT U1550 ( .A1(\ram[0][188] ), .A3(\ram[2][188] ), .A2(
        \ram[1][188] ), .A4(\ram[3][188] ), .S0(n524), .S1(n431), .Y(n1360) );
  MUX41X1_HVT U1551 ( .A1(n1360), .A3(n1358), .A2(n1359), .A4(n1357), .S0(n595), .S1(n562), .Y(q[188]) );
  MUX41X1_HVT U1552 ( .A1(\ram[12][189] ), .A3(\ram[14][189] ), .A2(
        \ram[13][189] ), .A4(\ram[15][189] ), .S0(n525), .S1(n432), .Y(n1361)
         );
  MUX41X1_HVT U1553 ( .A1(\ram[8][189] ), .A3(\ram[10][189] ), .A2(
        \ram[9][189] ), .A4(\ram[11][189] ), .S0(n525), .S1(n432), .Y(n1362)
         );
  MUX41X1_HVT U1554 ( .A1(\ram[4][189] ), .A3(\ram[6][189] ), .A2(
        \ram[5][189] ), .A4(\ram[7][189] ), .S0(n525), .S1(n432), .Y(n1363) );
  MUX41X1_HVT U1555 ( .A1(\ram[0][189] ), .A3(\ram[2][189] ), .A2(
        \ram[1][189] ), .A4(\ram[3][189] ), .S0(n525), .S1(n432), .Y(n1364) );
  MUX41X1_HVT U1556 ( .A1(n1364), .A3(n1362), .A2(n1363), .A4(n1361), .S0(n595), .S1(n562), .Y(q[189]) );
  MUX41X1_HVT U1557 ( .A1(\ram[12][190] ), .A3(\ram[14][190] ), .A2(
        \ram[13][190] ), .A4(\ram[15][190] ), .S0(n525), .S1(n432), .Y(n1365)
         );
  MUX41X1_HVT U1558 ( .A1(\ram[8][190] ), .A3(\ram[10][190] ), .A2(
        \ram[9][190] ), .A4(\ram[11][190] ), .S0(n525), .S1(n432), .Y(n1366)
         );
  MUX41X1_HVT U1559 ( .A1(\ram[4][190] ), .A3(\ram[6][190] ), .A2(
        \ram[5][190] ), .A4(\ram[7][190] ), .S0(n525), .S1(n432), .Y(n1367) );
  MUX41X1_HVT U1560 ( .A1(\ram[0][190] ), .A3(\ram[2][190] ), .A2(
        \ram[1][190] ), .A4(\ram[3][190] ), .S0(n525), .S1(n432), .Y(n1368) );
  MUX41X1_HVT U1561 ( .A1(n1368), .A3(n1366), .A2(n1367), .A4(n1365), .S0(n595), .S1(n562), .Y(q[190]) );
  MUX41X1_HVT U1562 ( .A1(\ram[12][191] ), .A3(\ram[14][191] ), .A2(
        \ram[13][191] ), .A4(\ram[15][191] ), .S0(n525), .S1(n432), .Y(n1369)
         );
  MUX41X1_HVT U1563 ( .A1(\ram[8][191] ), .A3(\ram[10][191] ), .A2(
        \ram[9][191] ), .A4(\ram[11][191] ), .S0(n525), .S1(n432), .Y(n1370)
         );
  MUX41X1_HVT U1564 ( .A1(\ram[4][191] ), .A3(\ram[6][191] ), .A2(
        \ram[5][191] ), .A4(\ram[7][191] ), .S0(n525), .S1(n432), .Y(n1371) );
  MUX41X1_HVT U1565 ( .A1(\ram[0][191] ), .A3(\ram[2][191] ), .A2(
        \ram[1][191] ), .A4(\ram[3][191] ), .S0(n525), .S1(n432), .Y(n1372) );
  MUX41X1_HVT U1566 ( .A1(n1372), .A3(n1370), .A2(n1371), .A4(n1369), .S0(n595), .S1(n562), .Y(q[191]) );
  MUX41X1_HVT U1567 ( .A1(\ram[12][192] ), .A3(\ram[14][192] ), .A2(
        \ram[13][192] ), .A4(\ram[15][192] ), .S0(n526), .S1(n433), .Y(n1373)
         );
  MUX41X1_HVT U1568 ( .A1(\ram[8][192] ), .A3(\ram[10][192] ), .A2(
        \ram[9][192] ), .A4(\ram[11][192] ), .S0(n526), .S1(n433), .Y(n1374)
         );
  MUX41X1_HVT U1569 ( .A1(\ram[4][192] ), .A3(\ram[6][192] ), .A2(
        \ram[5][192] ), .A4(\ram[7][192] ), .S0(n526), .S1(n433), .Y(n1375) );
  MUX41X1_HVT U1570 ( .A1(\ram[0][192] ), .A3(\ram[2][192] ), .A2(
        \ram[1][192] ), .A4(\ram[3][192] ), .S0(n526), .S1(n433), .Y(n1376) );
  MUX41X1_HVT U1571 ( .A1(n1376), .A3(n1374), .A2(n1375), .A4(n1373), .S0(n596), .S1(n562), .Y(q[192]) );
  MUX41X1_HVT U1572 ( .A1(\ram[12][193] ), .A3(\ram[14][193] ), .A2(
        \ram[13][193] ), .A4(\ram[15][193] ), .S0(n526), .S1(n433), .Y(n1377)
         );
  MUX41X1_HVT U1573 ( .A1(\ram[8][193] ), .A3(\ram[10][193] ), .A2(
        \ram[9][193] ), .A4(\ram[11][193] ), .S0(n526), .S1(n433), .Y(n1378)
         );
  MUX41X1_HVT U1574 ( .A1(\ram[4][193] ), .A3(\ram[6][193] ), .A2(
        \ram[5][193] ), .A4(\ram[7][193] ), .S0(n526), .S1(n433), .Y(n1379) );
  MUX41X1_HVT U1575 ( .A1(\ram[0][193] ), .A3(\ram[2][193] ), .A2(
        \ram[1][193] ), .A4(\ram[3][193] ), .S0(n526), .S1(n433), .Y(n1380) );
  MUX41X1_HVT U1576 ( .A1(n1380), .A3(n1378), .A2(n1379), .A4(n1377), .S0(n596), .S1(n567), .Y(q[193]) );
  MUX41X1_HVT U1577 ( .A1(\ram[12][194] ), .A3(\ram[14][194] ), .A2(
        \ram[13][194] ), .A4(\ram[15][194] ), .S0(n526), .S1(n433), .Y(n1381)
         );
  MUX41X1_HVT U1578 ( .A1(\ram[8][194] ), .A3(\ram[10][194] ), .A2(
        \ram[9][194] ), .A4(\ram[11][194] ), .S0(n526), .S1(n433), .Y(n1382)
         );
  MUX41X1_HVT U1579 ( .A1(\ram[4][194] ), .A3(\ram[6][194] ), .A2(
        \ram[5][194] ), .A4(\ram[7][194] ), .S0(n526), .S1(n433), .Y(n1383) );
  MUX41X1_HVT U1580 ( .A1(\ram[0][194] ), .A3(\ram[2][194] ), .A2(
        \ram[1][194] ), .A4(\ram[3][194] ), .S0(n526), .S1(n433), .Y(n1384) );
  MUX41X1_HVT U1581 ( .A1(n1384), .A3(n1382), .A2(n1383), .A4(n1381), .S0(n596), .S1(n562), .Y(q[194]) );
  MUX41X1_HVT U1582 ( .A1(\ram[12][195] ), .A3(\ram[14][195] ), .A2(
        \ram[13][195] ), .A4(\ram[15][195] ), .S0(n527), .S1(n434), .Y(n1385)
         );
  MUX41X1_HVT U1583 ( .A1(\ram[8][195] ), .A3(\ram[10][195] ), .A2(
        \ram[9][195] ), .A4(\ram[11][195] ), .S0(n527), .S1(n434), .Y(n1386)
         );
  MUX41X1_HVT U1584 ( .A1(\ram[4][195] ), .A3(\ram[6][195] ), .A2(
        \ram[5][195] ), .A4(\ram[7][195] ), .S0(n527), .S1(n434), .Y(n1387) );
  MUX41X1_HVT U1585 ( .A1(\ram[0][195] ), .A3(\ram[2][195] ), .A2(
        \ram[1][195] ), .A4(\ram[3][195] ), .S0(n527), .S1(n434), .Y(n1388) );
  MUX41X1_HVT U1586 ( .A1(n1388), .A3(n1386), .A2(n1387), .A4(n1385), .S0(n596), .S1(n562), .Y(q[195]) );
  MUX41X1_HVT U1587 ( .A1(\ram[12][196] ), .A3(\ram[14][196] ), .A2(
        \ram[13][196] ), .A4(\ram[15][196] ), .S0(n527), .S1(n434), .Y(n1389)
         );
  MUX41X1_HVT U1588 ( .A1(\ram[8][196] ), .A3(\ram[10][196] ), .A2(
        \ram[9][196] ), .A4(\ram[11][196] ), .S0(n527), .S1(n434), .Y(n1390)
         );
  MUX41X1_HVT U1589 ( .A1(\ram[4][196] ), .A3(\ram[6][196] ), .A2(
        \ram[5][196] ), .A4(\ram[7][196] ), .S0(n527), .S1(n434), .Y(n1391) );
  MUX41X1_HVT U1590 ( .A1(\ram[0][196] ), .A3(\ram[2][196] ), .A2(
        \ram[1][196] ), .A4(\ram[3][196] ), .S0(n527), .S1(n434), .Y(n1392) );
  MUX41X1_HVT U1591 ( .A1(n1392), .A3(n1390), .A2(n1391), .A4(n1389), .S0(n596), .S1(n562), .Y(q[196]) );
  MUX41X1_HVT U1592 ( .A1(\ram[12][197] ), .A3(\ram[14][197] ), .A2(
        \ram[13][197] ), .A4(\ram[15][197] ), .S0(n527), .S1(n434), .Y(n1393)
         );
  MUX41X1_HVT U1593 ( .A1(\ram[8][197] ), .A3(\ram[10][197] ), .A2(
        \ram[9][197] ), .A4(\ram[11][197] ), .S0(n527), .S1(n434), .Y(n1394)
         );
  MUX41X1_HVT U1594 ( .A1(\ram[4][197] ), .A3(\ram[6][197] ), .A2(
        \ram[5][197] ), .A4(\ram[7][197] ), .S0(n527), .S1(n434), .Y(n1395) );
  MUX41X1_HVT U1595 ( .A1(\ram[0][197] ), .A3(\ram[2][197] ), .A2(
        \ram[1][197] ), .A4(\ram[3][197] ), .S0(n527), .S1(n434), .Y(n1396) );
  MUX41X1_HVT U1596 ( .A1(n1396), .A3(n1394), .A2(n1395), .A4(n1393), .S0(n596), .S1(n562), .Y(q[197]) );
  MUX41X1_HVT U1597 ( .A1(\ram[12][198] ), .A3(\ram[14][198] ), .A2(
        \ram[13][198] ), .A4(\ram[15][198] ), .S0(n528), .S1(n435), .Y(n1397)
         );
  MUX41X1_HVT U1598 ( .A1(\ram[8][198] ), .A3(\ram[10][198] ), .A2(
        \ram[9][198] ), .A4(\ram[11][198] ), .S0(n528), .S1(n435), .Y(n1398)
         );
  MUX41X1_HVT U1599 ( .A1(\ram[4][198] ), .A3(\ram[6][198] ), .A2(
        \ram[5][198] ), .A4(\ram[7][198] ), .S0(n528), .S1(n435), .Y(n1399) );
  MUX41X1_HVT U1600 ( .A1(\ram[0][198] ), .A3(\ram[2][198] ), .A2(
        \ram[1][198] ), .A4(\ram[3][198] ), .S0(n528), .S1(n435), .Y(n1400) );
  MUX41X1_HVT U1601 ( .A1(n1400), .A3(n1398), .A2(n1399), .A4(n1397), .S0(n596), .S1(n562), .Y(q[198]) );
  MUX41X1_HVT U1602 ( .A1(\ram[12][199] ), .A3(\ram[14][199] ), .A2(
        \ram[13][199] ), .A4(\ram[15][199] ), .S0(n528), .S1(n435), .Y(n1401)
         );
  MUX41X1_HVT U1603 ( .A1(\ram[8][199] ), .A3(\ram[10][199] ), .A2(
        \ram[9][199] ), .A4(\ram[11][199] ), .S0(n528), .S1(n435), .Y(n1402)
         );
  MUX41X1_HVT U1604 ( .A1(\ram[4][199] ), .A3(\ram[6][199] ), .A2(
        \ram[5][199] ), .A4(\ram[7][199] ), .S0(n528), .S1(n435), .Y(n1403) );
  MUX41X1_HVT U1605 ( .A1(\ram[0][199] ), .A3(\ram[2][199] ), .A2(
        \ram[1][199] ), .A4(\ram[3][199] ), .S0(n528), .S1(n435), .Y(n1404) );
  MUX41X1_HVT U1606 ( .A1(n1404), .A3(n1402), .A2(n1403), .A4(n1401), .S0(n596), .S1(n562), .Y(q[199]) );
  MUX41X1_HVT U1607 ( .A1(\ram[12][200] ), .A3(\ram[14][200] ), .A2(
        \ram[13][200] ), .A4(\ram[15][200] ), .S0(n528), .S1(n435), .Y(n1405)
         );
  MUX41X1_HVT U1608 ( .A1(\ram[8][200] ), .A3(\ram[10][200] ), .A2(
        \ram[9][200] ), .A4(\ram[11][200] ), .S0(n528), .S1(n435), .Y(n1406)
         );
  MUX41X1_HVT U1609 ( .A1(\ram[4][200] ), .A3(\ram[6][200] ), .A2(
        \ram[5][200] ), .A4(\ram[7][200] ), .S0(n528), .S1(n435), .Y(n1407) );
  MUX41X1_HVT U1610 ( .A1(\ram[0][200] ), .A3(\ram[2][200] ), .A2(
        \ram[1][200] ), .A4(\ram[3][200] ), .S0(n528), .S1(n435), .Y(n1408) );
  MUX41X1_HVT U1611 ( .A1(n1408), .A3(n1406), .A2(n1407), .A4(n1405), .S0(n596), .S1(n563), .Y(q[200]) );
  MUX41X1_HVT U1612 ( .A1(\ram[12][201] ), .A3(\ram[14][201] ), .A2(
        \ram[13][201] ), .A4(\ram[15][201] ), .S0(n529), .S1(n436), .Y(n1409)
         );
  MUX41X1_HVT U1613 ( .A1(\ram[8][201] ), .A3(\ram[10][201] ), .A2(
        \ram[9][201] ), .A4(\ram[11][201] ), .S0(n529), .S1(n436), .Y(n1410)
         );
  MUX41X1_HVT U1614 ( .A1(\ram[4][201] ), .A3(\ram[6][201] ), .A2(
        \ram[5][201] ), .A4(\ram[7][201] ), .S0(n529), .S1(n436), .Y(n1411) );
  MUX41X1_HVT U1615 ( .A1(\ram[0][201] ), .A3(\ram[2][201] ), .A2(
        \ram[1][201] ), .A4(\ram[3][201] ), .S0(n529), .S1(n436), .Y(n1412) );
  MUX41X1_HVT U1616 ( .A1(n1412), .A3(n1410), .A2(n1411), .A4(n1409), .S0(n596), .S1(n563), .Y(q[201]) );
  MUX41X1_HVT U1617 ( .A1(\ram[12][202] ), .A3(\ram[14][202] ), .A2(
        \ram[13][202] ), .A4(\ram[15][202] ), .S0(n529), .S1(n436), .Y(n1413)
         );
  MUX41X1_HVT U1618 ( .A1(\ram[8][202] ), .A3(\ram[10][202] ), .A2(
        \ram[9][202] ), .A4(\ram[11][202] ), .S0(n529), .S1(n436), .Y(n1414)
         );
  MUX41X1_HVT U1619 ( .A1(\ram[4][202] ), .A3(\ram[6][202] ), .A2(
        \ram[5][202] ), .A4(\ram[7][202] ), .S0(n529), .S1(n436), .Y(n1415) );
  MUX41X1_HVT U1620 ( .A1(\ram[0][202] ), .A3(\ram[2][202] ), .A2(
        \ram[1][202] ), .A4(\ram[3][202] ), .S0(n529), .S1(n436), .Y(n1416) );
  MUX41X1_HVT U1621 ( .A1(n1416), .A3(n1414), .A2(n1415), .A4(n1413), .S0(n596), .S1(n563), .Y(q[202]) );
  MUX41X1_HVT U1622 ( .A1(\ram[12][203] ), .A3(\ram[14][203] ), .A2(
        \ram[13][203] ), .A4(\ram[15][203] ), .S0(n529), .S1(n436), .Y(n1417)
         );
  MUX41X1_HVT U1623 ( .A1(\ram[8][203] ), .A3(\ram[10][203] ), .A2(
        \ram[9][203] ), .A4(\ram[11][203] ), .S0(n529), .S1(n436), .Y(n1418)
         );
  MUX41X1_HVT U1624 ( .A1(\ram[4][203] ), .A3(\ram[6][203] ), .A2(
        \ram[5][203] ), .A4(\ram[7][203] ), .S0(n529), .S1(n436), .Y(n1419) );
  MUX41X1_HVT U1625 ( .A1(\ram[0][203] ), .A3(\ram[2][203] ), .A2(
        \ram[1][203] ), .A4(\ram[3][203] ), .S0(n529), .S1(n436), .Y(n1420) );
  MUX41X1_HVT U1626 ( .A1(n1420), .A3(n1418), .A2(n1419), .A4(n1417), .S0(n596), .S1(n563), .Y(q[203]) );
  MUX41X1_HVT U1627 ( .A1(\ram[12][204] ), .A3(\ram[14][204] ), .A2(
        \ram[13][204] ), .A4(\ram[15][204] ), .S0(n530), .S1(n437), .Y(n1421)
         );
  MUX41X1_HVT U1628 ( .A1(\ram[8][204] ), .A3(\ram[10][204] ), .A2(
        \ram[9][204] ), .A4(\ram[11][204] ), .S0(n530), .S1(n437), .Y(n1422)
         );
  MUX41X1_HVT U1629 ( .A1(\ram[4][204] ), .A3(\ram[6][204] ), .A2(
        \ram[5][204] ), .A4(\ram[7][204] ), .S0(n530), .S1(n437), .Y(n1423) );
  MUX41X1_HVT U1630 ( .A1(\ram[0][204] ), .A3(\ram[2][204] ), .A2(
        \ram[1][204] ), .A4(\ram[3][204] ), .S0(n530), .S1(n437), .Y(n1424) );
  MUX41X1_HVT U1631 ( .A1(n1424), .A3(n1422), .A2(n1423), .A4(n1421), .S0(n597), .S1(n563), .Y(q[204]) );
  MUX41X1_HVT U1632 ( .A1(\ram[12][205] ), .A3(\ram[14][205] ), .A2(
        \ram[13][205] ), .A4(\ram[15][205] ), .S0(n530), .S1(n437), .Y(n1425)
         );
  MUX41X1_HVT U1633 ( .A1(\ram[8][205] ), .A3(\ram[10][205] ), .A2(
        \ram[9][205] ), .A4(\ram[11][205] ), .S0(n530), .S1(n437), .Y(n1426)
         );
  MUX41X1_HVT U1634 ( .A1(\ram[4][205] ), .A3(\ram[6][205] ), .A2(
        \ram[5][205] ), .A4(\ram[7][205] ), .S0(n530), .S1(n437), .Y(n1427) );
  MUX41X1_HVT U1635 ( .A1(\ram[0][205] ), .A3(\ram[2][205] ), .A2(
        \ram[1][205] ), .A4(\ram[3][205] ), .S0(n530), .S1(n437), .Y(n1428) );
  MUX41X1_HVT U1636 ( .A1(n1428), .A3(n1426), .A2(n1427), .A4(n1425), .S0(n597), .S1(n563), .Y(q[205]) );
  MUX41X1_HVT U1637 ( .A1(\ram[12][206] ), .A3(\ram[14][206] ), .A2(
        \ram[13][206] ), .A4(\ram[15][206] ), .S0(n530), .S1(n437), .Y(n1429)
         );
  MUX41X1_HVT U1638 ( .A1(\ram[8][206] ), .A3(\ram[10][206] ), .A2(
        \ram[9][206] ), .A4(\ram[11][206] ), .S0(n530), .S1(n437), .Y(n1430)
         );
  MUX41X1_HVT U1639 ( .A1(\ram[4][206] ), .A3(\ram[6][206] ), .A2(
        \ram[5][206] ), .A4(\ram[7][206] ), .S0(n530), .S1(n437), .Y(n1431) );
  MUX41X1_HVT U1640 ( .A1(\ram[0][206] ), .A3(\ram[2][206] ), .A2(
        \ram[1][206] ), .A4(\ram[3][206] ), .S0(n530), .S1(n437), .Y(n1432) );
  MUX41X1_HVT U1641 ( .A1(n1432), .A3(n1430), .A2(n1431), .A4(n1429), .S0(n597), .S1(n563), .Y(q[206]) );
  MUX41X1_HVT U1642 ( .A1(\ram[12][207] ), .A3(\ram[14][207] ), .A2(
        \ram[13][207] ), .A4(\ram[15][207] ), .S0(n531), .S1(n438), .Y(n1433)
         );
  MUX41X1_HVT U1643 ( .A1(\ram[8][207] ), .A3(\ram[10][207] ), .A2(
        \ram[9][207] ), .A4(\ram[11][207] ), .S0(n531), .S1(n438), .Y(n1434)
         );
  MUX41X1_HVT U1644 ( .A1(\ram[4][207] ), .A3(\ram[6][207] ), .A2(
        \ram[5][207] ), .A4(\ram[7][207] ), .S0(n531), .S1(n438), .Y(n1435) );
  MUX41X1_HVT U1645 ( .A1(\ram[0][207] ), .A3(\ram[2][207] ), .A2(
        \ram[1][207] ), .A4(\ram[3][207] ), .S0(n531), .S1(n438), .Y(n1436) );
  MUX41X1_HVT U1646 ( .A1(n1436), .A3(n1434), .A2(n1435), .A4(n1433), .S0(n597), .S1(n563), .Y(q[207]) );
  MUX41X1_HVT U1647 ( .A1(\ram[12][208] ), .A3(\ram[14][208] ), .A2(
        \ram[13][208] ), .A4(\ram[15][208] ), .S0(n531), .S1(n438), .Y(n1437)
         );
  MUX41X1_HVT U1648 ( .A1(\ram[8][208] ), .A3(\ram[10][208] ), .A2(
        \ram[9][208] ), .A4(\ram[11][208] ), .S0(n531), .S1(n438), .Y(n1438)
         );
  MUX41X1_HVT U1649 ( .A1(\ram[4][208] ), .A3(\ram[6][208] ), .A2(
        \ram[5][208] ), .A4(\ram[7][208] ), .S0(n531), .S1(n438), .Y(n1439) );
  MUX41X1_HVT U1650 ( .A1(\ram[0][208] ), .A3(\ram[2][208] ), .A2(
        \ram[1][208] ), .A4(\ram[3][208] ), .S0(n531), .S1(n438), .Y(n1440) );
  MUX41X1_HVT U1651 ( .A1(n1440), .A3(n1438), .A2(n1439), .A4(n1437), .S0(n597), .S1(n563), .Y(q[208]) );
  MUX41X1_HVT U1652 ( .A1(\ram[12][209] ), .A3(\ram[14][209] ), .A2(
        \ram[13][209] ), .A4(\ram[15][209] ), .S0(n531), .S1(n438), .Y(n1441)
         );
  MUX41X1_HVT U1653 ( .A1(\ram[8][209] ), .A3(\ram[10][209] ), .A2(
        \ram[9][209] ), .A4(\ram[11][209] ), .S0(n531), .S1(n438), .Y(n1442)
         );
  MUX41X1_HVT U1654 ( .A1(\ram[4][209] ), .A3(\ram[6][209] ), .A2(
        \ram[5][209] ), .A4(\ram[7][209] ), .S0(n531), .S1(n438), .Y(n1443) );
  MUX41X1_HVT U1655 ( .A1(\ram[0][209] ), .A3(\ram[2][209] ), .A2(
        \ram[1][209] ), .A4(\ram[3][209] ), .S0(n531), .S1(n438), .Y(n1444) );
  MUX41X1_HVT U1656 ( .A1(n1444), .A3(n1442), .A2(n1443), .A4(n1441), .S0(n597), .S1(n563), .Y(q[209]) );
  MUX41X1_HVT U1657 ( .A1(\ram[12][210] ), .A3(\ram[14][210] ), .A2(
        \ram[13][210] ), .A4(\ram[15][210] ), .S0(n532), .S1(n439), .Y(n1445)
         );
  MUX41X1_HVT U1658 ( .A1(\ram[8][210] ), .A3(\ram[10][210] ), .A2(
        \ram[9][210] ), .A4(\ram[11][210] ), .S0(n532), .S1(n439), .Y(n1446)
         );
  MUX41X1_HVT U1659 ( .A1(\ram[4][210] ), .A3(\ram[6][210] ), .A2(
        \ram[5][210] ), .A4(\ram[7][210] ), .S0(n532), .S1(n439), .Y(n1447) );
  MUX41X1_HVT U1660 ( .A1(\ram[0][210] ), .A3(\ram[2][210] ), .A2(
        \ram[1][210] ), .A4(\ram[3][210] ), .S0(n532), .S1(n439), .Y(n1448) );
  MUX41X1_HVT U1661 ( .A1(n1448), .A3(n1446), .A2(n1447), .A4(n1445), .S0(n597), .S1(n563), .Y(q[210]) );
  MUX41X1_HVT U1662 ( .A1(\ram[12][211] ), .A3(\ram[14][211] ), .A2(
        \ram[13][211] ), .A4(\ram[15][211] ), .S0(n532), .S1(n439), .Y(n1449)
         );
  MUX41X1_HVT U1663 ( .A1(\ram[8][211] ), .A3(\ram[10][211] ), .A2(
        \ram[9][211] ), .A4(\ram[11][211] ), .S0(n532), .S1(n439), .Y(n1450)
         );
  MUX41X1_HVT U1664 ( .A1(\ram[4][211] ), .A3(\ram[6][211] ), .A2(
        \ram[5][211] ), .A4(\ram[7][211] ), .S0(n532), .S1(n439), .Y(n1451) );
  MUX41X1_HVT U1665 ( .A1(\ram[0][211] ), .A3(\ram[2][211] ), .A2(
        \ram[1][211] ), .A4(\ram[3][211] ), .S0(n532), .S1(n439), .Y(n1452) );
  MUX41X1_HVT U1666 ( .A1(n1452), .A3(n1450), .A2(n1451), .A4(n1449), .S0(n597), .S1(n563), .Y(q[211]) );
  MUX41X1_HVT U1667 ( .A1(\ram[12][212] ), .A3(\ram[14][212] ), .A2(
        \ram[13][212] ), .A4(\ram[15][212] ), .S0(n532), .S1(n439), .Y(n1453)
         );
  MUX41X1_HVT U1668 ( .A1(\ram[8][212] ), .A3(\ram[10][212] ), .A2(
        \ram[9][212] ), .A4(\ram[11][212] ), .S0(n532), .S1(n439), .Y(n1454)
         );
  MUX41X1_HVT U1669 ( .A1(\ram[4][212] ), .A3(\ram[6][212] ), .A2(
        \ram[5][212] ), .A4(\ram[7][212] ), .S0(n532), .S1(n439), .Y(n1455) );
  MUX41X1_HVT U1670 ( .A1(\ram[0][212] ), .A3(\ram[2][212] ), .A2(
        \ram[1][212] ), .A4(\ram[3][212] ), .S0(n532), .S1(n439), .Y(n1456) );
  MUX41X1_HVT U1671 ( .A1(n1456), .A3(n1454), .A2(n1455), .A4(n1453), .S0(n597), .S1(n564), .Y(q[212]) );
  MUX41X1_HVT U1672 ( .A1(\ram[12][213] ), .A3(\ram[14][213] ), .A2(
        \ram[13][213] ), .A4(\ram[15][213] ), .S0(n533), .S1(n440), .Y(n1457)
         );
  MUX41X1_HVT U1673 ( .A1(\ram[8][213] ), .A3(\ram[10][213] ), .A2(
        \ram[9][213] ), .A4(\ram[11][213] ), .S0(n533), .S1(n440), .Y(n1458)
         );
  MUX41X1_HVT U1674 ( .A1(\ram[4][213] ), .A3(\ram[6][213] ), .A2(
        \ram[5][213] ), .A4(\ram[7][213] ), .S0(n533), .S1(n440), .Y(n1459) );
  MUX41X1_HVT U1675 ( .A1(\ram[0][213] ), .A3(\ram[2][213] ), .A2(
        \ram[1][213] ), .A4(\ram[3][213] ), .S0(n533), .S1(n440), .Y(n1460) );
  MUX41X1_HVT U1676 ( .A1(n1460), .A3(n1458), .A2(n1459), .A4(n1457), .S0(n597), .S1(n564), .Y(q[213]) );
  MUX41X1_HVT U1677 ( .A1(\ram[12][214] ), .A3(\ram[14][214] ), .A2(
        \ram[13][214] ), .A4(\ram[15][214] ), .S0(n533), .S1(n440), .Y(n1461)
         );
  MUX41X1_HVT U1678 ( .A1(\ram[8][214] ), .A3(\ram[10][214] ), .A2(
        \ram[9][214] ), .A4(\ram[11][214] ), .S0(n533), .S1(n440), .Y(n1462)
         );
  MUX41X1_HVT U1679 ( .A1(\ram[4][214] ), .A3(\ram[6][214] ), .A2(
        \ram[5][214] ), .A4(\ram[7][214] ), .S0(n533), .S1(n440), .Y(n1463) );
  MUX41X1_HVT U1680 ( .A1(\ram[0][214] ), .A3(\ram[2][214] ), .A2(
        \ram[1][214] ), .A4(\ram[3][214] ), .S0(n533), .S1(n440), .Y(n1464) );
  MUX41X1_HVT U1681 ( .A1(n1464), .A3(n1462), .A2(n1463), .A4(n1461), .S0(n597), .S1(n564), .Y(q[214]) );
  MUX41X1_HVT U1682 ( .A1(\ram[12][215] ), .A3(\ram[14][215] ), .A2(
        \ram[13][215] ), .A4(\ram[15][215] ), .S0(n533), .S1(n440), .Y(n1465)
         );
  MUX41X1_HVT U1683 ( .A1(\ram[8][215] ), .A3(\ram[10][215] ), .A2(
        \ram[9][215] ), .A4(\ram[11][215] ), .S0(n533), .S1(n440), .Y(n1466)
         );
  MUX41X1_HVT U1684 ( .A1(\ram[4][215] ), .A3(\ram[6][215] ), .A2(
        \ram[5][215] ), .A4(\ram[7][215] ), .S0(n533), .S1(n440), .Y(n1467) );
  MUX41X1_HVT U1685 ( .A1(\ram[0][215] ), .A3(\ram[2][215] ), .A2(
        \ram[1][215] ), .A4(\ram[3][215] ), .S0(n533), .S1(n440), .Y(n1468) );
  MUX41X1_HVT U1686 ( .A1(n1468), .A3(n1466), .A2(n1467), .A4(n1465), .S0(n597), .S1(n564), .Y(q[215]) );
  MUX41X1_HVT U1687 ( .A1(\ram[12][216] ), .A3(\ram[14][216] ), .A2(
        \ram[13][216] ), .A4(\ram[15][216] ), .S0(n534), .S1(n441), .Y(n1469)
         );
  MUX41X1_HVT U1688 ( .A1(\ram[8][216] ), .A3(\ram[10][216] ), .A2(
        \ram[9][216] ), .A4(\ram[11][216] ), .S0(n534), .S1(n441), .Y(n1470)
         );
  MUX41X1_HVT U1689 ( .A1(\ram[4][216] ), .A3(\ram[6][216] ), .A2(
        \ram[5][216] ), .A4(\ram[7][216] ), .S0(n534), .S1(n441), .Y(n1471) );
  MUX41X1_HVT U1690 ( .A1(\ram[0][216] ), .A3(\ram[2][216] ), .A2(
        \ram[1][216] ), .A4(\ram[3][216] ), .S0(n534), .S1(n441), .Y(n1472) );
  MUX41X1_HVT U1691 ( .A1(n1472), .A3(n1470), .A2(n1471), .A4(n1469), .S0(n598), .S1(n564), .Y(q[216]) );
  MUX41X1_HVT U1692 ( .A1(\ram[12][217] ), .A3(\ram[14][217] ), .A2(
        \ram[13][217] ), .A4(\ram[15][217] ), .S0(n534), .S1(n441), .Y(n1473)
         );
  MUX41X1_HVT U1693 ( .A1(\ram[8][217] ), .A3(\ram[10][217] ), .A2(
        \ram[9][217] ), .A4(\ram[11][217] ), .S0(n534), .S1(n441), .Y(n1474)
         );
  MUX41X1_HVT U1694 ( .A1(\ram[4][217] ), .A3(\ram[6][217] ), .A2(
        \ram[5][217] ), .A4(\ram[7][217] ), .S0(n534), .S1(n441), .Y(n1475) );
  MUX41X1_HVT U1695 ( .A1(\ram[0][217] ), .A3(\ram[2][217] ), .A2(
        \ram[1][217] ), .A4(\ram[3][217] ), .S0(n534), .S1(n441), .Y(n1476) );
  MUX41X1_HVT U1696 ( .A1(n1476), .A3(n1474), .A2(n1475), .A4(n1473), .S0(n598), .S1(n564), .Y(q[217]) );
  MUX41X1_HVT U1697 ( .A1(\ram[12][218] ), .A3(\ram[14][218] ), .A2(
        \ram[13][218] ), .A4(\ram[15][218] ), .S0(n534), .S1(n441), .Y(n1477)
         );
  MUX41X1_HVT U1698 ( .A1(\ram[8][218] ), .A3(\ram[10][218] ), .A2(
        \ram[9][218] ), .A4(\ram[11][218] ), .S0(n534), .S1(n441), .Y(n1478)
         );
  MUX41X1_HVT U1699 ( .A1(\ram[4][218] ), .A3(\ram[6][218] ), .A2(
        \ram[5][218] ), .A4(\ram[7][218] ), .S0(n534), .S1(n441), .Y(n1479) );
  MUX41X1_HVT U1700 ( .A1(\ram[0][218] ), .A3(\ram[2][218] ), .A2(
        \ram[1][218] ), .A4(\ram[3][218] ), .S0(n534), .S1(n441), .Y(n1480) );
  MUX41X1_HVT U1701 ( .A1(n1480), .A3(n1478), .A2(n1479), .A4(n1477), .S0(n598), .S1(n564), .Y(q[218]) );
  MUX41X1_HVT U1702 ( .A1(\ram[12][219] ), .A3(\ram[14][219] ), .A2(
        \ram[13][219] ), .A4(\ram[15][219] ), .S0(n535), .S1(n442), .Y(n1481)
         );
  MUX41X1_HVT U1703 ( .A1(\ram[8][219] ), .A3(\ram[10][219] ), .A2(
        \ram[9][219] ), .A4(\ram[11][219] ), .S0(n535), .S1(n442), .Y(n1482)
         );
  MUX41X1_HVT U1704 ( .A1(\ram[4][219] ), .A3(\ram[6][219] ), .A2(
        \ram[5][219] ), .A4(\ram[7][219] ), .S0(n535), .S1(n442), .Y(n1483) );
  MUX41X1_HVT U1705 ( .A1(\ram[0][219] ), .A3(\ram[2][219] ), .A2(
        \ram[1][219] ), .A4(\ram[3][219] ), .S0(n535), .S1(n442), .Y(n1484) );
  MUX41X1_HVT U1706 ( .A1(n1484), .A3(n1482), .A2(n1483), .A4(n1481), .S0(n598), .S1(n564), .Y(q[219]) );
  MUX41X1_HVT U1707 ( .A1(\ram[12][220] ), .A3(\ram[14][220] ), .A2(
        \ram[13][220] ), .A4(\ram[15][220] ), .S0(n535), .S1(n442), .Y(n1485)
         );
  MUX41X1_HVT U1708 ( .A1(\ram[8][220] ), .A3(\ram[10][220] ), .A2(
        \ram[9][220] ), .A4(\ram[11][220] ), .S0(n535), .S1(n442), .Y(n1486)
         );
  MUX41X1_HVT U1709 ( .A1(\ram[4][220] ), .A3(\ram[6][220] ), .A2(
        \ram[5][220] ), .A4(\ram[7][220] ), .S0(n535), .S1(n442), .Y(n1487) );
  MUX41X1_HVT U1710 ( .A1(\ram[0][220] ), .A3(\ram[2][220] ), .A2(
        \ram[1][220] ), .A4(\ram[3][220] ), .S0(n535), .S1(n442), .Y(n1488) );
  MUX41X1_HVT U1711 ( .A1(n1488), .A3(n1486), .A2(n1487), .A4(n1485), .S0(n598), .S1(n564), .Y(q[220]) );
  MUX41X1_HVT U1712 ( .A1(\ram[12][221] ), .A3(\ram[14][221] ), .A2(
        \ram[13][221] ), .A4(\ram[15][221] ), .S0(n535), .S1(n442), .Y(n1489)
         );
  MUX41X1_HVT U1713 ( .A1(\ram[8][221] ), .A3(\ram[10][221] ), .A2(
        \ram[9][221] ), .A4(\ram[11][221] ), .S0(n535), .S1(n442), .Y(n1490)
         );
  MUX41X1_HVT U1714 ( .A1(\ram[4][221] ), .A3(\ram[6][221] ), .A2(
        \ram[5][221] ), .A4(\ram[7][221] ), .S0(n535), .S1(n442), .Y(n1491) );
  MUX41X1_HVT U1715 ( .A1(\ram[0][221] ), .A3(\ram[2][221] ), .A2(
        \ram[1][221] ), .A4(\ram[3][221] ), .S0(n535), .S1(n442), .Y(n1492) );
  MUX41X1_HVT U1716 ( .A1(n1492), .A3(n1490), .A2(n1491), .A4(n1489), .S0(n598), .S1(n564), .Y(q[221]) );
  MUX41X1_HVT U1717 ( .A1(\ram[12][222] ), .A3(\ram[14][222] ), .A2(
        \ram[13][222] ), .A4(\ram[15][222] ), .S0(n536), .S1(n443), .Y(n1493)
         );
  MUX41X1_HVT U1718 ( .A1(\ram[8][222] ), .A3(\ram[10][222] ), .A2(
        \ram[9][222] ), .A4(\ram[11][222] ), .S0(n536), .S1(n443), .Y(n1494)
         );
  MUX41X1_HVT U1719 ( .A1(\ram[4][222] ), .A3(\ram[6][222] ), .A2(
        \ram[5][222] ), .A4(\ram[7][222] ), .S0(n536), .S1(n443), .Y(n1495) );
  MUX41X1_HVT U1720 ( .A1(\ram[0][222] ), .A3(\ram[2][222] ), .A2(
        \ram[1][222] ), .A4(\ram[3][222] ), .S0(n536), .S1(n443), .Y(n1496) );
  MUX41X1_HVT U1721 ( .A1(n1496), .A3(n1494), .A2(n1495), .A4(n1493), .S0(n598), .S1(n564), .Y(q[222]) );
  MUX41X1_HVT U1722 ( .A1(\ram[12][223] ), .A3(\ram[14][223] ), .A2(
        \ram[13][223] ), .A4(\ram[15][223] ), .S0(n536), .S1(n443), .Y(n1497)
         );
  MUX41X1_HVT U1723 ( .A1(\ram[8][223] ), .A3(\ram[10][223] ), .A2(
        \ram[9][223] ), .A4(\ram[11][223] ), .S0(n536), .S1(n443), .Y(n1498)
         );
  MUX41X1_HVT U1724 ( .A1(\ram[4][223] ), .A3(\ram[6][223] ), .A2(
        \ram[5][223] ), .A4(\ram[7][223] ), .S0(n536), .S1(n443), .Y(n1499) );
  MUX41X1_HVT U1725 ( .A1(\ram[0][223] ), .A3(\ram[2][223] ), .A2(
        \ram[1][223] ), .A4(\ram[3][223] ), .S0(n536), .S1(n443), .Y(n1500) );
  MUX41X1_HVT U1726 ( .A1(n1500), .A3(n1498), .A2(n1499), .A4(n1497), .S0(n598), .S1(n564), .Y(q[223]) );
  MUX41X1_HVT U1727 ( .A1(\ram[12][224] ), .A3(\ram[14][224] ), .A2(
        \ram[13][224] ), .A4(\ram[15][224] ), .S0(n536), .S1(n443), .Y(n1501)
         );
  MUX41X1_HVT U1728 ( .A1(\ram[8][224] ), .A3(\ram[10][224] ), .A2(
        \ram[9][224] ), .A4(\ram[11][224] ), .S0(n536), .S1(n443), .Y(n1502)
         );
  MUX41X1_HVT U1729 ( .A1(\ram[4][224] ), .A3(\ram[6][224] ), .A2(
        \ram[5][224] ), .A4(\ram[7][224] ), .S0(n536), .S1(n443), .Y(n1503) );
  MUX41X1_HVT U1730 ( .A1(\ram[0][224] ), .A3(\ram[2][224] ), .A2(
        \ram[1][224] ), .A4(\ram[3][224] ), .S0(n536), .S1(n443), .Y(n1504) );
  MUX41X1_HVT U1731 ( .A1(n1504), .A3(n1502), .A2(n1503), .A4(n1501), .S0(n598), .S1(n565), .Y(q[224]) );
  MUX41X1_HVT U1732 ( .A1(\ram[12][225] ), .A3(\ram[14][225] ), .A2(
        \ram[13][225] ), .A4(\ram[15][225] ), .S0(n537), .S1(n444), .Y(n1505)
         );
  MUX41X1_HVT U1733 ( .A1(\ram[8][225] ), .A3(\ram[10][225] ), .A2(
        \ram[9][225] ), .A4(\ram[11][225] ), .S0(n537), .S1(n444), .Y(n1506)
         );
  MUX41X1_HVT U1734 ( .A1(\ram[4][225] ), .A3(\ram[6][225] ), .A2(
        \ram[5][225] ), .A4(\ram[7][225] ), .S0(n537), .S1(n444), .Y(n1507) );
  MUX41X1_HVT U1735 ( .A1(\ram[0][225] ), .A3(\ram[2][225] ), .A2(
        \ram[1][225] ), .A4(\ram[3][225] ), .S0(n537), .S1(n444), .Y(n1508) );
  MUX41X1_HVT U1736 ( .A1(n1508), .A3(n1506), .A2(n1507), .A4(n1505), .S0(n598), .S1(n565), .Y(q[225]) );
  MUX41X1_HVT U1737 ( .A1(\ram[12][226] ), .A3(\ram[14][226] ), .A2(
        \ram[13][226] ), .A4(\ram[15][226] ), .S0(n537), .S1(n444), .Y(n1509)
         );
  MUX41X1_HVT U1738 ( .A1(\ram[8][226] ), .A3(\ram[10][226] ), .A2(
        \ram[9][226] ), .A4(\ram[11][226] ), .S0(n537), .S1(n444), .Y(n1510)
         );
  MUX41X1_HVT U1739 ( .A1(\ram[4][226] ), .A3(\ram[6][226] ), .A2(
        \ram[5][226] ), .A4(\ram[7][226] ), .S0(n537), .S1(n444), .Y(n1511) );
  MUX41X1_HVT U1740 ( .A1(\ram[0][226] ), .A3(\ram[2][226] ), .A2(
        \ram[1][226] ), .A4(\ram[3][226] ), .S0(n537), .S1(n444), .Y(n1512) );
  MUX41X1_HVT U1741 ( .A1(n1512), .A3(n1510), .A2(n1511), .A4(n1509), .S0(n598), .S1(n565), .Y(q[226]) );
  MUX41X1_HVT U1742 ( .A1(\ram[12][227] ), .A3(\ram[14][227] ), .A2(
        \ram[13][227] ), .A4(\ram[15][227] ), .S0(n537), .S1(n444), .Y(n1513)
         );
  MUX41X1_HVT U1743 ( .A1(\ram[8][227] ), .A3(\ram[10][227] ), .A2(
        \ram[9][227] ), .A4(\ram[11][227] ), .S0(n537), .S1(n444), .Y(n1514)
         );
  MUX41X1_HVT U1744 ( .A1(\ram[4][227] ), .A3(\ram[6][227] ), .A2(
        \ram[5][227] ), .A4(\ram[7][227] ), .S0(n537), .S1(n444), .Y(n1515) );
  MUX41X1_HVT U1745 ( .A1(\ram[0][227] ), .A3(\ram[2][227] ), .A2(
        \ram[1][227] ), .A4(\ram[3][227] ), .S0(n537), .S1(n444), .Y(n1516) );
  MUX41X1_HVT U1746 ( .A1(n1516), .A3(n1514), .A2(n1515), .A4(n1513), .S0(n598), .S1(n565), .Y(q[227]) );
  MUX41X1_HVT U1747 ( .A1(\ram[12][228] ), .A3(\ram[14][228] ), .A2(
        \ram[13][228] ), .A4(\ram[15][228] ), .S0(n538), .S1(n445), .Y(n1517)
         );
  MUX41X1_HVT U1748 ( .A1(\ram[8][228] ), .A3(\ram[10][228] ), .A2(
        \ram[9][228] ), .A4(\ram[11][228] ), .S0(n538), .S1(n445), .Y(n1518)
         );
  MUX41X1_HVT U1749 ( .A1(\ram[4][228] ), .A3(\ram[6][228] ), .A2(
        \ram[5][228] ), .A4(\ram[7][228] ), .S0(n538), .S1(n445), .Y(n1519) );
  MUX41X1_HVT U1750 ( .A1(\ram[0][228] ), .A3(\ram[2][228] ), .A2(
        \ram[1][228] ), .A4(\ram[3][228] ), .S0(n538), .S1(n445), .Y(n1520) );
  MUX41X1_HVT U1751 ( .A1(n1520), .A3(n1518), .A2(n1519), .A4(n1517), .S0(n599), .S1(n565), .Y(q[228]) );
  MUX41X1_HVT U1752 ( .A1(\ram[12][229] ), .A3(\ram[14][229] ), .A2(
        \ram[13][229] ), .A4(\ram[15][229] ), .S0(n538), .S1(n445), .Y(n1521)
         );
  MUX41X1_HVT U1753 ( .A1(\ram[8][229] ), .A3(\ram[10][229] ), .A2(
        \ram[9][229] ), .A4(\ram[11][229] ), .S0(n538), .S1(n445), .Y(n1522)
         );
  MUX41X1_HVT U1754 ( .A1(\ram[4][229] ), .A3(\ram[6][229] ), .A2(
        \ram[5][229] ), .A4(\ram[7][229] ), .S0(n538), .S1(n445), .Y(n1523) );
  MUX41X1_HVT U1755 ( .A1(\ram[0][229] ), .A3(\ram[2][229] ), .A2(
        \ram[1][229] ), .A4(\ram[3][229] ), .S0(n538), .S1(n445), .Y(n1524) );
  MUX41X1_HVT U1756 ( .A1(n1524), .A3(n1522), .A2(n1523), .A4(n1521), .S0(n599), .S1(n565), .Y(q[229]) );
  MUX41X1_HVT U1757 ( .A1(\ram[12][230] ), .A3(\ram[14][230] ), .A2(
        \ram[13][230] ), .A4(\ram[15][230] ), .S0(n538), .S1(n445), .Y(n1525)
         );
  MUX41X1_HVT U1758 ( .A1(\ram[8][230] ), .A3(\ram[10][230] ), .A2(
        \ram[9][230] ), .A4(\ram[11][230] ), .S0(n538), .S1(n445), .Y(n1526)
         );
  MUX41X1_HVT U1759 ( .A1(\ram[4][230] ), .A3(\ram[6][230] ), .A2(
        \ram[5][230] ), .A4(\ram[7][230] ), .S0(n538), .S1(n445), .Y(n1527) );
  MUX41X1_HVT U1760 ( .A1(\ram[0][230] ), .A3(\ram[2][230] ), .A2(
        \ram[1][230] ), .A4(\ram[3][230] ), .S0(n538), .S1(n445), .Y(n1528) );
  MUX41X1_HVT U1761 ( .A1(n1528), .A3(n1526), .A2(n1527), .A4(n1525), .S0(n599), .S1(n565), .Y(q[230]) );
  MUX41X1_HVT U1762 ( .A1(\ram[12][231] ), .A3(\ram[14][231] ), .A2(
        \ram[13][231] ), .A4(\ram[15][231] ), .S0(n539), .S1(n446), .Y(n1529)
         );
  MUX41X1_HVT U1763 ( .A1(\ram[8][231] ), .A3(\ram[10][231] ), .A2(
        \ram[9][231] ), .A4(\ram[11][231] ), .S0(n539), .S1(n446), .Y(n1530)
         );
  MUX41X1_HVT U1764 ( .A1(\ram[4][231] ), .A3(\ram[6][231] ), .A2(
        \ram[5][231] ), .A4(\ram[7][231] ), .S0(n539), .S1(n446), .Y(n1531) );
  MUX41X1_HVT U1765 ( .A1(\ram[0][231] ), .A3(\ram[2][231] ), .A2(
        \ram[1][231] ), .A4(\ram[3][231] ), .S0(n539), .S1(n446), .Y(n1532) );
  MUX41X1_HVT U1766 ( .A1(n1532), .A3(n1530), .A2(n1531), .A4(n1529), .S0(n599), .S1(n565), .Y(q[231]) );
  MUX41X1_HVT U1767 ( .A1(\ram[12][232] ), .A3(\ram[14][232] ), .A2(
        \ram[13][232] ), .A4(\ram[15][232] ), .S0(n539), .S1(n446), .Y(n1533)
         );
  MUX41X1_HVT U1768 ( .A1(\ram[8][232] ), .A3(\ram[10][232] ), .A2(
        \ram[9][232] ), .A4(\ram[11][232] ), .S0(n539), .S1(n446), .Y(n1534)
         );
  MUX41X1_HVT U1769 ( .A1(\ram[4][232] ), .A3(\ram[6][232] ), .A2(
        \ram[5][232] ), .A4(\ram[7][232] ), .S0(n539), .S1(n446), .Y(n1535) );
  MUX41X1_HVT U1770 ( .A1(\ram[0][232] ), .A3(\ram[2][232] ), .A2(
        \ram[1][232] ), .A4(\ram[3][232] ), .S0(n539), .S1(n446), .Y(n1536) );
  MUX41X1_HVT U1771 ( .A1(n1536), .A3(n1534), .A2(n1535), .A4(n1533), .S0(n599), .S1(n565), .Y(q[232]) );
  MUX41X1_HVT U1772 ( .A1(\ram[12][233] ), .A3(\ram[14][233] ), .A2(
        \ram[13][233] ), .A4(\ram[15][233] ), .S0(n539), .S1(n446), .Y(n1537)
         );
  MUX41X1_HVT U1773 ( .A1(\ram[8][233] ), .A3(\ram[10][233] ), .A2(
        \ram[9][233] ), .A4(\ram[11][233] ), .S0(n539), .S1(n446), .Y(n1538)
         );
  MUX41X1_HVT U1774 ( .A1(\ram[4][233] ), .A3(\ram[6][233] ), .A2(
        \ram[5][233] ), .A4(\ram[7][233] ), .S0(n539), .S1(n446), .Y(n1539) );
  MUX41X1_HVT U1775 ( .A1(\ram[0][233] ), .A3(\ram[2][233] ), .A2(
        \ram[1][233] ), .A4(\ram[3][233] ), .S0(n539), .S1(n446), .Y(n1540) );
  MUX41X1_HVT U1776 ( .A1(n1540), .A3(n1538), .A2(n1539), .A4(n1537), .S0(n599), .S1(n565), .Y(q[233]) );
  MUX41X1_HVT U1777 ( .A1(\ram[12][234] ), .A3(\ram[14][234] ), .A2(
        \ram[13][234] ), .A4(\ram[15][234] ), .S0(n540), .S1(n447), .Y(n1541)
         );
  MUX41X1_HVT U1778 ( .A1(\ram[8][234] ), .A3(\ram[10][234] ), .A2(
        \ram[9][234] ), .A4(\ram[11][234] ), .S0(n540), .S1(n447), .Y(n1542)
         );
  MUX41X1_HVT U1779 ( .A1(\ram[4][234] ), .A3(\ram[6][234] ), .A2(
        \ram[5][234] ), .A4(\ram[7][234] ), .S0(n540), .S1(n447), .Y(n1543) );
  MUX41X1_HVT U1780 ( .A1(\ram[0][234] ), .A3(\ram[2][234] ), .A2(
        \ram[1][234] ), .A4(\ram[3][234] ), .S0(n540), .S1(n447), .Y(n1544) );
  MUX41X1_HVT U1781 ( .A1(n1544), .A3(n1542), .A2(n1543), .A4(n1541), .S0(n599), .S1(n565), .Y(q[234]) );
  MUX41X1_HVT U1782 ( .A1(\ram[12][235] ), .A3(\ram[14][235] ), .A2(
        \ram[13][235] ), .A4(\ram[15][235] ), .S0(n540), .S1(n447), .Y(n1545)
         );
  MUX41X1_HVT U1783 ( .A1(\ram[8][235] ), .A3(\ram[10][235] ), .A2(
        \ram[9][235] ), .A4(\ram[11][235] ), .S0(n540), .S1(n447), .Y(n1546)
         );
  MUX41X1_HVT U1784 ( .A1(\ram[4][235] ), .A3(\ram[6][235] ), .A2(
        \ram[5][235] ), .A4(\ram[7][235] ), .S0(n540), .S1(n447), .Y(n1547) );
  MUX41X1_HVT U1785 ( .A1(\ram[0][235] ), .A3(\ram[2][235] ), .A2(
        \ram[1][235] ), .A4(\ram[3][235] ), .S0(n540), .S1(n447), .Y(n1548) );
  MUX41X1_HVT U1786 ( .A1(n1548), .A3(n1546), .A2(n1547), .A4(n1545), .S0(n599), .S1(n565), .Y(q[235]) );
  MUX41X1_HVT U1787 ( .A1(\ram[12][236] ), .A3(\ram[14][236] ), .A2(
        \ram[13][236] ), .A4(\ram[15][236] ), .S0(n540), .S1(n447), .Y(n1549)
         );
  MUX41X1_HVT U1788 ( .A1(\ram[8][236] ), .A3(\ram[10][236] ), .A2(
        \ram[9][236] ), .A4(\ram[11][236] ), .S0(n540), .S1(n447), .Y(n1550)
         );
  MUX41X1_HVT U1789 ( .A1(\ram[4][236] ), .A3(\ram[6][236] ), .A2(
        \ram[5][236] ), .A4(\ram[7][236] ), .S0(n540), .S1(n447), .Y(n1551) );
  MUX41X1_HVT U1790 ( .A1(\ram[0][236] ), .A3(\ram[2][236] ), .A2(
        \ram[1][236] ), .A4(\ram[3][236] ), .S0(n540), .S1(n447), .Y(n1552) );
  MUX41X1_HVT U1791 ( .A1(n1552), .A3(n1550), .A2(n1551), .A4(n1549), .S0(n599), .S1(n566), .Y(q[236]) );
  MUX41X1_HVT U1792 ( .A1(\ram[12][237] ), .A3(\ram[14][237] ), .A2(
        \ram[13][237] ), .A4(\ram[15][237] ), .S0(n541), .S1(n448), .Y(n1553)
         );
  MUX41X1_HVT U1793 ( .A1(\ram[8][237] ), .A3(\ram[10][237] ), .A2(
        \ram[9][237] ), .A4(\ram[11][237] ), .S0(n541), .S1(n448), .Y(n1554)
         );
  MUX41X1_HVT U1794 ( .A1(\ram[4][237] ), .A3(\ram[6][237] ), .A2(
        \ram[5][237] ), .A4(\ram[7][237] ), .S0(n541), .S1(n448), .Y(n1555) );
  MUX41X1_HVT U1795 ( .A1(\ram[0][237] ), .A3(\ram[2][237] ), .A2(
        \ram[1][237] ), .A4(\ram[3][237] ), .S0(n541), .S1(n448), .Y(n1556) );
  MUX41X1_HVT U1796 ( .A1(n1556), .A3(n1554), .A2(n1555), .A4(n1553), .S0(n599), .S1(n566), .Y(q[237]) );
  MUX41X1_HVT U1797 ( .A1(\ram[12][238] ), .A3(\ram[14][238] ), .A2(
        \ram[13][238] ), .A4(\ram[15][238] ), .S0(n541), .S1(n448), .Y(n1557)
         );
  MUX41X1_HVT U1798 ( .A1(\ram[8][238] ), .A3(\ram[10][238] ), .A2(
        \ram[9][238] ), .A4(\ram[11][238] ), .S0(n541), .S1(n448), .Y(n1558)
         );
  MUX41X1_HVT U1799 ( .A1(\ram[4][238] ), .A3(\ram[6][238] ), .A2(
        \ram[5][238] ), .A4(\ram[7][238] ), .S0(n541), .S1(n448), .Y(n1559) );
  MUX41X1_HVT U1800 ( .A1(\ram[0][238] ), .A3(\ram[2][238] ), .A2(
        \ram[1][238] ), .A4(\ram[3][238] ), .S0(n541), .S1(n448), .Y(n1560) );
  MUX41X1_HVT U1801 ( .A1(n1560), .A3(n1558), .A2(n1559), .A4(n1557), .S0(n599), .S1(n566), .Y(q[238]) );
  MUX41X1_HVT U1802 ( .A1(\ram[12][239] ), .A3(\ram[14][239] ), .A2(
        \ram[13][239] ), .A4(\ram[15][239] ), .S0(n541), .S1(n448), .Y(n1561)
         );
  MUX41X1_HVT U1803 ( .A1(\ram[8][239] ), .A3(\ram[10][239] ), .A2(
        \ram[9][239] ), .A4(\ram[11][239] ), .S0(n541), .S1(n448), .Y(n1562)
         );
  MUX41X1_HVT U1804 ( .A1(\ram[4][239] ), .A3(\ram[6][239] ), .A2(
        \ram[5][239] ), .A4(\ram[7][239] ), .S0(n541), .S1(n448), .Y(n1563) );
  MUX41X1_HVT U1805 ( .A1(\ram[0][239] ), .A3(\ram[2][239] ), .A2(
        \ram[1][239] ), .A4(\ram[3][239] ), .S0(n541), .S1(n448), .Y(n1564) );
  MUX41X1_HVT U1806 ( .A1(n1564), .A3(n1562), .A2(n1563), .A4(n1561), .S0(n599), .S1(n566), .Y(q[239]) );
  MUX41X1_HVT U1807 ( .A1(\ram[12][240] ), .A3(\ram[14][240] ), .A2(
        \ram[13][240] ), .A4(\ram[15][240] ), .S0(n542), .S1(n449), .Y(n1565)
         );
  MUX41X1_HVT U1808 ( .A1(\ram[8][240] ), .A3(\ram[10][240] ), .A2(
        \ram[9][240] ), .A4(\ram[11][240] ), .S0(n542), .S1(n449), .Y(n1566)
         );
  MUX41X1_HVT U1809 ( .A1(\ram[4][240] ), .A3(\ram[6][240] ), .A2(
        \ram[5][240] ), .A4(\ram[7][240] ), .S0(n542), .S1(n449), .Y(n1567) );
  MUX41X1_HVT U1810 ( .A1(\ram[0][240] ), .A3(\ram[2][240] ), .A2(
        \ram[1][240] ), .A4(\ram[3][240] ), .S0(n542), .S1(n449), .Y(n1568) );
  MUX41X1_HVT U1811 ( .A1(n1568), .A3(n1566), .A2(n1567), .A4(n1565), .S0(n600), .S1(n566), .Y(q[240]) );
  MUX41X1_HVT U1812 ( .A1(\ram[12][241] ), .A3(\ram[14][241] ), .A2(
        \ram[13][241] ), .A4(\ram[15][241] ), .S0(n542), .S1(n449), .Y(n1569)
         );
  MUX41X1_HVT U1813 ( .A1(\ram[8][241] ), .A3(\ram[10][241] ), .A2(
        \ram[9][241] ), .A4(\ram[11][241] ), .S0(n542), .S1(n449), .Y(n1570)
         );
  MUX41X1_HVT U1814 ( .A1(\ram[4][241] ), .A3(\ram[6][241] ), .A2(
        \ram[5][241] ), .A4(\ram[7][241] ), .S0(n542), .S1(n449), .Y(n1571) );
  MUX41X1_HVT U1815 ( .A1(\ram[0][241] ), .A3(\ram[2][241] ), .A2(
        \ram[1][241] ), .A4(\ram[3][241] ), .S0(n542), .S1(n449), .Y(n1572) );
  MUX41X1_HVT U1816 ( .A1(n1572), .A3(n1570), .A2(n1571), .A4(n1569), .S0(n600), .S1(n566), .Y(q[241]) );
  MUX41X1_HVT U1817 ( .A1(\ram[12][242] ), .A3(\ram[14][242] ), .A2(
        \ram[13][242] ), .A4(\ram[15][242] ), .S0(n542), .S1(n449), .Y(n1573)
         );
  MUX41X1_HVT U1818 ( .A1(\ram[8][242] ), .A3(\ram[10][242] ), .A2(
        \ram[9][242] ), .A4(\ram[11][242] ), .S0(n542), .S1(n449), .Y(n1574)
         );
  MUX41X1_HVT U1819 ( .A1(\ram[4][242] ), .A3(\ram[6][242] ), .A2(
        \ram[5][242] ), .A4(\ram[7][242] ), .S0(n542), .S1(n449), .Y(n1575) );
  MUX41X1_HVT U1820 ( .A1(\ram[0][242] ), .A3(\ram[2][242] ), .A2(
        \ram[1][242] ), .A4(\ram[3][242] ), .S0(n542), .S1(n449), .Y(n1576) );
  MUX41X1_HVT U1821 ( .A1(n1576), .A3(n1574), .A2(n1575), .A4(n1573), .S0(n600), .S1(n566), .Y(q[242]) );
  MUX41X1_HVT U1822 ( .A1(\ram[12][243] ), .A3(\ram[14][243] ), .A2(
        \ram[13][243] ), .A4(\ram[15][243] ), .S0(n543), .S1(n450), .Y(n1577)
         );
  MUX41X1_HVT U1823 ( .A1(\ram[8][243] ), .A3(\ram[10][243] ), .A2(
        \ram[9][243] ), .A4(\ram[11][243] ), .S0(n543), .S1(n450), .Y(n1578)
         );
  MUX41X1_HVT U1824 ( .A1(\ram[4][243] ), .A3(\ram[6][243] ), .A2(
        \ram[5][243] ), .A4(\ram[7][243] ), .S0(n543), .S1(n450), .Y(n1579) );
  MUX41X1_HVT U1825 ( .A1(\ram[0][243] ), .A3(\ram[2][243] ), .A2(
        \ram[1][243] ), .A4(\ram[3][243] ), .S0(n543), .S1(n450), .Y(n1580) );
  MUX41X1_HVT U1826 ( .A1(n1580), .A3(n1578), .A2(n1579), .A4(n1577), .S0(n600), .S1(n566), .Y(q[243]) );
  MUX41X1_HVT U1827 ( .A1(\ram[12][244] ), .A3(\ram[14][244] ), .A2(
        \ram[13][244] ), .A4(\ram[15][244] ), .S0(n543), .S1(n450), .Y(n1581)
         );
  MUX41X1_HVT U1828 ( .A1(\ram[8][244] ), .A3(\ram[10][244] ), .A2(
        \ram[9][244] ), .A4(\ram[11][244] ), .S0(n543), .S1(n450), .Y(n1582)
         );
  MUX41X1_HVT U1829 ( .A1(\ram[4][244] ), .A3(\ram[6][244] ), .A2(
        \ram[5][244] ), .A4(\ram[7][244] ), .S0(n543), .S1(n450), .Y(n1583) );
  MUX41X1_HVT U1830 ( .A1(\ram[0][244] ), .A3(\ram[2][244] ), .A2(
        \ram[1][244] ), .A4(\ram[3][244] ), .S0(n543), .S1(n450), .Y(n1584) );
  MUX41X1_HVT U1831 ( .A1(n1584), .A3(n1582), .A2(n1583), .A4(n1581), .S0(n600), .S1(n566), .Y(q[244]) );
  MUX41X1_HVT U1832 ( .A1(\ram[12][245] ), .A3(\ram[14][245] ), .A2(
        \ram[13][245] ), .A4(\ram[15][245] ), .S0(n543), .S1(n450), .Y(n1585)
         );
  MUX41X1_HVT U1833 ( .A1(\ram[8][245] ), .A3(\ram[10][245] ), .A2(
        \ram[9][245] ), .A4(\ram[11][245] ), .S0(n543), .S1(n450), .Y(n1586)
         );
  MUX41X1_HVT U1834 ( .A1(\ram[4][245] ), .A3(\ram[6][245] ), .A2(
        \ram[5][245] ), .A4(\ram[7][245] ), .S0(n543), .S1(n450), .Y(n1587) );
  MUX41X1_HVT U1835 ( .A1(\ram[0][245] ), .A3(\ram[2][245] ), .A2(
        \ram[1][245] ), .A4(\ram[3][245] ), .S0(n543), .S1(n450), .Y(n1588) );
  MUX41X1_HVT U1836 ( .A1(n1588), .A3(n1586), .A2(n1587), .A4(n1585), .S0(n600), .S1(n566), .Y(q[245]) );
  MUX41X1_HVT U1837 ( .A1(\ram[12][246] ), .A3(\ram[14][246] ), .A2(
        \ram[13][246] ), .A4(\ram[15][246] ), .S0(n544), .S1(n451), .Y(n1589)
         );
  MUX41X1_HVT U1838 ( .A1(\ram[8][246] ), .A3(\ram[10][246] ), .A2(
        \ram[9][246] ), .A4(\ram[11][246] ), .S0(n544), .S1(n451), .Y(n1590)
         );
  MUX41X1_HVT U1839 ( .A1(\ram[4][246] ), .A3(\ram[6][246] ), .A2(
        \ram[5][246] ), .A4(\ram[7][246] ), .S0(n544), .S1(n451), .Y(n1591) );
  MUX41X1_HVT U1840 ( .A1(\ram[0][246] ), .A3(\ram[2][246] ), .A2(
        \ram[1][246] ), .A4(\ram[3][246] ), .S0(n544), .S1(n451), .Y(n1592) );
  MUX41X1_HVT U1841 ( .A1(n1592), .A3(n1590), .A2(n1591), .A4(n1589), .S0(n600), .S1(n566), .Y(q[246]) );
  MUX41X1_HVT U1842 ( .A1(\ram[12][247] ), .A3(\ram[14][247] ), .A2(
        \ram[13][247] ), .A4(\ram[15][247] ), .S0(n544), .S1(n451), .Y(n1593)
         );
  MUX41X1_HVT U1843 ( .A1(\ram[8][247] ), .A3(\ram[10][247] ), .A2(
        \ram[9][247] ), .A4(\ram[11][247] ), .S0(n544), .S1(n451), .Y(n1594)
         );
  MUX41X1_HVT U1844 ( .A1(\ram[4][247] ), .A3(\ram[6][247] ), .A2(
        \ram[5][247] ), .A4(\ram[7][247] ), .S0(n544), .S1(n451), .Y(n1595) );
  MUX41X1_HVT U1845 ( .A1(\ram[0][247] ), .A3(\ram[2][247] ), .A2(
        \ram[1][247] ), .A4(\ram[3][247] ), .S0(n544), .S1(n451), .Y(n1596) );
  MUX41X1_HVT U1846 ( .A1(n1596), .A3(n1594), .A2(n1595), .A4(n1593), .S0(n600), .S1(n566), .Y(q[247]) );
  MUX41X1_HVT U1847 ( .A1(\ram[12][248] ), .A3(\ram[14][248] ), .A2(
        \ram[13][248] ), .A4(\ram[15][248] ), .S0(n544), .S1(n451), .Y(n1597)
         );
  MUX41X1_HVT U1848 ( .A1(\ram[8][248] ), .A3(\ram[10][248] ), .A2(
        \ram[9][248] ), .A4(\ram[11][248] ), .S0(n544), .S1(n451), .Y(n1598)
         );
  MUX41X1_HVT U1849 ( .A1(\ram[4][248] ), .A3(\ram[6][248] ), .A2(
        \ram[5][248] ), .A4(\ram[7][248] ), .S0(n544), .S1(n451), .Y(n1599) );
  MUX41X1_HVT U1850 ( .A1(\ram[0][248] ), .A3(\ram[2][248] ), .A2(
        \ram[1][248] ), .A4(\ram[3][248] ), .S0(n544), .S1(n451), .Y(n1600) );
  MUX41X1_HVT U1851 ( .A1(n1600), .A3(n1598), .A2(n1599), .A4(n1597), .S0(n600), .S1(n567), .Y(q[248]) );
  MUX41X1_HVT U1852 ( .A1(\ram[12][249] ), .A3(\ram[14][249] ), .A2(
        \ram[13][249] ), .A4(\ram[15][249] ), .S0(n545), .S1(n452), .Y(n1601)
         );
  MUX41X1_HVT U1853 ( .A1(\ram[8][249] ), .A3(\ram[10][249] ), .A2(
        \ram[9][249] ), .A4(\ram[11][249] ), .S0(n545), .S1(n452), .Y(n1602)
         );
  MUX41X1_HVT U1854 ( .A1(\ram[4][249] ), .A3(\ram[6][249] ), .A2(
        \ram[5][249] ), .A4(\ram[7][249] ), .S0(n545), .S1(n452), .Y(n1603) );
  MUX41X1_HVT U1855 ( .A1(\ram[0][249] ), .A3(\ram[2][249] ), .A2(
        \ram[1][249] ), .A4(\ram[3][249] ), .S0(n545), .S1(n452), .Y(n1604) );
  MUX41X1_HVT U1856 ( .A1(n1604), .A3(n1602), .A2(n1603), .A4(n1601), .S0(n600), .S1(n567), .Y(q[249]) );
  MUX41X1_HVT U1857 ( .A1(\ram[12][250] ), .A3(\ram[14][250] ), .A2(
        \ram[13][250] ), .A4(\ram[15][250] ), .S0(n545), .S1(n452), .Y(n1605)
         );
  MUX41X1_HVT U1858 ( .A1(\ram[8][250] ), .A3(\ram[10][250] ), .A2(
        \ram[9][250] ), .A4(\ram[11][250] ), .S0(n545), .S1(n452), .Y(n1606)
         );
  MUX41X1_HVT U1859 ( .A1(\ram[4][250] ), .A3(\ram[6][250] ), .A2(
        \ram[5][250] ), .A4(\ram[7][250] ), .S0(n545), .S1(n452), .Y(n1607) );
  MUX41X1_HVT U1860 ( .A1(\ram[0][250] ), .A3(\ram[2][250] ), .A2(
        \ram[1][250] ), .A4(\ram[3][250] ), .S0(n545), .S1(n452), .Y(n1608) );
  MUX41X1_HVT U1861 ( .A1(n1608), .A3(n1606), .A2(n1607), .A4(n1605), .S0(n600), .S1(n567), .Y(q[250]) );
  MUX41X1_HVT U1862 ( .A1(\ram[12][251] ), .A3(\ram[14][251] ), .A2(
        \ram[13][251] ), .A4(\ram[15][251] ), .S0(n545), .S1(n452), .Y(n1609)
         );
  MUX41X1_HVT U1863 ( .A1(\ram[8][251] ), .A3(\ram[10][251] ), .A2(
        \ram[9][251] ), .A4(\ram[11][251] ), .S0(n545), .S1(n452), .Y(n1610)
         );
  MUX41X1_HVT U1864 ( .A1(\ram[4][251] ), .A3(\ram[6][251] ), .A2(
        \ram[5][251] ), .A4(\ram[7][251] ), .S0(n545), .S1(n452), .Y(n1611) );
  MUX41X1_HVT U1865 ( .A1(\ram[0][251] ), .A3(\ram[2][251] ), .A2(
        \ram[1][251] ), .A4(\ram[3][251] ), .S0(n545), .S1(n452), .Y(n1612) );
  MUX41X1_HVT U1866 ( .A1(n1612), .A3(n1610), .A2(n1611), .A4(n1609), .S0(n600), .S1(n567), .Y(q[251]) );
  MUX41X1_HVT U1867 ( .A1(\ram[12][252] ), .A3(\ram[14][252] ), .A2(
        \ram[13][252] ), .A4(\ram[15][252] ), .S0(n546), .S1(n453), .Y(n1613)
         );
  MUX41X1_HVT U1868 ( .A1(\ram[8][252] ), .A3(\ram[10][252] ), .A2(
        \ram[9][252] ), .A4(\ram[11][252] ), .S0(n546), .S1(n453), .Y(n1614)
         );
  MUX41X1_HVT U1869 ( .A1(\ram[4][252] ), .A3(\ram[6][252] ), .A2(
        \ram[5][252] ), .A4(\ram[7][252] ), .S0(n546), .S1(n453), .Y(n1615) );
  MUX41X1_HVT U1870 ( .A1(\ram[0][252] ), .A3(\ram[2][252] ), .A2(
        \ram[1][252] ), .A4(\ram[3][252] ), .S0(n546), .S1(n453), .Y(n1616) );
  MUX41X1_HVT U1871 ( .A1(n1616), .A3(n1614), .A2(n1615), .A4(n1613), .S0(n601), .S1(n567), .Y(q[252]) );
  MUX41X1_HVT U1872 ( .A1(\ram[12][253] ), .A3(\ram[14][253] ), .A2(
        \ram[13][253] ), .A4(\ram[15][253] ), .S0(n546), .S1(n453), .Y(n1617)
         );
  MUX41X1_HVT U1873 ( .A1(\ram[8][253] ), .A3(\ram[10][253] ), .A2(
        \ram[9][253] ), .A4(\ram[11][253] ), .S0(n546), .S1(n453), .Y(n1618)
         );
  MUX41X1_HVT U1874 ( .A1(\ram[4][253] ), .A3(\ram[6][253] ), .A2(
        \ram[5][253] ), .A4(\ram[7][253] ), .S0(n546), .S1(n453), .Y(n1619) );
  MUX41X1_HVT U1875 ( .A1(\ram[0][253] ), .A3(\ram[2][253] ), .A2(
        \ram[1][253] ), .A4(\ram[3][253] ), .S0(n546), .S1(n453), .Y(n1620) );
  MUX41X1_HVT U1876 ( .A1(n1620), .A3(n1618), .A2(n1619), .A4(n1617), .S0(n601), .S1(n567), .Y(q[253]) );
  MUX41X1_HVT U1877 ( .A1(\ram[12][254] ), .A3(\ram[14][254] ), .A2(
        \ram[13][254] ), .A4(\ram[15][254] ), .S0(n546), .S1(n453), .Y(n1621)
         );
  MUX41X1_HVT U1878 ( .A1(\ram[8][254] ), .A3(\ram[10][254] ), .A2(
        \ram[9][254] ), .A4(\ram[11][254] ), .S0(n546), .S1(n453), .Y(n1622)
         );
  MUX41X1_HVT U1879 ( .A1(\ram[4][254] ), .A3(\ram[6][254] ), .A2(
        \ram[5][254] ), .A4(\ram[7][254] ), .S0(n546), .S1(n453), .Y(n1623) );
  MUX41X1_HVT U1880 ( .A1(\ram[0][254] ), .A3(\ram[2][254] ), .A2(
        \ram[1][254] ), .A4(\ram[3][254] ), .S0(n546), .S1(n453), .Y(n1624) );
  MUX41X1_HVT U1881 ( .A1(n1624), .A3(n1622), .A2(n1623), .A4(n1621), .S0(n601), .S1(n567), .Y(q[254]) );
  MUX41X1_HVT U1882 ( .A1(\ram[12][255] ), .A3(\ram[14][255] ), .A2(
        \ram[13][255] ), .A4(\ram[15][255] ), .S0(n547), .S1(n454), .Y(n1625)
         );
  MUX41X1_HVT U1883 ( .A1(\ram[8][255] ), .A3(\ram[10][255] ), .A2(
        \ram[9][255] ), .A4(\ram[11][255] ), .S0(n547), .S1(n454), .Y(n1626)
         );
  MUX41X1_HVT U1884 ( .A1(\ram[4][255] ), .A3(\ram[6][255] ), .A2(
        \ram[5][255] ), .A4(\ram[7][255] ), .S0(n547), .S1(n454), .Y(n1627) );
  MUX41X1_HVT U1885 ( .A1(\ram[0][255] ), .A3(\ram[2][255] ), .A2(
        \ram[1][255] ), .A4(\ram[3][255] ), .S0(n547), .S1(n454), .Y(n1628) );
  MUX41X1_HVT U1886 ( .A1(n1628), .A3(n1626), .A2(n1627), .A4(n1625), .S0(n601), .S1(n567), .Y(q[255]) );
  AND2X1_HVT U1887 ( .A1(data[83]), .A2(n1629), .Y(N99) );
  AND2X1_HVT U1888 ( .A1(data[82]), .A2(n1629), .Y(N98) );
  AND2X1_HVT U1889 ( .A1(data[81]), .A2(n1629), .Y(N97) );
  AND2X1_HVT U1890 ( .A1(data[80]), .A2(n1629), .Y(N96) );
  AND2X1_HVT U1891 ( .A1(data[79]), .A2(n1629), .Y(N95) );
  AND2X1_HVT U1892 ( .A1(data[78]), .A2(n1629), .Y(N94) );
  AND2X1_HVT U1893 ( .A1(data[77]), .A2(n1629), .Y(N93) );
  AND2X1_HVT U1894 ( .A1(data[76]), .A2(n1629), .Y(N92) );
  AND2X1_HVT U1895 ( .A1(data[75]), .A2(n1629), .Y(N91) );
  AND2X1_HVT U1896 ( .A1(data[74]), .A2(n1629), .Y(N90) );
  AND2X1_HVT U1897 ( .A1(data[73]), .A2(n1629), .Y(N89) );
  AND2X1_HVT U1898 ( .A1(data[72]), .A2(n1629), .Y(N88) );
  AND2X1_HVT U1899 ( .A1(data[71]), .A2(n1629), .Y(N87) );
  AND2X1_HVT U1900 ( .A1(data[70]), .A2(n1629), .Y(N86) );
  AND2X1_HVT U1901 ( .A1(data[69]), .A2(n1629), .Y(N85) );
  AND2X1_HVT U1902 ( .A1(data[68]), .A2(n1629), .Y(N84) );
  AND2X1_HVT U1903 ( .A1(data[67]), .A2(n1629), .Y(N83) );
  AND2X1_HVT U1904 ( .A1(data[66]), .A2(n1629), .Y(N82) );
  AND2X1_HVT U1905 ( .A1(data[65]), .A2(n1629), .Y(N81) );
  AND2X1_HVT U1906 ( .A1(data[64]), .A2(n1629), .Y(N80) );
  AND2X1_HVT U1907 ( .A1(data[63]), .A2(n1629), .Y(N79) );
  AND2X1_HVT U1908 ( .A1(data[62]), .A2(n1629), .Y(N78) );
  AND2X1_HVT U1909 ( .A1(data[61]), .A2(n1629), .Y(N77) );
  AND2X1_HVT U1910 ( .A1(data[60]), .A2(n1629), .Y(N76) );
  AND2X1_HVT U1911 ( .A1(data[59]), .A2(n1629), .Y(N75) );
  AND2X1_HVT U1912 ( .A1(data[58]), .A2(n1629), .Y(N74) );
  AND2X1_HVT U1913 ( .A1(data[57]), .A2(n1629), .Y(N73) );
  AND2X1_HVT U1914 ( .A1(data[56]), .A2(n1629), .Y(N72) );
  AND2X1_HVT U1915 ( .A1(data[55]), .A2(n1629), .Y(N71) );
  AND2X1_HVT U1916 ( .A1(data[54]), .A2(n1629), .Y(N70) );
  AND2X1_HVT U1917 ( .A1(data[53]), .A2(n1629), .Y(N69) );
  AND2X1_HVT U1918 ( .A1(data[52]), .A2(n1629), .Y(N68) );
  AND2X1_HVT U1919 ( .A1(data[51]), .A2(n1629), .Y(N67) );
  AND2X1_HVT U1920 ( .A1(data[50]), .A2(n1629), .Y(N66) );
  AND2X1_HVT U1921 ( .A1(data[49]), .A2(n1629), .Y(N65) );
  AND2X1_HVT U1922 ( .A1(data[48]), .A2(n1629), .Y(N64) );
  AND2X1_HVT U1923 ( .A1(data[47]), .A2(n1629), .Y(N63) );
  AND2X1_HVT U1924 ( .A1(data[46]), .A2(n1629), .Y(N62) );
  AND2X1_HVT U1925 ( .A1(data[45]), .A2(n1629), .Y(N61) );
  AND2X1_HVT U1926 ( .A1(data[44]), .A2(n1629), .Y(N60) );
  AND2X1_HVT U1927 ( .A1(data[43]), .A2(n1629), .Y(N59) );
  AND2X1_HVT U1928 ( .A1(data[42]), .A2(n1629), .Y(N58) );
  AND2X1_HVT U1929 ( .A1(data[41]), .A2(n1629), .Y(N57) );
  AND2X1_HVT U1930 ( .A1(data[40]), .A2(n1629), .Y(N56) );
  AND2X1_HVT U1931 ( .A1(data[39]), .A2(n1629), .Y(N55) );
  AND2X1_HVT U1932 ( .A1(data[38]), .A2(n1629), .Y(N54) );
  AND2X1_HVT U1933 ( .A1(data[37]), .A2(n1629), .Y(N53) );
  AND2X1_HVT U1934 ( .A1(data[36]), .A2(n1629), .Y(N52) );
  AND2X1_HVT U1935 ( .A1(data[35]), .A2(n1629), .Y(N51) );
  AND2X1_HVT U1936 ( .A1(data[34]), .A2(n1629), .Y(N50) );
  AND2X1_HVT U1937 ( .A1(data[33]), .A2(n1629), .Y(N49) );
  AND2X1_HVT U1938 ( .A1(data[32]), .A2(n1629), .Y(N48) );
  AND2X1_HVT U1939 ( .A1(data[31]), .A2(n1629), .Y(N47) );
  AND2X1_HVT U1940 ( .A1(data[30]), .A2(n1629), .Y(N46) );
  AND2X1_HVT U1941 ( .A1(data[29]), .A2(n1629), .Y(N45) );
  AND2X1_HVT U1942 ( .A1(data[28]), .A2(n1629), .Y(N44) );
  AND2X1_HVT U1943 ( .A1(data[27]), .A2(n1629), .Y(N43) );
  AND2X1_HVT U1944 ( .A1(data[26]), .A2(n1629), .Y(N42) );
  AND2X1_HVT U1945 ( .A1(data[25]), .A2(n1629), .Y(N41) );
  AND2X1_HVT U1946 ( .A1(data[24]), .A2(n1629), .Y(N40) );
  AND2X1_HVT U1947 ( .A1(data[23]), .A2(n1629), .Y(N39) );
  AND2X1_HVT U1948 ( .A1(data[22]), .A2(n1629), .Y(N38) );
  AND2X1_HVT U1949 ( .A1(data[21]), .A2(n1629), .Y(N37) );
  AND2X1_HVT U1950 ( .A1(data[20]), .A2(n1629), .Y(N36) );
  AND2X1_HVT U1951 ( .A1(data[19]), .A2(n1629), .Y(N35) );
  AND2X1_HVT U1952 ( .A1(data[18]), .A2(n1629), .Y(N34) );
  AND2X1_HVT U1953 ( .A1(data[17]), .A2(n1629), .Y(N33) );
  AND2X1_HVT U1954 ( .A1(data[16]), .A2(n1629), .Y(N32) );
  AO21X1_HVT U1955 ( .A1(n1630), .A2(n1631), .A3(rst), .Y(N318) );
  AO21X1_HVT U1956 ( .A1(n1632), .A2(n1630), .A3(rst), .Y(N315) );
  AO21X1_HVT U1957 ( .A1(n1633), .A2(n1630), .A3(rst), .Y(N312) );
  AND2X1_HVT U1958 ( .A1(data[15]), .A2(n1629), .Y(N31) );
  AO21X1_HVT U1959 ( .A1(n1634), .A2(n1630), .A3(rst), .Y(N309) );
  AND2X1_HVT U1960 ( .A1(n601), .A2(N11), .Y(n1630) );
  AO21X1_HVT U1961 ( .A1(n1635), .A2(n1631), .A3(rst), .Y(N306) );
  AO21X1_HVT U1962 ( .A1(n1635), .A2(n1632), .A3(rst), .Y(N303) );
  AO21X1_HVT U1963 ( .A1(n1635), .A2(n1633), .A3(rst), .Y(N300) );
  AND2X1_HVT U1964 ( .A1(data[14]), .A2(n1629), .Y(N30) );
  AO21X1_HVT U1965 ( .A1(n1635), .A2(n1634), .A3(rst), .Y(N297) );
  AND2X1_HVT U1966 ( .A1(n601), .A2(n578), .Y(n1635) );
  AO21X1_HVT U1967 ( .A1(n1636), .A2(n1631), .A3(rst), .Y(N294) );
  AO21X1_HVT U1968 ( .A1(n1636), .A2(n1632), .A3(rst), .Y(N291) );
  AND2X1_HVT U1969 ( .A1(data[13]), .A2(n1629), .Y(N29) );
  AO21X1_HVT U1970 ( .A1(n1636), .A2(n1633), .A3(rst), .Y(N288) );
  AO21X1_HVT U1971 ( .A1(n1636), .A2(n1634), .A3(rst), .Y(N285) );
  AND2X1_HVT U1972 ( .A1(N11), .A2(n603), .Y(n1636) );
  AO21X1_HVT U1973 ( .A1(n1637), .A2(n1631), .A3(rst), .Y(N282) );
  AND2X1_HVT U1974 ( .A1(n547), .A2(n1638), .Y(n1631) );
  AND2X1_HVT U1975 ( .A1(data[12]), .A2(n1629), .Y(N28) );
  AO21X1_HVT U1976 ( .A1(n1637), .A2(n1632), .A3(rst), .Y(N279) );
  AND2X1_HVT U1977 ( .A1(n1639), .A2(n547), .Y(n1632) );
  AO21X1_HVT U1978 ( .A1(n1637), .A2(n1633), .A3(rst), .Y(N276) );
  AND2X1_HVT U1979 ( .A1(n1638), .A2(n554), .Y(n1633) );
  AND2X1_HVT U1980 ( .A1(n454), .A2(n1629), .Y(n1638) );
  AND2X1_HVT U1981 ( .A1(data[255]), .A2(n1629), .Y(N273) );
  AND2X1_HVT U1982 ( .A1(data[254]), .A2(n1629), .Y(N272) );
  AND2X1_HVT U1983 ( .A1(data[253]), .A2(n1629), .Y(N271) );
  AND2X1_HVT U1984 ( .A1(data[252]), .A2(n1629), .Y(N270) );
  AND2X1_HVT U1985 ( .A1(data[11]), .A2(n1629), .Y(N27) );
  AND2X1_HVT U1986 ( .A1(data[251]), .A2(n1629), .Y(N269) );
  AND2X1_HVT U1987 ( .A1(data[250]), .A2(n1629), .Y(N268) );
  AND2X1_HVT U1988 ( .A1(data[249]), .A2(n1629), .Y(N267) );
  AND2X1_HVT U1989 ( .A1(data[248]), .A2(n1629), .Y(N266) );
  AND2X1_HVT U1990 ( .A1(data[247]), .A2(n1629), .Y(N265) );
  AND2X1_HVT U1991 ( .A1(data[246]), .A2(n1629), .Y(N264) );
  AND2X1_HVT U1992 ( .A1(data[245]), .A2(n1629), .Y(N263) );
  AND2X1_HVT U1993 ( .A1(data[244]), .A2(n1629), .Y(N262) );
  AND2X1_HVT U1994 ( .A1(data[243]), .A2(n1629), .Y(N261) );
  AND2X1_HVT U1995 ( .A1(data[242]), .A2(n1629), .Y(N260) );
  AND2X1_HVT U1996 ( .A1(data[10]), .A2(n1629), .Y(N26) );
  AND2X1_HVT U1997 ( .A1(data[241]), .A2(n1629), .Y(N259) );
  AND2X1_HVT U1998 ( .A1(data[240]), .A2(n1629), .Y(N258) );
  AND2X1_HVT U1999 ( .A1(data[239]), .A2(n1629), .Y(N257) );
  AND2X1_HVT U2000 ( .A1(data[238]), .A2(n1629), .Y(N256) );
  AND2X1_HVT U2001 ( .A1(data[237]), .A2(n1629), .Y(N255) );
  AND2X1_HVT U2002 ( .A1(data[236]), .A2(n1629), .Y(N254) );
  AND2X1_HVT U2003 ( .A1(data[235]), .A2(n1629), .Y(N253) );
  AND2X1_HVT U2004 ( .A1(data[234]), .A2(n1629), .Y(N252) );
  AND2X1_HVT U2005 ( .A1(data[233]), .A2(n1629), .Y(N251) );
  AND2X1_HVT U2006 ( .A1(data[232]), .A2(n1629), .Y(N250) );
  AND2X1_HVT U2007 ( .A1(data[9]), .A2(n1629), .Y(N25) );
  AND2X1_HVT U2008 ( .A1(data[231]), .A2(n1629), .Y(N249) );
  AND2X1_HVT U2009 ( .A1(data[230]), .A2(n1629), .Y(N248) );
  AND2X1_HVT U2010 ( .A1(data[229]), .A2(n1629), .Y(N247) );
  AND2X1_HVT U2011 ( .A1(data[228]), .A2(n1629), .Y(N246) );
  AND2X1_HVT U2012 ( .A1(data[227]), .A2(n1629), .Y(N245) );
  AND2X1_HVT U2013 ( .A1(data[226]), .A2(n1629), .Y(N244) );
  AND2X1_HVT U2014 ( .A1(data[225]), .A2(n1629), .Y(N243) );
  AND2X1_HVT U2015 ( .A1(data[224]), .A2(n1629), .Y(N242) );
  AND2X1_HVT U2016 ( .A1(data[223]), .A2(n1629), .Y(N241) );
  AND2X1_HVT U2017 ( .A1(data[222]), .A2(n1629), .Y(N240) );
  AND2X1_HVT U2018 ( .A1(data[8]), .A2(n1629), .Y(N24) );
  AND2X1_HVT U2019 ( .A1(data[221]), .A2(n1629), .Y(N239) );
  AND2X1_HVT U2020 ( .A1(data[220]), .A2(n1629), .Y(N238) );
  AND2X1_HVT U2021 ( .A1(data[219]), .A2(n1629), .Y(N237) );
  AND2X1_HVT U2022 ( .A1(data[218]), .A2(n1629), .Y(N236) );
  AND2X1_HVT U2023 ( .A1(data[217]), .A2(n1629), .Y(N235) );
  AND2X1_HVT U2024 ( .A1(data[216]), .A2(n1629), .Y(N234) );
  AND2X1_HVT U2025 ( .A1(data[215]), .A2(n1629), .Y(N233) );
  AND2X1_HVT U2026 ( .A1(data[214]), .A2(n1629), .Y(N232) );
  AND2X1_HVT U2027 ( .A1(data[213]), .A2(n1629), .Y(N231) );
  AND2X1_HVT U2028 ( .A1(data[212]), .A2(n1629), .Y(N230) );
  AND2X1_HVT U2029 ( .A1(data[7]), .A2(n1629), .Y(N23) );
  AND2X1_HVT U2030 ( .A1(data[211]), .A2(n1629), .Y(N229) );
  AND2X1_HVT U2031 ( .A1(data[210]), .A2(n1629), .Y(N228) );
  AND2X1_HVT U2032 ( .A1(data[209]), .A2(n1629), .Y(N227) );
  AND2X1_HVT U2033 ( .A1(data[208]), .A2(n1629), .Y(N226) );
  AND2X1_HVT U2034 ( .A1(data[207]), .A2(n1629), .Y(N225) );
  AND2X1_HVT U2035 ( .A1(data[206]), .A2(n1629), .Y(N224) );
  AND2X1_HVT U2036 ( .A1(data[205]), .A2(n1629), .Y(N223) );
  AND2X1_HVT U2037 ( .A1(data[204]), .A2(n1629), .Y(N222) );
  AND2X1_HVT U2038 ( .A1(data[203]), .A2(n1629), .Y(N221) );
  AND2X1_HVT U2039 ( .A1(data[202]), .A2(n1629), .Y(N220) );
  AND2X1_HVT U2040 ( .A1(data[6]), .A2(n1629), .Y(N22) );
  AND2X1_HVT U2041 ( .A1(data[201]), .A2(n1629), .Y(N219) );
  AND2X1_HVT U2042 ( .A1(data[200]), .A2(n1629), .Y(N218) );
  AND2X1_HVT U2043 ( .A1(data[199]), .A2(n1629), .Y(N217) );
  AND2X1_HVT U2044 ( .A1(data[198]), .A2(n1629), .Y(N216) );
  AO21X1_HVT U2045 ( .A1(n1637), .A2(n1634), .A3(rst), .Y(N215) );
  AND2X1_HVT U2046 ( .A1(n1639), .A2(n553), .Y(n1634) );
  AND2X1_HVT U2047 ( .A1(n1629), .A2(n455), .Y(n1639) );
  AND2X1_HVT U2048 ( .A1(n578), .A2(n602), .Y(n1637) );
  AND2X1_HVT U2049 ( .A1(data[197]), .A2(n1629), .Y(N214) );
  AND2X1_HVT U2050 ( .A1(data[196]), .A2(n1629), .Y(N213) );
  AND2X1_HVT U2051 ( .A1(data[195]), .A2(n1629), .Y(N212) );
  AND2X1_HVT U2052 ( .A1(data[194]), .A2(n1629), .Y(N211) );
  AND2X1_HVT U2053 ( .A1(data[193]), .A2(n1629), .Y(N210) );
  AND2X1_HVT U2054 ( .A1(data[5]), .A2(n1629), .Y(N21) );
  AND2X1_HVT U2055 ( .A1(data[192]), .A2(n1629), .Y(N209) );
  AND2X1_HVT U2056 ( .A1(data[191]), .A2(n1629), .Y(N208) );
  AND2X1_HVT U2057 ( .A1(data[190]), .A2(n1629), .Y(N207) );
  AND2X1_HVT U2058 ( .A1(data[189]), .A2(n1629), .Y(N206) );
  AND2X1_HVT U2059 ( .A1(data[188]), .A2(n1629), .Y(N205) );
  AND2X1_HVT U2060 ( .A1(data[187]), .A2(n1629), .Y(N204) );
  AND2X1_HVT U2061 ( .A1(data[186]), .A2(n1629), .Y(N203) );
  AND2X1_HVT U2062 ( .A1(data[185]), .A2(n1629), .Y(N202) );
  AND2X1_HVT U2063 ( .A1(data[184]), .A2(n1629), .Y(N201) );
  AND2X1_HVT U2064 ( .A1(data[183]), .A2(n1629), .Y(N200) );
  AND2X1_HVT U2065 ( .A1(data[4]), .A2(n1629), .Y(N20) );
  AND2X1_HVT U2066 ( .A1(data[182]), .A2(n1629), .Y(N199) );
  AND2X1_HVT U2067 ( .A1(data[181]), .A2(n1629), .Y(N198) );
  AND2X1_HVT U2068 ( .A1(data[180]), .A2(n1629), .Y(N197) );
  AND2X1_HVT U2069 ( .A1(data[179]), .A2(n1629), .Y(N196) );
  AND2X1_HVT U2070 ( .A1(data[178]), .A2(n1629), .Y(N195) );
  AND2X1_HVT U2071 ( .A1(data[177]), .A2(n1629), .Y(N194) );
  AND2X1_HVT U2072 ( .A1(data[176]), .A2(n1629), .Y(N193) );
  AND2X1_HVT U2073 ( .A1(data[175]), .A2(n1629), .Y(N192) );
  AND2X1_HVT U2074 ( .A1(data[174]), .A2(n1629), .Y(N191) );
  AND2X1_HVT U2075 ( .A1(data[173]), .A2(n1629), .Y(N190) );
  AND2X1_HVT U2076 ( .A1(data[3]), .A2(n1629), .Y(N19) );
  AND2X1_HVT U2077 ( .A1(data[172]), .A2(n1629), .Y(N189) );
  AND2X1_HVT U2078 ( .A1(data[171]), .A2(n1629), .Y(N188) );
  AND2X1_HVT U2079 ( .A1(data[170]), .A2(n1629), .Y(N187) );
  AND2X1_HVT U2080 ( .A1(data[169]), .A2(n1629), .Y(N186) );
  AND2X1_HVT U2081 ( .A1(data[168]), .A2(n1629), .Y(N185) );
  AND2X1_HVT U2082 ( .A1(data[167]), .A2(n1629), .Y(N184) );
  AND2X1_HVT U2083 ( .A1(data[166]), .A2(n1629), .Y(N183) );
  AND2X1_HVT U2084 ( .A1(data[165]), .A2(n1629), .Y(N182) );
  AND2X1_HVT U2085 ( .A1(data[164]), .A2(n1629), .Y(N181) );
  AND2X1_HVT U2086 ( .A1(data[163]), .A2(n1629), .Y(N180) );
  AND2X1_HVT U2087 ( .A1(data[2]), .A2(n1629), .Y(N18) );
  AND2X1_HVT U2088 ( .A1(data[162]), .A2(n1629), .Y(N179) );
  AND2X1_HVT U2089 ( .A1(data[161]), .A2(n1629), .Y(N178) );
  AND2X1_HVT U2090 ( .A1(data[160]), .A2(n1629), .Y(N177) );
  AND2X1_HVT U2091 ( .A1(data[159]), .A2(n1629), .Y(N176) );
  AND2X1_HVT U2092 ( .A1(data[158]), .A2(n1629), .Y(N175) );
  AND2X1_HVT U2093 ( .A1(data[157]), .A2(n1629), .Y(N174) );
  AND2X1_HVT U2094 ( .A1(data[156]), .A2(n1629), .Y(N173) );
  AND2X1_HVT U2095 ( .A1(data[155]), .A2(n1629), .Y(N172) );
  AND2X1_HVT U2096 ( .A1(data[154]), .A2(n1629), .Y(N171) );
  AND2X1_HVT U2097 ( .A1(data[153]), .A2(n1629), .Y(N170) );
  AND2X1_HVT U2098 ( .A1(data[1]), .A2(n1629), .Y(N17) );
  AND2X1_HVT U2099 ( .A1(data[152]), .A2(n1629), .Y(N169) );
  AND2X1_HVT U2100 ( .A1(data[151]), .A2(n1629), .Y(N168) );
  AND2X1_HVT U2101 ( .A1(data[150]), .A2(n1629), .Y(N167) );
  AND2X1_HVT U2102 ( .A1(data[149]), .A2(n1629), .Y(N166) );
  AND2X1_HVT U2103 ( .A1(data[148]), .A2(n1629), .Y(N165) );
  AND2X1_HVT U2104 ( .A1(data[147]), .A2(n1629), .Y(N164) );
  AND2X1_HVT U2105 ( .A1(data[146]), .A2(n1629), .Y(N163) );
  AND2X1_HVT U2106 ( .A1(data[145]), .A2(n1629), .Y(N162) );
  AND2X1_HVT U2107 ( .A1(data[144]), .A2(n1629), .Y(N161) );
  AND2X1_HVT U2108 ( .A1(data[143]), .A2(n1629), .Y(N160) );
  AND2X1_HVT U2109 ( .A1(data[0]), .A2(n1629), .Y(N16) );
  AND2X1_HVT U2110 ( .A1(data[142]), .A2(n1629), .Y(N159) );
  AND2X1_HVT U2111 ( .A1(data[141]), .A2(n1629), .Y(N158) );
  AND2X1_HVT U2112 ( .A1(data[140]), .A2(n1629), .Y(N157) );
  AND2X1_HVT U2113 ( .A1(data[139]), .A2(n1629), .Y(N156) );
  AND2X1_HVT U2114 ( .A1(data[138]), .A2(n1629), .Y(N155) );
  AND2X1_HVT U2115 ( .A1(data[137]), .A2(n1629), .Y(N154) );
  AND2X1_HVT U2116 ( .A1(data[136]), .A2(n1629), .Y(N153) );
  AND2X1_HVT U2117 ( .A1(data[135]), .A2(n1629), .Y(N152) );
  AND2X1_HVT U2118 ( .A1(data[134]), .A2(n1629), .Y(N151) );
  AND2X1_HVT U2119 ( .A1(data[133]), .A2(n1629), .Y(N150) );
  AND2X1_HVT U2120 ( .A1(data[132]), .A2(n1629), .Y(N149) );
  AND2X1_HVT U2121 ( .A1(data[131]), .A2(n1629), .Y(N148) );
  AND2X1_HVT U2122 ( .A1(data[130]), .A2(n1629), .Y(N147) );
  AND2X1_HVT U2123 ( .A1(data[129]), .A2(n1629), .Y(N146) );
  AND2X1_HVT U2124 ( .A1(data[128]), .A2(n1629), .Y(N145) );
  AND2X1_HVT U2125 ( .A1(data[127]), .A2(n1629), .Y(N144) );
  AND2X1_HVT U2126 ( .A1(data[126]), .A2(n1629), .Y(N143) );
  AND2X1_HVT U2127 ( .A1(data[125]), .A2(n1629), .Y(N142) );
  AND2X1_HVT U2128 ( .A1(data[124]), .A2(n1629), .Y(N141) );
  AND2X1_HVT U2129 ( .A1(data[123]), .A2(n1629), .Y(N140) );
  AND2X1_HVT U2130 ( .A1(data[122]), .A2(n1629), .Y(N139) );
  AND2X1_HVT U2131 ( .A1(data[121]), .A2(n1629), .Y(N138) );
  AND2X1_HVT U2132 ( .A1(data[120]), .A2(n1629), .Y(N137) );
  AND2X1_HVT U2133 ( .A1(data[119]), .A2(n1629), .Y(N136) );
  AND2X1_HVT U2134 ( .A1(data[118]), .A2(n1629), .Y(N135) );
  AND2X1_HVT U2135 ( .A1(data[117]), .A2(n1629), .Y(N134) );
  AND2X1_HVT U2136 ( .A1(data[116]), .A2(n1629), .Y(N133) );
  AND2X1_HVT U2137 ( .A1(data[115]), .A2(n1629), .Y(N132) );
  AND2X1_HVT U2138 ( .A1(data[114]), .A2(n1629), .Y(N131) );
  AND2X1_HVT U2139 ( .A1(data[113]), .A2(n1629), .Y(N130) );
  AND2X1_HVT U2140 ( .A1(data[112]), .A2(n1629), .Y(N129) );
  AND2X1_HVT U2141 ( .A1(data[111]), .A2(n1629), .Y(N128) );
  AND2X1_HVT U2142 ( .A1(data[110]), .A2(n1629), .Y(N127) );
  AND2X1_HVT U2143 ( .A1(data[109]), .A2(n1629), .Y(N126) );
  AND2X1_HVT U2144 ( .A1(data[108]), .A2(n1629), .Y(N125) );
  AND2X1_HVT U2145 ( .A1(data[107]), .A2(n1629), .Y(N124) );
  AND2X1_HVT U2146 ( .A1(data[106]), .A2(n1629), .Y(N123) );
  AND2X1_HVT U2147 ( .A1(data[105]), .A2(n1629), .Y(N122) );
  AND2X1_HVT U2148 ( .A1(data[104]), .A2(n1629), .Y(N121) );
  AND2X1_HVT U2149 ( .A1(data[103]), .A2(n1629), .Y(N120) );
  AND2X1_HVT U2150 ( .A1(data[102]), .A2(n1629), .Y(N119) );
  AND2X1_HVT U2151 ( .A1(data[101]), .A2(n1629), .Y(N118) );
  AND2X1_HVT U2152 ( .A1(data[100]), .A2(n1629), .Y(N117) );
  AND2X1_HVT U2153 ( .A1(data[99]), .A2(n1629), .Y(N116) );
  AND2X1_HVT U2154 ( .A1(data[98]), .A2(n1629), .Y(N114) );
  AND2X1_HVT U2155 ( .A1(data[97]), .A2(n1629), .Y(N113) );
  AND2X1_HVT U2156 ( .A1(data[96]), .A2(n1629), .Y(N112) );
  AND2X1_HVT U2157 ( .A1(data[95]), .A2(n1629), .Y(N111) );
  AND2X1_HVT U2158 ( .A1(data[94]), .A2(n1629), .Y(N110) );
  AND2X1_HVT U2159 ( .A1(data[93]), .A2(n1629), .Y(N109) );
  AND2X1_HVT U2160 ( .A1(data[92]), .A2(n1629), .Y(N108) );
  AND2X1_HVT U2161 ( .A1(data[91]), .A2(n1629), .Y(N107) );
  AND2X1_HVT U2162 ( .A1(data[90]), .A2(n1629), .Y(N106) );
  AND2X1_HVT U2163 ( .A1(data[89]), .A2(n1629), .Y(N105) );
  AND2X1_HVT U2164 ( .A1(data[88]), .A2(n1629), .Y(N104) );
  AND2X1_HVT U2165 ( .A1(data[87]), .A2(n1629), .Y(N103) );
  AND2X1_HVT U2166 ( .A1(data[86]), .A2(n1629), .Y(N102) );
  AND2X1_HVT U2167 ( .A1(data[85]), .A2(n1629), .Y(N101) );
  AND2X1_HVT U2168 ( .A1(data[84]), .A2(n1629), .Y(N100) );
  AND2X1_HVT U2169 ( .A1(we), .A2(n1640), .Y(n1629) );
  INVX0_HVT U2170 ( .A(rst), .Y(n1640) );
endmodule

