
module inv_sbox_8 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n36, n196, n197, n198, n199, n200, n201, n202, n203, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626;

  NAND2X0_HVT U3 ( .A1(n282), .A2(n284), .Y(n624) );
  NAND2X0_HVT U5 ( .A1(n623), .A2(n303), .Y(n622) );
  NAND2X0_HVT U6 ( .A1(n351), .A2(n626), .Y(n620) );
  NAND2X0_HVT U7 ( .A1(n351), .A2(n346), .Y(n619) );
  NAND2X0_HVT U8 ( .A1(n354), .A2(n621), .Y(n618) );
  NAND2X0_HVT U9 ( .A1(n349), .A2(n618), .Y(n617) );
  NAND2X0_HVT U10 ( .A1(n349), .A2(n615), .Y(n616) );
  NAND2X0_HVT U12 ( .A1(n260), .A2(n337), .Y(n613) );
  NAND2X0_HVT U13 ( .A1(n347), .A2(n295), .Y(n612) );
  NAND2X0_HVT U15 ( .A1(n343), .A2(n352), .Y(n610) );
  NAND2X0_HVT U19 ( .A1(n259), .A2(n416), .Y(n605) );
  NAND2X0_HVT U25 ( .A1(in[6]), .A2(n414), .Y(n621) );
  NAND2X0_HVT U32 ( .A1(n326), .A2(n356), .Y(n593) );
  NAND2X0_HVT U35 ( .A1(n618), .A2(n417), .Y(n591) );
  NAND2X0_HVT U38 ( .A1(n337), .A2(n263), .Y(n588) );
  OA21X1_HVT U53 ( .A1(n362), .A2(n576), .A3(n387), .Y(n574) );
  NAND2X0_HVT U55 ( .A1(n347), .A2(n623), .Y(n572) );
  MUX41X1_HVT U56 ( .A1(n311), .A3(n293), .A2(n385), .A4(n306), .S0(n332), 
        .S1(n272), .Y(n571) );
  AO21X1_HVT U60 ( .A1(n566), .A2(n334), .A3(n604), .Y(n567) );
  MUX41X1_HVT U65 ( .A1(n378), .A3(n380), .A2(n379), .A4(n588), .S0(n330), 
        .S1(n227), .Y(n561) );
  NAND2X0_HVT U66 ( .A1(n353), .A2(n284), .Y(n560) );
  MUX41X1_HVT U67 ( .A1(n375), .A3(n398), .A2(n377), .A4(n560), .S0(n336), 
        .S1(n329), .Y(n559) );
  MUX41X1_HVT U68 ( .A1(n375), .A3(n282), .A2(n376), .A4(n349), .S0(n330), 
        .S1(n359), .Y(n558) );
  MUX41X1_HVT U71 ( .A1(n620), .A3(n415), .A2(n614), .A4(n371), .S0(n330), 
        .S1(n359), .Y(n556) );
  NAND2X0_HVT U72 ( .A1(n344), .A2(n619), .Y(n555) );
  MUX41X1_HVT U73 ( .A1(n598), .A3(n555), .A2(n399), .A4(n337), .S0(n335), 
        .S1(n328), .Y(n554) );
  NAND2X0_HVT U81 ( .A1(n220), .A2(n619), .Y(n546) );
  AND2X1_HVT U82 ( .A1(n620), .A2(n347), .Y(n545) );
  MUX41X1_HVT U84 ( .A1(n319), .A3(n388), .A2(n403), .A4(n600), .S0(n330), 
        .S1(n299), .Y(n543) );
  MUX41X1_HVT U87 ( .A1(n366), .A3(n319), .A2(n404), .A4(n385), .S0(n357), 
        .S1(n272), .Y(n541) );
  MUX41X1_HVT U88 ( .A1(n377), .A3(n363), .A2(n595), .A4(n580), .S0(n330), 
        .S1(n272), .Y(n540) );
  NAND2X0_HVT U89 ( .A1(n356), .A2(n413), .Y(n539) );
  MUX41X1_HVT U90 ( .A1(n415), .A3(n619), .A2(n579), .A4(n539), .S0(n330), 
        .S1(n272), .Y(n538) );
  MUX41X1_HVT U95 ( .A1(n534), .A3(n540), .A2(n538), .A4(n541), .S0(n341), 
        .S1(n310), .Y(n533) );
  MUX41X1_HVT U99 ( .A1(n593), .A3(n379), .A2(n578), .A4(n344), .S0(n334), 
        .S1(n329), .Y(n529) );
  NAND2X0_HVT U100 ( .A1(n263), .A2(n203), .Y(n528) );
  MUX41X1_HVT U101 ( .A1(n407), .A3(n613), .A2(n323), .A4(n528), .S0(n359), 
        .S1(n327), .Y(n527) );
  MUX41X1_HVT U102 ( .A1(n527), .A3(n530), .A2(n529), .A4(n532), .S0(n341), 
        .S1(n310), .Y(n526) );
  AND2X1_HVT U104 ( .A1(n619), .A2(n303), .Y(n525) );
  MUX41X1_HVT U107 ( .A1(n407), .A3(n624), .A2(n523), .A4(n368), .S0(n330), 
        .S1(n227), .Y(n522) );
  MUX41X1_HVT U108 ( .A1(n381), .A3(n293), .A2(n385), .A4(n222), .S0(n283), 
        .S1(n360), .Y(n521) );
  MUX41X1_HVT U109 ( .A1(n406), .A3(n363), .A2(n403), .A4(n396), .S0(n330), 
        .S1(n272), .Y(n520) );
  NAND2X0_HVT U114 ( .A1(n349), .A2(n619), .Y(n515) );
  MUX41X1_HVT U115 ( .A1(n515), .A3(n614), .A2(n393), .A4(n347), .S0(n227), 
        .S1(n329), .Y(n514) );
  MUX41X1_HVT U116 ( .A1(n392), .A3(n388), .A2(n363), .A4(n610), .S0(n327), 
        .S1(n360), .Y(n513) );
  NAND2X0_HVT U118 ( .A1(n356), .A2(n282), .Y(n511) );
  MUX41X1_HVT U119 ( .A1(n409), .A3(n512), .A2(n589), .A4(n511), .S0(n283), 
        .S1(n359), .Y(n510) );
  MUX41X1_HVT U122 ( .A1(n397), .A3(n314), .A2(n580), .A4(n400), .S0(n357), 
        .S1(n227), .Y(n508) );
  MUX41X1_HVT U124 ( .A1(n317), .A3(n507), .A2(n266), .A4(n383), .S0(n334), 
        .S1(n327), .Y(n506) );
  AOI21X1_HVT U127 ( .A1(n333), .A2(n502), .A3(n369), .Y(n503) );
  NAND2X0_HVT U129 ( .A1(n332), .A2(n349), .Y(n500) );
  MUX41X1_HVT U130 ( .A1(n500), .A3(n501), .A2(n504), .A4(n503), .S0(n336), 
        .S1(n339), .Y(n499) );
  AND2X1_HVT U131 ( .A1(n325), .A2(n263), .Y(n498) );
  MUX41X1_HVT U132 ( .A1(n367), .A3(n498), .A2(n411), .A4(n375), .S0(n335), 
        .S1(n328), .Y(n497) );
  MUX41X1_HVT U133 ( .A1(n412), .A3(n368), .A2(n306), .A4(n312), .S0(n334), 
        .S1(n327), .Y(n496) );
  MUX41X1_HVT U136 ( .A1(n577), .A3(n528), .A2(n494), .A4(n373), .S0(n332), 
        .S1(n227), .Y(n493) );
  MUX41X1_HVT U137 ( .A1(n295), .A3(n596), .A2(n600), .A4(n405), .S0(n336), 
        .S1(n327), .Y(n492) );
  MUX41X1_HVT U139 ( .A1(n491), .A3(n495), .A2(n499), .A4(n505), .S0(in[5]), 
        .S1(n281), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n390), .A3(n315), .A2(n304), .A4(n614), .S0(n335), 
        .S1(n329), .Y(n490) );
  NAND2X0_HVT U141 ( .A1(n293), .A2(n263), .Y(n489) );
  MUX41X1_HVT U142 ( .A1(n489), .A3(n587), .A2(n410), .A4(n307), .S0(n333), 
        .S1(n227), .Y(n488) );
  MUX41X1_HVT U143 ( .A1(n413), .A3(n394), .A2(n605), .A4(n602), .S0(n331), 
        .S1(n272), .Y(n487) );
  MUX41X1_HVT U145 ( .A1(n594), .A3(n408), .A2(n486), .A4(n546), .S0(n333), 
        .S1(n272), .Y(n485) );
  AO21X1_HVT U148 ( .A1(n336), .A2(n370), .A3(n203), .Y(n482) );
  MUX41X1_HVT U151 ( .A1(n402), .A3(n391), .A2(n382), .A4(n480), .S0(n334), 
        .S1(n327), .Y(n479) );
  MUX41X1_HVT U155 ( .A1(n304), .A3(n614), .A2(n606), .A4(n386), .S0(n331), 
        .S1(n359), .Y(n475) );
  NAND2X0_HVT U159 ( .A1(n471), .A2(n470), .Y(n472) );
  NAND2X0_HVT U163 ( .A1(n354), .A2(n413), .Y(n466) );
  MUX41X1_HVT U164 ( .A1(n617), .A3(n466), .A2(n589), .A4(n381), .S0(n327), 
        .S1(n336), .Y(n465) );
  NAND2X0_HVT U166 ( .A1(n615), .A2(n462), .Y(n463) );
  MUX41X1_HVT U173 ( .A1(n349), .A3(n415), .A2(n220), .A4(n590), .S0(n331), 
        .S1(n227), .Y(n455) );
  NAND2X0_HVT U177 ( .A1(n260), .A2(n282), .Y(n452) );
  MUX41X1_HVT U178 ( .A1(n318), .A3(n452), .A2(n415), .A4(n582), .S0(n331), 
        .S1(n359), .Y(n451) );
  AND2X1_HVT U179 ( .A1(n620), .A2(n345), .Y(n450) );
  MUX41X1_HVT U180 ( .A1(n593), .A3(n287), .A2(n450), .A4(n581), .S0(n331), 
        .S1(n336), .Y(n449) );
  AND2X1_HVT U185 ( .A1(n417), .A2(n263), .Y(n444) );
  MUX41X1_HVT U190 ( .A1(n441), .A3(n442), .A2(n440), .A4(n443), .S0(n280), 
        .S1(n328), .Y(n439) );
  NAND2X0_HVT U191 ( .A1(n362), .A2(n374), .Y(n438) );
  AND2X1_HVT U192 ( .A1(n297), .A2(n436), .Y(n437) );
  NAND2X0_HVT U194 ( .A1(n584), .A2(n436), .Y(n434) );
  MUX41X1_HVT U195 ( .A1(n435), .A3(n434), .A2(n437), .A4(n438), .S0(n330), 
        .S1(n280), .Y(n433) );
  NAND2X0_HVT U198 ( .A1(n353), .A2(n292), .Y(n615) );
  NAND2X0_HVT U200 ( .A1(n345), .A2(n356), .Y(n502) );
  NAND2X0_HVT U207 ( .A1(n263), .A2(n415), .Y(n566) );
  MUX21X2_HVT U1 ( .A1(n536), .A2(n535), .S0(n36), .Y(n534) );
  IBUFFX16_HVT U2 ( .A(n332), .Y(n36) );
  XNOR2X1_HVT U4 ( .A1(n196), .A2(n325), .Y(n609) );
  IBUFFX16_HVT U11 ( .A(n414), .Y(n196) );
  INVX1_HVT U14 ( .A(n225), .Y(n459) );
  MUX41X1_HVT U16 ( .A1(n454), .A3(n456), .A2(n455), .A4(n458), .S0(n250), 
        .S1(n197), .Y(n453) );
  IBUFFX16_HVT U17 ( .A(n251), .Y(n197) );
  MUX21X1_HVT U18 ( .A1(n282), .A2(n345), .S0(n324), .Y(n531) );
  IBUFFX2_HVT U20 ( .A(n355), .Y(n354) );
  MUX21X2_HVT U21 ( .A1(n472), .A2(n473), .S0(n333), .Y(n469) );
  MUX41X1_HVT U22 ( .A1(n404), .A3(n412), .A2(n572), .A4(n296), .S0(n227), 
        .S1(n283), .Y(n454) );
  INVX0_HVT U23 ( .A(n426), .Y(n404) );
  MUX21X2_HVT U24 ( .A1(n258), .A2(n348), .S0(n260), .Y(n257) );
  NBUFFX2_HVT U26 ( .A(n609), .Y(n343) );
  MUX21X1_HVT U27 ( .A1(n417), .A2(n345), .S0(n352), .Y(n297) );
  INVX1_HVT U28 ( .A(n355), .Y(n352) );
  AO21X2_HVT U29 ( .A1(n354), .A2(n202), .A3(n362), .Y(n436) );
  XNOR2X1_HVT U30 ( .A1(n222), .A2(n354), .Y(n315) );
  MUX21X2_HVT U31 ( .A1(n446), .A2(n447), .S0(n310), .Y(n445) );
  NBUFFX4_HVT U33 ( .A(n414), .Y(n337) );
  INVX0_HVT U34 ( .A(n366), .Y(n198) );
  INVX1_HVT U36 ( .A(n298), .Y(n199) );
  INVX1_HVT U37 ( .A(n298), .Y(n200) );
  INVX1_HVT U39 ( .A(n298), .Y(n201) );
  INVX1_HVT U40 ( .A(n199), .Y(n202) );
  INVX1_HVT U41 ( .A(n200), .Y(n203) );
  INVX1_HVT U42 ( .A(n201), .Y(n218) );
  IBUFFX2_HVT U43 ( .A(n625), .Y(n219) );
  INVX1_HVT U44 ( .A(n219), .Y(n220) );
  INVX0_HVT U45 ( .A(n219), .Y(n221) );
  INVX0_HVT U46 ( .A(n219), .Y(n222) );
  MUX21X2_HVT U47 ( .A1(n497), .A2(n496), .S0(n338), .Y(n495) );
  INVX0_HVT U48 ( .A(n623), .Y(n366) );
  NAND2X0_HVT U49 ( .A1(n414), .A2(n418), .Y(n625) );
  IBUFFX2_HVT U50 ( .A(n625), .Y(n298) );
  INVX1_HVT U51 ( .A(n338), .Y(n339) );
  INVX1_HVT U52 ( .A(n604), .Y(n381) );
  OA21X1_HVT U54 ( .A1(n365), .A2(n362), .A3(n604), .Y(n551) );
  INVX0_HVT U57 ( .A(n583), .Y(n394) );
  INVX1_HVT U58 ( .A(n355), .Y(n259) );
  INVX1_HVT U59 ( .A(n287), .Y(n614) );
  MUX41X1_HVT U61 ( .A1(n571), .A3(n565), .A2(n573), .A4(n569), .S0(n223), 
        .S1(n224), .Y(n564) );
  IBUFFX16_HVT U62 ( .A(n341), .Y(n223) );
  IBUFFX16_HVT U63 ( .A(n309), .Y(n224) );
  INVX1_HVT U64 ( .A(n418), .Y(n325) );
  INVX1_HVT U69 ( .A(in[6]), .Y(n418) );
  MUX21X1_HVT U70 ( .A1(n626), .A2(n226), .S0(n350), .Y(n225) );
  IBUFFX16_HVT U74 ( .A(n416), .Y(n226) );
  INVX1_HVT U75 ( .A(n348), .Y(n415) );
  MUX21X1_HVT U76 ( .A1(n284), .A2(n345), .S0(n356), .Y(n596) );
  IBUFFX2_HVT U77 ( .A(in[0]), .Y(n356) );
  IBUFFX2_HVT U78 ( .A(n361), .Y(n227) );
  INVX1_HVT U79 ( .A(n361), .Y(n299) );
  NAND2X1_HVT U80 ( .A1(n519), .A2(n228), .Y(n229) );
  NAND2X0_HVT U83 ( .A1(n509), .A2(n268), .Y(n230) );
  NAND2X0_HVT U85 ( .A1(n229), .A2(n230), .Y(out[3]) );
  IBUFFX2_HVT U86 ( .A(n268), .Y(n228) );
  MUX41X1_HVT U91 ( .A1(n556), .A3(n553), .A2(n554), .A4(n550), .S0(n340), 
        .S1(n232), .Y(n549) );
  IBUFFX2_HVT U92 ( .A(n260), .Y(n247) );
  INVX1_HVT U93 ( .A(n597), .Y(n387) );
  MUX21X2_HVT U94 ( .A1(n552), .A2(n551), .S0(n333), .Y(n550) );
  INVX0_HVT U96 ( .A(in[5]), .Y(n340) );
  INVX1_HVT U97 ( .A(n267), .Y(n232) );
  MUX41X1_HVT U98 ( .A1(n521), .A3(n524), .A2(n520), .A4(n522), .S0(n231), 
        .S1(n253), .Y(n519) );
  IBUFFX16_HVT U103 ( .A(n252), .Y(n231) );
  MUX41X1_HVT U105 ( .A1(n516), .A3(n513), .A2(n514), .A4(n510), .S0(n233), 
        .S1(n234), .Y(n509) );
  IBUFFX16_HVT U106 ( .A(n341), .Y(n233) );
  IBUFFX16_HVT U110 ( .A(n339), .Y(n234) );
  AO21X2_HVT U111 ( .A1(n393), .A2(n335), .A3(n601), .Y(n517) );
  MUX41X1_HVT U112 ( .A1(n544), .A3(n543), .A2(n548), .A4(n547), .S0(n240), 
        .S1(n239), .Y(n542) );
  MUX41X1_HVT U113 ( .A1(n388), .A3(n257), .A2(n607), .A4(n608), .S0(n359), 
        .S1(n357), .Y(n548) );
  IBUFFX2_HVT U117 ( .A(n340), .Y(n239) );
  IBUFFX2_HVT U120 ( .A(n280), .Y(n240) );
  INVX1_HVT U121 ( .A(n596), .Y(n388) );
  IBUFFX2_HVT U123 ( .A(n361), .Y(n272) );
  IBUFFX4_HVT U125 ( .A(n361), .Y(n360) );
  MUX41X1_HVT U126 ( .A1(n461), .A3(n467), .A2(n465), .A4(n469), .S0(n341), 
        .S1(n267), .Y(n460) );
  NAND2X0_HVT U128 ( .A1(n463), .A2(n235), .Y(n236) );
  NAND2X0_HVT U134 ( .A1(n464), .A2(n332), .Y(n237) );
  NAND2X0_HVT U135 ( .A1(n236), .A2(n237), .Y(n461) );
  IBUFFX2_HVT U138 ( .A(n332), .Y(n235) );
  INVX1_HVT U144 ( .A(n248), .Y(n457) );
  MUX41X1_HVT U146 ( .A1(n316), .A3(n459), .A2(n318), .A4(n317), .S0(n238), 
        .S1(n322), .Y(n458) );
  IBUFFX16_HVT U147 ( .A(n242), .Y(n238) );
  NAND2X0_HVT U149 ( .A1(n449), .A2(n254), .Y(n255) );
  MUX41X1_HVT U150 ( .A1(n389), .A3(n545), .A2(n546), .A4(n402), .S0(n241), 
        .S1(n272), .Y(n544) );
  IBUFFX16_HVT U152 ( .A(n330), .Y(n241) );
  NBUFFX2_HVT U153 ( .A(n308), .Y(n242) );
  INVX1_HVT U154 ( .A(n335), .Y(n308) );
  INVX0_HVT U156 ( .A(n293), .Y(n258) );
  INVX0_HVT U157 ( .A(n257), .Y(n594) );
  NAND2X0_HVT U158 ( .A1(n349), .A2(n243), .Y(n244) );
  NAND2X0_HVT U160 ( .A1(n244), .A2(n198), .Y(n611) );
  IBUFFX2_HVT U161 ( .A(n260), .Y(n243) );
  INVX1_HVT U162 ( .A(n355), .Y(n260) );
  MUX41X1_HVT U165 ( .A1(n490), .A3(n488), .A2(n487), .A4(n485), .S0(n245), 
        .S1(n246), .Y(n484) );
  IBUFFX16_HVT U167 ( .A(n310), .Y(n245) );
  IBUFFX16_HVT U168 ( .A(n341), .Y(n246) );
  MUX21X1_HVT U169 ( .A1(n413), .A2(n415), .S0(n247), .Y(n597) );
  MUX41X1_HVT U170 ( .A1(n313), .A3(n591), .A2(n380), .A4(n468), .S0(n359), 
        .S1(n331), .Y(n467) );
  MUX21X1_HVT U171 ( .A1(n348), .A2(n249), .S0(n352), .Y(n248) );
  IBUFFX16_HVT U172 ( .A(n321), .Y(n249) );
  MUX41X1_HVT U174 ( .A1(n316), .A3(n603), .A2(n539), .A4(n457), .S0(n357), 
        .S1(n242), .Y(n456) );
  IBUFFX16_HVT U175 ( .A(n340), .Y(n250) );
  IBUFFX16_HVT U176 ( .A(n280), .Y(n251) );
  NAND2X0_HVT U181 ( .A1(n557), .A2(n268), .Y(n285) );
  IBUFFX16_HVT U182 ( .A(in[5]), .Y(n252) );
  IBUFFX16_HVT U183 ( .A(n339), .Y(n253) );
  NAND2X0_HVT U184 ( .A1(n451), .A2(n339), .Y(n256) );
  NAND2X0_HVT U186 ( .A1(n255), .A2(n256), .Y(n448) );
  IBUFFX2_HVT U187 ( .A(n339), .Y(n254) );
  INVX2_HVT U188 ( .A(n357), .Y(n322) );
  AO21X1_HVT U189 ( .A1(n263), .A2(n349), .A3(n362), .Y(n470) );
  INVX2_HVT U193 ( .A(n418), .Y(n284) );
  INVX1_HVT U196 ( .A(in[4]), .Y(n361) );
  INVX1_HVT U197 ( .A(in[4]), .Y(n362) );
  MUX41X1_HVT U199 ( .A1(n584), .A3(n381), .A2(n311), .A4(n394), .S0(n261), 
        .S1(n262), .Y(n446) );
  IBUFFX16_HVT U201 ( .A(n334), .Y(n261) );
  IBUFFX16_HVT U202 ( .A(n328), .Y(n262) );
  INVX0_HVT U203 ( .A(n355), .Y(n351) );
  INVX1_HVT U204 ( .A(n355), .Y(n353) );
  INVX1_HVT U205 ( .A(n355), .Y(n350) );
  INVX1_HVT U206 ( .A(n584), .Y(n368) );
  INVX0_HVT U208 ( .A(in[0]), .Y(n263) );
  INVX0_HVT U209 ( .A(in[0]), .Y(n355) );
  NBUFFX16_HVT U210 ( .A(n299), .Y(n336) );
  MUX21X1_HVT U211 ( .A1(n386), .A2(n376), .S0(n336), .Y(n575) );
  NBUFFX2_HVT U212 ( .A(n299), .Y(n334) );
  MUX21X1_HVT U213 ( .A1(n369), .A2(n585), .S0(n336), .Y(n518) );
  MUX21X2_HVT U214 ( .A1(n517), .A2(n518), .S0(n333), .Y(n516) );
  OA21X2_HVT U215 ( .A1(n388), .A2(n362), .A3(n566), .Y(n440) );
  OA21X2_HVT U216 ( .A1(n364), .A2(n362), .A3(n372), .Y(n477) );
  AO21X2_HVT U217 ( .A1(n344), .A2(n623), .A3(n362), .Y(n462) );
  MUX21X1_HVT U218 ( .A1(n444), .A2(n401), .S0(n334), .Y(n443) );
  MUX21X1_HVT U219 ( .A1(n411), .A2(n367), .S0(n334), .Y(n483) );
  NAND2X0_HVT U220 ( .A1(n453), .A2(n268), .Y(n269) );
  INVX1_HVT U221 ( .A(n339), .Y(n271) );
  MUX21X1_HVT U222 ( .A1(n585), .A2(n399), .S0(n308), .Y(n441) );
  INVX1_HVT U223 ( .A(n361), .Y(n359) );
  INVX0_HVT U224 ( .A(n608), .Y(n377) );
  INVX1_HVT U225 ( .A(n268), .Y(n281) );
  INVX1_HVT U226 ( .A(in[7]), .Y(n268) );
  INVX1_HVT U227 ( .A(in[3]), .Y(n414) );
  INVX0_HVT U228 ( .A(n292), .Y(n293) );
  INVX1_HVT U229 ( .A(n343), .Y(n292) );
  INVX1_HVT U230 ( .A(n325), .Y(n326) );
  INVX1_HVT U231 ( .A(n336), .Y(n273) );
  INVX1_HVT U232 ( .A(n322), .Y(n283) );
  INVX1_HVT U233 ( .A(n309), .Y(n267) );
  MUX21X2_HVT U234 ( .A1(n568), .A2(n567), .S0(n332), .Y(n565) );
  MUX21X2_HVT U235 ( .A1(n574), .A2(n575), .S0(n322), .Y(n573) );
  INVX1_HVT U236 ( .A(n598), .Y(n386) );
  NAND2X0_HVT U237 ( .A1(n474), .A2(n268), .Y(n264) );
  NAND2X0_HVT U238 ( .A1(n484), .A2(n281), .Y(n265) );
  NAND2X0_HVT U239 ( .A1(n264), .A2(n265), .Y(out[5]) );
  INVX0_HVT U240 ( .A(n383), .Y(n266) );
  INVX1_HVT U241 ( .A(n602), .Y(n383) );
  MUX41X1_HVT U242 ( .A1(n448), .A3(n445), .A2(n439), .A4(n433), .S0(n340), 
        .S1(n268), .Y(out[7]) );
  NAND2X0_HVT U243 ( .A1(n460), .A2(n281), .Y(n270) );
  NAND2X0_HVT U244 ( .A1(n269), .A2(n270), .Y(out[6]) );
  MUX41X1_HVT U245 ( .A1(n481), .A3(n476), .A2(n479), .A4(n475), .S0(n340), 
        .S1(n271), .Y(n474) );
  MUX21X2_HVT U246 ( .A1(n483), .A2(n482), .S0(n332), .Y(n481) );
  NAND2X0_HVT U247 ( .A1(n319), .A2(n273), .Y(n274) );
  NAND2X0_HVT U248 ( .A1(n578), .A2(n336), .Y(n275) );
  NAND2X0_HVT U249 ( .A1(n274), .A2(n275), .Y(n442) );
  XOR2X1_HVT U250 ( .A1(n303), .A2(n259), .Y(n578) );
  MUX41X1_HVT U251 ( .A1(n611), .A3(n546), .A2(n408), .A4(n525), .S0(n227), 
        .S1(n283), .Y(n524) );
  INVX1_HVT U252 ( .A(n422), .Y(n408) );
  NAND2X0_HVT U253 ( .A1(n506), .A2(n309), .Y(n276) );
  NAND2X0_HVT U254 ( .A1(n508), .A2(n280), .Y(n277) );
  NAND2X0_HVT U255 ( .A1(n276), .A2(n277), .Y(n505) );
  IBUFFX2_HVT U256 ( .A(n338), .Y(n280) );
  NAND2X2_HVT U257 ( .A1(n526), .A2(n268), .Y(n278) );
  NAND2X0_HVT U258 ( .A1(n533), .A2(n281), .Y(n279) );
  NAND2X0_HVT U259 ( .A1(n278), .A2(n279), .Y(out[2]) );
  MUX21X1_HVT U260 ( .A1(n202), .A2(n282), .S0(n350), .Y(n602) );
  MUX21X1_HVT U261 ( .A1(n621), .A2(n321), .S0(n356), .Y(n311) );
  MUX41X1_HVT U262 ( .A1(n405), .A3(n386), .A2(n612), .A4(n398), .S0(n322), 
        .S1(n362), .Y(n532) );
  NAND2X0_HVT U263 ( .A1(n220), .A2(n351), .Y(n623) );
  MUX21X1_HVT U264 ( .A1(n384), .A2(n570), .S0(n320), .Y(n569) );
  MUX21X1_HVT U265 ( .A1(n337), .A2(n416), .S0(n351), .Y(n583) );
  XOR2X1_HVT U266 ( .A1(n348), .A2(n353), .Y(n589) );
  MUX21X1_HVT U267 ( .A1(n284), .A2(n415), .S0(n350), .Y(n601) );
  INVX1_HVT U268 ( .A(n294), .Y(n585) );
  MUX21X1_HVT U269 ( .A1(n347), .A2(n222), .S0(n353), .Y(n607) );
  MUX21X1_HVT U270 ( .A1(n307), .A2(n622), .S0(n333), .Y(n570) );
  MUX21X1_HVT U271 ( .A1(n395), .A2(n317), .S0(n334), .Y(n435) );
  MUX21X1_HVT U272 ( .A1(n346), .A2(n345), .S0(n263), .Y(n468) );
  INVX0_HVT U273 ( .A(n338), .Y(n310) );
  INVX1_HVT U274 ( .A(n310), .Y(n309) );
  MUX21X1_HVT U275 ( .A1(n337), .A2(n343), .S0(n263), .Y(n604) );
  NBUFFX2_HVT U276 ( .A(in[3]), .Y(n282) );
  MUX21X1_HVT U277 ( .A1(n344), .A2(n415), .S0(n356), .Y(n426) );
  OR2X1_HVT U278 ( .A1(n414), .A2(n284), .Y(n626) );
  INVX1_HVT U279 ( .A(n419), .Y(n412) );
  NAND2X0_HVT U280 ( .A1(n564), .A2(n281), .Y(n286) );
  NAND2X0_HVT U281 ( .A1(n285), .A2(n286), .Y(out[0]) );
  INVX1_HVT U282 ( .A(n313), .Y(n582) );
  MUX21X1_HVT U283 ( .A1(n348), .A2(n303), .S0(n324), .Y(n313) );
  AND2X1_HVT U284 ( .A1(n356), .A2(n221), .Y(n287) );
  NAND2X0_HVT U285 ( .A1(n417), .A2(n356), .Y(n288) );
  NAND2X0_HVT U286 ( .A1(n218), .A2(n350), .Y(n289) );
  NAND2X0_HVT U287 ( .A1(n288), .A2(n289), .Y(n603) );
  INVX0_HVT U288 ( .A(n603), .Y(n382) );
  NAND2X0_HVT U289 ( .A1(n549), .A2(n281), .Y(n290) );
  NAND2X0_HVT U290 ( .A1(n542), .A2(n268), .Y(n291) );
  NAND2X0_HVT U291 ( .A1(n290), .A2(n291), .Y(out[1]) );
  INVX0_HVT U292 ( .A(n622), .Y(n367) );
  MUX21X1_HVT U293 ( .A1(n417), .A2(n202), .S0(n324), .Y(n592) );
  INVX1_HVT U294 ( .A(n429), .Y(n401) );
  MUX21X1_HVT U295 ( .A1(n346), .A2(n321), .S0(n324), .Y(n294) );
  INVX0_HVT U296 ( .A(n370), .Y(n295) );
  INVX0_HVT U297 ( .A(n618), .Y(n370) );
  INVX0_HVT U298 ( .A(n344), .Y(n296) );
  INVX1_HVT U299 ( .A(n302), .Y(n552) );
  INVX1_HVT U300 ( .A(n340), .Y(n341) );
  MUX21X1_HVT U301 ( .A1(n623), .A2(n382), .S0(n322), .Y(n563) );
  NAND2X0_HVT U302 ( .A1(n359), .A2(n602), .Y(n300) );
  NAND2X0_HVT U303 ( .A1(n599), .A2(n273), .Y(n301) );
  NAND2X0_HVT U304 ( .A1(n300), .A2(n301), .Y(n464) );
  MUX21X2_HVT U305 ( .A1(n400), .A2(n583), .S0(n308), .Y(n473) );
  IBUFFX2_HVT U306 ( .A(n607), .Y(n378) );
  MUX21X1_HVT U307 ( .A1(n593), .A2(n430), .S0(n308), .Y(n302) );
  INVX1_HVT U308 ( .A(n342), .Y(n417) );
  IBUFFX2_HVT U309 ( .A(n601), .Y(n384) );
  INVX1_HVT U310 ( .A(n624), .Y(n416) );
  MUX41X1_HVT U311 ( .A1(n597), .A3(n391), .A2(n406), .A4(n531), .S0(n322), 
        .S1(n273), .Y(n530) );
  MUX21X1_HVT U312 ( .A1(n337), .A2(n416), .S0(n356), .Y(n430) );
  NBUFFX2_HVT U313 ( .A(n621), .Y(n303) );
  MUX41X1_HVT U314 ( .A1(n381), .A3(n297), .A2(n390), .A4(n616), .S0(n362), 
        .S1(n322), .Y(n553) );
  INVX1_HVT U315 ( .A(n600), .Y(n304) );
  INVX1_HVT U316 ( .A(n307), .Y(n600) );
  MUX41X1_HVT U317 ( .A1(n622), .A3(n617), .A2(n311), .A4(n401), .S0(n322), 
        .S1(n242), .Y(n547) );
  INVX0_HVT U318 ( .A(n572), .Y(n305) );
  INVX1_HVT U319 ( .A(n305), .Y(n306) );
  MUX21X1_HVT U320 ( .A1(n292), .A2(n284), .S0(n351), .Y(n307) );
  INVX1_HVT U321 ( .A(n621), .Y(n413) );
  INVX1_HVT U322 ( .A(n431), .Y(n399) );
  INVX1_HVT U323 ( .A(n592), .Y(n390) );
  MUX41X1_HVT U324 ( .A1(n562), .A3(n559), .A2(n561), .A4(n558), .S0(n340), 
        .S1(n309), .Y(n557) );
  INVX0_HVT U325 ( .A(n620), .Y(n312) );
  OR2X1_HVT U326 ( .A1(n312), .A2(n342), .Y(n584) );
  MUX21X2_HVT U327 ( .A1(n477), .A2(n478), .S0(n333), .Y(n476) );
  MUX21X2_HVT U328 ( .A1(n381), .A2(n563), .S0(n320), .Y(n562) );
  MUX21X1_HVT U329 ( .A1(n600), .A2(n319), .S0(n335), .Y(n478) );
  INVX0_HVT U330 ( .A(n351), .Y(n324) );
  INVX0_HVT U331 ( .A(in[1]), .Y(n338) );
  AND2X1_HVT U332 ( .A1(n221), .A2(n610), .Y(n314) );
  MUX21X1_HVT U333 ( .A1(n296), .A2(n337), .S0(n354), .Y(n587) );
  MUX21X1_HVT U334 ( .A1(n537), .A2(n346), .S0(n350), .Y(n536) );
  MUX21X1_HVT U335 ( .A1(n371), .A2(n293), .S0(n336), .Y(n535) );
  MUX21X1_HVT U336 ( .A1(n343), .A2(n326), .S0(n335), .Y(n537) );
  MUX21X1_HVT U337 ( .A1(n326), .A2(n413), .S0(n259), .Y(n480) );
  MUX21X1_HVT U338 ( .A1(n321), .A2(n221), .S0(n352), .Y(n523) );
  MUX21X1_HVT U339 ( .A1(n296), .A2(n326), .S0(n260), .Y(n421) );
  MUX21X1_HVT U340 ( .A1(n321), .A2(n344), .S0(n259), .Y(n586) );
  MUX21X1_HVT U341 ( .A1(n383), .A2(n306), .S0(n335), .Y(n568) );
  XOR2X1_HVT U342 ( .A1(n342), .A2(n353), .Y(n580) );
  MUX21X1_HVT U343 ( .A1(n592), .A2(n314), .S0(n333), .Y(n501) );
  MUX21X1_HVT U344 ( .A1(n410), .A2(n315), .S0(n332), .Y(n504) );
  MUX21X1_HVT U345 ( .A1(n303), .A2(n220), .S0(n260), .Y(n420) );
  MUX21X1_HVT U346 ( .A1(n337), .A2(n221), .S0(n259), .Y(n429) );
  MUX21X1_HVT U347 ( .A1(n321), .A2(n218), .S0(n352), .Y(n599) );
  MUX21X1_HVT U348 ( .A1(n346), .A2(n337), .S0(n350), .Y(n606) );
  MUX21X1_HVT U349 ( .A1(n337), .A2(n202), .S0(n352), .Y(n595) );
  INVX0_HVT U350 ( .A(n323), .Y(n590) );
  XOR2X1_HVT U351 ( .A1(n347), .A2(n352), .Y(n579) );
  AND2X1_HVT U352 ( .A1(n620), .A2(n222), .Y(n316) );
  MUX21X1_HVT U353 ( .A1(n337), .A2(n346), .S0(n259), .Y(n423) );
  AND2X1_HVT U354 ( .A1(n353), .A2(n321), .Y(n317) );
  NBUFFX2_HVT U355 ( .A(n299), .Y(n335) );
  NBUFFX2_HVT U356 ( .A(n609), .Y(n344) );
  NBUFFX2_HVT U357 ( .A(n609), .Y(n342) );
  AND2X1_HVT U358 ( .A1(n416), .A2(n356), .Y(n318) );
  MUX21X1_HVT U359 ( .A1(n203), .A2(n416), .S0(n354), .Y(n576) );
  AND2X1_HVT U360 ( .A1(n347), .A2(n263), .Y(n319) );
  MUX21X1_HVT U361 ( .A1(n220), .A2(n303), .S0(n259), .Y(n486) );
  NBUFFX2_HVT U362 ( .A(n624), .Y(n347) );
  NBUFFX2_HVT U363 ( .A(n624), .Y(n346) );
  NBUFFX2_HVT U364 ( .A(n621), .Y(n345) );
  NBUFFX2_HVT U365 ( .A(n358), .Y(n331) );
  NBUFFX2_HVT U366 ( .A(n358), .Y(n333) );
  NBUFFX2_HVT U367 ( .A(n358), .Y(n332) );
  XNOR2X1_HVT U368 ( .A1(n362), .A2(n357), .Y(n320) );
  NBUFFX2_HVT U369 ( .A(n358), .Y(n328) );
  NBUFFX2_HVT U370 ( .A(n357), .Y(n330) );
  NBUFFX2_HVT U371 ( .A(n328), .Y(n329) );
  NBUFFX2_HVT U372 ( .A(n358), .Y(n327) );
  MUX21X1_HVT U373 ( .A1(n416), .A2(n413), .S0(n259), .Y(n512) );
  MUX21X1_HVT U374 ( .A1(n415), .A2(n282), .S0(n354), .Y(n419) );
  MUX21X1_HVT U375 ( .A1(n321), .A2(n282), .S0(n260), .Y(n598) );
  MUX21X1_HVT U376 ( .A1(n492), .A2(n493), .S0(n310), .Y(n491) );
  MUX21X1_HVT U377 ( .A1(n282), .A2(n349), .S0(n352), .Y(n425) );
  MUX21X1_HVT U378 ( .A1(n282), .A2(n303), .S0(n354), .Y(n424) );
  MUX21X1_HVT U379 ( .A1(n349), .A2(n282), .S0(n350), .Y(n471) );
  NBUFFX2_HVT U380 ( .A(in[2]), .Y(n358) );
  NBUFFX2_HVT U381 ( .A(in[2]), .Y(n357) );
  NBUFFX2_HVT U382 ( .A(n326), .Y(n321) );
  NBUFFX2_HVT U383 ( .A(n626), .Y(n349) );
  NBUFFX2_HVT U384 ( .A(n626), .Y(n348) );
  MUX41X1_HVT U385 ( .A1(n402), .A3(n366), .A2(n623), .A4(n368), .S0(n322), 
        .S1(n242), .Y(n447) );
  MUX21X1_HVT U386 ( .A1(n344), .A2(n284), .S0(n324), .Y(n323) );
  MUX21X1_HVT U387 ( .A1(n337), .A2(n292), .S0(n352), .Y(n428) );
  INVX1_HVT U388 ( .A(n428), .Y(n402) );
  MUX21X1_HVT U389 ( .A1(n337), .A2(n321), .S0(n351), .Y(n581) );
  MUX21X1_HVT U390 ( .A1(n203), .A2(n321), .S0(n353), .Y(n431) );
  MUX21X1_HVT U391 ( .A1(n347), .A2(n321), .S0(n350), .Y(n507) );
  MUX21X1_HVT U392 ( .A1(n218), .A2(n325), .S0(n353), .Y(n494) );
  XOR2X1_HVT U393 ( .A1(n354), .A2(n325), .Y(n577) );
  MUX21X1_HVT U394 ( .A1(n325), .A2(n347), .S0(n260), .Y(n432) );
  MUX21X1_HVT U395 ( .A1(n346), .A2(n284), .S0(n350), .Y(n427) );
  MUX21X1_HVT U396 ( .A1(n337), .A2(n284), .S0(n353), .Y(n422) );
  MUX21X1_HVT U397 ( .A1(n284), .A2(n348), .S0(n259), .Y(n608) );
  INVX0_HVT U398 ( .A(n588), .Y(n363) );
  INVX0_HVT U399 ( .A(n528), .Y(n364) );
  INVX0_HVT U400 ( .A(n489), .Y(n365) );
  INVX0_HVT U401 ( .A(n619), .Y(n369) );
  INVX0_HVT U402 ( .A(n591), .Y(n371) );
  INVX0_HVT U403 ( .A(n612), .Y(n372) );
  INVX0_HVT U404 ( .A(n617), .Y(n373) );
  INVX0_HVT U405 ( .A(n613), .Y(n374) );
  INVX0_HVT U406 ( .A(n611), .Y(n375) );
  INVX0_HVT U407 ( .A(n610), .Y(n376) );
  INVX0_HVT U408 ( .A(n606), .Y(n379) );
  INVX0_HVT U409 ( .A(n605), .Y(n380) );
  INVX0_HVT U410 ( .A(n599), .Y(n385) );
  INVX0_HVT U411 ( .A(n595), .Y(n389) );
  INVX0_HVT U412 ( .A(n589), .Y(n391) );
  INVX0_HVT U413 ( .A(n587), .Y(n392) );
  INVX0_HVT U414 ( .A(n586), .Y(n393) );
  INVX0_HVT U415 ( .A(n581), .Y(n395) );
  INVX0_HVT U416 ( .A(n580), .Y(n396) );
  INVX0_HVT U417 ( .A(n616), .Y(n397) );
  INVX0_HVT U418 ( .A(n432), .Y(n398) );
  INVX0_HVT U419 ( .A(n430), .Y(n400) );
  INVX0_HVT U420 ( .A(n427), .Y(n403) );
  INVX0_HVT U421 ( .A(n425), .Y(n405) );
  INVX0_HVT U422 ( .A(n424), .Y(n406) );
  INVX0_HVT U423 ( .A(n423), .Y(n407) );
  INVX0_HVT U424 ( .A(n471), .Y(n409) );
  INVX0_HVT U425 ( .A(n421), .Y(n410) );
  INVX0_HVT U426 ( .A(n420), .Y(n411) );
endmodule

