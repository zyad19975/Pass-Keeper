
module inv_sbox_10 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n196, n197, n198, n199, n200, n201, n202, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638;

  NAND2X0_HVT U1 ( .A1(n291), .A2(n344), .Y(n638) );
  NAND2X0_HVT U5 ( .A1(n635), .A2(n299), .Y(n634) );
  NAND2X0_HVT U7 ( .A1(n359), .A2(n636), .Y(n631) );
  NAND2X0_HVT U8 ( .A1(n270), .A2(n351), .Y(n630) );
  NAND2X0_HVT U9 ( .A1(n355), .A2(n630), .Y(n629) );
  NAND2X0_HVT U10 ( .A1(n354), .A2(n627), .Y(n628) );
  NAND2X0_HVT U11 ( .A1(n294), .A2(n313), .Y(n626) );
  NAND2X0_HVT U12 ( .A1(n270), .A2(n341), .Y(n625) );
  NAND2X0_HVT U13 ( .A1(n353), .A2(n305), .Y(n624) );
  NAND2X0_HVT U15 ( .A1(n300), .A2(n271), .Y(n622) );
  NAND2X0_HVT U19 ( .A1(n267), .A2(n301), .Y(n617) );
  NAND2X0_HVT U32 ( .A1(n344), .A2(n277), .Y(n605) );
  NAND2X0_HVT U35 ( .A1(n630), .A2(n322), .Y(n602) );
  NAND2X0_HVT U38 ( .A1(n341), .A2(n277), .Y(n599) );
  NAND2X0_HVT U42 ( .A1(n632), .A2(n428), .Y(n595) );
  OA21X1_HVT U53 ( .A1(n279), .A2(n587), .A3(n395), .Y(n585) );
  NAND2X0_HVT U55 ( .A1(n353), .A2(n635), .Y(n583) );
  MUX41X1_HVT U56 ( .A1(n408), .A3(n298), .A2(n393), .A4(n583), .S0(n336), 
        .S1(n366), .Y(n582) );
  MUX41X1_HVT U62 ( .A1(n576), .A3(n582), .A2(n580), .A4(n584), .S0(n350), 
        .S1(n347), .Y(n575) );
  MUX41X1_HVT U65 ( .A1(n386), .A3(n388), .A2(n387), .A4(n599), .S0(n336), 
        .S1(n297), .Y(n572) );
  NAND2X0_HVT U66 ( .A1(n271), .A2(n310), .Y(n571) );
  MUX41X1_HVT U67 ( .A1(n383), .A3(n409), .A2(n385), .A4(n571), .S0(n297), 
        .S1(n333), .Y(n570) );
  MUX41X1_HVT U68 ( .A1(n383), .A3(n291), .A2(n384), .A4(n355), .S0(n335), 
        .S1(n366), .Y(n569) );
  NAND2X0_HVT U72 ( .A1(n298), .A2(n631), .Y(n566) );
  MUX41X1_HVT U73 ( .A1(n610), .A3(n566), .A2(n410), .A4(n341), .S0(n340), 
        .S1(n332), .Y(n565) );
  MUX41X1_HVT U74 ( .A1(n628), .A3(n400), .A2(n399), .A4(n276), .S0(n336), 
        .S1(n266), .Y(n564) );
  MUX41X1_HVT U78 ( .A1(n561), .A3(n565), .A2(n564), .A4(n567), .S0(n350), 
        .S1(n347), .Y(n560) );
  MUX41X1_HVT U79 ( .A1(n396), .A3(n619), .A2(n398), .A4(n620), .S0(n336), 
        .S1(n363), .Y(n559) );
  NAND2X0_HVT U81 ( .A1(n314), .A2(n631), .Y(n557) );
  AND2X1_HVT U82 ( .A1(n632), .A2(n352), .Y(n556) );
  MUX41X1_HVT U83 ( .A1(n556), .A3(n397), .A2(n413), .A4(n557), .S0(n335), 
        .S1(n366), .Y(n555) );
  MUX41X1_HVT U84 ( .A1(n320), .A3(n396), .A2(n414), .A4(n612), .S0(n336), 
        .S1(n266), .Y(n554) );
  MUX41X1_HVT U85 ( .A1(n554), .A3(n558), .A2(n555), .A4(n559), .S0(n350), 
        .S1(n347), .Y(n553) );
  NAND2X0_HVT U89 ( .A1(n277), .A2(n308), .Y(n550) );
  MUX41X1_HVT U99 ( .A1(n605), .A3(n387), .A2(n589), .A4(n298), .S0(n266), 
        .S1(n333), .Y(n540) );
  NAND2X0_HVT U100 ( .A1(n294), .A2(n424), .Y(n539) );
  MUX41X1_HVT U101 ( .A1(n418), .A3(n625), .A2(n401), .A4(n539), .S0(n366), 
        .S1(n331), .Y(n538) );
  MUX41X1_HVT U102 ( .A1(n538), .A3(n541), .A2(n540), .A4(n543), .S0(n350), 
        .S1(n347), .Y(n537) );
  AND2X1_HVT U104 ( .A1(n631), .A2(n304), .Y(n536) );
  MUX41X1_HVT U105 ( .A1(n623), .A3(n419), .A2(n557), .A4(n536), .S0(n336), 
        .S1(n366), .Y(n535) );
  MUX41X1_HVT U107 ( .A1(n418), .A3(n352), .A2(n534), .A4(n376), .S0(n335), 
        .S1(n297), .Y(n533) );
  MUX41X1_HVT U108 ( .A1(n276), .A3(n300), .A2(n393), .A4(n314), .S0(n336), 
        .S1(n363), .Y(n532) );
  MUX41X1_HVT U109 ( .A1(n417), .A3(n370), .A2(n414), .A4(n197), .S0(n335), 
        .S1(n266), .Y(n531) );
  MUX41X1_HVT U110 ( .A1(n531), .A3(n533), .A2(n532), .A4(n535), .S0(n350), 
        .S1(n348), .Y(n530) );
  NAND2X0_HVT U114 ( .A1(n355), .A2(n631), .Y(n526) );
  MUX41X1_HVT U115 ( .A1(n526), .A3(n626), .A2(n403), .A4(n352), .S0(n365), 
        .S1(n333), .Y(n525) );
  MUX41X1_HVT U116 ( .A1(n402), .A3(n396), .A2(n370), .A4(n622), .S0(n334), 
        .S1(n363), .Y(n524) );
  NAND2X0_HVT U118 ( .A1(n294), .A2(n291), .Y(n522) );
  MUX41X1_HVT U119 ( .A1(n420), .A3(n523), .A2(n600), .A4(n522), .S0(n334), 
        .S1(n365), .Y(n521) );
  MUX41X1_HVT U120 ( .A1(n521), .A3(n525), .A2(n524), .A4(n527), .S0(in[5]), 
        .S1(in[1]), .Y(n520) );
  MUX41X1_HVT U122 ( .A1(n407), .A3(n316), .A2(n591), .A4(n411), .S0(n334), 
        .S1(n366), .Y(n519) );
  MUX41X1_HVT U124 ( .A1(n318), .A3(n518), .A2(n614), .A4(n390), .S0(n266), 
        .S1(n334), .Y(n517) );
  AOI21X1_HVT U127 ( .A1(n339), .A2(n513), .A3(n377), .Y(n514) );
  NAND2X0_HVT U129 ( .A1(n338), .A2(n354), .Y(n511) );
  MUX41X1_HVT U130 ( .A1(n511), .A3(n512), .A2(n515), .A4(n514), .S0(n365), 
        .S1(n347), .Y(n510) );
  AND2X1_HVT U131 ( .A1(n310), .A2(n277), .Y(n509) );
  MUX41X1_HVT U132 ( .A1(n374), .A3(n509), .A2(n422), .A4(n383), .S0(n340), 
        .S1(n332), .Y(n508) );
  MUX41X1_HVT U133 ( .A1(n423), .A3(n376), .A2(n583), .A4(n375), .S0(n266), 
        .S1(n331), .Y(n507) );
  MUX41X1_HVT U136 ( .A1(n588), .A3(n539), .A2(n505), .A4(n381), .S0(n338), 
        .S1(n297), .Y(n504) );
  MUX41X1_HVT U137 ( .A1(n305), .A3(n608), .A2(n612), .A4(n416), .S0(n297), 
        .S1(n331), .Y(n503) );
  MUX41X1_HVT U139 ( .A1(n502), .A3(n506), .A2(n510), .A4(n516), .S0(in[5]), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n399), .A3(n317), .A2(n392), .A4(n626), .S0(n340), 
        .S1(n333), .Y(n501) );
  NAND2X0_HVT U141 ( .A1(n298), .A2(n277), .Y(n500) );
  MUX41X1_HVT U142 ( .A1(n500), .A3(n598), .A2(n421), .A4(n392), .S0(n339), 
        .S1(n365), .Y(n499) );
  MUX41X1_HVT U143 ( .A1(n425), .A3(n404), .A2(n617), .A4(n614), .S0(n337), 
        .S1(n297), .Y(n498) );
  MUX41X1_HVT U145 ( .A1(n606), .A3(n419), .A2(n497), .A4(n557), .S0(n339), 
        .S1(n363), .Y(n496) );
  MUX41X1_HVT U146 ( .A1(n496), .A3(n498), .A2(n499), .A4(n501), .S0(n348), 
        .S1(n350), .Y(n495) );
  MUX41X1_HVT U151 ( .A1(n413), .A3(n272), .A2(n324), .A4(n491), .S0(n365), 
        .S1(n331), .Y(n490) );
  MUX41X1_HVT U155 ( .A1(n392), .A3(n626), .A2(n618), .A4(n394), .S0(n337), 
        .S1(n363), .Y(n486) );
  NAND2X0_HVT U159 ( .A1(n482), .A2(n481), .Y(n483) );
  MUX41X1_HVT U162 ( .A1(n405), .A3(n388), .A2(n602), .A4(n479), .S0(n337), 
        .S1(n365), .Y(n478) );
  NAND2X0_HVT U163 ( .A1(n358), .A2(n425), .Y(n477) );
  NAND2X0_HVT U166 ( .A1(n627), .A2(n473), .Y(n474) );
  NAND2X0_HVT U177 ( .A1(n270), .A2(n291), .Y(n463) );
  AND2X1_HVT U179 ( .A1(n632), .A2(n304), .Y(n461) );
  AND2X1_HVT U185 ( .A1(n322), .A2(n294), .Y(n455) );
  MUX41X1_HVT U190 ( .A1(n452), .A3(n453), .A2(n451), .A4(n454), .S0(n348), 
        .S1(n332), .Y(n450) );
  NAND2X0_HVT U191 ( .A1(n303), .A2(n382), .Y(n449) );
  AND2X1_HVT U192 ( .A1(n400), .A2(n447), .Y(n448) );
  NAND2X0_HVT U194 ( .A1(n595), .A2(n447), .Y(n445) );
  MUX41X1_HVT U195 ( .A1(n446), .A3(n445), .A2(n448), .A4(n449), .S0(n335), 
        .S1(n348), .Y(n444) );
  NAND2X0_HVT U198 ( .A1(n271), .A2(n322), .Y(n627) );
  NAND2X0_HVT U200 ( .A1(n299), .A2(n277), .Y(n513) );
  NAND2X0_HVT U207 ( .A1(n277), .A2(n330), .Y(n577) );
  MUX21X2_HVT U2 ( .A1(n530), .A2(n520), .S0(n196), .Y(out[3]) );
  IBUFFX16_HVT U3 ( .A(in[7]), .Y(n196) );
  INVX0_HVT U4 ( .A(n611), .Y(n393) );
  XNOR2X1_HVT U6 ( .A1(n323), .A2(n358), .Y(n197) );
  INVX8_HVT U14 ( .A(n197), .Y(n591) );
  MUX41X1_HVT U16 ( .A1(n572), .A3(n569), .A2(n573), .A4(n570), .S0(n349), 
        .S1(n198), .Y(n568) );
  IBUFFX16_HVT U17 ( .A(n346), .Y(n198) );
  NAND2X0_HVT U18 ( .A1(n568), .A2(n199), .Y(n200) );
  NAND2X0_HVT U20 ( .A1(n575), .A2(n231), .Y(n201) );
  NAND2X0_HVT U21 ( .A1(n200), .A2(n201), .Y(out[0]) );
  INVX0_HVT U22 ( .A(n231), .Y(n199) );
  INVX1_HVT U23 ( .A(n249), .Y(n231) );
  NAND2X0_HVT U24 ( .A1(n563), .A2(n202), .Y(n218) );
  NAND2X0_HVT U25 ( .A1(n562), .A2(n339), .Y(n219) );
  NAND2X0_HVT U26 ( .A1(n218), .A2(n219), .Y(n561) );
  IBUFFX2_HVT U27 ( .A(n339), .Y(n202) );
  OA21X2_HVT U28 ( .A1(n372), .A2(n303), .A3(n616), .Y(n562) );
  IBUFFX2_HVT U29 ( .A(n349), .Y(n224) );
  INVX0_HVT U30 ( .A(in[5]), .Y(n349) );
  NAND2X0_HVT U31 ( .A1(n546), .A2(n220), .Y(n221) );
  NAND2X0_HVT U33 ( .A1(n547), .A2(n228), .Y(n222) );
  NAND2X0_HVT U34 ( .A1(n221), .A2(n222), .Y(n545) );
  INVX0_HVT U36 ( .A(n228), .Y(n220) );
  MUX21X1_HVT U37 ( .A1(n353), .A2(n548), .S0(n294), .Y(n547) );
  INVX1_HVT U39 ( .A(n229), .Y(n228) );
  INVX1_HVT U40 ( .A(n366), .Y(n284) );
  MUX21X2_HVT U41 ( .A1(n585), .A2(n586), .S0(n223), .Y(n584) );
  IBUFFX16_HVT U43 ( .A(n338), .Y(n223) );
  AO21X2_HVT U44 ( .A1(n403), .A2(n340), .A3(n613), .Y(n528) );
  MUX41X1_HVT U45 ( .A1(n466), .A3(n465), .A2(n469), .A4(n467), .S0(n346), 
        .S1(n224), .Y(n464) );
  NAND2X0_HVT U46 ( .A1(n495), .A2(n225), .Y(n226) );
  NAND2X0_HVT U47 ( .A1(n485), .A2(n290), .Y(n227) );
  NAND2X0_HVT U48 ( .A1(n226), .A2(n227), .Y(out[5]) );
  IBUFFX2_HVT U49 ( .A(n290), .Y(n225) );
  IBUFFX2_HVT U50 ( .A(in[7]), .Y(n290) );
  MUX41X1_HVT U51 ( .A1(n545), .A3(n551), .A2(n549), .A4(n552), .S0(n350), 
        .S1(n347), .Y(n544) );
  IBUFFX16_HVT U52 ( .A(n338), .Y(n229) );
  INVX1_HVT U54 ( .A(n346), .Y(n347) );
  INVX1_HVT U57 ( .A(n349), .Y(n350) );
  MUX41X1_HVT U58 ( .A1(n315), .A3(n615), .A2(n550), .A4(n468), .S0(n230), 
        .S1(n327), .Y(n467) );
  IBUFFX16_HVT U59 ( .A(n280), .Y(n230) );
  MUX21X2_HVT U60 ( .A1(n300), .A2(n427), .S0(n360), .Y(n606) );
  INVX1_HVT U61 ( .A(n429), .Y(n423) );
  INVX1_HVT U63 ( .A(n354), .Y(n427) );
  MUX41X1_HVT U64 ( .A1(n459), .A3(n456), .A2(n450), .A4(n444), .S0(n232), 
        .S1(n290), .Y(out[7]) );
  IBUFFX16_HVT U69 ( .A(in[5]), .Y(n232) );
  INVX0_HVT U70 ( .A(n632), .Y(n375) );
  NAND2X2_HVT U71 ( .A1(n359), .A2(n355), .Y(n632) );
  INVX0_HVT U75 ( .A(n274), .Y(n359) );
  INVX2_HVT U76 ( .A(n274), .Y(n358) );
  MUX21X2_HVT U77 ( .A1(n528), .A2(n529), .S0(n339), .Y(n527) );
  MUX21X2_HVT U80 ( .A1(n394), .A2(n384), .S0(n364), .Y(n586) );
  NAND2X0_HVT U86 ( .A1(n345), .A2(n233), .Y(n234) );
  NAND2X0_HVT U87 ( .A1(n427), .A2(n245), .Y(n235) );
  NAND2X0_HVT U88 ( .A1(n234), .A2(n235), .Y(n468) );
  INVX0_HVT U90 ( .A(n245), .Y(n233) );
  IBUFFX2_HVT U91 ( .A(n271), .Y(n245) );
  INVX0_HVT U92 ( .A(n321), .Y(n246) );
  INVX0_HVT U93 ( .A(n321), .Y(n253) );
  NBUFFX4_HVT U94 ( .A(n364), .Y(n340) );
  NAND2X0_HVT U95 ( .A1(n493), .A2(n236), .Y(n237) );
  NAND2X0_HVT U96 ( .A1(n494), .A2(n281), .Y(n238) );
  NAND2X0_HVT U97 ( .A1(n237), .A2(n238), .Y(n492) );
  IBUFFX2_HVT U98 ( .A(n281), .Y(n236) );
  NAND2X0_HVT U103 ( .A1(n304), .A2(n239), .Y(n240) );
  NAND2X0_HVT U106 ( .A1(n313), .A2(n278), .Y(n241) );
  NAND2X0_HVT U111 ( .A1(n240), .A2(n241), .Y(n430) );
  INVX1_HVT U112 ( .A(n278), .Y(n239) );
  AO21X2_HVT U113 ( .A1(n363), .A2(n378), .A3(n302), .Y(n493) );
  MUX21X1_HVT U117 ( .A1(n422), .A2(n374), .S0(n363), .Y(n494) );
  INVX1_HVT U121 ( .A(n311), .Y(n313) );
  IBUFFX2_HVT U123 ( .A(n277), .Y(n278) );
  INVX0_HVT U125 ( .A(n430), .Y(n422) );
  INVX2_HVT U126 ( .A(n621), .Y(n428) );
  NBUFFX4_HVT U128 ( .A(n309), .Y(n343) );
  MUX41X1_HVT U134 ( .A1(n470), .A3(n318), .A2(n315), .A4(n319), .S0(n242), 
        .S1(n243), .Y(n469) );
  IBUFFX16_HVT U135 ( .A(n337), .Y(n242) );
  IBUFFX16_HVT U138 ( .A(n266), .Y(n243) );
  IBUFFX16_HVT U144 ( .A(n367), .Y(n365) );
  MUX21X2_HVT U147 ( .A1(n537), .A2(n544), .S0(n244), .Y(out[2]) );
  IBUFFX16_HVT U148 ( .A(n290), .Y(n244) );
  NAND2X0_HVT U149 ( .A1(n391), .A2(n246), .Y(n247) );
  NAND2X0_HVT U150 ( .A1(n581), .A2(n321), .Y(n248) );
  NAND2X0_HVT U152 ( .A1(n247), .A2(n248), .Y(n580) );
  IBUFFX16_HVT U153 ( .A(in[7]), .Y(n249) );
  XNOR2X1_HVT U154 ( .A1(n303), .A2(n334), .Y(n321) );
  IBUFFX2_HVT U156 ( .A(n327), .Y(n251) );
  MUX41X1_HVT U157 ( .A1(n415), .A3(n583), .A2(n423), .A4(n428), .S0(n250), 
        .S1(n251), .Y(n465) );
  IBUFFX16_HVT U158 ( .A(n281), .Y(n250) );
  IBUFFX2_HVT U160 ( .A(n638), .Y(n330) );
  INVX1_HVT U161 ( .A(n262), .Y(n252) );
  INVX1_HVT U164 ( .A(n270), .Y(n262) );
  MUX21X1_HVT U165 ( .A1(n507), .A2(n508), .S0(n347), .Y(n506) );
  NAND2X0_HVT U167 ( .A1(n276), .A2(n253), .Y(n254) );
  NAND2X0_HVT U168 ( .A1(n574), .A2(n321), .Y(n255) );
  NAND2X0_HVT U169 ( .A1(n254), .A2(n255), .Y(n573) );
  INVX0_HVT U170 ( .A(n616), .Y(n276) );
  MUX21X1_HVT U171 ( .A1(n635), .A2(n324), .S0(n280), .Y(n574) );
  INVX1_HVT U172 ( .A(n272), .Y(n600) );
  INVX1_HVT U173 ( .A(in[6]), .Y(n309) );
  XNOR2X2_HVT U174 ( .A1(n343), .A2(n426), .Y(n621) );
  INVX0_HVT U175 ( .A(n322), .Y(n323) );
  INVX1_HVT U176 ( .A(n436), .Y(n415) );
  MUX41X1_HVT U178 ( .A1(n492), .A3(n490), .A2(n487), .A4(n486), .S0(n346), 
        .S1(n349), .Y(n485) );
  INVX0_HVT U180 ( .A(n324), .Y(n615) );
  IBUFFX2_HVT U181 ( .A(n364), .Y(n327) );
  IBUFFX2_HVT U182 ( .A(n364), .Y(n279) );
  IBUFFX2_HVT U183 ( .A(n367), .Y(n266) );
  IBUFFX2_HVT U184 ( .A(n367), .Y(n297) );
  IBUFFX16_HVT U186 ( .A(n364), .Y(n303) );
  MUX21X1_HVT U187 ( .A1(n425), .A2(n427), .S0(n358), .Y(n593) );
  IBUFFX2_HVT U188 ( .A(n359), .Y(n294) );
  MUX41X1_HVT U189 ( .A1(n592), .A3(n368), .A2(n461), .A4(n605), .S0(n284), 
        .S1(n287), .Y(n460) );
  NAND2X0_HVT U193 ( .A1(n462), .A2(n256), .Y(n257) );
  NAND2X0_HVT U196 ( .A1(n460), .A2(n263), .Y(n258) );
  NAND2X0_HVT U197 ( .A1(n257), .A2(n258), .Y(n459) );
  INVX0_HVT U199 ( .A(n263), .Y(n256) );
  IBUFFX2_HVT U201 ( .A(n626), .Y(n368) );
  INVX1_HVT U202 ( .A(n265), .Y(n263) );
  INVX0_HVT U203 ( .A(n593), .Y(n405) );
  NAND2X0_HVT U204 ( .A1(n457), .A2(n259), .Y(n260) );
  NAND2X0_HVT U205 ( .A1(n458), .A2(n348), .Y(n261) );
  NAND2X0_HVT U206 ( .A1(n261), .A2(n260), .Y(n456) );
  IBUFFX2_HVT U208 ( .A(n348), .Y(n259) );
  INVX2_HVT U209 ( .A(n346), .Y(n348) );
  MUX21X2_HVT U210 ( .A1(n301), .A2(n427), .S0(n262), .Y(n470) );
  INVX2_HVT U211 ( .A(n426), .Y(n291) );
  MUX21X1_HVT U212 ( .A1(n312), .A2(n323), .S0(n274), .Y(n324) );
  INVX1_HVT U213 ( .A(in[0]), .Y(n274) );
  INVX0_HVT U214 ( .A(n595), .Y(n376) );
  OR2X1_HVT U215 ( .A1(n309), .A2(n264), .Y(n633) );
  IBUFFX16_HVT U216 ( .A(n342), .Y(n264) );
  IBUFFX2_HVT U217 ( .A(n309), .Y(n310) );
  IBUFFX2_HVT U218 ( .A(n633), .Y(n308) );
  IBUFFX16_HVT U219 ( .A(n346), .Y(n265) );
  INVX1_HVT U220 ( .A(n351), .Y(n425) );
  INVX0_HVT U221 ( .A(n351), .Y(n275) );
  INVX1_HVT U222 ( .A(n273), .Y(n267) );
  INVX0_HVT U223 ( .A(n356), .Y(n273) );
  MUX21X1_HVT U224 ( .A1(n269), .A2(n637), .S0(n274), .Y(n268) );
  IBUFFX16_HVT U225 ( .A(n268), .Y(n614) );
  IBUFFX16_HVT U226 ( .A(n291), .Y(n269) );
  INVX1_HVT U227 ( .A(n637), .Y(n424) );
  INVX1_HVT U228 ( .A(n361), .Y(n270) );
  INVX1_HVT U229 ( .A(n361), .Y(n271) );
  XOR2X2_HVT U230 ( .A1(n354), .A2(n273), .Y(n272) );
  INVX0_HVT U231 ( .A(in[0]), .Y(n361) );
  INVX1_HVT U232 ( .A(n361), .Y(n357) );
  INVX1_HVT U233 ( .A(n361), .Y(n360) );
  INVX1_HVT U234 ( .A(n361), .Y(n356) );
  XNOR2X1_HVT U235 ( .A1(n275), .A2(n271), .Y(n589) );
  OA21X1_HVT U236 ( .A1(n396), .A2(n279), .A3(n577), .Y(n451) );
  MUX21X1_HVT U237 ( .A1(n323), .A2(n345), .S0(n340), .Y(n548) );
  OA21X1_HVT U238 ( .A1(n371), .A2(n279), .A3(n380), .Y(n488) );
  NAND2X0_HVT U239 ( .A1(n298), .A2(n340), .Y(n285) );
  INVX1_HVT U240 ( .A(n336), .Y(n287) );
  INVX1_HVT U241 ( .A(n332), .Y(n280) );
  INVX0_HVT U242 ( .A(n428), .Y(n300) );
  INVX0_HVT U243 ( .A(n428), .Y(n298) );
  INVX1_HVT U244 ( .A(in[1]), .Y(n346) );
  INVX1_HVT U245 ( .A(n338), .Y(n281) );
  INVX1_HVT U246 ( .A(n359), .Y(n277) );
  IBUFFX2_HVT U247 ( .A(n635), .Y(n373) );
  MUX41X1_HVT U248 ( .A1(n595), .A3(n389), .A2(n408), .A4(n404), .S0(n279), 
        .S1(n280), .Y(n457) );
  NAND2X0_HVT U249 ( .A1(n320), .A2(n279), .Y(n282) );
  NAND2X0_HVT U250 ( .A1(n589), .A2(n365), .Y(n283) );
  NAND2X0_HVT U251 ( .A1(n282), .A2(n283), .Y(n453) );
  MUX41X1_HVT U252 ( .A1(n330), .A3(n631), .A2(n590), .A4(n550), .S0(n331), 
        .S1(n266), .Y(n549) );
  INVX1_HVT U253 ( .A(n367), .Y(n364) );
  IBUFFX2_HVT U254 ( .A(n367), .Y(n366) );
  IBUFFX2_HVT U255 ( .A(n592), .Y(n406) );
  MUX41X1_HVT U256 ( .A1(n373), .A3(n413), .A2(n376), .A4(n635), .S0(n337), 
        .S1(n303), .Y(n458) );
  AO21X1_HVT U257 ( .A1(n298), .A2(n635), .A3(n279), .Y(n473) );
  NAND2X0_HVT U258 ( .A1(n379), .A2(n327), .Y(n286) );
  NAND2X0_HVT U259 ( .A1(n285), .A2(n286), .Y(n546) );
  MUX21X1_HVT U260 ( .A1(n455), .A2(n412), .S0(n363), .Y(n454) );
  MUX41X1_HVT U261 ( .A1(n417), .A3(n542), .A2(n609), .A4(n272), .S0(n287), 
        .S1(n365), .Y(n541) );
  NAND2X0_HVT U262 ( .A1(n483), .A2(n281), .Y(n288) );
  NAND2X0_HVT U263 ( .A1(n484), .A2(n339), .Y(n289) );
  NAND2X0_HVT U264 ( .A1(n288), .A2(n289), .Y(n480) );
  MUX21X1_HVT U265 ( .A1(n411), .A2(n594), .S0(n327), .Y(n484) );
  INVX0_HVT U266 ( .A(n594), .Y(n404) );
  INVX1_HVT U267 ( .A(in[4]), .Y(n367) );
  AO21X2_HVT U268 ( .A1(n277), .A2(n354), .A3(n279), .Y(n481) );
  MUX41X1_HVT U269 ( .A1(n379), .A3(n626), .A2(n330), .A4(n632), .S0(n287), 
        .S1(n279), .Y(n567) );
  MUX21X2_HVT U270 ( .A1(n560), .A2(n553), .S0(n290), .Y(out[1]) );
  AO21X2_HVT U271 ( .A1(n358), .A2(n424), .A3(n279), .Y(n447) );
  MUX21X1_HVT U272 ( .A1(n341), .A2(n301), .S0(n270), .Y(n594) );
  MUX21X1_HVT U273 ( .A1(n351), .A2(n353), .S0(n360), .Y(n479) );
  MUX21X1_HVT U274 ( .A1(n330), .A2(n308), .S0(n360), .Y(n609) );
  MUX21X1_HVT U275 ( .A1(n345), .A2(n621), .S0(n274), .Y(n612) );
  INVX1_HVT U276 ( .A(in[3]), .Y(n426) );
  INVX1_HVT U277 ( .A(n292), .Y(n542) );
  NBUFFX2_HVT U278 ( .A(n426), .Y(n342) );
  IBUFFX2_HVT U279 ( .A(n304), .Y(n293) );
  MUX21X1_HVT U280 ( .A1(n341), .A2(n293), .S0(n294), .Y(n292) );
  NAND2X0_HVT U281 ( .A1(n390), .A2(n303), .Y(n295) );
  NAND2X0_HVT U282 ( .A1(n583), .A2(n340), .Y(n296) );
  NAND2X0_HVT U283 ( .A1(n295), .A2(n296), .Y(n579) );
  MUX21X1_HVT U284 ( .A1(n579), .A2(n578), .S0(n338), .Y(n576) );
  IBUFFX2_HVT U285 ( .A(n624), .Y(n380) );
  MUX41X1_HVT U286 ( .A1(n624), .A3(n409), .A2(n416), .A4(n394), .S0(n281), 
        .S1(n297), .Y(n543) );
  MUX41X1_HVT U287 ( .A1(n415), .A3(n393), .A2(n373), .A4(n320), .S0(n334), 
        .S1(n327), .Y(n552) );
  MUX21X1_HVT U288 ( .A1(n323), .A2(n341), .S0(n356), .Y(n616) );
  INVX0_HVT U289 ( .A(n308), .Y(n299) );
  IBUFFX2_HVT U290 ( .A(n609), .Y(n395) );
  MUX21X1_HVT U291 ( .A1(n344), .A2(n302), .S0(n277), .Y(n441) );
  IBUFFX2_HVT U292 ( .A(n629), .Y(n381) );
  MUX41X1_HVT U293 ( .A1(n478), .A3(n480), .A2(n472), .A4(n476), .S0(n348), 
        .S1(n349), .Y(n471) );
  INVX1_HVT U294 ( .A(n636), .Y(n301) );
  INVX1_HVT U295 ( .A(n440), .Y(n411) );
  OR2X1_HVT U296 ( .A1(n426), .A2(n309), .Y(n636) );
  IBUFFX2_HVT U297 ( .A(n367), .Y(n363) );
  INVX0_HVT U298 ( .A(n312), .Y(n302) );
  INVX1_HVT U299 ( .A(n608), .Y(n396) );
  AO21X1_HVT U300 ( .A1(n577), .A2(n366), .A3(n616), .Y(n578) );
  MUX41X1_HVT U301 ( .A1(n591), .A3(n607), .A2(n370), .A4(n385), .S0(n281), 
        .S1(n303), .Y(n551) );
  MUX21X2_HVT U302 ( .A1(n474), .A2(n475), .S0(n338), .Y(n472) );
  MUX41X1_HVT U303 ( .A1(n389), .A3(n600), .A2(n477), .A4(n629), .S0(n281), 
        .S1(n303), .Y(n476) );
  INVX1_HVT U304 ( .A(n441), .Y(n410) );
  INVX1_HVT U305 ( .A(n311), .Y(n312) );
  NBUFFX2_HVT U306 ( .A(n633), .Y(n304) );
  INVX1_HVT U307 ( .A(n616), .Y(n389) );
  NAND2X0_HVT U308 ( .A1(n359), .A2(n637), .Y(n635) );
  INVX1_HVT U309 ( .A(n378), .Y(n305) );
  INVX1_HVT U310 ( .A(n637), .Y(n311) );
  NAND2X0_HVT U311 ( .A1(n464), .A2(n290), .Y(n306) );
  NAND2X0_HVT U312 ( .A1(n471), .A2(in[7]), .Y(n307) );
  NAND2X0_HVT U313 ( .A1(n307), .A2(n306), .Y(out[6]) );
  MUX41X1_HVT U314 ( .A1(n634), .A3(n629), .A2(n408), .A4(n412), .S0(n281), 
        .S1(n284), .Y(n558) );
  INVX1_HVT U315 ( .A(n443), .Y(n408) );
  MUX21X1_HVT U316 ( .A1(n517), .A2(n519), .S0(n348), .Y(n516) );
  INVX0_HVT U317 ( .A(n311), .Y(n314) );
  MUX21X2_HVT U318 ( .A1(n410), .A2(n596), .S0(n340), .Y(n452) );
  MUX21X2_HVT U319 ( .A1(n503), .A2(n504), .S0(n348), .Y(n502) );
  AND2X1_HVT U320 ( .A1(n632), .A2(n312), .Y(n315) );
  AND2X1_HVT U321 ( .A1(n313), .A2(n622), .Y(n316) );
  MUX21X1_HVT U322 ( .A1(n406), .A2(n318), .S0(n297), .Y(n446) );
  NAND2X0_HVT U323 ( .A1(n342), .A2(n343), .Y(n637) );
  MUX21X1_HVT U324 ( .A1(n342), .A2(n424), .S0(n357), .Y(n607) );
  MUX21X1_HVT U325 ( .A1(n301), .A2(n341), .S0(n356), .Y(n440) );
  MUX21X1_HVT U326 ( .A1(n427), .A2(n298), .S0(n270), .Y(n436) );
  MUX21X1_HVT U327 ( .A1(n353), .A2(n314), .S0(n359), .Y(n619) );
  MUX21X1_HVT U328 ( .A1(n604), .A2(n316), .S0(n339), .Y(n512) );
  MUX21X1_HVT U329 ( .A1(n424), .A2(n301), .S0(n360), .Y(n587) );
  MUX21X1_HVT U330 ( .A1(n421), .A2(n317), .S0(n338), .Y(n515) );
  MUX21X1_HVT U331 ( .A1(n300), .A2(n308), .S0(n267), .Y(n603) );
  XOR2X1_HVT U332 ( .A1(n352), .A2(n271), .Y(n590) );
  MUX21X1_HVT U333 ( .A1(n341), .A2(n314), .S0(n359), .Y(n439) );
  MUX21X1_HVT U334 ( .A1(n343), .A2(n300), .S0(n270), .Y(n597) );
  MUX21X1_HVT U335 ( .A1(n343), .A2(n312), .S0(n356), .Y(n534) );
  XNOR2X1_HVT U336 ( .A1(n313), .A2(n270), .Y(n317) );
  MUX21X1_HVT U337 ( .A1(n353), .A2(n342), .S0(n356), .Y(n618) );
  MUX21X1_HVT U338 ( .A1(n353), .A2(n344), .S0(n358), .Y(n518) );
  MUX21X1_HVT U339 ( .A1(n341), .A2(n636), .S0(n357), .Y(n433) );
  AND2X1_HVT U340 ( .A1(n267), .A2(n345), .Y(n318) );
  INVX0_HVT U341 ( .A(n614), .Y(n390) );
  MUX21X1_HVT U342 ( .A1(n411), .A2(n369), .S0(n365), .Y(n563) );
  NBUFFX2_HVT U343 ( .A(n636), .Y(n352) );
  AND2X1_HVT U344 ( .A1(n301), .A2(n294), .Y(n319) );
  MUX21X1_HVT U345 ( .A1(n392), .A2(n634), .S0(n339), .Y(n581) );
  NBUFFX2_HVT U346 ( .A(n633), .Y(n351) );
  AND2X1_HVT U347 ( .A1(n353), .A2(n294), .Y(n320) );
  NBUFFX2_HVT U348 ( .A(n636), .Y(n353) );
  MUX21X1_HVT U349 ( .A1(n377), .A2(n596), .S0(n366), .Y(n529) );
  NBUFFX2_HVT U350 ( .A(n309), .Y(n345) );
  NBUFFX2_HVT U351 ( .A(n426), .Y(n341) );
  NBUFFX2_HVT U352 ( .A(n362), .Y(n338) );
  NBUFFX2_HVT U353 ( .A(n362), .Y(n334) );
  NBUFFX2_HVT U354 ( .A(n362), .Y(n335) );
  NBUFFX2_HVT U355 ( .A(n362), .Y(n336) );
  NBUFFX2_HVT U356 ( .A(n362), .Y(n339) );
  NBUFFX2_HVT U357 ( .A(n362), .Y(n337) );
  NBUFFX2_HVT U358 ( .A(n362), .Y(n332) );
  NBUFFX2_HVT U359 ( .A(n335), .Y(n333) );
  NBUFFX2_HVT U360 ( .A(n337), .Y(n331) );
  MUX21X1_HVT U361 ( .A1(n427), .A2(n291), .S0(n358), .Y(n429) );
  MUX21X1_HVT U362 ( .A1(n355), .A2(n291), .S0(n360), .Y(n482) );
  MUX21X1_HVT U363 ( .A1(n291), .A2(n355), .S0(n357), .Y(n435) );
  MUX21X1_HVT U364 ( .A1(n345), .A2(n291), .S0(n357), .Y(n610) );
  MUX21X1_HVT U365 ( .A1(n301), .A2(n425), .S0(n271), .Y(n523) );
  MUX21X1_HVT U366 ( .A1(n291), .A2(n304), .S0(n252), .Y(n434) );
  NBUFFX2_HVT U367 ( .A(in[2]), .Y(n362) );
  INVX1_HVT U368 ( .A(n621), .Y(n322) );
  INVX1_HVT U369 ( .A(n438), .Y(n413) );
  MUX21X1_HVT U370 ( .A1(n312), .A2(n299), .S0(n356), .Y(n497) );
  NAND2X0_HVT U371 ( .A1(n489), .A2(n335), .Y(n325) );
  NAND2X0_HVT U372 ( .A1(n488), .A2(n287), .Y(n326) );
  NAND2X0_HVT U373 ( .A1(n325), .A2(n326), .Y(n487) );
  MUX21X1_HVT U374 ( .A1(n612), .A2(n320), .S0(n340), .Y(n489) );
  MUX41X1_HVT U375 ( .A1(n601), .A3(n314), .A2(n330), .A4(n355), .S0(n281), 
        .S1(n303), .Y(n466) );
  MUX21X1_HVT U376 ( .A1(n343), .A2(n308), .S0(n360), .Y(n491) );
  NAND2X0_HVT U377 ( .A1(n327), .A2(n611), .Y(n328) );
  NAND2X0_HVT U378 ( .A1(n614), .A2(n340), .Y(n329) );
  NAND2X0_HVT U379 ( .A1(n328), .A2(n329), .Y(n475) );
  MUX21X1_HVT U380 ( .A1(n322), .A2(n345), .S0(n358), .Y(n431) );
  MUX21X1_HVT U381 ( .A1(n424), .A2(n428), .S0(n267), .Y(n604) );
  MUX21X1_HVT U382 ( .A1(n428), .A2(n342), .S0(n271), .Y(n598) );
  MUX21X1_HVT U383 ( .A1(n354), .A2(n313), .S0(n358), .Y(n623) );
  MUX21X1_HVT U384 ( .A1(n343), .A2(n322), .S0(n358), .Y(n601) );
  MUX21X1_HVT U385 ( .A1(n424), .A2(n310), .S0(n357), .Y(n505) );
  XOR2X1_HVT U386 ( .A1(n267), .A2(n310), .Y(n588) );
  MUX21X1_HVT U387 ( .A1(n310), .A2(n330), .S0(n252), .Y(n613) );
  MUX21X1_HVT U388 ( .A1(n636), .A2(n310), .S0(n356), .Y(n437) );
  MUX21X1_HVT U389 ( .A1(n310), .A2(n353), .S0(n356), .Y(n442) );
  MUX21X1_HVT U390 ( .A1(n310), .A2(n354), .S0(n357), .Y(n620) );
  MUX21X1_HVT U391 ( .A1(n341), .A2(n310), .S0(n360), .Y(n432) );
  MUX21X1_HVT U392 ( .A1(n304), .A2(n310), .S0(n357), .Y(n608) );
  MUX41X1_HVT U393 ( .A1(n593), .A3(n330), .A2(n463), .A4(n319), .S0(n287), 
        .S1(n303), .Y(n462) );
  NBUFFX2_HVT U394 ( .A(n309), .Y(n344) );
  MUX21X1_HVT U395 ( .A1(n342), .A2(n344), .S0(n359), .Y(n592) );
  MUX21X1_HVT U396 ( .A1(n344), .A2(n424), .S0(n358), .Y(n611) );
  MUX21X1_HVT U397 ( .A1(n310), .A2(n301), .S0(n360), .Y(n596) );
  MUX21X1_HVT U398 ( .A1(n310), .A2(n308), .S0(n357), .Y(n443) );
  MUX21X1_HVT U399 ( .A1(n341), .A2(n428), .S0(n358), .Y(n438) );
  NBUFFX2_HVT U400 ( .A(n638), .Y(n354) );
  NBUFFX2_HVT U401 ( .A(n638), .Y(n355) );
  INVX0_HVT U402 ( .A(n605), .Y(n369) );
  INVX0_HVT U403 ( .A(n599), .Y(n370) );
  INVX0_HVT U404 ( .A(n539), .Y(n371) );
  INVX0_HVT U405 ( .A(n500), .Y(n372) );
  INVX0_HVT U406 ( .A(n634), .Y(n374) );
  INVX0_HVT U407 ( .A(n631), .Y(n377) );
  INVX0_HVT U408 ( .A(n630), .Y(n378) );
  INVX0_HVT U409 ( .A(n602), .Y(n379) );
  INVX0_HVT U410 ( .A(n625), .Y(n382) );
  INVX0_HVT U411 ( .A(n623), .Y(n383) );
  INVX0_HVT U412 ( .A(n622), .Y(n384) );
  INVX0_HVT U413 ( .A(n620), .Y(n385) );
  INVX0_HVT U414 ( .A(n619), .Y(n386) );
  INVX0_HVT U415 ( .A(n618), .Y(n387) );
  INVX0_HVT U416 ( .A(n617), .Y(n388) );
  INVX0_HVT U417 ( .A(n613), .Y(n391) );
  INVX0_HVT U418 ( .A(n612), .Y(n392) );
  INVX0_HVT U419 ( .A(n610), .Y(n394) );
  INVX0_HVT U420 ( .A(n607), .Y(n397) );
  INVX0_HVT U421 ( .A(n606), .Y(n398) );
  INVX0_HVT U422 ( .A(n604), .Y(n399) );
  INVX0_HVT U423 ( .A(n603), .Y(n400) );
  INVX0_HVT U424 ( .A(n601), .Y(n401) );
  INVX0_HVT U425 ( .A(n598), .Y(n402) );
  INVX0_HVT U426 ( .A(n597), .Y(n403) );
  INVX0_HVT U427 ( .A(n628), .Y(n407) );
  INVX0_HVT U428 ( .A(n442), .Y(n409) );
  INVX0_HVT U429 ( .A(n439), .Y(n412) );
  INVX0_HVT U430 ( .A(n437), .Y(n414) );
  INVX0_HVT U431 ( .A(n435), .Y(n416) );
  INVX0_HVT U432 ( .A(n434), .Y(n417) );
  INVX0_HVT U433 ( .A(n433), .Y(n418) );
  INVX0_HVT U434 ( .A(n432), .Y(n419) );
  INVX0_HVT U435 ( .A(n482), .Y(n420) );
  INVX0_HVT U436 ( .A(n431), .Y(n421) );
endmodule

