
module round ( in, round_num, keyin, keyout, out );
  input [127:0] in;
  input [3:0] round_num;
  input [127:0] keyin;
  output [127:0] keyout;
  output [127:0] out;
  wire   \_0_net_[127] , \_0_net_[126] , \_0_net_[125] , \_0_net_[124] ,
         \_0_net_[123] , \_0_net_[122] , \_0_net_[121] , \_0_net_[120] ,
         \_0_net_[119] , \_0_net_[118] , \_0_net_[117] , \_0_net_[116] ,
         \_0_net_[115] , \_0_net_[114] , \_0_net_[113] , \_0_net_[112] ,
         \_0_net_[111] , \_0_net_[110] , \_0_net_[109] , \_0_net_[108] ,
         \_0_net_[107] , \_0_net_[106] , \_0_net_[105] , \_0_net_[104] ,
         \_0_net_[103] , \_0_net_[102] , \_0_net_[101] , \_0_net_[100] ,
         \_0_net_[99] , \_0_net_[98] , \_0_net_[97] , \_0_net_[96] ,
         \_0_net_[95] , \_0_net_[94] , \_0_net_[93] , \_0_net_[92] ,
         \_0_net_[91] , \_0_net_[90] , \_0_net_[89] , \_0_net_[88] ,
         \_0_net_[87] , \_0_net_[86] , \_0_net_[85] , \_0_net_[84] ,
         \_0_net_[83] , \_0_net_[82] , \_0_net_[81] , \_0_net_[80] ,
         \_0_net_[79] , \_0_net_[78] , \_0_net_[77] , \_0_net_[76] ,
         \_0_net_[75] , \_0_net_[74] , \_0_net_[73] , \_0_net_[72] ,
         \_0_net_[71] , \_0_net_[70] , \_0_net_[69] , \_0_net_[68] ,
         \_0_net_[67] , \_0_net_[66] , \_0_net_[65] , \_0_net_[64] ,
         \_0_net_[63] , \_0_net_[62] , \_0_net_[61] , \_0_net_[60] ,
         \_0_net_[59] , \_0_net_[58] , \_0_net_[57] , \_0_net_[56] ,
         \_0_net_[55] , \_0_net_[54] , \_0_net_[53] , \_0_net_[52] ,
         \_0_net_[51] , \_0_net_[50] , \_0_net_[49] , \_0_net_[48] ,
         \_0_net_[47] , \_0_net_[46] , \_0_net_[45] , \_0_net_[44] ,
         \_0_net_[43] , \_0_net_[42] , \_0_net_[41] , \_0_net_[40] ,
         \_0_net_[39] , \_0_net_[38] , \_0_net_[37] , \_0_net_[36] ,
         \_0_net_[35] , \_0_net_[34] , \_0_net_[33] , \_0_net_[32] ,
         \_0_net_[31] , \_0_net_[30] , \_0_net_[29] , \_0_net_[28] ,
         \_0_net_[27] , \_0_net_[26] , \_0_net_[25] , \_0_net_[24] ,
         \_0_net_[23] , \_0_net_[22] , \_0_net_[21] , \_0_net_[20] ,
         \_0_net_[19] , \_0_net_[18] , \_0_net_[17] , \_0_net_[16] ,
         \_0_net_[15] , \_0_net_[14] , \_0_net_[13] , \_0_net_[12] ,
         \_0_net_[11] , \_0_net_[10] , \_0_net_[9] , \_0_net_[8] ,
         \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] , \_0_net_[3] ,
         \_0_net_[2] , \_0_net_[1] , \_0_net_[0] , n1, n2;
  wire   [127:0] sb_out;
  wire   [127:0] sr_out;
  wire   [127:0] mc_out;

  keygen_0 x ( .round_num(round_num), .keyin(keyin), .keyout(keyout) );
  subbytes sb ( .in(in), .out(sb_out) );
  shift_rows sr ( .in(sb_out), .out(sr_out) );
  Mix_Column mc ( .in(sr_out), .out(mc_out) );
  add_round_keys_1 adk ( .state({\_0_net_[127] , \_0_net_[126] , 
        \_0_net_[125] , \_0_net_[124] , \_0_net_[123] , \_0_net_[122] , 
        \_0_net_[121] , \_0_net_[120] , \_0_net_[119] , \_0_net_[118] , 
        \_0_net_[117] , \_0_net_[116] , \_0_net_[115] , \_0_net_[114] , 
        \_0_net_[113] , \_0_net_[112] , \_0_net_[111] , \_0_net_[110] , 
        \_0_net_[109] , \_0_net_[108] , \_0_net_[107] , \_0_net_[106] , 
        \_0_net_[105] , \_0_net_[104] , \_0_net_[103] , \_0_net_[102] , 
        \_0_net_[101] , \_0_net_[100] , \_0_net_[99] , \_0_net_[98] , 
        \_0_net_[97] , \_0_net_[96] , \_0_net_[95] , \_0_net_[94] , 
        \_0_net_[93] , \_0_net_[92] , \_0_net_[91] , \_0_net_[90] , 
        \_0_net_[89] , \_0_net_[88] , \_0_net_[87] , \_0_net_[86] , 
        \_0_net_[85] , \_0_net_[84] , \_0_net_[83] , \_0_net_[82] , 
        \_0_net_[81] , \_0_net_[80] , \_0_net_[79] , \_0_net_[78] , 
        \_0_net_[77] , \_0_net_[76] , \_0_net_[75] , \_0_net_[74] , 
        \_0_net_[73] , \_0_net_[72] , \_0_net_[71] , \_0_net_[70] , 
        \_0_net_[69] , \_0_net_[68] , \_0_net_[67] , \_0_net_[66] , 
        \_0_net_[65] , \_0_net_[64] , \_0_net_[63] , \_0_net_[62] , 
        \_0_net_[61] , \_0_net_[60] , \_0_net_[59] , \_0_net_[58] , 
        \_0_net_[57] , \_0_net_[56] , \_0_net_[55] , \_0_net_[54] , 
        \_0_net_[53] , \_0_net_[52] , \_0_net_[51] , \_0_net_[50] , 
        \_0_net_[49] , \_0_net_[48] , \_0_net_[47] , \_0_net_[46] , 
        \_0_net_[45] , \_0_net_[44] , \_0_net_[43] , \_0_net_[42] , 
        \_0_net_[41] , \_0_net_[40] , \_0_net_[39] , \_0_net_[38] , 
        \_0_net_[37] , \_0_net_[36] , \_0_net_[35] , \_0_net_[34] , 
        \_0_net_[33] , \_0_net_[32] , \_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_0_net_[0] }), 
        .subkey(keyout), .out(out) );
  MUX21X1_HVT U1 ( .A1(mc_out[9]), .A2(sr_out[9]), .S0(n1), .Y(\_0_net_[9] )
         );
  MUX21X1_HVT U2 ( .A1(mc_out[99]), .A2(sr_out[99]), .S0(n1), .Y(\_0_net_[99] ) );
  MUX21X1_HVT U3 ( .A1(mc_out[98]), .A2(sr_out[98]), .S0(n1), .Y(\_0_net_[98] ) );
  MUX21X1_HVT U4 ( .A1(mc_out[97]), .A2(sr_out[97]), .S0(n1), .Y(\_0_net_[97] ) );
  MUX21X1_HVT U5 ( .A1(mc_out[96]), .A2(sr_out[96]), .S0(n1), .Y(\_0_net_[96] ) );
  MUX21X1_HVT U6 ( .A1(mc_out[95]), .A2(sr_out[95]), .S0(n1), .Y(\_0_net_[95] ) );
  MUX21X1_HVT U7 ( .A1(mc_out[94]), .A2(sr_out[94]), .S0(n1), .Y(\_0_net_[94] ) );
  MUX21X1_HVT U8 ( .A1(mc_out[93]), .A2(sr_out[93]), .S0(n1), .Y(\_0_net_[93] ) );
  MUX21X1_HVT U9 ( .A1(mc_out[92]), .A2(sr_out[92]), .S0(n1), .Y(\_0_net_[92] ) );
  MUX21X1_HVT U10 ( .A1(mc_out[91]), .A2(sr_out[91]), .S0(n1), .Y(
        \_0_net_[91] ) );
  MUX21X1_HVT U11 ( .A1(mc_out[90]), .A2(sr_out[90]), .S0(n1), .Y(
        \_0_net_[90] ) );
  MUX21X1_HVT U12 ( .A1(mc_out[8]), .A2(sr_out[8]), .S0(n1), .Y(\_0_net_[8] )
         );
  MUX21X1_HVT U13 ( .A1(mc_out[89]), .A2(sr_out[89]), .S0(n1), .Y(
        \_0_net_[89] ) );
  MUX21X1_HVT U14 ( .A1(mc_out[88]), .A2(sr_out[88]), .S0(n1), .Y(
        \_0_net_[88] ) );
  MUX21X1_HVT U15 ( .A1(mc_out[87]), .A2(sr_out[87]), .S0(n1), .Y(
        \_0_net_[87] ) );
  MUX21X1_HVT U16 ( .A1(mc_out[86]), .A2(sr_out[86]), .S0(n1), .Y(
        \_0_net_[86] ) );
  MUX21X1_HVT U17 ( .A1(mc_out[85]), .A2(sr_out[85]), .S0(n1), .Y(
        \_0_net_[85] ) );
  MUX21X1_HVT U18 ( .A1(mc_out[84]), .A2(sr_out[84]), .S0(n1), .Y(
        \_0_net_[84] ) );
  MUX21X1_HVT U19 ( .A1(mc_out[83]), .A2(sr_out[83]), .S0(n1), .Y(
        \_0_net_[83] ) );
  MUX21X1_HVT U20 ( .A1(mc_out[82]), .A2(sr_out[82]), .S0(n1), .Y(
        \_0_net_[82] ) );
  MUX21X1_HVT U21 ( .A1(mc_out[81]), .A2(sr_out[81]), .S0(n1), .Y(
        \_0_net_[81] ) );
  MUX21X1_HVT U22 ( .A1(mc_out[80]), .A2(sr_out[80]), .S0(n1), .Y(
        \_0_net_[80] ) );
  MUX21X1_HVT U23 ( .A1(mc_out[7]), .A2(sr_out[7]), .S0(n1), .Y(\_0_net_[7] )
         );
  MUX21X1_HVT U24 ( .A1(mc_out[79]), .A2(sr_out[79]), .S0(n1), .Y(
        \_0_net_[79] ) );
  MUX21X1_HVT U25 ( .A1(mc_out[78]), .A2(sr_out[78]), .S0(n1), .Y(
        \_0_net_[78] ) );
  MUX21X1_HVT U26 ( .A1(mc_out[77]), .A2(sr_out[77]), .S0(n1), .Y(
        \_0_net_[77] ) );
  MUX21X1_HVT U27 ( .A1(mc_out[76]), .A2(sr_out[76]), .S0(n1), .Y(
        \_0_net_[76] ) );
  MUX21X1_HVT U28 ( .A1(mc_out[75]), .A2(sr_out[75]), .S0(n1), .Y(
        \_0_net_[75] ) );
  MUX21X1_HVT U29 ( .A1(mc_out[74]), .A2(sr_out[74]), .S0(n1), .Y(
        \_0_net_[74] ) );
  MUX21X1_HVT U30 ( .A1(mc_out[73]), .A2(sr_out[73]), .S0(n1), .Y(
        \_0_net_[73] ) );
  MUX21X1_HVT U31 ( .A1(mc_out[72]), .A2(sr_out[72]), .S0(n1), .Y(
        \_0_net_[72] ) );
  MUX21X1_HVT U32 ( .A1(mc_out[71]), .A2(sr_out[71]), .S0(n1), .Y(
        \_0_net_[71] ) );
  MUX21X1_HVT U33 ( .A1(mc_out[70]), .A2(sr_out[70]), .S0(n1), .Y(
        \_0_net_[70] ) );
  MUX21X1_HVT U34 ( .A1(mc_out[6]), .A2(sr_out[6]), .S0(n1), .Y(\_0_net_[6] )
         );
  MUX21X1_HVT U35 ( .A1(mc_out[69]), .A2(sr_out[69]), .S0(n1), .Y(
        \_0_net_[69] ) );
  MUX21X1_HVT U36 ( .A1(mc_out[68]), .A2(sr_out[68]), .S0(n1), .Y(
        \_0_net_[68] ) );
  MUX21X1_HVT U37 ( .A1(mc_out[67]), .A2(sr_out[67]), .S0(n1), .Y(
        \_0_net_[67] ) );
  MUX21X1_HVT U38 ( .A1(mc_out[66]), .A2(sr_out[66]), .S0(n1), .Y(
        \_0_net_[66] ) );
  MUX21X1_HVT U39 ( .A1(mc_out[65]), .A2(sr_out[65]), .S0(n1), .Y(
        \_0_net_[65] ) );
  MUX21X1_HVT U40 ( .A1(mc_out[64]), .A2(sr_out[64]), .S0(n1), .Y(
        \_0_net_[64] ) );
  MUX21X1_HVT U41 ( .A1(mc_out[63]), .A2(sr_out[63]), .S0(n1), .Y(
        \_0_net_[63] ) );
  MUX21X1_HVT U42 ( .A1(mc_out[62]), .A2(sr_out[62]), .S0(n1), .Y(
        \_0_net_[62] ) );
  MUX21X1_HVT U43 ( .A1(mc_out[61]), .A2(sr_out[61]), .S0(n1), .Y(
        \_0_net_[61] ) );
  MUX21X1_HVT U44 ( .A1(mc_out[60]), .A2(sr_out[60]), .S0(n1), .Y(
        \_0_net_[60] ) );
  MUX21X1_HVT U45 ( .A1(mc_out[5]), .A2(sr_out[5]), .S0(n1), .Y(\_0_net_[5] )
         );
  MUX21X1_HVT U46 ( .A1(mc_out[59]), .A2(sr_out[59]), .S0(n1), .Y(
        \_0_net_[59] ) );
  MUX21X1_HVT U47 ( .A1(mc_out[58]), .A2(sr_out[58]), .S0(n1), .Y(
        \_0_net_[58] ) );
  MUX21X1_HVT U48 ( .A1(mc_out[57]), .A2(sr_out[57]), .S0(n1), .Y(
        \_0_net_[57] ) );
  MUX21X1_HVT U49 ( .A1(mc_out[56]), .A2(sr_out[56]), .S0(n1), .Y(
        \_0_net_[56] ) );
  MUX21X1_HVT U50 ( .A1(mc_out[55]), .A2(sr_out[55]), .S0(n1), .Y(
        \_0_net_[55] ) );
  MUX21X1_HVT U51 ( .A1(mc_out[54]), .A2(sr_out[54]), .S0(n1), .Y(
        \_0_net_[54] ) );
  MUX21X1_HVT U52 ( .A1(mc_out[53]), .A2(sr_out[53]), .S0(n1), .Y(
        \_0_net_[53] ) );
  MUX21X1_HVT U53 ( .A1(mc_out[52]), .A2(sr_out[52]), .S0(n1), .Y(
        \_0_net_[52] ) );
  MUX21X1_HVT U54 ( .A1(mc_out[51]), .A2(sr_out[51]), .S0(n1), .Y(
        \_0_net_[51] ) );
  MUX21X1_HVT U55 ( .A1(mc_out[50]), .A2(sr_out[50]), .S0(n1), .Y(
        \_0_net_[50] ) );
  MUX21X1_HVT U56 ( .A1(mc_out[4]), .A2(sr_out[4]), .S0(n1), .Y(\_0_net_[4] )
         );
  MUX21X1_HVT U57 ( .A1(mc_out[49]), .A2(sr_out[49]), .S0(n1), .Y(
        \_0_net_[49] ) );
  MUX21X1_HVT U58 ( .A1(mc_out[48]), .A2(sr_out[48]), .S0(n1), .Y(
        \_0_net_[48] ) );
  MUX21X1_HVT U59 ( .A1(mc_out[47]), .A2(sr_out[47]), .S0(n1), .Y(
        \_0_net_[47] ) );
  MUX21X1_HVT U60 ( .A1(mc_out[46]), .A2(sr_out[46]), .S0(n1), .Y(
        \_0_net_[46] ) );
  MUX21X1_HVT U61 ( .A1(mc_out[45]), .A2(sr_out[45]), .S0(n1), .Y(
        \_0_net_[45] ) );
  MUX21X1_HVT U62 ( .A1(mc_out[44]), .A2(sr_out[44]), .S0(n1), .Y(
        \_0_net_[44] ) );
  MUX21X1_HVT U63 ( .A1(mc_out[43]), .A2(sr_out[43]), .S0(n1), .Y(
        \_0_net_[43] ) );
  MUX21X1_HVT U64 ( .A1(mc_out[42]), .A2(sr_out[42]), .S0(n1), .Y(
        \_0_net_[42] ) );
  MUX21X1_HVT U65 ( .A1(mc_out[41]), .A2(sr_out[41]), .S0(n1), .Y(
        \_0_net_[41] ) );
  MUX21X1_HVT U66 ( .A1(mc_out[40]), .A2(sr_out[40]), .S0(n1), .Y(
        \_0_net_[40] ) );
  MUX21X1_HVT U67 ( .A1(mc_out[3]), .A2(sr_out[3]), .S0(n1), .Y(\_0_net_[3] )
         );
  MUX21X1_HVT U68 ( .A1(mc_out[39]), .A2(sr_out[39]), .S0(n1), .Y(
        \_0_net_[39] ) );
  MUX21X1_HVT U69 ( .A1(mc_out[38]), .A2(sr_out[38]), .S0(n1), .Y(
        \_0_net_[38] ) );
  MUX21X1_HVT U70 ( .A1(mc_out[37]), .A2(sr_out[37]), .S0(n1), .Y(
        \_0_net_[37] ) );
  MUX21X1_HVT U71 ( .A1(mc_out[36]), .A2(sr_out[36]), .S0(n1), .Y(
        \_0_net_[36] ) );
  MUX21X1_HVT U72 ( .A1(mc_out[35]), .A2(sr_out[35]), .S0(n1), .Y(
        \_0_net_[35] ) );
  MUX21X1_HVT U73 ( .A1(mc_out[34]), .A2(sr_out[34]), .S0(n1), .Y(
        \_0_net_[34] ) );
  MUX21X1_HVT U74 ( .A1(mc_out[33]), .A2(sr_out[33]), .S0(n1), .Y(
        \_0_net_[33] ) );
  MUX21X1_HVT U75 ( .A1(mc_out[32]), .A2(sr_out[32]), .S0(n1), .Y(
        \_0_net_[32] ) );
  MUX21X1_HVT U76 ( .A1(mc_out[31]), .A2(sr_out[31]), .S0(n1), .Y(
        \_0_net_[31] ) );
  MUX21X1_HVT U77 ( .A1(mc_out[30]), .A2(sr_out[30]), .S0(n1), .Y(
        \_0_net_[30] ) );
  MUX21X1_HVT U78 ( .A1(mc_out[2]), .A2(sr_out[2]), .S0(n1), .Y(\_0_net_[2] )
         );
  MUX21X1_HVT U79 ( .A1(mc_out[29]), .A2(sr_out[29]), .S0(n1), .Y(
        \_0_net_[29] ) );
  MUX21X1_HVT U80 ( .A1(mc_out[28]), .A2(sr_out[28]), .S0(n1), .Y(
        \_0_net_[28] ) );
  MUX21X1_HVT U81 ( .A1(mc_out[27]), .A2(sr_out[27]), .S0(n1), .Y(
        \_0_net_[27] ) );
  MUX21X1_HVT U82 ( .A1(mc_out[26]), .A2(sr_out[26]), .S0(n1), .Y(
        \_0_net_[26] ) );
  MUX21X1_HVT U83 ( .A1(mc_out[25]), .A2(sr_out[25]), .S0(n1), .Y(
        \_0_net_[25] ) );
  MUX21X1_HVT U84 ( .A1(mc_out[24]), .A2(sr_out[24]), .S0(n1), .Y(
        \_0_net_[24] ) );
  MUX21X1_HVT U85 ( .A1(mc_out[23]), .A2(sr_out[23]), .S0(n1), .Y(
        \_0_net_[23] ) );
  MUX21X1_HVT U86 ( .A1(mc_out[22]), .A2(sr_out[22]), .S0(n1), .Y(
        \_0_net_[22] ) );
  MUX21X1_HVT U87 ( .A1(mc_out[21]), .A2(sr_out[21]), .S0(n1), .Y(
        \_0_net_[21] ) );
  MUX21X1_HVT U88 ( .A1(mc_out[20]), .A2(sr_out[20]), .S0(n1), .Y(
        \_0_net_[20] ) );
  MUX21X1_HVT U89 ( .A1(mc_out[1]), .A2(sr_out[1]), .S0(n1), .Y(\_0_net_[1] )
         );
  MUX21X1_HVT U90 ( .A1(mc_out[19]), .A2(sr_out[19]), .S0(n1), .Y(
        \_0_net_[19] ) );
  MUX21X1_HVT U91 ( .A1(mc_out[18]), .A2(sr_out[18]), .S0(n1), .Y(
        \_0_net_[18] ) );
  MUX21X1_HVT U92 ( .A1(mc_out[17]), .A2(sr_out[17]), .S0(n1), .Y(
        \_0_net_[17] ) );
  MUX21X1_HVT U93 ( .A1(mc_out[16]), .A2(sr_out[16]), .S0(n1), .Y(
        \_0_net_[16] ) );
  MUX21X1_HVT U94 ( .A1(mc_out[15]), .A2(sr_out[15]), .S0(n1), .Y(
        \_0_net_[15] ) );
  MUX21X1_HVT U95 ( .A1(mc_out[14]), .A2(sr_out[14]), .S0(n1), .Y(
        \_0_net_[14] ) );
  MUX21X1_HVT U96 ( .A1(mc_out[13]), .A2(sr_out[13]), .S0(n1), .Y(
        \_0_net_[13] ) );
  MUX21X1_HVT U97 ( .A1(mc_out[12]), .A2(sr_out[12]), .S0(n1), .Y(
        \_0_net_[12] ) );
  MUX21X1_HVT U98 ( .A1(mc_out[127]), .A2(sr_out[127]), .S0(n1), .Y(
        \_0_net_[127] ) );
  MUX21X1_HVT U99 ( .A1(mc_out[126]), .A2(sr_out[126]), .S0(n1), .Y(
        \_0_net_[126] ) );
  MUX21X1_HVT U100 ( .A1(mc_out[125]), .A2(sr_out[125]), .S0(n1), .Y(
        \_0_net_[125] ) );
  MUX21X1_HVT U101 ( .A1(mc_out[124]), .A2(sr_out[124]), .S0(n1), .Y(
        \_0_net_[124] ) );
  MUX21X1_HVT U102 ( .A1(mc_out[123]), .A2(sr_out[123]), .S0(n1), .Y(
        \_0_net_[123] ) );
  MUX21X1_HVT U103 ( .A1(mc_out[122]), .A2(sr_out[122]), .S0(n1), .Y(
        \_0_net_[122] ) );
  MUX21X1_HVT U104 ( .A1(mc_out[121]), .A2(sr_out[121]), .S0(n1), .Y(
        \_0_net_[121] ) );
  MUX21X1_HVT U105 ( .A1(mc_out[120]), .A2(sr_out[120]), .S0(n1), .Y(
        \_0_net_[120] ) );
  MUX21X1_HVT U106 ( .A1(mc_out[11]), .A2(sr_out[11]), .S0(n1), .Y(
        \_0_net_[11] ) );
  MUX21X1_HVT U107 ( .A1(mc_out[119]), .A2(sr_out[119]), .S0(n1), .Y(
        \_0_net_[119] ) );
  MUX21X1_HVT U108 ( .A1(mc_out[118]), .A2(sr_out[118]), .S0(n1), .Y(
        \_0_net_[118] ) );
  MUX21X1_HVT U109 ( .A1(mc_out[117]), .A2(sr_out[117]), .S0(n1), .Y(
        \_0_net_[117] ) );
  MUX21X1_HVT U110 ( .A1(mc_out[116]), .A2(sr_out[116]), .S0(n1), .Y(
        \_0_net_[116] ) );
  MUX21X1_HVT U111 ( .A1(mc_out[115]), .A2(sr_out[115]), .S0(n1), .Y(
        \_0_net_[115] ) );
  MUX21X1_HVT U112 ( .A1(mc_out[114]), .A2(sr_out[114]), .S0(n1), .Y(
        \_0_net_[114] ) );
  MUX21X1_HVT U113 ( .A1(mc_out[113]), .A2(sr_out[113]), .S0(n1), .Y(
        \_0_net_[113] ) );
  MUX21X1_HVT U114 ( .A1(mc_out[112]), .A2(sr_out[112]), .S0(n1), .Y(
        \_0_net_[112] ) );
  MUX21X1_HVT U115 ( .A1(mc_out[111]), .A2(sr_out[111]), .S0(n1), .Y(
        \_0_net_[111] ) );
  MUX21X1_HVT U116 ( .A1(mc_out[110]), .A2(sr_out[110]), .S0(n1), .Y(
        \_0_net_[110] ) );
  MUX21X1_HVT U117 ( .A1(mc_out[10]), .A2(sr_out[10]), .S0(n1), .Y(
        \_0_net_[10] ) );
  MUX21X1_HVT U118 ( .A1(mc_out[109]), .A2(sr_out[109]), .S0(n1), .Y(
        \_0_net_[109] ) );
  MUX21X1_HVT U119 ( .A1(mc_out[108]), .A2(sr_out[108]), .S0(n1), .Y(
        \_0_net_[108] ) );
  MUX21X1_HVT U120 ( .A1(mc_out[107]), .A2(sr_out[107]), .S0(n1), .Y(
        \_0_net_[107] ) );
  MUX21X1_HVT U121 ( .A1(mc_out[106]), .A2(sr_out[106]), .S0(n1), .Y(
        \_0_net_[106] ) );
  MUX21X1_HVT U122 ( .A1(mc_out[105]), .A2(sr_out[105]), .S0(n1), .Y(
        \_0_net_[105] ) );
  MUX21X1_HVT U123 ( .A1(mc_out[104]), .A2(sr_out[104]), .S0(n1), .Y(
        \_0_net_[104] ) );
  MUX21X1_HVT U124 ( .A1(mc_out[103]), .A2(sr_out[103]), .S0(n1), .Y(
        \_0_net_[103] ) );
  MUX21X1_HVT U125 ( .A1(mc_out[102]), .A2(sr_out[102]), .S0(n1), .Y(
        \_0_net_[102] ) );
  MUX21X1_HVT U126 ( .A1(mc_out[101]), .A2(sr_out[101]), .S0(n1), .Y(
        \_0_net_[101] ) );
  MUX21X1_HVT U127 ( .A1(mc_out[100]), .A2(sr_out[100]), .S0(n1), .Y(
        \_0_net_[100] ) );
  MUX21X1_HVT U128 ( .A1(mc_out[0]), .A2(sr_out[0]), .S0(n1), .Y(\_0_net_[0] )
         );
  NOR3X0_HVT U129 ( .A1(round_num[2]), .A2(round_num[0]), .A3(n2), .Y(n1) );
  NAND2X0_HVT U130 ( .A1(round_num[3]), .A2(round_num[1]), .Y(n2) );
endmodule

