
module cam_DATA_WIDTH128_ADDR_WIDTH4 ( clk, rst, start, write_enable, din, 
        write_addr, match, match_addr );
  input [127:0] din;
  input [3:0] write_addr;
  output [3:0] match_addr;
  input clk, rst, start, write_enable;
  output match;
  wire   \match_addr_unencoded_raw[31][15] ,
         \match_addr_unencoded_raw[31][14] ,
         \match_addr_unencoded_raw[31][13] ,
         \match_addr_unencoded_raw[31][12] ,
         \match_addr_unencoded_raw[31][11] ,
         \match_addr_unencoded_raw[31][10] , \match_addr_unencoded_raw[31][9] ,
         \match_addr_unencoded_raw[31][8] , \match_addr_unencoded_raw[31][7] ,
         \match_addr_unencoded_raw[31][6] , \match_addr_unencoded_raw[31][5] ,
         \match_addr_unencoded_raw[31][4] , \match_addr_unencoded_raw[31][3] ,
         \match_addr_unencoded_raw[31][2] , \match_addr_unencoded_raw[31][1] ,
         \match_addr_unencoded_raw[31][0] , \match_addr_unencoded_raw[30][15] ,
         \match_addr_unencoded_raw[30][14] ,
         \match_addr_unencoded_raw[30][13] ,
         \match_addr_unencoded_raw[30][12] ,
         \match_addr_unencoded_raw[30][11] ,
         \match_addr_unencoded_raw[30][10] , \match_addr_unencoded_raw[30][9] ,
         \match_addr_unencoded_raw[30][8] , \match_addr_unencoded_raw[30][7] ,
         \match_addr_unencoded_raw[30][6] , \match_addr_unencoded_raw[30][5] ,
         \match_addr_unencoded_raw[30][4] , \match_addr_unencoded_raw[30][3] ,
         \match_addr_unencoded_raw[30][2] , \match_addr_unencoded_raw[30][1] ,
         \match_addr_unencoded_raw[30][0] , \match_addr_unencoded_raw[29][15] ,
         \match_addr_unencoded_raw[29][14] ,
         \match_addr_unencoded_raw[29][13] ,
         \match_addr_unencoded_raw[29][12] ,
         \match_addr_unencoded_raw[29][11] ,
         \match_addr_unencoded_raw[29][10] , \match_addr_unencoded_raw[29][9] ,
         \match_addr_unencoded_raw[29][8] , \match_addr_unencoded_raw[29][7] ,
         \match_addr_unencoded_raw[29][6] , \match_addr_unencoded_raw[29][5] ,
         \match_addr_unencoded_raw[29][4] , \match_addr_unencoded_raw[29][3] ,
         \match_addr_unencoded_raw[29][2] , \match_addr_unencoded_raw[29][1] ,
         \match_addr_unencoded_raw[29][0] , \match_addr_unencoded_raw[28][15] ,
         \match_addr_unencoded_raw[28][14] ,
         \match_addr_unencoded_raw[28][13] ,
         \match_addr_unencoded_raw[28][12] ,
         \match_addr_unencoded_raw[28][11] ,
         \match_addr_unencoded_raw[28][10] , \match_addr_unencoded_raw[28][9] ,
         \match_addr_unencoded_raw[28][8] , \match_addr_unencoded_raw[28][7] ,
         \match_addr_unencoded_raw[28][6] , \match_addr_unencoded_raw[28][5] ,
         \match_addr_unencoded_raw[28][4] , \match_addr_unencoded_raw[28][3] ,
         \match_addr_unencoded_raw[28][2] , \match_addr_unencoded_raw[28][1] ,
         \match_addr_unencoded_raw[28][0] , \match_addr_unencoded_raw[27][15] ,
         \match_addr_unencoded_raw[27][14] ,
         \match_addr_unencoded_raw[27][13] ,
         \match_addr_unencoded_raw[27][12] ,
         \match_addr_unencoded_raw[27][11] ,
         \match_addr_unencoded_raw[27][10] , \match_addr_unencoded_raw[27][9] ,
         \match_addr_unencoded_raw[27][8] , \match_addr_unencoded_raw[27][7] ,
         \match_addr_unencoded_raw[27][6] , \match_addr_unencoded_raw[27][5] ,
         \match_addr_unencoded_raw[27][4] , \match_addr_unencoded_raw[27][3] ,
         \match_addr_unencoded_raw[27][2] , \match_addr_unencoded_raw[27][1] ,
         \match_addr_unencoded_raw[27][0] , \match_addr_unencoded_raw[26][15] ,
         \match_addr_unencoded_raw[26][14] ,
         \match_addr_unencoded_raw[26][13] ,
         \match_addr_unencoded_raw[26][12] ,
         \match_addr_unencoded_raw[26][11] ,
         \match_addr_unencoded_raw[26][10] , \match_addr_unencoded_raw[26][9] ,
         \match_addr_unencoded_raw[26][8] , \match_addr_unencoded_raw[26][7] ,
         \match_addr_unencoded_raw[26][6] , \match_addr_unencoded_raw[26][5] ,
         \match_addr_unencoded_raw[26][4] , \match_addr_unencoded_raw[26][3] ,
         \match_addr_unencoded_raw[26][2] , \match_addr_unencoded_raw[26][1] ,
         \match_addr_unencoded_raw[26][0] , \match_addr_unencoded_raw[25][15] ,
         \match_addr_unencoded_raw[25][14] ,
         \match_addr_unencoded_raw[25][13] ,
         \match_addr_unencoded_raw[25][12] ,
         \match_addr_unencoded_raw[25][11] ,
         \match_addr_unencoded_raw[25][10] , \match_addr_unencoded_raw[25][9] ,
         \match_addr_unencoded_raw[25][8] , \match_addr_unencoded_raw[25][7] ,
         \match_addr_unencoded_raw[25][6] , \match_addr_unencoded_raw[25][5] ,
         \match_addr_unencoded_raw[25][4] , \match_addr_unencoded_raw[25][3] ,
         \match_addr_unencoded_raw[25][2] , \match_addr_unencoded_raw[25][1] ,
         \match_addr_unencoded_raw[25][0] , \match_addr_unencoded_raw[24][15] ,
         \match_addr_unencoded_raw[24][14] ,
         \match_addr_unencoded_raw[24][13] ,
         \match_addr_unencoded_raw[24][12] ,
         \match_addr_unencoded_raw[24][11] ,
         \match_addr_unencoded_raw[24][10] , \match_addr_unencoded_raw[24][9] ,
         \match_addr_unencoded_raw[24][8] , \match_addr_unencoded_raw[24][7] ,
         \match_addr_unencoded_raw[24][6] , \match_addr_unencoded_raw[24][5] ,
         \match_addr_unencoded_raw[24][4] , \match_addr_unencoded_raw[24][3] ,
         \match_addr_unencoded_raw[24][2] , \match_addr_unencoded_raw[24][1] ,
         \match_addr_unencoded_raw[24][0] , \match_addr_unencoded_raw[23][15] ,
         \match_addr_unencoded_raw[23][14] ,
         \match_addr_unencoded_raw[23][13] ,
         \match_addr_unencoded_raw[23][12] ,
         \match_addr_unencoded_raw[23][11] ,
         \match_addr_unencoded_raw[23][10] , \match_addr_unencoded_raw[23][9] ,
         \match_addr_unencoded_raw[23][8] , \match_addr_unencoded_raw[23][7] ,
         \match_addr_unencoded_raw[23][6] , \match_addr_unencoded_raw[23][5] ,
         \match_addr_unencoded_raw[23][4] , \match_addr_unencoded_raw[23][3] ,
         \match_addr_unencoded_raw[23][2] , \match_addr_unencoded_raw[23][1] ,
         \match_addr_unencoded_raw[23][0] , \match_addr_unencoded_raw[22][15] ,
         \match_addr_unencoded_raw[22][14] ,
         \match_addr_unencoded_raw[22][13] ,
         \match_addr_unencoded_raw[22][12] ,
         \match_addr_unencoded_raw[22][11] ,
         \match_addr_unencoded_raw[22][10] , \match_addr_unencoded_raw[22][9] ,
         \match_addr_unencoded_raw[22][8] , \match_addr_unencoded_raw[22][7] ,
         \match_addr_unencoded_raw[22][6] , \match_addr_unencoded_raw[22][5] ,
         \match_addr_unencoded_raw[22][4] , \match_addr_unencoded_raw[22][3] ,
         \match_addr_unencoded_raw[22][2] , \match_addr_unencoded_raw[22][1] ,
         \match_addr_unencoded_raw[22][0] , \match_addr_unencoded_raw[21][15] ,
         \match_addr_unencoded_raw[21][14] ,
         \match_addr_unencoded_raw[21][13] ,
         \match_addr_unencoded_raw[21][12] ,
         \match_addr_unencoded_raw[21][11] ,
         \match_addr_unencoded_raw[21][10] , \match_addr_unencoded_raw[21][9] ,
         \match_addr_unencoded_raw[21][8] , \match_addr_unencoded_raw[21][7] ,
         \match_addr_unencoded_raw[21][6] , \match_addr_unencoded_raw[21][5] ,
         \match_addr_unencoded_raw[21][4] , \match_addr_unencoded_raw[21][3] ,
         \match_addr_unencoded_raw[21][2] , \match_addr_unencoded_raw[21][1] ,
         \match_addr_unencoded_raw[21][0] , \match_addr_unencoded_raw[20][15] ,
         \match_addr_unencoded_raw[20][14] ,
         \match_addr_unencoded_raw[20][13] ,
         \match_addr_unencoded_raw[20][12] ,
         \match_addr_unencoded_raw[20][11] ,
         \match_addr_unencoded_raw[20][10] , \match_addr_unencoded_raw[20][9] ,
         \match_addr_unencoded_raw[20][8] , \match_addr_unencoded_raw[20][7] ,
         \match_addr_unencoded_raw[20][6] , \match_addr_unencoded_raw[20][5] ,
         \match_addr_unencoded_raw[20][4] , \match_addr_unencoded_raw[20][3] ,
         \match_addr_unencoded_raw[20][2] , \match_addr_unencoded_raw[20][1] ,
         \match_addr_unencoded_raw[20][0] , \match_addr_unencoded_raw[19][15] ,
         \match_addr_unencoded_raw[19][14] ,
         \match_addr_unencoded_raw[19][13] ,
         \match_addr_unencoded_raw[19][12] ,
         \match_addr_unencoded_raw[19][11] ,
         \match_addr_unencoded_raw[19][10] , \match_addr_unencoded_raw[19][9] ,
         \match_addr_unencoded_raw[19][8] , \match_addr_unencoded_raw[19][7] ,
         \match_addr_unencoded_raw[19][6] , \match_addr_unencoded_raw[19][5] ,
         \match_addr_unencoded_raw[19][4] , \match_addr_unencoded_raw[19][3] ,
         \match_addr_unencoded_raw[19][2] , \match_addr_unencoded_raw[19][1] ,
         \match_addr_unencoded_raw[19][0] , \match_addr_unencoded_raw[18][15] ,
         \match_addr_unencoded_raw[18][14] ,
         \match_addr_unencoded_raw[18][13] ,
         \match_addr_unencoded_raw[18][12] ,
         \match_addr_unencoded_raw[18][11] ,
         \match_addr_unencoded_raw[18][10] , \match_addr_unencoded_raw[18][9] ,
         \match_addr_unencoded_raw[18][8] , \match_addr_unencoded_raw[18][7] ,
         \match_addr_unencoded_raw[18][6] , \match_addr_unencoded_raw[18][5] ,
         \match_addr_unencoded_raw[18][4] , \match_addr_unencoded_raw[18][3] ,
         \match_addr_unencoded_raw[18][2] , \match_addr_unencoded_raw[18][1] ,
         \match_addr_unencoded_raw[18][0] , \match_addr_unencoded_raw[17][15] ,
         \match_addr_unencoded_raw[17][14] ,
         \match_addr_unencoded_raw[17][13] ,
         \match_addr_unencoded_raw[17][12] ,
         \match_addr_unencoded_raw[17][11] ,
         \match_addr_unencoded_raw[17][10] , \match_addr_unencoded_raw[17][9] ,
         \match_addr_unencoded_raw[17][8] , \match_addr_unencoded_raw[17][7] ,
         \match_addr_unencoded_raw[17][6] , \match_addr_unencoded_raw[17][5] ,
         \match_addr_unencoded_raw[17][4] , \match_addr_unencoded_raw[17][3] ,
         \match_addr_unencoded_raw[17][2] , \match_addr_unencoded_raw[17][1] ,
         \match_addr_unencoded_raw[17][0] , \match_addr_unencoded_raw[16][15] ,
         \match_addr_unencoded_raw[16][14] ,
         \match_addr_unencoded_raw[16][13] ,
         \match_addr_unencoded_raw[16][12] ,
         \match_addr_unencoded_raw[16][11] ,
         \match_addr_unencoded_raw[16][10] , \match_addr_unencoded_raw[16][9] ,
         \match_addr_unencoded_raw[16][8] , \match_addr_unencoded_raw[16][7] ,
         \match_addr_unencoded_raw[16][6] , \match_addr_unencoded_raw[16][5] ,
         \match_addr_unencoded_raw[16][4] , \match_addr_unencoded_raw[16][3] ,
         \match_addr_unencoded_raw[16][2] , \match_addr_unencoded_raw[16][1] ,
         \match_addr_unencoded_raw[16][0] , \match_addr_unencoded_raw[15][15] ,
         \match_addr_unencoded_raw[15][14] ,
         \match_addr_unencoded_raw[15][13] ,
         \match_addr_unencoded_raw[15][12] ,
         \match_addr_unencoded_raw[15][11] ,
         \match_addr_unencoded_raw[15][10] , \match_addr_unencoded_raw[15][9] ,
         \match_addr_unencoded_raw[15][8] , \match_addr_unencoded_raw[15][7] ,
         \match_addr_unencoded_raw[15][6] , \match_addr_unencoded_raw[15][5] ,
         \match_addr_unencoded_raw[15][4] , \match_addr_unencoded_raw[15][3] ,
         \match_addr_unencoded_raw[15][2] , \match_addr_unencoded_raw[15][1] ,
         \match_addr_unencoded_raw[15][0] , \match_addr_unencoded_raw[14][15] ,
         \match_addr_unencoded_raw[14][14] ,
         \match_addr_unencoded_raw[14][13] ,
         \match_addr_unencoded_raw[14][12] ,
         \match_addr_unencoded_raw[14][11] ,
         \match_addr_unencoded_raw[14][10] , \match_addr_unencoded_raw[14][9] ,
         \match_addr_unencoded_raw[14][8] , \match_addr_unencoded_raw[14][7] ,
         \match_addr_unencoded_raw[14][6] , \match_addr_unencoded_raw[14][5] ,
         \match_addr_unencoded_raw[14][4] , \match_addr_unencoded_raw[14][3] ,
         \match_addr_unencoded_raw[14][2] , \match_addr_unencoded_raw[14][1] ,
         \match_addr_unencoded_raw[14][0] , \match_addr_unencoded_raw[13][15] ,
         \match_addr_unencoded_raw[13][14] ,
         \match_addr_unencoded_raw[13][13] ,
         \match_addr_unencoded_raw[13][12] ,
         \match_addr_unencoded_raw[13][11] ,
         \match_addr_unencoded_raw[13][10] , \match_addr_unencoded_raw[13][9] ,
         \match_addr_unencoded_raw[13][8] , \match_addr_unencoded_raw[13][7] ,
         \match_addr_unencoded_raw[13][6] , \match_addr_unencoded_raw[13][5] ,
         \match_addr_unencoded_raw[13][4] , \match_addr_unencoded_raw[13][3] ,
         \match_addr_unencoded_raw[13][2] , \match_addr_unencoded_raw[13][1] ,
         \match_addr_unencoded_raw[13][0] , \match_addr_unencoded_raw[12][15] ,
         \match_addr_unencoded_raw[12][14] ,
         \match_addr_unencoded_raw[12][13] ,
         \match_addr_unencoded_raw[12][12] ,
         \match_addr_unencoded_raw[12][11] ,
         \match_addr_unencoded_raw[12][10] , \match_addr_unencoded_raw[12][9] ,
         \match_addr_unencoded_raw[12][8] , \match_addr_unencoded_raw[12][7] ,
         \match_addr_unencoded_raw[12][6] , \match_addr_unencoded_raw[12][5] ,
         \match_addr_unencoded_raw[12][4] , \match_addr_unencoded_raw[12][3] ,
         \match_addr_unencoded_raw[12][2] , \match_addr_unencoded_raw[12][1] ,
         \match_addr_unencoded_raw[12][0] , \match_addr_unencoded_raw[11][15] ,
         \match_addr_unencoded_raw[11][14] ,
         \match_addr_unencoded_raw[11][13] ,
         \match_addr_unencoded_raw[11][12] ,
         \match_addr_unencoded_raw[11][11] ,
         \match_addr_unencoded_raw[11][10] , \match_addr_unencoded_raw[11][9] ,
         \match_addr_unencoded_raw[11][8] , \match_addr_unencoded_raw[11][7] ,
         \match_addr_unencoded_raw[11][6] , \match_addr_unencoded_raw[11][5] ,
         \match_addr_unencoded_raw[11][4] , \match_addr_unencoded_raw[11][3] ,
         \match_addr_unencoded_raw[11][2] , \match_addr_unencoded_raw[11][1] ,
         \match_addr_unencoded_raw[11][0] , \match_addr_unencoded_raw[10][15] ,
         \match_addr_unencoded_raw[10][14] ,
         \match_addr_unencoded_raw[10][13] ,
         \match_addr_unencoded_raw[10][12] ,
         \match_addr_unencoded_raw[10][11] ,
         \match_addr_unencoded_raw[10][10] , \match_addr_unencoded_raw[10][9] ,
         \match_addr_unencoded_raw[10][8] , \match_addr_unencoded_raw[10][7] ,
         \match_addr_unencoded_raw[10][6] , \match_addr_unencoded_raw[10][5] ,
         \match_addr_unencoded_raw[10][4] , \match_addr_unencoded_raw[10][3] ,
         \match_addr_unencoded_raw[10][2] , \match_addr_unencoded_raw[10][1] ,
         \match_addr_unencoded_raw[10][0] , \match_addr_unencoded_raw[9][15] ,
         \match_addr_unencoded_raw[9][14] , \match_addr_unencoded_raw[9][13] ,
         \match_addr_unencoded_raw[9][12] , \match_addr_unencoded_raw[9][11] ,
         \match_addr_unencoded_raw[9][10] , \match_addr_unencoded_raw[9][9] ,
         \match_addr_unencoded_raw[9][8] , \match_addr_unencoded_raw[9][7] ,
         \match_addr_unencoded_raw[9][6] , \match_addr_unencoded_raw[9][5] ,
         \match_addr_unencoded_raw[9][4] , \match_addr_unencoded_raw[9][3] ,
         \match_addr_unencoded_raw[9][2] , \match_addr_unencoded_raw[9][1] ,
         \match_addr_unencoded_raw[9][0] , \match_addr_unencoded_raw[8][15] ,
         \match_addr_unencoded_raw[8][14] , \match_addr_unencoded_raw[8][13] ,
         \match_addr_unencoded_raw[8][12] , \match_addr_unencoded_raw[8][11] ,
         \match_addr_unencoded_raw[8][10] , \match_addr_unencoded_raw[8][9] ,
         \match_addr_unencoded_raw[8][8] , \match_addr_unencoded_raw[8][7] ,
         \match_addr_unencoded_raw[8][6] , \match_addr_unencoded_raw[8][5] ,
         \match_addr_unencoded_raw[8][4] , \match_addr_unencoded_raw[8][3] ,
         \match_addr_unencoded_raw[8][2] , \match_addr_unencoded_raw[8][1] ,
         \match_addr_unencoded_raw[8][0] , \match_addr_unencoded_raw[7][15] ,
         \match_addr_unencoded_raw[7][14] , \match_addr_unencoded_raw[7][13] ,
         \match_addr_unencoded_raw[7][12] , \match_addr_unencoded_raw[7][11] ,
         \match_addr_unencoded_raw[7][10] , \match_addr_unencoded_raw[7][9] ,
         \match_addr_unencoded_raw[7][8] , \match_addr_unencoded_raw[7][7] ,
         \match_addr_unencoded_raw[7][6] , \match_addr_unencoded_raw[7][5] ,
         \match_addr_unencoded_raw[7][4] , \match_addr_unencoded_raw[7][3] ,
         \match_addr_unencoded_raw[7][2] , \match_addr_unencoded_raw[7][1] ,
         \match_addr_unencoded_raw[7][0] , \match_addr_unencoded_raw[6][15] ,
         \match_addr_unencoded_raw[6][14] , \match_addr_unencoded_raw[6][13] ,
         \match_addr_unencoded_raw[6][12] , \match_addr_unencoded_raw[6][11] ,
         \match_addr_unencoded_raw[6][10] , \match_addr_unencoded_raw[6][9] ,
         \match_addr_unencoded_raw[6][8] , \match_addr_unencoded_raw[6][7] ,
         \match_addr_unencoded_raw[6][6] , \match_addr_unencoded_raw[6][5] ,
         \match_addr_unencoded_raw[6][4] , \match_addr_unencoded_raw[6][3] ,
         \match_addr_unencoded_raw[6][2] , \match_addr_unencoded_raw[6][1] ,
         \match_addr_unencoded_raw[6][0] , \match_addr_unencoded_raw[5][15] ,
         \match_addr_unencoded_raw[5][14] , \match_addr_unencoded_raw[5][13] ,
         \match_addr_unencoded_raw[5][12] , \match_addr_unencoded_raw[5][11] ,
         \match_addr_unencoded_raw[5][10] , \match_addr_unencoded_raw[5][9] ,
         \match_addr_unencoded_raw[5][8] , \match_addr_unencoded_raw[5][7] ,
         \match_addr_unencoded_raw[5][6] , \match_addr_unencoded_raw[5][5] ,
         \match_addr_unencoded_raw[5][4] , \match_addr_unencoded_raw[5][3] ,
         \match_addr_unencoded_raw[5][2] , \match_addr_unencoded_raw[5][1] ,
         \match_addr_unencoded_raw[5][0] , \match_addr_unencoded_raw[4][15] ,
         \match_addr_unencoded_raw[4][14] , \match_addr_unencoded_raw[4][13] ,
         \match_addr_unencoded_raw[4][12] , \match_addr_unencoded_raw[4][11] ,
         \match_addr_unencoded_raw[4][10] , \match_addr_unencoded_raw[4][9] ,
         \match_addr_unencoded_raw[4][8] , \match_addr_unencoded_raw[4][7] ,
         \match_addr_unencoded_raw[4][6] , \match_addr_unencoded_raw[4][5] ,
         \match_addr_unencoded_raw[4][4] , \match_addr_unencoded_raw[4][3] ,
         \match_addr_unencoded_raw[4][2] , \match_addr_unencoded_raw[4][1] ,
         \match_addr_unencoded_raw[4][0] , \match_addr_unencoded_raw[3][15] ,
         \match_addr_unencoded_raw[3][14] , \match_addr_unencoded_raw[3][13] ,
         \match_addr_unencoded_raw[3][12] , \match_addr_unencoded_raw[3][11] ,
         \match_addr_unencoded_raw[3][10] , \match_addr_unencoded_raw[3][9] ,
         \match_addr_unencoded_raw[3][8] , \match_addr_unencoded_raw[3][7] ,
         \match_addr_unencoded_raw[3][6] , \match_addr_unencoded_raw[3][5] ,
         \match_addr_unencoded_raw[3][4] , \match_addr_unencoded_raw[3][3] ,
         \match_addr_unencoded_raw[3][2] , \match_addr_unencoded_raw[3][1] ,
         \match_addr_unencoded_raw[3][0] , \match_addr_unencoded_raw[2][15] ,
         \match_addr_unencoded_raw[2][14] , \match_addr_unencoded_raw[2][13] ,
         \match_addr_unencoded_raw[2][12] , \match_addr_unencoded_raw[2][11] ,
         \match_addr_unencoded_raw[2][10] , \match_addr_unencoded_raw[2][9] ,
         \match_addr_unencoded_raw[2][8] , \match_addr_unencoded_raw[2][7] ,
         \match_addr_unencoded_raw[2][6] , \match_addr_unencoded_raw[2][5] ,
         \match_addr_unencoded_raw[2][4] , \match_addr_unencoded_raw[2][3] ,
         \match_addr_unencoded_raw[2][2] , \match_addr_unencoded_raw[2][1] ,
         \match_addr_unencoded_raw[2][0] , \match_addr_unencoded_raw[1][15] ,
         \match_addr_unencoded_raw[1][14] , \match_addr_unencoded_raw[1][13] ,
         \match_addr_unencoded_raw[1][12] , \match_addr_unencoded_raw[1][11] ,
         \match_addr_unencoded_raw[1][10] , \match_addr_unencoded_raw[1][9] ,
         \match_addr_unencoded_raw[1][8] , \match_addr_unencoded_raw[1][7] ,
         \match_addr_unencoded_raw[1][6] , \match_addr_unencoded_raw[1][5] ,
         \match_addr_unencoded_raw[1][4] , \match_addr_unencoded_raw[1][3] ,
         \match_addr_unencoded_raw[1][2] , \match_addr_unencoded_raw[1][1] ,
         \match_addr_unencoded_raw[1][0] , \match_addr_unencoded_raw[0][15] ,
         \match_addr_unencoded_raw[0][14] , \match_addr_unencoded_raw[0][13] ,
         \match_addr_unencoded_raw[0][12] , \match_addr_unencoded_raw[0][11] ,
         \match_addr_unencoded_raw[0][10] , \match_addr_unencoded_raw[0][9] ,
         \match_addr_unencoded_raw[0][8] , \match_addr_unencoded_raw[0][7] ,
         \match_addr_unencoded_raw[0][6] , \match_addr_unencoded_raw[0][5] ,
         \match_addr_unencoded_raw[0][4] , \match_addr_unencoded_raw[0][3] ,
         \match_addr_unencoded_raw[0][2] , \match_addr_unencoded_raw[0][1] ,
         \match_addr_unencoded_raw[0][0] , N3, N4, N5, N6, N7, n1, n2, n3, n4,
         n5, n6, n11, n12, n13, n14, n15, n16, n25, n26, n27, n31, n32, n33,
         n34, n35, n36, n45, n46, n47, n51, n52, n53, n54, n55, n56, n65, n66,
         n67, n71, n72, n73, n74, n75, n76, n85, n86, n87, n91, n92, n93, n94,
         n95, n96, n101, n102, n103, n104, n105, n106, n111, n112, n113, n114,
         n115, n116, n121, n122, n123, n124, n125, n126, n131, n132, n133,
         n134, n135, n136, n141, n142, n143, n144, n145, n146, n151, n152,
         n153, n154, n155, n156, n7, n8, n9, n10, n17, n18, n19, n20, n21, n22,
         n23, n24, n28, n29, n30, n37, n38, n39, n40, n41, n42, n43, n44, n48,
         n49, n50, n57, n58, n59, n60, n61, n62, n63, n64, n68, n69, n70, n77,
         n78, n79, n80, n81, n82, n83, n84, n88, n89, n90, n97, n98, n99, n100,
         n107, n108, n109, n110, n117, n118, n119, n120, n127, n128, n129,
         n130, n137, n138, n139, n140, n147, n148, n149, n150, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196;
  wire   [15:0] match_addr_unencoded;
  wire   [3:0] match_addr_w;

  LATCHX1_HVT \match_addr_reg[3]  ( .CLK(N3), .D(N7), .Q(match_addr[3]) );
  LATCHX1_HVT \match_addr_reg[2]  ( .CLK(N3), .D(N6), .Q(match_addr[2]) );
  LATCHX1_HVT \match_addr_reg[1]  ( .CLK(N3), .D(N5), .Q(match_addr[1]) );
  LATCHX1_HVT \match_addr_reg[0]  ( .CLK(N3), .D(N4), .Q(match_addr[0]) );
  NOR4X1_HVT U2 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .Y(
        match_addr_unencoded[9]) );
  NOR4X1_HVT U4 ( .A1(n11), .A2(n12), .A3(n13), .A4(n14), .Y(
        match_addr_unencoded[8]) );
  NOR4X1_HVT U8 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .Y(
        match_addr_unencoded[6]) );
  NOR4X1_HVT U12 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .Y(
        match_addr_unencoded[4]) );
  NOR4X1_HVT U16 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .Y(
        match_addr_unencoded[2]) );
  NOR4X1_HVT U20 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .Y(
        match_addr_unencoded[15]) );
  NOR4X1_HVT U22 ( .A1(n101), .A2(n102), .A3(n103), .A4(n104), .Y(
        match_addr_unencoded[14]) );
  NOR4X1_HVT U24 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .Y(
        match_addr_unencoded[13]) );
  NOR4X1_HVT U26 ( .A1(n121), .A2(n122), .A3(n123), .A4(n124), .Y(
        match_addr_unencoded[12]) );
  NOR4X1_HVT U28 ( .A1(n131), .A2(n132), .A3(n133), .A4(n134), .Y(
        match_addr_unencoded[11]) );
  NOR4X1_HVT U30 ( .A1(n141), .A2(n142), .A3(n143), .A4(n144), .Y(
        match_addr_unencoded[10]) );
  NOR4X1_HVT U32 ( .A1(n151), .A2(n152), .A3(n153), .A4(n154), .Y(
        match_addr_unencoded[0]) );
  NAND4X0_HVT U34 ( .A1(\match_addr_unencoded_raw[24][9] ), .A2(
        \match_addr_unencoded_raw[23][9] ), .A3(
        \match_addr_unencoded_raw[22][9] ), .A4(
        \match_addr_unencoded_raw[21][9] ), .Y(n4) );
  NAND4X0_HVT U35 ( .A1(\match_addr_unencoded_raw[20][9] ), .A2(
        \match_addr_unencoded_raw[1][9] ), .A3(
        \match_addr_unencoded_raw[19][9] ), .A4(
        \match_addr_unencoded_raw[18][9] ), .Y(n3) );
  NAND4X0_HVT U36 ( .A1(\match_addr_unencoded_raw[13][9] ), .A2(
        \match_addr_unencoded_raw[12][9] ), .A3(n5), .A4(n6), .Y(n2) );
  AND4X1_HVT U37 ( .A1(\match_addr_unencoded_raw[17][9] ), .A2(
        \match_addr_unencoded_raw[16][9] ), .A3(
        \match_addr_unencoded_raw[15][9] ), .A4(
        \match_addr_unencoded_raw[14][9] ), .Y(n6) );
  AND3X1_HVT U38 ( .A1(\match_addr_unencoded_raw[10][9] ), .A2(
        \match_addr_unencoded_raw[0][9] ), .A3(
        \match_addr_unencoded_raw[11][9] ), .Y(n5) );
  NAND4X0_HVT U43 ( .A1(\match_addr_unencoded_raw[23][8] ), .A2(
        \match_addr_unencoded_raw[22][8] ), .A3(
        \match_addr_unencoded_raw[21][8] ), .A4(
        \match_addr_unencoded_raw[20][8] ), .Y(n14) );
  NAND4X0_HVT U44 ( .A1(\match_addr_unencoded_raw[1][8] ), .A2(
        \match_addr_unencoded_raw[19][8] ), .A3(
        \match_addr_unencoded_raw[18][8] ), .A4(
        \match_addr_unencoded_raw[17][8] ), .Y(n13) );
  NAND4X0_HVT U45 ( .A1(\match_addr_unencoded_raw[12][8] ), .A2(
        \match_addr_unencoded_raw[11][8] ), .A3(n15), .A4(n16), .Y(n12) );
  AND4X1_HVT U46 ( .A1(\match_addr_unencoded_raw[16][8] ), .A2(
        \match_addr_unencoded_raw[15][8] ), .A3(
        \match_addr_unencoded_raw[14][8] ), .A4(
        \match_addr_unencoded_raw[13][8] ), .Y(n16) );
  AND3X1_HVT U47 ( .A1(\match_addr_unencoded_raw[0][8] ), .A2(start), .A3(
        \match_addr_unencoded_raw[10][8] ), .Y(n15) );
  AND4X1_HVT U55 ( .A1(\match_addr_unencoded_raw[16][7] ), .A2(
        \match_addr_unencoded_raw[15][7] ), .A3(
        \match_addr_unencoded_raw[14][7] ), .A4(
        \match_addr_unencoded_raw[13][7] ), .Y(n26) );
  AND3X1_HVT U56 ( .A1(\match_addr_unencoded_raw[0][7] ), .A2(n175), .A3(
        \match_addr_unencoded_raw[10][7] ), .Y(n25) );
  NAND4X0_HVT U60 ( .A1(\match_addr_unencoded_raw[5][7] ), .A2(
        \match_addr_unencoded_raw[4][7] ), .A3(
        \match_addr_unencoded_raw[3][7] ), .A4(
        \match_addr_unencoded_raw[31][7] ), .Y(n27) );
  NAND4X0_HVT U61 ( .A1(\match_addr_unencoded_raw[23][6] ), .A2(
        \match_addr_unencoded_raw[22][6] ), .A3(
        \match_addr_unencoded_raw[21][6] ), .A4(
        \match_addr_unencoded_raw[20][6] ), .Y(n34) );
  NAND4X0_HVT U62 ( .A1(\match_addr_unencoded_raw[1][6] ), .A2(
        \match_addr_unencoded_raw[19][6] ), .A3(
        \match_addr_unencoded_raw[18][6] ), .A4(
        \match_addr_unencoded_raw[17][6] ), .Y(n33) );
  NAND4X0_HVT U63 ( .A1(\match_addr_unencoded_raw[12][6] ), .A2(
        \match_addr_unencoded_raw[11][6] ), .A3(n35), .A4(n36), .Y(n32) );
  AND4X1_HVT U64 ( .A1(\match_addr_unencoded_raw[16][6] ), .A2(
        \match_addr_unencoded_raw[15][6] ), .A3(
        \match_addr_unencoded_raw[14][6] ), .A4(
        \match_addr_unencoded_raw[13][6] ), .Y(n36) );
  AND3X1_HVT U65 ( .A1(\match_addr_unencoded_raw[0][6] ), .A2(n176), .A3(
        \match_addr_unencoded_raw[10][6] ), .Y(n35) );
  AND4X1_HVT U73 ( .A1(\match_addr_unencoded_raw[16][5] ), .A2(
        \match_addr_unencoded_raw[15][5] ), .A3(
        \match_addr_unencoded_raw[14][5] ), .A4(
        \match_addr_unencoded_raw[13][5] ), .Y(n46) );
  AND3X1_HVT U74 ( .A1(\match_addr_unencoded_raw[0][5] ), .A2(start), .A3(
        \match_addr_unencoded_raw[10][5] ), .Y(n45) );
  NAND4X0_HVT U78 ( .A1(\match_addr_unencoded_raw[5][5] ), .A2(
        \match_addr_unencoded_raw[4][5] ), .A3(
        \match_addr_unencoded_raw[3][5] ), .A4(
        \match_addr_unencoded_raw[31][5] ), .Y(n47) );
  NAND4X0_HVT U79 ( .A1(\match_addr_unencoded_raw[23][4] ), .A2(
        \match_addr_unencoded_raw[22][4] ), .A3(
        \match_addr_unencoded_raw[21][4] ), .A4(
        \match_addr_unencoded_raw[20][4] ), .Y(n54) );
  NAND4X0_HVT U80 ( .A1(\match_addr_unencoded_raw[1][4] ), .A2(
        \match_addr_unencoded_raw[19][4] ), .A3(
        \match_addr_unencoded_raw[18][4] ), .A4(
        \match_addr_unencoded_raw[17][4] ), .Y(n53) );
  NAND4X0_HVT U81 ( .A1(\match_addr_unencoded_raw[12][4] ), .A2(
        \match_addr_unencoded_raw[11][4] ), .A3(n55), .A4(n56), .Y(n52) );
  AND4X1_HVT U82 ( .A1(\match_addr_unencoded_raw[16][4] ), .A2(
        \match_addr_unencoded_raw[15][4] ), .A3(
        \match_addr_unencoded_raw[14][4] ), .A4(
        \match_addr_unencoded_raw[13][4] ), .Y(n56) );
  AND3X1_HVT U83 ( .A1(\match_addr_unencoded_raw[0][4] ), .A2(n175), .A3(
        \match_addr_unencoded_raw[10][4] ), .Y(n55) );
  AND4X1_HVT U91 ( .A1(\match_addr_unencoded_raw[16][3] ), .A2(
        \match_addr_unencoded_raw[15][3] ), .A3(
        \match_addr_unencoded_raw[14][3] ), .A4(
        \match_addr_unencoded_raw[13][3] ), .Y(n66) );
  AND3X1_HVT U92 ( .A1(\match_addr_unencoded_raw[0][3] ), .A2(n176), .A3(
        \match_addr_unencoded_raw[10][3] ), .Y(n65) );
  NAND4X0_HVT U96 ( .A1(\match_addr_unencoded_raw[5][3] ), .A2(
        \match_addr_unencoded_raw[4][3] ), .A3(
        \match_addr_unencoded_raw[3][3] ), .A4(
        \match_addr_unencoded_raw[31][3] ), .Y(n67) );
  NAND4X0_HVT U97 ( .A1(\match_addr_unencoded_raw[23][2] ), .A2(
        \match_addr_unencoded_raw[22][2] ), .A3(
        \match_addr_unencoded_raw[21][2] ), .A4(
        \match_addr_unencoded_raw[20][2] ), .Y(n74) );
  NAND4X0_HVT U98 ( .A1(\match_addr_unencoded_raw[1][2] ), .A2(
        \match_addr_unencoded_raw[19][2] ), .A3(
        \match_addr_unencoded_raw[18][2] ), .A4(
        \match_addr_unencoded_raw[17][2] ), .Y(n73) );
  NAND4X0_HVT U99 ( .A1(\match_addr_unencoded_raw[12][2] ), .A2(
        \match_addr_unencoded_raw[11][2] ), .A3(n75), .A4(n76), .Y(n72) );
  AND4X1_HVT U100 ( .A1(\match_addr_unencoded_raw[16][2] ), .A2(
        \match_addr_unencoded_raw[15][2] ), .A3(
        \match_addr_unencoded_raw[14][2] ), .A4(
        \match_addr_unencoded_raw[13][2] ), .Y(n76) );
  AND3X1_HVT U101 ( .A1(\match_addr_unencoded_raw[0][2] ), .A2(start), .A3(
        \match_addr_unencoded_raw[10][2] ), .Y(n75) );
  AND4X1_HVT U109 ( .A1(\match_addr_unencoded_raw[16][1] ), .A2(
        \match_addr_unencoded_raw[15][1] ), .A3(
        \match_addr_unencoded_raw[14][1] ), .A4(
        \match_addr_unencoded_raw[13][1] ), .Y(n86) );
  AND3X1_HVT U110 ( .A1(\match_addr_unencoded_raw[0][1] ), .A2(n175), .A3(
        \match_addr_unencoded_raw[10][1] ), .Y(n85) );
  NAND4X0_HVT U114 ( .A1(\match_addr_unencoded_raw[5][1] ), .A2(
        \match_addr_unencoded_raw[4][1] ), .A3(
        \match_addr_unencoded_raw[3][1] ), .A4(
        \match_addr_unencoded_raw[31][1] ), .Y(n87) );
  NAND4X0_HVT U115 ( .A1(\match_addr_unencoded_raw[23][15] ), .A2(
        \match_addr_unencoded_raw[22][15] ), .A3(
        \match_addr_unencoded_raw[21][15] ), .A4(
        \match_addr_unencoded_raw[20][15] ), .Y(n94) );
  NAND4X0_HVT U116 ( .A1(\match_addr_unencoded_raw[1][15] ), .A2(
        \match_addr_unencoded_raw[19][15] ), .A3(
        \match_addr_unencoded_raw[18][15] ), .A4(
        \match_addr_unencoded_raw[17][15] ), .Y(n93) );
  NAND4X0_HVT U117 ( .A1(\match_addr_unencoded_raw[12][15] ), .A2(
        \match_addr_unencoded_raw[11][15] ), .A3(n95), .A4(n96), .Y(n92) );
  AND4X1_HVT U118 ( .A1(\match_addr_unencoded_raw[16][15] ), .A2(
        \match_addr_unencoded_raw[15][15] ), .A3(
        \match_addr_unencoded_raw[14][15] ), .A4(
        \match_addr_unencoded_raw[13][15] ), .Y(n96) );
  AND3X1_HVT U119 ( .A1(\match_addr_unencoded_raw[0][15] ), .A2(n176), .A3(
        \match_addr_unencoded_raw[10][15] ), .Y(n95) );
  NAND4X0_HVT U124 ( .A1(\match_addr_unencoded_raw[23][14] ), .A2(
        \match_addr_unencoded_raw[22][14] ), .A3(
        \match_addr_unencoded_raw[21][14] ), .A4(
        \match_addr_unencoded_raw[20][14] ), .Y(n104) );
  NAND4X0_HVT U125 ( .A1(\match_addr_unencoded_raw[1][14] ), .A2(
        \match_addr_unencoded_raw[19][14] ), .A3(
        \match_addr_unencoded_raw[18][14] ), .A4(
        \match_addr_unencoded_raw[17][14] ), .Y(n103) );
  NAND4X0_HVT U126 ( .A1(\match_addr_unencoded_raw[12][14] ), .A2(
        \match_addr_unencoded_raw[11][14] ), .A3(n105), .A4(n106), .Y(n102) );
  AND4X1_HVT U127 ( .A1(\match_addr_unencoded_raw[16][14] ), .A2(
        \match_addr_unencoded_raw[15][14] ), .A3(
        \match_addr_unencoded_raw[14][14] ), .A4(
        \match_addr_unencoded_raw[13][14] ), .Y(n106) );
  AND3X1_HVT U128 ( .A1(\match_addr_unencoded_raw[0][14] ), .A2(n175), .A3(
        \match_addr_unencoded_raw[10][14] ), .Y(n105) );
  NAND4X0_HVT U133 ( .A1(\match_addr_unencoded_raw[23][13] ), .A2(
        \match_addr_unencoded_raw[22][13] ), .A3(
        \match_addr_unencoded_raw[21][13] ), .A4(
        \match_addr_unencoded_raw[20][13] ), .Y(n114) );
  NAND4X0_HVT U134 ( .A1(\match_addr_unencoded_raw[1][13] ), .A2(
        \match_addr_unencoded_raw[19][13] ), .A3(
        \match_addr_unencoded_raw[18][13] ), .A4(
        \match_addr_unencoded_raw[17][13] ), .Y(n113) );
  NAND4X0_HVT U135 ( .A1(\match_addr_unencoded_raw[12][13] ), .A2(
        \match_addr_unencoded_raw[11][13] ), .A3(n115), .A4(n116), .Y(n112) );
  AND4X1_HVT U136 ( .A1(\match_addr_unencoded_raw[16][13] ), .A2(
        \match_addr_unencoded_raw[15][13] ), .A3(
        \match_addr_unencoded_raw[14][13] ), .A4(
        \match_addr_unencoded_raw[13][13] ), .Y(n116) );
  AND3X1_HVT U137 ( .A1(\match_addr_unencoded_raw[0][13] ), .A2(n175), .A3(
        \match_addr_unencoded_raw[10][13] ), .Y(n115) );
  NAND4X0_HVT U142 ( .A1(\match_addr_unencoded_raw[23][12] ), .A2(
        \match_addr_unencoded_raw[22][12] ), .A3(
        \match_addr_unencoded_raw[21][12] ), .A4(
        \match_addr_unencoded_raw[20][12] ), .Y(n124) );
  NAND4X0_HVT U143 ( .A1(\match_addr_unencoded_raw[1][12] ), .A2(
        \match_addr_unencoded_raw[19][12] ), .A3(
        \match_addr_unencoded_raw[18][12] ), .A4(
        \match_addr_unencoded_raw[17][12] ), .Y(n123) );
  NAND4X0_HVT U144 ( .A1(\match_addr_unencoded_raw[12][12] ), .A2(
        \match_addr_unencoded_raw[11][12] ), .A3(n125), .A4(n126), .Y(n122) );
  AND4X1_HVT U145 ( .A1(\match_addr_unencoded_raw[16][12] ), .A2(
        \match_addr_unencoded_raw[15][12] ), .A3(
        \match_addr_unencoded_raw[14][12] ), .A4(
        \match_addr_unencoded_raw[13][12] ), .Y(n126) );
  AND3X1_HVT U146 ( .A1(\match_addr_unencoded_raw[0][12] ), .A2(n176), .A3(
        \match_addr_unencoded_raw[10][12] ), .Y(n125) );
  NAND4X0_HVT U151 ( .A1(\match_addr_unencoded_raw[23][11] ), .A2(
        \match_addr_unencoded_raw[22][11] ), .A3(
        \match_addr_unencoded_raw[21][11] ), .A4(
        \match_addr_unencoded_raw[20][11] ), .Y(n134) );
  NAND4X0_HVT U152 ( .A1(\match_addr_unencoded_raw[1][11] ), .A2(
        \match_addr_unencoded_raw[19][11] ), .A3(
        \match_addr_unencoded_raw[18][11] ), .A4(
        \match_addr_unencoded_raw[17][11] ), .Y(n133) );
  NAND4X0_HVT U153 ( .A1(\match_addr_unencoded_raw[12][11] ), .A2(
        \match_addr_unencoded_raw[11][11] ), .A3(n135), .A4(n136), .Y(n132) );
  AND4X1_HVT U154 ( .A1(\match_addr_unencoded_raw[16][11] ), .A2(
        \match_addr_unencoded_raw[15][11] ), .A3(
        \match_addr_unencoded_raw[14][11] ), .A4(
        \match_addr_unencoded_raw[13][11] ), .Y(n136) );
  AND3X1_HVT U155 ( .A1(\match_addr_unencoded_raw[0][11] ), .A2(n176), .A3(
        \match_addr_unencoded_raw[10][11] ), .Y(n135) );
  NAND4X0_HVT U160 ( .A1(\match_addr_unencoded_raw[23][10] ), .A2(
        \match_addr_unencoded_raw[22][10] ), .A3(
        \match_addr_unencoded_raw[21][10] ), .A4(
        \match_addr_unencoded_raw[20][10] ), .Y(n144) );
  NAND4X0_HVT U161 ( .A1(\match_addr_unencoded_raw[1][10] ), .A2(
        \match_addr_unencoded_raw[19][10] ), .A3(
        \match_addr_unencoded_raw[18][10] ), .A4(
        \match_addr_unencoded_raw[17][10] ), .Y(n143) );
  NAND4X0_HVT U162 ( .A1(\match_addr_unencoded_raw[12][10] ), .A2(
        \match_addr_unencoded_raw[11][10] ), .A3(n145), .A4(n146), .Y(n142) );
  AND4X1_HVT U163 ( .A1(\match_addr_unencoded_raw[16][10] ), .A2(
        \match_addr_unencoded_raw[15][10] ), .A3(
        \match_addr_unencoded_raw[14][10] ), .A4(
        \match_addr_unencoded_raw[13][10] ), .Y(n146) );
  AND3X1_HVT U164 ( .A1(\match_addr_unencoded_raw[0][10] ), .A2(n175), .A3(
        \match_addr_unencoded_raw[10][10] ), .Y(n145) );
  NAND4X0_HVT U169 ( .A1(\match_addr_unencoded_raw[23][0] ), .A2(
        \match_addr_unencoded_raw[22][0] ), .A3(
        \match_addr_unencoded_raw[21][0] ), .A4(
        \match_addr_unencoded_raw[20][0] ), .Y(n154) );
  NAND4X0_HVT U170 ( .A1(\match_addr_unencoded_raw[1][0] ), .A2(
        \match_addr_unencoded_raw[19][0] ), .A3(
        \match_addr_unencoded_raw[18][0] ), .A4(
        \match_addr_unencoded_raw[17][0] ), .Y(n153) );
  NAND4X0_HVT U171 ( .A1(\match_addr_unencoded_raw[12][0] ), .A2(
        \match_addr_unencoded_raw[11][0] ), .A3(n155), .A4(n156), .Y(n152) );
  AND4X1_HVT U172 ( .A1(\match_addr_unencoded_raw[16][0] ), .A2(
        \match_addr_unencoded_raw[15][0] ), .A3(
        \match_addr_unencoded_raw[14][0] ), .A4(
        \match_addr_unencoded_raw[13][0] ), .Y(n156) );
  AND3X1_HVT U173 ( .A1(\match_addr_unencoded_raw[0][0] ), .A2(n176), .A3(
        \match_addr_unencoded_raw[10][0] ), .Y(n155) );
  AND2X1_HVT U178 ( .A1(match_addr_w[3]), .A2(n176), .Y(N7) );
  AND2X1_HVT U179 ( .A1(match_addr_w[2]), .A2(start), .Y(N6) );
  AND2X1_HVT U180 ( .A1(match_addr_w[1]), .A2(n175), .Y(N5) );
  AND2X1_HVT U181 ( .A1(match_addr_w[0]), .A2(n176), .Y(N4) );
  OR2X1_HVT U182 ( .A1(n193), .A2(start), .Y(N3) );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_0 \slice[0].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n189), .a_addr({n185, n183, n179, n177}), .a_din(
        din[3:0]), .b_din(din[3:0]), .b_dout({
        \match_addr_unencoded_raw[0][15] , \match_addr_unencoded_raw[0][14] , 
        \match_addr_unencoded_raw[0][13] , \match_addr_unencoded_raw[0][12] , 
        \match_addr_unencoded_raw[0][11] , \match_addr_unencoded_raw[0][10] , 
        \match_addr_unencoded_raw[0][9] , \match_addr_unencoded_raw[0][8] , 
        \match_addr_unencoded_raw[0][7] , \match_addr_unencoded_raw[0][6] , 
        \match_addr_unencoded_raw[0][5] , \match_addr_unencoded_raw[0][4] , 
        \match_addr_unencoded_raw[0][3] , \match_addr_unencoded_raw[0][2] , 
        \match_addr_unencoded_raw[0][1] , \match_addr_unencoded_raw[0][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_31 \slice[1].ram_dp_inst  ( .clk(clk), .rst(
        n195), .write(n189), .a_addr({n187, n184, n181, write_addr[0]}), 
        .a_din(din[7:4]), .b_din(din[7:4]), .b_dout({
        \match_addr_unencoded_raw[1][15] , \match_addr_unencoded_raw[1][14] , 
        \match_addr_unencoded_raw[1][13] , \match_addr_unencoded_raw[1][12] , 
        \match_addr_unencoded_raw[1][11] , \match_addr_unencoded_raw[1][10] , 
        \match_addr_unencoded_raw[1][9] , \match_addr_unencoded_raw[1][8] , 
        \match_addr_unencoded_raw[1][7] , \match_addr_unencoded_raw[1][6] , 
        \match_addr_unencoded_raw[1][5] , \match_addr_unencoded_raw[1][4] , 
        \match_addr_unencoded_raw[1][3] , \match_addr_unencoded_raw[1][2] , 
        \match_addr_unencoded_raw[1][1] , \match_addr_unencoded_raw[1][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_30 \slice[2].ram_dp_inst  ( .clk(clk), .rst(
        n195), .write(n189), .a_addr({n187, write_addr[2], n181, n177}), 
        .a_din(din[11:8]), .b_din(din[11:8]), .b_dout({
        \match_addr_unencoded_raw[2][15] , \match_addr_unencoded_raw[2][14] , 
        \match_addr_unencoded_raw[2][13] , \match_addr_unencoded_raw[2][12] , 
        \match_addr_unencoded_raw[2][11] , \match_addr_unencoded_raw[2][10] , 
        \match_addr_unencoded_raw[2][9] , \match_addr_unencoded_raw[2][8] , 
        \match_addr_unencoded_raw[2][7] , \match_addr_unencoded_raw[2][6] , 
        \match_addr_unencoded_raw[2][5] , \match_addr_unencoded_raw[2][4] , 
        \match_addr_unencoded_raw[2][3] , \match_addr_unencoded_raw[2][2] , 
        \match_addr_unencoded_raw[2][1] , \match_addr_unencoded_raw[2][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_29 \slice[3].ram_dp_inst  ( .clk(clk), .rst(
        n195), .write(n191), .a_addr({n187, n183, n181, write_addr[0]}), 
        .a_din(din[15:12]), .b_din(din[15:12]), .b_dout({
        \match_addr_unencoded_raw[3][15] , \match_addr_unencoded_raw[3][14] , 
        \match_addr_unencoded_raw[3][13] , \match_addr_unencoded_raw[3][12] , 
        \match_addr_unencoded_raw[3][11] , \match_addr_unencoded_raw[3][10] , 
        \match_addr_unencoded_raw[3][9] , \match_addr_unencoded_raw[3][8] , 
        \match_addr_unencoded_raw[3][7] , \match_addr_unencoded_raw[3][6] , 
        \match_addr_unencoded_raw[3][5] , \match_addr_unencoded_raw[3][4] , 
        \match_addr_unencoded_raw[3][3] , \match_addr_unencoded_raw[3][2] , 
        \match_addr_unencoded_raw[3][1] , \match_addr_unencoded_raw[3][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_28 \slice[4].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n191), .a_addr({n187, n184, n181, n178}), .a_din(
        din[19:16]), .b_din(din[19:16]), .b_dout({
        \match_addr_unencoded_raw[4][15] , \match_addr_unencoded_raw[4][14] , 
        \match_addr_unencoded_raw[4][13] , \match_addr_unencoded_raw[4][12] , 
        \match_addr_unencoded_raw[4][11] , \match_addr_unencoded_raw[4][10] , 
        \match_addr_unencoded_raw[4][9] , \match_addr_unencoded_raw[4][8] , 
        \match_addr_unencoded_raw[4][7] , \match_addr_unencoded_raw[4][6] , 
        \match_addr_unencoded_raw[4][5] , \match_addr_unencoded_raw[4][4] , 
        \match_addr_unencoded_raw[4][3] , \match_addr_unencoded_raw[4][2] , 
        \match_addr_unencoded_raw[4][1] , \match_addr_unencoded_raw[4][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_27 \slice[5].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n191), .a_addr({n187, write_addr[2], n181, n177}), 
        .a_din(din[23:20]), .b_din(din[23:20]), .b_dout({
        \match_addr_unencoded_raw[5][15] , \match_addr_unencoded_raw[5][14] , 
        \match_addr_unencoded_raw[5][13] , \match_addr_unencoded_raw[5][12] , 
        \match_addr_unencoded_raw[5][11] , \match_addr_unencoded_raw[5][10] , 
        \match_addr_unencoded_raw[5][9] , \match_addr_unencoded_raw[5][8] , 
        \match_addr_unencoded_raw[5][7] , \match_addr_unencoded_raw[5][6] , 
        \match_addr_unencoded_raw[5][5] , \match_addr_unencoded_raw[5][4] , 
        \match_addr_unencoded_raw[5][3] , \match_addr_unencoded_raw[5][2] , 
        \match_addr_unencoded_raw[5][1] , \match_addr_unencoded_raw[5][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_26 \slice[6].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n191), .a_addr({n187, n183, n181, write_addr[0]}), 
        .a_din(din[27:24]), .b_din(din[27:24]), .b_dout({
        \match_addr_unencoded_raw[6][15] , \match_addr_unencoded_raw[6][14] , 
        \match_addr_unencoded_raw[6][13] , \match_addr_unencoded_raw[6][12] , 
        \match_addr_unencoded_raw[6][11] , \match_addr_unencoded_raw[6][10] , 
        \match_addr_unencoded_raw[6][9] , \match_addr_unencoded_raw[6][8] , 
        \match_addr_unencoded_raw[6][7] , \match_addr_unencoded_raw[6][6] , 
        \match_addr_unencoded_raw[6][5] , \match_addr_unencoded_raw[6][4] , 
        \match_addr_unencoded_raw[6][3] , \match_addr_unencoded_raw[6][2] , 
        \match_addr_unencoded_raw[6][1] , \match_addr_unencoded_raw[6][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_25 \slice[7].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n40), .a_addr({n187, n184, n181, n178}), .a_din(
        din[31:28]), .b_din(din[31:28]), .b_dout({
        \match_addr_unencoded_raw[7][15] , \match_addr_unencoded_raw[7][14] , 
        \match_addr_unencoded_raw[7][13] , \match_addr_unencoded_raw[7][12] , 
        \match_addr_unencoded_raw[7][11] , \match_addr_unencoded_raw[7][10] , 
        \match_addr_unencoded_raw[7][9] , \match_addr_unencoded_raw[7][8] , 
        \match_addr_unencoded_raw[7][7] , \match_addr_unencoded_raw[7][6] , 
        \match_addr_unencoded_raw[7][5] , \match_addr_unencoded_raw[7][4] , 
        \match_addr_unencoded_raw[7][3] , \match_addr_unencoded_raw[7][2] , 
        \match_addr_unencoded_raw[7][1] , \match_addr_unencoded_raw[7][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_24 \slice[8].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n39), .a_addr({n187, n172, n181, n167}), .a_din(
        din[35:32]), .b_din(din[35:32]), .b_dout({
        \match_addr_unencoded_raw[8][15] , \match_addr_unencoded_raw[8][14] , 
        \match_addr_unencoded_raw[8][13] , \match_addr_unencoded_raw[8][12] , 
        \match_addr_unencoded_raw[8][11] , \match_addr_unencoded_raw[8][10] , 
        \match_addr_unencoded_raw[8][9] , \match_addr_unencoded_raw[8][8] , 
        \match_addr_unencoded_raw[8][7] , \match_addr_unencoded_raw[8][6] , 
        \match_addr_unencoded_raw[8][5] , \match_addr_unencoded_raw[8][4] , 
        \match_addr_unencoded_raw[8][3] , \match_addr_unencoded_raw[8][2] , 
        \match_addr_unencoded_raw[8][1] , \match_addr_unencoded_raw[8][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_23 \slice[9].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n40), .a_addr({n186, n172, n180, n167}), .a_din(
        din[39:36]), .b_din(din[39:36]), .b_dout({
        \match_addr_unencoded_raw[9][15] , \match_addr_unencoded_raw[9][14] , 
        \match_addr_unencoded_raw[9][13] , \match_addr_unencoded_raw[9][12] , 
        \match_addr_unencoded_raw[9][11] , \match_addr_unencoded_raw[9][10] , 
        \match_addr_unencoded_raw[9][9] , \match_addr_unencoded_raw[9][8] , 
        \match_addr_unencoded_raw[9][7] , \match_addr_unencoded_raw[9][6] , 
        \match_addr_unencoded_raw[9][5] , \match_addr_unencoded_raw[9][4] , 
        \match_addr_unencoded_raw[9][3] , \match_addr_unencoded_raw[9][2] , 
        \match_addr_unencoded_raw[9][1] , \match_addr_unencoded_raw[9][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_22 \slice[10].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n190), .a_addr({n186, n172, n180, n167}), .a_din(
        din[43:40]), .b_din(din[43:40]), .b_dout({
        \match_addr_unencoded_raw[10][15] , \match_addr_unencoded_raw[10][14] , 
        \match_addr_unencoded_raw[10][13] , \match_addr_unencoded_raw[10][12] , 
        \match_addr_unencoded_raw[10][11] , \match_addr_unencoded_raw[10][10] , 
        \match_addr_unencoded_raw[10][9] , \match_addr_unencoded_raw[10][8] , 
        \match_addr_unencoded_raw[10][7] , \match_addr_unencoded_raw[10][6] , 
        \match_addr_unencoded_raw[10][5] , \match_addr_unencoded_raw[10][4] , 
        \match_addr_unencoded_raw[10][3] , \match_addr_unencoded_raw[10][2] , 
        \match_addr_unencoded_raw[10][1] , \match_addr_unencoded_raw[10][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_21 \slice[11].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n191), .a_addr({n186, n172, n180, n167}), .a_din(
        din[47:44]), .b_din(din[47:44]), .b_dout({
        \match_addr_unencoded_raw[11][15] , \match_addr_unencoded_raw[11][14] , 
        \match_addr_unencoded_raw[11][13] , \match_addr_unencoded_raw[11][12] , 
        \match_addr_unencoded_raw[11][11] , \match_addr_unencoded_raw[11][10] , 
        \match_addr_unencoded_raw[11][9] , \match_addr_unencoded_raw[11][8] , 
        \match_addr_unencoded_raw[11][7] , \match_addr_unencoded_raw[11][6] , 
        \match_addr_unencoded_raw[11][5] , \match_addr_unencoded_raw[11][4] , 
        \match_addr_unencoded_raw[11][3] , \match_addr_unencoded_raw[11][2] , 
        \match_addr_unencoded_raw[11][1] , \match_addr_unencoded_raw[11][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_20 \slice[12].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n40), .a_addr({n186, n172, n180, n167}), .a_din(
        din[51:48]), .b_din(din[51:48]), .b_dout({
        \match_addr_unencoded_raw[12][15] , \match_addr_unencoded_raw[12][14] , 
        \match_addr_unencoded_raw[12][13] , \match_addr_unencoded_raw[12][12] , 
        \match_addr_unencoded_raw[12][11] , \match_addr_unencoded_raw[12][10] , 
        \match_addr_unencoded_raw[12][9] , \match_addr_unencoded_raw[12][8] , 
        \match_addr_unencoded_raw[12][7] , \match_addr_unencoded_raw[12][6] , 
        \match_addr_unencoded_raw[12][5] , \match_addr_unencoded_raw[12][4] , 
        \match_addr_unencoded_raw[12][3] , \match_addr_unencoded_raw[12][2] , 
        \match_addr_unencoded_raw[12][1] , \match_addr_unencoded_raw[12][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_19 \slice[13].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n189), .a_addr({n186, n174, n180, n169}), .a_din(
        din[55:52]), .b_din(din[55:52]), .b_dout({
        \match_addr_unencoded_raw[13][15] , \match_addr_unencoded_raw[13][14] , 
        \match_addr_unencoded_raw[13][13] , \match_addr_unencoded_raw[13][12] , 
        \match_addr_unencoded_raw[13][11] , \match_addr_unencoded_raw[13][10] , 
        \match_addr_unencoded_raw[13][9] , \match_addr_unencoded_raw[13][8] , 
        \match_addr_unencoded_raw[13][7] , \match_addr_unencoded_raw[13][6] , 
        \match_addr_unencoded_raw[13][5] , \match_addr_unencoded_raw[13][4] , 
        \match_addr_unencoded_raw[13][3] , \match_addr_unencoded_raw[13][2] , 
        \match_addr_unencoded_raw[13][1] , \match_addr_unencoded_raw[13][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_18 \slice[14].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n190), .a_addr({n186, n173, n180, n168}), .a_din(
        din[59:56]), .b_din(din[59:56]), .b_dout({
        \match_addr_unencoded_raw[14][15] , \match_addr_unencoded_raw[14][14] , 
        \match_addr_unencoded_raw[14][13] , \match_addr_unencoded_raw[14][12] , 
        \match_addr_unencoded_raw[14][11] , \match_addr_unencoded_raw[14][10] , 
        \match_addr_unencoded_raw[14][9] , \match_addr_unencoded_raw[14][8] , 
        \match_addr_unencoded_raw[14][7] , \match_addr_unencoded_raw[14][6] , 
        \match_addr_unencoded_raw[14][5] , \match_addr_unencoded_raw[14][4] , 
        \match_addr_unencoded_raw[14][3] , \match_addr_unencoded_raw[14][2] , 
        \match_addr_unencoded_raw[14][1] , \match_addr_unencoded_raw[14][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_17 \slice[15].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n38), .a_addr({n186, n174, n180, n169}), .a_din(
        din[63:60]), .b_din(din[63:60]), .b_dout({
        \match_addr_unencoded_raw[15][15] , \match_addr_unencoded_raw[15][14] , 
        \match_addr_unencoded_raw[15][13] , \match_addr_unencoded_raw[15][12] , 
        \match_addr_unencoded_raw[15][11] , \match_addr_unencoded_raw[15][10] , 
        \match_addr_unencoded_raw[15][9] , \match_addr_unencoded_raw[15][8] , 
        \match_addr_unencoded_raw[15][7] , \match_addr_unencoded_raw[15][6] , 
        \match_addr_unencoded_raw[15][5] , \match_addr_unencoded_raw[15][4] , 
        \match_addr_unencoded_raw[15][3] , \match_addr_unencoded_raw[15][2] , 
        \match_addr_unencoded_raw[15][1] , \match_addr_unencoded_raw[15][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_16 \slice[16].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n189), .a_addr({n186, n173, n180, n168}), .a_din(
        din[67:64]), .b_din(din[67:64]), .b_dout({
        \match_addr_unencoded_raw[16][15] , \match_addr_unencoded_raw[16][14] , 
        \match_addr_unencoded_raw[16][13] , \match_addr_unencoded_raw[16][12] , 
        \match_addr_unencoded_raw[16][11] , \match_addr_unencoded_raw[16][10] , 
        \match_addr_unencoded_raw[16][9] , \match_addr_unencoded_raw[16][8] , 
        \match_addr_unencoded_raw[16][7] , \match_addr_unencoded_raw[16][6] , 
        \match_addr_unencoded_raw[16][5] , \match_addr_unencoded_raw[16][4] , 
        \match_addr_unencoded_raw[16][3] , \match_addr_unencoded_raw[16][2] , 
        \match_addr_unencoded_raw[16][1] , \match_addr_unencoded_raw[16][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_15 \slice[17].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n189), .a_addr({n186, n174, n180, n169}), .a_din(
        din[71:68]), .b_din(din[71:68]), .b_dout({
        \match_addr_unencoded_raw[17][15] , \match_addr_unencoded_raw[17][14] , 
        \match_addr_unencoded_raw[17][13] , \match_addr_unencoded_raw[17][12] , 
        \match_addr_unencoded_raw[17][11] , \match_addr_unencoded_raw[17][10] , 
        \match_addr_unencoded_raw[17][9] , \match_addr_unencoded_raw[17][8] , 
        \match_addr_unencoded_raw[17][7] , \match_addr_unencoded_raw[17][6] , 
        \match_addr_unencoded_raw[17][5] , \match_addr_unencoded_raw[17][4] , 
        \match_addr_unencoded_raw[17][3] , \match_addr_unencoded_raw[17][2] , 
        \match_addr_unencoded_raw[17][1] , \match_addr_unencoded_raw[17][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_14 \slice[18].ram_dp_inst  ( .clk(clk), .rst(
        n194), .write(n40), .a_addr({n186, n173, n180, n168}), .a_din(
        din[75:72]), .b_din(din[75:72]), .b_dout({
        \match_addr_unencoded_raw[18][15] , \match_addr_unencoded_raw[18][14] , 
        \match_addr_unencoded_raw[18][13] , \match_addr_unencoded_raw[18][12] , 
        \match_addr_unencoded_raw[18][11] , \match_addr_unencoded_raw[18][10] , 
        \match_addr_unencoded_raw[18][9] , \match_addr_unencoded_raw[18][8] , 
        \match_addr_unencoded_raw[18][7] , \match_addr_unencoded_raw[18][6] , 
        \match_addr_unencoded_raw[18][5] , \match_addr_unencoded_raw[18][4] , 
        \match_addr_unencoded_raw[18][3] , \match_addr_unencoded_raw[18][2] , 
        \match_addr_unencoded_raw[18][1] , \match_addr_unencoded_raw[18][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_13 \slice[19].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n40), .a_addr({n186, n174, n180, n169}), .a_din(
        din[79:76]), .b_din(din[79:76]), .b_dout({
        \match_addr_unencoded_raw[19][15] , \match_addr_unencoded_raw[19][14] , 
        \match_addr_unencoded_raw[19][13] , \match_addr_unencoded_raw[19][12] , 
        \match_addr_unencoded_raw[19][11] , \match_addr_unencoded_raw[19][10] , 
        \match_addr_unencoded_raw[19][9] , \match_addr_unencoded_raw[19][8] , 
        \match_addr_unencoded_raw[19][7] , \match_addr_unencoded_raw[19][6] , 
        \match_addr_unencoded_raw[19][5] , \match_addr_unencoded_raw[19][4] , 
        \match_addr_unencoded_raw[19][3] , \match_addr_unencoded_raw[19][2] , 
        \match_addr_unencoded_raw[19][1] , \match_addr_unencoded_raw[19][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_12 \slice[20].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n39), .a_addr({n186, n173, n180, n168}), .a_din(
        din[83:80]), .b_din(din[83:80]), .b_dout({
        \match_addr_unencoded_raw[20][15] , \match_addr_unencoded_raw[20][14] , 
        \match_addr_unencoded_raw[20][13] , \match_addr_unencoded_raw[20][12] , 
        \match_addr_unencoded_raw[20][11] , \match_addr_unencoded_raw[20][10] , 
        \match_addr_unencoded_raw[20][9] , \match_addr_unencoded_raw[20][8] , 
        \match_addr_unencoded_raw[20][7] , \match_addr_unencoded_raw[20][6] , 
        \match_addr_unencoded_raw[20][5] , \match_addr_unencoded_raw[20][4] , 
        \match_addr_unencoded_raw[20][3] , \match_addr_unencoded_raw[20][2] , 
        \match_addr_unencoded_raw[20][1] , \match_addr_unencoded_raw[20][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_11 \slice[21].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n38), .a_addr({n185, n170, n179, n165}), .a_din(
        din[87:84]), .b_din(din[87:84]), .b_dout({
        \match_addr_unencoded_raw[21][15] , \match_addr_unencoded_raw[21][14] , 
        \match_addr_unencoded_raw[21][13] , \match_addr_unencoded_raw[21][12] , 
        \match_addr_unencoded_raw[21][11] , \match_addr_unencoded_raw[21][10] , 
        \match_addr_unencoded_raw[21][9] , \match_addr_unencoded_raw[21][8] , 
        \match_addr_unencoded_raw[21][7] , \match_addr_unencoded_raw[21][6] , 
        \match_addr_unencoded_raw[21][5] , \match_addr_unencoded_raw[21][4] , 
        \match_addr_unencoded_raw[21][3] , \match_addr_unencoded_raw[21][2] , 
        \match_addr_unencoded_raw[21][1] , \match_addr_unencoded_raw[21][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_10 \slice[22].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n39), .a_addr({n185, n170, n179, n165}), .a_din(
        din[91:88]), .b_din(din[91:88]), .b_dout({
        \match_addr_unencoded_raw[22][15] , \match_addr_unencoded_raw[22][14] , 
        \match_addr_unencoded_raw[22][13] , \match_addr_unencoded_raw[22][12] , 
        \match_addr_unencoded_raw[22][11] , \match_addr_unencoded_raw[22][10] , 
        \match_addr_unencoded_raw[22][9] , \match_addr_unencoded_raw[22][8] , 
        \match_addr_unencoded_raw[22][7] , \match_addr_unencoded_raw[22][6] , 
        \match_addr_unencoded_raw[22][5] , \match_addr_unencoded_raw[22][4] , 
        \match_addr_unencoded_raw[22][3] , \match_addr_unencoded_raw[22][2] , 
        \match_addr_unencoded_raw[22][1] , \match_addr_unencoded_raw[22][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_9 \slice[23].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n190), .a_addr({n185, n170, n179, n165}), .a_din(
        din[95:92]), .b_din(din[95:92]), .b_dout({
        \match_addr_unencoded_raw[23][15] , \match_addr_unencoded_raw[23][14] , 
        \match_addr_unencoded_raw[23][13] , \match_addr_unencoded_raw[23][12] , 
        \match_addr_unencoded_raw[23][11] , \match_addr_unencoded_raw[23][10] , 
        \match_addr_unencoded_raw[23][9] , \match_addr_unencoded_raw[23][8] , 
        \match_addr_unencoded_raw[23][7] , \match_addr_unencoded_raw[23][6] , 
        \match_addr_unencoded_raw[23][5] , \match_addr_unencoded_raw[23][4] , 
        \match_addr_unencoded_raw[23][3] , \match_addr_unencoded_raw[23][2] , 
        \match_addr_unencoded_raw[23][1] , \match_addr_unencoded_raw[23][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_8 \slice[24].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n190), .a_addr({n185, n170, n179, n165}), .a_din(
        din[99:96]), .b_din(din[99:96]), .b_dout({
        \match_addr_unencoded_raw[24][15] , \match_addr_unencoded_raw[24][14] , 
        \match_addr_unencoded_raw[24][13] , \match_addr_unencoded_raw[24][12] , 
        \match_addr_unencoded_raw[24][11] , \match_addr_unencoded_raw[24][10] , 
        \match_addr_unencoded_raw[24][9] , \match_addr_unencoded_raw[24][8] , 
        \match_addr_unencoded_raw[24][7] , \match_addr_unencoded_raw[24][6] , 
        \match_addr_unencoded_raw[24][5] , \match_addr_unencoded_raw[24][4] , 
        \match_addr_unencoded_raw[24][3] , \match_addr_unencoded_raw[24][2] , 
        \match_addr_unencoded_raw[24][1] , \match_addr_unencoded_raw[24][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_7 \slice[25].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n39), .a_addr({n185, n171, n179, n166}), .a_din(
        din[103:100]), .b_din(din[103:100]), .b_dout({
        \match_addr_unencoded_raw[25][15] , \match_addr_unencoded_raw[25][14] , 
        \match_addr_unencoded_raw[25][13] , \match_addr_unencoded_raw[25][12] , 
        \match_addr_unencoded_raw[25][11] , \match_addr_unencoded_raw[25][10] , 
        \match_addr_unencoded_raw[25][9] , \match_addr_unencoded_raw[25][8] , 
        \match_addr_unencoded_raw[25][7] , \match_addr_unencoded_raw[25][6] , 
        \match_addr_unencoded_raw[25][5] , \match_addr_unencoded_raw[25][4] , 
        \match_addr_unencoded_raw[25][3] , \match_addr_unencoded_raw[25][2] , 
        \match_addr_unencoded_raw[25][1] , \match_addr_unencoded_raw[25][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_6 \slice[26].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n190), .a_addr({n185, write_addr[2], n179, n178}), 
        .a_din(din[107:104]), .b_din(din[107:104]), .b_dout({
        \match_addr_unencoded_raw[26][15] , \match_addr_unencoded_raw[26][14] , 
        \match_addr_unencoded_raw[26][13] , \match_addr_unencoded_raw[26][12] , 
        \match_addr_unencoded_raw[26][11] , \match_addr_unencoded_raw[26][10] , 
        \match_addr_unencoded_raw[26][9] , \match_addr_unencoded_raw[26][8] , 
        \match_addr_unencoded_raw[26][7] , \match_addr_unencoded_raw[26][6] , 
        \match_addr_unencoded_raw[26][5] , \match_addr_unencoded_raw[26][4] , 
        \match_addr_unencoded_raw[26][3] , \match_addr_unencoded_raw[26][2] , 
        \match_addr_unencoded_raw[26][1] , \match_addr_unencoded_raw[26][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_5 \slice[27].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n38), .a_addr({n185, n171, n179, n166}), .a_din(
        din[111:108]), .b_din(din[111:108]), .b_dout({
        \match_addr_unencoded_raw[27][15] , \match_addr_unencoded_raw[27][14] , 
        \match_addr_unencoded_raw[27][13] , \match_addr_unencoded_raw[27][12] , 
        \match_addr_unencoded_raw[27][11] , \match_addr_unencoded_raw[27][10] , 
        \match_addr_unencoded_raw[27][9] , \match_addr_unencoded_raw[27][8] , 
        \match_addr_unencoded_raw[27][7] , \match_addr_unencoded_raw[27][6] , 
        \match_addr_unencoded_raw[27][5] , \match_addr_unencoded_raw[27][4] , 
        \match_addr_unencoded_raw[27][3] , \match_addr_unencoded_raw[27][2] , 
        \match_addr_unencoded_raw[27][1] , \match_addr_unencoded_raw[27][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_4 \slice[28].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n39), .a_addr({n185, n183, n179, n177}), .a_din(
        din[115:112]), .b_din(din[115:112]), .b_dout({
        \match_addr_unencoded_raw[28][15] , \match_addr_unencoded_raw[28][14] , 
        \match_addr_unencoded_raw[28][13] , \match_addr_unencoded_raw[28][12] , 
        \match_addr_unencoded_raw[28][11] , \match_addr_unencoded_raw[28][10] , 
        \match_addr_unencoded_raw[28][9] , \match_addr_unencoded_raw[28][8] , 
        \match_addr_unencoded_raw[28][7] , \match_addr_unencoded_raw[28][6] , 
        \match_addr_unencoded_raw[28][5] , \match_addr_unencoded_raw[28][4] , 
        \match_addr_unencoded_raw[28][3] , \match_addr_unencoded_raw[28][2] , 
        \match_addr_unencoded_raw[28][1] , \match_addr_unencoded_raw[28][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_3 \slice[29].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n38), .a_addr({n185, n171, n179, n166}), .a_din(
        din[119:116]), .b_din(din[119:116]), .b_dout({
        \match_addr_unencoded_raw[29][15] , \match_addr_unencoded_raw[29][14] , 
        \match_addr_unencoded_raw[29][13] , \match_addr_unencoded_raw[29][12] , 
        \match_addr_unencoded_raw[29][11] , \match_addr_unencoded_raw[29][10] , 
        \match_addr_unencoded_raw[29][9] , \match_addr_unencoded_raw[29][8] , 
        \match_addr_unencoded_raw[29][7] , \match_addr_unencoded_raw[29][6] , 
        \match_addr_unencoded_raw[29][5] , \match_addr_unencoded_raw[29][4] , 
        \match_addr_unencoded_raw[29][3] , \match_addr_unencoded_raw[29][2] , 
        \match_addr_unencoded_raw[29][1] , \match_addr_unencoded_raw[29][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_2 \slice[30].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n39), .a_addr({n185, n184, n179, n178}), .a_din(
        din[123:120]), .b_din(din[123:120]), .b_dout({
        \match_addr_unencoded_raw[30][15] , \match_addr_unencoded_raw[30][14] , 
        \match_addr_unencoded_raw[30][13] , \match_addr_unencoded_raw[30][12] , 
        \match_addr_unencoded_raw[30][11] , \match_addr_unencoded_raw[30][10] , 
        \match_addr_unencoded_raw[30][9] , \match_addr_unencoded_raw[30][8] , 
        \match_addr_unencoded_raw[30][7] , \match_addr_unencoded_raw[30][6] , 
        \match_addr_unencoded_raw[30][5] , \match_addr_unencoded_raw[30][4] , 
        \match_addr_unencoded_raw[30][3] , \match_addr_unencoded_raw[30][2] , 
        \match_addr_unencoded_raw[30][1] , \match_addr_unencoded_raw[30][0] })
         );
  ram_dp_DATA_WIDTH4_ADDR_WIDTH4_1 \slice[31].ram_dp_inst  ( .clk(clk), .rst(
        n193), .write(n38), .a_addr({n185, n171, n179, n166}), .a_din(
        din[127:124]), .b_din(din[127:124]), .b_dout({
        \match_addr_unencoded_raw[31][15] , \match_addr_unencoded_raw[31][14] , 
        \match_addr_unencoded_raw[31][13] , \match_addr_unencoded_raw[31][12] , 
        \match_addr_unencoded_raw[31][11] , \match_addr_unencoded_raw[31][10] , 
        \match_addr_unencoded_raw[31][9] , \match_addr_unencoded_raw[31][8] , 
        \match_addr_unencoded_raw[31][7] , \match_addr_unencoded_raw[31][6] , 
        \match_addr_unencoded_raw[31][5] , \match_addr_unencoded_raw[31][4] , 
        \match_addr_unencoded_raw[31][3] , \match_addr_unencoded_raw[31][2] , 
        \match_addr_unencoded_raw[31][1] , \match_addr_unencoded_raw[31][0] })
         );
  encoder_WIDTH16 encoder_inst1 ( .clk(clk), .input_unencoded(
        match_addr_unencoded), .output_valid(match), .output_encoded(
        match_addr_w) );
  INVX0_HVT U3 ( .A(write_enable), .Y(n192) );
  INVX1_HVT U5 ( .A(n41), .Y(n39) );
  NOR4X1_HVT U6 ( .A1(n67), .A2(n42), .A3(n43), .A4(n44), .Y(n7) );
  AND4X1_HVT U7 ( .A1(\match_addr_unencoded_raw[5][2] ), .A2(
        \match_addr_unencoded_raw[4][2] ), .A3(
        \match_addr_unencoded_raw[3][2] ), .A4(
        \match_addr_unencoded_raw[31][2] ), .Y(n8) );
  NOR4X1_HVT U9 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .Y(n9) );
  NOR4X1_HVT U10 ( .A1(n87), .A2(n57), .A3(n58), .A4(n59), .Y(n10) );
  AND4X1_HVT U11 ( .A1(\match_addr_unencoded_raw[5][4] ), .A2(
        \match_addr_unencoded_raw[4][4] ), .A3(
        \match_addr_unencoded_raw[3][4] ), .A4(
        \match_addr_unencoded_raw[31][4] ), .Y(n17) );
  AND4X1_HVT U13 ( .A1(\match_addr_unencoded_raw[5][13] ), .A2(
        \match_addr_unencoded_raw[4][13] ), .A3(
        \match_addr_unencoded_raw[3][13] ), .A4(
        \match_addr_unencoded_raw[31][13] ), .Y(n18) );
  AND4X1_HVT U14 ( .A1(\match_addr_unencoded_raw[5][15] ), .A2(
        \match_addr_unencoded_raw[4][15] ), .A3(
        \match_addr_unencoded_raw[3][15] ), .A4(
        \match_addr_unencoded_raw[31][15] ), .Y(n19) );
  NOR4X1_HVT U15 ( .A1(n27), .A2(n60), .A3(n61), .A4(n62), .Y(n20) );
  AND4X1_HVT U17 ( .A1(\match_addr_unencoded_raw[5][6] ), .A2(
        \match_addr_unencoded_raw[4][6] ), .A3(
        \match_addr_unencoded_raw[3][6] ), .A4(
        \match_addr_unencoded_raw[31][6] ), .Y(n21) );
  AND4X1_HVT U18 ( .A1(\match_addr_unencoded_raw[5][12] ), .A2(
        \match_addr_unencoded_raw[4][12] ), .A3(
        \match_addr_unencoded_raw[3][12] ), .A4(
        \match_addr_unencoded_raw[31][12] ), .Y(n22) );
  AND4X1_HVT U19 ( .A1(\match_addr_unencoded_raw[5][14] ), .A2(
        \match_addr_unencoded_raw[4][14] ), .A3(
        \match_addr_unencoded_raw[3][14] ), .A4(
        \match_addr_unencoded_raw[31][14] ), .Y(n23) );
  AND4X1_HVT U21 ( .A1(\match_addr_unencoded_raw[6][9] ), .A2(
        \match_addr_unencoded_raw[5][9] ), .A3(
        \match_addr_unencoded_raw[4][9] ), .A4(
        \match_addr_unencoded_raw[3][9] ), .Y(n24) );
  AND4X1_HVT U23 ( .A1(\match_addr_unencoded_raw[5][11] ), .A2(
        \match_addr_unencoded_raw[4][11] ), .A3(
        \match_addr_unencoded_raw[3][11] ), .A4(
        \match_addr_unencoded_raw[31][11] ), .Y(n28) );
  AND4X1_HVT U25 ( .A1(\match_addr_unencoded_raw[5][8] ), .A2(
        \match_addr_unencoded_raw[4][8] ), .A3(
        \match_addr_unencoded_raw[3][8] ), .A4(
        \match_addr_unencoded_raw[31][8] ), .Y(n29) );
  AND4X1_HVT U27 ( .A1(\match_addr_unencoded_raw[5][10] ), .A2(
        \match_addr_unencoded_raw[4][10] ), .A3(
        \match_addr_unencoded_raw[3][10] ), .A4(
        \match_addr_unencoded_raw[31][10] ), .Y(n30) );
  AND4X1_HVT U29 ( .A1(\match_addr_unencoded_raw[5][0] ), .A2(
        \match_addr_unencoded_raw[4][0] ), .A3(
        \match_addr_unencoded_raw[3][0] ), .A4(
        \match_addr_unencoded_raw[31][0] ), .Y(n37) );
  INVX0_HVT U31 ( .A(n41), .Y(n38) );
  INVX0_HVT U33 ( .A(n41), .Y(n190) );
  IBUFFX2_HVT U39 ( .A(write_enable), .Y(n41) );
  INVX1_HVT U40 ( .A(n192), .Y(n40) );
  IBUFFX2_HVT U41 ( .A(n192), .Y(n191) );
  NAND4X0_HVT U42 ( .A1(\match_addr_unencoded_raw[9][3] ), .A2(
        \match_addr_unencoded_raw[8][3] ), .A3(
        \match_addr_unencoded_raw[7][3] ), .A4(
        \match_addr_unencoded_raw[6][3] ), .Y(n42) );
  NAND4X0_HVT U48 ( .A1(\match_addr_unencoded_raw[27][3] ), .A2(
        \match_addr_unencoded_raw[26][3] ), .A3(
        \match_addr_unencoded_raw[25][3] ), .A4(
        \match_addr_unencoded_raw[24][3] ), .Y(n43) );
  NAND4X0_HVT U49 ( .A1(\match_addr_unencoded_raw[30][3] ), .A2(
        \match_addr_unencoded_raw[2][3] ), .A3(
        \match_addr_unencoded_raw[29][3] ), .A4(
        \match_addr_unencoded_raw[28][3] ), .Y(n44) );
  NAND4X0_HVT U50 ( .A1(\match_addr_unencoded_raw[9][5] ), .A2(
        \match_addr_unencoded_raw[8][5] ), .A3(
        \match_addr_unencoded_raw[7][5] ), .A4(
        \match_addr_unencoded_raw[6][5] ), .Y(n48) );
  NAND4X0_HVT U51 ( .A1(\match_addr_unencoded_raw[27][5] ), .A2(
        \match_addr_unencoded_raw[26][5] ), .A3(
        \match_addr_unencoded_raw[25][5] ), .A4(
        \match_addr_unencoded_raw[24][5] ), .Y(n49) );
  NAND4X0_HVT U52 ( .A1(\match_addr_unencoded_raw[30][5] ), .A2(
        \match_addr_unencoded_raw[2][5] ), .A3(
        \match_addr_unencoded_raw[29][5] ), .A4(
        \match_addr_unencoded_raw[28][5] ), .Y(n50) );
  NAND4X0_HVT U53 ( .A1(\match_addr_unencoded_raw[9][1] ), .A2(
        \match_addr_unencoded_raw[8][1] ), .A3(
        \match_addr_unencoded_raw[7][1] ), .A4(
        \match_addr_unencoded_raw[6][1] ), .Y(n57) );
  NAND4X0_HVT U54 ( .A1(\match_addr_unencoded_raw[27][1] ), .A2(
        \match_addr_unencoded_raw[26][1] ), .A3(
        \match_addr_unencoded_raw[25][1] ), .A4(
        \match_addr_unencoded_raw[24][1] ), .Y(n58) );
  NAND4X0_HVT U57 ( .A1(\match_addr_unencoded_raw[30][1] ), .A2(
        \match_addr_unencoded_raw[2][1] ), .A3(
        \match_addr_unencoded_raw[29][1] ), .A4(
        \match_addr_unencoded_raw[28][1] ), .Y(n59) );
  NAND4X0_HVT U58 ( .A1(\match_addr_unencoded_raw[9][7] ), .A2(
        \match_addr_unencoded_raw[8][7] ), .A3(
        \match_addr_unencoded_raw[7][7] ), .A4(
        \match_addr_unencoded_raw[6][7] ), .Y(n60) );
  NAND4X0_HVT U59 ( .A1(\match_addr_unencoded_raw[27][7] ), .A2(
        \match_addr_unencoded_raw[26][7] ), .A3(
        \match_addr_unencoded_raw[25][7] ), .A4(
        \match_addr_unencoded_raw[24][7] ), .Y(n61) );
  NAND4X0_HVT U66 ( .A1(\match_addr_unencoded_raw[30][7] ), .A2(
        \match_addr_unencoded_raw[2][7] ), .A3(
        \match_addr_unencoded_raw[29][7] ), .A4(
        \match_addr_unencoded_raw[28][7] ), .Y(n62) );
  INVX1_HVT U67 ( .A(n192), .Y(n189) );
  INVX1_HVT U68 ( .A(n196), .Y(n194) );
  INVX1_HVT U69 ( .A(n196), .Y(n193) );
  INVX1_HVT U70 ( .A(n196), .Y(n195) );
  INVX1_HVT U71 ( .A(rst), .Y(n196) );
  INVX1_HVT U72 ( .A(n188), .Y(n186) );
  INVX1_HVT U75 ( .A(n188), .Y(n185) );
  INVX1_HVT U76 ( .A(n188), .Y(n187) );
  NBUFFX2_HVT U77 ( .A(n178), .Y(n167) );
  NBUFFX2_HVT U84 ( .A(n178), .Y(n169) );
  NBUFFX2_HVT U85 ( .A(n178), .Y(n168) );
  NBUFFX2_HVT U86 ( .A(n177), .Y(n165) );
  NBUFFX2_HVT U87 ( .A(n177), .Y(n166) );
  NBUFFX2_HVT U88 ( .A(n184), .Y(n172) );
  NBUFFX2_HVT U89 ( .A(n184), .Y(n174) );
  NBUFFX2_HVT U90 ( .A(n184), .Y(n173) );
  NBUFFX2_HVT U93 ( .A(n183), .Y(n170) );
  NBUFFX2_HVT U94 ( .A(n183), .Y(n171) );
  INVX1_HVT U95 ( .A(n182), .Y(n180) );
  INVX1_HVT U102 ( .A(n182), .Y(n179) );
  INVX1_HVT U103 ( .A(n182), .Y(n181) );
  AND4X1_HVT U104 ( .A1(n7), .A2(n63), .A3(n64), .A4(n68), .Y(
        match_addr_unencoded[3]) );
  AND4X1_HVT U105 ( .A1(\match_addr_unencoded_raw[12][3] ), .A2(
        \match_addr_unencoded_raw[11][3] ), .A3(n65), .A4(n66), .Y(n63) );
  AND4X1_HVT U106 ( .A1(\match_addr_unencoded_raw[1][3] ), .A2(
        \match_addr_unencoded_raw[19][3] ), .A3(
        \match_addr_unencoded_raw[18][3] ), .A4(
        \match_addr_unencoded_raw[17][3] ), .Y(n64) );
  AND4X1_HVT U107 ( .A1(\match_addr_unencoded_raw[23][3] ), .A2(
        \match_addr_unencoded_raw[22][3] ), .A3(
        \match_addr_unencoded_raw[21][3] ), .A4(
        \match_addr_unencoded_raw[20][3] ), .Y(n68) );
  AND4X1_HVT U108 ( .A1(n9), .A2(n69), .A3(n70), .A4(n77), .Y(
        match_addr_unencoded[5]) );
  AND4X1_HVT U111 ( .A1(\match_addr_unencoded_raw[12][5] ), .A2(
        \match_addr_unencoded_raw[11][5] ), .A3(n45), .A4(n46), .Y(n69) );
  AND4X1_HVT U112 ( .A1(\match_addr_unencoded_raw[1][5] ), .A2(
        \match_addr_unencoded_raw[19][5] ), .A3(
        \match_addr_unencoded_raw[18][5] ), .A4(
        \match_addr_unencoded_raw[17][5] ), .Y(n70) );
  AND4X1_HVT U113 ( .A1(\match_addr_unencoded_raw[23][5] ), .A2(
        \match_addr_unencoded_raw[22][5] ), .A3(
        \match_addr_unencoded_raw[21][5] ), .A4(
        \match_addr_unencoded_raw[20][5] ), .Y(n77) );
  NAND4X0_HVT U120 ( .A1(n8), .A2(n78), .A3(n79), .A4(n80), .Y(n71) );
  AND4X1_HVT U121 ( .A1(\match_addr_unencoded_raw[9][2] ), .A2(
        \match_addr_unencoded_raw[8][2] ), .A3(
        \match_addr_unencoded_raw[7][2] ), .A4(
        \match_addr_unencoded_raw[6][2] ), .Y(n78) );
  AND4X1_HVT U122 ( .A1(\match_addr_unencoded_raw[27][2] ), .A2(
        \match_addr_unencoded_raw[26][2] ), .A3(
        \match_addr_unencoded_raw[25][2] ), .A4(
        \match_addr_unencoded_raw[24][2] ), .Y(n79) );
  AND4X1_HVT U123 ( .A1(\match_addr_unencoded_raw[30][2] ), .A2(
        \match_addr_unencoded_raw[2][2] ), .A3(
        \match_addr_unencoded_raw[29][2] ), .A4(
        \match_addr_unencoded_raw[28][2] ), .Y(n80) );
  AND4X1_HVT U129 ( .A1(n10), .A2(n81), .A3(n82), .A4(n83), .Y(
        match_addr_unencoded[1]) );
  AND4X1_HVT U130 ( .A1(\match_addr_unencoded_raw[12][1] ), .A2(
        \match_addr_unencoded_raw[11][1] ), .A3(n85), .A4(n86), .Y(n81) );
  AND4X1_HVT U131 ( .A1(\match_addr_unencoded_raw[1][1] ), .A2(
        \match_addr_unencoded_raw[19][1] ), .A3(
        \match_addr_unencoded_raw[18][1] ), .A4(
        \match_addr_unencoded_raw[17][1] ), .Y(n82) );
  AND4X1_HVT U132 ( .A1(\match_addr_unencoded_raw[23][1] ), .A2(
        \match_addr_unencoded_raw[22][1] ), .A3(
        \match_addr_unencoded_raw[21][1] ), .A4(
        \match_addr_unencoded_raw[20][1] ), .Y(n83) );
  AND4X1_HVT U138 ( .A1(n20), .A2(n84), .A3(n88), .A4(n89), .Y(
        match_addr_unencoded[7]) );
  AND4X1_HVT U139 ( .A1(\match_addr_unencoded_raw[12][7] ), .A2(
        \match_addr_unencoded_raw[11][7] ), .A3(n25), .A4(n26), .Y(n84) );
  AND4X1_HVT U140 ( .A1(\match_addr_unencoded_raw[1][7] ), .A2(
        \match_addr_unencoded_raw[19][7] ), .A3(
        \match_addr_unencoded_raw[18][7] ), .A4(
        \match_addr_unencoded_raw[17][7] ), .Y(n88) );
  AND4X1_HVT U141 ( .A1(\match_addr_unencoded_raw[23][7] ), .A2(
        \match_addr_unencoded_raw[22][7] ), .A3(
        \match_addr_unencoded_raw[21][7] ), .A4(
        \match_addr_unencoded_raw[20][7] ), .Y(n89) );
  NAND4X0_HVT U147 ( .A1(n17), .A2(n90), .A3(n97), .A4(n98), .Y(n51) );
  AND4X1_HVT U148 ( .A1(\match_addr_unencoded_raw[9][4] ), .A2(
        \match_addr_unencoded_raw[8][4] ), .A3(
        \match_addr_unencoded_raw[7][4] ), .A4(
        \match_addr_unencoded_raw[6][4] ), .Y(n90) );
  AND4X1_HVT U149 ( .A1(\match_addr_unencoded_raw[27][4] ), .A2(
        \match_addr_unencoded_raw[26][4] ), .A3(
        \match_addr_unencoded_raw[25][4] ), .A4(
        \match_addr_unencoded_raw[24][4] ), .Y(n97) );
  AND4X1_HVT U150 ( .A1(\match_addr_unencoded_raw[30][4] ), .A2(
        \match_addr_unencoded_raw[2][4] ), .A3(
        \match_addr_unencoded_raw[29][4] ), .A4(
        \match_addr_unencoded_raw[28][4] ), .Y(n98) );
  NAND4X0_HVT U156 ( .A1(n18), .A2(n99), .A3(n100), .A4(n107), .Y(n111) );
  AND4X1_HVT U157 ( .A1(\match_addr_unencoded_raw[9][13] ), .A2(
        \match_addr_unencoded_raw[8][13] ), .A3(
        \match_addr_unencoded_raw[7][13] ), .A4(
        \match_addr_unencoded_raw[6][13] ), .Y(n99) );
  AND4X1_HVT U158 ( .A1(\match_addr_unencoded_raw[27][13] ), .A2(
        \match_addr_unencoded_raw[26][13] ), .A3(
        \match_addr_unencoded_raw[25][13] ), .A4(
        \match_addr_unencoded_raw[24][13] ), .Y(n100) );
  AND4X1_HVT U159 ( .A1(\match_addr_unencoded_raw[30][13] ), .A2(
        \match_addr_unencoded_raw[2][13] ), .A3(
        \match_addr_unencoded_raw[29][13] ), .A4(
        \match_addr_unencoded_raw[28][13] ), .Y(n107) );
  NAND4X0_HVT U165 ( .A1(n19), .A2(n108), .A3(n109), .A4(n110), .Y(n91) );
  AND4X1_HVT U166 ( .A1(\match_addr_unencoded_raw[9][15] ), .A2(
        \match_addr_unencoded_raw[8][15] ), .A3(
        \match_addr_unencoded_raw[7][15] ), .A4(
        \match_addr_unencoded_raw[6][15] ), .Y(n108) );
  AND4X1_HVT U167 ( .A1(\match_addr_unencoded_raw[27][15] ), .A2(
        \match_addr_unencoded_raw[26][15] ), .A3(
        \match_addr_unencoded_raw[25][15] ), .A4(
        \match_addr_unencoded_raw[24][15] ), .Y(n109) );
  AND4X1_HVT U168 ( .A1(\match_addr_unencoded_raw[30][15] ), .A2(
        \match_addr_unencoded_raw[2][15] ), .A3(
        \match_addr_unencoded_raw[29][15] ), .A4(
        \match_addr_unencoded_raw[28][15] ), .Y(n110) );
  NAND4X0_HVT U174 ( .A1(n21), .A2(n117), .A3(n118), .A4(n119), .Y(n31) );
  AND4X1_HVT U175 ( .A1(\match_addr_unencoded_raw[9][6] ), .A2(
        \match_addr_unencoded_raw[8][6] ), .A3(
        \match_addr_unencoded_raw[7][6] ), .A4(
        \match_addr_unencoded_raw[6][6] ), .Y(n117) );
  AND4X1_HVT U176 ( .A1(\match_addr_unencoded_raw[27][6] ), .A2(
        \match_addr_unencoded_raw[26][6] ), .A3(
        \match_addr_unencoded_raw[25][6] ), .A4(
        \match_addr_unencoded_raw[24][6] ), .Y(n118) );
  AND4X1_HVT U177 ( .A1(\match_addr_unencoded_raw[30][6] ), .A2(
        \match_addr_unencoded_raw[2][6] ), .A3(
        \match_addr_unencoded_raw[29][6] ), .A4(
        \match_addr_unencoded_raw[28][6] ), .Y(n119) );
  NAND4X0_HVT U183 ( .A1(n22), .A2(n120), .A3(n127), .A4(n128), .Y(n121) );
  AND4X1_HVT U184 ( .A1(\match_addr_unencoded_raw[9][12] ), .A2(
        \match_addr_unencoded_raw[8][12] ), .A3(
        \match_addr_unencoded_raw[7][12] ), .A4(
        \match_addr_unencoded_raw[6][12] ), .Y(n120) );
  AND4X1_HVT U185 ( .A1(\match_addr_unencoded_raw[27][12] ), .A2(
        \match_addr_unencoded_raw[26][12] ), .A3(
        \match_addr_unencoded_raw[25][12] ), .A4(
        \match_addr_unencoded_raw[24][12] ), .Y(n127) );
  AND4X1_HVT U186 ( .A1(\match_addr_unencoded_raw[30][12] ), .A2(
        \match_addr_unencoded_raw[2][12] ), .A3(
        \match_addr_unencoded_raw[29][12] ), .A4(
        \match_addr_unencoded_raw[28][12] ), .Y(n128) );
  NAND4X0_HVT U187 ( .A1(n23), .A2(n129), .A3(n130), .A4(n137), .Y(n101) );
  AND4X1_HVT U188 ( .A1(\match_addr_unencoded_raw[9][14] ), .A2(
        \match_addr_unencoded_raw[8][14] ), .A3(
        \match_addr_unencoded_raw[7][14] ), .A4(
        \match_addr_unencoded_raw[6][14] ), .Y(n129) );
  AND4X1_HVT U189 ( .A1(\match_addr_unencoded_raw[27][14] ), .A2(
        \match_addr_unencoded_raw[26][14] ), .A3(
        \match_addr_unencoded_raw[25][14] ), .A4(
        \match_addr_unencoded_raw[24][14] ), .Y(n130) );
  AND4X1_HVT U190 ( .A1(\match_addr_unencoded_raw[30][14] ), .A2(
        \match_addr_unencoded_raw[2][14] ), .A3(
        \match_addr_unencoded_raw[29][14] ), .A4(
        \match_addr_unencoded_raw[28][14] ), .Y(n137) );
  NAND4X0_HVT U191 ( .A1(n24), .A2(n138), .A3(n139), .A4(n140), .Y(n1) );
  AND4X1_HVT U192 ( .A1(n175), .A2(\match_addr_unencoded_raw[9][9] ), .A3(
        \match_addr_unencoded_raw[8][9] ), .A4(
        \match_addr_unencoded_raw[7][9] ), .Y(n138) );
  AND4X1_HVT U193 ( .A1(\match_addr_unencoded_raw[28][9] ), .A2(
        \match_addr_unencoded_raw[27][9] ), .A3(
        \match_addr_unencoded_raw[26][9] ), .A4(
        \match_addr_unencoded_raw[25][9] ), .Y(n139) );
  AND4X1_HVT U194 ( .A1(\match_addr_unencoded_raw[31][9] ), .A2(
        \match_addr_unencoded_raw[30][9] ), .A3(
        \match_addr_unencoded_raw[2][9] ), .A4(
        \match_addr_unencoded_raw[29][9] ), .Y(n140) );
  NAND4X0_HVT U195 ( .A1(n28), .A2(n147), .A3(n148), .A4(n149), .Y(n131) );
  AND4X1_HVT U196 ( .A1(\match_addr_unencoded_raw[9][11] ), .A2(
        \match_addr_unencoded_raw[8][11] ), .A3(
        \match_addr_unencoded_raw[7][11] ), .A4(
        \match_addr_unencoded_raw[6][11] ), .Y(n147) );
  AND4X1_HVT U197 ( .A1(\match_addr_unencoded_raw[27][11] ), .A2(
        \match_addr_unencoded_raw[26][11] ), .A3(
        \match_addr_unencoded_raw[25][11] ), .A4(
        \match_addr_unencoded_raw[24][11] ), .Y(n148) );
  AND4X1_HVT U198 ( .A1(\match_addr_unencoded_raw[30][11] ), .A2(
        \match_addr_unencoded_raw[2][11] ), .A3(
        \match_addr_unencoded_raw[29][11] ), .A4(
        \match_addr_unencoded_raw[28][11] ), .Y(n149) );
  NAND4X0_HVT U199 ( .A1(n29), .A2(n150), .A3(n157), .A4(n158), .Y(n11) );
  AND4X1_HVT U200 ( .A1(\match_addr_unencoded_raw[9][8] ), .A2(
        \match_addr_unencoded_raw[8][8] ), .A3(
        \match_addr_unencoded_raw[7][8] ), .A4(
        \match_addr_unencoded_raw[6][8] ), .Y(n150) );
  AND4X1_HVT U201 ( .A1(\match_addr_unencoded_raw[27][8] ), .A2(
        \match_addr_unencoded_raw[26][8] ), .A3(
        \match_addr_unencoded_raw[25][8] ), .A4(
        \match_addr_unencoded_raw[24][8] ), .Y(n157) );
  AND4X1_HVT U202 ( .A1(\match_addr_unencoded_raw[30][8] ), .A2(
        \match_addr_unencoded_raw[2][8] ), .A3(
        \match_addr_unencoded_raw[29][8] ), .A4(
        \match_addr_unencoded_raw[28][8] ), .Y(n158) );
  NAND4X0_HVT U203 ( .A1(n30), .A2(n159), .A3(n160), .A4(n161), .Y(n141) );
  AND4X1_HVT U204 ( .A1(\match_addr_unencoded_raw[9][10] ), .A2(
        \match_addr_unencoded_raw[8][10] ), .A3(
        \match_addr_unencoded_raw[7][10] ), .A4(
        \match_addr_unencoded_raw[6][10] ), .Y(n159) );
  AND4X1_HVT U205 ( .A1(\match_addr_unencoded_raw[27][10] ), .A2(
        \match_addr_unencoded_raw[26][10] ), .A3(
        \match_addr_unencoded_raw[25][10] ), .A4(
        \match_addr_unencoded_raw[24][10] ), .Y(n160) );
  AND4X1_HVT U206 ( .A1(\match_addr_unencoded_raw[30][10] ), .A2(
        \match_addr_unencoded_raw[2][10] ), .A3(
        \match_addr_unencoded_raw[29][10] ), .A4(
        \match_addr_unencoded_raw[28][10] ), .Y(n161) );
  NAND4X0_HVT U207 ( .A1(n37), .A2(n162), .A3(n163), .A4(n164), .Y(n151) );
  AND4X1_HVT U208 ( .A1(\match_addr_unencoded_raw[9][0] ), .A2(
        \match_addr_unencoded_raw[8][0] ), .A3(
        \match_addr_unencoded_raw[7][0] ), .A4(
        \match_addr_unencoded_raw[6][0] ), .Y(n162) );
  AND4X1_HVT U209 ( .A1(\match_addr_unencoded_raw[27][0] ), .A2(
        \match_addr_unencoded_raw[26][0] ), .A3(
        \match_addr_unencoded_raw[25][0] ), .A4(
        \match_addr_unencoded_raw[24][0] ), .Y(n163) );
  AND4X1_HVT U210 ( .A1(\match_addr_unencoded_raw[30][0] ), .A2(
        \match_addr_unencoded_raw[2][0] ), .A3(
        \match_addr_unencoded_raw[29][0] ), .A4(
        \match_addr_unencoded_raw[28][0] ), .Y(n164) );
  INVX1_HVT U211 ( .A(write_addr[1]), .Y(n182) );
  INVX1_HVT U212 ( .A(write_addr[3]), .Y(n188) );
  NBUFFX2_HVT U213 ( .A(start), .Y(n176) );
  NBUFFX2_HVT U214 ( .A(start), .Y(n175) );
  NBUFFX2_HVT U215 ( .A(write_addr[0]), .Y(n178) );
  NBUFFX2_HVT U216 ( .A(write_addr[0]), .Y(n177) );
  NBUFFX2_HVT U217 ( .A(write_addr[2]), .Y(n184) );
  NBUFFX2_HVT U218 ( .A(write_addr[2]), .Y(n183) );
endmodule

