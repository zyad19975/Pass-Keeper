
module inv_sbox_6 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n184, n196, n197, n198, n199, n200, n201, n202, n208, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672;

  NAND2X0_HVT U3 ( .A1(n344), .A2(n359), .Y(n670) );
  NAND2X0_HVT U5 ( .A1(n669), .A2(n384), .Y(n668) );
  NAND2X0_HVT U7 ( .A1(n331), .A2(n386), .Y(n665) );
  NAND2X0_HVT U8 ( .A1(n332), .A2(n384), .Y(n664) );
  NAND2X0_HVT U9 ( .A1(n390), .A2(n664), .Y(n663) );
  NAND2X0_HVT U10 ( .A1(n672), .A2(n661), .Y(n662) );
  NAND2X0_HVT U11 ( .A1(n262), .A2(n388), .Y(n660) );
  NAND2X0_HVT U12 ( .A1(n393), .A2(n281), .Y(n659) );
  NAND2X0_HVT U13 ( .A1(n387), .A2(n664), .Y(n658) );
  NAND2X0_HVT U15 ( .A1(n381), .A2(n392), .Y(n656) );
  NAND2X0_HVT U19 ( .A1(n394), .A2(n315), .Y(n651) );
  NAND2X0_HVT U25 ( .A1(n197), .A2(n373), .Y(n667) );
  NAND2X0_HVT U32 ( .A1(n374), .A2(n397), .Y(n639) );
  NAND2X0_HVT U35 ( .A1(n664), .A2(n463), .Y(n636) );
  NAND2X0_HVT U38 ( .A1(n281), .A2(n397), .Y(n633) );
  NAND2X0_HVT U42 ( .A1(n666), .A2(n463), .Y(n629) );
  OA21X1_HVT U53 ( .A1(n347), .A2(n621), .A3(n430), .Y(n619) );
  NAND2X0_HVT U55 ( .A1(n387), .A2(n669), .Y(n617) );
  NAND2X0_HVT U66 ( .A1(n265), .A2(n280), .Y(n605) );
  MUX41X1_HVT U67 ( .A1(n420), .A3(n444), .A2(n422), .A4(n605), .S0(n370), 
        .S1(n362), .Y(n604) );
  MUX41X1_HVT U69 ( .A1(n603), .A3(n606), .A2(n604), .A4(n607), .S0(n327), 
        .S1(n379), .Y(n602) );
  MUX41X1_HVT U71 ( .A1(n314), .A3(n222), .A2(n324), .A4(n416), .S0(n364), 
        .S1(n254), .Y(n601) );
  NAND2X0_HVT U72 ( .A1(n382), .A2(n233), .Y(n600) );
  MUX41X1_HVT U73 ( .A1(n644), .A3(n600), .A2(n445), .A4(n371), .S0(n369), 
        .S1(n361), .Y(n599) );
  MUX41X1_HVT U74 ( .A1(n662), .A3(n435), .A2(n434), .A4(n426), .S0(n365), 
        .S1(n254), .Y(n598) );
  MUX41X1_HVT U78 ( .A1(n595), .A3(n599), .A2(n598), .A4(n601), .S0(n327), 
        .S1(n378), .Y(n594) );
  MUX41X1_HVT U79 ( .A1(n250), .A3(n653), .A2(n433), .A4(n654), .S0(n365), 
        .S1(n400), .Y(n593) );
  MUX41X1_HVT U80 ( .A1(n447), .A3(n443), .A2(n663), .A4(n668), .S0(n364), 
        .S1(n254), .Y(n592) );
  NAND2X0_HVT U81 ( .A1(n389), .A2(n665), .Y(n591) );
  AND2X1_HVT U82 ( .A1(n314), .A2(n316), .Y(n590) );
  MUX41X1_HVT U83 ( .A1(n590), .A3(n432), .A2(n304), .A4(n591), .S0(n364), 
        .S1(n254), .Y(n589) );
  MUX41X1_HVT U84 ( .A1(n357), .A3(n250), .A2(n448), .A4(n271), .S0(n365), 
        .S1(n400), .Y(n588) );
  MUX41X1_HVT U85 ( .A1(n588), .A3(n592), .A2(n589), .A4(n593), .S0(n327), 
        .S1(in[1]), .Y(n587) );
  MUX41X1_HVT U87 ( .A1(n410), .A3(n357), .A2(n449), .A4(n350), .S0(n363), 
        .S1(n403), .Y(n586) );
  MUX41X1_HVT U88 ( .A1(n422), .A3(n407), .A2(n641), .A4(n625), .S0(n364), 
        .S1(n403), .Y(n585) );
  NAND2X0_HVT U89 ( .A1(n262), .A2(n459), .Y(n584) );
  MUX41X1_HVT U90 ( .A1(n222), .A3(n233), .A2(n624), .A4(n584), .S0(n364), 
        .S1(n326), .Y(n583) );
  MUX41X1_HVT U96 ( .A1(n444), .A3(n658), .A2(n429), .A4(n450), .S0(n365), 
        .S1(n400), .Y(n577) );
  MUX41X1_HVT U99 ( .A1(n639), .A3(n424), .A2(n623), .A4(n380), .S0(n403), 
        .S1(n362), .Y(n574) );
  NAND2X0_HVT U100 ( .A1(n397), .A2(n458), .Y(n573) );
  MUX41X1_HVT U101 ( .A1(n452), .A3(n659), .A2(n436), .A4(n573), .S0(n326), 
        .S1(n360), .Y(n572) );
  AND2X1_HVT U104 ( .A1(n233), .A2(n383), .Y(n570) );
  MUX41X1_HVT U105 ( .A1(n657), .A3(n453), .A2(n591), .A4(n570), .S0(n365), 
        .S1(n403), .Y(n569) );
  MUX41X1_HVT U107 ( .A1(n452), .A3(n316), .A2(n568), .A4(n298), .S0(n364), 
        .S1(n400), .Y(n567) );
  MUX41X1_HVT U108 ( .A1(n426), .A3(n380), .A2(n350), .A4(n348), .S0(n365), 
        .S1(n254), .Y(n566) );
  MUX41X1_HVT U109 ( .A1(n451), .A3(n407), .A2(n448), .A4(n441), .S0(n364), 
        .S1(n403), .Y(n565) );
  MUX41X1_HVT U110 ( .A1(n565), .A3(n567), .A2(n566), .A4(n569), .S0(n337), 
        .S1(n379), .Y(n564) );
  AO21X1_HVT U112 ( .A1(n439), .A2(n369), .A3(n647), .Y(n562) );
  NAND2X0_HVT U114 ( .A1(n390), .A2(n233), .Y(n560) );
  MUX41X1_HVT U115 ( .A1(n560), .A3(n324), .A2(n439), .A4(n316), .S0(n403), 
        .S1(n362), .Y(n559) );
  MUX41X1_HVT U116 ( .A1(n438), .A3(n431), .A2(n407), .A4(n656), .S0(n363), 
        .S1(n401), .Y(n558) );
  NAND2X0_HVT U118 ( .A1(n262), .A2(n344), .Y(n556) );
  MUX41X1_HVT U119 ( .A1(n454), .A3(n557), .A2(n634), .A4(n556), .S0(n363), 
        .S1(n400), .Y(n555) );
  MUX41X1_HVT U120 ( .A1(n555), .A3(n559), .A2(n558), .A4(n561), .S0(n337), 
        .S1(n379), .Y(n554) );
  MUX41X1_HVT U122 ( .A1(n442), .A3(n353), .A2(n625), .A4(n446), .S0(n363), 
        .S1(n400), .Y(n553) );
  MUX41X1_HVT U124 ( .A1(n355), .A3(n552), .A2(n341), .A4(n340), .S0(n368), 
        .S1(n363), .Y(n551) );
  AOI21X1_HVT U127 ( .A1(n366), .A2(n547), .A3(n414), .Y(n548) );
  NAND2X0_HVT U129 ( .A1(n367), .A2(n672), .Y(n545) );
  MUX41X1_HVT U130 ( .A1(n545), .A3(n546), .A2(n549), .A4(n548), .S0(n370), 
        .S1(n379), .Y(n544) );
  AND2X1_HVT U131 ( .A1(n280), .A2(n322), .Y(n543) );
  MUX41X1_HVT U132 ( .A1(n411), .A3(n543), .A2(n456), .A4(n420), .S0(n369), 
        .S1(n361), .Y(n542) );
  MUX41X1_HVT U133 ( .A1(n457), .A3(n298), .A2(n617), .A4(n412), .S0(n368), 
        .S1(n360), .Y(n541) );
  MUX41X1_HVT U136 ( .A1(n622), .A3(n573), .A2(n539), .A4(n418), .S0(n367), 
        .S1(n403), .Y(n538) );
  MUX41X1_HVT U137 ( .A1(n664), .A3(n239), .A2(n271), .A4(n450), .S0(n370), 
        .S1(n360), .Y(n537) );
  MUX41X1_HVT U139 ( .A1(n536), .A3(n540), .A2(n544), .A4(n550), .S0(n327), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n434), .A3(n354), .A2(n428), .A4(n660), .S0(n369), 
        .S1(n362), .Y(n535) );
  NAND2X0_HVT U141 ( .A1(n381), .A2(n262), .Y(n534) );
  AO21X1_HVT U148 ( .A1(n370), .A2(n415), .A3(n458), .Y(n527) );
  MUX41X1_HVT U155 ( .A1(n428), .A3(n324), .A2(n652), .A4(n429), .S0(n366), 
        .S1(n403), .Y(n520) );
  NAND2X0_HVT U159 ( .A1(n516), .A2(n515), .Y(n517) );
  MUX41X1_HVT U162 ( .A1(n345), .A3(n425), .A2(n636), .A4(n513), .S0(n366), 
        .S1(n401), .Y(n512) );
  NAND2X0_HVT U163 ( .A1(n265), .A2(n459), .Y(n511) );
  MUX41X1_HVT U164 ( .A1(n663), .A3(n511), .A2(n634), .A4(n426), .S0(n363), 
        .S1(n401), .Y(n510) );
  NAND2X0_HVT U166 ( .A1(n661), .A2(n507), .Y(n508) );
  MUX41X1_HVT U174 ( .A1(n449), .A3(n617), .A2(n457), .A4(n463), .S0(n366), 
        .S1(n402), .Y(n499) );
  NAND2X0_HVT U177 ( .A1(n227), .A2(n344), .Y(n497) );
  AND2X1_HVT U179 ( .A1(n314), .A2(n383), .Y(n495) );
  MUX41X1_HVT U183 ( .A1(n440), .A3(n443), .A2(n426), .A4(n629), .S0(n368), 
        .S1(n361), .Y(n491) );
  NAND2X0_HVT U191 ( .A1(n347), .A2(n419), .Y(n484) );
  AND2X1_HVT U192 ( .A1(n435), .A2(n482), .Y(n483) );
  NAND2X0_HVT U194 ( .A1(n297), .A2(n482), .Y(n480) );
  NAND2X0_HVT U198 ( .A1(n392), .A2(n463), .Y(n661) );
  NAND2X0_HVT U200 ( .A1(n384), .A2(n262), .Y(n547) );
  NAND2X0_HVT U207 ( .A1(n262), .A2(n222), .Y(n611) );
  NAND2X0_HVT U1 ( .A1(in[3]), .A2(n375), .Y(n672) );
  INVX2_HVT U2 ( .A(n385), .Y(n315) );
  MUX21X2_HVT U4 ( .A1(n581), .A2(n580), .S0(n261), .Y(n579) );
  MUX21X1_HVT U6 ( .A1(n374), .A2(n463), .S0(n331), .Y(n635) );
  MUX21X2_HVT U14 ( .A1(n597), .A2(n596), .S0(n362), .Y(n595) );
  INVX1_HVT U16 ( .A(n638), .Y(n434) );
  INVX2_HVT U17 ( .A(n404), .Y(n400) );
  IBUFFX2_HVT U18 ( .A(n396), .Y(n395) );
  IBUFFX2_HVT U20 ( .A(n396), .Y(n392) );
  MUX41X1_HVT U21 ( .A1(n635), .A3(n388), .A2(n222), .A4(n390), .S0(n184), 
        .S1(n196), .Y(n500) );
  IBUFFX16_HVT U22 ( .A(n366), .Y(n184) );
  IBUFFX16_HVT U23 ( .A(n401), .Y(n196) );
  INVX1_HVT U24 ( .A(n431), .Y(n235) );
  INVX0_HVT U26 ( .A(n376), .Y(n197) );
  NBUFFX2_HVT U27 ( .A(n464), .Y(n376) );
  INVX0_HVT U28 ( .A(n666), .Y(n412) );
  INVX0_HVT U29 ( .A(n646), .Y(n428) );
  MUX21X1_HVT U30 ( .A1(n459), .A2(n374), .S0(n198), .Y(n525) );
  IBUFFX16_HVT U31 ( .A(n393), .Y(n198) );
  MUX41X1_HVT U33 ( .A1(n525), .A3(n346), .A2(n437), .A4(n304), .S0(n199), 
        .S1(n200), .Y(n524) );
  IBUFFX16_HVT U34 ( .A(n368), .Y(n199) );
  IBUFFX16_HVT U36 ( .A(n360), .Y(n200) );
  NAND2X0_HVT U37 ( .A1(n630), .A2(n201), .Y(n202) );
  NAND2X0_HVT U39 ( .A1(n445), .A2(n320), .Y(n208) );
  NAND2X0_HVT U40 ( .A1(n202), .A2(n208), .Y(n487) );
  IBUFFX2_HVT U41 ( .A(n320), .Y(n201) );
  NAND2X0_HVT U43 ( .A1(n458), .A2(n218), .Y(n219) );
  NAND2X0_HVT U44 ( .A1(n374), .A2(n395), .Y(n220) );
  NAND2X0_HVT U45 ( .A1(n219), .A2(n220), .Y(n476) );
  IBUFFX2_HVT U46 ( .A(n395), .Y(n218) );
  INVX0_HVT U47 ( .A(n369), .Y(n320) );
  INVX0_HVT U48 ( .A(n476), .Y(n445) );
  INVX1_HVT U49 ( .A(n461), .Y(n221) );
  INVX2_HVT U50 ( .A(n221), .Y(n222) );
  MUX21X2_HVT U51 ( .A1(n357), .A2(n646), .S0(n334), .Y(n523) );
  INVX0_HVT U52 ( .A(n646), .Y(n270) );
  INVX1_HVT U54 ( .A(n647), .Y(n427) );
  MUX21X2_HVT U56 ( .A1(n359), .A2(n461), .S0(n227), .Y(n647) );
  MUX21X2_HVT U57 ( .A1(n669), .A2(n346), .S0(n223), .Y(n608) );
  IBUFFX16_HVT U58 ( .A(n367), .Y(n223) );
  MUX41X1_HVT U59 ( .A1(n579), .A3(n583), .A2(n585), .A4(n586), .S0(n379), 
        .S1(n327), .Y(n578) );
  INVX0_HVT U60 ( .A(n635), .Y(n436) );
  MUX21X2_HVT U61 ( .A1(n562), .A2(n563), .S0(n366), .Y(n561) );
  INVX0_HVT U62 ( .A(n331), .Y(n285) );
  INVX1_HVT U63 ( .A(n650), .Y(n426) );
  NAND2X0_HVT U64 ( .A1(n381), .A2(n224), .Y(n225) );
  NAND2X0_HVT U65 ( .A1(n222), .A2(n391), .Y(n226) );
  NAND2X0_HVT U68 ( .A1(n225), .A2(n226), .Y(n640) );
  IBUFFX2_HVT U70 ( .A(n391), .Y(n224) );
  INVX0_HVT U75 ( .A(n640), .Y(n433) );
  NBUFFX2_HVT U76 ( .A(n395), .Y(n227) );
  MUX41X1_HVT U77 ( .A1(n575), .A3(n572), .A2(n577), .A4(n574), .S0(n313), 
        .S1(n378), .Y(n571) );
  INVX0_HVT U86 ( .A(n347), .Y(n229) );
  INVX2_HVT U91 ( .A(n404), .Y(n402) );
  MUX41X1_HVT U92 ( .A1(n437), .A3(n643), .A2(n576), .A4(n451), .S0(n228), 
        .S1(n310), .Y(n575) );
  IBUFFX16_HVT U93 ( .A(n309), .Y(n228) );
  MUX21X1_HVT U94 ( .A1(n374), .A2(n373), .S0(n322), .Y(n626) );
  INVX1_HVT U95 ( .A(n322), .Y(n394) );
  INVX1_HVT U97 ( .A(n465), .Y(n457) );
  NAND2X0_HVT U98 ( .A1(n242), .A2(n243), .Y(n610) );
  MUX21X1_HVT U102 ( .A1(n350), .A2(n340), .S0(n229), .Y(n349) );
  MUX21X2_HVT U103 ( .A1(n382), .A2(n374), .S0(n395), .Y(n646) );
  NBUFFX2_HVT U106 ( .A(n464), .Y(n374) );
  MUX41X1_HVT U111 ( .A1(n618), .A3(n616), .A2(n614), .A4(n610), .S0(n377), 
        .S1(n351), .Y(n609) );
  NAND2X0_HVT U113 ( .A1(n619), .A2(n230), .Y(n231) );
  NAND2X0_HVT U117 ( .A1(n620), .A2(n249), .Y(n232) );
  NAND2X0_HVT U121 ( .A1(n231), .A2(n232), .Y(n618) );
  INVX0_HVT U123 ( .A(n249), .Y(n230) );
  IBUFFX2_HVT U125 ( .A(n367), .Y(n249) );
  INVX1_HVT U126 ( .A(n414), .Y(n233) );
  MUX21X1_HVT U128 ( .A1(n517), .A2(n518), .S0(n360), .Y(n514) );
  MUX21X2_HVT U134 ( .A1(n508), .A2(n509), .S0(n362), .Y(n506) );
  MUX41X1_HVT U135 ( .A1(n632), .A3(n534), .A2(n428), .A4(n455), .S0(n234), 
        .S1(n400), .Y(n533) );
  IBUFFX16_HVT U138 ( .A(n360), .Y(n234) );
  AO21X2_HVT U142 ( .A1(n394), .A2(n343), .A3(n347), .Y(n482) );
  NAND2X0_HVT U143 ( .A1(n235), .A2(n236), .Y(n237) );
  AND2X1_HVT U144 ( .A1(n237), .A2(n611), .Y(n486) );
  INVX0_HVT U145 ( .A(n323), .Y(n236) );
  INVX0_HVT U146 ( .A(n370), .Y(n323) );
  INVX0_HVT U147 ( .A(n642), .Y(n238) );
  INVX0_HVT U149 ( .A(n238), .Y(n239) );
  MUX21X1_HVT U150 ( .A1(n429), .A2(n421), .S0(n370), .Y(n620) );
  MUX41X1_HVT U151 ( .A1(n352), .A3(n356), .A2(n504), .A4(n355), .S0(n240), 
        .S1(n403), .Y(n503) );
  IBUFFX16_HVT U152 ( .A(n366), .Y(n240) );
  NAND2X0_HVT U153 ( .A1(n612), .A2(n241), .Y(n242) );
  NAND2X0_HVT U154 ( .A1(n613), .A2(n248), .Y(n243) );
  INVX0_HVT U156 ( .A(n248), .Y(n241) );
  MUX21X1_HVT U157 ( .A1(n340), .A2(n617), .S0(n369), .Y(n613) );
  IBUFFX2_HVT U158 ( .A(n367), .Y(n248) );
  NAND2X0_HVT U160 ( .A1(n393), .A2(n671), .Y(n669) );
  INVX2_HVT U161 ( .A(n369), .Y(n334) );
  MUX21X2_HVT U165 ( .A1(n357), .A2(n623), .S0(n370), .Y(n488) );
  NAND2X0_HVT U167 ( .A1(n375), .A2(n373), .Y(n246) );
  NAND2X0_HVT U168 ( .A1(n244), .A2(n245), .Y(n247) );
  NAND2X0_HVT U169 ( .A1(n247), .A2(n246), .Y(n655) );
  INVX0_HVT U170 ( .A(n375), .Y(n244) );
  INVX0_HVT U171 ( .A(n373), .Y(n245) );
  NBUFFX2_HVT U172 ( .A(n464), .Y(n375) );
  IBUFFX2_HVT U173 ( .A(n632), .Y(n438) );
  INVX1_HVT U175 ( .A(n380), .Y(n463) );
  INVX1_HVT U176 ( .A(n672), .Y(n461) );
  MUX21X2_HVT U178 ( .A1(n554), .A2(n564), .S0(in[7]), .Y(out[3]) );
  MUX21X1_HVT U180 ( .A1(n416), .A2(n381), .S0(n370), .Y(n580) );
  IBUFFX2_HVT U181 ( .A(n346), .Y(n649) );
  MUX21X2_HVT U182 ( .A1(n300), .A2(n626), .S0(n301), .Y(n299) );
  NBUFFX2_HVT U184 ( .A(n431), .Y(n250) );
  NAND2X0_HVT U185 ( .A1(n587), .A2(n251), .Y(n252) );
  NAND2X0_HVT U186 ( .A1(n594), .A2(in[7]), .Y(n253) );
  NAND2X0_HVT U187 ( .A1(n252), .A2(n253), .Y(out[1]) );
  IBUFFX2_HVT U188 ( .A(in[7]), .Y(n251) );
  NBUFFX2_HVT U189 ( .A(n401), .Y(n254) );
  IBUFFX2_HVT U190 ( .A(n404), .Y(n401) );
  IBUFFX2_HVT U193 ( .A(n400), .Y(n263) );
  INVX1_HVT U195 ( .A(n644), .Y(n429) );
  NAND2X0_HVT U196 ( .A1(n578), .A2(n255), .Y(n256) );
  NAND2X0_HVT U197 ( .A1(n571), .A2(n312), .Y(n257) );
  NAND2X0_HVT U199 ( .A1(n256), .A2(n257), .Y(out[2]) );
  INVX1_HVT U201 ( .A(n312), .Y(n255) );
  IBUFFX2_HVT U202 ( .A(in[7]), .Y(n312) );
  INVX1_HVT U203 ( .A(n322), .Y(n331) );
  NAND2X0_HVT U204 ( .A1(n505), .A2(n292), .Y(n293) );
  XOR2X1_HVT U205 ( .A1(n383), .A2(n395), .Y(n623) );
  INVX2_HVT U206 ( .A(n404), .Y(n403) );
  NAND2X0_HVT U208 ( .A1(n386), .A2(n258), .Y(n259) );
  NAND2X0_HVT U209 ( .A1(n582), .A2(n266), .Y(n260) );
  NAND2X0_HVT U210 ( .A1(n259), .A2(n260), .Y(n581) );
  INVX0_HVT U211 ( .A(n266), .Y(n258) );
  IBUFFX16_HVT U212 ( .A(n367), .Y(n261) );
  INVX1_HVT U213 ( .A(n332), .Y(n262) );
  MUX41X1_HVT U214 ( .A1(n626), .A3(n405), .A2(n495), .A4(n639), .S0(n263), 
        .S1(n291), .Y(n494) );
  INVX0_HVT U215 ( .A(n394), .Y(n295) );
  INVX1_HVT U216 ( .A(n642), .Y(n431) );
  MUX41X1_HVT U217 ( .A1(n627), .A3(n222), .A2(n497), .A4(n356), .S0(n264), 
        .S1(n310), .Y(n496) );
  IBUFFX16_HVT U218 ( .A(n366), .Y(n264) );
  INVX2_HVT U219 ( .A(n326), .Y(n310) );
  INVX2_HVT U220 ( .A(n302), .Y(n265) );
  MUX21X2_HVT U221 ( .A1(n426), .A2(n608), .S0(n358), .Y(n607) );
  MUX21X2_HVT U222 ( .A1(n348), .A2(n381), .S0(n322), .Y(n346) );
  IBUFFX2_HVT U223 ( .A(n393), .Y(n308) );
  IBUFFX2_HVT U224 ( .A(n391), .Y(n266) );
  INVX1_HVT U225 ( .A(n265), .Y(n306) );
  INVX1_HVT U226 ( .A(n332), .Y(n302) );
  NAND2X0_HVT U227 ( .A1(n427), .A2(n267), .Y(n268) );
  NAND2X0_HVT U228 ( .A1(n615), .A2(n358), .Y(n269) );
  NAND2X0_HVT U229 ( .A1(n268), .A2(n269), .Y(n614) );
  INVX0_HVT U230 ( .A(n358), .Y(n267) );
  INVX1_HVT U231 ( .A(n270), .Y(n271) );
  MUX21X1_HVT U232 ( .A1(n668), .A2(n428), .S0(n325), .Y(n615) );
  MUX41X1_HVT U233 ( .A1(n487), .A3(n486), .A2(n488), .A4(n489), .S0(n361), 
        .S1(n378), .Y(n485) );
  MUX41X1_HVT U234 ( .A1(n493), .A3(n490), .A2(n485), .A4(n479), .S0(n351), 
        .S1(n328), .Y(out[7]) );
  INVX0_HVT U235 ( .A(n272), .Y(n489) );
  MUX41X1_HVT U236 ( .A1(n481), .A3(n480), .A2(n483), .A4(n484), .S0(n364), 
        .S1(n378), .Y(n479) );
  INVX1_HVT U237 ( .A(in[7]), .Y(n328) );
  INVX1_HVT U238 ( .A(in[6]), .Y(n464) );
  INVX0_HVT U239 ( .A(n464), .Y(n359) );
  MUX21X1_HVT U240 ( .A1(n273), .A2(n474), .S0(n368), .Y(n272) );
  NAND2X0_HVT U241 ( .A1(n463), .A2(n322), .Y(n273) );
  IBUFFX2_HVT U242 ( .A(n474), .Y(n447) );
  NAND2X0_HVT U243 ( .A1(n611), .A2(n368), .Y(n274) );
  INVX0_HVT U244 ( .A(n650), .Y(n275) );
  NAND2X0_HVT U245 ( .A1(n274), .A2(n275), .Y(n612) );
  NBUFFX4_HVT U246 ( .A(n460), .Y(n373) );
  INVX1_HVT U247 ( .A(n299), .Y(n481) );
  NAND2X0_HVT U248 ( .A1(n459), .A2(n276), .Y(n277) );
  NAND2X0_HVT U249 ( .A1(n222), .A2(n285), .Y(n278) );
  NAND2X0_HVT U250 ( .A1(n277), .A2(n278), .Y(n643) );
  INVX0_HVT U251 ( .A(n285), .Y(n276) );
  INVX0_HVT U252 ( .A(n359), .Y(n279) );
  INVX1_HVT U253 ( .A(n279), .Y(n280) );
  INVX1_HVT U254 ( .A(n305), .Y(n281) );
  INVX0_HVT U255 ( .A(n371), .Y(n305) );
  NBUFFX2_HVT U256 ( .A(n460), .Y(n372) );
  NAND2X0_HVT U257 ( .A1(n492), .A2(n282), .Y(n283) );
  NAND2X0_HVT U258 ( .A1(n491), .A2(n296), .Y(n284) );
  NAND2X0_HVT U259 ( .A1(n283), .A2(n284), .Y(n490) );
  INVX0_HVT U260 ( .A(n296), .Y(n282) );
  IBUFFX2_HVT U261 ( .A(n378), .Y(n296) );
  NAND2X0_HVT U262 ( .A1(n519), .A2(n286), .Y(n287) );
  NAND2X0_HVT U263 ( .A1(n529), .A2(n311), .Y(n288) );
  NAND2X0_HVT U264 ( .A1(n287), .A2(n288), .Y(out[5]) );
  INVX1_HVT U265 ( .A(n311), .Y(n286) );
  IBUFFX2_HVT U266 ( .A(n328), .Y(n311) );
  MUX21X1_HVT U267 ( .A1(n385), .A2(n464), .S0(n308), .Y(n319) );
  NAND2X0_HVT U268 ( .A1(n382), .A2(n289), .Y(n290) );
  NAND2X0_HVT U269 ( .A1(n278), .A2(n290), .Y(n472) );
  INVX0_HVT U270 ( .A(n295), .Y(n289) );
  INVX0_HVT U271 ( .A(n472), .Y(n449) );
  INVX2_HVT U272 ( .A(n372), .Y(n344) );
  IBUFFX2_HVT U273 ( .A(n366), .Y(n291) );
  MUX21X2_HVT U274 ( .A1(n522), .A2(n523), .S0(n361), .Y(n521) );
  NAND2X0_HVT U275 ( .A1(n498), .A2(n328), .Y(n294) );
  NAND2X0_HVT U276 ( .A1(n293), .A2(n294), .Y(out[6]) );
  INVX0_HVT U277 ( .A(n328), .Y(n292) );
  INVX0_HVT U278 ( .A(n355), .Y(n300) );
  INVX0_HVT U279 ( .A(n413), .Y(n297) );
  INVX0_HVT U280 ( .A(n297), .Y(n298) );
  IBUFFX16_HVT U281 ( .A(n368), .Y(n301) );
  MUX21X1_HVT U282 ( .A1(n462), .A2(n222), .S0(n302), .Y(n504) );
  MUX41X1_HVT U283 ( .A1(n531), .A3(n591), .A2(n640), .A4(n453), .S0(n303), 
        .S1(n320), .Y(n530) );
  IBUFFX16_HVT U284 ( .A(n325), .Y(n303) );
  MUX21X1_HVT U285 ( .A1(n305), .A2(n380), .S0(n332), .Y(n304) );
  MUX21X1_HVT U286 ( .A1(n374), .A2(n461), .S0(n306), .Y(n502) );
  MUX41X1_HVT U287 ( .A1(n502), .A3(n584), .A2(n649), .A4(n352), .S0(n307), 
        .S1(n400), .Y(n501) );
  IBUFFX16_HVT U288 ( .A(n366), .Y(n307) );
  MUX21X1_HVT U289 ( .A1(n462), .A2(n281), .S0(n308), .Y(n628) );
  INVX1_HVT U290 ( .A(n385), .Y(n462) );
  IBUFFX16_HVT U291 ( .A(n365), .Y(n309) );
  INVX1_HVT U292 ( .A(in[4]), .Y(n404) );
  IBUFFX16_HVT U293 ( .A(n337), .Y(n313) );
  INVX1_HVT U294 ( .A(n412), .Y(n314) );
  NAND2X0_HVT U295 ( .A1(n391), .A2(n390), .Y(n666) );
  INVX0_HVT U296 ( .A(n629), .Y(n413) );
  INVX0_HVT U297 ( .A(n396), .Y(n321) );
  INVX1_HVT U298 ( .A(n315), .Y(n316) );
  INVX1_HVT U299 ( .A(n628), .Y(n440) );
  AO21X1_HVT U300 ( .A1(n322), .A2(n672), .A3(n347), .Y(n515) );
  MUX41X1_HVT U301 ( .A1(n514), .A3(n512), .A2(n510), .A4(n506), .S0(n317), 
        .S1(n318), .Y(n505) );
  IBUFFX16_HVT U302 ( .A(n378), .Y(n317) );
  IBUFFX16_HVT U303 ( .A(n337), .Y(n318) );
  INVX1_HVT U304 ( .A(n319), .Y(n630) );
  NAND2X0_HVT U305 ( .A1(n602), .A2(n328), .Y(n338) );
  OA21X1_HVT U306 ( .A1(n408), .A2(n347), .A3(n417), .Y(n522) );
  NBUFFX2_HVT U307 ( .A(n402), .Y(n369) );
  INVX1_HVT U308 ( .A(n645), .Y(n350) );
  INVX1_HVT U309 ( .A(n351), .Y(n327) );
  INVX1_HVT U310 ( .A(n648), .Y(n340) );
  INVX1_HVT U311 ( .A(n351), .Y(n337) );
  INVX0_HVT U312 ( .A(n365), .Y(n325) );
  INVX0_HVT U313 ( .A(n363), .Y(n333) );
  INVX0_HVT U314 ( .A(n364), .Y(n342) );
  INVX1_HVT U315 ( .A(in[1]), .Y(n377) );
  INVX2_HVT U316 ( .A(n321), .Y(n322) );
  INVX1_HVT U317 ( .A(in[0]), .Y(n396) );
  MUX21X2_HVT U318 ( .A1(n528), .A2(n527), .S0(n367), .Y(n526) );
  MUX21X2_HVT U319 ( .A1(n456), .A2(n411), .S0(n368), .Y(n528) );
  AO21X1_HVT U320 ( .A1(n382), .A2(n669), .A3(n334), .Y(n507) );
  INVX1_HVT U321 ( .A(n405), .Y(n324) );
  INVX0_HVT U322 ( .A(n660), .Y(n405) );
  INVX1_HVT U323 ( .A(n396), .Y(n393) );
  INVX1_HVT U324 ( .A(n392), .Y(n397) );
  INVX1_HVT U325 ( .A(n396), .Y(n391) );
  MUX41X1_HVT U326 ( .A1(n617), .A3(n350), .A2(n380), .A4(n443), .S0(n325), 
        .S1(n347), .Y(n616) );
  MUX41X1_HVT U327 ( .A1(n530), .A3(n532), .A2(n533), .A4(n535), .S0(n379), 
        .S1(n327), .Y(n529) );
  NBUFFX2_HVT U328 ( .A(n402), .Y(n326) );
  INVX1_HVT U329 ( .A(n402), .Y(n347) );
  NAND2X0_HVT U330 ( .A1(n496), .A2(n379), .Y(n329) );
  NAND2X0_HVT U331 ( .A1(n494), .A2(n377), .Y(n330) );
  NAND2X0_HVT U332 ( .A1(n329), .A2(n330), .Y(n493) );
  IBUFFX2_HVT U333 ( .A(n396), .Y(n332) );
  MUX41X1_HVT U334 ( .A1(n304), .A3(n410), .A2(n669), .A4(n413), .S0(n333), 
        .S1(n323), .Y(n492) );
  NAND2X0_HVT U335 ( .A1(n628), .A2(n334), .Y(n335) );
  NAND2X0_HVT U336 ( .A1(n446), .A2(n369), .Y(n336) );
  NAND2X0_HVT U337 ( .A1(n335), .A2(n336), .Y(n518) );
  INVX1_HVT U338 ( .A(n377), .Y(n378) );
  MUX41X1_HVT U339 ( .A1(n521), .A3(n526), .A2(n520), .A4(n524), .S0(n337), 
        .S1(n377), .Y(n519) );
  NAND2X0_HVT U340 ( .A1(n609), .A2(in[7]), .Y(n339) );
  NAND2X0_HVT U341 ( .A1(n338), .A2(n339), .Y(out[0]) );
  INVX1_HVT U342 ( .A(n340), .Y(n341) );
  OA21X2_HVT U343 ( .A1(n409), .A2(n334), .A3(n650), .Y(n596) );
  MUX41X1_HVT U344 ( .A1(n390), .A3(n421), .A2(n344), .A4(n420), .S0(n342), 
        .S1(n334), .Y(n603) );
  INVX0_HVT U345 ( .A(n345), .Y(n627) );
  INVX1_HVT U346 ( .A(in[5]), .Y(n351) );
  INVX1_HVT U347 ( .A(n475), .Y(n446) );
  MUX21X1_HVT U348 ( .A1(n381), .A2(n281), .S0(n395), .Y(n650) );
  MUX41X1_HVT U349 ( .A1(n633), .A3(n424), .A2(n425), .A4(n423), .S0(n342), 
        .S1(n334), .Y(n606) );
  INVX1_HVT U350 ( .A(n348), .Y(n343) );
  INVX0_HVT U351 ( .A(n348), .Y(n458) );
  NAND2X0_HVT U352 ( .A1(n371), .A2(n375), .Y(n348) );
  INVX0_HVT U353 ( .A(n349), .Y(n509) );
  MUX21X1_HVT U354 ( .A1(n672), .A2(n383), .S0(n322), .Y(n345) );
  MUX41X1_HVT U355 ( .A1(n341), .A3(n651), .A2(n440), .A4(n459), .S0(n333), 
        .S1(n347), .Y(n532) );
  NBUFFX2_HVT U356 ( .A(n460), .Y(n371) );
  MUX41X1_HVT U357 ( .A1(n503), .A3(n501), .A2(n500), .A4(n499), .S0(n377), 
        .S1(n351), .Y(n498) );
  INVX0_HVT U358 ( .A(n573), .Y(n408) );
  NBUFFX2_HVT U359 ( .A(n671), .Y(n388) );
  NBUFFX2_HVT U360 ( .A(n671), .Y(n389) );
  AND2X1_HVT U361 ( .A1(n666), .A2(n388), .Y(n352) );
  AND2X1_HVT U362 ( .A1(n388), .A2(n656), .Y(n353) );
  NAND2X0_HVT U363 ( .A1(n371), .A2(n375), .Y(n671) );
  MUX21X1_HVT U364 ( .A1(n458), .A2(n463), .S0(n394), .Y(n638) );
  MUX21X1_HVT U365 ( .A1(n376), .A2(n458), .S0(n393), .Y(n645) );
  INVX1_HVT U366 ( .A(n383), .Y(n459) );
  MUX21X1_HVT U367 ( .A1(n463), .A2(n373), .S0(n331), .Y(n632) );
  MUX21X1_HVT U368 ( .A1(n373), .A2(n343), .S0(n331), .Y(n641) );
  MUX21X1_HVT U369 ( .A1(n458), .A2(n315), .S0(n391), .Y(n621) );
  MUX21X1_HVT U370 ( .A1(n383), .A2(n386), .S0(n392), .Y(n513) );
  MUX21X1_HVT U371 ( .A1(n389), .A2(n384), .S0(n392), .Y(n531) );
  MUX21X1_HVT U372 ( .A1(n382), .A2(n459), .S0(n265), .Y(n637) );
  MUX21X1_HVT U373 ( .A1(n383), .A2(n348), .S0(n265), .Y(n466) );
  MUX21X1_HVT U374 ( .A1(n463), .A2(n374), .S0(n392), .Y(n467) );
  XNOR2X1_HVT U375 ( .A1(n389), .A2(n393), .Y(n354) );
  MUX21X1_HVT U376 ( .A1(n638), .A2(n353), .S0(n361), .Y(n546) );
  MUX21X1_HVT U377 ( .A1(n381), .A2(n374), .S0(n369), .Y(n582) );
  MUX21X1_HVT U378 ( .A1(n455), .A2(n354), .S0(n367), .Y(n549) );
  XOR2X1_HVT U379 ( .A1(n385), .A2(n391), .Y(n624) );
  MUX21X1_HVT U380 ( .A1(n315), .A2(n281), .S0(n265), .Y(n475) );
  MUX21X1_HVT U381 ( .A1(n281), .A2(n388), .S0(n391), .Y(n474) );
  MUX21X1_HVT U382 ( .A1(n387), .A2(n388), .S0(n332), .Y(n653) );
  MUX21X1_HVT U383 ( .A1(n414), .A2(n630), .S0(n370), .Y(n563) );
  XOR2X1_HVT U384 ( .A1(n380), .A2(n391), .Y(n625) );
  MUX21X1_HVT U385 ( .A1(n672), .A2(n389), .S0(n391), .Y(n657) );
  MUX21X1_HVT U386 ( .A1(n386), .A2(n373), .S0(n392), .Y(n652) );
  MUX21X1_HVT U387 ( .A1(n374), .A2(n389), .S0(n394), .Y(n568) );
  XOR2X1_HVT U388 ( .A1(n390), .A2(n391), .Y(n634) );
  MUX21X1_HVT U389 ( .A1(n374), .A2(n382), .S0(n331), .Y(n631) );
  MUX21X1_HVT U390 ( .A1(n387), .A2(n374), .S0(n227), .Y(n552) );
  MUX21X1_HVT U391 ( .A1(n371), .A2(n386), .S0(n394), .Y(n469) );
  NBUFFX2_HVT U392 ( .A(n402), .Y(n368) );
  NBUFFX2_HVT U393 ( .A(n402), .Y(n370) );
  AND2X1_HVT U394 ( .A1(n392), .A2(n374), .Y(n355) );
  NBUFFX2_HVT U395 ( .A(n667), .Y(n383) );
  NBUFFX2_HVT U396 ( .A(n655), .Y(n380) );
  AND2X1_HVT U397 ( .A1(n462), .A2(n262), .Y(n356) );
  MUX21X1_HVT U398 ( .A1(n551), .A2(n553), .S0(n378), .Y(n550) );
  NBUFFX2_HVT U399 ( .A(n670), .Y(n385) );
  NBUFFX2_HVT U400 ( .A(n655), .Y(n381) );
  NBUFFX2_HVT U401 ( .A(n655), .Y(n382) );
  AND2X1_HVT U402 ( .A1(n387), .A2(n397), .Y(n357) );
  NBUFFX2_HVT U403 ( .A(n667), .Y(n384) );
  NBUFFX2_HVT U404 ( .A(n670), .Y(n387) );
  MUX21X1_HVT U405 ( .A1(n446), .A2(n406), .S0(n370), .Y(n597) );
  NBUFFX2_HVT U406 ( .A(n670), .Y(n386) );
  NBUFFX2_HVT U407 ( .A(n399), .Y(n366) );
  NBUFFX2_HVT U408 ( .A(n399), .Y(n367) );
  XNOR2X1_HVT U409 ( .A1(n347), .A2(n363), .Y(n358) );
  NBUFFX2_HVT U410 ( .A(n398), .Y(n363) );
  NBUFFX2_HVT U411 ( .A(n399), .Y(n364) );
  NBUFFX2_HVT U412 ( .A(n399), .Y(n365) );
  NBUFFX2_HVT U413 ( .A(n398), .Y(n361) );
  NBUFFX2_HVT U414 ( .A(n398), .Y(n362) );
  NBUFFX2_HVT U415 ( .A(n398), .Y(n360) );
  INVX1_HVT U416 ( .A(n377), .Y(n379) );
  INVX0_HVT U417 ( .A(in[3]), .Y(n460) );
  MUX21X1_HVT U418 ( .A1(n343), .A2(n344), .S0(n395), .Y(n648) );
  MUX21X1_HVT U419 ( .A1(n541), .A2(n542), .S0(n379), .Y(n540) );
  MUX21X1_HVT U420 ( .A1(n537), .A2(n538), .S0(n378), .Y(n536) );
  MUX21X1_HVT U421 ( .A1(n384), .A2(n344), .S0(n331), .Y(n576) );
  MUX21X1_HVT U422 ( .A1(n461), .A2(n344), .S0(n394), .Y(n465) );
  MUX21X1_HVT U423 ( .A1(n315), .A2(n459), .S0(n393), .Y(n557) );
  MUX21X1_HVT U424 ( .A1(n344), .A2(n384), .S0(n394), .Y(n470) );
  MUX21X1_HVT U425 ( .A1(n390), .A2(n344), .S0(n393), .Y(n516) );
  MUX21X1_HVT U426 ( .A1(n344), .A2(n390), .S0(n331), .Y(n471) );
  MUX21X1_HVT U427 ( .A1(n374), .A2(n344), .S0(n227), .Y(n644) );
  NBUFFX2_HVT U428 ( .A(in[2]), .Y(n399) );
  NBUFFX2_HVT U429 ( .A(in[2]), .Y(n398) );
  NBUFFX2_HVT U430 ( .A(n672), .Y(n390) );
  MUX21X1_HVT U431 ( .A1(n343), .A2(n280), .S0(n391), .Y(n539) );
  XOR2X1_HVT U432 ( .A1(n393), .A2(n280), .Y(n622) );
  MUX21X1_HVT U433 ( .A1(n386), .A2(n280), .S0(n331), .Y(n473) );
  MUX21X1_HVT U434 ( .A1(n359), .A2(n387), .S0(n393), .Y(n477) );
  MUX21X1_HVT U435 ( .A1(n359), .A2(n672), .S0(n332), .Y(n654) );
  MUX21X1_HVT U436 ( .A1(n371), .A2(n280), .S0(n392), .Y(n468) );
  MUX21X1_HVT U437 ( .A1(n384), .A2(n359), .S0(n394), .Y(n642) );
  MUX21X1_HVT U438 ( .A1(n359), .A2(n459), .S0(n227), .Y(n478) );
  INVX0_HVT U439 ( .A(n639), .Y(n406) );
  INVX0_HVT U440 ( .A(n633), .Y(n407) );
  INVX0_HVT U441 ( .A(n534), .Y(n409) );
  INVX0_HVT U442 ( .A(n669), .Y(n410) );
  INVX0_HVT U443 ( .A(n668), .Y(n411) );
  INVX0_HVT U444 ( .A(n665), .Y(n414) );
  INVX0_HVT U445 ( .A(n664), .Y(n415) );
  INVX0_HVT U446 ( .A(n636), .Y(n416) );
  INVX0_HVT U447 ( .A(n658), .Y(n417) );
  INVX0_HVT U448 ( .A(n663), .Y(n418) );
  INVX0_HVT U449 ( .A(n659), .Y(n419) );
  INVX0_HVT U450 ( .A(n657), .Y(n420) );
  INVX0_HVT U451 ( .A(n656), .Y(n421) );
  INVX0_HVT U452 ( .A(n654), .Y(n422) );
  INVX0_HVT U453 ( .A(n653), .Y(n423) );
  INVX0_HVT U454 ( .A(n652), .Y(n424) );
  INVX0_HVT U455 ( .A(n651), .Y(n425) );
  INVX0_HVT U456 ( .A(n643), .Y(n430) );
  INVX0_HVT U457 ( .A(n641), .Y(n432) );
  INVX0_HVT U458 ( .A(n637), .Y(n435) );
  INVX0_HVT U459 ( .A(n634), .Y(n437) );
  INVX0_HVT U460 ( .A(n631), .Y(n439) );
  INVX0_HVT U461 ( .A(n625), .Y(n441) );
  INVX0_HVT U462 ( .A(n662), .Y(n442) );
  INVX0_HVT U463 ( .A(n478), .Y(n443) );
  INVX0_HVT U464 ( .A(n477), .Y(n444) );
  INVX0_HVT U465 ( .A(n473), .Y(n448) );
  INVX0_HVT U466 ( .A(n471), .Y(n450) );
  INVX0_HVT U467 ( .A(n470), .Y(n451) );
  INVX0_HVT U468 ( .A(n469), .Y(n452) );
  INVX0_HVT U469 ( .A(n468), .Y(n453) );
  INVX0_HVT U470 ( .A(n516), .Y(n454) );
  INVX0_HVT U471 ( .A(n467), .Y(n455) );
  INVX0_HVT U472 ( .A(n466), .Y(n456) );
endmodule

