
module ram_dp_DATA_WIDTH4_ADDR_WIDTH4_5 ( clk, rst, write, a_addr, a_din, 
        b_din, b_dout );
  input [3:0] a_addr;
  input [3:0] a_din;
  input [3:0] b_din;
  output [15:0] b_dout;
  input clk, rst, write;
  wire   N17, N18, N19, N20, \mem[15][15] , \mem[15][14] , \mem[15][13] ,
         \mem[15][12] , \mem[15][11] , \mem[15][10] , \mem[15][9] ,
         \mem[15][8] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][15] ,
         \mem[14][14] , \mem[14][13] , \mem[14][12] , \mem[14][11] ,
         \mem[14][10] , \mem[14][9] , \mem[14][8] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][15] , \mem[13][14] , \mem[13][13] ,
         \mem[13][12] , \mem[13][11] , \mem[13][10] , \mem[13][9] ,
         \mem[13][8] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][15] ,
         \mem[12][14] , \mem[12][13] , \mem[12][12] , \mem[12][11] ,
         \mem[12][10] , \mem[12][9] , \mem[12][8] , \mem[12][7] , \mem[12][6] ,
         \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] , \mem[12][1] ,
         \mem[12][0] , \mem[11][15] , \mem[11][14] , \mem[11][13] ,
         \mem[11][12] , \mem[11][11] , \mem[11][10] , \mem[11][9] ,
         \mem[11][8] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][15] , \mem[9][14] , \mem[9][13] , \mem[9][12] ,
         \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] , \mem[9][7] ,
         \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] ,
         \mem[9][1] , \mem[9][0] , \mem[8][15] , \mem[8][14] , \mem[8][13] ,
         \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] , \mem[8][8] ,
         \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] , \mem[8][3] ,
         \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][15] , \mem[7][14] ,
         \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] ,
         \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][15] ,
         \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] ,
         \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][15] , \mem[3][14] , \mem[3][13] ,
         \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] ,
         \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] ,
         \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][15] ,
         \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N539, N540, N541, N542, N543, N544, N545, N546, N547,
         N548, N549, N550, N551, N552, N553, N554, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n302, n320, n338, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580;
  assign N17 = b_din[0];
  assign N18 = b_din[1];
  assign N19 = b_din[2];
  assign N20 = b_din[3];

  DFFNX1_HVT \b_dout_reg[15]  ( .D(N539), .CLK(clk), .Q(b_dout[15]) );
  DFFNX1_HVT \b_dout_reg[14]  ( .D(N540), .CLK(clk), .Q(b_dout[14]) );
  DFFNX1_HVT \b_dout_reg[13]  ( .D(N541), .CLK(clk), .Q(b_dout[13]) );
  DFFNX1_HVT \b_dout_reg[12]  ( .D(N542), .CLK(clk), .Q(b_dout[12]) );
  DFFNX1_HVT \b_dout_reg[11]  ( .D(N543), .CLK(clk), .Q(b_dout[11]) );
  DFFNX1_HVT \b_dout_reg[10]  ( .D(N544), .CLK(clk), .Q(b_dout[10]) );
  DFFNX1_HVT \b_dout_reg[9]  ( .D(N545), .CLK(clk), .Q(b_dout[9]) );
  DFFNX1_HVT \b_dout_reg[8]  ( .D(N546), .CLK(clk), .Q(b_dout[8]) );
  DFFNX1_HVT \b_dout_reg[7]  ( .D(N547), .CLK(clk), .Q(b_dout[7]) );
  DFFNX1_HVT \b_dout_reg[6]  ( .D(N548), .CLK(clk), .Q(b_dout[6]) );
  DFFNX1_HVT \b_dout_reg[5]  ( .D(N549), .CLK(clk), .Q(b_dout[5]) );
  DFFNX1_HVT \b_dout_reg[4]  ( .D(N550), .CLK(clk), .Q(b_dout[4]) );
  DFFNX1_HVT \b_dout_reg[3]  ( .D(N551), .CLK(clk), .Q(b_dout[3]) );
  DFFNX1_HVT \b_dout_reg[2]  ( .D(N552), .CLK(clk), .Q(b_dout[2]) );
  DFFNX1_HVT \b_dout_reg[1]  ( .D(N553), .CLK(clk), .Q(b_dout[1]) );
  DFFNX1_HVT \b_dout_reg[0]  ( .D(N554), .CLK(clk), .Q(b_dout[0]) );
  DFFNX1_HVT \mem_reg[15][15]  ( .D(n1024), .CLK(clk), .Q(\mem[15][15] ) );
  DFFNX1_HVT \mem_reg[15][14]  ( .D(n1025), .CLK(clk), .Q(\mem[15][14] ) );
  DFFNX1_HVT \mem_reg[15][13]  ( .D(n1026), .CLK(clk), .Q(\mem[15][13] ) );
  DFFNX1_HVT \mem_reg[15][12]  ( .D(n1027), .CLK(clk), .Q(\mem[15][12] ) );
  DFFNX1_HVT \mem_reg[15][11]  ( .D(n1028), .CLK(clk), .Q(\mem[15][11] ) );
  DFFNX1_HVT \mem_reg[15][10]  ( .D(n1029), .CLK(clk), .Q(\mem[15][10] ) );
  DFFNX1_HVT \mem_reg[15][9]  ( .D(n1030), .CLK(clk), .Q(\mem[15][9] ) );
  DFFNX1_HVT \mem_reg[15][8]  ( .D(n1031), .CLK(clk), .Q(\mem[15][8] ) );
  DFFNX1_HVT \mem_reg[15][7]  ( .D(n1032), .CLK(clk), .Q(\mem[15][7] ) );
  DFFNX1_HVT \mem_reg[15][6]  ( .D(n1033), .CLK(clk), .Q(\mem[15][6] ) );
  DFFNX1_HVT \mem_reg[15][5]  ( .D(n1034), .CLK(clk), .Q(\mem[15][5] ) );
  DFFNX1_HVT \mem_reg[15][4]  ( .D(n1035), .CLK(clk), .Q(\mem[15][4] ) );
  DFFNX1_HVT \mem_reg[15][3]  ( .D(n1036), .CLK(clk), .Q(\mem[15][3] ) );
  DFFNX1_HVT \mem_reg[15][2]  ( .D(n1037), .CLK(clk), .Q(\mem[15][2] ) );
  DFFNX1_HVT \mem_reg[15][1]  ( .D(n1038), .CLK(clk), .Q(\mem[15][1] ) );
  DFFNX1_HVT \mem_reg[15][0]  ( .D(n1039), .CLK(clk), .Q(\mem[15][0] ) );
  DFFNX1_HVT \mem_reg[14][15]  ( .D(n1040), .CLK(clk), .Q(\mem[14][15] ) );
  DFFNX1_HVT \mem_reg[14][14]  ( .D(n1041), .CLK(clk), .Q(\mem[14][14] ) );
  DFFNX1_HVT \mem_reg[14][13]  ( .D(n1042), .CLK(clk), .Q(\mem[14][13] ) );
  DFFNX1_HVT \mem_reg[14][12]  ( .D(n1043), .CLK(clk), .Q(\mem[14][12] ) );
  DFFNX1_HVT \mem_reg[14][11]  ( .D(n1044), .CLK(clk), .Q(\mem[14][11] ) );
  DFFNX1_HVT \mem_reg[14][10]  ( .D(n1045), .CLK(clk), .Q(\mem[14][10] ) );
  DFFNX1_HVT \mem_reg[14][9]  ( .D(n1046), .CLK(clk), .Q(\mem[14][9] ) );
  DFFNX1_HVT \mem_reg[14][8]  ( .D(n1047), .CLK(clk), .Q(\mem[14][8] ) );
  DFFNX1_HVT \mem_reg[14][7]  ( .D(n1048), .CLK(clk), .Q(\mem[14][7] ) );
  DFFNX1_HVT \mem_reg[14][6]  ( .D(n1049), .CLK(clk), .Q(\mem[14][6] ) );
  DFFNX1_HVT \mem_reg[14][5]  ( .D(n1050), .CLK(clk), .Q(\mem[14][5] ) );
  DFFNX1_HVT \mem_reg[14][4]  ( .D(n1051), .CLK(clk), .Q(\mem[14][4] ) );
  DFFNX1_HVT \mem_reg[14][3]  ( .D(n1052), .CLK(clk), .Q(\mem[14][3] ) );
  DFFNX1_HVT \mem_reg[14][2]  ( .D(n1053), .CLK(clk), .Q(\mem[14][2] ) );
  DFFNX1_HVT \mem_reg[14][1]  ( .D(n1054), .CLK(clk), .Q(\mem[14][1] ) );
  DFFNX1_HVT \mem_reg[14][0]  ( .D(n1055), .CLK(clk), .Q(\mem[14][0] ) );
  DFFNX1_HVT \mem_reg[13][15]  ( .D(n1056), .CLK(clk), .Q(\mem[13][15] ) );
  DFFNX1_HVT \mem_reg[13][14]  ( .D(n1057), .CLK(clk), .Q(\mem[13][14] ) );
  DFFNX1_HVT \mem_reg[13][13]  ( .D(n1058), .CLK(clk), .Q(\mem[13][13] ) );
  DFFNX1_HVT \mem_reg[13][12]  ( .D(n1059), .CLK(clk), .Q(\mem[13][12] ) );
  DFFNX1_HVT \mem_reg[13][11]  ( .D(n1060), .CLK(clk), .Q(\mem[13][11] ) );
  DFFNX1_HVT \mem_reg[13][10]  ( .D(n1061), .CLK(clk), .Q(\mem[13][10] ) );
  DFFNX1_HVT \mem_reg[13][9]  ( .D(n1062), .CLK(clk), .Q(\mem[13][9] ) );
  DFFNX1_HVT \mem_reg[13][8]  ( .D(n1063), .CLK(clk), .Q(\mem[13][8] ) );
  DFFNX1_HVT \mem_reg[13][7]  ( .D(n1064), .CLK(clk), .Q(\mem[13][7] ) );
  DFFNX1_HVT \mem_reg[13][6]  ( .D(n1065), .CLK(clk), .Q(\mem[13][6] ) );
  DFFNX1_HVT \mem_reg[13][5]  ( .D(n1066), .CLK(clk), .Q(\mem[13][5] ) );
  DFFNX1_HVT \mem_reg[13][4]  ( .D(n1067), .CLK(clk), .Q(\mem[13][4] ) );
  DFFNX1_HVT \mem_reg[13][3]  ( .D(n1068), .CLK(clk), .Q(\mem[13][3] ) );
  DFFNX1_HVT \mem_reg[13][2]  ( .D(n1069), .CLK(clk), .Q(\mem[13][2] ) );
  DFFNX1_HVT \mem_reg[13][1]  ( .D(n1070), .CLK(clk), .Q(\mem[13][1] ) );
  DFFNX1_HVT \mem_reg[13][0]  ( .D(n1071), .CLK(clk), .Q(\mem[13][0] ) );
  DFFNX1_HVT \mem_reg[12][15]  ( .D(n1072), .CLK(clk), .Q(\mem[12][15] ) );
  DFFNX1_HVT \mem_reg[12][14]  ( .D(n1073), .CLK(clk), .Q(\mem[12][14] ) );
  DFFNX1_HVT \mem_reg[12][13]  ( .D(n1074), .CLK(clk), .Q(\mem[12][13] ) );
  DFFNX1_HVT \mem_reg[12][12]  ( .D(n1075), .CLK(clk), .Q(\mem[12][12] ) );
  DFFNX1_HVT \mem_reg[12][11]  ( .D(n1076), .CLK(clk), .Q(\mem[12][11] ) );
  DFFNX1_HVT \mem_reg[12][10]  ( .D(n1077), .CLK(clk), .Q(\mem[12][10] ) );
  DFFNX1_HVT \mem_reg[12][9]  ( .D(n1078), .CLK(clk), .Q(\mem[12][9] ) );
  DFFNX1_HVT \mem_reg[12][8]  ( .D(n1079), .CLK(clk), .Q(\mem[12][8] ) );
  DFFNX1_HVT \mem_reg[12][7]  ( .D(n1080), .CLK(clk), .Q(\mem[12][7] ) );
  DFFNX1_HVT \mem_reg[12][6]  ( .D(n1081), .CLK(clk), .Q(\mem[12][6] ) );
  DFFNX1_HVT \mem_reg[12][5]  ( .D(n1082), .CLK(clk), .Q(\mem[12][5] ) );
  DFFNX1_HVT \mem_reg[12][4]  ( .D(n1083), .CLK(clk), .Q(\mem[12][4] ) );
  DFFNX1_HVT \mem_reg[12][3]  ( .D(n1084), .CLK(clk), .Q(\mem[12][3] ) );
  DFFNX1_HVT \mem_reg[12][2]  ( .D(n1085), .CLK(clk), .Q(\mem[12][2] ) );
  DFFNX1_HVT \mem_reg[12][1]  ( .D(n1086), .CLK(clk), .Q(\mem[12][1] ) );
  DFFNX1_HVT \mem_reg[12][0]  ( .D(n1087), .CLK(clk), .Q(\mem[12][0] ) );
  DFFNX1_HVT \mem_reg[11][15]  ( .D(n1088), .CLK(clk), .Q(\mem[11][15] ) );
  DFFNX1_HVT \mem_reg[11][14]  ( .D(n1089), .CLK(clk), .Q(\mem[11][14] ) );
  DFFNX1_HVT \mem_reg[11][13]  ( .D(n1090), .CLK(clk), .Q(\mem[11][13] ) );
  DFFNX1_HVT \mem_reg[11][12]  ( .D(n1091), .CLK(clk), .Q(\mem[11][12] ) );
  DFFNX1_HVT \mem_reg[11][11]  ( .D(n1092), .CLK(clk), .Q(\mem[11][11] ) );
  DFFNX1_HVT \mem_reg[11][10]  ( .D(n1093), .CLK(clk), .Q(\mem[11][10] ) );
  DFFNX1_HVT \mem_reg[11][9]  ( .D(n1094), .CLK(clk), .Q(\mem[11][9] ) );
  DFFNX1_HVT \mem_reg[11][8]  ( .D(n1095), .CLK(clk), .Q(\mem[11][8] ) );
  DFFNX1_HVT \mem_reg[11][7]  ( .D(n1096), .CLK(clk), .Q(\mem[11][7] ) );
  DFFNX1_HVT \mem_reg[11][6]  ( .D(n1097), .CLK(clk), .Q(\mem[11][6] ) );
  DFFNX1_HVT \mem_reg[11][5]  ( .D(n1098), .CLK(clk), .Q(\mem[11][5] ) );
  DFFNX1_HVT \mem_reg[11][4]  ( .D(n1099), .CLK(clk), .Q(\mem[11][4] ) );
  DFFNX1_HVT \mem_reg[11][3]  ( .D(n1100), .CLK(clk), .Q(\mem[11][3] ) );
  DFFNX1_HVT \mem_reg[11][2]  ( .D(n1101), .CLK(clk), .Q(\mem[11][2] ) );
  DFFNX1_HVT \mem_reg[11][1]  ( .D(n1102), .CLK(clk), .Q(\mem[11][1] ) );
  DFFNX1_HVT \mem_reg[11][0]  ( .D(n1103), .CLK(clk), .Q(\mem[11][0] ) );
  DFFNX1_HVT \mem_reg[10][15]  ( .D(n1104), .CLK(clk), .Q(\mem[10][15] ) );
  DFFNX1_HVT \mem_reg[10][14]  ( .D(n1105), .CLK(clk), .Q(\mem[10][14] ) );
  DFFNX1_HVT \mem_reg[10][13]  ( .D(n1106), .CLK(clk), .Q(\mem[10][13] ) );
  DFFNX1_HVT \mem_reg[10][12]  ( .D(n1107), .CLK(clk), .Q(\mem[10][12] ) );
  DFFNX1_HVT \mem_reg[10][11]  ( .D(n1108), .CLK(clk), .Q(\mem[10][11] ) );
  DFFNX1_HVT \mem_reg[10][10]  ( .D(n1109), .CLK(clk), .Q(\mem[10][10] ) );
  DFFNX1_HVT \mem_reg[10][9]  ( .D(n1110), .CLK(clk), .Q(\mem[10][9] ) );
  DFFNX1_HVT \mem_reg[10][8]  ( .D(n1111), .CLK(clk), .Q(\mem[10][8] ) );
  DFFNX1_HVT \mem_reg[10][7]  ( .D(n1112), .CLK(clk), .Q(\mem[10][7] ) );
  DFFNX1_HVT \mem_reg[10][6]  ( .D(n1113), .CLK(clk), .Q(\mem[10][6] ) );
  DFFNX1_HVT \mem_reg[10][5]  ( .D(n1114), .CLK(clk), .Q(\mem[10][5] ) );
  DFFNX1_HVT \mem_reg[10][4]  ( .D(n1115), .CLK(clk), .Q(\mem[10][4] ) );
  DFFNX1_HVT \mem_reg[10][3]  ( .D(n1116), .CLK(clk), .Q(\mem[10][3] ) );
  DFFNX1_HVT \mem_reg[10][2]  ( .D(n1117), .CLK(clk), .Q(\mem[10][2] ) );
  DFFNX1_HVT \mem_reg[10][1]  ( .D(n1118), .CLK(clk), .Q(\mem[10][1] ) );
  DFFNX1_HVT \mem_reg[10][0]  ( .D(n1119), .CLK(clk), .Q(\mem[10][0] ) );
  DFFNX1_HVT \mem_reg[9][15]  ( .D(n1120), .CLK(clk), .Q(\mem[9][15] ) );
  DFFNX1_HVT \mem_reg[9][14]  ( .D(n1121), .CLK(clk), .Q(\mem[9][14] ) );
  DFFNX1_HVT \mem_reg[9][13]  ( .D(n1122), .CLK(clk), .Q(\mem[9][13] ) );
  DFFNX1_HVT \mem_reg[9][12]  ( .D(n1123), .CLK(clk), .Q(\mem[9][12] ) );
  DFFNX1_HVT \mem_reg[9][11]  ( .D(n1124), .CLK(clk), .Q(\mem[9][11] ) );
  DFFNX1_HVT \mem_reg[9][10]  ( .D(n1125), .CLK(clk), .Q(\mem[9][10] ) );
  DFFNX1_HVT \mem_reg[9][9]  ( .D(n1126), .CLK(clk), .Q(\mem[9][9] ) );
  DFFNX1_HVT \mem_reg[9][8]  ( .D(n1127), .CLK(clk), .Q(\mem[9][8] ) );
  DFFNX1_HVT \mem_reg[9][7]  ( .D(n1128), .CLK(clk), .Q(\mem[9][7] ) );
  DFFNX1_HVT \mem_reg[9][6]  ( .D(n1129), .CLK(clk), .Q(\mem[9][6] ) );
  DFFNX1_HVT \mem_reg[9][5]  ( .D(n1130), .CLK(clk), .Q(\mem[9][5] ) );
  DFFNX1_HVT \mem_reg[9][4]  ( .D(n1131), .CLK(clk), .Q(\mem[9][4] ) );
  DFFNX1_HVT \mem_reg[9][3]  ( .D(n1132), .CLK(clk), .Q(\mem[9][3] ) );
  DFFNX1_HVT \mem_reg[9][2]  ( .D(n1133), .CLK(clk), .Q(\mem[9][2] ) );
  DFFNX1_HVT \mem_reg[9][1]  ( .D(n1134), .CLK(clk), .Q(\mem[9][1] ) );
  DFFNX1_HVT \mem_reg[9][0]  ( .D(n1135), .CLK(clk), .Q(\mem[9][0] ) );
  DFFNX1_HVT \mem_reg[8][15]  ( .D(n1136), .CLK(clk), .Q(\mem[8][15] ) );
  DFFNX1_HVT \mem_reg[8][14]  ( .D(n1137), .CLK(clk), .Q(\mem[8][14] ) );
  DFFNX1_HVT \mem_reg[8][13]  ( .D(n1138), .CLK(clk), .Q(\mem[8][13] ) );
  DFFNX1_HVT \mem_reg[8][12]  ( .D(n1139), .CLK(clk), .Q(\mem[8][12] ) );
  DFFNX1_HVT \mem_reg[8][11]  ( .D(n1140), .CLK(clk), .Q(\mem[8][11] ) );
  DFFNX1_HVT \mem_reg[8][10]  ( .D(n1141), .CLK(clk), .Q(\mem[8][10] ) );
  DFFNX1_HVT \mem_reg[8][9]  ( .D(n1142), .CLK(clk), .Q(\mem[8][9] ) );
  DFFNX1_HVT \mem_reg[8][8]  ( .D(n1143), .CLK(clk), .Q(\mem[8][8] ) );
  DFFNX1_HVT \mem_reg[8][7]  ( .D(n1144), .CLK(clk), .Q(\mem[8][7] ) );
  DFFNX1_HVT \mem_reg[8][6]  ( .D(n1145), .CLK(clk), .Q(\mem[8][6] ) );
  DFFNX1_HVT \mem_reg[8][5]  ( .D(n1146), .CLK(clk), .Q(\mem[8][5] ) );
  DFFNX1_HVT \mem_reg[8][4]  ( .D(n1147), .CLK(clk), .Q(\mem[8][4] ) );
  DFFNX1_HVT \mem_reg[8][3]  ( .D(n1148), .CLK(clk), .Q(\mem[8][3] ) );
  DFFNX1_HVT \mem_reg[8][2]  ( .D(n1149), .CLK(clk), .Q(\mem[8][2] ) );
  DFFNX1_HVT \mem_reg[8][1]  ( .D(n1150), .CLK(clk), .Q(\mem[8][1] ) );
  DFFNX1_HVT \mem_reg[8][0]  ( .D(n1151), .CLK(clk), .Q(\mem[8][0] ) );
  DFFNX1_HVT \mem_reg[7][15]  ( .D(n1152), .CLK(clk), .Q(\mem[7][15] ) );
  DFFNX1_HVT \mem_reg[7][14]  ( .D(n1153), .CLK(clk), .Q(\mem[7][14] ) );
  DFFNX1_HVT \mem_reg[7][13]  ( .D(n1154), .CLK(clk), .Q(\mem[7][13] ) );
  DFFNX1_HVT \mem_reg[7][12]  ( .D(n1155), .CLK(clk), .Q(\mem[7][12] ) );
  DFFNX1_HVT \mem_reg[7][11]  ( .D(n1156), .CLK(clk), .Q(\mem[7][11] ) );
  DFFNX1_HVT \mem_reg[7][10]  ( .D(n1157), .CLK(clk), .Q(\mem[7][10] ) );
  DFFNX1_HVT \mem_reg[7][9]  ( .D(n1158), .CLK(clk), .Q(\mem[7][9] ) );
  DFFNX1_HVT \mem_reg[7][8]  ( .D(n1159), .CLK(clk), .Q(\mem[7][8] ) );
  DFFNX1_HVT \mem_reg[7][7]  ( .D(n1160), .CLK(clk), .Q(\mem[7][7] ) );
  DFFNX1_HVT \mem_reg[7][6]  ( .D(n1161), .CLK(clk), .Q(\mem[7][6] ) );
  DFFNX1_HVT \mem_reg[7][5]  ( .D(n1162), .CLK(clk), .Q(\mem[7][5] ) );
  DFFNX1_HVT \mem_reg[7][4]  ( .D(n1163), .CLK(clk), .Q(\mem[7][4] ) );
  DFFNX1_HVT \mem_reg[7][3]  ( .D(n1164), .CLK(clk), .Q(\mem[7][3] ) );
  DFFNX1_HVT \mem_reg[7][2]  ( .D(n1165), .CLK(clk), .Q(\mem[7][2] ) );
  DFFNX1_HVT \mem_reg[7][1]  ( .D(n1166), .CLK(clk), .Q(\mem[7][1] ) );
  DFFNX1_HVT \mem_reg[7][0]  ( .D(n1167), .CLK(clk), .Q(\mem[7][0] ) );
  DFFNX1_HVT \mem_reg[6][15]  ( .D(n1168), .CLK(clk), .Q(\mem[6][15] ) );
  DFFNX1_HVT \mem_reg[6][14]  ( .D(n1169), .CLK(clk), .Q(\mem[6][14] ) );
  DFFNX1_HVT \mem_reg[6][13]  ( .D(n1170), .CLK(clk), .Q(\mem[6][13] ) );
  DFFNX1_HVT \mem_reg[6][12]  ( .D(n1171), .CLK(clk), .Q(\mem[6][12] ) );
  DFFNX1_HVT \mem_reg[6][11]  ( .D(n1172), .CLK(clk), .Q(\mem[6][11] ) );
  DFFNX1_HVT \mem_reg[6][10]  ( .D(n1173), .CLK(clk), .Q(\mem[6][10] ) );
  DFFNX1_HVT \mem_reg[6][9]  ( .D(n1174), .CLK(clk), .Q(\mem[6][9] ) );
  DFFNX1_HVT \mem_reg[6][8]  ( .D(n1175), .CLK(clk), .Q(\mem[6][8] ) );
  DFFNX1_HVT \mem_reg[6][7]  ( .D(n1176), .CLK(clk), .Q(\mem[6][7] ) );
  DFFNX1_HVT \mem_reg[6][6]  ( .D(n1177), .CLK(clk), .Q(\mem[6][6] ) );
  DFFNX1_HVT \mem_reg[6][5]  ( .D(n1178), .CLK(clk), .Q(\mem[6][5] ) );
  DFFNX1_HVT \mem_reg[6][4]  ( .D(n1179), .CLK(clk), .Q(\mem[6][4] ) );
  DFFNX1_HVT \mem_reg[6][3]  ( .D(n1180), .CLK(clk), .Q(\mem[6][3] ) );
  DFFNX1_HVT \mem_reg[6][2]  ( .D(n1181), .CLK(clk), .Q(\mem[6][2] ) );
  DFFNX1_HVT \mem_reg[6][1]  ( .D(n1182), .CLK(clk), .Q(\mem[6][1] ) );
  DFFNX1_HVT \mem_reg[6][0]  ( .D(n1183), .CLK(clk), .Q(\mem[6][0] ) );
  DFFNX1_HVT \mem_reg[5][15]  ( .D(n1184), .CLK(clk), .Q(\mem[5][15] ) );
  DFFNX1_HVT \mem_reg[5][14]  ( .D(n1185), .CLK(clk), .Q(\mem[5][14] ) );
  DFFNX1_HVT \mem_reg[5][13]  ( .D(n1186), .CLK(clk), .Q(\mem[5][13] ) );
  DFFNX1_HVT \mem_reg[5][12]  ( .D(n1187), .CLK(clk), .Q(\mem[5][12] ) );
  DFFNX1_HVT \mem_reg[5][11]  ( .D(n1188), .CLK(clk), .Q(\mem[5][11] ) );
  DFFNX1_HVT \mem_reg[5][10]  ( .D(n1189), .CLK(clk), .Q(\mem[5][10] ) );
  DFFNX1_HVT \mem_reg[5][9]  ( .D(n1190), .CLK(clk), .Q(\mem[5][9] ) );
  DFFNX1_HVT \mem_reg[5][8]  ( .D(n1191), .CLK(clk), .Q(\mem[5][8] ) );
  DFFNX1_HVT \mem_reg[5][7]  ( .D(n1192), .CLK(clk), .Q(\mem[5][7] ) );
  DFFNX1_HVT \mem_reg[5][6]  ( .D(n1193), .CLK(clk), .Q(\mem[5][6] ) );
  DFFNX1_HVT \mem_reg[5][5]  ( .D(n1194), .CLK(clk), .Q(\mem[5][5] ) );
  DFFNX1_HVT \mem_reg[5][4]  ( .D(n1195), .CLK(clk), .Q(\mem[5][4] ) );
  DFFNX1_HVT \mem_reg[5][3]  ( .D(n1196), .CLK(clk), .Q(\mem[5][3] ) );
  DFFNX1_HVT \mem_reg[5][2]  ( .D(n1197), .CLK(clk), .Q(\mem[5][2] ) );
  DFFNX1_HVT \mem_reg[5][1]  ( .D(n1198), .CLK(clk), .Q(\mem[5][1] ) );
  DFFNX1_HVT \mem_reg[5][0]  ( .D(n1199), .CLK(clk), .Q(\mem[5][0] ) );
  DFFNX1_HVT \mem_reg[4][15]  ( .D(n1200), .CLK(clk), .Q(\mem[4][15] ) );
  DFFNX1_HVT \mem_reg[4][14]  ( .D(n1201), .CLK(clk), .Q(\mem[4][14] ) );
  DFFNX1_HVT \mem_reg[4][13]  ( .D(n1202), .CLK(clk), .Q(\mem[4][13] ) );
  DFFNX1_HVT \mem_reg[4][12]  ( .D(n1203), .CLK(clk), .Q(\mem[4][12] ) );
  DFFNX1_HVT \mem_reg[4][11]  ( .D(n1204), .CLK(clk), .Q(\mem[4][11] ) );
  DFFNX1_HVT \mem_reg[4][10]  ( .D(n1205), .CLK(clk), .Q(\mem[4][10] ) );
  DFFNX1_HVT \mem_reg[4][9]  ( .D(n1206), .CLK(clk), .Q(\mem[4][9] ) );
  DFFNX1_HVT \mem_reg[4][8]  ( .D(n1207), .CLK(clk), .Q(\mem[4][8] ) );
  DFFNX1_HVT \mem_reg[4][7]  ( .D(n1208), .CLK(clk), .Q(\mem[4][7] ) );
  DFFNX1_HVT \mem_reg[4][6]  ( .D(n1209), .CLK(clk), .Q(\mem[4][6] ) );
  DFFNX1_HVT \mem_reg[4][5]  ( .D(n1210), .CLK(clk), .Q(\mem[4][5] ) );
  DFFNX1_HVT \mem_reg[4][4]  ( .D(n1211), .CLK(clk), .Q(\mem[4][4] ) );
  DFFNX1_HVT \mem_reg[4][3]  ( .D(n1212), .CLK(clk), .Q(\mem[4][3] ) );
  DFFNX1_HVT \mem_reg[4][2]  ( .D(n1213), .CLK(clk), .Q(\mem[4][2] ) );
  DFFNX1_HVT \mem_reg[4][1]  ( .D(n1214), .CLK(clk), .Q(\mem[4][1] ) );
  DFFNX1_HVT \mem_reg[4][0]  ( .D(n1215), .CLK(clk), .Q(\mem[4][0] ) );
  DFFNX1_HVT \mem_reg[3][15]  ( .D(n1216), .CLK(clk), .Q(\mem[3][15] ) );
  DFFNX1_HVT \mem_reg[3][14]  ( .D(n1217), .CLK(clk), .Q(\mem[3][14] ) );
  DFFNX1_HVT \mem_reg[3][13]  ( .D(n1218), .CLK(clk), .Q(\mem[3][13] ) );
  DFFNX1_HVT \mem_reg[3][12]  ( .D(n1219), .CLK(clk), .Q(\mem[3][12] ) );
  DFFNX1_HVT \mem_reg[3][11]  ( .D(n1220), .CLK(clk), .Q(\mem[3][11] ) );
  DFFNX1_HVT \mem_reg[3][10]  ( .D(n1221), .CLK(clk), .Q(\mem[3][10] ) );
  DFFNX1_HVT \mem_reg[3][9]  ( .D(n1222), .CLK(clk), .Q(\mem[3][9] ) );
  DFFNX1_HVT \mem_reg[3][8]  ( .D(n1223), .CLK(clk), .Q(\mem[3][8] ) );
  DFFNX1_HVT \mem_reg[3][7]  ( .D(n1224), .CLK(clk), .Q(\mem[3][7] ) );
  DFFNX1_HVT \mem_reg[3][6]  ( .D(n1225), .CLK(clk), .Q(\mem[3][6] ) );
  DFFNX1_HVT \mem_reg[3][5]  ( .D(n1226), .CLK(clk), .Q(\mem[3][5] ) );
  DFFNX1_HVT \mem_reg[3][4]  ( .D(n1227), .CLK(clk), .Q(\mem[3][4] ) );
  DFFNX1_HVT \mem_reg[3][3]  ( .D(n1228), .CLK(clk), .Q(\mem[3][3] ) );
  DFFNX1_HVT \mem_reg[3][2]  ( .D(n1229), .CLK(clk), .Q(\mem[3][2] ) );
  DFFNX1_HVT \mem_reg[3][1]  ( .D(n1230), .CLK(clk), .Q(\mem[3][1] ) );
  DFFNX1_HVT \mem_reg[3][0]  ( .D(n1231), .CLK(clk), .Q(\mem[3][0] ) );
  DFFNX1_HVT \mem_reg[2][15]  ( .D(n1232), .CLK(clk), .Q(\mem[2][15] ) );
  DFFNX1_HVT \mem_reg[2][14]  ( .D(n1233), .CLK(clk), .Q(\mem[2][14] ) );
  DFFNX1_HVT \mem_reg[2][13]  ( .D(n1234), .CLK(clk), .Q(\mem[2][13] ) );
  DFFNX1_HVT \mem_reg[2][12]  ( .D(n1235), .CLK(clk), .Q(\mem[2][12] ) );
  DFFNX1_HVT \mem_reg[2][11]  ( .D(n1236), .CLK(clk), .Q(\mem[2][11] ) );
  DFFNX1_HVT \mem_reg[2][10]  ( .D(n1237), .CLK(clk), .Q(\mem[2][10] ) );
  DFFNX1_HVT \mem_reg[2][9]  ( .D(n1238), .CLK(clk), .Q(\mem[2][9] ) );
  DFFNX1_HVT \mem_reg[2][8]  ( .D(n1239), .CLK(clk), .Q(\mem[2][8] ) );
  DFFNX1_HVT \mem_reg[2][7]  ( .D(n1240), .CLK(clk), .Q(\mem[2][7] ) );
  DFFNX1_HVT \mem_reg[2][6]  ( .D(n1241), .CLK(clk), .Q(\mem[2][6] ) );
  DFFNX1_HVT \mem_reg[2][5]  ( .D(n1242), .CLK(clk), .Q(\mem[2][5] ) );
  DFFNX1_HVT \mem_reg[2][4]  ( .D(n1243), .CLK(clk), .Q(\mem[2][4] ) );
  DFFNX1_HVT \mem_reg[2][3]  ( .D(n1244), .CLK(clk), .Q(\mem[2][3] ) );
  DFFNX1_HVT \mem_reg[2][2]  ( .D(n1245), .CLK(clk), .Q(\mem[2][2] ) );
  DFFNX1_HVT \mem_reg[2][1]  ( .D(n1246), .CLK(clk), .Q(\mem[2][1] ) );
  DFFNX1_HVT \mem_reg[2][0]  ( .D(n1247), .CLK(clk), .Q(\mem[2][0] ) );
  DFFNX1_HVT \mem_reg[1][15]  ( .D(n1248), .CLK(clk), .Q(\mem[1][15] ) );
  DFFNX1_HVT \mem_reg[1][14]  ( .D(n1249), .CLK(clk), .Q(\mem[1][14] ) );
  DFFNX1_HVT \mem_reg[1][13]  ( .D(n1250), .CLK(clk), .Q(\mem[1][13] ) );
  DFFNX1_HVT \mem_reg[1][12]  ( .D(n1251), .CLK(clk), .Q(\mem[1][12] ) );
  DFFNX1_HVT \mem_reg[1][11]  ( .D(n1252), .CLK(clk), .Q(\mem[1][11] ) );
  DFFNX1_HVT \mem_reg[1][10]  ( .D(n1253), .CLK(clk), .Q(\mem[1][10] ) );
  DFFNX1_HVT \mem_reg[1][9]  ( .D(n1254), .CLK(clk), .Q(\mem[1][9] ) );
  DFFNX1_HVT \mem_reg[1][8]  ( .D(n1255), .CLK(clk), .Q(\mem[1][8] ) );
  DFFNX1_HVT \mem_reg[1][7]  ( .D(n1256), .CLK(clk), .Q(\mem[1][7] ) );
  DFFNX1_HVT \mem_reg[1][6]  ( .D(n1257), .CLK(clk), .Q(\mem[1][6] ) );
  DFFNX1_HVT \mem_reg[1][5]  ( .D(n1258), .CLK(clk), .Q(\mem[1][5] ) );
  DFFNX1_HVT \mem_reg[1][4]  ( .D(n1259), .CLK(clk), .Q(\mem[1][4] ) );
  DFFNX1_HVT \mem_reg[1][3]  ( .D(n1260), .CLK(clk), .Q(\mem[1][3] ) );
  DFFNX1_HVT \mem_reg[1][2]  ( .D(n1261), .CLK(clk), .Q(\mem[1][2] ) );
  DFFNX1_HVT \mem_reg[1][1]  ( .D(n1262), .CLK(clk), .Q(\mem[1][1] ) );
  DFFNX1_HVT \mem_reg[1][0]  ( .D(n1263), .CLK(clk), .Q(\mem[1][0] ) );
  DFFNX1_HVT \mem_reg[0][15]  ( .D(n1264), .CLK(clk), .Q(\mem[0][15] ) );
  DFFNX1_HVT \mem_reg[0][14]  ( .D(n1265), .CLK(clk), .Q(\mem[0][14] ) );
  DFFNX1_HVT \mem_reg[0][13]  ( .D(n1266), .CLK(clk), .Q(\mem[0][13] ) );
  DFFNX1_HVT \mem_reg[0][12]  ( .D(n1267), .CLK(clk), .Q(\mem[0][12] ) );
  DFFNX1_HVT \mem_reg[0][11]  ( .D(n1268), .CLK(clk), .Q(\mem[0][11] ) );
  DFFNX1_HVT \mem_reg[0][10]  ( .D(n1269), .CLK(clk), .Q(\mem[0][10] ) );
  DFFNX1_HVT \mem_reg[0][9]  ( .D(n1270), .CLK(clk), .Q(\mem[0][9] ) );
  DFFNX1_HVT \mem_reg[0][8]  ( .D(n1271), .CLK(clk), .Q(\mem[0][8] ) );
  DFFNX1_HVT \mem_reg[0][7]  ( .D(n1272), .CLK(clk), .Q(\mem[0][7] ) );
  DFFNX1_HVT \mem_reg[0][6]  ( .D(n1273), .CLK(clk), .Q(\mem[0][6] ) );
  DFFNX1_HVT \mem_reg[0][5]  ( .D(n1274), .CLK(clk), .Q(\mem[0][5] ) );
  DFFNX1_HVT \mem_reg[0][4]  ( .D(n1275), .CLK(clk), .Q(\mem[0][4] ) );
  DFFNX1_HVT \mem_reg[0][3]  ( .D(n1276), .CLK(clk), .Q(\mem[0][3] ) );
  DFFNX1_HVT \mem_reg[0][2]  ( .D(n1277), .CLK(clk), .Q(\mem[0][2] ) );
  DFFNX1_HVT \mem_reg[0][1]  ( .D(n1278), .CLK(clk), .Q(\mem[0][1] ) );
  DFFNX1_HVT \mem_reg[0][0]  ( .D(n1279), .CLK(clk), .Q(\mem[0][0] ) );
  AO22X1_HVT U268 ( .A1(n1580), .A2(n189), .A3(\mem[0][0] ), .A4(n893), .Y(
        n1279) );
  AO21X1_HVT U269 ( .A1(n1579), .A2(n150), .A3(n165), .Y(n1580) );
  AO22X1_HVT U270 ( .A1(n1577), .A2(n189), .A3(\mem[0][1] ), .A4(n892), .Y(
        n1278) );
  AO21X1_HVT U271 ( .A1(n1576), .A2(n152), .A3(n166), .Y(n1577) );
  AO22X1_HVT U272 ( .A1(n1575), .A2(n189), .A3(\mem[0][2] ), .A4(n891), .Y(
        n1277) );
  AO21X1_HVT U273 ( .A1(n1574), .A2(n151), .A3(n183), .Y(n1575) );
  AO22X1_HVT U274 ( .A1(n1573), .A2(n189), .A3(\mem[0][3] ), .A4(n890), .Y(
        n1276) );
  AO21X1_HVT U275 ( .A1(n1572), .A2(n150), .A3(n166), .Y(n1573) );
  AO22X1_HVT U276 ( .A1(n1571), .A2(n189), .A3(\mem[0][4] ), .A4(n889), .Y(
        n1275) );
  AO21X1_HVT U277 ( .A1(n1570), .A2(n152), .A3(n166), .Y(n1571) );
  AO22X1_HVT U278 ( .A1(n1569), .A2(n189), .A3(\mem[0][5] ), .A4(n888), .Y(
        n1274) );
  AO21X1_HVT U279 ( .A1(n1568), .A2(n151), .A3(n166), .Y(n1569) );
  AO22X1_HVT U280 ( .A1(n1567), .A2(n189), .A3(\mem[0][6] ), .A4(n887), .Y(
        n1273) );
  AO21X1_HVT U281 ( .A1(n1566), .A2(n150), .A3(n166), .Y(n1567) );
  AO22X1_HVT U282 ( .A1(n1565), .A2(n189), .A3(\mem[0][7] ), .A4(n886), .Y(
        n1272) );
  AO21X1_HVT U283 ( .A1(n1564), .A2(n152), .A3(n166), .Y(n1565) );
  AO22X1_HVT U284 ( .A1(n1563), .A2(n189), .A3(\mem[0][8] ), .A4(n885), .Y(
        n1271) );
  AO21X1_HVT U285 ( .A1(n1562), .A2(n151), .A3(n166), .Y(n1563) );
  AO22X1_HVT U286 ( .A1(n1561), .A2(n189), .A3(\mem[0][9] ), .A4(n884), .Y(
        n1270) );
  AO21X1_HVT U287 ( .A1(n1560), .A2(n150), .A3(n167), .Y(n1561) );
  AO22X1_HVT U288 ( .A1(n1559), .A2(n189), .A3(\mem[0][10] ), .A4(n883), .Y(
        n1269) );
  AO21X1_HVT U289 ( .A1(n1558), .A2(n152), .A3(n167), .Y(n1559) );
  AO22X1_HVT U290 ( .A1(n1557), .A2(n189), .A3(\mem[0][11] ), .A4(n882), .Y(
        n1268) );
  AO21X1_HVT U291 ( .A1(n1556), .A2(n151), .A3(n167), .Y(n1557) );
  AO22X1_HVT U292 ( .A1(n1555), .A2(n190), .A3(\mem[0][12] ), .A4(n881), .Y(
        n1267) );
  AO21X1_HVT U293 ( .A1(n1554), .A2(n150), .A3(n167), .Y(n1555) );
  AO22X1_HVT U294 ( .A1(n1553), .A2(n190), .A3(\mem[0][13] ), .A4(n880), .Y(
        n1266) );
  AO21X1_HVT U295 ( .A1(n1552), .A2(n152), .A3(n167), .Y(n1553) );
  AO22X1_HVT U296 ( .A1(n1551), .A2(n190), .A3(\mem[0][14] ), .A4(n879), .Y(
        n1265) );
  AO21X1_HVT U297 ( .A1(n1550), .A2(n151), .A3(n167), .Y(n1551) );
  AO22X1_HVT U298 ( .A1(n1549), .A2(n190), .A3(\mem[0][15] ), .A4(n878), .Y(
        n1264) );
  AO21X1_HVT U299 ( .A1(n1548), .A2(n150), .A3(n167), .Y(n1549) );
  AND3X1_HVT U300 ( .A1(n1547), .A2(n163), .A3(n1546), .Y(n1578) );
  AO22X1_HVT U301 ( .A1(n1545), .A2(n190), .A3(\mem[1][0] ), .A4(n877), .Y(
        n1263) );
  AO21X1_HVT U302 ( .A1(n149), .A2(n1579), .A3(n167), .Y(n1545) );
  AO22X1_HVT U303 ( .A1(n1544), .A2(n190), .A3(\mem[1][1] ), .A4(n876), .Y(
        n1262) );
  AO21X1_HVT U304 ( .A1(n149), .A2(n1576), .A3(n167), .Y(n1544) );
  AO22X1_HVT U305 ( .A1(n1543), .A2(n190), .A3(\mem[1][2] ), .A4(n875), .Y(
        n1261) );
  AO21X1_HVT U306 ( .A1(n149), .A2(n1574), .A3(n167), .Y(n1543) );
  AO22X1_HVT U307 ( .A1(n1542), .A2(n190), .A3(\mem[1][3] ), .A4(n874), .Y(
        n1260) );
  AO21X1_HVT U308 ( .A1(n149), .A2(n1572), .A3(n167), .Y(n1542) );
  AO22X1_HVT U309 ( .A1(n1541), .A2(n190), .A3(\mem[1][4] ), .A4(n873), .Y(
        n1259) );
  AO21X1_HVT U310 ( .A1(n149), .A2(n1570), .A3(n167), .Y(n1541) );
  AO22X1_HVT U311 ( .A1(n1540), .A2(n190), .A3(\mem[1][5] ), .A4(n872), .Y(
        n1258) );
  AO21X1_HVT U312 ( .A1(n149), .A2(n1568), .A3(n167), .Y(n1540) );
  AO22X1_HVT U313 ( .A1(n1539), .A2(n190), .A3(\mem[1][6] ), .A4(n871), .Y(
        n1257) );
  AO21X1_HVT U314 ( .A1(n149), .A2(n1566), .A3(n167), .Y(n1539) );
  AO22X1_HVT U315 ( .A1(n1538), .A2(n190), .A3(\mem[1][7] ), .A4(n870), .Y(
        n1256) );
  AO21X1_HVT U316 ( .A1(n149), .A2(n1564), .A3(n167), .Y(n1538) );
  AO22X1_HVT U317 ( .A1(n1537), .A2(n191), .A3(\mem[1][8] ), .A4(n869), .Y(
        n1255) );
  AO21X1_HVT U318 ( .A1(n148), .A2(n1562), .A3(n168), .Y(n1537) );
  AO22X1_HVT U319 ( .A1(n1536), .A2(n191), .A3(\mem[1][9] ), .A4(n868), .Y(
        n1254) );
  AO21X1_HVT U320 ( .A1(n148), .A2(n1560), .A3(n168), .Y(n1536) );
  AO22X1_HVT U321 ( .A1(n1535), .A2(n191), .A3(\mem[1][10] ), .A4(n867), .Y(
        n1253) );
  AO21X1_HVT U322 ( .A1(n148), .A2(n1558), .A3(n168), .Y(n1535) );
  AO22X1_HVT U323 ( .A1(n1534), .A2(n191), .A3(\mem[1][11] ), .A4(n866), .Y(
        n1252) );
  AO21X1_HVT U324 ( .A1(n148), .A2(n1556), .A3(n168), .Y(n1534) );
  AO22X1_HVT U325 ( .A1(n1533), .A2(n191), .A3(\mem[1][12] ), .A4(n865), .Y(
        n1251) );
  AO21X1_HVT U326 ( .A1(n148), .A2(n1554), .A3(n168), .Y(n1533) );
  AO22X1_HVT U327 ( .A1(n1532), .A2(n191), .A3(\mem[1][13] ), .A4(n864), .Y(
        n1250) );
  AO21X1_HVT U328 ( .A1(n148), .A2(n1552), .A3(n168), .Y(n1532) );
  AO22X1_HVT U329 ( .A1(n1531), .A2(n191), .A3(\mem[1][14] ), .A4(n863), .Y(
        n1249) );
  AO21X1_HVT U330 ( .A1(n148), .A2(n1550), .A3(n168), .Y(n1531) );
  AO22X1_HVT U331 ( .A1(n1530), .A2(n191), .A3(\mem[1][15] ), .A4(n862), .Y(
        n1248) );
  AO21X1_HVT U332 ( .A1(n148), .A2(n1548), .A3(n168), .Y(n1530) );
  AO22X1_HVT U334 ( .A1(n1528), .A2(n191), .A3(\mem[2][0] ), .A4(n861), .Y(
        n1247) );
  AO21X1_HVT U335 ( .A1(n5), .A2(n1579), .A3(n168), .Y(n1528) );
  AO22X1_HVT U336 ( .A1(n1527), .A2(n191), .A3(\mem[2][1] ), .A4(n860), .Y(
        n1246) );
  AO21X1_HVT U337 ( .A1(n146), .A2(n1576), .A3(n168), .Y(n1527) );
  AO22X1_HVT U338 ( .A1(n1526), .A2(n191), .A3(\mem[2][2] ), .A4(n859), .Y(
        n1245) );
  AO21X1_HVT U339 ( .A1(n5), .A2(n1574), .A3(n168), .Y(n1526) );
  AO22X1_HVT U340 ( .A1(n1525), .A2(n191), .A3(\mem[2][3] ), .A4(n858), .Y(
        n1244) );
  AO21X1_HVT U341 ( .A1(n146), .A2(n1572), .A3(n168), .Y(n1525) );
  AO22X1_HVT U342 ( .A1(n1524), .A2(n192), .A3(\mem[2][4] ), .A4(n857), .Y(
        n1243) );
  AO21X1_HVT U343 ( .A1(n5), .A2(n1570), .A3(n168), .Y(n1524) );
  AO22X1_HVT U344 ( .A1(n1523), .A2(n192), .A3(\mem[2][5] ), .A4(n856), .Y(
        n1242) );
  AO21X1_HVT U345 ( .A1(n146), .A2(n1568), .A3(n168), .Y(n1523) );
  AO22X1_HVT U346 ( .A1(n1522), .A2(n192), .A3(\mem[2][6] ), .A4(n855), .Y(
        n1241) );
  AO21X1_HVT U347 ( .A1(n5), .A2(n1566), .A3(n168), .Y(n1522) );
  AO22X1_HVT U348 ( .A1(n1521), .A2(n192), .A3(\mem[2][7] ), .A4(n854), .Y(
        n1240) );
  AO21X1_HVT U349 ( .A1(n146), .A2(n1564), .A3(n169), .Y(n1521) );
  AO22X1_HVT U350 ( .A1(n1520), .A2(n192), .A3(\mem[2][8] ), .A4(n853), .Y(
        n1239) );
  AO21X1_HVT U351 ( .A1(n147), .A2(n1562), .A3(n169), .Y(n1520) );
  AO22X1_HVT U352 ( .A1(n1519), .A2(n192), .A3(\mem[2][9] ), .A4(n852), .Y(
        n1238) );
  AO21X1_HVT U353 ( .A1(n147), .A2(n1560), .A3(n169), .Y(n1519) );
  AO22X1_HVT U354 ( .A1(n1518), .A2(n192), .A3(\mem[2][10] ), .A4(n851), .Y(
        n1237) );
  AO21X1_HVT U355 ( .A1(n147), .A2(n1558), .A3(n169), .Y(n1518) );
  AO22X1_HVT U356 ( .A1(n1517), .A2(n192), .A3(\mem[2][11] ), .A4(n850), .Y(
        n1236) );
  AO21X1_HVT U357 ( .A1(n147), .A2(n1556), .A3(n169), .Y(n1517) );
  AO22X1_HVT U358 ( .A1(n1516), .A2(n192), .A3(\mem[2][12] ), .A4(n849), .Y(
        n1235) );
  AO21X1_HVT U359 ( .A1(n147), .A2(n1554), .A3(n169), .Y(n1516) );
  AO22X1_HVT U360 ( .A1(n1515), .A2(n192), .A3(\mem[2][13] ), .A4(n848), .Y(
        n1234) );
  AO21X1_HVT U361 ( .A1(n147), .A2(n1552), .A3(n169), .Y(n1515) );
  AO22X1_HVT U362 ( .A1(n1514), .A2(n192), .A3(\mem[2][14] ), .A4(n847), .Y(
        n1233) );
  AO21X1_HVT U363 ( .A1(n5), .A2(n1550), .A3(n169), .Y(n1514) );
  AO22X1_HVT U364 ( .A1(n1513), .A2(n192), .A3(\mem[2][15] ), .A4(n846), .Y(
        n1232) );
  AO21X1_HVT U365 ( .A1(n146), .A2(n1548), .A3(n169), .Y(n1513) );
  AO22X1_HVT U367 ( .A1(n1511), .A2(n188), .A3(\mem[3][0] ), .A4(n845), .Y(
        n1231) );
  AO21X1_HVT U368 ( .A1(n145), .A2(n1579), .A3(n169), .Y(n1511) );
  AO22X1_HVT U369 ( .A1(n1510), .A2(n208), .A3(\mem[3][1] ), .A4(n844), .Y(
        n1230) );
  AO21X1_HVT U370 ( .A1(n145), .A2(n1576), .A3(n169), .Y(n1510) );
  AO22X1_HVT U371 ( .A1(n1509), .A2(n184), .A3(\mem[3][2] ), .A4(n843), .Y(
        n1229) );
  AO21X1_HVT U372 ( .A1(n145), .A2(n1574), .A3(n169), .Y(n1509) );
  AO22X1_HVT U373 ( .A1(n1508), .A2(n185), .A3(\mem[3][3] ), .A4(n842), .Y(
        n1228) );
  AO21X1_HVT U374 ( .A1(n145), .A2(n1572), .A3(n169), .Y(n1508) );
  AO22X1_HVT U375 ( .A1(n1507), .A2(n186), .A3(\mem[3][4] ), .A4(n841), .Y(
        n1227) );
  AO21X1_HVT U376 ( .A1(n145), .A2(n1570), .A3(n169), .Y(n1507) );
  AO22X1_HVT U377 ( .A1(n1506), .A2(n188), .A3(\mem[3][5] ), .A4(n840), .Y(
        n1226) );
  AO21X1_HVT U378 ( .A1(n145), .A2(n1568), .A3(n169), .Y(n1506) );
  AO22X1_HVT U379 ( .A1(n1505), .A2(n208), .A3(\mem[3][6] ), .A4(n839), .Y(
        n1225) );
  AO21X1_HVT U380 ( .A1(n145), .A2(n1566), .A3(n170), .Y(n1505) );
  AO22X1_HVT U381 ( .A1(n1504), .A2(n188), .A3(\mem[3][7] ), .A4(n838), .Y(
        n1224) );
  AO21X1_HVT U382 ( .A1(n145), .A2(n1564), .A3(n170), .Y(n1504) );
  AO22X1_HVT U383 ( .A1(n1503), .A2(n208), .A3(\mem[3][8] ), .A4(n837), .Y(
        n1223) );
  AO21X1_HVT U384 ( .A1(n144), .A2(n1562), .A3(n170), .Y(n1503) );
  AO22X1_HVT U385 ( .A1(n1502), .A2(n188), .A3(\mem[3][9] ), .A4(n836), .Y(
        n1222) );
  AO21X1_HVT U386 ( .A1(n144), .A2(n1560), .A3(n170), .Y(n1502) );
  AO22X1_HVT U387 ( .A1(n1501), .A2(n208), .A3(\mem[3][10] ), .A4(n835), .Y(
        n1221) );
  AO21X1_HVT U388 ( .A1(n144), .A2(n1558), .A3(n170), .Y(n1501) );
  AO22X1_HVT U389 ( .A1(n1500), .A2(n208), .A3(\mem[3][11] ), .A4(n834), .Y(
        n1220) );
  AO21X1_HVT U390 ( .A1(n144), .A2(n1556), .A3(n170), .Y(n1500) );
  AO22X1_HVT U391 ( .A1(n1499), .A2(n193), .A3(\mem[3][12] ), .A4(n833), .Y(
        n1219) );
  AO21X1_HVT U392 ( .A1(n144), .A2(n1554), .A3(n170), .Y(n1499) );
  AO22X1_HVT U393 ( .A1(n1498), .A2(n193), .A3(\mem[3][13] ), .A4(n832), .Y(
        n1218) );
  AO21X1_HVT U394 ( .A1(n144), .A2(n1552), .A3(n170), .Y(n1498) );
  AO22X1_HVT U395 ( .A1(n1497), .A2(n193), .A3(\mem[3][14] ), .A4(n831), .Y(
        n1217) );
  AO21X1_HVT U396 ( .A1(n144), .A2(n1550), .A3(n170), .Y(n1497) );
  AO22X1_HVT U397 ( .A1(n1496), .A2(n193), .A3(\mem[3][15] ), .A4(n830), .Y(
        n1216) );
  AO21X1_HVT U398 ( .A1(n144), .A2(n1548), .A3(n170), .Y(n1496) );
  AND2X1_HVT U400 ( .A1(n1023), .A2(n894), .Y(n1546) );
  AO22X1_HVT U401 ( .A1(n1494), .A2(n193), .A3(\mem[4][0] ), .A4(n829), .Y(
        n1215) );
  AO21X1_HVT U402 ( .A1(n141), .A2(n1579), .A3(n170), .Y(n1494) );
  AO22X1_HVT U403 ( .A1(n1492), .A2(n193), .A3(\mem[4][1] ), .A4(n828), .Y(
        n1214) );
  AO21X1_HVT U404 ( .A1(n143), .A2(n1576), .A3(n170), .Y(n1492) );
  AO22X1_HVT U405 ( .A1(n1491), .A2(n193), .A3(\mem[4][2] ), .A4(n827), .Y(
        n1213) );
  AO21X1_HVT U406 ( .A1(n142), .A2(n1574), .A3(n170), .Y(n1491) );
  AO22X1_HVT U407 ( .A1(n1490), .A2(n193), .A3(\mem[4][3] ), .A4(n826), .Y(
        n1212) );
  AO21X1_HVT U408 ( .A1(n141), .A2(n1572), .A3(n170), .Y(n1490) );
  AO22X1_HVT U409 ( .A1(n1489), .A2(n193), .A3(\mem[4][4] ), .A4(n338), .Y(
        n1211) );
  AO21X1_HVT U410 ( .A1(n143), .A2(n1570), .A3(n170), .Y(n1489) );
  AO22X1_HVT U411 ( .A1(n1488), .A2(n193), .A3(\mem[4][5] ), .A4(n320), .Y(
        n1210) );
  AO21X1_HVT U412 ( .A1(n142), .A2(n1568), .A3(n171), .Y(n1488) );
  AO22X1_HVT U413 ( .A1(n1487), .A2(n193), .A3(\mem[4][6] ), .A4(n302), .Y(
        n1209) );
  AO21X1_HVT U414 ( .A1(n141), .A2(n1566), .A3(n171), .Y(n1487) );
  AO22X1_HVT U415 ( .A1(n1486), .A2(n193), .A3(\mem[4][7] ), .A4(n265), .Y(
        n1208) );
  AO21X1_HVT U416 ( .A1(n143), .A2(n1564), .A3(n171), .Y(n1486) );
  AO22X1_HVT U417 ( .A1(n1485), .A2(n194), .A3(\mem[4][8] ), .A4(n264), .Y(
        n1207) );
  AO21X1_HVT U418 ( .A1(n142), .A2(n1562), .A3(n171), .Y(n1485) );
  AO22X1_HVT U419 ( .A1(n1484), .A2(n194), .A3(\mem[4][9] ), .A4(n263), .Y(
        n1206) );
  AO21X1_HVT U420 ( .A1(n141), .A2(n1560), .A3(n171), .Y(n1484) );
  AO22X1_HVT U421 ( .A1(n1483), .A2(n194), .A3(\mem[4][10] ), .A4(n262), .Y(
        n1205) );
  AO21X1_HVT U422 ( .A1(n143), .A2(n1558), .A3(n171), .Y(n1483) );
  AO22X1_HVT U423 ( .A1(n1482), .A2(n194), .A3(\mem[4][11] ), .A4(n261), .Y(
        n1204) );
  AO21X1_HVT U424 ( .A1(n142), .A2(n1556), .A3(n171), .Y(n1482) );
  AO22X1_HVT U425 ( .A1(n1481), .A2(n194), .A3(\mem[4][12] ), .A4(n260), .Y(
        n1203) );
  AO21X1_HVT U426 ( .A1(n141), .A2(n1554), .A3(n171), .Y(n1481) );
  AO22X1_HVT U427 ( .A1(n1480), .A2(n194), .A3(\mem[4][13] ), .A4(n259), .Y(
        n1202) );
  AO21X1_HVT U428 ( .A1(n143), .A2(n1552), .A3(n171), .Y(n1480) );
  AO22X1_HVT U429 ( .A1(n1479), .A2(n194), .A3(\mem[4][14] ), .A4(n258), .Y(
        n1201) );
  AO21X1_HVT U430 ( .A1(n142), .A2(n1550), .A3(n171), .Y(n1479) );
  AO22X1_HVT U431 ( .A1(n1478), .A2(n194), .A3(\mem[4][15] ), .A4(n257), .Y(
        n1200) );
  AO21X1_HVT U432 ( .A1(n141), .A2(n1548), .A3(n171), .Y(n1478) );
  AND3X1_HVT U433 ( .A1(n1547), .A2(n162), .A3(n1477), .Y(n1493) );
  AO22X1_HVT U434 ( .A1(n1476), .A2(n194), .A3(\mem[5][0] ), .A4(n256), .Y(
        n1199) );
  AO21X1_HVT U435 ( .A1(n138), .A2(n1579), .A3(n171), .Y(n1476) );
  AO22X1_HVT U436 ( .A1(n1474), .A2(n194), .A3(\mem[5][1] ), .A4(n255), .Y(
        n1198) );
  AO21X1_HVT U437 ( .A1(n140), .A2(n1576), .A3(n171), .Y(n1474) );
  AO22X1_HVT U438 ( .A1(n1473), .A2(n194), .A3(\mem[5][2] ), .A4(n254), .Y(
        n1197) );
  AO21X1_HVT U439 ( .A1(n139), .A2(n1574), .A3(n171), .Y(n1473) );
  AO22X1_HVT U440 ( .A1(n1472), .A2(n194), .A3(\mem[5][3] ), .A4(n253), .Y(
        n1196) );
  AO21X1_HVT U441 ( .A1(n138), .A2(n1572), .A3(n171), .Y(n1472) );
  AO22X1_HVT U442 ( .A1(n1471), .A2(n195), .A3(\mem[5][4] ), .A4(n252), .Y(
        n1195) );
  AO21X1_HVT U443 ( .A1(n140), .A2(n1570), .A3(n172), .Y(n1471) );
  AO22X1_HVT U444 ( .A1(n1470), .A2(n195), .A3(\mem[5][5] ), .A4(n251), .Y(
        n1194) );
  AO21X1_HVT U445 ( .A1(n139), .A2(n1568), .A3(n172), .Y(n1470) );
  AO22X1_HVT U446 ( .A1(n1469), .A2(n195), .A3(\mem[5][6] ), .A4(n250), .Y(
        n1193) );
  AO21X1_HVT U447 ( .A1(n138), .A2(n1566), .A3(n172), .Y(n1469) );
  AO22X1_HVT U448 ( .A1(n1468), .A2(n195), .A3(\mem[5][7] ), .A4(n249), .Y(
        n1192) );
  AO21X1_HVT U449 ( .A1(n140), .A2(n1564), .A3(n172), .Y(n1468) );
  AO22X1_HVT U450 ( .A1(n1467), .A2(n195), .A3(\mem[5][8] ), .A4(n248), .Y(
        n1191) );
  AO21X1_HVT U451 ( .A1(n139), .A2(n1562), .A3(n172), .Y(n1467) );
  AO22X1_HVT U452 ( .A1(n1466), .A2(n195), .A3(\mem[5][9] ), .A4(n247), .Y(
        n1190) );
  AO21X1_HVT U453 ( .A1(n138), .A2(n1560), .A3(n172), .Y(n1466) );
  AO22X1_HVT U454 ( .A1(n1465), .A2(n195), .A3(\mem[5][10] ), .A4(n246), .Y(
        n1189) );
  AO21X1_HVT U455 ( .A1(n140), .A2(n1558), .A3(n172), .Y(n1465) );
  AO22X1_HVT U456 ( .A1(n1464), .A2(n195), .A3(\mem[5][11] ), .A4(n245), .Y(
        n1188) );
  AO21X1_HVT U457 ( .A1(n139), .A2(n1556), .A3(n172), .Y(n1464) );
  AO22X1_HVT U458 ( .A1(n1463), .A2(n195), .A3(\mem[5][12] ), .A4(n244), .Y(
        n1187) );
  AO21X1_HVT U459 ( .A1(n138), .A2(n1554), .A3(n172), .Y(n1463) );
  AO22X1_HVT U460 ( .A1(n1462), .A2(n195), .A3(\mem[5][13] ), .A4(n243), .Y(
        n1186) );
  AO21X1_HVT U461 ( .A1(n140), .A2(n1552), .A3(n172), .Y(n1462) );
  AO22X1_HVT U462 ( .A1(n1461), .A2(n195), .A3(\mem[5][14] ), .A4(n242), .Y(
        n1185) );
  AO21X1_HVT U463 ( .A1(n139), .A2(n1550), .A3(n172), .Y(n1461) );
  AO22X1_HVT U464 ( .A1(n1460), .A2(n195), .A3(\mem[5][15] ), .A4(n241), .Y(
        n1184) );
  AO21X1_HVT U465 ( .A1(n138), .A2(n1548), .A3(n172), .Y(n1460) );
  AND3X1_HVT U466 ( .A1(n1529), .A2(n4), .A3(n1477), .Y(n1475) );
  AO22X1_HVT U467 ( .A1(n1459), .A2(n208), .A3(\mem[6][0] ), .A4(n240), .Y(
        n1183) );
  AO21X1_HVT U468 ( .A1(n135), .A2(n1579), .A3(n172), .Y(n1459) );
  AO22X1_HVT U469 ( .A1(n1457), .A2(n184), .A3(\mem[6][1] ), .A4(n239), .Y(
        n1182) );
  AO21X1_HVT U470 ( .A1(n137), .A2(n1576), .A3(n172), .Y(n1457) );
  AO22X1_HVT U471 ( .A1(n1456), .A2(n185), .A3(\mem[6][2] ), .A4(n238), .Y(
        n1181) );
  AO21X1_HVT U472 ( .A1(n136), .A2(n1574), .A3(n172), .Y(n1456) );
  AO22X1_HVT U473 ( .A1(n1455), .A2(n186), .A3(\mem[6][3] ), .A4(n237), .Y(
        n1180) );
  AO21X1_HVT U474 ( .A1(n135), .A2(n1572), .A3(n173), .Y(n1455) );
  AO22X1_HVT U475 ( .A1(n1454), .A2(n188), .A3(\mem[6][4] ), .A4(n236), .Y(
        n1179) );
  AO21X1_HVT U476 ( .A1(n137), .A2(n1570), .A3(n173), .Y(n1454) );
  AO22X1_HVT U477 ( .A1(n1453), .A2(n208), .A3(\mem[6][5] ), .A4(n235), .Y(
        n1178) );
  AO21X1_HVT U478 ( .A1(n136), .A2(n1568), .A3(n173), .Y(n1453) );
  AO22X1_HVT U479 ( .A1(n1452), .A2(n184), .A3(\mem[6][6] ), .A4(n234), .Y(
        n1177) );
  AO21X1_HVT U480 ( .A1(n135), .A2(n1566), .A3(n173), .Y(n1452) );
  AO22X1_HVT U481 ( .A1(n1451), .A2(n185), .A3(\mem[6][7] ), .A4(n233), .Y(
        n1176) );
  AO21X1_HVT U482 ( .A1(n137), .A2(n1564), .A3(n173), .Y(n1451) );
  AO22X1_HVT U483 ( .A1(n1450), .A2(n186), .A3(\mem[6][8] ), .A4(n232), .Y(
        n1175) );
  AO21X1_HVT U484 ( .A1(n136), .A2(n1562), .A3(n173), .Y(n1450) );
  AO22X1_HVT U485 ( .A1(n1449), .A2(n188), .A3(\mem[6][9] ), .A4(n231), .Y(
        n1174) );
  AO21X1_HVT U486 ( .A1(n135), .A2(n1560), .A3(n173), .Y(n1449) );
  AO22X1_HVT U487 ( .A1(n1448), .A2(n188), .A3(\mem[6][10] ), .A4(n230), .Y(
        n1173) );
  AO21X1_HVT U488 ( .A1(n137), .A2(n1558), .A3(n173), .Y(n1448) );
  AO22X1_HVT U489 ( .A1(n1447), .A2(n188), .A3(\mem[6][11] ), .A4(n229), .Y(
        n1172) );
  AO21X1_HVT U490 ( .A1(n136), .A2(n1556), .A3(n173), .Y(n1447) );
  AO22X1_HVT U491 ( .A1(n1446), .A2(n196), .A3(\mem[6][12] ), .A4(n228), .Y(
        n1171) );
  AO21X1_HVT U492 ( .A1(n135), .A2(n1554), .A3(n173), .Y(n1446) );
  AO22X1_HVT U493 ( .A1(n1445), .A2(n196), .A3(\mem[6][13] ), .A4(n227), .Y(
        n1170) );
  AO21X1_HVT U494 ( .A1(n137), .A2(n1552), .A3(n173), .Y(n1445) );
  AO22X1_HVT U495 ( .A1(n1444), .A2(n196), .A3(\mem[6][14] ), .A4(n226), .Y(
        n1169) );
  AO21X1_HVT U496 ( .A1(n136), .A2(n1550), .A3(n173), .Y(n1444) );
  AO22X1_HVT U497 ( .A1(n1443), .A2(n196), .A3(\mem[6][15] ), .A4(n225), .Y(
        n1168) );
  AO21X1_HVT U498 ( .A1(n135), .A2(n1548), .A3(n173), .Y(n1443) );
  AND3X1_HVT U499 ( .A1(n1512), .A2(n163), .A3(n1477), .Y(n1458) );
  AO22X1_HVT U500 ( .A1(n1442), .A2(n196), .A3(\mem[7][0] ), .A4(n224), .Y(
        n1167) );
  AO21X1_HVT U501 ( .A1(n132), .A2(n1579), .A3(n173), .Y(n1442) );
  AO22X1_HVT U502 ( .A1(n1440), .A2(n196), .A3(\mem[7][1] ), .A4(n223), .Y(
        n1166) );
  AO21X1_HVT U503 ( .A1(n134), .A2(n1576), .A3(n173), .Y(n1440) );
  AO22X1_HVT U504 ( .A1(n1439), .A2(n196), .A3(\mem[7][2] ), .A4(n222), .Y(
        n1165) );
  AO21X1_HVT U505 ( .A1(n133), .A2(n1574), .A3(n174), .Y(n1439) );
  AO22X1_HVT U506 ( .A1(n1438), .A2(n196), .A3(\mem[7][3] ), .A4(n221), .Y(
        n1164) );
  AO21X1_HVT U507 ( .A1(n132), .A2(n1572), .A3(n174), .Y(n1438) );
  AO22X1_HVT U508 ( .A1(n1437), .A2(n196), .A3(\mem[7][4] ), .A4(n220), .Y(
        n1163) );
  AO21X1_HVT U509 ( .A1(n134), .A2(n1570), .A3(n174), .Y(n1437) );
  AO22X1_HVT U510 ( .A1(n1436), .A2(n196), .A3(\mem[7][5] ), .A4(n219), .Y(
        n1162) );
  AO21X1_HVT U511 ( .A1(n133), .A2(n1568), .A3(n174), .Y(n1436) );
  AO22X1_HVT U512 ( .A1(n1435), .A2(n196), .A3(\mem[7][6] ), .A4(n218), .Y(
        n1161) );
  AO21X1_HVT U513 ( .A1(n132), .A2(n1566), .A3(n174), .Y(n1435) );
  AO22X1_HVT U514 ( .A1(n1434), .A2(n196), .A3(\mem[7][7] ), .A4(n217), .Y(
        n1160) );
  AO21X1_HVT U515 ( .A1(n134), .A2(n1564), .A3(n174), .Y(n1434) );
  AO22X1_HVT U516 ( .A1(n1433), .A2(n197), .A3(\mem[7][8] ), .A4(n216), .Y(
        n1159) );
  AO21X1_HVT U517 ( .A1(n133), .A2(n1562), .A3(n174), .Y(n1433) );
  AO22X1_HVT U518 ( .A1(n1432), .A2(n197), .A3(\mem[7][9] ), .A4(n215), .Y(
        n1158) );
  AO21X1_HVT U519 ( .A1(n132), .A2(n1560), .A3(n174), .Y(n1432) );
  AO22X1_HVT U520 ( .A1(n1431), .A2(n197), .A3(\mem[7][10] ), .A4(n214), .Y(
        n1157) );
  AO21X1_HVT U521 ( .A1(n134), .A2(n1558), .A3(n174), .Y(n1431) );
  AO22X1_HVT U522 ( .A1(n1430), .A2(n197), .A3(\mem[7][11] ), .A4(n213), .Y(
        n1156) );
  AO21X1_HVT U523 ( .A1(n133), .A2(n1556), .A3(n174), .Y(n1430) );
  AO22X1_HVT U524 ( .A1(n1429), .A2(n197), .A3(\mem[7][12] ), .A4(n212), .Y(
        n1155) );
  AO21X1_HVT U525 ( .A1(n132), .A2(n1554), .A3(n174), .Y(n1429) );
  AO22X1_HVT U526 ( .A1(n1428), .A2(n197), .A3(\mem[7][13] ), .A4(n211), .Y(
        n1154) );
  AO21X1_HVT U527 ( .A1(n134), .A2(n1552), .A3(n174), .Y(n1428) );
  AO22X1_HVT U528 ( .A1(n1427), .A2(n197), .A3(\mem[7][14] ), .A4(n210), .Y(
        n1153) );
  AO21X1_HVT U529 ( .A1(n133), .A2(n1550), .A3(n174), .Y(n1427) );
  AO22X1_HVT U530 ( .A1(n1426), .A2(n197), .A3(\mem[7][15] ), .A4(n209), .Y(
        n1152) );
  AO21X1_HVT U531 ( .A1(n132), .A2(n1548), .A3(n174), .Y(n1426) );
  AND3X1_HVT U532 ( .A1(n1495), .A2(n162), .A3(n1477), .Y(n1441) );
  AND2X1_HVT U533 ( .A1(a_din[2]), .A2(n894), .Y(n1477) );
  AO22X1_HVT U534 ( .A1(n1425), .A2(n197), .A3(\mem[8][0] ), .A4(n958), .Y(
        n1151) );
  AO21X1_HVT U535 ( .A1(n129), .A2(n1579), .A3(n174), .Y(n1425) );
  AO22X1_HVT U536 ( .A1(n1423), .A2(n197), .A3(\mem[8][1] ), .A4(n957), .Y(
        n1150) );
  AO21X1_HVT U537 ( .A1(n131), .A2(n1576), .A3(n175), .Y(n1423) );
  AO22X1_HVT U538 ( .A1(n1422), .A2(n197), .A3(\mem[8][2] ), .A4(n956), .Y(
        n1149) );
  AO21X1_HVT U539 ( .A1(n130), .A2(n1574), .A3(n175), .Y(n1422) );
  AO22X1_HVT U540 ( .A1(n1421), .A2(n197), .A3(\mem[8][3] ), .A4(n955), .Y(
        n1148) );
  AO21X1_HVT U541 ( .A1(n129), .A2(n1572), .A3(n175), .Y(n1421) );
  AO22X1_HVT U542 ( .A1(n1420), .A2(n198), .A3(\mem[8][4] ), .A4(n954), .Y(
        n1147) );
  AO21X1_HVT U543 ( .A1(n131), .A2(n1570), .A3(n175), .Y(n1420) );
  AO22X1_HVT U544 ( .A1(n1419), .A2(n198), .A3(\mem[8][5] ), .A4(n953), .Y(
        n1146) );
  AO21X1_HVT U545 ( .A1(n130), .A2(n1568), .A3(n175), .Y(n1419) );
  AO22X1_HVT U546 ( .A1(n1418), .A2(n198), .A3(\mem[8][6] ), .A4(n952), .Y(
        n1145) );
  AO21X1_HVT U547 ( .A1(n129), .A2(n1566), .A3(n175), .Y(n1418) );
  AO22X1_HVT U548 ( .A1(n1417), .A2(n198), .A3(\mem[8][7] ), .A4(n951), .Y(
        n1144) );
  AO21X1_HVT U549 ( .A1(n131), .A2(n1564), .A3(n175), .Y(n1417) );
  AO22X1_HVT U550 ( .A1(n1416), .A2(n198), .A3(\mem[8][8] ), .A4(n950), .Y(
        n1143) );
  AO21X1_HVT U551 ( .A1(n130), .A2(n1562), .A3(n175), .Y(n1416) );
  AO22X1_HVT U552 ( .A1(n1415), .A2(n198), .A3(\mem[8][9] ), .A4(n949), .Y(
        n1142) );
  AO21X1_HVT U553 ( .A1(n129), .A2(n1560), .A3(n175), .Y(n1415) );
  AO22X1_HVT U554 ( .A1(n1414), .A2(n198), .A3(\mem[8][10] ), .A4(n948), .Y(
        n1141) );
  AO21X1_HVT U555 ( .A1(n131), .A2(n1558), .A3(n175), .Y(n1414) );
  AO22X1_HVT U556 ( .A1(n1413), .A2(n198), .A3(\mem[8][11] ), .A4(n947), .Y(
        n1140) );
  AO21X1_HVT U557 ( .A1(n130), .A2(n1556), .A3(n175), .Y(n1413) );
  AO22X1_HVT U558 ( .A1(n1412), .A2(n198), .A3(\mem[8][12] ), .A4(n946), .Y(
        n1139) );
  AO21X1_HVT U559 ( .A1(n129), .A2(n1554), .A3(n175), .Y(n1412) );
  AO22X1_HVT U560 ( .A1(n1411), .A2(n198), .A3(\mem[8][13] ), .A4(n945), .Y(
        n1138) );
  AO21X1_HVT U561 ( .A1(n131), .A2(n1552), .A3(n175), .Y(n1411) );
  AO22X1_HVT U562 ( .A1(n1410), .A2(n198), .A3(\mem[8][14] ), .A4(n944), .Y(
        n1137) );
  AO21X1_HVT U563 ( .A1(n130), .A2(n1550), .A3(n175), .Y(n1410) );
  AO22X1_HVT U564 ( .A1(n1409), .A2(n198), .A3(\mem[8][15] ), .A4(n943), .Y(
        n1136) );
  AO21X1_HVT U565 ( .A1(n129), .A2(n1548), .A3(n175), .Y(n1409) );
  AND3X1_HVT U566 ( .A1(n1547), .A2(n4), .A3(n1408), .Y(n1424) );
  AO22X1_HVT U567 ( .A1(n1407), .A2(n199), .A3(\mem[9][0] ), .A4(n942), .Y(
        n1135) );
  AO21X1_HVT U568 ( .A1(n126), .A2(n1579), .A3(n176), .Y(n1407) );
  AO22X1_HVT U569 ( .A1(n1405), .A2(n199), .A3(\mem[9][1] ), .A4(n941), .Y(
        n1134) );
  AO21X1_HVT U570 ( .A1(n128), .A2(n1576), .A3(n176), .Y(n1405) );
  AO22X1_HVT U571 ( .A1(n1404), .A2(n199), .A3(\mem[9][2] ), .A4(n940), .Y(
        n1133) );
  AO21X1_HVT U572 ( .A1(n127), .A2(n1574), .A3(n176), .Y(n1404) );
  AO22X1_HVT U573 ( .A1(n1403), .A2(n199), .A3(\mem[9][3] ), .A4(n939), .Y(
        n1132) );
  AO21X1_HVT U574 ( .A1(n126), .A2(n1572), .A3(n176), .Y(n1403) );
  AO22X1_HVT U575 ( .A1(n1402), .A2(n199), .A3(\mem[9][4] ), .A4(n938), .Y(
        n1131) );
  AO21X1_HVT U576 ( .A1(n128), .A2(n1570), .A3(n176), .Y(n1402) );
  AO22X1_HVT U577 ( .A1(n1401), .A2(n199), .A3(\mem[9][5] ), .A4(n937), .Y(
        n1130) );
  AO21X1_HVT U578 ( .A1(n127), .A2(n1568), .A3(n176), .Y(n1401) );
  AO22X1_HVT U579 ( .A1(n1400), .A2(n199), .A3(\mem[9][6] ), .A4(n936), .Y(
        n1129) );
  AO21X1_HVT U580 ( .A1(n126), .A2(n1566), .A3(n176), .Y(n1400) );
  AO22X1_HVT U581 ( .A1(n1399), .A2(n199), .A3(\mem[9][7] ), .A4(n935), .Y(
        n1128) );
  AO21X1_HVT U582 ( .A1(n128), .A2(n1564), .A3(n176), .Y(n1399) );
  AO22X1_HVT U583 ( .A1(n1398), .A2(n199), .A3(\mem[9][8] ), .A4(n934), .Y(
        n1127) );
  AO21X1_HVT U584 ( .A1(n127), .A2(n1562), .A3(n176), .Y(n1398) );
  AO22X1_HVT U585 ( .A1(n1397), .A2(n199), .A3(\mem[9][9] ), .A4(n933), .Y(
        n1126) );
  AO21X1_HVT U586 ( .A1(n126), .A2(n1560), .A3(n176), .Y(n1397) );
  AO22X1_HVT U587 ( .A1(n1396), .A2(n199), .A3(\mem[9][10] ), .A4(n932), .Y(
        n1125) );
  AO21X1_HVT U588 ( .A1(n128), .A2(n1558), .A3(n176), .Y(n1396) );
  AO22X1_HVT U589 ( .A1(n1395), .A2(n199), .A3(\mem[9][11] ), .A4(n931), .Y(
        n1124) );
  AO21X1_HVT U590 ( .A1(n127), .A2(n1556), .A3(n176), .Y(n1395) );
  AO22X1_HVT U591 ( .A1(n1394), .A2(n200), .A3(\mem[9][12] ), .A4(n930), .Y(
        n1123) );
  AO21X1_HVT U592 ( .A1(n126), .A2(n1554), .A3(n176), .Y(n1394) );
  AO22X1_HVT U593 ( .A1(n1393), .A2(n200), .A3(\mem[9][13] ), .A4(n929), .Y(
        n1122) );
  AO21X1_HVT U594 ( .A1(n128), .A2(n1552), .A3(n176), .Y(n1393) );
  AO22X1_HVT U595 ( .A1(n1392), .A2(n200), .A3(\mem[9][14] ), .A4(n928), .Y(
        n1121) );
  AO21X1_HVT U596 ( .A1(n127), .A2(n1550), .A3(n176), .Y(n1392) );
  AO22X1_HVT U597 ( .A1(n1391), .A2(n200), .A3(\mem[9][15] ), .A4(n927), .Y(
        n1120) );
  AO21X1_HVT U598 ( .A1(n126), .A2(n1548), .A3(n177), .Y(n1391) );
  AND3X1_HVT U599 ( .A1(n1529), .A2(n163), .A3(n1408), .Y(n1406) );
  AO22X1_HVT U600 ( .A1(n1390), .A2(n200), .A3(\mem[10][0] ), .A4(n926), .Y(
        n1119) );
  AO21X1_HVT U601 ( .A1(n123), .A2(n1579), .A3(n177), .Y(n1390) );
  AO22X1_HVT U602 ( .A1(n1388), .A2(n200), .A3(\mem[10][1] ), .A4(n925), .Y(
        n1118) );
  AO21X1_HVT U603 ( .A1(n125), .A2(n1576), .A3(n177), .Y(n1388) );
  AO22X1_HVT U604 ( .A1(n1387), .A2(n200), .A3(\mem[10][2] ), .A4(n924), .Y(
        n1117) );
  AO21X1_HVT U605 ( .A1(n124), .A2(n1574), .A3(n177), .Y(n1387) );
  AO22X1_HVT U606 ( .A1(n1386), .A2(n200), .A3(\mem[10][3] ), .A4(n923), .Y(
        n1116) );
  AO21X1_HVT U607 ( .A1(n123), .A2(n1572), .A3(n177), .Y(n1386) );
  AO22X1_HVT U608 ( .A1(n1385), .A2(n200), .A3(\mem[10][4] ), .A4(n922), .Y(
        n1115) );
  AO21X1_HVT U609 ( .A1(n125), .A2(n1570), .A3(n177), .Y(n1385) );
  AO22X1_HVT U610 ( .A1(n1384), .A2(n200), .A3(\mem[10][5] ), .A4(n921), .Y(
        n1114) );
  AO21X1_HVT U611 ( .A1(n124), .A2(n1568), .A3(n177), .Y(n1384) );
  AO22X1_HVT U612 ( .A1(n1383), .A2(n200), .A3(\mem[10][6] ), .A4(n920), .Y(
        n1113) );
  AO21X1_HVT U613 ( .A1(n123), .A2(n1566), .A3(n177), .Y(n1383) );
  AO22X1_HVT U614 ( .A1(n1382), .A2(n200), .A3(\mem[10][7] ), .A4(n919), .Y(
        n1112) );
  AO21X1_HVT U615 ( .A1(n125), .A2(n1564), .A3(n177), .Y(n1382) );
  AO22X1_HVT U616 ( .A1(n1381), .A2(n201), .A3(\mem[10][8] ), .A4(n918), .Y(
        n1111) );
  AO21X1_HVT U617 ( .A1(n124), .A2(n1562), .A3(n177), .Y(n1381) );
  AO22X1_HVT U618 ( .A1(n1380), .A2(n201), .A3(\mem[10][9] ), .A4(n917), .Y(
        n1110) );
  AO21X1_HVT U619 ( .A1(n123), .A2(n1560), .A3(n177), .Y(n1380) );
  AO22X1_HVT U620 ( .A1(n1379), .A2(n201), .A3(\mem[10][10] ), .A4(n916), .Y(
        n1109) );
  AO21X1_HVT U621 ( .A1(n125), .A2(n1558), .A3(n177), .Y(n1379) );
  AO22X1_HVT U622 ( .A1(n1378), .A2(n201), .A3(\mem[10][11] ), .A4(n915), .Y(
        n1108) );
  AO21X1_HVT U623 ( .A1(n124), .A2(n1556), .A3(n177), .Y(n1378) );
  AO22X1_HVT U624 ( .A1(n1377), .A2(n201), .A3(\mem[10][12] ), .A4(n914), .Y(
        n1107) );
  AO21X1_HVT U625 ( .A1(n123), .A2(n1554), .A3(n177), .Y(n1377) );
  AO22X1_HVT U626 ( .A1(n1376), .A2(n201), .A3(\mem[10][13] ), .A4(n913), .Y(
        n1106) );
  AO21X1_HVT U627 ( .A1(n125), .A2(n1552), .A3(n177), .Y(n1376) );
  AO22X1_HVT U628 ( .A1(n1375), .A2(n201), .A3(\mem[10][14] ), .A4(n912), .Y(
        n1105) );
  AO21X1_HVT U629 ( .A1(n124), .A2(n1550), .A3(n178), .Y(n1375) );
  AO22X1_HVT U630 ( .A1(n1374), .A2(n201), .A3(\mem[10][15] ), .A4(n911), .Y(
        n1104) );
  AO21X1_HVT U631 ( .A1(n123), .A2(n1548), .A3(n178), .Y(n1374) );
  AND3X1_HVT U632 ( .A1(n1512), .A2(n162), .A3(n1408), .Y(n1389) );
  AO22X1_HVT U633 ( .A1(n1373), .A2(n201), .A3(\mem[11][0] ), .A4(n910), .Y(
        n1103) );
  AO21X1_HVT U634 ( .A1(n120), .A2(n1579), .A3(n178), .Y(n1373) );
  AO22X1_HVT U635 ( .A1(n1371), .A2(n201), .A3(\mem[11][1] ), .A4(n909), .Y(
        n1102) );
  AO21X1_HVT U636 ( .A1(n122), .A2(n1576), .A3(n178), .Y(n1371) );
  AO22X1_HVT U637 ( .A1(n1370), .A2(n201), .A3(\mem[11][2] ), .A4(n908), .Y(
        n1101) );
  AO21X1_HVT U638 ( .A1(n121), .A2(n1574), .A3(n178), .Y(n1370) );
  AO22X1_HVT U639 ( .A1(n1369), .A2(n201), .A3(\mem[11][3] ), .A4(n907), .Y(
        n1100) );
  AO21X1_HVT U640 ( .A1(n120), .A2(n1572), .A3(n178), .Y(n1369) );
  AO22X1_HVT U641 ( .A1(n1368), .A2(n202), .A3(\mem[11][4] ), .A4(n906), .Y(
        n1099) );
  AO21X1_HVT U642 ( .A1(n122), .A2(n1570), .A3(n178), .Y(n1368) );
  AO22X1_HVT U643 ( .A1(n1367), .A2(n202), .A3(\mem[11][5] ), .A4(n905), .Y(
        n1098) );
  AO21X1_HVT U644 ( .A1(n121), .A2(n1568), .A3(n178), .Y(n1367) );
  AO22X1_HVT U645 ( .A1(n1366), .A2(n202), .A3(\mem[11][6] ), .A4(n904), .Y(
        n1097) );
  AO21X1_HVT U646 ( .A1(n120), .A2(n1566), .A3(n178), .Y(n1366) );
  AO22X1_HVT U647 ( .A1(n1365), .A2(n202), .A3(\mem[11][7] ), .A4(n903), .Y(
        n1096) );
  AO21X1_HVT U648 ( .A1(n122), .A2(n1564), .A3(n178), .Y(n1365) );
  AO22X1_HVT U649 ( .A1(n1364), .A2(n202), .A3(\mem[11][8] ), .A4(n902), .Y(
        n1095) );
  AO21X1_HVT U650 ( .A1(n121), .A2(n1562), .A3(n178), .Y(n1364) );
  AO22X1_HVT U651 ( .A1(n1363), .A2(n202), .A3(\mem[11][9] ), .A4(n901), .Y(
        n1094) );
  AO21X1_HVT U652 ( .A1(n120), .A2(n1560), .A3(n178), .Y(n1363) );
  AO22X1_HVT U653 ( .A1(n1362), .A2(n202), .A3(\mem[11][10] ), .A4(n900), .Y(
        n1093) );
  AO21X1_HVT U654 ( .A1(n122), .A2(n1558), .A3(n178), .Y(n1362) );
  AO22X1_HVT U655 ( .A1(n1361), .A2(n202), .A3(\mem[11][11] ), .A4(n899), .Y(
        n1092) );
  AO21X1_HVT U656 ( .A1(n121), .A2(n1556), .A3(n178), .Y(n1361) );
  AO22X1_HVT U657 ( .A1(n1360), .A2(n202), .A3(\mem[11][12] ), .A4(n898), .Y(
        n1091) );
  AO21X1_HVT U658 ( .A1(n120), .A2(n1554), .A3(n178), .Y(n1360) );
  AO22X1_HVT U659 ( .A1(n1359), .A2(n202), .A3(\mem[11][13] ), .A4(n897), .Y(
        n1090) );
  AO21X1_HVT U660 ( .A1(n122), .A2(n1552), .A3(n179), .Y(n1359) );
  AO22X1_HVT U661 ( .A1(n1358), .A2(n202), .A3(\mem[11][14] ), .A4(n896), .Y(
        n1089) );
  AO21X1_HVT U662 ( .A1(n121), .A2(n1550), .A3(n179), .Y(n1358) );
  AO22X1_HVT U663 ( .A1(n1357), .A2(n202), .A3(\mem[11][15] ), .A4(n895), .Y(
        n1088) );
  AO21X1_HVT U664 ( .A1(n120), .A2(n1548), .A3(n179), .Y(n1357) );
  AND3X1_HVT U665 ( .A1(n1495), .A2(n4), .A3(n1408), .Y(n1372) );
  AND2X1_HVT U666 ( .A1(a_din[3]), .A2(n1023), .Y(n1408) );
  AO22X1_HVT U667 ( .A1(n1356), .A2(n203), .A3(\mem[12][0] ), .A4(n1022), .Y(
        n1087) );
  AO21X1_HVT U668 ( .A1(n117), .A2(n1579), .A3(n179), .Y(n1356) );
  AO22X1_HVT U669 ( .A1(n1354), .A2(n203), .A3(\mem[12][1] ), .A4(n1021), .Y(
        n1086) );
  AO21X1_HVT U670 ( .A1(n119), .A2(n1576), .A3(n179), .Y(n1354) );
  AO22X1_HVT U671 ( .A1(n1353), .A2(n203), .A3(\mem[12][2] ), .A4(n1020), .Y(
        n1085) );
  AO21X1_HVT U672 ( .A1(n118), .A2(n1574), .A3(n179), .Y(n1353) );
  AO22X1_HVT U673 ( .A1(n1352), .A2(n203), .A3(\mem[12][3] ), .A4(n1019), .Y(
        n1084) );
  AO21X1_HVT U674 ( .A1(n117), .A2(n1572), .A3(n179), .Y(n1352) );
  AO22X1_HVT U675 ( .A1(n1351), .A2(n203), .A3(\mem[12][4] ), .A4(n1018), .Y(
        n1083) );
  AO21X1_HVT U676 ( .A1(n119), .A2(n1570), .A3(n179), .Y(n1351) );
  AO22X1_HVT U677 ( .A1(n1350), .A2(n203), .A3(\mem[12][5] ), .A4(n1017), .Y(
        n1082) );
  AO21X1_HVT U678 ( .A1(n118), .A2(n1568), .A3(n179), .Y(n1350) );
  AO22X1_HVT U679 ( .A1(n1349), .A2(n203), .A3(\mem[12][6] ), .A4(n1016), .Y(
        n1081) );
  AO21X1_HVT U680 ( .A1(n117), .A2(n1566), .A3(n179), .Y(n1349) );
  AO22X1_HVT U681 ( .A1(n1348), .A2(n203), .A3(\mem[12][7] ), .A4(n1015), .Y(
        n1080) );
  AO21X1_HVT U682 ( .A1(n119), .A2(n1564), .A3(n179), .Y(n1348) );
  AO22X1_HVT U683 ( .A1(n1347), .A2(n203), .A3(\mem[12][8] ), .A4(n1014), .Y(
        n1079) );
  AO21X1_HVT U684 ( .A1(n118), .A2(n1562), .A3(n179), .Y(n1347) );
  AO22X1_HVT U685 ( .A1(n1346), .A2(n203), .A3(\mem[12][9] ), .A4(n1013), .Y(
        n1078) );
  AO21X1_HVT U686 ( .A1(n117), .A2(n1560), .A3(n179), .Y(n1346) );
  AO22X1_HVT U687 ( .A1(n1345), .A2(n203), .A3(\mem[12][10] ), .A4(n1012), .Y(
        n1077) );
  AO21X1_HVT U688 ( .A1(n119), .A2(n1558), .A3(n179), .Y(n1345) );
  AO22X1_HVT U689 ( .A1(n1344), .A2(n203), .A3(\mem[12][11] ), .A4(n1011), .Y(
        n1076) );
  AO21X1_HVT U690 ( .A1(n118), .A2(n1556), .A3(n179), .Y(n1344) );
  AO22X1_HVT U691 ( .A1(n1343), .A2(n204), .A3(\mem[12][12] ), .A4(n1010), .Y(
        n1075) );
  AO21X1_HVT U692 ( .A1(n117), .A2(n1554), .A3(n180), .Y(n1343) );
  AO22X1_HVT U693 ( .A1(n1342), .A2(n204), .A3(\mem[12][13] ), .A4(n1009), .Y(
        n1074) );
  AO21X1_HVT U694 ( .A1(n119), .A2(n1552), .A3(n180), .Y(n1342) );
  AO22X1_HVT U695 ( .A1(n1341), .A2(n204), .A3(\mem[12][14] ), .A4(n1008), .Y(
        n1073) );
  AO21X1_HVT U696 ( .A1(n118), .A2(n1550), .A3(n180), .Y(n1341) );
  AO22X1_HVT U697 ( .A1(n1340), .A2(n204), .A3(\mem[12][15] ), .A4(n1007), .Y(
        n1072) );
  AO21X1_HVT U698 ( .A1(n117), .A2(n1548), .A3(n180), .Y(n1340) );
  AND3X1_HVT U699 ( .A1(n1547), .A2(n4), .A3(n1339), .Y(n1355) );
  AND2X1_HVT U700 ( .A1(n153), .A2(n155), .Y(n1547) );
  AO22X1_HVT U701 ( .A1(n1338), .A2(n204), .A3(\mem[13][0] ), .A4(n1006), .Y(
        n1071) );
  AO21X1_HVT U702 ( .A1(n114), .A2(n1579), .A3(n180), .Y(n1338) );
  AO22X1_HVT U703 ( .A1(n1336), .A2(n204), .A3(\mem[13][1] ), .A4(n1005), .Y(
        n1070) );
  AO21X1_HVT U704 ( .A1(n116), .A2(n1576), .A3(n180), .Y(n1336) );
  AO22X1_HVT U705 ( .A1(n1335), .A2(n204), .A3(\mem[13][2] ), .A4(n1004), .Y(
        n1069) );
  AO21X1_HVT U706 ( .A1(n115), .A2(n1574), .A3(n180), .Y(n1335) );
  AO22X1_HVT U707 ( .A1(n1334), .A2(n204), .A3(\mem[13][3] ), .A4(n1003), .Y(
        n1068) );
  AO21X1_HVT U708 ( .A1(n114), .A2(n1572), .A3(n180), .Y(n1334) );
  AO22X1_HVT U709 ( .A1(n1333), .A2(n204), .A3(\mem[13][4] ), .A4(n1002), .Y(
        n1067) );
  AO21X1_HVT U710 ( .A1(n116), .A2(n1570), .A3(n180), .Y(n1333) );
  AO22X1_HVT U711 ( .A1(n1332), .A2(n204), .A3(\mem[13][5] ), .A4(n1001), .Y(
        n1066) );
  AO21X1_HVT U712 ( .A1(n115), .A2(n1568), .A3(n180), .Y(n1332) );
  AO22X1_HVT U713 ( .A1(n1331), .A2(n204), .A3(\mem[13][6] ), .A4(n1000), .Y(
        n1065) );
  AO21X1_HVT U714 ( .A1(n114), .A2(n1566), .A3(n180), .Y(n1331) );
  AO22X1_HVT U715 ( .A1(n1330), .A2(n204), .A3(\mem[13][7] ), .A4(n999), .Y(
        n1064) );
  AO21X1_HVT U716 ( .A1(n116), .A2(n1564), .A3(n180), .Y(n1330) );
  AO22X1_HVT U717 ( .A1(n1329), .A2(n205), .A3(\mem[13][8] ), .A4(n998), .Y(
        n1063) );
  AO21X1_HVT U718 ( .A1(n115), .A2(n1562), .A3(n180), .Y(n1329) );
  AO22X1_HVT U719 ( .A1(n1328), .A2(n205), .A3(\mem[13][9] ), .A4(n997), .Y(
        n1062) );
  AO21X1_HVT U720 ( .A1(n114), .A2(n1560), .A3(n180), .Y(n1328) );
  AO22X1_HVT U721 ( .A1(n1327), .A2(n205), .A3(\mem[13][10] ), .A4(n996), .Y(
        n1061) );
  AO21X1_HVT U722 ( .A1(n116), .A2(n1558), .A3(n180), .Y(n1327) );
  AO22X1_HVT U723 ( .A1(n1326), .A2(n205), .A3(\mem[13][11] ), .A4(n995), .Y(
        n1060) );
  AO21X1_HVT U724 ( .A1(n115), .A2(n1556), .A3(n181), .Y(n1326) );
  AO22X1_HVT U725 ( .A1(n1325), .A2(n205), .A3(\mem[13][12] ), .A4(n994), .Y(
        n1059) );
  AO21X1_HVT U726 ( .A1(n114), .A2(n1554), .A3(n181), .Y(n1325) );
  AO22X1_HVT U727 ( .A1(n1324), .A2(n205), .A3(\mem[13][13] ), .A4(n993), .Y(
        n1058) );
  AO21X1_HVT U728 ( .A1(n116), .A2(n1552), .A3(n181), .Y(n1324) );
  AO22X1_HVT U729 ( .A1(n1323), .A2(n205), .A3(\mem[13][14] ), .A4(n992), .Y(
        n1057) );
  AO21X1_HVT U730 ( .A1(n115), .A2(n1550), .A3(n181), .Y(n1323) );
  AO22X1_HVT U731 ( .A1(n1322), .A2(n205), .A3(\mem[13][15] ), .A4(n991), .Y(
        n1056) );
  AO21X1_HVT U732 ( .A1(n114), .A2(n1548), .A3(n181), .Y(n1322) );
  AND3X1_HVT U733 ( .A1(n1529), .A2(n162), .A3(n1339), .Y(n1337) );
  AND2X1_HVT U734 ( .A1(a_din[0]), .A2(n155), .Y(n1529) );
  AO22X1_HVT U735 ( .A1(n1321), .A2(n205), .A3(\mem[14][0] ), .A4(n990), .Y(
        n1055) );
  AO21X1_HVT U736 ( .A1(n111), .A2(n1579), .A3(n181), .Y(n1321) );
  AO22X1_HVT U737 ( .A1(n1319), .A2(n205), .A3(\mem[14][1] ), .A4(n989), .Y(
        n1054) );
  AO21X1_HVT U738 ( .A1(n113), .A2(n1576), .A3(n181), .Y(n1319) );
  AO22X1_HVT U739 ( .A1(n1318), .A2(n205), .A3(\mem[14][2] ), .A4(n988), .Y(
        n1053) );
  AO21X1_HVT U740 ( .A1(n112), .A2(n1574), .A3(n181), .Y(n1318) );
  AO22X1_HVT U741 ( .A1(n1317), .A2(n205), .A3(\mem[14][3] ), .A4(n987), .Y(
        n1052) );
  AO21X1_HVT U742 ( .A1(n111), .A2(n1572), .A3(n181), .Y(n1317) );
  AO22X1_HVT U743 ( .A1(n1316), .A2(n206), .A3(\mem[14][4] ), .A4(n986), .Y(
        n1051) );
  AO21X1_HVT U744 ( .A1(n113), .A2(n1570), .A3(n181), .Y(n1316) );
  AO22X1_HVT U745 ( .A1(n1315), .A2(n206), .A3(\mem[14][5] ), .A4(n985), .Y(
        n1050) );
  AO21X1_HVT U746 ( .A1(n112), .A2(n1568), .A3(n181), .Y(n1315) );
  AO22X1_HVT U747 ( .A1(n1314), .A2(n206), .A3(\mem[14][6] ), .A4(n984), .Y(
        n1049) );
  AO21X1_HVT U748 ( .A1(n111), .A2(n1566), .A3(n181), .Y(n1314) );
  AO22X1_HVT U749 ( .A1(n1313), .A2(n206), .A3(\mem[14][7] ), .A4(n983), .Y(
        n1048) );
  AO21X1_HVT U750 ( .A1(n113), .A2(n1564), .A3(n181), .Y(n1313) );
  AO22X1_HVT U751 ( .A1(n1312), .A2(n206), .A3(\mem[14][8] ), .A4(n982), .Y(
        n1047) );
  AO21X1_HVT U752 ( .A1(n112), .A2(n1562), .A3(n181), .Y(n1312) );
  AO22X1_HVT U753 ( .A1(n1311), .A2(n206), .A3(\mem[14][9] ), .A4(n981), .Y(
        n1046) );
  AO21X1_HVT U754 ( .A1(n111), .A2(n1560), .A3(n181), .Y(n1311) );
  AO22X1_HVT U755 ( .A1(n1310), .A2(n206), .A3(\mem[14][10] ), .A4(n980), .Y(
        n1045) );
  AO21X1_HVT U756 ( .A1(n113), .A2(n1558), .A3(n182), .Y(n1310) );
  AO22X1_HVT U757 ( .A1(n1309), .A2(n206), .A3(\mem[14][11] ), .A4(n979), .Y(
        n1044) );
  AO21X1_HVT U758 ( .A1(n112), .A2(n1556), .A3(n182), .Y(n1309) );
  AO22X1_HVT U759 ( .A1(n1308), .A2(n206), .A3(\mem[14][12] ), .A4(n978), .Y(
        n1043) );
  AO21X1_HVT U760 ( .A1(n111), .A2(n1554), .A3(n182), .Y(n1308) );
  AO22X1_HVT U761 ( .A1(n1307), .A2(n206), .A3(\mem[14][13] ), .A4(n977), .Y(
        n1042) );
  AO21X1_HVT U762 ( .A1(n113), .A2(n1552), .A3(n182), .Y(n1307) );
  AO22X1_HVT U763 ( .A1(n1306), .A2(n206), .A3(\mem[14][14] ), .A4(n976), .Y(
        n1041) );
  AO21X1_HVT U764 ( .A1(n112), .A2(n1550), .A3(n182), .Y(n1306) );
  AO22X1_HVT U765 ( .A1(n1305), .A2(n206), .A3(\mem[14][15] ), .A4(n975), .Y(
        n1040) );
  AO21X1_HVT U766 ( .A1(n111), .A2(n1548), .A3(n182), .Y(n1305) );
  AND3X1_HVT U767 ( .A1(n1512), .A2(n162), .A3(n1339), .Y(n1320) );
  AND2X1_HVT U768 ( .A1(n154), .A2(n153), .Y(n1512) );
  AO22X1_HVT U769 ( .A1(n1304), .A2(n207), .A3(\mem[15][0] ), .A4(n974), .Y(
        n1039) );
  AO21X1_HVT U770 ( .A1(n108), .A2(n1579), .A3(n182), .Y(n1304) );
  AND2X1_HVT U771 ( .A1(n1302), .A2(n1301), .Y(n1579) );
  AO22X1_HVT U772 ( .A1(n1300), .A2(n207), .A3(\mem[15][1] ), .A4(n973), .Y(
        n1038) );
  AO21X1_HVT U773 ( .A1(n110), .A2(n1576), .A3(n182), .Y(n1300) );
  AND2X1_HVT U774 ( .A1(n1299), .A2(n1302), .Y(n1576) );
  AO22X1_HVT U775 ( .A1(n1298), .A2(n207), .A3(\mem[15][2] ), .A4(n972), .Y(
        n1037) );
  AO21X1_HVT U776 ( .A1(n109), .A2(n1574), .A3(n182), .Y(n1298) );
  AND2X1_HVT U777 ( .A1(n1297), .A2(n1302), .Y(n1574) );
  AO22X1_HVT U778 ( .A1(n1296), .A2(n207), .A3(\mem[15][3] ), .A4(n971), .Y(
        n1036) );
  AO21X1_HVT U779 ( .A1(n108), .A2(n1572), .A3(n182), .Y(n1296) );
  AND2X1_HVT U780 ( .A1(n1295), .A2(n1302), .Y(n1572) );
  AND2X1_HVT U781 ( .A1(n159), .A2(n161), .Y(n1302) );
  AO22X1_HVT U782 ( .A1(n1294), .A2(n207), .A3(\mem[15][4] ), .A4(n970), .Y(
        n1035) );
  AO21X1_HVT U783 ( .A1(n110), .A2(n1570), .A3(n182), .Y(n1294) );
  AND2X1_HVT U784 ( .A1(n1293), .A2(n1301), .Y(n1570) );
  AO22X1_HVT U785 ( .A1(n1292), .A2(n207), .A3(\mem[15][5] ), .A4(n969), .Y(
        n1034) );
  AO21X1_HVT U786 ( .A1(n109), .A2(n1568), .A3(n182), .Y(n1292) );
  AND2X1_HVT U787 ( .A1(n1293), .A2(n1299), .Y(n1568) );
  AO22X1_HVT U788 ( .A1(n1291), .A2(n207), .A3(\mem[15][6] ), .A4(n968), .Y(
        n1033) );
  AO21X1_HVT U789 ( .A1(n108), .A2(n1566), .A3(n182), .Y(n1291) );
  AND2X1_HVT U790 ( .A1(n1293), .A2(n1297), .Y(n1566) );
  AO22X1_HVT U791 ( .A1(n1290), .A2(n207), .A3(\mem[15][7] ), .A4(n967), .Y(
        n1032) );
  AO21X1_HVT U792 ( .A1(n110), .A2(n1564), .A3(n182), .Y(n1290) );
  AND2X1_HVT U793 ( .A1(n1293), .A2(n1295), .Y(n1564) );
  AND2X1_HVT U794 ( .A1(a_addr[2]), .A2(n161), .Y(n1293) );
  AO22X1_HVT U795 ( .A1(n1289), .A2(n207), .A3(\mem[15][8] ), .A4(n966), .Y(
        n1031) );
  AO21X1_HVT U796 ( .A1(n109), .A2(n1562), .A3(n182), .Y(n1289) );
  AND2X1_HVT U797 ( .A1(n1288), .A2(n1301), .Y(n1562) );
  AO22X1_HVT U798 ( .A1(n1287), .A2(n207), .A3(\mem[15][9] ), .A4(n965), .Y(
        n1030) );
  AO21X1_HVT U799 ( .A1(n108), .A2(n1560), .A3(n183), .Y(n1287) );
  AND2X1_HVT U800 ( .A1(n1288), .A2(n1299), .Y(n1560) );
  AO22X1_HVT U801 ( .A1(n1286), .A2(n207), .A3(\mem[15][10] ), .A4(n964), .Y(
        n1029) );
  AO21X1_HVT U802 ( .A1(n110), .A2(n1558), .A3(n183), .Y(n1286) );
  AND2X1_HVT U803 ( .A1(n1288), .A2(n1297), .Y(n1558) );
  AO22X1_HVT U804 ( .A1(n1285), .A2(n207), .A3(\mem[15][11] ), .A4(n963), .Y(
        n1028) );
  AO21X1_HVT U805 ( .A1(n109), .A2(n1556), .A3(n183), .Y(n1285) );
  AND2X1_HVT U806 ( .A1(n1288), .A2(n1295), .Y(n1556) );
  AND2X1_HVT U807 ( .A1(n160), .A2(n159), .Y(n1288) );
  AO22X1_HVT U808 ( .A1(n1284), .A2(n208), .A3(\mem[15][12] ), .A4(n962), .Y(
        n1027) );
  AO21X1_HVT U809 ( .A1(n108), .A2(n1554), .A3(n183), .Y(n1284) );
  AND2X1_HVT U810 ( .A1(n1283), .A2(n1301), .Y(n1554) );
  AND2X1_HVT U811 ( .A1(n156), .A2(n158), .Y(n1301) );
  AO22X1_HVT U812 ( .A1(n1282), .A2(n208), .A3(\mem[15][13] ), .A4(n961), .Y(
        n1026) );
  AO21X1_HVT U813 ( .A1(n110), .A2(n1552), .A3(n183), .Y(n1282) );
  AND2X1_HVT U814 ( .A1(n1283), .A2(n1299), .Y(n1552) );
  AND2X1_HVT U815 ( .A1(a_addr[0]), .A2(n158), .Y(n1299) );
  AO22X1_HVT U816 ( .A1(n1281), .A2(n208), .A3(\mem[15][14] ), .A4(n960), .Y(
        n1025) );
  AO21X1_HVT U817 ( .A1(n109), .A2(n1550), .A3(n183), .Y(n1281) );
  AND2X1_HVT U818 ( .A1(n1283), .A2(n1297), .Y(n1550) );
  AND2X1_HVT U819 ( .A1(n157), .A2(n156), .Y(n1297) );
  AO22X1_HVT U820 ( .A1(n1280), .A2(n208), .A3(\mem[15][15] ), .A4(n959), .Y(
        n1024) );
  AO21X1_HVT U821 ( .A1(n108), .A2(n1548), .A3(n183), .Y(n1280) );
  AND2X1_HVT U822 ( .A1(n1283), .A2(n1295), .Y(n1548) );
  AND2X1_HVT U823 ( .A1(n157), .A2(a_addr[0]), .Y(n1295) );
  AND2X1_HVT U824 ( .A1(n160), .A2(a_addr[2]), .Y(n1283) );
  AND3X1_HVT U825 ( .A1(n1495), .A2(n163), .A3(n1339), .Y(n1303) );
  AND2X1_HVT U826 ( .A1(a_din[3]), .A2(a_din[2]), .Y(n1339) );
  AND2X1_HVT U827 ( .A1(n154), .A2(a_din[0]), .Y(n1495) );
  AND2X1_HVT U3 ( .A1(n1546), .A2(n1512), .Y(n1) );
  INVX0_HVT U4 ( .A(n1529), .Y(n7) );
  INVX0_HVT U5 ( .A(n1546), .Y(n6) );
  INVX0_HVT U6 ( .A(N17), .Y(n2) );
  INVX1_HVT U7 ( .A(n2), .Y(n3) );
  INVX1_HVT U8 ( .A(n164), .Y(n4) );
  INVX0_HVT U9 ( .A(n8), .Y(n5) );
  NAND2X0_HVT U10 ( .A1(n1), .A2(n4), .Y(n8) );
  INVX0_HVT U11 ( .A(n8), .Y(n147) );
  INVX0_HVT U12 ( .A(n8), .Y(n146) );
  OR3X1_HVT U13 ( .A1(n6), .A2(n164), .A3(n7), .Y(n10) );
  INVX1_HVT U14 ( .A(n164), .Y(n163) );
  IBUFFX2_HVT U15 ( .A(write), .Y(n164) );
  INVX1_HVT U16 ( .A(n187), .Y(n193) );
  INVX1_HVT U17 ( .A(n187), .Y(n194) );
  INVX1_HVT U18 ( .A(n187), .Y(n195) );
  INVX1_HVT U19 ( .A(n187), .Y(n196) );
  INVX1_HVT U20 ( .A(n165), .Y(n197) );
  INVX1_HVT U21 ( .A(n187), .Y(n198) );
  INVX1_HVT U22 ( .A(n183), .Y(n199) );
  INVX1_HVT U23 ( .A(n165), .Y(n200) );
  INVX1_HVT U24 ( .A(n187), .Y(n201) );
  INVX1_HVT U25 ( .A(n183), .Y(n202) );
  INVX1_HVT U26 ( .A(n165), .Y(n203) );
  INVX1_HVT U27 ( .A(n165), .Y(n204) );
  INVX1_HVT U28 ( .A(n165), .Y(n205) );
  INVX1_HVT U29 ( .A(n165), .Y(n206) );
  INVX1_HVT U30 ( .A(n165), .Y(n207) );
  INVX1_HVT U31 ( .A(n165), .Y(n208) );
  INVX1_HVT U32 ( .A(n166), .Y(n189) );
  INVX1_HVT U33 ( .A(n166), .Y(n190) );
  INVX1_HVT U34 ( .A(n166), .Y(n191) );
  INVX1_HVT U35 ( .A(n166), .Y(n192) );
  INVX1_HVT U36 ( .A(n164), .Y(n162) );
  INVX1_HVT U37 ( .A(n188), .Y(n165) );
  INVX1_HVT U38 ( .A(n186), .Y(n171) );
  INVX1_HVT U39 ( .A(n185), .Y(n177) );
  INVX1_HVT U40 ( .A(n184), .Y(n182) );
  INVX1_HVT U41 ( .A(n186), .Y(n167) );
  INVX1_HVT U42 ( .A(n186), .Y(n168) );
  INVX1_HVT U43 ( .A(n186), .Y(n169) );
  INVX1_HVT U44 ( .A(n186), .Y(n170) );
  INVX1_HVT U45 ( .A(n185), .Y(n172) );
  INVX1_HVT U46 ( .A(n185), .Y(n173) );
  INVX1_HVT U47 ( .A(n185), .Y(n174) );
  INVX1_HVT U48 ( .A(n185), .Y(n175) );
  INVX1_HVT U49 ( .A(n185), .Y(n176) );
  INVX1_HVT U50 ( .A(n184), .Y(n178) );
  INVX1_HVT U51 ( .A(n184), .Y(n179) );
  INVX1_HVT U52 ( .A(n184), .Y(n180) );
  INVX1_HVT U53 ( .A(n184), .Y(n181) );
  INVX1_HVT U54 ( .A(n186), .Y(n166) );
  INVX1_HVT U55 ( .A(n184), .Y(n183) );
  INVX1_HVT U56 ( .A(n187), .Y(n186) );
  INVX1_HVT U57 ( .A(n187), .Y(n185) );
  INVX1_HVT U58 ( .A(n187), .Y(n184) );
  NBUFFX2_HVT U59 ( .A(n1578), .Y(n150) );
  NBUFFX2_HVT U60 ( .A(n1578), .Y(n152) );
  NBUFFX2_HVT U61 ( .A(n1578), .Y(n151) );
  INVX1_HVT U62 ( .A(n188), .Y(n187) );
  INVX1_HVT U63 ( .A(rst), .Y(n188) );
  INVX1_HVT U64 ( .A(n161), .Y(n160) );
  INVX1_HVT U65 ( .A(n158), .Y(n157) );
  NBUFFX2_HVT U66 ( .A(n1389), .Y(n123) );
  NBUFFX2_HVT U67 ( .A(n1320), .Y(n111) );
  NBUFFX2_HVT U68 ( .A(n1493), .Y(n141) );
  NBUFFX2_HVT U69 ( .A(n1458), .Y(n135) );
  NBUFFX2_HVT U70 ( .A(n1424), .Y(n129) );
  NBUFFX2_HVT U71 ( .A(n1355), .Y(n117) );
  NBUFFX2_HVT U72 ( .A(n1389), .Y(n125) );
  NBUFFX2_HVT U73 ( .A(n1389), .Y(n124) );
  NBUFFX2_HVT U74 ( .A(n1320), .Y(n113) );
  NBUFFX2_HVT U75 ( .A(n1320), .Y(n112) );
  NBUFFX2_HVT U76 ( .A(n1493), .Y(n143) );
  NBUFFX2_HVT U77 ( .A(n1493), .Y(n142) );
  NBUFFX2_HVT U78 ( .A(n1458), .Y(n137) );
  NBUFFX2_HVT U79 ( .A(n1458), .Y(n136) );
  NBUFFX2_HVT U80 ( .A(n1424), .Y(n131) );
  NBUFFX2_HVT U81 ( .A(n1424), .Y(n130) );
  NBUFFX2_HVT U82 ( .A(n1355), .Y(n119) );
  NBUFFX2_HVT U83 ( .A(n1355), .Y(n118) );
  NBUFFX2_HVT U84 ( .A(n1303), .Y(n108) );
  NBUFFX2_HVT U85 ( .A(n1475), .Y(n138) );
  NBUFFX2_HVT U86 ( .A(n1406), .Y(n126) );
  NBUFFX2_HVT U87 ( .A(n1441), .Y(n132) );
  NBUFFX2_HVT U88 ( .A(n1372), .Y(n120) );
  NBUFFX2_HVT U89 ( .A(n1337), .Y(n114) );
  NBUFFX2_HVT U90 ( .A(n1303), .Y(n110) );
  NBUFFX2_HVT U91 ( .A(n1303), .Y(n109) );
  NBUFFX2_HVT U92 ( .A(n1475), .Y(n140) );
  NBUFFX2_HVT U93 ( .A(n1475), .Y(n139) );
  NBUFFX2_HVT U94 ( .A(n1441), .Y(n134) );
  NBUFFX2_HVT U95 ( .A(n1441), .Y(n133) );
  NBUFFX2_HVT U96 ( .A(n1372), .Y(n122) );
  NBUFFX2_HVT U97 ( .A(n1372), .Y(n121) );
  NBUFFX2_HVT U98 ( .A(n1406), .Y(n128) );
  NBUFFX2_HVT U99 ( .A(n1406), .Y(n127) );
  NBUFFX2_HVT U100 ( .A(n1337), .Y(n116) );
  NBUFFX2_HVT U101 ( .A(n1337), .Y(n115) );
  INVX1_HVT U102 ( .A(n9), .Y(n145) );
  INVX1_HVT U103 ( .A(n9), .Y(n144) );
  INVX1_HVT U104 ( .A(n10), .Y(n149) );
  INVX1_HVT U105 ( .A(n10), .Y(n148) );
  INVX1_HVT U106 ( .A(a_addr[1]), .Y(n158) );
  INVX1_HVT U107 ( .A(a_addr[3]), .Y(n161) );
  INVX1_HVT U108 ( .A(a_addr[2]), .Y(n159) );
  INVX1_HVT U109 ( .A(a_addr[0]), .Y(n156) );
  NBUFFX2_HVT U110 ( .A(n86), .Y(n106) );
  NBUFFX2_HVT U111 ( .A(n86), .Y(n103) );
  NBUFFX2_HVT U112 ( .A(n85), .Y(n100) );
  NBUFFX2_HVT U113 ( .A(n84), .Y(n97) );
  NBUFFX2_HVT U114 ( .A(n83), .Y(n94) );
  NBUFFX2_HVT U115 ( .A(n85), .Y(n107) );
  NBUFFX2_HVT U116 ( .A(n86), .Y(n104) );
  NBUFFX2_HVT U117 ( .A(n85), .Y(n101) );
  NBUFFX2_HVT U118 ( .A(n84), .Y(n98) );
  NBUFFX2_HVT U119 ( .A(n83), .Y(n95) );
  NBUFFX2_HVT U120 ( .A(n84), .Y(n105) );
  NBUFFX2_HVT U121 ( .A(n86), .Y(n102) );
  NBUFFX2_HVT U122 ( .A(n85), .Y(n99) );
  NBUFFX2_HVT U123 ( .A(n84), .Y(n96) );
  NBUFFX2_HVT U124 ( .A(n83), .Y(n93) );
  NAND3X0_HVT U125 ( .A1(n1546), .A2(n163), .A3(n1495), .Y(n9) );
  INVX1_HVT U126 ( .A(n75), .Y(n81) );
  INVX1_HVT U127 ( .A(n75), .Y(n80) );
  INVX1_HVT U128 ( .A(n75), .Y(n79) );
  INVX1_HVT U129 ( .A(n75), .Y(n78) );
  INVX1_HVT U130 ( .A(n75), .Y(n77) );
  INVX1_HVT U131 ( .A(n75), .Y(n76) );
  INVX1_HVT U132 ( .A(n89), .Y(n87) );
  INVX1_HVT U133 ( .A(n89), .Y(n88) );
  INVX1_HVT U134 ( .A(n155), .Y(n154) );
  INVX1_HVT U135 ( .A(n92), .Y(n90) );
  INVX1_HVT U136 ( .A(n92), .Y(n91) );
  INVX0_HVT U137 ( .A(a_din[0]), .Y(n153) );
  NBUFFX2_HVT U138 ( .A(n3), .Y(n86) );
  NBUFFX2_HVT U139 ( .A(n3), .Y(n85) );
  NBUFFX2_HVT U140 ( .A(n3), .Y(n84) );
  NBUFFX2_HVT U141 ( .A(n3), .Y(n83) );
  NBUFFX2_HVT U142 ( .A(n3), .Y(n82) );
  INVX1_HVT U143 ( .A(N18), .Y(n75) );
  INVX0_HVT U144 ( .A(N19), .Y(n89) );
  INVX0_HVT U145 ( .A(a_din[1]), .Y(n155) );
  INVX0_HVT U146 ( .A(N20), .Y(n92) );
  MUX41X1_HVT U147 ( .A1(\mem[12][0] ), .A3(\mem[14][0] ), .A2(\mem[13][0] ), 
        .A4(\mem[15][0] ), .S0(n81), .S1(n106), .Y(n11) );
  MUX41X1_HVT U148 ( .A1(\mem[8][0] ), .A3(\mem[10][0] ), .A2(\mem[9][0] ), 
        .A4(\mem[11][0] ), .S0(n81), .S1(n105), .Y(n12) );
  MUX41X1_HVT U149 ( .A1(\mem[4][0] ), .A3(\mem[6][0] ), .A2(\mem[5][0] ), 
        .A4(\mem[7][0] ), .S0(n81), .S1(n106), .Y(n13) );
  MUX41X1_HVT U150 ( .A1(\mem[0][0] ), .A3(\mem[2][0] ), .A2(\mem[1][0] ), 
        .A4(\mem[3][0] ), .S0(n81), .S1(n105), .Y(n14) );
  MUX41X1_HVT U151 ( .A1(n14), .A3(n12), .A2(n13), .A4(n11), .S0(n90), .S1(n87), .Y(N554) );
  MUX41X1_HVT U152 ( .A1(\mem[12][1] ), .A3(\mem[14][1] ), .A2(\mem[13][1] ), 
        .A4(\mem[15][1] ), .S0(n81), .S1(n106), .Y(n15) );
  MUX41X1_HVT U153 ( .A1(\mem[8][1] ), .A3(\mem[10][1] ), .A2(\mem[9][1] ), 
        .A4(\mem[11][1] ), .S0(n81), .S1(n105), .Y(n16) );
  MUX41X1_HVT U154 ( .A1(\mem[4][1] ), .A3(\mem[6][1] ), .A2(\mem[5][1] ), 
        .A4(\mem[7][1] ), .S0(n81), .S1(n106), .Y(n17) );
  MUX41X1_HVT U155 ( .A1(\mem[0][1] ), .A3(\mem[2][1] ), .A2(\mem[1][1] ), 
        .A4(\mem[3][1] ), .S0(n81), .S1(n105), .Y(n18) );
  MUX41X1_HVT U156 ( .A1(n18), .A3(n16), .A2(n17), .A4(n15), .S0(n90), .S1(n87), .Y(N553) );
  MUX41X1_HVT U157 ( .A1(\mem[12][2] ), .A3(\mem[14][2] ), .A2(\mem[13][2] ), 
        .A4(\mem[15][2] ), .S0(n81), .S1(n107), .Y(n19) );
  MUX41X1_HVT U158 ( .A1(\mem[8][2] ), .A3(\mem[10][2] ), .A2(\mem[9][2] ), 
        .A4(\mem[11][2] ), .S0(n81), .S1(n107), .Y(n20) );
  MUX41X1_HVT U159 ( .A1(\mem[4][2] ), .A3(\mem[6][2] ), .A2(\mem[5][2] ), 
        .A4(\mem[7][2] ), .S0(n81), .S1(n107), .Y(n21) );
  MUX41X1_HVT U160 ( .A1(\mem[0][2] ), .A3(\mem[2][2] ), .A2(\mem[1][2] ), 
        .A4(\mem[3][2] ), .S0(n81), .S1(n107), .Y(n22) );
  MUX41X1_HVT U161 ( .A1(n22), .A3(n20), .A2(n21), .A4(n19), .S0(n90), .S1(n87), .Y(N552) );
  MUX41X1_HVT U162 ( .A1(\mem[12][3] ), .A3(\mem[14][3] ), .A2(\mem[13][3] ), 
        .A4(\mem[15][3] ), .S0(n80), .S1(n103), .Y(n23) );
  MUX41X1_HVT U163 ( .A1(\mem[8][3] ), .A3(\mem[10][3] ), .A2(\mem[9][3] ), 
        .A4(\mem[11][3] ), .S0(n80), .S1(n102), .Y(n24) );
  MUX41X1_HVT U164 ( .A1(\mem[4][3] ), .A3(\mem[6][3] ), .A2(\mem[5][3] ), 
        .A4(\mem[7][3] ), .S0(n80), .S1(n103), .Y(n25) );
  MUX41X1_HVT U165 ( .A1(\mem[0][3] ), .A3(\mem[2][3] ), .A2(\mem[1][3] ), 
        .A4(\mem[3][3] ), .S0(n80), .S1(n102), .Y(n26) );
  MUX41X1_HVT U166 ( .A1(n26), .A3(n24), .A2(n25), .A4(n23), .S0(n90), .S1(n87), .Y(N551) );
  MUX41X1_HVT U167 ( .A1(\mem[12][4] ), .A3(\mem[14][4] ), .A2(\mem[13][4] ), 
        .A4(\mem[15][4] ), .S0(n80), .S1(n103), .Y(n27) );
  MUX41X1_HVT U168 ( .A1(\mem[8][4] ), .A3(\mem[10][4] ), .A2(\mem[9][4] ), 
        .A4(\mem[11][4] ), .S0(n80), .S1(n102), .Y(n28) );
  MUX41X1_HVT U169 ( .A1(\mem[4][4] ), .A3(\mem[6][4] ), .A2(\mem[5][4] ), 
        .A4(\mem[7][4] ), .S0(n80), .S1(n103), .Y(n29) );
  MUX41X1_HVT U170 ( .A1(\mem[0][4] ), .A3(\mem[2][4] ), .A2(\mem[1][4] ), 
        .A4(\mem[3][4] ), .S0(n80), .S1(n102), .Y(n30) );
  MUX41X1_HVT U171 ( .A1(n30), .A3(n28), .A2(n29), .A4(n27), .S0(n90), .S1(n87), .Y(N550) );
  MUX41X1_HVT U172 ( .A1(\mem[12][5] ), .A3(\mem[14][5] ), .A2(\mem[13][5] ), 
        .A4(\mem[15][5] ), .S0(n80), .S1(n104), .Y(n31) );
  MUX41X1_HVT U173 ( .A1(\mem[8][5] ), .A3(\mem[10][5] ), .A2(\mem[9][5] ), 
        .A4(\mem[11][5] ), .S0(n80), .S1(n104), .Y(n32) );
  MUX41X1_HVT U174 ( .A1(\mem[4][5] ), .A3(\mem[6][5] ), .A2(\mem[5][5] ), 
        .A4(\mem[7][5] ), .S0(n80), .S1(n104), .Y(n33) );
  MUX41X1_HVT U175 ( .A1(\mem[0][5] ), .A3(\mem[2][5] ), .A2(\mem[1][5] ), 
        .A4(\mem[3][5] ), .S0(n80), .S1(n104), .Y(n34) );
  MUX41X1_HVT U176 ( .A1(n34), .A3(n32), .A2(n33), .A4(n31), .S0(n90), .S1(n87), .Y(N549) );
  MUX41X1_HVT U177 ( .A1(\mem[12][6] ), .A3(\mem[14][6] ), .A2(\mem[13][6] ), 
        .A4(\mem[15][6] ), .S0(n79), .S1(n100), .Y(n35) );
  MUX41X1_HVT U178 ( .A1(\mem[8][6] ), .A3(\mem[10][6] ), .A2(\mem[9][6] ), 
        .A4(\mem[11][6] ), .S0(n79), .S1(n99), .Y(n36) );
  MUX41X1_HVT U179 ( .A1(\mem[4][6] ), .A3(\mem[6][6] ), .A2(\mem[5][6] ), 
        .A4(\mem[7][6] ), .S0(n79), .S1(n100), .Y(n37) );
  MUX41X1_HVT U180 ( .A1(\mem[0][6] ), .A3(\mem[2][6] ), .A2(\mem[1][6] ), 
        .A4(\mem[3][6] ), .S0(n79), .S1(n99), .Y(n38) );
  MUX41X1_HVT U181 ( .A1(n38), .A3(n36), .A2(n37), .A4(n35), .S0(n90), .S1(n87), .Y(N548) );
  MUX41X1_HVT U182 ( .A1(\mem[12][7] ), .A3(\mem[14][7] ), .A2(\mem[13][7] ), 
        .A4(\mem[15][7] ), .S0(n79), .S1(n100), .Y(n39) );
  MUX41X1_HVT U183 ( .A1(\mem[8][7] ), .A3(\mem[10][7] ), .A2(\mem[9][7] ), 
        .A4(\mem[11][7] ), .S0(n79), .S1(n99), .Y(n40) );
  MUX41X1_HVT U184 ( .A1(\mem[4][7] ), .A3(\mem[6][7] ), .A2(\mem[5][7] ), 
        .A4(\mem[7][7] ), .S0(n79), .S1(n100), .Y(n41) );
  MUX41X1_HVT U185 ( .A1(\mem[0][7] ), .A3(\mem[2][7] ), .A2(\mem[1][7] ), 
        .A4(\mem[3][7] ), .S0(n79), .S1(n99), .Y(n42) );
  MUX41X1_HVT U186 ( .A1(n42), .A3(n40), .A2(n41), .A4(n39), .S0(n90), .S1(n87), .Y(N547) );
  MUX41X1_HVT U187 ( .A1(\mem[12][8] ), .A3(\mem[14][8] ), .A2(\mem[13][8] ), 
        .A4(\mem[15][8] ), .S0(n79), .S1(n101), .Y(n43) );
  MUX41X1_HVT U188 ( .A1(\mem[8][8] ), .A3(\mem[10][8] ), .A2(\mem[9][8] ), 
        .A4(\mem[11][8] ), .S0(n79), .S1(n101), .Y(n44) );
  MUX41X1_HVT U189 ( .A1(\mem[4][8] ), .A3(\mem[6][8] ), .A2(\mem[5][8] ), 
        .A4(\mem[7][8] ), .S0(n79), .S1(n101), .Y(n45) );
  MUX41X1_HVT U190 ( .A1(\mem[0][8] ), .A3(\mem[2][8] ), .A2(\mem[1][8] ), 
        .A4(\mem[3][8] ), .S0(n79), .S1(n101), .Y(n46) );
  MUX41X1_HVT U191 ( .A1(n46), .A3(n44), .A2(n45), .A4(n43), .S0(n91), .S1(n88), .Y(N546) );
  MUX41X1_HVT U192 ( .A1(\mem[12][9] ), .A3(\mem[14][9] ), .A2(\mem[13][9] ), 
        .A4(\mem[15][9] ), .S0(n78), .S1(n97), .Y(n47) );
  MUX41X1_HVT U193 ( .A1(\mem[8][9] ), .A3(\mem[10][9] ), .A2(\mem[9][9] ), 
        .A4(\mem[11][9] ), .S0(n78), .S1(n96), .Y(n48) );
  MUX41X1_HVT U194 ( .A1(\mem[4][9] ), .A3(\mem[6][9] ), .A2(\mem[5][9] ), 
        .A4(\mem[7][9] ), .S0(n78), .S1(n97), .Y(n49) );
  MUX41X1_HVT U195 ( .A1(\mem[0][9] ), .A3(\mem[2][9] ), .A2(\mem[1][9] ), 
        .A4(\mem[3][9] ), .S0(n78), .S1(n96), .Y(n50) );
  MUX41X1_HVT U196 ( .A1(n50), .A3(n48), .A2(n49), .A4(n47), .S0(n91), .S1(n88), .Y(N545) );
  MUX41X1_HVT U197 ( .A1(\mem[12][10] ), .A3(\mem[14][10] ), .A2(\mem[13][10] ), .A4(\mem[15][10] ), .S0(n78), .S1(n97), .Y(n51) );
  MUX41X1_HVT U198 ( .A1(\mem[8][10] ), .A3(\mem[10][10] ), .A2(\mem[9][10] ), 
        .A4(\mem[11][10] ), .S0(n78), .S1(n96), .Y(n52) );
  MUX41X1_HVT U199 ( .A1(\mem[4][10] ), .A3(\mem[6][10] ), .A2(\mem[5][10] ), 
        .A4(\mem[7][10] ), .S0(n78), .S1(n97), .Y(n53) );
  MUX41X1_HVT U200 ( .A1(\mem[0][10] ), .A3(\mem[2][10] ), .A2(\mem[1][10] ), 
        .A4(\mem[3][10] ), .S0(n78), .S1(n96), .Y(n54) );
  MUX41X1_HVT U201 ( .A1(n54), .A3(n52), .A2(n53), .A4(n51), .S0(n91), .S1(n88), .Y(N544) );
  MUX41X1_HVT U202 ( .A1(\mem[12][11] ), .A3(\mem[14][11] ), .A2(\mem[13][11] ), .A4(\mem[15][11] ), .S0(n78), .S1(n98), .Y(n55) );
  MUX41X1_HVT U203 ( .A1(\mem[8][11] ), .A3(\mem[10][11] ), .A2(\mem[9][11] ), 
        .A4(\mem[11][11] ), .S0(n78), .S1(n98), .Y(n56) );
  MUX41X1_HVT U204 ( .A1(\mem[4][11] ), .A3(\mem[6][11] ), .A2(\mem[5][11] ), 
        .A4(\mem[7][11] ), .S0(n78), .S1(n98), .Y(n57) );
  MUX41X1_HVT U205 ( .A1(\mem[0][11] ), .A3(\mem[2][11] ), .A2(\mem[1][11] ), 
        .A4(\mem[3][11] ), .S0(n78), .S1(n98), .Y(n58) );
  MUX41X1_HVT U206 ( .A1(n58), .A3(n56), .A2(n57), .A4(n55), .S0(n91), .S1(n88), .Y(N543) );
  MUX41X1_HVT U207 ( .A1(\mem[12][12] ), .A3(\mem[14][12] ), .A2(\mem[13][12] ), .A4(\mem[15][12] ), .S0(n77), .S1(n94), .Y(n59) );
  MUX41X1_HVT U208 ( .A1(\mem[8][12] ), .A3(\mem[10][12] ), .A2(\mem[9][12] ), 
        .A4(\mem[11][12] ), .S0(n77), .S1(n93), .Y(n60) );
  MUX41X1_HVT U209 ( .A1(\mem[4][12] ), .A3(\mem[6][12] ), .A2(\mem[5][12] ), 
        .A4(\mem[7][12] ), .S0(n77), .S1(n94), .Y(n61) );
  MUX41X1_HVT U210 ( .A1(\mem[0][12] ), .A3(\mem[2][12] ), .A2(\mem[1][12] ), 
        .A4(\mem[3][12] ), .S0(n77), .S1(n93), .Y(n62) );
  MUX41X1_HVT U211 ( .A1(n62), .A3(n60), .A2(n61), .A4(n59), .S0(n91), .S1(n88), .Y(N542) );
  MUX41X1_HVT U212 ( .A1(\mem[12][13] ), .A3(\mem[14][13] ), .A2(\mem[13][13] ), .A4(\mem[15][13] ), .S0(n77), .S1(n94), .Y(n63) );
  MUX41X1_HVT U213 ( .A1(\mem[8][13] ), .A3(\mem[10][13] ), .A2(\mem[9][13] ), 
        .A4(\mem[11][13] ), .S0(n77), .S1(n93), .Y(n64) );
  MUX41X1_HVT U214 ( .A1(\mem[4][13] ), .A3(\mem[6][13] ), .A2(\mem[5][13] ), 
        .A4(\mem[7][13] ), .S0(n77), .S1(n94), .Y(n65) );
  MUX41X1_HVT U215 ( .A1(\mem[0][13] ), .A3(\mem[2][13] ), .A2(\mem[1][13] ), 
        .A4(\mem[3][13] ), .S0(n77), .S1(n93), .Y(n66) );
  MUX41X1_HVT U216 ( .A1(n66), .A3(n64), .A2(n65), .A4(n63), .S0(n91), .S1(n88), .Y(N541) );
  MUX41X1_HVT U217 ( .A1(\mem[12][14] ), .A3(\mem[14][14] ), .A2(\mem[13][14] ), .A4(\mem[15][14] ), .S0(n77), .S1(n95), .Y(n67) );
  MUX41X1_HVT U218 ( .A1(\mem[8][14] ), .A3(\mem[10][14] ), .A2(\mem[9][14] ), 
        .A4(\mem[11][14] ), .S0(n77), .S1(n95), .Y(n68) );
  MUX41X1_HVT U219 ( .A1(\mem[4][14] ), .A3(\mem[6][14] ), .A2(\mem[5][14] ), 
        .A4(\mem[7][14] ), .S0(n77), .S1(n95), .Y(n69) );
  MUX41X1_HVT U220 ( .A1(\mem[0][14] ), .A3(\mem[2][14] ), .A2(\mem[1][14] ), 
        .A4(\mem[3][14] ), .S0(n77), .S1(n95), .Y(n70) );
  MUX41X1_HVT U221 ( .A1(n70), .A3(n68), .A2(n69), .A4(n67), .S0(n91), .S1(n88), .Y(N540) );
  MUX41X1_HVT U222 ( .A1(\mem[12][15] ), .A3(\mem[14][15] ), .A2(\mem[13][15] ), .A4(\mem[15][15] ), .S0(n76), .S1(n82), .Y(n71) );
  MUX41X1_HVT U223 ( .A1(\mem[8][15] ), .A3(\mem[10][15] ), .A2(\mem[9][15] ), 
        .A4(\mem[11][15] ), .S0(n76), .S1(n82), .Y(n72) );
  MUX41X1_HVT U224 ( .A1(\mem[4][15] ), .A3(\mem[6][15] ), .A2(\mem[5][15] ), 
        .A4(\mem[7][15] ), .S0(n76), .S1(n82), .Y(n73) );
  MUX41X1_HVT U225 ( .A1(\mem[0][15] ), .A3(\mem[2][15] ), .A2(\mem[1][15] ), 
        .A4(\mem[3][15] ), .S0(n76), .S1(n82), .Y(n74) );
  MUX41X1_HVT U226 ( .A1(n74), .A3(n72), .A2(n73), .A4(n71), .S0(n91), .S1(n88), .Y(N539) );
  INVX0_HVT U227 ( .A(n1426), .Y(n209) );
  INVX0_HVT U228 ( .A(n1427), .Y(n210) );
  INVX0_HVT U229 ( .A(n1428), .Y(n211) );
  INVX0_HVT U230 ( .A(n1429), .Y(n212) );
  INVX0_HVT U231 ( .A(n1430), .Y(n213) );
  INVX0_HVT U232 ( .A(n1431), .Y(n214) );
  INVX0_HVT U233 ( .A(n1432), .Y(n215) );
  INVX0_HVT U234 ( .A(n1433), .Y(n216) );
  INVX0_HVT U235 ( .A(n1434), .Y(n217) );
  INVX0_HVT U236 ( .A(n1435), .Y(n218) );
  INVX0_HVT U237 ( .A(n1436), .Y(n219) );
  INVX0_HVT U238 ( .A(n1437), .Y(n220) );
  INVX0_HVT U239 ( .A(n1438), .Y(n221) );
  INVX0_HVT U240 ( .A(n1439), .Y(n222) );
  INVX0_HVT U241 ( .A(n1440), .Y(n223) );
  INVX0_HVT U242 ( .A(n1442), .Y(n224) );
  INVX0_HVT U243 ( .A(n1443), .Y(n225) );
  INVX0_HVT U244 ( .A(n1444), .Y(n226) );
  INVX0_HVT U245 ( .A(n1445), .Y(n227) );
  INVX0_HVT U246 ( .A(n1446), .Y(n228) );
  INVX0_HVT U247 ( .A(n1447), .Y(n229) );
  INVX0_HVT U248 ( .A(n1448), .Y(n230) );
  INVX0_HVT U249 ( .A(n1449), .Y(n231) );
  INVX0_HVT U250 ( .A(n1450), .Y(n232) );
  INVX0_HVT U251 ( .A(n1451), .Y(n233) );
  INVX0_HVT U252 ( .A(n1452), .Y(n234) );
  INVX0_HVT U253 ( .A(n1453), .Y(n235) );
  INVX0_HVT U254 ( .A(n1454), .Y(n236) );
  INVX0_HVT U255 ( .A(n1455), .Y(n237) );
  INVX0_HVT U256 ( .A(n1456), .Y(n238) );
  INVX0_HVT U257 ( .A(n1457), .Y(n239) );
  INVX0_HVT U258 ( .A(n1459), .Y(n240) );
  INVX0_HVT U259 ( .A(n1460), .Y(n241) );
  INVX0_HVT U260 ( .A(n1461), .Y(n242) );
  INVX0_HVT U261 ( .A(n1462), .Y(n243) );
  INVX0_HVT U262 ( .A(n1463), .Y(n244) );
  INVX0_HVT U263 ( .A(n1464), .Y(n245) );
  INVX0_HVT U264 ( .A(n1465), .Y(n246) );
  INVX0_HVT U265 ( .A(n1466), .Y(n247) );
  INVX0_HVT U266 ( .A(n1467), .Y(n248) );
  INVX0_HVT U267 ( .A(n1468), .Y(n249) );
  INVX0_HVT U333 ( .A(n1469), .Y(n250) );
  INVX0_HVT U366 ( .A(n1470), .Y(n251) );
  INVX0_HVT U399 ( .A(n1471), .Y(n252) );
  INVX0_HVT U828 ( .A(n1472), .Y(n253) );
  INVX0_HVT U829 ( .A(n1473), .Y(n254) );
  INVX0_HVT U830 ( .A(n1474), .Y(n255) );
  INVX0_HVT U831 ( .A(n1476), .Y(n256) );
  INVX0_HVT U832 ( .A(n1478), .Y(n257) );
  INVX0_HVT U833 ( .A(n1479), .Y(n258) );
  INVX0_HVT U834 ( .A(n1480), .Y(n259) );
  INVX0_HVT U835 ( .A(n1481), .Y(n260) );
  INVX0_HVT U836 ( .A(n1482), .Y(n261) );
  INVX0_HVT U837 ( .A(n1483), .Y(n262) );
  INVX0_HVT U838 ( .A(n1484), .Y(n263) );
  INVX0_HVT U839 ( .A(n1485), .Y(n264) );
  INVX0_HVT U840 ( .A(n1486), .Y(n265) );
  INVX0_HVT U841 ( .A(n1487), .Y(n302) );
  INVX0_HVT U842 ( .A(n1488), .Y(n320) );
  INVX0_HVT U843 ( .A(n1489), .Y(n338) );
  INVX0_HVT U844 ( .A(n1490), .Y(n826) );
  INVX0_HVT U845 ( .A(n1491), .Y(n827) );
  INVX0_HVT U846 ( .A(n1492), .Y(n828) );
  INVX0_HVT U847 ( .A(n1494), .Y(n829) );
  INVX0_HVT U848 ( .A(n1496), .Y(n830) );
  INVX0_HVT U849 ( .A(n1497), .Y(n831) );
  INVX0_HVT U850 ( .A(n1498), .Y(n832) );
  INVX0_HVT U851 ( .A(n1499), .Y(n833) );
  INVX0_HVT U852 ( .A(n1500), .Y(n834) );
  INVX0_HVT U853 ( .A(n1501), .Y(n835) );
  INVX0_HVT U854 ( .A(n1502), .Y(n836) );
  INVX0_HVT U855 ( .A(n1503), .Y(n837) );
  INVX0_HVT U856 ( .A(n1504), .Y(n838) );
  INVX0_HVT U857 ( .A(n1505), .Y(n839) );
  INVX0_HVT U858 ( .A(n1506), .Y(n840) );
  INVX0_HVT U859 ( .A(n1507), .Y(n841) );
  INVX0_HVT U860 ( .A(n1508), .Y(n842) );
  INVX0_HVT U861 ( .A(n1509), .Y(n843) );
  INVX0_HVT U862 ( .A(n1510), .Y(n844) );
  INVX0_HVT U863 ( .A(n1511), .Y(n845) );
  INVX0_HVT U864 ( .A(n1513), .Y(n846) );
  INVX0_HVT U865 ( .A(n1514), .Y(n847) );
  INVX0_HVT U866 ( .A(n1515), .Y(n848) );
  INVX0_HVT U867 ( .A(n1516), .Y(n849) );
  INVX0_HVT U868 ( .A(n1517), .Y(n850) );
  INVX0_HVT U869 ( .A(n1518), .Y(n851) );
  INVX0_HVT U870 ( .A(n1519), .Y(n852) );
  INVX0_HVT U871 ( .A(n1520), .Y(n853) );
  INVX0_HVT U872 ( .A(n1521), .Y(n854) );
  INVX0_HVT U873 ( .A(n1522), .Y(n855) );
  INVX0_HVT U874 ( .A(n1523), .Y(n856) );
  INVX0_HVT U875 ( .A(n1524), .Y(n857) );
  INVX0_HVT U876 ( .A(n1525), .Y(n858) );
  INVX0_HVT U877 ( .A(n1526), .Y(n859) );
  INVX0_HVT U878 ( .A(n1527), .Y(n860) );
  INVX0_HVT U879 ( .A(n1528), .Y(n861) );
  INVX0_HVT U880 ( .A(n1530), .Y(n862) );
  INVX0_HVT U881 ( .A(n1531), .Y(n863) );
  INVX0_HVT U882 ( .A(n1532), .Y(n864) );
  INVX0_HVT U883 ( .A(n1533), .Y(n865) );
  INVX0_HVT U884 ( .A(n1534), .Y(n866) );
  INVX0_HVT U885 ( .A(n1535), .Y(n867) );
  INVX0_HVT U886 ( .A(n1536), .Y(n868) );
  INVX0_HVT U887 ( .A(n1537), .Y(n869) );
  INVX0_HVT U888 ( .A(n1538), .Y(n870) );
  INVX0_HVT U889 ( .A(n1539), .Y(n871) );
  INVX0_HVT U890 ( .A(n1540), .Y(n872) );
  INVX0_HVT U891 ( .A(n1541), .Y(n873) );
  INVX0_HVT U892 ( .A(n1542), .Y(n874) );
  INVX0_HVT U893 ( .A(n1543), .Y(n875) );
  INVX0_HVT U894 ( .A(n1544), .Y(n876) );
  INVX0_HVT U895 ( .A(n1545), .Y(n877) );
  INVX0_HVT U896 ( .A(n1549), .Y(n878) );
  INVX0_HVT U897 ( .A(n1551), .Y(n879) );
  INVX0_HVT U898 ( .A(n1553), .Y(n880) );
  INVX0_HVT U899 ( .A(n1555), .Y(n881) );
  INVX0_HVT U900 ( .A(n1557), .Y(n882) );
  INVX0_HVT U901 ( .A(n1559), .Y(n883) );
  INVX0_HVT U902 ( .A(n1561), .Y(n884) );
  INVX0_HVT U903 ( .A(n1563), .Y(n885) );
  INVX0_HVT U904 ( .A(n1565), .Y(n886) );
  INVX0_HVT U905 ( .A(n1567), .Y(n887) );
  INVX0_HVT U906 ( .A(n1569), .Y(n888) );
  INVX0_HVT U907 ( .A(n1571), .Y(n889) );
  INVX0_HVT U908 ( .A(n1573), .Y(n890) );
  INVX0_HVT U909 ( .A(n1575), .Y(n891) );
  INVX0_HVT U910 ( .A(n1577), .Y(n892) );
  INVX0_HVT U911 ( .A(n1580), .Y(n893) );
  INVX0_HVT U912 ( .A(a_din[3]), .Y(n894) );
  INVX0_HVT U913 ( .A(n1357), .Y(n895) );
  INVX0_HVT U914 ( .A(n1358), .Y(n896) );
  INVX0_HVT U915 ( .A(n1359), .Y(n897) );
  INVX0_HVT U916 ( .A(n1360), .Y(n898) );
  INVX0_HVT U917 ( .A(n1361), .Y(n899) );
  INVX0_HVT U918 ( .A(n1362), .Y(n900) );
  INVX0_HVT U919 ( .A(n1363), .Y(n901) );
  INVX0_HVT U920 ( .A(n1364), .Y(n902) );
  INVX0_HVT U921 ( .A(n1365), .Y(n903) );
  INVX0_HVT U922 ( .A(n1366), .Y(n904) );
  INVX0_HVT U923 ( .A(n1367), .Y(n905) );
  INVX0_HVT U924 ( .A(n1368), .Y(n906) );
  INVX0_HVT U925 ( .A(n1369), .Y(n907) );
  INVX0_HVT U926 ( .A(n1370), .Y(n908) );
  INVX0_HVT U927 ( .A(n1371), .Y(n909) );
  INVX0_HVT U928 ( .A(n1373), .Y(n910) );
  INVX0_HVT U929 ( .A(n1374), .Y(n911) );
  INVX0_HVT U930 ( .A(n1375), .Y(n912) );
  INVX0_HVT U931 ( .A(n1376), .Y(n913) );
  INVX0_HVT U932 ( .A(n1377), .Y(n914) );
  INVX0_HVT U933 ( .A(n1378), .Y(n915) );
  INVX0_HVT U934 ( .A(n1379), .Y(n916) );
  INVX0_HVT U935 ( .A(n1380), .Y(n917) );
  INVX0_HVT U936 ( .A(n1381), .Y(n918) );
  INVX0_HVT U937 ( .A(n1382), .Y(n919) );
  INVX0_HVT U938 ( .A(n1383), .Y(n920) );
  INVX0_HVT U939 ( .A(n1384), .Y(n921) );
  INVX0_HVT U940 ( .A(n1385), .Y(n922) );
  INVX0_HVT U941 ( .A(n1386), .Y(n923) );
  INVX0_HVT U942 ( .A(n1387), .Y(n924) );
  INVX0_HVT U943 ( .A(n1388), .Y(n925) );
  INVX0_HVT U944 ( .A(n1390), .Y(n926) );
  INVX0_HVT U945 ( .A(n1391), .Y(n927) );
  INVX0_HVT U946 ( .A(n1392), .Y(n928) );
  INVX0_HVT U947 ( .A(n1393), .Y(n929) );
  INVX0_HVT U948 ( .A(n1394), .Y(n930) );
  INVX0_HVT U949 ( .A(n1395), .Y(n931) );
  INVX0_HVT U950 ( .A(n1396), .Y(n932) );
  INVX0_HVT U951 ( .A(n1397), .Y(n933) );
  INVX0_HVT U952 ( .A(n1398), .Y(n934) );
  INVX0_HVT U953 ( .A(n1399), .Y(n935) );
  INVX0_HVT U954 ( .A(n1400), .Y(n936) );
  INVX0_HVT U955 ( .A(n1401), .Y(n937) );
  INVX0_HVT U956 ( .A(n1402), .Y(n938) );
  INVX0_HVT U957 ( .A(n1403), .Y(n939) );
  INVX0_HVT U958 ( .A(n1404), .Y(n940) );
  INVX0_HVT U959 ( .A(n1405), .Y(n941) );
  INVX0_HVT U960 ( .A(n1407), .Y(n942) );
  INVX0_HVT U961 ( .A(n1409), .Y(n943) );
  INVX0_HVT U962 ( .A(n1410), .Y(n944) );
  INVX0_HVT U963 ( .A(n1411), .Y(n945) );
  INVX0_HVT U964 ( .A(n1412), .Y(n946) );
  INVX0_HVT U965 ( .A(n1413), .Y(n947) );
  INVX0_HVT U966 ( .A(n1414), .Y(n948) );
  INVX0_HVT U967 ( .A(n1415), .Y(n949) );
  INVX0_HVT U968 ( .A(n1416), .Y(n950) );
  INVX0_HVT U969 ( .A(n1417), .Y(n951) );
  INVX0_HVT U970 ( .A(n1418), .Y(n952) );
  INVX0_HVT U971 ( .A(n1419), .Y(n953) );
  INVX0_HVT U972 ( .A(n1420), .Y(n954) );
  INVX0_HVT U973 ( .A(n1421), .Y(n955) );
  INVX0_HVT U974 ( .A(n1422), .Y(n956) );
  INVX0_HVT U975 ( .A(n1423), .Y(n957) );
  INVX0_HVT U976 ( .A(n1425), .Y(n958) );
  INVX0_HVT U977 ( .A(n1280), .Y(n959) );
  INVX0_HVT U978 ( .A(n1281), .Y(n960) );
  INVX0_HVT U979 ( .A(n1282), .Y(n961) );
  INVX0_HVT U980 ( .A(n1284), .Y(n962) );
  INVX0_HVT U981 ( .A(n1285), .Y(n963) );
  INVX0_HVT U982 ( .A(n1286), .Y(n964) );
  INVX0_HVT U983 ( .A(n1287), .Y(n965) );
  INVX0_HVT U984 ( .A(n1289), .Y(n966) );
  INVX0_HVT U985 ( .A(n1290), .Y(n967) );
  INVX0_HVT U986 ( .A(n1291), .Y(n968) );
  INVX0_HVT U987 ( .A(n1292), .Y(n969) );
  INVX0_HVT U988 ( .A(n1294), .Y(n970) );
  INVX0_HVT U989 ( .A(n1296), .Y(n971) );
  INVX0_HVT U990 ( .A(n1298), .Y(n972) );
  INVX0_HVT U991 ( .A(n1300), .Y(n973) );
  INVX0_HVT U992 ( .A(n1304), .Y(n974) );
  INVX0_HVT U993 ( .A(n1305), .Y(n975) );
  INVX0_HVT U994 ( .A(n1306), .Y(n976) );
  INVX0_HVT U995 ( .A(n1307), .Y(n977) );
  INVX0_HVT U996 ( .A(n1308), .Y(n978) );
  INVX0_HVT U997 ( .A(n1309), .Y(n979) );
  INVX0_HVT U998 ( .A(n1310), .Y(n980) );
  INVX0_HVT U999 ( .A(n1311), .Y(n981) );
  INVX0_HVT U1000 ( .A(n1312), .Y(n982) );
  INVX0_HVT U1001 ( .A(n1313), .Y(n983) );
  INVX0_HVT U1002 ( .A(n1314), .Y(n984) );
  INVX0_HVT U1003 ( .A(n1315), .Y(n985) );
  INVX0_HVT U1004 ( .A(n1316), .Y(n986) );
  INVX0_HVT U1005 ( .A(n1317), .Y(n987) );
  INVX0_HVT U1006 ( .A(n1318), .Y(n988) );
  INVX0_HVT U1007 ( .A(n1319), .Y(n989) );
  INVX0_HVT U1008 ( .A(n1321), .Y(n990) );
  INVX0_HVT U1009 ( .A(n1322), .Y(n991) );
  INVX0_HVT U1010 ( .A(n1323), .Y(n992) );
  INVX0_HVT U1011 ( .A(n1324), .Y(n993) );
  INVX0_HVT U1012 ( .A(n1325), .Y(n994) );
  INVX0_HVT U1013 ( .A(n1326), .Y(n995) );
  INVX0_HVT U1014 ( .A(n1327), .Y(n996) );
  INVX0_HVT U1015 ( .A(n1328), .Y(n997) );
  INVX0_HVT U1016 ( .A(n1329), .Y(n998) );
  INVX0_HVT U1017 ( .A(n1330), .Y(n999) );
  INVX0_HVT U1018 ( .A(n1331), .Y(n1000) );
  INVX0_HVT U1019 ( .A(n1332), .Y(n1001) );
  INVX0_HVT U1020 ( .A(n1333), .Y(n1002) );
  INVX0_HVT U1021 ( .A(n1334), .Y(n1003) );
  INVX0_HVT U1022 ( .A(n1335), .Y(n1004) );
  INVX0_HVT U1023 ( .A(n1336), .Y(n1005) );
  INVX0_HVT U1024 ( .A(n1338), .Y(n1006) );
  INVX0_HVT U1025 ( .A(n1340), .Y(n1007) );
  INVX0_HVT U1026 ( .A(n1341), .Y(n1008) );
  INVX0_HVT U1027 ( .A(n1342), .Y(n1009) );
  INVX0_HVT U1028 ( .A(n1343), .Y(n1010) );
  INVX0_HVT U1029 ( .A(n1344), .Y(n1011) );
  INVX0_HVT U1030 ( .A(n1345), .Y(n1012) );
  INVX0_HVT U1031 ( .A(n1346), .Y(n1013) );
  INVX0_HVT U1032 ( .A(n1347), .Y(n1014) );
  INVX0_HVT U1033 ( .A(n1348), .Y(n1015) );
  INVX0_HVT U1034 ( .A(n1349), .Y(n1016) );
  INVX0_HVT U1035 ( .A(n1350), .Y(n1017) );
  INVX0_HVT U1036 ( .A(n1351), .Y(n1018) );
  INVX0_HVT U1037 ( .A(n1352), .Y(n1019) );
  INVX0_HVT U1038 ( .A(n1353), .Y(n1020) );
  INVX0_HVT U1039 ( .A(n1354), .Y(n1021) );
  INVX0_HVT U1040 ( .A(n1356), .Y(n1022) );
  INVX0_HVT U1041 ( .A(a_din[2]), .Y(n1023) );
endmodule

