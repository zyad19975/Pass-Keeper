
module Get_key ( clk, rest, local_key, rount_no, key_round, done );
  input [127:0] local_key;
  input [3:0] rount_no;
  output [127:0] key_round;
  input clk, rest;
  output done;
  wire   n1994, n1996, n1998, n2000, n2002, n2004, n2006, n2008, n2010, n2012,
         n2014, n2016, n2018, n2020, n2022, n2024, n2026, n2028, n2030, n2032,
         n2034, n2036, n2038, n2040, n2042, n2044, n2046, n2048, n2050, n2052,
         n2054, n2056, n2058, n2060, n2062, n2064, n2066, n2068, n2070, n2072,
         n2074, n2076, n2078, n2080, n2082, n2084, n2086, n2088, n2090, n2092,
         n2094, n2096, n2098, n2100, n2102, n2104, n2106, n2108, n2110, n2112,
         n2114, n2116, n2118, n2120, n2122, n2124, n2126, n2128, n2130, n2132,
         n2134, n2136, n2138, n2140, n2142, n2144, n2146, n2148, n2150, n2152,
         n2154, n2156, n2158, n2160, n2162, n2164, n2166, n2168, n2170, n2172,
         n2174, n2176, n2178, n2180, n2182, n2184, n2186, n2188, n2190, n2192,
         n2194, n2196, n2198, n2200, n2202, n2204, n2206, n2208, n2210, n2212,
         n2214, n2216, n2218, n2220, n2222, n2224, n2226, n2228, n2230, n2232,
         n2234, n2236, n2238, n2240, n2242, n2244, n2246, n2248, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1995, n1997, n1999, n2001, n2003, n2005, n2007, n2009,
         n2011, n2013, n2015, n2017, n2019, n2021, n2023, n2025, n2027, n2029,
         n2031, n2033, n2035, n2037, n2039, n2041, n2043, n2045, n2047, n2049,
         n2051, n2053, n2055, n2057, n2059, n2061, n2063, n2065, n2067, n2069,
         n2071, n2073, n2075, n2077, n2079, n2081, n2083, n2085, n2087, n2089,
         n2091, n2093, n2095, n2097, n2099, n2101, n2103, n2105, n2107, n2109,
         n2111, n2113, n2115, n2117, n2119, n2121, n2123, n2125, n2127, n2129,
         n2131, n2133, n2135, n2137, n2139, n2141, n2143, n2145, n2147, n2149,
         n2151, n2153, n2155, n2157, n2159, n2161, n2163, n2165, n2167, n2169,
         n2171, n2173, n2175, n2177, n2179, n2181, n2183, n2185, n2187, n2189,
         n2191, n2193, n2195, n2197, n2199, n2201, n2203, n2205, n2207, n2209,
         n2211, n2213, n2215, n2217, n2219, n2221, n2223, n2225, n2227, n2229,
         n2231, n2233, n2235, n2237, n2239, n2241, n2243, n2245, n2247, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528;
  wire   [3:0] round_number;
  wire   [127:0] prev_key;
  wire   [127:0] keyout;
  wire   [3:0] state;

  DFFARX1_HVT \state_reg[0]  ( .D(n5205), .CLK(clk), .RSTB(n3528), .Q(state[0]), .QN(n385) );
  DFFARX1_HVT \state_reg[2]  ( .D(n5202), .CLK(clk), .RSTB(n3528), .Q(state[2]), .QN(n899) );
  DFFX1_HVT \keys_reg[0][99]  ( .D(n5068), .CLK(clk), .Q(n3527), .QN(n642) );
  DFFX1_HVT \keys_reg[0][100]  ( .D(n5067), .CLK(clk), .Q(n3526), .QN(n645) );
  DFFX1_HVT \keys_reg[0][101]  ( .D(n5066), .CLK(clk), .Q(n3525), .QN(n647) );
  DFFX1_HVT \keys_reg[0][102]  ( .D(n5065), .CLK(clk), .Q(n3524), .QN(n649) );
  DFFX1_HVT \keys_reg[0][103]  ( .D(n5064), .CLK(clk), .Q(n3523), .QN(n651) );
  DFFX1_HVT \keys_reg[0][104]  ( .D(n5063), .CLK(clk), .Q(n3522), .QN(n653) );
  DFFX1_HVT \keys_reg[0][105]  ( .D(n5062), .CLK(clk), .Q(n3521), .QN(n655) );
  DFFX1_HVT \keys_reg[0][106]  ( .D(n5061), .CLK(clk), .Q(n3520), .QN(n657) );
  DFFX1_HVT \keys_reg[0][107]  ( .D(n5060), .CLK(clk), .Q(n3519), .QN(n659) );
  DFFX1_HVT \keys_reg[0][108]  ( .D(n5059), .CLK(clk), .Q(n3518), .QN(n661) );
  DFFX1_HVT \keys_reg[0][109]  ( .D(n5058), .CLK(clk), .Q(n3517), .QN(n663) );
  DFFX1_HVT \keys_reg[0][110]  ( .D(n5057), .CLK(clk), .Q(n3516), .QN(n665) );
  DFFX1_HVT \keys_reg[0][111]  ( .D(n5056), .CLK(clk), .Q(n3515), .QN(n667) );
  DFFX1_HVT \keys_reg[0][112]  ( .D(n5055), .CLK(clk), .Q(n3514), .QN(n669) );
  DFFX1_HVT \keys_reg[0][113]  ( .D(n5054), .CLK(clk), .Q(n3513), .QN(n671) );
  DFFX1_HVT \keys_reg[0][114]  ( .D(n5053), .CLK(clk), .Q(n3512), .QN(n673) );
  DFFX1_HVT \keys_reg[0][115]  ( .D(n5052), .CLK(clk), .Q(n3511), .QN(n675) );
  DFFX1_HVT \keys_reg[0][116]  ( .D(n5051), .CLK(clk), .Q(n3510), .QN(n677) );
  DFFX1_HVT \keys_reg[0][117]  ( .D(n5050), .CLK(clk), .Q(n3509), .QN(n679) );
  DFFX1_HVT \keys_reg[0][118]  ( .D(n5049), .CLK(clk), .Q(n3508), .QN(n681) );
  DFFX1_HVT \keys_reg[0][119]  ( .D(n5048), .CLK(clk), .Q(n3507), .QN(n683) );
  DFFX1_HVT \keys_reg[0][120]  ( .D(n5047), .CLK(clk), .Q(n3506), .QN(n685) );
  DFFX1_HVT \keys_reg[0][121]  ( .D(n5046), .CLK(clk), .Q(n3505), .QN(n687) );
  DFFX1_HVT \keys_reg[0][122]  ( .D(n5045), .CLK(clk), .Q(n3504), .QN(n689) );
  DFFX1_HVT \keys_reg[0][123]  ( .D(n5044), .CLK(clk), .Q(n3503), .QN(n691) );
  DFFX1_HVT \keys_reg[0][124]  ( .D(n5043), .CLK(clk), .Q(n3502), .QN(n693) );
  DFFX1_HVT \keys_reg[0][125]  ( .D(n5042), .CLK(clk), .Q(n3501), .QN(n695) );
  DFFX1_HVT \keys_reg[0][126]  ( .D(n5041), .CLK(clk), .Q(n3500), .QN(n697) );
  DFFX1_HVT \keys_reg[0][127]  ( .D(n5040), .CLK(clk), .Q(n3499), .QN(n699) );
  DFFX1_HVT \keys_reg[0][77]  ( .D(n5039), .CLK(clk), .Q(n3498), .QN(n839) );
  DFFX1_HVT \keys_reg[0][78]  ( .D(n5038), .CLK(clk), .Q(n3497), .QN(n837) );
  DFFX1_HVT \keys_reg[0][79]  ( .D(n5037), .CLK(clk), .Q(n3496), .QN(n835) );
  DFFX1_HVT \keys_reg[0][80]  ( .D(n5036), .CLK(clk), .Q(n3495), .QN(n833) );
  DFFX1_HVT \keys_reg[0][81]  ( .D(n5035), .CLK(clk), .Q(n3494), .QN(n831) );
  DFFX1_HVT \keys_reg[0][82]  ( .D(n5034), .CLK(clk), .Q(n3493), .QN(n701) );
  DFFX1_HVT \keys_reg[0][83]  ( .D(n5033), .CLK(clk), .Q(n3492), .QN(n703) );
  DFFX1_HVT \keys_reg[0][84]  ( .D(n5032), .CLK(clk), .Q(n3491), .QN(n705) );
  DFFX1_HVT \keys_reg[0][85]  ( .D(n5031), .CLK(clk), .Q(n3490), .QN(n707) );
  DFFX1_HVT \keys_reg[0][86]  ( .D(n5030), .CLK(clk), .Q(n3489), .QN(n709) );
  DFFX1_HVT \keys_reg[0][87]  ( .D(n5029), .CLK(clk), .Q(n3488), .QN(n711) );
  DFFX1_HVT \keys_reg[0][88]  ( .D(n5028), .CLK(clk), .Q(n3487), .QN(n713) );
  DFFX1_HVT \keys_reg[0][89]  ( .D(n5027), .CLK(clk), .Q(n3486), .QN(n715) );
  DFFX1_HVT \keys_reg[0][90]  ( .D(n5026), .CLK(clk), .Q(n3485), .QN(n717) );
  DFFX1_HVT \keys_reg[0][91]  ( .D(n5025), .CLK(clk), .Q(n3484), .QN(n719) );
  DFFX1_HVT \keys_reg[0][92]  ( .D(n5024), .CLK(clk), .Q(n3483), .QN(n721) );
  DFFX1_HVT \keys_reg[0][93]  ( .D(n5023), .CLK(clk), .Q(n3482), .QN(n723) );
  DFFX1_HVT \keys_reg[0][94]  ( .D(n5022), .CLK(clk), .Q(n3481), .QN(n725) );
  DFFX1_HVT \keys_reg[0][95]  ( .D(n5021), .CLK(clk), .Q(n3480), .QN(n727) );
  DFFX1_HVT \keys_reg[0][96]  ( .D(n5020), .CLK(clk), .Q(n3479), .QN(n729) );
  DFFX1_HVT \keys_reg[0][97]  ( .D(n5019), .CLK(clk), .Q(n3478), .QN(n731) );
  DFFX1_HVT \keys_reg[0][0]  ( .D(n5018), .CLK(clk), .Q(n3477), .QN(n733) );
  DFFX1_HVT \keys_reg[0][1]  ( .D(n5017), .CLK(clk), .Q(n3476), .QN(n735) );
  DFFX1_HVT \keys_reg[0][2]  ( .D(n5016), .CLK(clk), .Q(n3475), .QN(n737) );
  DFFX1_HVT \keys_reg[0][3]  ( .D(n5015), .CLK(clk), .Q(n3474), .QN(n739) );
  DFFX1_HVT \keys_reg[0][4]  ( .D(n5014), .CLK(clk), .Q(n3473), .QN(n741) );
  DFFX1_HVT \keys_reg[0][5]  ( .D(n5013), .CLK(clk), .Q(n3472), .QN(n743) );
  DFFX1_HVT \keys_reg[0][6]  ( .D(n5012), .CLK(clk), .Q(n3471), .QN(n745) );
  DFFX1_HVT \keys_reg[0][7]  ( .D(n5011), .CLK(clk), .Q(n3470), .QN(n747) );
  DFFX1_HVT \keys_reg[0][8]  ( .D(n5010), .CLK(clk), .Q(n3469), .QN(n749) );
  DFFX1_HVT \keys_reg[0][9]  ( .D(n5009), .CLK(clk), .Q(n3468), .QN(n751) );
  DFFX1_HVT \keys_reg[0][10]  ( .D(n5008), .CLK(clk), .Q(n3467), .QN(n753) );
  DFFX1_HVT \keys_reg[0][11]  ( .D(n5007), .CLK(clk), .Q(n3466), .QN(n755) );
  DFFX1_HVT \keys_reg[0][12]  ( .D(n5006), .CLK(clk), .Q(n3465), .QN(n757) );
  DFFX1_HVT \keys_reg[0][13]  ( .D(n5005), .CLK(clk), .Q(n3464), .QN(n759) );
  DFFX1_HVT \keys_reg[0][14]  ( .D(n5004), .CLK(clk), .Q(n3463), .QN(n761) );
  DFFX1_HVT \keys_reg[0][15]  ( .D(n5003), .CLK(clk), .Q(n3462), .QN(n763) );
  DFFX1_HVT \keys_reg[0][16]  ( .D(n5002), .CLK(clk), .Q(n3461), .QN(n765) );
  DFFX1_HVT \keys_reg[0][17]  ( .D(n5001), .CLK(clk), .Q(n3460), .QN(n767) );
  DFFX1_HVT \keys_reg[0][18]  ( .D(n5000), .CLK(clk), .Q(n3459), .QN(n769) );
  DFFX1_HVT \keys_reg[0][19]  ( .D(n4999), .CLK(clk), .Q(n3458), .QN(n771) );
  DFFX1_HVT \keys_reg[0][20]  ( .D(n4998), .CLK(clk), .Q(n3457), .QN(n773) );
  DFFX1_HVT \keys_reg[0][21]  ( .D(n4997), .CLK(clk), .Q(n3456), .QN(n775) );
  DFFX1_HVT \keys_reg[0][22]  ( .D(n4996), .CLK(clk), .Q(n3455), .QN(n777) );
  DFFX1_HVT \keys_reg[0][23]  ( .D(n4995), .CLK(clk), .Q(n3454), .QN(n779) );
  DFFX1_HVT \keys_reg[0][24]  ( .D(n4994), .CLK(clk), .Q(n3453), .QN(n781) );
  DFFX1_HVT \keys_reg[0][25]  ( .D(n4993), .CLK(clk), .Q(n3452), .QN(n783) );
  DFFX1_HVT \keys_reg[0][26]  ( .D(n4992), .CLK(clk), .Q(n3451), .QN(n785) );
  DFFX1_HVT \keys_reg[0][27]  ( .D(n4991), .CLK(clk), .Q(n3450), .QN(n787) );
  DFFX1_HVT \keys_reg[0][28]  ( .D(n4990), .CLK(clk), .Q(n3449), .QN(n789) );
  DFFX1_HVT \keys_reg[0][29]  ( .D(n4989), .CLK(clk), .Q(n3448), .QN(n791) );
  DFFX1_HVT \keys_reg[0][30]  ( .D(n4988), .CLK(clk), .Q(n3447), .QN(n793) );
  DFFX1_HVT \keys_reg[0][31]  ( .D(n4987), .CLK(clk), .Q(n3446), .QN(n795) );
  DFFX1_HVT \keys_reg[0][32]  ( .D(n4986), .CLK(clk), .Q(n3445), .QN(n797) );
  DFFX1_HVT \keys_reg[0][33]  ( .D(n4985), .CLK(clk), .Q(n3444), .QN(n799) );
  DFFX1_HVT \keys_reg[0][34]  ( .D(n4984), .CLK(clk), .Q(n3443), .QN(n801) );
  DFFX1_HVT \keys_reg[0][35]  ( .D(n4983), .CLK(clk), .Q(n3442), .QN(n803) );
  DFFX1_HVT \keys_reg[0][36]  ( .D(n4982), .CLK(clk), .Q(n3441), .QN(n805) );
  DFFX1_HVT \keys_reg[0][37]  ( .D(n4981), .CLK(clk), .Q(n3440), .QN(n807) );
  DFFX1_HVT \keys_reg[0][38]  ( .D(n4980), .CLK(clk), .Q(n3439), .QN(n809) );
  DFFX1_HVT \keys_reg[0][39]  ( .D(n4979), .CLK(clk), .Q(n3438), .QN(n811) );
  DFFX1_HVT \keys_reg[0][40]  ( .D(n4978), .CLK(clk), .Q(n3437), .QN(n813) );
  DFFX1_HVT \keys_reg[0][41]  ( .D(n4977), .CLK(clk), .Q(n3436), .QN(n815) );
  DFFX1_HVT \keys_reg[0][42]  ( .D(n4976), .CLK(clk), .Q(n3435), .QN(n817) );
  DFFX1_HVT \keys_reg[0][43]  ( .D(n4975), .CLK(clk), .Q(n3434), .QN(n819) );
  DFFX1_HVT \keys_reg[0][44]  ( .D(n4974), .CLK(clk), .Q(n3433), .QN(n821) );
  DFFX1_HVT \keys_reg[0][45]  ( .D(n4973), .CLK(clk), .Q(n3432), .QN(n823) );
  DFFX1_HVT \keys_reg[0][46]  ( .D(n4972), .CLK(clk), .Q(n3431), .QN(n825) );
  DFFX1_HVT \keys_reg[0][47]  ( .D(n4971), .CLK(clk), .Q(n3430), .QN(n827) );
  DFFX1_HVT \keys_reg[0][48]  ( .D(n4970), .CLK(clk), .Q(n3429), .QN(n829) );
  DFFX1_HVT \keys_reg[0][76]  ( .D(n4969), .CLK(clk), .Q(n3428), .QN(n841) );
  DFFX1_HVT \keys_reg[0][75]  ( .D(n4968), .CLK(clk), .Q(n3427), .QN(n843) );
  DFFX1_HVT \keys_reg[0][74]  ( .D(n4967), .CLK(clk), .Q(n3426), .QN(n845) );
  DFFX1_HVT \keys_reg[0][73]  ( .D(n4966), .CLK(clk), .Q(n3425), .QN(n847) );
  DFFX1_HVT \keys_reg[0][72]  ( .D(n4965), .CLK(clk), .Q(n3424), .QN(n849) );
  DFFX1_HVT \keys_reg[0][71]  ( .D(n4964), .CLK(clk), .Q(n3423), .QN(n851) );
  DFFX1_HVT \keys_reg[0][70]  ( .D(n4963), .CLK(clk), .Q(n3422), .QN(n853) );
  DFFX1_HVT \keys_reg[0][69]  ( .D(n4962), .CLK(clk), .Q(n3421), .QN(n855) );
  DFFX1_HVT \keys_reg[0][68]  ( .D(n4961), .CLK(clk), .Q(n3420), .QN(n857) );
  DFFX1_HVT \keys_reg[0][67]  ( .D(n4960), .CLK(clk), .Q(n3419), .QN(n859) );
  DFFX1_HVT \keys_reg[0][66]  ( .D(n4959), .CLK(clk), .Q(n3418), .QN(n861) );
  DFFX1_HVT \keys_reg[0][65]  ( .D(n4958), .CLK(clk), .Q(n3417), .QN(n863) );
  DFFX1_HVT \keys_reg[0][64]  ( .D(n4957), .CLK(clk), .Q(n3416), .QN(n865) );
  DFFX1_HVT \keys_reg[0][63]  ( .D(n4956), .CLK(clk), .Q(n3415), .QN(n867) );
  DFFX1_HVT \keys_reg[0][62]  ( .D(n4955), .CLK(clk), .Q(n3414), .QN(n869) );
  DFFX1_HVT \keys_reg[0][61]  ( .D(n4954), .CLK(clk), .Q(n3413), .QN(n871) );
  DFFX1_HVT \keys_reg[0][60]  ( .D(n4953), .CLK(clk), .Q(n3412), .QN(n873) );
  DFFX1_HVT \keys_reg[0][59]  ( .D(n4952), .CLK(clk), .Q(n3411), .QN(n875) );
  DFFX1_HVT \keys_reg[0][58]  ( .D(n4951), .CLK(clk), .Q(n3410), .QN(n877) );
  DFFX1_HVT \keys_reg[0][57]  ( .D(n4950), .CLK(clk), .Q(n3409), .QN(n879) );
  DFFX1_HVT \keys_reg[0][56]  ( .D(n4949), .CLK(clk), .Q(n3408), .QN(n881) );
  DFFX1_HVT \keys_reg[0][55]  ( .D(n4948), .CLK(clk), .Q(n3407), .QN(n883) );
  DFFX1_HVT \keys_reg[0][54]  ( .D(n4947), .CLK(clk), .Q(n3406), .QN(n885) );
  DFFX1_HVT \keys_reg[0][53]  ( .D(n4946), .CLK(clk), .Q(n3405), .QN(n887) );
  DFFX1_HVT \keys_reg[0][52]  ( .D(n4945), .CLK(clk), .Q(n3404), .QN(n889) );
  DFFX1_HVT \keys_reg[0][51]  ( .D(n4944), .CLK(clk), .Q(n3403), .QN(n891) );
  DFFX1_HVT \keys_reg[0][50]  ( .D(n4943), .CLK(clk), .Q(n3402), .QN(n893) );
  DFFX1_HVT \keys_reg[0][49]  ( .D(n4942), .CLK(clk), .Q(n3401), .QN(n895) );
  DFFX1_HVT \keys_reg[0][98]  ( .D(n4941), .CLK(clk), .Q(n3400), .QN(n897) );
  DFFARX1_HVT \state_reg[1]  ( .D(n5203), .CLK(clk), .RSTB(n3528), .Q(n898), 
        .QN(n3399) );
  DFFARX1_HVT \state_reg[3]  ( .D(n5204), .CLK(clk), .RSTB(n3528), .QN(n3398)
         );
  DFFARX1_HVT done_reg ( .D(n4940), .CLK(clk), .RSTB(n3528), .Q(done), .QN(
        n1988) );
  DFFX1_HVT \round_number_reg[3]  ( .D(n5198), .CLK(clk), .Q(round_number[3])
         );
  DFFX1_HVT \round_number_reg[2]  ( .D(n5199), .CLK(clk), .Q(round_number[2])
         );
  DFFX1_HVT \round_number_reg[1]  ( .D(n5200), .CLK(clk), .Q(round_number[1])
         );
  DFFX1_HVT \round_number_reg[0]  ( .D(n5201), .CLK(clk), .Q(round_number[0]), 
        .QN(n1989) );
  DFFX1_HVT \keys_reg[10][0]  ( .D(n4939), .CLK(clk), .Q(n3397), .QN(n945) );
  DFFX1_HVT \keys_reg[9][0]  ( .D(n4938), .CLK(clk), .Q(n3396), .QN(n476) );
  DFFX1_HVT \keys_reg[8][0]  ( .D(n4937), .CLK(clk), .Q(n3395), .QN(n1165) );
  DFFX1_HVT \keys_reg[6][0]  ( .D(n4936), .CLK(clk), .Q(n3394), .QN(n475) );
  DFFX1_HVT \keys_reg[5][0]  ( .D(n4935), .CLK(clk), .Q(n3393), .QN(n1164) );
  DFFX1_HVT \keys_reg[4][0]  ( .D(n4934), .CLK(clk), .Q(n3392), .QN(n219) );
  DFFX1_HVT \keys_reg[3][0]  ( .D(n4933), .CLK(clk), .Q(n3391), .QN(n1163) );
  DFFX1_HVT \keys_reg[1][0]  ( .D(n4932), .CLK(clk), .Q(n3390), .QN(n220) );
  DFFX1_HVT \prev_key_reg[0]  ( .D(n5197), .CLK(clk), .Q(prev_key[0]) );
  DFFX1_HVT \keys_reg[10][1]  ( .D(n4931), .CLK(clk), .Q(n3389), .QN(n946) );
  DFFX1_HVT \keys_reg[9][1]  ( .D(n4930), .CLK(clk), .Q(n3388), .QN(n478) );
  DFFX1_HVT \keys_reg[8][1]  ( .D(n4929), .CLK(clk), .Q(n3387), .QN(n1168) );
  DFFX1_HVT \keys_reg[6][1]  ( .D(n4928), .CLK(clk), .Q(n3386), .QN(n477) );
  DFFX1_HVT \keys_reg[5][1]  ( .D(n4927), .CLK(clk), .Q(n3385), .QN(n1167) );
  DFFX1_HVT \keys_reg[4][1]  ( .D(n4926), .CLK(clk), .Q(n3384), .QN(n221) );
  DFFX1_HVT \keys_reg[3][1]  ( .D(n4925), .CLK(clk), .Q(n3383), .QN(n1166) );
  DFFX1_HVT \keys_reg[1][1]  ( .D(n4924), .CLK(clk), .Q(n3382), .QN(n222) );
  DFFX1_HVT \prev_key_reg[1]  ( .D(n5196), .CLK(clk), .Q(prev_key[1]) );
  DFFX1_HVT \keys_reg[10][2]  ( .D(n4923), .CLK(clk), .Q(n3381), .QN(n947) );
  DFFX1_HVT \keys_reg[9][2]  ( .D(n4922), .CLK(clk), .Q(n3380), .QN(n480) );
  DFFX1_HVT \keys_reg[8][2]  ( .D(n4921), .CLK(clk), .Q(n3379), .QN(n1171) );
  DFFX1_HVT \keys_reg[6][2]  ( .D(n4920), .CLK(clk), .Q(n3378), .QN(n479) );
  DFFX1_HVT \keys_reg[5][2]  ( .D(n4919), .CLK(clk), .Q(n3377), .QN(n1170) );
  DFFX1_HVT \keys_reg[4][2]  ( .D(n4918), .CLK(clk), .Q(n3376), .QN(n223) );
  DFFX1_HVT \keys_reg[3][2]  ( .D(n4917), .CLK(clk), .Q(n3375), .QN(n1169) );
  DFFX1_HVT \keys_reg[1][2]  ( .D(n4916), .CLK(clk), .Q(n3374), .QN(n224) );
  DFFX1_HVT \prev_key_reg[2]  ( .D(n5195), .CLK(clk), .Q(prev_key[2]) );
  DFFX1_HVT \keys_reg[10][3]  ( .D(n4915), .CLK(clk), .Q(n3373), .QN(n948) );
  DFFX1_HVT \keys_reg[9][3]  ( .D(n4914), .CLK(clk), .Q(n3372), .QN(n482) );
  DFFX1_HVT \keys_reg[8][3]  ( .D(n4913), .CLK(clk), .Q(n3371), .QN(n1174) );
  DFFX1_HVT \keys_reg[6][3]  ( .D(n4912), .CLK(clk), .Q(n3370), .QN(n481) );
  DFFX1_HVT \keys_reg[5][3]  ( .D(n4911), .CLK(clk), .Q(n3369), .QN(n1173) );
  DFFX1_HVT \keys_reg[4][3]  ( .D(n4910), .CLK(clk), .Q(n3368), .QN(n225) );
  DFFX1_HVT \keys_reg[3][3]  ( .D(n4909), .CLK(clk), .Q(n3367), .QN(n1172) );
  DFFX1_HVT \keys_reg[1][3]  ( .D(n4908), .CLK(clk), .Q(n3366), .QN(n226) );
  DFFX1_HVT \prev_key_reg[3]  ( .D(n5194), .CLK(clk), .Q(prev_key[3]) );
  DFFX1_HVT \keys_reg[10][4]  ( .D(n4907), .CLK(clk), .Q(n3365), .QN(n949) );
  DFFX1_HVT \keys_reg[9][4]  ( .D(n4906), .CLK(clk), .Q(n3364), .QN(n484) );
  DFFX1_HVT \keys_reg[8][4]  ( .D(n4905), .CLK(clk), .Q(n3363), .QN(n1177) );
  DFFX1_HVT \keys_reg[6][4]  ( .D(n4904), .CLK(clk), .Q(n3362), .QN(n483) );
  DFFX1_HVT \keys_reg[5][4]  ( .D(n4903), .CLK(clk), .Q(n3361), .QN(n1176) );
  DFFX1_HVT \keys_reg[4][4]  ( .D(n4902), .CLK(clk), .Q(n3360), .QN(n227) );
  DFFX1_HVT \keys_reg[3][4]  ( .D(n4901), .CLK(clk), .Q(n3359), .QN(n1175) );
  DFFX1_HVT \keys_reg[1][4]  ( .D(n4900), .CLK(clk), .Q(n3358), .QN(n228) );
  DFFX1_HVT \prev_key_reg[4]  ( .D(n5193), .CLK(clk), .Q(prev_key[4]) );
  DFFX1_HVT \keys_reg[10][5]  ( .D(n4899), .CLK(clk), .Q(n3357), .QN(n950) );
  DFFX1_HVT \keys_reg[9][5]  ( .D(n4898), .CLK(clk), .Q(n3356), .QN(n486) );
  DFFX1_HVT \keys_reg[8][5]  ( .D(n4897), .CLK(clk), .Q(n3355), .QN(n1180) );
  DFFX1_HVT \keys_reg[6][5]  ( .D(n4896), .CLK(clk), .Q(n3354), .QN(n485) );
  DFFX1_HVT \keys_reg[5][5]  ( .D(n4895), .CLK(clk), .Q(n3353), .QN(n1179) );
  DFFX1_HVT \keys_reg[4][5]  ( .D(n4894), .CLK(clk), .Q(n3352), .QN(n229) );
  DFFX1_HVT \keys_reg[3][5]  ( .D(n4893), .CLK(clk), .Q(n3351), .QN(n1178) );
  DFFX1_HVT \keys_reg[1][5]  ( .D(n4892), .CLK(clk), .Q(n3350), .QN(n230) );
  DFFX1_HVT \prev_key_reg[5]  ( .D(n5192), .CLK(clk), .Q(prev_key[5]) );
  DFFX1_HVT \keys_reg[10][6]  ( .D(n4891), .CLK(clk), .Q(n3349), .QN(n951) );
  DFFX1_HVT \keys_reg[9][6]  ( .D(n4890), .CLK(clk), .Q(n3348), .QN(n488) );
  DFFX1_HVT \keys_reg[8][6]  ( .D(n4889), .CLK(clk), .Q(n3347), .QN(n1183) );
  DFFX1_HVT \keys_reg[6][6]  ( .D(n4888), .CLK(clk), .Q(n3346), .QN(n487) );
  DFFX1_HVT \keys_reg[5][6]  ( .D(n4887), .CLK(clk), .Q(n3345), .QN(n1182) );
  DFFX1_HVT \keys_reg[4][6]  ( .D(n4886), .CLK(clk), .Q(n3344), .QN(n231) );
  DFFX1_HVT \keys_reg[3][6]  ( .D(n4885), .CLK(clk), .Q(n3343), .QN(n1181) );
  DFFX1_HVT \keys_reg[1][6]  ( .D(n4884), .CLK(clk), .Q(n3342), .QN(n232) );
  DFFX1_HVT \prev_key_reg[6]  ( .D(n5191), .CLK(clk), .Q(prev_key[6]) );
  DFFX1_HVT \keys_reg[10][7]  ( .D(n4883), .CLK(clk), .Q(n3341), .QN(n952) );
  DFFX1_HVT \keys_reg[9][7]  ( .D(n4882), .CLK(clk), .Q(n3340), .QN(n490) );
  DFFX1_HVT \keys_reg[8][7]  ( .D(n4881), .CLK(clk), .Q(n3339), .QN(n1186) );
  DFFX1_HVT \keys_reg[6][7]  ( .D(n4880), .CLK(clk), .Q(n3338), .QN(n489) );
  DFFX1_HVT \keys_reg[5][7]  ( .D(n4879), .CLK(clk), .Q(n3337), .QN(n1185) );
  DFFX1_HVT \keys_reg[4][7]  ( .D(n4878), .CLK(clk), .Q(n3336), .QN(n233) );
  DFFX1_HVT \keys_reg[3][7]  ( .D(n4877), .CLK(clk), .Q(n3335), .QN(n1184) );
  DFFX1_HVT \keys_reg[1][7]  ( .D(n4876), .CLK(clk), .Q(n3334), .QN(n234) );
  DFFX1_HVT \prev_key_reg[7]  ( .D(n5190), .CLK(clk), .Q(prev_key[7]) );
  DFFX1_HVT \keys_reg[10][8]  ( .D(n4875), .CLK(clk), .Q(n3333), .QN(n953) );
  DFFX1_HVT \keys_reg[9][8]  ( .D(n4874), .CLK(clk), .Q(n3332), .QN(n492) );
  DFFX1_HVT \keys_reg[8][8]  ( .D(n4873), .CLK(clk), .Q(n3331), .QN(n1189) );
  DFFX1_HVT \keys_reg[6][8]  ( .D(n4872), .CLK(clk), .Q(n3330), .QN(n491) );
  DFFX1_HVT \keys_reg[5][8]  ( .D(n4871), .CLK(clk), .Q(n3329), .QN(n1188) );
  DFFX1_HVT \keys_reg[4][8]  ( .D(n4870), .CLK(clk), .Q(n3328), .QN(n235) );
  DFFX1_HVT \keys_reg[3][8]  ( .D(n4869), .CLK(clk), .Q(n3327), .QN(n1187) );
  DFFX1_HVT \keys_reg[1][8]  ( .D(n4868), .CLK(clk), .Q(n3326), .QN(n236) );
  DFFX1_HVT \prev_key_reg[8]  ( .D(n5189), .CLK(clk), .Q(prev_key[8]) );
  DFFX1_HVT \keys_reg[10][9]  ( .D(n4867), .CLK(clk), .Q(n3325), .QN(n954) );
  DFFX1_HVT \keys_reg[9][9]  ( .D(n4866), .CLK(clk), .Q(n3324), .QN(n494) );
  DFFX1_HVT \keys_reg[8][9]  ( .D(n4865), .CLK(clk), .Q(n3323), .QN(n1192) );
  DFFX1_HVT \keys_reg[6][9]  ( .D(n4864), .CLK(clk), .Q(n3322), .QN(n493) );
  DFFX1_HVT \keys_reg[5][9]  ( .D(n4863), .CLK(clk), .Q(n3321), .QN(n1191) );
  DFFX1_HVT \keys_reg[4][9]  ( .D(n4862), .CLK(clk), .Q(n3320), .QN(n237) );
  DFFX1_HVT \keys_reg[3][9]  ( .D(n4861), .CLK(clk), .Q(n3319), .QN(n1190) );
  DFFX1_HVT \keys_reg[1][9]  ( .D(n4860), .CLK(clk), .Q(n3318), .QN(n238) );
  DFFX1_HVT \prev_key_reg[9]  ( .D(n5188), .CLK(clk), .Q(prev_key[9]) );
  DFFX1_HVT \keys_reg[10][10]  ( .D(n4859), .CLK(clk), .Q(n3317), .QN(n955) );
  DFFX1_HVT \keys_reg[9][10]  ( .D(n4858), .CLK(clk), .Q(n3316), .QN(n496) );
  DFFX1_HVT \keys_reg[8][10]  ( .D(n4857), .CLK(clk), .Q(n3315), .QN(n1195) );
  DFFX1_HVT \keys_reg[6][10]  ( .D(n4856), .CLK(clk), .Q(n3314), .QN(n495) );
  DFFX1_HVT \keys_reg[5][10]  ( .D(n4855), .CLK(clk), .Q(n3313), .QN(n1194) );
  DFFX1_HVT \keys_reg[4][10]  ( .D(n4854), .CLK(clk), .Q(n3312), .QN(n239) );
  DFFX1_HVT \keys_reg[3][10]  ( .D(n4853), .CLK(clk), .Q(n3311), .QN(n1193) );
  DFFX1_HVT \keys_reg[1][10]  ( .D(n4852), .CLK(clk), .Q(n3310), .QN(n240) );
  DFFX1_HVT \prev_key_reg[10]  ( .D(n5187), .CLK(clk), .Q(prev_key[10]) );
  DFFX1_HVT \keys_reg[10][11]  ( .D(n4851), .CLK(clk), .Q(n3309), .QN(n956) );
  DFFX1_HVT \keys_reg[9][11]  ( .D(n4850), .CLK(clk), .Q(n3308), .QN(n498) );
  DFFX1_HVT \keys_reg[8][11]  ( .D(n4849), .CLK(clk), .Q(n3307), .QN(n1198) );
  DFFX1_HVT \keys_reg[6][11]  ( .D(n4848), .CLK(clk), .Q(n3306), .QN(n497) );
  DFFX1_HVT \keys_reg[5][11]  ( .D(n4847), .CLK(clk), .Q(n3305), .QN(n1197) );
  DFFX1_HVT \keys_reg[4][11]  ( .D(n4846), .CLK(clk), .Q(n3304), .QN(n241) );
  DFFX1_HVT \keys_reg[3][11]  ( .D(n4845), .CLK(clk), .Q(n3303), .QN(n1196) );
  DFFX1_HVT \keys_reg[1][11]  ( .D(n4844), .CLK(clk), .Q(n3302), .QN(n242) );
  DFFX1_HVT \prev_key_reg[11]  ( .D(n5186), .CLK(clk), .Q(prev_key[11]) );
  DFFX1_HVT \keys_reg[10][12]  ( .D(n4843), .CLK(clk), .Q(n3301), .QN(n957) );
  DFFX1_HVT \keys_reg[9][12]  ( .D(n4842), .CLK(clk), .Q(n3300), .QN(n500) );
  DFFX1_HVT \keys_reg[8][12]  ( .D(n4841), .CLK(clk), .Q(n3299), .QN(n1201) );
  DFFX1_HVT \keys_reg[6][12]  ( .D(n4840), .CLK(clk), .Q(n3298), .QN(n499) );
  DFFX1_HVT \keys_reg[5][12]  ( .D(n4839), .CLK(clk), .Q(n3297), .QN(n1200) );
  DFFX1_HVT \keys_reg[4][12]  ( .D(n4838), .CLK(clk), .Q(n3296), .QN(n243) );
  DFFX1_HVT \keys_reg[3][12]  ( .D(n4837), .CLK(clk), .Q(n3295), .QN(n1199) );
  DFFX1_HVT \keys_reg[1][12]  ( .D(n4836), .CLK(clk), .Q(n3294), .QN(n244) );
  DFFX1_HVT \prev_key_reg[12]  ( .D(n5185), .CLK(clk), .Q(prev_key[12]) );
  DFFX1_HVT \keys_reg[10][13]  ( .D(n4835), .CLK(clk), .Q(n3293), .QN(n958) );
  DFFX1_HVT \keys_reg[9][13]  ( .D(n4834), .CLK(clk), .Q(n3292), .QN(n502) );
  DFFX1_HVT \keys_reg[8][13]  ( .D(n4833), .CLK(clk), .Q(n3291), .QN(n1204) );
  DFFX1_HVT \keys_reg[6][13]  ( .D(n4832), .CLK(clk), .Q(n3290), .QN(n501) );
  DFFX1_HVT \keys_reg[5][13]  ( .D(n4831), .CLK(clk), .Q(n3289), .QN(n1203) );
  DFFX1_HVT \keys_reg[4][13]  ( .D(n4830), .CLK(clk), .Q(n3288), .QN(n245) );
  DFFX1_HVT \keys_reg[3][13]  ( .D(n4829), .CLK(clk), .Q(n3287), .QN(n1202) );
  DFFX1_HVT \keys_reg[1][13]  ( .D(n4828), .CLK(clk), .Q(n3286), .QN(n246) );
  DFFX1_HVT \prev_key_reg[13]  ( .D(n5184), .CLK(clk), .Q(prev_key[13]) );
  DFFX1_HVT \keys_reg[10][14]  ( .D(n4827), .CLK(clk), .Q(n3285), .QN(n959) );
  DFFX1_HVT \keys_reg[9][14]  ( .D(n4826), .CLK(clk), .Q(n3284), .QN(n504) );
  DFFX1_HVT \keys_reg[8][14]  ( .D(n4825), .CLK(clk), .Q(n3283), .QN(n1207) );
  DFFX1_HVT \keys_reg[6][14]  ( .D(n4824), .CLK(clk), .Q(n3282), .QN(n503) );
  DFFX1_HVT \keys_reg[5][14]  ( .D(n4823), .CLK(clk), .Q(n3281), .QN(n1206) );
  DFFX1_HVT \keys_reg[4][14]  ( .D(n4822), .CLK(clk), .Q(n3280), .QN(n247) );
  DFFX1_HVT \keys_reg[3][14]  ( .D(n4821), .CLK(clk), .Q(n3279), .QN(n1205) );
  DFFX1_HVT \keys_reg[1][14]  ( .D(n4820), .CLK(clk), .Q(n3278), .QN(n248) );
  DFFX1_HVT \prev_key_reg[14]  ( .D(n5183), .CLK(clk), .Q(prev_key[14]) );
  DFFX1_HVT \keys_reg[10][15]  ( .D(n4819), .CLK(clk), .Q(n3277), .QN(n960) );
  DFFX1_HVT \keys_reg[9][15]  ( .D(n4818), .CLK(clk), .Q(n3276), .QN(n506) );
  DFFX1_HVT \keys_reg[8][15]  ( .D(n4817), .CLK(clk), .Q(n3275), .QN(n1210) );
  DFFX1_HVT \keys_reg[6][15]  ( .D(n4816), .CLK(clk), .Q(n3274), .QN(n505) );
  DFFX1_HVT \keys_reg[5][15]  ( .D(n4815), .CLK(clk), .Q(n3273), .QN(n1209) );
  DFFX1_HVT \keys_reg[4][15]  ( .D(n4814), .CLK(clk), .Q(n3272), .QN(n249) );
  DFFX1_HVT \keys_reg[3][15]  ( .D(n4813), .CLK(clk), .Q(n3271), .QN(n1208) );
  DFFX1_HVT \keys_reg[1][15]  ( .D(n4812), .CLK(clk), .Q(n3270), .QN(n250) );
  DFFX1_HVT \prev_key_reg[15]  ( .D(n5182), .CLK(clk), .Q(prev_key[15]) );
  DFFX1_HVT \keys_reg[10][16]  ( .D(n4811), .CLK(clk), .Q(n3269), .QN(n961) );
  DFFX1_HVT \keys_reg[9][16]  ( .D(n4810), .CLK(clk), .Q(n3268), .QN(n508) );
  DFFX1_HVT \keys_reg[8][16]  ( .D(n4809), .CLK(clk), .Q(n3267), .QN(n1213) );
  DFFX1_HVT \keys_reg[6][16]  ( .D(n4808), .CLK(clk), .Q(n3266), .QN(n507) );
  DFFX1_HVT \keys_reg[5][16]  ( .D(n4807), .CLK(clk), .Q(n3265), .QN(n1212) );
  DFFX1_HVT \keys_reg[4][16]  ( .D(n4806), .CLK(clk), .Q(n3264), .QN(n251) );
  DFFX1_HVT \keys_reg[3][16]  ( .D(n4805), .CLK(clk), .Q(n3263), .QN(n1211) );
  DFFX1_HVT \keys_reg[1][16]  ( .D(n4804), .CLK(clk), .Q(n3262), .QN(n252) );
  DFFX1_HVT \prev_key_reg[16]  ( .D(n5181), .CLK(clk), .Q(prev_key[16]) );
  DFFX1_HVT \keys_reg[10][17]  ( .D(n4803), .CLK(clk), .Q(n3261), .QN(n962) );
  DFFX1_HVT \keys_reg[9][17]  ( .D(n4802), .CLK(clk), .Q(n3260), .QN(n510) );
  DFFX1_HVT \keys_reg[8][17]  ( .D(n4801), .CLK(clk), .Q(n3259), .QN(n1216) );
  DFFX1_HVT \keys_reg[6][17]  ( .D(n4800), .CLK(clk), .Q(n3258), .QN(n509) );
  DFFX1_HVT \keys_reg[5][17]  ( .D(n4799), .CLK(clk), .Q(n3257), .QN(n1215) );
  DFFX1_HVT \keys_reg[4][17]  ( .D(n4798), .CLK(clk), .Q(n3256), .QN(n253) );
  DFFX1_HVT \keys_reg[3][17]  ( .D(n4797), .CLK(clk), .Q(n3255), .QN(n1214) );
  DFFX1_HVT \keys_reg[1][17]  ( .D(n4796), .CLK(clk), .Q(n3254), .QN(n254) );
  DFFX1_HVT \prev_key_reg[17]  ( .D(n5180), .CLK(clk), .Q(prev_key[17]) );
  DFFX1_HVT \keys_reg[10][18]  ( .D(n4795), .CLK(clk), .Q(n3253), .QN(n963) );
  DFFX1_HVT \keys_reg[9][18]  ( .D(n4794), .CLK(clk), .Q(n3252), .QN(n512) );
  DFFX1_HVT \keys_reg[8][18]  ( .D(n4793), .CLK(clk), .Q(n3251), .QN(n1219) );
  DFFX1_HVT \keys_reg[6][18]  ( .D(n4792), .CLK(clk), .Q(n3250), .QN(n511) );
  DFFX1_HVT \keys_reg[5][18]  ( .D(n4791), .CLK(clk), .Q(n3249), .QN(n1218) );
  DFFX1_HVT \keys_reg[4][18]  ( .D(n4790), .CLK(clk), .Q(n3248), .QN(n255) );
  DFFX1_HVT \keys_reg[3][18]  ( .D(n4789), .CLK(clk), .Q(n3247), .QN(n1217) );
  DFFX1_HVT \keys_reg[1][18]  ( .D(n4788), .CLK(clk), .Q(n3246), .QN(n256) );
  DFFX1_HVT \prev_key_reg[18]  ( .D(n5179), .CLK(clk), .Q(prev_key[18]) );
  DFFX1_HVT \keys_reg[10][19]  ( .D(n4787), .CLK(clk), .Q(n3245), .QN(n964) );
  DFFX1_HVT \keys_reg[9][19]  ( .D(n4786), .CLK(clk), .Q(n3244), .QN(n514) );
  DFFX1_HVT \keys_reg[8][19]  ( .D(n4785), .CLK(clk), .Q(n3243), .QN(n1222) );
  DFFX1_HVT \keys_reg[6][19]  ( .D(n4784), .CLK(clk), .Q(n3242), .QN(n513) );
  DFFX1_HVT \keys_reg[5][19]  ( .D(n4783), .CLK(clk), .Q(n3241), .QN(n1221) );
  DFFX1_HVT \keys_reg[4][19]  ( .D(n4782), .CLK(clk), .Q(n3240), .QN(n257) );
  DFFX1_HVT \keys_reg[3][19]  ( .D(n4781), .CLK(clk), .Q(n3239), .QN(n1220) );
  DFFX1_HVT \keys_reg[1][19]  ( .D(n4780), .CLK(clk), .Q(n3238), .QN(n258) );
  DFFX1_HVT \prev_key_reg[19]  ( .D(n5178), .CLK(clk), .Q(prev_key[19]) );
  DFFX1_HVT \keys_reg[10][20]  ( .D(n4779), .CLK(clk), .Q(n3237), .QN(n965) );
  DFFX1_HVT \keys_reg[9][20]  ( .D(n4778), .CLK(clk), .Q(n3236), .QN(n516) );
  DFFX1_HVT \keys_reg[8][20]  ( .D(n4777), .CLK(clk), .Q(n3235), .QN(n1225) );
  DFFX1_HVT \keys_reg[6][20]  ( .D(n4776), .CLK(clk), .Q(n3234), .QN(n515) );
  DFFX1_HVT \keys_reg[5][20]  ( .D(n4775), .CLK(clk), .Q(n3233), .QN(n1224) );
  DFFX1_HVT \keys_reg[4][20]  ( .D(n4774), .CLK(clk), .Q(n3232), .QN(n259) );
  DFFX1_HVT \keys_reg[3][20]  ( .D(n4773), .CLK(clk), .Q(n3231), .QN(n1223) );
  DFFX1_HVT \keys_reg[1][20]  ( .D(n4772), .CLK(clk), .Q(n3230), .QN(n260) );
  DFFX1_HVT \prev_key_reg[20]  ( .D(n5177), .CLK(clk), .Q(prev_key[20]) );
  DFFX1_HVT \keys_reg[10][21]  ( .D(n4771), .CLK(clk), .Q(n3229), .QN(n966) );
  DFFX1_HVT \keys_reg[9][21]  ( .D(n4770), .CLK(clk), .Q(n3228), .QN(n518) );
  DFFX1_HVT \keys_reg[8][21]  ( .D(n4769), .CLK(clk), .Q(n3227), .QN(n1228) );
  DFFX1_HVT \keys_reg[6][21]  ( .D(n4768), .CLK(clk), .Q(n3226), .QN(n517) );
  DFFX1_HVT \keys_reg[5][21]  ( .D(n4767), .CLK(clk), .Q(n3225), .QN(n1227) );
  DFFX1_HVT \keys_reg[4][21]  ( .D(n4766), .CLK(clk), .Q(n3224), .QN(n261) );
  DFFX1_HVT \keys_reg[3][21]  ( .D(n4765), .CLK(clk), .Q(n3223), .QN(n1226) );
  DFFX1_HVT \keys_reg[1][21]  ( .D(n4764), .CLK(clk), .Q(n3222), .QN(n262) );
  DFFX1_HVT \prev_key_reg[21]  ( .D(n5176), .CLK(clk), .Q(prev_key[21]) );
  DFFX1_HVT \keys_reg[10][22]  ( .D(n4763), .CLK(clk), .Q(n3221), .QN(n967) );
  DFFX1_HVT \keys_reg[9][22]  ( .D(n4762), .CLK(clk), .Q(n3220), .QN(n520) );
  DFFX1_HVT \keys_reg[8][22]  ( .D(n4761), .CLK(clk), .Q(n3219), .QN(n1231) );
  DFFX1_HVT \keys_reg[6][22]  ( .D(n4760), .CLK(clk), .Q(n3218), .QN(n519) );
  DFFX1_HVT \keys_reg[5][22]  ( .D(n4759), .CLK(clk), .Q(n3217), .QN(n1230) );
  DFFX1_HVT \keys_reg[4][22]  ( .D(n4758), .CLK(clk), .Q(n3216), .QN(n263) );
  DFFX1_HVT \keys_reg[3][22]  ( .D(n4757), .CLK(clk), .Q(n3215), .QN(n1229) );
  DFFX1_HVT \keys_reg[1][22]  ( .D(n4756), .CLK(clk), .Q(n3214), .QN(n264) );
  DFFX1_HVT \prev_key_reg[22]  ( .D(n5175), .CLK(clk), .Q(prev_key[22]) );
  DFFX1_HVT \keys_reg[10][23]  ( .D(n4755), .CLK(clk), .Q(n3213), .QN(n968) );
  DFFX1_HVT \keys_reg[9][23]  ( .D(n4754), .CLK(clk), .Q(n3212), .QN(n522) );
  DFFX1_HVT \keys_reg[8][23]  ( .D(n4753), .CLK(clk), .Q(n3211), .QN(n1234) );
  DFFX1_HVT \keys_reg[6][23]  ( .D(n4752), .CLK(clk), .Q(n3210), .QN(n521) );
  DFFX1_HVT \keys_reg[5][23]  ( .D(n4751), .CLK(clk), .Q(n3209), .QN(n1233) );
  DFFX1_HVT \keys_reg[4][23]  ( .D(n4750), .CLK(clk), .Q(n3208), .QN(n265) );
  DFFX1_HVT \keys_reg[3][23]  ( .D(n4749), .CLK(clk), .Q(n3207), .QN(n1232) );
  DFFX1_HVT \keys_reg[1][23]  ( .D(n4748), .CLK(clk), .Q(n3206), .QN(n266) );
  DFFX1_HVT \prev_key_reg[23]  ( .D(n5174), .CLK(clk), .Q(prev_key[23]) );
  DFFX1_HVT \keys_reg[10][24]  ( .D(n4747), .CLK(clk), .Q(n3205), .QN(n969) );
  DFFX1_HVT \keys_reg[9][24]  ( .D(n4746), .CLK(clk), .Q(n3204), .QN(n524) );
  DFFX1_HVT \keys_reg[8][24]  ( .D(n4745), .CLK(clk), .Q(n3203), .QN(n1237) );
  DFFX1_HVT \keys_reg[6][24]  ( .D(n4744), .CLK(clk), .Q(n3202), .QN(n523) );
  DFFX1_HVT \keys_reg[5][24]  ( .D(n4743), .CLK(clk), .Q(n3201), .QN(n1236) );
  DFFX1_HVT \keys_reg[4][24]  ( .D(n4742), .CLK(clk), .Q(n3200), .QN(n267) );
  DFFX1_HVT \keys_reg[3][24]  ( .D(n4741), .CLK(clk), .Q(n3199), .QN(n1235) );
  DFFX1_HVT \keys_reg[1][24]  ( .D(n4740), .CLK(clk), .Q(n3198), .QN(n268) );
  DFFX1_HVT \prev_key_reg[24]  ( .D(n5173), .CLK(clk), .Q(prev_key[24]) );
  DFFX1_HVT \keys_reg[10][25]  ( .D(n4739), .CLK(clk), .Q(n3197), .QN(n970) );
  DFFX1_HVT \keys_reg[9][25]  ( .D(n4738), .CLK(clk), .Q(n3196), .QN(n526) );
  DFFX1_HVT \keys_reg[8][25]  ( .D(n4737), .CLK(clk), .Q(n3195), .QN(n1240) );
  DFFX1_HVT \keys_reg[6][25]  ( .D(n4736), .CLK(clk), .Q(n3194), .QN(n525) );
  DFFX1_HVT \keys_reg[5][25]  ( .D(n4735), .CLK(clk), .Q(n3193), .QN(n1239) );
  DFFX1_HVT \keys_reg[4][25]  ( .D(n4734), .CLK(clk), .Q(n3192), .QN(n269) );
  DFFX1_HVT \keys_reg[3][25]  ( .D(n4733), .CLK(clk), .Q(n3191), .QN(n1238) );
  DFFX1_HVT \keys_reg[1][25]  ( .D(n4732), .CLK(clk), .Q(n3190), .QN(n270) );
  DFFX1_HVT \prev_key_reg[25]  ( .D(n5172), .CLK(clk), .Q(prev_key[25]) );
  DFFX1_HVT \keys_reg[10][26]  ( .D(n4731), .CLK(clk), .Q(n3189), .QN(n971) );
  DFFX1_HVT \keys_reg[9][26]  ( .D(n4730), .CLK(clk), .Q(n3188), .QN(n528) );
  DFFX1_HVT \keys_reg[8][26]  ( .D(n4729), .CLK(clk), .Q(n3187), .QN(n1243) );
  DFFX1_HVT \keys_reg[6][26]  ( .D(n4728), .CLK(clk), .Q(n3186), .QN(n527) );
  DFFX1_HVT \keys_reg[5][26]  ( .D(n4727), .CLK(clk), .Q(n3185), .QN(n1242) );
  DFFX1_HVT \keys_reg[4][26]  ( .D(n4726), .CLK(clk), .Q(n3184), .QN(n271) );
  DFFX1_HVT \keys_reg[3][26]  ( .D(n4725), .CLK(clk), .Q(n3183), .QN(n1241) );
  DFFX1_HVT \keys_reg[1][26]  ( .D(n4724), .CLK(clk), .Q(n3182), .QN(n272) );
  DFFX1_HVT \prev_key_reg[26]  ( .D(n5171), .CLK(clk), .Q(prev_key[26]) );
  DFFX1_HVT \keys_reg[10][27]  ( .D(n4723), .CLK(clk), .Q(n3181), .QN(n972) );
  DFFX1_HVT \keys_reg[9][27]  ( .D(n4722), .CLK(clk), .Q(n3180), .QN(n530) );
  DFFX1_HVT \keys_reg[8][27]  ( .D(n4721), .CLK(clk), .Q(n3179), .QN(n1246) );
  DFFX1_HVT \keys_reg[6][27]  ( .D(n4720), .CLK(clk), .Q(n3178), .QN(n529) );
  DFFX1_HVT \keys_reg[5][27]  ( .D(n4719), .CLK(clk), .Q(n3177), .QN(n1245) );
  DFFX1_HVT \keys_reg[4][27]  ( .D(n4718), .CLK(clk), .Q(n3176), .QN(n273) );
  DFFX1_HVT \keys_reg[3][27]  ( .D(n4717), .CLK(clk), .Q(n3175), .QN(n1244) );
  DFFX1_HVT \keys_reg[1][27]  ( .D(n4716), .CLK(clk), .Q(n3174), .QN(n274) );
  DFFX1_HVT \prev_key_reg[27]  ( .D(n5170), .CLK(clk), .Q(prev_key[27]) );
  DFFX1_HVT \keys_reg[10][28]  ( .D(n4715), .CLK(clk), .Q(n3173), .QN(n973) );
  DFFX1_HVT \keys_reg[9][28]  ( .D(n4714), .CLK(clk), .Q(n3172), .QN(n532) );
  DFFX1_HVT \keys_reg[8][28]  ( .D(n4713), .CLK(clk), .Q(n3171), .QN(n1249) );
  DFFX1_HVT \keys_reg[6][28]  ( .D(n4712), .CLK(clk), .Q(n3170), .QN(n531) );
  DFFX1_HVT \keys_reg[5][28]  ( .D(n4711), .CLK(clk), .Q(n3169), .QN(n1248) );
  DFFX1_HVT \keys_reg[4][28]  ( .D(n4710), .CLK(clk), .Q(n3168), .QN(n275) );
  DFFX1_HVT \keys_reg[3][28]  ( .D(n4709), .CLK(clk), .Q(n3167), .QN(n1247) );
  DFFX1_HVT \keys_reg[1][28]  ( .D(n4708), .CLK(clk), .Q(n3166), .QN(n276) );
  DFFX1_HVT \prev_key_reg[28]  ( .D(n5169), .CLK(clk), .Q(prev_key[28]) );
  DFFX1_HVT \keys_reg[10][29]  ( .D(n4707), .CLK(clk), .Q(n3165), .QN(n974) );
  DFFX1_HVT \keys_reg[9][29]  ( .D(n4706), .CLK(clk), .Q(n3164), .QN(n534) );
  DFFX1_HVT \keys_reg[8][29]  ( .D(n4705), .CLK(clk), .Q(n3163), .QN(n1252) );
  DFFX1_HVT \keys_reg[6][29]  ( .D(n4704), .CLK(clk), .Q(n3162), .QN(n533) );
  DFFX1_HVT \keys_reg[5][29]  ( .D(n4703), .CLK(clk), .Q(n3161), .QN(n1251) );
  DFFX1_HVT \keys_reg[4][29]  ( .D(n4702), .CLK(clk), .Q(n3160), .QN(n277) );
  DFFX1_HVT \keys_reg[3][29]  ( .D(n4701), .CLK(clk), .Q(n3159), .QN(n1250) );
  DFFX1_HVT \keys_reg[1][29]  ( .D(n4700), .CLK(clk), .Q(n3158), .QN(n278) );
  DFFX1_HVT \prev_key_reg[29]  ( .D(n5168), .CLK(clk), .Q(prev_key[29]) );
  DFFX1_HVT \keys_reg[10][30]  ( .D(n4699), .CLK(clk), .Q(n3157), .QN(n975) );
  DFFX1_HVT \keys_reg[9][30]  ( .D(n4698), .CLK(clk), .Q(n3156), .QN(n536) );
  DFFX1_HVT \keys_reg[8][30]  ( .D(n4697), .CLK(clk), .Q(n3155), .QN(n1255) );
  DFFX1_HVT \keys_reg[6][30]  ( .D(n4696), .CLK(clk), .Q(n3154), .QN(n535) );
  DFFX1_HVT \keys_reg[5][30]  ( .D(n4695), .CLK(clk), .Q(n3153), .QN(n1254) );
  DFFX1_HVT \keys_reg[4][30]  ( .D(n4694), .CLK(clk), .Q(n3152), .QN(n279) );
  DFFX1_HVT \keys_reg[3][30]  ( .D(n4693), .CLK(clk), .Q(n3151), .QN(n1253) );
  DFFX1_HVT \keys_reg[1][30]  ( .D(n4692), .CLK(clk), .Q(n3150), .QN(n280) );
  DFFX1_HVT \prev_key_reg[30]  ( .D(n5167), .CLK(clk), .Q(prev_key[30]) );
  DFFX1_HVT \keys_reg[10][31]  ( .D(n4691), .CLK(clk), .Q(n3149), .QN(n976) );
  DFFX1_HVT \keys_reg[9][31]  ( .D(n4690), .CLK(clk), .Q(n3148), .QN(n538) );
  DFFX1_HVT \keys_reg[8][31]  ( .D(n4689), .CLK(clk), .Q(n3147), .QN(n1258) );
  DFFX1_HVT \keys_reg[6][31]  ( .D(n4688), .CLK(clk), .Q(n3146), .QN(n537) );
  DFFX1_HVT \keys_reg[5][31]  ( .D(n4687), .CLK(clk), .Q(n3145), .QN(n1257) );
  DFFX1_HVT \keys_reg[4][31]  ( .D(n4686), .CLK(clk), .Q(n3144), .QN(n281) );
  DFFX1_HVT \keys_reg[3][31]  ( .D(n4685), .CLK(clk), .Q(n3143), .QN(n1256) );
  DFFX1_HVT \keys_reg[1][31]  ( .D(n4684), .CLK(clk), .Q(n3142), .QN(n282) );
  DFFX1_HVT \prev_key_reg[31]  ( .D(n5166), .CLK(clk), .Q(prev_key[31]) );
  DFFX1_HVT \keys_reg[10][32]  ( .D(n4683), .CLK(clk), .Q(n3141), .QN(n977) );
  DFFX1_HVT \keys_reg[9][32]  ( .D(n4682), .CLK(clk), .Q(n3140), .QN(n540) );
  DFFX1_HVT \keys_reg[8][32]  ( .D(n4681), .CLK(clk), .Q(n3139), .QN(n1261) );
  DFFX1_HVT \keys_reg[6][32]  ( .D(n4680), .CLK(clk), .Q(n3138), .QN(n539) );
  DFFX1_HVT \keys_reg[5][32]  ( .D(n4679), .CLK(clk), .Q(n3137), .QN(n1260) );
  DFFX1_HVT \keys_reg[4][32]  ( .D(n4678), .CLK(clk), .Q(n3136), .QN(n283) );
  DFFX1_HVT \keys_reg[3][32]  ( .D(n4677), .CLK(clk), .Q(n3135), .QN(n1259) );
  DFFX1_HVT \keys_reg[1][32]  ( .D(n4676), .CLK(clk), .Q(n3134), .QN(n284) );
  DFFX1_HVT \prev_key_reg[32]  ( .D(n5165), .CLK(clk), .Q(prev_key[32]) );
  DFFX1_HVT \keys_reg[10][33]  ( .D(n4675), .CLK(clk), .Q(n3133), .QN(n978) );
  DFFX1_HVT \keys_reg[9][33]  ( .D(n4674), .CLK(clk), .Q(n3132), .QN(n542) );
  DFFX1_HVT \keys_reg[8][33]  ( .D(n4673), .CLK(clk), .Q(n3131), .QN(n1264) );
  DFFX1_HVT \keys_reg[6][33]  ( .D(n4672), .CLK(clk), .Q(n3130), .QN(n541) );
  DFFX1_HVT \keys_reg[5][33]  ( .D(n4671), .CLK(clk), .Q(n3129), .QN(n1263) );
  DFFX1_HVT \keys_reg[4][33]  ( .D(n4670), .CLK(clk), .Q(n3128), .QN(n285) );
  DFFX1_HVT \keys_reg[3][33]  ( .D(n4669), .CLK(clk), .Q(n3127), .QN(n1262) );
  DFFX1_HVT \keys_reg[1][33]  ( .D(n4668), .CLK(clk), .Q(n3126), .QN(n286) );
  DFFX1_HVT \prev_key_reg[33]  ( .D(n5164), .CLK(clk), .Q(prev_key[33]) );
  DFFX1_HVT \keys_reg[10][34]  ( .D(n4667), .CLK(clk), .Q(n3125), .QN(n979) );
  DFFX1_HVT \keys_reg[9][34]  ( .D(n4666), .CLK(clk), .Q(n3124), .QN(n544) );
  DFFX1_HVT \keys_reg[8][34]  ( .D(n4665), .CLK(clk), .Q(n3123), .QN(n1267) );
  DFFX1_HVT \keys_reg[6][34]  ( .D(n4664), .CLK(clk), .Q(n3122), .QN(n543) );
  DFFX1_HVT \keys_reg[5][34]  ( .D(n4663), .CLK(clk), .Q(n3121), .QN(n1266) );
  DFFX1_HVT \keys_reg[4][34]  ( .D(n4662), .CLK(clk), .Q(n3120), .QN(n287) );
  DFFX1_HVT \keys_reg[3][34]  ( .D(n4661), .CLK(clk), .Q(n3119), .QN(n1265) );
  DFFX1_HVT \keys_reg[1][34]  ( .D(n4660), .CLK(clk), .Q(n3118), .QN(n288) );
  DFFX1_HVT \prev_key_reg[34]  ( .D(n5163), .CLK(clk), .Q(prev_key[34]) );
  DFFX1_HVT \keys_reg[10][35]  ( .D(n4659), .CLK(clk), .Q(n3117), .QN(n980) );
  DFFX1_HVT \keys_reg[9][35]  ( .D(n4658), .CLK(clk), .Q(n3116), .QN(n546) );
  DFFX1_HVT \keys_reg[8][35]  ( .D(n4657), .CLK(clk), .Q(n3115), .QN(n1270) );
  DFFX1_HVT \keys_reg[6][35]  ( .D(n4656), .CLK(clk), .Q(n3114), .QN(n545) );
  DFFX1_HVT \keys_reg[5][35]  ( .D(n4655), .CLK(clk), .Q(n3113), .QN(n1269) );
  DFFX1_HVT \keys_reg[4][35]  ( .D(n4654), .CLK(clk), .Q(n3112), .QN(n289) );
  DFFX1_HVT \keys_reg[3][35]  ( .D(n4653), .CLK(clk), .Q(n3111), .QN(n1268) );
  DFFX1_HVT \keys_reg[1][35]  ( .D(n4652), .CLK(clk), .Q(n3110), .QN(n290) );
  DFFX1_HVT \prev_key_reg[35]  ( .D(n5162), .CLK(clk), .Q(prev_key[35]) );
  DFFX1_HVT \keys_reg[10][36]  ( .D(n4651), .CLK(clk), .Q(n3109), .QN(n981) );
  DFFX1_HVT \keys_reg[9][36]  ( .D(n4650), .CLK(clk), .Q(n3108), .QN(n548) );
  DFFX1_HVT \keys_reg[8][36]  ( .D(n4649), .CLK(clk), .Q(n3107), .QN(n1273) );
  DFFX1_HVT \keys_reg[6][36]  ( .D(n4648), .CLK(clk), .Q(n3106), .QN(n547) );
  DFFX1_HVT \keys_reg[5][36]  ( .D(n4647), .CLK(clk), .Q(n3105), .QN(n1272) );
  DFFX1_HVT \keys_reg[4][36]  ( .D(n4646), .CLK(clk), .Q(n3104), .QN(n291) );
  DFFX1_HVT \keys_reg[3][36]  ( .D(n4645), .CLK(clk), .Q(n3103), .QN(n1271) );
  DFFX1_HVT \keys_reg[1][36]  ( .D(n4644), .CLK(clk), .Q(n3102), .QN(n292) );
  DFFX1_HVT \prev_key_reg[36]  ( .D(n5161), .CLK(clk), .Q(prev_key[36]) );
  DFFX1_HVT \keys_reg[10][37]  ( .D(n4643), .CLK(clk), .Q(n3101), .QN(n982) );
  DFFX1_HVT \keys_reg[9][37]  ( .D(n4642), .CLK(clk), .Q(n3100), .QN(n550) );
  DFFX1_HVT \keys_reg[8][37]  ( .D(n4641), .CLK(clk), .Q(n3099), .QN(n1276) );
  DFFX1_HVT \keys_reg[6][37]  ( .D(n4640), .CLK(clk), .Q(n3098), .QN(n549) );
  DFFX1_HVT \keys_reg[5][37]  ( .D(n4639), .CLK(clk), .Q(n3097), .QN(n1275) );
  DFFX1_HVT \keys_reg[4][37]  ( .D(n4638), .CLK(clk), .Q(n3096), .QN(n293) );
  DFFX1_HVT \keys_reg[3][37]  ( .D(n4637), .CLK(clk), .Q(n3095), .QN(n1274) );
  DFFX1_HVT \keys_reg[1][37]  ( .D(n4636), .CLK(clk), .Q(n3094), .QN(n294) );
  DFFX1_HVT \prev_key_reg[37]  ( .D(n5160), .CLK(clk), .Q(prev_key[37]) );
  DFFX1_HVT \keys_reg[10][38]  ( .D(n4635), .CLK(clk), .Q(n3093), .QN(n983) );
  DFFX1_HVT \keys_reg[9][38]  ( .D(n4634), .CLK(clk), .Q(n3092), .QN(n552) );
  DFFX1_HVT \keys_reg[8][38]  ( .D(n4633), .CLK(clk), .Q(n3091), .QN(n1279) );
  DFFX1_HVT \keys_reg[6][38]  ( .D(n4632), .CLK(clk), .Q(n3090), .QN(n551) );
  DFFX1_HVT \keys_reg[5][38]  ( .D(n4631), .CLK(clk), .Q(n3089), .QN(n1278) );
  DFFX1_HVT \keys_reg[4][38]  ( .D(n4630), .CLK(clk), .Q(n3088), .QN(n295) );
  DFFX1_HVT \keys_reg[3][38]  ( .D(n4629), .CLK(clk), .Q(n3087), .QN(n1277) );
  DFFX1_HVT \keys_reg[1][38]  ( .D(n4628), .CLK(clk), .Q(n3086), .QN(n296) );
  DFFX1_HVT \prev_key_reg[38]  ( .D(n5159), .CLK(clk), .Q(prev_key[38]) );
  DFFX1_HVT \keys_reg[10][39]  ( .D(n4627), .CLK(clk), .Q(n3085), .QN(n984) );
  DFFX1_HVT \keys_reg[9][39]  ( .D(n4626), .CLK(clk), .Q(n3084), .QN(n554) );
  DFFX1_HVT \keys_reg[8][39]  ( .D(n4625), .CLK(clk), .Q(n3083), .QN(n1282) );
  DFFX1_HVT \keys_reg[6][39]  ( .D(n4624), .CLK(clk), .Q(n3082), .QN(n553) );
  DFFX1_HVT \keys_reg[5][39]  ( .D(n4623), .CLK(clk), .Q(n3081), .QN(n1281) );
  DFFX1_HVT \keys_reg[4][39]  ( .D(n4622), .CLK(clk), .Q(n3080), .QN(n297) );
  DFFX1_HVT \keys_reg[3][39]  ( .D(n4621), .CLK(clk), .Q(n3079), .QN(n1280) );
  DFFX1_HVT \keys_reg[1][39]  ( .D(n4620), .CLK(clk), .Q(n3078), .QN(n298) );
  DFFX1_HVT \prev_key_reg[39]  ( .D(n5158), .CLK(clk), .Q(prev_key[39]) );
  DFFX1_HVT \keys_reg[10][40]  ( .D(n4619), .CLK(clk), .Q(n3077), .QN(n985) );
  DFFX1_HVT \keys_reg[9][40]  ( .D(n4618), .CLK(clk), .Q(n3076), .QN(n556) );
  DFFX1_HVT \keys_reg[8][40]  ( .D(n4617), .CLK(clk), .Q(n3075), .QN(n1285) );
  DFFX1_HVT \keys_reg[6][40]  ( .D(n4616), .CLK(clk), .Q(n3074), .QN(n555) );
  DFFX1_HVT \keys_reg[5][40]  ( .D(n4615), .CLK(clk), .Q(n3073), .QN(n1284) );
  DFFX1_HVT \keys_reg[4][40]  ( .D(n4614), .CLK(clk), .Q(n3072), .QN(n299) );
  DFFX1_HVT \keys_reg[3][40]  ( .D(n4613), .CLK(clk), .Q(n3071), .QN(n1283) );
  DFFX1_HVT \keys_reg[1][40]  ( .D(n4612), .CLK(clk), .Q(n3070), .QN(n300) );
  DFFX1_HVT \prev_key_reg[40]  ( .D(n5157), .CLK(clk), .Q(prev_key[40]) );
  DFFX1_HVT \keys_reg[10][41]  ( .D(n4611), .CLK(clk), .Q(n3069), .QN(n986) );
  DFFX1_HVT \keys_reg[9][41]  ( .D(n4610), .CLK(clk), .Q(n3068), .QN(n558) );
  DFFX1_HVT \keys_reg[8][41]  ( .D(n4609), .CLK(clk), .Q(n3067), .QN(n1288) );
  DFFX1_HVT \keys_reg[6][41]  ( .D(n4608), .CLK(clk), .Q(n3066), .QN(n557) );
  DFFX1_HVT \keys_reg[5][41]  ( .D(n4607), .CLK(clk), .Q(n3065), .QN(n1287) );
  DFFX1_HVT \keys_reg[4][41]  ( .D(n4606), .CLK(clk), .Q(n3064), .QN(n301) );
  DFFX1_HVT \keys_reg[3][41]  ( .D(n4605), .CLK(clk), .Q(n3063), .QN(n1286) );
  DFFX1_HVT \keys_reg[1][41]  ( .D(n4604), .CLK(clk), .Q(n3062), .QN(n302) );
  DFFX1_HVT \prev_key_reg[41]  ( .D(n5156), .CLK(clk), .Q(prev_key[41]) );
  DFFX1_HVT \keys_reg[10][42]  ( .D(n4603), .CLK(clk), .Q(n3061), .QN(n987) );
  DFFX1_HVT \keys_reg[9][42]  ( .D(n4602), .CLK(clk), .Q(n3060), .QN(n560) );
  DFFX1_HVT \keys_reg[8][42]  ( .D(n4601), .CLK(clk), .Q(n3059), .QN(n1291) );
  DFFX1_HVT \keys_reg[6][42]  ( .D(n4600), .CLK(clk), .Q(n3058), .QN(n559) );
  DFFX1_HVT \keys_reg[5][42]  ( .D(n4599), .CLK(clk), .Q(n3057), .QN(n1290) );
  DFFX1_HVT \keys_reg[4][42]  ( .D(n4598), .CLK(clk), .Q(n3056), .QN(n303) );
  DFFX1_HVT \keys_reg[3][42]  ( .D(n4597), .CLK(clk), .Q(n3055), .QN(n1289) );
  DFFX1_HVT \keys_reg[1][42]  ( .D(n4596), .CLK(clk), .Q(n3054), .QN(n304) );
  DFFX1_HVT \prev_key_reg[42]  ( .D(n5155), .CLK(clk), .Q(prev_key[42]) );
  DFFX1_HVT \keys_reg[10][43]  ( .D(n4595), .CLK(clk), .Q(n3053), .QN(n988) );
  DFFX1_HVT \keys_reg[9][43]  ( .D(n4594), .CLK(clk), .Q(n3052), .QN(n562) );
  DFFX1_HVT \keys_reg[8][43]  ( .D(n4593), .CLK(clk), .Q(n3051), .QN(n1294) );
  DFFX1_HVT \keys_reg[6][43]  ( .D(n4592), .CLK(clk), .Q(n3050), .QN(n561) );
  DFFX1_HVT \keys_reg[5][43]  ( .D(n4591), .CLK(clk), .Q(n3049), .QN(n1293) );
  DFFX1_HVT \keys_reg[4][43]  ( .D(n4590), .CLK(clk), .Q(n3048), .QN(n305) );
  DFFX1_HVT \keys_reg[3][43]  ( .D(n4589), .CLK(clk), .Q(n3047), .QN(n1292) );
  DFFX1_HVT \keys_reg[1][43]  ( .D(n4588), .CLK(clk), .Q(n3046), .QN(n306) );
  DFFX1_HVT \prev_key_reg[43]  ( .D(n5154), .CLK(clk), .Q(prev_key[43]) );
  DFFX1_HVT \keys_reg[10][44]  ( .D(n4587), .CLK(clk), .Q(n3045), .QN(n989) );
  DFFX1_HVT \keys_reg[9][44]  ( .D(n4586), .CLK(clk), .Q(n3044), .QN(n564) );
  DFFX1_HVT \keys_reg[8][44]  ( .D(n4585), .CLK(clk), .Q(n3043), .QN(n1297) );
  DFFX1_HVT \keys_reg[6][44]  ( .D(n4584), .CLK(clk), .Q(n3042), .QN(n563) );
  DFFX1_HVT \keys_reg[5][44]  ( .D(n4583), .CLK(clk), .Q(n3041), .QN(n1296) );
  DFFX1_HVT \keys_reg[4][44]  ( .D(n4582), .CLK(clk), .Q(n3040), .QN(n307) );
  DFFX1_HVT \keys_reg[3][44]  ( .D(n4581), .CLK(clk), .Q(n3039), .QN(n1295) );
  DFFX1_HVT \keys_reg[1][44]  ( .D(n4580), .CLK(clk), .Q(n3038), .QN(n308) );
  DFFX1_HVT \prev_key_reg[44]  ( .D(n5153), .CLK(clk), .Q(prev_key[44]) );
  DFFX1_HVT \keys_reg[10][45]  ( .D(n4579), .CLK(clk), .Q(n3037), .QN(n990) );
  DFFX1_HVT \keys_reg[9][45]  ( .D(n4578), .CLK(clk), .Q(n3036), .QN(n566) );
  DFFX1_HVT \keys_reg[8][45]  ( .D(n4577), .CLK(clk), .Q(n3035), .QN(n1300) );
  DFFX1_HVT \keys_reg[6][45]  ( .D(n4576), .CLK(clk), .Q(n3034), .QN(n565) );
  DFFX1_HVT \keys_reg[5][45]  ( .D(n4575), .CLK(clk), .Q(n3033), .QN(n1299) );
  DFFX1_HVT \keys_reg[4][45]  ( .D(n4574), .CLK(clk), .Q(n3032), .QN(n309) );
  DFFX1_HVT \keys_reg[3][45]  ( .D(n4573), .CLK(clk), .Q(n3031), .QN(n1298) );
  DFFX1_HVT \keys_reg[1][45]  ( .D(n4572), .CLK(clk), .Q(n3030), .QN(n310) );
  DFFX1_HVT \prev_key_reg[45]  ( .D(n5152), .CLK(clk), .Q(prev_key[45]) );
  DFFX1_HVT \keys_reg[10][46]  ( .D(n4571), .CLK(clk), .Q(n3029), .QN(n991) );
  DFFX1_HVT \keys_reg[9][46]  ( .D(n4570), .CLK(clk), .Q(n3028), .QN(n568) );
  DFFX1_HVT \keys_reg[8][46]  ( .D(n4569), .CLK(clk), .Q(n3027), .QN(n1303) );
  DFFX1_HVT \keys_reg[6][46]  ( .D(n4568), .CLK(clk), .Q(n3026), .QN(n567) );
  DFFX1_HVT \keys_reg[5][46]  ( .D(n4567), .CLK(clk), .Q(n3025), .QN(n1302) );
  DFFX1_HVT \keys_reg[4][46]  ( .D(n4566), .CLK(clk), .Q(n3024), .QN(n311) );
  DFFX1_HVT \keys_reg[3][46]  ( .D(n4565), .CLK(clk), .Q(n3023), .QN(n1301) );
  DFFX1_HVT \keys_reg[1][46]  ( .D(n4564), .CLK(clk), .Q(n3022), .QN(n312) );
  DFFX1_HVT \prev_key_reg[46]  ( .D(n5151), .CLK(clk), .Q(prev_key[46]) );
  DFFX1_HVT \keys_reg[10][47]  ( .D(n4563), .CLK(clk), .Q(n3021), .QN(n992) );
  DFFX1_HVT \keys_reg[9][47]  ( .D(n4562), .CLK(clk), .Q(n3020), .QN(n570) );
  DFFX1_HVT \keys_reg[8][47]  ( .D(n4561), .CLK(clk), .Q(n3019), .QN(n1306) );
  DFFX1_HVT \keys_reg[6][47]  ( .D(n4560), .CLK(clk), .Q(n3018), .QN(n569) );
  DFFX1_HVT \keys_reg[5][47]  ( .D(n4559), .CLK(clk), .Q(n3017), .QN(n1305) );
  DFFX1_HVT \keys_reg[4][47]  ( .D(n4558), .CLK(clk), .Q(n3016), .QN(n313) );
  DFFX1_HVT \keys_reg[3][47]  ( .D(n4557), .CLK(clk), .Q(n3015), .QN(n1304) );
  DFFX1_HVT \keys_reg[1][47]  ( .D(n4556), .CLK(clk), .Q(n3014), .QN(n314) );
  DFFX1_HVT \prev_key_reg[47]  ( .D(n5150), .CLK(clk), .Q(prev_key[47]) );
  DFFX1_HVT \keys_reg[10][48]  ( .D(n4555), .CLK(clk), .Q(n3013), .QN(n993) );
  DFFX1_HVT \keys_reg[9][48]  ( .D(n4554), .CLK(clk), .Q(n3012), .QN(n572) );
  DFFX1_HVT \keys_reg[8][48]  ( .D(n4553), .CLK(clk), .Q(n3011), .QN(n1309) );
  DFFX1_HVT \keys_reg[6][48]  ( .D(n4552), .CLK(clk), .Q(n3010), .QN(n571) );
  DFFX1_HVT \keys_reg[5][48]  ( .D(n4551), .CLK(clk), .Q(n3009), .QN(n1308) );
  DFFX1_HVT \keys_reg[4][48]  ( .D(n4550), .CLK(clk), .Q(n3008), .QN(n315) );
  DFFX1_HVT \keys_reg[3][48]  ( .D(n4549), .CLK(clk), .Q(n3007), .QN(n1307) );
  DFFX1_HVT \keys_reg[1][48]  ( .D(n4548), .CLK(clk), .Q(n3006), .QN(n316) );
  DFFX1_HVT \prev_key_reg[48]  ( .D(n5149), .CLK(clk), .Q(prev_key[48]) );
  DFFX1_HVT \keys_reg[10][49]  ( .D(n4547), .CLK(clk), .Q(n3005), .QN(n1026)
         );
  DFFX1_HVT \keys_reg[9][49]  ( .D(n4546), .CLK(clk), .Q(n3004), .QN(n638) );
  DFFX1_HVT \keys_reg[8][49]  ( .D(n4545), .CLK(clk), .Q(n3003), .QN(n1408) );
  DFFX1_HVT \keys_reg[6][49]  ( .D(n4544), .CLK(clk), .Q(n3002), .QN(n637) );
  DFFX1_HVT \keys_reg[5][49]  ( .D(n4543), .CLK(clk), .Q(n3001), .QN(n1407) );
  DFFX1_HVT \keys_reg[4][49]  ( .D(n4542), .CLK(clk), .Q(n3000), .QN(n381) );
  DFFX1_HVT \keys_reg[3][49]  ( .D(n4541), .CLK(clk), .Q(n2999), .QN(n1406) );
  DFFX1_HVT \keys_reg[1][49]  ( .D(n4540), .CLK(clk), .Q(n2998), .QN(n382) );
  DFFX1_HVT \prev_key_reg[49]  ( .D(n5148), .CLK(clk), .Q(prev_key[49]) );
  DFFX1_HVT \keys_reg[10][50]  ( .D(n4539), .CLK(clk), .Q(n2997), .QN(n1025)
         );
  DFFX1_HVT \keys_reg[9][50]  ( .D(n4538), .CLK(clk), .Q(n2996), .QN(n636) );
  DFFX1_HVT \keys_reg[8][50]  ( .D(n4537), .CLK(clk), .Q(n2995), .QN(n1405) );
  DFFX1_HVT \keys_reg[6][50]  ( .D(n4536), .CLK(clk), .Q(n2994), .QN(n635) );
  DFFX1_HVT \keys_reg[5][50]  ( .D(n4535), .CLK(clk), .Q(n2993), .QN(n1404) );
  DFFX1_HVT \keys_reg[4][50]  ( .D(n4534), .CLK(clk), .Q(n2992), .QN(n379) );
  DFFX1_HVT \keys_reg[3][50]  ( .D(n4533), .CLK(clk), .Q(n2991), .QN(n1403) );
  DFFX1_HVT \keys_reg[1][50]  ( .D(n4532), .CLK(clk), .Q(n2990), .QN(n380) );
  DFFX1_HVT \prev_key_reg[50]  ( .D(n5147), .CLK(clk), .Q(prev_key[50]) );
  DFFX1_HVT \keys_reg[10][51]  ( .D(n4531), .CLK(clk), .Q(n2989), .QN(n1024)
         );
  DFFX1_HVT \keys_reg[9][51]  ( .D(n4530), .CLK(clk), .Q(n2988), .QN(n634) );
  DFFX1_HVT \keys_reg[8][51]  ( .D(n4529), .CLK(clk), .Q(n2987), .QN(n1402) );
  DFFX1_HVT \keys_reg[6][51]  ( .D(n4528), .CLK(clk), .Q(n2986), .QN(n633) );
  DFFX1_HVT \keys_reg[5][51]  ( .D(n4527), .CLK(clk), .Q(n2985), .QN(n1401) );
  DFFX1_HVT \keys_reg[4][51]  ( .D(n4526), .CLK(clk), .Q(n2984), .QN(n377) );
  DFFX1_HVT \keys_reg[3][51]  ( .D(n4525), .CLK(clk), .Q(n2983), .QN(n1400) );
  DFFX1_HVT \keys_reg[1][51]  ( .D(n4524), .CLK(clk), .Q(n2982), .QN(n378) );
  DFFX1_HVT \prev_key_reg[51]  ( .D(n5146), .CLK(clk), .Q(prev_key[51]) );
  DFFX1_HVT \keys_reg[10][52]  ( .D(n4523), .CLK(clk), .Q(n2981), .QN(n1023)
         );
  DFFX1_HVT \keys_reg[9][52]  ( .D(n4522), .CLK(clk), .Q(n2980), .QN(n632) );
  DFFX1_HVT \keys_reg[8][52]  ( .D(n4521), .CLK(clk), .Q(n2979), .QN(n1399) );
  DFFX1_HVT \keys_reg[6][52]  ( .D(n4520), .CLK(clk), .Q(n2978), .QN(n631) );
  DFFX1_HVT \keys_reg[5][52]  ( .D(n4519), .CLK(clk), .Q(n2977), .QN(n1398) );
  DFFX1_HVT \keys_reg[4][52]  ( .D(n4518), .CLK(clk), .Q(n2976), .QN(n375) );
  DFFX1_HVT \keys_reg[3][52]  ( .D(n4517), .CLK(clk), .Q(n2975), .QN(n1397) );
  DFFX1_HVT \keys_reg[1][52]  ( .D(n4516), .CLK(clk), .Q(n2974), .QN(n376) );
  DFFX1_HVT \prev_key_reg[52]  ( .D(n5145), .CLK(clk), .Q(prev_key[52]) );
  DFFX1_HVT \keys_reg[10][53]  ( .D(n4515), .CLK(clk), .Q(n2973), .QN(n1022)
         );
  DFFX1_HVT \keys_reg[9][53]  ( .D(n4514), .CLK(clk), .Q(n2972), .QN(n630) );
  DFFX1_HVT \keys_reg[8][53]  ( .D(n4513), .CLK(clk), .Q(n2971), .QN(n1396) );
  DFFX1_HVT \keys_reg[6][53]  ( .D(n4512), .CLK(clk), .Q(n2970), .QN(n629) );
  DFFX1_HVT \keys_reg[5][53]  ( .D(n4511), .CLK(clk), .Q(n2969), .QN(n1395) );
  DFFX1_HVT \keys_reg[4][53]  ( .D(n4510), .CLK(clk), .Q(n2968), .QN(n373) );
  DFFX1_HVT \keys_reg[3][53]  ( .D(n4509), .CLK(clk), .Q(n2967), .QN(n1394) );
  DFFX1_HVT \keys_reg[1][53]  ( .D(n4508), .CLK(clk), .Q(n2966), .QN(n374) );
  DFFX1_HVT \prev_key_reg[53]  ( .D(n5144), .CLK(clk), .Q(prev_key[53]) );
  DFFX1_HVT \keys_reg[10][54]  ( .D(n4507), .CLK(clk), .Q(n2965), .QN(n1021)
         );
  DFFX1_HVT \keys_reg[9][54]  ( .D(n4506), .CLK(clk), .Q(n2964), .QN(n628) );
  DFFX1_HVT \keys_reg[8][54]  ( .D(n4505), .CLK(clk), .Q(n2963), .QN(n1393) );
  DFFX1_HVT \keys_reg[6][54]  ( .D(n4504), .CLK(clk), .Q(n2962), .QN(n627) );
  DFFX1_HVT \keys_reg[5][54]  ( .D(n4503), .CLK(clk), .Q(n2961), .QN(n1392) );
  DFFX1_HVT \keys_reg[4][54]  ( .D(n4502), .CLK(clk), .Q(n2960), .QN(n371) );
  DFFX1_HVT \keys_reg[3][54]  ( .D(n4501), .CLK(clk), .Q(n2959), .QN(n1391) );
  DFFX1_HVT \keys_reg[1][54]  ( .D(n4500), .CLK(clk), .Q(n2958), .QN(n372) );
  DFFX1_HVT \prev_key_reg[54]  ( .D(n5143), .CLK(clk), .Q(prev_key[54]) );
  DFFX1_HVT \keys_reg[10][55]  ( .D(n4499), .CLK(clk), .Q(n2957), .QN(n1020)
         );
  DFFX1_HVT \keys_reg[9][55]  ( .D(n4498), .CLK(clk), .Q(n2956), .QN(n626) );
  DFFX1_HVT \keys_reg[8][55]  ( .D(n4497), .CLK(clk), .Q(n2955), .QN(n1390) );
  DFFX1_HVT \keys_reg[6][55]  ( .D(n4496), .CLK(clk), .Q(n2954), .QN(n625) );
  DFFX1_HVT \keys_reg[5][55]  ( .D(n4495), .CLK(clk), .Q(n2953), .QN(n1389) );
  DFFX1_HVT \keys_reg[4][55]  ( .D(n4494), .CLK(clk), .Q(n2952), .QN(n369) );
  DFFX1_HVT \keys_reg[3][55]  ( .D(n4493), .CLK(clk), .Q(n2951), .QN(n1388) );
  DFFX1_HVT \keys_reg[1][55]  ( .D(n4492), .CLK(clk), .Q(n2950), .QN(n370) );
  DFFX1_HVT \prev_key_reg[55]  ( .D(n5142), .CLK(clk), .Q(prev_key[55]) );
  DFFX1_HVT \keys_reg[10][56]  ( .D(n4491), .CLK(clk), .Q(n2949), .QN(n1019)
         );
  DFFX1_HVT \keys_reg[9][56]  ( .D(n4490), .CLK(clk), .Q(n2948), .QN(n624) );
  DFFX1_HVT \keys_reg[8][56]  ( .D(n4489), .CLK(clk), .Q(n2947), .QN(n1387) );
  DFFX1_HVT \keys_reg[6][56]  ( .D(n4488), .CLK(clk), .Q(n2946), .QN(n623) );
  DFFX1_HVT \keys_reg[5][56]  ( .D(n4487), .CLK(clk), .Q(n2945), .QN(n1386) );
  DFFX1_HVT \keys_reg[4][56]  ( .D(n4486), .CLK(clk), .Q(n2944), .QN(n367) );
  DFFX1_HVT \keys_reg[3][56]  ( .D(n4485), .CLK(clk), .Q(n2943), .QN(n1385) );
  DFFX1_HVT \keys_reg[1][56]  ( .D(n4484), .CLK(clk), .Q(n2942), .QN(n368) );
  DFFX1_HVT \prev_key_reg[56]  ( .D(n5141), .CLK(clk), .Q(prev_key[56]) );
  DFFX1_HVT \keys_reg[10][57]  ( .D(n4483), .CLK(clk), .Q(n2941), .QN(n1018)
         );
  DFFX1_HVT \keys_reg[9][57]  ( .D(n4482), .CLK(clk), .Q(n2940), .QN(n622) );
  DFFX1_HVT \keys_reg[8][57]  ( .D(n4481), .CLK(clk), .Q(n2939), .QN(n1384) );
  DFFX1_HVT \keys_reg[6][57]  ( .D(n4480), .CLK(clk), .Q(n2938), .QN(n621) );
  DFFX1_HVT \keys_reg[5][57]  ( .D(n4479), .CLK(clk), .Q(n2937), .QN(n1383) );
  DFFX1_HVT \keys_reg[4][57]  ( .D(n4478), .CLK(clk), .Q(n2936), .QN(n365) );
  DFFX1_HVT \keys_reg[3][57]  ( .D(n4477), .CLK(clk), .Q(n2935), .QN(n1382) );
  DFFX1_HVT \keys_reg[1][57]  ( .D(n4476), .CLK(clk), .Q(n2934), .QN(n366) );
  DFFX1_HVT \prev_key_reg[57]  ( .D(n5140), .CLK(clk), .Q(prev_key[57]) );
  DFFX1_HVT \keys_reg[10][58]  ( .D(n4475), .CLK(clk), .Q(n2933), .QN(n1017)
         );
  DFFX1_HVT \keys_reg[9][58]  ( .D(n4474), .CLK(clk), .Q(n2932), .QN(n620) );
  DFFX1_HVT \keys_reg[8][58]  ( .D(n4473), .CLK(clk), .Q(n2931), .QN(n1381) );
  DFFX1_HVT \keys_reg[6][58]  ( .D(n4472), .CLK(clk), .Q(n2930), .QN(n619) );
  DFFX1_HVT \keys_reg[5][58]  ( .D(n4471), .CLK(clk), .Q(n2929), .QN(n1380) );
  DFFX1_HVT \keys_reg[4][58]  ( .D(n4470), .CLK(clk), .Q(n2928), .QN(n363) );
  DFFX1_HVT \keys_reg[3][58]  ( .D(n4469), .CLK(clk), .Q(n2927), .QN(n1379) );
  DFFX1_HVT \keys_reg[1][58]  ( .D(n4468), .CLK(clk), .Q(n2926), .QN(n364) );
  DFFX1_HVT \prev_key_reg[58]  ( .D(n5139), .CLK(clk), .Q(prev_key[58]) );
  DFFX1_HVT \keys_reg[10][59]  ( .D(n4467), .CLK(clk), .Q(n2925), .QN(n1016)
         );
  DFFX1_HVT \keys_reg[9][59]  ( .D(n4466), .CLK(clk), .Q(n2924), .QN(n618) );
  DFFX1_HVT \keys_reg[8][59]  ( .D(n4465), .CLK(clk), .Q(n2923), .QN(n1378) );
  DFFX1_HVT \keys_reg[6][59]  ( .D(n4464), .CLK(clk), .Q(n2922), .QN(n617) );
  DFFX1_HVT \keys_reg[5][59]  ( .D(n4463), .CLK(clk), .Q(n2921), .QN(n1377) );
  DFFX1_HVT \keys_reg[4][59]  ( .D(n4462), .CLK(clk), .Q(n2920), .QN(n361) );
  DFFX1_HVT \keys_reg[3][59]  ( .D(n4461), .CLK(clk), .Q(n2919), .QN(n1376) );
  DFFX1_HVT \keys_reg[1][59]  ( .D(n4460), .CLK(clk), .Q(n2918), .QN(n362) );
  DFFX1_HVT \prev_key_reg[59]  ( .D(n5138), .CLK(clk), .Q(prev_key[59]) );
  DFFX1_HVT \keys_reg[10][60]  ( .D(n4459), .CLK(clk), .Q(n2917), .QN(n1015)
         );
  DFFX1_HVT \keys_reg[9][60]  ( .D(n4458), .CLK(clk), .Q(n2916), .QN(n616) );
  DFFX1_HVT \keys_reg[8][60]  ( .D(n4457), .CLK(clk), .Q(n2915), .QN(n1375) );
  DFFX1_HVT \keys_reg[6][60]  ( .D(n4456), .CLK(clk), .Q(n2914), .QN(n615) );
  DFFX1_HVT \keys_reg[5][60]  ( .D(n4455), .CLK(clk), .Q(n2913), .QN(n1374) );
  DFFX1_HVT \keys_reg[4][60]  ( .D(n4454), .CLK(clk), .Q(n2912), .QN(n359) );
  DFFX1_HVT \keys_reg[3][60]  ( .D(n4453), .CLK(clk), .Q(n2911), .QN(n1373) );
  DFFX1_HVT \keys_reg[1][60]  ( .D(n4452), .CLK(clk), .Q(n2910), .QN(n360) );
  DFFX1_HVT \prev_key_reg[60]  ( .D(n5137), .CLK(clk), .Q(prev_key[60]) );
  DFFX1_HVT \keys_reg[10][61]  ( .D(n4451), .CLK(clk), .Q(n2909), .QN(n1014)
         );
  DFFX1_HVT \keys_reg[9][61]  ( .D(n4450), .CLK(clk), .Q(n2908), .QN(n614) );
  DFFX1_HVT \keys_reg[8][61]  ( .D(n4449), .CLK(clk), .Q(n2907), .QN(n1372) );
  DFFX1_HVT \keys_reg[6][61]  ( .D(n4448), .CLK(clk), .Q(n2906), .QN(n613) );
  DFFX1_HVT \keys_reg[5][61]  ( .D(n4447), .CLK(clk), .Q(n2905), .QN(n1371) );
  DFFX1_HVT \keys_reg[4][61]  ( .D(n4446), .CLK(clk), .Q(n2904), .QN(n357) );
  DFFX1_HVT \keys_reg[3][61]  ( .D(n4445), .CLK(clk), .Q(n2903), .QN(n1370) );
  DFFX1_HVT \keys_reg[1][61]  ( .D(n4444), .CLK(clk), .Q(n2902), .QN(n358) );
  DFFX1_HVT \prev_key_reg[61]  ( .D(n5136), .CLK(clk), .Q(prev_key[61]) );
  DFFX1_HVT \keys_reg[10][62]  ( .D(n4443), .CLK(clk), .Q(n2901), .QN(n1013)
         );
  DFFX1_HVT \keys_reg[9][62]  ( .D(n4442), .CLK(clk), .Q(n2900), .QN(n612) );
  DFFX1_HVT \keys_reg[8][62]  ( .D(n4441), .CLK(clk), .Q(n2899), .QN(n1369) );
  DFFX1_HVT \keys_reg[6][62]  ( .D(n4440), .CLK(clk), .Q(n2898), .QN(n611) );
  DFFX1_HVT \keys_reg[5][62]  ( .D(n4439), .CLK(clk), .Q(n2897), .QN(n1368) );
  DFFX1_HVT \keys_reg[4][62]  ( .D(n4438), .CLK(clk), .Q(n2896), .QN(n355) );
  DFFX1_HVT \keys_reg[3][62]  ( .D(n4437), .CLK(clk), .Q(n2895), .QN(n1367) );
  DFFX1_HVT \keys_reg[1][62]  ( .D(n4436), .CLK(clk), .Q(n2894), .QN(n356) );
  DFFX1_HVT \prev_key_reg[62]  ( .D(n5135), .CLK(clk), .Q(prev_key[62]) );
  DFFX1_HVT \keys_reg[10][63]  ( .D(n4435), .CLK(clk), .Q(n2893), .QN(n1012)
         );
  DFFX1_HVT \keys_reg[9][63]  ( .D(n4434), .CLK(clk), .Q(n2892), .QN(n610) );
  DFFX1_HVT \keys_reg[8][63]  ( .D(n4433), .CLK(clk), .Q(n2891), .QN(n1366) );
  DFFX1_HVT \keys_reg[6][63]  ( .D(n4432), .CLK(clk), .Q(n2890), .QN(n609) );
  DFFX1_HVT \keys_reg[5][63]  ( .D(n4431), .CLK(clk), .Q(n2889), .QN(n1365) );
  DFFX1_HVT \keys_reg[4][63]  ( .D(n4430), .CLK(clk), .Q(n2888), .QN(n353) );
  DFFX1_HVT \keys_reg[3][63]  ( .D(n4429), .CLK(clk), .Q(n2887), .QN(n1364) );
  DFFX1_HVT \keys_reg[1][63]  ( .D(n4428), .CLK(clk), .Q(n2886), .QN(n354) );
  DFFX1_HVT \prev_key_reg[63]  ( .D(n5134), .CLK(clk), .Q(prev_key[63]) );
  DFFX1_HVT \keys_reg[10][64]  ( .D(n4427), .CLK(clk), .Q(n2885), .QN(n1011)
         );
  DFFX1_HVT \keys_reg[9][64]  ( .D(n4426), .CLK(clk), .Q(n2884), .QN(n608) );
  DFFX1_HVT \keys_reg[8][64]  ( .D(n4425), .CLK(clk), .Q(n2883), .QN(n1363) );
  DFFX1_HVT \keys_reg[6][64]  ( .D(n4424), .CLK(clk), .Q(n2882), .QN(n607) );
  DFFX1_HVT \keys_reg[5][64]  ( .D(n4423), .CLK(clk), .Q(n2881), .QN(n1362) );
  DFFX1_HVT \keys_reg[4][64]  ( .D(n4422), .CLK(clk), .Q(n2880), .QN(n351) );
  DFFX1_HVT \keys_reg[3][64]  ( .D(n4421), .CLK(clk), .Q(n2879), .QN(n1361) );
  DFFX1_HVT \keys_reg[1][64]  ( .D(n4420), .CLK(clk), .Q(n2878), .QN(n352) );
  DFFX1_HVT \prev_key_reg[64]  ( .D(n5133), .CLK(clk), .Q(prev_key[64]) );
  DFFX1_HVT \keys_reg[10][65]  ( .D(n4419), .CLK(clk), .Q(n2877), .QN(n1010)
         );
  DFFX1_HVT \keys_reg[9][65]  ( .D(n4418), .CLK(clk), .Q(n2876), .QN(n606) );
  DFFX1_HVT \keys_reg[8][65]  ( .D(n4417), .CLK(clk), .Q(n2875), .QN(n1360) );
  DFFX1_HVT \keys_reg[6][65]  ( .D(n4416), .CLK(clk), .Q(n2874), .QN(n605) );
  DFFX1_HVT \keys_reg[5][65]  ( .D(n4415), .CLK(clk), .Q(n2873), .QN(n1359) );
  DFFX1_HVT \keys_reg[4][65]  ( .D(n4414), .CLK(clk), .Q(n2872), .QN(n349) );
  DFFX1_HVT \keys_reg[3][65]  ( .D(n4413), .CLK(clk), .Q(n2871), .QN(n1358) );
  DFFX1_HVT \keys_reg[1][65]  ( .D(n4412), .CLK(clk), .Q(n2870), .QN(n350) );
  DFFX1_HVT \prev_key_reg[65]  ( .D(n5132), .CLK(clk), .Q(prev_key[65]) );
  DFFX1_HVT \keys_reg[10][66]  ( .D(n4411), .CLK(clk), .Q(n2869), .QN(n1009)
         );
  DFFX1_HVT \keys_reg[9][66]  ( .D(n4410), .CLK(clk), .Q(n2868), .QN(n604) );
  DFFX1_HVT \keys_reg[8][66]  ( .D(n4409), .CLK(clk), .Q(n2867), .QN(n1357) );
  DFFX1_HVT \keys_reg[6][66]  ( .D(n4408), .CLK(clk), .Q(n2866), .QN(n603) );
  DFFX1_HVT \keys_reg[5][66]  ( .D(n4407), .CLK(clk), .Q(n2865), .QN(n1356) );
  DFFX1_HVT \keys_reg[4][66]  ( .D(n4406), .CLK(clk), .Q(n2864), .QN(n347) );
  DFFX1_HVT \keys_reg[3][66]  ( .D(n4405), .CLK(clk), .Q(n2863), .QN(n1355) );
  DFFX1_HVT \keys_reg[1][66]  ( .D(n4404), .CLK(clk), .Q(n2862), .QN(n348) );
  DFFX1_HVT \prev_key_reg[66]  ( .D(n5131), .CLK(clk), .Q(prev_key[66]) );
  DFFX1_HVT \keys_reg[10][67]  ( .D(n4403), .CLK(clk), .Q(n2861), .QN(n1008)
         );
  DFFX1_HVT \keys_reg[9][67]  ( .D(n4402), .CLK(clk), .Q(n2860), .QN(n602) );
  DFFX1_HVT \keys_reg[8][67]  ( .D(n4401), .CLK(clk), .Q(n2859), .QN(n1354) );
  DFFX1_HVT \keys_reg[6][67]  ( .D(n4400), .CLK(clk), .Q(n2858), .QN(n601) );
  DFFX1_HVT \keys_reg[5][67]  ( .D(n4399), .CLK(clk), .Q(n2857), .QN(n1353) );
  DFFX1_HVT \keys_reg[4][67]  ( .D(n4398), .CLK(clk), .Q(n2856), .QN(n345) );
  DFFX1_HVT \keys_reg[3][67]  ( .D(n4397), .CLK(clk), .Q(n2855), .QN(n1352) );
  DFFX1_HVT \keys_reg[1][67]  ( .D(n4396), .CLK(clk), .Q(n2854), .QN(n346) );
  DFFX1_HVT \prev_key_reg[67]  ( .D(n5130), .CLK(clk), .Q(prev_key[67]) );
  DFFX1_HVT \keys_reg[10][68]  ( .D(n4395), .CLK(clk), .Q(n2853), .QN(n1007)
         );
  DFFX1_HVT \keys_reg[9][68]  ( .D(n4394), .CLK(clk), .Q(n2852), .QN(n600) );
  DFFX1_HVT \keys_reg[8][68]  ( .D(n4393), .CLK(clk), .Q(n2851), .QN(n1351) );
  DFFX1_HVT \keys_reg[6][68]  ( .D(n4392), .CLK(clk), .Q(n2850), .QN(n599) );
  DFFX1_HVT \keys_reg[5][68]  ( .D(n4391), .CLK(clk), .Q(n2849), .QN(n1350) );
  DFFX1_HVT \keys_reg[4][68]  ( .D(n4390), .CLK(clk), .Q(n2848), .QN(n343) );
  DFFX1_HVT \keys_reg[3][68]  ( .D(n4389), .CLK(clk), .Q(n2847), .QN(n1349) );
  DFFX1_HVT \keys_reg[1][68]  ( .D(n4388), .CLK(clk), .Q(n2846), .QN(n344) );
  DFFX1_HVT \prev_key_reg[68]  ( .D(n5129), .CLK(clk), .Q(prev_key[68]) );
  DFFX1_HVT \keys_reg[10][69]  ( .D(n4387), .CLK(clk), .Q(n2845), .QN(n1006)
         );
  DFFX1_HVT \keys_reg[9][69]  ( .D(n4386), .CLK(clk), .Q(n2844), .QN(n598) );
  DFFX1_HVT \keys_reg[8][69]  ( .D(n4385), .CLK(clk), .Q(n2843), .QN(n1348) );
  DFFX1_HVT \keys_reg[6][69]  ( .D(n4384), .CLK(clk), .Q(n2842), .QN(n597) );
  DFFX1_HVT \keys_reg[5][69]  ( .D(n4383), .CLK(clk), .Q(n2841), .QN(n1347) );
  DFFX1_HVT \keys_reg[4][69]  ( .D(n4382), .CLK(clk), .Q(n2840), .QN(n341) );
  DFFX1_HVT \keys_reg[3][69]  ( .D(n4381), .CLK(clk), .Q(n2839), .QN(n1346) );
  DFFX1_HVT \keys_reg[1][69]  ( .D(n4380), .CLK(clk), .Q(n2838), .QN(n342) );
  DFFX1_HVT \prev_key_reg[69]  ( .D(n5128), .CLK(clk), .Q(prev_key[69]) );
  DFFX1_HVT \keys_reg[10][70]  ( .D(n4379), .CLK(clk), .Q(n2837), .QN(n1005)
         );
  DFFX1_HVT \keys_reg[9][70]  ( .D(n4378), .CLK(clk), .Q(n2836), .QN(n596) );
  DFFX1_HVT \keys_reg[8][70]  ( .D(n4377), .CLK(clk), .Q(n2835), .QN(n1345) );
  DFFX1_HVT \keys_reg[6][70]  ( .D(n4376), .CLK(clk), .Q(n2834), .QN(n595) );
  DFFX1_HVT \keys_reg[5][70]  ( .D(n4375), .CLK(clk), .Q(n2833), .QN(n1344) );
  DFFX1_HVT \keys_reg[4][70]  ( .D(n4374), .CLK(clk), .Q(n2832), .QN(n339) );
  DFFX1_HVT \keys_reg[3][70]  ( .D(n4373), .CLK(clk), .Q(n2831), .QN(n1343) );
  DFFX1_HVT \keys_reg[1][70]  ( .D(n4372), .CLK(clk), .Q(n2830), .QN(n340) );
  DFFX1_HVT \prev_key_reg[70]  ( .D(n5127), .CLK(clk), .Q(prev_key[70]) );
  DFFX1_HVT \keys_reg[10][71]  ( .D(n4371), .CLK(clk), .Q(n2829), .QN(n1004)
         );
  DFFX1_HVT \keys_reg[9][71]  ( .D(n4370), .CLK(clk), .Q(n2828), .QN(n594) );
  DFFX1_HVT \keys_reg[8][71]  ( .D(n4369), .CLK(clk), .Q(n2827), .QN(n1342) );
  DFFX1_HVT \keys_reg[6][71]  ( .D(n4368), .CLK(clk), .Q(n2826), .QN(n593) );
  DFFX1_HVT \keys_reg[5][71]  ( .D(n4367), .CLK(clk), .Q(n2825), .QN(n1341) );
  DFFX1_HVT \keys_reg[4][71]  ( .D(n4366), .CLK(clk), .Q(n2824), .QN(n337) );
  DFFX1_HVT \keys_reg[3][71]  ( .D(n4365), .CLK(clk), .Q(n2823), .QN(n1340) );
  DFFX1_HVT \keys_reg[1][71]  ( .D(n4364), .CLK(clk), .Q(n2822), .QN(n338) );
  DFFX1_HVT \prev_key_reg[71]  ( .D(n5126), .CLK(clk), .Q(prev_key[71]) );
  DFFX1_HVT \keys_reg[10][72]  ( .D(n4363), .CLK(clk), .Q(n2821), .QN(n1003)
         );
  DFFX1_HVT \keys_reg[9][72]  ( .D(n4362), .CLK(clk), .Q(n2820), .QN(n592) );
  DFFX1_HVT \keys_reg[8][72]  ( .D(n4361), .CLK(clk), .Q(n2819), .QN(n1339) );
  DFFX1_HVT \keys_reg[6][72]  ( .D(n4360), .CLK(clk), .Q(n2818), .QN(n591) );
  DFFX1_HVT \keys_reg[5][72]  ( .D(n4359), .CLK(clk), .Q(n2817), .QN(n1338) );
  DFFX1_HVT \keys_reg[4][72]  ( .D(n4358), .CLK(clk), .Q(n2816), .QN(n335) );
  DFFX1_HVT \keys_reg[3][72]  ( .D(n4357), .CLK(clk), .Q(n2815), .QN(n1337) );
  DFFX1_HVT \keys_reg[1][72]  ( .D(n4356), .CLK(clk), .Q(n2814), .QN(n336) );
  DFFX1_HVT \prev_key_reg[72]  ( .D(n5125), .CLK(clk), .Q(prev_key[72]) );
  DFFX1_HVT \keys_reg[10][73]  ( .D(n4355), .CLK(clk), .Q(n2813), .QN(n1002)
         );
  DFFX1_HVT \keys_reg[9][73]  ( .D(n4354), .CLK(clk), .Q(n2812), .QN(n590) );
  DFFX1_HVT \keys_reg[8][73]  ( .D(n4353), .CLK(clk), .Q(n2811), .QN(n1336) );
  DFFX1_HVT \keys_reg[6][73]  ( .D(n4352), .CLK(clk), .Q(n2810), .QN(n589) );
  DFFX1_HVT \keys_reg[5][73]  ( .D(n4351), .CLK(clk), .Q(n2809), .QN(n1335) );
  DFFX1_HVT \keys_reg[4][73]  ( .D(n4350), .CLK(clk), .Q(n2808), .QN(n333) );
  DFFX1_HVT \keys_reg[3][73]  ( .D(n4349), .CLK(clk), .Q(n2807), .QN(n1334) );
  DFFX1_HVT \keys_reg[1][73]  ( .D(n4348), .CLK(clk), .Q(n2806), .QN(n334) );
  DFFX1_HVT \prev_key_reg[73]  ( .D(n5124), .CLK(clk), .Q(prev_key[73]) );
  DFFX1_HVT \keys_reg[10][74]  ( .D(n4347), .CLK(clk), .Q(n2805), .QN(n1001)
         );
  DFFX1_HVT \keys_reg[9][74]  ( .D(n4346), .CLK(clk), .Q(n2804), .QN(n588) );
  DFFX1_HVT \keys_reg[8][74]  ( .D(n4345), .CLK(clk), .Q(n2803), .QN(n1333) );
  DFFX1_HVT \keys_reg[6][74]  ( .D(n4344), .CLK(clk), .Q(n2802), .QN(n587) );
  DFFX1_HVT \keys_reg[5][74]  ( .D(n4343), .CLK(clk), .Q(n2801), .QN(n1332) );
  DFFX1_HVT \keys_reg[4][74]  ( .D(n4342), .CLK(clk), .Q(n2800), .QN(n331) );
  DFFX1_HVT \keys_reg[3][74]  ( .D(n4341), .CLK(clk), .Q(n2799), .QN(n1331) );
  DFFX1_HVT \keys_reg[1][74]  ( .D(n4340), .CLK(clk), .Q(n2798), .QN(n332) );
  DFFX1_HVT \prev_key_reg[74]  ( .D(n5123), .CLK(clk), .Q(prev_key[74]) );
  DFFX1_HVT \keys_reg[10][75]  ( .D(n4339), .CLK(clk), .Q(n2797), .QN(n1000)
         );
  DFFX1_HVT \keys_reg[9][75]  ( .D(n4338), .CLK(clk), .Q(n2796), .QN(n586) );
  DFFX1_HVT \keys_reg[8][75]  ( .D(n4337), .CLK(clk), .Q(n2795), .QN(n1330) );
  DFFX1_HVT \keys_reg[6][75]  ( .D(n4336), .CLK(clk), .Q(n2794), .QN(n585) );
  DFFX1_HVT \keys_reg[5][75]  ( .D(n4335), .CLK(clk), .Q(n2793), .QN(n1329) );
  DFFX1_HVT \keys_reg[4][75]  ( .D(n4334), .CLK(clk), .Q(n2792), .QN(n329) );
  DFFX1_HVT \keys_reg[3][75]  ( .D(n4333), .CLK(clk), .Q(n2791), .QN(n1328) );
  DFFX1_HVT \keys_reg[1][75]  ( .D(n4332), .CLK(clk), .Q(n2790), .QN(n330) );
  DFFX1_HVT \prev_key_reg[75]  ( .D(n5122), .CLK(clk), .Q(prev_key[75]) );
  DFFX1_HVT \keys_reg[10][76]  ( .D(n4331), .CLK(clk), .Q(n2789), .QN(n999) );
  DFFX1_HVT \keys_reg[9][76]  ( .D(n4330), .CLK(clk), .Q(n2788), .QN(n584) );
  DFFX1_HVT \keys_reg[8][76]  ( .D(n4329), .CLK(clk), .Q(n2787), .QN(n1327) );
  DFFX1_HVT \keys_reg[6][76]  ( .D(n4328), .CLK(clk), .Q(n2786), .QN(n583) );
  DFFX1_HVT \keys_reg[5][76]  ( .D(n4327), .CLK(clk), .Q(n2785), .QN(n1326) );
  DFFX1_HVT \keys_reg[4][76]  ( .D(n4326), .CLK(clk), .Q(n2784), .QN(n327) );
  DFFX1_HVT \keys_reg[3][76]  ( .D(n4325), .CLK(clk), .Q(n2783), .QN(n1325) );
  DFFX1_HVT \keys_reg[1][76]  ( .D(n4324), .CLK(clk), .Q(n2782), .QN(n328) );
  DFFX1_HVT \prev_key_reg[76]  ( .D(n5121), .CLK(clk), .Q(prev_key[76]) );
  DFFX1_HVT \keys_reg[10][77]  ( .D(n4323), .CLK(clk), .Q(n2781), .QN(n998) );
  DFFX1_HVT \keys_reg[9][77]  ( .D(n4322), .CLK(clk), .Q(n2780), .QN(n582) );
  DFFX1_HVT \keys_reg[8][77]  ( .D(n4321), .CLK(clk), .Q(n2779), .QN(n1324) );
  DFFX1_HVT \keys_reg[6][77]  ( .D(n4320), .CLK(clk), .Q(n2778), .QN(n581) );
  DFFX1_HVT \keys_reg[5][77]  ( .D(n4319), .CLK(clk), .Q(n2777), .QN(n1323) );
  DFFX1_HVT \keys_reg[4][77]  ( .D(n4318), .CLK(clk), .Q(n2776), .QN(n325) );
  DFFX1_HVT \keys_reg[3][77]  ( .D(n4317), .CLK(clk), .Q(n2775), .QN(n1322) );
  DFFX1_HVT \keys_reg[1][77]  ( .D(n4316), .CLK(clk), .Q(n2774), .QN(n326) );
  DFFX1_HVT \prev_key_reg[77]  ( .D(n5120), .CLK(clk), .Q(prev_key[77]) );
  DFFX1_HVT \keys_reg[10][78]  ( .D(n4315), .CLK(clk), .Q(n2773), .QN(n997) );
  DFFX1_HVT \keys_reg[9][78]  ( .D(n4314), .CLK(clk), .Q(n2772), .QN(n580) );
  DFFX1_HVT \keys_reg[8][78]  ( .D(n4313), .CLK(clk), .Q(n2771), .QN(n1321) );
  DFFX1_HVT \keys_reg[6][78]  ( .D(n4312), .CLK(clk), .Q(n2770), .QN(n579) );
  DFFX1_HVT \keys_reg[5][78]  ( .D(n4311), .CLK(clk), .Q(n2769), .QN(n1320) );
  DFFX1_HVT \keys_reg[4][78]  ( .D(n4310), .CLK(clk), .Q(n2768), .QN(n323) );
  DFFX1_HVT \keys_reg[3][78]  ( .D(n4309), .CLK(clk), .Q(n2767), .QN(n1319) );
  DFFX1_HVT \keys_reg[1][78]  ( .D(n4308), .CLK(clk), .Q(n2766), .QN(n324) );
  DFFX1_HVT \prev_key_reg[78]  ( .D(n5119), .CLK(clk), .Q(prev_key[78]) );
  DFFX1_HVT \keys_reg[10][79]  ( .D(n4307), .CLK(clk), .Q(n2765), .QN(n996) );
  DFFX1_HVT \keys_reg[9][79]  ( .D(n4306), .CLK(clk), .Q(n2764), .QN(n578) );
  DFFX1_HVT \keys_reg[8][79]  ( .D(n4305), .CLK(clk), .Q(n2763), .QN(n1318) );
  DFFX1_HVT \keys_reg[6][79]  ( .D(n4304), .CLK(clk), .Q(n2762), .QN(n577) );
  DFFX1_HVT \keys_reg[5][79]  ( .D(n4303), .CLK(clk), .Q(n2761), .QN(n1317) );
  DFFX1_HVT \keys_reg[4][79]  ( .D(n4302), .CLK(clk), .Q(n2760), .QN(n321) );
  DFFX1_HVT \keys_reg[3][79]  ( .D(n4301), .CLK(clk), .Q(n2759), .QN(n1316) );
  DFFX1_HVT \keys_reg[1][79]  ( .D(n4300), .CLK(clk), .Q(n2758), .QN(n322) );
  DFFX1_HVT \prev_key_reg[79]  ( .D(n5118), .CLK(clk), .Q(prev_key[79]) );
  DFFX1_HVT \keys_reg[10][80]  ( .D(n4299), .CLK(clk), .Q(n2757), .QN(n995) );
  DFFX1_HVT \keys_reg[9][80]  ( .D(n4298), .CLK(clk), .Q(n2756), .QN(n576) );
  DFFX1_HVT \keys_reg[8][80]  ( .D(n4297), .CLK(clk), .Q(n2755), .QN(n1315) );
  DFFX1_HVT \keys_reg[6][80]  ( .D(n4296), .CLK(clk), .Q(n2754), .QN(n575) );
  DFFX1_HVT \keys_reg[5][80]  ( .D(n4295), .CLK(clk), .Q(n2753), .QN(n1314) );
  DFFX1_HVT \keys_reg[4][80]  ( .D(n4294), .CLK(clk), .Q(n2752), .QN(n319) );
  DFFX1_HVT \keys_reg[3][80]  ( .D(n4293), .CLK(clk), .Q(n2751), .QN(n1313) );
  DFFX1_HVT \keys_reg[1][80]  ( .D(n4292), .CLK(clk), .Q(n2750), .QN(n320) );
  DFFX1_HVT \prev_key_reg[80]  ( .D(n5117), .CLK(clk), .Q(prev_key[80]) );
  DFFX1_HVT \keys_reg[10][81]  ( .D(n4291), .CLK(clk), .Q(n2749), .QN(n994) );
  DFFX1_HVT \keys_reg[9][81]  ( .D(n4290), .CLK(clk), .Q(n2748), .QN(n574) );
  DFFX1_HVT \keys_reg[8][81]  ( .D(n4289), .CLK(clk), .Q(n2747), .QN(n1312) );
  DFFX1_HVT \keys_reg[6][81]  ( .D(n4288), .CLK(clk), .Q(n2746), .QN(n573) );
  DFFX1_HVT \keys_reg[5][81]  ( .D(n4287), .CLK(clk), .Q(n2745), .QN(n1311) );
  DFFX1_HVT \keys_reg[4][81]  ( .D(n4286), .CLK(clk), .Q(n2744), .QN(n317) );
  DFFX1_HVT \keys_reg[3][81]  ( .D(n4285), .CLK(clk), .Q(n2743), .QN(n1310) );
  DFFX1_HVT \keys_reg[1][81]  ( .D(n4284), .CLK(clk), .Q(n2742), .QN(n318) );
  DFFX1_HVT \prev_key_reg[81]  ( .D(n5116), .CLK(clk), .Q(prev_key[81]) );
  DFFX1_HVT \keys_reg[10][82]  ( .D(n4283), .CLK(clk), .Q(n2741), .QN(n929) );
  DFFX1_HVT \keys_reg[9][82]  ( .D(n4282), .CLK(clk), .Q(n2740), .QN(n444) );
  DFFX1_HVT \keys_reg[8][82]  ( .D(n4281), .CLK(clk), .Q(n2739), .QN(n1117) );
  DFFX1_HVT \keys_reg[6][82]  ( .D(n4280), .CLK(clk), .Q(n2738), .QN(n443) );
  DFFX1_HVT \keys_reg[5][82]  ( .D(n4279), .CLK(clk), .Q(n2737), .QN(n1116) );
  DFFX1_HVT \keys_reg[4][82]  ( .D(n4278), .CLK(clk), .Q(n2736), .QN(n187) );
  DFFX1_HVT \keys_reg[3][82]  ( .D(n4277), .CLK(clk), .Q(n2735), .QN(n1115) );
  DFFX1_HVT \keys_reg[1][82]  ( .D(n4276), .CLK(clk), .Q(n2734), .QN(n188) );
  DFFX1_HVT \prev_key_reg[82]  ( .D(n5115), .CLK(clk), .Q(prev_key[82]) );
  DFFX1_HVT \keys_reg[10][83]  ( .D(n4275), .CLK(clk), .Q(n2733), .QN(n930) );
  DFFX1_HVT \keys_reg[9][83]  ( .D(n4274), .CLK(clk), .Q(n2732), .QN(n446) );
  DFFX1_HVT \keys_reg[8][83]  ( .D(n4273), .CLK(clk), .Q(n2731), .QN(n1120) );
  DFFX1_HVT \keys_reg[6][83]  ( .D(n4272), .CLK(clk), .Q(n2730), .QN(n445) );
  DFFX1_HVT \keys_reg[5][83]  ( .D(n4271), .CLK(clk), .Q(n2729), .QN(n1119) );
  DFFX1_HVT \keys_reg[4][83]  ( .D(n4270), .CLK(clk), .Q(n2728), .QN(n189) );
  DFFX1_HVT \keys_reg[3][83]  ( .D(n4269), .CLK(clk), .Q(n2727), .QN(n1118) );
  DFFX1_HVT \keys_reg[1][83]  ( .D(n4268), .CLK(clk), .Q(n2726), .QN(n190) );
  DFFX1_HVT \prev_key_reg[83]  ( .D(n5114), .CLK(clk), .Q(prev_key[83]) );
  DFFX1_HVT \keys_reg[10][84]  ( .D(n4267), .CLK(clk), .Q(n2725), .QN(n931) );
  DFFX1_HVT \keys_reg[9][84]  ( .D(n4266), .CLK(clk), .Q(n2724), .QN(n448) );
  DFFX1_HVT \keys_reg[8][84]  ( .D(n4265), .CLK(clk), .Q(n2723), .QN(n1123) );
  DFFX1_HVT \keys_reg[6][84]  ( .D(n4264), .CLK(clk), .Q(n2722), .QN(n447) );
  DFFX1_HVT \keys_reg[5][84]  ( .D(n4263), .CLK(clk), .Q(n2721), .QN(n1122) );
  DFFX1_HVT \keys_reg[4][84]  ( .D(n4262), .CLK(clk), .Q(n2720), .QN(n191) );
  DFFX1_HVT \keys_reg[3][84]  ( .D(n4261), .CLK(clk), .Q(n2719), .QN(n1121) );
  DFFX1_HVT \keys_reg[1][84]  ( .D(n4260), .CLK(clk), .Q(n2718), .QN(n192) );
  DFFX1_HVT \prev_key_reg[84]  ( .D(n5113), .CLK(clk), .Q(prev_key[84]) );
  DFFX1_HVT \keys_reg[10][85]  ( .D(n4259), .CLK(clk), .Q(n2717), .QN(n932) );
  DFFX1_HVT \keys_reg[9][85]  ( .D(n4258), .CLK(clk), .Q(n2716), .QN(n450) );
  DFFX1_HVT \keys_reg[8][85]  ( .D(n4257), .CLK(clk), .Q(n2715), .QN(n1126) );
  DFFX1_HVT \keys_reg[6][85]  ( .D(n4256), .CLK(clk), .Q(n2714), .QN(n449) );
  DFFX1_HVT \keys_reg[5][85]  ( .D(n4255), .CLK(clk), .Q(n2713), .QN(n1125) );
  DFFX1_HVT \keys_reg[4][85]  ( .D(n4254), .CLK(clk), .Q(n2712), .QN(n193) );
  DFFX1_HVT \keys_reg[3][85]  ( .D(n4253), .CLK(clk), .Q(n2711), .QN(n1124) );
  DFFX1_HVT \keys_reg[1][85]  ( .D(n4252), .CLK(clk), .Q(n2710), .QN(n194) );
  DFFX1_HVT \prev_key_reg[85]  ( .D(n5112), .CLK(clk), .Q(prev_key[85]) );
  DFFX1_HVT \keys_reg[10][86]  ( .D(n4251), .CLK(clk), .Q(n2709), .QN(n933) );
  DFFX1_HVT \keys_reg[9][86]  ( .D(n4250), .CLK(clk), .Q(n2708), .QN(n452) );
  DFFX1_HVT \keys_reg[8][86]  ( .D(n4249), .CLK(clk), .Q(n2707), .QN(n1129) );
  DFFX1_HVT \keys_reg[6][86]  ( .D(n4248), .CLK(clk), .Q(n2706), .QN(n451) );
  DFFX1_HVT \keys_reg[5][86]  ( .D(n4247), .CLK(clk), .Q(n2705), .QN(n1128) );
  DFFX1_HVT \keys_reg[4][86]  ( .D(n4246), .CLK(clk), .Q(n2704), .QN(n195) );
  DFFX1_HVT \keys_reg[3][86]  ( .D(n4245), .CLK(clk), .Q(n2703), .QN(n1127) );
  DFFX1_HVT \keys_reg[1][86]  ( .D(n4244), .CLK(clk), .Q(n2702), .QN(n196) );
  DFFX1_HVT \prev_key_reg[86]  ( .D(n5111), .CLK(clk), .Q(prev_key[86]) );
  DFFX1_HVT \keys_reg[10][87]  ( .D(n4243), .CLK(clk), .Q(n2701), .QN(n934) );
  DFFX1_HVT \keys_reg[9][87]  ( .D(n4242), .CLK(clk), .Q(n2700), .QN(n454) );
  DFFX1_HVT \keys_reg[8][87]  ( .D(n4241), .CLK(clk), .Q(n2699), .QN(n1132) );
  DFFX1_HVT \keys_reg[6][87]  ( .D(n4240), .CLK(clk), .Q(n2698), .QN(n453) );
  DFFX1_HVT \keys_reg[5][87]  ( .D(n4239), .CLK(clk), .Q(n2697), .QN(n1131) );
  DFFX1_HVT \keys_reg[4][87]  ( .D(n4238), .CLK(clk), .Q(n2696), .QN(n197) );
  DFFX1_HVT \keys_reg[3][87]  ( .D(n4237), .CLK(clk), .Q(n2695), .QN(n1130) );
  DFFX1_HVT \keys_reg[1][87]  ( .D(n4236), .CLK(clk), .Q(n2694), .QN(n198) );
  DFFX1_HVT \prev_key_reg[87]  ( .D(n5110), .CLK(clk), .Q(prev_key[87]) );
  DFFX1_HVT \keys_reg[10][88]  ( .D(n4235), .CLK(clk), .Q(n2693), .QN(n935) );
  DFFX1_HVT \keys_reg[9][88]  ( .D(n4234), .CLK(clk), .Q(n2692), .QN(n456) );
  DFFX1_HVT \keys_reg[8][88]  ( .D(n4233), .CLK(clk), .Q(n2691), .QN(n1135) );
  DFFX1_HVT \keys_reg[6][88]  ( .D(n4232), .CLK(clk), .Q(n2690), .QN(n455) );
  DFFX1_HVT \keys_reg[5][88]  ( .D(n4231), .CLK(clk), .Q(n2689), .QN(n1134) );
  DFFX1_HVT \keys_reg[4][88]  ( .D(n4230), .CLK(clk), .Q(n2688), .QN(n199) );
  DFFX1_HVT \keys_reg[3][88]  ( .D(n4229), .CLK(clk), .Q(n2687), .QN(n1133) );
  DFFX1_HVT \keys_reg[1][88]  ( .D(n4228), .CLK(clk), .Q(n2686), .QN(n200) );
  DFFX1_HVT \prev_key_reg[88]  ( .D(n5109), .CLK(clk), .Q(prev_key[88]) );
  DFFX1_HVT \keys_reg[10][89]  ( .D(n4227), .CLK(clk), .Q(n2685), .QN(n936) );
  DFFX1_HVT \keys_reg[9][89]  ( .D(n4226), .CLK(clk), .Q(n2684), .QN(n458) );
  DFFX1_HVT \keys_reg[8][89]  ( .D(n4225), .CLK(clk), .Q(n2683), .QN(n1138) );
  DFFX1_HVT \keys_reg[6][89]  ( .D(n4224), .CLK(clk), .Q(n2682), .QN(n457) );
  DFFX1_HVT \keys_reg[5][89]  ( .D(n4223), .CLK(clk), .Q(n2681), .QN(n1137) );
  DFFX1_HVT \keys_reg[4][89]  ( .D(n4222), .CLK(clk), .Q(n2680), .QN(n201) );
  DFFX1_HVT \keys_reg[3][89]  ( .D(n4221), .CLK(clk), .Q(n2679), .QN(n1136) );
  DFFX1_HVT \keys_reg[1][89]  ( .D(n4220), .CLK(clk), .Q(n2678), .QN(n202) );
  DFFX1_HVT \prev_key_reg[89]  ( .D(n5108), .CLK(clk), .Q(prev_key[89]) );
  DFFX1_HVT \keys_reg[10][90]  ( .D(n4219), .CLK(clk), .Q(n2677), .QN(n937) );
  DFFX1_HVT \keys_reg[9][90]  ( .D(n4218), .CLK(clk), .Q(n2676), .QN(n460) );
  DFFX1_HVT \keys_reg[8][90]  ( .D(n4217), .CLK(clk), .Q(n2675), .QN(n1141) );
  DFFX1_HVT \keys_reg[6][90]  ( .D(n4216), .CLK(clk), .Q(n2674), .QN(n459) );
  DFFX1_HVT \keys_reg[5][90]  ( .D(n4215), .CLK(clk), .Q(n2673), .QN(n1140) );
  DFFX1_HVT \keys_reg[4][90]  ( .D(n4214), .CLK(clk), .Q(n2672), .QN(n203) );
  DFFX1_HVT \keys_reg[3][90]  ( .D(n4213), .CLK(clk), .Q(n2671), .QN(n1139) );
  DFFX1_HVT \keys_reg[1][90]  ( .D(n4212), .CLK(clk), .Q(n2670), .QN(n204) );
  DFFX1_HVT \prev_key_reg[90]  ( .D(n5107), .CLK(clk), .Q(prev_key[90]) );
  DFFX1_HVT \keys_reg[10][91]  ( .D(n4211), .CLK(clk), .Q(n2669), .QN(n938) );
  DFFX1_HVT \keys_reg[9][91]  ( .D(n4210), .CLK(clk), .Q(n2668), .QN(n462) );
  DFFX1_HVT \keys_reg[8][91]  ( .D(n4209), .CLK(clk), .Q(n2667), .QN(n1144) );
  DFFX1_HVT \keys_reg[6][91]  ( .D(n4208), .CLK(clk), .Q(n2666), .QN(n461) );
  DFFX1_HVT \keys_reg[5][91]  ( .D(n4207), .CLK(clk), .Q(n2665), .QN(n1143) );
  DFFX1_HVT \keys_reg[4][91]  ( .D(n4206), .CLK(clk), .Q(n2664), .QN(n205) );
  DFFX1_HVT \keys_reg[3][91]  ( .D(n4205), .CLK(clk), .Q(n2663), .QN(n1142) );
  DFFX1_HVT \keys_reg[1][91]  ( .D(n4204), .CLK(clk), .Q(n2662), .QN(n206) );
  DFFX1_HVT \prev_key_reg[91]  ( .D(n5106), .CLK(clk), .Q(prev_key[91]) );
  DFFX1_HVT \keys_reg[10][92]  ( .D(n4203), .CLK(clk), .Q(n2661), .QN(n939) );
  DFFX1_HVT \keys_reg[9][92]  ( .D(n4202), .CLK(clk), .Q(n2660), .QN(n464) );
  DFFX1_HVT \keys_reg[8][92]  ( .D(n4201), .CLK(clk), .Q(n2659), .QN(n1147) );
  DFFX1_HVT \keys_reg[6][92]  ( .D(n4200), .CLK(clk), .Q(n2658), .QN(n463) );
  DFFX1_HVT \keys_reg[5][92]  ( .D(n4199), .CLK(clk), .Q(n2657), .QN(n1146) );
  DFFX1_HVT \keys_reg[4][92]  ( .D(n4198), .CLK(clk), .Q(n2656), .QN(n207) );
  DFFX1_HVT \keys_reg[3][92]  ( .D(n4197), .CLK(clk), .Q(n2655), .QN(n1145) );
  DFFX1_HVT \keys_reg[1][92]  ( .D(n4196), .CLK(clk), .Q(n2654), .QN(n208) );
  DFFX1_HVT \prev_key_reg[92]  ( .D(n5105), .CLK(clk), .Q(prev_key[92]) );
  DFFX1_HVT \keys_reg[10][93]  ( .D(n4195), .CLK(clk), .Q(n2653), .QN(n940) );
  DFFX1_HVT \keys_reg[9][93]  ( .D(n4194), .CLK(clk), .Q(n2652), .QN(n466) );
  DFFX1_HVT \keys_reg[8][93]  ( .D(n4193), .CLK(clk), .Q(n2651), .QN(n1150) );
  DFFX1_HVT \keys_reg[6][93]  ( .D(n4192), .CLK(clk), .Q(n2650), .QN(n465) );
  DFFX1_HVT \keys_reg[5][93]  ( .D(n4191), .CLK(clk), .Q(n2649), .QN(n1149) );
  DFFX1_HVT \keys_reg[4][93]  ( .D(n4190), .CLK(clk), .Q(n2648), .QN(n209) );
  DFFX1_HVT \keys_reg[3][93]  ( .D(n4189), .CLK(clk), .Q(n2647), .QN(n1148) );
  DFFX1_HVT \keys_reg[1][93]  ( .D(n4188), .CLK(clk), .Q(n2646), .QN(n210) );
  DFFX1_HVT \prev_key_reg[93]  ( .D(n5104), .CLK(clk), .Q(prev_key[93]) );
  DFFX1_HVT \keys_reg[10][94]  ( .D(n4187), .CLK(clk), .Q(n2645), .QN(n941) );
  DFFX1_HVT \keys_reg[9][94]  ( .D(n4186), .CLK(clk), .Q(n2644), .QN(n468) );
  DFFX1_HVT \keys_reg[8][94]  ( .D(n4185), .CLK(clk), .Q(n2643), .QN(n1153) );
  DFFX1_HVT \keys_reg[6][94]  ( .D(n4184), .CLK(clk), .Q(n2642), .QN(n467) );
  DFFX1_HVT \keys_reg[5][94]  ( .D(n4183), .CLK(clk), .Q(n2641), .QN(n1152) );
  DFFX1_HVT \keys_reg[4][94]  ( .D(n4182), .CLK(clk), .Q(n2640), .QN(n211) );
  DFFX1_HVT \keys_reg[3][94]  ( .D(n4181), .CLK(clk), .Q(n2639), .QN(n1151) );
  DFFX1_HVT \keys_reg[1][94]  ( .D(n4180), .CLK(clk), .Q(n2638), .QN(n212) );
  DFFX1_HVT \prev_key_reg[94]  ( .D(n5103), .CLK(clk), .Q(prev_key[94]) );
  DFFX1_HVT \keys_reg[10][95]  ( .D(n4179), .CLK(clk), .Q(n2637), .QN(n942) );
  DFFX1_HVT \keys_reg[9][95]  ( .D(n4178), .CLK(clk), .Q(n2636), .QN(n470) );
  DFFX1_HVT \keys_reg[8][95]  ( .D(n4177), .CLK(clk), .Q(n2635), .QN(n1156) );
  DFFX1_HVT \keys_reg[6][95]  ( .D(n4176), .CLK(clk), .Q(n2634), .QN(n469) );
  DFFX1_HVT \keys_reg[5][95]  ( .D(n4175), .CLK(clk), .Q(n2633), .QN(n1155) );
  DFFX1_HVT \keys_reg[4][95]  ( .D(n4174), .CLK(clk), .Q(n2632), .QN(n213) );
  DFFX1_HVT \keys_reg[3][95]  ( .D(n4173), .CLK(clk), .Q(n2631), .QN(n1154) );
  DFFX1_HVT \keys_reg[1][95]  ( .D(n4172), .CLK(clk), .Q(n2630), .QN(n214) );
  DFFX1_HVT \prev_key_reg[95]  ( .D(n5102), .CLK(clk), .Q(prev_key[95]) );
  DFFX1_HVT \keys_reg[10][96]  ( .D(n4171), .CLK(clk), .Q(n2629), .QN(n943) );
  DFFX1_HVT \keys_reg[9][96]  ( .D(n4170), .CLK(clk), .Q(n2628), .QN(n472) );
  DFFX1_HVT \keys_reg[8][96]  ( .D(n4169), .CLK(clk), .Q(n2627), .QN(n1159) );
  DFFX1_HVT \keys_reg[6][96]  ( .D(n4168), .CLK(clk), .Q(n2626), .QN(n471) );
  DFFX1_HVT \keys_reg[5][96]  ( .D(n4167), .CLK(clk), .Q(n2625), .QN(n1158) );
  DFFX1_HVT \keys_reg[4][96]  ( .D(n4166), .CLK(clk), .Q(n2624), .QN(n215) );
  DFFX1_HVT \keys_reg[3][96]  ( .D(n4165), .CLK(clk), .Q(n2623), .QN(n1157) );
  DFFX1_HVT \keys_reg[1][96]  ( .D(n4164), .CLK(clk), .Q(n2622), .QN(n216) );
  DFFX1_HVT \prev_key_reg[96]  ( .D(n5101), .CLK(clk), .Q(prev_key[96]) );
  DFFX1_HVT \keys_reg[10][97]  ( .D(n4163), .CLK(clk), .Q(n2621), .QN(n944) );
  DFFX1_HVT \keys_reg[9][97]  ( .D(n4162), .CLK(clk), .Q(n2620), .QN(n474) );
  DFFX1_HVT \keys_reg[8][97]  ( .D(n4161), .CLK(clk), .Q(n2619), .QN(n1162) );
  DFFX1_HVT \keys_reg[6][97]  ( .D(n4160), .CLK(clk), .Q(n2618), .QN(n473) );
  DFFX1_HVT \keys_reg[5][97]  ( .D(n4159), .CLK(clk), .Q(n2617), .QN(n1161) );
  DFFX1_HVT \keys_reg[4][97]  ( .D(n4158), .CLK(clk), .Q(n2616), .QN(n217) );
  DFFX1_HVT \keys_reg[3][97]  ( .D(n4157), .CLK(clk), .Q(n2615), .QN(n1160) );
  DFFX1_HVT \keys_reg[1][97]  ( .D(n4156), .CLK(clk), .Q(n2614), .QN(n218) );
  DFFX1_HVT \prev_key_reg[97]  ( .D(n5100), .CLK(clk), .Q(prev_key[97]) );
  DFFX1_HVT \keys_reg[10][98]  ( .D(n4155), .CLK(clk), .Q(n2613), .QN(n1027)
         );
  DFFX1_HVT \keys_reg[9][98]  ( .D(n4154), .CLK(clk), .Q(n2612), .QN(n640) );
  DFFX1_HVT \keys_reg[8][98]  ( .D(n4153), .CLK(clk), .Q(n2611), .QN(n1411) );
  DFFX1_HVT \keys_reg[6][98]  ( .D(n4152), .CLK(clk), .Q(n2610), .QN(n639) );
  DFFX1_HVT \keys_reg[5][98]  ( .D(n4151), .CLK(clk), .Q(n2609), .QN(n1410) );
  DFFX1_HVT \keys_reg[4][98]  ( .D(n4150), .CLK(clk), .Q(n2608), .QN(n383) );
  DFFX1_HVT \keys_reg[3][98]  ( .D(n4149), .CLK(clk), .Q(n2607), .QN(n1409) );
  DFFX1_HVT \keys_reg[1][98]  ( .D(n4148), .CLK(clk), .Q(n2606), .QN(n384) );
  DFFX1_HVT \prev_key_reg[98]  ( .D(n5099), .CLK(clk), .Q(prev_key[98]) );
  DFFX1_HVT \keys_reg[10][99]  ( .D(n4147), .CLK(clk), .Q(n2605), .QN(n900) );
  DFFX1_HVT \keys_reg[9][99]  ( .D(n4146), .CLK(clk), .Q(n2604), .QN(n386) );
  DFFX1_HVT \keys_reg[8][99]  ( .D(n4145), .CLK(clk), .Q(n2603), .QN(n1030) );
  DFFX1_HVT \keys_reg[6][99]  ( .D(n4144), .CLK(clk), .Q(n2602), .QN(n130) );
  DFFX1_HVT \keys_reg[5][99]  ( .D(n4143), .CLK(clk), .Q(n2601), .QN(n1029) );
  DFFX1_HVT \keys_reg[4][99]  ( .D(n4142), .CLK(clk), .Q(n2600), .QN(n128) );
  DFFX1_HVT \keys_reg[3][99]  ( .D(n4141), .CLK(clk), .Q(n2599), .QN(n1028) );
  DFFX1_HVT \keys_reg[1][99]  ( .D(n4140), .CLK(clk), .Q(n2598), .QN(n129) );
  DFFX1_HVT \prev_key_reg[99]  ( .D(n5098), .CLK(clk), .Q(prev_key[99]) );
  DFFX1_HVT \keys_reg[10][100]  ( .D(n4139), .CLK(clk), .Q(n2597), .QN(n901)
         );
  DFFX1_HVT \keys_reg[9][100]  ( .D(n4138), .CLK(clk), .Q(n2596), .QN(n388) );
  DFFX1_HVT \keys_reg[8][100]  ( .D(n4137), .CLK(clk), .Q(n2595), .QN(n1033)
         );
  DFFX1_HVT \keys_reg[6][100]  ( .D(n4136), .CLK(clk), .Q(n2594), .QN(n387) );
  DFFX1_HVT \keys_reg[5][100]  ( .D(n4135), .CLK(clk), .Q(n2593), .QN(n1032)
         );
  DFFX1_HVT \keys_reg[4][100]  ( .D(n4134), .CLK(clk), .Q(n2592), .QN(n131) );
  DFFX1_HVT \keys_reg[3][100]  ( .D(n4133), .CLK(clk), .Q(n2591), .QN(n1031)
         );
  DFFX1_HVT \keys_reg[1][100]  ( .D(n4132), .CLK(clk), .Q(n2590), .QN(n132) );
  DFFX1_HVT \prev_key_reg[100]  ( .D(n5097), .CLK(clk), .Q(prev_key[100]) );
  DFFX1_HVT \keys_reg[10][101]  ( .D(n4131), .CLK(clk), .Q(n2589), .QN(n902)
         );
  DFFX1_HVT \keys_reg[9][101]  ( .D(n4130), .CLK(clk), .Q(n2588), .QN(n390) );
  DFFX1_HVT \keys_reg[8][101]  ( .D(n4129), .CLK(clk), .Q(n2587), .QN(n1036)
         );
  DFFX1_HVT \keys_reg[6][101]  ( .D(n4128), .CLK(clk), .Q(n2586), .QN(n389) );
  DFFX1_HVT \keys_reg[5][101]  ( .D(n4127), .CLK(clk), .Q(n2585), .QN(n1035)
         );
  DFFX1_HVT \keys_reg[4][101]  ( .D(n4126), .CLK(clk), .Q(n2584), .QN(n133) );
  DFFX1_HVT \keys_reg[3][101]  ( .D(n4125), .CLK(clk), .Q(n2583), .QN(n1034)
         );
  DFFX1_HVT \keys_reg[1][101]  ( .D(n4124), .CLK(clk), .Q(n2582), .QN(n134) );
  DFFX1_HVT \prev_key_reg[101]  ( .D(n5096), .CLK(clk), .Q(prev_key[101]) );
  DFFX1_HVT \keys_reg[10][102]  ( .D(n4123), .CLK(clk), .Q(n2581), .QN(n903)
         );
  DFFX1_HVT \keys_reg[9][102]  ( .D(n4122), .CLK(clk), .Q(n2580), .QN(n392) );
  DFFX1_HVT \keys_reg[8][102]  ( .D(n4121), .CLK(clk), .Q(n2579), .QN(n1039)
         );
  DFFX1_HVT \keys_reg[6][102]  ( .D(n4120), .CLK(clk), .Q(n2578), .QN(n391) );
  DFFX1_HVT \keys_reg[5][102]  ( .D(n4119), .CLK(clk), .Q(n2577), .QN(n1038)
         );
  DFFX1_HVT \keys_reg[4][102]  ( .D(n4118), .CLK(clk), .Q(n2576), .QN(n135) );
  DFFX1_HVT \keys_reg[3][102]  ( .D(n4117), .CLK(clk), .Q(n2575), .QN(n1037)
         );
  DFFX1_HVT \keys_reg[1][102]  ( .D(n4116), .CLK(clk), .Q(n2574), .QN(n136) );
  DFFX1_HVT \prev_key_reg[102]  ( .D(n5095), .CLK(clk), .Q(prev_key[102]) );
  DFFX1_HVT \keys_reg[10][103]  ( .D(n4115), .CLK(clk), .Q(n2573), .QN(n904)
         );
  DFFX1_HVT \keys_reg[9][103]  ( .D(n4114), .CLK(clk), .Q(n2572), .QN(n394) );
  DFFX1_HVT \keys_reg[8][103]  ( .D(n4113), .CLK(clk), .Q(n2571), .QN(n1042)
         );
  DFFX1_HVT \keys_reg[6][103]  ( .D(n4112), .CLK(clk), .Q(n2570), .QN(n393) );
  DFFX1_HVT \keys_reg[5][103]  ( .D(n4111), .CLK(clk), .Q(n2569), .QN(n1041)
         );
  DFFX1_HVT \keys_reg[4][103]  ( .D(n4110), .CLK(clk), .Q(n2568), .QN(n137) );
  DFFX1_HVT \keys_reg[3][103]  ( .D(n4109), .CLK(clk), .Q(n2567), .QN(n1040)
         );
  DFFX1_HVT \keys_reg[1][103]  ( .D(n4108), .CLK(clk), .Q(n2566), .QN(n138) );
  DFFX1_HVT \prev_key_reg[103]  ( .D(n5094), .CLK(clk), .Q(prev_key[103]) );
  DFFX1_HVT \keys_reg[10][104]  ( .D(n4107), .CLK(clk), .Q(n2565), .QN(n905)
         );
  DFFX1_HVT \keys_reg[9][104]  ( .D(n4106), .CLK(clk), .Q(n2564), .QN(n396) );
  DFFX1_HVT \keys_reg[8][104]  ( .D(n4105), .CLK(clk), .Q(n2563), .QN(n1045)
         );
  DFFX1_HVT \keys_reg[6][104]  ( .D(n4104), .CLK(clk), .Q(n2562), .QN(n395) );
  DFFX1_HVT \keys_reg[5][104]  ( .D(n4103), .CLK(clk), .Q(n2561), .QN(n1044)
         );
  DFFX1_HVT \keys_reg[4][104]  ( .D(n4102), .CLK(clk), .Q(n2560), .QN(n139) );
  DFFX1_HVT \keys_reg[3][104]  ( .D(n4101), .CLK(clk), .Q(n2559), .QN(n1043)
         );
  DFFX1_HVT \keys_reg[1][104]  ( .D(n4100), .CLK(clk), .Q(n2558), .QN(n140) );
  DFFX1_HVT \prev_key_reg[104]  ( .D(n5093), .CLK(clk), .Q(prev_key[104]) );
  DFFX1_HVT \keys_reg[10][105]  ( .D(n4099), .CLK(clk), .Q(n2557), .QN(n906)
         );
  DFFX1_HVT \keys_reg[9][105]  ( .D(n4098), .CLK(clk), .Q(n2556), .QN(n398) );
  DFFX1_HVT \keys_reg[8][105]  ( .D(n4097), .CLK(clk), .Q(n2555), .QN(n1048)
         );
  DFFX1_HVT \keys_reg[6][105]  ( .D(n4096), .CLK(clk), .Q(n2554), .QN(n397) );
  DFFX1_HVT \keys_reg[5][105]  ( .D(n4095), .CLK(clk), .Q(n2553), .QN(n1047)
         );
  DFFX1_HVT \keys_reg[4][105]  ( .D(n4094), .CLK(clk), .Q(n2552), .QN(n141) );
  DFFX1_HVT \keys_reg[3][105]  ( .D(n4093), .CLK(clk), .Q(n2551), .QN(n1046)
         );
  DFFX1_HVT \keys_reg[1][105]  ( .D(n4092), .CLK(clk), .Q(n2550), .QN(n142) );
  DFFX1_HVT \prev_key_reg[105]  ( .D(n5092), .CLK(clk), .Q(prev_key[105]) );
  DFFX1_HVT \keys_reg[10][106]  ( .D(n4091), .CLK(clk), .Q(n2549), .QN(n907)
         );
  DFFX1_HVT \keys_reg[9][106]  ( .D(n4090), .CLK(clk), .Q(n2548), .QN(n400) );
  DFFX1_HVT \keys_reg[8][106]  ( .D(n4089), .CLK(clk), .Q(n2547), .QN(n1051)
         );
  DFFX1_HVT \keys_reg[6][106]  ( .D(n4088), .CLK(clk), .Q(n2546), .QN(n399) );
  DFFX1_HVT \keys_reg[5][106]  ( .D(n4087), .CLK(clk), .Q(n2545), .QN(n1050)
         );
  DFFX1_HVT \keys_reg[4][106]  ( .D(n4086), .CLK(clk), .Q(n2544), .QN(n143) );
  DFFX1_HVT \keys_reg[3][106]  ( .D(n4085), .CLK(clk), .Q(n2543), .QN(n1049)
         );
  DFFX1_HVT \keys_reg[1][106]  ( .D(n4084), .CLK(clk), .Q(n2542), .QN(n144) );
  DFFX1_HVT \prev_key_reg[106]  ( .D(n5091), .CLK(clk), .Q(prev_key[106]) );
  DFFX1_HVT \keys_reg[10][107]  ( .D(n4083), .CLK(clk), .Q(n2541), .QN(n908)
         );
  DFFX1_HVT \keys_reg[9][107]  ( .D(n4082), .CLK(clk), .Q(n2540), .QN(n402) );
  DFFX1_HVT \keys_reg[8][107]  ( .D(n4081), .CLK(clk), .Q(n2539), .QN(n1054)
         );
  DFFX1_HVT \keys_reg[6][107]  ( .D(n4080), .CLK(clk), .Q(n2538), .QN(n401) );
  DFFX1_HVT \keys_reg[5][107]  ( .D(n4079), .CLK(clk), .Q(n2537), .QN(n1053)
         );
  DFFX1_HVT \keys_reg[4][107]  ( .D(n4078), .CLK(clk), .Q(n2536), .QN(n145) );
  DFFX1_HVT \keys_reg[3][107]  ( .D(n4077), .CLK(clk), .Q(n2535), .QN(n1052)
         );
  DFFX1_HVT \keys_reg[1][107]  ( .D(n4076), .CLK(clk), .Q(n2534), .QN(n146) );
  DFFX1_HVT \prev_key_reg[107]  ( .D(n5090), .CLK(clk), .Q(prev_key[107]) );
  DFFX1_HVT \keys_reg[10][108]  ( .D(n4075), .CLK(clk), .Q(n2533), .QN(n909)
         );
  DFFX1_HVT \keys_reg[9][108]  ( .D(n4074), .CLK(clk), .Q(n2532), .QN(n404) );
  DFFX1_HVT \keys_reg[8][108]  ( .D(n4073), .CLK(clk), .Q(n2531), .QN(n1057)
         );
  DFFX1_HVT \keys_reg[6][108]  ( .D(n4072), .CLK(clk), .Q(n2530), .QN(n403) );
  DFFX1_HVT \keys_reg[5][108]  ( .D(n4071), .CLK(clk), .Q(n2529), .QN(n1056)
         );
  DFFX1_HVT \keys_reg[4][108]  ( .D(n4070), .CLK(clk), .Q(n2528), .QN(n147) );
  DFFX1_HVT \keys_reg[3][108]  ( .D(n4069), .CLK(clk), .Q(n2527), .QN(n1055)
         );
  DFFX1_HVT \keys_reg[1][108]  ( .D(n4068), .CLK(clk), .Q(n2526), .QN(n148) );
  DFFX1_HVT \prev_key_reg[108]  ( .D(n5089), .CLK(clk), .Q(prev_key[108]) );
  DFFX1_HVT \keys_reg[10][109]  ( .D(n4067), .CLK(clk), .Q(n2525), .QN(n910)
         );
  DFFX1_HVT \keys_reg[9][109]  ( .D(n4066), .CLK(clk), .Q(n2524), .QN(n406) );
  DFFX1_HVT \keys_reg[8][109]  ( .D(n4065), .CLK(clk), .Q(n2523), .QN(n1060)
         );
  DFFX1_HVT \keys_reg[6][109]  ( .D(n4064), .CLK(clk), .Q(n2522), .QN(n405) );
  DFFX1_HVT \keys_reg[5][109]  ( .D(n4063), .CLK(clk), .Q(n2521), .QN(n1059)
         );
  DFFX1_HVT \keys_reg[4][109]  ( .D(n4062), .CLK(clk), .Q(n2520), .QN(n149) );
  DFFX1_HVT \keys_reg[3][109]  ( .D(n4061), .CLK(clk), .Q(n2519), .QN(n1058)
         );
  DFFX1_HVT \keys_reg[1][109]  ( .D(n4060), .CLK(clk), .Q(n2518), .QN(n150) );
  DFFX1_HVT \prev_key_reg[109]  ( .D(n5088), .CLK(clk), .Q(prev_key[109]) );
  DFFX1_HVT \keys_reg[10][110]  ( .D(n4059), .CLK(clk), .Q(n2517), .QN(n911)
         );
  DFFX1_HVT \keys_reg[9][110]  ( .D(n4058), .CLK(clk), .Q(n2516), .QN(n408) );
  DFFX1_HVT \keys_reg[8][110]  ( .D(n4057), .CLK(clk), .Q(n2515), .QN(n1063)
         );
  DFFX1_HVT \keys_reg[6][110]  ( .D(n4056), .CLK(clk), .Q(n2514), .QN(n407) );
  DFFX1_HVT \keys_reg[5][110]  ( .D(n4055), .CLK(clk), .Q(n2513), .QN(n1062)
         );
  DFFX1_HVT \keys_reg[4][110]  ( .D(n4054), .CLK(clk), .Q(n2512), .QN(n151) );
  DFFX1_HVT \keys_reg[3][110]  ( .D(n4053), .CLK(clk), .Q(n2511), .QN(n1061)
         );
  DFFX1_HVT \keys_reg[1][110]  ( .D(n4052), .CLK(clk), .Q(n2510), .QN(n152) );
  DFFX1_HVT \prev_key_reg[110]  ( .D(n5087), .CLK(clk), .Q(prev_key[110]) );
  DFFX1_HVT \keys_reg[10][111]  ( .D(n4051), .CLK(clk), .Q(n2509), .QN(n912)
         );
  DFFX1_HVT \keys_reg[9][111]  ( .D(n4050), .CLK(clk), .Q(n2508), .QN(n410) );
  DFFX1_HVT \keys_reg[8][111]  ( .D(n4049), .CLK(clk), .Q(n2507), .QN(n1066)
         );
  DFFX1_HVT \keys_reg[6][111]  ( .D(n4048), .CLK(clk), .Q(n2506), .QN(n409) );
  DFFX1_HVT \keys_reg[5][111]  ( .D(n4047), .CLK(clk), .Q(n2505), .QN(n1065)
         );
  DFFX1_HVT \keys_reg[4][111]  ( .D(n4046), .CLK(clk), .Q(n2504), .QN(n153) );
  DFFX1_HVT \keys_reg[3][111]  ( .D(n4045), .CLK(clk), .Q(n2503), .QN(n1064)
         );
  DFFX1_HVT \keys_reg[1][111]  ( .D(n4044), .CLK(clk), .Q(n2502), .QN(n154) );
  DFFX1_HVT \prev_key_reg[111]  ( .D(n5086), .CLK(clk), .Q(prev_key[111]) );
  DFFX1_HVT \keys_reg[10][112]  ( .D(n4043), .CLK(clk), .Q(n2501), .QN(n913)
         );
  DFFX1_HVT \keys_reg[9][112]  ( .D(n4042), .CLK(clk), .Q(n2500), .QN(n412) );
  DFFX1_HVT \keys_reg[8][112]  ( .D(n4041), .CLK(clk), .Q(n2499), .QN(n1069)
         );
  DFFX1_HVT \keys_reg[6][112]  ( .D(n4040), .CLK(clk), .Q(n2498), .QN(n411) );
  DFFX1_HVT \keys_reg[5][112]  ( .D(n4039), .CLK(clk), .Q(n2497), .QN(n1068)
         );
  DFFX1_HVT \keys_reg[4][112]  ( .D(n4038), .CLK(clk), .Q(n2496), .QN(n155) );
  DFFX1_HVT \keys_reg[3][112]  ( .D(n4037), .CLK(clk), .Q(n2495), .QN(n1067)
         );
  DFFX1_HVT \keys_reg[1][112]  ( .D(n4036), .CLK(clk), .Q(n2494), .QN(n156) );
  DFFX1_HVT \prev_key_reg[112]  ( .D(n5085), .CLK(clk), .Q(prev_key[112]) );
  DFFX1_HVT \keys_reg[10][113]  ( .D(n4035), .CLK(clk), .Q(n2493), .QN(n914)
         );
  DFFX1_HVT \keys_reg[9][113]  ( .D(n4034), .CLK(clk), .Q(n2492), .QN(n414) );
  DFFX1_HVT \keys_reg[8][113]  ( .D(n4033), .CLK(clk), .Q(n2491), .QN(n1072)
         );
  DFFX1_HVT \keys_reg[6][113]  ( .D(n4032), .CLK(clk), .Q(n2490), .QN(n413) );
  DFFX1_HVT \keys_reg[5][113]  ( .D(n4031), .CLK(clk), .Q(n2489), .QN(n1071)
         );
  DFFX1_HVT \keys_reg[4][113]  ( .D(n4030), .CLK(clk), .Q(n2488), .QN(n157) );
  DFFX1_HVT \keys_reg[3][113]  ( .D(n4029), .CLK(clk), .Q(n2487), .QN(n1070)
         );
  DFFX1_HVT \keys_reg[1][113]  ( .D(n4028), .CLK(clk), .Q(n2486), .QN(n158) );
  DFFX1_HVT \prev_key_reg[113]  ( .D(n5084), .CLK(clk), .Q(prev_key[113]) );
  DFFX1_HVT \keys_reg[10][114]  ( .D(n4027), .CLK(clk), .Q(n2485), .QN(n915)
         );
  DFFX1_HVT \keys_reg[9][114]  ( .D(n4026), .CLK(clk), .Q(n2484), .QN(n416) );
  DFFX1_HVT \keys_reg[8][114]  ( .D(n4025), .CLK(clk), .Q(n2483), .QN(n1075)
         );
  DFFX1_HVT \keys_reg[6][114]  ( .D(n4024), .CLK(clk), .Q(n2482), .QN(n415) );
  DFFX1_HVT \keys_reg[5][114]  ( .D(n4023), .CLK(clk), .Q(n2481), .QN(n1074)
         );
  DFFX1_HVT \keys_reg[4][114]  ( .D(n4022), .CLK(clk), .Q(n2480), .QN(n159) );
  DFFX1_HVT \keys_reg[3][114]  ( .D(n4021), .CLK(clk), .Q(n2479), .QN(n1073)
         );
  DFFX1_HVT \keys_reg[1][114]  ( .D(n4020), .CLK(clk), .Q(n2478), .QN(n160) );
  DFFX1_HVT \prev_key_reg[114]  ( .D(n5083), .CLK(clk), .Q(prev_key[114]) );
  DFFX1_HVT \keys_reg[10][115]  ( .D(n4019), .CLK(clk), .Q(n2477), .QN(n916)
         );
  DFFX1_HVT \keys_reg[9][115]  ( .D(n4018), .CLK(clk), .Q(n2476), .QN(n418) );
  DFFX1_HVT \keys_reg[8][115]  ( .D(n4017), .CLK(clk), .Q(n2475), .QN(n1078)
         );
  DFFX1_HVT \keys_reg[6][115]  ( .D(n4016), .CLK(clk), .Q(n2474), .QN(n417) );
  DFFX1_HVT \keys_reg[5][115]  ( .D(n4015), .CLK(clk), .Q(n2473), .QN(n1077)
         );
  DFFX1_HVT \keys_reg[4][115]  ( .D(n4014), .CLK(clk), .Q(n2472), .QN(n161) );
  DFFX1_HVT \keys_reg[3][115]  ( .D(n4013), .CLK(clk), .Q(n2471), .QN(n1076)
         );
  DFFX1_HVT \keys_reg[1][115]  ( .D(n4012), .CLK(clk), .Q(n2470), .QN(n162) );
  DFFX1_HVT \prev_key_reg[115]  ( .D(n5082), .CLK(clk), .Q(prev_key[115]) );
  DFFX1_HVT \keys_reg[10][116]  ( .D(n4011), .CLK(clk), .Q(n2469), .QN(n917)
         );
  DFFX1_HVT \keys_reg[9][116]  ( .D(n4010), .CLK(clk), .Q(n2468), .QN(n420) );
  DFFX1_HVT \keys_reg[8][116]  ( .D(n4009), .CLK(clk), .Q(n2467), .QN(n1081)
         );
  DFFX1_HVT \keys_reg[6][116]  ( .D(n4008), .CLK(clk), .Q(n2466), .QN(n419) );
  DFFX1_HVT \keys_reg[5][116]  ( .D(n4007), .CLK(clk), .Q(n2465), .QN(n1080)
         );
  DFFX1_HVT \keys_reg[4][116]  ( .D(n4006), .CLK(clk), .Q(n2464), .QN(n163) );
  DFFX1_HVT \keys_reg[3][116]  ( .D(n4005), .CLK(clk), .Q(n2463), .QN(n1079)
         );
  DFFX1_HVT \keys_reg[1][116]  ( .D(n4004), .CLK(clk), .Q(n2462), .QN(n164) );
  DFFX1_HVT \prev_key_reg[116]  ( .D(n5081), .CLK(clk), .Q(prev_key[116]) );
  DFFX1_HVT \keys_reg[10][117]  ( .D(n4003), .CLK(clk), .Q(n2461), .QN(n918)
         );
  DFFX1_HVT \keys_reg[9][117]  ( .D(n4002), .CLK(clk), .Q(n2460), .QN(n422) );
  DFFX1_HVT \keys_reg[8][117]  ( .D(n4001), .CLK(clk), .Q(n2459), .QN(n1084)
         );
  DFFX1_HVT \keys_reg[6][117]  ( .D(n4000), .CLK(clk), .Q(n2458), .QN(n421) );
  DFFX1_HVT \keys_reg[5][117]  ( .D(n3999), .CLK(clk), .Q(n2457), .QN(n1083)
         );
  DFFX1_HVT \keys_reg[4][117]  ( .D(n3998), .CLK(clk), .Q(n2456), .QN(n165) );
  DFFX1_HVT \keys_reg[3][117]  ( .D(n3997), .CLK(clk), .Q(n2455), .QN(n1082)
         );
  DFFX1_HVT \keys_reg[1][117]  ( .D(n3996), .CLK(clk), .Q(n2454), .QN(n166) );
  DFFX1_HVT \prev_key_reg[117]  ( .D(n5080), .CLK(clk), .Q(prev_key[117]) );
  DFFX1_HVT \keys_reg[10][118]  ( .D(n3995), .CLK(clk), .Q(n2453), .QN(n919)
         );
  DFFX1_HVT \keys_reg[9][118]  ( .D(n3994), .CLK(clk), .Q(n2452), .QN(n424) );
  DFFX1_HVT \keys_reg[8][118]  ( .D(n3993), .CLK(clk), .Q(n2451), .QN(n1087)
         );
  DFFX1_HVT \keys_reg[6][118]  ( .D(n3992), .CLK(clk), .Q(n2450), .QN(n423) );
  DFFX1_HVT \keys_reg[5][118]  ( .D(n3991), .CLK(clk), .Q(n2449), .QN(n1086)
         );
  DFFX1_HVT \keys_reg[4][118]  ( .D(n3990), .CLK(clk), .Q(n2448), .QN(n167) );
  DFFX1_HVT \keys_reg[3][118]  ( .D(n3989), .CLK(clk), .Q(n2447), .QN(n1085)
         );
  DFFX1_HVT \keys_reg[1][118]  ( .D(n3988), .CLK(clk), .Q(n2446), .QN(n168) );
  DFFX1_HVT \prev_key_reg[118]  ( .D(n5079), .CLK(clk), .Q(prev_key[118]) );
  DFFX1_HVT \keys_reg[10][119]  ( .D(n3987), .CLK(clk), .Q(n2445), .QN(n920)
         );
  DFFX1_HVT \keys_reg[9][119]  ( .D(n3986), .CLK(clk), .Q(n2444), .QN(n426) );
  DFFX1_HVT \keys_reg[8][119]  ( .D(n3985), .CLK(clk), .Q(n2443), .QN(n1090)
         );
  DFFX1_HVT \keys_reg[6][119]  ( .D(n3984), .CLK(clk), .Q(n2442), .QN(n425) );
  DFFX1_HVT \keys_reg[5][119]  ( .D(n3983), .CLK(clk), .Q(n2441), .QN(n1089)
         );
  DFFX1_HVT \keys_reg[4][119]  ( .D(n3982), .CLK(clk), .Q(n2440), .QN(n169) );
  DFFX1_HVT \keys_reg[3][119]  ( .D(n3981), .CLK(clk), .Q(n2439), .QN(n1088)
         );
  DFFX1_HVT \keys_reg[1][119]  ( .D(n3980), .CLK(clk), .Q(n2438), .QN(n170) );
  DFFX1_HVT \prev_key_reg[119]  ( .D(n5078), .CLK(clk), .Q(prev_key[119]) );
  DFFX1_HVT \keys_reg[10][120]  ( .D(n3979), .CLK(clk), .Q(n2437), .QN(n921)
         );
  DFFX1_HVT \keys_reg[9][120]  ( .D(n3978), .CLK(clk), .Q(n2436), .QN(n428) );
  DFFX1_HVT \keys_reg[8][120]  ( .D(n3977), .CLK(clk), .Q(n2435), .QN(n1093)
         );
  DFFX1_HVT \keys_reg[6][120]  ( .D(n3976), .CLK(clk), .Q(n2434), .QN(n427) );
  DFFX1_HVT \keys_reg[5][120]  ( .D(n3975), .CLK(clk), .Q(n2433), .QN(n1092)
         );
  DFFX1_HVT \keys_reg[4][120]  ( .D(n3974), .CLK(clk), .Q(n2432), .QN(n171) );
  DFFX1_HVT \keys_reg[3][120]  ( .D(n3973), .CLK(clk), .Q(n2431), .QN(n1091)
         );
  DFFX1_HVT \keys_reg[1][120]  ( .D(n3972), .CLK(clk), .Q(n2430), .QN(n172) );
  DFFX1_HVT \prev_key_reg[120]  ( .D(n5077), .CLK(clk), .Q(prev_key[120]) );
  DFFX1_HVT \keys_reg[10][121]  ( .D(n3971), .CLK(clk), .Q(n2429), .QN(n922)
         );
  DFFX1_HVT \keys_reg[9][121]  ( .D(n3970), .CLK(clk), .Q(n2428), .QN(n430) );
  DFFX1_HVT \keys_reg[8][121]  ( .D(n3969), .CLK(clk), .Q(n2427), .QN(n1096)
         );
  DFFX1_HVT \keys_reg[6][121]  ( .D(n3968), .CLK(clk), .Q(n2426), .QN(n429) );
  DFFX1_HVT \keys_reg[5][121]  ( .D(n3967), .CLK(clk), .Q(n2425), .QN(n1095)
         );
  DFFX1_HVT \keys_reg[4][121]  ( .D(n3966), .CLK(clk), .Q(n2424), .QN(n173) );
  DFFX1_HVT \keys_reg[3][121]  ( .D(n3965), .CLK(clk), .Q(n2423), .QN(n1094)
         );
  DFFX1_HVT \keys_reg[1][121]  ( .D(n3964), .CLK(clk), .Q(n2422), .QN(n174) );
  DFFX1_HVT \prev_key_reg[121]  ( .D(n5076), .CLK(clk), .Q(prev_key[121]) );
  DFFX1_HVT \keys_reg[10][122]  ( .D(n3963), .CLK(clk), .Q(n2421), .QN(n923)
         );
  DFFX1_HVT \keys_reg[9][122]  ( .D(n3962), .CLK(clk), .Q(n2420), .QN(n432) );
  DFFX1_HVT \keys_reg[8][122]  ( .D(n3961), .CLK(clk), .Q(n2419), .QN(n1099)
         );
  DFFX1_HVT \keys_reg[6][122]  ( .D(n3960), .CLK(clk), .Q(n2418), .QN(n431) );
  DFFX1_HVT \keys_reg[5][122]  ( .D(n3959), .CLK(clk), .Q(n2417), .QN(n1098)
         );
  DFFX1_HVT \keys_reg[4][122]  ( .D(n3958), .CLK(clk), .Q(n2416), .QN(n175) );
  DFFX1_HVT \keys_reg[3][122]  ( .D(n3957), .CLK(clk), .Q(n2415), .QN(n1097)
         );
  DFFX1_HVT \keys_reg[1][122]  ( .D(n3956), .CLK(clk), .Q(n2414), .QN(n176) );
  DFFX1_HVT \prev_key_reg[122]  ( .D(n5075), .CLK(clk), .Q(prev_key[122]) );
  DFFX1_HVT \keys_reg[10][123]  ( .D(n3955), .CLK(clk), .Q(n2413), .QN(n924)
         );
  DFFX1_HVT \keys_reg[9][123]  ( .D(n3954), .CLK(clk), .Q(n2412), .QN(n434) );
  DFFX1_HVT \keys_reg[8][123]  ( .D(n3953), .CLK(clk), .Q(n2411), .QN(n1102)
         );
  DFFX1_HVT \keys_reg[6][123]  ( .D(n3952), .CLK(clk), .Q(n2410), .QN(n433) );
  DFFX1_HVT \keys_reg[5][123]  ( .D(n3951), .CLK(clk), .Q(n2409), .QN(n1101)
         );
  DFFX1_HVT \keys_reg[4][123]  ( .D(n3950), .CLK(clk), .Q(n2408), .QN(n177) );
  DFFX1_HVT \keys_reg[3][123]  ( .D(n3949), .CLK(clk), .Q(n2407), .QN(n1100)
         );
  DFFX1_HVT \keys_reg[1][123]  ( .D(n3948), .CLK(clk), .Q(n2406), .QN(n178) );
  DFFX1_HVT \prev_key_reg[123]  ( .D(n5074), .CLK(clk), .Q(prev_key[123]) );
  DFFX1_HVT \keys_reg[10][124]  ( .D(n3947), .CLK(clk), .Q(n2405), .QN(n925)
         );
  DFFX1_HVT \keys_reg[9][124]  ( .D(n3946), .CLK(clk), .Q(n2404), .QN(n436) );
  DFFX1_HVT \keys_reg[8][124]  ( .D(n3945), .CLK(clk), .Q(n2403), .QN(n1105)
         );
  DFFX1_HVT \keys_reg[6][124]  ( .D(n3944), .CLK(clk), .Q(n2402), .QN(n435) );
  DFFX1_HVT \keys_reg[5][124]  ( .D(n3943), .CLK(clk), .Q(n2401), .QN(n1104)
         );
  DFFX1_HVT \keys_reg[4][124]  ( .D(n3942), .CLK(clk), .Q(n2400), .QN(n179) );
  DFFX1_HVT \keys_reg[3][124]  ( .D(n3941), .CLK(clk), .Q(n2399), .QN(n1103)
         );
  DFFX1_HVT \keys_reg[1][124]  ( .D(n3940), .CLK(clk), .Q(n2398), .QN(n180) );
  DFFX1_HVT \prev_key_reg[124]  ( .D(n5073), .CLK(clk), .Q(prev_key[124]) );
  DFFX1_HVT \keys_reg[10][125]  ( .D(n3939), .CLK(clk), .Q(n2397), .QN(n926)
         );
  DFFX1_HVT \keys_reg[9][125]  ( .D(n3938), .CLK(clk), .Q(n2396), .QN(n438) );
  DFFX1_HVT \keys_reg[8][125]  ( .D(n3937), .CLK(clk), .Q(n2395), .QN(n1108)
         );
  DFFX1_HVT \keys_reg[6][125]  ( .D(n3936), .CLK(clk), .Q(n2394), .QN(n437) );
  DFFX1_HVT \keys_reg[5][125]  ( .D(n3935), .CLK(clk), .Q(n2393), .QN(n1107)
         );
  DFFX1_HVT \keys_reg[4][125]  ( .D(n3934), .CLK(clk), .Q(n2392), .QN(n181) );
  DFFX1_HVT \keys_reg[3][125]  ( .D(n3933), .CLK(clk), .Q(n2391), .QN(n1106)
         );
  DFFX1_HVT \keys_reg[1][125]  ( .D(n3932), .CLK(clk), .Q(n2390), .QN(n182) );
  DFFX1_HVT \prev_key_reg[125]  ( .D(n5072), .CLK(clk), .Q(prev_key[125]) );
  DFFX1_HVT \keys_reg[10][126]  ( .D(n3931), .CLK(clk), .Q(n2389), .QN(n927)
         );
  DFFX1_HVT \keys_reg[9][126]  ( .D(n3930), .CLK(clk), .Q(n2388), .QN(n440) );
  DFFX1_HVT \keys_reg[8][126]  ( .D(n3929), .CLK(clk), .Q(n2387), .QN(n1111)
         );
  DFFX1_HVT \keys_reg[6][126]  ( .D(n3928), .CLK(clk), .Q(n2386), .QN(n439) );
  DFFX1_HVT \keys_reg[5][126]  ( .D(n3927), .CLK(clk), .Q(n2385), .QN(n1110)
         );
  DFFX1_HVT \keys_reg[4][126]  ( .D(n3926), .CLK(clk), .Q(n2384), .QN(n183) );
  DFFX1_HVT \keys_reg[3][126]  ( .D(n3925), .CLK(clk), .Q(n2383), .QN(n1109)
         );
  DFFX1_HVT \keys_reg[1][126]  ( .D(n3924), .CLK(clk), .Q(n2382), .QN(n184) );
  DFFX1_HVT \prev_key_reg[126]  ( .D(n5071), .CLK(clk), .Q(prev_key[126]) );
  DFFX1_HVT \keys_reg[10][127]  ( .D(n3923), .CLK(clk), .Q(n2381), .QN(n928)
         );
  DFFX1_HVT \keys_reg[9][127]  ( .D(n3922), .CLK(clk), .Q(n2380), .QN(n442) );
  DFFX1_HVT \keys_reg[8][127]  ( .D(n3921), .CLK(clk), .Q(n2379), .QN(n1114)
         );
  DFFX1_HVT \keys_reg[6][127]  ( .D(n3920), .CLK(clk), .Q(n2378), .QN(n441) );
  DFFX1_HVT \keys_reg[5][127]  ( .D(n3919), .CLK(clk), .Q(n2377), .QN(n1113)
         );
  DFFX1_HVT \keys_reg[4][127]  ( .D(n3918), .CLK(clk), .Q(n2376), .QN(n185) );
  DFFX1_HVT \keys_reg[3][127]  ( .D(n3917), .CLK(clk), .Q(n2375), .QN(n1112)
         );
  DFFX1_HVT \keys_reg[1][127]  ( .D(n3916), .CLK(clk), .Q(n2374), .QN(n186) );
  DFFX1_HVT \prev_key_reg[127]  ( .D(n5070), .CLK(clk), .Q(prev_key[127]) );
  DFFX1_HVT \keys_reg[2][99]  ( .D(n3915), .CLK(clk), .Q(n2373), .QN(n641) );
  DFFX1_HVT \keys_reg[2][100]  ( .D(n3914), .CLK(clk), .Q(n2372), .QN(n644) );
  DFFX1_HVT \keys_reg[2][101]  ( .D(n3913), .CLK(clk), .Q(n2371), .QN(n646) );
  DFFX1_HVT \keys_reg[2][102]  ( .D(n3912), .CLK(clk), .Q(n2370), .QN(n648) );
  DFFX1_HVT \keys_reg[2][103]  ( .D(n3911), .CLK(clk), .Q(n2369), .QN(n650) );
  DFFX1_HVT \keys_reg[2][104]  ( .D(n3910), .CLK(clk), .Q(n2368), .QN(n652) );
  DFFX1_HVT \keys_reg[2][105]  ( .D(n3909), .CLK(clk), .Q(n2367), .QN(n654) );
  DFFX1_HVT \keys_reg[2][106]  ( .D(n3908), .CLK(clk), .Q(n2366), .QN(n656) );
  DFFX1_HVT \keys_reg[2][107]  ( .D(n3907), .CLK(clk), .Q(n2365), .QN(n658) );
  DFFX1_HVT \keys_reg[2][108]  ( .D(n3906), .CLK(clk), .Q(n2364), .QN(n660) );
  DFFX1_HVT \keys_reg[2][109]  ( .D(n3905), .CLK(clk), .Q(n2363), .QN(n662) );
  DFFX1_HVT \keys_reg[2][110]  ( .D(n3904), .CLK(clk), .Q(n2362), .QN(n664) );
  DFFX1_HVT \keys_reg[2][111]  ( .D(n3903), .CLK(clk), .Q(n2361), .QN(n666) );
  DFFX1_HVT \keys_reg[2][112]  ( .D(n3902), .CLK(clk), .Q(n2360), .QN(n668) );
  DFFX1_HVT \keys_reg[2][113]  ( .D(n3901), .CLK(clk), .Q(n2359), .QN(n670) );
  DFFX1_HVT \keys_reg[2][114]  ( .D(n3900), .CLK(clk), .Q(n2358), .QN(n672) );
  DFFX1_HVT \keys_reg[2][115]  ( .D(n3899), .CLK(clk), .Q(n2357), .QN(n674) );
  DFFX1_HVT \keys_reg[2][116]  ( .D(n3898), .CLK(clk), .Q(n2356), .QN(n676) );
  DFFX1_HVT \keys_reg[2][117]  ( .D(n3897), .CLK(clk), .Q(n2355), .QN(n678) );
  DFFX1_HVT \keys_reg[2][118]  ( .D(n3896), .CLK(clk), .Q(n2354), .QN(n680) );
  DFFX1_HVT \keys_reg[2][119]  ( .D(n3895), .CLK(clk), .Q(n2353), .QN(n682) );
  DFFX1_HVT \keys_reg[2][120]  ( .D(n3894), .CLK(clk), .Q(n2352), .QN(n684) );
  DFFX1_HVT \keys_reg[2][121]  ( .D(n3893), .CLK(clk), .Q(n2351), .QN(n686) );
  DFFX1_HVT \keys_reg[2][122]  ( .D(n3892), .CLK(clk), .Q(n2350), .QN(n688) );
  DFFX1_HVT \keys_reg[2][123]  ( .D(n3891), .CLK(clk), .Q(n2349), .QN(n690) );
  DFFX1_HVT \keys_reg[2][124]  ( .D(n3890), .CLK(clk), .Q(n2348), .QN(n692) );
  DFFX1_HVT \keys_reg[2][125]  ( .D(n3889), .CLK(clk), .Q(n2347), .QN(n694) );
  DFFX1_HVT \keys_reg[2][126]  ( .D(n3888), .CLK(clk), .Q(n2346), .QN(n696) );
  DFFX1_HVT \keys_reg[2][127]  ( .D(n3887), .CLK(clk), .Q(n2345), .QN(n698) );
  DFFX1_HVT \keys_reg[2][49]  ( .D(n3886), .CLK(clk), .Q(n2344), .QN(n894) );
  DFFX1_HVT \keys_reg[2][50]  ( .D(n3885), .CLK(clk), .Q(n2343), .QN(n892) );
  DFFX1_HVT \keys_reg[2][51]  ( .D(n3884), .CLK(clk), .Q(n2342), .QN(n890) );
  DFFX1_HVT \keys_reg[2][52]  ( .D(n3883), .CLK(clk), .Q(n2341), .QN(n888) );
  DFFX1_HVT \keys_reg[2][53]  ( .D(n3882), .CLK(clk), .Q(n2340), .QN(n886) );
  DFFX1_HVT \keys_reg[2][54]  ( .D(n3881), .CLK(clk), .Q(n2339), .QN(n884) );
  DFFX1_HVT \keys_reg[2][55]  ( .D(n3880), .CLK(clk), .Q(n2338), .QN(n882) );
  DFFX1_HVT \keys_reg[2][56]  ( .D(n3879), .CLK(clk), .Q(n2337), .QN(n880) );
  DFFX1_HVT \keys_reg[2][57]  ( .D(n3878), .CLK(clk), .Q(n2336), .QN(n878) );
  DFFX1_HVT \keys_reg[2][58]  ( .D(n3877), .CLK(clk), .Q(n2335), .QN(n876) );
  DFFX1_HVT \keys_reg[2][59]  ( .D(n3876), .CLK(clk), .Q(n2334), .QN(n874) );
  DFFX1_HVT \keys_reg[2][60]  ( .D(n3875), .CLK(clk), .Q(n2333), .QN(n872) );
  DFFX1_HVT \keys_reg[2][61]  ( .D(n3874), .CLK(clk), .Q(n2332), .QN(n870) );
  DFFX1_HVT \keys_reg[2][62]  ( .D(n3873), .CLK(clk), .Q(n2331), .QN(n868) );
  DFFX1_HVT \keys_reg[2][63]  ( .D(n3872), .CLK(clk), .Q(n2330), .QN(n866) );
  DFFX1_HVT \keys_reg[2][64]  ( .D(n3871), .CLK(clk), .Q(n2329), .QN(n864) );
  DFFX1_HVT \keys_reg[2][65]  ( .D(n3870), .CLK(clk), .Q(n2328), .QN(n862) );
  DFFX1_HVT \keys_reg[2][66]  ( .D(n3869), .CLK(clk), .Q(n2327), .QN(n860) );
  DFFX1_HVT \keys_reg[2][67]  ( .D(n3868), .CLK(clk), .Q(n2326), .QN(n858) );
  DFFX1_HVT \keys_reg[2][68]  ( .D(n3867), .CLK(clk), .Q(n2325), .QN(n856) );
  DFFX1_HVT \keys_reg[2][69]  ( .D(n3866), .CLK(clk), .Q(n2324), .QN(n854) );
  DFFX1_HVT \keys_reg[2][70]  ( .D(n3865), .CLK(clk), .Q(n2323), .QN(n852) );
  DFFX1_HVT \keys_reg[2][71]  ( .D(n3864), .CLK(clk), .Q(n2322), .QN(n850) );
  DFFX1_HVT \keys_reg[2][72]  ( .D(n3863), .CLK(clk), .Q(n2321), .QN(n848) );
  DFFX1_HVT \keys_reg[2][73]  ( .D(n3862), .CLK(clk), .Q(n2320), .QN(n846) );
  DFFX1_HVT \keys_reg[2][74]  ( .D(n3861), .CLK(clk), .Q(n2319), .QN(n844) );
  DFFX1_HVT \keys_reg[2][75]  ( .D(n3860), .CLK(clk), .Q(n2318), .QN(n842) );
  DFFX1_HVT \keys_reg[2][76]  ( .D(n3859), .CLK(clk), .Q(n2317), .QN(n840) );
  DFFX1_HVT \keys_reg[2][77]  ( .D(n3858), .CLK(clk), .Q(n2316), .QN(n838) );
  DFFX1_HVT \keys_reg[2][78]  ( .D(n3857), .CLK(clk), .Q(n2315), .QN(n836) );
  DFFX1_HVT \keys_reg[2][79]  ( .D(n3856), .CLK(clk), .Q(n2314), .QN(n834) );
  DFFX1_HVT \keys_reg[2][80]  ( .D(n3855), .CLK(clk), .Q(n2313), .QN(n832) );
  DFFX1_HVT \keys_reg[2][81]  ( .D(n3854), .CLK(clk), .Q(n2312), .QN(n830) );
  DFFX1_HVT \keys_reg[2][82]  ( .D(n3853), .CLK(clk), .Q(n2311), .QN(n700) );
  DFFX1_HVT \keys_reg[2][83]  ( .D(n3852), .CLK(clk), .Q(n2310), .QN(n702) );
  DFFX1_HVT \keys_reg[2][84]  ( .D(n3851), .CLK(clk), .Q(n2309), .QN(n704) );
  DFFX1_HVT \keys_reg[2][85]  ( .D(n3850), .CLK(clk), .Q(n2308), .QN(n706) );
  DFFX1_HVT \keys_reg[2][86]  ( .D(n3849), .CLK(clk), .Q(n2307), .QN(n708) );
  DFFX1_HVT \keys_reg[2][87]  ( .D(n3848), .CLK(clk), .Q(n2306), .QN(n710) );
  DFFX1_HVT \keys_reg[2][88]  ( .D(n3847), .CLK(clk), .Q(n2305), .QN(n712) );
  DFFX1_HVT \keys_reg[2][89]  ( .D(n3846), .CLK(clk), .Q(n2304), .QN(n714) );
  DFFX1_HVT \keys_reg[2][90]  ( .D(n3845), .CLK(clk), .Q(n2303), .QN(n716) );
  DFFX1_HVT \keys_reg[2][91]  ( .D(n3844), .CLK(clk), .Q(n2302), .QN(n718) );
  DFFX1_HVT \keys_reg[2][92]  ( .D(n3843), .CLK(clk), .Q(n2301), .QN(n720) );
  DFFX1_HVT \keys_reg[2][93]  ( .D(n3842), .CLK(clk), .Q(n2300), .QN(n722) );
  DFFX1_HVT \keys_reg[2][94]  ( .D(n3841), .CLK(clk), .Q(n2299), .QN(n724) );
  DFFX1_HVT \keys_reg[2][95]  ( .D(n3840), .CLK(clk), .Q(n2298), .QN(n726) );
  DFFX1_HVT \keys_reg[2][96]  ( .D(n3839), .CLK(clk), .Q(n2297), .QN(n728) );
  DFFX1_HVT \keys_reg[2][97]  ( .D(n3838), .CLK(clk), .Q(n2296), .QN(n730) );
  DFFX1_HVT \keys_reg[2][0]  ( .D(n3837), .CLK(clk), .Q(n2295), .QN(n732) );
  DFFX1_HVT \keys_reg[2][1]  ( .D(n3836), .CLK(clk), .Q(n2294), .QN(n734) );
  DFFX1_HVT \keys_reg[2][2]  ( .D(n3835), .CLK(clk), .Q(n2293), .QN(n736) );
  DFFX1_HVT \keys_reg[2][3]  ( .D(n3834), .CLK(clk), .Q(n2292), .QN(n738) );
  DFFX1_HVT \keys_reg[2][4]  ( .D(n3833), .CLK(clk), .Q(n2291), .QN(n740) );
  DFFX1_HVT \keys_reg[2][5]  ( .D(n3832), .CLK(clk), .Q(n2290), .QN(n742) );
  DFFX1_HVT \keys_reg[2][6]  ( .D(n3831), .CLK(clk), .Q(n2289), .QN(n744) );
  DFFX1_HVT \keys_reg[2][7]  ( .D(n3830), .CLK(clk), .Q(n2288), .QN(n746) );
  DFFX1_HVT \keys_reg[2][8]  ( .D(n3829), .CLK(clk), .Q(n2287), .QN(n748) );
  DFFX1_HVT \keys_reg[2][9]  ( .D(n3828), .CLK(clk), .Q(n2286), .QN(n750) );
  DFFX1_HVT \keys_reg[2][10]  ( .D(n3827), .CLK(clk), .Q(n2285), .QN(n752) );
  DFFX1_HVT \keys_reg[2][11]  ( .D(n3826), .CLK(clk), .Q(n2284), .QN(n754) );
  DFFX1_HVT \keys_reg[2][12]  ( .D(n3825), .CLK(clk), .Q(n2283), .QN(n756) );
  DFFX1_HVT \keys_reg[2][13]  ( .D(n3824), .CLK(clk), .Q(n2282), .QN(n758) );
  DFFX1_HVT \keys_reg[2][14]  ( .D(n3823), .CLK(clk), .Q(n2281), .QN(n760) );
  DFFX1_HVT \keys_reg[2][15]  ( .D(n3822), .CLK(clk), .Q(n2280), .QN(n762) );
  DFFX1_HVT \keys_reg[2][16]  ( .D(n3821), .CLK(clk), .Q(n2279), .QN(n764) );
  DFFX1_HVT \keys_reg[2][17]  ( .D(n3820), .CLK(clk), .Q(n2278), .QN(n766) );
  DFFX1_HVT \keys_reg[2][18]  ( .D(n3819), .CLK(clk), .Q(n2277), .QN(n768) );
  DFFX1_HVT \keys_reg[2][19]  ( .D(n3818), .CLK(clk), .Q(n2276), .QN(n770) );
  DFFX1_HVT \keys_reg[2][20]  ( .D(n3817), .CLK(clk), .Q(n2275), .QN(n772) );
  DFFX1_HVT \keys_reg[2][21]  ( .D(n3816), .CLK(clk), .Q(n2274), .QN(n774) );
  DFFX1_HVT \keys_reg[2][22]  ( .D(n3815), .CLK(clk), .Q(n2273), .QN(n776) );
  DFFX1_HVT \keys_reg[2][23]  ( .D(n3814), .CLK(clk), .Q(n2272), .QN(n778) );
  DFFX1_HVT \keys_reg[2][24]  ( .D(n3813), .CLK(clk), .Q(n2271), .QN(n780) );
  DFFX1_HVT \keys_reg[2][25]  ( .D(n3812), .CLK(clk), .Q(n2270), .QN(n782) );
  DFFX1_HVT \keys_reg[2][26]  ( .D(n3811), .CLK(clk), .Q(n2269), .QN(n784) );
  DFFX1_HVT \keys_reg[2][27]  ( .D(n3810), .CLK(clk), .Q(n2268), .QN(n786) );
  DFFX1_HVT \keys_reg[2][28]  ( .D(n3809), .CLK(clk), .Q(n2267), .QN(n788) );
  DFFX1_HVT \keys_reg[2][29]  ( .D(n3808), .CLK(clk), .Q(n2266), .QN(n790) );
  DFFX1_HVT \keys_reg[2][30]  ( .D(n3807), .CLK(clk), .Q(n2265), .QN(n792) );
  DFFX1_HVT \keys_reg[2][31]  ( .D(n3806), .CLK(clk), .Q(n2264), .QN(n794) );
  DFFX1_HVT \keys_reg[2][32]  ( .D(n3805), .CLK(clk), .Q(n2263), .QN(n796) );
  DFFX1_HVT \keys_reg[2][33]  ( .D(n3804), .CLK(clk), .Q(n2262), .QN(n798) );
  DFFX1_HVT \keys_reg[2][34]  ( .D(n3803), .CLK(clk), .Q(n2261), .QN(n800) );
  DFFX1_HVT \keys_reg[2][35]  ( .D(n3802), .CLK(clk), .Q(n2260), .QN(n802) );
  DFFX1_HVT \keys_reg[2][48]  ( .D(n3801), .CLK(clk), .Q(n2259), .QN(n828) );
  DFFX1_HVT \keys_reg[2][47]  ( .D(n3800), .CLK(clk), .Q(n2258), .QN(n826) );
  DFFX1_HVT \keys_reg[2][46]  ( .D(n3799), .CLK(clk), .Q(n2257), .QN(n824) );
  DFFX1_HVT \keys_reg[2][45]  ( .D(n3798), .CLK(clk), .Q(n2256), .QN(n822) );
  DFFX1_HVT \keys_reg[2][44]  ( .D(n3797), .CLK(clk), .Q(n2255), .QN(n820) );
  DFFX1_HVT \keys_reg[2][43]  ( .D(n3796), .CLK(clk), .Q(n2254), .QN(n818) );
  DFFX1_HVT \keys_reg[2][42]  ( .D(n3795), .CLK(clk), .Q(n2253), .QN(n816) );
  DFFX1_HVT \keys_reg[2][41]  ( .D(n3794), .CLK(clk), .Q(n2252), .QN(n814) );
  DFFX1_HVT \keys_reg[2][40]  ( .D(n3793), .CLK(clk), .Q(n2251), .QN(n812) );
  DFFX1_HVT \keys_reg[2][39]  ( .D(n3792), .CLK(clk), .Q(n2250), .QN(n810) );
  DFFX1_HVT \keys_reg[2][38]  ( .D(n3791), .CLK(clk), .Q(n2249), .QN(n808) );
  DFFX1_HVT \keys_reg[2][37]  ( .D(n3790), .CLK(clk), .Q(n2247), .QN(n806) );
  DFFX1_HVT \keys_reg[2][36]  ( .D(n3789), .CLK(clk), .Q(n2245), .QN(n804) );
  DFFX1_HVT \keys_reg[2][98]  ( .D(n3788), .CLK(clk), .Q(n2243), .QN(n896) );
  DFFX1_HVT \keys_reg[7][99]  ( .D(n3787), .CLK(clk), .Q(n2241), .QN(n643) );
  DFFX1_HVT \key_round_reg[99]  ( .D(n3786), .CLK(clk), .Q(key_round[99]), 
        .QN(n2248) );
  DFFX1_HVT \keys_reg[7][100]  ( .D(n3785), .CLK(clk), .Q(n2239), .QN(n1) );
  DFFX1_HVT \key_round_reg[100]  ( .D(n3784), .CLK(clk), .Q(key_round[100]), 
        .QN(n2246) );
  DFFX1_HVT \keys_reg[7][101]  ( .D(n3783), .CLK(clk), .Q(n2237), .QN(n2) );
  DFFX1_HVT \key_round_reg[101]  ( .D(n3782), .CLK(clk), .Q(key_round[101]), 
        .QN(n2244) );
  DFFX1_HVT \keys_reg[7][102]  ( .D(n3781), .CLK(clk), .Q(n2235), .QN(n3) );
  DFFX1_HVT \key_round_reg[102]  ( .D(n3780), .CLK(clk), .Q(key_round[102]), 
        .QN(n2242) );
  DFFX1_HVT \keys_reg[7][103]  ( .D(n3779), .CLK(clk), .Q(n2233), .QN(n4) );
  DFFX1_HVT \key_round_reg[103]  ( .D(n3778), .CLK(clk), .Q(key_round[103]), 
        .QN(n2240) );
  DFFX1_HVT \keys_reg[7][104]  ( .D(n3777), .CLK(clk), .Q(n2231), .QN(n5) );
  DFFX1_HVT \key_round_reg[104]  ( .D(n3776), .CLK(clk), .Q(key_round[104]), 
        .QN(n2238) );
  DFFX1_HVT \keys_reg[7][105]  ( .D(n3775), .CLK(clk), .Q(n2229), .QN(n6) );
  DFFX1_HVT \key_round_reg[105]  ( .D(n3774), .CLK(clk), .Q(key_round[105]), 
        .QN(n2236) );
  DFFX1_HVT \keys_reg[7][106]  ( .D(n3773), .CLK(clk), .Q(n2227), .QN(n7) );
  DFFX1_HVT \key_round_reg[106]  ( .D(n3772), .CLK(clk), .Q(key_round[106]), 
        .QN(n2234) );
  DFFX1_HVT \keys_reg[7][107]  ( .D(n3771), .CLK(clk), .Q(n2225), .QN(n8) );
  DFFX1_HVT \key_round_reg[107]  ( .D(n3770), .CLK(clk), .Q(key_round[107]), 
        .QN(n2232) );
  DFFX1_HVT \keys_reg[7][108]  ( .D(n3769), .CLK(clk), .Q(n2223), .QN(n9) );
  DFFX1_HVT \key_round_reg[108]  ( .D(n3768), .CLK(clk), .Q(key_round[108]), 
        .QN(n2230) );
  DFFX1_HVT \keys_reg[7][109]  ( .D(n3767), .CLK(clk), .Q(n2221), .QN(n10) );
  DFFX1_HVT \key_round_reg[109]  ( .D(n3766), .CLK(clk), .Q(key_round[109]), 
        .QN(n2228) );
  DFFX1_HVT \keys_reg[7][110]  ( .D(n3765), .CLK(clk), .Q(n2219), .QN(n11) );
  DFFX1_HVT \key_round_reg[110]  ( .D(n3764), .CLK(clk), .Q(key_round[110]), 
        .QN(n2226) );
  DFFX1_HVT \keys_reg[7][111]  ( .D(n3763), .CLK(clk), .Q(n2217), .QN(n12) );
  DFFX1_HVT \key_round_reg[111]  ( .D(n3762), .CLK(clk), .Q(key_round[111]), 
        .QN(n2224) );
  DFFX1_HVT \keys_reg[7][112]  ( .D(n3761), .CLK(clk), .Q(n2215), .QN(n13) );
  DFFX1_HVT \key_round_reg[112]  ( .D(n3760), .CLK(clk), .Q(key_round[112]), 
        .QN(n2222) );
  DFFX1_HVT \keys_reg[7][113]  ( .D(n3759), .CLK(clk), .Q(n2213), .QN(n14) );
  DFFX1_HVT \key_round_reg[113]  ( .D(n3758), .CLK(clk), .Q(key_round[113]), 
        .QN(n2220) );
  DFFX1_HVT \keys_reg[7][114]  ( .D(n3757), .CLK(clk), .Q(n2211), .QN(n15) );
  DFFX1_HVT \key_round_reg[114]  ( .D(n3756), .CLK(clk), .Q(key_round[114]), 
        .QN(n2218) );
  DFFX1_HVT \keys_reg[7][115]  ( .D(n3755), .CLK(clk), .Q(n2209), .QN(n16) );
  DFFX1_HVT \key_round_reg[115]  ( .D(n3754), .CLK(clk), .Q(key_round[115]), 
        .QN(n2216) );
  DFFX1_HVT \keys_reg[7][116]  ( .D(n3753), .CLK(clk), .Q(n2207), .QN(n17) );
  DFFX1_HVT \key_round_reg[116]  ( .D(n3752), .CLK(clk), .Q(key_round[116]), 
        .QN(n2214) );
  DFFX1_HVT \keys_reg[7][117]  ( .D(n3751), .CLK(clk), .Q(n2205), .QN(n18) );
  DFFX1_HVT \key_round_reg[117]  ( .D(n3750), .CLK(clk), .Q(key_round[117]), 
        .QN(n2212) );
  DFFX1_HVT \keys_reg[7][118]  ( .D(n3749), .CLK(clk), .Q(n2203), .QN(n19) );
  DFFX1_HVT \key_round_reg[118]  ( .D(n3748), .CLK(clk), .Q(key_round[118]), 
        .QN(n2210) );
  DFFX1_HVT \keys_reg[7][119]  ( .D(n3747), .CLK(clk), .Q(n2201), .QN(n20) );
  DFFX1_HVT \key_round_reg[119]  ( .D(n3746), .CLK(clk), .Q(key_round[119]), 
        .QN(n2208) );
  DFFX1_HVT \keys_reg[7][120]  ( .D(n3745), .CLK(clk), .Q(n2199), .QN(n21) );
  DFFX1_HVT \key_round_reg[120]  ( .D(n3744), .CLK(clk), .Q(key_round[120]), 
        .QN(n2206) );
  DFFX1_HVT \keys_reg[7][121]  ( .D(n3743), .CLK(clk), .Q(n2197), .QN(n22) );
  DFFX1_HVT \key_round_reg[121]  ( .D(n3742), .CLK(clk), .Q(key_round[121]), 
        .QN(n2204) );
  DFFX1_HVT \keys_reg[7][122]  ( .D(n3741), .CLK(clk), .Q(n2195), .QN(n23) );
  DFFX1_HVT \key_round_reg[122]  ( .D(n3740), .CLK(clk), .Q(key_round[122]), 
        .QN(n2202) );
  DFFX1_HVT \keys_reg[7][123]  ( .D(n3739), .CLK(clk), .Q(n2193), .QN(n24) );
  DFFX1_HVT \key_round_reg[123]  ( .D(n3738), .CLK(clk), .Q(key_round[123]), 
        .QN(n2200) );
  DFFX1_HVT \keys_reg[7][124]  ( .D(n3737), .CLK(clk), .Q(n2191), .QN(n25) );
  DFFX1_HVT \key_round_reg[124]  ( .D(n3736), .CLK(clk), .Q(key_round[124]), 
        .QN(n2198) );
  DFFX1_HVT \keys_reg[7][125]  ( .D(n3735), .CLK(clk), .Q(n2189), .QN(n26) );
  DFFX1_HVT \key_round_reg[125]  ( .D(n3734), .CLK(clk), .Q(key_round[125]), 
        .QN(n2196) );
  DFFX1_HVT \keys_reg[7][126]  ( .D(n3733), .CLK(clk), .Q(n2187), .QN(n27) );
  DFFX1_HVT \key_round_reg[126]  ( .D(n3732), .CLK(clk), .Q(key_round[126]), 
        .QN(n2194) );
  DFFX1_HVT \keys_reg[7][127]  ( .D(n3731), .CLK(clk), .Q(n2185), .QN(n28) );
  DFFX1_HVT \key_round_reg[127]  ( .D(n3730), .CLK(clk), .Q(key_round[127]), 
        .QN(n2192) );
  DFFX1_HVT \keys_reg[7][82]  ( .D(n3729), .CLK(clk), .Q(n2183), .QN(n29) );
  DFFX1_HVT \key_round_reg[82]  ( .D(n3728), .CLK(clk), .Q(key_round[82]), 
        .QN(n2190) );
  DFFX1_HVT \keys_reg[7][83]  ( .D(n3727), .CLK(clk), .Q(n2181), .QN(n30) );
  DFFX1_HVT \key_round_reg[83]  ( .D(n3726), .CLK(clk), .Q(key_round[83]), 
        .QN(n2188) );
  DFFX1_HVT \keys_reg[7][84]  ( .D(n3725), .CLK(clk), .Q(n2179), .QN(n31) );
  DFFX1_HVT \key_round_reg[84]  ( .D(n3724), .CLK(clk), .Q(key_round[84]), 
        .QN(n2186) );
  DFFX1_HVT \keys_reg[7][85]  ( .D(n3723), .CLK(clk), .Q(n2177), .QN(n32) );
  DFFX1_HVT \key_round_reg[85]  ( .D(n3722), .CLK(clk), .Q(key_round[85]), 
        .QN(n2184) );
  DFFX1_HVT \keys_reg[7][86]  ( .D(n3721), .CLK(clk), .Q(n2175), .QN(n33) );
  DFFX1_HVT \key_round_reg[86]  ( .D(n3720), .CLK(clk), .Q(key_round[86]), 
        .QN(n2182) );
  DFFX1_HVT \keys_reg[7][87]  ( .D(n3719), .CLK(clk), .Q(n2173), .QN(n34) );
  DFFX1_HVT \key_round_reg[87]  ( .D(n3718), .CLK(clk), .Q(key_round[87]), 
        .QN(n2180) );
  DFFX1_HVT \keys_reg[7][88]  ( .D(n3717), .CLK(clk), .Q(n2171), .QN(n35) );
  DFFX1_HVT \key_round_reg[88]  ( .D(n3716), .CLK(clk), .Q(key_round[88]), 
        .QN(n2178) );
  DFFX1_HVT \keys_reg[7][89]  ( .D(n3715), .CLK(clk), .Q(n2169), .QN(n36) );
  DFFX1_HVT \key_round_reg[89]  ( .D(n3714), .CLK(clk), .Q(key_round[89]), 
        .QN(n2176) );
  DFFX1_HVT \keys_reg[7][90]  ( .D(n3713), .CLK(clk), .Q(n2167), .QN(n37) );
  DFFX1_HVT \key_round_reg[90]  ( .D(n3712), .CLK(clk), .Q(key_round[90]), 
        .QN(n2174) );
  DFFX1_HVT \keys_reg[7][91]  ( .D(n3711), .CLK(clk), .Q(n2165), .QN(n38) );
  DFFX1_HVT \key_round_reg[91]  ( .D(n3710), .CLK(clk), .Q(key_round[91]), 
        .QN(n2172) );
  DFFX1_HVT \keys_reg[7][92]  ( .D(n3709), .CLK(clk), .Q(n2163), .QN(n39) );
  DFFX1_HVT \key_round_reg[92]  ( .D(n3708), .CLK(clk), .Q(key_round[92]), 
        .QN(n2170) );
  DFFX1_HVT \keys_reg[7][93]  ( .D(n3707), .CLK(clk), .Q(n2161), .QN(n40) );
  DFFX1_HVT \key_round_reg[93]  ( .D(n3706), .CLK(clk), .Q(key_round[93]), 
        .QN(n2168) );
  DFFX1_HVT \keys_reg[7][94]  ( .D(n3705), .CLK(clk), .Q(n2159), .QN(n41) );
  DFFX1_HVT \key_round_reg[94]  ( .D(n3704), .CLK(clk), .Q(key_round[94]), 
        .QN(n2166) );
  DFFX1_HVT \keys_reg[7][95]  ( .D(n3703), .CLK(clk), .Q(n2157), .QN(n42) );
  DFFX1_HVT \key_round_reg[95]  ( .D(n3702), .CLK(clk), .Q(key_round[95]), 
        .QN(n2164) );
  DFFX1_HVT \keys_reg[7][96]  ( .D(n3701), .CLK(clk), .Q(n2155), .QN(n43) );
  DFFX1_HVT \key_round_reg[96]  ( .D(n3700), .CLK(clk), .Q(key_round[96]), 
        .QN(n2162) );
  DFFX1_HVT \keys_reg[7][97]  ( .D(n3699), .CLK(clk), .Q(n2153), .QN(n44) );
  DFFX1_HVT \key_round_reg[97]  ( .D(n3698), .CLK(clk), .Q(key_round[97]), 
        .QN(n2160) );
  DFFX1_HVT \keys_reg[7][0]  ( .D(n3697), .CLK(clk), .Q(n2151), .QN(n45) );
  DFFX1_HVT \key_round_reg[0]  ( .D(n3696), .CLK(clk), .Q(key_round[0]), .QN(
        n2158) );
  DFFX1_HVT \keys_reg[7][1]  ( .D(n3695), .CLK(clk), .Q(n2149), .QN(n46) );
  DFFX1_HVT \key_round_reg[1]  ( .D(n3694), .CLK(clk), .Q(key_round[1]), .QN(
        n2156) );
  DFFX1_HVT \keys_reg[7][2]  ( .D(n3693), .CLK(clk), .Q(n2147), .QN(n47) );
  DFFX1_HVT \key_round_reg[2]  ( .D(n3692), .CLK(clk), .Q(key_round[2]), .QN(
        n2154) );
  DFFX1_HVT \keys_reg[7][3]  ( .D(n3691), .CLK(clk), .Q(n2145), .QN(n48) );
  DFFX1_HVT \key_round_reg[3]  ( .D(n3690), .CLK(clk), .Q(key_round[3]), .QN(
        n2152) );
  DFFX1_HVT \keys_reg[7][4]  ( .D(n3689), .CLK(clk), .Q(n2143), .QN(n49) );
  DFFX1_HVT \key_round_reg[4]  ( .D(n3688), .CLK(clk), .Q(key_round[4]), .QN(
        n2150) );
  DFFX1_HVT \keys_reg[7][5]  ( .D(n3687), .CLK(clk), .Q(n2141), .QN(n50) );
  DFFX1_HVT \key_round_reg[5]  ( .D(n3686), .CLK(clk), .Q(key_round[5]), .QN(
        n2148) );
  DFFX1_HVT \keys_reg[7][6]  ( .D(n3685), .CLK(clk), .Q(n2139), .QN(n51) );
  DFFX1_HVT \key_round_reg[6]  ( .D(n3684), .CLK(clk), .Q(key_round[6]), .QN(
        n2146) );
  DFFX1_HVT \keys_reg[7][7]  ( .D(n3683), .CLK(clk), .Q(n2137), .QN(n52) );
  DFFX1_HVT \key_round_reg[7]  ( .D(n3682), .CLK(clk), .Q(key_round[7]), .QN(
        n2144) );
  DFFX1_HVT \keys_reg[7][8]  ( .D(n3681), .CLK(clk), .Q(n2135), .QN(n53) );
  DFFX1_HVT \key_round_reg[8]  ( .D(n3680), .CLK(clk), .Q(key_round[8]), .QN(
        n2142) );
  DFFX1_HVT \keys_reg[7][9]  ( .D(n3679), .CLK(clk), .Q(n2133), .QN(n54) );
  DFFX1_HVT \key_round_reg[9]  ( .D(n3678), .CLK(clk), .Q(key_round[9]), .QN(
        n2140) );
  DFFX1_HVT \keys_reg[7][10]  ( .D(n3677), .CLK(clk), .Q(n2131), .QN(n55) );
  DFFX1_HVT \key_round_reg[10]  ( .D(n3676), .CLK(clk), .Q(key_round[10]), 
        .QN(n2138) );
  DFFX1_HVT \keys_reg[7][11]  ( .D(n3675), .CLK(clk), .Q(n2129), .QN(n56) );
  DFFX1_HVT \key_round_reg[11]  ( .D(n3674), .CLK(clk), .Q(key_round[11]), 
        .QN(n2136) );
  DFFX1_HVT \keys_reg[7][12]  ( .D(n3673), .CLK(clk), .Q(n2127), .QN(n57) );
  DFFX1_HVT \key_round_reg[12]  ( .D(n3672), .CLK(clk), .Q(key_round[12]), 
        .QN(n2134) );
  DFFX1_HVT \keys_reg[7][13]  ( .D(n3671), .CLK(clk), .Q(n2125), .QN(n58) );
  DFFX1_HVT \key_round_reg[13]  ( .D(n3670), .CLK(clk), .Q(key_round[13]), 
        .QN(n2132) );
  DFFX1_HVT \keys_reg[7][14]  ( .D(n3669), .CLK(clk), .Q(n2123), .QN(n59) );
  DFFX1_HVT \key_round_reg[14]  ( .D(n3668), .CLK(clk), .Q(key_round[14]), 
        .QN(n2130) );
  DFFX1_HVT \keys_reg[7][15]  ( .D(n3667), .CLK(clk), .Q(n2121), .QN(n60) );
  DFFX1_HVT \key_round_reg[15]  ( .D(n3666), .CLK(clk), .Q(key_round[15]), 
        .QN(n2128) );
  DFFX1_HVT \keys_reg[7][16]  ( .D(n3665), .CLK(clk), .Q(n2119), .QN(n61) );
  DFFX1_HVT \key_round_reg[16]  ( .D(n3664), .CLK(clk), .Q(key_round[16]), 
        .QN(n2126) );
  DFFX1_HVT \keys_reg[7][17]  ( .D(n3663), .CLK(clk), .Q(n2117), .QN(n62) );
  DFFX1_HVT \key_round_reg[17]  ( .D(n3662), .CLK(clk), .Q(key_round[17]), 
        .QN(n2124) );
  DFFX1_HVT \keys_reg[7][18]  ( .D(n3661), .CLK(clk), .Q(n2115), .QN(n63) );
  DFFX1_HVT \key_round_reg[18]  ( .D(n3660), .CLK(clk), .Q(key_round[18]), 
        .QN(n2122) );
  DFFX1_HVT \keys_reg[7][19]  ( .D(n3659), .CLK(clk), .Q(n2113), .QN(n64) );
  DFFX1_HVT \key_round_reg[19]  ( .D(n3658), .CLK(clk), .Q(key_round[19]), 
        .QN(n2120) );
  DFFX1_HVT \keys_reg[7][20]  ( .D(n3657), .CLK(clk), .Q(n2111), .QN(n65) );
  DFFX1_HVT \key_round_reg[20]  ( .D(n3656), .CLK(clk), .Q(key_round[20]), 
        .QN(n2118) );
  DFFX1_HVT \keys_reg[7][21]  ( .D(n3655), .CLK(clk), .Q(n2109), .QN(n66) );
  DFFX1_HVT \key_round_reg[21]  ( .D(n3654), .CLK(clk), .Q(key_round[21]), 
        .QN(n2116) );
  DFFX1_HVT \keys_reg[7][22]  ( .D(n3653), .CLK(clk), .Q(n2107), .QN(n67) );
  DFFX1_HVT \key_round_reg[22]  ( .D(n3652), .CLK(clk), .Q(key_round[22]), 
        .QN(n2114) );
  DFFX1_HVT \keys_reg[7][23]  ( .D(n3651), .CLK(clk), .Q(n2105), .QN(n68) );
  DFFX1_HVT \key_round_reg[23]  ( .D(n3650), .CLK(clk), .Q(key_round[23]), 
        .QN(n2112) );
  DFFX1_HVT \keys_reg[7][24]  ( .D(n3649), .CLK(clk), .Q(n2103), .QN(n69) );
  DFFX1_HVT \key_round_reg[24]  ( .D(n3648), .CLK(clk), .Q(key_round[24]), 
        .QN(n2110) );
  DFFX1_HVT \keys_reg[7][25]  ( .D(n3647), .CLK(clk), .Q(n2101), .QN(n70) );
  DFFX1_HVT \key_round_reg[25]  ( .D(n3646), .CLK(clk), .Q(key_round[25]), 
        .QN(n2108) );
  DFFX1_HVT \keys_reg[7][26]  ( .D(n3645), .CLK(clk), .Q(n2099), .QN(n71) );
  DFFX1_HVT \key_round_reg[26]  ( .D(n3644), .CLK(clk), .Q(key_round[26]), 
        .QN(n2106) );
  DFFX1_HVT \keys_reg[7][27]  ( .D(n3643), .CLK(clk), .Q(n2097), .QN(n72) );
  DFFX1_HVT \key_round_reg[27]  ( .D(n3642), .CLK(clk), .Q(key_round[27]), 
        .QN(n2104) );
  DFFX1_HVT \keys_reg[7][28]  ( .D(n3641), .CLK(clk), .Q(n2095), .QN(n73) );
  DFFX1_HVT \key_round_reg[28]  ( .D(n3640), .CLK(clk), .Q(key_round[28]), 
        .QN(n2102) );
  DFFX1_HVT \keys_reg[7][29]  ( .D(n3639), .CLK(clk), .Q(n2093), .QN(n74) );
  DFFX1_HVT \key_round_reg[29]  ( .D(n3638), .CLK(clk), .Q(key_round[29]), 
        .QN(n2100) );
  DFFX1_HVT \keys_reg[7][30]  ( .D(n3637), .CLK(clk), .Q(n2091), .QN(n75) );
  DFFX1_HVT \key_round_reg[30]  ( .D(n3636), .CLK(clk), .Q(key_round[30]), 
        .QN(n2098) );
  DFFX1_HVT \keys_reg[7][31]  ( .D(n3635), .CLK(clk), .Q(n2089), .QN(n76) );
  DFFX1_HVT \key_round_reg[31]  ( .D(n3634), .CLK(clk), .Q(key_round[31]), 
        .QN(n2096) );
  DFFX1_HVT \keys_reg[7][32]  ( .D(n3633), .CLK(clk), .Q(n2087), .QN(n77) );
  DFFX1_HVT \key_round_reg[32]  ( .D(n3632), .CLK(clk), .Q(key_round[32]), 
        .QN(n2094) );
  DFFX1_HVT \keys_reg[7][33]  ( .D(n3631), .CLK(clk), .Q(n2085), .QN(n78) );
  DFFX1_HVT \key_round_reg[33]  ( .D(n3630), .CLK(clk), .Q(key_round[33]), 
        .QN(n2092) );
  DFFX1_HVT \keys_reg[7][34]  ( .D(n3629), .CLK(clk), .Q(n2083), .QN(n79) );
  DFFX1_HVT \key_round_reg[34]  ( .D(n3628), .CLK(clk), .Q(key_round[34]), 
        .QN(n2090) );
  DFFX1_HVT \keys_reg[7][35]  ( .D(n3627), .CLK(clk), .Q(n2081), .QN(n80) );
  DFFX1_HVT \key_round_reg[35]  ( .D(n3626), .CLK(clk), .Q(key_round[35]), 
        .QN(n2088) );
  DFFX1_HVT \keys_reg[7][36]  ( .D(n3625), .CLK(clk), .Q(n2079), .QN(n81) );
  DFFX1_HVT \key_round_reg[36]  ( .D(n3624), .CLK(clk), .Q(key_round[36]), 
        .QN(n2086) );
  DFFX1_HVT \keys_reg[7][37]  ( .D(n3623), .CLK(clk), .Q(n2077), .QN(n82) );
  DFFX1_HVT \key_round_reg[37]  ( .D(n3622), .CLK(clk), .Q(key_round[37]), 
        .QN(n2084) );
  DFFX1_HVT \keys_reg[7][38]  ( .D(n3621), .CLK(clk), .Q(n2075), .QN(n83) );
  DFFX1_HVT \key_round_reg[38]  ( .D(n3620), .CLK(clk), .Q(key_round[38]), 
        .QN(n2082) );
  DFFX1_HVT \keys_reg[7][39]  ( .D(n3619), .CLK(clk), .Q(n2073), .QN(n84) );
  DFFX1_HVT \key_round_reg[39]  ( .D(n3618), .CLK(clk), .Q(key_round[39]), 
        .QN(n2080) );
  DFFX1_HVT \keys_reg[7][40]  ( .D(n3617), .CLK(clk), .Q(n2071), .QN(n85) );
  DFFX1_HVT \key_round_reg[40]  ( .D(n3616), .CLK(clk), .Q(key_round[40]), 
        .QN(n2078) );
  DFFX1_HVT \keys_reg[7][41]  ( .D(n3615), .CLK(clk), .Q(n2069), .QN(n86) );
  DFFX1_HVT \key_round_reg[41]  ( .D(n3614), .CLK(clk), .Q(key_round[41]), 
        .QN(n2076) );
  DFFX1_HVT \keys_reg[7][42]  ( .D(n3613), .CLK(clk), .Q(n2067), .QN(n87) );
  DFFX1_HVT \key_round_reg[42]  ( .D(n3612), .CLK(clk), .Q(key_round[42]), 
        .QN(n2074) );
  DFFX1_HVT \keys_reg[7][43]  ( .D(n3611), .CLK(clk), .Q(n2065), .QN(n88) );
  DFFX1_HVT \key_round_reg[43]  ( .D(n3610), .CLK(clk), .Q(key_round[43]), 
        .QN(n2072) );
  DFFX1_HVT \keys_reg[7][44]  ( .D(n3609), .CLK(clk), .Q(n2063), .QN(n89) );
  DFFX1_HVT \key_round_reg[44]  ( .D(n3608), .CLK(clk), .Q(key_round[44]), 
        .QN(n2070) );
  DFFX1_HVT \keys_reg[7][45]  ( .D(n3607), .CLK(clk), .Q(n2061), .QN(n90) );
  DFFX1_HVT \key_round_reg[45]  ( .D(n3606), .CLK(clk), .Q(key_round[45]), 
        .QN(n2068) );
  DFFX1_HVT \keys_reg[7][46]  ( .D(n3605), .CLK(clk), .Q(n2059), .QN(n91) );
  DFFX1_HVT \key_round_reg[46]  ( .D(n3604), .CLK(clk), .Q(key_round[46]), 
        .QN(n2066) );
  DFFX1_HVT \keys_reg[7][47]  ( .D(n3603), .CLK(clk), .Q(n2057), .QN(n92) );
  DFFX1_HVT \key_round_reg[47]  ( .D(n3602), .CLK(clk), .Q(key_round[47]), 
        .QN(n2064) );
  DFFX1_HVT \keys_reg[7][48]  ( .D(n3601), .CLK(clk), .Q(n2055), .QN(n93) );
  DFFX1_HVT \key_round_reg[48]  ( .D(n3600), .CLK(clk), .Q(key_round[48]), 
        .QN(n2062) );
  DFFX1_HVT \keys_reg[7][81]  ( .D(n3599), .CLK(clk), .Q(n2053), .QN(n94) );
  DFFX1_HVT \key_round_reg[81]  ( .D(n3598), .CLK(clk), .Q(key_round[81]), 
        .QN(n2060) );
  DFFX1_HVT \keys_reg[7][80]  ( .D(n3597), .CLK(clk), .Q(n2051), .QN(n95) );
  DFFX1_HVT \key_round_reg[80]  ( .D(n3596), .CLK(clk), .Q(key_round[80]), 
        .QN(n2058) );
  DFFX1_HVT \keys_reg[7][79]  ( .D(n3595), .CLK(clk), .Q(n2049), .QN(n96) );
  DFFX1_HVT \key_round_reg[79]  ( .D(n3594), .CLK(clk), .Q(key_round[79]), 
        .QN(n2056) );
  DFFX1_HVT \keys_reg[7][78]  ( .D(n3593), .CLK(clk), .Q(n2047), .QN(n97) );
  DFFX1_HVT \key_round_reg[78]  ( .D(n3592), .CLK(clk), .Q(key_round[78]), 
        .QN(n2054) );
  DFFX1_HVT \keys_reg[7][77]  ( .D(n3591), .CLK(clk), .Q(n2045), .QN(n98) );
  DFFX1_HVT \key_round_reg[77]  ( .D(n3590), .CLK(clk), .Q(key_round[77]), 
        .QN(n2052) );
  DFFX1_HVT \keys_reg[7][76]  ( .D(n3589), .CLK(clk), .Q(n2043), .QN(n99) );
  DFFX1_HVT \key_round_reg[76]  ( .D(n3588), .CLK(clk), .Q(key_round[76]), 
        .QN(n2050) );
  DFFX1_HVT \keys_reg[7][75]  ( .D(n3587), .CLK(clk), .Q(n2041), .QN(n100) );
  DFFX1_HVT \key_round_reg[75]  ( .D(n3586), .CLK(clk), .Q(key_round[75]), 
        .QN(n2048) );
  DFFX1_HVT \keys_reg[7][74]  ( .D(n3585), .CLK(clk), .Q(n2039), .QN(n101) );
  DFFX1_HVT \key_round_reg[74]  ( .D(n3584), .CLK(clk), .Q(key_round[74]), 
        .QN(n2046) );
  DFFX1_HVT \keys_reg[7][73]  ( .D(n3583), .CLK(clk), .Q(n2037), .QN(n102) );
  DFFX1_HVT \key_round_reg[73]  ( .D(n3582), .CLK(clk), .Q(key_round[73]), 
        .QN(n2044) );
  DFFX1_HVT \keys_reg[7][72]  ( .D(n3581), .CLK(clk), .Q(n2035), .QN(n103) );
  DFFX1_HVT \key_round_reg[72]  ( .D(n3580), .CLK(clk), .Q(key_round[72]), 
        .QN(n2042) );
  DFFX1_HVT \keys_reg[7][71]  ( .D(n3579), .CLK(clk), .Q(n2033), .QN(n104) );
  DFFX1_HVT \key_round_reg[71]  ( .D(n3578), .CLK(clk), .Q(key_round[71]), 
        .QN(n2040) );
  DFFX1_HVT \keys_reg[7][70]  ( .D(n3577), .CLK(clk), .Q(n2031), .QN(n105) );
  DFFX1_HVT \key_round_reg[70]  ( .D(n3576), .CLK(clk), .Q(key_round[70]), 
        .QN(n2038) );
  DFFX1_HVT \keys_reg[7][69]  ( .D(n3575), .CLK(clk), .Q(n2029), .QN(n106) );
  DFFX1_HVT \key_round_reg[69]  ( .D(n3574), .CLK(clk), .Q(key_round[69]), 
        .QN(n2036) );
  DFFX1_HVT \keys_reg[7][68]  ( .D(n3573), .CLK(clk), .Q(n2027), .QN(n107) );
  DFFX1_HVT \key_round_reg[68]  ( .D(n3572), .CLK(clk), .Q(key_round[68]), 
        .QN(n2034) );
  DFFX1_HVT \keys_reg[7][67]  ( .D(n3571), .CLK(clk), .Q(n2025), .QN(n108) );
  DFFX1_HVT \key_round_reg[67]  ( .D(n3570), .CLK(clk), .Q(key_round[67]), 
        .QN(n2032) );
  DFFX1_HVT \keys_reg[7][66]  ( .D(n3569), .CLK(clk), .Q(n2023), .QN(n109) );
  DFFX1_HVT \key_round_reg[66]  ( .D(n3568), .CLK(clk), .Q(key_round[66]), 
        .QN(n2030) );
  DFFX1_HVT \keys_reg[7][65]  ( .D(n3567), .CLK(clk), .Q(n2021), .QN(n110) );
  DFFX1_HVT \key_round_reg[65]  ( .D(n3566), .CLK(clk), .Q(key_round[65]), 
        .QN(n2028) );
  DFFX1_HVT \keys_reg[7][64]  ( .D(n3565), .CLK(clk), .Q(n2019), .QN(n111) );
  DFFX1_HVT \key_round_reg[64]  ( .D(n3564), .CLK(clk), .Q(key_round[64]), 
        .QN(n2026) );
  DFFX1_HVT \keys_reg[7][63]  ( .D(n3563), .CLK(clk), .Q(n2017), .QN(n112) );
  DFFX1_HVT \key_round_reg[63]  ( .D(n3562), .CLK(clk), .Q(key_round[63]), 
        .QN(n2024) );
  DFFX1_HVT \keys_reg[7][62]  ( .D(n3561), .CLK(clk), .Q(n2015), .QN(n113) );
  DFFX1_HVT \key_round_reg[62]  ( .D(n3560), .CLK(clk), .Q(key_round[62]), 
        .QN(n2022) );
  DFFX1_HVT \keys_reg[7][61]  ( .D(n3559), .CLK(clk), .Q(n2013), .QN(n114) );
  DFFX1_HVT \key_round_reg[61]  ( .D(n3558), .CLK(clk), .Q(key_round[61]), 
        .QN(n2020) );
  DFFX1_HVT \keys_reg[7][60]  ( .D(n3557), .CLK(clk), .Q(n2011), .QN(n115) );
  DFFX1_HVT \key_round_reg[60]  ( .D(n3556), .CLK(clk), .Q(key_round[60]), 
        .QN(n2018) );
  DFFX1_HVT \keys_reg[7][59]  ( .D(n3555), .CLK(clk), .Q(n2009), .QN(n116) );
  DFFX1_HVT \key_round_reg[59]  ( .D(n3554), .CLK(clk), .Q(key_round[59]), 
        .QN(n2016) );
  DFFX1_HVT \keys_reg[7][58]  ( .D(n3553), .CLK(clk), .Q(n2007), .QN(n117) );
  DFFX1_HVT \key_round_reg[58]  ( .D(n3552), .CLK(clk), .Q(key_round[58]), 
        .QN(n2014) );
  DFFX1_HVT \keys_reg[7][57]  ( .D(n3551), .CLK(clk), .Q(n2005), .QN(n118) );
  DFFX1_HVT \key_round_reg[57]  ( .D(n3550), .CLK(clk), .Q(key_round[57]), 
        .QN(n2012) );
  DFFX1_HVT \keys_reg[7][56]  ( .D(n3549), .CLK(clk), .Q(n2003), .QN(n119) );
  DFFX1_HVT \key_round_reg[56]  ( .D(n3548), .CLK(clk), .Q(key_round[56]), 
        .QN(n2010) );
  DFFX1_HVT \keys_reg[7][55]  ( .D(n3547), .CLK(clk), .Q(n2001), .QN(n120) );
  DFFX1_HVT \key_round_reg[55]  ( .D(n3546), .CLK(clk), .Q(key_round[55]), 
        .QN(n2008) );
  DFFX1_HVT \keys_reg[7][54]  ( .D(n3545), .CLK(clk), .Q(n1999), .QN(n121) );
  DFFX1_HVT \key_round_reg[54]  ( .D(n3544), .CLK(clk), .Q(key_round[54]), 
        .QN(n2006) );
  DFFX1_HVT \keys_reg[7][53]  ( .D(n3543), .CLK(clk), .Q(n1997), .QN(n122) );
  DFFX1_HVT \key_round_reg[53]  ( .D(n3542), .CLK(clk), .Q(key_round[53]), 
        .QN(n2004) );
  DFFX1_HVT \keys_reg[7][52]  ( .D(n3541), .CLK(clk), .Q(n1995), .QN(n123) );
  DFFX1_HVT \key_round_reg[52]  ( .D(n3540), .CLK(clk), .Q(key_round[52]), 
        .QN(n2002) );
  DFFX1_HVT \keys_reg[7][51]  ( .D(n3539), .CLK(clk), .Q(n1993), .QN(n124) );
  DFFX1_HVT \key_round_reg[51]  ( .D(n3538), .CLK(clk), .Q(key_round[51]), 
        .QN(n2000) );
  DFFX1_HVT \keys_reg[7][50]  ( .D(n3537), .CLK(clk), .Q(n1992), .QN(n125) );
  DFFX1_HVT \key_round_reg[50]  ( .D(n3536), .CLK(clk), .Q(key_round[50]), 
        .QN(n1998) );
  DFFX1_HVT \keys_reg[7][49]  ( .D(n3535), .CLK(clk), .Q(n1991), .QN(n126) );
  DFFX1_HVT \key_round_reg[49]  ( .D(n3534), .CLK(clk), .Q(key_round[49]), 
        .QN(n1996) );
  DFFX1_HVT \keys_reg[7][98]  ( .D(n3533), .CLK(clk), .Q(n1990), .QN(n127) );
  DFFX1_HVT \key_round_reg[98]  ( .D(n3532), .CLK(clk), .Q(key_round[98]), 
        .QN(n1994) );
  keygen_1 key ( .round_num(round_number), .keyin(prev_key), .keyout(keyout)
         );
  AO21X1_HVT U3 ( .A1(n1412), .A2(state[0]), .A3(n1413), .Y(n5205) );
  NAND2X0_HVT U4 ( .A1(n3398), .A2(n1414), .Y(n5204) );
  NAND4X0_HVT U5 ( .A1(n1415), .A2(n1416), .A3(n1417), .A4(n1418), .Y(n5203)
         );
  OA21X1_HVT U6 ( .A1(n3399), .A2(n1419), .A3(n1420), .Y(n1418) );
  NAND3X0_HVT U7 ( .A1(n1421), .A2(n1422), .A3(n1423), .Y(n5202) );
  NAND2X0_HVT U8 ( .A1(n1412), .A2(state[2]), .Y(n1421) );
  INVX0_HVT U9 ( .A(n1424), .Y(n1412) );
  NAND2X0_HVT U10 ( .A1(n1425), .A2(n1426), .Y(n5201) );
  MUX21X1_HVT U11 ( .A1(n1427), .A2(n1989), .S0(n1428), .Y(n1425) );
  MUX21X1_HVT U12 ( .A1(n1429), .A2(round_number[1]), .S0(n1428), .Y(n5200) );
  NAND2X0_HVT U13 ( .A1(n1430), .A2(n1420), .Y(n1429) );
  MUX21X1_HVT U14 ( .A1(n1431), .A2(round_number[2]), .S0(n1428), .Y(n5199) );
  NAND2X0_HVT U15 ( .A1(n1423), .A2(n1414), .Y(n1431) );
  AND3X1_HVT U16 ( .A1(n1432), .A2(n1433), .A3(n1415), .Y(n1423) );
  MUX21X1_HVT U17 ( .A1(n1434), .A2(round_number[3]), .S0(n1428), .Y(n5198) );
  NAND3X0_HVT U18 ( .A1(n1435), .A2(n1436), .A3(n1417), .Y(n1434) );
  AO222X1_HVT U19 ( .A1(local_key[0]), .A2(n1437), .A3(keyout[0]), .A4(n1438), 
        .A5(prev_key[0]), .A6(n1428), .Y(n5197) );
  AO222X1_HVT U20 ( .A1(local_key[1]), .A2(n1437), .A3(keyout[1]), .A4(n1438), 
        .A5(prev_key[1]), .A6(n1428), .Y(n5196) );
  AO222X1_HVT U21 ( .A1(local_key[2]), .A2(n1437), .A3(keyout[2]), .A4(n1438), 
        .A5(prev_key[2]), .A6(n1428), .Y(n5195) );
  AO222X1_HVT U22 ( .A1(local_key[3]), .A2(n1437), .A3(keyout[3]), .A4(n1438), 
        .A5(prev_key[3]), .A6(n1428), .Y(n5194) );
  AO222X1_HVT U23 ( .A1(local_key[4]), .A2(n1437), .A3(keyout[4]), .A4(n1438), 
        .A5(prev_key[4]), .A6(n1428), .Y(n5193) );
  AO222X1_HVT U24 ( .A1(local_key[5]), .A2(n1437), .A3(keyout[5]), .A4(n1438), 
        .A5(prev_key[5]), .A6(n1428), .Y(n5192) );
  AO222X1_HVT U25 ( .A1(local_key[6]), .A2(n1437), .A3(keyout[6]), .A4(n1438), 
        .A5(prev_key[6]), .A6(n1428), .Y(n5191) );
  AO222X1_HVT U26 ( .A1(local_key[7]), .A2(n1437), .A3(keyout[7]), .A4(n1438), 
        .A5(prev_key[7]), .A6(n1428), .Y(n5190) );
  AO222X1_HVT U27 ( .A1(local_key[8]), .A2(n1437), .A3(keyout[8]), .A4(n1438), 
        .A5(prev_key[8]), .A6(n1428), .Y(n5189) );
  AO222X1_HVT U28 ( .A1(local_key[9]), .A2(n1437), .A3(keyout[9]), .A4(n1438), 
        .A5(prev_key[9]), .A6(n1428), .Y(n5188) );
  AO222X1_HVT U29 ( .A1(local_key[10]), .A2(n1437), .A3(keyout[10]), .A4(n1438), .A5(prev_key[10]), .A6(n1428), .Y(n5187) );
  AO222X1_HVT U30 ( .A1(local_key[11]), .A2(n1437), .A3(keyout[11]), .A4(n1438), .A5(prev_key[11]), .A6(n1428), .Y(n5186) );
  AO222X1_HVT U31 ( .A1(local_key[12]), .A2(n1437), .A3(keyout[12]), .A4(n1438), .A5(prev_key[12]), .A6(n1428), .Y(n5185) );
  AO222X1_HVT U32 ( .A1(local_key[13]), .A2(n1437), .A3(keyout[13]), .A4(n1438), .A5(prev_key[13]), .A6(n1428), .Y(n5184) );
  AO222X1_HVT U33 ( .A1(local_key[14]), .A2(n1437), .A3(keyout[14]), .A4(n1438), .A5(prev_key[14]), .A6(n1428), .Y(n5183) );
  AO222X1_HVT U34 ( .A1(local_key[15]), .A2(n1437), .A3(keyout[15]), .A4(n1438), .A5(prev_key[15]), .A6(n1428), .Y(n5182) );
  AO222X1_HVT U35 ( .A1(local_key[16]), .A2(n1437), .A3(keyout[16]), .A4(n1438), .A5(prev_key[16]), .A6(n1428), .Y(n5181) );
  AO222X1_HVT U36 ( .A1(local_key[17]), .A2(n1437), .A3(keyout[17]), .A4(n1438), .A5(prev_key[17]), .A6(n1428), .Y(n5180) );
  AO222X1_HVT U37 ( .A1(local_key[18]), .A2(n1437), .A3(keyout[18]), .A4(n1438), .A5(prev_key[18]), .A6(n1428), .Y(n5179) );
  AO222X1_HVT U38 ( .A1(local_key[19]), .A2(n1437), .A3(keyout[19]), .A4(n1438), .A5(prev_key[19]), .A6(n1428), .Y(n5178) );
  AO222X1_HVT U39 ( .A1(local_key[20]), .A2(n1437), .A3(keyout[20]), .A4(n1438), .A5(prev_key[20]), .A6(n1428), .Y(n5177) );
  AO222X1_HVT U40 ( .A1(local_key[21]), .A2(n1437), .A3(keyout[21]), .A4(n1438), .A5(prev_key[21]), .A6(n1428), .Y(n5176) );
  AO222X1_HVT U41 ( .A1(local_key[22]), .A2(n1437), .A3(keyout[22]), .A4(n1438), .A5(prev_key[22]), .A6(n1428), .Y(n5175) );
  AO222X1_HVT U42 ( .A1(local_key[23]), .A2(n1437), .A3(keyout[23]), .A4(n1438), .A5(prev_key[23]), .A6(n1428), .Y(n5174) );
  AO222X1_HVT U43 ( .A1(local_key[24]), .A2(n1437), .A3(keyout[24]), .A4(n1438), .A5(prev_key[24]), .A6(n1428), .Y(n5173) );
  AO222X1_HVT U44 ( .A1(local_key[25]), .A2(n1437), .A3(keyout[25]), .A4(n1438), .A5(prev_key[25]), .A6(n1428), .Y(n5172) );
  AO222X1_HVT U45 ( .A1(local_key[26]), .A2(n1437), .A3(keyout[26]), .A4(n1438), .A5(prev_key[26]), .A6(n1428), .Y(n5171) );
  AO222X1_HVT U46 ( .A1(local_key[27]), .A2(n1437), .A3(keyout[27]), .A4(n1438), .A5(prev_key[27]), .A6(n1428), .Y(n5170) );
  AO222X1_HVT U47 ( .A1(local_key[28]), .A2(n1437), .A3(keyout[28]), .A4(n1438), .A5(prev_key[28]), .A6(n1428), .Y(n5169) );
  AO222X1_HVT U48 ( .A1(local_key[29]), .A2(n1437), .A3(keyout[29]), .A4(n1438), .A5(prev_key[29]), .A6(n1428), .Y(n5168) );
  AO222X1_HVT U49 ( .A1(local_key[30]), .A2(n1437), .A3(keyout[30]), .A4(n1438), .A5(prev_key[30]), .A6(n1428), .Y(n5167) );
  AO222X1_HVT U50 ( .A1(local_key[31]), .A2(n1437), .A3(keyout[31]), .A4(n1438), .A5(prev_key[31]), .A6(n1428), .Y(n5166) );
  AO222X1_HVT U51 ( .A1(local_key[32]), .A2(n1437), .A3(keyout[32]), .A4(n1438), .A5(prev_key[32]), .A6(n1428), .Y(n5165) );
  AO222X1_HVT U52 ( .A1(local_key[33]), .A2(n1437), .A3(keyout[33]), .A4(n1438), .A5(prev_key[33]), .A6(n1428), .Y(n5164) );
  AO222X1_HVT U53 ( .A1(local_key[34]), .A2(n1437), .A3(keyout[34]), .A4(n1438), .A5(prev_key[34]), .A6(n1428), .Y(n5163) );
  AO222X1_HVT U54 ( .A1(local_key[35]), .A2(n1437), .A3(keyout[35]), .A4(n1438), .A5(prev_key[35]), .A6(n1428), .Y(n5162) );
  AO222X1_HVT U55 ( .A1(local_key[36]), .A2(n1437), .A3(keyout[36]), .A4(n1438), .A5(prev_key[36]), .A6(n1428), .Y(n5161) );
  AO222X1_HVT U56 ( .A1(local_key[37]), .A2(n1437), .A3(keyout[37]), .A4(n1438), .A5(prev_key[37]), .A6(n1428), .Y(n5160) );
  AO222X1_HVT U57 ( .A1(local_key[38]), .A2(n1437), .A3(keyout[38]), .A4(n1438), .A5(prev_key[38]), .A6(n1428), .Y(n5159) );
  AO222X1_HVT U58 ( .A1(local_key[39]), .A2(n1437), .A3(keyout[39]), .A4(n1438), .A5(prev_key[39]), .A6(n1428), .Y(n5158) );
  AO222X1_HVT U59 ( .A1(local_key[40]), .A2(n1437), .A3(keyout[40]), .A4(n1438), .A5(prev_key[40]), .A6(n1428), .Y(n5157) );
  AO222X1_HVT U60 ( .A1(local_key[41]), .A2(n1437), .A3(keyout[41]), .A4(n1438), .A5(prev_key[41]), .A6(n1428), .Y(n5156) );
  AO222X1_HVT U61 ( .A1(local_key[42]), .A2(n1437), .A3(keyout[42]), .A4(n1438), .A5(prev_key[42]), .A6(n1428), .Y(n5155) );
  AO222X1_HVT U62 ( .A1(local_key[43]), .A2(n1437), .A3(keyout[43]), .A4(n1438), .A5(prev_key[43]), .A6(n1428), .Y(n5154) );
  AO222X1_HVT U63 ( .A1(local_key[44]), .A2(n1437), .A3(keyout[44]), .A4(n1438), .A5(prev_key[44]), .A6(n1428), .Y(n5153) );
  AO222X1_HVT U64 ( .A1(local_key[45]), .A2(n1437), .A3(keyout[45]), .A4(n1438), .A5(prev_key[45]), .A6(n1428), .Y(n5152) );
  AO222X1_HVT U65 ( .A1(local_key[46]), .A2(n1437), .A3(keyout[46]), .A4(n1438), .A5(prev_key[46]), .A6(n1428), .Y(n5151) );
  AO222X1_HVT U66 ( .A1(local_key[47]), .A2(n1437), .A3(keyout[47]), .A4(n1438), .A5(prev_key[47]), .A6(n1428), .Y(n5150) );
  AO222X1_HVT U67 ( .A1(local_key[48]), .A2(n1437), .A3(keyout[48]), .A4(n1438), .A5(prev_key[48]), .A6(n1428), .Y(n5149) );
  AO222X1_HVT U68 ( .A1(local_key[49]), .A2(n1437), .A3(keyout[49]), .A4(n1438), .A5(prev_key[49]), .A6(n1428), .Y(n5148) );
  AO222X1_HVT U69 ( .A1(local_key[50]), .A2(n1437), .A3(keyout[50]), .A4(n1438), .A5(prev_key[50]), .A6(n1428), .Y(n5147) );
  AO222X1_HVT U70 ( .A1(local_key[51]), .A2(n1437), .A3(keyout[51]), .A4(n1438), .A5(prev_key[51]), .A6(n1428), .Y(n5146) );
  AO222X1_HVT U71 ( .A1(local_key[52]), .A2(n1437), .A3(keyout[52]), .A4(n1438), .A5(prev_key[52]), .A6(n1428), .Y(n5145) );
  AO222X1_HVT U72 ( .A1(local_key[53]), .A2(n1437), .A3(keyout[53]), .A4(n1438), .A5(prev_key[53]), .A6(n1428), .Y(n5144) );
  AO222X1_HVT U73 ( .A1(local_key[54]), .A2(n1437), .A3(keyout[54]), .A4(n1438), .A5(prev_key[54]), .A6(n1428), .Y(n5143) );
  AO222X1_HVT U74 ( .A1(local_key[55]), .A2(n1437), .A3(keyout[55]), .A4(n1438), .A5(prev_key[55]), .A6(n1428), .Y(n5142) );
  AO222X1_HVT U75 ( .A1(local_key[56]), .A2(n1437), .A3(keyout[56]), .A4(n1438), .A5(prev_key[56]), .A6(n1428), .Y(n5141) );
  AO222X1_HVT U76 ( .A1(local_key[57]), .A2(n1437), .A3(keyout[57]), .A4(n1438), .A5(prev_key[57]), .A6(n1428), .Y(n5140) );
  AO222X1_HVT U77 ( .A1(local_key[58]), .A2(n1437), .A3(keyout[58]), .A4(n1438), .A5(prev_key[58]), .A6(n1428), .Y(n5139) );
  AO222X1_HVT U78 ( .A1(local_key[59]), .A2(n1437), .A3(keyout[59]), .A4(n1438), .A5(prev_key[59]), .A6(n1428), .Y(n5138) );
  AO222X1_HVT U79 ( .A1(local_key[60]), .A2(n1437), .A3(keyout[60]), .A4(n1438), .A5(prev_key[60]), .A6(n1428), .Y(n5137) );
  AO222X1_HVT U80 ( .A1(local_key[61]), .A2(n1437), .A3(keyout[61]), .A4(n1438), .A5(prev_key[61]), .A6(n1428), .Y(n5136) );
  AO222X1_HVT U81 ( .A1(local_key[62]), .A2(n1437), .A3(keyout[62]), .A4(n1438), .A5(prev_key[62]), .A6(n1428), .Y(n5135) );
  AO222X1_HVT U82 ( .A1(local_key[63]), .A2(n1437), .A3(keyout[63]), .A4(n1438), .A5(prev_key[63]), .A6(n1428), .Y(n5134) );
  AO222X1_HVT U83 ( .A1(local_key[64]), .A2(n1437), .A3(keyout[64]), .A4(n1438), .A5(prev_key[64]), .A6(n1428), .Y(n5133) );
  AO222X1_HVT U84 ( .A1(local_key[65]), .A2(n1437), .A3(keyout[65]), .A4(n1438), .A5(prev_key[65]), .A6(n1428), .Y(n5132) );
  AO222X1_HVT U85 ( .A1(local_key[66]), .A2(n1437), .A3(keyout[66]), .A4(n1438), .A5(prev_key[66]), .A6(n1428), .Y(n5131) );
  AO222X1_HVT U86 ( .A1(local_key[67]), .A2(n1437), .A3(keyout[67]), .A4(n1438), .A5(prev_key[67]), .A6(n1428), .Y(n5130) );
  AO222X1_HVT U87 ( .A1(local_key[68]), .A2(n1437), .A3(keyout[68]), .A4(n1438), .A5(prev_key[68]), .A6(n1428), .Y(n5129) );
  AO222X1_HVT U88 ( .A1(local_key[69]), .A2(n1437), .A3(keyout[69]), .A4(n1438), .A5(prev_key[69]), .A6(n1428), .Y(n5128) );
  AO222X1_HVT U89 ( .A1(local_key[70]), .A2(n1437), .A3(keyout[70]), .A4(n1438), .A5(prev_key[70]), .A6(n1428), .Y(n5127) );
  AO222X1_HVT U90 ( .A1(local_key[71]), .A2(n1437), .A3(keyout[71]), .A4(n1438), .A5(prev_key[71]), .A6(n1428), .Y(n5126) );
  AO222X1_HVT U91 ( .A1(local_key[72]), .A2(n1437), .A3(keyout[72]), .A4(n1438), .A5(prev_key[72]), .A6(n1428), .Y(n5125) );
  AO222X1_HVT U92 ( .A1(local_key[73]), .A2(n1437), .A3(keyout[73]), .A4(n1438), .A5(prev_key[73]), .A6(n1428), .Y(n5124) );
  AO222X1_HVT U93 ( .A1(local_key[74]), .A2(n1437), .A3(keyout[74]), .A4(n1438), .A5(prev_key[74]), .A6(n1428), .Y(n5123) );
  AO222X1_HVT U94 ( .A1(local_key[75]), .A2(n1437), .A3(keyout[75]), .A4(n1438), .A5(prev_key[75]), .A6(n1428), .Y(n5122) );
  AO222X1_HVT U95 ( .A1(local_key[76]), .A2(n1437), .A3(keyout[76]), .A4(n1438), .A5(prev_key[76]), .A6(n1428), .Y(n5121) );
  AO222X1_HVT U96 ( .A1(local_key[77]), .A2(n1437), .A3(keyout[77]), .A4(n1438), .A5(prev_key[77]), .A6(n1428), .Y(n5120) );
  AO222X1_HVT U97 ( .A1(local_key[78]), .A2(n1437), .A3(keyout[78]), .A4(n1438), .A5(prev_key[78]), .A6(n1428), .Y(n5119) );
  AO222X1_HVT U98 ( .A1(local_key[79]), .A2(n1437), .A3(keyout[79]), .A4(n1438), .A5(prev_key[79]), .A6(n1428), .Y(n5118) );
  AO222X1_HVT U99 ( .A1(local_key[80]), .A2(n1437), .A3(keyout[80]), .A4(n1438), .A5(prev_key[80]), .A6(n1428), .Y(n5117) );
  AO222X1_HVT U100 ( .A1(local_key[81]), .A2(n1437), .A3(keyout[81]), .A4(
        n1438), .A5(prev_key[81]), .A6(n1428), .Y(n5116) );
  AO222X1_HVT U101 ( .A1(local_key[82]), .A2(n1437), .A3(keyout[82]), .A4(
        n1438), .A5(prev_key[82]), .A6(n1428), .Y(n5115) );
  AO222X1_HVT U102 ( .A1(local_key[83]), .A2(n1437), .A3(keyout[83]), .A4(
        n1438), .A5(prev_key[83]), .A6(n1428), .Y(n5114) );
  AO222X1_HVT U103 ( .A1(local_key[84]), .A2(n1437), .A3(keyout[84]), .A4(
        n1438), .A5(prev_key[84]), .A6(n1428), .Y(n5113) );
  AO222X1_HVT U104 ( .A1(local_key[85]), .A2(n1437), .A3(keyout[85]), .A4(
        n1438), .A5(prev_key[85]), .A6(n1428), .Y(n5112) );
  AO222X1_HVT U105 ( .A1(local_key[86]), .A2(n1437), .A3(keyout[86]), .A4(
        n1438), .A5(prev_key[86]), .A6(n1428), .Y(n5111) );
  AO222X1_HVT U106 ( .A1(local_key[87]), .A2(n1437), .A3(keyout[87]), .A4(
        n1438), .A5(prev_key[87]), .A6(n1428), .Y(n5110) );
  AO222X1_HVT U107 ( .A1(local_key[88]), .A2(n1437), .A3(keyout[88]), .A4(
        n1438), .A5(prev_key[88]), .A6(n1428), .Y(n5109) );
  AO222X1_HVT U108 ( .A1(local_key[89]), .A2(n1437), .A3(keyout[89]), .A4(
        n1438), .A5(prev_key[89]), .A6(n1428), .Y(n5108) );
  AO222X1_HVT U109 ( .A1(local_key[90]), .A2(n1437), .A3(keyout[90]), .A4(
        n1438), .A5(prev_key[90]), .A6(n1428), .Y(n5107) );
  AO222X1_HVT U110 ( .A1(local_key[91]), .A2(n1437), .A3(keyout[91]), .A4(
        n1438), .A5(prev_key[91]), .A6(n1428), .Y(n5106) );
  AO222X1_HVT U111 ( .A1(local_key[92]), .A2(n1437), .A3(keyout[92]), .A4(
        n1438), .A5(prev_key[92]), .A6(n1428), .Y(n5105) );
  AO222X1_HVT U112 ( .A1(local_key[93]), .A2(n1437), .A3(keyout[93]), .A4(
        n1438), .A5(prev_key[93]), .A6(n1428), .Y(n5104) );
  AO222X1_HVT U113 ( .A1(local_key[94]), .A2(n1437), .A3(keyout[94]), .A4(
        n1438), .A5(prev_key[94]), .A6(n1428), .Y(n5103) );
  AO222X1_HVT U114 ( .A1(local_key[95]), .A2(n1437), .A3(keyout[95]), .A4(
        n1438), .A5(prev_key[95]), .A6(n1428), .Y(n5102) );
  AO222X1_HVT U115 ( .A1(local_key[96]), .A2(n1437), .A3(keyout[96]), .A4(
        n1438), .A5(prev_key[96]), .A6(n1428), .Y(n5101) );
  AO222X1_HVT U116 ( .A1(local_key[97]), .A2(n1437), .A3(keyout[97]), .A4(
        n1438), .A5(prev_key[97]), .A6(n1428), .Y(n5100) );
  AO222X1_HVT U117 ( .A1(local_key[98]), .A2(n1437), .A3(keyout[98]), .A4(
        n1438), .A5(prev_key[98]), .A6(n1428), .Y(n5099) );
  AO222X1_HVT U118 ( .A1(local_key[99]), .A2(n1437), .A3(keyout[99]), .A4(
        n1438), .A5(prev_key[99]), .A6(n1428), .Y(n5098) );
  AO222X1_HVT U119 ( .A1(local_key[100]), .A2(n1437), .A3(keyout[100]), .A4(
        n1438), .A5(prev_key[100]), .A6(n1428), .Y(n5097) );
  AO222X1_HVT U120 ( .A1(local_key[101]), .A2(n1437), .A3(keyout[101]), .A4(
        n1438), .A5(prev_key[101]), .A6(n1428), .Y(n5096) );
  AO222X1_HVT U121 ( .A1(local_key[102]), .A2(n1437), .A3(keyout[102]), .A4(
        n1438), .A5(prev_key[102]), .A6(n1428), .Y(n5095) );
  AO222X1_HVT U122 ( .A1(local_key[103]), .A2(n1437), .A3(keyout[103]), .A4(
        n1438), .A5(prev_key[103]), .A6(n1428), .Y(n5094) );
  AO222X1_HVT U123 ( .A1(local_key[104]), .A2(n1437), .A3(keyout[104]), .A4(
        n1438), .A5(prev_key[104]), .A6(n1428), .Y(n5093) );
  AO222X1_HVT U124 ( .A1(local_key[105]), .A2(n1437), .A3(keyout[105]), .A4(
        n1438), .A5(prev_key[105]), .A6(n1428), .Y(n5092) );
  AO222X1_HVT U125 ( .A1(local_key[106]), .A2(n1437), .A3(keyout[106]), .A4(
        n1438), .A5(prev_key[106]), .A6(n1428), .Y(n5091) );
  AO222X1_HVT U126 ( .A1(local_key[107]), .A2(n1437), .A3(keyout[107]), .A4(
        n1438), .A5(prev_key[107]), .A6(n1428), .Y(n5090) );
  AO222X1_HVT U127 ( .A1(local_key[108]), .A2(n1437), .A3(keyout[108]), .A4(
        n1438), .A5(prev_key[108]), .A6(n1428), .Y(n5089) );
  AO222X1_HVT U128 ( .A1(local_key[109]), .A2(n1437), .A3(keyout[109]), .A4(
        n1438), .A5(prev_key[109]), .A6(n1428), .Y(n5088) );
  AO222X1_HVT U129 ( .A1(local_key[110]), .A2(n1437), .A3(keyout[110]), .A4(
        n1438), .A5(prev_key[110]), .A6(n1428), .Y(n5087) );
  AO222X1_HVT U130 ( .A1(local_key[111]), .A2(n1437), .A3(keyout[111]), .A4(
        n1438), .A5(prev_key[111]), .A6(n1428), .Y(n5086) );
  AO222X1_HVT U131 ( .A1(local_key[112]), .A2(n1437), .A3(keyout[112]), .A4(
        n1438), .A5(prev_key[112]), .A6(n1428), .Y(n5085) );
  AO222X1_HVT U132 ( .A1(local_key[113]), .A2(n1437), .A3(keyout[113]), .A4(
        n1438), .A5(prev_key[113]), .A6(n1428), .Y(n5084) );
  AO222X1_HVT U133 ( .A1(local_key[114]), .A2(n1437), .A3(keyout[114]), .A4(
        n1438), .A5(prev_key[114]), .A6(n1428), .Y(n5083) );
  AO222X1_HVT U134 ( .A1(local_key[115]), .A2(n1437), .A3(keyout[115]), .A4(
        n1438), .A5(prev_key[115]), .A6(n1428), .Y(n5082) );
  AO222X1_HVT U135 ( .A1(local_key[116]), .A2(n1437), .A3(keyout[116]), .A4(
        n1438), .A5(prev_key[116]), .A6(n1428), .Y(n5081) );
  AO222X1_HVT U136 ( .A1(local_key[117]), .A2(n1437), .A3(keyout[117]), .A4(
        n1438), .A5(prev_key[117]), .A6(n1428), .Y(n5080) );
  AO222X1_HVT U137 ( .A1(local_key[118]), .A2(n1437), .A3(keyout[118]), .A4(
        n1438), .A5(prev_key[118]), .A6(n1428), .Y(n5079) );
  AO222X1_HVT U138 ( .A1(local_key[119]), .A2(n1437), .A3(keyout[119]), .A4(
        n1438), .A5(prev_key[119]), .A6(n1428), .Y(n5078) );
  AO222X1_HVT U139 ( .A1(local_key[120]), .A2(n1437), .A3(keyout[120]), .A4(
        n1438), .A5(prev_key[120]), .A6(n1428), .Y(n5077) );
  AO222X1_HVT U140 ( .A1(local_key[121]), .A2(n1437), .A3(keyout[121]), .A4(
        n1438), .A5(prev_key[121]), .A6(n1428), .Y(n5076) );
  AO222X1_HVT U141 ( .A1(local_key[122]), .A2(n1437), .A3(keyout[122]), .A4(
        n1438), .A5(prev_key[122]), .A6(n1428), .Y(n5075) );
  AO222X1_HVT U142 ( .A1(local_key[123]), .A2(n1437), .A3(keyout[123]), .A4(
        n1438), .A5(prev_key[123]), .A6(n1428), .Y(n5074) );
  AO222X1_HVT U143 ( .A1(local_key[124]), .A2(n1437), .A3(keyout[124]), .A4(
        n1438), .A5(prev_key[124]), .A6(n1428), .Y(n5073) );
  AO222X1_HVT U144 ( .A1(local_key[125]), .A2(n1437), .A3(keyout[125]), .A4(
        n1438), .A5(prev_key[125]), .A6(n1428), .Y(n5072) );
  AO222X1_HVT U145 ( .A1(local_key[126]), .A2(n1437), .A3(keyout[126]), .A4(
        n1438), .A5(prev_key[126]), .A6(n1428), .Y(n5071) );
  AO222X1_HVT U146 ( .A1(local_key[127]), .A2(n1437), .A3(keyout[127]), .A4(
        n1438), .A5(prev_key[127]), .A6(n1428), .Y(n5070) );
  AND2X1_HVT U147 ( .A1(n1439), .A2(n1419), .Y(n1438) );
  INVX0_HVT U148 ( .A(n1426), .Y(n1437) );
  NAND2X0_HVT U149 ( .A1(n1440), .A2(n1439), .Y(n1426) );
  INVX0_HVT U150 ( .A(n1428), .Y(n1439) );
  NAND2X0_HVT U151 ( .A1(n3528), .A2(n1424), .Y(n1428) );
  OR2X1_HVT U152 ( .A1(n1419), .A2(n1440), .Y(n1424) );
  NAND2X0_HVT U153 ( .A1(n1441), .A2(n1427), .Y(n1419) );
  AND3X1_HVT U154 ( .A1(n1417), .A2(n1415), .A3(n1430), .Y(n1427) );
  AND2X1_HVT U155 ( .A1(n1422), .A2(n1414), .Y(n1430) );
  INVX0_HVT U156 ( .A(n1413), .Y(n1441) );
  NAND3X0_HVT U157 ( .A1(n1433), .A2(n1436), .A3(n1420), .Y(n1413) );
  AND3X1_HVT U158 ( .A1(n1432), .A2(n1442), .A3(n1435), .Y(n1420) );
  MUX21X1_HVT U159 ( .A1(n3527), .A2(local_key[99]), .S0(n1443), .Y(n5068) );
  MUX21X1_HVT U160 ( .A1(n3526), .A2(local_key[100]), .S0(n1443), .Y(n5067) );
  MUX21X1_HVT U161 ( .A1(n3525), .A2(local_key[101]), .S0(n1443), .Y(n5066) );
  MUX21X1_HVT U162 ( .A1(n3524), .A2(local_key[102]), .S0(n1443), .Y(n5065) );
  MUX21X1_HVT U163 ( .A1(n3523), .A2(local_key[103]), .S0(n1443), .Y(n5064) );
  MUX21X1_HVT U164 ( .A1(n3522), .A2(local_key[104]), .S0(n1443), .Y(n5063) );
  MUX21X1_HVT U165 ( .A1(n3521), .A2(local_key[105]), .S0(n1443), .Y(n5062) );
  MUX21X1_HVT U166 ( .A1(n3520), .A2(local_key[106]), .S0(n1443), .Y(n5061) );
  MUX21X1_HVT U167 ( .A1(n3519), .A2(local_key[107]), .S0(n1443), .Y(n5060) );
  MUX21X1_HVT U168 ( .A1(n3518), .A2(local_key[108]), .S0(n1443), .Y(n5059) );
  MUX21X1_HVT U169 ( .A1(n3517), .A2(local_key[109]), .S0(n1443), .Y(n5058) );
  MUX21X1_HVT U170 ( .A1(n3516), .A2(local_key[110]), .S0(n1443), .Y(n5057) );
  MUX21X1_HVT U171 ( .A1(n3515), .A2(local_key[111]), .S0(n1443), .Y(n5056) );
  MUX21X1_HVT U172 ( .A1(n3514), .A2(local_key[112]), .S0(n1443), .Y(n5055) );
  MUX21X1_HVT U173 ( .A1(n3513), .A2(local_key[113]), .S0(n1443), .Y(n5054) );
  MUX21X1_HVT U174 ( .A1(n3512), .A2(local_key[114]), .S0(n1443), .Y(n5053) );
  MUX21X1_HVT U175 ( .A1(n3511), .A2(local_key[115]), .S0(n1443), .Y(n5052) );
  MUX21X1_HVT U176 ( .A1(n3510), .A2(local_key[116]), .S0(n1443), .Y(n5051) );
  MUX21X1_HVT U177 ( .A1(n3509), .A2(local_key[117]), .S0(n1443), .Y(n5050) );
  MUX21X1_HVT U178 ( .A1(n3508), .A2(local_key[118]), .S0(n1443), .Y(n5049) );
  MUX21X1_HVT U179 ( .A1(n3507), .A2(local_key[119]), .S0(n1443), .Y(n5048) );
  MUX21X1_HVT U180 ( .A1(n3506), .A2(local_key[120]), .S0(n1443), .Y(n5047) );
  MUX21X1_HVT U181 ( .A1(n3505), .A2(local_key[121]), .S0(n1443), .Y(n5046) );
  MUX21X1_HVT U182 ( .A1(n3504), .A2(local_key[122]), .S0(n1443), .Y(n5045) );
  MUX21X1_HVT U183 ( .A1(n3503), .A2(local_key[123]), .S0(n1443), .Y(n5044) );
  MUX21X1_HVT U184 ( .A1(n3502), .A2(local_key[124]), .S0(n1443), .Y(n5043) );
  MUX21X1_HVT U185 ( .A1(n3501), .A2(local_key[125]), .S0(n1443), .Y(n5042) );
  MUX21X1_HVT U186 ( .A1(n3500), .A2(local_key[126]), .S0(n1443), .Y(n5041) );
  MUX21X1_HVT U187 ( .A1(n3499), .A2(local_key[127]), .S0(n1443), .Y(n5040) );
  MUX21X1_HVT U188 ( .A1(n3498), .A2(local_key[77]), .S0(n1443), .Y(n5039) );
  MUX21X1_HVT U189 ( .A1(n3497), .A2(local_key[78]), .S0(n1443), .Y(n5038) );
  MUX21X1_HVT U190 ( .A1(n3496), .A2(local_key[79]), .S0(n1443), .Y(n5037) );
  MUX21X1_HVT U191 ( .A1(n3495), .A2(local_key[80]), .S0(n1443), .Y(n5036) );
  MUX21X1_HVT U192 ( .A1(n3494), .A2(local_key[81]), .S0(n1443), .Y(n5035) );
  MUX21X1_HVT U193 ( .A1(n3493), .A2(local_key[82]), .S0(n1443), .Y(n5034) );
  MUX21X1_HVT U194 ( .A1(n3492), .A2(local_key[83]), .S0(n1443), .Y(n5033) );
  MUX21X1_HVT U195 ( .A1(n3491), .A2(local_key[84]), .S0(n1443), .Y(n5032) );
  MUX21X1_HVT U196 ( .A1(n3490), .A2(local_key[85]), .S0(n1443), .Y(n5031) );
  MUX21X1_HVT U197 ( .A1(n3489), .A2(local_key[86]), .S0(n1443), .Y(n5030) );
  MUX21X1_HVT U198 ( .A1(n3488), .A2(local_key[87]), .S0(n1443), .Y(n5029) );
  MUX21X1_HVT U199 ( .A1(n3487), .A2(local_key[88]), .S0(n1443), .Y(n5028) );
  MUX21X1_HVT U200 ( .A1(n3486), .A2(local_key[89]), .S0(n1443), .Y(n5027) );
  MUX21X1_HVT U201 ( .A1(n3485), .A2(local_key[90]), .S0(n1443), .Y(n5026) );
  MUX21X1_HVT U202 ( .A1(n3484), .A2(local_key[91]), .S0(n1443), .Y(n5025) );
  MUX21X1_HVT U203 ( .A1(n3483), .A2(local_key[92]), .S0(n1443), .Y(n5024) );
  MUX21X1_HVT U204 ( .A1(n3482), .A2(local_key[93]), .S0(n1443), .Y(n5023) );
  MUX21X1_HVT U205 ( .A1(n3481), .A2(local_key[94]), .S0(n1443), .Y(n5022) );
  MUX21X1_HVT U206 ( .A1(n3480), .A2(local_key[95]), .S0(n1443), .Y(n5021) );
  MUX21X1_HVT U207 ( .A1(n3479), .A2(local_key[96]), .S0(n1443), .Y(n5020) );
  MUX21X1_HVT U208 ( .A1(n3478), .A2(local_key[97]), .S0(n1443), .Y(n5019) );
  MUX21X1_HVT U209 ( .A1(n3477), .A2(local_key[0]), .S0(n1443), .Y(n5018) );
  MUX21X1_HVT U210 ( .A1(n3476), .A2(local_key[1]), .S0(n1443), .Y(n5017) );
  MUX21X1_HVT U211 ( .A1(n3475), .A2(local_key[2]), .S0(n1443), .Y(n5016) );
  MUX21X1_HVT U212 ( .A1(n3474), .A2(local_key[3]), .S0(n1443), .Y(n5015) );
  MUX21X1_HVT U213 ( .A1(n3473), .A2(local_key[4]), .S0(n1443), .Y(n5014) );
  MUX21X1_HVT U214 ( .A1(n3472), .A2(local_key[5]), .S0(n1443), .Y(n5013) );
  MUX21X1_HVT U215 ( .A1(n3471), .A2(local_key[6]), .S0(n1443), .Y(n5012) );
  MUX21X1_HVT U216 ( .A1(n3470), .A2(local_key[7]), .S0(n1443), .Y(n5011) );
  MUX21X1_HVT U217 ( .A1(n3469), .A2(local_key[8]), .S0(n1443), .Y(n5010) );
  MUX21X1_HVT U218 ( .A1(n3468), .A2(local_key[9]), .S0(n1443), .Y(n5009) );
  MUX21X1_HVT U219 ( .A1(n3467), .A2(local_key[10]), .S0(n1443), .Y(n5008) );
  MUX21X1_HVT U220 ( .A1(n3466), .A2(local_key[11]), .S0(n1443), .Y(n5007) );
  MUX21X1_HVT U221 ( .A1(n3465), .A2(local_key[12]), .S0(n1443), .Y(n5006) );
  MUX21X1_HVT U222 ( .A1(n3464), .A2(local_key[13]), .S0(n1443), .Y(n5005) );
  MUX21X1_HVT U223 ( .A1(n3463), .A2(local_key[14]), .S0(n1443), .Y(n5004) );
  MUX21X1_HVT U224 ( .A1(n3462), .A2(local_key[15]), .S0(n1443), .Y(n5003) );
  MUX21X1_HVT U225 ( .A1(n3461), .A2(local_key[16]), .S0(n1443), .Y(n5002) );
  MUX21X1_HVT U226 ( .A1(n3460), .A2(local_key[17]), .S0(n1443), .Y(n5001) );
  MUX21X1_HVT U227 ( .A1(n3459), .A2(local_key[18]), .S0(n1443), .Y(n5000) );
  MUX21X1_HVT U228 ( .A1(n3458), .A2(local_key[19]), .S0(n1443), .Y(n4999) );
  MUX21X1_HVT U229 ( .A1(n3457), .A2(local_key[20]), .S0(n1443), .Y(n4998) );
  MUX21X1_HVT U230 ( .A1(n3456), .A2(local_key[21]), .S0(n1443), .Y(n4997) );
  MUX21X1_HVT U231 ( .A1(n3455), .A2(local_key[22]), .S0(n1443), .Y(n4996) );
  MUX21X1_HVT U232 ( .A1(n3454), .A2(local_key[23]), .S0(n1443), .Y(n4995) );
  MUX21X1_HVT U233 ( .A1(n3453), .A2(local_key[24]), .S0(n1443), .Y(n4994) );
  MUX21X1_HVT U234 ( .A1(n3452), .A2(local_key[25]), .S0(n1443), .Y(n4993) );
  MUX21X1_HVT U235 ( .A1(n3451), .A2(local_key[26]), .S0(n1443), .Y(n4992) );
  MUX21X1_HVT U236 ( .A1(n3450), .A2(local_key[27]), .S0(n1443), .Y(n4991) );
  MUX21X1_HVT U237 ( .A1(n3449), .A2(local_key[28]), .S0(n1443), .Y(n4990) );
  MUX21X1_HVT U238 ( .A1(n3448), .A2(local_key[29]), .S0(n1443), .Y(n4989) );
  MUX21X1_HVT U239 ( .A1(n3447), .A2(local_key[30]), .S0(n1443), .Y(n4988) );
  MUX21X1_HVT U240 ( .A1(n3446), .A2(local_key[31]), .S0(n1443), .Y(n4987) );
  MUX21X1_HVT U241 ( .A1(n3445), .A2(local_key[32]), .S0(n1443), .Y(n4986) );
  MUX21X1_HVT U242 ( .A1(n3444), .A2(local_key[33]), .S0(n1443), .Y(n4985) );
  MUX21X1_HVT U243 ( .A1(n3443), .A2(local_key[34]), .S0(n1443), .Y(n4984) );
  MUX21X1_HVT U244 ( .A1(n3442), .A2(local_key[35]), .S0(n1443), .Y(n4983) );
  MUX21X1_HVT U245 ( .A1(n3441), .A2(local_key[36]), .S0(n1443), .Y(n4982) );
  MUX21X1_HVT U246 ( .A1(n3440), .A2(local_key[37]), .S0(n1443), .Y(n4981) );
  MUX21X1_HVT U247 ( .A1(n3439), .A2(local_key[38]), .S0(n1443), .Y(n4980) );
  MUX21X1_HVT U248 ( .A1(n3438), .A2(local_key[39]), .S0(n1443), .Y(n4979) );
  MUX21X1_HVT U249 ( .A1(n3437), .A2(local_key[40]), .S0(n1443), .Y(n4978) );
  MUX21X1_HVT U250 ( .A1(n3436), .A2(local_key[41]), .S0(n1443), .Y(n4977) );
  MUX21X1_HVT U251 ( .A1(n3435), .A2(local_key[42]), .S0(n1443), .Y(n4976) );
  MUX21X1_HVT U252 ( .A1(n3434), .A2(local_key[43]), .S0(n1443), .Y(n4975) );
  MUX21X1_HVT U253 ( .A1(n3433), .A2(local_key[44]), .S0(n1443), .Y(n4974) );
  MUX21X1_HVT U254 ( .A1(n3432), .A2(local_key[45]), .S0(n1443), .Y(n4973) );
  MUX21X1_HVT U255 ( .A1(n3431), .A2(local_key[46]), .S0(n1443), .Y(n4972) );
  MUX21X1_HVT U256 ( .A1(n3430), .A2(local_key[47]), .S0(n1443), .Y(n4971) );
  MUX21X1_HVT U257 ( .A1(n3429), .A2(local_key[48]), .S0(n1443), .Y(n4970) );
  MUX21X1_HVT U258 ( .A1(n3428), .A2(local_key[76]), .S0(n1443), .Y(n4969) );
  MUX21X1_HVT U259 ( .A1(n3427), .A2(local_key[75]), .S0(n1443), .Y(n4968) );
  MUX21X1_HVT U260 ( .A1(n3426), .A2(local_key[74]), .S0(n1443), .Y(n4967) );
  MUX21X1_HVT U261 ( .A1(n3425), .A2(local_key[73]), .S0(n1443), .Y(n4966) );
  MUX21X1_HVT U262 ( .A1(n3424), .A2(local_key[72]), .S0(n1443), .Y(n4965) );
  MUX21X1_HVT U263 ( .A1(n3423), .A2(local_key[71]), .S0(n1443), .Y(n4964) );
  MUX21X1_HVT U264 ( .A1(n3422), .A2(local_key[70]), .S0(n1443), .Y(n4963) );
  MUX21X1_HVT U265 ( .A1(n3421), .A2(local_key[69]), .S0(n1443), .Y(n4962) );
  MUX21X1_HVT U266 ( .A1(n3420), .A2(local_key[68]), .S0(n1443), .Y(n4961) );
  MUX21X1_HVT U267 ( .A1(n3419), .A2(local_key[67]), .S0(n1443), .Y(n4960) );
  MUX21X1_HVT U268 ( .A1(n3418), .A2(local_key[66]), .S0(n1443), .Y(n4959) );
  MUX21X1_HVT U269 ( .A1(n3417), .A2(local_key[65]), .S0(n1443), .Y(n4958) );
  MUX21X1_HVT U270 ( .A1(n3416), .A2(local_key[64]), .S0(n1443), .Y(n4957) );
  MUX21X1_HVT U271 ( .A1(n3415), .A2(local_key[63]), .S0(n1443), .Y(n4956) );
  MUX21X1_HVT U272 ( .A1(n3414), .A2(local_key[62]), .S0(n1443), .Y(n4955) );
  MUX21X1_HVT U273 ( .A1(n3413), .A2(local_key[61]), .S0(n1443), .Y(n4954) );
  MUX21X1_HVT U274 ( .A1(n3412), .A2(local_key[60]), .S0(n1443), .Y(n4953) );
  MUX21X1_HVT U275 ( .A1(n3411), .A2(local_key[59]), .S0(n1443), .Y(n4952) );
  MUX21X1_HVT U276 ( .A1(n3410), .A2(local_key[58]), .S0(n1443), .Y(n4951) );
  MUX21X1_HVT U277 ( .A1(n3409), .A2(local_key[57]), .S0(n1443), .Y(n4950) );
  MUX21X1_HVT U278 ( .A1(n3408), .A2(local_key[56]), .S0(n1443), .Y(n4949) );
  MUX21X1_HVT U279 ( .A1(n3407), .A2(local_key[55]), .S0(n1443), .Y(n4948) );
  MUX21X1_HVT U280 ( .A1(n3406), .A2(local_key[54]), .S0(n1443), .Y(n4947) );
  MUX21X1_HVT U281 ( .A1(n3405), .A2(local_key[53]), .S0(n1443), .Y(n4946) );
  MUX21X1_HVT U282 ( .A1(n3404), .A2(local_key[52]), .S0(n1443), .Y(n4945) );
  MUX21X1_HVT U283 ( .A1(n3403), .A2(local_key[51]), .S0(n1443), .Y(n4944) );
  MUX21X1_HVT U284 ( .A1(n3402), .A2(local_key[50]), .S0(n1443), .Y(n4943) );
  MUX21X1_HVT U285 ( .A1(n3401), .A2(local_key[49]), .S0(n1443), .Y(n4942) );
  MUX21X1_HVT U286 ( .A1(n3400), .A2(local_key[98]), .S0(n1443), .Y(n4941) );
  AND2X1_HVT U287 ( .A1(n1440), .A2(n3528), .Y(n1443) );
  INVX0_HVT U288 ( .A(n1416), .Y(n1440) );
  NAND2X0_HVT U289 ( .A1(n1444), .A2(n899), .Y(n1416) );
  NAND2X0_HVT U290 ( .A1(n1988), .A2(n1445), .Y(n4940) );
  NAND3X0_HVT U291 ( .A1(n1446), .A2(n898), .A3(state[0]), .Y(n1445) );
  MUX21X1_HVT U292 ( .A1(n3397), .A2(keyout[0]), .S0(n1447), .Y(n4939) );
  MUX21X1_HVT U293 ( .A1(n3396), .A2(keyout[0]), .S0(n1448), .Y(n4938) );
  MUX21X1_HVT U294 ( .A1(n3395), .A2(keyout[0]), .S0(n1449), .Y(n4937) );
  MUX21X1_HVT U295 ( .A1(n3394), .A2(keyout[0]), .S0(n1450), .Y(n4936) );
  MUX21X1_HVT U296 ( .A1(n3393), .A2(keyout[0]), .S0(n1451), .Y(n4935) );
  MUX21X1_HVT U297 ( .A1(n3392), .A2(keyout[0]), .S0(n1452), .Y(n4934) );
  MUX21X1_HVT U298 ( .A1(n3391), .A2(keyout[0]), .S0(n1453), .Y(n4933) );
  MUX21X1_HVT U299 ( .A1(n3390), .A2(keyout[0]), .S0(n1454), .Y(n4932) );
  MUX21X1_HVT U300 ( .A1(n3389), .A2(keyout[1]), .S0(n1447), .Y(n4931) );
  MUX21X1_HVT U301 ( .A1(n3388), .A2(keyout[1]), .S0(n1448), .Y(n4930) );
  MUX21X1_HVT U302 ( .A1(n3387), .A2(keyout[1]), .S0(n1449), .Y(n4929) );
  MUX21X1_HVT U303 ( .A1(n3386), .A2(keyout[1]), .S0(n1450), .Y(n4928) );
  MUX21X1_HVT U304 ( .A1(n3385), .A2(keyout[1]), .S0(n1451), .Y(n4927) );
  MUX21X1_HVT U305 ( .A1(n3384), .A2(keyout[1]), .S0(n1452), .Y(n4926) );
  MUX21X1_HVT U306 ( .A1(n3383), .A2(keyout[1]), .S0(n1453), .Y(n4925) );
  MUX21X1_HVT U307 ( .A1(n3382), .A2(keyout[1]), .S0(n1454), .Y(n4924) );
  MUX21X1_HVT U308 ( .A1(n3381), .A2(keyout[2]), .S0(n1447), .Y(n4923) );
  MUX21X1_HVT U309 ( .A1(n3380), .A2(keyout[2]), .S0(n1448), .Y(n4922) );
  MUX21X1_HVT U310 ( .A1(n3379), .A2(keyout[2]), .S0(n1449), .Y(n4921) );
  MUX21X1_HVT U311 ( .A1(n3378), .A2(keyout[2]), .S0(n1450), .Y(n4920) );
  MUX21X1_HVT U312 ( .A1(n3377), .A2(keyout[2]), .S0(n1451), .Y(n4919) );
  MUX21X1_HVT U313 ( .A1(n3376), .A2(keyout[2]), .S0(n1452), .Y(n4918) );
  MUX21X1_HVT U314 ( .A1(n3375), .A2(keyout[2]), .S0(n1453), .Y(n4917) );
  MUX21X1_HVT U315 ( .A1(n3374), .A2(keyout[2]), .S0(n1454), .Y(n4916) );
  MUX21X1_HVT U316 ( .A1(n3373), .A2(keyout[3]), .S0(n1447), .Y(n4915) );
  MUX21X1_HVT U317 ( .A1(n3372), .A2(keyout[3]), .S0(n1448), .Y(n4914) );
  MUX21X1_HVT U318 ( .A1(n3371), .A2(keyout[3]), .S0(n1449), .Y(n4913) );
  MUX21X1_HVT U319 ( .A1(n3370), .A2(keyout[3]), .S0(n1450), .Y(n4912) );
  MUX21X1_HVT U320 ( .A1(n3369), .A2(keyout[3]), .S0(n1451), .Y(n4911) );
  MUX21X1_HVT U321 ( .A1(n3368), .A2(keyout[3]), .S0(n1452), .Y(n4910) );
  MUX21X1_HVT U322 ( .A1(n3367), .A2(keyout[3]), .S0(n1453), .Y(n4909) );
  MUX21X1_HVT U323 ( .A1(n3366), .A2(keyout[3]), .S0(n1454), .Y(n4908) );
  MUX21X1_HVT U324 ( .A1(n3365), .A2(keyout[4]), .S0(n1447), .Y(n4907) );
  MUX21X1_HVT U325 ( .A1(n3364), .A2(keyout[4]), .S0(n1448), .Y(n4906) );
  MUX21X1_HVT U326 ( .A1(n3363), .A2(keyout[4]), .S0(n1449), .Y(n4905) );
  MUX21X1_HVT U327 ( .A1(n3362), .A2(keyout[4]), .S0(n1450), .Y(n4904) );
  MUX21X1_HVT U328 ( .A1(n3361), .A2(keyout[4]), .S0(n1451), .Y(n4903) );
  MUX21X1_HVT U329 ( .A1(n3360), .A2(keyout[4]), .S0(n1452), .Y(n4902) );
  MUX21X1_HVT U330 ( .A1(n3359), .A2(keyout[4]), .S0(n1453), .Y(n4901) );
  MUX21X1_HVT U331 ( .A1(n3358), .A2(keyout[4]), .S0(n1454), .Y(n4900) );
  MUX21X1_HVT U332 ( .A1(n3357), .A2(keyout[5]), .S0(n1447), .Y(n4899) );
  MUX21X1_HVT U333 ( .A1(n3356), .A2(keyout[5]), .S0(n1448), .Y(n4898) );
  MUX21X1_HVT U334 ( .A1(n3355), .A2(keyout[5]), .S0(n1449), .Y(n4897) );
  MUX21X1_HVT U335 ( .A1(n3354), .A2(keyout[5]), .S0(n1450), .Y(n4896) );
  MUX21X1_HVT U336 ( .A1(n3353), .A2(keyout[5]), .S0(n1451), .Y(n4895) );
  MUX21X1_HVT U337 ( .A1(n3352), .A2(keyout[5]), .S0(n1452), .Y(n4894) );
  MUX21X1_HVT U338 ( .A1(n3351), .A2(keyout[5]), .S0(n1453), .Y(n4893) );
  MUX21X1_HVT U339 ( .A1(n3350), .A2(keyout[5]), .S0(n1454), .Y(n4892) );
  MUX21X1_HVT U340 ( .A1(n3349), .A2(keyout[6]), .S0(n1447), .Y(n4891) );
  MUX21X1_HVT U341 ( .A1(n3348), .A2(keyout[6]), .S0(n1448), .Y(n4890) );
  MUX21X1_HVT U342 ( .A1(n3347), .A2(keyout[6]), .S0(n1449), .Y(n4889) );
  MUX21X1_HVT U343 ( .A1(n3346), .A2(keyout[6]), .S0(n1450), .Y(n4888) );
  MUX21X1_HVT U344 ( .A1(n3345), .A2(keyout[6]), .S0(n1451), .Y(n4887) );
  MUX21X1_HVT U345 ( .A1(n3344), .A2(keyout[6]), .S0(n1452), .Y(n4886) );
  MUX21X1_HVT U346 ( .A1(n3343), .A2(keyout[6]), .S0(n1453), .Y(n4885) );
  MUX21X1_HVT U347 ( .A1(n3342), .A2(keyout[6]), .S0(n1454), .Y(n4884) );
  MUX21X1_HVT U348 ( .A1(n3341), .A2(keyout[7]), .S0(n1447), .Y(n4883) );
  MUX21X1_HVT U349 ( .A1(n3340), .A2(keyout[7]), .S0(n1448), .Y(n4882) );
  MUX21X1_HVT U350 ( .A1(n3339), .A2(keyout[7]), .S0(n1449), .Y(n4881) );
  MUX21X1_HVT U351 ( .A1(n3338), .A2(keyout[7]), .S0(n1450), .Y(n4880) );
  MUX21X1_HVT U352 ( .A1(n3337), .A2(keyout[7]), .S0(n1451), .Y(n4879) );
  MUX21X1_HVT U353 ( .A1(n3336), .A2(keyout[7]), .S0(n1452), .Y(n4878) );
  MUX21X1_HVT U354 ( .A1(n3335), .A2(keyout[7]), .S0(n1453), .Y(n4877) );
  MUX21X1_HVT U355 ( .A1(n3334), .A2(keyout[7]), .S0(n1454), .Y(n4876) );
  MUX21X1_HVT U356 ( .A1(n3333), .A2(keyout[8]), .S0(n1447), .Y(n4875) );
  MUX21X1_HVT U357 ( .A1(n3332), .A2(keyout[8]), .S0(n1448), .Y(n4874) );
  MUX21X1_HVT U358 ( .A1(n3331), .A2(keyout[8]), .S0(n1449), .Y(n4873) );
  MUX21X1_HVT U359 ( .A1(n3330), .A2(keyout[8]), .S0(n1450), .Y(n4872) );
  MUX21X1_HVT U360 ( .A1(n3329), .A2(keyout[8]), .S0(n1451), .Y(n4871) );
  MUX21X1_HVT U361 ( .A1(n3328), .A2(keyout[8]), .S0(n1452), .Y(n4870) );
  MUX21X1_HVT U362 ( .A1(n3327), .A2(keyout[8]), .S0(n1453), .Y(n4869) );
  MUX21X1_HVT U363 ( .A1(n3326), .A2(keyout[8]), .S0(n1454), .Y(n4868) );
  MUX21X1_HVT U364 ( .A1(n3325), .A2(keyout[9]), .S0(n1447), .Y(n4867) );
  MUX21X1_HVT U365 ( .A1(n3324), .A2(keyout[9]), .S0(n1448), .Y(n4866) );
  MUX21X1_HVT U366 ( .A1(n3323), .A2(keyout[9]), .S0(n1449), .Y(n4865) );
  MUX21X1_HVT U367 ( .A1(n3322), .A2(keyout[9]), .S0(n1450), .Y(n4864) );
  MUX21X1_HVT U368 ( .A1(n3321), .A2(keyout[9]), .S0(n1451), .Y(n4863) );
  MUX21X1_HVT U369 ( .A1(n3320), .A2(keyout[9]), .S0(n1452), .Y(n4862) );
  MUX21X1_HVT U370 ( .A1(n3319), .A2(keyout[9]), .S0(n1453), .Y(n4861) );
  MUX21X1_HVT U371 ( .A1(n3318), .A2(keyout[9]), .S0(n1454), .Y(n4860) );
  MUX21X1_HVT U372 ( .A1(n3317), .A2(keyout[10]), .S0(n1447), .Y(n4859) );
  MUX21X1_HVT U373 ( .A1(n3316), .A2(keyout[10]), .S0(n1448), .Y(n4858) );
  MUX21X1_HVT U374 ( .A1(n3315), .A2(keyout[10]), .S0(n1449), .Y(n4857) );
  MUX21X1_HVT U375 ( .A1(n3314), .A2(keyout[10]), .S0(n1450), .Y(n4856) );
  MUX21X1_HVT U376 ( .A1(n3313), .A2(keyout[10]), .S0(n1451), .Y(n4855) );
  MUX21X1_HVT U377 ( .A1(n3312), .A2(keyout[10]), .S0(n1452), .Y(n4854) );
  MUX21X1_HVT U378 ( .A1(n3311), .A2(keyout[10]), .S0(n1453), .Y(n4853) );
  MUX21X1_HVT U379 ( .A1(n3310), .A2(keyout[10]), .S0(n1454), .Y(n4852) );
  MUX21X1_HVT U380 ( .A1(n3309), .A2(keyout[11]), .S0(n1447), .Y(n4851) );
  MUX21X1_HVT U381 ( .A1(n3308), .A2(keyout[11]), .S0(n1448), .Y(n4850) );
  MUX21X1_HVT U382 ( .A1(n3307), .A2(keyout[11]), .S0(n1449), .Y(n4849) );
  MUX21X1_HVT U383 ( .A1(n3306), .A2(keyout[11]), .S0(n1450), .Y(n4848) );
  MUX21X1_HVT U384 ( .A1(n3305), .A2(keyout[11]), .S0(n1451), .Y(n4847) );
  MUX21X1_HVT U385 ( .A1(n3304), .A2(keyout[11]), .S0(n1452), .Y(n4846) );
  MUX21X1_HVT U386 ( .A1(n3303), .A2(keyout[11]), .S0(n1453), .Y(n4845) );
  MUX21X1_HVT U387 ( .A1(n3302), .A2(keyout[11]), .S0(n1454), .Y(n4844) );
  MUX21X1_HVT U388 ( .A1(n3301), .A2(keyout[12]), .S0(n1447), .Y(n4843) );
  MUX21X1_HVT U389 ( .A1(n3300), .A2(keyout[12]), .S0(n1448), .Y(n4842) );
  MUX21X1_HVT U390 ( .A1(n3299), .A2(keyout[12]), .S0(n1449), .Y(n4841) );
  MUX21X1_HVT U391 ( .A1(n3298), .A2(keyout[12]), .S0(n1450), .Y(n4840) );
  MUX21X1_HVT U392 ( .A1(n3297), .A2(keyout[12]), .S0(n1451), .Y(n4839) );
  MUX21X1_HVT U393 ( .A1(n3296), .A2(keyout[12]), .S0(n1452), .Y(n4838) );
  MUX21X1_HVT U394 ( .A1(n3295), .A2(keyout[12]), .S0(n1453), .Y(n4837) );
  MUX21X1_HVT U395 ( .A1(n3294), .A2(keyout[12]), .S0(n1454), .Y(n4836) );
  MUX21X1_HVT U396 ( .A1(n3293), .A2(keyout[13]), .S0(n1447), .Y(n4835) );
  MUX21X1_HVT U397 ( .A1(n3292), .A2(keyout[13]), .S0(n1448), .Y(n4834) );
  MUX21X1_HVT U398 ( .A1(n3291), .A2(keyout[13]), .S0(n1449), .Y(n4833) );
  MUX21X1_HVT U399 ( .A1(n3290), .A2(keyout[13]), .S0(n1450), .Y(n4832) );
  MUX21X1_HVT U400 ( .A1(n3289), .A2(keyout[13]), .S0(n1451), .Y(n4831) );
  MUX21X1_HVT U401 ( .A1(n3288), .A2(keyout[13]), .S0(n1452), .Y(n4830) );
  MUX21X1_HVT U402 ( .A1(n3287), .A2(keyout[13]), .S0(n1453), .Y(n4829) );
  MUX21X1_HVT U403 ( .A1(n3286), .A2(keyout[13]), .S0(n1454), .Y(n4828) );
  MUX21X1_HVT U404 ( .A1(n3285), .A2(keyout[14]), .S0(n1447), .Y(n4827) );
  MUX21X1_HVT U405 ( .A1(n3284), .A2(keyout[14]), .S0(n1448), .Y(n4826) );
  MUX21X1_HVT U406 ( .A1(n3283), .A2(keyout[14]), .S0(n1449), .Y(n4825) );
  MUX21X1_HVT U407 ( .A1(n3282), .A2(keyout[14]), .S0(n1450), .Y(n4824) );
  MUX21X1_HVT U408 ( .A1(n3281), .A2(keyout[14]), .S0(n1451), .Y(n4823) );
  MUX21X1_HVT U409 ( .A1(n3280), .A2(keyout[14]), .S0(n1452), .Y(n4822) );
  MUX21X1_HVT U410 ( .A1(n3279), .A2(keyout[14]), .S0(n1453), .Y(n4821) );
  MUX21X1_HVT U411 ( .A1(n3278), .A2(keyout[14]), .S0(n1454), .Y(n4820) );
  MUX21X1_HVT U412 ( .A1(n3277), .A2(keyout[15]), .S0(n1447), .Y(n4819) );
  MUX21X1_HVT U413 ( .A1(n3276), .A2(keyout[15]), .S0(n1448), .Y(n4818) );
  MUX21X1_HVT U414 ( .A1(n3275), .A2(keyout[15]), .S0(n1449), .Y(n4817) );
  MUX21X1_HVT U415 ( .A1(n3274), .A2(keyout[15]), .S0(n1450), .Y(n4816) );
  MUX21X1_HVT U416 ( .A1(n3273), .A2(keyout[15]), .S0(n1451), .Y(n4815) );
  MUX21X1_HVT U417 ( .A1(n3272), .A2(keyout[15]), .S0(n1452), .Y(n4814) );
  MUX21X1_HVT U418 ( .A1(n3271), .A2(keyout[15]), .S0(n1453), .Y(n4813) );
  MUX21X1_HVT U419 ( .A1(n3270), .A2(keyout[15]), .S0(n1454), .Y(n4812) );
  MUX21X1_HVT U420 ( .A1(n3269), .A2(keyout[16]), .S0(n1447), .Y(n4811) );
  MUX21X1_HVT U421 ( .A1(n3268), .A2(keyout[16]), .S0(n1448), .Y(n4810) );
  MUX21X1_HVT U422 ( .A1(n3267), .A2(keyout[16]), .S0(n1449), .Y(n4809) );
  MUX21X1_HVT U423 ( .A1(n3266), .A2(keyout[16]), .S0(n1450), .Y(n4808) );
  MUX21X1_HVT U424 ( .A1(n3265), .A2(keyout[16]), .S0(n1451), .Y(n4807) );
  MUX21X1_HVT U425 ( .A1(n3264), .A2(keyout[16]), .S0(n1452), .Y(n4806) );
  MUX21X1_HVT U426 ( .A1(n3263), .A2(keyout[16]), .S0(n1453), .Y(n4805) );
  MUX21X1_HVT U427 ( .A1(n3262), .A2(keyout[16]), .S0(n1454), .Y(n4804) );
  MUX21X1_HVT U428 ( .A1(n3261), .A2(keyout[17]), .S0(n1447), .Y(n4803) );
  MUX21X1_HVT U429 ( .A1(n3260), .A2(keyout[17]), .S0(n1448), .Y(n4802) );
  MUX21X1_HVT U430 ( .A1(n3259), .A2(keyout[17]), .S0(n1449), .Y(n4801) );
  MUX21X1_HVT U431 ( .A1(n3258), .A2(keyout[17]), .S0(n1450), .Y(n4800) );
  MUX21X1_HVT U432 ( .A1(n3257), .A2(keyout[17]), .S0(n1451), .Y(n4799) );
  MUX21X1_HVT U433 ( .A1(n3256), .A2(keyout[17]), .S0(n1452), .Y(n4798) );
  MUX21X1_HVT U434 ( .A1(n3255), .A2(keyout[17]), .S0(n1453), .Y(n4797) );
  MUX21X1_HVT U435 ( .A1(n3254), .A2(keyout[17]), .S0(n1454), .Y(n4796) );
  MUX21X1_HVT U436 ( .A1(n3253), .A2(keyout[18]), .S0(n1447), .Y(n4795) );
  MUX21X1_HVT U437 ( .A1(n3252), .A2(keyout[18]), .S0(n1448), .Y(n4794) );
  MUX21X1_HVT U438 ( .A1(n3251), .A2(keyout[18]), .S0(n1449), .Y(n4793) );
  MUX21X1_HVT U439 ( .A1(n3250), .A2(keyout[18]), .S0(n1450), .Y(n4792) );
  MUX21X1_HVT U440 ( .A1(n3249), .A2(keyout[18]), .S0(n1451), .Y(n4791) );
  MUX21X1_HVT U441 ( .A1(n3248), .A2(keyout[18]), .S0(n1452), .Y(n4790) );
  MUX21X1_HVT U442 ( .A1(n3247), .A2(keyout[18]), .S0(n1453), .Y(n4789) );
  MUX21X1_HVT U443 ( .A1(n3246), .A2(keyout[18]), .S0(n1454), .Y(n4788) );
  MUX21X1_HVT U444 ( .A1(n3245), .A2(keyout[19]), .S0(n1447), .Y(n4787) );
  MUX21X1_HVT U445 ( .A1(n3244), .A2(keyout[19]), .S0(n1448), .Y(n4786) );
  MUX21X1_HVT U446 ( .A1(n3243), .A2(keyout[19]), .S0(n1449), .Y(n4785) );
  MUX21X1_HVT U447 ( .A1(n3242), .A2(keyout[19]), .S0(n1450), .Y(n4784) );
  MUX21X1_HVT U448 ( .A1(n3241), .A2(keyout[19]), .S0(n1451), .Y(n4783) );
  MUX21X1_HVT U449 ( .A1(n3240), .A2(keyout[19]), .S0(n1452), .Y(n4782) );
  MUX21X1_HVT U450 ( .A1(n3239), .A2(keyout[19]), .S0(n1453), .Y(n4781) );
  MUX21X1_HVT U451 ( .A1(n3238), .A2(keyout[19]), .S0(n1454), .Y(n4780) );
  MUX21X1_HVT U452 ( .A1(n3237), .A2(keyout[20]), .S0(n1447), .Y(n4779) );
  MUX21X1_HVT U453 ( .A1(n3236), .A2(keyout[20]), .S0(n1448), .Y(n4778) );
  MUX21X1_HVT U454 ( .A1(n3235), .A2(keyout[20]), .S0(n1449), .Y(n4777) );
  MUX21X1_HVT U455 ( .A1(n3234), .A2(keyout[20]), .S0(n1450), .Y(n4776) );
  MUX21X1_HVT U456 ( .A1(n3233), .A2(keyout[20]), .S0(n1451), .Y(n4775) );
  MUX21X1_HVT U457 ( .A1(n3232), .A2(keyout[20]), .S0(n1452), .Y(n4774) );
  MUX21X1_HVT U458 ( .A1(n3231), .A2(keyout[20]), .S0(n1453), .Y(n4773) );
  MUX21X1_HVT U459 ( .A1(n3230), .A2(keyout[20]), .S0(n1454), .Y(n4772) );
  MUX21X1_HVT U460 ( .A1(n3229), .A2(keyout[21]), .S0(n1447), .Y(n4771) );
  MUX21X1_HVT U461 ( .A1(n3228), .A2(keyout[21]), .S0(n1448), .Y(n4770) );
  MUX21X1_HVT U462 ( .A1(n3227), .A2(keyout[21]), .S0(n1449), .Y(n4769) );
  MUX21X1_HVT U463 ( .A1(n3226), .A2(keyout[21]), .S0(n1450), .Y(n4768) );
  MUX21X1_HVT U464 ( .A1(n3225), .A2(keyout[21]), .S0(n1451), .Y(n4767) );
  MUX21X1_HVT U465 ( .A1(n3224), .A2(keyout[21]), .S0(n1452), .Y(n4766) );
  MUX21X1_HVT U466 ( .A1(n3223), .A2(keyout[21]), .S0(n1453), .Y(n4765) );
  MUX21X1_HVT U467 ( .A1(n3222), .A2(keyout[21]), .S0(n1454), .Y(n4764) );
  MUX21X1_HVT U468 ( .A1(n3221), .A2(keyout[22]), .S0(n1447), .Y(n4763) );
  MUX21X1_HVT U469 ( .A1(n3220), .A2(keyout[22]), .S0(n1448), .Y(n4762) );
  MUX21X1_HVT U470 ( .A1(n3219), .A2(keyout[22]), .S0(n1449), .Y(n4761) );
  MUX21X1_HVT U471 ( .A1(n3218), .A2(keyout[22]), .S0(n1450), .Y(n4760) );
  MUX21X1_HVT U472 ( .A1(n3217), .A2(keyout[22]), .S0(n1451), .Y(n4759) );
  MUX21X1_HVT U473 ( .A1(n3216), .A2(keyout[22]), .S0(n1452), .Y(n4758) );
  MUX21X1_HVT U474 ( .A1(n3215), .A2(keyout[22]), .S0(n1453), .Y(n4757) );
  MUX21X1_HVT U475 ( .A1(n3214), .A2(keyout[22]), .S0(n1454), .Y(n4756) );
  MUX21X1_HVT U476 ( .A1(n3213), .A2(keyout[23]), .S0(n1447), .Y(n4755) );
  MUX21X1_HVT U477 ( .A1(n3212), .A2(keyout[23]), .S0(n1448), .Y(n4754) );
  MUX21X1_HVT U478 ( .A1(n3211), .A2(keyout[23]), .S0(n1449), .Y(n4753) );
  MUX21X1_HVT U479 ( .A1(n3210), .A2(keyout[23]), .S0(n1450), .Y(n4752) );
  MUX21X1_HVT U480 ( .A1(n3209), .A2(keyout[23]), .S0(n1451), .Y(n4751) );
  MUX21X1_HVT U481 ( .A1(n3208), .A2(keyout[23]), .S0(n1452), .Y(n4750) );
  MUX21X1_HVT U482 ( .A1(n3207), .A2(keyout[23]), .S0(n1453), .Y(n4749) );
  MUX21X1_HVT U483 ( .A1(n3206), .A2(keyout[23]), .S0(n1454), .Y(n4748) );
  MUX21X1_HVT U484 ( .A1(n3205), .A2(keyout[24]), .S0(n1447), .Y(n4747) );
  MUX21X1_HVT U485 ( .A1(n3204), .A2(keyout[24]), .S0(n1448), .Y(n4746) );
  MUX21X1_HVT U486 ( .A1(n3203), .A2(keyout[24]), .S0(n1449), .Y(n4745) );
  MUX21X1_HVT U487 ( .A1(n3202), .A2(keyout[24]), .S0(n1450), .Y(n4744) );
  MUX21X1_HVT U488 ( .A1(n3201), .A2(keyout[24]), .S0(n1451), .Y(n4743) );
  MUX21X1_HVT U489 ( .A1(n3200), .A2(keyout[24]), .S0(n1452), .Y(n4742) );
  MUX21X1_HVT U490 ( .A1(n3199), .A2(keyout[24]), .S0(n1453), .Y(n4741) );
  MUX21X1_HVT U491 ( .A1(n3198), .A2(keyout[24]), .S0(n1454), .Y(n4740) );
  MUX21X1_HVT U492 ( .A1(n3197), .A2(keyout[25]), .S0(n1447), .Y(n4739) );
  MUX21X1_HVT U493 ( .A1(n3196), .A2(keyout[25]), .S0(n1448), .Y(n4738) );
  MUX21X1_HVT U494 ( .A1(n3195), .A2(keyout[25]), .S0(n1449), .Y(n4737) );
  MUX21X1_HVT U495 ( .A1(n3194), .A2(keyout[25]), .S0(n1450), .Y(n4736) );
  MUX21X1_HVT U496 ( .A1(n3193), .A2(keyout[25]), .S0(n1451), .Y(n4735) );
  MUX21X1_HVT U497 ( .A1(n3192), .A2(keyout[25]), .S0(n1452), .Y(n4734) );
  MUX21X1_HVT U498 ( .A1(n3191), .A2(keyout[25]), .S0(n1453), .Y(n4733) );
  MUX21X1_HVT U499 ( .A1(n3190), .A2(keyout[25]), .S0(n1454), .Y(n4732) );
  MUX21X1_HVT U500 ( .A1(n3189), .A2(keyout[26]), .S0(n1447), .Y(n4731) );
  MUX21X1_HVT U501 ( .A1(n3188), .A2(keyout[26]), .S0(n1448), .Y(n4730) );
  MUX21X1_HVT U502 ( .A1(n3187), .A2(keyout[26]), .S0(n1449), .Y(n4729) );
  MUX21X1_HVT U503 ( .A1(n3186), .A2(keyout[26]), .S0(n1450), .Y(n4728) );
  MUX21X1_HVT U504 ( .A1(n3185), .A2(keyout[26]), .S0(n1451), .Y(n4727) );
  MUX21X1_HVT U505 ( .A1(n3184), .A2(keyout[26]), .S0(n1452), .Y(n4726) );
  MUX21X1_HVT U506 ( .A1(n3183), .A2(keyout[26]), .S0(n1453), .Y(n4725) );
  MUX21X1_HVT U507 ( .A1(n3182), .A2(keyout[26]), .S0(n1454), .Y(n4724) );
  MUX21X1_HVT U508 ( .A1(n3181), .A2(keyout[27]), .S0(n1447), .Y(n4723) );
  MUX21X1_HVT U509 ( .A1(n3180), .A2(keyout[27]), .S0(n1448), .Y(n4722) );
  MUX21X1_HVT U510 ( .A1(n3179), .A2(keyout[27]), .S0(n1449), .Y(n4721) );
  MUX21X1_HVT U511 ( .A1(n3178), .A2(keyout[27]), .S0(n1450), .Y(n4720) );
  MUX21X1_HVT U512 ( .A1(n3177), .A2(keyout[27]), .S0(n1451), .Y(n4719) );
  MUX21X1_HVT U513 ( .A1(n3176), .A2(keyout[27]), .S0(n1452), .Y(n4718) );
  MUX21X1_HVT U514 ( .A1(n3175), .A2(keyout[27]), .S0(n1453), .Y(n4717) );
  MUX21X1_HVT U515 ( .A1(n3174), .A2(keyout[27]), .S0(n1454), .Y(n4716) );
  MUX21X1_HVT U516 ( .A1(n3173), .A2(keyout[28]), .S0(n1447), .Y(n4715) );
  MUX21X1_HVT U517 ( .A1(n3172), .A2(keyout[28]), .S0(n1448), .Y(n4714) );
  MUX21X1_HVT U518 ( .A1(n3171), .A2(keyout[28]), .S0(n1449), .Y(n4713) );
  MUX21X1_HVT U519 ( .A1(n3170), .A2(keyout[28]), .S0(n1450), .Y(n4712) );
  MUX21X1_HVT U520 ( .A1(n3169), .A2(keyout[28]), .S0(n1451), .Y(n4711) );
  MUX21X1_HVT U521 ( .A1(n3168), .A2(keyout[28]), .S0(n1452), .Y(n4710) );
  MUX21X1_HVT U522 ( .A1(n3167), .A2(keyout[28]), .S0(n1453), .Y(n4709) );
  MUX21X1_HVT U523 ( .A1(n3166), .A2(keyout[28]), .S0(n1454), .Y(n4708) );
  MUX21X1_HVT U524 ( .A1(n3165), .A2(keyout[29]), .S0(n1447), .Y(n4707) );
  MUX21X1_HVT U525 ( .A1(n3164), .A2(keyout[29]), .S0(n1448), .Y(n4706) );
  MUX21X1_HVT U526 ( .A1(n3163), .A2(keyout[29]), .S0(n1449), .Y(n4705) );
  MUX21X1_HVT U527 ( .A1(n3162), .A2(keyout[29]), .S0(n1450), .Y(n4704) );
  MUX21X1_HVT U528 ( .A1(n3161), .A2(keyout[29]), .S0(n1451), .Y(n4703) );
  MUX21X1_HVT U529 ( .A1(n3160), .A2(keyout[29]), .S0(n1452), .Y(n4702) );
  MUX21X1_HVT U530 ( .A1(n3159), .A2(keyout[29]), .S0(n1453), .Y(n4701) );
  MUX21X1_HVT U531 ( .A1(n3158), .A2(keyout[29]), .S0(n1454), .Y(n4700) );
  MUX21X1_HVT U532 ( .A1(n3157), .A2(keyout[30]), .S0(n1447), .Y(n4699) );
  MUX21X1_HVT U533 ( .A1(n3156), .A2(keyout[30]), .S0(n1448), .Y(n4698) );
  MUX21X1_HVT U534 ( .A1(n3155), .A2(keyout[30]), .S0(n1449), .Y(n4697) );
  MUX21X1_HVT U535 ( .A1(n3154), .A2(keyout[30]), .S0(n1450), .Y(n4696) );
  MUX21X1_HVT U536 ( .A1(n3153), .A2(keyout[30]), .S0(n1451), .Y(n4695) );
  MUX21X1_HVT U537 ( .A1(n3152), .A2(keyout[30]), .S0(n1452), .Y(n4694) );
  MUX21X1_HVT U538 ( .A1(n3151), .A2(keyout[30]), .S0(n1453), .Y(n4693) );
  MUX21X1_HVT U539 ( .A1(n3150), .A2(keyout[30]), .S0(n1454), .Y(n4692) );
  MUX21X1_HVT U540 ( .A1(n3149), .A2(keyout[31]), .S0(n1447), .Y(n4691) );
  MUX21X1_HVT U541 ( .A1(n3148), .A2(keyout[31]), .S0(n1448), .Y(n4690) );
  MUX21X1_HVT U542 ( .A1(n3147), .A2(keyout[31]), .S0(n1449), .Y(n4689) );
  MUX21X1_HVT U543 ( .A1(n3146), .A2(keyout[31]), .S0(n1450), .Y(n4688) );
  MUX21X1_HVT U544 ( .A1(n3145), .A2(keyout[31]), .S0(n1451), .Y(n4687) );
  MUX21X1_HVT U545 ( .A1(n3144), .A2(keyout[31]), .S0(n1452), .Y(n4686) );
  MUX21X1_HVT U546 ( .A1(n3143), .A2(keyout[31]), .S0(n1453), .Y(n4685) );
  MUX21X1_HVT U547 ( .A1(n3142), .A2(keyout[31]), .S0(n1454), .Y(n4684) );
  MUX21X1_HVT U548 ( .A1(n3141), .A2(keyout[32]), .S0(n1447), .Y(n4683) );
  MUX21X1_HVT U549 ( .A1(n3140), .A2(keyout[32]), .S0(n1448), .Y(n4682) );
  MUX21X1_HVT U550 ( .A1(n3139), .A2(keyout[32]), .S0(n1449), .Y(n4681) );
  MUX21X1_HVT U551 ( .A1(n3138), .A2(keyout[32]), .S0(n1450), .Y(n4680) );
  MUX21X1_HVT U552 ( .A1(n3137), .A2(keyout[32]), .S0(n1451), .Y(n4679) );
  MUX21X1_HVT U553 ( .A1(n3136), .A2(keyout[32]), .S0(n1452), .Y(n4678) );
  MUX21X1_HVT U554 ( .A1(n3135), .A2(keyout[32]), .S0(n1453), .Y(n4677) );
  MUX21X1_HVT U555 ( .A1(n3134), .A2(keyout[32]), .S0(n1454), .Y(n4676) );
  MUX21X1_HVT U556 ( .A1(n3133), .A2(keyout[33]), .S0(n1447), .Y(n4675) );
  MUX21X1_HVT U557 ( .A1(n3132), .A2(keyout[33]), .S0(n1448), .Y(n4674) );
  MUX21X1_HVT U558 ( .A1(n3131), .A2(keyout[33]), .S0(n1449), .Y(n4673) );
  MUX21X1_HVT U559 ( .A1(n3130), .A2(keyout[33]), .S0(n1450), .Y(n4672) );
  MUX21X1_HVT U560 ( .A1(n3129), .A2(keyout[33]), .S0(n1451), .Y(n4671) );
  MUX21X1_HVT U561 ( .A1(n3128), .A2(keyout[33]), .S0(n1452), .Y(n4670) );
  MUX21X1_HVT U562 ( .A1(n3127), .A2(keyout[33]), .S0(n1453), .Y(n4669) );
  MUX21X1_HVT U563 ( .A1(n3126), .A2(keyout[33]), .S0(n1454), .Y(n4668) );
  MUX21X1_HVT U564 ( .A1(n3125), .A2(keyout[34]), .S0(n1447), .Y(n4667) );
  MUX21X1_HVT U565 ( .A1(n3124), .A2(keyout[34]), .S0(n1448), .Y(n4666) );
  MUX21X1_HVT U566 ( .A1(n3123), .A2(keyout[34]), .S0(n1449), .Y(n4665) );
  MUX21X1_HVT U567 ( .A1(n3122), .A2(keyout[34]), .S0(n1450), .Y(n4664) );
  MUX21X1_HVT U568 ( .A1(n3121), .A2(keyout[34]), .S0(n1451), .Y(n4663) );
  MUX21X1_HVT U569 ( .A1(n3120), .A2(keyout[34]), .S0(n1452), .Y(n4662) );
  MUX21X1_HVT U570 ( .A1(n3119), .A2(keyout[34]), .S0(n1453), .Y(n4661) );
  MUX21X1_HVT U571 ( .A1(n3118), .A2(keyout[34]), .S0(n1454), .Y(n4660) );
  MUX21X1_HVT U572 ( .A1(n3117), .A2(keyout[35]), .S0(n1447), .Y(n4659) );
  MUX21X1_HVT U573 ( .A1(n3116), .A2(keyout[35]), .S0(n1448), .Y(n4658) );
  MUX21X1_HVT U574 ( .A1(n3115), .A2(keyout[35]), .S0(n1449), .Y(n4657) );
  MUX21X1_HVT U575 ( .A1(n3114), .A2(keyout[35]), .S0(n1450), .Y(n4656) );
  MUX21X1_HVT U576 ( .A1(n3113), .A2(keyout[35]), .S0(n1451), .Y(n4655) );
  MUX21X1_HVT U577 ( .A1(n3112), .A2(keyout[35]), .S0(n1452), .Y(n4654) );
  MUX21X1_HVT U578 ( .A1(n3111), .A2(keyout[35]), .S0(n1453), .Y(n4653) );
  MUX21X1_HVT U579 ( .A1(n3110), .A2(keyout[35]), .S0(n1454), .Y(n4652) );
  MUX21X1_HVT U580 ( .A1(n3109), .A2(keyout[36]), .S0(n1447), .Y(n4651) );
  MUX21X1_HVT U581 ( .A1(n3108), .A2(keyout[36]), .S0(n1448), .Y(n4650) );
  MUX21X1_HVT U582 ( .A1(n3107), .A2(keyout[36]), .S0(n1449), .Y(n4649) );
  MUX21X1_HVT U583 ( .A1(n3106), .A2(keyout[36]), .S0(n1450), .Y(n4648) );
  MUX21X1_HVT U584 ( .A1(n3105), .A2(keyout[36]), .S0(n1451), .Y(n4647) );
  MUX21X1_HVT U585 ( .A1(n3104), .A2(keyout[36]), .S0(n1452), .Y(n4646) );
  MUX21X1_HVT U586 ( .A1(n3103), .A2(keyout[36]), .S0(n1453), .Y(n4645) );
  MUX21X1_HVT U587 ( .A1(n3102), .A2(keyout[36]), .S0(n1454), .Y(n4644) );
  MUX21X1_HVT U588 ( .A1(n3101), .A2(keyout[37]), .S0(n1447), .Y(n4643) );
  MUX21X1_HVT U589 ( .A1(n3100), .A2(keyout[37]), .S0(n1448), .Y(n4642) );
  MUX21X1_HVT U590 ( .A1(n3099), .A2(keyout[37]), .S0(n1449), .Y(n4641) );
  MUX21X1_HVT U591 ( .A1(n3098), .A2(keyout[37]), .S0(n1450), .Y(n4640) );
  MUX21X1_HVT U592 ( .A1(n3097), .A2(keyout[37]), .S0(n1451), .Y(n4639) );
  MUX21X1_HVT U593 ( .A1(n3096), .A2(keyout[37]), .S0(n1452), .Y(n4638) );
  MUX21X1_HVT U594 ( .A1(n3095), .A2(keyout[37]), .S0(n1453), .Y(n4637) );
  MUX21X1_HVT U595 ( .A1(n3094), .A2(keyout[37]), .S0(n1454), .Y(n4636) );
  MUX21X1_HVT U596 ( .A1(n3093), .A2(keyout[38]), .S0(n1447), .Y(n4635) );
  MUX21X1_HVT U597 ( .A1(n3092), .A2(keyout[38]), .S0(n1448), .Y(n4634) );
  MUX21X1_HVT U598 ( .A1(n3091), .A2(keyout[38]), .S0(n1449), .Y(n4633) );
  MUX21X1_HVT U599 ( .A1(n3090), .A2(keyout[38]), .S0(n1450), .Y(n4632) );
  MUX21X1_HVT U600 ( .A1(n3089), .A2(keyout[38]), .S0(n1451), .Y(n4631) );
  MUX21X1_HVT U601 ( .A1(n3088), .A2(keyout[38]), .S0(n1452), .Y(n4630) );
  MUX21X1_HVT U602 ( .A1(n3087), .A2(keyout[38]), .S0(n1453), .Y(n4629) );
  MUX21X1_HVT U603 ( .A1(n3086), .A2(keyout[38]), .S0(n1454), .Y(n4628) );
  MUX21X1_HVT U604 ( .A1(n3085), .A2(keyout[39]), .S0(n1447), .Y(n4627) );
  MUX21X1_HVT U605 ( .A1(n3084), .A2(keyout[39]), .S0(n1448), .Y(n4626) );
  MUX21X1_HVT U606 ( .A1(n3083), .A2(keyout[39]), .S0(n1449), .Y(n4625) );
  MUX21X1_HVT U607 ( .A1(n3082), .A2(keyout[39]), .S0(n1450), .Y(n4624) );
  MUX21X1_HVT U608 ( .A1(n3081), .A2(keyout[39]), .S0(n1451), .Y(n4623) );
  MUX21X1_HVT U609 ( .A1(n3080), .A2(keyout[39]), .S0(n1452), .Y(n4622) );
  MUX21X1_HVT U610 ( .A1(n3079), .A2(keyout[39]), .S0(n1453), .Y(n4621) );
  MUX21X1_HVT U611 ( .A1(n3078), .A2(keyout[39]), .S0(n1454), .Y(n4620) );
  MUX21X1_HVT U612 ( .A1(n3077), .A2(keyout[40]), .S0(n1447), .Y(n4619) );
  MUX21X1_HVT U613 ( .A1(n3076), .A2(keyout[40]), .S0(n1448), .Y(n4618) );
  MUX21X1_HVT U614 ( .A1(n3075), .A2(keyout[40]), .S0(n1449), .Y(n4617) );
  MUX21X1_HVT U615 ( .A1(n3074), .A2(keyout[40]), .S0(n1450), .Y(n4616) );
  MUX21X1_HVT U616 ( .A1(n3073), .A2(keyout[40]), .S0(n1451), .Y(n4615) );
  MUX21X1_HVT U617 ( .A1(n3072), .A2(keyout[40]), .S0(n1452), .Y(n4614) );
  MUX21X1_HVT U618 ( .A1(n3071), .A2(keyout[40]), .S0(n1453), .Y(n4613) );
  MUX21X1_HVT U619 ( .A1(n3070), .A2(keyout[40]), .S0(n1454), .Y(n4612) );
  MUX21X1_HVT U620 ( .A1(n3069), .A2(keyout[41]), .S0(n1447), .Y(n4611) );
  MUX21X1_HVT U621 ( .A1(n3068), .A2(keyout[41]), .S0(n1448), .Y(n4610) );
  MUX21X1_HVT U622 ( .A1(n3067), .A2(keyout[41]), .S0(n1449), .Y(n4609) );
  MUX21X1_HVT U623 ( .A1(n3066), .A2(keyout[41]), .S0(n1450), .Y(n4608) );
  MUX21X1_HVT U624 ( .A1(n3065), .A2(keyout[41]), .S0(n1451), .Y(n4607) );
  MUX21X1_HVT U625 ( .A1(n3064), .A2(keyout[41]), .S0(n1452), .Y(n4606) );
  MUX21X1_HVT U626 ( .A1(n3063), .A2(keyout[41]), .S0(n1453), .Y(n4605) );
  MUX21X1_HVT U627 ( .A1(n3062), .A2(keyout[41]), .S0(n1454), .Y(n4604) );
  MUX21X1_HVT U628 ( .A1(n3061), .A2(keyout[42]), .S0(n1447), .Y(n4603) );
  MUX21X1_HVT U629 ( .A1(n3060), .A2(keyout[42]), .S0(n1448), .Y(n4602) );
  MUX21X1_HVT U630 ( .A1(n3059), .A2(keyout[42]), .S0(n1449), .Y(n4601) );
  MUX21X1_HVT U631 ( .A1(n3058), .A2(keyout[42]), .S0(n1450), .Y(n4600) );
  MUX21X1_HVT U632 ( .A1(n3057), .A2(keyout[42]), .S0(n1451), .Y(n4599) );
  MUX21X1_HVT U633 ( .A1(n3056), .A2(keyout[42]), .S0(n1452), .Y(n4598) );
  MUX21X1_HVT U634 ( .A1(n3055), .A2(keyout[42]), .S0(n1453), .Y(n4597) );
  MUX21X1_HVT U635 ( .A1(n3054), .A2(keyout[42]), .S0(n1454), .Y(n4596) );
  MUX21X1_HVT U636 ( .A1(n3053), .A2(keyout[43]), .S0(n1447), .Y(n4595) );
  MUX21X1_HVT U637 ( .A1(n3052), .A2(keyout[43]), .S0(n1448), .Y(n4594) );
  MUX21X1_HVT U638 ( .A1(n3051), .A2(keyout[43]), .S0(n1449), .Y(n4593) );
  MUX21X1_HVT U639 ( .A1(n3050), .A2(keyout[43]), .S0(n1450), .Y(n4592) );
  MUX21X1_HVT U640 ( .A1(n3049), .A2(keyout[43]), .S0(n1451), .Y(n4591) );
  MUX21X1_HVT U641 ( .A1(n3048), .A2(keyout[43]), .S0(n1452), .Y(n4590) );
  MUX21X1_HVT U642 ( .A1(n3047), .A2(keyout[43]), .S0(n1453), .Y(n4589) );
  MUX21X1_HVT U643 ( .A1(n3046), .A2(keyout[43]), .S0(n1454), .Y(n4588) );
  MUX21X1_HVT U644 ( .A1(n3045), .A2(keyout[44]), .S0(n1447), .Y(n4587) );
  MUX21X1_HVT U645 ( .A1(n3044), .A2(keyout[44]), .S0(n1448), .Y(n4586) );
  MUX21X1_HVT U646 ( .A1(n3043), .A2(keyout[44]), .S0(n1449), .Y(n4585) );
  MUX21X1_HVT U647 ( .A1(n3042), .A2(keyout[44]), .S0(n1450), .Y(n4584) );
  MUX21X1_HVT U648 ( .A1(n3041), .A2(keyout[44]), .S0(n1451), .Y(n4583) );
  MUX21X1_HVT U649 ( .A1(n3040), .A2(keyout[44]), .S0(n1452), .Y(n4582) );
  MUX21X1_HVT U650 ( .A1(n3039), .A2(keyout[44]), .S0(n1453), .Y(n4581) );
  MUX21X1_HVT U651 ( .A1(n3038), .A2(keyout[44]), .S0(n1454), .Y(n4580) );
  MUX21X1_HVT U652 ( .A1(n3037), .A2(keyout[45]), .S0(n1447), .Y(n4579) );
  MUX21X1_HVT U653 ( .A1(n3036), .A2(keyout[45]), .S0(n1448), .Y(n4578) );
  MUX21X1_HVT U654 ( .A1(n3035), .A2(keyout[45]), .S0(n1449), .Y(n4577) );
  MUX21X1_HVT U655 ( .A1(n3034), .A2(keyout[45]), .S0(n1450), .Y(n4576) );
  MUX21X1_HVT U656 ( .A1(n3033), .A2(keyout[45]), .S0(n1451), .Y(n4575) );
  MUX21X1_HVT U657 ( .A1(n3032), .A2(keyout[45]), .S0(n1452), .Y(n4574) );
  MUX21X1_HVT U658 ( .A1(n3031), .A2(keyout[45]), .S0(n1453), .Y(n4573) );
  MUX21X1_HVT U659 ( .A1(n3030), .A2(keyout[45]), .S0(n1454), .Y(n4572) );
  MUX21X1_HVT U660 ( .A1(n3029), .A2(keyout[46]), .S0(n1447), .Y(n4571) );
  MUX21X1_HVT U661 ( .A1(n3028), .A2(keyout[46]), .S0(n1448), .Y(n4570) );
  MUX21X1_HVT U662 ( .A1(n3027), .A2(keyout[46]), .S0(n1449), .Y(n4569) );
  MUX21X1_HVT U663 ( .A1(n3026), .A2(keyout[46]), .S0(n1450), .Y(n4568) );
  MUX21X1_HVT U664 ( .A1(n3025), .A2(keyout[46]), .S0(n1451), .Y(n4567) );
  MUX21X1_HVT U665 ( .A1(n3024), .A2(keyout[46]), .S0(n1452), .Y(n4566) );
  MUX21X1_HVT U666 ( .A1(n3023), .A2(keyout[46]), .S0(n1453), .Y(n4565) );
  MUX21X1_HVT U667 ( .A1(n3022), .A2(keyout[46]), .S0(n1454), .Y(n4564) );
  MUX21X1_HVT U668 ( .A1(n3021), .A2(keyout[47]), .S0(n1447), .Y(n4563) );
  MUX21X1_HVT U669 ( .A1(n3020), .A2(keyout[47]), .S0(n1448), .Y(n4562) );
  MUX21X1_HVT U670 ( .A1(n3019), .A2(keyout[47]), .S0(n1449), .Y(n4561) );
  MUX21X1_HVT U671 ( .A1(n3018), .A2(keyout[47]), .S0(n1450), .Y(n4560) );
  MUX21X1_HVT U672 ( .A1(n3017), .A2(keyout[47]), .S0(n1451), .Y(n4559) );
  MUX21X1_HVT U673 ( .A1(n3016), .A2(keyout[47]), .S0(n1452), .Y(n4558) );
  MUX21X1_HVT U674 ( .A1(n3015), .A2(keyout[47]), .S0(n1453), .Y(n4557) );
  MUX21X1_HVT U675 ( .A1(n3014), .A2(keyout[47]), .S0(n1454), .Y(n4556) );
  MUX21X1_HVT U676 ( .A1(n3013), .A2(keyout[48]), .S0(n1447), .Y(n4555) );
  MUX21X1_HVT U677 ( .A1(n3012), .A2(keyout[48]), .S0(n1448), .Y(n4554) );
  MUX21X1_HVT U678 ( .A1(n3011), .A2(keyout[48]), .S0(n1449), .Y(n4553) );
  MUX21X1_HVT U679 ( .A1(n3010), .A2(keyout[48]), .S0(n1450), .Y(n4552) );
  MUX21X1_HVT U680 ( .A1(n3009), .A2(keyout[48]), .S0(n1451), .Y(n4551) );
  MUX21X1_HVT U681 ( .A1(n3008), .A2(keyout[48]), .S0(n1452), .Y(n4550) );
  MUX21X1_HVT U682 ( .A1(n3007), .A2(keyout[48]), .S0(n1453), .Y(n4549) );
  MUX21X1_HVT U683 ( .A1(n3006), .A2(keyout[48]), .S0(n1454), .Y(n4548) );
  MUX21X1_HVT U684 ( .A1(n3005), .A2(keyout[49]), .S0(n1447), .Y(n4547) );
  MUX21X1_HVT U685 ( .A1(n3004), .A2(keyout[49]), .S0(n1448), .Y(n4546) );
  MUX21X1_HVT U686 ( .A1(n3003), .A2(keyout[49]), .S0(n1449), .Y(n4545) );
  MUX21X1_HVT U687 ( .A1(n3002), .A2(keyout[49]), .S0(n1450), .Y(n4544) );
  MUX21X1_HVT U688 ( .A1(n3001), .A2(keyout[49]), .S0(n1451), .Y(n4543) );
  MUX21X1_HVT U689 ( .A1(n3000), .A2(keyout[49]), .S0(n1452), .Y(n4542) );
  MUX21X1_HVT U690 ( .A1(n2999), .A2(keyout[49]), .S0(n1453), .Y(n4541) );
  MUX21X1_HVT U691 ( .A1(n2998), .A2(keyout[49]), .S0(n1454), .Y(n4540) );
  MUX21X1_HVT U692 ( .A1(n2997), .A2(keyout[50]), .S0(n1447), .Y(n4539) );
  MUX21X1_HVT U693 ( .A1(n2996), .A2(keyout[50]), .S0(n1448), .Y(n4538) );
  MUX21X1_HVT U694 ( .A1(n2995), .A2(keyout[50]), .S0(n1449), .Y(n4537) );
  MUX21X1_HVT U695 ( .A1(n2994), .A2(keyout[50]), .S0(n1450), .Y(n4536) );
  MUX21X1_HVT U696 ( .A1(n2993), .A2(keyout[50]), .S0(n1451), .Y(n4535) );
  MUX21X1_HVT U697 ( .A1(n2992), .A2(keyout[50]), .S0(n1452), .Y(n4534) );
  MUX21X1_HVT U698 ( .A1(n2991), .A2(keyout[50]), .S0(n1453), .Y(n4533) );
  MUX21X1_HVT U699 ( .A1(n2990), .A2(keyout[50]), .S0(n1454), .Y(n4532) );
  MUX21X1_HVT U700 ( .A1(n2989), .A2(keyout[51]), .S0(n1447), .Y(n4531) );
  MUX21X1_HVT U701 ( .A1(n2988), .A2(keyout[51]), .S0(n1448), .Y(n4530) );
  MUX21X1_HVT U702 ( .A1(n2987), .A2(keyout[51]), .S0(n1449), .Y(n4529) );
  MUX21X1_HVT U703 ( .A1(n2986), .A2(keyout[51]), .S0(n1450), .Y(n4528) );
  MUX21X1_HVT U704 ( .A1(n2985), .A2(keyout[51]), .S0(n1451), .Y(n4527) );
  MUX21X1_HVT U705 ( .A1(n2984), .A2(keyout[51]), .S0(n1452), .Y(n4526) );
  MUX21X1_HVT U706 ( .A1(n2983), .A2(keyout[51]), .S0(n1453), .Y(n4525) );
  MUX21X1_HVT U707 ( .A1(n2982), .A2(keyout[51]), .S0(n1454), .Y(n4524) );
  MUX21X1_HVT U708 ( .A1(n2981), .A2(keyout[52]), .S0(n1447), .Y(n4523) );
  MUX21X1_HVT U709 ( .A1(n2980), .A2(keyout[52]), .S0(n1448), .Y(n4522) );
  MUX21X1_HVT U710 ( .A1(n2979), .A2(keyout[52]), .S0(n1449), .Y(n4521) );
  MUX21X1_HVT U711 ( .A1(n2978), .A2(keyout[52]), .S0(n1450), .Y(n4520) );
  MUX21X1_HVT U712 ( .A1(n2977), .A2(keyout[52]), .S0(n1451), .Y(n4519) );
  MUX21X1_HVT U713 ( .A1(n2976), .A2(keyout[52]), .S0(n1452), .Y(n4518) );
  MUX21X1_HVT U714 ( .A1(n2975), .A2(keyout[52]), .S0(n1453), .Y(n4517) );
  MUX21X1_HVT U715 ( .A1(n2974), .A2(keyout[52]), .S0(n1454), .Y(n4516) );
  MUX21X1_HVT U716 ( .A1(n2973), .A2(keyout[53]), .S0(n1447), .Y(n4515) );
  MUX21X1_HVT U717 ( .A1(n2972), .A2(keyout[53]), .S0(n1448), .Y(n4514) );
  MUX21X1_HVT U718 ( .A1(n2971), .A2(keyout[53]), .S0(n1449), .Y(n4513) );
  MUX21X1_HVT U719 ( .A1(n2970), .A2(keyout[53]), .S0(n1450), .Y(n4512) );
  MUX21X1_HVT U720 ( .A1(n2969), .A2(keyout[53]), .S0(n1451), .Y(n4511) );
  MUX21X1_HVT U721 ( .A1(n2968), .A2(keyout[53]), .S0(n1452), .Y(n4510) );
  MUX21X1_HVT U722 ( .A1(n2967), .A2(keyout[53]), .S0(n1453), .Y(n4509) );
  MUX21X1_HVT U723 ( .A1(n2966), .A2(keyout[53]), .S0(n1454), .Y(n4508) );
  MUX21X1_HVT U724 ( .A1(n2965), .A2(keyout[54]), .S0(n1447), .Y(n4507) );
  MUX21X1_HVT U725 ( .A1(n2964), .A2(keyout[54]), .S0(n1448), .Y(n4506) );
  MUX21X1_HVT U726 ( .A1(n2963), .A2(keyout[54]), .S0(n1449), .Y(n4505) );
  MUX21X1_HVT U727 ( .A1(n2962), .A2(keyout[54]), .S0(n1450), .Y(n4504) );
  MUX21X1_HVT U728 ( .A1(n2961), .A2(keyout[54]), .S0(n1451), .Y(n4503) );
  MUX21X1_HVT U729 ( .A1(n2960), .A2(keyout[54]), .S0(n1452), .Y(n4502) );
  MUX21X1_HVT U730 ( .A1(n2959), .A2(keyout[54]), .S0(n1453), .Y(n4501) );
  MUX21X1_HVT U731 ( .A1(n2958), .A2(keyout[54]), .S0(n1454), .Y(n4500) );
  MUX21X1_HVT U732 ( .A1(n2957), .A2(keyout[55]), .S0(n1447), .Y(n4499) );
  MUX21X1_HVT U733 ( .A1(n2956), .A2(keyout[55]), .S0(n1448), .Y(n4498) );
  MUX21X1_HVT U734 ( .A1(n2955), .A2(keyout[55]), .S0(n1449), .Y(n4497) );
  MUX21X1_HVT U735 ( .A1(n2954), .A2(keyout[55]), .S0(n1450), .Y(n4496) );
  MUX21X1_HVT U736 ( .A1(n2953), .A2(keyout[55]), .S0(n1451), .Y(n4495) );
  MUX21X1_HVT U737 ( .A1(n2952), .A2(keyout[55]), .S0(n1452), .Y(n4494) );
  MUX21X1_HVT U738 ( .A1(n2951), .A2(keyout[55]), .S0(n1453), .Y(n4493) );
  MUX21X1_HVT U739 ( .A1(n2950), .A2(keyout[55]), .S0(n1454), .Y(n4492) );
  MUX21X1_HVT U740 ( .A1(n2949), .A2(keyout[56]), .S0(n1447), .Y(n4491) );
  MUX21X1_HVT U741 ( .A1(n2948), .A2(keyout[56]), .S0(n1448), .Y(n4490) );
  MUX21X1_HVT U742 ( .A1(n2947), .A2(keyout[56]), .S0(n1449), .Y(n4489) );
  MUX21X1_HVT U743 ( .A1(n2946), .A2(keyout[56]), .S0(n1450), .Y(n4488) );
  MUX21X1_HVT U744 ( .A1(n2945), .A2(keyout[56]), .S0(n1451), .Y(n4487) );
  MUX21X1_HVT U745 ( .A1(n2944), .A2(keyout[56]), .S0(n1452), .Y(n4486) );
  MUX21X1_HVT U746 ( .A1(n2943), .A2(keyout[56]), .S0(n1453), .Y(n4485) );
  MUX21X1_HVT U747 ( .A1(n2942), .A2(keyout[56]), .S0(n1454), .Y(n4484) );
  MUX21X1_HVT U748 ( .A1(n2941), .A2(keyout[57]), .S0(n1447), .Y(n4483) );
  MUX21X1_HVT U749 ( .A1(n2940), .A2(keyout[57]), .S0(n1448), .Y(n4482) );
  MUX21X1_HVT U750 ( .A1(n2939), .A2(keyout[57]), .S0(n1449), .Y(n4481) );
  MUX21X1_HVT U751 ( .A1(n2938), .A2(keyout[57]), .S0(n1450), .Y(n4480) );
  MUX21X1_HVT U752 ( .A1(n2937), .A2(keyout[57]), .S0(n1451), .Y(n4479) );
  MUX21X1_HVT U753 ( .A1(n2936), .A2(keyout[57]), .S0(n1452), .Y(n4478) );
  MUX21X1_HVT U754 ( .A1(n2935), .A2(keyout[57]), .S0(n1453), .Y(n4477) );
  MUX21X1_HVT U755 ( .A1(n2934), .A2(keyout[57]), .S0(n1454), .Y(n4476) );
  MUX21X1_HVT U756 ( .A1(n2933), .A2(keyout[58]), .S0(n1447), .Y(n4475) );
  MUX21X1_HVT U757 ( .A1(n2932), .A2(keyout[58]), .S0(n1448), .Y(n4474) );
  MUX21X1_HVT U758 ( .A1(n2931), .A2(keyout[58]), .S0(n1449), .Y(n4473) );
  MUX21X1_HVT U759 ( .A1(n2930), .A2(keyout[58]), .S0(n1450), .Y(n4472) );
  MUX21X1_HVT U760 ( .A1(n2929), .A2(keyout[58]), .S0(n1451), .Y(n4471) );
  MUX21X1_HVT U761 ( .A1(n2928), .A2(keyout[58]), .S0(n1452), .Y(n4470) );
  MUX21X1_HVT U762 ( .A1(n2927), .A2(keyout[58]), .S0(n1453), .Y(n4469) );
  MUX21X1_HVT U763 ( .A1(n2926), .A2(keyout[58]), .S0(n1454), .Y(n4468) );
  MUX21X1_HVT U764 ( .A1(n2925), .A2(keyout[59]), .S0(n1447), .Y(n4467) );
  MUX21X1_HVT U765 ( .A1(n2924), .A2(keyout[59]), .S0(n1448), .Y(n4466) );
  MUX21X1_HVT U766 ( .A1(n2923), .A2(keyout[59]), .S0(n1449), .Y(n4465) );
  MUX21X1_HVT U767 ( .A1(n2922), .A2(keyout[59]), .S0(n1450), .Y(n4464) );
  MUX21X1_HVT U768 ( .A1(n2921), .A2(keyout[59]), .S0(n1451), .Y(n4463) );
  MUX21X1_HVT U769 ( .A1(n2920), .A2(keyout[59]), .S0(n1452), .Y(n4462) );
  MUX21X1_HVT U770 ( .A1(n2919), .A2(keyout[59]), .S0(n1453), .Y(n4461) );
  MUX21X1_HVT U771 ( .A1(n2918), .A2(keyout[59]), .S0(n1454), .Y(n4460) );
  MUX21X1_HVT U772 ( .A1(n2917), .A2(keyout[60]), .S0(n1447), .Y(n4459) );
  MUX21X1_HVT U773 ( .A1(n2916), .A2(keyout[60]), .S0(n1448), .Y(n4458) );
  MUX21X1_HVT U774 ( .A1(n2915), .A2(keyout[60]), .S0(n1449), .Y(n4457) );
  MUX21X1_HVT U775 ( .A1(n2914), .A2(keyout[60]), .S0(n1450), .Y(n4456) );
  MUX21X1_HVT U776 ( .A1(n2913), .A2(keyout[60]), .S0(n1451), .Y(n4455) );
  MUX21X1_HVT U777 ( .A1(n2912), .A2(keyout[60]), .S0(n1452), .Y(n4454) );
  MUX21X1_HVT U778 ( .A1(n2911), .A2(keyout[60]), .S0(n1453), .Y(n4453) );
  MUX21X1_HVT U779 ( .A1(n2910), .A2(keyout[60]), .S0(n1454), .Y(n4452) );
  MUX21X1_HVT U780 ( .A1(n2909), .A2(keyout[61]), .S0(n1447), .Y(n4451) );
  MUX21X1_HVT U781 ( .A1(n2908), .A2(keyout[61]), .S0(n1448), .Y(n4450) );
  MUX21X1_HVT U782 ( .A1(n2907), .A2(keyout[61]), .S0(n1449), .Y(n4449) );
  MUX21X1_HVT U783 ( .A1(n2906), .A2(keyout[61]), .S0(n1450), .Y(n4448) );
  MUX21X1_HVT U784 ( .A1(n2905), .A2(keyout[61]), .S0(n1451), .Y(n4447) );
  MUX21X1_HVT U785 ( .A1(n2904), .A2(keyout[61]), .S0(n1452), .Y(n4446) );
  MUX21X1_HVT U786 ( .A1(n2903), .A2(keyout[61]), .S0(n1453), .Y(n4445) );
  MUX21X1_HVT U787 ( .A1(n2902), .A2(keyout[61]), .S0(n1454), .Y(n4444) );
  MUX21X1_HVT U788 ( .A1(n2901), .A2(keyout[62]), .S0(n1447), .Y(n4443) );
  MUX21X1_HVT U789 ( .A1(n2900), .A2(keyout[62]), .S0(n1448), .Y(n4442) );
  MUX21X1_HVT U790 ( .A1(n2899), .A2(keyout[62]), .S0(n1449), .Y(n4441) );
  MUX21X1_HVT U791 ( .A1(n2898), .A2(keyout[62]), .S0(n1450), .Y(n4440) );
  MUX21X1_HVT U792 ( .A1(n2897), .A2(keyout[62]), .S0(n1451), .Y(n4439) );
  MUX21X1_HVT U793 ( .A1(n2896), .A2(keyout[62]), .S0(n1452), .Y(n4438) );
  MUX21X1_HVT U794 ( .A1(n2895), .A2(keyout[62]), .S0(n1453), .Y(n4437) );
  MUX21X1_HVT U795 ( .A1(n2894), .A2(keyout[62]), .S0(n1454), .Y(n4436) );
  MUX21X1_HVT U796 ( .A1(n2893), .A2(keyout[63]), .S0(n1447), .Y(n4435) );
  MUX21X1_HVT U797 ( .A1(n2892), .A2(keyout[63]), .S0(n1448), .Y(n4434) );
  MUX21X1_HVT U798 ( .A1(n2891), .A2(keyout[63]), .S0(n1449), .Y(n4433) );
  MUX21X1_HVT U799 ( .A1(n2890), .A2(keyout[63]), .S0(n1450), .Y(n4432) );
  MUX21X1_HVT U800 ( .A1(n2889), .A2(keyout[63]), .S0(n1451), .Y(n4431) );
  MUX21X1_HVT U801 ( .A1(n2888), .A2(keyout[63]), .S0(n1452), .Y(n4430) );
  MUX21X1_HVT U802 ( .A1(n2887), .A2(keyout[63]), .S0(n1453), .Y(n4429) );
  MUX21X1_HVT U803 ( .A1(n2886), .A2(keyout[63]), .S0(n1454), .Y(n4428) );
  MUX21X1_HVT U804 ( .A1(n2885), .A2(keyout[64]), .S0(n1447), .Y(n4427) );
  MUX21X1_HVT U805 ( .A1(n2884), .A2(keyout[64]), .S0(n1448), .Y(n4426) );
  MUX21X1_HVT U806 ( .A1(n2883), .A2(keyout[64]), .S0(n1449), .Y(n4425) );
  MUX21X1_HVT U807 ( .A1(n2882), .A2(keyout[64]), .S0(n1450), .Y(n4424) );
  MUX21X1_HVT U808 ( .A1(n2881), .A2(keyout[64]), .S0(n1451), .Y(n4423) );
  MUX21X1_HVT U809 ( .A1(n2880), .A2(keyout[64]), .S0(n1452), .Y(n4422) );
  MUX21X1_HVT U810 ( .A1(n2879), .A2(keyout[64]), .S0(n1453), .Y(n4421) );
  MUX21X1_HVT U811 ( .A1(n2878), .A2(keyout[64]), .S0(n1454), .Y(n4420) );
  MUX21X1_HVT U812 ( .A1(n2877), .A2(keyout[65]), .S0(n1447), .Y(n4419) );
  MUX21X1_HVT U813 ( .A1(n2876), .A2(keyout[65]), .S0(n1448), .Y(n4418) );
  MUX21X1_HVT U814 ( .A1(n2875), .A2(keyout[65]), .S0(n1449), .Y(n4417) );
  MUX21X1_HVT U815 ( .A1(n2874), .A2(keyout[65]), .S0(n1450), .Y(n4416) );
  MUX21X1_HVT U816 ( .A1(n2873), .A2(keyout[65]), .S0(n1451), .Y(n4415) );
  MUX21X1_HVT U817 ( .A1(n2872), .A2(keyout[65]), .S0(n1452), .Y(n4414) );
  MUX21X1_HVT U818 ( .A1(n2871), .A2(keyout[65]), .S0(n1453), .Y(n4413) );
  MUX21X1_HVT U819 ( .A1(n2870), .A2(keyout[65]), .S0(n1454), .Y(n4412) );
  MUX21X1_HVT U820 ( .A1(n2869), .A2(keyout[66]), .S0(n1447), .Y(n4411) );
  MUX21X1_HVT U821 ( .A1(n2868), .A2(keyout[66]), .S0(n1448), .Y(n4410) );
  MUX21X1_HVT U822 ( .A1(n2867), .A2(keyout[66]), .S0(n1449), .Y(n4409) );
  MUX21X1_HVT U823 ( .A1(n2866), .A2(keyout[66]), .S0(n1450), .Y(n4408) );
  MUX21X1_HVT U824 ( .A1(n2865), .A2(keyout[66]), .S0(n1451), .Y(n4407) );
  MUX21X1_HVT U825 ( .A1(n2864), .A2(keyout[66]), .S0(n1452), .Y(n4406) );
  MUX21X1_HVT U826 ( .A1(n2863), .A2(keyout[66]), .S0(n1453), .Y(n4405) );
  MUX21X1_HVT U827 ( .A1(n2862), .A2(keyout[66]), .S0(n1454), .Y(n4404) );
  MUX21X1_HVT U828 ( .A1(n2861), .A2(keyout[67]), .S0(n1447), .Y(n4403) );
  MUX21X1_HVT U829 ( .A1(n2860), .A2(keyout[67]), .S0(n1448), .Y(n4402) );
  MUX21X1_HVT U830 ( .A1(n2859), .A2(keyout[67]), .S0(n1449), .Y(n4401) );
  MUX21X1_HVT U831 ( .A1(n2858), .A2(keyout[67]), .S0(n1450), .Y(n4400) );
  MUX21X1_HVT U832 ( .A1(n2857), .A2(keyout[67]), .S0(n1451), .Y(n4399) );
  MUX21X1_HVT U833 ( .A1(n2856), .A2(keyout[67]), .S0(n1452), .Y(n4398) );
  MUX21X1_HVT U834 ( .A1(n2855), .A2(keyout[67]), .S0(n1453), .Y(n4397) );
  MUX21X1_HVT U835 ( .A1(n2854), .A2(keyout[67]), .S0(n1454), .Y(n4396) );
  MUX21X1_HVT U836 ( .A1(n2853), .A2(keyout[68]), .S0(n1447), .Y(n4395) );
  MUX21X1_HVT U837 ( .A1(n2852), .A2(keyout[68]), .S0(n1448), .Y(n4394) );
  MUX21X1_HVT U838 ( .A1(n2851), .A2(keyout[68]), .S0(n1449), .Y(n4393) );
  MUX21X1_HVT U839 ( .A1(n2850), .A2(keyout[68]), .S0(n1450), .Y(n4392) );
  MUX21X1_HVT U840 ( .A1(n2849), .A2(keyout[68]), .S0(n1451), .Y(n4391) );
  MUX21X1_HVT U841 ( .A1(n2848), .A2(keyout[68]), .S0(n1452), .Y(n4390) );
  MUX21X1_HVT U842 ( .A1(n2847), .A2(keyout[68]), .S0(n1453), .Y(n4389) );
  MUX21X1_HVT U843 ( .A1(n2846), .A2(keyout[68]), .S0(n1454), .Y(n4388) );
  MUX21X1_HVT U844 ( .A1(n2845), .A2(keyout[69]), .S0(n1447), .Y(n4387) );
  MUX21X1_HVT U845 ( .A1(n2844), .A2(keyout[69]), .S0(n1448), .Y(n4386) );
  MUX21X1_HVT U846 ( .A1(n2843), .A2(keyout[69]), .S0(n1449), .Y(n4385) );
  MUX21X1_HVT U847 ( .A1(n2842), .A2(keyout[69]), .S0(n1450), .Y(n4384) );
  MUX21X1_HVT U848 ( .A1(n2841), .A2(keyout[69]), .S0(n1451), .Y(n4383) );
  MUX21X1_HVT U849 ( .A1(n2840), .A2(keyout[69]), .S0(n1452), .Y(n4382) );
  MUX21X1_HVT U850 ( .A1(n2839), .A2(keyout[69]), .S0(n1453), .Y(n4381) );
  MUX21X1_HVT U851 ( .A1(n2838), .A2(keyout[69]), .S0(n1454), .Y(n4380) );
  MUX21X1_HVT U852 ( .A1(n2837), .A2(keyout[70]), .S0(n1447), .Y(n4379) );
  MUX21X1_HVT U853 ( .A1(n2836), .A2(keyout[70]), .S0(n1448), .Y(n4378) );
  MUX21X1_HVT U854 ( .A1(n2835), .A2(keyout[70]), .S0(n1449), .Y(n4377) );
  MUX21X1_HVT U855 ( .A1(n2834), .A2(keyout[70]), .S0(n1450), .Y(n4376) );
  MUX21X1_HVT U856 ( .A1(n2833), .A2(keyout[70]), .S0(n1451), .Y(n4375) );
  MUX21X1_HVT U857 ( .A1(n2832), .A2(keyout[70]), .S0(n1452), .Y(n4374) );
  MUX21X1_HVT U858 ( .A1(n2831), .A2(keyout[70]), .S0(n1453), .Y(n4373) );
  MUX21X1_HVT U859 ( .A1(n2830), .A2(keyout[70]), .S0(n1454), .Y(n4372) );
  MUX21X1_HVT U860 ( .A1(n2829), .A2(keyout[71]), .S0(n1447), .Y(n4371) );
  MUX21X1_HVT U861 ( .A1(n2828), .A2(keyout[71]), .S0(n1448), .Y(n4370) );
  MUX21X1_HVT U862 ( .A1(n2827), .A2(keyout[71]), .S0(n1449), .Y(n4369) );
  MUX21X1_HVT U863 ( .A1(n2826), .A2(keyout[71]), .S0(n1450), .Y(n4368) );
  MUX21X1_HVT U864 ( .A1(n2825), .A2(keyout[71]), .S0(n1451), .Y(n4367) );
  MUX21X1_HVT U865 ( .A1(n2824), .A2(keyout[71]), .S0(n1452), .Y(n4366) );
  MUX21X1_HVT U866 ( .A1(n2823), .A2(keyout[71]), .S0(n1453), .Y(n4365) );
  MUX21X1_HVT U867 ( .A1(n2822), .A2(keyout[71]), .S0(n1454), .Y(n4364) );
  MUX21X1_HVT U868 ( .A1(n2821), .A2(keyout[72]), .S0(n1447), .Y(n4363) );
  MUX21X1_HVT U869 ( .A1(n2820), .A2(keyout[72]), .S0(n1448), .Y(n4362) );
  MUX21X1_HVT U870 ( .A1(n2819), .A2(keyout[72]), .S0(n1449), .Y(n4361) );
  MUX21X1_HVT U871 ( .A1(n2818), .A2(keyout[72]), .S0(n1450), .Y(n4360) );
  MUX21X1_HVT U872 ( .A1(n2817), .A2(keyout[72]), .S0(n1451), .Y(n4359) );
  MUX21X1_HVT U873 ( .A1(n2816), .A2(keyout[72]), .S0(n1452), .Y(n4358) );
  MUX21X1_HVT U874 ( .A1(n2815), .A2(keyout[72]), .S0(n1453), .Y(n4357) );
  MUX21X1_HVT U875 ( .A1(n2814), .A2(keyout[72]), .S0(n1454), .Y(n4356) );
  MUX21X1_HVT U876 ( .A1(n2813), .A2(keyout[73]), .S0(n1447), .Y(n4355) );
  MUX21X1_HVT U877 ( .A1(n2812), .A2(keyout[73]), .S0(n1448), .Y(n4354) );
  MUX21X1_HVT U878 ( .A1(n2811), .A2(keyout[73]), .S0(n1449), .Y(n4353) );
  MUX21X1_HVT U879 ( .A1(n2810), .A2(keyout[73]), .S0(n1450), .Y(n4352) );
  MUX21X1_HVT U880 ( .A1(n2809), .A2(keyout[73]), .S0(n1451), .Y(n4351) );
  MUX21X1_HVT U881 ( .A1(n2808), .A2(keyout[73]), .S0(n1452), .Y(n4350) );
  MUX21X1_HVT U882 ( .A1(n2807), .A2(keyout[73]), .S0(n1453), .Y(n4349) );
  MUX21X1_HVT U883 ( .A1(n2806), .A2(keyout[73]), .S0(n1454), .Y(n4348) );
  MUX21X1_HVT U884 ( .A1(n2805), .A2(keyout[74]), .S0(n1447), .Y(n4347) );
  MUX21X1_HVT U885 ( .A1(n2804), .A2(keyout[74]), .S0(n1448), .Y(n4346) );
  MUX21X1_HVT U886 ( .A1(n2803), .A2(keyout[74]), .S0(n1449), .Y(n4345) );
  MUX21X1_HVT U887 ( .A1(n2802), .A2(keyout[74]), .S0(n1450), .Y(n4344) );
  MUX21X1_HVT U888 ( .A1(n2801), .A2(keyout[74]), .S0(n1451), .Y(n4343) );
  MUX21X1_HVT U889 ( .A1(n2800), .A2(keyout[74]), .S0(n1452), .Y(n4342) );
  MUX21X1_HVT U890 ( .A1(n2799), .A2(keyout[74]), .S0(n1453), .Y(n4341) );
  MUX21X1_HVT U891 ( .A1(n2798), .A2(keyout[74]), .S0(n1454), .Y(n4340) );
  MUX21X1_HVT U892 ( .A1(n2797), .A2(keyout[75]), .S0(n1447), .Y(n4339) );
  MUX21X1_HVT U893 ( .A1(n2796), .A2(keyout[75]), .S0(n1448), .Y(n4338) );
  MUX21X1_HVT U894 ( .A1(n2795), .A2(keyout[75]), .S0(n1449), .Y(n4337) );
  MUX21X1_HVT U895 ( .A1(n2794), .A2(keyout[75]), .S0(n1450), .Y(n4336) );
  MUX21X1_HVT U896 ( .A1(n2793), .A2(keyout[75]), .S0(n1451), .Y(n4335) );
  MUX21X1_HVT U897 ( .A1(n2792), .A2(keyout[75]), .S0(n1452), .Y(n4334) );
  MUX21X1_HVT U898 ( .A1(n2791), .A2(keyout[75]), .S0(n1453), .Y(n4333) );
  MUX21X1_HVT U899 ( .A1(n2790), .A2(keyout[75]), .S0(n1454), .Y(n4332) );
  MUX21X1_HVT U900 ( .A1(n2789), .A2(keyout[76]), .S0(n1447), .Y(n4331) );
  MUX21X1_HVT U901 ( .A1(n2788), .A2(keyout[76]), .S0(n1448), .Y(n4330) );
  MUX21X1_HVT U902 ( .A1(n2787), .A2(keyout[76]), .S0(n1449), .Y(n4329) );
  MUX21X1_HVT U903 ( .A1(n2786), .A2(keyout[76]), .S0(n1450), .Y(n4328) );
  MUX21X1_HVT U904 ( .A1(n2785), .A2(keyout[76]), .S0(n1451), .Y(n4327) );
  MUX21X1_HVT U905 ( .A1(n2784), .A2(keyout[76]), .S0(n1452), .Y(n4326) );
  MUX21X1_HVT U906 ( .A1(n2783), .A2(keyout[76]), .S0(n1453), .Y(n4325) );
  MUX21X1_HVT U907 ( .A1(n2782), .A2(keyout[76]), .S0(n1454), .Y(n4324) );
  MUX21X1_HVT U908 ( .A1(n2781), .A2(keyout[77]), .S0(n1447), .Y(n4323) );
  MUX21X1_HVT U909 ( .A1(n2780), .A2(keyout[77]), .S0(n1448), .Y(n4322) );
  MUX21X1_HVT U910 ( .A1(n2779), .A2(keyout[77]), .S0(n1449), .Y(n4321) );
  MUX21X1_HVT U911 ( .A1(n2778), .A2(keyout[77]), .S0(n1450), .Y(n4320) );
  MUX21X1_HVT U912 ( .A1(n2777), .A2(keyout[77]), .S0(n1451), .Y(n4319) );
  MUX21X1_HVT U913 ( .A1(n2776), .A2(keyout[77]), .S0(n1452), .Y(n4318) );
  MUX21X1_HVT U914 ( .A1(n2775), .A2(keyout[77]), .S0(n1453), .Y(n4317) );
  MUX21X1_HVT U915 ( .A1(n2774), .A2(keyout[77]), .S0(n1454), .Y(n4316) );
  MUX21X1_HVT U916 ( .A1(n2773), .A2(keyout[78]), .S0(n1447), .Y(n4315) );
  MUX21X1_HVT U917 ( .A1(n2772), .A2(keyout[78]), .S0(n1448), .Y(n4314) );
  MUX21X1_HVT U918 ( .A1(n2771), .A2(keyout[78]), .S0(n1449), .Y(n4313) );
  MUX21X1_HVT U919 ( .A1(n2770), .A2(keyout[78]), .S0(n1450), .Y(n4312) );
  MUX21X1_HVT U920 ( .A1(n2769), .A2(keyout[78]), .S0(n1451), .Y(n4311) );
  MUX21X1_HVT U921 ( .A1(n2768), .A2(keyout[78]), .S0(n1452), .Y(n4310) );
  MUX21X1_HVT U922 ( .A1(n2767), .A2(keyout[78]), .S0(n1453), .Y(n4309) );
  MUX21X1_HVT U923 ( .A1(n2766), .A2(keyout[78]), .S0(n1454), .Y(n4308) );
  MUX21X1_HVT U924 ( .A1(n2765), .A2(keyout[79]), .S0(n1447), .Y(n4307) );
  MUX21X1_HVT U925 ( .A1(n2764), .A2(keyout[79]), .S0(n1448), .Y(n4306) );
  MUX21X1_HVT U926 ( .A1(n2763), .A2(keyout[79]), .S0(n1449), .Y(n4305) );
  MUX21X1_HVT U927 ( .A1(n2762), .A2(keyout[79]), .S0(n1450), .Y(n4304) );
  MUX21X1_HVT U928 ( .A1(n2761), .A2(keyout[79]), .S0(n1451), .Y(n4303) );
  MUX21X1_HVT U929 ( .A1(n2760), .A2(keyout[79]), .S0(n1452), .Y(n4302) );
  MUX21X1_HVT U930 ( .A1(n2759), .A2(keyout[79]), .S0(n1453), .Y(n4301) );
  MUX21X1_HVT U931 ( .A1(n2758), .A2(keyout[79]), .S0(n1454), .Y(n4300) );
  MUX21X1_HVT U932 ( .A1(n2757), .A2(keyout[80]), .S0(n1447), .Y(n4299) );
  MUX21X1_HVT U933 ( .A1(n2756), .A2(keyout[80]), .S0(n1448), .Y(n4298) );
  MUX21X1_HVT U934 ( .A1(n2755), .A2(keyout[80]), .S0(n1449), .Y(n4297) );
  MUX21X1_HVT U935 ( .A1(n2754), .A2(keyout[80]), .S0(n1450), .Y(n4296) );
  MUX21X1_HVT U936 ( .A1(n2753), .A2(keyout[80]), .S0(n1451), .Y(n4295) );
  MUX21X1_HVT U937 ( .A1(n2752), .A2(keyout[80]), .S0(n1452), .Y(n4294) );
  MUX21X1_HVT U938 ( .A1(n2751), .A2(keyout[80]), .S0(n1453), .Y(n4293) );
  MUX21X1_HVT U939 ( .A1(n2750), .A2(keyout[80]), .S0(n1454), .Y(n4292) );
  MUX21X1_HVT U940 ( .A1(n2749), .A2(keyout[81]), .S0(n1447), .Y(n4291) );
  MUX21X1_HVT U941 ( .A1(n2748), .A2(keyout[81]), .S0(n1448), .Y(n4290) );
  MUX21X1_HVT U942 ( .A1(n2747), .A2(keyout[81]), .S0(n1449), .Y(n4289) );
  MUX21X1_HVT U943 ( .A1(n2746), .A2(keyout[81]), .S0(n1450), .Y(n4288) );
  MUX21X1_HVT U944 ( .A1(n2745), .A2(keyout[81]), .S0(n1451), .Y(n4287) );
  MUX21X1_HVT U945 ( .A1(n2744), .A2(keyout[81]), .S0(n1452), .Y(n4286) );
  MUX21X1_HVT U946 ( .A1(n2743), .A2(keyout[81]), .S0(n1453), .Y(n4285) );
  MUX21X1_HVT U947 ( .A1(n2742), .A2(keyout[81]), .S0(n1454), .Y(n4284) );
  MUX21X1_HVT U948 ( .A1(n2741), .A2(keyout[82]), .S0(n1447), .Y(n4283) );
  MUX21X1_HVT U949 ( .A1(n2740), .A2(keyout[82]), .S0(n1448), .Y(n4282) );
  MUX21X1_HVT U950 ( .A1(n2739), .A2(keyout[82]), .S0(n1449), .Y(n4281) );
  MUX21X1_HVT U951 ( .A1(n2738), .A2(keyout[82]), .S0(n1450), .Y(n4280) );
  MUX21X1_HVT U952 ( .A1(n2737), .A2(keyout[82]), .S0(n1451), .Y(n4279) );
  MUX21X1_HVT U953 ( .A1(n2736), .A2(keyout[82]), .S0(n1452), .Y(n4278) );
  MUX21X1_HVT U954 ( .A1(n2735), .A2(keyout[82]), .S0(n1453), .Y(n4277) );
  MUX21X1_HVT U955 ( .A1(n2734), .A2(keyout[82]), .S0(n1454), .Y(n4276) );
  MUX21X1_HVT U956 ( .A1(n2733), .A2(keyout[83]), .S0(n1447), .Y(n4275) );
  MUX21X1_HVT U957 ( .A1(n2732), .A2(keyout[83]), .S0(n1448), .Y(n4274) );
  MUX21X1_HVT U958 ( .A1(n2731), .A2(keyout[83]), .S0(n1449), .Y(n4273) );
  MUX21X1_HVT U959 ( .A1(n2730), .A2(keyout[83]), .S0(n1450), .Y(n4272) );
  MUX21X1_HVT U960 ( .A1(n2729), .A2(keyout[83]), .S0(n1451), .Y(n4271) );
  MUX21X1_HVT U961 ( .A1(n2728), .A2(keyout[83]), .S0(n1452), .Y(n4270) );
  MUX21X1_HVT U962 ( .A1(n2727), .A2(keyout[83]), .S0(n1453), .Y(n4269) );
  MUX21X1_HVT U963 ( .A1(n2726), .A2(keyout[83]), .S0(n1454), .Y(n4268) );
  MUX21X1_HVT U964 ( .A1(n2725), .A2(keyout[84]), .S0(n1447), .Y(n4267) );
  MUX21X1_HVT U965 ( .A1(n2724), .A2(keyout[84]), .S0(n1448), .Y(n4266) );
  MUX21X1_HVT U966 ( .A1(n2723), .A2(keyout[84]), .S0(n1449), .Y(n4265) );
  MUX21X1_HVT U967 ( .A1(n2722), .A2(keyout[84]), .S0(n1450), .Y(n4264) );
  MUX21X1_HVT U968 ( .A1(n2721), .A2(keyout[84]), .S0(n1451), .Y(n4263) );
  MUX21X1_HVT U969 ( .A1(n2720), .A2(keyout[84]), .S0(n1452), .Y(n4262) );
  MUX21X1_HVT U970 ( .A1(n2719), .A2(keyout[84]), .S0(n1453), .Y(n4261) );
  MUX21X1_HVT U971 ( .A1(n2718), .A2(keyout[84]), .S0(n1454), .Y(n4260) );
  MUX21X1_HVT U972 ( .A1(n2717), .A2(keyout[85]), .S0(n1447), .Y(n4259) );
  MUX21X1_HVT U973 ( .A1(n2716), .A2(keyout[85]), .S0(n1448), .Y(n4258) );
  MUX21X1_HVT U974 ( .A1(n2715), .A2(keyout[85]), .S0(n1449), .Y(n4257) );
  MUX21X1_HVT U975 ( .A1(n2714), .A2(keyout[85]), .S0(n1450), .Y(n4256) );
  MUX21X1_HVT U976 ( .A1(n2713), .A2(keyout[85]), .S0(n1451), .Y(n4255) );
  MUX21X1_HVT U977 ( .A1(n2712), .A2(keyout[85]), .S0(n1452), .Y(n4254) );
  MUX21X1_HVT U978 ( .A1(n2711), .A2(keyout[85]), .S0(n1453), .Y(n4253) );
  MUX21X1_HVT U979 ( .A1(n2710), .A2(keyout[85]), .S0(n1454), .Y(n4252) );
  MUX21X1_HVT U980 ( .A1(n2709), .A2(keyout[86]), .S0(n1447), .Y(n4251) );
  MUX21X1_HVT U981 ( .A1(n2708), .A2(keyout[86]), .S0(n1448), .Y(n4250) );
  MUX21X1_HVT U982 ( .A1(n2707), .A2(keyout[86]), .S0(n1449), .Y(n4249) );
  MUX21X1_HVT U983 ( .A1(n2706), .A2(keyout[86]), .S0(n1450), .Y(n4248) );
  MUX21X1_HVT U984 ( .A1(n2705), .A2(keyout[86]), .S0(n1451), .Y(n4247) );
  MUX21X1_HVT U985 ( .A1(n2704), .A2(keyout[86]), .S0(n1452), .Y(n4246) );
  MUX21X1_HVT U986 ( .A1(n2703), .A2(keyout[86]), .S0(n1453), .Y(n4245) );
  MUX21X1_HVT U987 ( .A1(n2702), .A2(keyout[86]), .S0(n1454), .Y(n4244) );
  MUX21X1_HVT U988 ( .A1(n2701), .A2(keyout[87]), .S0(n1447), .Y(n4243) );
  MUX21X1_HVT U989 ( .A1(n2700), .A2(keyout[87]), .S0(n1448), .Y(n4242) );
  MUX21X1_HVT U990 ( .A1(n2699), .A2(keyout[87]), .S0(n1449), .Y(n4241) );
  MUX21X1_HVT U991 ( .A1(n2698), .A2(keyout[87]), .S0(n1450), .Y(n4240) );
  MUX21X1_HVT U992 ( .A1(n2697), .A2(keyout[87]), .S0(n1451), .Y(n4239) );
  MUX21X1_HVT U993 ( .A1(n2696), .A2(keyout[87]), .S0(n1452), .Y(n4238) );
  MUX21X1_HVT U994 ( .A1(n2695), .A2(keyout[87]), .S0(n1453), .Y(n4237) );
  MUX21X1_HVT U995 ( .A1(n2694), .A2(keyout[87]), .S0(n1454), .Y(n4236) );
  MUX21X1_HVT U996 ( .A1(n2693), .A2(keyout[88]), .S0(n1447), .Y(n4235) );
  MUX21X1_HVT U997 ( .A1(n2692), .A2(keyout[88]), .S0(n1448), .Y(n4234) );
  MUX21X1_HVT U998 ( .A1(n2691), .A2(keyout[88]), .S0(n1449), .Y(n4233) );
  MUX21X1_HVT U999 ( .A1(n2690), .A2(keyout[88]), .S0(n1450), .Y(n4232) );
  MUX21X1_HVT U1000 ( .A1(n2689), .A2(keyout[88]), .S0(n1451), .Y(n4231) );
  MUX21X1_HVT U1001 ( .A1(n2688), .A2(keyout[88]), .S0(n1452), .Y(n4230) );
  MUX21X1_HVT U1002 ( .A1(n2687), .A2(keyout[88]), .S0(n1453), .Y(n4229) );
  MUX21X1_HVT U1003 ( .A1(n2686), .A2(keyout[88]), .S0(n1454), .Y(n4228) );
  MUX21X1_HVT U1004 ( .A1(n2685), .A2(keyout[89]), .S0(n1447), .Y(n4227) );
  MUX21X1_HVT U1005 ( .A1(n2684), .A2(keyout[89]), .S0(n1448), .Y(n4226) );
  MUX21X1_HVT U1006 ( .A1(n2683), .A2(keyout[89]), .S0(n1449), .Y(n4225) );
  MUX21X1_HVT U1007 ( .A1(n2682), .A2(keyout[89]), .S0(n1450), .Y(n4224) );
  MUX21X1_HVT U1008 ( .A1(n2681), .A2(keyout[89]), .S0(n1451), .Y(n4223) );
  MUX21X1_HVT U1009 ( .A1(n2680), .A2(keyout[89]), .S0(n1452), .Y(n4222) );
  MUX21X1_HVT U1010 ( .A1(n2679), .A2(keyout[89]), .S0(n1453), .Y(n4221) );
  MUX21X1_HVT U1011 ( .A1(n2678), .A2(keyout[89]), .S0(n1454), .Y(n4220) );
  MUX21X1_HVT U1012 ( .A1(n2677), .A2(keyout[90]), .S0(n1447), .Y(n4219) );
  MUX21X1_HVT U1013 ( .A1(n2676), .A2(keyout[90]), .S0(n1448), .Y(n4218) );
  MUX21X1_HVT U1014 ( .A1(n2675), .A2(keyout[90]), .S0(n1449), .Y(n4217) );
  MUX21X1_HVT U1015 ( .A1(n2674), .A2(keyout[90]), .S0(n1450), .Y(n4216) );
  MUX21X1_HVT U1016 ( .A1(n2673), .A2(keyout[90]), .S0(n1451), .Y(n4215) );
  MUX21X1_HVT U1017 ( .A1(n2672), .A2(keyout[90]), .S0(n1452), .Y(n4214) );
  MUX21X1_HVT U1018 ( .A1(n2671), .A2(keyout[90]), .S0(n1453), .Y(n4213) );
  MUX21X1_HVT U1019 ( .A1(n2670), .A2(keyout[90]), .S0(n1454), .Y(n4212) );
  MUX21X1_HVT U1020 ( .A1(n2669), .A2(keyout[91]), .S0(n1447), .Y(n4211) );
  MUX21X1_HVT U1021 ( .A1(n2668), .A2(keyout[91]), .S0(n1448), .Y(n4210) );
  MUX21X1_HVT U1022 ( .A1(n2667), .A2(keyout[91]), .S0(n1449), .Y(n4209) );
  MUX21X1_HVT U1023 ( .A1(n2666), .A2(keyout[91]), .S0(n1450), .Y(n4208) );
  MUX21X1_HVT U1024 ( .A1(n2665), .A2(keyout[91]), .S0(n1451), .Y(n4207) );
  MUX21X1_HVT U1025 ( .A1(n2664), .A2(keyout[91]), .S0(n1452), .Y(n4206) );
  MUX21X1_HVT U1026 ( .A1(n2663), .A2(keyout[91]), .S0(n1453), .Y(n4205) );
  MUX21X1_HVT U1027 ( .A1(n2662), .A2(keyout[91]), .S0(n1454), .Y(n4204) );
  MUX21X1_HVT U1028 ( .A1(n2661), .A2(keyout[92]), .S0(n1447), .Y(n4203) );
  MUX21X1_HVT U1029 ( .A1(n2660), .A2(keyout[92]), .S0(n1448), .Y(n4202) );
  MUX21X1_HVT U1030 ( .A1(n2659), .A2(keyout[92]), .S0(n1449), .Y(n4201) );
  MUX21X1_HVT U1031 ( .A1(n2658), .A2(keyout[92]), .S0(n1450), .Y(n4200) );
  MUX21X1_HVT U1032 ( .A1(n2657), .A2(keyout[92]), .S0(n1451), .Y(n4199) );
  MUX21X1_HVT U1033 ( .A1(n2656), .A2(keyout[92]), .S0(n1452), .Y(n4198) );
  MUX21X1_HVT U1034 ( .A1(n2655), .A2(keyout[92]), .S0(n1453), .Y(n4197) );
  MUX21X1_HVT U1035 ( .A1(n2654), .A2(keyout[92]), .S0(n1454), .Y(n4196) );
  MUX21X1_HVT U1036 ( .A1(n2653), .A2(keyout[93]), .S0(n1447), .Y(n4195) );
  MUX21X1_HVT U1037 ( .A1(n2652), .A2(keyout[93]), .S0(n1448), .Y(n4194) );
  MUX21X1_HVT U1038 ( .A1(n2651), .A2(keyout[93]), .S0(n1449), .Y(n4193) );
  MUX21X1_HVT U1039 ( .A1(n2650), .A2(keyout[93]), .S0(n1450), .Y(n4192) );
  MUX21X1_HVT U1040 ( .A1(n2649), .A2(keyout[93]), .S0(n1451), .Y(n4191) );
  MUX21X1_HVT U1041 ( .A1(n2648), .A2(keyout[93]), .S0(n1452), .Y(n4190) );
  MUX21X1_HVT U1042 ( .A1(n2647), .A2(keyout[93]), .S0(n1453), .Y(n4189) );
  MUX21X1_HVT U1043 ( .A1(n2646), .A2(keyout[93]), .S0(n1454), .Y(n4188) );
  MUX21X1_HVT U1044 ( .A1(n2645), .A2(keyout[94]), .S0(n1447), .Y(n4187) );
  MUX21X1_HVT U1045 ( .A1(n2644), .A2(keyout[94]), .S0(n1448), .Y(n4186) );
  MUX21X1_HVT U1046 ( .A1(n2643), .A2(keyout[94]), .S0(n1449), .Y(n4185) );
  MUX21X1_HVT U1047 ( .A1(n2642), .A2(keyout[94]), .S0(n1450), .Y(n4184) );
  MUX21X1_HVT U1048 ( .A1(n2641), .A2(keyout[94]), .S0(n1451), .Y(n4183) );
  MUX21X1_HVT U1049 ( .A1(n2640), .A2(keyout[94]), .S0(n1452), .Y(n4182) );
  MUX21X1_HVT U1050 ( .A1(n2639), .A2(keyout[94]), .S0(n1453), .Y(n4181) );
  MUX21X1_HVT U1051 ( .A1(n2638), .A2(keyout[94]), .S0(n1454), .Y(n4180) );
  MUX21X1_HVT U1052 ( .A1(n2637), .A2(keyout[95]), .S0(n1447), .Y(n4179) );
  MUX21X1_HVT U1053 ( .A1(n2636), .A2(keyout[95]), .S0(n1448), .Y(n4178) );
  MUX21X1_HVT U1054 ( .A1(n2635), .A2(keyout[95]), .S0(n1449), .Y(n4177) );
  MUX21X1_HVT U1055 ( .A1(n2634), .A2(keyout[95]), .S0(n1450), .Y(n4176) );
  MUX21X1_HVT U1056 ( .A1(n2633), .A2(keyout[95]), .S0(n1451), .Y(n4175) );
  MUX21X1_HVT U1057 ( .A1(n2632), .A2(keyout[95]), .S0(n1452), .Y(n4174) );
  MUX21X1_HVT U1058 ( .A1(n2631), .A2(keyout[95]), .S0(n1453), .Y(n4173) );
  MUX21X1_HVT U1059 ( .A1(n2630), .A2(keyout[95]), .S0(n1454), .Y(n4172) );
  MUX21X1_HVT U1060 ( .A1(n2629), .A2(keyout[96]), .S0(n1447), .Y(n4171) );
  MUX21X1_HVT U1061 ( .A1(n2628), .A2(keyout[96]), .S0(n1448), .Y(n4170) );
  MUX21X1_HVT U1062 ( .A1(n2627), .A2(keyout[96]), .S0(n1449), .Y(n4169) );
  MUX21X1_HVT U1063 ( .A1(n2626), .A2(keyout[96]), .S0(n1450), .Y(n4168) );
  MUX21X1_HVT U1064 ( .A1(n2625), .A2(keyout[96]), .S0(n1451), .Y(n4167) );
  MUX21X1_HVT U1065 ( .A1(n2624), .A2(keyout[96]), .S0(n1452), .Y(n4166) );
  MUX21X1_HVT U1066 ( .A1(n2623), .A2(keyout[96]), .S0(n1453), .Y(n4165) );
  MUX21X1_HVT U1067 ( .A1(n2622), .A2(keyout[96]), .S0(n1454), .Y(n4164) );
  MUX21X1_HVT U1068 ( .A1(n2621), .A2(keyout[97]), .S0(n1447), .Y(n4163) );
  MUX21X1_HVT U1069 ( .A1(n2620), .A2(keyout[97]), .S0(n1448), .Y(n4162) );
  MUX21X1_HVT U1070 ( .A1(n2619), .A2(keyout[97]), .S0(n1449), .Y(n4161) );
  MUX21X1_HVT U1071 ( .A1(n2618), .A2(keyout[97]), .S0(n1450), .Y(n4160) );
  MUX21X1_HVT U1072 ( .A1(n2617), .A2(keyout[97]), .S0(n1451), .Y(n4159) );
  MUX21X1_HVT U1073 ( .A1(n2616), .A2(keyout[97]), .S0(n1452), .Y(n4158) );
  MUX21X1_HVT U1074 ( .A1(n2615), .A2(keyout[97]), .S0(n1453), .Y(n4157) );
  MUX21X1_HVT U1075 ( .A1(n2614), .A2(keyout[97]), .S0(n1454), .Y(n4156) );
  MUX21X1_HVT U1076 ( .A1(n2613), .A2(keyout[98]), .S0(n1447), .Y(n4155) );
  MUX21X1_HVT U1077 ( .A1(n2612), .A2(keyout[98]), .S0(n1448), .Y(n4154) );
  MUX21X1_HVT U1078 ( .A1(n2611), .A2(keyout[98]), .S0(n1449), .Y(n4153) );
  MUX21X1_HVT U1079 ( .A1(n2610), .A2(keyout[98]), .S0(n1450), .Y(n4152) );
  MUX21X1_HVT U1080 ( .A1(n2609), .A2(keyout[98]), .S0(n1451), .Y(n4151) );
  MUX21X1_HVT U1081 ( .A1(n2608), .A2(keyout[98]), .S0(n1452), .Y(n4150) );
  MUX21X1_HVT U1082 ( .A1(n2607), .A2(keyout[98]), .S0(n1453), .Y(n4149) );
  MUX21X1_HVT U1083 ( .A1(n2606), .A2(keyout[98]), .S0(n1454), .Y(n4148) );
  MUX21X1_HVT U1084 ( .A1(n2605), .A2(keyout[99]), .S0(n1447), .Y(n4147) );
  MUX21X1_HVT U1085 ( .A1(n2604), .A2(keyout[99]), .S0(n1448), .Y(n4146) );
  MUX21X1_HVT U1086 ( .A1(n2603), .A2(keyout[99]), .S0(n1449), .Y(n4145) );
  MUX21X1_HVT U1087 ( .A1(n2602), .A2(keyout[99]), .S0(n1450), .Y(n4144) );
  MUX21X1_HVT U1088 ( .A1(n2601), .A2(keyout[99]), .S0(n1451), .Y(n4143) );
  MUX21X1_HVT U1089 ( .A1(n2600), .A2(keyout[99]), .S0(n1452), .Y(n4142) );
  MUX21X1_HVT U1090 ( .A1(n2599), .A2(keyout[99]), .S0(n1453), .Y(n4141) );
  MUX21X1_HVT U1091 ( .A1(n2598), .A2(keyout[99]), .S0(n1454), .Y(n4140) );
  MUX21X1_HVT U1092 ( .A1(n2597), .A2(keyout[100]), .S0(n1447), .Y(n4139) );
  MUX21X1_HVT U1093 ( .A1(n2596), .A2(keyout[100]), .S0(n1448), .Y(n4138) );
  MUX21X1_HVT U1094 ( .A1(n2595), .A2(keyout[100]), .S0(n1449), .Y(n4137) );
  MUX21X1_HVT U1095 ( .A1(n2594), .A2(keyout[100]), .S0(n1450), .Y(n4136) );
  MUX21X1_HVT U1096 ( .A1(n2593), .A2(keyout[100]), .S0(n1451), .Y(n4135) );
  MUX21X1_HVT U1097 ( .A1(n2592), .A2(keyout[100]), .S0(n1452), .Y(n4134) );
  MUX21X1_HVT U1098 ( .A1(n2591), .A2(keyout[100]), .S0(n1453), .Y(n4133) );
  MUX21X1_HVT U1099 ( .A1(n2590), .A2(keyout[100]), .S0(n1454), .Y(n4132) );
  MUX21X1_HVT U1100 ( .A1(n2589), .A2(keyout[101]), .S0(n1447), .Y(n4131) );
  MUX21X1_HVT U1101 ( .A1(n2588), .A2(keyout[101]), .S0(n1448), .Y(n4130) );
  MUX21X1_HVT U1102 ( .A1(n2587), .A2(keyout[101]), .S0(n1449), .Y(n4129) );
  MUX21X1_HVT U1103 ( .A1(n2586), .A2(keyout[101]), .S0(n1450), .Y(n4128) );
  MUX21X1_HVT U1104 ( .A1(n2585), .A2(keyout[101]), .S0(n1451), .Y(n4127) );
  MUX21X1_HVT U1105 ( .A1(n2584), .A2(keyout[101]), .S0(n1452), .Y(n4126) );
  MUX21X1_HVT U1106 ( .A1(n2583), .A2(keyout[101]), .S0(n1453), .Y(n4125) );
  MUX21X1_HVT U1107 ( .A1(n2582), .A2(keyout[101]), .S0(n1454), .Y(n4124) );
  MUX21X1_HVT U1108 ( .A1(n2581), .A2(keyout[102]), .S0(n1447), .Y(n4123) );
  MUX21X1_HVT U1109 ( .A1(n2580), .A2(keyout[102]), .S0(n1448), .Y(n4122) );
  MUX21X1_HVT U1110 ( .A1(n2579), .A2(keyout[102]), .S0(n1449), .Y(n4121) );
  MUX21X1_HVT U1111 ( .A1(n2578), .A2(keyout[102]), .S0(n1450), .Y(n4120) );
  MUX21X1_HVT U1112 ( .A1(n2577), .A2(keyout[102]), .S0(n1451), .Y(n4119) );
  MUX21X1_HVT U1113 ( .A1(n2576), .A2(keyout[102]), .S0(n1452), .Y(n4118) );
  MUX21X1_HVT U1114 ( .A1(n2575), .A2(keyout[102]), .S0(n1453), .Y(n4117) );
  MUX21X1_HVT U1115 ( .A1(n2574), .A2(keyout[102]), .S0(n1454), .Y(n4116) );
  MUX21X1_HVT U1116 ( .A1(n2573), .A2(keyout[103]), .S0(n1447), .Y(n4115) );
  MUX21X1_HVT U1117 ( .A1(n2572), .A2(keyout[103]), .S0(n1448), .Y(n4114) );
  MUX21X1_HVT U1118 ( .A1(n2571), .A2(keyout[103]), .S0(n1449), .Y(n4113) );
  MUX21X1_HVT U1119 ( .A1(n2570), .A2(keyout[103]), .S0(n1450), .Y(n4112) );
  MUX21X1_HVT U1120 ( .A1(n2569), .A2(keyout[103]), .S0(n1451), .Y(n4111) );
  MUX21X1_HVT U1121 ( .A1(n2568), .A2(keyout[103]), .S0(n1452), .Y(n4110) );
  MUX21X1_HVT U1122 ( .A1(n2567), .A2(keyout[103]), .S0(n1453), .Y(n4109) );
  MUX21X1_HVT U1123 ( .A1(n2566), .A2(keyout[103]), .S0(n1454), .Y(n4108) );
  MUX21X1_HVT U1124 ( .A1(n2565), .A2(keyout[104]), .S0(n1447), .Y(n4107) );
  MUX21X1_HVT U1125 ( .A1(n2564), .A2(keyout[104]), .S0(n1448), .Y(n4106) );
  MUX21X1_HVT U1126 ( .A1(n2563), .A2(keyout[104]), .S0(n1449), .Y(n4105) );
  MUX21X1_HVT U1127 ( .A1(n2562), .A2(keyout[104]), .S0(n1450), .Y(n4104) );
  MUX21X1_HVT U1128 ( .A1(n2561), .A2(keyout[104]), .S0(n1451), .Y(n4103) );
  MUX21X1_HVT U1129 ( .A1(n2560), .A2(keyout[104]), .S0(n1452), .Y(n4102) );
  MUX21X1_HVT U1130 ( .A1(n2559), .A2(keyout[104]), .S0(n1453), .Y(n4101) );
  MUX21X1_HVT U1131 ( .A1(n2558), .A2(keyout[104]), .S0(n1454), .Y(n4100) );
  MUX21X1_HVT U1132 ( .A1(n2557), .A2(keyout[105]), .S0(n1447), .Y(n4099) );
  MUX21X1_HVT U1133 ( .A1(n2556), .A2(keyout[105]), .S0(n1448), .Y(n4098) );
  MUX21X1_HVT U1134 ( .A1(n2555), .A2(keyout[105]), .S0(n1449), .Y(n4097) );
  MUX21X1_HVT U1135 ( .A1(n2554), .A2(keyout[105]), .S0(n1450), .Y(n4096) );
  MUX21X1_HVT U1136 ( .A1(n2553), .A2(keyout[105]), .S0(n1451), .Y(n4095) );
  MUX21X1_HVT U1137 ( .A1(n2552), .A2(keyout[105]), .S0(n1452), .Y(n4094) );
  MUX21X1_HVT U1138 ( .A1(n2551), .A2(keyout[105]), .S0(n1453), .Y(n4093) );
  MUX21X1_HVT U1139 ( .A1(n2550), .A2(keyout[105]), .S0(n1454), .Y(n4092) );
  MUX21X1_HVT U1140 ( .A1(n2549), .A2(keyout[106]), .S0(n1447), .Y(n4091) );
  MUX21X1_HVT U1141 ( .A1(n2548), .A2(keyout[106]), .S0(n1448), .Y(n4090) );
  MUX21X1_HVT U1142 ( .A1(n2547), .A2(keyout[106]), .S0(n1449), .Y(n4089) );
  MUX21X1_HVT U1143 ( .A1(n2546), .A2(keyout[106]), .S0(n1450), .Y(n4088) );
  MUX21X1_HVT U1144 ( .A1(n2545), .A2(keyout[106]), .S0(n1451), .Y(n4087) );
  MUX21X1_HVT U1145 ( .A1(n2544), .A2(keyout[106]), .S0(n1452), .Y(n4086) );
  MUX21X1_HVT U1146 ( .A1(n2543), .A2(keyout[106]), .S0(n1453), .Y(n4085) );
  MUX21X1_HVT U1147 ( .A1(n2542), .A2(keyout[106]), .S0(n1454), .Y(n4084) );
  MUX21X1_HVT U1148 ( .A1(n2541), .A2(keyout[107]), .S0(n1447), .Y(n4083) );
  MUX21X1_HVT U1149 ( .A1(n2540), .A2(keyout[107]), .S0(n1448), .Y(n4082) );
  MUX21X1_HVT U1150 ( .A1(n2539), .A2(keyout[107]), .S0(n1449), .Y(n4081) );
  MUX21X1_HVT U1151 ( .A1(n2538), .A2(keyout[107]), .S0(n1450), .Y(n4080) );
  MUX21X1_HVT U1152 ( .A1(n2537), .A2(keyout[107]), .S0(n1451), .Y(n4079) );
  MUX21X1_HVT U1153 ( .A1(n2536), .A2(keyout[107]), .S0(n1452), .Y(n4078) );
  MUX21X1_HVT U1154 ( .A1(n2535), .A2(keyout[107]), .S0(n1453), .Y(n4077) );
  MUX21X1_HVT U1155 ( .A1(n2534), .A2(keyout[107]), .S0(n1454), .Y(n4076) );
  MUX21X1_HVT U1156 ( .A1(n2533), .A2(keyout[108]), .S0(n1447), .Y(n4075) );
  MUX21X1_HVT U1157 ( .A1(n2532), .A2(keyout[108]), .S0(n1448), .Y(n4074) );
  MUX21X1_HVT U1158 ( .A1(n2531), .A2(keyout[108]), .S0(n1449), .Y(n4073) );
  MUX21X1_HVT U1159 ( .A1(n2530), .A2(keyout[108]), .S0(n1450), .Y(n4072) );
  MUX21X1_HVT U1160 ( .A1(n2529), .A2(keyout[108]), .S0(n1451), .Y(n4071) );
  MUX21X1_HVT U1161 ( .A1(n2528), .A2(keyout[108]), .S0(n1452), .Y(n4070) );
  MUX21X1_HVT U1162 ( .A1(n2527), .A2(keyout[108]), .S0(n1453), .Y(n4069) );
  MUX21X1_HVT U1163 ( .A1(n2526), .A2(keyout[108]), .S0(n1454), .Y(n4068) );
  MUX21X1_HVT U1164 ( .A1(n2525), .A2(keyout[109]), .S0(n1447), .Y(n4067) );
  MUX21X1_HVT U1165 ( .A1(n2524), .A2(keyout[109]), .S0(n1448), .Y(n4066) );
  MUX21X1_HVT U1166 ( .A1(n2523), .A2(keyout[109]), .S0(n1449), .Y(n4065) );
  MUX21X1_HVT U1167 ( .A1(n2522), .A2(keyout[109]), .S0(n1450), .Y(n4064) );
  MUX21X1_HVT U1168 ( .A1(n2521), .A2(keyout[109]), .S0(n1451), .Y(n4063) );
  MUX21X1_HVT U1169 ( .A1(n2520), .A2(keyout[109]), .S0(n1452), .Y(n4062) );
  MUX21X1_HVT U1170 ( .A1(n2519), .A2(keyout[109]), .S0(n1453), .Y(n4061) );
  MUX21X1_HVT U1171 ( .A1(n2518), .A2(keyout[109]), .S0(n1454), .Y(n4060) );
  MUX21X1_HVT U1172 ( .A1(n2517), .A2(keyout[110]), .S0(n1447), .Y(n4059) );
  MUX21X1_HVT U1173 ( .A1(n2516), .A2(keyout[110]), .S0(n1448), .Y(n4058) );
  MUX21X1_HVT U1174 ( .A1(n2515), .A2(keyout[110]), .S0(n1449), .Y(n4057) );
  MUX21X1_HVT U1175 ( .A1(n2514), .A2(keyout[110]), .S0(n1450), .Y(n4056) );
  MUX21X1_HVT U1176 ( .A1(n2513), .A2(keyout[110]), .S0(n1451), .Y(n4055) );
  MUX21X1_HVT U1177 ( .A1(n2512), .A2(keyout[110]), .S0(n1452), .Y(n4054) );
  MUX21X1_HVT U1178 ( .A1(n2511), .A2(keyout[110]), .S0(n1453), .Y(n4053) );
  MUX21X1_HVT U1179 ( .A1(n2510), .A2(keyout[110]), .S0(n1454), .Y(n4052) );
  MUX21X1_HVT U1180 ( .A1(n2509), .A2(keyout[111]), .S0(n1447), .Y(n4051) );
  MUX21X1_HVT U1181 ( .A1(n2508), .A2(keyout[111]), .S0(n1448), .Y(n4050) );
  MUX21X1_HVT U1182 ( .A1(n2507), .A2(keyout[111]), .S0(n1449), .Y(n4049) );
  MUX21X1_HVT U1183 ( .A1(n2506), .A2(keyout[111]), .S0(n1450), .Y(n4048) );
  MUX21X1_HVT U1184 ( .A1(n2505), .A2(keyout[111]), .S0(n1451), .Y(n4047) );
  MUX21X1_HVT U1185 ( .A1(n2504), .A2(keyout[111]), .S0(n1452), .Y(n4046) );
  MUX21X1_HVT U1186 ( .A1(n2503), .A2(keyout[111]), .S0(n1453), .Y(n4045) );
  MUX21X1_HVT U1187 ( .A1(n2502), .A2(keyout[111]), .S0(n1454), .Y(n4044) );
  MUX21X1_HVT U1188 ( .A1(n2501), .A2(keyout[112]), .S0(n1447), .Y(n4043) );
  MUX21X1_HVT U1189 ( .A1(n2500), .A2(keyout[112]), .S0(n1448), .Y(n4042) );
  MUX21X1_HVT U1190 ( .A1(n2499), .A2(keyout[112]), .S0(n1449), .Y(n4041) );
  MUX21X1_HVT U1191 ( .A1(n2498), .A2(keyout[112]), .S0(n1450), .Y(n4040) );
  MUX21X1_HVT U1192 ( .A1(n2497), .A2(keyout[112]), .S0(n1451), .Y(n4039) );
  MUX21X1_HVT U1193 ( .A1(n2496), .A2(keyout[112]), .S0(n1452), .Y(n4038) );
  MUX21X1_HVT U1194 ( .A1(n2495), .A2(keyout[112]), .S0(n1453), .Y(n4037) );
  MUX21X1_HVT U1195 ( .A1(n2494), .A2(keyout[112]), .S0(n1454), .Y(n4036) );
  MUX21X1_HVT U1196 ( .A1(n2493), .A2(keyout[113]), .S0(n1447), .Y(n4035) );
  MUX21X1_HVT U1197 ( .A1(n2492), .A2(keyout[113]), .S0(n1448), .Y(n4034) );
  MUX21X1_HVT U1198 ( .A1(n2491), .A2(keyout[113]), .S0(n1449), .Y(n4033) );
  MUX21X1_HVT U1199 ( .A1(n2490), .A2(keyout[113]), .S0(n1450), .Y(n4032) );
  MUX21X1_HVT U1200 ( .A1(n2489), .A2(keyout[113]), .S0(n1451), .Y(n4031) );
  MUX21X1_HVT U1201 ( .A1(n2488), .A2(keyout[113]), .S0(n1452), .Y(n4030) );
  MUX21X1_HVT U1202 ( .A1(n2487), .A2(keyout[113]), .S0(n1453), .Y(n4029) );
  MUX21X1_HVT U1203 ( .A1(n2486), .A2(keyout[113]), .S0(n1454), .Y(n4028) );
  MUX21X1_HVT U1204 ( .A1(n2485), .A2(keyout[114]), .S0(n1447), .Y(n4027) );
  MUX21X1_HVT U1205 ( .A1(n2484), .A2(keyout[114]), .S0(n1448), .Y(n4026) );
  MUX21X1_HVT U1206 ( .A1(n2483), .A2(keyout[114]), .S0(n1449), .Y(n4025) );
  MUX21X1_HVT U1207 ( .A1(n2482), .A2(keyout[114]), .S0(n1450), .Y(n4024) );
  MUX21X1_HVT U1208 ( .A1(n2481), .A2(keyout[114]), .S0(n1451), .Y(n4023) );
  MUX21X1_HVT U1209 ( .A1(n2480), .A2(keyout[114]), .S0(n1452), .Y(n4022) );
  MUX21X1_HVT U1210 ( .A1(n2479), .A2(keyout[114]), .S0(n1453), .Y(n4021) );
  MUX21X1_HVT U1211 ( .A1(n2478), .A2(keyout[114]), .S0(n1454), .Y(n4020) );
  MUX21X1_HVT U1212 ( .A1(n2477), .A2(keyout[115]), .S0(n1447), .Y(n4019) );
  MUX21X1_HVT U1213 ( .A1(n2476), .A2(keyout[115]), .S0(n1448), .Y(n4018) );
  MUX21X1_HVT U1214 ( .A1(n2475), .A2(keyout[115]), .S0(n1449), .Y(n4017) );
  MUX21X1_HVT U1215 ( .A1(n2474), .A2(keyout[115]), .S0(n1450), .Y(n4016) );
  MUX21X1_HVT U1216 ( .A1(n2473), .A2(keyout[115]), .S0(n1451), .Y(n4015) );
  MUX21X1_HVT U1217 ( .A1(n2472), .A2(keyout[115]), .S0(n1452), .Y(n4014) );
  MUX21X1_HVT U1218 ( .A1(n2471), .A2(keyout[115]), .S0(n1453), .Y(n4013) );
  MUX21X1_HVT U1219 ( .A1(n2470), .A2(keyout[115]), .S0(n1454), .Y(n4012) );
  MUX21X1_HVT U1220 ( .A1(n2469), .A2(keyout[116]), .S0(n1447), .Y(n4011) );
  MUX21X1_HVT U1221 ( .A1(n2468), .A2(keyout[116]), .S0(n1448), .Y(n4010) );
  MUX21X1_HVT U1222 ( .A1(n2467), .A2(keyout[116]), .S0(n1449), .Y(n4009) );
  MUX21X1_HVT U1223 ( .A1(n2466), .A2(keyout[116]), .S0(n1450), .Y(n4008) );
  MUX21X1_HVT U1224 ( .A1(n2465), .A2(keyout[116]), .S0(n1451), .Y(n4007) );
  MUX21X1_HVT U1225 ( .A1(n2464), .A2(keyout[116]), .S0(n1452), .Y(n4006) );
  MUX21X1_HVT U1226 ( .A1(n2463), .A2(keyout[116]), .S0(n1453), .Y(n4005) );
  MUX21X1_HVT U1227 ( .A1(n2462), .A2(keyout[116]), .S0(n1454), .Y(n4004) );
  MUX21X1_HVT U1228 ( .A1(n2461), .A2(keyout[117]), .S0(n1447), .Y(n4003) );
  MUX21X1_HVT U1229 ( .A1(n2460), .A2(keyout[117]), .S0(n1448), .Y(n4002) );
  MUX21X1_HVT U1230 ( .A1(n2459), .A2(keyout[117]), .S0(n1449), .Y(n4001) );
  MUX21X1_HVT U1231 ( .A1(n2458), .A2(keyout[117]), .S0(n1450), .Y(n4000) );
  MUX21X1_HVT U1232 ( .A1(n2457), .A2(keyout[117]), .S0(n1451), .Y(n3999) );
  MUX21X1_HVT U1233 ( .A1(n2456), .A2(keyout[117]), .S0(n1452), .Y(n3998) );
  MUX21X1_HVT U1234 ( .A1(n2455), .A2(keyout[117]), .S0(n1453), .Y(n3997) );
  MUX21X1_HVT U1235 ( .A1(n2454), .A2(keyout[117]), .S0(n1454), .Y(n3996) );
  MUX21X1_HVT U1236 ( .A1(n2453), .A2(keyout[118]), .S0(n1447), .Y(n3995) );
  MUX21X1_HVT U1237 ( .A1(n2452), .A2(keyout[118]), .S0(n1448), .Y(n3994) );
  MUX21X1_HVT U1238 ( .A1(n2451), .A2(keyout[118]), .S0(n1449), .Y(n3993) );
  MUX21X1_HVT U1239 ( .A1(n2450), .A2(keyout[118]), .S0(n1450), .Y(n3992) );
  MUX21X1_HVT U1240 ( .A1(n2449), .A2(keyout[118]), .S0(n1451), .Y(n3991) );
  MUX21X1_HVT U1241 ( .A1(n2448), .A2(keyout[118]), .S0(n1452), .Y(n3990) );
  MUX21X1_HVT U1242 ( .A1(n2447), .A2(keyout[118]), .S0(n1453), .Y(n3989) );
  MUX21X1_HVT U1243 ( .A1(n2446), .A2(keyout[118]), .S0(n1454), .Y(n3988) );
  MUX21X1_HVT U1244 ( .A1(n2445), .A2(keyout[119]), .S0(n1447), .Y(n3987) );
  MUX21X1_HVT U1245 ( .A1(n2444), .A2(keyout[119]), .S0(n1448), .Y(n3986) );
  MUX21X1_HVT U1246 ( .A1(n2443), .A2(keyout[119]), .S0(n1449), .Y(n3985) );
  MUX21X1_HVT U1247 ( .A1(n2442), .A2(keyout[119]), .S0(n1450), .Y(n3984) );
  MUX21X1_HVT U1248 ( .A1(n2441), .A2(keyout[119]), .S0(n1451), .Y(n3983) );
  MUX21X1_HVT U1249 ( .A1(n2440), .A2(keyout[119]), .S0(n1452), .Y(n3982) );
  MUX21X1_HVT U1250 ( .A1(n2439), .A2(keyout[119]), .S0(n1453), .Y(n3981) );
  MUX21X1_HVT U1251 ( .A1(n2438), .A2(keyout[119]), .S0(n1454), .Y(n3980) );
  MUX21X1_HVT U1252 ( .A1(n2437), .A2(keyout[120]), .S0(n1447), .Y(n3979) );
  MUX21X1_HVT U1253 ( .A1(n2436), .A2(keyout[120]), .S0(n1448), .Y(n3978) );
  MUX21X1_HVT U1254 ( .A1(n2435), .A2(keyout[120]), .S0(n1449), .Y(n3977) );
  MUX21X1_HVT U1255 ( .A1(n2434), .A2(keyout[120]), .S0(n1450), .Y(n3976) );
  MUX21X1_HVT U1256 ( .A1(n2433), .A2(keyout[120]), .S0(n1451), .Y(n3975) );
  MUX21X1_HVT U1257 ( .A1(n2432), .A2(keyout[120]), .S0(n1452), .Y(n3974) );
  MUX21X1_HVT U1258 ( .A1(n2431), .A2(keyout[120]), .S0(n1453), .Y(n3973) );
  MUX21X1_HVT U1259 ( .A1(n2430), .A2(keyout[120]), .S0(n1454), .Y(n3972) );
  MUX21X1_HVT U1260 ( .A1(n2429), .A2(keyout[121]), .S0(n1447), .Y(n3971) );
  MUX21X1_HVT U1261 ( .A1(n2428), .A2(keyout[121]), .S0(n1448), .Y(n3970) );
  MUX21X1_HVT U1262 ( .A1(n2427), .A2(keyout[121]), .S0(n1449), .Y(n3969) );
  MUX21X1_HVT U1263 ( .A1(n2426), .A2(keyout[121]), .S0(n1450), .Y(n3968) );
  MUX21X1_HVT U1264 ( .A1(n2425), .A2(keyout[121]), .S0(n1451), .Y(n3967) );
  MUX21X1_HVT U1265 ( .A1(n2424), .A2(keyout[121]), .S0(n1452), .Y(n3966) );
  MUX21X1_HVT U1266 ( .A1(n2423), .A2(keyout[121]), .S0(n1453), .Y(n3965) );
  MUX21X1_HVT U1267 ( .A1(n2422), .A2(keyout[121]), .S0(n1454), .Y(n3964) );
  MUX21X1_HVT U1268 ( .A1(n2421), .A2(keyout[122]), .S0(n1447), .Y(n3963) );
  MUX21X1_HVT U1269 ( .A1(n2420), .A2(keyout[122]), .S0(n1448), .Y(n3962) );
  MUX21X1_HVT U1270 ( .A1(n2419), .A2(keyout[122]), .S0(n1449), .Y(n3961) );
  MUX21X1_HVT U1271 ( .A1(n2418), .A2(keyout[122]), .S0(n1450), .Y(n3960) );
  MUX21X1_HVT U1272 ( .A1(n2417), .A2(keyout[122]), .S0(n1451), .Y(n3959) );
  MUX21X1_HVT U1273 ( .A1(n2416), .A2(keyout[122]), .S0(n1452), .Y(n3958) );
  MUX21X1_HVT U1274 ( .A1(n2415), .A2(keyout[122]), .S0(n1453), .Y(n3957) );
  MUX21X1_HVT U1275 ( .A1(n2414), .A2(keyout[122]), .S0(n1454), .Y(n3956) );
  MUX21X1_HVT U1276 ( .A1(n2413), .A2(keyout[123]), .S0(n1447), .Y(n3955) );
  MUX21X1_HVT U1277 ( .A1(n2412), .A2(keyout[123]), .S0(n1448), .Y(n3954) );
  MUX21X1_HVT U1278 ( .A1(n2411), .A2(keyout[123]), .S0(n1449), .Y(n3953) );
  MUX21X1_HVT U1279 ( .A1(n2410), .A2(keyout[123]), .S0(n1450), .Y(n3952) );
  MUX21X1_HVT U1280 ( .A1(n2409), .A2(keyout[123]), .S0(n1451), .Y(n3951) );
  MUX21X1_HVT U1281 ( .A1(n2408), .A2(keyout[123]), .S0(n1452), .Y(n3950) );
  MUX21X1_HVT U1282 ( .A1(n2407), .A2(keyout[123]), .S0(n1453), .Y(n3949) );
  MUX21X1_HVT U1283 ( .A1(n2406), .A2(keyout[123]), .S0(n1454), .Y(n3948) );
  MUX21X1_HVT U1284 ( .A1(n2405), .A2(keyout[124]), .S0(n1447), .Y(n3947) );
  MUX21X1_HVT U1285 ( .A1(n2404), .A2(keyout[124]), .S0(n1448), .Y(n3946) );
  MUX21X1_HVT U1286 ( .A1(n2403), .A2(keyout[124]), .S0(n1449), .Y(n3945) );
  MUX21X1_HVT U1287 ( .A1(n2402), .A2(keyout[124]), .S0(n1450), .Y(n3944) );
  MUX21X1_HVT U1288 ( .A1(n2401), .A2(keyout[124]), .S0(n1451), .Y(n3943) );
  MUX21X1_HVT U1289 ( .A1(n2400), .A2(keyout[124]), .S0(n1452), .Y(n3942) );
  MUX21X1_HVT U1290 ( .A1(n2399), .A2(keyout[124]), .S0(n1453), .Y(n3941) );
  MUX21X1_HVT U1291 ( .A1(n2398), .A2(keyout[124]), .S0(n1454), .Y(n3940) );
  MUX21X1_HVT U1292 ( .A1(n2397), .A2(keyout[125]), .S0(n1447), .Y(n3939) );
  MUX21X1_HVT U1293 ( .A1(n2396), .A2(keyout[125]), .S0(n1448), .Y(n3938) );
  MUX21X1_HVT U1294 ( .A1(n2395), .A2(keyout[125]), .S0(n1449), .Y(n3937) );
  MUX21X1_HVT U1295 ( .A1(n2394), .A2(keyout[125]), .S0(n1450), .Y(n3936) );
  MUX21X1_HVT U1296 ( .A1(n2393), .A2(keyout[125]), .S0(n1451), .Y(n3935) );
  MUX21X1_HVT U1297 ( .A1(n2392), .A2(keyout[125]), .S0(n1452), .Y(n3934) );
  MUX21X1_HVT U1298 ( .A1(n2391), .A2(keyout[125]), .S0(n1453), .Y(n3933) );
  MUX21X1_HVT U1299 ( .A1(n2390), .A2(keyout[125]), .S0(n1454), .Y(n3932) );
  MUX21X1_HVT U1300 ( .A1(n2389), .A2(keyout[126]), .S0(n1447), .Y(n3931) );
  MUX21X1_HVT U1301 ( .A1(n2388), .A2(keyout[126]), .S0(n1448), .Y(n3930) );
  MUX21X1_HVT U1302 ( .A1(n2387), .A2(keyout[126]), .S0(n1449), .Y(n3929) );
  MUX21X1_HVT U1303 ( .A1(n2386), .A2(keyout[126]), .S0(n1450), .Y(n3928) );
  MUX21X1_HVT U1304 ( .A1(n2385), .A2(keyout[126]), .S0(n1451), .Y(n3927) );
  MUX21X1_HVT U1305 ( .A1(n2384), .A2(keyout[126]), .S0(n1452), .Y(n3926) );
  MUX21X1_HVT U1306 ( .A1(n2383), .A2(keyout[126]), .S0(n1453), .Y(n3925) );
  MUX21X1_HVT U1307 ( .A1(n2382), .A2(keyout[126]), .S0(n1454), .Y(n3924) );
  MUX21X1_HVT U1308 ( .A1(n2381), .A2(keyout[127]), .S0(n1447), .Y(n3923) );
  MUX21X1_HVT U1309 ( .A1(n2380), .A2(keyout[127]), .S0(n1448), .Y(n3922) );
  NOR2X0_HVT U1310 ( .A1(n1435), .A2(rest), .Y(n1448) );
  NAND3X0_HVT U1311 ( .A1(n898), .A2(n385), .A3(n1446), .Y(n1435) );
  MUX21X1_HVT U1312 ( .A1(n2379), .A2(keyout[127]), .S0(n1449), .Y(n3921) );
  NOR2X0_HVT U1313 ( .A1(n1417), .A2(rest), .Y(n1449) );
  NAND3X0_HVT U1314 ( .A1(n3399), .A2(n1446), .A3(state[0]), .Y(n1417) );
  MUX21X1_HVT U1315 ( .A1(n2378), .A2(keyout[127]), .S0(n1450), .Y(n3920) );
  NOR2X0_HVT U1316 ( .A1(n1414), .A2(rest), .Y(n1450) );
  NAND3X0_HVT U1317 ( .A1(state[2]), .A2(n1455), .A3(state[0]), .Y(n1414) );
  MUX21X1_HVT U1318 ( .A1(n2377), .A2(keyout[127]), .S0(n1451), .Y(n3919) );
  NOR2X0_HVT U1319 ( .A1(n1432), .A2(rest), .Y(n1451) );
  NAND3X0_HVT U1320 ( .A1(n1455), .A2(n385), .A3(state[2]), .Y(n1432) );
  MUX21X1_HVT U1321 ( .A1(n2376), .A2(keyout[127]), .S0(n1452), .Y(n3918) );
  NOR2X0_HVT U1322 ( .A1(n1415), .A2(rest), .Y(n1452) );
  NAND4X0_HVT U1323 ( .A1(state[0]), .A2(n3399), .A3(state[2]), .A4(n3398), 
        .Y(n1415) );
  MUX21X1_HVT U1324 ( .A1(n2375), .A2(keyout[127]), .S0(n1453), .Y(n3917) );
  NOR2X0_HVT U1325 ( .A1(n1433), .A2(rest), .Y(n1453) );
  NAND2X0_HVT U1326 ( .A1(n1444), .A2(state[2]), .Y(n1433) );
  AND3X1_HVT U1327 ( .A1(n3398), .A2(n385), .A3(n3399), .Y(n1444) );
  MUX21X1_HVT U1328 ( .A1(n2374), .A2(keyout[127]), .S0(n1454), .Y(n3916) );
  NOR2X0_HVT U1329 ( .A1(n1442), .A2(rest), .Y(n1454) );
  NAND3X0_HVT U1330 ( .A1(n385), .A2(n899), .A3(n1455), .Y(n1442) );
  MUX21X1_HVT U1331 ( .A1(n2373), .A2(keyout[99]), .S0(n1456), .Y(n3915) );
  MUX21X1_HVT U1332 ( .A1(n2372), .A2(keyout[100]), .S0(n1456), .Y(n3914) );
  MUX21X1_HVT U1333 ( .A1(n2371), .A2(keyout[101]), .S0(n1456), .Y(n3913) );
  MUX21X1_HVT U1334 ( .A1(n2370), .A2(keyout[102]), .S0(n1456), .Y(n3912) );
  MUX21X1_HVT U1335 ( .A1(n2369), .A2(keyout[103]), .S0(n1456), .Y(n3911) );
  MUX21X1_HVT U1336 ( .A1(n2368), .A2(keyout[104]), .S0(n1456), .Y(n3910) );
  MUX21X1_HVT U1337 ( .A1(n2367), .A2(keyout[105]), .S0(n1456), .Y(n3909) );
  MUX21X1_HVT U1338 ( .A1(n2366), .A2(keyout[106]), .S0(n1456), .Y(n3908) );
  MUX21X1_HVT U1339 ( .A1(n2365), .A2(keyout[107]), .S0(n1456), .Y(n3907) );
  MUX21X1_HVT U1340 ( .A1(n2364), .A2(keyout[108]), .S0(n1456), .Y(n3906) );
  MUX21X1_HVT U1341 ( .A1(n2363), .A2(keyout[109]), .S0(n1456), .Y(n3905) );
  MUX21X1_HVT U1342 ( .A1(n2362), .A2(keyout[110]), .S0(n1456), .Y(n3904) );
  MUX21X1_HVT U1343 ( .A1(n2361), .A2(keyout[111]), .S0(n1456), .Y(n3903) );
  MUX21X1_HVT U1344 ( .A1(n2360), .A2(keyout[112]), .S0(n1456), .Y(n3902) );
  MUX21X1_HVT U1345 ( .A1(n2359), .A2(keyout[113]), .S0(n1456), .Y(n3901) );
  MUX21X1_HVT U1346 ( .A1(n2358), .A2(keyout[114]), .S0(n1456), .Y(n3900) );
  MUX21X1_HVT U1347 ( .A1(n2357), .A2(keyout[115]), .S0(n1456), .Y(n3899) );
  MUX21X1_HVT U1348 ( .A1(n2356), .A2(keyout[116]), .S0(n1456), .Y(n3898) );
  MUX21X1_HVT U1349 ( .A1(n2355), .A2(keyout[117]), .S0(n1456), .Y(n3897) );
  MUX21X1_HVT U1350 ( .A1(n2354), .A2(keyout[118]), .S0(n1456), .Y(n3896) );
  MUX21X1_HVT U1351 ( .A1(n2353), .A2(keyout[119]), .S0(n1456), .Y(n3895) );
  MUX21X1_HVT U1352 ( .A1(n2352), .A2(keyout[120]), .S0(n1456), .Y(n3894) );
  MUX21X1_HVT U1353 ( .A1(n2351), .A2(keyout[121]), .S0(n1456), .Y(n3893) );
  MUX21X1_HVT U1354 ( .A1(n2350), .A2(keyout[122]), .S0(n1456), .Y(n3892) );
  MUX21X1_HVT U1355 ( .A1(n2349), .A2(keyout[123]), .S0(n1456), .Y(n3891) );
  MUX21X1_HVT U1356 ( .A1(n2348), .A2(keyout[124]), .S0(n1456), .Y(n3890) );
  MUX21X1_HVT U1357 ( .A1(n2347), .A2(keyout[125]), .S0(n1456), .Y(n3889) );
  MUX21X1_HVT U1358 ( .A1(n2346), .A2(keyout[126]), .S0(n1456), .Y(n3888) );
  MUX21X1_HVT U1359 ( .A1(n2345), .A2(keyout[127]), .S0(n1456), .Y(n3887) );
  MUX21X1_HVT U1360 ( .A1(n2344), .A2(keyout[49]), .S0(n1456), .Y(n3886) );
  MUX21X1_HVT U1361 ( .A1(n2343), .A2(keyout[50]), .S0(n1456), .Y(n3885) );
  MUX21X1_HVT U1362 ( .A1(n2342), .A2(keyout[51]), .S0(n1456), .Y(n3884) );
  MUX21X1_HVT U1363 ( .A1(n2341), .A2(keyout[52]), .S0(n1456), .Y(n3883) );
  MUX21X1_HVT U1364 ( .A1(n2340), .A2(keyout[53]), .S0(n1456), .Y(n3882) );
  MUX21X1_HVT U1365 ( .A1(n2339), .A2(keyout[54]), .S0(n1456), .Y(n3881) );
  MUX21X1_HVT U1366 ( .A1(n2338), .A2(keyout[55]), .S0(n1456), .Y(n3880) );
  MUX21X1_HVT U1367 ( .A1(n2337), .A2(keyout[56]), .S0(n1456), .Y(n3879) );
  MUX21X1_HVT U1368 ( .A1(n2336), .A2(keyout[57]), .S0(n1456), .Y(n3878) );
  MUX21X1_HVT U1369 ( .A1(n2335), .A2(keyout[58]), .S0(n1456), .Y(n3877) );
  MUX21X1_HVT U1370 ( .A1(n2334), .A2(keyout[59]), .S0(n1456), .Y(n3876) );
  MUX21X1_HVT U1371 ( .A1(n2333), .A2(keyout[60]), .S0(n1456), .Y(n3875) );
  MUX21X1_HVT U1372 ( .A1(n2332), .A2(keyout[61]), .S0(n1456), .Y(n3874) );
  MUX21X1_HVT U1373 ( .A1(n2331), .A2(keyout[62]), .S0(n1456), .Y(n3873) );
  MUX21X1_HVT U1374 ( .A1(n2330), .A2(keyout[63]), .S0(n1456), .Y(n3872) );
  MUX21X1_HVT U1375 ( .A1(n2329), .A2(keyout[64]), .S0(n1456), .Y(n3871) );
  MUX21X1_HVT U1376 ( .A1(n2328), .A2(keyout[65]), .S0(n1456), .Y(n3870) );
  MUX21X1_HVT U1377 ( .A1(n2327), .A2(keyout[66]), .S0(n1456), .Y(n3869) );
  MUX21X1_HVT U1378 ( .A1(n2326), .A2(keyout[67]), .S0(n1456), .Y(n3868) );
  MUX21X1_HVT U1379 ( .A1(n2325), .A2(keyout[68]), .S0(n1456), .Y(n3867) );
  MUX21X1_HVT U1380 ( .A1(n2324), .A2(keyout[69]), .S0(n1456), .Y(n3866) );
  MUX21X1_HVT U1381 ( .A1(n2323), .A2(keyout[70]), .S0(n1456), .Y(n3865) );
  MUX21X1_HVT U1382 ( .A1(n2322), .A2(keyout[71]), .S0(n1456), .Y(n3864) );
  MUX21X1_HVT U1383 ( .A1(n2321), .A2(keyout[72]), .S0(n1456), .Y(n3863) );
  MUX21X1_HVT U1384 ( .A1(n2320), .A2(keyout[73]), .S0(n1456), .Y(n3862) );
  MUX21X1_HVT U1385 ( .A1(n2319), .A2(keyout[74]), .S0(n1456), .Y(n3861) );
  MUX21X1_HVT U1386 ( .A1(n2318), .A2(keyout[75]), .S0(n1456), .Y(n3860) );
  MUX21X1_HVT U1387 ( .A1(n2317), .A2(keyout[76]), .S0(n1456), .Y(n3859) );
  MUX21X1_HVT U1388 ( .A1(n2316), .A2(keyout[77]), .S0(n1456), .Y(n3858) );
  MUX21X1_HVT U1389 ( .A1(n2315), .A2(keyout[78]), .S0(n1456), .Y(n3857) );
  MUX21X1_HVT U1390 ( .A1(n2314), .A2(keyout[79]), .S0(n1456), .Y(n3856) );
  MUX21X1_HVT U1391 ( .A1(n2313), .A2(keyout[80]), .S0(n1456), .Y(n3855) );
  MUX21X1_HVT U1392 ( .A1(n2312), .A2(keyout[81]), .S0(n1456), .Y(n3854) );
  MUX21X1_HVT U1393 ( .A1(n2311), .A2(keyout[82]), .S0(n1456), .Y(n3853) );
  MUX21X1_HVT U1394 ( .A1(n2310), .A2(keyout[83]), .S0(n1456), .Y(n3852) );
  MUX21X1_HVT U1395 ( .A1(n2309), .A2(keyout[84]), .S0(n1456), .Y(n3851) );
  MUX21X1_HVT U1396 ( .A1(n2308), .A2(keyout[85]), .S0(n1456), .Y(n3850) );
  MUX21X1_HVT U1397 ( .A1(n2307), .A2(keyout[86]), .S0(n1456), .Y(n3849) );
  MUX21X1_HVT U1398 ( .A1(n2306), .A2(keyout[87]), .S0(n1456), .Y(n3848) );
  MUX21X1_HVT U1399 ( .A1(n2305), .A2(keyout[88]), .S0(n1456), .Y(n3847) );
  MUX21X1_HVT U1400 ( .A1(n2304), .A2(keyout[89]), .S0(n1456), .Y(n3846) );
  MUX21X1_HVT U1401 ( .A1(n2303), .A2(keyout[90]), .S0(n1456), .Y(n3845) );
  MUX21X1_HVT U1402 ( .A1(n2302), .A2(keyout[91]), .S0(n1456), .Y(n3844) );
  MUX21X1_HVT U1403 ( .A1(n2301), .A2(keyout[92]), .S0(n1456), .Y(n3843) );
  MUX21X1_HVT U1404 ( .A1(n2300), .A2(keyout[93]), .S0(n1456), .Y(n3842) );
  MUX21X1_HVT U1405 ( .A1(n2299), .A2(keyout[94]), .S0(n1456), .Y(n3841) );
  MUX21X1_HVT U1406 ( .A1(n2298), .A2(keyout[95]), .S0(n1456), .Y(n3840) );
  MUX21X1_HVT U1407 ( .A1(n2297), .A2(keyout[96]), .S0(n1456), .Y(n3839) );
  MUX21X1_HVT U1408 ( .A1(n2296), .A2(keyout[97]), .S0(n1456), .Y(n3838) );
  MUX21X1_HVT U1409 ( .A1(n2295), .A2(keyout[0]), .S0(n1456), .Y(n3837) );
  MUX21X1_HVT U1410 ( .A1(n2294), .A2(keyout[1]), .S0(n1456), .Y(n3836) );
  MUX21X1_HVT U1411 ( .A1(n2293), .A2(keyout[2]), .S0(n1456), .Y(n3835) );
  MUX21X1_HVT U1412 ( .A1(n2292), .A2(keyout[3]), .S0(n1456), .Y(n3834) );
  MUX21X1_HVT U1413 ( .A1(n2291), .A2(keyout[4]), .S0(n1456), .Y(n3833) );
  MUX21X1_HVT U1414 ( .A1(n2290), .A2(keyout[5]), .S0(n1456), .Y(n3832) );
  MUX21X1_HVT U1415 ( .A1(n2289), .A2(keyout[6]), .S0(n1456), .Y(n3831) );
  MUX21X1_HVT U1416 ( .A1(n2288), .A2(keyout[7]), .S0(n1456), .Y(n3830) );
  MUX21X1_HVT U1417 ( .A1(n2287), .A2(keyout[8]), .S0(n1456), .Y(n3829) );
  MUX21X1_HVT U1418 ( .A1(n2286), .A2(keyout[9]), .S0(n1456), .Y(n3828) );
  MUX21X1_HVT U1419 ( .A1(n2285), .A2(keyout[10]), .S0(n1456), .Y(n3827) );
  MUX21X1_HVT U1420 ( .A1(n2284), .A2(keyout[11]), .S0(n1456), .Y(n3826) );
  MUX21X1_HVT U1421 ( .A1(n2283), .A2(keyout[12]), .S0(n1456), .Y(n3825) );
  MUX21X1_HVT U1422 ( .A1(n2282), .A2(keyout[13]), .S0(n1456), .Y(n3824) );
  MUX21X1_HVT U1423 ( .A1(n2281), .A2(keyout[14]), .S0(n1456), .Y(n3823) );
  MUX21X1_HVT U1424 ( .A1(n2280), .A2(keyout[15]), .S0(n1456), .Y(n3822) );
  MUX21X1_HVT U1425 ( .A1(n2279), .A2(keyout[16]), .S0(n1456), .Y(n3821) );
  MUX21X1_HVT U1426 ( .A1(n2278), .A2(keyout[17]), .S0(n1456), .Y(n3820) );
  MUX21X1_HVT U1427 ( .A1(n2277), .A2(keyout[18]), .S0(n1456), .Y(n3819) );
  MUX21X1_HVT U1428 ( .A1(n2276), .A2(keyout[19]), .S0(n1456), .Y(n3818) );
  MUX21X1_HVT U1429 ( .A1(n2275), .A2(keyout[20]), .S0(n1456), .Y(n3817) );
  MUX21X1_HVT U1430 ( .A1(n2274), .A2(keyout[21]), .S0(n1456), .Y(n3816) );
  MUX21X1_HVT U1431 ( .A1(n2273), .A2(keyout[22]), .S0(n1456), .Y(n3815) );
  MUX21X1_HVT U1432 ( .A1(n2272), .A2(keyout[23]), .S0(n1456), .Y(n3814) );
  MUX21X1_HVT U1433 ( .A1(n2271), .A2(keyout[24]), .S0(n1456), .Y(n3813) );
  MUX21X1_HVT U1434 ( .A1(n2270), .A2(keyout[25]), .S0(n1456), .Y(n3812) );
  MUX21X1_HVT U1435 ( .A1(n2269), .A2(keyout[26]), .S0(n1456), .Y(n3811) );
  MUX21X1_HVT U1436 ( .A1(n2268), .A2(keyout[27]), .S0(n1456), .Y(n3810) );
  MUX21X1_HVT U1437 ( .A1(n2267), .A2(keyout[28]), .S0(n1456), .Y(n3809) );
  MUX21X1_HVT U1438 ( .A1(n2266), .A2(keyout[29]), .S0(n1456), .Y(n3808) );
  MUX21X1_HVT U1439 ( .A1(n2265), .A2(keyout[30]), .S0(n1456), .Y(n3807) );
  MUX21X1_HVT U1440 ( .A1(n2264), .A2(keyout[31]), .S0(n1456), .Y(n3806) );
  MUX21X1_HVT U1441 ( .A1(n2263), .A2(keyout[32]), .S0(n1456), .Y(n3805) );
  MUX21X1_HVT U1442 ( .A1(n2262), .A2(keyout[33]), .S0(n1456), .Y(n3804) );
  MUX21X1_HVT U1443 ( .A1(n2261), .A2(keyout[34]), .S0(n1456), .Y(n3803) );
  MUX21X1_HVT U1444 ( .A1(n2260), .A2(keyout[35]), .S0(n1456), .Y(n3802) );
  MUX21X1_HVT U1445 ( .A1(n2259), .A2(keyout[48]), .S0(n1456), .Y(n3801) );
  MUX21X1_HVT U1446 ( .A1(n2258), .A2(keyout[47]), .S0(n1456), .Y(n3800) );
  MUX21X1_HVT U1447 ( .A1(n2257), .A2(keyout[46]), .S0(n1456), .Y(n3799) );
  MUX21X1_HVT U1448 ( .A1(n2256), .A2(keyout[45]), .S0(n1456), .Y(n3798) );
  MUX21X1_HVT U1449 ( .A1(n2255), .A2(keyout[44]), .S0(n1456), .Y(n3797) );
  MUX21X1_HVT U1450 ( .A1(n2254), .A2(keyout[43]), .S0(n1456), .Y(n3796) );
  MUX21X1_HVT U1451 ( .A1(n2253), .A2(keyout[42]), .S0(n1456), .Y(n3795) );
  MUX21X1_HVT U1452 ( .A1(n2252), .A2(keyout[41]), .S0(n1456), .Y(n3794) );
  MUX21X1_HVT U1453 ( .A1(n2251), .A2(keyout[40]), .S0(n1456), .Y(n3793) );
  MUX21X1_HVT U1454 ( .A1(n2250), .A2(keyout[39]), .S0(n1456), .Y(n3792) );
  MUX21X1_HVT U1455 ( .A1(n2249), .A2(keyout[38]), .S0(n1456), .Y(n3791) );
  MUX21X1_HVT U1456 ( .A1(n2247), .A2(keyout[37]), .S0(n1456), .Y(n3790) );
  MUX21X1_HVT U1457 ( .A1(n2245), .A2(keyout[36]), .S0(n1456), .Y(n3789) );
  MUX21X1_HVT U1458 ( .A1(n2243), .A2(keyout[98]), .S0(n1456), .Y(n3788) );
  NOR2X0_HVT U1459 ( .A1(n1422), .A2(rest), .Y(n1456) );
  NAND3X0_HVT U1460 ( .A1(n1455), .A2(n899), .A3(state[0]), .Y(n1422) );
  AND2X1_HVT U1461 ( .A1(n3398), .A2(n898), .Y(n1455) );
  MUX21X1_HVT U1462 ( .A1(n2241), .A2(keyout[99]), .S0(n1457), .Y(n3787) );
  NAND4X0_HVT U1463 ( .A1(n1458), .A2(n1459), .A3(n1460), .A4(n1461), .Y(n3786) );
  OA222X1_HVT U1464 ( .A1(n1028), .A2(n1462), .A3(n128), .A4(n1463), .A5(n641), 
        .A6(n1464), .Y(n1461) );
  OA222X1_HVT U1465 ( .A1(n1029), .A2(n1465), .A3(n129), .A4(n1466), .A5(n642), 
        .A6(n1467), .Y(n1460) );
  OA222X1_HVT U1466 ( .A1(n1030), .A2(n1468), .A3(n130), .A4(n1469), .A5(n643), 
        .A6(n1470), .Y(n1459) );
  OA222X1_HVT U1467 ( .A1(n2248), .A2(n1447), .A3(n386), .A4(n1471), .A5(n900), 
        .A6(n1472), .Y(n1458) );
  MUX21X1_HVT U1468 ( .A1(n2239), .A2(keyout[100]), .S0(n1457), .Y(n3785) );
  NAND4X0_HVT U1469 ( .A1(n1473), .A2(n1474), .A3(n1475), .A4(n1476), .Y(n3784) );
  OA222X1_HVT U1470 ( .A1(n1031), .A2(n1462), .A3(n131), .A4(n1463), .A5(n644), 
        .A6(n1464), .Y(n1476) );
  OA222X1_HVT U1471 ( .A1(n1032), .A2(n1465), .A3(n132), .A4(n1466), .A5(n645), 
        .A6(n1467), .Y(n1475) );
  OA222X1_HVT U1472 ( .A1(n1033), .A2(n1468), .A3(n387), .A4(n1469), .A5(n1470), .A6(n1), .Y(n1474) );
  OA222X1_HVT U1473 ( .A1(n2246), .A2(n1447), .A3(n388), .A4(n1471), .A5(n901), 
        .A6(n1472), .Y(n1473) );
  MUX21X1_HVT U1474 ( .A1(n2237), .A2(keyout[101]), .S0(n1457), .Y(n3783) );
  NAND4X0_HVT U1475 ( .A1(n1477), .A2(n1478), .A3(n1479), .A4(n1480), .Y(n3782) );
  OA222X1_HVT U1476 ( .A1(n1034), .A2(n1462), .A3(n133), .A4(n1463), .A5(n646), 
        .A6(n1464), .Y(n1480) );
  OA222X1_HVT U1477 ( .A1(n1035), .A2(n1465), .A3(n134), .A4(n1466), .A5(n647), 
        .A6(n1467), .Y(n1479) );
  OA222X1_HVT U1478 ( .A1(n1036), .A2(n1468), .A3(n389), .A4(n1469), .A5(n1470), .A6(n2), .Y(n1478) );
  OA222X1_HVT U1479 ( .A1(n2244), .A2(n1447), .A3(n390), .A4(n1471), .A5(n902), 
        .A6(n1472), .Y(n1477) );
  MUX21X1_HVT U1480 ( .A1(n2235), .A2(keyout[102]), .S0(n1457), .Y(n3781) );
  NAND4X0_HVT U1481 ( .A1(n1481), .A2(n1482), .A3(n1483), .A4(n1484), .Y(n3780) );
  OA222X1_HVT U1482 ( .A1(n1037), .A2(n1462), .A3(n135), .A4(n1463), .A5(n648), 
        .A6(n1464), .Y(n1484) );
  OA222X1_HVT U1483 ( .A1(n1038), .A2(n1465), .A3(n136), .A4(n1466), .A5(n649), 
        .A6(n1467), .Y(n1483) );
  OA222X1_HVT U1484 ( .A1(n1039), .A2(n1468), .A3(n391), .A4(n1469), .A5(n1470), .A6(n3), .Y(n1482) );
  OA222X1_HVT U1485 ( .A1(n2242), .A2(n1447), .A3(n392), .A4(n1471), .A5(n903), 
        .A6(n1472), .Y(n1481) );
  MUX21X1_HVT U1486 ( .A1(n2233), .A2(keyout[103]), .S0(n1457), .Y(n3779) );
  NAND4X0_HVT U1487 ( .A1(n1485), .A2(n1486), .A3(n1487), .A4(n1488), .Y(n3778) );
  OA222X1_HVT U1488 ( .A1(n1040), .A2(n1462), .A3(n137), .A4(n1463), .A5(n650), 
        .A6(n1464), .Y(n1488) );
  OA222X1_HVT U1489 ( .A1(n1041), .A2(n1465), .A3(n138), .A4(n1466), .A5(n651), 
        .A6(n1467), .Y(n1487) );
  OA222X1_HVT U1490 ( .A1(n1042), .A2(n1468), .A3(n393), .A4(n1469), .A5(n1470), .A6(n4), .Y(n1486) );
  OA222X1_HVT U1491 ( .A1(n2240), .A2(n1447), .A3(n394), .A4(n1471), .A5(n904), 
        .A6(n1472), .Y(n1485) );
  MUX21X1_HVT U1492 ( .A1(n2231), .A2(keyout[104]), .S0(n1457), .Y(n3777) );
  NAND4X0_HVT U1493 ( .A1(n1489), .A2(n1490), .A3(n1491), .A4(n1492), .Y(n3776) );
  OA222X1_HVT U1494 ( .A1(n1043), .A2(n1462), .A3(n139), .A4(n1463), .A5(n652), 
        .A6(n1464), .Y(n1492) );
  OA222X1_HVT U1495 ( .A1(n1044), .A2(n1465), .A3(n140), .A4(n1466), .A5(n653), 
        .A6(n1467), .Y(n1491) );
  OA222X1_HVT U1496 ( .A1(n1045), .A2(n1468), .A3(n395), .A4(n1469), .A5(n1470), .A6(n5), .Y(n1490) );
  OA222X1_HVT U1497 ( .A1(n2238), .A2(n1447), .A3(n396), .A4(n1471), .A5(n905), 
        .A6(n1472), .Y(n1489) );
  MUX21X1_HVT U1498 ( .A1(n2229), .A2(keyout[105]), .S0(n1457), .Y(n3775) );
  NAND4X0_HVT U1499 ( .A1(n1493), .A2(n1494), .A3(n1495), .A4(n1496), .Y(n3774) );
  OA222X1_HVT U1500 ( .A1(n1046), .A2(n1462), .A3(n141), .A4(n1463), .A5(n654), 
        .A6(n1464), .Y(n1496) );
  OA222X1_HVT U1501 ( .A1(n1047), .A2(n1465), .A3(n142), .A4(n1466), .A5(n655), 
        .A6(n1467), .Y(n1495) );
  OA222X1_HVT U1502 ( .A1(n1048), .A2(n1468), .A3(n397), .A4(n1469), .A5(n1470), .A6(n6), .Y(n1494) );
  OA222X1_HVT U1503 ( .A1(n2236), .A2(n1447), .A3(n398), .A4(n1471), .A5(n906), 
        .A6(n1472), .Y(n1493) );
  MUX21X1_HVT U1504 ( .A1(n2227), .A2(keyout[106]), .S0(n1457), .Y(n3773) );
  NAND4X0_HVT U1505 ( .A1(n1497), .A2(n1498), .A3(n1499), .A4(n1500), .Y(n3772) );
  OA222X1_HVT U1506 ( .A1(n1049), .A2(n1462), .A3(n143), .A4(n1463), .A5(n656), 
        .A6(n1464), .Y(n1500) );
  OA222X1_HVT U1507 ( .A1(n1050), .A2(n1465), .A3(n144), .A4(n1466), .A5(n657), 
        .A6(n1467), .Y(n1499) );
  OA222X1_HVT U1508 ( .A1(n1051), .A2(n1468), .A3(n399), .A4(n1469), .A5(n1470), .A6(n7), .Y(n1498) );
  OA222X1_HVT U1509 ( .A1(n2234), .A2(n1447), .A3(n400), .A4(n1471), .A5(n907), 
        .A6(n1472), .Y(n1497) );
  MUX21X1_HVT U1510 ( .A1(n2225), .A2(keyout[107]), .S0(n1457), .Y(n3771) );
  NAND4X0_HVT U1511 ( .A1(n1501), .A2(n1502), .A3(n1503), .A4(n1504), .Y(n3770) );
  OA222X1_HVT U1512 ( .A1(n1052), .A2(n1462), .A3(n145), .A4(n1463), .A5(n658), 
        .A6(n1464), .Y(n1504) );
  OA222X1_HVT U1513 ( .A1(n1053), .A2(n1465), .A3(n146), .A4(n1466), .A5(n659), 
        .A6(n1467), .Y(n1503) );
  OA222X1_HVT U1514 ( .A1(n1054), .A2(n1468), .A3(n401), .A4(n1469), .A5(n1470), .A6(n8), .Y(n1502) );
  OA222X1_HVT U1515 ( .A1(n2232), .A2(n1447), .A3(n402), .A4(n1471), .A5(n908), 
        .A6(n1472), .Y(n1501) );
  MUX21X1_HVT U1516 ( .A1(n2223), .A2(keyout[108]), .S0(n1457), .Y(n3769) );
  NAND4X0_HVT U1517 ( .A1(n1505), .A2(n1506), .A3(n1507), .A4(n1508), .Y(n3768) );
  OA222X1_HVT U1518 ( .A1(n1055), .A2(n1462), .A3(n147), .A4(n1463), .A5(n660), 
        .A6(n1464), .Y(n1508) );
  OA222X1_HVT U1519 ( .A1(n1056), .A2(n1465), .A3(n148), .A4(n1466), .A5(n661), 
        .A6(n1467), .Y(n1507) );
  OA222X1_HVT U1520 ( .A1(n1057), .A2(n1468), .A3(n403), .A4(n1469), .A5(n1470), .A6(n9), .Y(n1506) );
  OA222X1_HVT U1521 ( .A1(n2230), .A2(n1447), .A3(n404), .A4(n1471), .A5(n909), 
        .A6(n1472), .Y(n1505) );
  MUX21X1_HVT U1522 ( .A1(n2221), .A2(keyout[109]), .S0(n1457), .Y(n3767) );
  NAND4X0_HVT U1523 ( .A1(n1509), .A2(n1510), .A3(n1511), .A4(n1512), .Y(n3766) );
  OA222X1_HVT U1524 ( .A1(n1058), .A2(n1462), .A3(n149), .A4(n1463), .A5(n662), 
        .A6(n1464), .Y(n1512) );
  OA222X1_HVT U1525 ( .A1(n1059), .A2(n1465), .A3(n150), .A4(n1466), .A5(n663), 
        .A6(n1467), .Y(n1511) );
  OA222X1_HVT U1526 ( .A1(n1060), .A2(n1468), .A3(n405), .A4(n1469), .A5(n1470), .A6(n10), .Y(n1510) );
  OA222X1_HVT U1527 ( .A1(n2228), .A2(n1447), .A3(n406), .A4(n1471), .A5(n910), 
        .A6(n1472), .Y(n1509) );
  MUX21X1_HVT U1528 ( .A1(n2219), .A2(keyout[110]), .S0(n1457), .Y(n3765) );
  NAND4X0_HVT U1529 ( .A1(n1513), .A2(n1514), .A3(n1515), .A4(n1516), .Y(n3764) );
  OA222X1_HVT U1530 ( .A1(n1061), .A2(n1462), .A3(n151), .A4(n1463), .A5(n664), 
        .A6(n1464), .Y(n1516) );
  OA222X1_HVT U1531 ( .A1(n1062), .A2(n1465), .A3(n152), .A4(n1466), .A5(n665), 
        .A6(n1467), .Y(n1515) );
  OA222X1_HVT U1532 ( .A1(n1063), .A2(n1468), .A3(n407), .A4(n1469), .A5(n1470), .A6(n11), .Y(n1514) );
  OA222X1_HVT U1533 ( .A1(n2226), .A2(n1447), .A3(n408), .A4(n1471), .A5(n911), 
        .A6(n1472), .Y(n1513) );
  MUX21X1_HVT U1534 ( .A1(n2217), .A2(keyout[111]), .S0(n1457), .Y(n3763) );
  NAND4X0_HVT U1535 ( .A1(n1517), .A2(n1518), .A3(n1519), .A4(n1520), .Y(n3762) );
  OA222X1_HVT U1536 ( .A1(n1064), .A2(n1462), .A3(n153), .A4(n1463), .A5(n666), 
        .A6(n1464), .Y(n1520) );
  OA222X1_HVT U1537 ( .A1(n1065), .A2(n1465), .A3(n154), .A4(n1466), .A5(n667), 
        .A6(n1467), .Y(n1519) );
  OA222X1_HVT U1538 ( .A1(n1066), .A2(n1468), .A3(n409), .A4(n1469), .A5(n1470), .A6(n12), .Y(n1518) );
  OA222X1_HVT U1539 ( .A1(n2224), .A2(n1447), .A3(n410), .A4(n1471), .A5(n912), 
        .A6(n1472), .Y(n1517) );
  MUX21X1_HVT U1540 ( .A1(n2215), .A2(keyout[112]), .S0(n1457), .Y(n3761) );
  NAND4X0_HVT U1541 ( .A1(n1521), .A2(n1522), .A3(n1523), .A4(n1524), .Y(n3760) );
  OA222X1_HVT U1542 ( .A1(n1067), .A2(n1462), .A3(n155), .A4(n1463), .A5(n668), 
        .A6(n1464), .Y(n1524) );
  OA222X1_HVT U1543 ( .A1(n1068), .A2(n1465), .A3(n156), .A4(n1466), .A5(n669), 
        .A6(n1467), .Y(n1523) );
  OA222X1_HVT U1544 ( .A1(n1069), .A2(n1468), .A3(n411), .A4(n1469), .A5(n1470), .A6(n13), .Y(n1522) );
  OA222X1_HVT U1545 ( .A1(n2222), .A2(n1447), .A3(n412), .A4(n1471), .A5(n913), 
        .A6(n1472), .Y(n1521) );
  MUX21X1_HVT U1546 ( .A1(n2213), .A2(keyout[113]), .S0(n1457), .Y(n3759) );
  NAND4X0_HVT U1547 ( .A1(n1525), .A2(n1526), .A3(n1527), .A4(n1528), .Y(n3758) );
  OA222X1_HVT U1548 ( .A1(n1070), .A2(n1462), .A3(n157), .A4(n1463), .A5(n670), 
        .A6(n1464), .Y(n1528) );
  OA222X1_HVT U1549 ( .A1(n1071), .A2(n1465), .A3(n158), .A4(n1466), .A5(n671), 
        .A6(n1467), .Y(n1527) );
  OA222X1_HVT U1550 ( .A1(n1072), .A2(n1468), .A3(n413), .A4(n1469), .A5(n1470), .A6(n14), .Y(n1526) );
  OA222X1_HVT U1551 ( .A1(n2220), .A2(n1447), .A3(n414), .A4(n1471), .A5(n914), 
        .A6(n1472), .Y(n1525) );
  MUX21X1_HVT U1552 ( .A1(n2211), .A2(keyout[114]), .S0(n1457), .Y(n3757) );
  NAND4X0_HVT U1553 ( .A1(n1529), .A2(n1530), .A3(n1531), .A4(n1532), .Y(n3756) );
  OA222X1_HVT U1554 ( .A1(n1073), .A2(n1462), .A3(n159), .A4(n1463), .A5(n672), 
        .A6(n1464), .Y(n1532) );
  OA222X1_HVT U1555 ( .A1(n1074), .A2(n1465), .A3(n160), .A4(n1466), .A5(n673), 
        .A6(n1467), .Y(n1531) );
  OA222X1_HVT U1556 ( .A1(n1075), .A2(n1468), .A3(n415), .A4(n1469), .A5(n1470), .A6(n15), .Y(n1530) );
  OA222X1_HVT U1557 ( .A1(n2218), .A2(n1447), .A3(n416), .A4(n1471), .A5(n915), 
        .A6(n1472), .Y(n1529) );
  MUX21X1_HVT U1558 ( .A1(n2209), .A2(keyout[115]), .S0(n1457), .Y(n3755) );
  NAND4X0_HVT U1559 ( .A1(n1533), .A2(n1534), .A3(n1535), .A4(n1536), .Y(n3754) );
  OA222X1_HVT U1560 ( .A1(n1076), .A2(n1462), .A3(n161), .A4(n1463), .A5(n674), 
        .A6(n1464), .Y(n1536) );
  OA222X1_HVT U1561 ( .A1(n1077), .A2(n1465), .A3(n162), .A4(n1466), .A5(n675), 
        .A6(n1467), .Y(n1535) );
  OA222X1_HVT U1562 ( .A1(n1078), .A2(n1468), .A3(n417), .A4(n1469), .A5(n1470), .A6(n16), .Y(n1534) );
  OA222X1_HVT U1563 ( .A1(n2216), .A2(n1447), .A3(n418), .A4(n1471), .A5(n916), 
        .A6(n1472), .Y(n1533) );
  MUX21X1_HVT U1564 ( .A1(n2207), .A2(keyout[116]), .S0(n1457), .Y(n3753) );
  NAND4X0_HVT U1565 ( .A1(n1537), .A2(n1538), .A3(n1539), .A4(n1540), .Y(n3752) );
  OA222X1_HVT U1566 ( .A1(n1079), .A2(n1462), .A3(n163), .A4(n1463), .A5(n676), 
        .A6(n1464), .Y(n1540) );
  OA222X1_HVT U1567 ( .A1(n1080), .A2(n1465), .A3(n164), .A4(n1466), .A5(n677), 
        .A6(n1467), .Y(n1539) );
  OA222X1_HVT U1568 ( .A1(n1081), .A2(n1468), .A3(n419), .A4(n1469), .A5(n1470), .A6(n17), .Y(n1538) );
  OA222X1_HVT U1569 ( .A1(n2214), .A2(n1447), .A3(n420), .A4(n1471), .A5(n917), 
        .A6(n1472), .Y(n1537) );
  MUX21X1_HVT U1570 ( .A1(n2205), .A2(keyout[117]), .S0(n1457), .Y(n3751) );
  NAND4X0_HVT U1571 ( .A1(n1541), .A2(n1542), .A3(n1543), .A4(n1544), .Y(n3750) );
  OA222X1_HVT U1572 ( .A1(n1082), .A2(n1462), .A3(n165), .A4(n1463), .A5(n678), 
        .A6(n1464), .Y(n1544) );
  OA222X1_HVT U1573 ( .A1(n1083), .A2(n1465), .A3(n166), .A4(n1466), .A5(n679), 
        .A6(n1467), .Y(n1543) );
  OA222X1_HVT U1574 ( .A1(n1084), .A2(n1468), .A3(n421), .A4(n1469), .A5(n1470), .A6(n18), .Y(n1542) );
  OA222X1_HVT U1575 ( .A1(n2212), .A2(n1447), .A3(n422), .A4(n1471), .A5(n918), 
        .A6(n1472), .Y(n1541) );
  MUX21X1_HVT U1576 ( .A1(n2203), .A2(keyout[118]), .S0(n1457), .Y(n3749) );
  NAND4X0_HVT U1577 ( .A1(n1545), .A2(n1546), .A3(n1547), .A4(n1548), .Y(n3748) );
  OA222X1_HVT U1578 ( .A1(n1085), .A2(n1462), .A3(n167), .A4(n1463), .A5(n680), 
        .A6(n1464), .Y(n1548) );
  OA222X1_HVT U1579 ( .A1(n1086), .A2(n1465), .A3(n168), .A4(n1466), .A5(n681), 
        .A6(n1467), .Y(n1547) );
  OA222X1_HVT U1580 ( .A1(n1087), .A2(n1468), .A3(n423), .A4(n1469), .A5(n1470), .A6(n19), .Y(n1546) );
  OA222X1_HVT U1581 ( .A1(n2210), .A2(n1447), .A3(n424), .A4(n1471), .A5(n919), 
        .A6(n1472), .Y(n1545) );
  MUX21X1_HVT U1582 ( .A1(n2201), .A2(keyout[119]), .S0(n1457), .Y(n3747) );
  NAND4X0_HVT U1583 ( .A1(n1549), .A2(n1550), .A3(n1551), .A4(n1552), .Y(n3746) );
  OA222X1_HVT U1584 ( .A1(n1088), .A2(n1462), .A3(n169), .A4(n1463), .A5(n682), 
        .A6(n1464), .Y(n1552) );
  OA222X1_HVT U1585 ( .A1(n1089), .A2(n1465), .A3(n170), .A4(n1466), .A5(n683), 
        .A6(n1467), .Y(n1551) );
  OA222X1_HVT U1586 ( .A1(n1090), .A2(n1468), .A3(n425), .A4(n1469), .A5(n1470), .A6(n20), .Y(n1550) );
  OA222X1_HVT U1587 ( .A1(n2208), .A2(n1447), .A3(n426), .A4(n1471), .A5(n920), 
        .A6(n1472), .Y(n1549) );
  MUX21X1_HVT U1588 ( .A1(n2199), .A2(keyout[120]), .S0(n1457), .Y(n3745) );
  NAND4X0_HVT U1589 ( .A1(n1553), .A2(n1554), .A3(n1555), .A4(n1556), .Y(n3744) );
  OA222X1_HVT U1590 ( .A1(n1091), .A2(n1462), .A3(n171), .A4(n1463), .A5(n684), 
        .A6(n1464), .Y(n1556) );
  OA222X1_HVT U1591 ( .A1(n1092), .A2(n1465), .A3(n172), .A4(n1466), .A5(n685), 
        .A6(n1467), .Y(n1555) );
  OA222X1_HVT U1592 ( .A1(n1093), .A2(n1468), .A3(n427), .A4(n1469), .A5(n1470), .A6(n21), .Y(n1554) );
  OA222X1_HVT U1593 ( .A1(n2206), .A2(n1447), .A3(n428), .A4(n1471), .A5(n921), 
        .A6(n1472), .Y(n1553) );
  MUX21X1_HVT U1594 ( .A1(n2197), .A2(keyout[121]), .S0(n1457), .Y(n3743) );
  NAND4X0_HVT U1595 ( .A1(n1557), .A2(n1558), .A3(n1559), .A4(n1560), .Y(n3742) );
  OA222X1_HVT U1596 ( .A1(n1094), .A2(n1462), .A3(n173), .A4(n1463), .A5(n686), 
        .A6(n1464), .Y(n1560) );
  OA222X1_HVT U1597 ( .A1(n1095), .A2(n1465), .A3(n174), .A4(n1466), .A5(n687), 
        .A6(n1467), .Y(n1559) );
  OA222X1_HVT U1598 ( .A1(n1096), .A2(n1468), .A3(n429), .A4(n1469), .A5(n1470), .A6(n22), .Y(n1558) );
  OA222X1_HVT U1599 ( .A1(n2204), .A2(n1447), .A3(n430), .A4(n1471), .A5(n922), 
        .A6(n1472), .Y(n1557) );
  MUX21X1_HVT U1600 ( .A1(n2195), .A2(keyout[122]), .S0(n1457), .Y(n3741) );
  NAND4X0_HVT U1601 ( .A1(n1561), .A2(n1562), .A3(n1563), .A4(n1564), .Y(n3740) );
  OA222X1_HVT U1602 ( .A1(n1097), .A2(n1462), .A3(n175), .A4(n1463), .A5(n688), 
        .A6(n1464), .Y(n1564) );
  OA222X1_HVT U1603 ( .A1(n1098), .A2(n1465), .A3(n176), .A4(n1466), .A5(n689), 
        .A6(n1467), .Y(n1563) );
  OA222X1_HVT U1604 ( .A1(n1099), .A2(n1468), .A3(n431), .A4(n1469), .A5(n1470), .A6(n23), .Y(n1562) );
  OA222X1_HVT U1605 ( .A1(n2202), .A2(n1447), .A3(n432), .A4(n1471), .A5(n923), 
        .A6(n1472), .Y(n1561) );
  MUX21X1_HVT U1606 ( .A1(n2193), .A2(keyout[123]), .S0(n1457), .Y(n3739) );
  NAND4X0_HVT U1607 ( .A1(n1565), .A2(n1566), .A3(n1567), .A4(n1568), .Y(n3738) );
  OA222X1_HVT U1608 ( .A1(n1100), .A2(n1462), .A3(n177), .A4(n1463), .A5(n690), 
        .A6(n1464), .Y(n1568) );
  OA222X1_HVT U1609 ( .A1(n1101), .A2(n1465), .A3(n178), .A4(n1466), .A5(n691), 
        .A6(n1467), .Y(n1567) );
  OA222X1_HVT U1610 ( .A1(n1102), .A2(n1468), .A3(n433), .A4(n1469), .A5(n1470), .A6(n24), .Y(n1566) );
  OA222X1_HVT U1611 ( .A1(n2200), .A2(n1447), .A3(n434), .A4(n1471), .A5(n924), 
        .A6(n1472), .Y(n1565) );
  MUX21X1_HVT U1612 ( .A1(n2191), .A2(keyout[124]), .S0(n1457), .Y(n3737) );
  NAND4X0_HVT U1613 ( .A1(n1569), .A2(n1570), .A3(n1571), .A4(n1572), .Y(n3736) );
  OA222X1_HVT U1614 ( .A1(n1103), .A2(n1462), .A3(n179), .A4(n1463), .A5(n692), 
        .A6(n1464), .Y(n1572) );
  OA222X1_HVT U1615 ( .A1(n1104), .A2(n1465), .A3(n180), .A4(n1466), .A5(n693), 
        .A6(n1467), .Y(n1571) );
  OA222X1_HVT U1616 ( .A1(n1105), .A2(n1468), .A3(n435), .A4(n1469), .A5(n1470), .A6(n25), .Y(n1570) );
  OA222X1_HVT U1617 ( .A1(n2198), .A2(n1447), .A3(n436), .A4(n1471), .A5(n925), 
        .A6(n1472), .Y(n1569) );
  MUX21X1_HVT U1618 ( .A1(n2189), .A2(keyout[125]), .S0(n1457), .Y(n3735) );
  NAND4X0_HVT U1619 ( .A1(n1573), .A2(n1574), .A3(n1575), .A4(n1576), .Y(n3734) );
  OA222X1_HVT U1620 ( .A1(n1106), .A2(n1462), .A3(n181), .A4(n1463), .A5(n694), 
        .A6(n1464), .Y(n1576) );
  OA222X1_HVT U1621 ( .A1(n1107), .A2(n1465), .A3(n182), .A4(n1466), .A5(n695), 
        .A6(n1467), .Y(n1575) );
  OA222X1_HVT U1622 ( .A1(n1108), .A2(n1468), .A3(n437), .A4(n1469), .A5(n1470), .A6(n26), .Y(n1574) );
  OA222X1_HVT U1623 ( .A1(n2196), .A2(n1447), .A3(n438), .A4(n1471), .A5(n926), 
        .A6(n1472), .Y(n1573) );
  MUX21X1_HVT U1624 ( .A1(n2187), .A2(keyout[126]), .S0(n1457), .Y(n3733) );
  NAND4X0_HVT U1625 ( .A1(n1577), .A2(n1578), .A3(n1579), .A4(n1580), .Y(n3732) );
  OA222X1_HVT U1626 ( .A1(n1109), .A2(n1462), .A3(n183), .A4(n1463), .A5(n696), 
        .A6(n1464), .Y(n1580) );
  OA222X1_HVT U1627 ( .A1(n1110), .A2(n1465), .A3(n184), .A4(n1466), .A5(n697), 
        .A6(n1467), .Y(n1579) );
  OA222X1_HVT U1628 ( .A1(n1111), .A2(n1468), .A3(n439), .A4(n1469), .A5(n1470), .A6(n27), .Y(n1578) );
  OA222X1_HVT U1629 ( .A1(n2194), .A2(n1447), .A3(n440), .A4(n1471), .A5(n927), 
        .A6(n1472), .Y(n1577) );
  MUX21X1_HVT U1630 ( .A1(n2185), .A2(keyout[127]), .S0(n1457), .Y(n3731) );
  NAND4X0_HVT U1631 ( .A1(n1581), .A2(n1582), .A3(n1583), .A4(n1584), .Y(n3730) );
  OA222X1_HVT U1632 ( .A1(n1112), .A2(n1462), .A3(n185), .A4(n1463), .A5(n698), 
        .A6(n1464), .Y(n1584) );
  OA222X1_HVT U1633 ( .A1(n1113), .A2(n1465), .A3(n186), .A4(n1466), .A5(n699), 
        .A6(n1467), .Y(n1583) );
  OA222X1_HVT U1634 ( .A1(n1114), .A2(n1468), .A3(n441), .A4(n1469), .A5(n1470), .A6(n28), .Y(n1582) );
  OA222X1_HVT U1635 ( .A1(n2192), .A2(n1447), .A3(n442), .A4(n1471), .A5(n928), 
        .A6(n1472), .Y(n1581) );
  MUX21X1_HVT U1636 ( .A1(n2183), .A2(keyout[82]), .S0(n1457), .Y(n3729) );
  NAND4X0_HVT U1637 ( .A1(n1585), .A2(n1586), .A3(n1587), .A4(n1588), .Y(n3728) );
  OA222X1_HVT U1638 ( .A1(n1115), .A2(n1462), .A3(n187), .A4(n1463), .A5(n700), 
        .A6(n1464), .Y(n1588) );
  OA222X1_HVT U1639 ( .A1(n1116), .A2(n1465), .A3(n188), .A4(n1466), .A5(n701), 
        .A6(n1467), .Y(n1587) );
  OA222X1_HVT U1640 ( .A1(n1117), .A2(n1468), .A3(n443), .A4(n1469), .A5(n1470), .A6(n29), .Y(n1586) );
  OA222X1_HVT U1641 ( .A1(n2190), .A2(n1447), .A3(n444), .A4(n1471), .A5(n929), 
        .A6(n1472), .Y(n1585) );
  MUX21X1_HVT U1642 ( .A1(n2181), .A2(keyout[83]), .S0(n1457), .Y(n3727) );
  NAND4X0_HVT U1643 ( .A1(n1589), .A2(n1590), .A3(n1591), .A4(n1592), .Y(n3726) );
  OA222X1_HVT U1644 ( .A1(n1118), .A2(n1462), .A3(n189), .A4(n1463), .A5(n702), 
        .A6(n1464), .Y(n1592) );
  OA222X1_HVT U1645 ( .A1(n1119), .A2(n1465), .A3(n190), .A4(n1466), .A5(n703), 
        .A6(n1467), .Y(n1591) );
  OA222X1_HVT U1646 ( .A1(n1120), .A2(n1468), .A3(n445), .A4(n1469), .A5(n1470), .A6(n30), .Y(n1590) );
  OA222X1_HVT U1647 ( .A1(n2188), .A2(n1447), .A3(n446), .A4(n1471), .A5(n930), 
        .A6(n1472), .Y(n1589) );
  MUX21X1_HVT U1648 ( .A1(n2179), .A2(keyout[84]), .S0(n1457), .Y(n3725) );
  NAND4X0_HVT U1649 ( .A1(n1593), .A2(n1594), .A3(n1595), .A4(n1596), .Y(n3724) );
  OA222X1_HVT U1650 ( .A1(n1121), .A2(n1462), .A3(n191), .A4(n1463), .A5(n704), 
        .A6(n1464), .Y(n1596) );
  OA222X1_HVT U1651 ( .A1(n1122), .A2(n1465), .A3(n192), .A4(n1466), .A5(n705), 
        .A6(n1467), .Y(n1595) );
  OA222X1_HVT U1652 ( .A1(n1123), .A2(n1468), .A3(n447), .A4(n1469), .A5(n1470), .A6(n31), .Y(n1594) );
  OA222X1_HVT U1653 ( .A1(n2186), .A2(n1447), .A3(n448), .A4(n1471), .A5(n931), 
        .A6(n1472), .Y(n1593) );
  MUX21X1_HVT U1654 ( .A1(n2177), .A2(keyout[85]), .S0(n1457), .Y(n3723) );
  NAND4X0_HVT U1655 ( .A1(n1597), .A2(n1598), .A3(n1599), .A4(n1600), .Y(n3722) );
  OA222X1_HVT U1656 ( .A1(n1124), .A2(n1462), .A3(n193), .A4(n1463), .A5(n706), 
        .A6(n1464), .Y(n1600) );
  OA222X1_HVT U1657 ( .A1(n1125), .A2(n1465), .A3(n194), .A4(n1466), .A5(n707), 
        .A6(n1467), .Y(n1599) );
  OA222X1_HVT U1658 ( .A1(n1126), .A2(n1468), .A3(n449), .A4(n1469), .A5(n1470), .A6(n32), .Y(n1598) );
  OA222X1_HVT U1659 ( .A1(n2184), .A2(n1447), .A3(n450), .A4(n1471), .A5(n932), 
        .A6(n1472), .Y(n1597) );
  MUX21X1_HVT U1660 ( .A1(n2175), .A2(keyout[86]), .S0(n1457), .Y(n3721) );
  NAND4X0_HVT U1661 ( .A1(n1601), .A2(n1602), .A3(n1603), .A4(n1604), .Y(n3720) );
  OA222X1_HVT U1662 ( .A1(n1127), .A2(n1462), .A3(n195), .A4(n1463), .A5(n708), 
        .A6(n1464), .Y(n1604) );
  OA222X1_HVT U1663 ( .A1(n1128), .A2(n1465), .A3(n196), .A4(n1466), .A5(n709), 
        .A6(n1467), .Y(n1603) );
  OA222X1_HVT U1664 ( .A1(n1129), .A2(n1468), .A3(n451), .A4(n1469), .A5(n1470), .A6(n33), .Y(n1602) );
  OA222X1_HVT U1665 ( .A1(n2182), .A2(n1447), .A3(n452), .A4(n1471), .A5(n933), 
        .A6(n1472), .Y(n1601) );
  MUX21X1_HVT U1666 ( .A1(n2173), .A2(keyout[87]), .S0(n1457), .Y(n3719) );
  NAND4X0_HVT U1667 ( .A1(n1605), .A2(n1606), .A3(n1607), .A4(n1608), .Y(n3718) );
  OA222X1_HVT U1668 ( .A1(n1130), .A2(n1462), .A3(n197), .A4(n1463), .A5(n710), 
        .A6(n1464), .Y(n1608) );
  OA222X1_HVT U1669 ( .A1(n1131), .A2(n1465), .A3(n198), .A4(n1466), .A5(n711), 
        .A6(n1467), .Y(n1607) );
  OA222X1_HVT U1670 ( .A1(n1132), .A2(n1468), .A3(n453), .A4(n1469), .A5(n1470), .A6(n34), .Y(n1606) );
  OA222X1_HVT U1671 ( .A1(n2180), .A2(n1447), .A3(n454), .A4(n1471), .A5(n934), 
        .A6(n1472), .Y(n1605) );
  MUX21X1_HVT U1672 ( .A1(n2171), .A2(keyout[88]), .S0(n1457), .Y(n3717) );
  NAND4X0_HVT U1673 ( .A1(n1609), .A2(n1610), .A3(n1611), .A4(n1612), .Y(n3716) );
  OA222X1_HVT U1674 ( .A1(n1133), .A2(n1462), .A3(n199), .A4(n1463), .A5(n712), 
        .A6(n1464), .Y(n1612) );
  OA222X1_HVT U1675 ( .A1(n1134), .A2(n1465), .A3(n200), .A4(n1466), .A5(n713), 
        .A6(n1467), .Y(n1611) );
  OA222X1_HVT U1676 ( .A1(n1135), .A2(n1468), .A3(n455), .A4(n1469), .A5(n1470), .A6(n35), .Y(n1610) );
  OA222X1_HVT U1677 ( .A1(n2178), .A2(n1447), .A3(n456), .A4(n1471), .A5(n935), 
        .A6(n1472), .Y(n1609) );
  MUX21X1_HVT U1678 ( .A1(n2169), .A2(keyout[89]), .S0(n1457), .Y(n3715) );
  NAND4X0_HVT U1679 ( .A1(n1613), .A2(n1614), .A3(n1615), .A4(n1616), .Y(n3714) );
  OA222X1_HVT U1680 ( .A1(n1136), .A2(n1462), .A3(n201), .A4(n1463), .A5(n714), 
        .A6(n1464), .Y(n1616) );
  OA222X1_HVT U1681 ( .A1(n1137), .A2(n1465), .A3(n202), .A4(n1466), .A5(n715), 
        .A6(n1467), .Y(n1615) );
  OA222X1_HVT U1682 ( .A1(n1138), .A2(n1468), .A3(n457), .A4(n1469), .A5(n1470), .A6(n36), .Y(n1614) );
  OA222X1_HVT U1683 ( .A1(n2176), .A2(n1447), .A3(n458), .A4(n1471), .A5(n936), 
        .A6(n1472), .Y(n1613) );
  MUX21X1_HVT U1684 ( .A1(n2167), .A2(keyout[90]), .S0(n1457), .Y(n3713) );
  NAND4X0_HVT U1685 ( .A1(n1617), .A2(n1618), .A3(n1619), .A4(n1620), .Y(n3712) );
  OA222X1_HVT U1686 ( .A1(n1139), .A2(n1462), .A3(n203), .A4(n1463), .A5(n716), 
        .A6(n1464), .Y(n1620) );
  OA222X1_HVT U1687 ( .A1(n1140), .A2(n1465), .A3(n204), .A4(n1466), .A5(n717), 
        .A6(n1467), .Y(n1619) );
  OA222X1_HVT U1688 ( .A1(n1141), .A2(n1468), .A3(n459), .A4(n1469), .A5(n1470), .A6(n37), .Y(n1618) );
  OA222X1_HVT U1689 ( .A1(n2174), .A2(n1447), .A3(n460), .A4(n1471), .A5(n937), 
        .A6(n1472), .Y(n1617) );
  MUX21X1_HVT U1690 ( .A1(n2165), .A2(keyout[91]), .S0(n1457), .Y(n3711) );
  NAND4X0_HVT U1691 ( .A1(n1621), .A2(n1622), .A3(n1623), .A4(n1624), .Y(n3710) );
  OA222X1_HVT U1692 ( .A1(n1142), .A2(n1462), .A3(n205), .A4(n1463), .A5(n718), 
        .A6(n1464), .Y(n1624) );
  OA222X1_HVT U1693 ( .A1(n1143), .A2(n1465), .A3(n206), .A4(n1466), .A5(n719), 
        .A6(n1467), .Y(n1623) );
  OA222X1_HVT U1694 ( .A1(n1144), .A2(n1468), .A3(n461), .A4(n1469), .A5(n1470), .A6(n38), .Y(n1622) );
  OA222X1_HVT U1695 ( .A1(n2172), .A2(n1447), .A3(n462), .A4(n1471), .A5(n938), 
        .A6(n1472), .Y(n1621) );
  MUX21X1_HVT U1696 ( .A1(n2163), .A2(keyout[92]), .S0(n1457), .Y(n3709) );
  NAND4X0_HVT U1697 ( .A1(n1625), .A2(n1626), .A3(n1627), .A4(n1628), .Y(n3708) );
  OA222X1_HVT U1698 ( .A1(n1145), .A2(n1462), .A3(n207), .A4(n1463), .A5(n720), 
        .A6(n1464), .Y(n1628) );
  OA222X1_HVT U1699 ( .A1(n1146), .A2(n1465), .A3(n208), .A4(n1466), .A5(n721), 
        .A6(n1467), .Y(n1627) );
  OA222X1_HVT U1700 ( .A1(n1147), .A2(n1468), .A3(n463), .A4(n1469), .A5(n1470), .A6(n39), .Y(n1626) );
  OA222X1_HVT U1701 ( .A1(n2170), .A2(n1447), .A3(n464), .A4(n1471), .A5(n939), 
        .A6(n1472), .Y(n1625) );
  MUX21X1_HVT U1702 ( .A1(n2161), .A2(keyout[93]), .S0(n1457), .Y(n3707) );
  NAND4X0_HVT U1703 ( .A1(n1629), .A2(n1630), .A3(n1631), .A4(n1632), .Y(n3706) );
  OA222X1_HVT U1704 ( .A1(n1148), .A2(n1462), .A3(n209), .A4(n1463), .A5(n722), 
        .A6(n1464), .Y(n1632) );
  OA222X1_HVT U1705 ( .A1(n1149), .A2(n1465), .A3(n210), .A4(n1466), .A5(n723), 
        .A6(n1467), .Y(n1631) );
  OA222X1_HVT U1706 ( .A1(n1150), .A2(n1468), .A3(n465), .A4(n1469), .A5(n1470), .A6(n40), .Y(n1630) );
  OA222X1_HVT U1707 ( .A1(n2168), .A2(n1447), .A3(n466), .A4(n1471), .A5(n940), 
        .A6(n1472), .Y(n1629) );
  MUX21X1_HVT U1708 ( .A1(n2159), .A2(keyout[94]), .S0(n1457), .Y(n3705) );
  NAND4X0_HVT U1709 ( .A1(n1633), .A2(n1634), .A3(n1635), .A4(n1636), .Y(n3704) );
  OA222X1_HVT U1710 ( .A1(n1151), .A2(n1462), .A3(n211), .A4(n1463), .A5(n724), 
        .A6(n1464), .Y(n1636) );
  OA222X1_HVT U1711 ( .A1(n1152), .A2(n1465), .A3(n212), .A4(n1466), .A5(n725), 
        .A6(n1467), .Y(n1635) );
  OA222X1_HVT U1712 ( .A1(n1153), .A2(n1468), .A3(n467), .A4(n1469), .A5(n1470), .A6(n41), .Y(n1634) );
  OA222X1_HVT U1713 ( .A1(n2166), .A2(n1447), .A3(n468), .A4(n1471), .A5(n941), 
        .A6(n1472), .Y(n1633) );
  MUX21X1_HVT U1714 ( .A1(n2157), .A2(keyout[95]), .S0(n1457), .Y(n3703) );
  NAND4X0_HVT U1715 ( .A1(n1637), .A2(n1638), .A3(n1639), .A4(n1640), .Y(n3702) );
  OA222X1_HVT U1716 ( .A1(n1154), .A2(n1462), .A3(n213), .A4(n1463), .A5(n726), 
        .A6(n1464), .Y(n1640) );
  OA222X1_HVT U1717 ( .A1(n1155), .A2(n1465), .A3(n214), .A4(n1466), .A5(n727), 
        .A6(n1467), .Y(n1639) );
  OA222X1_HVT U1718 ( .A1(n1156), .A2(n1468), .A3(n469), .A4(n1469), .A5(n1470), .A6(n42), .Y(n1638) );
  OA222X1_HVT U1719 ( .A1(n2164), .A2(n1447), .A3(n470), .A4(n1471), .A5(n942), 
        .A6(n1472), .Y(n1637) );
  MUX21X1_HVT U1720 ( .A1(n2155), .A2(keyout[96]), .S0(n1457), .Y(n3701) );
  NAND4X0_HVT U1721 ( .A1(n1641), .A2(n1642), .A3(n1643), .A4(n1644), .Y(n3700) );
  OA222X1_HVT U1722 ( .A1(n1157), .A2(n1462), .A3(n215), .A4(n1463), .A5(n728), 
        .A6(n1464), .Y(n1644) );
  OA222X1_HVT U1723 ( .A1(n1158), .A2(n1465), .A3(n216), .A4(n1466), .A5(n729), 
        .A6(n1467), .Y(n1643) );
  OA222X1_HVT U1724 ( .A1(n1159), .A2(n1468), .A3(n471), .A4(n1469), .A5(n1470), .A6(n43), .Y(n1642) );
  OA222X1_HVT U1725 ( .A1(n2162), .A2(n1447), .A3(n472), .A4(n1471), .A5(n943), 
        .A6(n1472), .Y(n1641) );
  MUX21X1_HVT U1726 ( .A1(n2153), .A2(keyout[97]), .S0(n1457), .Y(n3699) );
  NAND4X0_HVT U1727 ( .A1(n1645), .A2(n1646), .A3(n1647), .A4(n1648), .Y(n3698) );
  OA222X1_HVT U1728 ( .A1(n1160), .A2(n1462), .A3(n217), .A4(n1463), .A5(n730), 
        .A6(n1464), .Y(n1648) );
  OA222X1_HVT U1729 ( .A1(n1161), .A2(n1465), .A3(n218), .A4(n1466), .A5(n731), 
        .A6(n1467), .Y(n1647) );
  OA222X1_HVT U1730 ( .A1(n1162), .A2(n1468), .A3(n473), .A4(n1469), .A5(n1470), .A6(n44), .Y(n1646) );
  OA222X1_HVT U1731 ( .A1(n2160), .A2(n1447), .A3(n474), .A4(n1471), .A5(n944), 
        .A6(n1472), .Y(n1645) );
  MUX21X1_HVT U1732 ( .A1(n2151), .A2(keyout[0]), .S0(n1457), .Y(n3697) );
  NAND4X0_HVT U1733 ( .A1(n1649), .A2(n1650), .A3(n1651), .A4(n1652), .Y(n3696) );
  OA222X1_HVT U1734 ( .A1(n1163), .A2(n1462), .A3(n219), .A4(n1463), .A5(n732), 
        .A6(n1464), .Y(n1652) );
  OA222X1_HVT U1735 ( .A1(n1164), .A2(n1465), .A3(n220), .A4(n1466), .A5(n733), 
        .A6(n1467), .Y(n1651) );
  OA222X1_HVT U1736 ( .A1(n1165), .A2(n1468), .A3(n475), .A4(n1469), .A5(n1470), .A6(n45), .Y(n1650) );
  OA222X1_HVT U1737 ( .A1(n2158), .A2(n1447), .A3(n476), .A4(n1471), .A5(n945), 
        .A6(n1472), .Y(n1649) );
  MUX21X1_HVT U1738 ( .A1(n2149), .A2(keyout[1]), .S0(n1457), .Y(n3695) );
  NAND4X0_HVT U1739 ( .A1(n1653), .A2(n1654), .A3(n1655), .A4(n1656), .Y(n3694) );
  OA222X1_HVT U1740 ( .A1(n1166), .A2(n1462), .A3(n221), .A4(n1463), .A5(n734), 
        .A6(n1464), .Y(n1656) );
  OA222X1_HVT U1741 ( .A1(n1167), .A2(n1465), .A3(n222), .A4(n1466), .A5(n735), 
        .A6(n1467), .Y(n1655) );
  OA222X1_HVT U1742 ( .A1(n1168), .A2(n1468), .A3(n477), .A4(n1469), .A5(n1470), .A6(n46), .Y(n1654) );
  OA222X1_HVT U1743 ( .A1(n2156), .A2(n1447), .A3(n478), .A4(n1471), .A5(n946), 
        .A6(n1472), .Y(n1653) );
  MUX21X1_HVT U1744 ( .A1(n2147), .A2(keyout[2]), .S0(n1457), .Y(n3693) );
  NAND4X0_HVT U1745 ( .A1(n1657), .A2(n1658), .A3(n1659), .A4(n1660), .Y(n3692) );
  OA222X1_HVT U1746 ( .A1(n1169), .A2(n1462), .A3(n223), .A4(n1463), .A5(n736), 
        .A6(n1464), .Y(n1660) );
  OA222X1_HVT U1747 ( .A1(n1170), .A2(n1465), .A3(n224), .A4(n1466), .A5(n737), 
        .A6(n1467), .Y(n1659) );
  OA222X1_HVT U1748 ( .A1(n1171), .A2(n1468), .A3(n479), .A4(n1469), .A5(n1470), .A6(n47), .Y(n1658) );
  OA222X1_HVT U1749 ( .A1(n2154), .A2(n1447), .A3(n480), .A4(n1471), .A5(n947), 
        .A6(n1472), .Y(n1657) );
  MUX21X1_HVT U1750 ( .A1(n2145), .A2(keyout[3]), .S0(n1457), .Y(n3691) );
  NAND4X0_HVT U1751 ( .A1(n1661), .A2(n1662), .A3(n1663), .A4(n1664), .Y(n3690) );
  OA222X1_HVT U1752 ( .A1(n1172), .A2(n1462), .A3(n225), .A4(n1463), .A5(n738), 
        .A6(n1464), .Y(n1664) );
  OA222X1_HVT U1753 ( .A1(n1173), .A2(n1465), .A3(n226), .A4(n1466), .A5(n739), 
        .A6(n1467), .Y(n1663) );
  OA222X1_HVT U1754 ( .A1(n1174), .A2(n1468), .A3(n481), .A4(n1469), .A5(n1470), .A6(n48), .Y(n1662) );
  OA222X1_HVT U1755 ( .A1(n2152), .A2(n1447), .A3(n482), .A4(n1471), .A5(n948), 
        .A6(n1472), .Y(n1661) );
  MUX21X1_HVT U1756 ( .A1(n2143), .A2(keyout[4]), .S0(n1457), .Y(n3689) );
  NAND4X0_HVT U1757 ( .A1(n1665), .A2(n1666), .A3(n1667), .A4(n1668), .Y(n3688) );
  OA222X1_HVT U1758 ( .A1(n1175), .A2(n1462), .A3(n227), .A4(n1463), .A5(n740), 
        .A6(n1464), .Y(n1668) );
  OA222X1_HVT U1759 ( .A1(n1176), .A2(n1465), .A3(n228), .A4(n1466), .A5(n741), 
        .A6(n1467), .Y(n1667) );
  OA222X1_HVT U1760 ( .A1(n1177), .A2(n1468), .A3(n483), .A4(n1469), .A5(n1470), .A6(n49), .Y(n1666) );
  OA222X1_HVT U1761 ( .A1(n2150), .A2(n1447), .A3(n484), .A4(n1471), .A5(n949), 
        .A6(n1472), .Y(n1665) );
  MUX21X1_HVT U1762 ( .A1(n2141), .A2(keyout[5]), .S0(n1457), .Y(n3687) );
  NAND4X0_HVT U1763 ( .A1(n1669), .A2(n1670), .A3(n1671), .A4(n1672), .Y(n3686) );
  OA222X1_HVT U1764 ( .A1(n1178), .A2(n1462), .A3(n229), .A4(n1463), .A5(n742), 
        .A6(n1464), .Y(n1672) );
  OA222X1_HVT U1765 ( .A1(n1179), .A2(n1465), .A3(n230), .A4(n1466), .A5(n743), 
        .A6(n1467), .Y(n1671) );
  OA222X1_HVT U1766 ( .A1(n1180), .A2(n1468), .A3(n485), .A4(n1469), .A5(n1470), .A6(n50), .Y(n1670) );
  OA222X1_HVT U1767 ( .A1(n2148), .A2(n1447), .A3(n486), .A4(n1471), .A5(n950), 
        .A6(n1472), .Y(n1669) );
  MUX21X1_HVT U1768 ( .A1(n2139), .A2(keyout[6]), .S0(n1457), .Y(n3685) );
  NAND4X0_HVT U1769 ( .A1(n1673), .A2(n1674), .A3(n1675), .A4(n1676), .Y(n3684) );
  OA222X1_HVT U1770 ( .A1(n1181), .A2(n1462), .A3(n231), .A4(n1463), .A5(n744), 
        .A6(n1464), .Y(n1676) );
  OA222X1_HVT U1771 ( .A1(n1182), .A2(n1465), .A3(n232), .A4(n1466), .A5(n745), 
        .A6(n1467), .Y(n1675) );
  OA222X1_HVT U1772 ( .A1(n1183), .A2(n1468), .A3(n487), .A4(n1469), .A5(n1470), .A6(n51), .Y(n1674) );
  OA222X1_HVT U1773 ( .A1(n2146), .A2(n1447), .A3(n488), .A4(n1471), .A5(n951), 
        .A6(n1472), .Y(n1673) );
  MUX21X1_HVT U1774 ( .A1(n2137), .A2(keyout[7]), .S0(n1457), .Y(n3683) );
  NAND4X0_HVT U1775 ( .A1(n1677), .A2(n1678), .A3(n1679), .A4(n1680), .Y(n3682) );
  OA222X1_HVT U1776 ( .A1(n1184), .A2(n1462), .A3(n233), .A4(n1463), .A5(n746), 
        .A6(n1464), .Y(n1680) );
  OA222X1_HVT U1777 ( .A1(n1185), .A2(n1465), .A3(n234), .A4(n1466), .A5(n747), 
        .A6(n1467), .Y(n1679) );
  OA222X1_HVT U1778 ( .A1(n1186), .A2(n1468), .A3(n489), .A4(n1469), .A5(n1470), .A6(n52), .Y(n1678) );
  OA222X1_HVT U1779 ( .A1(n2144), .A2(n1447), .A3(n490), .A4(n1471), .A5(n952), 
        .A6(n1472), .Y(n1677) );
  MUX21X1_HVT U1780 ( .A1(n2135), .A2(keyout[8]), .S0(n1457), .Y(n3681) );
  NAND4X0_HVT U1781 ( .A1(n1681), .A2(n1682), .A3(n1683), .A4(n1684), .Y(n3680) );
  OA222X1_HVT U1782 ( .A1(n1187), .A2(n1462), .A3(n235), .A4(n1463), .A5(n748), 
        .A6(n1464), .Y(n1684) );
  OA222X1_HVT U1783 ( .A1(n1188), .A2(n1465), .A3(n236), .A4(n1466), .A5(n749), 
        .A6(n1467), .Y(n1683) );
  OA222X1_HVT U1784 ( .A1(n1189), .A2(n1468), .A3(n491), .A4(n1469), .A5(n1470), .A6(n53), .Y(n1682) );
  OA222X1_HVT U1785 ( .A1(n2142), .A2(n1447), .A3(n492), .A4(n1471), .A5(n953), 
        .A6(n1472), .Y(n1681) );
  MUX21X1_HVT U1786 ( .A1(n2133), .A2(keyout[9]), .S0(n1457), .Y(n3679) );
  NAND4X0_HVT U1787 ( .A1(n1685), .A2(n1686), .A3(n1687), .A4(n1688), .Y(n3678) );
  OA222X1_HVT U1788 ( .A1(n1190), .A2(n1462), .A3(n237), .A4(n1463), .A5(n750), 
        .A6(n1464), .Y(n1688) );
  OA222X1_HVT U1789 ( .A1(n1191), .A2(n1465), .A3(n238), .A4(n1466), .A5(n751), 
        .A6(n1467), .Y(n1687) );
  OA222X1_HVT U1790 ( .A1(n1192), .A2(n1468), .A3(n493), .A4(n1469), .A5(n1470), .A6(n54), .Y(n1686) );
  OA222X1_HVT U1791 ( .A1(n2140), .A2(n1447), .A3(n494), .A4(n1471), .A5(n954), 
        .A6(n1472), .Y(n1685) );
  MUX21X1_HVT U1792 ( .A1(n2131), .A2(keyout[10]), .S0(n1457), .Y(n3677) );
  NAND4X0_HVT U1793 ( .A1(n1689), .A2(n1690), .A3(n1691), .A4(n1692), .Y(n3676) );
  OA222X1_HVT U1794 ( .A1(n1193), .A2(n1462), .A3(n239), .A4(n1463), .A5(n752), 
        .A6(n1464), .Y(n1692) );
  OA222X1_HVT U1795 ( .A1(n1194), .A2(n1465), .A3(n240), .A4(n1466), .A5(n753), 
        .A6(n1467), .Y(n1691) );
  OA222X1_HVT U1796 ( .A1(n1195), .A2(n1468), .A3(n495), .A4(n1469), .A5(n1470), .A6(n55), .Y(n1690) );
  OA222X1_HVT U1797 ( .A1(n2138), .A2(n1447), .A3(n496), .A4(n1471), .A5(n955), 
        .A6(n1472), .Y(n1689) );
  MUX21X1_HVT U1798 ( .A1(n2129), .A2(keyout[11]), .S0(n1457), .Y(n3675) );
  NAND4X0_HVT U1799 ( .A1(n1693), .A2(n1694), .A3(n1695), .A4(n1696), .Y(n3674) );
  OA222X1_HVT U1800 ( .A1(n1196), .A2(n1462), .A3(n241), .A4(n1463), .A5(n754), 
        .A6(n1464), .Y(n1696) );
  OA222X1_HVT U1801 ( .A1(n1197), .A2(n1465), .A3(n242), .A4(n1466), .A5(n755), 
        .A6(n1467), .Y(n1695) );
  OA222X1_HVT U1802 ( .A1(n1198), .A2(n1468), .A3(n497), .A4(n1469), .A5(n1470), .A6(n56), .Y(n1694) );
  OA222X1_HVT U1803 ( .A1(n2136), .A2(n1447), .A3(n498), .A4(n1471), .A5(n956), 
        .A6(n1472), .Y(n1693) );
  MUX21X1_HVT U1804 ( .A1(n2127), .A2(keyout[12]), .S0(n1457), .Y(n3673) );
  NAND4X0_HVT U1805 ( .A1(n1697), .A2(n1698), .A3(n1699), .A4(n1700), .Y(n3672) );
  OA222X1_HVT U1806 ( .A1(n1199), .A2(n1462), .A3(n243), .A4(n1463), .A5(n756), 
        .A6(n1464), .Y(n1700) );
  OA222X1_HVT U1807 ( .A1(n1200), .A2(n1465), .A3(n244), .A4(n1466), .A5(n757), 
        .A6(n1467), .Y(n1699) );
  OA222X1_HVT U1808 ( .A1(n1201), .A2(n1468), .A3(n499), .A4(n1469), .A5(n1470), .A6(n57), .Y(n1698) );
  OA222X1_HVT U1809 ( .A1(n2134), .A2(n1447), .A3(n500), .A4(n1471), .A5(n957), 
        .A6(n1472), .Y(n1697) );
  MUX21X1_HVT U1810 ( .A1(n2125), .A2(keyout[13]), .S0(n1457), .Y(n3671) );
  NAND4X0_HVT U1811 ( .A1(n1701), .A2(n1702), .A3(n1703), .A4(n1704), .Y(n3670) );
  OA222X1_HVT U1812 ( .A1(n1202), .A2(n1462), .A3(n245), .A4(n1463), .A5(n758), 
        .A6(n1464), .Y(n1704) );
  OA222X1_HVT U1813 ( .A1(n1203), .A2(n1465), .A3(n246), .A4(n1466), .A5(n759), 
        .A6(n1467), .Y(n1703) );
  OA222X1_HVT U1814 ( .A1(n1204), .A2(n1468), .A3(n501), .A4(n1469), .A5(n1470), .A6(n58), .Y(n1702) );
  OA222X1_HVT U1815 ( .A1(n2132), .A2(n1447), .A3(n502), .A4(n1471), .A5(n958), 
        .A6(n1472), .Y(n1701) );
  MUX21X1_HVT U1816 ( .A1(n2123), .A2(keyout[14]), .S0(n1457), .Y(n3669) );
  NAND4X0_HVT U1817 ( .A1(n1705), .A2(n1706), .A3(n1707), .A4(n1708), .Y(n3668) );
  OA222X1_HVT U1818 ( .A1(n1205), .A2(n1462), .A3(n247), .A4(n1463), .A5(n760), 
        .A6(n1464), .Y(n1708) );
  OA222X1_HVT U1819 ( .A1(n1206), .A2(n1465), .A3(n248), .A4(n1466), .A5(n761), 
        .A6(n1467), .Y(n1707) );
  OA222X1_HVT U1820 ( .A1(n1207), .A2(n1468), .A3(n503), .A4(n1469), .A5(n1470), .A6(n59), .Y(n1706) );
  OA222X1_HVT U1821 ( .A1(n2130), .A2(n1447), .A3(n504), .A4(n1471), .A5(n959), 
        .A6(n1472), .Y(n1705) );
  MUX21X1_HVT U1822 ( .A1(n2121), .A2(keyout[15]), .S0(n1457), .Y(n3667) );
  NAND4X0_HVT U1823 ( .A1(n1709), .A2(n1710), .A3(n1711), .A4(n1712), .Y(n3666) );
  OA222X1_HVT U1824 ( .A1(n1208), .A2(n1462), .A3(n249), .A4(n1463), .A5(n762), 
        .A6(n1464), .Y(n1712) );
  OA222X1_HVT U1825 ( .A1(n1209), .A2(n1465), .A3(n250), .A4(n1466), .A5(n763), 
        .A6(n1467), .Y(n1711) );
  OA222X1_HVT U1826 ( .A1(n1210), .A2(n1468), .A3(n505), .A4(n1469), .A5(n1470), .A6(n60), .Y(n1710) );
  OA222X1_HVT U1827 ( .A1(n2128), .A2(n1447), .A3(n506), .A4(n1471), .A5(n960), 
        .A6(n1472), .Y(n1709) );
  MUX21X1_HVT U1828 ( .A1(n2119), .A2(keyout[16]), .S0(n1457), .Y(n3665) );
  NAND4X0_HVT U1829 ( .A1(n1713), .A2(n1714), .A3(n1715), .A4(n1716), .Y(n3664) );
  OA222X1_HVT U1830 ( .A1(n1211), .A2(n1462), .A3(n251), .A4(n1463), .A5(n764), 
        .A6(n1464), .Y(n1716) );
  OA222X1_HVT U1831 ( .A1(n1212), .A2(n1465), .A3(n252), .A4(n1466), .A5(n765), 
        .A6(n1467), .Y(n1715) );
  OA222X1_HVT U1832 ( .A1(n1213), .A2(n1468), .A3(n507), .A4(n1469), .A5(n1470), .A6(n61), .Y(n1714) );
  OA222X1_HVT U1833 ( .A1(n2126), .A2(n1447), .A3(n508), .A4(n1471), .A5(n961), 
        .A6(n1472), .Y(n1713) );
  MUX21X1_HVT U1834 ( .A1(n2117), .A2(keyout[17]), .S0(n1457), .Y(n3663) );
  NAND4X0_HVT U1835 ( .A1(n1717), .A2(n1718), .A3(n1719), .A4(n1720), .Y(n3662) );
  OA222X1_HVT U1836 ( .A1(n1214), .A2(n1462), .A3(n253), .A4(n1463), .A5(n766), 
        .A6(n1464), .Y(n1720) );
  OA222X1_HVT U1837 ( .A1(n1215), .A2(n1465), .A3(n254), .A4(n1466), .A5(n767), 
        .A6(n1467), .Y(n1719) );
  OA222X1_HVT U1838 ( .A1(n1216), .A2(n1468), .A3(n509), .A4(n1469), .A5(n1470), .A6(n62), .Y(n1718) );
  OA222X1_HVT U1839 ( .A1(n2124), .A2(n1447), .A3(n510), .A4(n1471), .A5(n962), 
        .A6(n1472), .Y(n1717) );
  MUX21X1_HVT U1840 ( .A1(n2115), .A2(keyout[18]), .S0(n1457), .Y(n3661) );
  NAND4X0_HVT U1841 ( .A1(n1721), .A2(n1722), .A3(n1723), .A4(n1724), .Y(n3660) );
  OA222X1_HVT U1842 ( .A1(n1217), .A2(n1462), .A3(n255), .A4(n1463), .A5(n768), 
        .A6(n1464), .Y(n1724) );
  OA222X1_HVT U1843 ( .A1(n1218), .A2(n1465), .A3(n256), .A4(n1466), .A5(n769), 
        .A6(n1467), .Y(n1723) );
  OA222X1_HVT U1844 ( .A1(n1219), .A2(n1468), .A3(n511), .A4(n1469), .A5(n1470), .A6(n63), .Y(n1722) );
  OA222X1_HVT U1845 ( .A1(n2122), .A2(n1447), .A3(n512), .A4(n1471), .A5(n963), 
        .A6(n1472), .Y(n1721) );
  MUX21X1_HVT U1846 ( .A1(n2113), .A2(keyout[19]), .S0(n1457), .Y(n3659) );
  NAND4X0_HVT U1847 ( .A1(n1725), .A2(n1726), .A3(n1727), .A4(n1728), .Y(n3658) );
  OA222X1_HVT U1848 ( .A1(n1220), .A2(n1462), .A3(n257), .A4(n1463), .A5(n770), 
        .A6(n1464), .Y(n1728) );
  OA222X1_HVT U1849 ( .A1(n1221), .A2(n1465), .A3(n258), .A4(n1466), .A5(n771), 
        .A6(n1467), .Y(n1727) );
  OA222X1_HVT U1850 ( .A1(n1222), .A2(n1468), .A3(n513), .A4(n1469), .A5(n1470), .A6(n64), .Y(n1726) );
  OA222X1_HVT U1851 ( .A1(n2120), .A2(n1447), .A3(n514), .A4(n1471), .A5(n964), 
        .A6(n1472), .Y(n1725) );
  MUX21X1_HVT U1852 ( .A1(n2111), .A2(keyout[20]), .S0(n1457), .Y(n3657) );
  NAND4X0_HVT U1853 ( .A1(n1729), .A2(n1730), .A3(n1731), .A4(n1732), .Y(n3656) );
  OA222X1_HVT U1854 ( .A1(n1223), .A2(n1462), .A3(n259), .A4(n1463), .A5(n772), 
        .A6(n1464), .Y(n1732) );
  OA222X1_HVT U1855 ( .A1(n1224), .A2(n1465), .A3(n260), .A4(n1466), .A5(n773), 
        .A6(n1467), .Y(n1731) );
  OA222X1_HVT U1856 ( .A1(n1225), .A2(n1468), .A3(n515), .A4(n1469), .A5(n1470), .A6(n65), .Y(n1730) );
  OA222X1_HVT U1857 ( .A1(n2118), .A2(n1447), .A3(n516), .A4(n1471), .A5(n965), 
        .A6(n1472), .Y(n1729) );
  MUX21X1_HVT U1858 ( .A1(n2109), .A2(keyout[21]), .S0(n1457), .Y(n3655) );
  NAND4X0_HVT U1859 ( .A1(n1733), .A2(n1734), .A3(n1735), .A4(n1736), .Y(n3654) );
  OA222X1_HVT U1860 ( .A1(n1226), .A2(n1462), .A3(n261), .A4(n1463), .A5(n774), 
        .A6(n1464), .Y(n1736) );
  OA222X1_HVT U1861 ( .A1(n1227), .A2(n1465), .A3(n262), .A4(n1466), .A5(n775), 
        .A6(n1467), .Y(n1735) );
  OA222X1_HVT U1862 ( .A1(n1228), .A2(n1468), .A3(n517), .A4(n1469), .A5(n1470), .A6(n66), .Y(n1734) );
  OA222X1_HVT U1863 ( .A1(n2116), .A2(n1447), .A3(n518), .A4(n1471), .A5(n966), 
        .A6(n1472), .Y(n1733) );
  MUX21X1_HVT U1864 ( .A1(n2107), .A2(keyout[22]), .S0(n1457), .Y(n3653) );
  NAND4X0_HVT U1865 ( .A1(n1737), .A2(n1738), .A3(n1739), .A4(n1740), .Y(n3652) );
  OA222X1_HVT U1866 ( .A1(n1229), .A2(n1462), .A3(n263), .A4(n1463), .A5(n776), 
        .A6(n1464), .Y(n1740) );
  OA222X1_HVT U1867 ( .A1(n1230), .A2(n1465), .A3(n264), .A4(n1466), .A5(n777), 
        .A6(n1467), .Y(n1739) );
  OA222X1_HVT U1868 ( .A1(n1231), .A2(n1468), .A3(n519), .A4(n1469), .A5(n1470), .A6(n67), .Y(n1738) );
  OA222X1_HVT U1869 ( .A1(n2114), .A2(n1447), .A3(n520), .A4(n1471), .A5(n967), 
        .A6(n1472), .Y(n1737) );
  MUX21X1_HVT U1870 ( .A1(n2105), .A2(keyout[23]), .S0(n1457), .Y(n3651) );
  NAND4X0_HVT U1871 ( .A1(n1741), .A2(n1742), .A3(n1743), .A4(n1744), .Y(n3650) );
  OA222X1_HVT U1872 ( .A1(n1232), .A2(n1462), .A3(n265), .A4(n1463), .A5(n778), 
        .A6(n1464), .Y(n1744) );
  OA222X1_HVT U1873 ( .A1(n1233), .A2(n1465), .A3(n266), .A4(n1466), .A5(n779), 
        .A6(n1467), .Y(n1743) );
  OA222X1_HVT U1874 ( .A1(n1234), .A2(n1468), .A3(n521), .A4(n1469), .A5(n1470), .A6(n68), .Y(n1742) );
  OA222X1_HVT U1875 ( .A1(n2112), .A2(n1447), .A3(n522), .A4(n1471), .A5(n968), 
        .A6(n1472), .Y(n1741) );
  MUX21X1_HVT U1876 ( .A1(n2103), .A2(keyout[24]), .S0(n1457), .Y(n3649) );
  NAND4X0_HVT U1877 ( .A1(n1745), .A2(n1746), .A3(n1747), .A4(n1748), .Y(n3648) );
  OA222X1_HVT U1878 ( .A1(n1235), .A2(n1462), .A3(n267), .A4(n1463), .A5(n780), 
        .A6(n1464), .Y(n1748) );
  OA222X1_HVT U1879 ( .A1(n1236), .A2(n1465), .A3(n268), .A4(n1466), .A5(n781), 
        .A6(n1467), .Y(n1747) );
  OA222X1_HVT U1880 ( .A1(n1237), .A2(n1468), .A3(n523), .A4(n1469), .A5(n1470), .A6(n69), .Y(n1746) );
  OA222X1_HVT U1881 ( .A1(n2110), .A2(n1447), .A3(n524), .A4(n1471), .A5(n969), 
        .A6(n1472), .Y(n1745) );
  MUX21X1_HVT U1882 ( .A1(n2101), .A2(keyout[25]), .S0(n1457), .Y(n3647) );
  NAND4X0_HVT U1883 ( .A1(n1749), .A2(n1750), .A3(n1751), .A4(n1752), .Y(n3646) );
  OA222X1_HVT U1884 ( .A1(n1238), .A2(n1462), .A3(n269), .A4(n1463), .A5(n782), 
        .A6(n1464), .Y(n1752) );
  OA222X1_HVT U1885 ( .A1(n1239), .A2(n1465), .A3(n270), .A4(n1466), .A5(n783), 
        .A6(n1467), .Y(n1751) );
  OA222X1_HVT U1886 ( .A1(n1240), .A2(n1468), .A3(n525), .A4(n1469), .A5(n1470), .A6(n70), .Y(n1750) );
  OA222X1_HVT U1887 ( .A1(n2108), .A2(n1447), .A3(n526), .A4(n1471), .A5(n970), 
        .A6(n1472), .Y(n1749) );
  MUX21X1_HVT U1888 ( .A1(n2099), .A2(keyout[26]), .S0(n1457), .Y(n3645) );
  NAND4X0_HVT U1889 ( .A1(n1753), .A2(n1754), .A3(n1755), .A4(n1756), .Y(n3644) );
  OA222X1_HVT U1890 ( .A1(n1241), .A2(n1462), .A3(n271), .A4(n1463), .A5(n784), 
        .A6(n1464), .Y(n1756) );
  OA222X1_HVT U1891 ( .A1(n1242), .A2(n1465), .A3(n272), .A4(n1466), .A5(n785), 
        .A6(n1467), .Y(n1755) );
  OA222X1_HVT U1892 ( .A1(n1243), .A2(n1468), .A3(n527), .A4(n1469), .A5(n1470), .A6(n71), .Y(n1754) );
  OA222X1_HVT U1893 ( .A1(n2106), .A2(n1447), .A3(n528), .A4(n1471), .A5(n971), 
        .A6(n1472), .Y(n1753) );
  MUX21X1_HVT U1894 ( .A1(n2097), .A2(keyout[27]), .S0(n1457), .Y(n3643) );
  NAND4X0_HVT U1895 ( .A1(n1757), .A2(n1758), .A3(n1759), .A4(n1760), .Y(n3642) );
  OA222X1_HVT U1896 ( .A1(n1244), .A2(n1462), .A3(n273), .A4(n1463), .A5(n786), 
        .A6(n1464), .Y(n1760) );
  OA222X1_HVT U1897 ( .A1(n1245), .A2(n1465), .A3(n274), .A4(n1466), .A5(n787), 
        .A6(n1467), .Y(n1759) );
  OA222X1_HVT U1898 ( .A1(n1246), .A2(n1468), .A3(n529), .A4(n1469), .A5(n1470), .A6(n72), .Y(n1758) );
  OA222X1_HVT U1899 ( .A1(n2104), .A2(n1447), .A3(n530), .A4(n1471), .A5(n972), 
        .A6(n1472), .Y(n1757) );
  MUX21X1_HVT U1900 ( .A1(n2095), .A2(keyout[28]), .S0(n1457), .Y(n3641) );
  NAND4X0_HVT U1901 ( .A1(n1761), .A2(n1762), .A3(n1763), .A4(n1764), .Y(n3640) );
  OA222X1_HVT U1902 ( .A1(n1247), .A2(n1462), .A3(n275), .A4(n1463), .A5(n788), 
        .A6(n1464), .Y(n1764) );
  OA222X1_HVT U1903 ( .A1(n1248), .A2(n1465), .A3(n276), .A4(n1466), .A5(n789), 
        .A6(n1467), .Y(n1763) );
  OA222X1_HVT U1904 ( .A1(n1249), .A2(n1468), .A3(n531), .A4(n1469), .A5(n1470), .A6(n73), .Y(n1762) );
  OA222X1_HVT U1905 ( .A1(n2102), .A2(n1447), .A3(n532), .A4(n1471), .A5(n973), 
        .A6(n1472), .Y(n1761) );
  MUX21X1_HVT U1906 ( .A1(n2093), .A2(keyout[29]), .S0(n1457), .Y(n3639) );
  NAND4X0_HVT U1907 ( .A1(n1765), .A2(n1766), .A3(n1767), .A4(n1768), .Y(n3638) );
  OA222X1_HVT U1908 ( .A1(n1250), .A2(n1462), .A3(n277), .A4(n1463), .A5(n790), 
        .A6(n1464), .Y(n1768) );
  OA222X1_HVT U1909 ( .A1(n1251), .A2(n1465), .A3(n278), .A4(n1466), .A5(n791), 
        .A6(n1467), .Y(n1767) );
  OA222X1_HVT U1910 ( .A1(n1252), .A2(n1468), .A3(n533), .A4(n1469), .A5(n1470), .A6(n74), .Y(n1766) );
  OA222X1_HVT U1911 ( .A1(n2100), .A2(n1447), .A3(n534), .A4(n1471), .A5(n974), 
        .A6(n1472), .Y(n1765) );
  MUX21X1_HVT U1912 ( .A1(n2091), .A2(keyout[30]), .S0(n1457), .Y(n3637) );
  NAND4X0_HVT U1913 ( .A1(n1769), .A2(n1770), .A3(n1771), .A4(n1772), .Y(n3636) );
  OA222X1_HVT U1914 ( .A1(n1253), .A2(n1462), .A3(n279), .A4(n1463), .A5(n792), 
        .A6(n1464), .Y(n1772) );
  OA222X1_HVT U1915 ( .A1(n1254), .A2(n1465), .A3(n280), .A4(n1466), .A5(n793), 
        .A6(n1467), .Y(n1771) );
  OA222X1_HVT U1916 ( .A1(n1255), .A2(n1468), .A3(n535), .A4(n1469), .A5(n1470), .A6(n75), .Y(n1770) );
  OA222X1_HVT U1917 ( .A1(n2098), .A2(n1447), .A3(n536), .A4(n1471), .A5(n975), 
        .A6(n1472), .Y(n1769) );
  MUX21X1_HVT U1918 ( .A1(n2089), .A2(keyout[31]), .S0(n1457), .Y(n3635) );
  NAND4X0_HVT U1919 ( .A1(n1773), .A2(n1774), .A3(n1775), .A4(n1776), .Y(n3634) );
  OA222X1_HVT U1920 ( .A1(n1256), .A2(n1462), .A3(n281), .A4(n1463), .A5(n794), 
        .A6(n1464), .Y(n1776) );
  OA222X1_HVT U1921 ( .A1(n1257), .A2(n1465), .A3(n282), .A4(n1466), .A5(n795), 
        .A6(n1467), .Y(n1775) );
  OA222X1_HVT U1922 ( .A1(n1258), .A2(n1468), .A3(n537), .A4(n1469), .A5(n1470), .A6(n76), .Y(n1774) );
  OA222X1_HVT U1923 ( .A1(n2096), .A2(n1447), .A3(n538), .A4(n1471), .A5(n976), 
        .A6(n1472), .Y(n1773) );
  MUX21X1_HVT U1924 ( .A1(n2087), .A2(keyout[32]), .S0(n1457), .Y(n3633) );
  NAND4X0_HVT U1925 ( .A1(n1777), .A2(n1778), .A3(n1779), .A4(n1780), .Y(n3632) );
  OA222X1_HVT U1926 ( .A1(n1259), .A2(n1462), .A3(n283), .A4(n1463), .A5(n796), 
        .A6(n1464), .Y(n1780) );
  OA222X1_HVT U1927 ( .A1(n1260), .A2(n1465), .A3(n284), .A4(n1466), .A5(n797), 
        .A6(n1467), .Y(n1779) );
  OA222X1_HVT U1928 ( .A1(n1261), .A2(n1468), .A3(n539), .A4(n1469), .A5(n1470), .A6(n77), .Y(n1778) );
  OA222X1_HVT U1929 ( .A1(n2094), .A2(n1447), .A3(n540), .A4(n1471), .A5(n977), 
        .A6(n1472), .Y(n1777) );
  MUX21X1_HVT U1930 ( .A1(n2085), .A2(keyout[33]), .S0(n1457), .Y(n3631) );
  NAND4X0_HVT U1931 ( .A1(n1781), .A2(n1782), .A3(n1783), .A4(n1784), .Y(n3630) );
  OA222X1_HVT U1932 ( .A1(n1262), .A2(n1462), .A3(n285), .A4(n1463), .A5(n798), 
        .A6(n1464), .Y(n1784) );
  OA222X1_HVT U1933 ( .A1(n1263), .A2(n1465), .A3(n286), .A4(n1466), .A5(n799), 
        .A6(n1467), .Y(n1783) );
  OA222X1_HVT U1934 ( .A1(n1264), .A2(n1468), .A3(n541), .A4(n1469), .A5(n1470), .A6(n78), .Y(n1782) );
  OA222X1_HVT U1935 ( .A1(n2092), .A2(n1447), .A3(n542), .A4(n1471), .A5(n978), 
        .A6(n1472), .Y(n1781) );
  MUX21X1_HVT U1936 ( .A1(n2083), .A2(keyout[34]), .S0(n1457), .Y(n3629) );
  NAND4X0_HVT U1937 ( .A1(n1785), .A2(n1786), .A3(n1787), .A4(n1788), .Y(n3628) );
  OA222X1_HVT U1938 ( .A1(n1265), .A2(n1462), .A3(n287), .A4(n1463), .A5(n800), 
        .A6(n1464), .Y(n1788) );
  OA222X1_HVT U1939 ( .A1(n1266), .A2(n1465), .A3(n288), .A4(n1466), .A5(n801), 
        .A6(n1467), .Y(n1787) );
  OA222X1_HVT U1940 ( .A1(n1267), .A2(n1468), .A3(n543), .A4(n1469), .A5(n1470), .A6(n79), .Y(n1786) );
  OA222X1_HVT U1941 ( .A1(n2090), .A2(n1447), .A3(n544), .A4(n1471), .A5(n979), 
        .A6(n1472), .Y(n1785) );
  MUX21X1_HVT U1942 ( .A1(n2081), .A2(keyout[35]), .S0(n1457), .Y(n3627) );
  NAND4X0_HVT U1943 ( .A1(n1789), .A2(n1790), .A3(n1791), .A4(n1792), .Y(n3626) );
  OA222X1_HVT U1944 ( .A1(n1268), .A2(n1462), .A3(n289), .A4(n1463), .A5(n802), 
        .A6(n1464), .Y(n1792) );
  OA222X1_HVT U1945 ( .A1(n1269), .A2(n1465), .A3(n290), .A4(n1466), .A5(n803), 
        .A6(n1467), .Y(n1791) );
  OA222X1_HVT U1946 ( .A1(n1270), .A2(n1468), .A3(n545), .A4(n1469), .A5(n1470), .A6(n80), .Y(n1790) );
  OA222X1_HVT U1947 ( .A1(n2088), .A2(n1447), .A3(n546), .A4(n1471), .A5(n980), 
        .A6(n1472), .Y(n1789) );
  MUX21X1_HVT U1948 ( .A1(n2079), .A2(keyout[36]), .S0(n1457), .Y(n3625) );
  NAND4X0_HVT U1949 ( .A1(n1793), .A2(n1794), .A3(n1795), .A4(n1796), .Y(n3624) );
  OA222X1_HVT U1950 ( .A1(n1271), .A2(n1462), .A3(n291), .A4(n1463), .A5(n804), 
        .A6(n1464), .Y(n1796) );
  OA222X1_HVT U1951 ( .A1(n1272), .A2(n1465), .A3(n292), .A4(n1466), .A5(n805), 
        .A6(n1467), .Y(n1795) );
  OA222X1_HVT U1952 ( .A1(n1273), .A2(n1468), .A3(n547), .A4(n1469), .A5(n1470), .A6(n81), .Y(n1794) );
  OA222X1_HVT U1953 ( .A1(n2086), .A2(n1447), .A3(n548), .A4(n1471), .A5(n981), 
        .A6(n1472), .Y(n1793) );
  MUX21X1_HVT U1954 ( .A1(n2077), .A2(keyout[37]), .S0(n1457), .Y(n3623) );
  NAND4X0_HVT U1955 ( .A1(n1797), .A2(n1798), .A3(n1799), .A4(n1800), .Y(n3622) );
  OA222X1_HVT U1956 ( .A1(n1274), .A2(n1462), .A3(n293), .A4(n1463), .A5(n806), 
        .A6(n1464), .Y(n1800) );
  OA222X1_HVT U1957 ( .A1(n1275), .A2(n1465), .A3(n294), .A4(n1466), .A5(n807), 
        .A6(n1467), .Y(n1799) );
  OA222X1_HVT U1958 ( .A1(n1276), .A2(n1468), .A3(n549), .A4(n1469), .A5(n1470), .A6(n82), .Y(n1798) );
  OA222X1_HVT U1959 ( .A1(n2084), .A2(n1447), .A3(n550), .A4(n1471), .A5(n982), 
        .A6(n1472), .Y(n1797) );
  MUX21X1_HVT U1960 ( .A1(n2075), .A2(keyout[38]), .S0(n1457), .Y(n3621) );
  NAND4X0_HVT U1961 ( .A1(n1801), .A2(n1802), .A3(n1803), .A4(n1804), .Y(n3620) );
  OA222X1_HVT U1962 ( .A1(n1277), .A2(n1462), .A3(n295), .A4(n1463), .A5(n808), 
        .A6(n1464), .Y(n1804) );
  OA222X1_HVT U1963 ( .A1(n1278), .A2(n1465), .A3(n296), .A4(n1466), .A5(n809), 
        .A6(n1467), .Y(n1803) );
  OA222X1_HVT U1964 ( .A1(n1279), .A2(n1468), .A3(n551), .A4(n1469), .A5(n1470), .A6(n83), .Y(n1802) );
  OA222X1_HVT U1965 ( .A1(n2082), .A2(n1447), .A3(n552), .A4(n1471), .A5(n983), 
        .A6(n1472), .Y(n1801) );
  MUX21X1_HVT U1966 ( .A1(n2073), .A2(keyout[39]), .S0(n1457), .Y(n3619) );
  NAND4X0_HVT U1967 ( .A1(n1805), .A2(n1806), .A3(n1807), .A4(n1808), .Y(n3618) );
  OA222X1_HVT U1968 ( .A1(n1280), .A2(n1462), .A3(n297), .A4(n1463), .A5(n810), 
        .A6(n1464), .Y(n1808) );
  OA222X1_HVT U1969 ( .A1(n1281), .A2(n1465), .A3(n298), .A4(n1466), .A5(n811), 
        .A6(n1467), .Y(n1807) );
  OA222X1_HVT U1970 ( .A1(n1282), .A2(n1468), .A3(n553), .A4(n1469), .A5(n1470), .A6(n84), .Y(n1806) );
  OA222X1_HVT U1971 ( .A1(n2080), .A2(n1447), .A3(n554), .A4(n1471), .A5(n984), 
        .A6(n1472), .Y(n1805) );
  MUX21X1_HVT U1972 ( .A1(n2071), .A2(keyout[40]), .S0(n1457), .Y(n3617) );
  NAND4X0_HVT U1973 ( .A1(n1809), .A2(n1810), .A3(n1811), .A4(n1812), .Y(n3616) );
  OA222X1_HVT U1974 ( .A1(n1283), .A2(n1462), .A3(n299), .A4(n1463), .A5(n812), 
        .A6(n1464), .Y(n1812) );
  OA222X1_HVT U1975 ( .A1(n1284), .A2(n1465), .A3(n300), .A4(n1466), .A5(n813), 
        .A6(n1467), .Y(n1811) );
  OA222X1_HVT U1976 ( .A1(n1285), .A2(n1468), .A3(n555), .A4(n1469), .A5(n1470), .A6(n85), .Y(n1810) );
  OA222X1_HVT U1977 ( .A1(n2078), .A2(n1447), .A3(n556), .A4(n1471), .A5(n985), 
        .A6(n1472), .Y(n1809) );
  MUX21X1_HVT U1978 ( .A1(n2069), .A2(keyout[41]), .S0(n1457), .Y(n3615) );
  NAND4X0_HVT U1979 ( .A1(n1813), .A2(n1814), .A3(n1815), .A4(n1816), .Y(n3614) );
  OA222X1_HVT U1980 ( .A1(n1286), .A2(n1462), .A3(n301), .A4(n1463), .A5(n814), 
        .A6(n1464), .Y(n1816) );
  OA222X1_HVT U1981 ( .A1(n1287), .A2(n1465), .A3(n302), .A4(n1466), .A5(n815), 
        .A6(n1467), .Y(n1815) );
  OA222X1_HVT U1982 ( .A1(n1288), .A2(n1468), .A3(n557), .A4(n1469), .A5(n1470), .A6(n86), .Y(n1814) );
  OA222X1_HVT U1983 ( .A1(n2076), .A2(n1447), .A3(n558), .A4(n1471), .A5(n986), 
        .A6(n1472), .Y(n1813) );
  MUX21X1_HVT U1984 ( .A1(n2067), .A2(keyout[42]), .S0(n1457), .Y(n3613) );
  NAND4X0_HVT U1985 ( .A1(n1817), .A2(n1818), .A3(n1819), .A4(n1820), .Y(n3612) );
  OA222X1_HVT U1986 ( .A1(n1289), .A2(n1462), .A3(n303), .A4(n1463), .A5(n816), 
        .A6(n1464), .Y(n1820) );
  OA222X1_HVT U1987 ( .A1(n1290), .A2(n1465), .A3(n304), .A4(n1466), .A5(n817), 
        .A6(n1467), .Y(n1819) );
  OA222X1_HVT U1988 ( .A1(n1291), .A2(n1468), .A3(n559), .A4(n1469), .A5(n1470), .A6(n87), .Y(n1818) );
  OA222X1_HVT U1989 ( .A1(n2074), .A2(n1447), .A3(n560), .A4(n1471), .A5(n987), 
        .A6(n1472), .Y(n1817) );
  MUX21X1_HVT U1990 ( .A1(n2065), .A2(keyout[43]), .S0(n1457), .Y(n3611) );
  NAND4X0_HVT U1991 ( .A1(n1821), .A2(n1822), .A3(n1823), .A4(n1824), .Y(n3610) );
  OA222X1_HVT U1992 ( .A1(n1292), .A2(n1462), .A3(n305), .A4(n1463), .A5(n818), 
        .A6(n1464), .Y(n1824) );
  OA222X1_HVT U1993 ( .A1(n1293), .A2(n1465), .A3(n306), .A4(n1466), .A5(n819), 
        .A6(n1467), .Y(n1823) );
  OA222X1_HVT U1994 ( .A1(n1294), .A2(n1468), .A3(n561), .A4(n1469), .A5(n1470), .A6(n88), .Y(n1822) );
  OA222X1_HVT U1995 ( .A1(n2072), .A2(n1447), .A3(n562), .A4(n1471), .A5(n988), 
        .A6(n1472), .Y(n1821) );
  MUX21X1_HVT U1996 ( .A1(n2063), .A2(keyout[44]), .S0(n1457), .Y(n3609) );
  NAND4X0_HVT U1997 ( .A1(n1825), .A2(n1826), .A3(n1827), .A4(n1828), .Y(n3608) );
  OA222X1_HVT U1998 ( .A1(n1295), .A2(n1462), .A3(n307), .A4(n1463), .A5(n820), 
        .A6(n1464), .Y(n1828) );
  OA222X1_HVT U1999 ( .A1(n1296), .A2(n1465), .A3(n308), .A4(n1466), .A5(n821), 
        .A6(n1467), .Y(n1827) );
  OA222X1_HVT U2000 ( .A1(n1297), .A2(n1468), .A3(n563), .A4(n1469), .A5(n1470), .A6(n89), .Y(n1826) );
  OA222X1_HVT U2001 ( .A1(n2070), .A2(n1447), .A3(n564), .A4(n1471), .A5(n989), 
        .A6(n1472), .Y(n1825) );
  MUX21X1_HVT U2002 ( .A1(n2061), .A2(keyout[45]), .S0(n1457), .Y(n3607) );
  NAND4X0_HVT U2003 ( .A1(n1829), .A2(n1830), .A3(n1831), .A4(n1832), .Y(n3606) );
  OA222X1_HVT U2004 ( .A1(n1298), .A2(n1462), .A3(n309), .A4(n1463), .A5(n822), 
        .A6(n1464), .Y(n1832) );
  OA222X1_HVT U2005 ( .A1(n1299), .A2(n1465), .A3(n310), .A4(n1466), .A5(n823), 
        .A6(n1467), .Y(n1831) );
  OA222X1_HVT U2006 ( .A1(n1300), .A2(n1468), .A3(n565), .A4(n1469), .A5(n1470), .A6(n90), .Y(n1830) );
  OA222X1_HVT U2007 ( .A1(n2068), .A2(n1447), .A3(n566), .A4(n1471), .A5(n990), 
        .A6(n1472), .Y(n1829) );
  MUX21X1_HVT U2008 ( .A1(n2059), .A2(keyout[46]), .S0(n1457), .Y(n3605) );
  NAND4X0_HVT U2009 ( .A1(n1833), .A2(n1834), .A3(n1835), .A4(n1836), .Y(n3604) );
  OA222X1_HVT U2010 ( .A1(n1301), .A2(n1462), .A3(n311), .A4(n1463), .A5(n824), 
        .A6(n1464), .Y(n1836) );
  OA222X1_HVT U2011 ( .A1(n1302), .A2(n1465), .A3(n312), .A4(n1466), .A5(n825), 
        .A6(n1467), .Y(n1835) );
  OA222X1_HVT U2012 ( .A1(n1303), .A2(n1468), .A3(n567), .A4(n1469), .A5(n1470), .A6(n91), .Y(n1834) );
  OA222X1_HVT U2013 ( .A1(n2066), .A2(n1447), .A3(n568), .A4(n1471), .A5(n991), 
        .A6(n1472), .Y(n1833) );
  MUX21X1_HVT U2014 ( .A1(n2057), .A2(keyout[47]), .S0(n1457), .Y(n3603) );
  NAND4X0_HVT U2015 ( .A1(n1837), .A2(n1838), .A3(n1839), .A4(n1840), .Y(n3602) );
  OA222X1_HVT U2016 ( .A1(n1304), .A2(n1462), .A3(n313), .A4(n1463), .A5(n826), 
        .A6(n1464), .Y(n1840) );
  OA222X1_HVT U2017 ( .A1(n1305), .A2(n1465), .A3(n314), .A4(n1466), .A5(n827), 
        .A6(n1467), .Y(n1839) );
  OA222X1_HVT U2018 ( .A1(n1306), .A2(n1468), .A3(n569), .A4(n1469), .A5(n1470), .A6(n92), .Y(n1838) );
  OA222X1_HVT U2019 ( .A1(n2064), .A2(n1447), .A3(n570), .A4(n1471), .A5(n992), 
        .A6(n1472), .Y(n1837) );
  MUX21X1_HVT U2020 ( .A1(n2055), .A2(keyout[48]), .S0(n1457), .Y(n3601) );
  NAND4X0_HVT U2021 ( .A1(n1841), .A2(n1842), .A3(n1843), .A4(n1844), .Y(n3600) );
  OA222X1_HVT U2022 ( .A1(n1307), .A2(n1462), .A3(n315), .A4(n1463), .A5(n828), 
        .A6(n1464), .Y(n1844) );
  OA222X1_HVT U2023 ( .A1(n1308), .A2(n1465), .A3(n316), .A4(n1466), .A5(n829), 
        .A6(n1467), .Y(n1843) );
  OA222X1_HVT U2024 ( .A1(n1309), .A2(n1468), .A3(n571), .A4(n1469), .A5(n1470), .A6(n93), .Y(n1842) );
  OA222X1_HVT U2025 ( .A1(n2062), .A2(n1447), .A3(n572), .A4(n1471), .A5(n993), 
        .A6(n1472), .Y(n1841) );
  MUX21X1_HVT U2026 ( .A1(n2053), .A2(keyout[81]), .S0(n1457), .Y(n3599) );
  NAND4X0_HVT U2027 ( .A1(n1845), .A2(n1846), .A3(n1847), .A4(n1848), .Y(n3598) );
  OA222X1_HVT U2028 ( .A1(n1310), .A2(n1462), .A3(n317), .A4(n1463), .A5(n830), 
        .A6(n1464), .Y(n1848) );
  OA222X1_HVT U2029 ( .A1(n1311), .A2(n1465), .A3(n318), .A4(n1466), .A5(n831), 
        .A6(n1467), .Y(n1847) );
  OA222X1_HVT U2030 ( .A1(n1312), .A2(n1468), .A3(n573), .A4(n1469), .A5(n1470), .A6(n94), .Y(n1846) );
  OA222X1_HVT U2031 ( .A1(n2060), .A2(n1447), .A3(n574), .A4(n1471), .A5(n994), 
        .A6(n1472), .Y(n1845) );
  MUX21X1_HVT U2032 ( .A1(n2051), .A2(keyout[80]), .S0(n1457), .Y(n3597) );
  NAND4X0_HVT U2033 ( .A1(n1849), .A2(n1850), .A3(n1851), .A4(n1852), .Y(n3596) );
  OA222X1_HVT U2034 ( .A1(n1313), .A2(n1462), .A3(n319), .A4(n1463), .A5(n832), 
        .A6(n1464), .Y(n1852) );
  OA222X1_HVT U2035 ( .A1(n1314), .A2(n1465), .A3(n320), .A4(n1466), .A5(n833), 
        .A6(n1467), .Y(n1851) );
  OA222X1_HVT U2036 ( .A1(n1315), .A2(n1468), .A3(n575), .A4(n1469), .A5(n1470), .A6(n95), .Y(n1850) );
  OA222X1_HVT U2037 ( .A1(n2058), .A2(n1447), .A3(n576), .A4(n1471), .A5(n995), 
        .A6(n1472), .Y(n1849) );
  MUX21X1_HVT U2038 ( .A1(n2049), .A2(keyout[79]), .S0(n1457), .Y(n3595) );
  NAND4X0_HVT U2039 ( .A1(n1853), .A2(n1854), .A3(n1855), .A4(n1856), .Y(n3594) );
  OA222X1_HVT U2040 ( .A1(n1316), .A2(n1462), .A3(n321), .A4(n1463), .A5(n834), 
        .A6(n1464), .Y(n1856) );
  OA222X1_HVT U2041 ( .A1(n1317), .A2(n1465), .A3(n322), .A4(n1466), .A5(n835), 
        .A6(n1467), .Y(n1855) );
  OA222X1_HVT U2042 ( .A1(n1318), .A2(n1468), .A3(n577), .A4(n1469), .A5(n1470), .A6(n96), .Y(n1854) );
  OA222X1_HVT U2043 ( .A1(n2056), .A2(n1447), .A3(n578), .A4(n1471), .A5(n996), 
        .A6(n1472), .Y(n1853) );
  MUX21X1_HVT U2044 ( .A1(n2047), .A2(keyout[78]), .S0(n1457), .Y(n3593) );
  NAND4X0_HVT U2045 ( .A1(n1857), .A2(n1858), .A3(n1859), .A4(n1860), .Y(n3592) );
  OA222X1_HVT U2046 ( .A1(n1319), .A2(n1462), .A3(n323), .A4(n1463), .A5(n836), 
        .A6(n1464), .Y(n1860) );
  OA222X1_HVT U2047 ( .A1(n1320), .A2(n1465), .A3(n324), .A4(n1466), .A5(n837), 
        .A6(n1467), .Y(n1859) );
  OA222X1_HVT U2048 ( .A1(n1321), .A2(n1468), .A3(n579), .A4(n1469), .A5(n1470), .A6(n97), .Y(n1858) );
  OA222X1_HVT U2049 ( .A1(n2054), .A2(n1447), .A3(n580), .A4(n1471), .A5(n997), 
        .A6(n1472), .Y(n1857) );
  MUX21X1_HVT U2050 ( .A1(n2045), .A2(keyout[77]), .S0(n1457), .Y(n3591) );
  NAND4X0_HVT U2051 ( .A1(n1861), .A2(n1862), .A3(n1863), .A4(n1864), .Y(n3590) );
  OA222X1_HVT U2052 ( .A1(n1322), .A2(n1462), .A3(n325), .A4(n1463), .A5(n838), 
        .A6(n1464), .Y(n1864) );
  OA222X1_HVT U2053 ( .A1(n1323), .A2(n1465), .A3(n326), .A4(n1466), .A5(n839), 
        .A6(n1467), .Y(n1863) );
  OA222X1_HVT U2054 ( .A1(n1324), .A2(n1468), .A3(n581), .A4(n1469), .A5(n1470), .A6(n98), .Y(n1862) );
  OA222X1_HVT U2055 ( .A1(n2052), .A2(n1447), .A3(n582), .A4(n1471), .A5(n998), 
        .A6(n1472), .Y(n1861) );
  MUX21X1_HVT U2056 ( .A1(n2043), .A2(keyout[76]), .S0(n1457), .Y(n3589) );
  NAND4X0_HVT U2057 ( .A1(n1865), .A2(n1866), .A3(n1867), .A4(n1868), .Y(n3588) );
  OA222X1_HVT U2058 ( .A1(n1325), .A2(n1462), .A3(n327), .A4(n1463), .A5(n840), 
        .A6(n1464), .Y(n1868) );
  OA222X1_HVT U2059 ( .A1(n1326), .A2(n1465), .A3(n328), .A4(n1466), .A5(n841), 
        .A6(n1467), .Y(n1867) );
  OA222X1_HVT U2060 ( .A1(n1327), .A2(n1468), .A3(n583), .A4(n1469), .A5(n1470), .A6(n99), .Y(n1866) );
  OA222X1_HVT U2061 ( .A1(n2050), .A2(n1447), .A3(n584), .A4(n1471), .A5(n999), 
        .A6(n1472), .Y(n1865) );
  MUX21X1_HVT U2062 ( .A1(n2041), .A2(keyout[75]), .S0(n1457), .Y(n3587) );
  NAND4X0_HVT U2063 ( .A1(n1869), .A2(n1870), .A3(n1871), .A4(n1872), .Y(n3586) );
  OA222X1_HVT U2064 ( .A1(n1328), .A2(n1462), .A3(n329), .A4(n1463), .A5(n842), 
        .A6(n1464), .Y(n1872) );
  OA222X1_HVT U2065 ( .A1(n1329), .A2(n1465), .A3(n330), .A4(n1466), .A5(n843), 
        .A6(n1467), .Y(n1871) );
  OA222X1_HVT U2066 ( .A1(n1330), .A2(n1468), .A3(n585), .A4(n1469), .A5(n1470), .A6(n100), .Y(n1870) );
  OA222X1_HVT U2067 ( .A1(n2048), .A2(n1447), .A3(n586), .A4(n1471), .A5(n1000), .A6(n1472), .Y(n1869) );
  MUX21X1_HVT U2068 ( .A1(n2039), .A2(keyout[74]), .S0(n1457), .Y(n3585) );
  NAND4X0_HVT U2069 ( .A1(n1873), .A2(n1874), .A3(n1875), .A4(n1876), .Y(n3584) );
  OA222X1_HVT U2070 ( .A1(n1331), .A2(n1462), .A3(n331), .A4(n1463), .A5(n844), 
        .A6(n1464), .Y(n1876) );
  OA222X1_HVT U2071 ( .A1(n1332), .A2(n1465), .A3(n332), .A4(n1466), .A5(n845), 
        .A6(n1467), .Y(n1875) );
  OA222X1_HVT U2072 ( .A1(n1333), .A2(n1468), .A3(n587), .A4(n1469), .A5(n1470), .A6(n101), .Y(n1874) );
  OA222X1_HVT U2073 ( .A1(n2046), .A2(n1447), .A3(n588), .A4(n1471), .A5(n1001), .A6(n1472), .Y(n1873) );
  MUX21X1_HVT U2074 ( .A1(n2037), .A2(keyout[73]), .S0(n1457), .Y(n3583) );
  NAND4X0_HVT U2075 ( .A1(n1877), .A2(n1878), .A3(n1879), .A4(n1880), .Y(n3582) );
  OA222X1_HVT U2076 ( .A1(n1334), .A2(n1462), .A3(n333), .A4(n1463), .A5(n846), 
        .A6(n1464), .Y(n1880) );
  OA222X1_HVT U2077 ( .A1(n1335), .A2(n1465), .A3(n334), .A4(n1466), .A5(n847), 
        .A6(n1467), .Y(n1879) );
  OA222X1_HVT U2078 ( .A1(n1336), .A2(n1468), .A3(n589), .A4(n1469), .A5(n1470), .A6(n102), .Y(n1878) );
  OA222X1_HVT U2079 ( .A1(n2044), .A2(n1447), .A3(n590), .A4(n1471), .A5(n1002), .A6(n1472), .Y(n1877) );
  MUX21X1_HVT U2080 ( .A1(n2035), .A2(keyout[72]), .S0(n1457), .Y(n3581) );
  NAND4X0_HVT U2081 ( .A1(n1881), .A2(n1882), .A3(n1883), .A4(n1884), .Y(n3580) );
  OA222X1_HVT U2082 ( .A1(n1337), .A2(n1462), .A3(n335), .A4(n1463), .A5(n848), 
        .A6(n1464), .Y(n1884) );
  OA222X1_HVT U2083 ( .A1(n1338), .A2(n1465), .A3(n336), .A4(n1466), .A5(n849), 
        .A6(n1467), .Y(n1883) );
  OA222X1_HVT U2084 ( .A1(n1339), .A2(n1468), .A3(n591), .A4(n1469), .A5(n1470), .A6(n103), .Y(n1882) );
  OA222X1_HVT U2085 ( .A1(n2042), .A2(n1447), .A3(n592), .A4(n1471), .A5(n1003), .A6(n1472), .Y(n1881) );
  MUX21X1_HVT U2086 ( .A1(n2033), .A2(keyout[71]), .S0(n1457), .Y(n3579) );
  NAND4X0_HVT U2087 ( .A1(n1885), .A2(n1886), .A3(n1887), .A4(n1888), .Y(n3578) );
  OA222X1_HVT U2088 ( .A1(n1340), .A2(n1462), .A3(n337), .A4(n1463), .A5(n850), 
        .A6(n1464), .Y(n1888) );
  OA222X1_HVT U2089 ( .A1(n1341), .A2(n1465), .A3(n338), .A4(n1466), .A5(n851), 
        .A6(n1467), .Y(n1887) );
  OA222X1_HVT U2090 ( .A1(n1342), .A2(n1468), .A3(n593), .A4(n1469), .A5(n1470), .A6(n104), .Y(n1886) );
  OA222X1_HVT U2091 ( .A1(n2040), .A2(n1447), .A3(n594), .A4(n1471), .A5(n1004), .A6(n1472), .Y(n1885) );
  MUX21X1_HVT U2092 ( .A1(n2031), .A2(keyout[70]), .S0(n1457), .Y(n3577) );
  NAND4X0_HVT U2093 ( .A1(n1889), .A2(n1890), .A3(n1891), .A4(n1892), .Y(n3576) );
  OA222X1_HVT U2094 ( .A1(n1343), .A2(n1462), .A3(n339), .A4(n1463), .A5(n852), 
        .A6(n1464), .Y(n1892) );
  OA222X1_HVT U2095 ( .A1(n1344), .A2(n1465), .A3(n340), .A4(n1466), .A5(n853), 
        .A6(n1467), .Y(n1891) );
  OA222X1_HVT U2096 ( .A1(n1345), .A2(n1468), .A3(n595), .A4(n1469), .A5(n1470), .A6(n105), .Y(n1890) );
  OA222X1_HVT U2097 ( .A1(n2038), .A2(n1447), .A3(n596), .A4(n1471), .A5(n1005), .A6(n1472), .Y(n1889) );
  MUX21X1_HVT U2098 ( .A1(n2029), .A2(keyout[69]), .S0(n1457), .Y(n3575) );
  NAND4X0_HVT U2099 ( .A1(n1893), .A2(n1894), .A3(n1895), .A4(n1896), .Y(n3574) );
  OA222X1_HVT U2100 ( .A1(n1346), .A2(n1462), .A3(n341), .A4(n1463), .A5(n854), 
        .A6(n1464), .Y(n1896) );
  OA222X1_HVT U2101 ( .A1(n1347), .A2(n1465), .A3(n342), .A4(n1466), .A5(n855), 
        .A6(n1467), .Y(n1895) );
  OA222X1_HVT U2102 ( .A1(n1348), .A2(n1468), .A3(n597), .A4(n1469), .A5(n1470), .A6(n106), .Y(n1894) );
  OA222X1_HVT U2103 ( .A1(n2036), .A2(n1447), .A3(n598), .A4(n1471), .A5(n1006), .A6(n1472), .Y(n1893) );
  MUX21X1_HVT U2104 ( .A1(n2027), .A2(keyout[68]), .S0(n1457), .Y(n3573) );
  NAND4X0_HVT U2105 ( .A1(n1897), .A2(n1898), .A3(n1899), .A4(n1900), .Y(n3572) );
  OA222X1_HVT U2106 ( .A1(n1349), .A2(n1462), .A3(n343), .A4(n1463), .A5(n856), 
        .A6(n1464), .Y(n1900) );
  OA222X1_HVT U2107 ( .A1(n1350), .A2(n1465), .A3(n344), .A4(n1466), .A5(n857), 
        .A6(n1467), .Y(n1899) );
  OA222X1_HVT U2108 ( .A1(n1351), .A2(n1468), .A3(n599), .A4(n1469), .A5(n1470), .A6(n107), .Y(n1898) );
  OA222X1_HVT U2109 ( .A1(n2034), .A2(n1447), .A3(n600), .A4(n1471), .A5(n1007), .A6(n1472), .Y(n1897) );
  MUX21X1_HVT U2110 ( .A1(n2025), .A2(keyout[67]), .S0(n1457), .Y(n3571) );
  NAND4X0_HVT U2111 ( .A1(n1901), .A2(n1902), .A3(n1903), .A4(n1904), .Y(n3570) );
  OA222X1_HVT U2112 ( .A1(n1352), .A2(n1462), .A3(n345), .A4(n1463), .A5(n858), 
        .A6(n1464), .Y(n1904) );
  OA222X1_HVT U2113 ( .A1(n1353), .A2(n1465), .A3(n346), .A4(n1466), .A5(n859), 
        .A6(n1467), .Y(n1903) );
  OA222X1_HVT U2114 ( .A1(n1354), .A2(n1468), .A3(n601), .A4(n1469), .A5(n1470), .A6(n108), .Y(n1902) );
  OA222X1_HVT U2115 ( .A1(n2032), .A2(n1447), .A3(n602), .A4(n1471), .A5(n1008), .A6(n1472), .Y(n1901) );
  MUX21X1_HVT U2116 ( .A1(n2023), .A2(keyout[66]), .S0(n1457), .Y(n3569) );
  NAND4X0_HVT U2117 ( .A1(n1905), .A2(n1906), .A3(n1907), .A4(n1908), .Y(n3568) );
  OA222X1_HVT U2118 ( .A1(n1355), .A2(n1462), .A3(n347), .A4(n1463), .A5(n860), 
        .A6(n1464), .Y(n1908) );
  OA222X1_HVT U2119 ( .A1(n1356), .A2(n1465), .A3(n348), .A4(n1466), .A5(n861), 
        .A6(n1467), .Y(n1907) );
  OA222X1_HVT U2120 ( .A1(n1357), .A2(n1468), .A3(n603), .A4(n1469), .A5(n1470), .A6(n109), .Y(n1906) );
  OA222X1_HVT U2121 ( .A1(n2030), .A2(n1447), .A3(n604), .A4(n1471), .A5(n1009), .A6(n1472), .Y(n1905) );
  MUX21X1_HVT U2122 ( .A1(n2021), .A2(keyout[65]), .S0(n1457), .Y(n3567) );
  NAND4X0_HVT U2123 ( .A1(n1909), .A2(n1910), .A3(n1911), .A4(n1912), .Y(n3566) );
  OA222X1_HVT U2124 ( .A1(n1358), .A2(n1462), .A3(n349), .A4(n1463), .A5(n862), 
        .A6(n1464), .Y(n1912) );
  OA222X1_HVT U2125 ( .A1(n1359), .A2(n1465), .A3(n350), .A4(n1466), .A5(n863), 
        .A6(n1467), .Y(n1911) );
  OA222X1_HVT U2126 ( .A1(n1360), .A2(n1468), .A3(n605), .A4(n1469), .A5(n1470), .A6(n110), .Y(n1910) );
  OA222X1_HVT U2127 ( .A1(n2028), .A2(n1447), .A3(n606), .A4(n1471), .A5(n1010), .A6(n1472), .Y(n1909) );
  MUX21X1_HVT U2128 ( .A1(n2019), .A2(keyout[64]), .S0(n1457), .Y(n3565) );
  NAND4X0_HVT U2129 ( .A1(n1913), .A2(n1914), .A3(n1915), .A4(n1916), .Y(n3564) );
  OA222X1_HVT U2130 ( .A1(n1361), .A2(n1462), .A3(n351), .A4(n1463), .A5(n864), 
        .A6(n1464), .Y(n1916) );
  OA222X1_HVT U2131 ( .A1(n1362), .A2(n1465), .A3(n352), .A4(n1466), .A5(n865), 
        .A6(n1467), .Y(n1915) );
  OA222X1_HVT U2132 ( .A1(n1363), .A2(n1468), .A3(n607), .A4(n1469), .A5(n1470), .A6(n111), .Y(n1914) );
  OA222X1_HVT U2133 ( .A1(n2026), .A2(n1447), .A3(n608), .A4(n1471), .A5(n1011), .A6(n1472), .Y(n1913) );
  MUX21X1_HVT U2134 ( .A1(n2017), .A2(keyout[63]), .S0(n1457), .Y(n3563) );
  NAND4X0_HVT U2135 ( .A1(n1917), .A2(n1918), .A3(n1919), .A4(n1920), .Y(n3562) );
  OA222X1_HVT U2136 ( .A1(n1364), .A2(n1462), .A3(n353), .A4(n1463), .A5(n866), 
        .A6(n1464), .Y(n1920) );
  OA222X1_HVT U2137 ( .A1(n1365), .A2(n1465), .A3(n354), .A4(n1466), .A5(n867), 
        .A6(n1467), .Y(n1919) );
  OA222X1_HVT U2138 ( .A1(n1366), .A2(n1468), .A3(n609), .A4(n1469), .A5(n1470), .A6(n112), .Y(n1918) );
  OA222X1_HVT U2139 ( .A1(n2024), .A2(n1447), .A3(n610), .A4(n1471), .A5(n1012), .A6(n1472), .Y(n1917) );
  MUX21X1_HVT U2140 ( .A1(n2015), .A2(keyout[62]), .S0(n1457), .Y(n3561) );
  NAND4X0_HVT U2141 ( .A1(n1921), .A2(n1922), .A3(n1923), .A4(n1924), .Y(n3560) );
  OA222X1_HVT U2142 ( .A1(n1367), .A2(n1462), .A3(n355), .A4(n1463), .A5(n868), 
        .A6(n1464), .Y(n1924) );
  OA222X1_HVT U2143 ( .A1(n1368), .A2(n1465), .A3(n356), .A4(n1466), .A5(n869), 
        .A6(n1467), .Y(n1923) );
  OA222X1_HVT U2144 ( .A1(n1369), .A2(n1468), .A3(n611), .A4(n1469), .A5(n1470), .A6(n113), .Y(n1922) );
  OA222X1_HVT U2145 ( .A1(n2022), .A2(n1447), .A3(n612), .A4(n1471), .A5(n1013), .A6(n1472), .Y(n1921) );
  MUX21X1_HVT U2146 ( .A1(n2013), .A2(keyout[61]), .S0(n1457), .Y(n3559) );
  NAND4X0_HVT U2147 ( .A1(n1925), .A2(n1926), .A3(n1927), .A4(n1928), .Y(n3558) );
  OA222X1_HVT U2148 ( .A1(n1370), .A2(n1462), .A3(n357), .A4(n1463), .A5(n870), 
        .A6(n1464), .Y(n1928) );
  OA222X1_HVT U2149 ( .A1(n1371), .A2(n1465), .A3(n358), .A4(n1466), .A5(n871), 
        .A6(n1467), .Y(n1927) );
  OA222X1_HVT U2150 ( .A1(n1372), .A2(n1468), .A3(n613), .A4(n1469), .A5(n1470), .A6(n114), .Y(n1926) );
  OA222X1_HVT U2151 ( .A1(n2020), .A2(n1447), .A3(n614), .A4(n1471), .A5(n1014), .A6(n1472), .Y(n1925) );
  MUX21X1_HVT U2152 ( .A1(n2011), .A2(keyout[60]), .S0(n1457), .Y(n3557) );
  NAND4X0_HVT U2153 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .Y(n3556) );
  OA222X1_HVT U2154 ( .A1(n1373), .A2(n1462), .A3(n359), .A4(n1463), .A5(n872), 
        .A6(n1464), .Y(n1932) );
  OA222X1_HVT U2155 ( .A1(n1374), .A2(n1465), .A3(n360), .A4(n1466), .A5(n873), 
        .A6(n1467), .Y(n1931) );
  OA222X1_HVT U2156 ( .A1(n1375), .A2(n1468), .A3(n615), .A4(n1469), .A5(n1470), .A6(n115), .Y(n1930) );
  OA222X1_HVT U2157 ( .A1(n2018), .A2(n1447), .A3(n616), .A4(n1471), .A5(n1015), .A6(n1472), .Y(n1929) );
  MUX21X1_HVT U2158 ( .A1(n2009), .A2(keyout[59]), .S0(n1457), .Y(n3555) );
  NAND4X0_HVT U2159 ( .A1(n1933), .A2(n1934), .A3(n1935), .A4(n1936), .Y(n3554) );
  OA222X1_HVT U2160 ( .A1(n1376), .A2(n1462), .A3(n361), .A4(n1463), .A5(n874), 
        .A6(n1464), .Y(n1936) );
  OA222X1_HVT U2161 ( .A1(n1377), .A2(n1465), .A3(n362), .A4(n1466), .A5(n875), 
        .A6(n1467), .Y(n1935) );
  OA222X1_HVT U2162 ( .A1(n1378), .A2(n1468), .A3(n617), .A4(n1469), .A5(n1470), .A6(n116), .Y(n1934) );
  OA222X1_HVT U2163 ( .A1(n2016), .A2(n1447), .A3(n618), .A4(n1471), .A5(n1016), .A6(n1472), .Y(n1933) );
  MUX21X1_HVT U2164 ( .A1(n2007), .A2(keyout[58]), .S0(n1457), .Y(n3553) );
  NAND4X0_HVT U2165 ( .A1(n1937), .A2(n1938), .A3(n1939), .A4(n1940), .Y(n3552) );
  OA222X1_HVT U2166 ( .A1(n1379), .A2(n1462), .A3(n363), .A4(n1463), .A5(n876), 
        .A6(n1464), .Y(n1940) );
  OA222X1_HVT U2167 ( .A1(n1380), .A2(n1465), .A3(n364), .A4(n1466), .A5(n877), 
        .A6(n1467), .Y(n1939) );
  OA222X1_HVT U2168 ( .A1(n1381), .A2(n1468), .A3(n619), .A4(n1469), .A5(n1470), .A6(n117), .Y(n1938) );
  OA222X1_HVT U2169 ( .A1(n2014), .A2(n1447), .A3(n620), .A4(n1471), .A5(n1017), .A6(n1472), .Y(n1937) );
  MUX21X1_HVT U2170 ( .A1(n2005), .A2(keyout[57]), .S0(n1457), .Y(n3551) );
  NAND4X0_HVT U2171 ( .A1(n1941), .A2(n1942), .A3(n1943), .A4(n1944), .Y(n3550) );
  OA222X1_HVT U2172 ( .A1(n1382), .A2(n1462), .A3(n365), .A4(n1463), .A5(n878), 
        .A6(n1464), .Y(n1944) );
  OA222X1_HVT U2173 ( .A1(n1383), .A2(n1465), .A3(n366), .A4(n1466), .A5(n879), 
        .A6(n1467), .Y(n1943) );
  OA222X1_HVT U2174 ( .A1(n1384), .A2(n1468), .A3(n621), .A4(n1469), .A5(n1470), .A6(n118), .Y(n1942) );
  OA222X1_HVT U2175 ( .A1(n2012), .A2(n1447), .A3(n622), .A4(n1471), .A5(n1018), .A6(n1472), .Y(n1941) );
  MUX21X1_HVT U2176 ( .A1(n2003), .A2(keyout[56]), .S0(n1457), .Y(n3549) );
  NAND4X0_HVT U2177 ( .A1(n1945), .A2(n1946), .A3(n1947), .A4(n1948), .Y(n3548) );
  OA222X1_HVT U2178 ( .A1(n1385), .A2(n1462), .A3(n367), .A4(n1463), .A5(n880), 
        .A6(n1464), .Y(n1948) );
  OA222X1_HVT U2179 ( .A1(n1386), .A2(n1465), .A3(n368), .A4(n1466), .A5(n881), 
        .A6(n1467), .Y(n1947) );
  OA222X1_HVT U2180 ( .A1(n1387), .A2(n1468), .A3(n623), .A4(n1469), .A5(n1470), .A6(n119), .Y(n1946) );
  OA222X1_HVT U2181 ( .A1(n2010), .A2(n1447), .A3(n624), .A4(n1471), .A5(n1019), .A6(n1472), .Y(n1945) );
  MUX21X1_HVT U2182 ( .A1(n2001), .A2(keyout[55]), .S0(n1457), .Y(n3547) );
  NAND4X0_HVT U2183 ( .A1(n1949), .A2(n1950), .A3(n1951), .A4(n1952), .Y(n3546) );
  OA222X1_HVT U2184 ( .A1(n1388), .A2(n1462), .A3(n369), .A4(n1463), .A5(n882), 
        .A6(n1464), .Y(n1952) );
  OA222X1_HVT U2185 ( .A1(n1389), .A2(n1465), .A3(n370), .A4(n1466), .A5(n883), 
        .A6(n1467), .Y(n1951) );
  OA222X1_HVT U2186 ( .A1(n1390), .A2(n1468), .A3(n625), .A4(n1469), .A5(n1470), .A6(n120), .Y(n1950) );
  OA222X1_HVT U2187 ( .A1(n2008), .A2(n1447), .A3(n626), .A4(n1471), .A5(n1020), .A6(n1472), .Y(n1949) );
  MUX21X1_HVT U2188 ( .A1(n1999), .A2(keyout[54]), .S0(n1457), .Y(n3545) );
  NAND4X0_HVT U2189 ( .A1(n1953), .A2(n1954), .A3(n1955), .A4(n1956), .Y(n3544) );
  OA222X1_HVT U2190 ( .A1(n1391), .A2(n1462), .A3(n371), .A4(n1463), .A5(n884), 
        .A6(n1464), .Y(n1956) );
  OA222X1_HVT U2191 ( .A1(n1392), .A2(n1465), .A3(n372), .A4(n1466), .A5(n885), 
        .A6(n1467), .Y(n1955) );
  OA222X1_HVT U2192 ( .A1(n1393), .A2(n1468), .A3(n627), .A4(n1469), .A5(n1470), .A6(n121), .Y(n1954) );
  OA222X1_HVT U2193 ( .A1(n2006), .A2(n1447), .A3(n628), .A4(n1471), .A5(n1021), .A6(n1472), .Y(n1953) );
  MUX21X1_HVT U2194 ( .A1(n1997), .A2(keyout[53]), .S0(n1457), .Y(n3543) );
  NAND4X0_HVT U2195 ( .A1(n1957), .A2(n1958), .A3(n1959), .A4(n1960), .Y(n3542) );
  OA222X1_HVT U2196 ( .A1(n1394), .A2(n1462), .A3(n373), .A4(n1463), .A5(n886), 
        .A6(n1464), .Y(n1960) );
  OA222X1_HVT U2197 ( .A1(n1395), .A2(n1465), .A3(n374), .A4(n1466), .A5(n887), 
        .A6(n1467), .Y(n1959) );
  OA222X1_HVT U2198 ( .A1(n1396), .A2(n1468), .A3(n629), .A4(n1469), .A5(n1470), .A6(n122), .Y(n1958) );
  OA222X1_HVT U2199 ( .A1(n2004), .A2(n1447), .A3(n630), .A4(n1471), .A5(n1022), .A6(n1472), .Y(n1957) );
  MUX21X1_HVT U2200 ( .A1(n1995), .A2(keyout[52]), .S0(n1457), .Y(n3541) );
  NAND4X0_HVT U2201 ( .A1(n1961), .A2(n1962), .A3(n1963), .A4(n1964), .Y(n3540) );
  OA222X1_HVT U2202 ( .A1(n1397), .A2(n1462), .A3(n375), .A4(n1463), .A5(n888), 
        .A6(n1464), .Y(n1964) );
  OA222X1_HVT U2203 ( .A1(n1398), .A2(n1465), .A3(n376), .A4(n1466), .A5(n889), 
        .A6(n1467), .Y(n1963) );
  OA222X1_HVT U2204 ( .A1(n1399), .A2(n1468), .A3(n631), .A4(n1469), .A5(n1470), .A6(n123), .Y(n1962) );
  OA222X1_HVT U2205 ( .A1(n2002), .A2(n1447), .A3(n632), .A4(n1471), .A5(n1023), .A6(n1472), .Y(n1961) );
  MUX21X1_HVT U2206 ( .A1(n1993), .A2(keyout[51]), .S0(n1457), .Y(n3539) );
  NAND4X0_HVT U2207 ( .A1(n1965), .A2(n1966), .A3(n1967), .A4(n1968), .Y(n3538) );
  OA222X1_HVT U2208 ( .A1(n1400), .A2(n1462), .A3(n377), .A4(n1463), .A5(n890), 
        .A6(n1464), .Y(n1968) );
  OA222X1_HVT U2209 ( .A1(n1401), .A2(n1465), .A3(n378), .A4(n1466), .A5(n891), 
        .A6(n1467), .Y(n1967) );
  OA222X1_HVT U2210 ( .A1(n1402), .A2(n1468), .A3(n633), .A4(n1469), .A5(n1470), .A6(n124), .Y(n1966) );
  OA222X1_HVT U2211 ( .A1(n2000), .A2(n1447), .A3(n634), .A4(n1471), .A5(n1024), .A6(n1472), .Y(n1965) );
  MUX21X1_HVT U2212 ( .A1(n1992), .A2(keyout[50]), .S0(n1457), .Y(n3537) );
  NAND4X0_HVT U2213 ( .A1(n1969), .A2(n1970), .A3(n1971), .A4(n1972), .Y(n3536) );
  OA222X1_HVT U2214 ( .A1(n1403), .A2(n1462), .A3(n379), .A4(n1463), .A5(n892), 
        .A6(n1464), .Y(n1972) );
  OA222X1_HVT U2215 ( .A1(n1404), .A2(n1465), .A3(n380), .A4(n1466), .A5(n893), 
        .A6(n1467), .Y(n1971) );
  OA222X1_HVT U2216 ( .A1(n1405), .A2(n1468), .A3(n635), .A4(n1469), .A5(n1470), .A6(n125), .Y(n1970) );
  OA222X1_HVT U2217 ( .A1(n1998), .A2(n1447), .A3(n636), .A4(n1471), .A5(n1025), .A6(n1472), .Y(n1969) );
  MUX21X1_HVT U2218 ( .A1(n1991), .A2(keyout[49]), .S0(n1457), .Y(n3535) );
  NAND4X0_HVT U2219 ( .A1(n1973), .A2(n1974), .A3(n1975), .A4(n1976), .Y(n3534) );
  OA222X1_HVT U2220 ( .A1(n1406), .A2(n1462), .A3(n381), .A4(n1463), .A5(n894), 
        .A6(n1464), .Y(n1976) );
  OA222X1_HVT U2221 ( .A1(n1407), .A2(n1465), .A3(n382), .A4(n1466), .A5(n895), 
        .A6(n1467), .Y(n1975) );
  OA222X1_HVT U2222 ( .A1(n1408), .A2(n1468), .A3(n637), .A4(n1469), .A5(n1470), .A6(n126), .Y(n1974) );
  OA222X1_HVT U2223 ( .A1(n1996), .A2(n1447), .A3(n638), .A4(n1471), .A5(n1026), .A6(n1472), .Y(n1973) );
  MUX21X1_HVT U2224 ( .A1(n1990), .A2(keyout[98]), .S0(n1457), .Y(n3533) );
  NOR2X0_HVT U2225 ( .A1(n1436), .A2(rest), .Y(n1457) );
  NAND3X0_HVT U2226 ( .A1(n1446), .A2(n385), .A3(n3399), .Y(n1436) );
  NAND4X0_HVT U2227 ( .A1(n1977), .A2(n1978), .A3(n1979), .A4(n1980), .Y(n3532) );
  OA222X1_HVT U2228 ( .A1(n1409), .A2(n1462), .A3(n383), .A4(n1463), .A5(n896), 
        .A6(n1464), .Y(n1980) );
  NAND2X0_HVT U2229 ( .A1(n1981), .A2(n1982), .Y(n1464) );
  NAND3X0_HVT U2230 ( .A1(n1983), .A2(n1984), .A3(rount_no[2]), .Y(n1463) );
  NAND3X0_HVT U2231 ( .A1(n1981), .A2(n1985), .A3(rount_no[0]), .Y(n1462) );
  OA222X1_HVT U2232 ( .A1(n1410), .A2(n1465), .A3(n384), .A4(n1466), .A5(n897), 
        .A6(n1467), .Y(n1979) );
  NAND2X0_HVT U2233 ( .A1(n1982), .A2(n1983), .Y(n1467) );
  AND3X1_HVT U2234 ( .A1(n1985), .A2(n1986), .A3(n1984), .Y(n1982) );
  NAND4X0_HVT U2235 ( .A1(rount_no[0]), .A2(n1983), .A3(n1985), .A4(n1986), 
        .Y(n1466) );
  INVX0_HVT U2236 ( .A(rount_no[3]), .Y(n1986) );
  INVX0_HVT U2237 ( .A(rount_no[2]), .Y(n1985) );
  NAND3X0_HVT U2238 ( .A1(rount_no[2]), .A2(n1983), .A3(rount_no[0]), .Y(n1465) );
  OA222X1_HVT U2239 ( .A1(n1411), .A2(n1468), .A3(n639), .A4(n1469), .A5(n1470), .A6(n127), .Y(n1978) );
  NAND3X0_HVT U2240 ( .A1(n1981), .A2(rount_no[2]), .A3(rount_no[0]), .Y(n1470) );
  NAND3X0_HVT U2241 ( .A1(rount_no[2]), .A2(n1984), .A3(n1981), .Y(n1469) );
  NAND3X0_HVT U2242 ( .A1(n1983), .A2(n1984), .A3(rount_no[3]), .Y(n1468) );
  INVX0_HVT U2243 ( .A(rount_no[0]), .Y(n1984) );
  AND2X1_HVT U2244 ( .A1(n1447), .A2(n1987), .Y(n1983) );
  INVX0_HVT U2245 ( .A(rount_no[1]), .Y(n1987) );
  OA222X1_HVT U2246 ( .A1(n1994), .A2(n1447), .A3(n640), .A4(n1471), .A5(n1027), .A6(n1472), .Y(n1977) );
  NAND2X0_HVT U2247 ( .A1(rount_no[3]), .A2(n1981), .Y(n1472) );
  AND2X1_HVT U2248 ( .A1(rount_no[1]), .A2(n1447), .Y(n1981) );
  NAND3X0_HVT U2249 ( .A1(rount_no[0]), .A2(n1447), .A3(rount_no[3]), .Y(n1471) );
  AND4X1_HVT U2250 ( .A1(state[0]), .A2(n1446), .A3(n898), .A4(n3528), .Y(
        n1447) );
  INVX0_HVT U2251 ( .A(rest), .Y(n3528) );
  NOR2X0_HVT U2252 ( .A1(state[2]), .A2(n3398), .Y(n1446) );
endmodule

