
module cde ( clk, rst, cam_start, pass, start_dec, start_enc, master_key, 
        account, data_flash, flash_pass_reg, flash_acc_reg, flash_or_acc_reg, 
        flash_or_acc_sel, pass_enc_reg, new_old_pass_sel, plain_reg, 
        local_master_reg, local_master_sel, out_reg, write_en, write_add, 
        boot_lood, match, dec_done, ready_encryption, write_data_flash, 
        add_flash, final_output );
  input [127:0] pass;
  input [127:0] master_key;
  input [127:0] account;
  input [255:0] data_flash;
  input [3:0] write_add;
  output [255:0] write_data_flash;
  output [3:0] add_flash;
  output [127:0] final_output;
  input clk, rst, cam_start, start_dec, start_enc, flash_pass_reg,
         flash_acc_reg, flash_or_acc_reg, flash_or_acc_sel, pass_enc_reg,
         new_old_pass_sel, plain_reg, local_master_reg, local_master_sel,
         out_reg, write_en, boot_lood;
  output match, dec_done, ready_encryption;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208;
  wire   [127:0] out_flash_or_acc_sel;
  wire   [127:0] out_new_old_pass_sel;
  wire   [127:0] out_decry;
  wire   [127:0] out_local_master_sel;
  wire   [127:0] out_encryption;
  wire   [127:0] out_reg_pass_enc;
  wire   [127:0] out_reg_plain_reg;
  wire   [127:0] out_local_master_reg;
  tri   clk;
  tri   rst;
  tri   cam_start;
  tri   write_en;
  tri   [3:0] write_add;
  tri   match;
  tri   [3:0] match_add;
  tri   [127:0] out_reg_flash_or_acc;

  AO22X1_HVT U6 ( .A1(out_decry[99]), .A2(n139), .A3(pass[99]), .A4(n124), .Y(
        out_new_old_pass_sel[99]) );
  AO22X1_HVT U7 ( .A1(out_decry[98]), .A2(n173), .A3(pass[98]), .A4(n123), .Y(
        out_new_old_pass_sel[98]) );
  AO22X1_HVT U8 ( .A1(out_decry[97]), .A2(n140), .A3(pass[97]), .A4(n37), .Y(
        out_new_old_pass_sel[97]) );
  AO22X1_HVT U9 ( .A1(out_decry[96]), .A2(n166), .A3(pass[96]), .A4(n182), .Y(
        out_new_old_pass_sel[96]) );
  AO22X1_HVT U10 ( .A1(out_decry[95]), .A2(n168), .A3(pass[95]), .A4(n178), 
        .Y(out_new_old_pass_sel[95]) );
  AO22X1_HVT U11 ( .A1(out_decry[94]), .A2(n141), .A3(pass[94]), .A4(n177), 
        .Y(out_new_old_pass_sel[94]) );
  AO22X1_HVT U12 ( .A1(out_decry[93]), .A2(n171), .A3(pass[93]), .A4(n176), 
        .Y(out_new_old_pass_sel[93]) );
  AO22X1_HVT U13 ( .A1(out_decry[92]), .A2(n141), .A3(pass[92]), .A4(n124), 
        .Y(out_new_old_pass_sel[92]) );
  AO22X1_HVT U14 ( .A1(out_decry[91]), .A2(n45), .A3(pass[91]), .A4(n123), .Y(
        out_new_old_pass_sel[91]) );
  AO22X1_HVT U15 ( .A1(out_decry[90]), .A2(n141), .A3(pass[90]), .A4(n180), 
        .Y(out_new_old_pass_sel[90]) );
  AO22X1_HVT U16 ( .A1(out_decry[8]), .A2(n174), .A3(pass[8]), .A4(n28), .Y(
        out_new_old_pass_sel[8]) );
  AO22X1_HVT U17 ( .A1(out_decry[89]), .A2(n167), .A3(pass[89]), .A4(n37), .Y(
        out_new_old_pass_sel[89]) );
  AO22X1_HVT U18 ( .A1(out_decry[88]), .A2(n142), .A3(pass[88]), .A4(n182), 
        .Y(out_new_old_pass_sel[88]) );
  AO22X1_HVT U19 ( .A1(out_decry[87]), .A2(n167), .A3(pass[87]), .A4(n178), 
        .Y(out_new_old_pass_sel[87]) );
  AO22X1_HVT U20 ( .A1(out_decry[86]), .A2(n169), .A3(pass[86]), .A4(n177), 
        .Y(out_new_old_pass_sel[86]) );
  AO22X1_HVT U21 ( .A1(out_decry[85]), .A2(n33), .A3(pass[85]), .A4(n176), .Y(
        out_new_old_pass_sel[85]) );
  AO22X1_HVT U22 ( .A1(out_decry[84]), .A2(n46), .A3(pass[84]), .A4(n124), .Y(
        out_new_old_pass_sel[84]) );
  AO22X1_HVT U23 ( .A1(out_decry[83]), .A2(n24), .A3(pass[83]), .A4(n123), .Y(
        out_new_old_pass_sel[83]) );
  AO22X1_HVT U24 ( .A1(out_decry[82]), .A2(n174), .A3(pass[82]), .A4(n180), 
        .Y(out_new_old_pass_sel[82]) );
  AO22X1_HVT U25 ( .A1(out_decry[81]), .A2(n166), .A3(pass[81]), .A4(n28), .Y(
        out_new_old_pass_sel[81]) );
  AO22X1_HVT U26 ( .A1(out_decry[80]), .A2(n170), .A3(pass[80]), .A4(n178), 
        .Y(out_new_old_pass_sel[80]) );
  AO22X1_HVT U27 ( .A1(out_decry[7]), .A2(n24), .A3(pass[7]), .A4(n182), .Y(
        out_new_old_pass_sel[7]) );
  AO22X1_HVT U28 ( .A1(out_decry[79]), .A2(n171), .A3(pass[79]), .A4(n176), 
        .Y(out_new_old_pass_sel[79]) );
  AO22X1_HVT U29 ( .A1(out_decry[78]), .A2(n166), .A3(pass[78]), .A4(n180), 
        .Y(out_new_old_pass_sel[78]) );
  AO22X1_HVT U30 ( .A1(out_decry[77]), .A2(n169), .A3(pass[77]), .A4(n177), 
        .Y(out_new_old_pass_sel[77]) );
  AO22X1_HVT U31 ( .A1(out_decry[76]), .A2(n138), .A3(pass[76]), .A4(n176), 
        .Y(out_new_old_pass_sel[76]) );
  AO22X1_HVT U32 ( .A1(out_decry[75]), .A2(n29), .A3(pass[75]), .A4(n124), .Y(
        out_new_old_pass_sel[75]) );
  AO22X1_HVT U33 ( .A1(out_decry[74]), .A2(n33), .A3(pass[74]), .A4(n123), .Y(
        out_new_old_pass_sel[74]) );
  AO22X1_HVT U34 ( .A1(out_decry[73]), .A2(n174), .A3(pass[73]), .A4(n185), 
        .Y(out_new_old_pass_sel[73]) );
  AO22X1_HVT U35 ( .A1(out_decry[72]), .A2(n24), .A3(pass[72]), .A4(n179), .Y(
        out_new_old_pass_sel[72]) );
  AO22X1_HVT U36 ( .A1(out_decry[71]), .A2(n140), .A3(pass[71]), .A4(n37), .Y(
        out_new_old_pass_sel[71]) );
  AO22X1_HVT U37 ( .A1(out_decry[70]), .A2(n166), .A3(pass[70]), .A4(n177), 
        .Y(out_new_old_pass_sel[70]) );
  AO22X1_HVT U39 ( .A1(out_decry[69]), .A2(n33), .A3(pass[69]), .A4(n124), .Y(
        out_new_old_pass_sel[69]) );
  AO22X1_HVT U40 ( .A1(out_decry[68]), .A2(n138), .A3(pass[68]), .A4(n123), 
        .Y(out_new_old_pass_sel[68]) );
  AO22X1_HVT U41 ( .A1(out_decry[67]), .A2(n138), .A3(pass[67]), .A4(n123), 
        .Y(out_new_old_pass_sel[67]) );
  AO22X1_HVT U42 ( .A1(out_decry[66]), .A2(n169), .A3(pass[66]), .A4(n180), 
        .Y(out_new_old_pass_sel[66]) );
  AO22X1_HVT U43 ( .A1(out_decry[65]), .A2(n143), .A3(pass[65]), .A4(n182), 
        .Y(out_new_old_pass_sel[65]) );
  AO22X1_HVT U44 ( .A1(out_decry[64]), .A2(n138), .A3(pass[64]), .A4(n178), 
        .Y(out_new_old_pass_sel[64]) );
  AO22X1_HVT U45 ( .A1(out_decry[63]), .A2(n24), .A3(pass[63]), .A4(n177), .Y(
        out_new_old_pass_sel[63]) );
  AO22X1_HVT U46 ( .A1(out_decry[62]), .A2(n173), .A3(pass[62]), .A4(n176), 
        .Y(out_new_old_pass_sel[62]) );
  AO22X1_HVT U47 ( .A1(out_decry[61]), .A2(n50), .A3(pass[61]), .A4(n124), .Y(
        out_new_old_pass_sel[61]) );
  AO22X1_HVT U48 ( .A1(out_decry[60]), .A2(n141), .A3(pass[60]), .A4(n123), 
        .Y(out_new_old_pass_sel[60]) );
  AO22X1_HVT U49 ( .A1(out_decry[5]), .A2(n24), .A3(pass[5]), .A4(n185), .Y(
        out_new_old_pass_sel[5]) );
  AO22X1_HVT U50 ( .A1(out_decry[59]), .A2(n139), .A3(pass[59]), .A4(n179), 
        .Y(out_new_old_pass_sel[59]) );
  AO22X1_HVT U51 ( .A1(out_decry[58]), .A2(n141), .A3(pass[58]), .A4(n178), 
        .Y(out_new_old_pass_sel[58]) );
  AO22X1_HVT U52 ( .A1(out_decry[57]), .A2(n138), .A3(pass[57]), .A4(n179), 
        .Y(out_new_old_pass_sel[57]) );
  AO22X1_HVT U53 ( .A1(out_decry[56]), .A2(n139), .A3(pass[56]), .A4(n178), 
        .Y(out_new_old_pass_sel[56]) );
  AO22X1_HVT U54 ( .A1(out_decry[55]), .A2(n141), .A3(pass[55]), .A4(n177), 
        .Y(out_new_old_pass_sel[55]) );
  AO22X1_HVT U56 ( .A1(out_decry[53]), .A2(n33), .A3(pass[53]), .A4(n124), .Y(
        out_new_old_pass_sel[53]) );
  AO22X1_HVT U57 ( .A1(out_decry[52]), .A2(n140), .A3(pass[52]), .A4(n123), 
        .Y(out_new_old_pass_sel[52]) );
  AO22X1_HVT U58 ( .A1(out_decry[51]), .A2(n143), .A3(pass[51]), .A4(n185), 
        .Y(out_new_old_pass_sel[51]) );
  AO22X1_HVT U59 ( .A1(out_decry[50]), .A2(n173), .A3(pass[50]), .A4(n28), .Y(
        out_new_old_pass_sel[50]) );
  AO22X1_HVT U61 ( .A1(out_decry[49]), .A2(n29), .A3(pass[49]), .A4(n178), .Y(
        out_new_old_pass_sel[49]) );
  AO22X1_HVT U62 ( .A1(out_decry[48]), .A2(n50), .A3(pass[48]), .A4(n177), .Y(
        out_new_old_pass_sel[48]) );
  AO22X1_HVT U63 ( .A1(out_decry[47]), .A2(n139), .A3(pass[47]), .A4(n176), 
        .Y(out_new_old_pass_sel[47]) );
  AO22X1_HVT U64 ( .A1(out_decry[46]), .A2(n170), .A3(pass[46]), .A4(n124), 
        .Y(out_new_old_pass_sel[46]) );
  AO22X1_HVT U65 ( .A1(out_decry[45]), .A2(n171), .A3(pass[45]), .A4(n126), 
        .Y(out_new_old_pass_sel[45]) );
  AO22X1_HVT U66 ( .A1(out_decry[44]), .A2(n170), .A3(pass[44]), .A4(n185), 
        .Y(out_new_old_pass_sel[44]) );
  AO22X1_HVT U67 ( .A1(out_decry[43]), .A2(n140), .A3(pass[43]), .A4(n179), 
        .Y(out_new_old_pass_sel[43]) );
  AO22X1_HVT U68 ( .A1(out_decry[42]), .A2(n141), .A3(pass[42]), .A4(n181), 
        .Y(out_new_old_pass_sel[42]) );
  AO22X1_HVT U69 ( .A1(out_decry[41]), .A2(n169), .A3(pass[41]), .A4(n183), 
        .Y(out_new_old_pass_sel[41]) );
  AO22X1_HVT U70 ( .A1(out_decry[40]), .A2(n50), .A3(pass[40]), .A4(n125), .Y(
        out_new_old_pass_sel[40]) );
  AO22X1_HVT U72 ( .A1(out_decry[39]), .A2(n167), .A3(pass[39]), .A4(n37), .Y(
        out_new_old_pass_sel[39]) );
  AO22X1_HVT U73 ( .A1(out_decry[38]), .A2(n174), .A3(pass[38]), .A4(n182), 
        .Y(out_new_old_pass_sel[38]) );
  AO22X1_HVT U74 ( .A1(out_decry[37]), .A2(n33), .A3(pass[37]), .A4(n181), .Y(
        out_new_old_pass_sel[37]) );
  AO22X1_HVT U75 ( .A1(out_decry[36]), .A2(n169), .A3(pass[36]), .A4(n183), 
        .Y(out_new_old_pass_sel[36]) );
  AO22X1_HVT U76 ( .A1(out_decry[35]), .A2(n167), .A3(pass[35]), .A4(n125), 
        .Y(out_new_old_pass_sel[35]) );
  AO22X1_HVT U77 ( .A1(n171), .A2(out_decry[34]), .A3(pass[34]), .A4(n126), 
        .Y(out_new_old_pass_sel[34]) );
  AO22X1_HVT U78 ( .A1(out_decry[33]), .A2(n143), .A3(pass[33]), .A4(n185), 
        .Y(out_new_old_pass_sel[33]) );
  AO22X1_HVT U79 ( .A1(out_decry[32]), .A2(n173), .A3(pass[32]), .A4(n28), .Y(
        out_new_old_pass_sel[32]) );
  AO22X1_HVT U80 ( .A1(out_decry[31]), .A2(n143), .A3(pass[31]), .A4(n181), 
        .Y(out_new_old_pass_sel[31]) );
  AO22X1_HVT U81 ( .A1(out_decry[30]), .A2(n29), .A3(pass[30]), .A4(n183), .Y(
        out_new_old_pass_sel[30]) );
  AO22X1_HVT U82 ( .A1(out_decry[2]), .A2(n167), .A3(pass[2]), .A4(n125), .Y(
        out_new_old_pass_sel[2]) );
  AO22X1_HVT U83 ( .A1(out_decry[29]), .A2(n143), .A3(pass[29]), .A4(n126), 
        .Y(out_new_old_pass_sel[29]) );
  AO22X1_HVT U84 ( .A1(out_decry[28]), .A2(n166), .A3(pass[28]), .A4(n180), 
        .Y(out_new_old_pass_sel[28]) );
  AO22X1_HVT U85 ( .A1(out_decry[27]), .A2(n29), .A3(pass[27]), .A4(n28), .Y(
        out_new_old_pass_sel[27]) );
  AO22X1_HVT U86 ( .A1(out_decry[26]), .A2(n172), .A3(pass[26]), .A4(n181), 
        .Y(out_new_old_pass_sel[26]) );
  AO22X1_HVT U87 ( .A1(out_decry[25]), .A2(n167), .A3(pass[25]), .A4(n183), 
        .Y(out_new_old_pass_sel[25]) );
  AO22X1_HVT U88 ( .A1(out_decry[24]), .A2(n143), .A3(pass[24]), .A4(n125), 
        .Y(out_new_old_pass_sel[24]) );
  AO22X1_HVT U89 ( .A1(out_decry[23]), .A2(n174), .A3(pass[23]), .A4(n126), 
        .Y(out_new_old_pass_sel[23]) );
  AO22X1_HVT U90 ( .A1(out_decry[22]), .A2(n29), .A3(pass[22]), .A4(n37), .Y(
        out_new_old_pass_sel[22]) );
  AO22X1_HVT U91 ( .A1(out_decry[21]), .A2(n167), .A3(pass[21]), .A4(n179), 
        .Y(out_new_old_pass_sel[21]) );
  AO22X1_HVT U92 ( .A1(out_decry[20]), .A2(n166), .A3(pass[20]), .A4(n181), 
        .Y(out_new_old_pass_sel[20]) );
  AO22X1_HVT U93 ( .A1(out_decry[1]), .A2(n140), .A3(pass[1]), .A4(n184), .Y(
        out_new_old_pass_sel[1]) );
  AO22X1_HVT U94 ( .A1(out_decry[19]), .A2(n169), .A3(pass[19]), .A4(n184), 
        .Y(out_new_old_pass_sel[19]) );
  AO22X1_HVT U95 ( .A1(out_decry[18]), .A2(n170), .A3(pass[18]), .A4(n184), 
        .Y(out_new_old_pass_sel[18]) );
  AO22X1_HVT U96 ( .A1(out_decry[17]), .A2(n50), .A3(pass[17]), .A4(n184), .Y(
        out_new_old_pass_sel[17]) );
  AO22X1_HVT U98 ( .A1(out_decry[15]), .A2(n33), .A3(pass[15]), .A4(n184), .Y(
        out_new_old_pass_sel[15]) );
  AO22X1_HVT U100 ( .A1(out_decry[13]), .A2(n140), .A3(pass[13]), .A4(n184), 
        .Y(out_new_old_pass_sel[13]) );
  AO22X1_HVT U103 ( .A1(out_decry[126]), .A2(n141), .A3(pass[126]), .A4(n179), 
        .Y(out_new_old_pass_sel[126]) );
  AO22X1_HVT U104 ( .A1(out_decry[125]), .A2(n29), .A3(pass[125]), .A4(n181), 
        .Y(out_new_old_pass_sel[125]) );
  AO22X1_HVT U105 ( .A1(out_decry[124]), .A2(n171), .A3(pass[124]), .A4(n183), 
        .Y(out_new_old_pass_sel[124]) );
  AO22X1_HVT U106 ( .A1(out_decry[123]), .A2(n170), .A3(pass[123]), .A4(n125), 
        .Y(out_new_old_pass_sel[123]) );
  AO22X1_HVT U107 ( .A1(out_decry[122]), .A2(n166), .A3(pass[122]), .A4(n126), 
        .Y(out_new_old_pass_sel[122]) );
  AO22X1_HVT U108 ( .A1(out_decry[121]), .A2(n171), .A3(pass[121]), .A4(n180), 
        .Y(out_new_old_pass_sel[121]) );
  AO22X1_HVT U109 ( .A1(out_decry[120]), .A2(n174), .A3(pass[120]), .A4(n182), 
        .Y(out_new_old_pass_sel[120]) );
  AO22X1_HVT U111 ( .A1(out_decry[119]), .A2(n166), .A3(pass[119]), .A4(n183), 
        .Y(out_new_old_pass_sel[119]) );
  AO22X1_HVT U112 ( .A1(out_decry[118]), .A2(n173), .A3(pass[118]), .A4(n125), 
        .Y(out_new_old_pass_sel[118]) );
  AO22X1_HVT U113 ( .A1(out_decry[117]), .A2(n170), .A3(pass[117]), .A4(n126), 
        .Y(out_new_old_pass_sel[117]) );
  AO22X1_HVT U114 ( .A1(out_decry[116]), .A2(n29), .A3(pass[116]), .A4(n37), 
        .Y(out_new_old_pass_sel[116]) );
  AO22X1_HVT U115 ( .A1(out_decry[115]), .A2(n167), .A3(pass[115]), .A4(n28), 
        .Y(out_new_old_pass_sel[115]) );
  AO22X1_HVT U116 ( .A1(out_decry[114]), .A2(n172), .A3(pass[114]), .A4(n181), 
        .Y(out_new_old_pass_sel[114]) );
  AO22X1_HVT U117 ( .A1(out_decry[113]), .A2(n50), .A3(pass[113]), .A4(n183), 
        .Y(out_new_old_pass_sel[113]) );
  AO22X1_HVT U118 ( .A1(out_decry[112]), .A2(n140), .A3(pass[112]), .A4(n125), 
        .Y(out_new_old_pass_sel[112]) );
  AO22X1_HVT U119 ( .A1(out_decry[111]), .A2(n33), .A3(pass[111]), .A4(n126), 
        .Y(out_new_old_pass_sel[111]) );
  AO22X1_HVT U120 ( .A1(out_decry[110]), .A2(n142), .A3(pass[110]), .A4(n185), 
        .Y(out_new_old_pass_sel[110]) );
  AO22X1_HVT U122 ( .A1(out_decry[109]), .A2(n139), .A3(pass[109]), .A4(n181), 
        .Y(out_new_old_pass_sel[109]) );
  AO22X1_HVT U123 ( .A1(out_decry[108]), .A2(n50), .A3(pass[108]), .A4(n183), 
        .Y(out_new_old_pass_sel[108]) );
  AO22X1_HVT U124 ( .A1(out_decry[107]), .A2(n168), .A3(pass[107]), .A4(n125), 
        .Y(out_new_old_pass_sel[107]) );
  AO22X1_HVT U125 ( .A1(out_decry[106]), .A2(n50), .A3(pass[106]), .A4(n82), 
        .Y(out_new_old_pass_sel[106]) );
  AO22X1_HVT U126 ( .A1(out_decry[105]), .A2(n173), .A3(pass[105]), .A4(n82), 
        .Y(out_new_old_pass_sel[105]) );
  AO22X1_HVT U127 ( .A1(out_decry[104]), .A2(n143), .A3(pass[104]), .A4(n82), 
        .Y(out_new_old_pass_sel[104]) );
  AO22X1_HVT U128 ( .A1(out_decry[103]), .A2(n139), .A3(pass[103]), .A4(n82), 
        .Y(out_new_old_pass_sel[103]) );
  AO22X1_HVT U129 ( .A1(out_decry[102]), .A2(n139), .A3(pass[102]), .A4(n82), 
        .Y(out_new_old_pass_sel[102]) );
  AO22X1_HVT U130 ( .A1(out_decry[101]), .A2(n33), .A3(pass[101]), .A4(n186), 
        .Y(out_new_old_pass_sel[101]) );
  AO22X1_HVT U131 ( .A1(out_decry[100]), .A2(n143), .A3(pass[100]), .A4(n186), 
        .Y(out_new_old_pass_sel[100]) );
  AO22X1_HVT U132 ( .A1(out_decry[0]), .A2(n173), .A3(pass[0]), .A4(n186), .Y(
        out_new_old_pass_sel[0]) );
  AND2X1_HVT U133 ( .A1(master_key[9]), .A2(n157), .Y(out_local_master_sel[9])
         );
  AND2X1_HVT U134 ( .A1(master_key[99]), .A2(n162), .Y(
        out_local_master_sel[99]) );
  AND2X1_HVT U135 ( .A1(master_key[98]), .A2(n156), .Y(
        out_local_master_sel[98]) );
  AND2X1_HVT U136 ( .A1(master_key[97]), .A2(n159), .Y(
        out_local_master_sel[97]) );
  AND2X1_HVT U137 ( .A1(master_key[96]), .A2(n161), .Y(
        out_local_master_sel[96]) );
  AND2X1_HVT U138 ( .A1(master_key[95]), .A2(n160), .Y(
        out_local_master_sel[95]) );
  AND2X1_HVT U139 ( .A1(master_key[94]), .A2(n155), .Y(
        out_local_master_sel[94]) );
  AND2X1_HVT U140 ( .A1(master_key[93]), .A2(n163), .Y(
        out_local_master_sel[93]) );
  AND2X1_HVT U141 ( .A1(master_key[92]), .A2(n76), .Y(out_local_master_sel[92]) );
  AND2X1_HVT U142 ( .A1(master_key[91]), .A2(n113), .Y(
        out_local_master_sel[91]) );
  AND2X1_HVT U143 ( .A1(master_key[90]), .A2(n76), .Y(out_local_master_sel[90]) );
  AND2X1_HVT U144 ( .A1(master_key[8]), .A2(n157), .Y(out_local_master_sel[8])
         );
  AND2X1_HVT U145 ( .A1(master_key[89]), .A2(n112), .Y(
        out_local_master_sel[89]) );
  AND2X1_HVT U146 ( .A1(master_key[88]), .A2(n162), .Y(
        out_local_master_sel[88]) );
  AND2X1_HVT U147 ( .A1(master_key[87]), .A2(n160), .Y(
        out_local_master_sel[87]) );
  AND2X1_HVT U148 ( .A1(master_key[86]), .A2(n155), .Y(
        out_local_master_sel[86]) );
  AND2X1_HVT U149 ( .A1(master_key[85]), .A2(n107), .Y(
        out_local_master_sel[85]) );
  AND2X1_HVT U150 ( .A1(master_key[84]), .A2(n160), .Y(
        out_local_master_sel[84]) );
  AND2X1_HVT U151 ( .A1(master_key[83]), .A2(n112), .Y(
        out_local_master_sel[83]) );
  AND2X1_HVT U152 ( .A1(master_key[82]), .A2(n108), .Y(
        out_local_master_sel[82]) );
  AND2X1_HVT U153 ( .A1(master_key[81]), .A2(n158), .Y(
        out_local_master_sel[81]) );
  AND2X1_HVT U154 ( .A1(master_key[80]), .A2(n158), .Y(
        out_local_master_sel[80]) );
  AND2X1_HVT U155 ( .A1(master_key[7]), .A2(n155), .Y(out_local_master_sel[7])
         );
  AND2X1_HVT U156 ( .A1(master_key[79]), .A2(n108), .Y(
        out_local_master_sel[79]) );
  AND2X1_HVT U157 ( .A1(master_key[78]), .A2(n107), .Y(
        out_local_master_sel[78]) );
  AND2X1_HVT U158 ( .A1(master_key[77]), .A2(n160), .Y(
        out_local_master_sel[77]) );
  AND2X1_HVT U159 ( .A1(master_key[76]), .A2(n155), .Y(
        out_local_master_sel[76]) );
  AND2X1_HVT U160 ( .A1(master_key[75]), .A2(n76), .Y(out_local_master_sel[75]) );
  AND2X1_HVT U161 ( .A1(master_key[74]), .A2(n162), .Y(
        out_local_master_sel[74]) );
  AND2X1_HVT U162 ( .A1(master_key[73]), .A2(n156), .Y(
        out_local_master_sel[73]) );
  AND2X1_HVT U163 ( .A1(master_key[72]), .A2(n77), .Y(out_local_master_sel[72]) );
  AND2X1_HVT U164 ( .A1(master_key[71]), .A2(n76), .Y(out_local_master_sel[71]) );
  AND2X1_HVT U165 ( .A1(master_key[70]), .A2(n162), .Y(
        out_local_master_sel[70]) );
  AND2X1_HVT U166 ( .A1(master_key[6]), .A2(n76), .Y(out_local_master_sel[6])
         );
  AND2X1_HVT U167 ( .A1(master_key[69]), .A2(n162), .Y(
        out_local_master_sel[69]) );
  AND2X1_HVT U168 ( .A1(master_key[68]), .A2(n161), .Y(
        out_local_master_sel[68]) );
  AND2X1_HVT U169 ( .A1(master_key[67]), .A2(n160), .Y(
        out_local_master_sel[67]) );
  AND2X1_HVT U170 ( .A1(master_key[66]), .A2(n108), .Y(
        out_local_master_sel[66]) );
  AND2X1_HVT U171 ( .A1(master_key[65]), .A2(n156), .Y(
        out_local_master_sel[65]) );
  AND2X1_HVT U172 ( .A1(master_key[64]), .A2(n159), .Y(
        out_local_master_sel[64]) );
  AND2X1_HVT U173 ( .A1(master_key[63]), .A2(n163), .Y(
        out_local_master_sel[63]) );
  AND2X1_HVT U174 ( .A1(master_key[62]), .A2(n107), .Y(
        out_local_master_sel[62]) );
  AND2X1_HVT U175 ( .A1(master_key[61]), .A2(n108), .Y(
        out_local_master_sel[61]) );
  AND2X1_HVT U176 ( .A1(master_key[60]), .A2(n112), .Y(
        out_local_master_sel[60]) );
  AND2X1_HVT U177 ( .A1(master_key[5]), .A2(n161), .Y(out_local_master_sel[5])
         );
  AND2X1_HVT U178 ( .A1(master_key[59]), .A2(n77), .Y(out_local_master_sel[59]) );
  AND2X1_HVT U179 ( .A1(master_key[58]), .A2(n159), .Y(
        out_local_master_sel[58]) );
  AND2X1_HVT U180 ( .A1(master_key[57]), .A2(n113), .Y(
        out_local_master_sel[57]) );
  AND2X1_HVT U181 ( .A1(master_key[56]), .A2(n163), .Y(
        out_local_master_sel[56]) );
  AND2X1_HVT U182 ( .A1(master_key[55]), .A2(n155), .Y(
        out_local_master_sel[55]) );
  AND2X1_HVT U183 ( .A1(master_key[54]), .A2(n159), .Y(
        out_local_master_sel[54]) );
  AND2X1_HVT U184 ( .A1(master_key[53]), .A2(n108), .Y(
        out_local_master_sel[53]) );
  AND2X1_HVT U185 ( .A1(master_key[52]), .A2(n77), .Y(out_local_master_sel[52]) );
  AND2X1_HVT U186 ( .A1(master_key[51]), .A2(n112), .Y(
        out_local_master_sel[51]) );
  AND2X1_HVT U187 ( .A1(master_key[50]), .A2(n113), .Y(
        out_local_master_sel[50]) );
  AND2X1_HVT U188 ( .A1(master_key[4]), .A2(n157), .Y(out_local_master_sel[4])
         );
  AND2X1_HVT U189 ( .A1(master_key[49]), .A2(n160), .Y(
        out_local_master_sel[49]) );
  AND2X1_HVT U190 ( .A1(master_key[48]), .A2(n159), .Y(
        out_local_master_sel[48]) );
  AND2X1_HVT U191 ( .A1(master_key[47]), .A2(n155), .Y(
        out_local_master_sel[47]) );
  AND2X1_HVT U192 ( .A1(master_key[46]), .A2(n156), .Y(
        out_local_master_sel[46]) );
  AND2X1_HVT U193 ( .A1(master_key[45]), .A2(n163), .Y(
        out_local_master_sel[45]) );
  AND2X1_HVT U194 ( .A1(master_key[44]), .A2(n159), .Y(
        out_local_master_sel[44]) );
  AND2X1_HVT U195 ( .A1(master_key[43]), .A2(n157), .Y(
        out_local_master_sel[43]) );
  AND2X1_HVT U196 ( .A1(master_key[42]), .A2(n156), .Y(
        out_local_master_sel[42]) );
  AND2X1_HVT U197 ( .A1(master_key[41]), .A2(n113), .Y(
        out_local_master_sel[41]) );
  AND2X1_HVT U198 ( .A1(master_key[40]), .A2(n107), .Y(
        out_local_master_sel[40]) );
  AND2X1_HVT U199 ( .A1(master_key[3]), .A2(n163), .Y(out_local_master_sel[3])
         );
  AND2X1_HVT U200 ( .A1(master_key[39]), .A2(n158), .Y(
        out_local_master_sel[39]) );
  AND2X1_HVT U201 ( .A1(master_key[38]), .A2(n157), .Y(
        out_local_master_sel[38]) );
  AND2X1_HVT U202 ( .A1(master_key[37]), .A2(n158), .Y(
        out_local_master_sel[37]) );
  AND2X1_HVT U203 ( .A1(master_key[36]), .A2(n158), .Y(
        out_local_master_sel[36]) );
  AND2X1_HVT U204 ( .A1(master_key[35]), .A2(n158), .Y(
        out_local_master_sel[35]) );
  AND2X1_HVT U205 ( .A1(master_key[34]), .A2(n157), .Y(
        out_local_master_sel[34]) );
  AND2X1_HVT U206 ( .A1(master_key[33]), .A2(n107), .Y(
        out_local_master_sel[33]) );
  AND2X1_HVT U207 ( .A1(master_key[32]), .A2(n107), .Y(
        out_local_master_sel[32]) );
  AND2X1_HVT U208 ( .A1(master_key[31]), .A2(n107), .Y(
        out_local_master_sel[31]) );
  AND2X1_HVT U209 ( .A1(master_key[30]), .A2(n108), .Y(
        out_local_master_sel[30]) );
  AND2X1_HVT U210 ( .A1(master_key[2]), .A2(n108), .Y(out_local_master_sel[2])
         );
  AND2X1_HVT U211 ( .A1(master_key[29]), .A2(n159), .Y(
        out_local_master_sel[29]) );
  AND2X1_HVT U212 ( .A1(master_key[28]), .A2(n157), .Y(
        out_local_master_sel[28]) );
  AND2X1_HVT U213 ( .A1(master_key[27]), .A2(n77), .Y(out_local_master_sel[27]) );
  AND2X1_HVT U214 ( .A1(master_key[26]), .A2(n161), .Y(
        out_local_master_sel[26]) );
  AND2X1_HVT U215 ( .A1(master_key[25]), .A2(n160), .Y(
        out_local_master_sel[25]) );
  AND2X1_HVT U216 ( .A1(master_key[24]), .A2(n76), .Y(out_local_master_sel[24]) );
  AND2X1_HVT U217 ( .A1(master_key[23]), .A2(n76), .Y(out_local_master_sel[23]) );
  AND2X1_HVT U218 ( .A1(master_key[22]), .A2(n161), .Y(
        out_local_master_sel[22]) );
  AND2X1_HVT U219 ( .A1(master_key[21]), .A2(n156), .Y(
        out_local_master_sel[21]) );
  AND2X1_HVT U220 ( .A1(master_key[20]), .A2(n77), .Y(out_local_master_sel[20]) );
  AND2X1_HVT U222 ( .A1(master_key[19]), .A2(n156), .Y(
        out_local_master_sel[19]) );
  AND2X1_HVT U223 ( .A1(master_key[18]), .A2(n161), .Y(
        out_local_master_sel[18]) );
  AND2X1_HVT U224 ( .A1(master_key[17]), .A2(n77), .Y(out_local_master_sel[17]) );
  AND2X1_HVT U225 ( .A1(master_key[16]), .A2(n113), .Y(
        out_local_master_sel[16]) );
  AND2X1_HVT U226 ( .A1(master_key[15]), .A2(n112), .Y(
        out_local_master_sel[15]) );
  AND2X1_HVT U227 ( .A1(master_key[14]), .A2(n162), .Y(
        out_local_master_sel[14]) );
  AND2X1_HVT U228 ( .A1(master_key[13]), .A2(n113), .Y(
        out_local_master_sel[13]) );
  AND2X1_HVT U229 ( .A1(master_key[12]), .A2(n112), .Y(
        out_local_master_sel[12]) );
  AND2X1_HVT U230 ( .A1(master_key[127]), .A2(n112), .Y(
        out_local_master_sel[127]) );
  AND2X1_HVT U231 ( .A1(master_key[126]), .A2(n162), .Y(
        out_local_master_sel[126]) );
  AND2X1_HVT U232 ( .A1(master_key[125]), .A2(n113), .Y(
        out_local_master_sel[125]) );
  AND2X1_HVT U233 ( .A1(master_key[124]), .A2(n155), .Y(
        out_local_master_sel[124]) );
  AND2X1_HVT U234 ( .A1(master_key[123]), .A2(n155), .Y(
        out_local_master_sel[123]) );
  AND2X1_HVT U235 ( .A1(master_key[122]), .A2(n163), .Y(
        out_local_master_sel[122]) );
  AND2X1_HVT U236 ( .A1(master_key[121]), .A2(n163), .Y(
        out_local_master_sel[121]) );
  AND2X1_HVT U237 ( .A1(master_key[120]), .A2(n104), .Y(
        out_local_master_sel[120]) );
  AND2X1_HVT U238 ( .A1(master_key[11]), .A2(n103), .Y(
        out_local_master_sel[11]) );
  AND2X1_HVT U239 ( .A1(master_key[119]), .A2(n154), .Y(
        out_local_master_sel[119]) );
  AND2X1_HVT U240 ( .A1(master_key[118]), .A2(n104), .Y(
        out_local_master_sel[118]) );
  AND2X1_HVT U241 ( .A1(master_key[117]), .A2(n103), .Y(
        out_local_master_sel[117]) );
  AND2X1_HVT U242 ( .A1(master_key[116]), .A2(n154), .Y(
        out_local_master_sel[116]) );
  AND2X1_HVT U243 ( .A1(master_key[115]), .A2(n104), .Y(
        out_local_master_sel[115]) );
  AND2X1_HVT U244 ( .A1(master_key[114]), .A2(n103), .Y(
        out_local_master_sel[114]) );
  AND2X1_HVT U245 ( .A1(master_key[113]), .A2(n154), .Y(
        out_local_master_sel[113]) );
  AND2X1_HVT U246 ( .A1(master_key[112]), .A2(n104), .Y(
        out_local_master_sel[112]) );
  AND2X1_HVT U247 ( .A1(master_key[111]), .A2(n103), .Y(
        out_local_master_sel[111]) );
  AND2X1_HVT U248 ( .A1(master_key[110]), .A2(n154), .Y(
        out_local_master_sel[110]) );
  AND2X1_HVT U249 ( .A1(master_key[10]), .A2(n153), .Y(
        out_local_master_sel[10]) );
  AND2X1_HVT U250 ( .A1(master_key[109]), .A2(n153), .Y(
        out_local_master_sel[109]) );
  AND2X1_HVT U251 ( .A1(master_key[108]), .A2(n153), .Y(
        out_local_master_sel[108]) );
  AND2X1_HVT U252 ( .A1(master_key[107]), .A2(n153), .Y(
        out_local_master_sel[107]) );
  AND2X1_HVT U253 ( .A1(master_key[106]), .A2(n153), .Y(
        out_local_master_sel[106]) );
  AND2X1_HVT U254 ( .A1(master_key[105]), .A2(n153), .Y(
        out_local_master_sel[105]) );
  AND2X1_HVT U255 ( .A1(master_key[104]), .A2(n104), .Y(
        out_local_master_sel[104]) );
  AND2X1_HVT U256 ( .A1(master_key[103]), .A2(n103), .Y(
        out_local_master_sel[103]) );
  AND2X1_HVT U257 ( .A1(master_key[102]), .A2(n154), .Y(
        out_local_master_sel[102]) );
  AND2X1_HVT U258 ( .A1(master_key[101]), .A2(n104), .Y(
        out_local_master_sel[101]) );
  AND2X1_HVT U259 ( .A1(master_key[100]), .A2(n103), .Y(
        out_local_master_sel[100]) );
  AND2X1_HVT U260 ( .A1(master_key[0]), .A2(n154), .Y(out_local_master_sel[0])
         );
  AO22X1_HVT U262 ( .A1(data_flash[227]), .A2(n18), .A3(account[99]), .A4(n128), .Y(out_flash_or_acc_sel[99]) );
  AO22X1_HVT U263 ( .A1(data_flash[226]), .A2(n40), .A3(account[98]), .A4(n128), .Y(out_flash_or_acc_sel[98]) );
  AO22X1_HVT U264 ( .A1(data_flash[225]), .A2(n40), .A3(account[97]), .A4(n128), .Y(out_flash_or_acc_sel[97]) );
  AO22X1_HVT U266 ( .A1(data_flash[223]), .A2(n198), .A3(account[95]), .A4(
        n128), .Y(out_flash_or_acc_sel[95]) );
  AO22X1_HVT U267 ( .A1(data_flash[222]), .A2(n202), .A3(account[94]), .A4(
        n128), .Y(out_flash_or_acc_sel[94]) );
  AO22X1_HVT U268 ( .A1(data_flash[221]), .A2(n147), .A3(account[93]), .A4(
        n128), .Y(out_flash_or_acc_sel[93]) );
  AO22X1_HVT U269 ( .A1(data_flash[220]), .A2(n119), .A3(account[92]), .A4(
        n197), .Y(out_flash_or_acc_sel[92]) );
  AO22X1_HVT U270 ( .A1(data_flash[219]), .A2(n18), .A3(account[91]), .A4(n197), .Y(out_flash_or_acc_sel[91]) );
  AO22X1_HVT U271 ( .A1(data_flash[218]), .A2(n145), .A3(account[90]), .A4(
        n197), .Y(out_flash_or_acc_sel[90]) );
  AO22X1_HVT U273 ( .A1(data_flash[217]), .A2(n19), .A3(account[89]), .A4(n106), .Y(out_flash_or_acc_sel[89]) );
  AO22X1_HVT U274 ( .A1(data_flash[216]), .A2(n129), .A3(account[88]), .A4(
        n106), .Y(out_flash_or_acc_sel[88]) );
  AO22X1_HVT U275 ( .A1(data_flash[215]), .A2(n129), .A3(account[87]), .A4(
        n106), .Y(out_flash_or_acc_sel[87]) );
  AO22X1_HVT U276 ( .A1(data_flash[214]), .A2(n19), .A3(account[86]), .A4(n106), .Y(out_flash_or_acc_sel[86]) );
  AO22X1_HVT U278 ( .A1(data_flash[212]), .A2(n129), .A3(account[84]), .A4(
        n197), .Y(out_flash_or_acc_sel[84]) );
  AO22X1_HVT U279 ( .A1(data_flash[211]), .A2(n206), .A3(account[83]), .A4(
        n106), .Y(out_flash_or_acc_sel[83]) );
  AO22X1_HVT U281 ( .A1(data_flash[209]), .A2(n206), .A3(account[81]), .A4(
        n196), .Y(out_flash_or_acc_sel[81]) );
  AO22X1_HVT U282 ( .A1(data_flash[208]), .A2(n201), .A3(account[80]), .A4(
        n189), .Y(out_flash_or_acc_sel[80]) );
  AO22X1_HVT U284 ( .A1(data_flash[207]), .A2(n146), .A3(account[79]), .A4(n44), .Y(out_flash_or_acc_sel[79]) );
  AO22X1_HVT U285 ( .A1(data_flash[206]), .A2(n68), .A3(account[78]), .A4(n43), 
        .Y(out_flash_or_acc_sel[78]) );
  AO22X1_HVT U287 ( .A1(data_flash[204]), .A2(n14), .A3(account[76]), .A4(n196), .Y(out_flash_or_acc_sel[76]) );
  AO22X1_HVT U288 ( .A1(data_flash[203]), .A2(n68), .A3(account[75]), .A4(n44), 
        .Y(out_flash_or_acc_sel[75]) );
  AO22X1_HVT U289 ( .A1(data_flash[202]), .A2(n18), .A3(account[74]), .A4(n44), 
        .Y(out_flash_or_acc_sel[74]) );
  AO22X1_HVT U290 ( .A1(data_flash[201]), .A2(n14), .A3(account[73]), .A4(n43), 
        .Y(out_flash_or_acc_sel[73]) );
  AO22X1_HVT U291 ( .A1(data_flash[200]), .A2(n39), .A3(account[72]), .A4(n189), .Y(out_flash_or_acc_sel[72]) );
  AO22X1_HVT U292 ( .A1(data_flash[199]), .A2(n199), .A3(account[71]), .A4(n43), .Y(out_flash_or_acc_sel[71]) );
  AO22X1_HVT U293 ( .A1(data_flash[198]), .A2(n198), .A3(account[70]), .A4(
        n114), .Y(out_flash_or_acc_sel[70]) );
  AO22X1_HVT U294 ( .A1(data_flash[134]), .A2(n201), .A3(account[6]), .A4(n195), .Y(out_flash_or_acc_sel[6]) );
  AO22X1_HVT U295 ( .A1(data_flash[197]), .A2(n204), .A3(account[69]), .A4(
        n115), .Y(out_flash_or_acc_sel[69]) );
  AO22X1_HVT U296 ( .A1(data_flash[196]), .A2(n144), .A3(account[68]), .A4(
        n195), .Y(out_flash_or_acc_sel[68]) );
  AO22X1_HVT U297 ( .A1(data_flash[195]), .A2(n145), .A3(account[67]), .A4(
        n191), .Y(out_flash_or_acc_sel[67]) );
  AO22X1_HVT U298 ( .A1(data_flash[194]), .A2(n206), .A3(account[66]), .A4(
        n195), .Y(out_flash_or_acc_sel[66]) );
  AO22X1_HVT U299 ( .A1(data_flash[193]), .A2(n145), .A3(account[65]), .A4(
        n195), .Y(out_flash_or_acc_sel[65]) );
  AO22X1_HVT U300 ( .A1(data_flash[192]), .A2(n201), .A3(account[64]), .A4(
        n195), .Y(out_flash_or_acc_sel[64]) );
  AO22X1_HVT U301 ( .A1(data_flash[191]), .A2(n204), .A3(account[63]), .A4(
        n114), .Y(out_flash_or_acc_sel[63]) );
  AO22X1_HVT U306 ( .A1(data_flash[187]), .A2(n201), .A3(account[59]), .A4(
        n101), .Y(out_flash_or_acc_sel[59]) );
  AO22X1_HVT U308 ( .A1(data_flash[185]), .A2(n40), .A3(account[57]), .A4(n101), .Y(out_flash_or_acc_sel[57]) );
  AO22X1_HVT U309 ( .A1(data_flash[184]), .A2(n144), .A3(account[56]), .A4(n89), .Y(out_flash_or_acc_sel[56]) );
  AO22X1_HVT U310 ( .A1(data_flash[183]), .A2(n205), .A3(account[55]), .A4(
        n101), .Y(out_flash_or_acc_sel[55]) );
  AO22X1_HVT U311 ( .A1(data_flash[182]), .A2(n68), .A3(account[54]), .A4(n101), .Y(out_flash_or_acc_sel[54]) );
  AO22X1_HVT U312 ( .A1(data_flash[181]), .A2(n199), .A3(account[53]), .A4(
        n101), .Y(out_flash_or_acc_sel[53]) );
  AO22X1_HVT U313 ( .A1(data_flash[180]), .A2(n18), .A3(account[52]), .A4(n86), 
        .Y(out_flash_or_acc_sel[52]) );
  AO22X1_HVT U314 ( .A1(data_flash[179]), .A2(n146), .A3(account[51]), .A4(n89), .Y(out_flash_or_acc_sel[51]) );
  AO22X1_HVT U315 ( .A1(data_flash[178]), .A2(n146), .A3(account[50]), .A4(
        n101), .Y(out_flash_or_acc_sel[50]) );
  AO22X1_HVT U317 ( .A1(data_flash[177]), .A2(n68), .A3(account[49]), .A4(n194), .Y(out_flash_or_acc_sel[49]) );
  AO22X1_HVT U318 ( .A1(data_flash[176]), .A2(n205), .A3(account[48]), .A4(n51), .Y(out_flash_or_acc_sel[48]) );
  AO22X1_HVT U319 ( .A1(data_flash[175]), .A2(n146), .A3(account[47]), .A4(n51), .Y(out_flash_or_acc_sel[47]) );
  AO22X1_HVT U320 ( .A1(data_flash[174]), .A2(n119), .A3(account[46]), .A4(
        n194), .Y(out_flash_or_acc_sel[46]) );
  AO22X1_HVT U321 ( .A1(data_flash[173]), .A2(n39), .A3(account[45]), .A4(n194), .Y(out_flash_or_acc_sel[45]) );
  AO22X1_HVT U322 ( .A1(data_flash[172]), .A2(n69), .A3(account[44]), .A4(n187), .Y(out_flash_or_acc_sel[44]) );
  AO22X1_HVT U325 ( .A1(data_flash[169]), .A2(n202), .A3(account[41]), .A4(
        n120), .Y(out_flash_or_acc_sel[41]) );
  AO22X1_HVT U326 ( .A1(data_flash[168]), .A2(n14), .A3(account[40]), .A4(n187), .Y(out_flash_or_acc_sel[40]) );
  AO22X1_HVT U327 ( .A1(data_flash[131]), .A2(n69), .A3(account[3]), .A4(n120), 
        .Y(out_flash_or_acc_sel[3]) );
  AO22X1_HVT U328 ( .A1(data_flash[167]), .A2(n198), .A3(account[39]), .A4(
        n120), .Y(out_flash_or_acc_sel[39]) );
  AO22X1_HVT U329 ( .A1(data_flash[166]), .A2(n201), .A3(account[38]), .A4(n42), .Y(out_flash_or_acc_sel[38]) );
  AO22X1_HVT U330 ( .A1(data_flash[165]), .A2(n39), .A3(account[37]), .A4(n192), .Y(out_flash_or_acc_sel[37]) );
  AO22X1_HVT U331 ( .A1(data_flash[164]), .A2(n205), .A3(account[36]), .A4(n42), .Y(out_flash_or_acc_sel[36]) );
  AO22X1_HVT U332 ( .A1(data_flash[163]), .A2(n202), .A3(account[35]), .A4(
        n192), .Y(out_flash_or_acc_sel[35]) );
  AO22X1_HVT U334 ( .A1(data_flash[161]), .A2(n206), .A3(account[33]), .A4(
        n190), .Y(out_flash_or_acc_sel[33]) );
  AO22X1_HVT U336 ( .A1(data_flash[159]), .A2(n144), .A3(account[31]), .A4(n41), .Y(out_flash_or_acc_sel[31]) );
  AO22X1_HVT U337 ( .A1(data_flash[158]), .A2(n202), .A3(account[30]), .A4(n41), .Y(out_flash_or_acc_sel[30]) );
  AO22X1_HVT U339 ( .A1(data_flash[157]), .A2(n119), .A3(account[29]), .A4(n41), .Y(out_flash_or_acc_sel[29]) );
  AO22X1_HVT U340 ( .A1(data_flash[156]), .A2(n15), .A3(account[28]), .A4(n190), .Y(out_flash_or_acc_sel[28]) );
  AO22X1_HVT U341 ( .A1(data_flash[155]), .A2(n199), .A3(account[27]), .A4(
        n191), .Y(out_flash_or_acc_sel[27]) );
  AO22X1_HVT U343 ( .A1(data_flash[153]), .A2(n146), .A3(account[25]), .A4(
        n191), .Y(out_flash_or_acc_sel[25]) );
  AO22X1_HVT U344 ( .A1(data_flash[152]), .A2(n15), .A3(account[24]), .A4(n191), .Y(out_flash_or_acc_sel[24]) );
  AO22X1_HVT U345 ( .A1(data_flash[151]), .A2(n144), .A3(account[23]), .A4(
        n114), .Y(out_flash_or_acc_sel[23]) );
  AO22X1_HVT U346 ( .A1(data_flash[150]), .A2(n40), .A3(account[22]), .A4(n195), .Y(out_flash_or_acc_sel[22]) );
  AO22X1_HVT U347 ( .A1(data_flash[149]), .A2(n145), .A3(account[21]), .A4(
        n195), .Y(out_flash_or_acc_sel[21]) );
  AO22X1_HVT U348 ( .A1(data_flash[148]), .A2(n204), .A3(account[20]), .A4(
        n195), .Y(out_flash_or_acc_sel[20]) );
  AO22X1_HVT U350 ( .A1(data_flash[147]), .A2(n68), .A3(account[19]), .A4(n115), .Y(out_flash_or_acc_sel[19]) );
  AO22X1_HVT U351 ( .A1(data_flash[146]), .A2(n198), .A3(account[18]), .A4(
        n191), .Y(out_flash_or_acc_sel[18]) );
  AO22X1_HVT U352 ( .A1(data_flash[145]), .A2(n69), .A3(account[17]), .A4(n114), .Y(out_flash_or_acc_sel[17]) );
  AO22X1_HVT U353 ( .A1(data_flash[144]), .A2(n119), .A3(account[16]), .A4(n41), .Y(out_flash_or_acc_sel[16]) );
  AO22X1_HVT U354 ( .A1(data_flash[143]), .A2(n204), .A3(account[15]), .A4(
        n192), .Y(out_flash_or_acc_sel[15]) );
  AO22X1_HVT U356 ( .A1(data_flash[141]), .A2(n202), .A3(account[13]), .A4(n42), .Y(out_flash_or_acc_sel[13]) );
  AO22X1_HVT U357 ( .A1(data_flash[140]), .A2(n205), .A3(account[12]), .A4(
        n190), .Y(out_flash_or_acc_sel[12]) );
  AO22X1_HVT U359 ( .A1(data_flash[254]), .A2(n15), .A3(account[126]), .A4(n42), .Y(out_flash_or_acc_sel[126]) );
  AO22X1_HVT U360 ( .A1(data_flash[253]), .A2(n206), .A3(account[125]), .A4(
        n192), .Y(out_flash_or_acc_sel[125]) );
  AO22X1_HVT U361 ( .A1(data_flash[252]), .A2(n39), .A3(account[124]), .A4(n41), .Y(out_flash_or_acc_sel[124]) );
  AO22X1_HVT U362 ( .A1(data_flash[251]), .A2(n15), .A3(account[123]), .A4(n42), .Y(out_flash_or_acc_sel[123]) );
  AO22X1_HVT U363 ( .A1(data_flash[250]), .A2(n119), .A3(account[122]), .A4(
        n190), .Y(out_flash_or_acc_sel[122]) );
  AO22X1_HVT U364 ( .A1(data_flash[249]), .A2(n14), .A3(account[121]), .A4(
        n192), .Y(out_flash_or_acc_sel[121]) );
  AO22X1_HVT U365 ( .A1(data_flash[248]), .A2(n146), .A3(account[120]), .A4(
        n114), .Y(out_flash_or_acc_sel[120]) );
  AO22X1_HVT U366 ( .A1(data_flash[139]), .A2(n145), .A3(account[11]), .A4(
        n115), .Y(out_flash_or_acc_sel[11]) );
  AO22X1_HVT U367 ( .A1(data_flash[247]), .A2(n69), .A3(account[119]), .A4(
        n191), .Y(out_flash_or_acc_sel[119]) );
  AO22X1_HVT U368 ( .A1(data_flash[246]), .A2(n206), .A3(account[118]), .A4(
        n191), .Y(out_flash_or_acc_sel[118]) );
  AO22X1_HVT U370 ( .A1(data_flash[244]), .A2(n119), .A3(account[116]), .A4(
        n115), .Y(out_flash_or_acc_sel[116]) );
  AO22X1_HVT U372 ( .A1(data_flash[242]), .A2(n69), .A3(account[114]), .A4(
        n191), .Y(out_flash_or_acc_sel[114]) );
  AO22X1_HVT U373 ( .A1(data_flash[241]), .A2(n69), .A3(account[113]), .A4(
        n128), .Y(out_flash_or_acc_sel[113]) );
  AO22X1_HVT U374 ( .A1(data_flash[240]), .A2(n201), .A3(account[112]), .A4(
        n114), .Y(out_flash_or_acc_sel[112]) );
  AO22X1_HVT U375 ( .A1(data_flash[239]), .A2(n199), .A3(account[111]), .A4(
        n114), .Y(out_flash_or_acc_sel[111]) );
  AO22X1_HVT U376 ( .A1(data_flash[238]), .A2(n205), .A3(account[110]), .A4(
        n115), .Y(out_flash_or_acc_sel[110]) );
  AO22X1_HVT U378 ( .A1(data_flash[237]), .A2(n14), .A3(account[109]), .A4(
        n196), .Y(out_flash_or_acc_sel[109]) );
  AO22X1_HVT U379 ( .A1(data_flash[236]), .A2(n144), .A3(account[108]), .A4(
        n196), .Y(out_flash_or_acc_sel[108]) );
  AO22X1_HVT U380 ( .A1(data_flash[235]), .A2(n206), .A3(account[107]), .A4(
        n189), .Y(out_flash_or_acc_sel[107]) );
  AO22X1_HVT U381 ( .A1(data_flash[234]), .A2(n144), .A3(account[106]), .A4(
        n189), .Y(out_flash_or_acc_sel[106]) );
  AO22X1_HVT U382 ( .A1(data_flash[233]), .A2(n40), .A3(account[105]), .A4(n44), .Y(out_flash_or_acc_sel[105]) );
  AO22X1_HVT U384 ( .A1(data_flash[231]), .A2(n68), .A3(account[103]), .A4(n44), .Y(out_flash_or_acc_sel[103]) );
  AO22X1_HVT U385 ( .A1(data_flash[230]), .A2(n201), .A3(account[102]), .A4(
        n43), .Y(out_flash_or_acc_sel[102]) );
  AO22X1_HVT U387 ( .A1(data_flash[228]), .A2(n144), .A3(account[100]), .A4(
        n43), .Y(out_flash_or_acc_sel[100]) );
  AO22X1_HVT U389 ( .A1(n102), .A2(match_add[3]), .A3(write_add[3]), .A4(n105), 
        .Y(add_flash[3]) );
  AO22X1_HVT U390 ( .A1(n127), .A2(match_add[2]), .A3(n208), .A4(write_add[2]), 
        .Y(add_flash[2]) );
  AO22X1_HVT U391 ( .A1(n150), .A2(match_add[1]), .A3(n208), .A4(write_add[1]), 
        .Y(add_flash[1]) );
  AO22X1_HVT U392 ( .A1(n150), .A2(match_add[0]), .A3(n208), .A4(write_add[0]), 
        .Y(add_flash[0]) );
  reg_D_0 reg_flash_or_acc ( .clk(clk), .rst(rst), .enable(flash_or_acc_reg), 
        .in({out_flash_or_acc_sel[127:43], n100, out_flash_or_acc_sel[41:33], 
        n20, out_flash_or_acc_sel[31:3], n80, out_flash_or_acc_sel[1:0]}), 
        .out(out_reg_flash_or_acc) );
  reg_D_6 reg_flash_account ( .clk(clk), .rst(rst), .enable(flash_acc_reg), 
        .in(out_reg_flash_or_acc), .out(write_data_flash[255:128]) );
  reg_D_5 reg_flash_pass ( .clk(clk), .rst(rst), .enable(flash_pass_reg), .in(
        out_encryption), .out(write_data_flash[127:0]) );
  reg_D_4 reg_pass_enc ( .clk(clk), .rst(rst), .enable(pass_enc_reg), .in(
        data_flash[127:0]), .out(out_reg_pass_enc) );
  reg_D_3 reg_plain_reg ( .clk(clk), .rst(rst), .enable(plain_reg), .in({
        out_new_old_pass_sel[127:5], n63, out_new_old_pass_sel[3:0]}), .out(
        out_reg_plain_reg) );
  reg_D_2 reg_local_master ( .clk(clk), .rst(rst), .enable(local_master_reg), 
        .in(out_local_master_sel), .out(out_local_master_reg) );
  reg_D_1 reg_out_reg ( .clk(clk), .rst(rst), .enable(out_reg), .in(
        out_encryption), .out(final_output) );
  cam cam_inst ( .clk(clk), .rst(rst), .start(cam_start), .write_enable(
        write_en), .din(out_reg_flash_or_acc), .write_addr(write_add), .match(
        match), .match_addr(match_add) );
  aes ENC ( .plaintext(out_reg_plain_reg), .key(out_local_master_reg), .clk(
        clk), .reset(rst), .start(start_enc), .cipher_text(out_encryption), 
        .ready(ready_encryption) );
  inv_aes DEC ( .clk(clk), .rest(rst), .start(start_dec), .plaintext1(
        out_reg_pass_enc), .local_key({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cipher_text(out_decry), .done(dec_done) );
  NAND2X0_HVT U2 ( .A1(data_flash[154]), .A2(n68), .Y(n1) );
  NAND2X0_HVT U3 ( .A1(account[26]), .A2(n191), .Y(n2) );
  NAND2X0_HVT U4 ( .A1(n1), .A2(n2), .Y(out_flash_or_acc_sel[26]) );
  NAND2X0_HVT U5 ( .A1(data_flash[162]), .A2(n198), .Y(n3) );
  NAND2X0_HVT U38 ( .A1(account[34]), .A2(n190), .Y(n4) );
  NAND2X0_HVT U55 ( .A1(n3), .A2(n4), .Y(out_flash_or_acc_sel[34]) );
  NAND2X0_HVT U60 ( .A1(data_flash[130]), .A2(n30), .Y(n5) );
  NAND2X0_HVT U71 ( .A1(account[2]), .A2(n101), .Y(n6) );
  NAND2X0_HVT U97 ( .A1(n5), .A2(n6), .Y(n80) );
  INVX0_HVT U99 ( .A(flash_or_acc_sel), .Y(n30) );
  INVX1_HVT U101 ( .A(n188), .Y(n101) );
  NAND2X0_HVT U102 ( .A1(data_flash[137]), .A2(n144), .Y(n7) );
  NAND2X0_HVT U110 ( .A1(n128), .A2(account[9]), .Y(n8) );
  NAND2X0_HVT U121 ( .A1(n7), .A2(n8), .Y(out_flash_or_acc_sel[9]) );
  IBUFFX2_HVT U221 ( .A(n203), .Y(n187) );
  NAND2X0_HVT U261 ( .A1(data_flash[132]), .A2(n207), .Y(n9) );
  NAND2X0_HVT U265 ( .A1(account[4]), .A2(n86), .Y(n10) );
  NAND2X0_HVT U272 ( .A1(n9), .A2(n10), .Y(out_flash_or_acc_sel[4]) );
  INVX0_HVT U277 ( .A(n207), .Y(n86) );
  NAND2X0_HVT U280 ( .A1(data_flash[243]), .A2(n205), .Y(n11) );
  NAND2X0_HVT U283 ( .A1(account[115]), .A2(n114), .Y(n12) );
  NAND2X0_HVT U286 ( .A1(n11), .A2(n12), .Y(out_flash_or_acc_sel[115]) );
  INVX0_HVT U302 ( .A(n137), .Y(n205) );
  INVX0_HVT U303 ( .A(n13), .Y(n114) );
  NBUFFX2_HVT U304 ( .A(n116), .Y(n13) );
  IBUFFX2_HVT U305 ( .A(flash_or_acc_sel), .Y(n116) );
  IBUFFX2_HVT U307 ( .A(n193), .Y(n202) );
  IBUFFX2_HVT U316 ( .A(n193), .Y(n40) );
  IBUFFX2_HVT U323 ( .A(n193), .Y(n119) );
  IBUFFX2_HVT U324 ( .A(n13), .Y(n115) );
  INVX0_HVT U333 ( .A(n13), .Y(n195) );
  IBUFFX2_HVT U335 ( .A(n137), .Y(n14) );
  IBUFFX2_HVT U338 ( .A(n137), .Y(n15) );
  NAND2X0_HVT U342 ( .A1(data_flash[245]), .A2(n145), .Y(n16) );
  NAND2X0_HVT U349 ( .A1(account[117]), .A2(n115), .Y(n17) );
  NAND2X0_HVT U355 ( .A1(n16), .A2(n17), .Y(out_flash_or_acc_sel[117]) );
  IBUFFX2_HVT U358 ( .A(n188), .Y(n120) );
  INVX0_HVT U369 ( .A(n137), .Y(n207) );
  INVX0_HVT U371 ( .A(n137), .Y(n145) );
  NBUFFX2_HVT U377 ( .A(n199), .Y(n18) );
  INVX1_HVT U383 ( .A(n116), .Y(n194) );
  INVX0_HVT U386 ( .A(n105), .Y(n102) );
  NBUFFX2_HVT U388 ( .A(n129), .Y(n19) );
  OAI22X1_HVT U393 ( .A1(n85), .A2(n86), .A3(n87), .A4(n200), .Y(n20) );
  IBUFFX2_HVT U394 ( .A(n207), .Y(n89) );
  NBUFFX2_HVT U395 ( .A(n38), .Y(n21) );
  OAI22X1_HVT U396 ( .A1(n22), .A2(n185), .A3(n23), .A4(n24), .Y(
        out_new_old_pass_sel[54]) );
  IBUFFX16_HVT U397 ( .A(out_decry[54]), .Y(n22) );
  IBUFFX16_HVT U398 ( .A(pass[54]), .Y(n23) );
  INVX0_HVT U399 ( .A(n54), .Y(out_new_old_pass_sel[11]) );
  NBUFFX2_HVT U400 ( .A(n138), .Y(n24) );
  INVX0_HVT U401 ( .A(n96), .Y(n138) );
  OA22X1_HVT U402 ( .A1(n26), .A2(n28), .A3(n27), .A4(n81), .Y(n25) );
  IBUFFX16_HVT U403 ( .A(n25), .Y(out_new_old_pass_sel[6]) );
  IBUFFX16_HVT U404 ( .A(out_decry[6]), .Y(n26) );
  IBUFFX16_HVT U405 ( .A(pass[6]), .Y(n27) );
  INVX0_HVT U406 ( .A(n142), .Y(n28) );
  INVX0_HVT U407 ( .A(n148), .Y(n142) );
  IBUFFX2_HVT U408 ( .A(n21), .Y(n29) );
  OAI22X1_HVT U409 ( .A1(n31), .A2(n184), .A3(n32), .A4(n81), .Y(
        out_new_old_pass_sel[3]) );
  IBUFFX16_HVT U410 ( .A(out_decry[3]), .Y(n31) );
  IBUFFX16_HVT U411 ( .A(pass[3]), .Y(n32) );
  NBUFFX2_HVT U412 ( .A(n97), .Y(n33) );
  INVX0_HVT U413 ( .A(n97), .Y(n175) );
  OA22X1_HVT U414 ( .A1(n35), .A2(n186), .A3(n36), .A4(n81), .Y(n34) );
  IBUFFX16_HVT U415 ( .A(n34), .Y(out_new_old_pass_sel[16]) );
  IBUFFX16_HVT U416 ( .A(out_decry[16]), .Y(n35) );
  IBUFFX16_HVT U417 ( .A(pass[16]), .Y(n36) );
  INVX0_HVT U418 ( .A(n172), .Y(n37) );
  INVX0_HVT U419 ( .A(n142), .Y(n177) );
  INVX0_HVT U420 ( .A(n172), .Y(n185) );
  INVX0_HVT U421 ( .A(n172), .Y(n178) );
  INVX0_HVT U422 ( .A(n172), .Y(n180) );
  NBUFFX2_HVT U423 ( .A(n96), .Y(n38) );
  INVX0_HVT U424 ( .A(n168), .Y(n176) );
  INVX0_HVT U425 ( .A(n148), .Y(n168) );
  NBUFFX2_HVT U426 ( .A(n204), .Y(n39) );
  INVX0_HVT U427 ( .A(n200), .Y(n41) );
  INVX0_HVT U428 ( .A(n200), .Y(n42) );
  AO22X1_HVT U429 ( .A1(data_flash[255]), .A2(n203), .A3(account[127]), .A4(
        n187), .Y(out_flash_or_acc_sel[127]) );
  INVX0_HVT U430 ( .A(n147), .Y(n43) );
  INVX0_HVT U431 ( .A(n147), .Y(n44) );
  INVX0_HVT U432 ( .A(n148), .Y(n45) );
  INVX0_HVT U433 ( .A(n148), .Y(n46) );
  OA22X1_HVT U434 ( .A1(n48), .A2(n56), .A3(n49), .A4(n50), .Y(n47) );
  IBUFFX16_HVT U435 ( .A(n47), .Y(out_new_old_pass_sel[14]) );
  IBUFFX16_HVT U436 ( .A(out_decry[14]), .Y(n48) );
  IBUFFX16_HVT U437 ( .A(pass[14]), .Y(n49) );
  IBUFFX4_HVT U438 ( .A(n170), .Y(n56) );
  NBUFFX2_HVT U439 ( .A(n97), .Y(n50) );
  INVX0_HVT U440 ( .A(n120), .Y(n204) );
  INVX0_HVT U441 ( .A(n203), .Y(n51) );
  INVX0_HVT U442 ( .A(new_old_pass_sel), .Y(n148) );
  INVX0_HVT U443 ( .A(n116), .Y(n193) );
  INVX0_HVT U444 ( .A(n175), .Y(n170) );
  IBUFFX2_HVT U445 ( .A(n175), .Y(n166) );
  INVX0_HVT U446 ( .A(n175), .Y(n167) );
  OAI22X1_HVT U447 ( .A1(n52), .A2(n59), .A3(n53), .A4(n174), .Y(
        out_new_old_pass_sel[12]) );
  IBUFFX16_HVT U448 ( .A(out_decry[12]), .Y(n52) );
  IBUFFX16_HVT U449 ( .A(pass[12]), .Y(n53) );
  IBUFFX2_HVT U450 ( .A(n21), .Y(n140) );
  IBUFFX4_HVT U451 ( .A(n170), .Y(n59) );
  OA22X1_HVT U452 ( .A1(n55), .A2(n56), .A3(n57), .A4(n171), .Y(n54) );
  IBUFFX16_HVT U453 ( .A(out_decry[11]), .Y(n55) );
  IBUFFX16_HVT U454 ( .A(pass[11]), .Y(n57) );
  OAI22X1_HVT U455 ( .A1(n58), .A2(n59), .A3(n60), .A4(n169), .Y(
        out_new_old_pass_sel[10]) );
  IBUFFX16_HVT U456 ( .A(out_decry[10]), .Y(n58) );
  IBUFFX16_HVT U457 ( .A(pass[10]), .Y(n60) );
  NAND2X0_HVT U458 ( .A1(out_decry[127]), .A2(n50), .Y(n61) );
  NAND2X0_HVT U459 ( .A1(pass[127]), .A2(n184), .Y(n62) );
  NAND2X0_HVT U460 ( .A1(n61), .A2(n62), .Y(out_new_old_pass_sel[127]) );
  AO22X1_HVT U461 ( .A1(out_decry[4]), .A2(n171), .A3(pass[4]), .A4(n186), .Y(
        n63) );
  IBUFFX2_HVT U462 ( .A(n45), .Y(n123) );
  NAND2X0_HVT U463 ( .A1(out_decry[9]), .A2(n33), .Y(n64) );
  NAND2X0_HVT U464 ( .A1(pass[9]), .A2(n176), .Y(n65) );
  NAND2X0_HVT U465 ( .A1(n64), .A2(n65), .Y(out_new_old_pass_sel[9]) );
  INVX0_HVT U466 ( .A(flash_or_acc_sel), .Y(n203) );
  INVX0_HVT U467 ( .A(n200), .Y(n190) );
  INVX0_HVT U468 ( .A(n148), .Y(n172) );
  INVX1_HVT U469 ( .A(account[7]), .Y(n91) );
  INVX1_HVT U470 ( .A(account[14]), .Y(n90) );
  INVX1_HVT U471 ( .A(account[32]), .Y(n87) );
  INVX1_HVT U472 ( .A(account[85]), .Y(n71) );
  INVX0_HVT U473 ( .A(data_flash[213]), .Y(n70) );
  INVX0_HVT U474 ( .A(n38), .Y(n171) );
  NAND2X0_HVT U475 ( .A1(data_flash[171]), .A2(n15), .Y(n66) );
  NAND2X0_HVT U476 ( .A1(account[43]), .A2(n194), .Y(n67) );
  NAND2X0_HVT U477 ( .A1(n66), .A2(n67), .Y(out_flash_or_acc_sel[43]) );
  INVX0_HVT U478 ( .A(n136), .Y(n68) );
  INVX0_HVT U479 ( .A(n136), .Y(n69) );
  INVX0_HVT U480 ( .A(new_old_pass_sel), .Y(n96) );
  IBUFFX2_HVT U481 ( .A(n21), .Y(n139) );
  IBUFFX2_HVT U482 ( .A(n38), .Y(n169) );
  OAI22X1_HVT U483 ( .A1(n70), .A2(n101), .A3(n71), .A4(n146), .Y(
        out_flash_or_acc_sel[85]) );
  NAND2X0_HVT U484 ( .A1(data_flash[136]), .A2(n19), .Y(n72) );
  NAND2X0_HVT U485 ( .A1(account[8]), .A2(n197), .Y(n73) );
  NAND2X0_HVT U486 ( .A1(n72), .A2(n73), .Y(out_flash_or_acc_sel[8]) );
  INVX0_HVT U487 ( .A(n136), .Y(n201) );
  NAND2X0_HVT U488 ( .A1(n69), .A2(data_flash[188]), .Y(n74) );
  NAND2X0_HVT U489 ( .A1(account[60]), .A2(n115), .Y(n75) );
  NAND2X0_HVT U490 ( .A1(n74), .A2(n75), .Y(out_flash_or_acc_sel[60]) );
  INVX0_HVT U491 ( .A(n122), .Y(n76) );
  INVX0_HVT U492 ( .A(n122), .Y(n77) );
  IBUFFX2_HVT U493 ( .A(local_master_sel), .Y(n122) );
  AO22X1_HVT U494 ( .A1(data_flash[205]), .A2(n69), .A3(account[77]), .A4(n194), .Y(out_flash_or_acc_sel[77]) );
  INVX0_HVT U495 ( .A(n122), .Y(n160) );
  INVX0_HVT U496 ( .A(n122), .Y(n161) );
  INVX0_HVT U497 ( .A(n122), .Y(n156) );
  INVX0_HVT U498 ( .A(data_flash[160]), .Y(n85) );
  NAND2X0_HVT U499 ( .A1(data_flash[210]), .A2(n40), .Y(n78) );
  NAND2X0_HVT U500 ( .A1(account[82]), .A2(n106), .Y(n79) );
  NAND2X0_HVT U501 ( .A1(n78), .A2(n79), .Y(out_flash_or_acc_sel[82]) );
  IBUFFX2_HVT U502 ( .A(flash_or_acc_sel), .Y(n188) );
  INVX0_HVT U503 ( .A(data_flash[142]), .Y(n88) );
  INVX0_HVT U504 ( .A(n186), .Y(n81) );
  INVX0_HVT U505 ( .A(n81), .Y(n82) );
  IBUFFX2_HVT U506 ( .A(n45), .Y(n184) );
  IBUFFX2_HVT U507 ( .A(n45), .Y(n125) );
  IBUFFX2_HVT U508 ( .A(n168), .Y(n126) );
  INVX1_HVT U509 ( .A(n188), .Y(n137) );
  NAND2X0_HVT U510 ( .A1(data_flash[229]), .A2(n206), .Y(n83) );
  NAND2X0_HVT U511 ( .A1(account[101]), .A2(n196), .Y(n84) );
  NAND2X0_HVT U512 ( .A1(n83), .A2(n84), .Y(out_flash_or_acc_sel[101]) );
  INVX0_HVT U513 ( .A(n136), .Y(n144) );
  INVX0_HVT U514 ( .A(n147), .Y(n189) );
  INVX0_HVT U515 ( .A(n200), .Y(n192) );
  INVX0_HVT U516 ( .A(n46), .Y(n186) );
  OAI22X1_HVT U517 ( .A1(n89), .A2(n88), .A3(n90), .A4(n68), .Y(
        out_flash_or_acc_sel[14]) );
  OR2X2_HVT U518 ( .A1(n91), .A2(n40), .Y(n118) );
  INVX0_HVT U519 ( .A(n187), .Y(n147) );
  NAND2X0_HVT U520 ( .A1(data_flash[224]), .A2(n18), .Y(n92) );
  NAND2X0_HVT U521 ( .A1(account[96]), .A2(n128), .Y(n93) );
  NAND2X0_HVT U522 ( .A1(n92), .A2(n93), .Y(out_flash_or_acc_sel[96]) );
  NAND2X0_HVT U523 ( .A1(data_flash[133]), .A2(n14), .Y(n94) );
  NAND2X0_HVT U524 ( .A1(account[5]), .A2(n89), .Y(n95) );
  NAND2X0_HVT U525 ( .A1(n94), .A2(n95), .Y(out_flash_or_acc_sel[5]) );
  INVX0_HVT U526 ( .A(local_master_sel), .Y(n164) );
  INVX0_HVT U527 ( .A(n121), .Y(n157) );
  INVX0_HVT U528 ( .A(n147), .Y(n196) );
  INVX1_HVT U529 ( .A(master_key[1]), .Y(n109) );
  INVX1_HVT U530 ( .A(account[10]), .Y(n99) );
  INVX0_HVT U531 ( .A(data_flash[138]), .Y(n98) );
  INVX0_HVT U532 ( .A(n137), .Y(n198) );
  INVX0_HVT U533 ( .A(n96), .Y(n97) );
  OAI22X1_HVT U534 ( .A1(n120), .A2(n98), .A3(n99), .A4(n147), .Y(
        out_flash_or_acc_sel[10]) );
  AO22X1_HVT U535 ( .A1(data_flash[232]), .A2(n15), .A3(account[104]), .A4(
        n120), .Y(out_flash_or_acc_sel[104]) );
  AO22X1_HVT U536 ( .A1(data_flash[170]), .A2(n202), .A3(account[42]), .A4(
        n137), .Y(n100) );
  INVX0_HVT U537 ( .A(n165), .Y(n103) );
  INVX0_HVT U538 ( .A(n165), .Y(n104) );
  INVX0_HVT U539 ( .A(n165), .Y(n153) );
  IBUFFX2_HVT U540 ( .A(local_master_sel), .Y(n165) );
  INVX0_HVT U541 ( .A(n127), .Y(n105) );
  NBUFFX2_HVT U542 ( .A(n197), .Y(n106) );
  IBUFFX2_HVT U543 ( .A(n30), .Y(n197) );
  INVX0_HVT U544 ( .A(n121), .Y(n107) );
  INVX0_HVT U545 ( .A(n121), .Y(n108) );
  INVX0_HVT U546 ( .A(n121), .Y(n159) );
  IBUFFX2_HVT U547 ( .A(local_master_sel), .Y(n121) );
  NOR2X4_HVT U548 ( .A1(n109), .A2(n164), .Y(out_local_master_sel[1]) );
  INVX0_HVT U549 ( .A(n149), .Y(n127) );
  NAND2X0_HVT U550 ( .A1(data_flash[190]), .A2(n201), .Y(n110) );
  NAND2X0_HVT U551 ( .A1(account[62]), .A2(n115), .Y(n111) );
  NAND2X0_HVT U552 ( .A1(n110), .A2(n111), .Y(out_flash_or_acc_sel[62]) );
  INVX0_HVT U553 ( .A(n136), .Y(n146) );
  INVX0_HVT U554 ( .A(n30), .Y(n136) );
  INVX0_HVT U555 ( .A(n164), .Y(n112) );
  INVX0_HVT U556 ( .A(n164), .Y(n113) );
  INVX0_HVT U557 ( .A(n13), .Y(n191) );
  INVX0_HVT U558 ( .A(n164), .Y(n155) );
  NAND2X0_HVT U559 ( .A1(data_flash[135]), .A2(n198), .Y(n117) );
  NAND2X0_HVT U560 ( .A1(n117), .A2(n118), .Y(out_flash_or_acc_sel[7]) );
  IBUFFX2_HVT U561 ( .A(n46), .Y(n124) );
  INVX0_HVT U562 ( .A(n164), .Y(n162) );
  INVX0_HVT U563 ( .A(n164), .Y(n163) );
  IBUFFX2_HVT U564 ( .A(n121), .Y(n158) );
  INVX0_HVT U565 ( .A(n149), .Y(n150) );
  IBUFFX2_HVT U566 ( .A(n21), .Y(n173) );
  IBUFFX2_HVT U567 ( .A(n175), .Y(n143) );
  IBUFFX2_HVT U568 ( .A(n38), .Y(n174) );
  IBUFFX2_HVT U569 ( .A(n175), .Y(n141) );
  NBUFFX2_HVT U570 ( .A(n51), .Y(n128) );
  INVX0_HVT U571 ( .A(n194), .Y(n199) );
  NBUFFX2_HVT U572 ( .A(n207), .Y(n129) );
  INVX0_HVT U573 ( .A(n51), .Y(n200) );
  NAND2X0_HVT U574 ( .A1(data_flash[129]), .A2(n146), .Y(n130) );
  NAND2X0_HVT U575 ( .A1(account[1]), .A2(n195), .Y(n131) );
  NAND2X0_HVT U576 ( .A1(n131), .A2(n130), .Y(out_flash_or_acc_sel[1]) );
  NAND2X0_HVT U577 ( .A1(data_flash[186]), .A2(n39), .Y(n132) );
  NAND2X0_HVT U578 ( .A1(account[58]), .A2(n86), .Y(n133) );
  NAND2X0_HVT U579 ( .A1(n133), .A2(n132), .Y(out_flash_or_acc_sel[58]) );
  NAND2X0_HVT U580 ( .A1(data_flash[189]), .A2(n19), .Y(n134) );
  NAND2X0_HVT U581 ( .A1(account[61]), .A2(n115), .Y(n135) );
  NAND2X0_HVT U582 ( .A1(n134), .A2(n135), .Y(out_flash_or_acc_sel[61]) );
  IBUFFX2_HVT U583 ( .A(n46), .Y(n181) );
  IBUFFX2_HVT U584 ( .A(n142), .Y(n182) );
  IBUFFX2_HVT U585 ( .A(n168), .Y(n183) );
  IBUFFX2_HVT U586 ( .A(n142), .Y(n179) );
  INVX0_HVT U587 ( .A(boot_lood), .Y(n208) );
  INVX0_HVT U588 ( .A(boot_lood), .Y(n149) );
  NAND2X0_HVT U589 ( .A1(data_flash[128]), .A2(n119), .Y(n151) );
  NAND2X0_HVT U590 ( .A1(account[0]), .A2(n189), .Y(n152) );
  NAND2X0_HVT U591 ( .A1(n151), .A2(n152), .Y(out_flash_or_acc_sel[0]) );
  INVX0_HVT U592 ( .A(n136), .Y(n206) );
  INVX1_HVT U593 ( .A(n165), .Y(n154) );
endmodule

