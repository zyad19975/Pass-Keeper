
module sbox_5 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n50, n168, n210, n211, n212, n213, n216, n217, n218, n219,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614;

  NAND2X0_HVT U3 ( .A1(n325), .A2(n321), .Y(n612) );
  NAND2X0_HVT U4 ( .A1(n319), .A2(n612), .Y(n611) );
  NAND2X0_HVT U5 ( .A1(n239), .A2(n309), .Y(n609) );
  NAND2X0_HVT U13 ( .A1(n601), .A2(n324), .Y(n602) );
  NAND2X0_HVT U15 ( .A1(n612), .A2(n311), .Y(n599) );
  NAND2X0_HVT U21 ( .A1(n319), .A2(n331), .Y(n593) );
  NAND2X0_HVT U24 ( .A1(n316), .A2(n331), .Y(n591) );
  NAND2X0_HVT U33 ( .A1(n391), .A2(n331), .Y(n582) );
  NAND2X0_HVT U35 ( .A1(n314), .A2(n331), .Y(n580) );
  NAND2X0_HVT U42 ( .A1(n239), .A2(n316), .Y(n573) );
  MUX41X1_HVT U51 ( .A1(n379), .A3(n339), .A2(n355), .A4(n356), .S0(n243), 
        .S1(n333), .Y(n566) );
  NAND2X0_HVT U53 ( .A1(n563), .A2(n572), .Y(n564) );
  NAND2X0_HVT U56 ( .A1(n319), .A2(n259), .Y(n560) );
  MUX41X1_HVT U57 ( .A1(n380), .A3(n595), .A2(n560), .A4(n604), .S0(n243), 
        .S1(n333), .Y(n558) );
  NAND2X0_HVT U58 ( .A1(n324), .A2(n612), .Y(n557) );
  MUX41X1_HVT U59 ( .A1(n297), .A3(n557), .A2(n295), .A4(n354), .S0(n243), 
        .S1(n333), .Y(n556) );
  MUX41X1_HVT U61 ( .A1(n293), .A3(n353), .A2(n264), .A4(n310), .S0(n243), 
        .S1(n333), .Y(n554) );
  NAND2X0_HVT U62 ( .A1(n331), .A2(n322), .Y(n553) );
  MUX41X1_HVT U63 ( .A1(n553), .A3(n346), .A2(n374), .A4(n352), .S0(n243), 
        .S1(n333), .Y(n552) );
  AO21X1_HVT U66 ( .A1(n350), .A2(n305), .A3(n373), .Y(n549) );
  MUX41X1_HVT U68 ( .A1(n348), .A3(n549), .A2(n548), .A4(n550), .S0(n298), 
        .S1(n281), .Y(n547) );
  MUX41X1_HVT U69 ( .A1(n547), .A3(n555), .A2(n551), .A4(n561), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n605), .A2(n542), .Y(n543) );
  MUX41X1_HVT U74 ( .A1(n544), .A3(n589), .A2(n543), .A4(n591), .S0(n299), 
        .S1(n335), .Y(n541) );
  MUX41X1_HVT U75 ( .A1(n377), .A3(n382), .A2(n395), .A4(n358), .S0(n298), 
        .S1(n335), .Y(n540) );
  MUX41X1_HVT U77 ( .A1(n606), .A3(n384), .A2(n539), .A4(n383), .S0(n306), 
        .S1(in[2]), .Y(n538) );
  AND2X1_HVT U83 ( .A1(n326), .A2(n282), .Y(n531) );
  NAND2X0_HVT U85 ( .A1(n331), .A2(n394), .Y(n529) );
  MUX41X1_HVT U86 ( .A1(n382), .A3(n529), .A2(n294), .A4(n290), .S0(n298), 
        .S1(n240), .Y(n528) );
  AO21X1_HVT U93 ( .A1(n308), .A2(n521), .A3(n378), .Y(n522) );
  MUX41X1_HVT U96 ( .A1(n340), .A3(n292), .A2(n381), .A4(n519), .S0(n298), 
        .S1(n240), .Y(n518) );
  MUX41X1_HVT U97 ( .A1(n377), .A3(n292), .A2(n327), .A4(n599), .S0(n298), 
        .S1(n240), .Y(n517) );
  MUX41X1_HVT U98 ( .A1(n517), .A3(n520), .A2(n518), .A4(n525), .S0(in[0]), 
        .S1(n303), .Y(n516) );
  NAND2X0_HVT U101 ( .A1(n512), .A2(n511), .Y(n513) );
  MUX41X1_HVT U103 ( .A1(n612), .A3(n349), .A2(n247), .A4(n580), .S0(n298), 
        .S1(n240), .Y(n509) );
  MUX41X1_HVT U105 ( .A1(n360), .A3(n568), .A2(n508), .A4(n376), .S0(n298), 
        .S1(n240), .Y(n507) );
  MUX41X1_HVT U106 ( .A1(n507), .A3(n510), .A2(n509), .A4(n514), .S0(in[0]), 
        .S1(n303), .Y(n506) );
  MUX21X2_HVT U107 ( .A1(n506), .A2(n516), .S0(in[6]), .Y(out[2]) );
  OA21X1_HVT U109 ( .A1(n367), .A2(n267), .A3(n354), .Y(n504) );
  NAND2X0_HVT U110 ( .A1(n321), .A2(n502), .Y(n503) );
  AND2X1_HVT U115 ( .A1(n328), .A2(n310), .Y(n497) );
  MUX41X1_HVT U116 ( .A1(n602), .A3(n497), .A2(n358), .A4(n584), .S0(n301), 
        .S1(n243), .Y(n496) );
  NAND2X0_HVT U123 ( .A1(n488), .A2(n487), .Y(n489) );
  MUX41X1_HVT U125 ( .A1(n593), .A3(n297), .A2(n348), .A4(n386), .S0(n302), 
        .S1(n243), .Y(n485) );
  AND3X1_HVT U128 ( .A1(n301), .A2(n331), .A3(n282), .Y(n482) );
  MUX41X1_HVT U131 ( .A1(n480), .A3(n482), .A2(n481), .A4(n483), .S0(n305), 
        .S1(n243), .Y(n479) );
  MUX41X1_HVT U132 ( .A1(n479), .A3(n492), .A2(n484), .A4(n498), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  AND2X1_HVT U140 ( .A1(n317), .A2(n330), .Y(n471) );
  MUX41X1_HVT U141 ( .A1(n590), .A3(n368), .A2(n471), .A4(n364), .S0(n299), 
        .S1(n243), .Y(n470) );
  NAND2X0_HVT U146 ( .A1(n327), .A2(n324), .Y(n542) );
  MUX41X1_HVT U147 ( .A1(n388), .A3(n542), .A2(n377), .A4(n569), .S0(n299), 
        .S1(n243), .Y(n465) );
  OA21X1_HVT U151 ( .A1(n575), .A2(n337), .A3(n461), .Y(n462) );
  MUX41X1_HVT U153 ( .A1(n503), .A3(n293), .A2(n320), .A4(n342), .S0(n298), 
        .S1(n240), .Y(n459) );
  AND2X1_HVT U154 ( .A1(n308), .A2(n316), .Y(n458) );
  NAND2X0_HVT U158 ( .A1(n239), .A2(n394), .Y(n454) );
  MUX41X1_HVT U165 ( .A1(n593), .A3(n361), .A2(n569), .A4(n449), .S0(n243), 
        .S1(n332), .Y(n448) );
  NAND2X0_HVT U166 ( .A1(n324), .A2(n259), .Y(n447) );
  NAND2X0_HVT U167 ( .A1(n395), .A2(n331), .Y(n446) );
  MUX41X1_HVT U168 ( .A1(n380), .A3(n317), .A2(n446), .A4(n447), .S0(n332), 
        .S1(n281), .Y(n445) );
  MUX41X1_HVT U172 ( .A1(n442), .A3(n448), .A2(n445), .A4(n450), .S0(in[0]), 
        .S1(n303), .Y(n441) );
  NAND2X0_HVT U174 ( .A1(n326), .A2(n608), .Y(n601) );
  NAND2X0_HVT U177 ( .A1(n325), .A2(n313), .Y(n438) );
  MUX41X1_HVT U179 ( .A1(n587), .A3(n390), .A2(n344), .A4(n389), .S0(n332), 
        .S1(n335), .Y(n436) );
  MUX41X1_HVT U180 ( .A1(n347), .A3(n606), .A2(n602), .A4(n289), .S0(n306), 
        .S1(n332), .Y(n435) );
  MUX41X1_HVT U181 ( .A1(n435), .A3(n437), .A2(n436), .A4(n439), .S0(in[0]), 
        .S1(n304), .Y(n434) );
  OA21X1_HVT U184 ( .A1(n581), .A2(n337), .A3(n357), .Y(n431) );
  MUX41X1_HVT U186 ( .A1(n292), .A3(n576), .A2(n542), .A4(n569), .S0(n332), 
        .S1(n335), .Y(n429) );
  MUX41X1_HVT U189 ( .A1(n427), .A3(n601), .A2(n428), .A4(n376), .S0(n306), 
        .S1(in[2]), .Y(n426) );
  MUX41X1_HVT U193 ( .A1(n573), .A3(n580), .A2(n567), .A4(n424), .S0(n332), 
        .S1(n281), .Y(n423) );
  MUX41X1_HVT U195 ( .A1(n608), .A3(n381), .A2(n323), .A4(n578), .S0(n332), 
        .S1(n335), .Y(n421) );
  AO21X1_HVT U197 ( .A1(n294), .A2(n307), .A3(n378), .Y(n419) );
  OA21X1_HVT U201 ( .A1(n607), .A2(n337), .A3(n368), .Y(n415) );
  MUX41X1_HVT U203 ( .A1(n579), .A3(n370), .A2(n603), .A4(n583), .S0(n332), 
        .S1(n335), .Y(n413) );
  MUX41X1_HVT U204 ( .A1(n560), .A3(n602), .A2(n365), .A4(n592), .S0(n332), 
        .S1(n335), .Y(n412) );
  MUX41X1_HVT U205 ( .A1(n282), .A3(n612), .A2(n390), .A4(n363), .S0(n332), 
        .S1(n281), .Y(n411) );
  NAND2X0_HVT U208 ( .A1(n238), .A2(n319), .Y(n502) );
  NAND2X0_HVT U212 ( .A1(n238), .A2(n318), .Y(n559) );
  NAND2X0_HVT U214 ( .A1(n608), .A2(n331), .Y(n409) );
  NAND2X0_HVT U215 ( .A1(n502), .A2(n318), .Y(n408) );
  AO21X1_HVT U216 ( .A1(n330), .A2(n392), .A3(n337), .Y(n512) );
  NAND2X0_HVT U218 ( .A1(n392), .A2(n327), .Y(n461) );
  NAND2X0_HVT U220 ( .A1(n307), .A2(n409), .Y(n534) );
  MUX41X1_HVT U1 ( .A1(n429), .A3(n426), .A2(n433), .A4(n430), .S0(n23), .S1(
        in[0]), .Y(n425) );
  IBUFFX16_HVT U2 ( .A(n304), .Y(n23) );
  MUX21X1_HVT U6 ( .A1(n415), .A2(n416), .S0(n300), .Y(n414) );
  MUX21X1_HVT U7 ( .A1(n266), .A2(n265), .S0(n233), .Y(n264) );
  INVX0_HVT U8 ( .A(n325), .Y(n233) );
  MUX21X1_HVT U9 ( .A1(n310), .A2(n357), .S0(n168), .Y(n48) );
  MUX21X1_HVT U10 ( .A1(n317), .A2(n375), .S0(n168), .Y(n50) );
  MUX21X1_HVT U11 ( .A1(n48), .A2(n50), .S0(n243), .Y(n469) );
  DELLN2X2_HVT U12 ( .A(n217), .Y(n310) );
  IBUFFX2_HVT U14 ( .A(n502), .Y(n375) );
  IBUFFX2_HVT U16 ( .A(n302), .Y(n168) );
  MUX21X2_HVT U17 ( .A1(n486), .A2(n485), .S0(n210), .Y(n484) );
  IBUFFX16_HVT U18 ( .A(n305), .Y(n210) );
  NBUFFX16_HVT U19 ( .A(in[7]), .Y(n243) );
  MUX41X1_HVT U20 ( .A1(n577), .A3(n389), .A2(n438), .A4(n597), .S0(n211), 
        .S1(n283), .Y(n437) );
  IBUFFX16_HVT U22 ( .A(n299), .Y(n211) );
  INVX0_HVT U23 ( .A(n306), .Y(n283) );
  NAND2X2_HVT U25 ( .A1(n236), .A2(n237), .Y(out[4]) );
  NAND2X0_HVT U26 ( .A1(n493), .A2(n212), .Y(n213) );
  NAND2X0_HVT U27 ( .A1(n496), .A2(n305), .Y(n216) );
  NAND2X0_HVT U28 ( .A1(n213), .A2(n216), .Y(n492) );
  IBUFFX2_HVT U29 ( .A(n305), .Y(n212) );
  XNOR2X2_HVT U30 ( .A1(n312), .A2(n315), .Y(n217) );
  IBUFFX16_HVT U31 ( .A(n217), .Y(n608) );
  INVX1_HVT U32 ( .A(n264), .Y(n598) );
  INVX4_HVT U34 ( .A(n245), .Y(n337) );
  MUX21X1_HVT U36 ( .A1(n291), .A2(n264), .S0(n301), .Y(n481) );
  INVX0_HVT U37 ( .A(in[7]), .Y(n244) );
  IBUFFX2_HVT U38 ( .A(in[7]), .Y(n338) );
  INVX2_HVT U39 ( .A(n337), .Y(n335) );
  MUX41X1_HVT U40 ( .A1(n385), .A3(n601), .A2(n312), .A4(n440), .S0(n218), 
        .S1(n267), .Y(n439) );
  IBUFFX16_HVT U41 ( .A(n338), .Y(n218) );
  NBUFFX4_HVT U43 ( .A(n396), .Y(n312) );
  AO21X2_HVT U44 ( .A1(n302), .A2(n317), .A3(n608), .Y(n494) );
  NAND2X0_HVT U45 ( .A1(n394), .A2(n219), .Y(n231) );
  NAND2X0_HVT U46 ( .A1(n310), .A2(n234), .Y(n232) );
  NAND2X0_HVT U47 ( .A1(n231), .A2(n232), .Y(n607) );
  INVX8_HVT U48 ( .A(n234), .Y(n219) );
  IBUFFX2_HVT U49 ( .A(n238), .Y(n234) );
  NAND2X0_HVT U50 ( .A1(n472), .A2(n235), .Y(n236) );
  NAND2X0_HVT U52 ( .A1(n464), .A2(n280), .Y(n237) );
  IBUFFX2_HVT U54 ( .A(n280), .Y(n235) );
  INVX0_HVT U55 ( .A(n311), .Y(n265) );
  INVX0_HVT U60 ( .A(n330), .Y(n238) );
  INVX0_HVT U64 ( .A(n330), .Y(n239) );
  INVX0_HVT U65 ( .A(n330), .Y(n328) );
  MUX21X1_HVT U67 ( .A1(n577), .A2(n384), .S0(n306), .Y(n456) );
  NBUFFX4_HVT U70 ( .A(n245), .Y(n240) );
  INVX2_HVT U71 ( .A(n244), .Y(n245) );
  MUX21X1_HVT U72 ( .A1(n598), .A2(n289), .S0(n306), .Y(n416) );
  MUX21X2_HVT U76 ( .A1(n434), .A2(n425), .S0(n241), .Y(out[6]) );
  IBUFFX16_HVT U78 ( .A(in[6]), .Y(n241) );
  MUX21X2_HVT U79 ( .A1(n441), .A2(n452), .S0(n242), .Y(out[5]) );
  IBUFFX16_HVT U80 ( .A(n280), .Y(n242) );
  INVX1_HVT U81 ( .A(n247), .Y(n586) );
  MUX21X1_HVT U82 ( .A1(n467), .A2(n468), .S0(n263), .Y(n466) );
  MUX21X2_HVT U84 ( .A1(n537), .A2(n527), .S0(n246), .Y(out[1]) );
  IBUFFX16_HVT U87 ( .A(in[6]), .Y(n246) );
  MUX21X2_HVT U88 ( .A1(n363), .A2(n600), .S0(n302), .Y(n515) );
  MUX21X1_HVT U89 ( .A1(n248), .A2(n610), .S0(n326), .Y(n247) );
  IBUFFX16_HVT U90 ( .A(n314), .Y(n248) );
  MUX41X1_HVT U91 ( .A1(n466), .A3(n470), .A2(n465), .A4(n469), .S0(in[0]), 
        .S1(n249), .Y(n464) );
  IBUFFX16_HVT U92 ( .A(n303), .Y(n249) );
  MUX41X1_HVT U94 ( .A1(n545), .A3(n540), .A2(n541), .A4(n538), .S0(n250), 
        .S1(n251), .Y(n537) );
  IBUFFX16_HVT U95 ( .A(in[0]), .Y(n250) );
  IBUFFX16_HVT U99 ( .A(n303), .Y(n251) );
  MUX21X1_HVT U100 ( .A1(n573), .A2(n569), .S0(n254), .Y(n252) );
  MUX21X2_HVT U102 ( .A1(n526), .A2(n379), .S0(n254), .Y(n253) );
  MUX21X1_HVT U104 ( .A1(n252), .A2(n253), .S0(n240), .Y(n525) );
  IBUFFX2_HVT U108 ( .A(n299), .Y(n254) );
  MUX21X2_HVT U111 ( .A1(n571), .A2(n546), .S0(n300), .Y(n545) );
  MUX41X1_HVT U112 ( .A1(n530), .A3(n533), .A2(n528), .A4(n532), .S0(in[0]), 
        .S1(n255), .Y(n527) );
  IBUFFX16_HVT U113 ( .A(n303), .Y(n255) );
  AND3X1_HVT U114 ( .A1(n321), .A2(n259), .A3(n534), .Y(n535) );
  MUX21X2_HVT U117 ( .A1(n536), .A2(n535), .S0(n302), .Y(n533) );
  NAND2X0_HVT U118 ( .A1(n417), .A2(n256), .Y(n257) );
  NAND2X0_HVT U119 ( .A1(n410), .A2(n280), .Y(n258) );
  NAND2X0_HVT U120 ( .A1(n257), .A2(n258), .Y(out[7]) );
  IBUFFX2_HVT U121 ( .A(n280), .Y(n256) );
  INVX1_HVT U122 ( .A(n377), .Y(n259) );
  INVX1_HVT U124 ( .A(n559), .Y(n377) );
  MUX21X2_HVT U126 ( .A1(n594), .A2(n318), .S0(n308), .Y(n536) );
  IBUFFX2_HVT U127 ( .A(n594), .Y(n356) );
  MUX41X1_HVT U129 ( .A1(n459), .A3(n460), .A2(n453), .A4(n455), .S0(n304), 
        .S1(n262), .Y(n452) );
  MUX41X1_HVT U130 ( .A1(n310), .A3(n602), .A2(n277), .A4(n454), .S0(n268), 
        .S1(n240), .Y(n453) );
  MUX21X1_HVT U133 ( .A1(n456), .A2(n457), .S0(n302), .Y(n455) );
  IBUFFX2_HVT U134 ( .A(in[0]), .Y(n262) );
  INVX2_HVT U135 ( .A(n268), .Y(n332) );
  MUX41X1_HVT U136 ( .A1(n473), .A3(n476), .A2(n475), .A4(n477), .S0(n260), 
        .S1(n261), .Y(n472) );
  IBUFFX16_HVT U137 ( .A(n269), .Y(n260) );
  IBUFFX16_HVT U138 ( .A(n270), .Y(n261) );
  MUX21X2_HVT U139 ( .A1(n474), .A2(n611), .S0(n302), .Y(n473) );
  IBUFFX16_HVT U142 ( .A(n330), .Y(n327) );
  IBUFFX16_HVT U143 ( .A(n301), .Y(n263) );
  IBUFFX2_HVT U144 ( .A(in[1]), .Y(n331) );
  INVX2_HVT U145 ( .A(in[1]), .Y(n330) );
  MUX21X2_HVT U148 ( .A1(n586), .A2(n345), .S0(n308), .Y(n468) );
  XOR2X2_HVT U149 ( .A1(n337), .A2(n588), .Y(n571) );
  IBUFFX16_HVT U150 ( .A(n309), .Y(n266) );
  INVX0_HVT U152 ( .A(n291), .Y(n273) );
  INVX0_HVT U155 ( .A(n271), .Y(n450) );
  INVX1_HVT U156 ( .A(n300), .Y(n268) );
  INVX0_HVT U157 ( .A(n301), .Y(n267) );
  INVX1_HVT U159 ( .A(n304), .Y(n270) );
  INVX1_HVT U160 ( .A(in[0]), .Y(n269) );
  MUX41X1_HVT U161 ( .A1(n357), .A3(n598), .A2(n608), .A4(n531), .S0(n240), 
        .S1(n298), .Y(n530) );
  MUX41X1_HVT U162 ( .A1(n579), .A3(n388), .A2(n582), .A4(n290), .S0(n267), 
        .S1(n338), .Y(n475) );
  IBUFFX2_HVT U163 ( .A(n330), .Y(n329) );
  OA21X2_HVT U164 ( .A1(n295), .A2(n337), .A3(n584), .Y(n443) );
  OA21X2_HVT U169 ( .A1(n343), .A2(n337), .A3(n584), .Y(n467) );
  MUX21X2_HVT U170 ( .A1(n419), .A2(n420), .S0(n268), .Y(n418) );
  INVX1_HVT U171 ( .A(n398), .Y(n389) );
  MUX41X1_HVT U173 ( .A1(n600), .A3(n340), .A2(n356), .A4(n570), .S0(n267), 
        .S1(n337), .Y(n532) );
  MUX41X1_HVT U175 ( .A1(n414), .A3(n412), .A2(n413), .A4(n411), .S0(n269), 
        .S1(n270), .Y(n410) );
  MUX21X2_HVT U176 ( .A1(n592), .A2(n369), .S0(n307), .Y(n474) );
  INVX0_HVT U178 ( .A(n353), .Y(n272) );
  INVX1_HVT U182 ( .A(n451), .Y(n274) );
  MUX41X1_HVT U183 ( .A1(n274), .A3(n273), .A2(n275), .A4(n272), .S0(n267), 
        .S1(n337), .Y(n271) );
  NAND2X0_HVT U185 ( .A1(n608), .A2(n542), .Y(n275) );
  INVX0_HVT U187 ( .A(n285), .Y(n288) );
  INVX0_HVT U188 ( .A(in[6]), .Y(n280) );
  NBUFFX2_HVT U190 ( .A(n217), .Y(n311) );
  INVX0_HVT U191 ( .A(n276), .Y(n476) );
  INVX0_HVT U192 ( .A(n299), .Y(n279) );
  INVX0_HVT U194 ( .A(n588), .Y(n278) );
  INVX0_HVT U196 ( .A(n609), .Y(n277) );
  MUX41X1_HVT U198 ( .A1(n278), .A3(n277), .A2(n317), .A4(n400), .S0(n279), 
        .S1(n338), .Y(n276) );
  INVX2_HVT U199 ( .A(n283), .Y(n281) );
  INVX1_HVT U200 ( .A(n314), .Y(n282) );
  MUX41X1_HVT U202 ( .A1(n317), .A3(n387), .A2(n588), .A4(n574), .S0(n283), 
        .S1(n279), .Y(n422) );
  MUX41X1_HVT U206 ( .A1(n423), .A3(n421), .A2(n422), .A4(n418), .S0(n269), 
        .S1(n270), .Y(n417) );
  MUX41X1_HVT U207 ( .A1(n359), .A3(n371), .A2(n610), .A4(n369), .S0(n338), 
        .S1(n267), .Y(n433) );
  XOR2X1_HVT U209 ( .A1(n279), .A2(n338), .Y(n284) );
  MUX21X2_HVT U210 ( .A1(n293), .A2(n515), .S0(n284), .Y(n514) );
  XOR2X1_HVT U211 ( .A1(n330), .A2(n279), .Y(n285) );
  IBUFFX2_HVT U213 ( .A(n330), .Y(n325) );
  MUX41X1_HVT U217 ( .A1(n499), .A3(n501), .A2(n505), .A4(n504), .S0(n240), 
        .S1(n305), .Y(n498) );
  NAND2X0_HVT U219 ( .A1(n322), .A2(n285), .Y(n286) );
  NAND2X0_HVT U221 ( .A1(n500), .A2(n288), .Y(n287) );
  NAND2X0_HVT U222 ( .A1(n286), .A2(n287), .Y(n499) );
  NBUFFX16_HVT U223 ( .A(n334), .Y(n305) );
  IBUFFX2_HVT U224 ( .A(n330), .Y(n326) );
  MUX21X2_HVT U225 ( .A1(n372), .A2(n389), .S0(n307), .Y(n420) );
  INVX0_HVT U226 ( .A(n338), .Y(n336) );
  INVX0_HVT U227 ( .A(n315), .Y(n393) );
  INVX1_HVT U228 ( .A(n610), .Y(n391) );
  AND2X1_HVT U229 ( .A1(n310), .A2(n559), .Y(n289) );
  INVX1_HVT U230 ( .A(n320), .Y(n395) );
  MUX21X1_HVT U231 ( .A1(n391), .A2(n394), .S0(n305), .Y(n563) );
  MUX21X1_HVT U232 ( .A1(n584), .A2(n503), .S0(n302), .Y(n501) );
  NBUFFX2_HVT U233 ( .A(n610), .Y(n319) );
  MUX21X1_HVT U234 ( .A1(n349), .A2(n392), .S0(n305), .Y(n548) );
  AND2X1_HVT U235 ( .A1(n321), .A2(n542), .Y(n290) );
  MUX21X1_HVT U236 ( .A1(n321), .A2(n311), .S0(n326), .Y(n574) );
  MUX21X1_HVT U237 ( .A1(n310), .A2(n314), .S0(n238), .Y(n511) );
  MUX21X1_HVT U238 ( .A1(n490), .A2(n489), .S0(n308), .Y(n486) );
  MUX21X1_HVT U239 ( .A1(n391), .A2(n395), .S0(n329), .Y(n440) );
  MUX21X1_HVT U240 ( .A1(n394), .A2(n311), .S0(n328), .Y(n451) );
  MUX21X1_HVT U241 ( .A1(n311), .A2(n391), .S0(n327), .Y(n519) );
  MUX21X1_HVT U242 ( .A1(n608), .A2(n392), .S0(n328), .Y(n400) );
  MUX21X1_HVT U243 ( .A1(n608), .A2(n395), .S0(n325), .Y(n590) );
  MUX21X1_HVT U244 ( .A1(n319), .A2(n608), .S0(n328), .Y(n578) );
  MUX21X1_HVT U245 ( .A1(n319), .A2(n318), .S0(n239), .Y(n526) );
  XOR2X1_HVT U246 ( .A1(n608), .A2(n326), .Y(n569) );
  MUX21X1_HVT U247 ( .A1(n309), .A2(n608), .S0(n325), .Y(n403) );
  MUX21X1_HVT U248 ( .A1(n395), .A2(n394), .S0(n238), .Y(n588) );
  MUX21X1_HVT U249 ( .A1(n394), .A2(n391), .S0(n329), .Y(n577) );
  MUX21X1_HVT U250 ( .A1(n309), .A2(n395), .S0(n327), .Y(n575) );
  MUX21X1_HVT U251 ( .A1(n494), .A2(n495), .S0(n307), .Y(n493) );
  MUX21X1_HVT U252 ( .A1(n342), .A2(n365), .S0(n301), .Y(n495) );
  MUX21X1_HVT U253 ( .A1(n362), .A2(n478), .S0(n301), .Y(n477) );
  MUX21X1_HVT U254 ( .A1(n386), .A2(n318), .S0(n307), .Y(n478) );
  MUX21X1_HVT U255 ( .A1(n608), .A2(n314), .S0(n239), .Y(n539) );
  NAND2X0_HVT U256 ( .A1(n312), .A2(n393), .Y(n610) );
  MUX21X1_HVT U257 ( .A1(n391), .A2(n313), .S0(n329), .Y(n401) );
  NBUFFX2_HVT U258 ( .A(n613), .Y(n320) );
  MUX21X1_HVT U259 ( .A1(n394), .A2(n309), .S0(n238), .Y(n581) );
  MUX21X1_HVT U260 ( .A1(n392), .A2(n391), .S0(n327), .Y(n596) );
  MUX21X1_HVT U261 ( .A1(n341), .A2(n491), .S0(n299), .Y(n490) );
  MUX21X1_HVT U262 ( .A1(n313), .A2(n309), .S0(n328), .Y(n491) );
  MUX21X1_HVT U263 ( .A1(n309), .A2(n324), .S0(n238), .Y(n427) );
  MUX21X1_HVT U264 ( .A1(n323), .A2(n321), .S0(n327), .Y(n428) );
  INVX1_HVT U265 ( .A(n317), .Y(n392) );
  INVX1_HVT U266 ( .A(n323), .Y(n394) );
  MUX21X1_HVT U267 ( .A1(n322), .A2(n318), .S0(n239), .Y(n600) );
  MUX21X1_HVT U268 ( .A1(n610), .A2(n324), .S0(n239), .Y(n521) );
  NBUFFX2_HVT U269 ( .A(n613), .Y(n321) );
  NBUFFX2_HVT U270 ( .A(n613), .Y(n322) );
  XOR2X1_HVT U271 ( .A1(n329), .A2(n392), .Y(n570) );
  MUX21X1_HVT U272 ( .A1(n309), .A2(n314), .S0(n325), .Y(n424) );
  XOR2X1_HVT U273 ( .A1(n320), .A2(n325), .Y(n567) );
  XNOR2X1_HVT U274 ( .A1(n610), .A2(n326), .Y(n291) );
  AND2X1_HVT U275 ( .A1(n329), .A2(n395), .Y(n292) );
  MUX21X1_HVT U276 ( .A1(n323), .A2(n318), .S0(n328), .Y(n584) );
  MUX21X1_HVT U277 ( .A1(n309), .A2(n394), .S0(n327), .Y(n604) );
  MUX21X1_HVT U278 ( .A1(n319), .A2(n309), .S0(n328), .Y(n603) );
  MUX21X1_HVT U279 ( .A1(n320), .A2(n313), .S0(n239), .Y(n407) );
  MUX21X1_HVT U280 ( .A1(n320), .A2(n319), .S0(n329), .Y(n399) );
  AND2X1_HVT U281 ( .A1(n324), .A2(n502), .Y(n293) );
  MUX21X1_HVT U282 ( .A1(n318), .A2(n309), .S0(n328), .Y(n405) );
  XNOR2X1_HVT U283 ( .A1(n323), .A2(n239), .Y(n294) );
  MUX21X1_HVT U284 ( .A1(n318), .A2(n324), .S0(n301), .Y(n488) );
  MUX21X1_HVT U285 ( .A1(n318), .A2(n313), .S0(n327), .Y(n544) );
  XOR2X1_HVT U286 ( .A1(n312), .A2(n326), .Y(n589) );
  NBUFFX2_HVT U287 ( .A(n336), .Y(n308) );
  NBUFFX2_HVT U288 ( .A(n336), .Y(n307) );
  NBUFFX2_HVT U289 ( .A(n336), .Y(n306) );
  NBUFFX2_HVT U290 ( .A(n393), .Y(n309) );
  NBUFFX2_HVT U291 ( .A(in[2]), .Y(n299) );
  NBUFFX2_HVT U292 ( .A(in[2]), .Y(n301) );
  NBUFFX2_HVT U293 ( .A(in[2]), .Y(n302) );
  NBUFFX2_HVT U294 ( .A(in[2]), .Y(n300) );
  NBUFFX2_HVT U295 ( .A(n334), .Y(n304) );
  NBUFFX2_HVT U296 ( .A(in[2]), .Y(n298) );
  NBUFFX2_HVT U297 ( .A(n333), .Y(n303) );
  MUX21X1_HVT U298 ( .A1(n217), .A2(n316), .S0(n328), .Y(n592) );
  MUX21X1_HVT U299 ( .A1(n513), .A2(n362), .S0(n301), .Y(n510) );
  MUX21X1_HVT U300 ( .A1(n431), .A2(n432), .S0(n300), .Y(n430) );
  MUX21X1_HVT U301 ( .A1(n529), .A2(n316), .S0(n307), .Y(n432) );
  MUX21X1_HVT U302 ( .A1(n552), .A2(n554), .S0(n300), .Y(n551) );
  XOR2X1_HVT U303 ( .A1(n327), .A2(n315), .Y(n568) );
  MUX21X1_HVT U304 ( .A1(n605), .A2(n217), .S0(n325), .Y(n508) );
  MUX21X1_HVT U305 ( .A1(n462), .A2(n463), .S0(n302), .Y(n460) );
  MUX21X1_HVT U306 ( .A1(n383), .A2(n392), .S0(n307), .Y(n463) );
  MUX21X1_HVT U307 ( .A1(n444), .A2(n443), .S0(n301), .Y(n442) );
  MUX21X1_HVT U308 ( .A1(n318), .A2(n381), .S0(n308), .Y(n444) );
  AND2X1_HVT U309 ( .A1(n217), .A2(n331), .Y(n295) );
  MUX21X1_HVT U310 ( .A1(n316), .A2(n391), .S0(n326), .Y(n576) );
  MUX21X1_HVT U311 ( .A1(n394), .A2(n381), .S0(n308), .Y(n546) );
  MUX21X1_HVT U312 ( .A1(n392), .A2(n395), .S0(n326), .Y(n449) );
  NAND2X0_HVT U313 ( .A1(n315), .A2(n314), .Y(n613) );
  NBUFFX2_HVT U314 ( .A(n396), .Y(n314) );
  MUX21X1_HVT U315 ( .A1(n366), .A2(n612), .S0(n299), .Y(n505) );
  MUX21X1_HVT U316 ( .A1(n458), .A2(n322), .S0(n296), .Y(n457) );
  MUX21X1_HVT U317 ( .A1(n597), .A2(n364), .S0(n299), .Y(n480) );
  NBUFFX2_HVT U318 ( .A(n614), .Y(n323) );
  NBUFFX2_HVT U319 ( .A(n605), .Y(n317) );
  MUX21X1_HVT U320 ( .A1(n395), .A2(n316), .S0(n325), .Y(n595) );
  MUX21X1_HVT U321 ( .A1(n564), .A2(n565), .S0(n306), .Y(n562) );
  MUX21X1_HVT U322 ( .A1(n316), .A2(n580), .S0(n305), .Y(n565) );
  XOR2X1_HVT U323 ( .A1(n326), .A2(n304), .Y(n572) );
  MUX21X1_HVT U324 ( .A1(n612), .A2(n330), .S0(n300), .Y(n487) );
  MUX21X1_HVT U325 ( .A1(n316), .A2(n392), .S0(n329), .Y(n404) );
  MUX21X1_HVT U326 ( .A1(n585), .A2(n408), .S0(n306), .Y(n402) );
  MUX21X1_HVT U327 ( .A1(n319), .A2(n316), .S0(n239), .Y(n606) );
  MUX21X1_HVT U328 ( .A1(n360), .A2(n585), .S0(n299), .Y(n483) );
  MUX21X1_HVT U329 ( .A1(n351), .A2(n331), .S0(n305), .Y(n550) );
  MUX21X1_HVT U330 ( .A1(n322), .A2(n524), .S0(n296), .Y(n523) );
  MUX21X1_HVT U331 ( .A1(n316), .A2(n313), .S0(n308), .Y(n524) );
  NBUFFX2_HVT U332 ( .A(n614), .Y(n324) );
  NBUFFX2_HVT U333 ( .A(n396), .Y(n313) );
  NBUFFX2_HVT U334 ( .A(n605), .Y(n318) );
  XNOR2X1_HVT U335 ( .A1(n337), .A2(n239), .Y(n296) );
  AND2X1_HVT U336 ( .A1(n309), .A2(n331), .Y(n297) );
  NBUFFX2_HVT U337 ( .A(in[5]), .Y(n334) );
  NBUFFX2_HVT U338 ( .A(in[5]), .Y(n333) );
  INVX0_HVT U339 ( .A(in[4]), .Y(n396) );
  MUX21X1_HVT U340 ( .A1(n522), .A2(n523), .S0(n302), .Y(n520) );
  MUX21X1_HVT U341 ( .A1(n562), .A2(n566), .S0(n301), .Y(n561) );
  MUX21X1_HVT U342 ( .A1(n556), .A2(n558), .S0(n300), .Y(n555) );
  MUX21X1_HVT U343 ( .A1(n391), .A2(n282), .S0(n329), .Y(n583) );
  MUX21X1_HVT U344 ( .A1(n282), .A2(n608), .S0(n238), .Y(n406) );
  MUX21X1_HVT U345 ( .A1(n282), .A2(n394), .S0(n329), .Y(n579) );
  MUX21X1_HVT U346 ( .A1(n282), .A2(n392), .S0(n325), .Y(n597) );
  NAND2X0_HVT U347 ( .A1(in[4]), .A2(n393), .Y(n605) );
  NAND2X0_HVT U348 ( .A1(n315), .A2(in[4]), .Y(n614) );
  MUX21X1_HVT U349 ( .A1(n282), .A2(n322), .S0(n238), .Y(n594) );
  MUX21X1_HVT U350 ( .A1(n324), .A2(n282), .S0(n328), .Y(n587) );
  MUX21X1_HVT U351 ( .A1(n316), .A2(n282), .S0(n302), .Y(n500) );
  MUX21X1_HVT U352 ( .A1(n282), .A2(n318), .S0(n329), .Y(n398) );
  MUX21X1_HVT U353 ( .A1(n282), .A2(n324), .S0(n238), .Y(n397) );
  MUX21X1_HVT U354 ( .A1(n309), .A2(n282), .S0(n327), .Y(n585) );
  NBUFFX2_HVT U355 ( .A(in[3]), .Y(n315) );
  NBUFFX2_HVT U356 ( .A(in[3]), .Y(n316) );
  INVX0_HVT U357 ( .A(n593), .Y(n339) );
  INVX0_HVT U358 ( .A(n591), .Y(n340) );
  INVX0_HVT U359 ( .A(n582), .Y(n341) );
  INVX0_HVT U360 ( .A(n580), .Y(n342) );
  INVX0_HVT U361 ( .A(n446), .Y(n343) );
  INVX0_HVT U362 ( .A(n409), .Y(n344) );
  INVX0_HVT U363 ( .A(n612), .Y(n345) );
  INVX0_HVT U364 ( .A(n599), .Y(n346) );
  INVX0_HVT U365 ( .A(n611), .Y(n347) );
  INVX0_HVT U366 ( .A(n607), .Y(n348) );
  INVX0_HVT U367 ( .A(n606), .Y(n349) );
  INVX0_HVT U368 ( .A(n604), .Y(n350) );
  INVX0_HVT U369 ( .A(n603), .Y(n351) );
  INVX0_HVT U370 ( .A(n600), .Y(n352) );
  INVX0_HVT U371 ( .A(n597), .Y(n353) );
  INVX0_HVT U372 ( .A(n596), .Y(n354) );
  INVX0_HVT U373 ( .A(n595), .Y(n355) );
  INVX0_HVT U374 ( .A(n592), .Y(n357) );
  INVX0_HVT U375 ( .A(n590), .Y(n358) );
  INVX0_HVT U376 ( .A(n589), .Y(n359) );
  INVX0_HVT U377 ( .A(n587), .Y(n360) );
  INVX0_HVT U378 ( .A(n585), .Y(n361) );
  INVX0_HVT U379 ( .A(n402), .Y(n362) );
  INVX0_HVT U380 ( .A(n584), .Y(n363) );
  INVX0_HVT U381 ( .A(n583), .Y(n364) );
  INVX0_HVT U382 ( .A(n581), .Y(n365) );
  INVX0_HVT U383 ( .A(n579), .Y(n366) );
  INVX0_HVT U384 ( .A(n578), .Y(n367) );
  INVX0_HVT U385 ( .A(n577), .Y(n368) );
  INVX0_HVT U386 ( .A(n576), .Y(n369) );
  INVX0_HVT U387 ( .A(n575), .Y(n370) );
  INVX0_HVT U388 ( .A(n574), .Y(n371) );
  INVX0_HVT U389 ( .A(n573), .Y(n372) );
  INVX0_HVT U390 ( .A(n542), .Y(n373) );
  INVX0_HVT U391 ( .A(n602), .Y(n374) );
  INVX0_HVT U392 ( .A(n408), .Y(n376) );
  INVX0_HVT U393 ( .A(n461), .Y(n378) );
  INVX0_HVT U394 ( .A(n407), .Y(n379) );
  INVX0_HVT U395 ( .A(n406), .Y(n380) );
  INVX0_HVT U396 ( .A(n405), .Y(n381) );
  INVX0_HVT U397 ( .A(n404), .Y(n382) );
  INVX0_HVT U398 ( .A(n403), .Y(n383) );
  INVX0_HVT U399 ( .A(n521), .Y(n384) );
  INVX0_HVT U400 ( .A(n511), .Y(n385) );
  INVX0_HVT U401 ( .A(n401), .Y(n386) );
  INVX0_HVT U402 ( .A(n400), .Y(n387) );
  INVX0_HVT U403 ( .A(n399), .Y(n388) );
  INVX0_HVT U404 ( .A(n397), .Y(n390) );
endmodule

