
module sbox_14 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n50, n210, n211, n212, n213, n216, n217, n218, n219, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588;

  NAND2X0_HVT U3 ( .A1(n299), .A2(n587), .Y(n586) );
  NAND2X0_HVT U4 ( .A1(n584), .A2(n586), .Y(n585) );
  NAND2X0_HVT U5 ( .A1(n298), .A2(n288), .Y(n583) );
  NAND2X0_HVT U13 ( .A1(n575), .A2(n297), .Y(n576) );
  NAND2X0_HVT U15 ( .A1(n586), .A2(n289), .Y(n573) );
  NAND2X0_HVT U21 ( .A1(n303), .A2(n584), .Y(n567) );
  NAND2X0_HVT U24 ( .A1(n292), .A2(n303), .Y(n565) );
  NAND2X0_HVT U33 ( .A1(n364), .A2(n303), .Y(n556) );
  NAND2X0_HVT U42 ( .A1(n301), .A2(n292), .Y(n547) );
  NAND2X0_HVT U53 ( .A1(n537), .A2(n546), .Y(n538) );
  NAND2X0_HVT U56 ( .A1(n584), .A2(n533), .Y(n534) );
  MUX41X1_HVT U57 ( .A1(n353), .A3(n569), .A2(n534), .A4(n578), .S0(n50), .S1(
        n306), .Y(n532) );
  NAND2X0_HVT U58 ( .A1(n297), .A2(n586), .Y(n531) );
  MUX41X1_HVT U59 ( .A1(n278), .A3(n531), .A2(n276), .A4(n327), .S0(n308), 
        .S1(n306), .Y(n530) );
  MUX41X1_HVT U61 ( .A1(n274), .A3(n326), .A2(n325), .A4(n289), .S0(n243), 
        .S1(n307), .Y(n528) );
  NAND2X0_HVT U62 ( .A1(n303), .A2(n587), .Y(n527) );
  MUX41X1_HVT U63 ( .A1(n527), .A3(n317), .A2(n347), .A4(n324), .S0(n50), .S1(
        n306), .Y(n526) );
  AO21X1_HVT U66 ( .A1(n322), .A2(n284), .A3(n346), .Y(n523) );
  MUX41X1_HVT U68 ( .A1(n320), .A3(n523), .A2(n522), .A4(n524), .S0(n238), 
        .S1(n217), .Y(n521) );
  MUX41X1_HVT U69 ( .A1(n521), .A3(n529), .A2(n525), .A4(n535), .S0(in[6]), 
        .S1(n260), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n294), .A2(n516), .Y(n517) );
  MUX41X1_HVT U74 ( .A1(n518), .A3(n563), .A2(n517), .A4(n565), .S0(n280), 
        .S1(n265), .Y(n515) );
  MUX41X1_HVT U75 ( .A1(n350), .A3(n355), .A2(n368), .A4(n331), .S0(n238), 
        .S1(n217), .Y(n514) );
  MUX41X1_HVT U77 ( .A1(n580), .A3(n357), .A2(n513), .A4(n356), .S0(n285), 
        .S1(n304), .Y(n512) );
  MUX41X1_HVT U78 ( .A1(n512), .A3(n515), .A2(n514), .A4(n519), .S0(n260), 
        .S1(in[5]), .Y(n511) );
  AND3X1_HVT U80 ( .A1(n587), .A2(n533), .A3(n508), .Y(n509) );
  MUX41X1_HVT U82 ( .A1(n544), .A3(n329), .A2(n312), .A4(n574), .S0(n246), 
        .S1(n50), .Y(n506) );
  AND2X1_HVT U83 ( .A1(n300), .A2(n266), .Y(n505) );
  MUX41X1_HVT U84 ( .A1(n330), .A3(n582), .A2(n572), .A4(n505), .S0(n246), 
        .S1(n48), .Y(n504) );
  NAND2X0_HVT U85 ( .A1(n303), .A2(n367), .Y(n503) );
  MUX41X1_HVT U86 ( .A1(n355), .A3(n503), .A2(n275), .A4(n271), .S0(n249), 
        .S1(n243), .Y(n502) );
  MUX41X1_HVT U87 ( .A1(n502), .A3(n506), .A2(n504), .A4(n507), .S0(n260), 
        .S1(n306), .Y(n501) );
  MUX41X1_HVT U90 ( .A1(n543), .A3(n547), .A2(n352), .A4(n500), .S0(n279), 
        .S1(n48), .Y(n499) );
  AO21X1_HVT U93 ( .A1(n287), .A2(n495), .A3(n351), .Y(n496) );
  MUX41X1_HVT U96 ( .A1(n312), .A3(n273), .A2(n354), .A4(n493), .S0(n249), 
        .S1(n308), .Y(n492) );
  MUX41X1_HVT U97 ( .A1(n350), .A3(n273), .A2(n301), .A4(n573), .S0(n249), 
        .S1(n243), .Y(n491) );
  NAND2X0_HVT U101 ( .A1(n486), .A2(n485), .Y(n487) );
  MUX41X1_HVT U103 ( .A1(n586), .A3(n321), .A2(n334), .A4(n554), .S0(n246), 
        .S1(n48), .Y(n483) );
  MUX41X1_HVT U105 ( .A1(n333), .A3(n542), .A2(n482), .A4(n349), .S0(n246), 
        .S1(n243), .Y(n481) );
  OA21X1_HVT U109 ( .A1(n340), .A2(n256), .A3(n327), .Y(n478) );
  NAND2X0_HVT U110 ( .A1(n587), .A2(n476), .Y(n477) );
  MUX41X1_HVT U114 ( .A1(n473), .A3(n479), .A2(n475), .A4(n478), .S0(n284), 
        .S1(n48), .Y(n472) );
  AND2X1_HVT U115 ( .A1(n211), .A2(n289), .Y(n471) );
  NAND2X0_HVT U123 ( .A1(n462), .A2(n461), .Y(n463) );
  MUX41X1_HVT U125 ( .A1(n567), .A3(n278), .A2(n320), .A4(n359), .S0(n279), 
        .S1(n48), .Y(n459) );
  AND3X1_HVT U128 ( .A1(n246), .A2(n303), .A3(n266), .Y(n456) );
  MUX41X1_HVT U131 ( .A1(n454), .A3(n456), .A2(n455), .A4(n457), .S0(n284), 
        .S1(n308), .Y(n453) );
  MUX41X1_HVT U135 ( .A1(n360), .A3(n365), .A2(n583), .A4(n562), .S0(n280), 
        .S1(n48), .Y(n450) );
  MUX41X1_HVT U136 ( .A1(n271), .A3(n556), .A2(n361), .A4(n553), .S0(n279), 
        .S1(n308), .Y(n449) );
  MUX41X1_HVT U139 ( .A1(n447), .A3(n450), .A2(n449), .A4(n451), .S0(n260), 
        .S1(n307), .Y(n446) );
  AND2X1_HVT U140 ( .A1(n293), .A2(n302), .Y(n445) );
  MUX41X1_HVT U141 ( .A1(n564), .A3(n341), .A2(n445), .A4(n338), .S0(n280), 
        .S1(n50), .Y(n444) );
  MUX41X1_HVT U142 ( .A1(n330), .A3(n289), .A2(n348), .A4(n293), .S0(n279), 
        .S1(n308), .Y(n443) );
  NAND2X0_HVT U146 ( .A1(n300), .A2(n297), .Y(n516) );
  MUX41X1_HVT U147 ( .A1(n361), .A3(n516), .A2(n350), .A4(n543), .S0(n280), 
        .S1(n308), .Y(n439) );
  MUX41X1_HVT U148 ( .A1(n439), .A3(n443), .A2(n440), .A4(n444), .S0(n260), 
        .S1(n306), .Y(n438) );
  OA21X1_HVT U151 ( .A1(n549), .A2(n239), .A3(n435), .Y(n436) );
  MUX41X1_HVT U153 ( .A1(n477), .A3(n274), .A2(n296), .A4(n245), .S0(n279), 
        .S1(n243), .Y(n433) );
  AND2X1_HVT U154 ( .A1(n287), .A2(n292), .Y(n432) );
  NAND2X0_HVT U158 ( .A1(n298), .A2(n367), .Y(n428) );
  MUX41X1_HVT U159 ( .A1(n576), .A3(n289), .A2(n428), .A4(n319), .S0(n304), 
        .S1(n50), .Y(n427) );
  MUX41X1_HVT U160 ( .A1(n427), .A3(n433), .A2(n429), .A4(n434), .S0(n244), 
        .S1(n283), .Y(n426) );
  AND2X1_HVT U162 ( .A1(n582), .A2(n516), .Y(n424) );
  NAND2X0_HVT U166 ( .A1(n297), .A2(n533), .Y(n420) );
  NAND2X0_HVT U167 ( .A1(n368), .A2(n303), .Y(n419) );
  MUX41X1_HVT U168 ( .A1(n353), .A3(n293), .A2(n419), .A4(n420), .S0(n304), 
        .S1(n265), .Y(n418) );
  MUX41X1_HVT U172 ( .A1(n415), .A3(n421), .A2(n418), .A4(n423), .S0(n244), 
        .S1(in[5]), .Y(n414) );
  MUX21X2_HVT U173 ( .A1(n414), .A2(n426), .S0(in[6]), .Y(out[5]) );
  NAND2X0_HVT U174 ( .A1(n301), .A2(n582), .Y(n575) );
  NAND2X0_HVT U177 ( .A1(n210), .A2(n291), .Y(n411) );
  MUX41X1_HVT U178 ( .A1(n571), .A3(n411), .A2(n362), .A4(n551), .S0(n280), 
        .S1(n265), .Y(n410) );
  MUX41X1_HVT U179 ( .A1(n561), .A3(n363), .A2(n315), .A4(n362), .S0(n304), 
        .S1(n265), .Y(n409) );
  MUX41X1_HVT U180 ( .A1(n318), .A3(n580), .A2(n576), .A4(n270), .S0(n285), 
        .S1(n304), .Y(n408) );
  MUX41X1_HVT U181 ( .A1(n408), .A3(n410), .A2(n409), .A4(n412), .S0(n260), 
        .S1(n283), .Y(n407) );
  OA21X1_HVT U184 ( .A1(n555), .A2(n239), .A3(n330), .Y(n404) );
  MUX41X1_HVT U186 ( .A1(n273), .A3(n550), .A2(n516), .A4(n543), .S0(n304), 
        .S1(n265), .Y(n402) );
  MUX41X1_HVT U189 ( .A1(n400), .A3(n575), .A2(n401), .A4(n349), .S0(n285), 
        .S1(n304), .Y(n399) );
  MUX41X1_HVT U190 ( .A1(n399), .A3(n402), .A2(n403), .A4(n406), .S0(n283), 
        .S1(n260), .Y(n398) );
  MUX41X1_HVT U193 ( .A1(n547), .A3(n554), .A2(n541), .A4(n397), .S0(n304), 
        .S1(n265), .Y(n396) );
  AO21X1_HVT U197 ( .A1(n275), .A2(n286), .A3(n351), .Y(n392) );
  OA21X1_HVT U201 ( .A1(n581), .A2(n242), .A3(n341), .Y(n388) );
  MUX41X1_HVT U204 ( .A1(n534), .A3(n576), .A2(n339), .A4(n566), .S0(n304), 
        .S1(n265), .Y(n385) );
  MUX41X1_HVT U205 ( .A1(n266), .A3(n586), .A2(n363), .A4(n337), .S0(n304), 
        .S1(n265), .Y(n384) );
  MUX41X1_HVT U206 ( .A1(n384), .A3(n386), .A2(n385), .A4(n387), .S0(n244), 
        .S1(n283), .Y(n383) );
  NAND2X0_HVT U208 ( .A1(n298), .A2(n584), .Y(n476) );
  NAND2X0_HVT U212 ( .A1(n210), .A2(n294), .Y(n533) );
  NAND2X0_HVT U214 ( .A1(n582), .A2(n303), .Y(n382) );
  NAND2X0_HVT U215 ( .A1(n476), .A2(n294), .Y(n381) );
  NAND2X0_HVT U218 ( .A1(n365), .A2(n211), .Y(n435) );
  NAND2X0_HVT U220 ( .A1(n286), .A2(n382), .Y(n508) );
  XOR2X2_HVT U1 ( .A1(n242), .A2(n562), .Y(n545) );
  XNOR2X1_HVT U2 ( .A1(n369), .A2(in[3]), .Y(n23) );
  IBUFFX16_HVT U6 ( .A(n23), .Y(n582) );
  AO21X2_HVT U7 ( .A1(n282), .A2(n293), .A3(n582), .Y(n468) );
  MUX21X2_HVT U8 ( .A1(n289), .A2(n364), .S0(n235), .Y(n493) );
  IBUFFX2_HVT U9 ( .A(n310), .Y(n48) );
  IBUFFX2_HVT U10 ( .A(n310), .Y(n50) );
  INVX0_HVT U11 ( .A(n310), .Y(n309) );
  XNOR2X2_HVT U12 ( .A1(n242), .A2(n299), .Y(n277) );
  MUX21X1_HVT U14 ( .A1(n496), .A2(n497), .S0(n282), .Y(n494) );
  NAND2X2_HVT U16 ( .A1(in[3]), .A2(n369), .Y(n587) );
  INVX2_HVT U17 ( .A(in[4]), .Y(n369) );
  IBUFFX2_HVT U18 ( .A(n302), .Y(n210) );
  IBUFFX2_HVT U19 ( .A(n302), .Y(n211) );
  NOR2X1_HVT U20 ( .A1(n266), .A2(n300), .Y(n245) );
  INVX1_HVT U22 ( .A(n302), .Y(n299) );
  MUX21X1_HVT U23 ( .A1(n388), .A2(n389), .S0(n281), .Y(n387) );
  MUX21X2_HVT U25 ( .A1(n404), .A2(n405), .S0(n212), .Y(n403) );
  IBUFFX16_HVT U26 ( .A(n256), .Y(n212) );
  NAND2X0_HVT U27 ( .A1(n501), .A2(n231), .Y(n232) );
  INVX2_HVT U28 ( .A(in[7]), .Y(n310) );
  INVX2_HVT U29 ( .A(n310), .Y(n308) );
  INVX1_HVT U30 ( .A(n310), .Y(n243) );
  MUX41X1_HVT U31 ( .A1(n458), .A3(n472), .A2(n453), .A4(n466), .S0(n213), 
        .S1(n216), .Y(out[3]) );
  IBUFFX16_HVT U32 ( .A(n268), .Y(n213) );
  IBUFFX16_HVT U34 ( .A(n244), .Y(n216) );
  INVX0_HVT U35 ( .A(n239), .Y(n217) );
  MUX21X1_HVT U36 ( .A1(n354), .A2(n582), .S0(n263), .Y(n218) );
  MUX21X1_HVT U37 ( .A1(n552), .A2(n588), .S0(n263), .Y(n219) );
  MUX21X1_HVT U38 ( .A1(n218), .A2(n219), .S0(n265), .Y(n394) );
  INVX2_HVT U39 ( .A(in[2]), .Y(n263) );
  NBUFFX2_HVT U40 ( .A(in[7]), .Y(n265) );
  IBUFFX2_HVT U41 ( .A(n263), .Y(n304) );
  NAND2X0_HVT U43 ( .A1(n511), .A2(in[6]), .Y(n233) );
  NAND2X0_HVT U44 ( .A1(n232), .A2(n233), .Y(out[1]) );
  IBUFFX2_HVT U45 ( .A(in[6]), .Y(n231) );
  MUX41X1_HVT U46 ( .A1(n396), .A3(n394), .A2(n395), .A4(n391), .S0(n257), 
        .S1(n234), .Y(n390) );
  IBUFFX16_HVT U47 ( .A(in[5]), .Y(n234) );
  INVX2_HVT U48 ( .A(n257), .Y(n260) );
  NBUFFX2_HVT U49 ( .A(n299), .Y(n235) );
  NBUFFX2_HVT U50 ( .A(n299), .Y(n236) );
  NBUFFX2_HVT U51 ( .A(n299), .Y(n237) );
  NAND2X0_HVT U52 ( .A1(n254), .A2(n255), .Y(out[6]) );
  INVX0_HVT U54 ( .A(n240), .Y(n430) );
  INVX0_HVT U55 ( .A(n357), .Y(n241) );
  MUX21X1_HVT U60 ( .A1(n558), .A2(n477), .S0(n279), .Y(n475) );
  MUX21X1_HVT U64 ( .A1(n587), .A2(n474), .S0(n269), .Y(n473) );
  INVX1_HVT U65 ( .A(n245), .Y(n554) );
  INVX1_HVT U67 ( .A(n282), .Y(n261) );
  INVX1_HVT U70 ( .A(n285), .Y(n242) );
  INVX0_HVT U71 ( .A(n50), .Y(n239) );
  INVX1_HVT U72 ( .A(in[0]), .Y(n257) );
  INVX1_HVT U76 ( .A(n257), .Y(n244) );
  INVX1_HVT U79 ( .A(n281), .Y(n256) );
  INVX1_HVT U81 ( .A(n261), .Y(n246) );
  INVX1_HVT U88 ( .A(n263), .Y(n238) );
  INVX0_HVT U89 ( .A(n306), .Y(n264) );
  INVX0_HVT U91 ( .A(n558), .Y(n337) );
  MUX21X1_HVT U92 ( .A1(n467), .A2(n470), .S0(n284), .Y(n466) );
  MUX21X2_HVT U94 ( .A1(n468), .A2(n469), .S0(n286), .Y(n467) );
  MUX41X1_HVT U95 ( .A1(n291), .A3(n413), .A2(n358), .A4(n575), .S0(n50), .S1(
        n238), .Y(n412) );
  MUX21X2_HVT U98 ( .A1(n356), .A2(n365), .S0(n286), .Y(n437) );
  MUX41X1_HVT U99 ( .A1(n311), .A3(n352), .A2(n329), .A4(n328), .S0(n239), 
        .S1(n306), .Y(n540) );
  INVX1_HVT U100 ( .A(n376), .Y(n356) );
  INVX1_HVT U102 ( .A(n299), .Y(n303) );
  MUX21X1_HVT U104 ( .A1(n241), .A2(n341), .S0(n242), .Y(n240) );
  MUX21X2_HVT U106 ( .A1(n438), .A2(n446), .S0(in[6]), .Y(out[4]) );
  MUX21X2_HVT U107 ( .A1(n437), .A2(n436), .S0(n256), .Y(n434) );
  OA21X1_HVT U108 ( .A1(n276), .A2(n242), .A3(n558), .Y(n416) );
  MUX41X1_HVT U111 ( .A1(n558), .A3(n331), .A2(n471), .A4(n576), .S0(n263), 
        .S1(n239), .Y(n470) );
  OA21X1_HVT U112 ( .A1(n314), .A2(n239), .A3(n558), .Y(n441) );
  NAND2X0_HVT U113 ( .A1(n431), .A2(n246), .Y(n247) );
  NAND2X0_HVT U116 ( .A1(n430), .A2(n261), .Y(n248) );
  NAND2X0_HVT U117 ( .A1(n247), .A2(n248), .Y(n429) );
  INVX1_HVT U118 ( .A(n551), .Y(n341) );
  MUX41X1_HVT U119 ( .A1(n488), .A3(n484), .A2(n483), .A4(n481), .S0(n264), 
        .S1(n257), .Y(n480) );
  NAND2X0_HVT U120 ( .A1(n574), .A2(n249), .Y(n250) );
  NAND2X0_HVT U121 ( .A1(n337), .A2(n261), .Y(n251) );
  NAND2X0_HVT U122 ( .A1(n250), .A2(n251), .Y(n489) );
  INVX1_HVT U124 ( .A(n261), .Y(n249) );
  MUX21X2_HVT U126 ( .A1(n367), .A2(n354), .S0(n287), .Y(n520) );
  MUX21X2_HVT U127 ( .A1(n538), .A2(n539), .S0(n285), .Y(n536) );
  NAND2X1_HVT U129 ( .A1(n463), .A2(n287), .Y(n252) );
  NAND2X0_HVT U130 ( .A1(n464), .A2(n242), .Y(n253) );
  NAND2X0_HVT U132 ( .A1(n252), .A2(n253), .Y(n460) );
  MUX21X2_HVT U133 ( .A1(n460), .A2(n459), .S0(n264), .Y(n458) );
  MUX21X1_HVT U134 ( .A1(n262), .A2(n586), .S0(n280), .Y(n479) );
  INVX1_HVT U137 ( .A(n262), .Y(n553) );
  NAND2X0_HVT U138 ( .A1(n398), .A2(n268), .Y(n254) );
  NAND2X0_HVT U143 ( .A1(n407), .A2(in[6]), .Y(n255) );
  INVX1_HVT U144 ( .A(n557), .Y(n338) );
  MUX21X2_HVT U145 ( .A1(n545), .A2(n520), .S0(n281), .Y(n519) );
  INVX1_HVT U149 ( .A(n378), .Y(n354) );
  NAND2X0_HVT U150 ( .A1(n383), .A2(n268), .Y(n258) );
  NAND2X0_HVT U152 ( .A1(n390), .A2(in[6]), .Y(n259) );
  NAND2X0_HVT U155 ( .A1(n258), .A2(n259), .Y(out[7]) );
  IBUFFX2_HVT U156 ( .A(n549), .Y(n343) );
  MUX21X1_HVT U157 ( .A1(n369), .A2(n588), .S0(n236), .Y(n262) );
  MUX41X1_HVT U161 ( .A1(n343), .A3(n553), .A2(n557), .A4(n577), .S0(n263), 
        .S1(n265), .Y(n386) );
  MUX21X2_HVT U163 ( .A1(n442), .A2(n441), .S0(n249), .Y(n440) );
  MUX21X2_HVT U164 ( .A1(n392), .A2(n393), .S0(n256), .Y(n391) );
  MUX21X2_HVT U165 ( .A1(n292), .A2(n554), .S0(n284), .Y(n539) );
  MUX21X2_HVT U169 ( .A1(n536), .A2(n540), .S0(n281), .Y(n535) );
  MUX41X1_HVT U170 ( .A1(n425), .A3(n272), .A2(n424), .A4(n326), .S0(n263), 
        .S1(n310), .Y(n423) );
  MUX21X2_HVT U171 ( .A1(n345), .A2(n362), .S0(n286), .Y(n393) );
  MUX21X2_HVT U175 ( .A1(n313), .A2(n465), .S0(n280), .Y(n464) );
  AO21X2_HVT U176 ( .A1(n302), .A2(n365), .A3(n242), .Y(n486) );
  IBUFFX2_HVT U182 ( .A(n302), .Y(n301) );
  MUX41X1_HVT U183 ( .A1(n492), .A3(n499), .A2(n491), .A4(n494), .S0(n260), 
        .S1(n264), .Y(n490) );
  INVX2_HVT U185 ( .A(in[1]), .Y(n302) );
  MUX21X2_HVT U187 ( .A1(n480), .A2(n490), .S0(in[6]), .Y(out[2]) );
  MUX41X1_HVT U188 ( .A1(n344), .A3(n332), .A2(n342), .A4(n295), .S0(n243), 
        .S1(n256), .Y(n406) );
  INVX0_HVT U191 ( .A(in[6]), .Y(n268) );
  IBUFFX2_HVT U192 ( .A(n369), .Y(n266) );
  MUX21X1_HVT U194 ( .A1(n288), .A2(n23), .S0(n302), .Y(n572) );
  IBUFFX2_HVT U195 ( .A(n302), .Y(n300) );
  MUX41X1_HVT U196 ( .A1(n293), .A3(n360), .A2(n562), .A4(n548), .S0(n242), 
        .S1(n261), .Y(n395) );
  MUX41X1_HVT U198 ( .A1(n422), .A3(n543), .A2(n335), .A4(n567), .S0(n310), 
        .S1(n256), .Y(n421) );
  XOR2X1_HVT U199 ( .A1(n261), .A2(n310), .Y(n267) );
  MUX21X2_HVT U200 ( .A1(n274), .A2(n489), .S0(n267), .Y(n488) );
  XNOR2X1_HVT U202 ( .A1(n302), .A2(n261), .Y(n269) );
  IBUFFX2_HVT U203 ( .A(n302), .Y(n298) );
  NBUFFX4_HVT U207 ( .A(n305), .Y(n279) );
  INVX0_HVT U209 ( .A(in[3]), .Y(n366) );
  INVX0_HVT U210 ( .A(n263), .Y(n305) );
  INVX1_HVT U211 ( .A(n295), .Y(n364) );
  MUX21X1_HVT U213 ( .A1(n272), .A2(n325), .S0(n279), .Y(n455) );
  NBUFFX2_HVT U216 ( .A(n23), .Y(n290) );
  NBUFFX2_HVT U217 ( .A(n23), .Y(n289) );
  AND2X1_HVT U219 ( .A1(n290), .A2(n533), .Y(n270) );
  NBUFFX2_HVT U221 ( .A(n584), .Y(n295) );
  INVX1_HVT U222 ( .A(n296), .Y(n368) );
  MUX21X1_HVT U223 ( .A1(n364), .A2(n367), .S0(n284), .Y(n537) );
  MUX21X1_HVT U224 ( .A1(n321), .A2(n365), .S0(n284), .Y(n522) );
  AND2X1_HVT U225 ( .A1(n587), .A2(n516), .Y(n271) );
  MUX21X1_HVT U226 ( .A1(n290), .A2(n367), .S0(n299), .Y(n581) );
  MUX21X1_HVT U227 ( .A1(n587), .A2(n289), .S0(n235), .Y(n548) );
  MUX21X1_HVT U228 ( .A1(n289), .A2(n291), .S0(n235), .Y(n485) );
  MUX21X1_HVT U229 ( .A1(n448), .A2(n585), .S0(n282), .Y(n447) );
  MUX21X1_HVT U230 ( .A1(n566), .A2(n342), .S0(n286), .Y(n448) );
  MUX21X1_HVT U231 ( .A1(n364), .A2(n368), .S0(n236), .Y(n413) );
  MUX21X1_HVT U232 ( .A1(n367), .A2(n23), .S0(n298), .Y(n425) );
  MUX21X1_HVT U233 ( .A1(n584), .A2(n582), .S0(n237), .Y(n552) );
  MUX21X1_HVT U234 ( .A1(n582), .A2(n365), .S0(n237), .Y(n373) );
  MUX21X1_HVT U235 ( .A1(n582), .A2(n368), .S0(n301), .Y(n564) );
  MUX21X1_HVT U236 ( .A1(n584), .A2(n294), .S0(n235), .Y(n500) );
  MUX21X1_HVT U237 ( .A1(n582), .A2(n291), .S0(n237), .Y(n513) );
  XOR2X1_HVT U238 ( .A1(n582), .A2(n210), .Y(n543) );
  MUX21X1_HVT U239 ( .A1(n288), .A2(n582), .S0(n211), .Y(n376) );
  MUX21X1_HVT U240 ( .A1(n368), .A2(n367), .S0(n211), .Y(n562) );
  MUX21X1_HVT U241 ( .A1(n367), .A2(n364), .S0(n237), .Y(n551) );
  MUX21X1_HVT U242 ( .A1(n367), .A2(n288), .S0(n235), .Y(n555) );
  MUX21X1_HVT U243 ( .A1(n288), .A2(n368), .S0(n236), .Y(n549) );
  MUX21X1_HVT U244 ( .A1(n291), .A2(n364), .S0(n298), .Y(n560) );
  MUX21X1_HVT U245 ( .A1(n336), .A2(n452), .S0(n281), .Y(n451) );
  MUX21X1_HVT U246 ( .A1(n359), .A2(n294), .S0(n286), .Y(n452) );
  MUX21X1_HVT U247 ( .A1(n245), .A2(n339), .S0(n279), .Y(n469) );
  NAND2X0_HVT U248 ( .A1(n369), .A2(n366), .Y(n584) );
  MUX21X1_HVT U249 ( .A1(n364), .A2(n291), .S0(n211), .Y(n374) );
  NBUFFX2_HVT U250 ( .A(n587), .Y(n296) );
  INVX1_HVT U251 ( .A(n588), .Y(n367) );
  MUX21X1_HVT U252 ( .A1(n587), .A2(n294), .S0(n298), .Y(n574) );
  MUX21X1_HVT U253 ( .A1(n295), .A2(n297), .S0(n300), .Y(n495) );
  MUX21X1_HVT U254 ( .A1(n291), .A2(n288), .S0(n237), .Y(n465) );
  MUX21X1_HVT U255 ( .A1(n288), .A2(n297), .S0(n300), .Y(n400) );
  MUX21X1_HVT U256 ( .A1(n588), .A2(n587), .S0(n236), .Y(n401) );
  MUX21X1_HVT U257 ( .A1(n365), .A2(n364), .S0(n301), .Y(n570) );
  INVX1_HVT U258 ( .A(n293), .Y(n365) );
  MUX21X1_HVT U259 ( .A1(n288), .A2(n367), .S0(n298), .Y(n578) );
  XOR2X1_HVT U260 ( .A1(n298), .A2(n365), .Y(n544) );
  MUX21X1_HVT U261 ( .A1(n288), .A2(n291), .S0(n300), .Y(n397) );
  XOR2X1_HVT U262 ( .A1(n296), .A2(n300), .Y(n541) );
  MUX21X1_HVT U263 ( .A1(n296), .A2(n291), .S0(n236), .Y(n380) );
  XNOR2X1_HVT U264 ( .A1(n295), .A2(n211), .Y(n272) );
  AND2X1_HVT U265 ( .A1(n211), .A2(n368), .Y(n273) );
  MUX21X1_HVT U266 ( .A1(n588), .A2(n294), .S0(n235), .Y(n558) );
  MUX21X1_HVT U267 ( .A1(n584), .A2(n288), .S0(n211), .Y(n577) );
  MUX21X1_HVT U268 ( .A1(n296), .A2(n584), .S0(n301), .Y(n372) );
  AND2X1_HVT U269 ( .A1(n297), .A2(n476), .Y(n274) );
  XNOR2X1_HVT U270 ( .A1(n588), .A2(n211), .Y(n275) );
  MUX21X1_HVT U271 ( .A1(n294), .A2(n288), .S0(n301), .Y(n378) );
  MUX21X1_HVT U272 ( .A1(n294), .A2(n291), .S0(n236), .Y(n518) );
  MUX21X1_HVT U273 ( .A1(n579), .A2(n297), .S0(n281), .Y(n462) );
  XOR2X1_HVT U274 ( .A1(n291), .A2(n298), .Y(n563) );
  NBUFFX2_HVT U275 ( .A(n309), .Y(n287) );
  NBUFFX2_HVT U276 ( .A(n309), .Y(n285) );
  NBUFFX2_HVT U277 ( .A(n243), .Y(n286) );
  NBUFFX2_HVT U278 ( .A(n366), .Y(n288) );
  NBUFFX2_HVT U279 ( .A(n307), .Y(n284) );
  NBUFFX2_HVT U280 ( .A(n305), .Y(n280) );
  NBUFFX2_HVT U281 ( .A(n307), .Y(n283) );
  NBUFFX2_HVT U282 ( .A(n238), .Y(n282) );
  NBUFFX2_HVT U283 ( .A(n238), .Y(n281) );
  MUX21X1_HVT U284 ( .A1(n572), .A2(n270), .S0(n285), .Y(n389) );
  MUX21X1_HVT U285 ( .A1(n290), .A2(n292), .S0(n301), .Y(n566) );
  MUX21X1_HVT U286 ( .A1(n487), .A2(n336), .S0(n249), .Y(n484) );
  MUX21X1_HVT U287 ( .A1(n503), .A2(n292), .S0(n286), .Y(n405) );
  MUX21X1_HVT U288 ( .A1(n526), .A2(n528), .S0(n281), .Y(n525) );
  XOR2X1_HVT U289 ( .A1(n301), .A2(n292), .Y(n542) );
  MUX21X1_HVT U290 ( .A1(n294), .A2(n290), .S0(n235), .Y(n482) );
  MUX21X1_HVT U291 ( .A1(n510), .A2(n509), .S0(n282), .Y(n507) );
  MUX21X1_HVT U292 ( .A1(n568), .A2(n294), .S0(n287), .Y(n510) );
  MUX21X1_HVT U293 ( .A1(n417), .A2(n416), .S0(n246), .Y(n415) );
  MUX21X1_HVT U294 ( .A1(n294), .A2(n354), .S0(n287), .Y(n417) );
  MUX21X1_HVT U295 ( .A1(n365), .A2(n368), .S0(n300), .Y(n422) );
  AND2X1_HVT U296 ( .A1(n290), .A2(n303), .Y(n276) );
  MUX21X1_HVT U297 ( .A1(n292), .A2(n364), .S0(n237), .Y(n550) );
  MUX21X1_HVT U298 ( .A1(n560), .A2(n316), .S0(n287), .Y(n442) );
  MUX21X1_HVT U299 ( .A1(n368), .A2(n292), .S0(n210), .Y(n569) );
  MUX21X1_HVT U300 ( .A1(n432), .A2(n587), .S0(n277), .Y(n431) );
  MUX21X1_HVT U301 ( .A1(n571), .A2(n338), .S0(n280), .Y(n454) );
  XOR2X1_HVT U302 ( .A1(n210), .A2(n283), .Y(n546) );
  MUX21X1_HVT U303 ( .A1(n586), .A2(n302), .S0(n281), .Y(n461) );
  NBUFFX2_HVT U304 ( .A(n579), .Y(n293) );
  MUX21X1_HVT U305 ( .A1(n292), .A2(n365), .S0(n210), .Y(n377) );
  MUX21X1_HVT U306 ( .A1(n559), .A2(n381), .S0(n285), .Y(n375) );
  MUX21X1_HVT U307 ( .A1(n584), .A2(n292), .S0(n211), .Y(n580) );
  MUX21X1_HVT U308 ( .A1(n323), .A2(n303), .S0(n284), .Y(n524) );
  NBUFFX2_HVT U309 ( .A(n579), .Y(n294) );
  MUX21X1_HVT U310 ( .A1(n333), .A2(n559), .S0(n280), .Y(n457) );
  MUX21X1_HVT U311 ( .A1(n587), .A2(n498), .S0(n277), .Y(n497) );
  MUX21X1_HVT U312 ( .A1(n292), .A2(n291), .S0(n287), .Y(n498) );
  NBUFFX2_HVT U313 ( .A(n588), .Y(n297) );
  NBUFFX2_HVT U314 ( .A(n369), .Y(n291) );
  AND2X1_HVT U315 ( .A1(n288), .A2(n303), .Y(n278) );
  NBUFFX2_HVT U316 ( .A(in[5]), .Y(n307) );
  NBUFFX2_HVT U317 ( .A(in[5]), .Y(n306) );
  MUX21X1_HVT U318 ( .A1(n530), .A2(n532), .S0(n281), .Y(n529) );
  MUX21X1_HVT U319 ( .A1(n364), .A2(n266), .S0(n237), .Y(n557) );
  NAND2X0_HVT U320 ( .A1(in[3]), .A2(in[4]), .Y(n588) );
  MUX21X1_HVT U321 ( .A1(n266), .A2(n582), .S0(n301), .Y(n379) );
  MUX21X1_HVT U322 ( .A1(n266), .A2(n365), .S0(n210), .Y(n571) );
  NAND2X0_HVT U323 ( .A1(in[4]), .A2(n366), .Y(n579) );
  MUX21X1_HVT U324 ( .A1(n266), .A2(n587), .S0(n300), .Y(n568) );
  MUX21X1_HVT U325 ( .A1(n297), .A2(n266), .S0(n210), .Y(n561) );
  MUX21X1_HVT U326 ( .A1(n292), .A2(n266), .S0(n279), .Y(n474) );
  MUX21X1_HVT U327 ( .A1(n266), .A2(n294), .S0(n210), .Y(n371) );
  MUX21X1_HVT U328 ( .A1(n266), .A2(n297), .S0(n236), .Y(n370) );
  MUX21X1_HVT U329 ( .A1(n288), .A2(n266), .S0(n298), .Y(n559) );
  NBUFFX2_HVT U330 ( .A(in[3]), .Y(n292) );
  INVX0_HVT U331 ( .A(n567), .Y(n311) );
  INVX0_HVT U332 ( .A(n565), .Y(n312) );
  INVX0_HVT U333 ( .A(n556), .Y(n313) );
  INVX0_HVT U334 ( .A(n419), .Y(n314) );
  INVX0_HVT U335 ( .A(n382), .Y(n315) );
  INVX0_HVT U336 ( .A(n586), .Y(n316) );
  INVX0_HVT U337 ( .A(n573), .Y(n317) );
  INVX0_HVT U338 ( .A(n585), .Y(n318) );
  INVX0_HVT U339 ( .A(n583), .Y(n319) );
  INVX0_HVT U340 ( .A(n581), .Y(n320) );
  INVX0_HVT U341 ( .A(n580), .Y(n321) );
  INVX0_HVT U342 ( .A(n578), .Y(n322) );
  INVX0_HVT U343 ( .A(n577), .Y(n323) );
  INVX0_HVT U344 ( .A(n574), .Y(n324) );
  INVX0_HVT U345 ( .A(n572), .Y(n325) );
  INVX0_HVT U346 ( .A(n571), .Y(n326) );
  INVX0_HVT U347 ( .A(n570), .Y(n327) );
  INVX0_HVT U348 ( .A(n569), .Y(n328) );
  INVX0_HVT U349 ( .A(n568), .Y(n329) );
  INVX0_HVT U350 ( .A(n566), .Y(n330) );
  INVX0_HVT U351 ( .A(n564), .Y(n331) );
  INVX0_HVT U352 ( .A(n563), .Y(n332) );
  INVX0_HVT U353 ( .A(n561), .Y(n333) );
  INVX0_HVT U354 ( .A(n560), .Y(n334) );
  INVX0_HVT U355 ( .A(n559), .Y(n335) );
  INVX0_HVT U356 ( .A(n375), .Y(n336) );
  INVX0_HVT U357 ( .A(n555), .Y(n339) );
  INVX0_HVT U358 ( .A(n552), .Y(n340) );
  INVX0_HVT U359 ( .A(n550), .Y(n342) );
  INVX0_HVT U360 ( .A(n548), .Y(n344) );
  INVX0_HVT U361 ( .A(n547), .Y(n345) );
  INVX0_HVT U362 ( .A(n516), .Y(n346) );
  INVX0_HVT U363 ( .A(n576), .Y(n347) );
  INVX0_HVT U364 ( .A(n476), .Y(n348) );
  INVX0_HVT U365 ( .A(n381), .Y(n349) );
  INVX0_HVT U366 ( .A(n533), .Y(n350) );
  INVX0_HVT U367 ( .A(n435), .Y(n351) );
  INVX0_HVT U368 ( .A(n380), .Y(n352) );
  INVX0_HVT U369 ( .A(n379), .Y(n353) );
  INVX0_HVT U370 ( .A(n377), .Y(n355) );
  INVX0_HVT U371 ( .A(n495), .Y(n357) );
  INVX0_HVT U372 ( .A(n485), .Y(n358) );
  INVX0_HVT U373 ( .A(n374), .Y(n359) );
  INVX0_HVT U374 ( .A(n373), .Y(n360) );
  INVX0_HVT U375 ( .A(n372), .Y(n361) );
  INVX0_HVT U376 ( .A(n371), .Y(n362) );
  INVX0_HVT U377 ( .A(n370), .Y(n363) );
endmodule

