
module inv_sbox_10 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n177, n196, n197, n198, n199, n200, n201, n202, n203, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609;

  NAND2X0_HVT U1 ( .A1(in[3]), .A2(n307), .Y(n609) );
  NAND2X0_HVT U3 ( .A1(in[3]), .A2(in[6]), .Y(n607) );
  NAND2X0_HVT U4 ( .A1(n328), .A2(n322), .Y(n606) );
  NAND2X0_HVT U5 ( .A1(n606), .A2(n318), .Y(n605) );
  NAND2X0_HVT U7 ( .A1(n326), .A2(n320), .Y(n602) );
  NAND2X0_HVT U8 ( .A1(n326), .A2(n318), .Y(n601) );
  NAND2X0_HVT U9 ( .A1(n275), .A2(n601), .Y(n600) );
  NAND2X0_HVT U10 ( .A1(n324), .A2(n598), .Y(n599) );
  NAND2X0_HVT U11 ( .A1(n330), .A2(n323), .Y(n597) );
  NAND2X0_HVT U12 ( .A1(n261), .A2(n281), .Y(n596) );
  NAND2X0_HVT U13 ( .A1(n320), .A2(n238), .Y(n595) );
  NAND2X0_HVT U15 ( .A1(n315), .A2(n326), .Y(n593) );
  NAND2X0_HVT U19 ( .A1(n274), .A2(n399), .Y(n588) );
  NAND2X0_HVT U32 ( .A1(n307), .A2(n330), .Y(n576) );
  NAND2X0_HVT U35 ( .A1(n601), .A2(n285), .Y(n573) );
  NAND2X0_HVT U38 ( .A1(n282), .A2(n330), .Y(n570) );
  NAND2X0_HVT U42 ( .A1(n603), .A2(n400), .Y(n566) );
  OA21X1_HVT U53 ( .A1(n231), .A2(n558), .A3(n367), .Y(n556) );
  NAND2X0_HVT U55 ( .A1(n320), .A2(n606), .Y(n554) );
  MUX41X1_HVT U56 ( .A1(n278), .A3(n314), .A2(n365), .A4(n554), .S0(n301), 
        .S1(n335), .Y(n553) );
  AO21X1_HVT U60 ( .A1(n548), .A2(n245), .A3(n587), .Y(n549) );
  MUX41X1_HVT U65 ( .A1(n357), .A3(n359), .A2(n358), .A4(n570), .S0(n301), 
        .S1(n335), .Y(n543) );
  NAND2X0_HVT U66 ( .A1(n274), .A2(n288), .Y(n542) );
  MUX41X1_HVT U67 ( .A1(n354), .A3(n381), .A2(n356), .A4(n542), .S0(n305), 
        .S1(n298), .Y(n541) );
  MUX41X1_HVT U71 ( .A1(n603), .A3(n277), .A2(n597), .A4(n350), .S0(n300), 
        .S1(n335), .Y(n538) );
  NAND2X0_HVT U72 ( .A1(n316), .A2(n602), .Y(n537) );
  MUX41X1_HVT U73 ( .A1(n581), .A3(n537), .A2(n382), .A4(n281), .S0(n245), 
        .S1(n297), .Y(n536) );
  MUX41X1_HVT U74 ( .A1(n599), .A3(n372), .A2(n371), .A4(n360), .S0(n301), 
        .S1(n304), .Y(n535) );
  MUX41X1_HVT U78 ( .A1(n532), .A3(n536), .A2(n535), .A4(n538), .S0(in[5]), 
        .S1(n310), .Y(n531) );
  MUX41X1_HVT U79 ( .A1(n368), .A3(n590), .A2(n370), .A4(n591), .S0(n301), 
        .S1(n335), .Y(n530) );
  MUX41X1_HVT U80 ( .A1(n384), .A3(n278), .A2(n600), .A4(n605), .S0(n300), 
        .S1(n335), .Y(n529) );
  NAND2X0_HVT U81 ( .A1(n321), .A2(n602), .Y(n528) );
  AND2X1_HVT U82 ( .A1(n603), .A2(n319), .Y(n527) );
  MUX41X1_HVT U83 ( .A1(n527), .A3(n369), .A2(n385), .A4(n528), .S0(n300), 
        .S1(n335), .Y(n526) );
  MUX41X1_HVT U84 ( .A1(n293), .A3(n368), .A2(n386), .A4(n583), .S0(n301), 
        .S1(n244), .Y(n525) );
  MUX41X1_HVT U85 ( .A1(n525), .A3(n529), .A2(n526), .A4(n530), .S0(in[5]), 
        .S1(n310), .Y(n524) );
  MUX41X1_HVT U87 ( .A1(n344), .A3(n293), .A2(n387), .A4(n365), .S0(n299), 
        .S1(n305), .Y(n523) );
  NAND2X0_HVT U89 ( .A1(n330), .A2(n397), .Y(n521) );
  MUX41X1_HVT U90 ( .A1(n277), .A3(n198), .A2(n561), .A4(n521), .S0(n300), 
        .S1(n245), .Y(n520) );
  MUX41X1_HVT U95 ( .A1(n516), .A3(n522), .A2(n520), .A4(n523), .S0(n313), 
        .S1(n310), .Y(n515) );
  MUX41X1_HVT U96 ( .A1(n381), .A3(n595), .A2(n366), .A4(n388), .S0(n301), 
        .S1(n250), .Y(n514) );
  MUX41X1_HVT U99 ( .A1(n576), .A3(n358), .A2(n560), .A4(n314), .S0(n305), 
        .S1(n298), .Y(n511) );
  NAND2X0_HVT U100 ( .A1(n330), .A2(n279), .Y(n510) );
  MUX41X1_HVT U101 ( .A1(n390), .A3(n596), .A2(n373), .A4(n510), .S0(n303), 
        .S1(n296), .Y(n509) );
  AND2X1_HVT U104 ( .A1(n198), .A2(n317), .Y(n507) );
  MUX41X1_HVT U105 ( .A1(n594), .A3(n391), .A2(n197), .A4(n507), .S0(n301), 
        .S1(n334), .Y(n506) );
  MUX41X1_HVT U107 ( .A1(n390), .A3(n319), .A2(n505), .A4(n347), .S0(n300), 
        .S1(n250), .Y(n504) );
  MUX41X1_HVT U108 ( .A1(n360), .A3(n314), .A2(n365), .A4(n323), .S0(n301), 
        .S1(n333), .Y(n503) );
  MUX41X1_HVT U109 ( .A1(n389), .A3(n341), .A2(n386), .A4(n379), .S0(n300), 
        .S1(n250), .Y(n502) );
  MUX41X1_HVT U110 ( .A1(n502), .A3(n504), .A2(n503), .A4(n506), .S0(n313), 
        .S1(n311), .Y(n501) );
  AO21X1_HVT U112 ( .A1(n376), .A2(n244), .A3(n584), .Y(n499) );
  NAND2X0_HVT U114 ( .A1(n276), .A2(n198), .Y(n497) );
  MUX41X1_HVT U115 ( .A1(n497), .A3(n597), .A2(n376), .A4(n319), .S0(n335), 
        .S1(n298), .Y(n496) );
  MUX41X1_HVT U116 ( .A1(n375), .A3(n368), .A2(n341), .A4(n593), .S0(n299), 
        .S1(n250), .Y(n495) );
  NAND2X0_HVT U118 ( .A1(n330), .A2(n273), .Y(n493) );
  MUX41X1_HVT U119 ( .A1(n392), .A3(n494), .A2(n571), .A4(n493), .S0(n299), 
        .S1(n334), .Y(n492) );
  MUX41X1_HVT U120 ( .A1(n492), .A3(n496), .A2(n495), .A4(n498), .S0(n313), 
        .S1(n310), .Y(n491) );
  MUX41X1_HVT U122 ( .A1(n380), .A3(n289), .A2(n562), .A4(n383), .S0(n299), 
        .S1(n334), .Y(n490) );
  MUX41X1_HVT U124 ( .A1(n292), .A3(n489), .A2(n585), .A4(n362), .S0(n305), 
        .S1(n299), .Y(n488) );
  AOI21X1_HVT U127 ( .A1(n296), .A2(n484), .A3(n348), .Y(n485) );
  NAND2X0_HVT U129 ( .A1(n302), .A2(n324), .Y(n482) );
  MUX41X1_HVT U130 ( .A1(n482), .A3(n483), .A2(n486), .A4(n485), .S0(n305), 
        .S1(n310), .Y(n481) );
  AND2X1_HVT U131 ( .A1(n288), .A2(n242), .Y(n480) );
  MUX41X1_HVT U132 ( .A1(n345), .A3(n480), .A2(n394), .A4(n354), .S0(n245), 
        .S1(n297), .Y(n479) );
  MUX41X1_HVT U133 ( .A1(n395), .A3(n347), .A2(n554), .A4(n346), .S0(n244), 
        .S1(n296), .Y(n478) );
  MUX41X1_HVT U136 ( .A1(n559), .A3(n510), .A2(n476), .A4(n352), .S0(n302), 
        .S1(n334), .Y(n475) );
  MUX41X1_HVT U137 ( .A1(n238), .A3(n579), .A2(n583), .A4(n388), .S0(n304), 
        .S1(n296), .Y(n474) );
  MUX41X1_HVT U139 ( .A1(n473), .A3(n477), .A2(n481), .A4(n487), .S0(n313), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n371), .A3(n290), .A2(n364), .A4(n597), .S0(n244), 
        .S1(n298), .Y(n472) );
  NAND2X0_HVT U141 ( .A1(n315), .A2(n330), .Y(n471) );
  MUX41X1_HVT U142 ( .A1(n471), .A3(n569), .A2(n393), .A4(n364), .S0(n235), 
        .S1(n333), .Y(n470) );
  MUX41X1_HVT U151 ( .A1(n385), .A3(n374), .A2(n361), .A4(n462), .S0(n304), 
        .S1(n296), .Y(n461) );
  MUX41X1_HVT U155 ( .A1(n364), .A3(n597), .A2(n589), .A4(n366), .S0(n271), 
        .S1(n333), .Y(n457) );
  MUX41X1_HVT U156 ( .A1(n457), .A3(n461), .A2(n458), .A4(n463), .S0(n313), 
        .S1(in[1]), .Y(n456) );
  NAND2X0_HVT U159 ( .A1(n453), .A2(n452), .Y(n454) );
  MUX41X1_HVT U162 ( .A1(n280), .A3(n359), .A2(n573), .A4(n450), .S0(n235), 
        .S1(n333), .Y(n449) );
  NAND2X0_HVT U163 ( .A1(n328), .A2(n397), .Y(n448) );
  MUX41X1_HVT U164 ( .A1(n600), .A3(n448), .A2(n571), .A4(n360), .S0(n299), 
        .S1(n333), .Y(n447) );
  NAND2X0_HVT U166 ( .A1(n598), .A2(n444), .Y(n445) );
  MUX41X1_HVT U172 ( .A1(n521), .A3(n439), .A2(n291), .A4(n586), .S0(n271), 
        .S1(n250), .Y(n438) );
  MUX41X1_HVT U173 ( .A1(n276), .A3(n277), .A2(n321), .A4(n572), .S0(n235), 
        .S1(n251), .Y(n437) );
  MUX41X1_HVT U174 ( .A1(n387), .A3(n554), .A2(n395), .A4(n285), .S0(n235), 
        .S1(n334), .Y(n436) );
  MUX41X1_HVT U175 ( .A1(n436), .A3(n437), .A2(n438), .A4(n440), .S0(n311), 
        .S1(n313), .Y(n435) );
  NAND2X0_HVT U177 ( .A1(n262), .A2(n273), .Y(n434) );
  AND2X1_HVT U179 ( .A1(n603), .A2(n317), .Y(n433) );
  MUX41X1_HVT U183 ( .A1(n377), .A3(n278), .A2(n360), .A4(n566), .S0(n304), 
        .S1(n297), .Y(n429) );
  AND2X1_HVT U185 ( .A1(n285), .A2(n242), .Y(n427) );
  NAND2X0_HVT U191 ( .A1(n231), .A2(n353), .Y(n421) );
  AND2X1_HVT U192 ( .A1(n372), .A2(n419), .Y(n420) );
  NAND2X0_HVT U194 ( .A1(n566), .A2(n419), .Y(n417) );
  MUX41X1_HVT U195 ( .A1(n418), .A3(n417), .A2(n420), .A4(n421), .S0(n300), 
        .S1(n311), .Y(n416) );
  NAND2X0_HVT U198 ( .A1(n327), .A2(n285), .Y(n598) );
  NAND2X0_HVT U200 ( .A1(n318), .A2(n330), .Y(n484) );
  NAND2X0_HVT U207 ( .A1(n330), .A2(n277), .Y(n548) );
  NBUFFX4_HVT U2 ( .A(n329), .Y(n233) );
  DELLN1X2_HVT U6 ( .A(n309), .Y(n177) );
  INVX0_HVT U14 ( .A(in[1]), .Y(n309) );
  MUX21X2_HVT U16 ( .A1(n565), .A2(n383), .S0(n305), .Y(n455) );
  INVX0_HVT U17 ( .A(n274), .Y(n330) );
  INVX0_HVT U18 ( .A(n274), .Y(n260) );
  INVX1_HVT U20 ( .A(n329), .Y(n274) );
  INVX0_HVT U21 ( .A(n528), .Y(n196) );
  INVX0_HVT U22 ( .A(n196), .Y(n197) );
  INVX1_HVT U23 ( .A(n348), .Y(n198) );
  MUX21X2_HVT U24 ( .A1(n348), .A2(n567), .S0(n245), .Y(n500) );
  MUX41X1_HVT U25 ( .A1(n416), .A3(n428), .A2(n422), .A4(n431), .S0(n199), 
        .S1(n200), .Y(out[7]) );
  IBUFFX16_HVT U26 ( .A(n272), .Y(n199) );
  IBUFFX16_HVT U27 ( .A(n312), .Y(n200) );
  INVX4_HVT U28 ( .A(n233), .Y(n327) );
  MUX21X2_HVT U29 ( .A1(n534), .A2(n533), .S0(n271), .Y(n532) );
  MUX41X1_HVT U30 ( .A1(n606), .A3(n347), .A2(n385), .A4(n344), .S0(n201), 
        .S1(n251), .Y(n430) );
  IBUFFX16_HVT U31 ( .A(n299), .Y(n201) );
  INVX0_HVT U33 ( .A(n398), .Y(n273) );
  MUX21X2_HVT U34 ( .A1(n499), .A2(n500), .S0(n271), .Y(n498) );
  INVX1_HVT U36 ( .A(n574), .Y(n372) );
  MUX21X2_HVT U37 ( .A1(n454), .A2(n455), .S0(n298), .Y(n451) );
  INVX2_HVT U39 ( .A(n233), .Y(n262) );
  MUX21X2_HVT U40 ( .A1(n293), .A2(n583), .S0(n202), .Y(n460) );
  IBUFFX16_HVT U41 ( .A(n244), .Y(n202) );
  OA21X2_HVT U43 ( .A1(n342), .A2(n231), .A3(n351), .Y(n459) );
  IBUFFX2_HVT U44 ( .A(n571), .Y(n374) );
  INVX0_HVT U45 ( .A(n583), .Y(n364) );
  NAND2X0_HVT U46 ( .A1(n360), .A2(n203), .Y(n218) );
  NAND2X0_HVT U47 ( .A1(n545), .A2(n295), .Y(n219) );
  NAND2X0_HVT U48 ( .A1(n218), .A2(n219), .Y(n544) );
  IBUFFX2_HVT U49 ( .A(n295), .Y(n203) );
  NAND2X0_HVT U50 ( .A1(n396), .A2(n220), .Y(n221) );
  NAND2X0_HVT U51 ( .A1(n400), .A2(n228), .Y(n222) );
  NAND2X0_HVT U52 ( .A1(n221), .A2(n222), .Y(n586) );
  INVX0_HVT U54 ( .A(n228), .Y(n220) );
  INVX1_HVT U57 ( .A(n587), .Y(n360) );
  MUX21X1_HVT U58 ( .A1(n606), .A2(n361), .S0(n227), .Y(n545) );
  INVX0_HVT U59 ( .A(n586), .Y(n361) );
  NAND2X0_HVT U61 ( .A1(n363), .A2(n223), .Y(n224) );
  NAND2X0_HVT U62 ( .A1(n552), .A2(n295), .Y(n225) );
  NAND2X0_HVT U63 ( .A1(n224), .A2(n225), .Y(n551) );
  INVX0_HVT U64 ( .A(n295), .Y(n223) );
  MUX21X1_HVT U68 ( .A1(n382), .A2(n567), .S0(n303), .Y(n424) );
  INVX1_HVT U69 ( .A(n229), .Y(n567) );
  INVX1_HVT U70 ( .A(n329), .Y(n325) );
  INVX0_HVT U75 ( .A(n592), .Y(n285) );
  IBUFFX16_HVT U76 ( .A(n309), .Y(n310) );
  MUX41X1_HVT U77 ( .A1(n423), .A3(n426), .A2(n424), .A4(n425), .S0(n311), 
        .S1(n226), .Y(n422) );
  IBUFFX16_HVT U86 ( .A(n297), .Y(n226) );
  INVX1_HVT U88 ( .A(n412), .Y(n384) );
  INVX2_HVT U91 ( .A(n309), .Y(n311) );
  MUX21X1_HVT U92 ( .A1(n306), .A2(n285), .S0(n261), .Y(n572) );
  AO21X1_HVT U93 ( .A1(n242), .A2(n276), .A3(n231), .Y(n452) );
  IBUFFX16_HVT U94 ( .A(n302), .Y(n227) );
  IBUFFX2_HVT U97 ( .A(n328), .Y(n228) );
  MUX21X2_HVT U98 ( .A1(n394), .A2(n345), .S0(n303), .Y(n465) );
  IBUFFX2_HVT U102 ( .A(n606), .Y(n344) );
  AO21X2_HVT U103 ( .A1(n316), .A2(n606), .A3(n231), .Y(n444) );
  AO21X2_HVT U106 ( .A1(n328), .A2(n279), .A3(n231), .Y(n419) );
  MUX21X1_HVT U111 ( .A1(n308), .A2(n319), .S0(n325), .Y(n229) );
  INVX0_HVT U113 ( .A(n308), .Y(n288) );
  INVX1_HVT U117 ( .A(n319), .Y(n399) );
  MUX21X1_HVT U121 ( .A1(n318), .A2(n275), .S0(n274), .Y(n280) );
  MUX21X2_HVT U123 ( .A1(n427), .A2(n384), .S0(n303), .Y(n426) );
  MUX21X2_HVT U125 ( .A1(n491), .A2(n501), .S0(in[7]), .Y(out[3]) );
  MUX21X2_HVT U126 ( .A1(n459), .A2(n460), .S0(n301), .Y(n458) );
  MUX21X2_HVT U128 ( .A1(n316), .A2(n308), .S0(n261), .Y(n583) );
  INVX2_HVT U134 ( .A(n233), .Y(n261) );
  IBUFFX2_HVT U135 ( .A(n338), .Y(n230) );
  INVX2_HVT U138 ( .A(n230), .Y(n231) );
  INVX0_HVT U143 ( .A(in[4]), .Y(n338) );
  INVX1_HVT U144 ( .A(n338), .Y(n336) );
  INVX0_HVT U145 ( .A(n337), .Y(n251) );
  INVX1_HVT U146 ( .A(n337), .Y(n333) );
  MUX21X2_HVT U147 ( .A1(n531), .A2(n524), .S0(n232), .Y(out[1]) );
  IBUFFX16_HVT U148 ( .A(in[7]), .Y(n232) );
  INVX1_HVT U149 ( .A(n304), .Y(n263) );
  INVX0_HVT U150 ( .A(n308), .Y(n249) );
  INVX1_HVT U152 ( .A(in[0]), .Y(n329) );
  INVX0_HVT U153 ( .A(n398), .Y(n234) );
  OA21X1_HVT U154 ( .A1(n368), .A2(n231), .A3(n548), .Y(n423) );
  NAND2X0_HVT U157 ( .A1(n607), .A2(n257), .Y(n258) );
  MUX21X1_HVT U158 ( .A1(n306), .A2(n397), .S0(n262), .Y(n462) );
  INVX1_HVT U160 ( .A(n603), .Y(n346) );
  INVX1_HVT U161 ( .A(n337), .Y(n334) );
  INVX1_HVT U165 ( .A(n336), .Y(n337) );
  NAND2X0_HVT U167 ( .A1(n328), .A2(n609), .Y(n603) );
  INVX0_HVT U168 ( .A(n563), .Y(n378) );
  NAND2X0_HVT U169 ( .A1(n518), .A2(n235), .Y(n236) );
  INVX1_HVT U170 ( .A(n312), .Y(n313) );
  INVX1_HVT U171 ( .A(in[5]), .Y(n312) );
  INVX0_HVT U176 ( .A(n296), .Y(n243) );
  INVX1_HVT U178 ( .A(n302), .Y(n241) );
  INVX1_HVT U180 ( .A(n266), .Y(n271) );
  INVX1_HVT U181 ( .A(n241), .Y(n235) );
  INVX0_HVT U182 ( .A(n272), .Y(n254) );
  OR2X1_HVT U184 ( .A1(n308), .A2(n234), .Y(n604) );
  NAND2X0_HVT U186 ( .A1(n517), .A2(n241), .Y(n237) );
  NAND2X0_HVT U187 ( .A1(n236), .A2(n237), .Y(n516) );
  INVX0_HVT U188 ( .A(n349), .Y(n238) );
  MUX21X1_HVT U189 ( .A1(n350), .A2(n315), .S0(n305), .Y(n517) );
  INVX0_HVT U190 ( .A(n601), .Y(n349) );
  INVX1_HVT U193 ( .A(n579), .Y(n368) );
  INVX1_HVT U196 ( .A(n317), .Y(n397) );
  MUX21X1_HVT U197 ( .A1(n465), .A2(n464), .S0(n302), .Y(n463) );
  AO21X1_HVT U199 ( .A1(n304), .A2(n349), .A3(n279), .Y(n464) );
  NAND2X0_HVT U201 ( .A1(n429), .A2(n177), .Y(n239) );
  NAND2X0_HVT U202 ( .A1(n430), .A2(n311), .Y(n240) );
  NAND2X0_HVT U203 ( .A1(n239), .A2(n240), .Y(n428) );
  MUX21X1_HVT U204 ( .A1(n308), .A2(n317), .S0(n262), .Y(n278) );
  INVX1_HVT U205 ( .A(n257), .Y(n242) );
  INVX1_HVT U206 ( .A(n260), .Y(n257) );
  MUX21X1_HVT U208 ( .A1(n605), .A2(n364), .S0(n266), .Y(n552) );
  MUX41X1_HVT U209 ( .A1(n391), .A3(n577), .A2(n197), .A4(n468), .S0(n243), 
        .S1(n251), .Y(n467) );
  NBUFFX2_HVT U210 ( .A(n336), .Y(n244) );
  NBUFFX2_HVT U211 ( .A(n336), .Y(n245) );
  INVX1_HVT U212 ( .A(n269), .Y(n557) );
  MUX41X1_HVT U213 ( .A1(n553), .A3(n547), .A2(n555), .A4(n551), .S0(n312), 
        .S1(n310), .Y(n546) );
  NBUFFX2_HVT U214 ( .A(n336), .Y(n305) );
  NBUFFX2_HVT U215 ( .A(n336), .Y(n303) );
  NAND2X0_HVT U216 ( .A1(n432), .A2(n177), .Y(n246) );
  NAND2X0_HVT U217 ( .A1(n286), .A2(n310), .Y(n247) );
  NAND2X0_HVT U218 ( .A1(n247), .A2(n246), .Y(n431) );
  NBUFFX2_HVT U219 ( .A(n336), .Y(n304) );
  INVX0_HVT U220 ( .A(n248), .Y(n519) );
  MUX21X1_HVT U221 ( .A1(n285), .A2(n249), .S0(n245), .Y(n248) );
  INVX1_HVT U222 ( .A(n337), .Y(n250) );
  MUX41X1_HVT U223 ( .A1(n339), .A3(n576), .A2(n563), .A4(n433), .S0(n241), 
        .S1(n251), .Y(n432) );
  OA21X2_HVT U224 ( .A1(n343), .A2(n231), .A3(n587), .Y(n533) );
  MUX21X1_HVT U225 ( .A1(n556), .A2(n557), .S0(n241), .Y(n555) );
  NAND2X0_HVT U226 ( .A1(n539), .A2(n272), .Y(n252) );
  NAND2X0_HVT U227 ( .A1(n546), .A2(n254), .Y(n253) );
  NAND2X0_HVT U228 ( .A1(n252), .A2(n253), .Y(out[0]) );
  MUX41X1_HVT U229 ( .A1(n441), .A3(n291), .A2(n292), .A4(n294), .S0(n263), 
        .S1(n266), .Y(n440) );
  NAND2X0_HVT U230 ( .A1(n442), .A2(n254), .Y(n255) );
  NAND2X0_HVT U231 ( .A1(n435), .A2(n272), .Y(n256) );
  NAND2X0_HVT U232 ( .A1(n255), .A2(n256), .Y(out[6]) );
  INVX0_HVT U233 ( .A(n331), .Y(n266) );
  NAND2X0_HVT U234 ( .A1(n519), .A2(n260), .Y(n259) );
  NAND2X0_HVT U235 ( .A1(n258), .A2(n259), .Y(n518) );
  MUX21X2_HVT U236 ( .A1(n508), .A2(n515), .S0(n254), .Y(out[2]) );
  INVX1_HVT U237 ( .A(n303), .Y(n270) );
  MUX41X1_HVT U238 ( .A1(n562), .A3(n578), .A2(n341), .A4(n356), .S0(n243), 
        .S1(n337), .Y(n522) );
  MUX21X2_HVT U239 ( .A1(n549), .A2(n550), .S0(n241), .Y(n547) );
  INVX1_HVT U240 ( .A(n329), .Y(n328) );
  NAND2X0_HVT U241 ( .A1(n293), .A2(n263), .Y(n264) );
  NAND2X0_HVT U242 ( .A1(n560), .A2(n245), .Y(n265) );
  NAND2X0_HVT U243 ( .A1(n264), .A2(n265), .Y(n425) );
  XOR2X1_HVT U244 ( .A1(n317), .A2(n325), .Y(n560) );
  MUX41X1_HVT U245 ( .A1(n451), .A3(n447), .A2(n449), .A4(n443), .S0(n312), 
        .S1(n177), .Y(n442) );
  NBUFFX2_HVT U246 ( .A(n401), .Y(n307) );
  INVX1_HVT U247 ( .A(n280), .Y(n564) );
  MUX21X1_HVT U248 ( .A1(n593), .A2(n581), .S0(n231), .Y(n269) );
  INVX0_HVT U249 ( .A(in[7]), .Y(n272) );
  NAND2X0_HVT U250 ( .A1(n456), .A2(n272), .Y(n267) );
  INVX1_HVT U251 ( .A(n581), .Y(n366) );
  IBUFFX2_HVT U252 ( .A(n338), .Y(n335) );
  MUX21X1_HVT U253 ( .A1(n273), .A2(n396), .S0(n242), .Y(n585) );
  INVX1_HVT U254 ( .A(n585), .Y(n362) );
  NAND2X0_HVT U255 ( .A1(n466), .A2(n254), .Y(n268) );
  NAND2X0_HVT U256 ( .A1(n267), .A2(n268), .Y(out[5]) );
  MUX41X1_HVT U257 ( .A1(n512), .A3(n509), .A2(n514), .A4(n511), .S0(n312), 
        .S1(n311), .Y(n508) );
  IBUFFX2_HVT U258 ( .A(n593), .Y(n355) );
  MUX41X1_HVT U259 ( .A1(n374), .A3(n580), .A2(n513), .A4(n389), .S0(n271), 
        .S1(n270), .Y(n512) );
  MUX41X1_HVT U260 ( .A1(n472), .A3(n470), .A2(n469), .A4(n467), .S0(n177), 
        .S1(n312), .Y(n466) );
  MUX41X1_HVT U261 ( .A1(n324), .A3(n355), .A2(n273), .A4(n354), .S0(n266), 
        .S1(n270), .Y(n540) );
  INVX0_HVT U262 ( .A(in[3]), .Y(n398) );
  MUX21X2_HVT U263 ( .A1(n362), .A2(n554), .S0(n244), .Y(n550) );
  MUX41X1_HVT U264 ( .A1(n544), .A3(n541), .A2(n543), .A4(n540), .S0(n312), 
        .S1(n177), .Y(n539) );
  IBUFFX2_HVT U265 ( .A(n608), .Y(n279) );
  NBUFFX2_HVT U266 ( .A(n609), .Y(n275) );
  NBUFFX2_HVT U267 ( .A(n609), .Y(n276) );
  INVX1_HVT U268 ( .A(n275), .Y(n277) );
  INVX1_HVT U269 ( .A(n324), .Y(n287) );
  MUX21X1_HVT U270 ( .A1(n287), .A2(n399), .S0(n327), .Y(n441) );
  IBUFFX2_HVT U271 ( .A(n329), .Y(n326) );
  NBUFFX2_HVT U272 ( .A(n609), .Y(n324) );
  INVX1_HVT U273 ( .A(n322), .Y(n396) );
  NBUFFX2_HVT U274 ( .A(n398), .Y(n281) );
  NBUFFX2_HVT U275 ( .A(n398), .Y(n282) );
  MUX21X2_HVT U276 ( .A1(n445), .A2(n446), .S0(n302), .Y(n443) );
  NAND2X0_HVT U277 ( .A1(n582), .A2(n270), .Y(n283) );
  NAND2X0_HVT U278 ( .A1(n585), .A2(n244), .Y(n284) );
  NAND2X0_HVT U279 ( .A1(n283), .A2(n284), .Y(n446) );
  INVX1_HVT U280 ( .A(n414), .Y(n382) );
  MUX41X1_HVT U281 ( .A1(n287), .A3(n564), .A2(n294), .A4(n434), .S0(n298), 
        .S1(n270), .Y(n286) );
  INVX1_HVT U282 ( .A(n411), .Y(n385) );
  MUX41X1_HVT U283 ( .A1(n585), .A3(n588), .A2(n377), .A4(n397), .S0(n266), 
        .S1(n263), .Y(n469) );
  NBUFFX4_HVT U284 ( .A(n401), .Y(n308) );
  XOR2X1_HVT U285 ( .A1(n306), .A2(in[3]), .Y(n592) );
  NBUFFX2_HVT U286 ( .A(n608), .Y(n321) );
  NBUFFX2_HVT U287 ( .A(n608), .Y(n323) );
  NBUFFX2_HVT U288 ( .A(n608), .Y(n322) );
  AND2X1_HVT U289 ( .A1(n321), .A2(n593), .Y(n289) );
  MUX21X1_HVT U290 ( .A1(n378), .A2(n292), .S0(n303), .Y(n418) );
  MUX21X1_HVT U291 ( .A1(n317), .A2(n320), .S0(n325), .Y(n450) );
  XOR2X1_HVT U292 ( .A1(n276), .A2(n262), .Y(n571) );
  MUX21X1_HVT U293 ( .A1(n287), .A2(n397), .S0(n262), .Y(n580) );
  MUX21X1_HVT U294 ( .A1(n400), .A2(n281), .S0(n261), .Y(n569) );
  MUX21X1_HVT U295 ( .A1(n279), .A2(n285), .S0(n327), .Y(n575) );
  MUX21X1_HVT U296 ( .A1(n396), .A2(n307), .S0(n261), .Y(n414) );
  MUX21X1_HVT U297 ( .A1(n287), .A2(n308), .S0(n327), .Y(n439) );
  INVX1_HVT U298 ( .A(n314), .Y(n400) );
  NAND2X0_HVT U299 ( .A1(n398), .A2(n306), .Y(n608) );
  MUX21X1_HVT U300 ( .A1(n277), .A2(n316), .S0(n328), .Y(n409) );
  MUX21X1_HVT U301 ( .A1(n315), .A2(n281), .S0(n327), .Y(n587) );
  MUX21X1_HVT U302 ( .A1(n276), .A2(n323), .S0(n328), .Y(n594) );
  MUX21X1_HVT U303 ( .A1(n315), .A2(n277), .S0(n328), .Y(n577) );
  MUX21X1_HVT U304 ( .A1(n307), .A2(n279), .S0(n261), .Y(n582) );
  MUX21X1_HVT U305 ( .A1(n285), .A2(n308), .S0(n274), .Y(n404) );
  MUX21X1_HVT U306 ( .A1(n282), .A2(n279), .S0(n326), .Y(n578) );
  XNOR2X1_HVT U307 ( .A1(n323), .A2(n327), .Y(n290) );
  MUX21X1_HVT U308 ( .A1(n575), .A2(n289), .S0(n271), .Y(n483) );
  MUX21X1_HVT U309 ( .A1(n393), .A2(n290), .S0(n302), .Y(n486) );
  MUX21X1_HVT U310 ( .A1(n306), .A2(n323), .S0(n325), .Y(n505) );
  MUX21X1_HVT U311 ( .A1(n316), .A2(n397), .S0(n326), .Y(n574) );
  MUX21X1_HVT U312 ( .A1(n281), .A2(n399), .S0(n327), .Y(n565) );
  MUX21X1_HVT U313 ( .A1(n281), .A2(n322), .S0(n326), .Y(n412) );
  XOR2X1_HVT U314 ( .A1(n319), .A2(n325), .Y(n561) );
  XOR2X1_HVT U315 ( .A1(n314), .A2(n328), .Y(n562) );
  MUX21X1_HVT U316 ( .A1(n399), .A2(n282), .S0(n326), .Y(n413) );
  MUX21X1_HVT U317 ( .A1(n317), .A2(n321), .S0(n326), .Y(n403) );
  MUX21X1_HVT U318 ( .A1(n306), .A2(n316), .S0(n261), .Y(n568) );
  AND2X1_HVT U319 ( .A1(n603), .A2(n323), .Y(n291) );
  MUX21X1_HVT U320 ( .A1(n320), .A2(n321), .S0(n325), .Y(n590) );
  MUX21X1_HVT U321 ( .A1(n320), .A2(n282), .S0(n262), .Y(n589) );
  MUX21X1_HVT U322 ( .A1(n282), .A2(n307), .S0(n328), .Y(n563) );
  AND2X1_HVT U323 ( .A1(n325), .A2(n308), .Y(n292) );
  MUX21X1_HVT U324 ( .A1(n320), .A2(n307), .S0(n326), .Y(n489) );
  MUX21X1_HVT U325 ( .A1(n282), .A2(n320), .S0(n274), .Y(n406) );
  NBUFFX2_HVT U326 ( .A(n401), .Y(n306) );
  NBUFFX2_HVT U327 ( .A(n592), .Y(n314) );
  MUX21X1_HVT U328 ( .A1(n396), .A2(n399), .S0(n325), .Y(n558) );
  NBUFFX2_HVT U329 ( .A(n592), .Y(n315) );
  NBUFFX2_HVT U330 ( .A(n592), .Y(n316) );
  MUX21X1_HVT U331 ( .A1(n321), .A2(n318), .S0(n262), .Y(n468) );
  MUX21X1_HVT U332 ( .A1(n488), .A2(n490), .S0(n311), .Y(n487) );
  AND2X1_HVT U333 ( .A1(n320), .A2(n330), .Y(n293) );
  AND2X1_HVT U334 ( .A1(n399), .A2(n330), .Y(n294) );
  MUX21X1_HVT U335 ( .A1(n383), .A2(n340), .S0(n304), .Y(n534) );
  NBUFFX2_HVT U336 ( .A(n604), .Y(n317) );
  NBUFFX2_HVT U337 ( .A(n607), .Y(n319) );
  NBUFFX2_HVT U338 ( .A(n607), .Y(n320) );
  NBUFFX2_HVT U339 ( .A(n604), .Y(n318) );
  XNOR2X1_HVT U340 ( .A1(n231), .A2(n299), .Y(n295) );
  NBUFFX2_HVT U341 ( .A(n331), .Y(n302) );
  NBUFFX2_HVT U342 ( .A(n332), .Y(n299) );
  NBUFFX2_HVT U343 ( .A(n331), .Y(n297) );
  NBUFFX2_HVT U344 ( .A(n331), .Y(n298) );
  NBUFFX2_HVT U345 ( .A(n331), .Y(n296) );
  NBUFFX2_HVT U346 ( .A(n332), .Y(n300) );
  NBUFFX2_HVT U347 ( .A(n332), .Y(n301) );
  MUX21X1_HVT U348 ( .A1(n287), .A2(n273), .S0(n262), .Y(n402) );
  MUX21X1_HVT U349 ( .A1(n318), .A2(n273), .S0(n262), .Y(n513) );
  MUX21X1_HVT U350 ( .A1(n474), .A2(n475), .S0(n311), .Y(n473) );
  MUX21X1_HVT U351 ( .A1(n478), .A2(n479), .S0(n310), .Y(n477) );
  MUX21X1_HVT U352 ( .A1(n273), .A2(n276), .S0(n274), .Y(n408) );
  MUX21X1_HVT U353 ( .A1(n399), .A2(n397), .S0(n261), .Y(n494) );
  MUX21X1_HVT U354 ( .A1(n276), .A2(n273), .S0(n326), .Y(n453) );
  MUX21X1_HVT U355 ( .A1(n308), .A2(n273), .S0(n262), .Y(n581) );
  MUX21X1_HVT U356 ( .A1(n273), .A2(n318), .S0(n326), .Y(n407) );
  NBUFFX2_HVT U357 ( .A(in[2]), .Y(n332) );
  NBUFFX2_HVT U358 ( .A(in[2]), .Y(n331) );
  MUX21X1_HVT U359 ( .A1(n279), .A2(n288), .S0(n327), .Y(n476) );
  XOR2X1_HVT U360 ( .A1(n274), .A2(n288), .Y(n559) );
  MUX21X1_HVT U361 ( .A1(n288), .A2(n277), .S0(n261), .Y(n584) );
  MUX21X1_HVT U362 ( .A1(n320), .A2(n288), .S0(n325), .Y(n410) );
  MUX21X1_HVT U363 ( .A1(n288), .A2(n320), .S0(n328), .Y(n415) );
  MUX21X1_HVT U364 ( .A1(n288), .A2(n324), .S0(n327), .Y(n591) );
  MUX21X1_HVT U365 ( .A1(n281), .A2(n288), .S0(n261), .Y(n405) );
  MUX21X1_HVT U366 ( .A1(n318), .A2(n288), .S0(n325), .Y(n579) );
  INVX0_HVT U367 ( .A(in[6]), .Y(n401) );
  MUX21X1_HVT U368 ( .A1(n281), .A2(n400), .S0(n327), .Y(n411) );
  INVX0_HVT U369 ( .A(n597), .Y(n339) );
  INVX0_HVT U370 ( .A(n576), .Y(n340) );
  INVX0_HVT U371 ( .A(n570), .Y(n341) );
  INVX0_HVT U372 ( .A(n510), .Y(n342) );
  INVX0_HVT U373 ( .A(n471), .Y(n343) );
  INVX0_HVT U374 ( .A(n605), .Y(n345) );
  INVX0_HVT U375 ( .A(n566), .Y(n347) );
  INVX0_HVT U376 ( .A(n602), .Y(n348) );
  INVX0_HVT U377 ( .A(n573), .Y(n350) );
  INVX0_HVT U378 ( .A(n595), .Y(n351) );
  INVX0_HVT U379 ( .A(n600), .Y(n352) );
  INVX0_HVT U380 ( .A(n596), .Y(n353) );
  INVX0_HVT U381 ( .A(n594), .Y(n354) );
  INVX0_HVT U382 ( .A(n591), .Y(n356) );
  INVX0_HVT U383 ( .A(n590), .Y(n357) );
  INVX0_HVT U384 ( .A(n589), .Y(n358) );
  INVX0_HVT U385 ( .A(n588), .Y(n359) );
  INVX0_HVT U386 ( .A(n584), .Y(n363) );
  INVX0_HVT U387 ( .A(n582), .Y(n365) );
  INVX0_HVT U388 ( .A(n580), .Y(n367) );
  INVX0_HVT U389 ( .A(n578), .Y(n369) );
  INVX0_HVT U390 ( .A(n577), .Y(n370) );
  INVX0_HVT U391 ( .A(n575), .Y(n371) );
  INVX0_HVT U392 ( .A(n572), .Y(n373) );
  INVX0_HVT U393 ( .A(n569), .Y(n375) );
  INVX0_HVT U394 ( .A(n568), .Y(n376) );
  INVX0_HVT U395 ( .A(n565), .Y(n377) );
  INVX0_HVT U396 ( .A(n562), .Y(n379) );
  INVX0_HVT U397 ( .A(n599), .Y(n380) );
  INVX0_HVT U398 ( .A(n415), .Y(n381) );
  INVX0_HVT U399 ( .A(n413), .Y(n383) );
  INVX0_HVT U400 ( .A(n410), .Y(n386) );
  INVX0_HVT U401 ( .A(n409), .Y(n387) );
  INVX0_HVT U402 ( .A(n408), .Y(n388) );
  INVX0_HVT U403 ( .A(n407), .Y(n389) );
  INVX0_HVT U404 ( .A(n406), .Y(n390) );
  INVX0_HVT U405 ( .A(n405), .Y(n391) );
  INVX0_HVT U406 ( .A(n453), .Y(n392) );
  INVX0_HVT U407 ( .A(n404), .Y(n393) );
  INVX0_HVT U408 ( .A(n403), .Y(n394) );
  INVX0_HVT U409 ( .A(n402), .Y(n395) );
endmodule

