
module inv_aes ( clk, rest, start, plaintext1, local_key, cipher_text, done, 
        busy );
  input [127:0] plaintext1;
  input [127:0] local_key;
  output [127:0] cipher_text;
  input clk, rest, start;
  output done, busy;
  wire   last, done_k, flag, n12, n13, n14, n15, n16, n17, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n18, n155, n207, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366;
  wire   [127:0] adk_out;
  wire   [127:0] keys1;
  wire   [127:0] out1;
  wire   [3:0] rount_no;
  wire   [127:0] key_round;
  wire   [3:0] state;
  tri   clk;
  tri   rest;

  DFFX1_HVT \rount_no_reg[0]  ( .D(n601), .CLK(clk), .Q(rount_no[0]) );
  DFFX1_HVT \state_reg[1]  ( .D(n596), .CLK(clk), .Q(state[1]), .QN(n14) );
  DFFX1_HVT \state_reg[3]  ( .D(n599), .CLK(clk), .Q(state[3]), .QN(n12) );
  DFFX1_HVT \state_reg[2]  ( .D(n597), .CLK(clk), .Q(state[2]), .QN(n13) );
  DFFX1_HVT done_reg ( .D(n591), .CLK(clk), .Q(done), .QN(n17) );
  DFFX1_HVT busy_reg ( .D(n600), .CLK(clk), .Q(busy), .QN(n16) );
  DFFX1_HVT \state_reg[0]  ( .D(n598), .CLK(clk), .Q(state[0]), .QN(n15) );
  DFFX1_HVT last_reg ( .D(n595), .CLK(clk), .Q(last) );
  DFFX1_HVT \rount_no_reg[3]  ( .D(n592), .CLK(clk), .Q(rount_no[3]) );
  DFFX1_HVT \rount_no_reg[2]  ( .D(n593), .CLK(clk), .Q(rount_no[2]) );
  DFFX1_HVT \rount_no_reg[1]  ( .D(n594), .CLK(clk), .Q(rount_no[1]) );
  DFFX1_HVT \keys1_reg[0]  ( .D(n590), .CLK(clk), .Q(keys1[0]) );
  DFFX1_HVT \keys1_reg[1]  ( .D(n589), .CLK(clk), .Q(keys1[1]) );
  DFFX1_HVT \keys1_reg[2]  ( .D(n588), .CLK(clk), .Q(keys1[2]) );
  DFFX1_HVT \keys1_reg[3]  ( .D(n587), .CLK(clk), .Q(keys1[3]) );
  DFFX1_HVT \keys1_reg[4]  ( .D(n586), .CLK(clk), .Q(keys1[4]) );
  DFFX1_HVT \keys1_reg[5]  ( .D(n585), .CLK(clk), .Q(keys1[5]) );
  DFFX1_HVT \keys1_reg[6]  ( .D(n584), .CLK(clk), .Q(keys1[6]) );
  DFFX1_HVT \keys1_reg[7]  ( .D(n583), .CLK(clk), .Q(keys1[7]) );
  DFFX1_HVT \keys1_reg[8]  ( .D(n582), .CLK(clk), .Q(keys1[8]) );
  DFFX1_HVT \keys1_reg[9]  ( .D(n581), .CLK(clk), .Q(keys1[9]) );
  DFFX1_HVT \keys1_reg[10]  ( .D(n580), .CLK(clk), .Q(keys1[10]) );
  DFFX1_HVT \keys1_reg[11]  ( .D(n579), .CLK(clk), .Q(keys1[11]) );
  DFFX1_HVT \keys1_reg[12]  ( .D(n578), .CLK(clk), .Q(keys1[12]) );
  DFFX1_HVT \keys1_reg[13]  ( .D(n577), .CLK(clk), .Q(keys1[13]) );
  DFFX1_HVT \keys1_reg[14]  ( .D(n576), .CLK(clk), .Q(keys1[14]) );
  DFFX1_HVT \keys1_reg[15]  ( .D(n575), .CLK(clk), .Q(keys1[15]) );
  DFFX1_HVT \keys1_reg[16]  ( .D(n574), .CLK(clk), .Q(keys1[16]) );
  DFFX1_HVT \keys1_reg[17]  ( .D(n573), .CLK(clk), .Q(keys1[17]) );
  DFFX1_HVT \keys1_reg[18]  ( .D(n572), .CLK(clk), .Q(keys1[18]) );
  DFFX1_HVT \keys1_reg[19]  ( .D(n571), .CLK(clk), .Q(keys1[19]) );
  DFFX1_HVT \keys1_reg[20]  ( .D(n570), .CLK(clk), .Q(keys1[20]) );
  DFFX1_HVT \keys1_reg[21]  ( .D(n569), .CLK(clk), .Q(keys1[21]) );
  DFFX1_HVT \keys1_reg[22]  ( .D(n568), .CLK(clk), .Q(keys1[22]) );
  DFFX1_HVT \keys1_reg[23]  ( .D(n567), .CLK(clk), .Q(keys1[23]) );
  DFFX1_HVT \keys1_reg[24]  ( .D(n566), .CLK(clk), .Q(keys1[24]) );
  DFFX1_HVT \keys1_reg[25]  ( .D(n565), .CLK(clk), .Q(keys1[25]) );
  DFFX1_HVT \keys1_reg[26]  ( .D(n564), .CLK(clk), .Q(keys1[26]) );
  DFFX1_HVT \keys1_reg[27]  ( .D(n563), .CLK(clk), .Q(keys1[27]) );
  DFFX1_HVT \keys1_reg[28]  ( .D(n562), .CLK(clk), .Q(keys1[28]) );
  DFFX1_HVT \keys1_reg[29]  ( .D(n561), .CLK(clk), .Q(keys1[29]) );
  DFFX1_HVT \keys1_reg[30]  ( .D(n560), .CLK(clk), .Q(keys1[30]) );
  DFFX1_HVT \keys1_reg[31]  ( .D(n559), .CLK(clk), .Q(keys1[31]) );
  DFFX1_HVT \keys1_reg[32]  ( .D(n558), .CLK(clk), .Q(keys1[32]) );
  DFFX1_HVT \keys1_reg[33]  ( .D(n557), .CLK(clk), .Q(keys1[33]) );
  DFFX1_HVT \keys1_reg[34]  ( .D(n556), .CLK(clk), .Q(keys1[34]) );
  DFFX1_HVT \keys1_reg[35]  ( .D(n555), .CLK(clk), .Q(keys1[35]) );
  DFFX1_HVT \keys1_reg[36]  ( .D(n554), .CLK(clk), .Q(keys1[36]) );
  DFFX1_HVT \keys1_reg[37]  ( .D(n553), .CLK(clk), .Q(keys1[37]) );
  DFFX1_HVT \keys1_reg[38]  ( .D(n552), .CLK(clk), .Q(keys1[38]) );
  DFFX1_HVT \keys1_reg[39]  ( .D(n551), .CLK(clk), .Q(keys1[39]) );
  DFFX1_HVT \keys1_reg[40]  ( .D(n550), .CLK(clk), .Q(keys1[40]) );
  DFFX1_HVT \keys1_reg[41]  ( .D(n549), .CLK(clk), .Q(keys1[41]) );
  DFFX1_HVT \keys1_reg[42]  ( .D(n548), .CLK(clk), .Q(keys1[42]) );
  DFFX1_HVT \keys1_reg[43]  ( .D(n547), .CLK(clk), .Q(keys1[43]) );
  DFFX1_HVT \keys1_reg[44]  ( .D(n546), .CLK(clk), .Q(keys1[44]) );
  DFFX1_HVT \keys1_reg[45]  ( .D(n545), .CLK(clk), .Q(keys1[45]) );
  DFFX1_HVT \keys1_reg[46]  ( .D(n544), .CLK(clk), .Q(keys1[46]) );
  DFFX1_HVT \keys1_reg[47]  ( .D(n543), .CLK(clk), .Q(keys1[47]) );
  DFFX1_HVT \keys1_reg[48]  ( .D(n542), .CLK(clk), .Q(keys1[48]) );
  DFFX1_HVT \keys1_reg[49]  ( .D(n541), .CLK(clk), .Q(keys1[49]) );
  DFFX1_HVT \keys1_reg[50]  ( .D(n540), .CLK(clk), .Q(keys1[50]) );
  DFFX1_HVT \keys1_reg[51]  ( .D(n539), .CLK(clk), .Q(keys1[51]) );
  DFFX1_HVT \keys1_reg[52]  ( .D(n538), .CLK(clk), .Q(keys1[52]) );
  DFFX1_HVT \keys1_reg[53]  ( .D(n537), .CLK(clk), .Q(keys1[53]) );
  DFFX1_HVT \keys1_reg[54]  ( .D(n536), .CLK(clk), .Q(keys1[54]) );
  DFFX1_HVT \keys1_reg[55]  ( .D(n535), .CLK(clk), .Q(keys1[55]) );
  DFFX1_HVT \keys1_reg[56]  ( .D(n534), .CLK(clk), .Q(keys1[56]) );
  DFFX1_HVT \keys1_reg[57]  ( .D(n533), .CLK(clk), .Q(keys1[57]) );
  DFFX1_HVT \keys1_reg[58]  ( .D(n532), .CLK(clk), .Q(keys1[58]) );
  DFFX1_HVT \keys1_reg[59]  ( .D(n531), .CLK(clk), .Q(keys1[59]) );
  DFFX1_HVT \keys1_reg[60]  ( .D(n530), .CLK(clk), .Q(keys1[60]) );
  DFFX1_HVT \keys1_reg[61]  ( .D(n529), .CLK(clk), .Q(keys1[61]) );
  DFFX1_HVT \keys1_reg[62]  ( .D(n528), .CLK(clk), .Q(keys1[62]) );
  DFFX1_HVT \keys1_reg[63]  ( .D(n527), .CLK(clk), .Q(keys1[63]) );
  DFFX1_HVT \keys1_reg[64]  ( .D(n526), .CLK(clk), .Q(keys1[64]) );
  DFFX1_HVT \keys1_reg[65]  ( .D(n525), .CLK(clk), .Q(keys1[65]) );
  DFFX1_HVT \keys1_reg[66]  ( .D(n524), .CLK(clk), .Q(keys1[66]) );
  DFFX1_HVT \keys1_reg[67]  ( .D(n523), .CLK(clk), .Q(keys1[67]) );
  DFFX1_HVT \keys1_reg[68]  ( .D(n522), .CLK(clk), .Q(keys1[68]) );
  DFFX1_HVT \keys1_reg[69]  ( .D(n521), .CLK(clk), .Q(keys1[69]) );
  DFFX1_HVT \keys1_reg[70]  ( .D(n520), .CLK(clk), .Q(keys1[70]) );
  DFFX1_HVT \keys1_reg[71]  ( .D(n519), .CLK(clk), .Q(keys1[71]) );
  DFFX1_HVT \keys1_reg[72]  ( .D(n518), .CLK(clk), .Q(keys1[72]) );
  DFFX1_HVT \keys1_reg[73]  ( .D(n517), .CLK(clk), .Q(keys1[73]) );
  DFFX1_HVT \keys1_reg[74]  ( .D(n516), .CLK(clk), .Q(keys1[74]) );
  DFFX1_HVT \keys1_reg[75]  ( .D(n515), .CLK(clk), .Q(keys1[75]) );
  DFFX1_HVT \keys1_reg[76]  ( .D(n514), .CLK(clk), .Q(keys1[76]) );
  DFFX1_HVT \keys1_reg[77]  ( .D(n513), .CLK(clk), .Q(keys1[77]) );
  DFFX1_HVT \keys1_reg[78]  ( .D(n512), .CLK(clk), .Q(keys1[78]) );
  DFFX1_HVT \keys1_reg[79]  ( .D(n511), .CLK(clk), .Q(keys1[79]) );
  DFFX1_HVT \keys1_reg[80]  ( .D(n510), .CLK(clk), .Q(keys1[80]) );
  DFFX1_HVT \keys1_reg[81]  ( .D(n509), .CLK(clk), .Q(keys1[81]) );
  DFFX1_HVT \keys1_reg[82]  ( .D(n508), .CLK(clk), .Q(keys1[82]) );
  DFFX1_HVT \keys1_reg[83]  ( .D(n507), .CLK(clk), .Q(keys1[83]) );
  DFFX1_HVT \keys1_reg[84]  ( .D(n506), .CLK(clk), .Q(keys1[84]) );
  DFFX1_HVT \keys1_reg[85]  ( .D(n505), .CLK(clk), .Q(keys1[85]) );
  DFFX1_HVT \keys1_reg[86]  ( .D(n504), .CLK(clk), .Q(keys1[86]) );
  DFFX1_HVT \keys1_reg[87]  ( .D(n503), .CLK(clk), .Q(keys1[87]) );
  DFFX1_HVT \keys1_reg[88]  ( .D(n502), .CLK(clk), .Q(keys1[88]) );
  DFFX1_HVT \keys1_reg[89]  ( .D(n501), .CLK(clk), .Q(keys1[89]), .QN(n991) );
  DFFX1_HVT \keys1_reg[90]  ( .D(n500), .CLK(clk), .Q(keys1[90]) );
  DFFX1_HVT \keys1_reg[91]  ( .D(n499), .CLK(clk), .Q(keys1[91]), .QN(n1167)
         );
  DFFX1_HVT \keys1_reg[92]  ( .D(n498), .CLK(clk), .Q(keys1[92]) );
  DFFX1_HVT \keys1_reg[93]  ( .D(n497), .CLK(clk), .Q(keys1[93]) );
  DFFX1_HVT \keys1_reg[94]  ( .D(n496), .CLK(clk), .Q(keys1[94]) );
  DFFX1_HVT \keys1_reg[95]  ( .D(n495), .CLK(clk), .Q(keys1[95]) );
  DFFX1_HVT \keys1_reg[96]  ( .D(n494), .CLK(clk), .Q(keys1[96]) );
  DFFX1_HVT \keys1_reg[97]  ( .D(n493), .CLK(clk), .Q(keys1[97]) );
  DFFX1_HVT \keys1_reg[98]  ( .D(n492), .CLK(clk), .Q(keys1[98]) );
  DFFX1_HVT \keys1_reg[99]  ( .D(n491), .CLK(clk), .Q(keys1[99]) );
  DFFX1_HVT \keys1_reg[100]  ( .D(n490), .CLK(clk), .Q(keys1[100]) );
  DFFX1_HVT \keys1_reg[101]  ( .D(n489), .CLK(clk), .Q(keys1[101]) );
  DFFX1_HVT \keys1_reg[102]  ( .D(n488), .CLK(clk), .Q(keys1[102]) );
  DFFX1_HVT \keys1_reg[103]  ( .D(n487), .CLK(clk), .Q(keys1[103]) );
  DFFX1_HVT \keys1_reg[104]  ( .D(n486), .CLK(clk), .Q(keys1[104]) );
  DFFX1_HVT \keys1_reg[105]  ( .D(n485), .CLK(clk), .Q(keys1[105]) );
  DFFX1_HVT \keys1_reg[106]  ( .D(n484), .CLK(clk), .Q(keys1[106]) );
  DFFX1_HVT \keys1_reg[107]  ( .D(n483), .CLK(clk), .Q(keys1[107]), .QN(n1170)
         );
  DFFX1_HVT \keys1_reg[108]  ( .D(n482), .CLK(clk), .Q(keys1[108]) );
  DFFX1_HVT \keys1_reg[109]  ( .D(n481), .CLK(clk), .Q(keys1[109]) );
  DFFX1_HVT \keys1_reg[110]  ( .D(n480), .CLK(clk), .Q(keys1[110]) );
  DFFX1_HVT \keys1_reg[111]  ( .D(n479), .CLK(clk), .Q(keys1[111]) );
  DFFX1_HVT \keys1_reg[112]  ( .D(n478), .CLK(clk), .Q(keys1[112]) );
  DFFX1_HVT \keys1_reg[113]  ( .D(n477), .CLK(clk), .Q(keys1[113]) );
  DFFX1_HVT \keys1_reg[114]  ( .D(n476), .CLK(clk), .Q(keys1[114]) );
  DFFX1_HVT \keys1_reg[115]  ( .D(n475), .CLK(clk), .Q(keys1[115]) );
  DFFX1_HVT \keys1_reg[116]  ( .D(n474), .CLK(clk), .Q(keys1[116]) );
  DFFX1_HVT \keys1_reg[117]  ( .D(n473), .CLK(clk), .Q(keys1[117]) );
  DFFX1_HVT \keys1_reg[118]  ( .D(n472), .CLK(clk), .Q(keys1[118]) );
  DFFX1_HVT \keys1_reg[119]  ( .D(n471), .CLK(clk), .Q(keys1[119]) );
  DFFX1_HVT \keys1_reg[120]  ( .D(n470), .CLK(clk), .Q(keys1[120]) );
  DFFX1_HVT \keys1_reg[121]  ( .D(n469), .CLK(clk), .Q(keys1[121]) );
  DFFX1_HVT \keys1_reg[122]  ( .D(n468), .CLK(clk), .Q(keys1[122]) );
  DFFX1_HVT \keys1_reg[123]  ( .D(n467), .CLK(clk), .Q(keys1[123]), .QN(n1172)
         );
  DFFX1_HVT \keys1_reg[124]  ( .D(n466), .CLK(clk), .Q(keys1[124]) );
  DFFX1_HVT \keys1_reg[125]  ( .D(n465), .CLK(clk), .Q(keys1[125]) );
  DFFX1_HVT \keys1_reg[126]  ( .D(n464), .CLK(clk), .Q(keys1[126]), .QN(n994)
         );
  DFFX1_HVT \keys1_reg[127]  ( .D(n463), .CLK(clk), .Q(keys1[127]) );
  DFFX1_HVT \adk_out_reg[127]  ( .D(n335), .CLK(clk), .Q(adk_out[127]), .QN(
        n666) );
  DFFX1_HVT \adk_out_reg[0]  ( .D(n462), .CLK(clk), .Q(adk_out[0]), .QN(n920)
         );
  DFFX1_HVT \cipher_text_reg[0]  ( .D(n334), .CLK(clk), .Q(cipher_text[0]) );
  DFFX1_HVT \adk_out_reg[1]  ( .D(n461), .CLK(clk), .Q(adk_out[1]) );
  DFFX1_HVT \cipher_text_reg[1]  ( .D(n333), .CLK(clk), .Q(cipher_text[1]) );
  DFFX1_HVT \adk_out_reg[2]  ( .D(n460), .CLK(clk), .Q(adk_out[2]) );
  DFFX1_HVT \cipher_text_reg[2]  ( .D(n332), .CLK(clk), .Q(cipher_text[2]) );
  DFFX1_HVT \adk_out_reg[3]  ( .D(n459), .CLK(clk), .Q(n1183), .QN(n632) );
  DFFX1_HVT \cipher_text_reg[3]  ( .D(n331), .CLK(clk), .Q(cipher_text[3]) );
  DFFX1_HVT \adk_out_reg[4]  ( .D(n458), .CLK(clk), .Q(adk_out[4]), .QN(n902)
         );
  DFFX1_HVT \cipher_text_reg[4]  ( .D(n330), .CLK(clk), .Q(cipher_text[4]) );
  DFFX1_HVT \adk_out_reg[5]  ( .D(n457), .CLK(clk), .Q(adk_out[5]) );
  DFFX1_HVT \cipher_text_reg[5]  ( .D(n329), .CLK(clk), .Q(cipher_text[5]) );
  DFFX1_HVT \adk_out_reg[6]  ( .D(n456), .CLK(clk), .Q(adk_out[6]), .QN(n656)
         );
  DFFX1_HVT \cipher_text_reg[6]  ( .D(n328), .CLK(clk), .Q(cipher_text[6]) );
  DFFX1_HVT \adk_out_reg[7]  ( .D(n455), .CLK(clk), .Q(adk_out[7]), .QN(n1036)
         );
  DFFX1_HVT \cipher_text_reg[7]  ( .D(n327), .CLK(clk), .Q(cipher_text[7]) );
  DFFX1_HVT \adk_out_reg[8]  ( .D(n454), .CLK(clk), .Q(adk_out[8]), .QN(n779)
         );
  DFFX1_HVT \cipher_text_reg[8]  ( .D(n326), .CLK(clk), .Q(cipher_text[8]) );
  DFFX1_HVT \adk_out_reg[9]  ( .D(n453), .CLK(clk), .Q(adk_out[9]) );
  DFFX1_HVT \cipher_text_reg[9]  ( .D(n325), .CLK(clk), .Q(cipher_text[9]) );
  DFFX1_HVT \adk_out_reg[10]  ( .D(n452), .CLK(clk), .Q(adk_out[10]) );
  DFFX1_HVT \cipher_text_reg[10]  ( .D(n324), .CLK(clk), .Q(cipher_text[10])
         );
  DFFX1_HVT \adk_out_reg[11]  ( .D(n451), .CLK(clk), .Q(adk_out[11]), .QN(n9)
         );
  DFFX1_HVT \cipher_text_reg[11]  ( .D(n323), .CLK(clk), .Q(cipher_text[11])
         );
  DFFX1_HVT \adk_out_reg[12]  ( .D(n450), .CLK(clk), .Q(adk_out[12]) );
  DFFX1_HVT \cipher_text_reg[12]  ( .D(n322), .CLK(clk), .Q(cipher_text[12])
         );
  DFFX1_HVT \adk_out_reg[13]  ( .D(n449), .CLK(clk), .Q(adk_out[13]) );
  DFFX1_HVT \cipher_text_reg[13]  ( .D(n321), .CLK(clk), .Q(cipher_text[13])
         );
  DFFX1_HVT \adk_out_reg[14]  ( .D(n448), .CLK(clk), .Q(n1207) );
  DFFX1_HVT \cipher_text_reg[14]  ( .D(n320), .CLK(clk), .Q(cipher_text[14])
         );
  DFFX1_HVT \adk_out_reg[15]  ( .D(n447), .CLK(clk), .Q(adk_out[15]) );
  DFFX1_HVT \cipher_text_reg[15]  ( .D(n319), .CLK(clk), .Q(cipher_text[15])
         );
  DFFX1_HVT \adk_out_reg[16]  ( .D(n446), .CLK(clk), .Q(adk_out[16]), .QN(n843) );
  DFFX1_HVT \cipher_text_reg[16]  ( .D(n318), .CLK(clk), .Q(cipher_text[16])
         );
  DFFX1_HVT \adk_out_reg[17]  ( .D(n445), .CLK(clk), .Q(adk_out[17]) );
  DFFX1_HVT \cipher_text_reg[17]  ( .D(n317), .CLK(clk), .Q(cipher_text[17])
         );
  DFFX1_HVT \adk_out_reg[18]  ( .D(n444), .CLK(clk), .Q(adk_out[18]) );
  DFFX1_HVT \cipher_text_reg[18]  ( .D(n316), .CLK(clk), .Q(cipher_text[18])
         );
  DFFX1_HVT \adk_out_reg[19]  ( .D(n443), .CLK(clk), .Q(adk_out[19]) );
  DFFX1_HVT \cipher_text_reg[19]  ( .D(n315), .CLK(clk), .Q(cipher_text[19])
         );
  DFFX1_HVT \adk_out_reg[20]  ( .D(n442), .CLK(clk), .Q(adk_out[20]), .QN(n685) );
  DFFX1_HVT \cipher_text_reg[20]  ( .D(n314), .CLK(clk), .Q(cipher_text[20])
         );
  DFFX1_HVT \adk_out_reg[21]  ( .D(n441), .CLK(clk), .Q(adk_out[21]) );
  DFFX1_HVT \cipher_text_reg[21]  ( .D(n313), .CLK(clk), .Q(cipher_text[21])
         );
  DFFX1_HVT \adk_out_reg[22]  ( .D(n440), .CLK(clk), .Q(adk_out[22]), .QN(n681) );
  DFFX1_HVT \cipher_text_reg[22]  ( .D(n312), .CLK(clk), .Q(cipher_text[22])
         );
  DFFX1_HVT \adk_out_reg[23]  ( .D(n439), .CLK(clk), .Q(adk_out[23]) );
  DFFX1_HVT \cipher_text_reg[23]  ( .D(n311), .CLK(clk), .Q(cipher_text[23])
         );
  DFFX1_HVT \adk_out_reg[24]  ( .D(n438), .CLK(clk), .Q(adk_out[24]), .QN(n922) );
  DFFX1_HVT \cipher_text_reg[24]  ( .D(n310), .CLK(clk), .Q(cipher_text[24])
         );
  DFFX1_HVT \adk_out_reg[25]  ( .D(n437), .CLK(clk), .Q(adk_out[25]) );
  DFFX1_HVT \cipher_text_reg[25]  ( .D(n309), .CLK(clk), .Q(cipher_text[25])
         );
  DFFX1_HVT \adk_out_reg[26]  ( .D(n436), .CLK(clk), .Q(adk_out[26]) );
  DFFX1_HVT \cipher_text_reg[26]  ( .D(n308), .CLK(clk), .Q(cipher_text[26])
         );
  DFFX1_HVT \adk_out_reg[27]  ( .D(n435), .CLK(clk), .Q(n1093) );
  DFFX1_HVT \cipher_text_reg[27]  ( .D(n307), .CLK(clk), .Q(cipher_text[27])
         );
  DFFX1_HVT \adk_out_reg[28]  ( .D(n434), .CLK(clk), .Q(adk_out[28]), .QN(n672) );
  DFFX1_HVT \cipher_text_reg[28]  ( .D(n306), .CLK(clk), .Q(cipher_text[28])
         );
  DFFX1_HVT \adk_out_reg[29]  ( .D(n433), .CLK(clk), .Q(adk_out[29]) );
  DFFX1_HVT \cipher_text_reg[29]  ( .D(n305), .CLK(clk), .Q(cipher_text[29])
         );
  DFFX1_HVT \adk_out_reg[30]  ( .D(n432), .CLK(clk), .Q(adk_out[30]) );
  DFFX1_HVT \cipher_text_reg[30]  ( .D(n304), .CLK(clk), .Q(cipher_text[30])
         );
  DFFX1_HVT \adk_out_reg[31]  ( .D(n431), .CLK(clk), .Q(adk_out[31]), .QN(
        n1039) );
  DFFX1_HVT \cipher_text_reg[31]  ( .D(n303), .CLK(clk), .Q(cipher_text[31])
         );
  DFFX1_HVT \adk_out_reg[32]  ( .D(n430), .CLK(clk), .Q(adk_out[32]), .QN(n904) );
  DFFX1_HVT \cipher_text_reg[32]  ( .D(n302), .CLK(clk), .Q(cipher_text[32])
         );
  DFFX1_HVT \adk_out_reg[33]  ( .D(n429), .CLK(clk), .Q(adk_out[33]) );
  DFFX1_HVT \cipher_text_reg[33]  ( .D(n301), .CLK(clk), .Q(cipher_text[33])
         );
  DFFX1_HVT \adk_out_reg[34]  ( .D(n428), .CLK(clk), .Q(adk_out[34]) );
  DFFX1_HVT \cipher_text_reg[34]  ( .D(n300), .CLK(clk), .Q(cipher_text[34])
         );
  DFFX1_HVT \adk_out_reg[35]  ( .D(n427), .CLK(clk), .Q(n1182), .QN(n11) );
  DFFX1_HVT \cipher_text_reg[35]  ( .D(n299), .CLK(clk), .Q(cipher_text[35])
         );
  DFFX1_HVT \adk_out_reg[36]  ( .D(n426), .CLK(clk), .Q(adk_out[36]), .QN(n813) );
  DFFX1_HVT \cipher_text_reg[36]  ( .D(n298), .CLK(clk), .Q(cipher_text[36])
         );
  DFFX1_HVT \adk_out_reg[37]  ( .D(n425), .CLK(clk), .Q(adk_out[37]) );
  DFFX1_HVT \cipher_text_reg[37]  ( .D(n297), .CLK(clk), .Q(cipher_text[37])
         );
  DFFX1_HVT \adk_out_reg[38]  ( .D(n424), .CLK(clk), .Q(adk_out[38]) );
  DFFX1_HVT \cipher_text_reg[38]  ( .D(n296), .CLK(clk), .Q(cipher_text[38])
         );
  DFFX1_HVT \adk_out_reg[39]  ( .D(n423), .CLK(clk), .Q(adk_out[39]) );
  DFFX1_HVT \cipher_text_reg[39]  ( .D(n295), .CLK(clk), .Q(cipher_text[39])
         );
  DFFX1_HVT \adk_out_reg[40]  ( .D(n422), .CLK(clk), .Q(adk_out[40]) );
  DFFX1_HVT \cipher_text_reg[40]  ( .D(n294), .CLK(clk), .Q(cipher_text[40])
         );
  DFFX1_HVT \adk_out_reg[41]  ( .D(n421), .CLK(clk), .Q(adk_out[41]) );
  DFFX1_HVT \cipher_text_reg[41]  ( .D(n293), .CLK(clk), .Q(cipher_text[41])
         );
  DFFX1_HVT \adk_out_reg[42]  ( .D(n420), .CLK(clk), .Q(adk_out[42]) );
  DFFX1_HVT \cipher_text_reg[42]  ( .D(n292), .CLK(clk), .Q(cipher_text[42])
         );
  DFFX1_HVT \adk_out_reg[43]  ( .D(n419), .CLK(clk), .Q(n1178) );
  DFFX1_HVT \cipher_text_reg[43]  ( .D(n291), .CLK(clk), .Q(cipher_text[43])
         );
  DFFX1_HVT \adk_out_reg[44]  ( .D(n418), .CLK(clk), .Q(adk_out[44]) );
  DFFX1_HVT \cipher_text_reg[44]  ( .D(n290), .CLK(clk), .Q(cipher_text[44])
         );
  DFFX1_HVT \adk_out_reg[45]  ( .D(n417), .CLK(clk), .Q(adk_out[45]) );
  DFFX1_HVT \cipher_text_reg[45]  ( .D(n289), .CLK(clk), .Q(cipher_text[45])
         );
  DFFX1_HVT \adk_out_reg[46]  ( .D(n416), .CLK(clk), .Q(adk_out[46]) );
  DFFX1_HVT \cipher_text_reg[46]  ( .D(n288), .CLK(clk), .Q(cipher_text[46])
         );
  DFFX1_HVT \adk_out_reg[47]  ( .D(n415), .CLK(clk), .Q(adk_out[47]) );
  DFFX1_HVT \cipher_text_reg[47]  ( .D(n287), .CLK(clk), .Q(cipher_text[47])
         );
  DFFX1_HVT \adk_out_reg[48]  ( .D(n414), .CLK(clk), .Q(adk_out[48]), .QN(n865) );
  DFFX1_HVT \cipher_text_reg[48]  ( .D(n286), .CLK(clk), .Q(cipher_text[48])
         );
  DFFX1_HVT \adk_out_reg[49]  ( .D(n413), .CLK(clk), .Q(adk_out[49]) );
  DFFX1_HVT \cipher_text_reg[49]  ( .D(n285), .CLK(clk), .Q(cipher_text[49])
         );
  DFFX1_HVT \adk_out_reg[50]  ( .D(n412), .CLK(clk), .Q(adk_out[50]) );
  DFFX1_HVT \cipher_text_reg[50]  ( .D(n284), .CLK(clk), .Q(cipher_text[50])
         );
  DFFX1_HVT \adk_out_reg[51]  ( .D(n411), .CLK(clk), .Q(n1173) );
  DFFX1_HVT \cipher_text_reg[51]  ( .D(n283), .CLK(clk), .Q(cipher_text[51])
         );
  DFFX1_HVT \adk_out_reg[52]  ( .D(n410), .CLK(clk), .Q(adk_out[52]), .QN(
        n1038) );
  DFFX1_HVT \cipher_text_reg[52]  ( .D(n282), .CLK(clk), .Q(cipher_text[52])
         );
  DFFX1_HVT \adk_out_reg[53]  ( .D(n409), .CLK(clk), .Q(adk_out[53]) );
  DFFX1_HVT \cipher_text_reg[53]  ( .D(n281), .CLK(clk), .Q(cipher_text[53])
         );
  DFFX1_HVT \adk_out_reg[54]  ( .D(n408), .CLK(clk), .Q(adk_out[54]) );
  DFFX1_HVT \cipher_text_reg[54]  ( .D(n280), .CLK(clk), .Q(cipher_text[54])
         );
  DFFX1_HVT \adk_out_reg[55]  ( .D(n407), .CLK(clk), .Q(adk_out[55]) );
  DFFX1_HVT \cipher_text_reg[55]  ( .D(n279), .CLK(clk), .Q(cipher_text[55])
         );
  DFFX1_HVT \adk_out_reg[56]  ( .D(n406), .CLK(clk), .Q(adk_out[56]) );
  DFFX1_HVT \cipher_text_reg[56]  ( .D(n278), .CLK(clk), .Q(cipher_text[56])
         );
  DFFX1_HVT \adk_out_reg[57]  ( .D(n405), .CLK(clk), .Q(adk_out[57]) );
  DFFX1_HVT \cipher_text_reg[57]  ( .D(n277), .CLK(clk), .Q(cipher_text[57])
         );
  DFFX1_HVT \adk_out_reg[58]  ( .D(n404), .CLK(clk), .Q(adk_out[58]) );
  DFFX1_HVT \cipher_text_reg[58]  ( .D(n276), .CLK(clk), .Q(cipher_text[58])
         );
  DFFX1_HVT \adk_out_reg[59]  ( .D(n403), .CLK(clk), .Q(adk_out[59]), .QN(
        n1156) );
  DFFX1_HVT \cipher_text_reg[59]  ( .D(n275), .CLK(clk), .Q(cipher_text[59])
         );
  DFFX1_HVT \adk_out_reg[60]  ( .D(n402), .CLK(clk), .Q(adk_out[60]) );
  DFFX1_HVT \cipher_text_reg[60]  ( .D(n274), .CLK(clk), .Q(cipher_text[60])
         );
  DFFX1_HVT \adk_out_reg[61]  ( .D(n401), .CLK(clk), .Q(adk_out[61]) );
  DFFX1_HVT \cipher_text_reg[61]  ( .D(n273), .CLK(clk), .Q(cipher_text[61])
         );
  DFFX1_HVT \adk_out_reg[62]  ( .D(n400), .CLK(clk), .Q(adk_out[62]) );
  DFFX1_HVT \cipher_text_reg[62]  ( .D(n272), .CLK(clk), .Q(cipher_text[62])
         );
  DFFX1_HVT \adk_out_reg[63]  ( .D(n399), .CLK(clk), .Q(adk_out[63]) );
  DFFX1_HVT \cipher_text_reg[63]  ( .D(n271), .CLK(clk), .Q(cipher_text[63])
         );
  DFFX1_HVT \adk_out_reg[64]  ( .D(n398), .CLK(clk), .Q(adk_out[64]) );
  DFFX1_HVT \cipher_text_reg[64]  ( .D(n270), .CLK(clk), .Q(cipher_text[64])
         );
  DFFX1_HVT \adk_out_reg[65]  ( .D(n397), .CLK(clk), .Q(adk_out[65]) );
  DFFX1_HVT \cipher_text_reg[65]  ( .D(n269), .CLK(clk), .Q(cipher_text[65])
         );
  DFFX1_HVT \adk_out_reg[66]  ( .D(n396), .CLK(clk), .Q(adk_out[66]) );
  DFFX1_HVT \cipher_text_reg[66]  ( .D(n268), .CLK(clk), .Q(cipher_text[66])
         );
  DFFX1_HVT \adk_out_reg[67]  ( .D(n395), .CLK(clk), .Q(n1177) );
  DFFX1_HVT \cipher_text_reg[67]  ( .D(n267), .CLK(clk), .Q(cipher_text[67])
         );
  DFFX1_HVT \adk_out_reg[68]  ( .D(n394), .CLK(clk), .Q(adk_out[68]), .QN(n997) );
  DFFX1_HVT \cipher_text_reg[68]  ( .D(n266), .CLK(clk), .Q(cipher_text[68])
         );
  DFFX1_HVT \adk_out_reg[69]  ( .D(n393), .CLK(clk), .Q(adk_out[69]) );
  DFFX1_HVT \cipher_text_reg[69]  ( .D(n265), .CLK(clk), .Q(cipher_text[69])
         );
  DFFX1_HVT \adk_out_reg[70]  ( .D(n392), .CLK(clk), .Q(adk_out[70]) );
  DFFX1_HVT \cipher_text_reg[70]  ( .D(n264), .CLK(clk), .Q(cipher_text[70])
         );
  DFFX1_HVT \adk_out_reg[71]  ( .D(n391), .CLK(clk), .Q(adk_out[71]) );
  DFFX1_HVT \cipher_text_reg[71]  ( .D(n263), .CLK(clk), .Q(cipher_text[71])
         );
  DFFX1_HVT \adk_out_reg[72]  ( .D(n390), .CLK(clk), .Q(adk_out[72]), .QN(n155) );
  DFFX1_HVT \cipher_text_reg[72]  ( .D(n262), .CLK(clk), .Q(cipher_text[72])
         );
  DFFX1_HVT \adk_out_reg[73]  ( .D(n389), .CLK(clk), .Q(adk_out[73]) );
  DFFX1_HVT \cipher_text_reg[73]  ( .D(n261), .CLK(clk), .Q(cipher_text[73])
         );
  DFFX1_HVT \adk_out_reg[74]  ( .D(n388), .CLK(clk), .Q(adk_out[74]) );
  DFFX1_HVT \cipher_text_reg[74]  ( .D(n260), .CLK(clk), .Q(cipher_text[74])
         );
  DFFX1_HVT \adk_out_reg[75]  ( .D(n387), .CLK(clk), .Q(n1188) );
  DFFX1_HVT \cipher_text_reg[75]  ( .D(n259), .CLK(clk), .Q(cipher_text[75])
         );
  DFFX1_HVT \adk_out_reg[76]  ( .D(n386), .CLK(clk), .Q(adk_out[76]), .QN(n690) );
  DFFX1_HVT \cipher_text_reg[76]  ( .D(n258), .CLK(clk), .Q(cipher_text[76])
         );
  DFFX1_HVT \adk_out_reg[77]  ( .D(n385), .CLK(clk), .Q(adk_out[77]) );
  DFFX1_HVT \cipher_text_reg[77]  ( .D(n257), .CLK(clk), .Q(cipher_text[77])
         );
  DFFX1_HVT \adk_out_reg[78]  ( .D(n384), .CLK(clk), .Q(adk_out[78]), .QN(n699) );
  DFFX1_HVT \cipher_text_reg[78]  ( .D(n256), .CLK(clk), .Q(cipher_text[78])
         );
  DFFX1_HVT \cipher_text_reg[79]  ( .D(n255), .CLK(clk), .Q(cipher_text[79])
         );
  DFFX1_HVT \adk_out_reg[80]  ( .D(n382), .CLK(clk), .Q(adk_out[80]), .QN(n789) );
  DFFX1_HVT \cipher_text_reg[80]  ( .D(n254), .CLK(clk), .Q(cipher_text[80])
         );
  DFFX1_HVT \adk_out_reg[81]  ( .D(n381), .CLK(clk), .Q(adk_out[81]) );
  DFFX1_HVT \cipher_text_reg[81]  ( .D(n253), .CLK(clk), .Q(cipher_text[81])
         );
  DFFX1_HVT \adk_out_reg[82]  ( .D(n380), .CLK(clk), .Q(adk_out[82]) );
  DFFX1_HVT \cipher_text_reg[82]  ( .D(n252), .CLK(clk), .Q(cipher_text[82])
         );
  DFFX1_HVT \adk_out_reg[83]  ( .D(n379), .CLK(clk), .Q(adk_out[83]) );
  DFFX1_HVT \cipher_text_reg[83]  ( .D(n251), .CLK(clk), .Q(cipher_text[83])
         );
  DFFX1_HVT \adk_out_reg[84]  ( .D(n378), .CLK(clk), .Q(adk_out[84]), .QN(n995) );
  DFFX1_HVT \cipher_text_reg[84]  ( .D(n250), .CLK(clk), .Q(cipher_text[84])
         );
  DFFX1_HVT \adk_out_reg[85]  ( .D(n377), .CLK(clk), .Q(adk_out[85]) );
  DFFX1_HVT \cipher_text_reg[85]  ( .D(n249), .CLK(clk), .Q(cipher_text[85])
         );
  DFFX1_HVT \adk_out_reg[86]  ( .D(n376), .CLK(clk), .Q(adk_out[86]) );
  DFFX1_HVT \cipher_text_reg[86]  ( .D(n248), .CLK(clk), .Q(cipher_text[86])
         );
  DFFX1_HVT \adk_out_reg[87]  ( .D(n375), .CLK(clk), .Q(adk_out[87]) );
  DFFX1_HVT \cipher_text_reg[87]  ( .D(n247), .CLK(clk), .Q(cipher_text[87])
         );
  DFFX1_HVT \adk_out_reg[88]  ( .D(n374), .CLK(clk), .Q(adk_out[88]) );
  DFFX1_HVT \cipher_text_reg[88]  ( .D(n246), .CLK(clk), .Q(cipher_text[88])
         );
  DFFX1_HVT \adk_out_reg[89]  ( .D(n373), .CLK(clk), .Q(adk_out[89]) );
  DFFX1_HVT \cipher_text_reg[89]  ( .D(n245), .CLK(clk), .Q(cipher_text[89])
         );
  DFFX1_HVT \adk_out_reg[90]  ( .D(n372), .CLK(clk), .Q(adk_out[90]) );
  DFFX1_HVT \cipher_text_reg[90]  ( .D(n244), .CLK(clk), .Q(cipher_text[90])
         );
  DFFX1_HVT \adk_out_reg[91]  ( .D(n371), .CLK(clk), .Q(adk_out[91]), .QN(n649) );
  DFFX1_HVT \cipher_text_reg[91]  ( .D(n243), .CLK(clk), .Q(cipher_text[91])
         );
  DFFX1_HVT \adk_out_reg[92]  ( .D(n370), .CLK(clk), .Q(adk_out[92]), .QN(n787) );
  DFFX1_HVT \cipher_text_reg[92]  ( .D(n242), .CLK(clk), .Q(cipher_text[92])
         );
  DFFX1_HVT \adk_out_reg[93]  ( .D(n369), .CLK(clk), .Q(adk_out[93]) );
  DFFX1_HVT \cipher_text_reg[93]  ( .D(n241), .CLK(clk), .Q(cipher_text[93])
         );
  DFFX1_HVT \adk_out_reg[94]  ( .D(n368), .CLK(clk), .Q(adk_out[94]) );
  DFFX1_HVT \cipher_text_reg[94]  ( .D(n240), .CLK(clk), .Q(cipher_text[94])
         );
  DFFX1_HVT \adk_out_reg[95]  ( .D(n367), .CLK(clk), .Q(adk_out[95]) );
  DFFX1_HVT \cipher_text_reg[95]  ( .D(n239), .CLK(clk), .Q(cipher_text[95])
         );
  DFFX1_HVT \adk_out_reg[96]  ( .D(n366), .CLK(clk), .Q(adk_out[96]), .QN(n944) );
  DFFX1_HVT \cipher_text_reg[96]  ( .D(n238), .CLK(clk), .Q(cipher_text[96])
         );
  DFFX1_HVT \adk_out_reg[97]  ( .D(n365), .CLK(clk), .Q(adk_out[97]) );
  DFFX1_HVT \cipher_text_reg[97]  ( .D(n237), .CLK(clk), .Q(cipher_text[97])
         );
  DFFX1_HVT \adk_out_reg[98]  ( .D(n364), .CLK(clk), .Q(adk_out[98]) );
  DFFX1_HVT \cipher_text_reg[98]  ( .D(n236), .CLK(clk), .Q(cipher_text[98])
         );
  DFFX1_HVT \adk_out_reg[99]  ( .D(n363), .CLK(clk), .Q(adk_out[99]) );
  DFFX1_HVT \cipher_text_reg[99]  ( .D(n235), .CLK(clk), .Q(cipher_text[99])
         );
  DFFX1_HVT \adk_out_reg[100]  ( .D(n362), .CLK(clk), .Q(adk_out[100]), .QN(
        n897) );
  DFFX1_HVT \cipher_text_reg[100]  ( .D(n234), .CLK(clk), .Q(cipher_text[100])
         );
  DFFX1_HVT \adk_out_reg[101]  ( .D(n361), .CLK(clk), .Q(adk_out[101]) );
  DFFX1_HVT \cipher_text_reg[101]  ( .D(n233), .CLK(clk), .Q(cipher_text[101])
         );
  DFFX1_HVT \adk_out_reg[102]  ( .D(n360), .CLK(clk), .Q(adk_out[102]) );
  DFFX1_HVT \cipher_text_reg[102]  ( .D(n232), .CLK(clk), .Q(cipher_text[102])
         );
  DFFX1_HVT \adk_out_reg[103]  ( .D(n359), .CLK(clk), .Q(adk_out[103]), .QN(
        n1032) );
  DFFX1_HVT \cipher_text_reg[103]  ( .D(n231), .CLK(clk), .Q(cipher_text[103])
         );
  DFFX1_HVT \adk_out_reg[104]  ( .D(n358), .CLK(clk), .Q(adk_out[104]), .QN(
        n939) );
  DFFX1_HVT \cipher_text_reg[104]  ( .D(n230), .CLK(clk), .Q(cipher_text[104])
         );
  DFFX1_HVT \adk_out_reg[105]  ( .D(n357), .CLK(clk), .Q(adk_out[105]) );
  DFFX1_HVT \cipher_text_reg[105]  ( .D(n229), .CLK(clk), .Q(cipher_text[105])
         );
  DFFX1_HVT \adk_out_reg[106]  ( .D(n356), .CLK(clk), .Q(adk_out[106]) );
  DFFX1_HVT \cipher_text_reg[106]  ( .D(n228), .CLK(clk), .Q(cipher_text[106])
         );
  DFFX1_HVT \adk_out_reg[107]  ( .D(n355), .CLK(clk), .Q(n1184), .QN(n692) );
  DFFX1_HVT \cipher_text_reg[107]  ( .D(n227), .CLK(clk), .Q(cipher_text[107])
         );
  DFFX1_HVT \adk_out_reg[108]  ( .D(n354), .CLK(clk), .Q(adk_out[108]), .QN(
        n845) );
  DFFX1_HVT \cipher_text_reg[108]  ( .D(n226), .CLK(clk), .Q(cipher_text[108])
         );
  DFFX1_HVT \adk_out_reg[109]  ( .D(n353), .CLK(clk), .Q(adk_out[109]) );
  DFFX1_HVT \cipher_text_reg[109]  ( .D(n225), .CLK(clk), .Q(cipher_text[109])
         );
  DFFX1_HVT \adk_out_reg[110]  ( .D(n352), .CLK(clk), .Q(adk_out[110]), .QN(
        n697) );
  DFFX1_HVT \cipher_text_reg[110]  ( .D(n224), .CLK(clk), .Q(cipher_text[110])
         );
  DFFX1_HVT \adk_out_reg[111]  ( .D(n351), .CLK(clk), .Q(adk_out[111]) );
  DFFX1_HVT \cipher_text_reg[111]  ( .D(n223), .CLK(clk), .Q(cipher_text[111])
         );
  DFFX1_HVT \adk_out_reg[112]  ( .D(n350), .CLK(clk), .Q(adk_out[112]), .QN(
        n893) );
  DFFX1_HVT \cipher_text_reg[112]  ( .D(n222), .CLK(clk), .Q(cipher_text[112])
         );
  DFFX1_HVT \adk_out_reg[113]  ( .D(n349), .CLK(clk), .Q(adk_out[113]) );
  DFFX1_HVT \cipher_text_reg[113]  ( .D(n221), .CLK(clk), .Q(cipher_text[113])
         );
  DFFX1_HVT \adk_out_reg[114]  ( .D(n348), .CLK(clk), .Q(adk_out[114]) );
  DFFX1_HVT \cipher_text_reg[114]  ( .D(n220), .CLK(clk), .Q(cipher_text[114])
         );
  DFFX1_HVT \adk_out_reg[115]  ( .D(n347), .CLK(clk), .Q(adk_out[115]), .QN(
        n1106) );
  DFFX1_HVT \cipher_text_reg[115]  ( .D(n219), .CLK(clk), .Q(cipher_text[115])
         );
  DFFX1_HVT \adk_out_reg[116]  ( .D(n346), .CLK(clk), .Q(adk_out[116]) );
  DFFX1_HVT \cipher_text_reg[116]  ( .D(n218), .CLK(clk), .Q(cipher_text[116])
         );
  DFFX1_HVT \adk_out_reg[117]  ( .D(n345), .CLK(clk), .Q(adk_out[117]) );
  DFFX1_HVT \cipher_text_reg[117]  ( .D(n217), .CLK(clk), .Q(cipher_text[117])
         );
  DFFX1_HVT \adk_out_reg[118]  ( .D(n344), .CLK(clk), .Q(adk_out[118]) );
  DFFX1_HVT \cipher_text_reg[118]  ( .D(n216), .CLK(clk), .Q(cipher_text[118])
         );
  DFFX1_HVT \cipher_text_reg[119]  ( .D(n215), .CLK(clk), .Q(cipher_text[119])
         );
  DFFX1_HVT \adk_out_reg[120]  ( .D(n342), .CLK(clk), .Q(adk_out[120]), .QN(
        n915) );
  DFFX1_HVT \cipher_text_reg[120]  ( .D(n214), .CLK(clk), .Q(cipher_text[120])
         );
  DFFX1_HVT \adk_out_reg[121]  ( .D(n341), .CLK(clk), .Q(adk_out[121]) );
  DFFX1_HVT \cipher_text_reg[121]  ( .D(n213), .CLK(clk), .Q(cipher_text[121])
         );
  DFFX1_HVT \adk_out_reg[122]  ( .D(n340), .CLK(clk), .Q(adk_out[122]) );
  DFFX1_HVT \cipher_text_reg[122]  ( .D(n212), .CLK(clk), .Q(cipher_text[122])
         );
  DFFX1_HVT \adk_out_reg[123]  ( .D(n339), .CLK(clk), .Q(adk_out[123]) );
  DFFX1_HVT \cipher_text_reg[123]  ( .D(n211), .CLK(clk), .Q(cipher_text[123])
         );
  DFFX1_HVT \adk_out_reg[124]  ( .D(n338), .CLK(clk), .Q(adk_out[124]), .QN(
        n1024) );
  DFFX1_HVT \cipher_text_reg[124]  ( .D(n210), .CLK(clk), .Q(cipher_text[124])
         );
  DFFX1_HVT \adk_out_reg[125]  ( .D(n337), .CLK(clk), .Q(adk_out[125]) );
  DFFX1_HVT \cipher_text_reg[125]  ( .D(n209), .CLK(clk), .Q(cipher_text[125])
         );
  DFFX1_HVT \adk_out_reg[126]  ( .D(n336), .CLK(clk), .Q(adk_out[126]) );
  DFFX1_HVT \cipher_text_reg[126]  ( .D(n208), .CLK(clk), .Q(cipher_text[126])
         );
  DFFX1_HVT \cipher_text_reg[127]  ( .D(n964), .CLK(clk), .Q(cipher_text[127]), 
        .QN(n1053) );
  AO22X1_HVT U144 ( .A1(cipher_text[126]), .A2(n1048), .A3(out1[126]), .A4(
        n1297), .Y(n208) );
  AO22X1_HVT U145 ( .A1(cipher_text[125]), .A2(n1328), .A3(out1[125]), .A4(
        n1296), .Y(n209) );
  AO22X1_HVT U146 ( .A1(cipher_text[124]), .A2(n1046), .A3(out1[124]), .A4(
        n1295), .Y(n210) );
  AO22X1_HVT U147 ( .A1(cipher_text[123]), .A2(n708), .A3(out1[123]), .A4(
        n1294), .Y(n211) );
  AO22X1_HVT U148 ( .A1(cipher_text[122]), .A2(n818), .A3(out1[122]), .A4(
        n1293), .Y(n212) );
  AO22X1_HVT U149 ( .A1(cipher_text[121]), .A2(n1336), .A3(out1[121]), .A4(
        n1292), .Y(n213) );
  AO22X1_HVT U150 ( .A1(cipher_text[120]), .A2(n704), .A3(out1[120]), .A4(
        n1291), .Y(n214) );
  AO22X1_HVT U151 ( .A1(cipher_text[119]), .A2(n1048), .A3(out1[119]), .A4(
        n1296), .Y(n215) );
  AO22X1_HVT U152 ( .A1(cipher_text[118]), .A2(n1332), .A3(out1[118]), .A4(
        n1295), .Y(n216) );
  AO22X1_HVT U153 ( .A1(cipher_text[117]), .A2(n707), .A3(out1[117]), .A4(
        n1294), .Y(n217) );
  AO22X1_HVT U154 ( .A1(cipher_text[116]), .A2(n1336), .A3(out1[116]), .A4(
        n1293), .Y(n218) );
  AO22X1_HVT U155 ( .A1(cipher_text[115]), .A2(n1045), .A3(out1[115]), .A4(
        n1292), .Y(n219) );
  AO22X1_HVT U156 ( .A1(cipher_text[114]), .A2(n704), .A3(out1[114]), .A4(
        n1291), .Y(n220) );
  AO22X1_HVT U157 ( .A1(cipher_text[113]), .A2(n704), .A3(out1[113]), .A4(
        n1302), .Y(n221) );
  AO22X1_HVT U158 ( .A1(cipher_text[112]), .A2(n1046), .A3(out1[112]), .A4(
        n1301), .Y(n222) );
  AO22X1_HVT U159 ( .A1(cipher_text[111]), .A2(n1327), .A3(out1[111]), .A4(
        n1300), .Y(n223) );
  AO22X1_HVT U160 ( .A1(cipher_text[110]), .A2(n1045), .A3(out1[110]), .A4(
        n1299), .Y(n224) );
  AO22X1_HVT U161 ( .A1(cipher_text[109]), .A2(n1047), .A3(out1[109]), .A4(
        n1298), .Y(n225) );
  AO22X1_HVT U162 ( .A1(cipher_text[108]), .A2(n705), .A3(out1[108]), .A4(
        n1297), .Y(n226) );
  AO22X1_HVT U163 ( .A1(cipher_text[107]), .A2(n1048), .A3(out1[107]), .A4(
        n1298), .Y(n227) );
  AO22X1_HVT U164 ( .A1(cipher_text[106]), .A2(n707), .A3(out1[106]), .A4(
        n1297), .Y(n228) );
  AO22X1_HVT U165 ( .A1(cipher_text[105]), .A2(n1327), .A3(out1[105]), .A4(
        n1296), .Y(n229) );
  AO22X1_HVT U166 ( .A1(cipher_text[104]), .A2(n1330), .A3(out1[104]), .A4(
        n1295), .Y(n230) );
  AO22X1_HVT U167 ( .A1(cipher_text[103]), .A2(n818), .A3(out1[103]), .A4(
        n1317), .Y(n231) );
  AO22X1_HVT U168 ( .A1(cipher_text[102]), .A2(n1328), .A3(out1[102]), .A4(
        n1316), .Y(n232) );
  AO22X1_HVT U169 ( .A1(cipher_text[101]), .A2(n705), .A3(out1[101]), .A4(
        n1315), .Y(n233) );
  AO22X1_HVT U170 ( .A1(cipher_text[100]), .A2(n1332), .A3(out1[100]), .A4(
        n1314), .Y(n234) );
  AO22X1_HVT U171 ( .A1(cipher_text[99]), .A2(n708), .A3(out1[99]), .A4(n1313), 
        .Y(n235) );
  AO22X1_HVT U172 ( .A1(cipher_text[98]), .A2(n1045), .A3(out1[98]), .A4(n1312), .Y(n236) );
  AO22X1_HVT U173 ( .A1(cipher_text[97]), .A2(n819), .A3(out1[97]), .A4(n1310), 
        .Y(n237) );
  AO22X1_HVT U174 ( .A1(cipher_text[96]), .A2(n1328), .A3(out1[96]), .A4(n1309), .Y(n238) );
  AO22X1_HVT U175 ( .A1(cipher_text[95]), .A2(n1329), .A3(out1[95]), .A4(n1317), .Y(n239) );
  AO22X1_HVT U176 ( .A1(cipher_text[94]), .A2(n708), .A3(out1[94]), .A4(n1316), 
        .Y(n240) );
  AO22X1_HVT U177 ( .A1(cipher_text[93]), .A2(n1332), .A3(out1[93]), .A4(n1315), .Y(n241) );
  AO22X1_HVT U178 ( .A1(cipher_text[92]), .A2(n818), .A3(out1[92]), .A4(n1314), 
        .Y(n242) );
  AO22X1_HVT U179 ( .A1(cipher_text[91]), .A2(n1336), .A3(out1[91]), .A4(n1313), .Y(n243) );
  AO22X1_HVT U180 ( .A1(cipher_text[90]), .A2(n705), .A3(out1[90]), .A4(n1312), 
        .Y(n244) );
  AO22X1_HVT U181 ( .A1(cipher_text[89]), .A2(n1329), .A3(out1[89]), .A4(n1296), .Y(n245) );
  AO22X1_HVT U182 ( .A1(cipher_text[88]), .A2(n1327), .A3(out1[88]), .A4(n1295), .Y(n246) );
  AO22X1_HVT U183 ( .A1(cipher_text[87]), .A2(n1046), .A3(out1[87]), .A4(n1294), .Y(n247) );
  AO22X1_HVT U184 ( .A1(cipher_text[86]), .A2(n819), .A3(out1[86]), .A4(n1293), 
        .Y(n248) );
  AO22X1_HVT U185 ( .A1(cipher_text[85]), .A2(n1330), .A3(out1[85]), .A4(n1292), .Y(n249) );
  AO22X1_HVT U186 ( .A1(cipher_text[84]), .A2(n1329), .A3(out1[84]), .A4(n1291), .Y(n250) );
  AO22X1_HVT U187 ( .A1(cipher_text[83]), .A2(n704), .A3(out1[83]), .A4(n1294), 
        .Y(n251) );
  AO22X1_HVT U188 ( .A1(cipher_text[82]), .A2(n707), .A3(out1[82]), .A4(n1293), 
        .Y(n252) );
  AO22X1_HVT U189 ( .A1(cipher_text[81]), .A2(n707), .A3(out1[81]), .A4(n1292), 
        .Y(n253) );
  AO22X1_HVT U190 ( .A1(cipher_text[80]), .A2(n1047), .A3(out1[80]), .A4(n1291), .Y(n254) );
  AO22X1_HVT U191 ( .A1(cipher_text[79]), .A2(n1047), .A3(out1[79]), .A4(n1308), .Y(n255) );
  AO22X1_HVT U192 ( .A1(cipher_text[78]), .A2(n1329), .A3(out1[78]), .A4(n1307), .Y(n256) );
  AO22X1_HVT U195 ( .A1(cipher_text[75]), .A2(n1335), .A3(out1[75]), .A4(n1302), .Y(n259) );
  AO22X1_HVT U196 ( .A1(cipher_text[74]), .A2(n708), .A3(out1[74]), .A4(n1301), 
        .Y(n260) );
  AO22X1_HVT U197 ( .A1(cipher_text[73]), .A2(n708), .A3(out1[73]), .A4(n1300), 
        .Y(n261) );
  AO22X1_HVT U198 ( .A1(cipher_text[72]), .A2(n1047), .A3(out1[72]), .A4(n1299), .Y(n262) );
  AO22X1_HVT U199 ( .A1(cipher_text[71]), .A2(n1335), .A3(out1[71]), .A4(n1310), .Y(n263) );
  AO22X1_HVT U200 ( .A1(cipher_text[70]), .A2(n1045), .A3(out1[70]), .A4(n1309), .Y(n264) );
  AO22X1_HVT U201 ( .A1(cipher_text[69]), .A2(n1045), .A3(out1[69]), .A4(n1308), .Y(n265) );
  AO22X1_HVT U202 ( .A1(cipher_text[68]), .A2(n835), .A3(out1[68]), .A4(n1307), 
        .Y(n266) );
  AO22X1_HVT U203 ( .A1(cipher_text[67]), .A2(n819), .A3(out1[67]), .A4(n1317), 
        .Y(n267) );
  AO22X1_HVT U204 ( .A1(cipher_text[66]), .A2(n1048), .A3(out1[66]), .A4(n1316), .Y(n268) );
  AO22X1_HVT U205 ( .A1(cipher_text[65]), .A2(n1334), .A3(out1[65]), .A4(n1315), .Y(n269) );
  AO22X1_HVT U206 ( .A1(cipher_text[64]), .A2(n819), .A3(out1[64]), .A4(n1314), 
        .Y(n270) );
  AO22X1_HVT U207 ( .A1(cipher_text[63]), .A2(n1336), .A3(out1[63]), .A4(n1317), .Y(n271) );
  AO22X1_HVT U208 ( .A1(cipher_text[62]), .A2(n1331), .A3(out1[62]), .A4(n1316), .Y(n272) );
  AO22X1_HVT U209 ( .A1(cipher_text[61]), .A2(n1331), .A3(out1[61]), .A4(n1315), .Y(n273) );
  AO22X1_HVT U210 ( .A1(cipher_text[60]), .A2(n818), .A3(out1[60]), .A4(n1314), 
        .Y(n274) );
  AO22X1_HVT U211 ( .A1(cipher_text[59]), .A2(n1335), .A3(out1[59]), .A4(n1313), .Y(n275) );
  AO22X1_HVT U212 ( .A1(cipher_text[58]), .A2(n835), .A3(out1[58]), .A4(n1312), 
        .Y(n276) );
  AO22X1_HVT U213 ( .A1(cipher_text[57]), .A2(n705), .A3(out1[57]), .A4(n1310), 
        .Y(n277) );
  AO22X1_HVT U214 ( .A1(cipher_text[56]), .A2(n1330), .A3(out1[56]), .A4(n1309), .Y(n278) );
  AO22X1_HVT U215 ( .A1(cipher_text[55]), .A2(n1333), .A3(out1[55]), .A4(n1302), .Y(n279) );
  AO22X1_HVT U216 ( .A1(cipher_text[54]), .A2(n1046), .A3(out1[54]), .A4(n1301), .Y(n280) );
  AO22X1_HVT U217 ( .A1(cipher_text[53]), .A2(n1047), .A3(n1300), .A4(out1[53]), .Y(n281) );
  AO22X1_HVT U218 ( .A1(cipher_text[52]), .A2(n1048), .A3(out1[52]), .A4(n1299), .Y(n282) );
  AO22X1_HVT U219 ( .A1(cipher_text[51]), .A2(n1336), .A3(out1[51]), .A4(n1298), .Y(n283) );
  AO22X1_HVT U220 ( .A1(cipher_text[50]), .A2(n1334), .A3(out1[50]), .A4(n1297), .Y(n284) );
  AO22X1_HVT U221 ( .A1(cipher_text[49]), .A2(n1335), .A3(out1[49]), .A4(n1310), .Y(n285) );
  AO22X1_HVT U222 ( .A1(cipher_text[48]), .A2(n1331), .A3(out1[48]), .A4(n1309), .Y(n286) );
  AO22X1_HVT U223 ( .A1(cipher_text[47]), .A2(n1047), .A3(out1[47]), .A4(n1308), .Y(n287) );
  AO22X1_HVT U224 ( .A1(cipher_text[46]), .A2(n1330), .A3(out1[46]), .A4(n1307), .Y(n288) );
  AO22X1_HVT U225 ( .A1(cipher_text[45]), .A2(n705), .A3(out1[45]), .A4(n1306), 
        .Y(n289) );
  AO22X1_HVT U226 ( .A1(cipher_text[44]), .A2(n1334), .A3(out1[44]), .A4(n1305), .Y(n290) );
  AO22X1_HVT U227 ( .A1(cipher_text[43]), .A2(n1333), .A3(out1[43]), .A4(n1313), .Y(n291) );
  AO22X1_HVT U228 ( .A1(cipher_text[42]), .A2(n1331), .A3(out1[42]), .A4(n1312), .Y(n292) );
  AO22X1_HVT U229 ( .A1(cipher_text[41]), .A2(n1330), .A3(out1[41]), .A4(n1310), .Y(n293) );
  AO22X1_HVT U230 ( .A1(cipher_text[40]), .A2(n1332), .A3(out1[40]), .A4(n1309), .Y(n294) );
  AO22X1_HVT U231 ( .A1(cipher_text[39]), .A2(n818), .A3(out1[39]), .A4(n1308), 
        .Y(n295) );
  AO22X1_HVT U232 ( .A1(cipher_text[38]), .A2(n1333), .A3(out1[38]), .A4(n1307), .Y(n296) );
  AO22X1_HVT U233 ( .A1(cipher_text[37]), .A2(n1046), .A3(out1[37]), .A4(n1306), .Y(n297) );
  AO22X1_HVT U234 ( .A1(cipher_text[36]), .A2(n835), .A3(out1[36]), .A4(n1305), 
        .Y(n298) );
  AO22X1_HVT U235 ( .A1(cipher_text[35]), .A2(n1328), .A3(out1[35]), .A4(n1302), .Y(n299) );
  AO22X1_HVT U236 ( .A1(cipher_text[34]), .A2(n1335), .A3(out1[34]), .A4(n1301), .Y(n300) );
  AO22X1_HVT U237 ( .A1(cipher_text[33]), .A2(n1332), .A3(out1[33]), .A4(n1300), .Y(n301) );
  AO22X1_HVT U238 ( .A1(cipher_text[32]), .A2(n818), .A3(out1[32]), .A4(n1299), 
        .Y(n302) );
  AO22X1_HVT U239 ( .A1(cipher_text[31]), .A2(n835), .A3(out1[31]), .A4(n1296), 
        .Y(n303) );
  AO22X1_HVT U240 ( .A1(cipher_text[30]), .A2(n835), .A3(out1[30]), .A4(n1295), 
        .Y(n304) );
  AO22X1_HVT U241 ( .A1(cipher_text[29]), .A2(n1045), .A3(out1[29]), .A4(n1294), .Y(n305) );
  AO22X1_HVT U242 ( .A1(cipher_text[28]), .A2(n1333), .A3(out1[28]), .A4(n1293), .Y(n306) );
  AO22X1_HVT U243 ( .A1(cipher_text[27]), .A2(n1333), .A3(out1[27]), .A4(n1292), .Y(n307) );
  AO22X1_HVT U244 ( .A1(cipher_text[26]), .A2(n1334), .A3(out1[26]), .A4(n1291), .Y(n308) );
  AO22X1_HVT U245 ( .A1(cipher_text[25]), .A2(n1334), .A3(out1[25]), .A4(n1302), .Y(n309) );
  AO22X1_HVT U246 ( .A1(cipher_text[24]), .A2(n819), .A3(out1[24]), .A4(n1301), 
        .Y(n310) );
  AO22X1_HVT U247 ( .A1(cipher_text[23]), .A2(n1327), .A3(out1[23]), .A4(n1300), .Y(n311) );
  AO22X1_HVT U248 ( .A1(cipher_text[22]), .A2(n835), .A3(out1[22]), .A4(n1299), 
        .Y(n312) );
  AO22X1_HVT U249 ( .A1(cipher_text[21]), .A2(n1045), .A3(out1[21]), .A4(n1298), .Y(n313) );
  AO22X1_HVT U250 ( .A1(cipher_text[20]), .A2(n818), .A3(out1[20]), .A4(n1297), 
        .Y(n314) );
  AO22X1_HVT U251 ( .A1(cipher_text[19]), .A2(n1333), .A3(out1[19]), .A4(n1308), .Y(n315) );
  AO22X1_HVT U252 ( .A1(cipher_text[18]), .A2(n1329), .A3(out1[18]), .A4(n1307), .Y(n316) );
  AO22X1_HVT U253 ( .A1(cipher_text[17]), .A2(n1335), .A3(out1[17]), .A4(n1306), .Y(n317) );
  AO22X1_HVT U254 ( .A1(cipher_text[16]), .A2(n1335), .A3(n1305), .A4(out1[16]), .Y(n318) );
  AO22X1_HVT U255 ( .A1(cipher_text[15]), .A2(n1328), .A3(out1[15]), .A4(n1298), .Y(n319) );
  AO22X1_HVT U256 ( .A1(cipher_text[14]), .A2(n704), .A3(out1[14]), .A4(n1297), 
        .Y(n320) );
  AO22X1_HVT U257 ( .A1(cipher_text[13]), .A2(n1331), .A3(out1[13]), .A4(n1296), .Y(n321) );
  AO22X1_HVT U258 ( .A1(cipher_text[12]), .A2(n1334), .A3(out1[12]), .A4(n1295), .Y(n322) );
  AO22X1_HVT U259 ( .A1(cipher_text[11]), .A2(n835), .A3(out1[11]), .A4(n1294), 
        .Y(n323) );
  AO22X1_HVT U260 ( .A1(cipher_text[10]), .A2(n1327), .A3(out1[10]), .A4(n1293), .Y(n324) );
  AO22X1_HVT U261 ( .A1(cipher_text[9]), .A2(n1331), .A3(out1[9]), .A4(n1292), 
        .Y(n325) );
  AO22X1_HVT U262 ( .A1(cipher_text[8]), .A2(n1336), .A3(out1[8]), .A4(n1291), 
        .Y(n326) );
  AO22X1_HVT U263 ( .A1(cipher_text[7]), .A2(n1047), .A3(out1[7]), .A4(n1306), 
        .Y(n327) );
  AO22X1_HVT U264 ( .A1(cipher_text[6]), .A2(n1330), .A3(out1[6]), .A4(n1305), 
        .Y(n328) );
  AO22X1_HVT U265 ( .A1(cipher_text[5]), .A2(n1333), .A3(out1[5]), .A4(n1317), 
        .Y(n329) );
  AO22X1_HVT U266 ( .A1(cipher_text[4]), .A2(n819), .A3(out1[4]), .A4(n1316), 
        .Y(n330) );
  AO22X1_HVT U267 ( .A1(cipher_text[3]), .A2(n1331), .A3(out1[3]), .A4(n1315), 
        .Y(n331) );
  AO22X1_HVT U268 ( .A1(cipher_text[2]), .A2(n707), .A3(out1[2]), .A4(n1314), 
        .Y(n332) );
  AO22X1_HVT U269 ( .A1(cipher_text[1]), .A2(n1329), .A3(out1[1]), .A4(n1313), 
        .Y(n333) );
  AO22X1_HVT U270 ( .A1(cipher_text[0]), .A2(n1330), .A3(out1[0]), .A4(n1312), 
        .Y(n334) );
  AND2X1_HVT U271 ( .A1(n999), .A2(n8), .Y(n19) );
  AO222X1_HVT U277 ( .A1(n1229), .A2(n29), .A3(n1270), .A4(out1[122]), .A5(
        adk_out[122]), .A6(n1323), .Y(n340) );
  AO222X1_HVT U285 ( .A1(n1214), .A2(n37), .A3(n1276), .A4(out1[114]), .A5(
        adk_out[114]), .A6(n677), .Y(n348) );
  AO222X1_HVT U295 ( .A1(n1228), .A2(n47), .A3(n1270), .A4(out1[104]), .A5(
        n940), .A6(n1349), .Y(n358) );
  AO222X1_HVT U296 ( .A1(n1227), .A2(n48), .A3(n1270), .A4(out1[103]), .A5(
        n1033), .A6(n1350), .Y(n359) );
  AO222X1_HVT U303 ( .A1(n1214), .A2(n55), .A3(n1259), .A4(out1[96]), .A5(n945), .A6(n1349), .Y(n366) );
  AO222X1_HVT U304 ( .A1(n1230), .A2(n56), .A3(n1276), .A4(out1[95]), .A5(
        adk_out[95]), .A6(n1240), .Y(n367) );
  AO222X1_HVT U310 ( .A1(n1215), .A2(n62), .A3(n1257), .A4(out1[89]), .A5(
        adk_out[89]), .A6(n1345), .Y(n373) );
  AO222X1_HVT U311 ( .A1(n1214), .A2(n63), .A3(n1258), .A4(out1[88]), .A5(
        adk_out[88]), .A6(n1353), .Y(n374) );
  AO222X1_HVT U312 ( .A1(n1215), .A2(n64), .A3(n1254), .A4(out1[87]), .A5(
        adk_out[87]), .A6(n1348), .Y(n375) );
  AO222X1_HVT U319 ( .A1(n1223), .A2(n71), .A3(n1256), .A4(out1[80]), .A5(n790), .A6(n678), .Y(n382) );
  AO222X1_HVT U321 ( .A1(n1229), .A2(n73), .A3(n1256), .A4(out1[78]), .A5(n700), .A6(n1240), .Y(n384) );
  AO222X1_HVT U326 ( .A1(n1234), .A2(n78), .A3(n1253), .A4(out1[73]), .A5(
        adk_out[73]), .A6(n1323), .Y(n389) );
  AO222X1_HVT U327 ( .A1(n1233), .A2(n79), .A3(n1252), .A4(out1[72]), .A5(n207), .A6(n1237), .Y(n390) );
  AO222X1_HVT U328 ( .A1(n1230), .A2(n80), .A3(n1253), .A4(out1[71]), .A5(
        adk_out[71]), .A6(n1345), .Y(n391) );
  AO222X1_HVT U333 ( .A1(n1235), .A2(n85), .A3(out1[66]), .A4(n1261), .A5(
        adk_out[66]), .A6(n1349), .Y(n396) );
  AO222X1_HVT U335 ( .A1(n1233), .A2(n87), .A3(n1257), .A4(out1[64]), .A5(
        adk_out[64]), .A6(n658), .Y(n398) );
  AO222X1_HVT U351 ( .A1(n1216), .A2(n103), .A3(n1262), .A4(out1[48]), .A5(
        n866), .A6(n1237), .Y(n414) );
  AO222X1_HVT U367 ( .A1(n1214), .A2(n119), .A3(n1262), .A4(out1[32]), .A5(
        n905), .A6(n668), .Y(n430) );
  AO222X1_HVT U383 ( .A1(n1222), .A2(n135), .A3(out1[16]), .A4(n1275), .A5(
        n844), .A6(n1351), .Y(n446) );
  AO222X1_HVT U384 ( .A1(n1221), .A2(n136), .A3(n1269), .A4(out1[15]), .A5(
        adk_out[15]), .A6(n658), .Y(n447) );
  AO222X1_HVT U391 ( .A1(n1224), .A2(n143), .A3(n1252), .A4(out1[8]), .A5(n780), .A6(n1346), .Y(n454) );
  AO222X1_HVT U392 ( .A1(n1236), .A2(n144), .A3(n1258), .A4(out1[7]), .A5(
        n1037), .A6(n1320), .Y(n455) );
  NAND2X0_HVT U402 ( .A1(n154), .A2(n999), .Y(n24) );
  AO22X1_HVT U403 ( .A1(n793), .A2(key_round[127]), .A3(keys1[127]), .A4(n1131), .Y(n463) );
  AO22X1_HVT U405 ( .A1(n985), .A2(key_round[125]), .A3(keys1[125]), .A4(n1140), .Y(n465) );
  AO22X1_HVT U406 ( .A1(n984), .A2(key_round[124]), .A3(keys1[124]), .A4(n1164), .Y(n466) );
  AO22X1_HVT U408 ( .A1(n984), .A2(key_round[122]), .A3(keys1[122]), .A4(n1122), .Y(n468) );
  AO22X1_HVT U409 ( .A1(n1147), .A2(key_round[121]), .A3(keys1[121]), .A4(
        n1164), .Y(n469) );
  AO22X1_HVT U410 ( .A1(n799), .A2(key_round[120]), .A3(keys1[120]), .A4(n1108), .Y(n470) );
  AO22X1_HVT U411 ( .A1(n799), .A2(key_round[119]), .A3(keys1[119]), .A4(n1122), .Y(n471) );
  AO22X1_HVT U412 ( .A1(n799), .A2(key_round[118]), .A3(keys1[118]), .A4(n1118), .Y(n472) );
  AO22X1_HVT U413 ( .A1(n1152), .A2(key_round[117]), .A3(keys1[117]), .A4(
        n1119), .Y(n473) );
  AO22X1_HVT U414 ( .A1(n1145), .A2(key_round[116]), .A3(keys1[116]), .A4(
        n1118), .Y(n474) );
  AO22X1_HVT U415 ( .A1(n983), .A2(key_round[115]), .A3(keys1[115]), .A4(n1119), .Y(n475) );
  AO22X1_HVT U416 ( .A1(n1146), .A2(key_round[114]), .A3(keys1[114]), .A4(
        n1128), .Y(n476) );
  AO22X1_HVT U417 ( .A1(n1146), .A2(key_round[113]), .A3(keys1[113]), .A4(
        n1134), .Y(n477) );
  AO22X1_HVT U418 ( .A1(n1148), .A2(key_round[112]), .A3(keys1[112]), .A4(
        n1124), .Y(n478) );
  AO22X1_HVT U419 ( .A1(n1145), .A2(key_round[111]), .A3(keys1[111]), .A4(
        n1125), .Y(n479) );
  AO22X1_HVT U420 ( .A1(n1148), .A2(key_round[110]), .A3(keys1[110]), .A4(
        n1127), .Y(n480) );
  AO22X1_HVT U421 ( .A1(n1146), .A2(key_round[109]), .A3(keys1[109]), .A4(
        n1128), .Y(n481) );
  AO22X1_HVT U424 ( .A1(n982), .A2(key_round[106]), .A3(keys1[106]), .A4(n1124), .Y(n484) );
  AO22X1_HVT U425 ( .A1(n1153), .A2(key_round[105]), .A3(keys1[105]), .A4(
        n1130), .Y(n485) );
  AO22X1_HVT U426 ( .A1(n1154), .A2(key_round[104]), .A3(keys1[104]), .A4(
        n1116), .Y(n486) );
  AO22X1_HVT U427 ( .A1(n985), .A2(key_round[103]), .A3(keys1[103]), .A4(n1117), .Y(n487) );
  AO22X1_HVT U428 ( .A1(n792), .A2(key_round[102]), .A3(keys1[102]), .A4(n1118), .Y(n488) );
  AO22X1_HVT U429 ( .A1(n1146), .A2(key_round[101]), .A3(keys1[101]), .A4(
        n1119), .Y(n489) );
  AO22X1_HVT U430 ( .A1(n1144), .A2(key_round[100]), .A3(keys1[100]), .A4(
        n1121), .Y(n490) );
  AO22X1_HVT U431 ( .A1(n1145), .A2(key_round[99]), .A3(keys1[99]), .A4(n1139), 
        .Y(n491) );
  AO22X1_HVT U432 ( .A1(n1143), .A2(key_round[98]), .A3(keys1[98]), .A4(n1124), 
        .Y(n492) );
  AO22X1_HVT U433 ( .A1(n985), .A2(key_round[97]), .A3(keys1[97]), .A4(n1125), 
        .Y(n493) );
  AO22X1_HVT U434 ( .A1(n984), .A2(key_round[96]), .A3(keys1[96]), .A4(n1127), 
        .Y(n494) );
  AO22X1_HVT U435 ( .A1(n798), .A2(key_round[95]), .A3(keys1[95]), .A4(n1115), 
        .Y(n495) );
  AO22X1_HVT U436 ( .A1(n792), .A2(key_round[94]), .A3(keys1[94]), .A4(n1116), 
        .Y(n496) );
  AO22X1_HVT U437 ( .A1(n792), .A2(key_round[93]), .A3(keys1[93]), .A4(n1117), 
        .Y(n497) );
  AO22X1_HVT U438 ( .A1(n1152), .A2(key_round[92]), .A3(keys1[92]), .A4(n1110), 
        .Y(n498) );
  AO22X1_HVT U440 ( .A1(n793), .A2(key_round[90]), .A3(keys1[90]), .A4(n1111), 
        .Y(n500) );
  AO22X1_HVT U442 ( .A1(n1147), .A2(key_round[88]), .A3(keys1[88]), .A4(n1137), 
        .Y(n502) );
  AO22X1_HVT U443 ( .A1(n984), .A2(key_round[87]), .A3(keys1[87]), .A4(n1133), 
        .Y(n503) );
  AO22X1_HVT U444 ( .A1(n1148), .A2(key_round[86]), .A3(keys1[86]), .A4(n1134), 
        .Y(n504) );
  AO22X1_HVT U445 ( .A1(n983), .A2(key_round[85]), .A3(keys1[85]), .A4(n1133), 
        .Y(n505) );
  AO22X1_HVT U446 ( .A1(n1152), .A2(key_round[84]), .A3(keys1[84]), .A4(n1134), 
        .Y(n506) );
  AO22X1_HVT U447 ( .A1(n1129), .A2(key_round[83]), .A3(keys1[83]), .A4(n1127), 
        .Y(n507) );
  AO22X1_HVT U448 ( .A1(n792), .A2(key_round[82]), .A3(keys1[82]), .A4(n1164), 
        .Y(n508) );
  AO22X1_HVT U449 ( .A1(n1151), .A2(key_round[81]), .A3(keys1[81]), .A4(n1122), 
        .Y(n509) );
  AO22X1_HVT U450 ( .A1(n1146), .A2(key_round[80]), .A3(keys1[80]), .A4(n1108), 
        .Y(n510) );
  AO22X1_HVT U451 ( .A1(n1147), .A2(key_round[79]), .A3(keys1[79]), .A4(n1108), 
        .Y(n511) );
  AO22X1_HVT U452 ( .A1(n1112), .A2(key_round[78]), .A3(keys1[78]), .A4(n1127), 
        .Y(n512) );
  AO22X1_HVT U453 ( .A1(n984), .A2(key_round[77]), .A3(keys1[77]), .A4(n1128), 
        .Y(n513) );
  AO22X1_HVT U454 ( .A1(n1143), .A2(key_round[76]), .A3(keys1[76]), .A4(n1136), 
        .Y(n514) );
  AO22X1_HVT U455 ( .A1(n1143), .A2(key_round[75]), .A3(keys1[75]), .A4(n1121), 
        .Y(n515) );
  AO22X1_HVT U456 ( .A1(n793), .A2(key_round[74]), .A3(keys1[74]), .A4(n1136), 
        .Y(n516) );
  AO22X1_HVT U457 ( .A1(n1132), .A2(key_round[73]), .A3(keys1[73]), .A4(n1137), 
        .Y(n517) );
  AO22X1_HVT U458 ( .A1(n982), .A2(key_round[72]), .A3(keys1[72]), .A4(n1128), 
        .Y(n518) );
  AO22X1_HVT U459 ( .A1(n1148), .A2(key_round[71]), .A3(keys1[71]), .A4(n1117), 
        .Y(n519) );
  AO22X1_HVT U460 ( .A1(n985), .A2(key_round[70]), .A3(keys1[70]), .A4(n1127), 
        .Y(n520) );
  AO22X1_HVT U461 ( .A1(n1147), .A2(key_round[69]), .A3(keys1[69]), .A4(n1133), 
        .Y(n521) );
  AO22X1_HVT U462 ( .A1(n798), .A2(key_round[68]), .A3(keys1[68]), .A4(n1164), 
        .Y(n522) );
  AO22X1_HVT U463 ( .A1(n799), .A2(key_round[67]), .A3(keys1[67]), .A4(n1108), 
        .Y(n523) );
  AO22X1_HVT U464 ( .A1(n983), .A2(key_round[66]), .A3(keys1[66]), .A4(n1110), 
        .Y(n524) );
  AO22X1_HVT U465 ( .A1(n982), .A2(key_round[65]), .A3(keys1[65]), .A4(n1111), 
        .Y(n525) );
  AO22X1_HVT U466 ( .A1(n1154), .A2(key_round[64]), .A3(keys1[64]), .A4(n1109), 
        .Y(n526) );
  AO22X1_HVT U467 ( .A1(n1151), .A2(key_round[63]), .A3(keys1[63]), .A4(n1121), 
        .Y(n527) );
  AO22X1_HVT U468 ( .A1(n1153), .A2(key_round[62]), .A3(keys1[62]), .A4(n1118), 
        .Y(n528) );
  AO22X1_HVT U469 ( .A1(n1154), .A2(key_round[61]), .A3(keys1[61]), .A4(n1119), 
        .Y(n529) );
  AO22X1_HVT U470 ( .A1(n1145), .A2(key_round[60]), .A3(keys1[60]), .A4(n1121), 
        .Y(n530) );
  AO22X1_HVT U471 ( .A1(n1154), .A2(key_round[59]), .A3(keys1[59]), .A4(n1109), 
        .Y(n531) );
  AO22X1_HVT U472 ( .A1(n798), .A2(key_round[58]), .A3(keys1[58]), .A4(n1111), 
        .Y(n532) );
  AO22X1_HVT U473 ( .A1(n1153), .A2(key_round[57]), .A3(keys1[57]), .A4(n1110), 
        .Y(n533) );
  AO22X1_HVT U474 ( .A1(n1126), .A2(key_round[56]), .A3(keys1[56]), .A4(n1108), 
        .Y(n534) );
  AO22X1_HVT U475 ( .A1(n798), .A2(key_round[55]), .A3(keys1[55]), .A4(n1108), 
        .Y(n535) );
  AO22X1_HVT U476 ( .A1(n1151), .A2(key_round[54]), .A3(keys1[54]), .A4(n1115), 
        .Y(n536) );
  AO22X1_HVT U477 ( .A1(n1143), .A2(key_round[53]), .A3(keys1[53]), .A4(n1114), 
        .Y(n537) );
  AO22X1_HVT U478 ( .A1(n1144), .A2(key_round[52]), .A3(keys1[52]), .A4(n1134), 
        .Y(n538) );
  AO22X1_HVT U479 ( .A1(n1153), .A2(key_round[51]), .A3(keys1[51]), .A4(n1133), 
        .Y(n539) );
  AO22X1_HVT U480 ( .A1(n1153), .A2(key_round[50]), .A3(keys1[50]), .A4(n1131), 
        .Y(n540) );
  AO22X1_HVT U481 ( .A1(n798), .A2(key_round[49]), .A3(keys1[49]), .A4(n1130), 
        .Y(n541) );
  AO22X1_HVT U482 ( .A1(n982), .A2(key_round[48]), .A3(keys1[48]), .A4(n1110), 
        .Y(n542) );
  AO22X1_HVT U483 ( .A1(n793), .A2(key_round[47]), .A3(keys1[47]), .A4(n1114), 
        .Y(n543) );
  AO22X1_HVT U484 ( .A1(n1129), .A2(key_round[46]), .A3(keys1[46]), .A4(n1111), 
        .Y(n544) );
  AO22X1_HVT U485 ( .A1(n1147), .A2(key_round[45]), .A3(keys1[45]), .A4(n1110), 
        .Y(n545) );
  AO22X1_HVT U486 ( .A1(n1147), .A2(key_round[44]), .A3(keys1[44]), .A4(n1111), 
        .Y(n546) );
  AO22X1_HVT U487 ( .A1(n1148), .A2(key_round[43]), .A3(keys1[43]), .A4(n1140), 
        .Y(n547) );
  AO22X1_HVT U488 ( .A1(n1144), .A2(key_round[42]), .A3(keys1[42]), .A4(n1124), 
        .Y(n548) );
  AO22X1_HVT U489 ( .A1(n983), .A2(key_round[41]), .A3(keys1[41]), .A4(n1125), 
        .Y(n549) );
  AO22X1_HVT U490 ( .A1(n1143), .A2(key_round[40]), .A3(keys1[40]), .A4(n1139), 
        .Y(n550) );
  AO22X1_HVT U491 ( .A1(n799), .A2(key_round[39]), .A3(keys1[39]), .A4(n1140), 
        .Y(n551) );
  AO22X1_HVT U492 ( .A1(n1155), .A2(key_round[38]), .A3(keys1[38]), .A4(n1116), 
        .Y(n552) );
  AO22X1_HVT U493 ( .A1(n1144), .A2(key_round[37]), .A3(keys1[37]), .A4(n1117), 
        .Y(n553) );
  AO22X1_HVT U494 ( .A1(n1147), .A2(key_round[36]), .A3(keys1[36]), .A4(n1116), 
        .Y(n554) );
  AO22X1_HVT U495 ( .A1(n1152), .A2(key_round[35]), .A3(keys1[35]), .A4(n1122), 
        .Y(n555) );
  AO22X1_HVT U496 ( .A1(n792), .A2(key_round[34]), .A3(keys1[34]), .A4(n1133), 
        .Y(n556) );
  AO22X1_HVT U497 ( .A1(n984), .A2(key_round[33]), .A3(keys1[33]), .A4(n1134), 
        .Y(n557) );
  AO22X1_HVT U498 ( .A1(n984), .A2(key_round[32]), .A3(keys1[32]), .A4(n1114), 
        .Y(n558) );
  AO22X1_HVT U499 ( .A1(n1145), .A2(key_round[31]), .A3(keys1[31]), .A4(n1115), 
        .Y(n559) );
  AO22X1_HVT U500 ( .A1(n983), .A2(key_round[30]), .A3(keys1[30]), .A4(n1116), 
        .Y(n560) );
  AO22X1_HVT U501 ( .A1(n1153), .A2(key_round[29]), .A3(keys1[29]), .A4(n1117), 
        .Y(n561) );
  AO22X1_HVT U502 ( .A1(n1152), .A2(key_round[28]), .A3(keys1[28]), .A4(n1124), 
        .Y(n562) );
  AO22X1_HVT U503 ( .A1(n1151), .A2(key_round[27]), .A3(keys1[27]), .A4(n1125), 
        .Y(n563) );
  AO22X1_HVT U504 ( .A1(n793), .A2(key_round[26]), .A3(keys1[26]), .A4(n1136), 
        .Y(n564) );
  AO22X1_HVT U505 ( .A1(n982), .A2(key_round[25]), .A3(keys1[25]), .A4(n1137), 
        .Y(n565) );
  AO22X1_HVT U506 ( .A1(n982), .A2(key_round[24]), .A3(keys1[24]), .A4(n1139), 
        .Y(n566) );
  AO22X1_HVT U507 ( .A1(n985), .A2(key_round[23]), .A3(keys1[23]), .A4(n1137), 
        .Y(n567) );
  AO22X1_HVT U508 ( .A1(n1143), .A2(key_round[22]), .A3(keys1[22]), .A4(n1114), 
        .Y(n568) );
  AO22X1_HVT U509 ( .A1(n1145), .A2(key_round[21]), .A3(keys1[21]), .A4(n1115), 
        .Y(n569) );
  AO22X1_HVT U510 ( .A1(n1145), .A2(key_round[20]), .A3(keys1[20]), .A4(n1114), 
        .Y(n570) );
  AO22X1_HVT U511 ( .A1(n1154), .A2(key_round[19]), .A3(keys1[19]), .A4(n1115), 
        .Y(n571) );
  AO22X1_HVT U512 ( .A1(n799), .A2(key_round[18]), .A3(keys1[18]), .A4(n1125), 
        .Y(n572) );
  AO22X1_HVT U513 ( .A1(n985), .A2(key_round[17]), .A3(keys1[17]), .A4(n1131), 
        .Y(n573) );
  AO22X1_HVT U514 ( .A1(n1146), .A2(key_round[16]), .A3(keys1[16]), .A4(n1136), 
        .Y(n574) );
  AO22X1_HVT U515 ( .A1(n1146), .A2(key_round[15]), .A3(keys1[15]), .A4(n1137), 
        .Y(n575) );
  AO22X1_HVT U516 ( .A1(n1144), .A2(key_round[14]), .A3(keys1[14]), .A4(n1139), 
        .Y(n576) );
  AO22X1_HVT U517 ( .A1(n1143), .A2(key_round[13]), .A3(keys1[13]), .A4(n1140), 
        .Y(n577) );
  AO22X1_HVT U518 ( .A1(n982), .A2(key_round[12]), .A3(keys1[12]), .A4(n1139), 
        .Y(n578) );
  AO22X1_HVT U519 ( .A1(n983), .A2(key_round[11]), .A3(keys1[11]), .A4(n1128), 
        .Y(n579) );
  AO22X1_HVT U520 ( .A1(n1154), .A2(key_round[10]), .A3(keys1[10]), .A4(n1130), 
        .Y(n580) );
  AO22X1_HVT U521 ( .A1(n1155), .A2(key_round[9]), .A3(keys1[9]), .A4(n1131), 
        .Y(n581) );
  AO22X1_HVT U522 ( .A1(n1155), .A2(key_round[8]), .A3(keys1[8]), .A4(n1109), 
        .Y(n582) );
  AO22X1_HVT U523 ( .A1(n792), .A2(key_round[7]), .A3(keys1[7]), .A4(n1109), 
        .Y(n583) );
  AO22X1_HVT U524 ( .A1(n1152), .A2(key_round[6]), .A3(keys1[6]), .A4(n1118), 
        .Y(n584) );
  AO22X1_HVT U525 ( .A1(n1151), .A2(key_round[5]), .A3(keys1[5]), .A4(n1119), 
        .Y(n585) );
  AO22X1_HVT U526 ( .A1(n1151), .A2(key_round[4]), .A3(keys1[4]), .A4(n1121), 
        .Y(n586) );
  AO22X1_HVT U527 ( .A1(n1123), .A2(key_round[3]), .A3(keys1[3]), .A4(n1122), 
        .Y(n587) );
  AO22X1_HVT U528 ( .A1(n1155), .A2(key_round[2]), .A3(keys1[2]), .A4(n1109), 
        .Y(n588) );
  AO22X1_HVT U529 ( .A1(n1155), .A2(key_round[1]), .A3(keys1[1]), .A4(n1164), 
        .Y(n589) );
  AO22X1_HVT U530 ( .A1(n1155), .A2(key_round[0]), .A3(keys1[0]), .A4(n1136), 
        .Y(n590) );
  AO21X1_HVT U532 ( .A1(done), .A2(n158), .A3(n1360), .Y(n591) );
  NAND2X0_HVT U534 ( .A1(n163), .A2(n153), .Y(n160) );
  AO22X1_HVT U535 ( .A1(rount_no[2]), .A2(n161), .A3(n663), .A4(n164), .Y(n593) );
  AND2X1_HVT U539 ( .A1(n156), .A2(n171), .Y(n167) );
  AO22X1_HVT U540 ( .A1(last), .A2(n908), .A3(n663), .A4(n1365), .Y(n595) );
  AO221X1_HVT U541 ( .A1(n1158), .A2(n173), .A3(n1359), .A4(n791), .A5(n1363), 
        .Y(n596) );
  NAND2X0_HVT U542 ( .A1(n174), .A2(n175), .Y(n173) );
  NAND2X0_HVT U545 ( .A1(n1359), .A2(n683), .Y(n176) );
  AO22X1_HVT U546 ( .A1(n1359), .A2(state[0]), .A3(n181), .A4(n182), .Y(n598)
         );
  NAND2X0_HVT U548 ( .A1(n1366), .A2(n159), .Y(n20) );
  NAND2X0_HVT U549 ( .A1(n1158), .A2(n185), .Y(n183) );
  AO221X1_HVT U551 ( .A1(n1158), .A2(n188), .A3(n1359), .A4(state[3]), .A5(
        n1325), .Y(n599) );
  OA21X1_HVT U554 ( .A1(n1364), .A2(n175), .A3(n637), .Y(n191) );
  NAND2X0_HVT U555 ( .A1(n1041), .A2(n153), .Y(n154) );
  AND3X1_HVT U557 ( .A1(n193), .A2(n170), .A3(n166), .Y(n192) );
  AND2X1_HVT U559 ( .A1(n195), .A2(n172), .Y(n194) );
  NAND2X0_HVT U566 ( .A1(n1366), .A2(n200), .Y(n199) );
  OR2X1_HVT U568 ( .A1(n157), .A2(n190), .Y(n159) );
  NAND2X0_HVT U569 ( .A1(n992), .A2(n989), .Y(n190) );
  AO22X1_HVT U571 ( .A1(rount_no[0]), .A2(n161), .A3(n663), .A4(n203), .Y(n601) );
  NAND2X0_HVT U572 ( .A1(n187), .A2(n163), .Y(n203) );
  AND2X1_HVT U576 ( .A1(n193), .A2(n153), .Y(n205) );
  AND3X1_HVT U579 ( .A1(n836), .A2(n166), .A3(n163), .Y(n179) );
  AND2X1_HVT U581 ( .A1(state[3]), .A2(n13), .Y(n197) );
  NAND2X0_HVT U583 ( .A1(n832), .A2(n202), .Y(n169) );
  AND2X1_HVT U584 ( .A1(state[0]), .A2(n12), .Y(n206) );
  AND3X1_HVT U585 ( .A1(n165), .A2(n156), .A3(n180), .Y(n187) );
  AND2X1_HVT U586 ( .A1(n170), .A2(n195), .Y(n180) );
  AND2X1_HVT U589 ( .A1(state[2]), .A2(n14), .Y(n202) );
  NAND3X0_HVT U591 ( .A1(n13), .A2(n12), .A3(n198), .Y(n165) );
  AND2X1_HVT U592 ( .A1(state[1]), .A2(n15), .Y(n198) );
  OR2X1_HVT U594 ( .A1(rest), .A2(n200), .Y(n162) );
  NAND2X0_HVT U595 ( .A1(n184), .A2(n178), .Y(n200) );
  inv_round r1 ( .in({adk_out[127:108], n1184, adk_out[106:76], n1188, 
        adk_out[74:68], n1177, adk_out[66:52], n1173, adk_out[50:44], n1178, 
        adk_out[42:36], n1182, adk_out[34:28], n1093, adk_out[26:15], n1207, 
        adk_out[13:4], n1183, adk_out[2:0]}), .last(last), .keyin(keys1), 
        .out(out1) );
  Get_key as1 ( .clk(clk), .rest(rest), .local_key(local_key), .rount_no(
        rount_no), .key_round(key_round), .done(done_k) );
  DFFSSRX1_HVT flag_reg ( .D(n663), .SETB(n199), .RSTB(1'b1), .CLK(clk), .Q(
        flag), .QN(n606) );
  DFFX1_HVT \adk_out_reg[79]  ( .D(n383), .CLK(clk), .Q(adk_out[79]) );
  DFFX1_HVT \adk_out_reg[119]  ( .D(n343), .CLK(clk), .Q(adk_out[119]), .QN(
        n1034) );
  NAND2X0_HVT U4 ( .A1(n712), .A2(n714), .Y(n673) );
  NAND3X2_HVT U5 ( .A1(n175), .A2(n186), .A3(n187), .Y(n185) );
  NAND3X2_HVT U6 ( .A1(n989), .A2(state[3]), .A3(state[2]), .Y(n175) );
  INVX0_HVT U7 ( .A(n24), .Y(n1318) );
  NAND3X2_HVT U8 ( .A1(state[3]), .A2(n684), .A3(n202), .Y(n153) );
  INVX0_HVT U9 ( .A(n1318), .Y(n1351) );
  NAND2X0_HVT U10 ( .A1(n1219), .A2(n127), .Y(n2) );
  NAND2X0_HVT U11 ( .A1(n1261), .A2(out1[24]), .Y(n3) );
  NAND2X0_HVT U12 ( .A1(n923), .A2(n1347), .Y(n4) );
  NAND3X0_HVT U13 ( .A1(n2), .A2(n3), .A3(n4), .Y(n438) );
  NAND2X0_HVT U14 ( .A1(n1220), .A2(n120), .Y(n5) );
  NAND2X0_HVT U15 ( .A1(n1260), .A2(out1[31]), .Y(n6) );
  NAND2X0_HVT U16 ( .A1(n1040), .A2(n1346), .Y(n7) );
  NAND3X0_HVT U17 ( .A1(n5), .A2(n6), .A3(n7), .Y(n431) );
  DELLN1X2_HVT U18 ( .A(n20), .Y(n8) );
  IBUFFX2_HVT U19 ( .A(n13), .Y(n683) );
  INVX0_HVT U20 ( .A(n24), .Y(n1319) );
  NAND3X0_HVT U21 ( .A1(n836), .A2(n170), .A3(n167), .Y(n168) );
  INVX1_HVT U22 ( .A(n9), .Y(n10) );
  IBUFFX2_HVT U23 ( .A(n987), .Y(n818) );
  IBUFFX2_HVT U24 ( .A(n987), .Y(n819) );
  NAND3X1_HVT U25 ( .A1(n791), .A2(n13), .A3(n206), .Y(n166) );
  INVX1_HVT U26 ( .A(n11), .Y(n18) );
  INVX1_HVT U27 ( .A(n155), .Y(n207) );
  NAND2X0_HVT U28 ( .A1(n815), .A2(n817), .Y(n602) );
  NAND2X0_HVT U29 ( .A1(n603), .A2(n816), .Y(n403) );
  INVX0_HVT U30 ( .A(n602), .Y(n603) );
  IBUFFX2_HVT U31 ( .A(n1318), .Y(n1240) );
  DELLN1X2_HVT U32 ( .A(n24), .Y(n658) );
  NAND2X0_HVT U33 ( .A1(n810), .A2(n812), .Y(n604) );
  NAND2X0_HVT U34 ( .A1(n605), .A2(n811), .Y(n456) );
  INVX0_HVT U35 ( .A(n604), .Y(n605) );
  OR2X1_HVT U36 ( .A1(n162), .A2(n606), .Y(n157) );
  INVX0_HVT U37 ( .A(n162), .Y(n1362) );
  INVX0_HVT U38 ( .A(n1212), .Y(n1217) );
  INVX0_HVT U39 ( .A(n21), .Y(n1212) );
  INVX0_HVT U40 ( .A(n1160), .Y(n1354) );
  NAND3X1_HVT U41 ( .A1(n684), .A2(n14), .A3(n988), .Y(n186) );
  DELLN2X2_HVT U42 ( .A(n178), .Y(n607) );
  IBUFFX2_HVT U43 ( .A(n987), .Y(n1047) );
  IBUFFX2_HVT U44 ( .A(n21), .Y(n1211) );
  AND3X2_HVT U45 ( .A1(n174), .A2(n192), .A3(n186), .Y(n152) );
  NAND2X0_HVT U46 ( .A1(n1217), .A2(n111), .Y(n608) );
  NAND2X0_HVT U47 ( .A1(n1263), .A2(out1[40]), .Y(n609) );
  NAND2X0_HVT U48 ( .A1(adk_out[40]), .A2(n1240), .Y(n610) );
  NAND3X0_HVT U49 ( .A1(n608), .A2(n609), .A3(n610), .Y(n422) );
  NAND2X0_HVT U50 ( .A1(n881), .A2(n879), .Y(n611) );
  NAND2X0_HVT U51 ( .A1(n612), .A2(n880), .Y(n376) );
  INVX0_HVT U52 ( .A(n611), .Y(n612) );
  NAND2X0_HVT U53 ( .A1(n1214), .A2(n65), .Y(n879) );
  IBUFFX2_HVT U54 ( .A(n1361), .Y(n1337) );
  IBUFFX2_HVT U55 ( .A(n1361), .Y(n986) );
  IBUFFX2_HVT U56 ( .A(n1361), .Y(n1338) );
  NAND2X0_HVT U57 ( .A1(n1219), .A2(n121), .Y(n613) );
  NAND2X0_HVT U58 ( .A1(n1259), .A2(out1[30]), .Y(n614) );
  NAND2X0_HVT U59 ( .A1(adk_out[30]), .A2(n1353), .Y(n615) );
  NAND3X0_HVT U60 ( .A1(n613), .A2(n614), .A3(n615), .Y(n432) );
  INVX0_HVT U61 ( .A(n1265), .Y(n1259) );
  AND2X1_HVT U62 ( .A1(n192), .A2(n186), .Y(n616) );
  AND2X1_HVT U63 ( .A1(n616), .A2(n174), .Y(n1041) );
  NAND2X0_HVT U64 ( .A1(n1220), .A2(n38), .Y(n617) );
  NAND2X0_HVT U65 ( .A1(n1276), .A2(out1[113]), .Y(n618) );
  NAND2X0_HVT U66 ( .A1(adk_out[113]), .A2(n677), .Y(n619) );
  NAND3X0_HVT U67 ( .A1(n617), .A2(n618), .A3(n619), .Y(n349) );
  NAND2X0_HVT U68 ( .A1(n1218), .A2(n32), .Y(n620) );
  NAND2X0_HVT U69 ( .A1(out1[119]), .A2(n1270), .Y(n621) );
  NAND2X0_HVT U70 ( .A1(n1035), .A2(n1348), .Y(n622) );
  NAND3X0_HVT U71 ( .A1(n620), .A2(n621), .A3(n622), .Y(n343) );
  INVX0_HVT U72 ( .A(n1355), .Y(n1348) );
  NAND3X4_HVT U73 ( .A1(n183), .A2(n1327), .A3(n184), .Y(n181) );
  AO21X2_HVT U74 ( .A1(n179), .A2(n180), .A3(n157), .Y(n177) );
  AOI21X2_HVT U75 ( .A1(n152), .A2(n156), .A3(n157), .Y(n1208) );
  NAND2X0_HVT U76 ( .A1(n1219), .A2(n39), .Y(n623) );
  NAND2X0_HVT U77 ( .A1(n1276), .A2(out1[112]), .Y(n624) );
  NAND2X0_HVT U78 ( .A1(n894), .A2(n658), .Y(n625) );
  NAND3X0_HVT U79 ( .A1(n623), .A2(n624), .A3(n625), .Y(n350) );
  NAND2X1_HVT U80 ( .A1(n1234), .A2(n88), .Y(n626) );
  NAND2X0_HVT U81 ( .A1(out1[63]), .A2(n1256), .Y(n627) );
  NAND2X1_HVT U82 ( .A1(adk_out[63]), .A2(n1352), .Y(n628) );
  NAND3X0_HVT U83 ( .A1(n626), .A2(n627), .A3(n628), .Y(n399) );
  IBUFFX32_HVT U84 ( .A(n1251), .Y(n1256) );
  NAND2X1_HVT U85 ( .A1(n1230), .A2(n72), .Y(n629) );
  NAND2X0_HVT U86 ( .A1(n1257), .A2(out1[79]), .Y(n630) );
  NAND2X1_HVT U87 ( .A1(adk_out[79]), .A2(n1352), .Y(n631) );
  NAND3X0_HVT U88 ( .A1(n629), .A2(n630), .A3(n631), .Y(n383) );
  INVX0_HVT U89 ( .A(n1319), .Y(n1352) );
  INVX1_HVT U90 ( .A(n632), .Y(n633) );
  NAND2X0_HVT U91 ( .A1(n1220), .A2(n30), .Y(n634) );
  NAND2X0_HVT U92 ( .A1(n1271), .A2(out1[121]), .Y(n635) );
  NAND2X0_HVT U93 ( .A1(adk_out[121]), .A2(n1350), .Y(n636) );
  NAND3X0_HVT U94 ( .A1(n634), .A2(n635), .A3(n636), .Y(n341) );
  AND2X1_HVT U95 ( .A1(n1041), .A2(n153), .Y(n637) );
  NAND2X0_HVT U96 ( .A1(n1222), .A2(n22), .Y(n638) );
  NAND2X0_HVT U97 ( .A1(n1273), .A2(out1[127]), .Y(n639) );
  NAND2X0_HVT U98 ( .A1(n667), .A2(n668), .Y(n640) );
  NAND3X0_HVT U99 ( .A1(n638), .A2(n639), .A3(n640), .Y(n335) );
  NAND2X1_HVT U100 ( .A1(n1224), .A2(n128), .Y(n641) );
  NAND2X0_HVT U101 ( .A1(n1260), .A2(out1[23]), .Y(n642) );
  NAND2X1_HVT U102 ( .A1(adk_out[23]), .A2(n1347), .Y(n643) );
  NAND3X0_HVT U103 ( .A1(n641), .A2(n642), .A3(n643), .Y(n439) );
  NAND2X0_HVT U104 ( .A1(n1218), .A2(n96), .Y(n644) );
  NAND2X0_HVT U105 ( .A1(n1252), .A2(out1[55]), .Y(n645) );
  NAND2X0_HVT U106 ( .A1(adk_out[55]), .A2(n678), .Y(n646) );
  NAND3X0_HVT U107 ( .A1(n644), .A2(n645), .A3(n646), .Y(n407) );
  NAND2X0_HVT U108 ( .A1(n717), .A2(n719), .Y(n647) );
  NAND2X0_HVT U109 ( .A1(n648), .A2(n718), .Y(n336) );
  INVX0_HVT U110 ( .A(n647), .Y(n648) );
  INVX1_HVT U111 ( .A(n649), .Y(n650) );
  NAND2X0_HVT U112 ( .A1(n1078), .A2(n1080), .Y(n651) );
  NAND2X0_HVT U113 ( .A1(n652), .A2(n1079), .Y(n386) );
  INVX0_HVT U114 ( .A(n651), .Y(n652) );
  NAND2X0_HVT U115 ( .A1(n1227), .A2(n75), .Y(n1078) );
  NAND2X0_HVT U116 ( .A1(n1217), .A2(n33), .Y(n653) );
  NAND2X0_HVT U117 ( .A1(n1269), .A2(out1[118]), .Y(n654) );
  NAND2X0_HVT U118 ( .A1(adk_out[118]), .A2(n1350), .Y(n655) );
  NAND3X0_HVT U119 ( .A1(n653), .A2(n654), .A3(n655), .Y(n344) );
  INVX1_HVT U120 ( .A(n656), .Y(n657) );
  NAND2X0_HVT U121 ( .A1(n1219), .A2(n31), .Y(n659) );
  NAND2X0_HVT U122 ( .A1(n1271), .A2(out1[120]), .Y(n660) );
  NAND2X0_HVT U123 ( .A1(n916), .A2(n1351), .Y(n661) );
  NAND3X0_HVT U124 ( .A1(n659), .A2(n660), .A3(n661), .Y(n342) );
  NAND2X0_HVT U125 ( .A1(n154), .A2(n999), .Y(n662) );
  AND2X1_HVT U126 ( .A1(n1362), .A2(flag), .Y(n663) );
  NAND2X0_HVT U127 ( .A1(n1220), .A2(n126), .Y(n946) );
  NAND2X0_HVT U128 ( .A1(n888), .A2(n890), .Y(n664) );
  NAND2X0_HVT U129 ( .A1(n665), .A2(n889), .Y(n395) );
  INVX0_HVT U130 ( .A(n664), .Y(n665) );
  NAND2X0_HVT U131 ( .A1(n1236), .A2(n84), .Y(n888) );
  NAND2X0_HVT U132 ( .A1(n1177), .A2(n1321), .Y(n890) );
  INVX1_HVT U133 ( .A(n666), .Y(n667) );
  NBUFFX2_HVT U134 ( .A(n1238), .Y(n668) );
  IBUFFX2_HVT U135 ( .A(n1355), .Y(n1320) );
  NAND2X0_HVT U136 ( .A1(n694), .A2(n696), .Y(n669) );
  NAND2X0_HVT U137 ( .A1(n670), .A2(n695), .Y(n451) );
  IBUFFX16_HVT U138 ( .A(n669), .Y(n670) );
  NOR2X4_HVT U139 ( .A1(n672), .A2(n1319), .Y(n671) );
  IBUFFX16_HVT U140 ( .A(n671), .Y(n1008) );
  IBUFFX2_HVT U141 ( .A(n1355), .Y(n1237) );
  NAND2X0_HVT U142 ( .A1(n674), .A2(n713), .Y(n441) );
  INVX1_HVT U143 ( .A(n673), .Y(n674) );
  NAND2X0_HVT U193 ( .A1(n1228), .A2(n130), .Y(n712) );
  NAND2X0_HVT U194 ( .A1(adk_out[21]), .A2(n1321), .Y(n714) );
  NAND2X0_HVT U272 ( .A1(n783), .A2(n781), .Y(n675) );
  NAND2X0_HVT U273 ( .A1(n676), .A2(n782), .Y(n435) );
  INVX0_HVT U274 ( .A(n675), .Y(n676) );
  INVX0_HVT U275 ( .A(n1319), .Y(n677) );
  INVX0_HVT U276 ( .A(n1319), .Y(n678) );
  INVX0_HVT U278 ( .A(n1319), .Y(n1322) );
  NAND2X0_HVT U279 ( .A1(n709), .A2(n711), .Y(n679) );
  NAND2X0_HVT U280 ( .A1(n680), .A2(n710), .Y(n405) );
  INVX1_HVT U281 ( .A(n679), .Y(n680) );
  NAND2X0_HVT U282 ( .A1(adk_out[57]), .A2(n1320), .Y(n711) );
  INVX0_HVT U283 ( .A(n722), .Y(n723) );
  DELLN2X2_HVT U284 ( .A(n169), .Y(n836) );
  INVX1_HVT U286 ( .A(n681), .Y(n682) );
  OR3X1_HVT U287 ( .A1(state[1]), .A2(n683), .A3(n831), .Y(n171) );
  INVX0_HVT U288 ( .A(n831), .Y(n832) );
  NAND3X4_HVT U289 ( .A1(n992), .A2(n791), .A3(state[0]), .Y(n163) );
  NBUFFX2_HVT U290 ( .A(n15), .Y(n684) );
  NAND3X2_HVT U291 ( .A1(n165), .A2(n166), .A3(n167), .Y(n164) );
  INVX1_HVT U292 ( .A(n685), .Y(n686) );
  NAND2X0_HVT U293 ( .A1(n1236), .A2(n49), .Y(n687) );
  NAND2X0_HVT U294 ( .A1(n1270), .A2(out1[102]), .Y(n688) );
  NAND2X0_HVT U297 ( .A1(adk_out[102]), .A2(n668), .Y(n689) );
  NAND3X0_HVT U298 ( .A1(n687), .A2(n688), .A3(n689), .Y(n360) );
  INVX1_HVT U299 ( .A(n690), .Y(n691) );
  AO21X2_HVT U300 ( .A1(n999), .A2(n189), .A3(n1325), .Y(n182) );
  DELLN2X2_HVT U301 ( .A(n999), .Y(n1158) );
  IBUFFX2_HVT U302 ( .A(n1318), .Y(n1349) );
  INVX1_HVT U305 ( .A(n1160), .Y(n1355) );
  INVX1_HVT U306 ( .A(n692), .Y(n693) );
  NAND2X0_HVT U307 ( .A1(adk_out[98]), .A2(n1353), .Y(n872) );
  NAND2X0_HVT U308 ( .A1(n1223), .A2(n140), .Y(n694) );
  NAND2X0_HVT U309 ( .A1(out1[11]), .A2(n1278), .Y(n695) );
  NAND2X0_HVT U313 ( .A1(n10), .A2(n1240), .Y(n696) );
  INVX1_HVT U314 ( .A(n697), .Y(n698) );
  INVX1_HVT U315 ( .A(n699), .Y(n700) );
  NAND2X1_HVT U316 ( .A1(n1235), .A2(n77), .Y(n701) );
  NAND2X0_HVT U317 ( .A1(out1[74]), .A2(n1254), .Y(n702) );
  NAND2X1_HVT U318 ( .A1(adk_out[74]), .A2(n1322), .Y(n703) );
  NAND3X0_HVT U320 ( .A1(n701), .A2(n702), .A3(n703), .Y(n388) );
  IBUFFX32_HVT U322 ( .A(n1250), .Y(n1254) );
  NAND2X0_HVT U323 ( .A1(adk_out[111]), .A2(n1351), .Y(n804) );
  INVX0_HVT U324 ( .A(n1338), .Y(n704) );
  INVX0_HVT U325 ( .A(n1338), .Y(n705) );
  INVX0_HVT U329 ( .A(n1338), .Y(n1048) );
  INVX0_HVT U330 ( .A(n1338), .Y(n1329) );
  AND2X1_HVT U331 ( .A1(n827), .A2(n825), .Y(n706) );
  OR2X1_HVT U332 ( .A1(n1038), .A2(n1159), .Y(n1281) );
  INVX0_HVT U334 ( .A(n715), .Y(n716) );
  NAND2X0_HVT U336 ( .A1(n657), .A2(n678), .Y(n812) );
  INVX0_HVT U337 ( .A(n986), .Y(n707) );
  INVX0_HVT U338 ( .A(n986), .Y(n708) );
  NAND2X0_HVT U339 ( .A1(adk_out[86]), .A2(n677), .Y(n881) );
  NAND2X1_HVT U340 ( .A1(n1224), .A2(n94), .Y(n709) );
  NAND2X0_HVT U341 ( .A1(n1253), .A2(out1[57]), .Y(n710) );
  NAND2X0_HVT U342 ( .A1(n706), .A2(n826), .Y(n423) );
  NAND2X0_HVT U343 ( .A1(n1220), .A2(n112), .Y(n825) );
  NAND2X0_HVT U344 ( .A1(adk_out[39]), .A2(n1351), .Y(n827) );
  NAND2X0_HVT U345 ( .A1(out1[21]), .A2(n1259), .Y(n713) );
  NAND2X0_HVT U346 ( .A1(n795), .A2(n797), .Y(n715) );
  NAND2X0_HVT U347 ( .A1(n716), .A2(n796), .Y(n420) );
  NAND2X0_HVT U348 ( .A1(n1219), .A2(n109), .Y(n795) );
  NAND2X0_HVT U349 ( .A1(adk_out[42]), .A2(n1237), .Y(n797) );
  NAND2X0_HVT U350 ( .A1(n1221), .A2(n25), .Y(n717) );
  NAND2X0_HVT U352 ( .A1(n1273), .A2(out1[126]), .Y(n718) );
  NAND2X0_HVT U353 ( .A1(adk_out[126]), .A2(n1350), .Y(n719) );
  NAND2X0_HVT U354 ( .A1(n784), .A2(n786), .Y(n720) );
  NAND2X0_HVT U355 ( .A1(n721), .A2(n785), .Y(n443) );
  IBUFFX16_HVT U356 ( .A(n720), .Y(n721) );
  NAND2X0_HVT U357 ( .A1(n822), .A2(n824), .Y(n722) );
  NAND2X0_HVT U358 ( .A1(n723), .A2(n823), .Y(n339) );
  NAND2X0_HVT U359 ( .A1(n1230), .A2(n28), .Y(n822) );
  NAND2X0_HVT U360 ( .A1(adk_out[123]), .A2(n1348), .Y(n824) );
  INVX0_HVT U361 ( .A(n23), .Y(n1356) );
  INVX1_HVT U362 ( .A(n1024), .Y(n1025) );
  INVX0_HVT U363 ( .A(n662), .Y(n1159) );
  INVX1_HVT U364 ( .A(n920), .Y(n921) );
  INVX0_HVT U365 ( .A(n1344), .Y(n1150) );
  NBUFFX2_HVT U366 ( .A(n198), .Y(n989) );
  NAND2X0_HVT U368 ( .A1(adk_out[34]), .A2(n668), .Y(n1102) );
  NAND2X0_HVT U369 ( .A1(n1221), .A2(n125), .Y(n930) );
  INVX0_HVT U370 ( .A(n986), .Y(n1332) );
  INVX0_HVT U371 ( .A(n199), .Y(n1363) );
  NAND2X0_HVT U372 ( .A1(n1216), .A2(n42), .Y(n917) );
  NAND2X0_HVT U373 ( .A1(n1220), .A2(n45), .Y(n853) );
  NAND2X0_HVT U374 ( .A1(n1215), .A2(n54), .Y(n1003) );
  NAND2X0_HVT U375 ( .A1(n1229), .A2(n57), .Y(n873) );
  NAND2X0_HVT U376 ( .A1(n1216), .A2(n60), .Y(n924) );
  NAND2X0_HVT U377 ( .A1(n1232), .A2(n61), .Y(n862) );
  NAND2X0_HVT U378 ( .A1(adk_out[90]), .A2(n1347), .Y(n864) );
  NAND2X0_HVT U379 ( .A1(n1233), .A2(n69), .Y(n885) );
  NAND2X0_HVT U380 ( .A1(n1228), .A2(n74), .Y(n1097) );
  NAND2X0_HVT U381 ( .A1(n1229), .A2(n81), .Y(n882) );
  NAND2X0_HVT U382 ( .A1(n1234), .A2(n86), .Y(n1066) );
  NAND2X0_HVT U385 ( .A1(n1233), .A2(n89), .Y(n1021) );
  NAND2X0_HVT U386 ( .A1(n1229), .A2(n93), .Y(n949) );
  NAND2X0_HVT U387 ( .A1(n1223), .A2(n95), .Y(n1057) );
  NAND2X0_HVT U388 ( .A1(n1217), .A2(n97), .Y(n837) );
  NAND2X0_HVT U389 ( .A1(n1235), .A2(n102), .Y(n1063) );
  NAND2X0_HVT U390 ( .A1(n1225), .A2(n104), .Y(n840) );
  NAND2X0_HVT U393 ( .A1(n1215), .A2(n105), .Y(n1195) );
  NAND2X0_HVT U394 ( .A1(n1220), .A2(n108), .Y(n1054) );
  NAND2X0_HVT U395 ( .A1(n1218), .A2(n110), .Y(n1060) );
  NAND2X0_HVT U396 ( .A1(n1223), .A2(n134), .Y(n1087) );
  NAND2X0_HVT U397 ( .A1(n1224), .A2(n137), .Y(n955) );
  NAND2X0_HVT U398 ( .A1(n1223), .A2(n138), .Y(n1204) );
  NAND2X0_HVT U399 ( .A1(n1221), .A2(n142), .Y(n1072) );
  NAND2X0_HVT U400 ( .A1(n1235), .A2(n145), .Y(n810) );
  NAND2X0_HVT U401 ( .A1(n1233), .A2(n151), .Y(n859) );
  AND2X1_HVT U404 ( .A1(n955), .A2(n957), .Y(n724) );
  AND2X1_HVT U407 ( .A1(n1163), .A2(n1161), .Y(n725) );
  INVX0_HVT U422 ( .A(n1251), .Y(n1258) );
  INVX0_HVT U423 ( .A(n1277), .Y(n1255) );
  INVX0_HVT U439 ( .A(n1277), .Y(n1257) );
  INVX0_HVT U441 ( .A(n1264), .Y(n1271) );
  INVX0_HVT U531 ( .A(n1265), .Y(n1272) );
  INVX0_HVT U533 ( .A(n1251), .Y(n1262) );
  INVX0_HVT U536 ( .A(n1250), .Y(n1263) );
  AND2X1_HVT U537 ( .A1(n16), .A2(n17), .Y(n726) );
  INVX0_HVT U538 ( .A(n1344), .Y(n1340) );
  INVX0_HVT U543 ( .A(n1135), .Y(n1136) );
  INVX0_HVT U544 ( .A(n1132), .Y(n1137) );
  INVX1_HVT U547 ( .A(n1341), .Y(n1132) );
  INVX0_HVT U550 ( .A(n1344), .Y(n1164) );
  AND2X1_HVT U552 ( .A1(state[2]), .A2(state[1]), .Y(n727) );
  INVX0_HVT U553 ( .A(n1325), .Y(n908) );
  AND2X1_HVT U556 ( .A1(n1192), .A2(n1194), .Y(n728) );
  AND2X1_HVT U558 ( .A1(n856), .A2(n858), .Y(n729) );
  AND2X1_HVT U560 ( .A1(n914), .A2(n912), .Y(n730) );
  AND2X1_HVT U561 ( .A1(n1012), .A2(n1014), .Y(n731) );
  AND2X1_HVT U562 ( .A1(n878), .A2(n876), .Y(n732) );
  AND2X1_HVT U563 ( .A1(n840), .A2(n842), .Y(n733) );
  AND2X1_HVT U564 ( .A1(n1015), .A2(n1017), .Y(n734) );
  AND2X1_HVT U565 ( .A1(n1195), .A2(n1197), .Y(n735) );
  AND2X1_HVT U567 ( .A1(n927), .A2(n929), .Y(n736) );
  AND2X1_HVT U570 ( .A1(n837), .A2(n839), .Y(n737) );
  AND2X1_HVT U573 ( .A1(n1042), .A2(n1044), .Y(n738) );
  AND2X1_HVT U574 ( .A1(n1244), .A2(n1246), .Y(n739) );
  AND2X1_HVT U575 ( .A1(n1021), .A2(n1023), .Y(n740) );
  AND2X1_HVT U577 ( .A1(n949), .A2(n951), .Y(n741) );
  AND2X1_HVT U578 ( .A1(n1198), .A2(n1200), .Y(n742) );
  AND2X1_HVT U580 ( .A1(n1087), .A2(n1089), .Y(n743) );
  AND2X1_HVT U582 ( .A1(n1063), .A2(n1065), .Y(n744) );
  AND2X1_HVT U587 ( .A1(n1029), .A2(n1031), .Y(n745) );
  AND2X1_HVT U588 ( .A1(n1060), .A2(n1062), .Y(n746) );
  AND2X1_HVT U590 ( .A1(n961), .A2(n963), .Y(n747) );
  AND2X1_HVT U593 ( .A1(n917), .A2(n919), .Y(n748) );
  AND2X1_HVT U596 ( .A1(n850), .A2(n852), .Y(n749) );
  AND2X1_HVT U597 ( .A1(n847), .A2(n849), .Y(n750) );
  AND2X1_HVT U598 ( .A1(n869), .A2(n867), .Y(n751) );
  AND2X1_HVT U599 ( .A1(n828), .A2(n830), .Y(n752) );
  AND2X1_HVT U600 ( .A1(n1179), .A2(n1181), .Y(n753) );
  AND2X1_HVT U601 ( .A1(n1072), .A2(n1074), .Y(n754) );
  AND2X1_HVT U602 ( .A1(n1009), .A2(n1011), .Y(n755) );
  AND2X1_HVT U603 ( .A1(n933), .A2(n935), .Y(n756) );
  AND2X1_HVT U604 ( .A1(n1204), .A2(n1206), .Y(n757) );
  AND2X1_HVT U605 ( .A1(n930), .A2(n932), .Y(n758) );
  AND2X1_HVT U606 ( .A1(n1006), .A2(n1008), .Y(n759) );
  AND2X1_HVT U607 ( .A1(n952), .A2(n954), .Y(n760) );
  AND2X1_HVT U608 ( .A1(n1090), .A2(n1092), .Y(n761) );
  AND2X1_HVT U609 ( .A1(n946), .A2(n948), .Y(n762) );
  AND2X1_HVT U610 ( .A1(n909), .A2(n911), .Y(n763) );
  AND2X1_HVT U611 ( .A1(n1003), .A2(n1005), .Y(n764) );
  AND2X1_HVT U612 ( .A1(n1000), .A2(n1002), .Y(n765) );
  AND2X1_HVT U613 ( .A1(n853), .A2(n855), .Y(n766) );
  AND2X1_HVT U614 ( .A1(n941), .A2(n943), .Y(n767) );
  AND2X1_HVT U615 ( .A1(n1102), .A2(n1100), .Y(n768) );
  AND2X1_HVT U616 ( .A1(n899), .A2(n901), .Y(n769) );
  AND2X1_HVT U617 ( .A1(n1054), .A2(n1056), .Y(n770) );
  AND2X1_HVT U618 ( .A1(n958), .A2(n960), .Y(n771) );
  AND2X1_HVT U619 ( .A1(n1097), .A2(n1099), .Y(n772) );
  AND2X1_HVT U620 ( .A1(n924), .A2(n926), .Y(n773) );
  AND2X1_HVT U621 ( .A1(n936), .A2(n938), .Y(n774) );
  AND2X1_HVT U622 ( .A1(n882), .A2(n884), .Y(n775) );
  AND2X1_HVT U623 ( .A1(n873), .A2(n875), .Y(n776) );
  AND2X1_HVT U624 ( .A1(n885), .A2(n887), .Y(n777) );
  AND2X1_HVT U625 ( .A1(n1066), .A2(n1068), .Y(n778) );
  NAND2X0_HVT U626 ( .A1(n763), .A2(n910), .Y(n412) );
  INVX1_HVT U627 ( .A(n779), .Y(n780) );
  NAND2X0_HVT U628 ( .A1(n1222), .A2(n124), .Y(n781) );
  NAND2X0_HVT U629 ( .A1(out1[27]), .A2(n1259), .Y(n782) );
  NAND2X0_HVT U630 ( .A1(n1093), .A2(n1345), .Y(n783) );
  NAND2X0_HVT U631 ( .A1(n1221), .A2(n132), .Y(n784) );
  NAND2X0_HVT U632 ( .A1(out1[19]), .A2(n1276), .Y(n785) );
  NAND2X0_HVT U633 ( .A1(adk_out[19]), .A2(n1238), .Y(n786) );
  NAND2X0_HVT U634 ( .A1(n738), .A2(n1043), .Y(n378) );
  NAND2X0_HVT U635 ( .A1(n743), .A2(n1088), .Y(n445) );
  INVX1_HVT U636 ( .A(n787), .Y(n788) );
  INVX1_HVT U637 ( .A(n789), .Y(n790) );
  NBUFFX2_HVT U638 ( .A(state[1]), .Y(n791) );
  INVX0_HVT U639 ( .A(n1149), .Y(n792) );
  INVX0_HVT U640 ( .A(n1149), .Y(n793) );
  AND3X1_HVT U641 ( .A1(n169), .A2(n165), .A3(n194), .Y(n794) );
  AND2X1_HVT U642 ( .A1(n794), .A2(n171), .Y(n174) );
  NAND2X0_HVT U643 ( .A1(n736), .A2(n928), .Y(n444) );
  NAND2X0_HVT U644 ( .A1(out1[42]), .A2(n1261), .Y(n796) );
  AND3X2_HVT U645 ( .A1(n190), .A2(n186), .A3(n193), .Y(n196) );
  NAND4X1_HVT U646 ( .A1(n190), .A2(n156), .A3(n163), .A4(n191), .Y(n189) );
  NAND2X0_HVT U647 ( .A1(n729), .A2(n857), .Y(n427) );
  NAND2X0_HVT U648 ( .A1(n1216), .A2(n116), .Y(n856) );
  NAND2X0_HVT U649 ( .A1(n18), .A2(n1320), .Y(n858) );
  NAND2X0_HVT U650 ( .A1(n756), .A2(n934), .Y(n440) );
  INVX0_HVT U651 ( .A(n1150), .Y(n798) );
  INVX0_HVT U652 ( .A(n1150), .Y(n799) );
  INVX0_HVT U653 ( .A(n1150), .Y(n1155) );
  NAND2X0_HVT U654 ( .A1(n749), .A2(n851), .Y(n461) );
  INVX0_HVT U655 ( .A(n1149), .Y(n1152) );
  NAND2X0_HVT U656 ( .A1(n770), .A2(n1055), .Y(n419) );
  NAND2X0_HVT U657 ( .A1(n12), .A2(state[2]), .Y(n800) );
  NAND2X0_HVT U658 ( .A1(n198), .A2(n801), .Y(n195) );
  INVX0_HVT U659 ( .A(n800), .Y(n801) );
  NAND2X1_HVT U660 ( .A1(n1218), .A2(n40), .Y(n802) );
  NAND2X0_HVT U661 ( .A1(n1274), .A2(out1[111]), .Y(n803) );
  NAND3X0_HVT U662 ( .A1(n802), .A2(n803), .A3(n804), .Y(n351) );
  NAND2X0_HVT U663 ( .A1(n753), .A2(n1180), .Y(n337) );
  NAND2X0_HVT U664 ( .A1(n1215), .A2(n26), .Y(n1179) );
  NAND2X0_HVT U665 ( .A1(n778), .A2(n1067), .Y(n397) );
  NAND2X0_HVT U666 ( .A1(n750), .A2(n848), .Y(n457) );
  NAND2X0_HVT U667 ( .A1(n1234), .A2(n146), .Y(n847) );
  NAND2X0_HVT U668 ( .A1(adk_out[5]), .A2(n1240), .Y(n849) );
  INVX0_HVT U669 ( .A(n1149), .Y(n1151) );
  INVX0_HVT U670 ( .A(n1343), .Y(n1149) );
  INVX0_HVT U671 ( .A(n1150), .Y(n1153) );
  INVX0_HVT U672 ( .A(n1150), .Y(n1154) );
  NAND2X0_HVT U673 ( .A1(n15), .A2(n12), .Y(n805) );
  NAND2X0_HVT U674 ( .A1(n806), .A2(n202), .Y(n170) );
  INVX0_HVT U675 ( .A(n805), .Y(n806) );
  NAND2X0_HVT U676 ( .A1(n793), .A2(key_round[108]), .Y(n807) );
  NAND2X0_HVT U677 ( .A1(keys1[108]), .A2(n1130), .Y(n808) );
  NAND2X0_HVT U678 ( .A1(n807), .A2(n808), .Y(n482) );
  INVX0_HVT U679 ( .A(n1365), .Y(n809) );
  INVX0_HVT U680 ( .A(n1129), .Y(n1130) );
  NAND2X0_HVT U681 ( .A1(n733), .A2(n841), .Y(n415) );
  NAND2X0_HVT U682 ( .A1(adk_out[47]), .A2(n1347), .Y(n842) );
  NAND2X0_HVT U683 ( .A1(n769), .A2(n900), .Y(n424) );
  NAND2X0_HVT U684 ( .A1(out1[6]), .A2(n1268), .Y(n811) );
  IBUFFX2_HVT U685 ( .A(n172), .Y(n1365) );
  NAND4X1_HVT U686 ( .A1(n163), .A2(n809), .A3(n175), .A4(n196), .Y(n188) );
  NAND2X0_HVT U687 ( .A1(n728), .A2(n1193), .Y(n426) );
  NAND2X0_HVT U688 ( .A1(n942), .A2(n767), .Y(n346) );
  NAND2X0_HVT U689 ( .A1(n1226), .A2(n35), .Y(n941) );
  INVX1_HVT U690 ( .A(n813), .Y(n814) );
  NAND2X0_HVT U691 ( .A1(n1230), .A2(n92), .Y(n815) );
  NAND2X0_HVT U692 ( .A1(out1[59]), .A2(n1254), .Y(n816) );
  NAND2X0_HVT U693 ( .A1(n1157), .A2(n658), .Y(n817) );
  NAND2X0_HVT U694 ( .A1(n959), .A2(n771), .Y(n411) );
  NAND2X0_HVT U695 ( .A1(n744), .A2(n1064), .Y(n413) );
  NAND2X0_HVT U696 ( .A1(n727), .A2(n832), .Y(n193) );
  NAND2X0_HVT U697 ( .A1(n755), .A2(n1010), .Y(n450) );
  NAND2X0_HVT U698 ( .A1(n1222), .A2(n139), .Y(n1009) );
  NAND2X0_HVT U699 ( .A1(n752), .A2(n829), .Y(n338) );
  NAND2X0_HVT U700 ( .A1(n1214), .A2(n27), .Y(n828) );
  NAND2X0_HVT U701 ( .A1(n766), .A2(n854), .Y(n356) );
  NAND2X0_HVT U702 ( .A1(adk_out[106]), .A2(n1348), .Y(n855) );
  NAND2X0_HVT U703 ( .A1(n14), .A2(state[0]), .Y(n820) );
  NAND2X0_HVT U704 ( .A1(n821), .A2(n197), .Y(n172) );
  INVX0_HVT U705 ( .A(n820), .Y(n821) );
  NAND2X0_HVT U706 ( .A1(n737), .A2(n838), .Y(n408) );
  NAND2X0_HVT U707 ( .A1(adk_out[54]), .A2(n1322), .Y(n839) );
  NAND2X0_HVT U708 ( .A1(n746), .A2(n1061), .Y(n421) );
  NAND2X0_HVT U709 ( .A1(n757), .A2(n1205), .Y(n449) );
  NAND2X0_HVT U710 ( .A1(out1[123]), .A2(n1271), .Y(n823) );
  NAND2X0_HVT U711 ( .A1(n730), .A2(n913), .Y(n460) );
  NAND2X0_HVT U712 ( .A1(n1235), .A2(n149), .Y(n912) );
  NAND2X0_HVT U713 ( .A1(adk_out[2]), .A2(n1320), .Y(n914) );
  NAND2X0_HVT U714 ( .A1(n1073), .A2(n754), .Y(n453) );
  NAND2X0_HVT U715 ( .A1(n1260), .A2(out1[39]), .Y(n826) );
  NAND2X0_HVT U716 ( .A1(out1[124]), .A2(n1272), .Y(n829) );
  NAND2X0_HVT U717 ( .A1(n1025), .A2(n1345), .Y(n830) );
  NAND2X0_HVT U718 ( .A1(n762), .A2(n947), .Y(n437) );
  NAND2X0_HVT U719 ( .A1(adk_out[25]), .A2(n1351), .Y(n948) );
  INVX0_HVT U720 ( .A(n206), .Y(n831) );
  NAND2X0_HVT U721 ( .A1(cipher_text[77]), .A2(n1334), .Y(n833) );
  NAND2X0_HVT U722 ( .A1(out1[77]), .A2(n1306), .Y(n834) );
  NAND2X0_HVT U723 ( .A1(n833), .A2(n834), .Y(n257) );
  INVX0_HVT U724 ( .A(n1337), .Y(n835) );
  NAND2X0_HVT U725 ( .A1(out1[54]), .A2(n1269), .Y(n838) );
  NAND2X0_HVT U726 ( .A1(n1273), .A2(out1[47]), .Y(n841) );
  INVX1_HVT U727 ( .A(n843), .Y(n844) );
  NAND2X0_HVT U728 ( .A1(adk_out[125]), .A2(n1323), .Y(n1181) );
  INVX1_HVT U729 ( .A(n845), .Y(n846) );
  NAND2X0_HVT U730 ( .A1(n742), .A2(n1199), .Y(n409) );
  NAND2X0_HVT U731 ( .A1(out1[5]), .A2(n1258), .Y(n848) );
  NAND2X0_HVT U732 ( .A1(n776), .A2(n874), .Y(n368) );
  NAND2X0_HVT U733 ( .A1(adk_out[94]), .A2(n1346), .Y(n875) );
  NAND2X0_HVT U734 ( .A1(n886), .A2(n777), .Y(n380) );
  NAND2X0_HVT U735 ( .A1(adk_out[82]), .A2(n658), .Y(n887) );
  INVX0_HVT U736 ( .A(n20), .Y(n1361) );
  NAND2X0_HVT U737 ( .A1(n1234), .A2(n150), .Y(n850) );
  NAND2X0_HVT U738 ( .A1(out1[1]), .A2(n1267), .Y(n851) );
  NAND2X0_HVT U739 ( .A1(adk_out[1]), .A2(n1352), .Y(n852) );
  NAND2X0_HVT U740 ( .A1(n1272), .A2(out1[106]), .Y(n854) );
  NAND2X0_HVT U741 ( .A1(n918), .A2(n748), .Y(n353) );
  NAND2X0_HVT U742 ( .A1(adk_out[109]), .A2(n1321), .Y(n919) );
  NAND2X0_HVT U743 ( .A1(n1091), .A2(n761), .Y(n370) );
  NAND2X0_HVT U744 ( .A1(n1227), .A2(n59), .Y(n1090) );
  NAND2X0_HVT U745 ( .A1(out1[35]), .A2(n1262), .Y(n857) );
  NAND2X0_HVT U746 ( .A1(n1263), .A2(out1[0]), .Y(n860) );
  NAND2X0_HVT U747 ( .A1(n921), .A2(n1349), .Y(n861) );
  NAND3X0_HVT U748 ( .A1(n859), .A2(n860), .A3(n861), .Y(n462) );
  NAND2X0_HVT U749 ( .A1(n745), .A2(n1030), .Y(n345) );
  NAND2X0_HVT U750 ( .A1(n1245), .A2(n739), .Y(n402) );
  NAND2X0_HVT U751 ( .A1(n868), .A2(n751), .Y(n387) );
  NAND2X0_HVT U752 ( .A1(n1236), .A2(n76), .Y(n867) );
  NAND2X0_HVT U753 ( .A1(n1188), .A2(n1351), .Y(n869) );
  NAND2X0_HVT U754 ( .A1(out1[90]), .A2(n1278), .Y(n863) );
  NAND3X0_HVT U755 ( .A1(n863), .A2(n862), .A3(n864), .Y(n372) );
  INVX1_HVT U756 ( .A(n865), .Y(n866) );
  NAND2X0_HVT U757 ( .A1(out1[75]), .A2(n1255), .Y(n868) );
  NAND2X1_HVT U758 ( .A1(n1231), .A2(n53), .Y(n870) );
  NAND2X0_HVT U759 ( .A1(n1268), .A2(out1[98]), .Y(n871) );
  NAND3X0_HVT U760 ( .A1(n870), .A2(n871), .A3(n872), .Y(n364) );
  NAND2X0_HVT U761 ( .A1(n877), .A2(n732), .Y(n418) );
  NAND2X0_HVT U762 ( .A1(n1214), .A2(n107), .Y(n876) );
  NAND2X0_HVT U763 ( .A1(out1[94]), .A2(n1271), .Y(n874) );
  NAND2X0_HVT U764 ( .A1(out1[44]), .A2(n1269), .Y(n877) );
  NAND2X0_HVT U765 ( .A1(adk_out[44]), .A2(n1350), .Y(n878) );
  NAND2X0_HVT U766 ( .A1(n775), .A2(n883), .Y(n392) );
  NAND2X0_HVT U767 ( .A1(adk_out[70]), .A2(n1350), .Y(n884) );
  NAND2X0_HVT U768 ( .A1(n1259), .A2(out1[86]), .Y(n880) );
  NAND2X0_HVT U769 ( .A1(n962), .A2(n747), .Y(n357) );
  NAND2X0_HVT U770 ( .A1(n1219), .A2(n46), .Y(n961) );
  NAND2X0_HVT U771 ( .A1(adk_out[105]), .A2(n1322), .Y(n963) );
  NAND2X0_HVT U772 ( .A1(n774), .A2(n937), .Y(n352) );
  NAND2X0_HVT U773 ( .A1(n1252), .A2(out1[70]), .Y(n883) );
  INVX0_HVT U774 ( .A(n1277), .Y(n1252) );
  NAND2X0_HVT U775 ( .A1(out1[82]), .A2(n1252), .Y(n886) );
  NAND2X0_HVT U776 ( .A1(out1[67]), .A2(n1261), .Y(n889) );
  NAND2X0_HVT U777 ( .A1(busy), .A2(n158), .Y(n891) );
  INVX0_HVT U778 ( .A(n1363), .Y(n892) );
  NAND2X0_HVT U779 ( .A1(n891), .A2(n892), .Y(n600) );
  NAND2X0_HVT U780 ( .A1(n758), .A2(n931), .Y(n436) );
  NAND2X0_HVT U781 ( .A1(adk_out[26]), .A2(n1351), .Y(n932) );
  INVX1_HVT U782 ( .A(n893), .Y(n894) );
  NAND2X0_HVT U783 ( .A1(n663), .A2(n168), .Y(n895) );
  NAND2X0_HVT U784 ( .A1(rount_no[1]), .A2(n161), .Y(n896) );
  NAND3X0_HVT U785 ( .A1(n895), .A2(n896), .A3(n908), .Y(n594) );
  INVX1_HVT U786 ( .A(n897), .Y(n898) );
  NAND2X0_HVT U787 ( .A1(n735), .A2(n1196), .Y(n416) );
  NAND2X0_HVT U788 ( .A1(adk_out[46]), .A2(n1322), .Y(n1197) );
  NAND2X0_HVT U789 ( .A1(n1219), .A2(n113), .Y(n899) );
  NAND2X0_HVT U790 ( .A1(out1[38]), .A2(n1253), .Y(n900) );
  NAND2X0_HVT U791 ( .A1(adk_out[38]), .A2(n1348), .Y(n901) );
  INVX1_HVT U792 ( .A(n902), .Y(n903) );
  INVX1_HVT U793 ( .A(n904), .Y(n905) );
  NAND2X0_HVT U794 ( .A1(n663), .A2(n160), .Y(n906) );
  NAND2X0_HVT U795 ( .A1(rount_no[3]), .A2(n161), .Y(n907) );
  NAND3X0_HVT U796 ( .A1(n906), .A2(n907), .A3(n908), .Y(n592) );
  AOI21X2_HVT U797 ( .A1(n1158), .A2(n204), .A3(n1325), .Y(n161) );
  NAND3X0_HVT U798 ( .A1(n1364), .A2(n726), .A3(start), .Y(n178) );
  NAND2X0_HVT U799 ( .A1(n1236), .A2(n101), .Y(n909) );
  NAND2X0_HVT U800 ( .A1(n1272), .A2(out1[50]), .Y(n910) );
  NAND2X0_HVT U801 ( .A1(adk_out[50]), .A2(n1240), .Y(n911) );
  NAND2X0_HVT U802 ( .A1(n764), .A2(n1004), .Y(n365) );
  NAND2X0_HVT U803 ( .A1(out1[2]), .A2(n1267), .Y(n913) );
  NAND2X0_HVT U804 ( .A1(n725), .A2(n1162), .Y(n377) );
  NAND2X0_HVT U805 ( .A1(n925), .A2(n773), .Y(n371) );
  NAND2X0_HVT U806 ( .A1(n650), .A2(n1322), .Y(n926) );
  NAND2X0_HVT U807 ( .A1(n765), .A2(n1001), .Y(n362) );
  INVX1_HVT U808 ( .A(n915), .Y(n916) );
  NAND2X0_HVT U809 ( .A1(out1[109]), .A2(n1273), .Y(n918) );
  INVX1_HVT U810 ( .A(n922), .Y(n923) );
  NAND2X0_HVT U811 ( .A1(n956), .A2(n724), .Y(n448) );
  NAND2X0_HVT U812 ( .A1(n1207), .A2(n1238), .Y(n957) );
  NAND2X0_HVT U813 ( .A1(n741), .A2(n950), .Y(n404) );
  NAND2X0_HVT U814 ( .A1(adk_out[58]), .A2(n658), .Y(n951) );
  NAND2X0_HVT U815 ( .A1(out1[91]), .A2(n1278), .Y(n925) );
  NAND2X0_HVT U816 ( .A1(n1224), .A2(n133), .Y(n927) );
  NAND2X0_HVT U817 ( .A1(n1275), .A2(out1[18]), .Y(n928) );
  NAND2X0_HVT U818 ( .A1(adk_out[18]), .A2(n1346), .Y(n929) );
  NAND2X0_HVT U819 ( .A1(n1268), .A2(out1[26]), .Y(n931) );
  NAND2X0_HVT U820 ( .A1(n1223), .A2(n129), .Y(n933) );
  NAND2X0_HVT U821 ( .A1(out1[22]), .A2(n1255), .Y(n934) );
  NAND2X0_HVT U822 ( .A1(n682), .A2(n1323), .Y(n935) );
  NAND2X0_HVT U823 ( .A1(n1217), .A2(n41), .Y(n936) );
  NAND2X0_HVT U824 ( .A1(n1273), .A2(out1[110]), .Y(n937) );
  NAND2X0_HVT U825 ( .A1(n698), .A2(n1353), .Y(n938) );
  NAND2X0_HVT U826 ( .A1(n772), .A2(n1098), .Y(n385) );
  INVX1_HVT U827 ( .A(n939), .Y(n940) );
  NAND2X0_HVT U828 ( .A1(out1[116]), .A2(n1268), .Y(n942) );
  NAND2X0_HVT U829 ( .A1(adk_out[116]), .A2(n678), .Y(n943) );
  INVX1_HVT U830 ( .A(n944), .Y(n945) );
  NAND2X0_HVT U831 ( .A1(n953), .A2(n760), .Y(n433) );
  NAND2X0_HVT U832 ( .A1(n1254), .A2(out1[25]), .Y(n947) );
  NAND2X0_HVT U833 ( .A1(out1[58]), .A2(n1253), .Y(n950) );
  INVX0_HVT U834 ( .A(n1357), .Y(n1253) );
  NAND2X0_HVT U835 ( .A1(n1218), .A2(n122), .Y(n952) );
  NAND2X0_HVT U836 ( .A1(out1[29]), .A2(n1258), .Y(n953) );
  NAND2X0_HVT U837 ( .A1(adk_out[29]), .A2(n1237), .Y(n954) );
  NAND2X0_HVT U838 ( .A1(n740), .A2(n1022), .Y(n400) );
  NAND2X0_HVT U839 ( .A1(out1[14]), .A2(n1267), .Y(n956) );
  NAND2X0_HVT U840 ( .A1(n731), .A2(n1013), .Y(n458) );
  NAND2X0_HVT U841 ( .A1(n1101), .A2(n768), .Y(n428) );
  NAND2X0_HVT U842 ( .A1(n1226), .A2(n117), .Y(n1100) );
  NAND2X0_HVT U843 ( .A1(n759), .A2(n1007), .Y(n434) );
  NAND2X0_HVT U844 ( .A1(n1221), .A2(n100), .Y(n958) );
  NAND2X0_HVT U845 ( .A1(out1[51]), .A2(n1272), .Y(n959) );
  NAND2X0_HVT U846 ( .A1(n1173), .A2(n1240), .Y(n960) );
  NAND2X0_HVT U847 ( .A1(n1016), .A2(n734), .Y(n354) );
  NAND2X0_HVT U848 ( .A1(out1[105]), .A2(n1271), .Y(n962) );
  NAND2X0_HVT U849 ( .A1(adk_out[81]), .A2(n1352), .Y(n1176) );
  INVX0_HVT U850 ( .A(n986), .Y(n1327) );
  INVX0_HVT U851 ( .A(n1338), .Y(n1328) );
  INVX1_HVT U852 ( .A(n1106), .Y(n1107) );
  INVX0_HVT U853 ( .A(n1319), .Y(n1323) );
  NAND2X0_HVT U854 ( .A1(adk_out[37]), .A2(n1348), .Y(n1203) );
  NAND2X0_HVT U855 ( .A1(adk_out[33]), .A2(n1346), .Y(n1071) );
  INVX0_HVT U856 ( .A(n1266), .Y(n1267) );
  INVX0_HVT U857 ( .A(n1319), .Y(n1345) );
  INVX0_HVT U858 ( .A(n1298), .Y(n1052) );
  NAND2X0_HVT U859 ( .A1(n1232), .A2(n43), .Y(n1015) );
  NAND2X0_HVT U860 ( .A1(n1218), .A2(n66), .Y(n1161) );
  NAND2X0_HVT U861 ( .A1(n1217), .A2(n67), .Y(n1042) );
  NAND2X0_HVT U862 ( .A1(n996), .A2(n1321), .Y(n1044) );
  NAND2X0_HVT U863 ( .A1(n1234), .A2(n68), .Y(n1094) );
  NAND2X0_HVT U864 ( .A1(n1224), .A2(n70), .Y(n1174) );
  NAND2X0_HVT U865 ( .A1(n1228), .A2(n82), .Y(n1075) );
  NAND2X0_HVT U866 ( .A1(n1222), .A2(n90), .Y(n1185) );
  NAND2X0_HVT U867 ( .A1(n1222), .A2(n98), .Y(n1198) );
  NAND2X0_HVT U868 ( .A1(adk_out[53]), .A2(n1347), .Y(n1200) );
  NAND2X0_HVT U869 ( .A1(n1217), .A2(n115), .Y(n1192) );
  NAND2X0_HVT U870 ( .A1(n1233), .A2(n147), .Y(n1012) );
  INVX1_HVT U871 ( .A(key_round[126]), .Y(n993) );
  INVX1_HVT U872 ( .A(key_round[123]), .Y(n1171) );
  INVX1_HVT U873 ( .A(key_round[107]), .Y(n1169) );
  INVX1_HVT U874 ( .A(key_round[91]), .Y(n1166) );
  INVX1_HVT U875 ( .A(key_round[89]), .Y(n990) );
  INVX0_HVT U876 ( .A(n1126), .Y(n1110) );
  INVX0_HVT U877 ( .A(n19), .Y(n1358) );
  INVX0_HVT U878 ( .A(n1358), .Y(n1304) );
  INVX0_HVT U879 ( .A(n1358), .Y(n1303) );
  INVX0_HVT U880 ( .A(n1123), .Y(n1111) );
  OAI22X1_HVT U881 ( .A1(n1053), .A2(n986), .A3(n1051), .A4(n1052), .Y(n964)
         );
  AND2X1_HVT U882 ( .A1(n1282), .A2(n1284), .Y(n965) );
  AND2X1_HVT U883 ( .A1(n1247), .A2(n1249), .Y(n966) );
  AND2X1_HVT U884 ( .A1(n1285), .A2(n1287), .Y(n967) );
  AND2X1_HVT U885 ( .A1(n1075), .A2(n1077), .Y(n968) );
  AND2X1_HVT U886 ( .A1(n1018), .A2(n1020), .Y(n969) );
  AND2X1_HVT U887 ( .A1(n1185), .A2(n1187), .Y(n970) );
  AND2X1_HVT U888 ( .A1(n1174), .A2(n1176), .Y(n971) );
  AND2X1_HVT U889 ( .A1(n1094), .A2(n1096), .Y(n972) );
  AND2X1_HVT U890 ( .A1(n1026), .A2(n1028), .Y(n973) );
  AND2X1_HVT U891 ( .A1(n1103), .A2(n1105), .Y(n974) );
  AND2X1_HVT U892 ( .A1(n1203), .A2(n1201), .Y(n975) );
  AND2X1_HVT U893 ( .A1(n1071), .A2(n1069), .Y(n976) );
  AND2X1_HVT U894 ( .A1(n1189), .A2(n1191), .Y(n977) );
  AND2X1_HVT U895 ( .A1(n1084), .A2(n1086), .Y(n978) );
  AND2X1_HVT U896 ( .A1(n1081), .A2(n1083), .Y(n979) );
  AND2X1_HVT U897 ( .A1(n1241), .A2(n1243), .Y(n980) );
  AND2X1_HVT U898 ( .A1(n1279), .A2(n1281), .Y(n981) );
  INVX0_HVT U899 ( .A(n1358), .Y(n1311) );
  INVX0_HVT U900 ( .A(n1135), .Y(n1108) );
  AND3X1_HVT U901 ( .A1(n201), .A2(n159), .A3(n908), .Y(n158) );
  INVX0_HVT U902 ( .A(n1141), .Y(n982) );
  INVX0_HVT U903 ( .A(n1141), .Y(n983) );
  IBUFFX2_HVT U904 ( .A(n1208), .Y(n1141) );
  INVX0_HVT U905 ( .A(n1142), .Y(n984) );
  INVX0_HVT U906 ( .A(n1142), .Y(n985) );
  IBUFFX2_HVT U907 ( .A(n1208), .Y(n1142) );
  INVX0_HVT U908 ( .A(n1141), .Y(n1145) );
  INVX0_HVT U909 ( .A(n1142), .Y(n1146) );
  INVX0_HVT U910 ( .A(n1361), .Y(n987) );
  NBUFFX2_HVT U911 ( .A(n197), .Y(n988) );
  INVX0_HVT U912 ( .A(n1165), .Y(n499) );
  INVX0_HVT U913 ( .A(n1168), .Y(n483) );
  OAI22X1_HVT U914 ( .A1(n1109), .A2(n990), .A3(n991), .A4(n1120), .Y(n501) );
  INVX0_HVT U915 ( .A(n1344), .Y(n1109) );
  INVX0_HVT U916 ( .A(n1120), .Y(n1121) );
  NAND4X1_HVT U917 ( .A1(state[0]), .A2(n202), .A3(n1158), .A4(state[3]), .Y(
        n201) );
  NAND4X1_HVT U918 ( .A1(n684), .A2(n14), .A3(n13), .A4(n12), .Y(n156) );
  NAND2X0_HVT U919 ( .A1(adk_out[65]), .A2(n1353), .Y(n1068) );
  NAND2X0_HVT U920 ( .A1(n903), .A2(n1349), .Y(n1014) );
  NAND4X1_HVT U921 ( .A1(n187), .A2(n179), .A3(n205), .A4(n171), .Y(n204) );
  INVX0_HVT U922 ( .A(out1[127]), .Y(n1051) );
  NBUFFX2_HVT U923 ( .A(n988), .Y(n992) );
  OAI22X1_HVT U924 ( .A1(n1164), .A2(n993), .A3(n994), .A4(n1112), .Y(n464) );
  INVX0_HVT U925 ( .A(n1138), .Y(n1139) );
  INVX1_HVT U926 ( .A(n995), .Y(n996) );
  IBUFFX2_HVT U927 ( .A(n1041), .Y(n1326) );
  IBUFFX2_HVT U928 ( .A(n987), .Y(n1330) );
  IBUFFX2_HVT U929 ( .A(n987), .Y(n1045) );
  IBUFFX2_HVT U930 ( .A(n986), .Y(n1046) );
  INVX1_HVT U931 ( .A(n997), .Y(n998) );
  AND2X1_HVT U932 ( .A1(n1362), .A2(flag), .Y(n999) );
  NAND2X0_HVT U933 ( .A1(adk_out[13]), .A2(n1346), .Y(n1206) );
  NAND2X0_HVT U934 ( .A1(n1216), .A2(n51), .Y(n1000) );
  NAND2X0_HVT U935 ( .A1(out1[100]), .A2(n1269), .Y(n1001) );
  NAND2X0_HVT U936 ( .A1(n898), .A2(n1345), .Y(n1002) );
  NAND2X0_HVT U937 ( .A1(out1[97]), .A2(n1267), .Y(n1004) );
  NAND2X0_HVT U938 ( .A1(adk_out[97]), .A2(n677), .Y(n1005) );
  NAND2X0_HVT U939 ( .A1(n1217), .A2(n123), .Y(n1006) );
  NAND2X0_HVT U940 ( .A1(out1[28]), .A2(n1261), .Y(n1007) );
  NAND2X0_HVT U941 ( .A1(out1[12]), .A2(n1260), .Y(n1010) );
  NAND2X0_HVT U942 ( .A1(adk_out[12]), .A2(n1323), .Y(n1011) );
  NAND2X0_HVT U943 ( .A1(n691), .A2(n1320), .Y(n1080) );
  NAND2X0_HVT U944 ( .A1(out1[4]), .A2(n1263), .Y(n1013) );
  NAND2X0_HVT U945 ( .A1(n1019), .A2(n969), .Y(n442) );
  NAND2X0_HVT U946 ( .A1(n1076), .A2(n968), .Y(n393) );
  NAND2X0_HVT U947 ( .A1(n1027), .A2(n973), .Y(n347) );
  NAND2X0_HVT U948 ( .A1(n1215), .A2(n36), .Y(n1026) );
  NAND2X0_HVT U949 ( .A1(out1[108]), .A2(n1274), .Y(n1016) );
  NAND2X0_HVT U950 ( .A1(n846), .A2(n1345), .Y(n1017) );
  NAND2X0_HVT U951 ( .A1(n1227), .A2(n131), .Y(n1018) );
  NAND2X0_HVT U952 ( .A1(out1[20]), .A2(n1258), .Y(n1019) );
  NAND2X0_HVT U953 ( .A1(n686), .A2(n1321), .Y(n1020) );
  NAND2X0_HVT U954 ( .A1(out1[62]), .A2(n1256), .Y(n1022) );
  NAND2X0_HVT U955 ( .A1(adk_out[62]), .A2(n1322), .Y(n1023) );
  NAND2X0_HVT U956 ( .A1(out1[115]), .A2(n1275), .Y(n1027) );
  NAND2X0_HVT U957 ( .A1(n1107), .A2(n1238), .Y(n1028) );
  NAND2X0_HVT U958 ( .A1(n1216), .A2(n34), .Y(n1029) );
  NAND2X0_HVT U959 ( .A1(out1[117]), .A2(n1268), .Y(n1030) );
  NAND2X0_HVT U960 ( .A1(adk_out[117]), .A2(n1323), .Y(n1031) );
  INVX1_HVT U961 ( .A(n1032), .Y(n1033) );
  INVX1_HVT U962 ( .A(n1034), .Y(n1035) );
  INVX1_HVT U963 ( .A(n1036), .Y(n1037) );
  INVX1_HVT U964 ( .A(n1039), .Y(n1040) );
  NAND2X0_HVT U965 ( .A1(n1085), .A2(n978), .Y(n361) );
  NAND2X0_HVT U966 ( .A1(n1235), .A2(n50), .Y(n1084) );
  NAND2X0_HVT U967 ( .A1(out1[84]), .A2(n1256), .Y(n1043) );
  INVX0_HVT U968 ( .A(n1318), .Y(n1350) );
  DELLN2X2_HVT U969 ( .A(n162), .Y(n1325) );
  IBUFFX2_HVT U970 ( .A(n987), .Y(n1336) );
  NAND2X0_HVT U971 ( .A1(cipher_text[76]), .A2(n819), .Y(n1049) );
  NAND2X0_HVT U972 ( .A1(out1[76]), .A2(n1305), .Y(n1050) );
  NAND2X0_HVT U973 ( .A1(n1049), .A2(n1050), .Y(n258) );
  IBUFFX2_HVT U974 ( .A(n159), .Y(n1360) );
  INVX0_HVT U975 ( .A(n1337), .Y(n1335) );
  INVX0_HVT U976 ( .A(n1337), .Y(n1331) );
  INVX0_HVT U977 ( .A(n1337), .Y(n1333) );
  INVX0_HVT U978 ( .A(n1337), .Y(n1334) );
  NAND2X0_HVT U979 ( .A1(n814), .A2(n1353), .Y(n1194) );
  NAND2X0_HVT U980 ( .A1(n976), .A2(n1070), .Y(n429) );
  NAND2X0_HVT U981 ( .A1(n1215), .A2(n118), .Y(n1069) );
  NAND2X0_HVT U982 ( .A1(n1278), .A2(out1[43]), .Y(n1055) );
  NAND2X0_HVT U983 ( .A1(n1178), .A2(n1237), .Y(n1056) );
  NAND2X0_HVT U984 ( .A1(n1254), .A2(out1[56]), .Y(n1058) );
  NAND2X0_HVT U985 ( .A1(adk_out[56]), .A2(n1351), .Y(n1059) );
  NAND3X0_HVT U986 ( .A1(n1057), .A2(n1058), .A3(n1059), .Y(n406) );
  NAND2X0_HVT U987 ( .A1(n970), .A2(n1186), .Y(n401) );
  NAND2X0_HVT U988 ( .A1(adk_out[61]), .A2(n1237), .Y(n1187) );
  NAND2X0_HVT U989 ( .A1(n1260), .A2(out1[41]), .Y(n1061) );
  NAND2X0_HVT U990 ( .A1(adk_out[41]), .A2(n678), .Y(n1062) );
  NAND2X0_HVT U991 ( .A1(out1[49]), .A2(n1262), .Y(n1064) );
  NAND2X0_HVT U992 ( .A1(adk_out[49]), .A2(n658), .Y(n1065) );
  NAND2X0_HVT U993 ( .A1(n1202), .A2(n975), .Y(n425) );
  NAND2X0_HVT U994 ( .A1(n1218), .A2(n114), .Y(n1201) );
  NAND2X0_HVT U995 ( .A1(out1[65]), .A2(n1269), .Y(n1067) );
  NAND2X0_HVT U996 ( .A1(out1[33]), .A2(n1262), .Y(n1070) );
  NAND2X0_HVT U997 ( .A1(n971), .A2(n1175), .Y(n381) );
  NAND2X0_HVT U998 ( .A1(out1[9]), .A2(n1261), .Y(n1073) );
  NAND2X0_HVT U999 ( .A1(adk_out[9]), .A2(n1321), .Y(n1074) );
  NAND2X0_HVT U1000 ( .A1(out1[69]), .A2(n1272), .Y(n1076) );
  NAND2X0_HVT U1001 ( .A1(adk_out[69]), .A2(n1321), .Y(n1077) );
  NAND2X0_HVT U1002 ( .A1(adk_out[85]), .A2(n658), .Y(n1163) );
  NAND2X0_HVT U1003 ( .A1(n1257), .A2(out1[76]), .Y(n1079) );
  NAND2X0_HVT U1004 ( .A1(n979), .A2(n1082), .Y(n369) );
  NAND2X0_HVT U1005 ( .A1(n1228), .A2(n58), .Y(n1081) );
  NAND2X0_HVT U1006 ( .A1(out1[93]), .A2(n1267), .Y(n1082) );
  NAND2X0_HVT U1007 ( .A1(adk_out[93]), .A2(n1350), .Y(n1083) );
  NAND2X0_HVT U1008 ( .A1(out1[101]), .A2(n1271), .Y(n1085) );
  NAND2X0_HVT U1009 ( .A1(adk_out[101]), .A2(n1349), .Y(n1086) );
  NAND2X0_HVT U1010 ( .A1(n1275), .A2(out1[17]), .Y(n1088) );
  NAND2X0_HVT U1011 ( .A1(adk_out[17]), .A2(n1352), .Y(n1089) );
  NAND2X0_HVT U1012 ( .A1(n974), .A2(n1104), .Y(n459) );
  NAND2X0_HVT U1013 ( .A1(n1236), .A2(n148), .Y(n1103) );
  NAND2X0_HVT U1014 ( .A1(out1[92]), .A2(n1255), .Y(n1091) );
  NAND2X0_HVT U1015 ( .A1(n788), .A2(n677), .Y(n1092) );
  NAND2X0_HVT U1016 ( .A1(n1095), .A2(n972), .Y(n379) );
  NAND2X0_HVT U1017 ( .A1(adk_out[83]), .A2(n1347), .Y(n1096) );
  NAND2X0_HVT U1018 ( .A1(out1[83]), .A2(n1253), .Y(n1095) );
  NAND2X0_HVT U1019 ( .A1(out1[77]), .A2(n1255), .Y(n1098) );
  NAND2X0_HVT U1020 ( .A1(adk_out[77]), .A2(n1350), .Y(n1099) );
  NAND2X0_HVT U1021 ( .A1(out1[34]), .A2(n1263), .Y(n1101) );
  NAND2X0_HVT U1022 ( .A1(n1272), .A2(out1[3]), .Y(n1104) );
  NAND2X0_HVT U1023 ( .A1(n633), .A2(n1320), .Y(n1105) );
  INVX0_HVT U1024 ( .A(n1341), .Y(n1112) );
  INVX0_HVT U1025 ( .A(n1340), .Y(n1113) );
  INVX1_HVT U1026 ( .A(n1112), .Y(n1114) );
  INVX1_HVT U1027 ( .A(n1113), .Y(n1115) );
  INVX1_HVT U1028 ( .A(n1112), .Y(n1116) );
  INVX1_HVT U1029 ( .A(n1113), .Y(n1117) );
  INVX1_HVT U1030 ( .A(n1138), .Y(n1118) );
  INVX1_HVT U1031 ( .A(n1138), .Y(n1119) );
  INVX0_HVT U1032 ( .A(n1340), .Y(n1120) );
  INVX1_HVT U1033 ( .A(n1120), .Y(n1122) );
  INVX0_HVT U1034 ( .A(n1341), .Y(n1123) );
  INVX1_HVT U1035 ( .A(n1132), .Y(n1124) );
  INVX1_HVT U1036 ( .A(n1123), .Y(n1125) );
  INVX0_HVT U1037 ( .A(n1342), .Y(n1126) );
  INVX1_HVT U1038 ( .A(n1126), .Y(n1127) );
  INVX1_HVT U1039 ( .A(n1126), .Y(n1128) );
  INVX0_HVT U1040 ( .A(n1342), .Y(n1129) );
  INVX1_HVT U1041 ( .A(n1129), .Y(n1131) );
  INVX1_HVT U1042 ( .A(n1132), .Y(n1133) );
  INVX1_HVT U1043 ( .A(n1123), .Y(n1134) );
  INVX0_HVT U1044 ( .A(n1342), .Y(n1135) );
  INVX0_HVT U1045 ( .A(n1340), .Y(n1138) );
  INVX1_HVT U1046 ( .A(n1113), .Y(n1140) );
  INVX0_HVT U1047 ( .A(n1141), .Y(n1143) );
  INVX0_HVT U1048 ( .A(n1141), .Y(n1144) );
  INVX0_HVT U1049 ( .A(n1142), .Y(n1147) );
  INVX0_HVT U1050 ( .A(n1142), .Y(n1148) );
  INVX0_HVT U1051 ( .A(n1343), .Y(n1342) );
  INVX0_HVT U1052 ( .A(n1343), .Y(n1341) );
  NAND2X0_HVT U1053 ( .A1(n1242), .A2(n980), .Y(n417) );
  INVX1_HVT U1054 ( .A(n1156), .Y(n1157) );
  INVX0_HVT U1055 ( .A(n1159), .Y(n1160) );
  NAND2X0_HVT U1056 ( .A1(out1[85]), .A2(n1257), .Y(n1162) );
  OA22X1_HVT U1057 ( .A1(n1130), .A2(n1166), .A3(n1167), .A4(n1144), .Y(n1165)
         );
  OA22X1_HVT U1058 ( .A1(n1131), .A2(n1169), .A3(n1170), .A4(n1148), .Y(n1168)
         );
  NAND4X1_HVT U1059 ( .A1(n1328), .A2(n176), .A3(n177), .A4(n607), .Y(n597) );
  OAI22X1_HVT U1060 ( .A1(n1109), .A2(n1171), .A3(n1172), .A4(n798), .Y(n467)
         );
  NAND2X0_HVT U1061 ( .A1(out1[81]), .A2(n1263), .Y(n1175) );
  NAND2X0_HVT U1062 ( .A1(out1[125]), .A2(n1274), .Y(n1180) );
  NAND2X0_HVT U1063 ( .A1(n1257), .A2(out1[61]), .Y(n1186) );
  NAND2X0_HVT U1064 ( .A1(n1280), .A2(n981), .Y(n410) );
  NAND2X0_HVT U1065 ( .A1(n1286), .A2(n967), .Y(n355) );
  NAND2X0_HVT U1066 ( .A1(n1190), .A2(n977), .Y(n394) );
  NAND2X0_HVT U1067 ( .A1(n1227), .A2(n83), .Y(n1189) );
  NAND2X0_HVT U1068 ( .A1(n998), .A2(n1238), .Y(n1191) );
  NAND2X0_HVT U1069 ( .A1(out1[68]), .A2(n1263), .Y(n1190) );
  NAND2X0_HVT U1070 ( .A1(out1[36]), .A2(n1255), .Y(n1193) );
  NAND2X0_HVT U1071 ( .A1(out1[46]), .A2(n1267), .Y(n1196) );
  NAND2X0_HVT U1072 ( .A1(out1[53]), .A2(n1274), .Y(n1199) );
  NAND2X0_HVT U1073 ( .A1(out1[37]), .A2(n1253), .Y(n1202) );
  INVX0_HVT U1074 ( .A(n1355), .Y(n1346) );
  NAND2X0_HVT U1075 ( .A1(out1[13]), .A2(n1278), .Y(n1205) );
  NAND2X0_HVT U1076 ( .A1(n966), .A2(n1248), .Y(n452) );
  NAND2X0_HVT U1077 ( .A1(n965), .A2(n1283), .Y(n363) );
  INVX0_HVT U1078 ( .A(n1318), .Y(n1321) );
  INVX0_HVT U1079 ( .A(n1339), .Y(n1344) );
  INVX0_HVT U1080 ( .A(n1339), .Y(n1343) );
  INVX0_HVT U1081 ( .A(n1208), .Y(n1339) );
  INVX0_HVT U1082 ( .A(n1355), .Y(n1347) );
  INVX0_HVT U1083 ( .A(n1211), .Y(n1215) );
  INVX0_HVT U1084 ( .A(n1211), .Y(n1214) );
  INVX0_HVT U1085 ( .A(n1212), .Y(n1218) );
  INVX0_HVT U1086 ( .A(n1212), .Y(n1220) );
  INVX0_HVT U1087 ( .A(n1212), .Y(n1219) );
  INVX0_HVT U1088 ( .A(n1211), .Y(n1216) );
  IBUFFX2_HVT U1089 ( .A(n21), .Y(n1213) );
  IBUFFX2_HVT U1090 ( .A(n23), .Y(n1277) );
  IBUFFX2_HVT U1091 ( .A(n19), .Y(n1290) );
  INVX0_HVT U1092 ( .A(n1250), .Y(n1261) );
  INVX0_HVT U1093 ( .A(n1251), .Y(n1260) );
  AND3X2_HVT U1094 ( .A1(n17), .A2(n16), .A3(done_k), .Y(n1209) );
  INVX0_HVT U1095 ( .A(n19), .Y(n1289) );
  INVX0_HVT U1096 ( .A(n19), .Y(n1288) );
  NAND2X0_HVT U1097 ( .A1(n1229), .A2(n106), .Y(n1241) );
  NAND2X0_HVT U1098 ( .A1(adk_out[45]), .A2(n1321), .Y(n1243) );
  NAND2X0_HVT U1099 ( .A1(n1227), .A2(n141), .Y(n1247) );
  NAND2X0_HVT U1100 ( .A1(adk_out[10]), .A2(n1349), .Y(n1249) );
  NAND2X0_HVT U1101 ( .A1(n1225), .A2(n52), .Y(n1282) );
  NAND2X0_HVT U1102 ( .A1(adk_out[99]), .A2(n1352), .Y(n1284) );
  NAND2X0_HVT U1103 ( .A1(n1230), .A2(n99), .Y(n1279) );
  NAND2X0_HVT U1104 ( .A1(n1228), .A2(n91), .Y(n1244) );
  NAND2X0_HVT U1105 ( .A1(adk_out[60]), .A2(n677), .Y(n1246) );
  XOR2X1_HVT U1106 ( .A1(plaintext1[68]), .A2(key_round[68]), .Y(n83) );
  XOR2X1_HVT U1107 ( .A1(plaintext1[5]), .A2(key_round[5]), .Y(n146) );
  XOR2X1_HVT U1108 ( .A1(plaintext1[92]), .A2(key_round[92]), .Y(n59) );
  XOR2X1_HVT U1109 ( .A1(plaintext1[123]), .A2(key_round[123]), .Y(n28) );
  XOR2X1_HVT U1110 ( .A1(plaintext1[83]), .A2(key_round[83]), .Y(n68) );
  XOR2X1_HVT U1111 ( .A1(plaintext1[101]), .A2(key_round[101]), .Y(n50) );
  XOR2X1_HVT U1112 ( .A1(plaintext1[93]), .A2(key_round[93]), .Y(n58) );
  XOR2X1_HVT U1113 ( .A1(plaintext1[59]), .A2(key_round[59]), .Y(n92) );
  XOR2X1_HVT U1114 ( .A1(plaintext1[124]), .A2(key_round[124]), .Y(n27) );
  XOR2X1_HVT U1115 ( .A1(plaintext1[98]), .A2(key_round[98]), .Y(n53) );
  XOR2X1_HVT U1116 ( .A1(plaintext1[117]), .A2(key_round[117]), .Y(n34) );
  XOR2X1_HVT U1117 ( .A1(plaintext1[44]), .A2(key_round[44]), .Y(n107) );
  XOR2X1_HVT U1118 ( .A1(plaintext1[36]), .A2(key_round[36]), .Y(n115) );
  XOR2X1_HVT U1119 ( .A1(plaintext1[116]), .A2(key_round[116]), .Y(n35) );
  XOR2X1_HVT U1120 ( .A1(plaintext1[97]), .A2(key_round[97]), .Y(n54) );
  XOR2X1_HVT U1121 ( .A1(plaintext1[25]), .A2(key_round[25]), .Y(n126) );
  XOR2X1_HVT U1122 ( .A1(plaintext1[108]), .A2(key_round[108]), .Y(n43) );
  XOR2X1_HVT U1123 ( .A1(plaintext1[100]), .A2(key_round[100]), .Y(n51) );
  XOR2X1_HVT U1124 ( .A1(plaintext1[85]), .A2(key_round[85]), .Y(n66) );
  XOR2X1_HVT U1125 ( .A1(plaintext1[19]), .A2(key_round[19]), .Y(n132) );
  XOR2X1_HVT U1126 ( .A1(plaintext1[27]), .A2(key_round[27]), .Y(n124) );
  XOR2X1_HVT U1127 ( .A1(plaintext1[57]), .A2(key_round[57]), .Y(n94) );
  XOR2X1_HVT U1128 ( .A1(plaintext1[13]), .A2(key_round[13]), .Y(n138) );
  XOR2X1_HVT U1129 ( .A1(plaintext1[11]), .A2(key_round[11]), .Y(n140) );
  XOR2X1_HVT U1130 ( .A1(plaintext1[20]), .A2(key_round[20]), .Y(n131) );
  XOR2X1_HVT U1131 ( .A1(plaintext1[4]), .A2(key_round[4]), .Y(n147) );
  XOR2X1_HVT U1132 ( .A1(plaintext1[75]), .A2(key_round[75]), .Y(n76) );
  XOR2X1_HVT U1133 ( .A1(plaintext1[76]), .A2(key_round[76]), .Y(n75) );
  XOR2X1_HVT U1134 ( .A1(plaintext1[69]), .A2(key_round[69]), .Y(n82) );
  XOR2X1_HVT U1135 ( .A1(plaintext1[122]), .A2(key_round[122]), .Y(n29) );
  XOR2X1_HVT U1136 ( .A1(plaintext1[82]), .A2(key_round[82]), .Y(n69) );
  XOR2X1_HVT U1137 ( .A1(plaintext1[67]), .A2(key_round[67]), .Y(n84) );
  XOR2X1_HVT U1138 ( .A1(plaintext1[1]), .A2(key_round[1]), .Y(n150) );
  XOR2X1_HVT U1139 ( .A1(plaintext1[73]), .A2(key_round[73]), .Y(n78) );
  XOR2X1_HVT U1140 ( .A1(plaintext1[0]), .A2(key_round[0]), .Y(n151) );
  XOR2X1_HVT U1141 ( .A1(plaintext1[2]), .A2(key_round[2]), .Y(n149) );
  XOR2X1_HVT U1142 ( .A1(plaintext1[74]), .A2(key_round[74]), .Y(n77) );
  XOR2X1_HVT U1143 ( .A1(plaintext1[77]), .A2(key_round[77]), .Y(n74) );
  XOR2X1_HVT U1144 ( .A1(plaintext1[94]), .A2(key_round[94]), .Y(n57) );
  XOR2X1_HVT U1145 ( .A1(plaintext1[70]), .A2(key_round[70]), .Y(n81) );
  XOR2X1_HVT U1146 ( .A1(plaintext1[125]), .A2(key_round[125]), .Y(n26) );
  XOR2X1_HVT U1147 ( .A1(plaintext1[115]), .A2(key_round[115]), .Y(n36) );
  XOR2X1_HVT U1148 ( .A1(plaintext1[84]), .A2(key_round[84]), .Y(n67) );
  XOR2X1_HVT U1149 ( .A1(plaintext1[46]), .A2(key_round[46]), .Y(n105) );
  XOR2X1_HVT U1150 ( .A1(plaintext1[29]), .A2(key_round[29]), .Y(n122) );
  XOR2X1_HVT U1151 ( .A1(plaintext1[28]), .A2(key_round[28]), .Y(n123) );
  XOR2X1_HVT U1152 ( .A1(plaintext1[38]), .A2(key_round[38]), .Y(n113) );
  XOR2X1_HVT U1153 ( .A1(plaintext1[114]), .A2(key_round[114]), .Y(n37) );
  XOR2X1_HVT U1154 ( .A1(plaintext1[41]), .A2(key_round[41]), .Y(n110) );
  XOR2X1_HVT U1155 ( .A1(plaintext1[91]), .A2(key_round[91]), .Y(n60) );
  XOR2X1_HVT U1156 ( .A1(plaintext1[43]), .A2(key_round[43]), .Y(n108) );
  XOR2X1_HVT U1157 ( .A1(plaintext1[113]), .A2(key_round[113]), .Y(n38) );
  XOR2X1_HVT U1158 ( .A1(plaintext1[33]), .A2(key_round[33]), .Y(n118) );
  XOR2X1_HVT U1159 ( .A1(plaintext1[86]), .A2(key_round[86]), .Y(n65) );
  XOR2X1_HVT U1160 ( .A1(plaintext1[121]), .A2(key_round[121]), .Y(n30) );
  XOR2X1_HVT U1161 ( .A1(plaintext1[109]), .A2(key_round[109]), .Y(n42) );
  XOR2X1_HVT U1162 ( .A1(plaintext1[37]), .A2(key_round[37]), .Y(n114) );
  XOR2X1_HVT U1163 ( .A1(plaintext1[42]), .A2(key_round[42]), .Y(n109) );
  XOR2X1_HVT U1164 ( .A1(plaintext1[35]), .A2(key_round[35]), .Y(n116) );
  XOR2X1_HVT U1165 ( .A1(plaintext1[118]), .A2(key_round[118]), .Y(n33) );
  XOR2X1_HVT U1166 ( .A1(plaintext1[61]), .A2(key_round[61]), .Y(n90) );
  XOR2X1_HVT U1167 ( .A1(plaintext1[14]), .A2(key_round[14]), .Y(n137) );
  XOR2X1_HVT U1168 ( .A1(plaintext1[17]), .A2(key_round[17]), .Y(n134) );
  XOR2X1_HVT U1169 ( .A1(plaintext1[12]), .A2(key_round[12]), .Y(n139) );
  XOR2X1_HVT U1170 ( .A1(plaintext1[126]), .A2(key_round[126]), .Y(n25) );
  XOR2X1_HVT U1171 ( .A1(plaintext1[53]), .A2(key_round[53]), .Y(n98) );
  XOR2X1_HVT U1172 ( .A1(plaintext1[81]), .A2(key_round[81]), .Y(n70) );
  XOR2X1_HVT U1173 ( .A1(plaintext1[18]), .A2(key_round[18]), .Y(n133) );
  XOR2X1_HVT U1174 ( .A1(plaintext1[51]), .A2(key_round[51]), .Y(n100) );
  XOR2X1_HVT U1175 ( .A1(plaintext1[26]), .A2(key_round[26]), .Y(n125) );
  NAND2X0_HVT U1176 ( .A1(n1216), .A2(n44), .Y(n1285) );
  NAND2X0_HVT U1177 ( .A1(n693), .A2(n678), .Y(n1287) );
  XOR2X1_HVT U1178 ( .A1(plaintext1[66]), .A2(key_round[66]), .Y(n85) );
  XOR2X1_HVT U1179 ( .A1(plaintext1[3]), .A2(key_round[3]), .Y(n148) );
  XOR2X1_HVT U1180 ( .A1(plaintext1[58]), .A2(key_round[58]), .Y(n93) );
  XOR2X1_HVT U1181 ( .A1(plaintext1[49]), .A2(key_round[49]), .Y(n102) );
  XOR2X1_HVT U1182 ( .A1(plaintext1[65]), .A2(key_round[65]), .Y(n86) );
  XOR2X1_HVT U1183 ( .A1(plaintext1[21]), .A2(key_round[21]), .Y(n130) );
  XOR2X1_HVT U1184 ( .A1(plaintext1[102]), .A2(key_round[102]), .Y(n49) );
  XOR2X1_HVT U1185 ( .A1(plaintext1[62]), .A2(key_round[62]), .Y(n89) );
  XOR2X1_HVT U1186 ( .A1(plaintext1[63]), .A2(key_round[63]), .Y(n88) );
  XOR2X1_HVT U1187 ( .A1(plaintext1[7]), .A2(key_round[7]), .Y(n144) );
  XOR2X1_HVT U1188 ( .A1(plaintext1[89]), .A2(key_round[89]), .Y(n62) );
  XOR2X1_HVT U1189 ( .A1(plaintext1[105]), .A2(key_round[105]), .Y(n46) );
  XOR2X1_HVT U1190 ( .A1(plaintext1[30]), .A2(key_round[30]), .Y(n121) );
  XOR2X1_HVT U1191 ( .A1(plaintext1[106]), .A2(key_round[106]), .Y(n45) );
  XOR2X1_HVT U1192 ( .A1(plaintext1[90]), .A2(key_round[90]), .Y(n61) );
  XOR2X1_HVT U1193 ( .A1(plaintext1[24]), .A2(key_round[24]), .Y(n127) );
  XOR2X1_HVT U1194 ( .A1(plaintext1[120]), .A2(key_round[120]), .Y(n31) );
  XOR2X1_HVT U1195 ( .A1(plaintext1[112]), .A2(key_round[112]), .Y(n39) );
  XOR2X1_HVT U1196 ( .A1(plaintext1[56]), .A2(key_round[56]), .Y(n95) );
  XOR2X1_HVT U1197 ( .A1(plaintext1[9]), .A2(key_round[9]), .Y(n142) );
  XOR2X1_HVT U1198 ( .A1(plaintext1[127]), .A2(key_round[127]), .Y(n22) );
  XOR2X1_HVT U1199 ( .A1(plaintext1[80]), .A2(key_round[80]), .Y(n71) );
  XOR2X1_HVT U1200 ( .A1(plaintext1[50]), .A2(key_round[50]), .Y(n101) );
  XOR2X1_HVT U1201 ( .A1(plaintext1[72]), .A2(key_round[72]), .Y(n79) );
  XOR2X1_HVT U1202 ( .A1(plaintext1[6]), .A2(key_round[6]), .Y(n145) );
  XOR2X1_HVT U1203 ( .A1(plaintext1[95]), .A2(key_round[95]), .Y(n56) );
  XOR2X1_HVT U1204 ( .A1(plaintext1[71]), .A2(key_round[71]), .Y(n80) );
  XOR2X1_HVT U1205 ( .A1(plaintext1[78]), .A2(key_round[78]), .Y(n73) );
  XOR2X1_HVT U1206 ( .A1(plaintext1[104]), .A2(key_round[104]), .Y(n47) );
  XOR2X1_HVT U1207 ( .A1(plaintext1[34]), .A2(key_round[34]), .Y(n117) );
  XOR2X1_HVT U1208 ( .A1(plaintext1[54]), .A2(key_round[54]), .Y(n97) );
  XOR2X1_HVT U1209 ( .A1(plaintext1[87]), .A2(key_round[87]), .Y(n64) );
  XOR2X1_HVT U1210 ( .A1(plaintext1[40]), .A2(key_round[40]), .Y(n111) );
  XOR2X1_HVT U1211 ( .A1(plaintext1[110]), .A2(key_round[110]), .Y(n41) );
  XOR2X1_HVT U1212 ( .A1(plaintext1[47]), .A2(key_round[47]), .Y(n104) );
  XOR2X1_HVT U1213 ( .A1(plaintext1[39]), .A2(key_round[39]), .Y(n112) );
  XOR2X1_HVT U1214 ( .A1(plaintext1[111]), .A2(key_round[111]), .Y(n40) );
  XOR2X1_HVT U1215 ( .A1(plaintext1[8]), .A2(key_round[8]), .Y(n143) );
  XOR2X1_HVT U1216 ( .A1(plaintext1[22]), .A2(key_round[22]), .Y(n129) );
  XOR2X1_HVT U1217 ( .A1(plaintext1[15]), .A2(key_round[15]), .Y(n136) );
  XOR2X1_HVT U1218 ( .A1(plaintext1[64]), .A2(key_round[64]), .Y(n87) );
  XOR2X1_HVT U1219 ( .A1(plaintext1[79]), .A2(key_round[79]), .Y(n72) );
  XOR2X1_HVT U1220 ( .A1(plaintext1[88]), .A2(key_round[88]), .Y(n63) );
  XOR2X1_HVT U1221 ( .A1(plaintext1[32]), .A2(key_round[32]), .Y(n119) );
  XOR2X1_HVT U1222 ( .A1(plaintext1[48]), .A2(key_round[48]), .Y(n103) );
  XOR2X1_HVT U1223 ( .A1(plaintext1[119]), .A2(key_round[119]), .Y(n32) );
  XOR2X1_HVT U1224 ( .A1(plaintext1[96]), .A2(key_round[96]), .Y(n55) );
  XOR2X1_HVT U1225 ( .A1(plaintext1[23]), .A2(key_round[23]), .Y(n128) );
  XOR2X1_HVT U1226 ( .A1(plaintext1[16]), .A2(key_round[16]), .Y(n135) );
  XOR2X1_HVT U1227 ( .A1(plaintext1[103]), .A2(key_round[103]), .Y(n48) );
  XOR2X1_HVT U1228 ( .A1(plaintext1[31]), .A2(key_round[31]), .Y(n120) );
  XOR2X1_HVT U1229 ( .A1(plaintext1[55]), .A2(key_round[55]), .Y(n96) );
  NAND2X0_HVT U1230 ( .A1(n1324), .A2(n1354), .Y(n1210) );
  INVX0_HVT U1231 ( .A(n1213), .Y(n1221) );
  INVX0_HVT U1232 ( .A(n1213), .Y(n1222) );
  INVX0_HVT U1233 ( .A(n1213), .Y(n1223) );
  INVX0_HVT U1234 ( .A(n1213), .Y(n1224) );
  INVX0_HVT U1235 ( .A(n1239), .Y(n1225) );
  INVX0_HVT U1236 ( .A(n1239), .Y(n1226) );
  NBUFFX2_HVT U1237 ( .A(n1225), .Y(n1227) );
  NBUFFX2_HVT U1238 ( .A(n1225), .Y(n1228) );
  NBUFFX2_HVT U1239 ( .A(n1226), .Y(n1229) );
  NBUFFX2_HVT U1240 ( .A(n1226), .Y(n1230) );
  INVX0_HVT U1241 ( .A(n1210), .Y(n1231) );
  INVX0_HVT U1242 ( .A(n1210), .Y(n1232) );
  NBUFFX2_HVT U1243 ( .A(n1231), .Y(n1233) );
  NBUFFX2_HVT U1244 ( .A(n1231), .Y(n1234) );
  NBUFFX2_HVT U1245 ( .A(n1232), .Y(n1235) );
  NBUFFX2_HVT U1246 ( .A(n1232), .Y(n1236) );
  INVX0_HVT U1247 ( .A(n1355), .Y(n1238) );
  NAND2X0_HVT U1248 ( .A1(n1324), .A2(n1354), .Y(n1239) );
  INVX0_HVT U1249 ( .A(n153), .Y(n1324) );
  NAND2X0_HVT U1250 ( .A1(out1[45]), .A2(n1275), .Y(n1242) );
  XOR2X1_HVT U1251 ( .A1(plaintext1[45]), .A2(key_round[45]), .Y(n106) );
  NAND2X0_HVT U1252 ( .A1(out1[60]), .A2(n1255), .Y(n1245) );
  XOR2X1_HVT U1253 ( .A1(plaintext1[60]), .A2(key_round[60]), .Y(n91) );
  NAND2X0_HVT U1254 ( .A1(n1278), .A2(out1[10]), .Y(n1248) );
  XOR2X1_HVT U1255 ( .A1(plaintext1[10]), .A2(key_round[10]), .Y(n141) );
  NBUFFX2_HVT U1256 ( .A(n1357), .Y(n1250) );
  NBUFFX2_HVT U1257 ( .A(n1357), .Y(n1251) );
  NBUFFX2_HVT U1258 ( .A(n1356), .Y(n1264) );
  NBUFFX2_HVT U1259 ( .A(n1356), .Y(n1265) );
  NBUFFX2_HVT U1260 ( .A(n1356), .Y(n1266) );
  INVX0_HVT U1261 ( .A(n1266), .Y(n1268) );
  INVX0_HVT U1262 ( .A(n1264), .Y(n1269) );
  INVX0_HVT U1263 ( .A(n1264), .Y(n1270) );
  INVX0_HVT U1264 ( .A(n1265), .Y(n1273) );
  INVX0_HVT U1265 ( .A(n1265), .Y(n1274) );
  INVX0_HVT U1266 ( .A(n1266), .Y(n1275) );
  INVX0_HVT U1267 ( .A(n1266), .Y(n1276) );
  INVX0_HVT U1268 ( .A(n1277), .Y(n1278) );
  INVX0_HVT U1269 ( .A(n23), .Y(n1357) );
  NAND2X0_HVT U1270 ( .A1(out1[52]), .A2(n1252), .Y(n1280) );
  XOR2X1_HVT U1271 ( .A1(plaintext1[52]), .A2(key_round[52]), .Y(n99) );
  NAND2X0_HVT U1272 ( .A1(n1274), .A2(out1[99]), .Y(n1283) );
  XOR2X1_HVT U1273 ( .A1(plaintext1[99]), .A2(key_round[99]), .Y(n52) );
  NAND2X0_HVT U1274 ( .A1(out1[107]), .A2(n1254), .Y(n1286) );
  XOR2X1_HVT U1275 ( .A1(plaintext1[107]), .A2(key_round[107]), .Y(n44) );
  INVX0_HVT U1276 ( .A(n1288), .Y(n1291) );
  INVX0_HVT U1277 ( .A(n1288), .Y(n1292) );
  INVX0_HVT U1278 ( .A(n1288), .Y(n1293) );
  INVX0_HVT U1279 ( .A(n1288), .Y(n1294) );
  INVX0_HVT U1280 ( .A(n1289), .Y(n1295) );
  INVX0_HVT U1281 ( .A(n1289), .Y(n1296) );
  INVX0_HVT U1282 ( .A(n1289), .Y(n1297) );
  INVX0_HVT U1283 ( .A(n1289), .Y(n1298) );
  INVX0_HVT U1284 ( .A(n1290), .Y(n1299) );
  INVX0_HVT U1285 ( .A(n1290), .Y(n1300) );
  INVX0_HVT U1286 ( .A(n1290), .Y(n1301) );
  INVX0_HVT U1287 ( .A(n1290), .Y(n1302) );
  NBUFFX2_HVT U1288 ( .A(n1303), .Y(n1305) );
  NBUFFX2_HVT U1289 ( .A(n1303), .Y(n1306) );
  NBUFFX2_HVT U1290 ( .A(n1304), .Y(n1307) );
  NBUFFX2_HVT U1291 ( .A(n1304), .Y(n1308) );
  NBUFFX2_HVT U1292 ( .A(n1303), .Y(n1309) );
  NBUFFX2_HVT U1293 ( .A(n1304), .Y(n1310) );
  NBUFFX2_HVT U1294 ( .A(n1311), .Y(n1312) );
  NBUFFX2_HVT U1295 ( .A(n1311), .Y(n1313) );
  NBUFFX2_HVT U1296 ( .A(n1304), .Y(n1314) );
  NBUFFX2_HVT U1297 ( .A(n1303), .Y(n1315) );
  NBUFFX2_HVT U1298 ( .A(n1311), .Y(n1316) );
  NBUFFX2_HVT U1299 ( .A(n1311), .Y(n1317) );
  AND2X1_HVT U1300 ( .A1(n1324), .A2(n1354), .Y(n21) );
  INVX0_HVT U1301 ( .A(n1355), .Y(n1353) );
  AND2X1_HVT U1302 ( .A1(n1354), .A2(n1326), .Y(n23) );
  NAND2X0_HVT U1303 ( .A1(n1209), .A2(start), .Y(n184) );
  INVX0_HVT U1304 ( .A(n182), .Y(n1359) );
  INVX0_HVT U1305 ( .A(done_k), .Y(n1364) );
  INVX0_HVT U1306 ( .A(rest), .Y(n1366) );
endmodule

