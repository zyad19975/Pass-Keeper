
module sbox_7 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n13, n23, n35, n50, n113, n114, n117, n119, n127, n210, n211, n212,
         n213, n216, n217, n218, n219, n222, n224, n225, n227, n229, n231,
         n232, n235, n236, n238, n241, n243, n245, n246, n252, n253, n259,
         n261, n264, n269, n270, n272, n273, n274, n275, n278, n279, n280,
         n282, n283, n284, n285, n291, n293, n297, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748;

  NAND2X0_HVT U4 ( .A1(n483), .A2(n746), .Y(n745) );
  NAND2X0_HVT U5 ( .A1(n393), .A2(n231), .Y(n743) );
  NAND2X0_HVT U15 ( .A1(n746), .A2(n478), .Y(n734) );
  NAND2X0_HVT U21 ( .A1(n229), .A2(n437), .Y(n728) );
  NAND2X0_HVT U24 ( .A1(n477), .A2(n344), .Y(n726) );
  NAND2X0_HVT U33 ( .A1(n519), .A2(n344), .Y(n717) );
  NAND2X0_HVT U35 ( .A1(n446), .A2(n344), .Y(n716) );
  NAND2X0_HVT U42 ( .A1(n409), .A2(n477), .Y(n709) );
  MUX41X1_HVT U51 ( .A1(n506), .A3(n523), .A2(n500), .A4(n348), .S0(n365), 
        .S1(n494), .Y(n701) );
  NAND2X0_HVT U53 ( .A1(n698), .A2(n708), .Y(n699) );
  NAND2X0_HVT U56 ( .A1(n229), .A2(n694), .Y(n695) );
  NAND2X0_HVT U58 ( .A1(n373), .A2(n314), .Y(n692) );
  MUX41X1_HVT U61 ( .A1(n459), .A3(n531), .A2(n238), .A4(n316), .S0(n365), 
        .S1(n493), .Y(n689) );
  NAND2X0_HVT U62 ( .A1(n114), .A2(n484), .Y(n688) );
  MUX41X1_HVT U63 ( .A1(n688), .A3(n510), .A2(n13), .A4(n508), .S0(n365), .S1(
        n493), .Y(n687) );
  AO21X1_HVT U66 ( .A1(n535), .A2(n494), .A3(n537), .Y(n684) );
  MUX41X1_HVT U68 ( .A1(n512), .A3(n684), .A2(n683), .A4(n685), .S0(n468), 
        .S1(n496), .Y(n682) );
  NAND2X0_HVT U73 ( .A1(n396), .A2(n335), .Y(n678) );
  MUX41X1_HVT U74 ( .A1(n679), .A3(n724), .A2(n678), .A4(n726), .S0(n468), 
        .S1(n350), .Y(n676) );
  AND2X1_HVT U83 ( .A1(n409), .A2(n436), .Y(n666) );
  NAND2X0_HVT U85 ( .A1(n437), .A2(n536), .Y(n664) );
  MUX41X1_HVT U90 ( .A1(n705), .A3(n709), .A2(n506), .A4(n661), .S0(n324), 
        .S1(n452), .Y(n660) );
  NAND2X0_HVT U101 ( .A1(n647), .A2(n646), .Y(n648) );
  NAND2X0_HVT U110 ( .A1(n484), .A2(n639), .Y(n640) );
  AND2X1_HVT U115 ( .A1(n409), .A2(n316), .Y(n636) );
  MUX41X1_HVT U116 ( .A1(n241), .A3(n636), .A2(n501), .A4(n719), .S0(n324), 
        .S1(n497), .Y(n635) );
  NAND2X0_HVT U123 ( .A1(n628), .A2(n627), .Y(n629) );
  AND2X1_HVT U140 ( .A1(n396), .A2(n303), .Y(n611) );
  MUX41X1_HVT U142 ( .A1(n351), .A3(n478), .A2(n521), .A4(n397), .S0(n280), 
        .S1(n365), .Y(n609) );
  MUX41X1_HVT U153 ( .A1(n640), .A3(n459), .A2(n264), .A4(n526), .S0(n469), 
        .S1(n451), .Y(n599) );
  AND2X1_HVT U154 ( .A1(n473), .A2(n477), .Y(n598) );
  NAND2X0_HVT U158 ( .A1(n353), .A2(n376), .Y(n594) );
  MUX41X1_HVT U159 ( .A1(n241), .A3(n360), .A2(n594), .A4(n538), .S0(n217), 
        .S1(n451), .Y(n593) );
  AND2X1_HVT U162 ( .A1(n447), .A2(n677), .Y(n590) );
  MUX41X1_HVT U163 ( .A1(n531), .A3(n590), .A2(n456), .A4(n591), .S0(n217), 
        .S1(n451), .Y(n589) );
  NAND2X0_HVT U166 ( .A1(n372), .A2(n694), .Y(n586) );
  NAND2X0_HVT U167 ( .A1(n504), .A2(n445), .Y(n585) );
  MUX41X1_HVT U168 ( .A1(n514), .A3(n480), .A2(n585), .A4(n586), .S0(n324), 
        .S1(n496), .Y(n584) );
  MUX41X1_HVT U176 ( .A1(n446), .A3(n579), .A2(n513), .A4(n736), .S0(n365), 
        .S1(n280), .Y(n578) );
  NAND2X0_HVT U177 ( .A1(n393), .A2(n306), .Y(n577) );
  MUX41X1_HVT U178 ( .A1(n732), .A3(n577), .A2(n414), .A4(n713), .S0(n471), 
        .S1(n452), .Y(n576) );
  MUX41X1_HVT U179 ( .A1(n722), .A3(n528), .A2(n515), .A4(n414), .S0(n469), 
        .S1(n452), .Y(n575) );
  MUX41X1_HVT U182 ( .A1(n517), .A3(n483), .A2(n507), .A4(n525), .S0(n365), 
        .S1(n354), .Y(n572) );
  NAND2X0_HVT U208 ( .A1(n318), .A2(n483), .Y(n639) );
  NAND2X0_HVT U212 ( .A1(n410), .A2(n397), .Y(n694) );
  NAND2X0_HVT U214 ( .A1(n447), .A2(n344), .Y(n548) );
  NAND2X0_HVT U215 ( .A1(n639), .A2(n398), .Y(n547) );
  NAND2X0_HVT U218 ( .A1(n415), .A2(n369), .Y(n601) );
  NAND2X0_HVT U220 ( .A1(n475), .A2(n548), .Y(n669) );
  INVX0_HVT U241 ( .A(n726), .Y(n540) );
  INVX0_HVT U245 ( .A(n743), .Y(n538) );
  INVX0_HVT U256 ( .A(n601), .Y(n532) );
  INVX0_HVT U268 ( .A(n728), .Y(n523) );
  INVX0_HVT U270 ( .A(n547), .Y(n522) );
  INVX0_HVT U271 ( .A(n639), .Y(n521) );
  INVX0_HVT U284 ( .A(n548), .Y(n515) );
  INVX0_HVT U296 ( .A(n734), .Y(n510) );
  INVX0_HVT U297 ( .A(n746), .Y(n509) );
  INVX0_HVT U298 ( .A(n735), .Y(n508) );
  INVX0_HVT U306 ( .A(n585), .Y(n503) );
  INVX0_HVT U307 ( .A(n711), .Y(n502) );
  INVX1_HVT U1 ( .A(n341), .Y(n231) );
  NBUFFX2_HVT U2 ( .A(n343), .Y(n477) );
  XOR2X1_HVT U3 ( .A1(n411), .A2(n396), .Y(n706) );
  AND3X1_HVT U6 ( .A1(n484), .A2(n694), .A3(n669), .Y(n670) );
  MUX21X1_HVT U7 ( .A1(n319), .A2(n735), .S0(n471), .Y(n650) );
  MUX21X1_HVT U8 ( .A1(n487), .A2(n481), .S0(n412), .Y(n210) );
  MUX21X1_HVT U9 ( .A1(n519), .A2(n477), .S0(n344), .Y(n712) );
  INVX1_HVT U10 ( .A(n416), .Y(n496) );
  MUX21X1_HVT U11 ( .A1(n482), .A2(n449), .S0(n488), .Y(n740) );
  MUX21X1_HVT U12 ( .A1(n482), .A2(n359), .S0(n318), .Y(n714) );
  INVX1_HVT U13 ( .A(n730), .Y(n500) );
  AND3X1_HVT U14 ( .A1(n470), .A2(n445), .A3(n436), .Y(n622) );
  MUX21X1_HVT U16 ( .A1(n633), .A2(n634), .S0(n473), .Y(n632) );
  INVX1_HVT U17 ( .A(n489), .Y(n442) );
  INVX1_HVT U18 ( .A(n442), .Y(n437) );
  AND2X1_HVT U19 ( .A1(n736), .A2(n373), .Y(n13) );
  AND2X1_HVT U20 ( .A1(n117), .A2(n119), .Y(n23) );
  INVX0_HVT U22 ( .A(n307), .Y(n306) );
  MUX41X1_HVT U23 ( .A1(n613), .A3(n616), .A2(n615), .A4(n617), .S0(n476), 
        .S1(n472), .Y(n612) );
  INVX1_HVT U25 ( .A(n742), .Y(n270) );
  NAND2X0_HVT U26 ( .A1(n583), .A2(n35), .Y(n50) );
  NAND2X0_HVT U27 ( .A1(n582), .A2(n470), .Y(n113) );
  NAND2X0_HVT U28 ( .A1(n50), .A2(n113), .Y(n581) );
  INVX0_HVT U29 ( .A(n470), .Y(n35) );
  NAND2X0_HVT U30 ( .A1(n397), .A2(n114), .Y(n117) );
  NAND2X0_HVT U31 ( .A1(n231), .A2(n409), .Y(n119) );
  INVX0_HVT U32 ( .A(n409), .Y(n114) );
  MUX21X1_HVT U34 ( .A1(n398), .A2(n23), .S0(n475), .Y(n583) );
  INVX1_HVT U36 ( .A(n489), .Y(n409) );
  MUX21X1_HVT U37 ( .A1(n381), .A2(n319), .S0(n450), .Y(n380) );
  INVX1_HVT U38 ( .A(n499), .Y(n498) );
  INVX1_HVT U39 ( .A(n416), .Y(n350) );
  INVX1_HVT U40 ( .A(n485), .Y(n504) );
  INVX1_HVT U41 ( .A(in[2]), .Y(n492) );
  INVX1_HVT U43 ( .A(n475), .Y(n304) );
  INVX1_HVT U44 ( .A(n488), .Y(n391) );
  INVX1_HVT U45 ( .A(n408), .Y(n217) );
  OA21X1_HVT U46 ( .A1(n503), .A2(n363), .A3(n719), .Y(n607) );
  MUX21X1_HVT U47 ( .A1(n598), .A2(n264), .S0(n461), .Y(n597) );
  OA21X1_HVT U48 ( .A1(n711), .A2(n374), .A3(n601), .Y(n602) );
  INVX1_HVT U49 ( .A(n720), .Y(n529) );
  MUX21X1_HVT U50 ( .A1(n376), .A2(n316), .S0(n392), .Y(n591) );
  INVX1_HVT U52 ( .A(n391), .Y(n392) );
  INVX1_HVT U54 ( .A(n469), .Y(n408) );
  MUX21X1_HVT U55 ( .A1(n436), .A2(n536), .S0(n305), .Y(n715) );
  AO21X1_HVT U57 ( .A1(n457), .A2(n473), .A3(n532), .Y(n558) );
  MUX21X1_HVT U59 ( .A1(n415), .A2(n524), .S0(n495), .Y(n683) );
  MUX21X1_HVT U60 ( .A1(n699), .A2(n700), .S0(n474), .Y(n697) );
  INVX1_HVT U64 ( .A(n461), .Y(n336) );
  MUX21X1_HVT U65 ( .A1(n396), .A2(n270), .S0(n392), .Y(n643) );
  NBUFFX2_HVT U67 ( .A(n491), .Y(n471) );
  MUX21X1_HVT U69 ( .A1(n127), .A2(n618), .S0(n470), .Y(n617) );
  MUX21X1_HVT U70 ( .A1(n360), .A2(n519), .S0(n305), .Y(n654) );
  INVX1_HVT U71 ( .A(in[5]), .Y(n495) );
  INVX1_HVT U72 ( .A(n493), .Y(n434) );
  INVX1_HVT U75 ( .A(n468), .Y(n269) );
  INVX0_HVT U76 ( .A(in[1]), .Y(n489) );
  INVX1_HVT U77 ( .A(n368), .Y(n488) );
  INVX0_HVT U78 ( .A(n391), .Y(n327) );
  INVX0_HVT U79 ( .A(n330), .Y(n318) );
  INVX0_HVT U80 ( .A(n480), .Y(n415) );
  INVX1_HVT U81 ( .A(n490), .Y(n450) );
  INVX1_HVT U82 ( .A(n476), .Y(n253) );
  AND2X1_HVT U84 ( .A1(n246), .A2(n252), .Y(n127) );
  INVX0_HVT U86 ( .A(n445), .Y(n393) );
  INVX1_HVT U87 ( .A(n487), .Y(n376) );
  INVX0_HVT U88 ( .A(n442), .Y(n236) );
  INVX0_HVT U89 ( .A(n442), .Y(n344) );
  INVX1_HVT U91 ( .A(n351), .Y(n727) );
  INVX1_HVT U92 ( .A(n212), .Y(n359) );
  INVX0_HVT U93 ( .A(n319), .Y(n719) );
  INVX0_HVT U94 ( .A(n725), .Y(n501) );
  XOR2X2_HVT U95 ( .A1(n446), .A2(n412), .Y(n724) );
  INVX0_HVT U96 ( .A(n395), .Y(n396) );
  INVX0_HVT U97 ( .A(n395), .Y(n398) );
  MUX21X2_HVT U98 ( .A1(n526), .A2(n379), .S0(n280), .Y(n634) );
  AO21X1_HVT U99 ( .A1(n303), .A2(n415), .A3(n333), .Y(n647) );
  INVX0_HVT U100 ( .A(n474), .Y(n333) );
  MUX41X1_HVT U102 ( .A1(n660), .A3(n653), .A2(n655), .A4(n652), .S0(n253), 
        .S1(n434), .Y(n651) );
  MUX21X1_HVT U103 ( .A1(n465), .A2(n477), .S0(n369), .Y(n730) );
  XOR2X1_HVT U104 ( .A1(n353), .A2(n477), .Y(n703) );
  INVX1_HVT U105 ( .A(n395), .Y(n397) );
  MUX41X1_HVT U106 ( .A1(n589), .A3(n584), .A2(n587), .A4(n581), .S0(n253), 
        .S1(n434), .Y(n580) );
  INVX1_HVT U107 ( .A(n315), .Y(n316) );
  INVX0_HVT U108 ( .A(n732), .Y(n531) );
  INVX0_HVT U109 ( .A(n210), .Y(n713) );
  INVX1_HVT U111 ( .A(n481), .Y(n519) );
  INVX0_HVT U112 ( .A(n741), .Y(n512) );
  INVX1_HVT U113 ( .A(n543), .Y(n518) );
  INVX0_HVT U114 ( .A(n302), .Y(n218) );
  INVX0_HVT U117 ( .A(n318), .Y(n303) );
  INVX0_HVT U118 ( .A(n13), .Y(n211) );
  MUX41X1_HVT U119 ( .A1(n712), .A3(n458), .A2(n705), .A4(n335), .S0(n492), 
        .S1(n496), .Y(n568) );
  INVX1_HVT U120 ( .A(n718), .Y(n516) );
  INVX1_HVT U121 ( .A(n13), .Y(n241) );
  MUX21X1_HVT U122 ( .A1(n444), .A2(n477), .S0(n492), .Y(n638) );
  INVX1_HVT U124 ( .A(n492), .Y(n491) );
  NAND2X0_HVT U125 ( .A1(n309), .A2(n310), .Y(n212) );
  INVX1_HVT U126 ( .A(n453), .Y(n447) );
  INVX0_HVT U127 ( .A(n742), .Y(n360) );
  INVX0_HVT U128 ( .A(n740), .Y(n524) );
  NAND2X0_HVT U129 ( .A1(n456), .A2(n450), .Y(n213) );
  NAND2X0_HVT U130 ( .A1(n238), .A2(n280), .Y(n216) );
  NAND2X0_HVT U131 ( .A1(n213), .A2(n216), .Y(n621) );
  XNOR2X1_HVT U132 ( .A1(n482), .A2(n412), .Y(n456) );
  MUX41X1_HVT U133 ( .A1(n725), .A3(n210), .A2(n611), .A4(n516), .S0(n217), 
        .S1(n365), .Y(n610) );
  MUX41X1_HVT U134 ( .A1(n675), .A3(n680), .A2(n673), .A4(n676), .S0(in[0]), 
        .S1(n434), .Y(n672) );
  NAND2X0_HVT U135 ( .A1(n480), .A2(n218), .Y(n219) );
  NAND2X0_HVT U136 ( .A1(n306), .A2(n302), .Y(n222) );
  NAND2X0_HVT U137 ( .A1(n219), .A2(n222), .Y(n679) );
  INVX0_HVT U138 ( .A(n330), .Y(n302) );
  INVX1_HVT U139 ( .A(n724), .Y(n525) );
  NAND2X0_HVT U141 ( .A1(n602), .A2(n269), .Y(n224) );
  NAND2X0_HVT U143 ( .A1(n603), .A2(n468), .Y(n225) );
  NAND2X0_HVT U144 ( .A1(n224), .A2(n225), .Y(n600) );
  MUX21X1_HVT U145 ( .A1(n448), .A2(n394), .S0(n475), .Y(n603) );
  INVX0_HVT U146 ( .A(n227), .Y(n685) );
  MUX21X1_HVT U147 ( .A1(n393), .A2(n737), .S0(n495), .Y(n227) );
  MUX41X1_HVT U148 ( .A1(n512), .A3(n518), .A2(n728), .A4(n462), .S0(n217), 
        .S1(n304), .Y(n625) );
  MUX21X1_HVT U149 ( .A1(n465), .A2(n359), .S0(n236), .Y(n725) );
  MUX21X1_HVT U150 ( .A1(n436), .A2(n519), .S0(n411), .Y(n718) );
  MUX21X1_HVT U151 ( .A1(n713), .A2(n520), .S0(n474), .Y(n596) );
  MUX21X1_HVT U152 ( .A1(n479), .A2(n465), .S0(n430), .Y(n711) );
  INVX0_HVT U155 ( .A(n284), .Y(n630) );
  MUX21X1_HVT U156 ( .A1(n373), .A2(n229), .S0(n411), .Y(n656) );
  INVX1_HVT U157 ( .A(n236), .Y(n353) );
  NBUFFX2_HVT U160 ( .A(n482), .Y(n229) );
  INVX1_HVT U161 ( .A(n342), .Y(n341) );
  INVX0_HVT U164 ( .A(in[4]), .Y(n527) );
  INVX1_HVT U165 ( .A(n656), .Y(n520) );
  MUX41X1_HVT U169 ( .A1(n514), .A3(n730), .A2(n695), .A4(n738), .S0(n370), 
        .S1(n493), .Y(n693) );
  MUX41X1_HVT U170 ( .A1(n505), .A3(n715), .A2(n455), .A4(n717), .S0(n324), 
        .S1(n374), .Y(n615) );
  MUX41X1_HVT U171 ( .A1(n457), .A3(n455), .A2(n533), .A4(n664), .S0(n468), 
        .S1(n363), .Y(n663) );
  MUX21X1_HVT U172 ( .A1(n436), .A2(n415), .S0(n392), .Y(n732) );
  NAND2X0_HVT U173 ( .A1(n509), .A2(n280), .Y(n232) );
  NAND2X0_HVT U174 ( .A1(n407), .A2(n715), .Y(n235) );
  NAND2X0_HVT U175 ( .A1(n232), .A2(n235), .Y(n334) );
  INVX1_HVT U180 ( .A(n490), .Y(n407) );
  INVX0_HVT U181 ( .A(n640), .Y(n381) );
  INVX0_HVT U183 ( .A(n238), .Y(n733) );
  XOR2X1_HVT U184 ( .A1(n485), .A2(n409), .Y(n702) );
  AND2X1_HVT U185 ( .A1(n328), .A2(n329), .Y(n238) );
  NAND2X0_HVT U186 ( .A1(n530), .A2(n450), .Y(n243) );
  NAND2X0_HVT U187 ( .A1(n720), .A2(n490), .Y(n245) );
  NAND2X0_HVT U188 ( .A1(n243), .A2(n245), .Y(n623) );
  MUX21X1_HVT U189 ( .A1(n231), .A2(n444), .S0(n410), .Y(n720) );
  INVX1_HVT U190 ( .A(n407), .Y(n280) );
  INVX1_HVT U191 ( .A(n236), .Y(n430) );
  NAND2X0_HVT U192 ( .A1(n547), .A2(n272), .Y(n246) );
  NAND2X0_HVT U193 ( .A1(n720), .A2(n304), .Y(n252) );
  MUX41X1_HVT U194 ( .A1(n737), .A3(n718), .A2(n715), .A4(n502), .S0(n470), 
        .S1(n363), .Y(n552) );
  INVX1_HVT U195 ( .A(n363), .Y(n452) );
  INVX0_HVT U196 ( .A(n738), .Y(n535) );
  MUX41X1_HVT U197 ( .A1(n696), .A3(n686), .A2(n690), .A4(n682), .S0(n311), 
        .S1(n253), .Y(out[0]) );
  MUX41X1_HVT U198 ( .A1(n710), .A3(n723), .A2(n317), .A4(n397), .S0(n473), 
        .S1(n468), .Y(n561) );
  NAND2X0_HVT U199 ( .A1(n440), .A2(n304), .Y(n259) );
  NAND2X0_HVT U200 ( .A1(n441), .A2(n382), .Y(n261) );
  NAND2X0_HVT U201 ( .A1(n259), .A2(n261), .Y(n550) );
  MUX21X1_HVT U202 ( .A1(n528), .A2(n319), .S0(n354), .Y(n441) );
  INVX1_HVT U203 ( .A(in[3]), .Y(n342) );
  MUX21X1_HVT U204 ( .A1(n479), .A2(n742), .S0(n430), .Y(n313) );
  NBUFFX2_HVT U205 ( .A(in[7]), .Y(n365) );
  INVX2_HVT U206 ( .A(n498), .Y(n416) );
  MUX41X1_HVT U207 ( .A1(n702), .A3(n563), .A2(n709), .A4(n355), .S0(n471), 
        .S1(n363), .Y(n562) );
  XOR2X2_HVT U209 ( .A1(n353), .A2(n354), .Y(n312) );
  INVX1_HVT U210 ( .A(n442), .Y(n411) );
  INVX0_HVT U211 ( .A(n466), .Y(n637) );
  NBUFFX2_HVT U213 ( .A(n486), .Y(n264) );
  INVX0_HVT U216 ( .A(n709), .Y(n539) );
  MUX41X1_HVT U217 ( .A1(n557), .A3(n561), .A2(n560), .A4(n562), .S0(n476), 
        .S1(n494), .Y(n556) );
  INVX0_HVT U219 ( .A(n712), .Y(n517) );
  MUX41X1_HVT U221 ( .A1(n23), .A3(n447), .A2(n714), .A4(n373), .S0(n269), 
        .S1(n497), .Y(n560) );
  INVX0_HVT U222 ( .A(n453), .Y(n742) );
  MUX41X1_HVT U223 ( .A1(n458), .A3(n540), .A2(n654), .A4(n23), .S0(n269), 
        .S1(n496), .Y(n653) );
  NBUFFX2_HVT U224 ( .A(n360), .Y(n478) );
  INVX1_HVT U225 ( .A(n485), .Y(n465) );
  NAND2X0_HVT U226 ( .A1(n278), .A2(n272), .Y(n273) );
  AND2X1_HVT U227 ( .A1(n273), .A2(n719), .Y(n582) );
  INVX0_HVT U228 ( .A(n304), .Y(n272) );
  INVX1_HVT U229 ( .A(n527), .Y(n436) );
  NAND2X0_HVT U230 ( .A1(n486), .A2(n218), .Y(n274) );
  NAND2X0_HVT U231 ( .A1(n270), .A2(n302), .Y(n275) );
  NAND2X0_HVT U232 ( .A1(n274), .A2(n275), .Y(n710) );
  INVX1_HVT U233 ( .A(n710), .Y(n507) );
  MUX41X1_HVT U234 ( .A1(n642), .A3(n645), .A2(n644), .A4(n649), .S0(n476), 
        .S1(n472), .Y(n641) );
  AO21X1_HVT U235 ( .A1(n473), .A2(n656), .A3(n532), .Y(n657) );
  NAND2X0_HVT U236 ( .A1(n270), .A2(n218), .Y(n278) );
  NAND2X0_HVT U237 ( .A1(n398), .A2(n327), .Y(n279) );
  NAND2X0_HVT U238 ( .A1(n278), .A2(n279), .Y(n317) );
  MUX41X1_HVT U239 ( .A1(n703), .A3(n530), .A2(n522), .A4(n643), .S0(n269), 
        .S1(n496), .Y(n642) );
  NAND2X0_HVT U240 ( .A1(n516), .A2(n280), .Y(n282) );
  NAND2X0_HVT U242 ( .A1(n732), .A2(n407), .Y(n283) );
  NAND2X0_HVT U243 ( .A1(n283), .A2(n282), .Y(n620) );
  MUX21X1_HVT U244 ( .A1(n285), .A2(n717), .S0(n408), .Y(n284) );
  AND2X1_HVT U246 ( .A1(n355), .A2(n356), .Y(n285) );
  NAND2X0_HVT U247 ( .A1(n464), .A2(n291), .Y(n293) );
  NAND2X0_HVT U248 ( .A1(n465), .A2(n312), .Y(n297) );
  NAND2X0_HVT U249 ( .A1(n293), .A2(n297), .Y(n463) );
  INVX0_HVT U250 ( .A(n312), .Y(n291) );
  XNOR2X1_HVT U251 ( .A1(n370), .A2(n347), .Y(n707) );
  MUX41X1_HVT U252 ( .A1(n578), .A3(n575), .A2(n576), .A4(n574), .S0(n253), 
        .S1(n495), .Y(n573) );
  MUX21X2_HVT U253 ( .A1(n394), .A2(n306), .S0(n437), .Y(n414) );
  INVX1_HVT U254 ( .A(n542), .Y(n505) );
  INVX1_HVT U255 ( .A(n437), .Y(n305) );
  INVX1_HVT U257 ( .A(n368), .Y(n410) );
  MUX21X2_HVT U258 ( .A1(n671), .A2(n670), .S0(n471), .Y(n668) );
  MUX41X1_HVT U259 ( .A1(n663), .A3(n665), .A2(n667), .A4(n668), .S0(n472), 
        .S1(n476), .Y(n662) );
  MUX21X1_HVT U260 ( .A1(n415), .A2(n477), .S0(n114), .Y(n544) );
  INVX0_HVT U261 ( .A(n306), .Y(n444) );
  INVX0_HVT U262 ( .A(n722), .Y(n530) );
  NAND2X0_HVT U263 ( .A1(n425), .A2(n424), .Y(out[2]) );
  NAND2X0_HVT U264 ( .A1(n364), .A2(n341), .Y(n309) );
  NAND2X0_HVT U265 ( .A1(n307), .A2(n308), .Y(n310) );
  NAND2X0_HVT U266 ( .A1(n309), .A2(n310), .Y(n453) );
  INVX0_HVT U267 ( .A(n364), .Y(n307) );
  INVX1_HVT U269 ( .A(n341), .Y(n308) );
  INVX0_HVT U272 ( .A(in[4]), .Y(n364) );
  INVX0_HVT U273 ( .A(n646), .Y(n513) );
  INVX1_HVT U274 ( .A(n313), .Y(n448) );
  OA21X1_HVT U275 ( .A1(n375), .A2(n413), .A3(n351), .Y(n570) );
  INVX0_HVT U276 ( .A(in[7]), .Y(n499) );
  INVX1_HVT U277 ( .A(n480), .Y(n394) );
  XOR2X2_HVT U278 ( .A1(n359), .A2(n327), .Y(n705) );
  MUX21X1_HVT U279 ( .A1(n539), .A2(n414), .S0(n474), .Y(n559) );
  INVX0_HVT U280 ( .A(in[6]), .Y(n311) );
  NAND2X0_HVT U281 ( .A1(n322), .A2(n323), .Y(out[1]) );
  MUX41X1_HVT U282 ( .A1(n622), .A3(n623), .A2(n620), .A4(n621), .S0(n382), 
        .S1(n495), .Y(n619) );
  MUX41X1_HVT U283 ( .A1(n533), .A3(n534), .A2(n501), .A4(n504), .S0(n407), 
        .S1(n350), .Y(n675) );
  INVX1_HVT U285 ( .A(n509), .Y(n314) );
  NBUFFX2_HVT U286 ( .A(n498), .Y(n473) );
  INVX1_HVT U287 ( .A(n473), .Y(n374) );
  INVX0_HVT U288 ( .A(n212), .Y(n315) );
  INVX1_HVT U289 ( .A(n541), .Y(n528) );
  INVX1_HVT U290 ( .A(n342), .Y(n343) );
  OA21X1_HVT U291 ( .A1(n304), .A2(n741), .A3(n210), .Y(n554) );
  AND2X1_HVT U292 ( .A1(n345), .A2(n346), .Y(n319) );
  NAND2X0_HVT U293 ( .A1(n454), .A2(n370), .Y(n320) );
  NAND2X0_HVT U294 ( .A1(n733), .A2(n333), .Y(n321) );
  NAND2X0_HVT U295 ( .A1(n320), .A2(n321), .Y(n555) );
  NBUFFX2_HVT U299 ( .A(in[5]), .Y(n494) );
  NAND2X0_HVT U300 ( .A1(n662), .A2(n311), .Y(n322) );
  NAND2X0_HVT U301 ( .A1(n672), .A2(in[6]), .Y(n323) );
  NAND2X0_HVT U302 ( .A1(n607), .A2(n324), .Y(n325) );
  NAND2X0_HVT U303 ( .A1(n608), .A2(n35), .Y(n326) );
  NAND2X0_HVT U304 ( .A1(n325), .A2(n326), .Y(n606) );
  INVX0_HVT U305 ( .A(n450), .Y(n324) );
  MUX41X1_HVT U308 ( .A1(n317), .A3(n394), .A2(n743), .A4(n347), .S0(n490), 
        .S1(n382), .Y(n616) );
  MUX41X1_HVT U309 ( .A1(n568), .A3(n565), .A2(n572), .A4(n569), .S0(n434), 
        .S1(n476), .Y(n564) );
  NAND2X0_HVT U310 ( .A1(n231), .A2(n327), .Y(n328) );
  NAND2X0_HVT U311 ( .A1(n360), .A2(n391), .Y(n329) );
  NBUFFX2_HVT U312 ( .A(n490), .Y(n468) );
  NBUFFX2_HVT U313 ( .A(n368), .Y(n330) );
  NBUFFX2_HVT U314 ( .A(n489), .Y(n368) );
  NAND2X0_HVT U315 ( .A1(n398), .A2(n272), .Y(n331) );
  NAND2X0_HVT U316 ( .A1(n518), .A2(n333), .Y(n332) );
  NAND2X0_HVT U317 ( .A1(n331), .A2(n332), .Y(n618) );
  INVX1_HVT U318 ( .A(n375), .Y(n379) );
  MUX21X1_HVT U319 ( .A1(n479), .A2(n376), .S0(n411), .Y(n375) );
  INVX0_HVT U320 ( .A(n348), .Y(n729) );
  INVX1_HVT U321 ( .A(n537), .Y(n335) );
  INVX1_HVT U322 ( .A(n677), .Y(n537) );
  INVX0_HVT U323 ( .A(n748), .Y(n371) );
  MUX21X1_HVT U324 ( .A1(n486), .A2(n480), .S0(n412), .Y(n735) );
  NAND2X0_HVT U325 ( .A1(n318), .A2(n486), .Y(n746) );
  MUX21X1_HVT U326 ( .A1(n372), .A2(n436), .S0(n411), .Y(n541) );
  MUX21X2_HVT U327 ( .A1(n231), .A2(n359), .S0(n391), .Y(n351) );
  NAND2X0_HVT U328 ( .A1(n486), .A2(n336), .Y(n337) );
  NAND2X0_HVT U329 ( .A1(n659), .A2(n461), .Y(n338) );
  NAND2X0_HVT U330 ( .A1(n337), .A2(n338), .Y(n658) );
  NAND2X0_HVT U331 ( .A1(n658), .A2(n491), .Y(n339) );
  NAND2X0_HVT U332 ( .A1(n657), .A2(n35), .Y(n340) );
  NAND2X0_HVT U333 ( .A1(n339), .A2(n340), .Y(n655) );
  MUX21X1_HVT U334 ( .A1(n477), .A2(n306), .S0(n473), .Y(n659) );
  INVX0_HVT U335 ( .A(n492), .Y(n490) );
  INVX1_HVT U336 ( .A(n745), .Y(n511) );
  INVX0_HVT U337 ( .A(n475), .Y(n413) );
  INVX0_HVT U338 ( .A(n484), .Y(n349) );
  MUX41X1_HVT U339 ( .A1(n740), .A3(n674), .A2(n520), .A4(n448), .S0(n470), 
        .S1(n370), .Y(n673) );
  NAND2X0_HVT U340 ( .A1(n372), .A2(n344), .Y(n345) );
  NAND2X0_HVT U341 ( .A1(n396), .A2(n430), .Y(n346) );
  INVX0_HVT U342 ( .A(n413), .Y(n370) );
  NBUFFX2_HVT U343 ( .A(in[1]), .Y(n412) );
  NAND2X0_HVT U344 ( .A1(n387), .A2(n388), .Y(n347) );
  MUX21X1_HVT U345 ( .A1(n349), .A2(n446), .S0(n236), .Y(n348) );
  INVX1_HVT U346 ( .A(n236), .Y(n369) );
  INVX1_HVT U347 ( .A(n371), .Y(n372) );
  INVX0_HVT U348 ( .A(n333), .Y(n497) );
  INVX0_HVT U349 ( .A(n527), .Y(n352) );
  INVX1_HVT U350 ( .A(n416), .Y(n451) );
  INVX1_HVT U351 ( .A(n739), .Y(n395) );
  NBUFFX2_HVT U352 ( .A(n491), .Y(n354) );
  NAND2X0_HVT U353 ( .A1(n446), .A2(n218), .Y(n355) );
  NAND2X0_HVT U354 ( .A1(n479), .A2(n393), .Y(n356) );
  MUX41X1_HVT U355 ( .A1(n566), .A3(n567), .A2(n736), .A4(n522), .S0(n468), 
        .S1(n474), .Y(n565) );
  OR2X1_HVT U356 ( .A1(n303), .A2(n270), .Y(n736) );
  NAND2X0_HVT U357 ( .A1(n433), .A2(n432), .Y(out[4]) );
  MUX21X1_HVT U358 ( .A1(n745), .A2(n614), .S0(n408), .Y(n613) );
  NAND2X0_HVT U359 ( .A1(n687), .A2(n450), .Y(n357) );
  NAND2X0_HVT U360 ( .A1(n689), .A2(n471), .Y(n358) );
  NAND2X0_HVT U361 ( .A1(n358), .A2(n357), .Y(n686) );
  MUX41X1_HVT U362 ( .A1(n211), .A3(n695), .A2(n727), .A4(n379), .S0(n408), 
        .S1(n350), .Y(n551) );
  MUX41X1_HVT U363 ( .A1(n454), .A3(n740), .A2(n241), .A4(n511), .S0(n35), 
        .S1(n374), .Y(n574) );
  NAND2X0_HVT U364 ( .A1(n691), .A2(n450), .Y(n361) );
  NAND2X0_HVT U365 ( .A1(n693), .A2(n324), .Y(n362) );
  NAND2X0_HVT U366 ( .A1(n361), .A2(n362), .Y(n690) );
  MUX41X1_HVT U367 ( .A1(n705), .A3(n588), .A2(n728), .A4(n529), .S0(n272), 
        .S1(n408), .Y(n587) );
  NBUFFX2_HVT U368 ( .A(n499), .Y(n363) );
  XNOR2X2_HVT U369 ( .A1(n413), .A2(n369), .Y(n461) );
  OR2X1_HVT U370 ( .A1(n330), .A2(n536), .Y(n677) );
  MUX41X1_HVT U371 ( .A1(n348), .A3(n706), .A2(n735), .A4(n540), .S0(n450), 
        .S1(n350), .Y(n667) );
  INVX1_HVT U372 ( .A(n544), .Y(n533) );
  NAND2X0_HVT U373 ( .A1(n517), .A2(n272), .Y(n366) );
  NAND2X0_HVT U374 ( .A1(n727), .A2(n333), .Y(n367) );
  NAND2X0_HVT U375 ( .A1(n366), .A2(n367), .Y(n614) );
  INVX1_HVT U376 ( .A(n716), .Y(n526) );
  INVX0_HVT U377 ( .A(n694), .Y(n534) );
  MUX21X1_HVT U378 ( .A1(n479), .A2(n536), .S0(n302), .Y(n738) );
  MUX41X1_HVT U379 ( .A1(n463), .A3(n334), .A2(n380), .A4(n467), .S0(n494), 
        .S1(n452), .Y(n466) );
  NAND2X0_HVT U380 ( .A1(n630), .A2(n304), .Y(n428) );
  INVX1_HVT U381 ( .A(n371), .Y(n373) );
  MUX41X1_HVT U382 ( .A1(n355), .A3(n443), .A2(n524), .A4(n314), .S0(n269), 
        .S1(n374), .Y(n644) );
  INVX0_HVT U383 ( .A(n435), .Y(n674) );
  INVX1_HVT U384 ( .A(n546), .Y(n506) );
  NBUFFX2_HVT U385 ( .A(n308), .Y(n479) );
  NAND2X0_HVT U386 ( .A1(n571), .A2(n469), .Y(n377) );
  NAND2X0_HVT U387 ( .A1(n570), .A2(n408), .Y(n378) );
  NAND2X0_HVT U388 ( .A1(n377), .A2(n378), .Y(n569) );
  INVX1_HVT U389 ( .A(n487), .Y(n536) );
  MUX41X1_HVT U390 ( .A1(n431), .A3(n460), .A2(n692), .A4(n462), .S0(n363), 
        .S1(n495), .Y(n691) );
  NAND2X0_HVT U391 ( .A1(n417), .A2(n418), .Y(out[5]) );
  NAND2X0_HVT U392 ( .A1(n397), .A2(n382), .Y(n383) );
  NAND2X0_HVT U393 ( .A1(n729), .A2(n413), .Y(n384) );
  NAND2X0_HVT U394 ( .A1(n384), .A2(n383), .Y(n671) );
  INVX0_HVT U395 ( .A(n413), .Y(n382) );
  NAND2X0_HVT U396 ( .A1(n556), .A2(in[6]), .Y(n385) );
  NAND2X0_HVT U397 ( .A1(n549), .A2(n311), .Y(n386) );
  NAND2X0_HVT U398 ( .A1(n385), .A2(n386), .Y(out[7]) );
  NAND2X0_HVT U399 ( .A1(n465), .A2(n344), .Y(n387) );
  NAND2X0_HVT U400 ( .A1(n376), .A2(n430), .Y(n388) );
  NAND2X0_HVT U401 ( .A1(n387), .A2(n388), .Y(n723) );
  NAND2X0_HVT U402 ( .A1(n422), .A2(n423), .Y(n624) );
  NAND2X0_HVT U403 ( .A1(n635), .A2(n472), .Y(n389) );
  NAND2X0_HVT U404 ( .A1(n632), .A2(n434), .Y(n390) );
  NAND2X0_HVT U405 ( .A1(n390), .A2(n389), .Y(n631) );
  MUX41X1_HVT U406 ( .A1(n631), .A3(n637), .A2(n619), .A4(n624), .S0(n476), 
        .S1(n311), .Y(out[3]) );
  INVX1_HVT U407 ( .A(n410), .Y(n445) );
  NBUFFX2_HVT U408 ( .A(n739), .Y(n480) );
  NAND2X0_HVT U409 ( .A1(n597), .A2(n324), .Y(n399) );
  NAND2X0_HVT U410 ( .A1(n596), .A2(n35), .Y(n400) );
  NAND2X0_HVT U411 ( .A1(n399), .A2(n400), .Y(n595) );
  INVX0_HVT U412 ( .A(n431), .Y(n731) );
  NAND2X0_HVT U413 ( .A1(n558), .A2(n471), .Y(n401) );
  NAND2X0_HVT U414 ( .A1(n559), .A2(n35), .Y(n402) );
  NAND2X0_HVT U415 ( .A1(n401), .A2(n402), .Y(n557) );
  NAND2X0_HVT U416 ( .A1(n564), .A2(n311), .Y(n403) );
  NAND2X0_HVT U417 ( .A1(n573), .A2(in[6]), .Y(n404) );
  NAND2X0_HVT U418 ( .A1(n404), .A2(n403), .Y(out[6]) );
  NAND2X0_HVT U419 ( .A1(n701), .A2(n490), .Y(n405) );
  NAND2X0_HVT U420 ( .A1(n697), .A2(n35), .Y(n406) );
  NAND2X0_HVT U421 ( .A1(n406), .A2(n405), .Y(n696) );
  INVX1_HVT U422 ( .A(n231), .Y(n449) );
  MUX41X1_HVT U423 ( .A1(n550), .A3(n551), .A2(n552), .A4(n553), .S0(n472), 
        .S1(n476), .Y(n549) );
  MUX41X1_HVT U424 ( .A1(n733), .A3(n666), .A2(n351), .A4(n447), .S0(n491), 
        .S1(n416), .Y(n665) );
  AO21X1_HVT U425 ( .A1(n714), .A2(n471), .A3(n731), .Y(n467) );
  NAND2X0_HVT U426 ( .A1(n580), .A2(n311), .Y(n417) );
  NAND2X0_HVT U427 ( .A1(n592), .A2(in[6]), .Y(n418) );
  MUX21X1_HVT U428 ( .A1(n482), .A2(n444), .S0(n437), .Y(n443) );
  NAND2X0_HVT U429 ( .A1(n459), .A2(n419), .Y(n420) );
  NAND2X0_HVT U430 ( .A1(n650), .A2(n704), .Y(n421) );
  NAND2X0_HVT U431 ( .A1(n420), .A2(n421), .Y(n649) );
  INVX0_HVT U432 ( .A(n704), .Y(n419) );
  NAND2X0_HVT U433 ( .A1(n625), .A2(n434), .Y(n422) );
  NAND2X0_HVT U434 ( .A1(n626), .A2(n472), .Y(n423) );
  MUX21X1_HVT U435 ( .A1(n444), .A2(n746), .S0(n354), .Y(n440) );
  AO21X1_HVT U436 ( .A1(n471), .A2(n398), .A3(n447), .Y(n633) );
  NAND2X0_HVT U437 ( .A1(n641), .A2(n311), .Y(n424) );
  NAND2X0_HVT U438 ( .A1(n651), .A2(in[6]), .Y(n425) );
  NAND2X0_HVT U439 ( .A1(n554), .A2(n450), .Y(n426) );
  NAND2X0_HVT U440 ( .A1(n555), .A2(n469), .Y(n427) );
  NAND2X0_HVT U441 ( .A1(n426), .A2(n427), .Y(n553) );
  MUX41X1_HVT U442 ( .A1(n458), .A3(n534), .A2(n734), .A4(n327), .S0(n269), 
        .S1(n451), .Y(n652) );
  NAND2X0_HVT U443 ( .A1(n604), .A2(n311), .Y(n432) );
  MUX41X1_HVT U444 ( .A1(n600), .A3(n595), .A2(n599), .A4(n593), .S0(n253), 
        .S1(n495), .Y(n592) );
  NAND2X0_HVT U445 ( .A1(n629), .A2(n370), .Y(n429) );
  NAND2X0_HVT U446 ( .A1(n428), .A2(n429), .Y(n626) );
  MUX21X1_HVT U447 ( .A1(n398), .A2(n229), .S0(n369), .Y(n431) );
  NAND2X0_HVT U448 ( .A1(n612), .A2(in[6]), .Y(n433) );
  MUX21X1_HVT U449 ( .A1(n436), .A2(n270), .S0(n344), .Y(n435) );
  NAND2X0_HVT U450 ( .A1(n681), .A2(n217), .Y(n438) );
  NAND2X0_HVT U451 ( .A1(n707), .A2(n35), .Y(n439) );
  NAND2X0_HVT U452 ( .A1(n439), .A2(n438), .Y(n680) );
  MUX21X1_HVT U453 ( .A1(n316), .A2(n536), .S0(n305), .Y(n741) );
  MUX21X1_HVT U454 ( .A1(n721), .A2(n509), .S0(n474), .Y(n608) );
  INVX0_HVT U455 ( .A(n443), .Y(n721) );
  NBUFFX2_HVT U456 ( .A(n364), .Y(n446) );
  MUX41X1_HVT U457 ( .A1(n606), .A3(n610), .A2(n605), .A4(n609), .S0(in[0]), 
        .S1(n434), .Y(n604) );
  MUX41X1_HVT U458 ( .A1(n705), .A3(n534), .A2(n335), .A4(n505), .S0(n450), 
        .S1(n416), .Y(n605) );
  INVX1_HVT U459 ( .A(n545), .Y(n514) );
  AND2X1_HVT U460 ( .A1(n316), .A2(n694), .Y(n454) );
  NBUFFX2_HVT U461 ( .A(n744), .Y(n481) );
  NBUFFX2_HVT U462 ( .A(n744), .Y(n482) );
  NBUFFX2_HVT U463 ( .A(n744), .Y(n483) );
  MUX21X1_HVT U464 ( .A1(n519), .A2(n376), .S0(n494), .Y(n698) );
  AND2X1_HVT U465 ( .A1(n264), .A2(n677), .Y(n455) );
  MUX21X1_HVT U466 ( .A1(n478), .A2(n306), .S0(n353), .Y(n646) );
  MUX21X1_HVT U467 ( .A1(n519), .A2(n504), .S0(n410), .Y(n579) );
  NAND2X0_HVT U468 ( .A1(n527), .A2(n342), .Y(n744) );
  MUX21X1_HVT U469 ( .A1(n519), .A2(n446), .S0(n412), .Y(n543) );
  NBUFFX2_HVT U470 ( .A(n747), .Y(n484) );
  MUX21X1_HVT U471 ( .A1(n483), .A2(n398), .S0(n412), .Y(n661) );
  NBUFFX2_HVT U472 ( .A(n747), .Y(n485) );
  MUX21X1_HVT U473 ( .A1(n479), .A2(n306), .S0(n488), .Y(n563) );
  MUX21X1_HVT U474 ( .A1(n483), .A2(n479), .S0(n412), .Y(n737) );
  MUX21X1_HVT U475 ( .A1(n484), .A2(n483), .S0(n302), .Y(n542) );
  NBUFFX2_HVT U476 ( .A(n747), .Y(n486) );
  MUX21X1_HVT U477 ( .A1(n231), .A2(n372), .S0(n392), .Y(n566) );
  MUX21X1_HVT U478 ( .A1(n373), .A2(n484), .S0(n305), .Y(n567) );
  XNOR2X1_HVT U479 ( .A1(n373), .A2(n409), .Y(n457) );
  AND2X1_HVT U480 ( .A1(n353), .A2(n504), .Y(n458) );
  MUX21X1_HVT U481 ( .A1(n486), .A2(n446), .S0(n353), .Y(n546) );
  AND2X1_HVT U482 ( .A1(n372), .A2(n639), .Y(n459) );
  MUX21X1_HVT U483 ( .A1(n398), .A2(n373), .S0(n470), .Y(n628) );
  NBUFFX2_HVT U484 ( .A(n498), .Y(n474) );
  NBUFFX2_HVT U485 ( .A(n498), .Y(n475) );
  NBUFFX2_HVT U486 ( .A(n493), .Y(n472) );
  MUX21X1_HVT U487 ( .A1(n648), .A2(n127), .S0(n470), .Y(n645) );
  MUX21X1_HVT U488 ( .A1(n664), .A2(n477), .S0(n473), .Y(n571) );
  NAND2X0_HVT U489 ( .A1(n343), .A2(n364), .Y(n747) );
  AND2X1_HVT U490 ( .A1(n478), .A2(n445), .Y(n460) );
  NBUFFX2_HVT U491 ( .A(n748), .Y(n487) );
  MUX21X1_HVT U492 ( .A1(n376), .A2(n23), .S0(n474), .Y(n681) );
  MUX21X1_HVT U493 ( .A1(n314), .A2(n303), .S0(n469), .Y(n627) );
  MUX21X1_HVT U494 ( .A1(n477), .A2(n716), .S0(n494), .Y(n700) );
  XOR2X1_HVT U495 ( .A1(n393), .A2(n494), .Y(n708) );
  AND2X1_HVT U496 ( .A1(n479), .A2(n445), .Y(n462) );
  NBUFFX2_HVT U497 ( .A(in[5]), .Y(n493) );
  MUX21X1_HVT U498 ( .A1(n415), .A2(n504), .S0(n410), .Y(n588) );
  INVX1_HVT U499 ( .A(n638), .Y(n464) );
  NBUFFX2_HVT U500 ( .A(in[0]), .Y(n476) );
  MUX21X1_HVT U501 ( .A1(n444), .A2(n447), .S0(n409), .Y(n545) );
  MUX21X1_HVT U502 ( .A1(n372), .A2(n444), .S0(n410), .Y(n722) );
  NAND2X0_HVT U503 ( .A1(n352), .A2(n308), .Y(n739) );
  NAND2X0_HVT U504 ( .A1(n343), .A2(n352), .Y(n748) );
  NBUFFX2_HVT U505 ( .A(n491), .Y(n470) );
  NBUFFX2_HVT U506 ( .A(n491), .Y(n469) );
  XOR2X1_HVT U507 ( .A1(n492), .A2(n416), .Y(n704) );
endmodule

