
module inv_Mix_Column ( in, out1 );
  input [127:0] in;
  output [127:0] out1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616;

  XNOR3X1_HVT U1 ( .A1(n1), .A2(n2), .A3(n3), .Y(out1[9]) );
  XNOR3X1_HVT U2 ( .A1(n4), .A2(n5), .A3(n6), .Y(n3) );
  XNOR3X1_HVT U3 ( .A1(n7), .A2(n8), .A3(n9), .Y(out1[99]) );
  XNOR3X1_HVT U4 ( .A1(n10), .A2(n11), .A3(n12), .Y(n7) );
  XNOR3X1_HVT U5 ( .A1(n13), .A2(n14), .A3(n15), .Y(out1[98]) );
  XNOR3X1_HVT U6 ( .A1(n16), .A2(in[121]), .A3(n17), .Y(n13) );
  XNOR3X1_HVT U7 ( .A1(n18), .A2(n19), .A3(n20), .Y(out1[97]) );
  XNOR3X1_HVT U8 ( .A1(n21), .A2(n22), .A3(n23), .Y(n18) );
  XNOR3X1_HVT U9 ( .A1(n24), .A2(n25), .A3(n26), .Y(out1[96]) );
  XNOR3X1_HVT U10 ( .A1(in[127]), .A2(n27), .A3(n28), .Y(n26) );
  XNOR3X1_HVT U11 ( .A1(n29), .A2(n30), .A3(n31), .Y(out1[95]) );
  XOR3X1_HVT U12 ( .A1(in[86]), .A2(n32), .A3(n33), .Y(n31) );
  XNOR3X1_HVT U13 ( .A1(n34), .A2(n35), .A3(n36), .Y(out1[94]) );
  XNOR3X1_HVT U14 ( .A1(n37), .A2(n30), .A3(n38), .Y(n34) );
  XOR2X1_HVT U15 ( .A1(in[92]), .A2(in[93]), .Y(n30) );
  XNOR3X1_HVT U16 ( .A1(n39), .A2(n40), .A3(n41), .Y(out1[93]) );
  XNOR3X1_HVT U17 ( .A1(in[84]), .A2(n42), .A3(n43), .Y(n39) );
  XOR2X1_HVT U18 ( .A1(n44), .A2(n45), .Y(out1[92]) );
  XNOR3X1_HVT U19 ( .A1(n46), .A2(n47), .A3(n48), .Y(n45) );
  XNOR3X1_HVT U20 ( .A1(n49), .A2(n50), .A3(n40), .Y(n44) );
  XNOR2X1_HVT U21 ( .A1(n51), .A2(n52), .Y(n40) );
  INVX0_HVT U22 ( .A(n53), .Y(n52) );
  XNOR3X1_HVT U23 ( .A1(n54), .A2(n55), .A3(n56), .Y(out1[91]) );
  XNOR3X1_HVT U24 ( .A1(n57), .A2(n58), .A3(n59), .Y(n54) );
  XNOR3X1_HVT U25 ( .A1(n60), .A2(n61), .A3(n62), .Y(out1[90]) );
  XNOR3X1_HVT U26 ( .A1(n63), .A2(in[89]), .A3(n64), .Y(n62) );
  XNOR3X1_HVT U27 ( .A1(n65), .A2(n66), .A3(n67), .Y(out1[8]) );
  XOR2X1_HVT U28 ( .A1(n68), .A2(n69), .Y(n65) );
  XNOR3X1_HVT U29 ( .A1(n70), .A2(n71), .A3(n72), .Y(out1[89]) );
  XNOR3X1_HVT U30 ( .A1(n73), .A2(n74), .A3(n75), .Y(n72) );
  XNOR3X1_HVT U31 ( .A1(n76), .A2(n77), .A3(n78), .Y(out1[88]) );
  XOR2X1_HVT U32 ( .A1(n79), .A2(n80), .Y(n76) );
  INVX0_HVT U33 ( .A(n60), .Y(n79) );
  XNOR3X1_HVT U34 ( .A1(n81), .A2(n82), .A3(n83), .Y(out1[87]) );
  XNOR3X1_HVT U35 ( .A1(in[78]), .A2(n84), .A3(n33), .Y(n83) );
  XOR2X1_HVT U36 ( .A1(n85), .A2(n86), .Y(n33) );
  XNOR3X1_HVT U37 ( .A1(n87), .A2(n88), .A3(n89), .Y(out1[86]) );
  XNOR3X1_HVT U38 ( .A1(n90), .A2(n82), .A3(n36), .Y(n89) );
  XOR2X1_HVT U39 ( .A1(n91), .A2(n92), .Y(n36) );
  XOR2X1_HVT U40 ( .A1(in[84]), .A2(in[85]), .Y(n82) );
  XNOR3X1_HVT U41 ( .A1(n93), .A2(n94), .A3(n95), .Y(out1[85]) );
  XNOR3X1_HVT U42 ( .A1(n96), .A2(n97), .A3(n41), .Y(n95) );
  XNOR2X1_HVT U43 ( .A1(n98), .A2(n99), .Y(n41) );
  INVX0_HVT U44 ( .A(n100), .Y(n97) );
  XOR2X1_HVT U45 ( .A1(n101), .A2(n102), .Y(out1[84]) );
  XNOR3X1_HVT U46 ( .A1(n103), .A2(n94), .A3(n48), .Y(n102) );
  XOR2X1_HVT U47 ( .A1(n104), .A2(n105), .Y(n48) );
  XOR2X1_HVT U48 ( .A1(n106), .A2(n50), .Y(n94) );
  XOR3X1_HVT U49 ( .A1(n107), .A2(n108), .A3(n109), .Y(n101) );
  XNOR3X1_HVT U50 ( .A1(n110), .A2(n111), .A3(n112), .Y(out1[83]) );
  XNOR3X1_HVT U51 ( .A1(n113), .A2(n114), .A3(n56), .Y(n112) );
  XNOR3X1_HVT U52 ( .A1(n115), .A2(n116), .A3(n117), .Y(n56) );
  XNOR3X1_HVT U53 ( .A1(n118), .A2(n119), .A3(n120), .Y(out1[82]) );
  XOR3X1_HVT U54 ( .A1(n121), .A2(in[73]), .A3(n61), .Y(n120) );
  XNOR3X1_HVT U55 ( .A1(n122), .A2(in[81]), .A3(n123), .Y(n61) );
  XNOR3X1_HVT U56 ( .A1(n124), .A2(n125), .A3(n126), .Y(out1[81]) );
  XNOR3X1_HVT U57 ( .A1(n127), .A2(n128), .A3(n71), .Y(n126) );
  XNOR3X1_HVT U58 ( .A1(n129), .A2(n130), .A3(n131), .Y(n71) );
  XOR3X1_HVT U59 ( .A1(n132), .A2(n133), .A3(n134), .Y(out1[80]) );
  XNOR3X1_HVT U60 ( .A1(in[86]), .A2(in[79]), .A3(n78), .Y(n134) );
  XNOR3X1_HVT U61 ( .A1(n135), .A2(in[87]), .A3(n136), .Y(n78) );
  XNOR3X1_HVT U62 ( .A1(n137), .A2(n138), .A3(n139), .Y(out1[7]) );
  XOR3X1_HVT U63 ( .A1(in[30]), .A2(n140), .A3(n141), .Y(n139) );
  XNOR3X1_HVT U64 ( .A1(n142), .A2(n143), .A3(n144), .Y(out1[79]) );
  XNOR3X1_HVT U65 ( .A1(n86), .A2(n145), .A3(n77), .Y(n144) );
  XNOR2X1_HVT U66 ( .A1(in[78]), .A2(in[93]), .Y(n77) );
  XOR2X1_HVT U67 ( .A1(in[68]), .A2(in[71]), .Y(n86) );
  XNOR3X1_HVT U68 ( .A1(n143), .A2(n146), .A3(n147), .Y(out1[78]) );
  XNOR3X1_HVT U69 ( .A1(n91), .A2(in[69]), .A3(n42), .Y(n147) );
  XOR2X1_HVT U70 ( .A1(n107), .A2(n148), .Y(n42) );
  INVX0_HVT U71 ( .A(in[92]), .Y(n148) );
  XOR2X1_HVT U72 ( .A1(n149), .A2(n145), .Y(n91) );
  XOR2X1_HVT U73 ( .A1(in[76]), .A2(in[77]), .Y(n143) );
  XNOR3X1_HVT U74 ( .A1(n150), .A2(n151), .A3(n152), .Y(out1[77]) );
  XNOR3X1_HVT U75 ( .A1(in[68]), .A2(n35), .A3(n99), .Y(n150) );
  XNOR2X1_HVT U76 ( .A1(n108), .A2(n153), .Y(n99) );
  XOR2X1_HVT U77 ( .A1(n53), .A2(n96), .Y(n35) );
  XOR2X1_HVT U78 ( .A1(n154), .A2(n155), .Y(out1[76]) );
  XNOR3X1_HVT U79 ( .A1(n105), .A2(n151), .A3(n156), .Y(n155) );
  XNOR2X1_HVT U80 ( .A1(n49), .A2(n107), .Y(n151) );
  XOR2X1_HVT U81 ( .A1(n157), .A2(in[68]), .Y(n105) );
  XNOR3X1_HVT U82 ( .A1(n51), .A2(n149), .A3(n158), .Y(n154) );
  XNOR3X1_HVT U83 ( .A1(n159), .A2(n160), .A3(n161), .Y(out1[75]) );
  XNOR3X1_HVT U84 ( .A1(n114), .A2(n55), .A3(n115), .Y(n159) );
  XOR2X1_HVT U85 ( .A1(n162), .A2(in[67]), .Y(n115) );
  XNOR2X1_HVT U86 ( .A1(n163), .A2(n164), .Y(n55) );
  XOR3X1_HVT U87 ( .A1(n165), .A2(n166), .A3(n167), .Y(out1[74]) );
  XNOR3X1_HVT U88 ( .A1(n63), .A2(in[73]), .A3(n122), .Y(n167) );
  XNOR2X1_HVT U89 ( .A1(n168), .A2(in[66]), .Y(n122) );
  XNOR2X1_HVT U90 ( .A1(n128), .A2(n74), .Y(n63) );
  XNOR3X1_HVT U91 ( .A1(n169), .A2(n170), .A3(n171), .Y(out1[73]) );
  XNOR3X1_HVT U92 ( .A1(n73), .A2(n128), .A3(n129), .Y(n171) );
  XNOR2X1_HVT U93 ( .A1(n172), .A2(in[65]), .Y(n129) );
  XOR2X1_HVT U94 ( .A1(n165), .A2(n60), .Y(n73) );
  XNOR3X1_HVT U95 ( .A1(n173), .A2(n135), .A3(n174), .Y(out1[72]) );
  XOR2X1_HVT U96 ( .A1(in[64]), .A2(in[69]), .Y(n135) );
  XOR2X1_HVT U97 ( .A1(n29), .A2(n165), .Y(n173) );
  XOR2X1_HVT U98 ( .A1(in[94]), .A2(in[77]), .Y(n29) );
  XNOR3X1_HVT U99 ( .A1(n142), .A2(n175), .A3(n176), .Y(out1[71]) );
  XNOR3X1_HVT U100 ( .A1(n85), .A2(n177), .A3(n133), .Y(n176) );
  XNOR2X1_HVT U101 ( .A1(n145), .A2(in[85]), .Y(n133) );
  XOR2X1_HVT U102 ( .A1(n96), .A2(in[79]), .Y(n85) );
  INVX0_HVT U103 ( .A(in[76]), .Y(n96) );
  XNOR2X1_HVT U104 ( .A1(n84), .A2(n32), .Y(n142) );
  XOR2X1_HVT U105 ( .A1(in[84]), .A2(in[87]), .Y(n32) );
  XNOR2X1_HVT U106 ( .A1(in[92]), .A2(in[95]), .Y(n84) );
  XNOR3X1_HVT U107 ( .A1(n146), .A2(n175), .A3(n178), .Y(out1[70]) );
  XNOR3X1_HVT U108 ( .A1(n92), .A2(in[93]), .A3(n93), .Y(n178) );
  XOR2X1_HVT U109 ( .A1(n149), .A2(in[84]), .Y(n93) );
  XOR2X1_HVT U110 ( .A1(n107), .A2(in[78]), .Y(n92) );
  XOR2X1_HVT U111 ( .A1(in[75]), .A2(in[79]), .Y(n107) );
  XNOR2X1_HVT U112 ( .A1(in[68]), .A2(n153), .Y(n175) );
  XOR2X1_HVT U113 ( .A1(n88), .A2(n38), .Y(n146) );
  XNOR2X1_HVT U114 ( .A1(n50), .A2(in[86]), .Y(n38) );
  INVX0_HVT U115 ( .A(n179), .Y(n50) );
  XOR2X1_HVT U116 ( .A1(n53), .A2(n177), .Y(n88) );
  XNOR3X1_HVT U117 ( .A1(n180), .A2(n181), .A3(n182), .Y(out1[6]) );
  XNOR3X1_HVT U118 ( .A1(in[29]), .A2(n138), .A3(n183), .Y(n182) );
  XOR2X1_HVT U119 ( .A1(in[4]), .A2(in[5]), .Y(n138) );
  XNOR3X1_HVT U120 ( .A1(n184), .A2(n185), .A3(n152), .Y(out1[69]) );
  XOR2X1_HVT U121 ( .A1(n100), .A2(n43), .Y(n152) );
  XNOR2X1_HVT U122 ( .A1(n106), .A2(in[85]), .Y(n43) );
  XOR2X1_HVT U123 ( .A1(n51), .A2(in[93]), .Y(n100) );
  XOR2X1_HVT U124 ( .A1(n57), .A2(in[94]), .Y(n51) );
  XNOR3X1_HVT U125 ( .A1(n87), .A2(in[92]), .A3(n98), .Y(n184) );
  XOR2X1_HVT U126 ( .A1(n49), .A2(in[77]), .Y(n98) );
  XNOR2X1_HVT U127 ( .A1(n114), .A2(in[78]), .Y(n49) );
  XOR2X1_HVT U128 ( .A1(in[74]), .A2(in[79]), .Y(n114) );
  XOR2X1_HVT U129 ( .A1(n179), .A2(in[68]), .Y(n87) );
  XOR2X1_HVT U130 ( .A1(in[83]), .A2(in[87]), .Y(n179) );
  XOR2X1_HVT U131 ( .A1(n186), .A2(n187), .Y(out1[68]) );
  XOR3X1_HVT U132 ( .A1(n185), .A2(n157), .A3(n156), .Y(n187) );
  XOR2X1_HVT U133 ( .A1(n103), .A2(n46), .Y(n156) );
  XOR2X1_HVT U134 ( .A1(n109), .A2(n188), .Y(n46) );
  INVX0_HVT U135 ( .A(in[84]), .Y(n188) );
  XOR2X1_HVT U136 ( .A1(n189), .A2(n37), .Y(n109) );
  XNOR2X1_HVT U137 ( .A1(n47), .A2(in[92]), .Y(n103) );
  XNOR2X1_HVT U138 ( .A1(n164), .A2(in[93]), .Y(n47) );
  XOR2X1_HVT U139 ( .A1(in[89]), .A2(in[94]), .Y(n164) );
  XNOR2X1_HVT U140 ( .A1(n190), .A2(in[69]), .Y(n157) );
  XNOR2X1_HVT U141 ( .A1(n108), .A2(n149), .Y(n185) );
  XOR2X1_HVT U142 ( .A1(in[67]), .A2(in[71]), .Y(n149) );
  XOR2X1_HVT U143 ( .A1(n191), .A2(n145), .Y(n108) );
  XNOR3X1_HVT U144 ( .A1(n53), .A2(n106), .A3(n104), .Y(n186) );
  XOR2X1_HVT U145 ( .A1(n158), .A2(in[76]), .Y(n104) );
  XOR2X1_HVT U146 ( .A1(n163), .A2(in[77]), .Y(n158) );
  XNOR2X1_HVT U147 ( .A1(in[73]), .A2(in[78]), .Y(n163) );
  XNOR2X1_HVT U148 ( .A1(n116), .A2(in[86]), .Y(n106) );
  XOR2X1_HVT U149 ( .A1(in[82]), .A2(in[87]), .Y(n116) );
  XNOR2X1_HVT U150 ( .A1(in[91]), .A2(in[95]), .Y(n53) );
  XNOR3X1_HVT U151 ( .A1(n192), .A2(n110), .A3(n161), .Y(out1[67]) );
  XOR3X1_HVT U152 ( .A1(n59), .A2(n191), .A3(n111), .Y(n161) );
  XNOR2X1_HVT U153 ( .A1(n58), .A2(in[91]), .Y(n111) );
  XNOR2X1_HVT U154 ( .A1(n74), .A2(in[93]), .Y(n58) );
  XOR2X1_HVT U155 ( .A1(in[66]), .A2(in[71]), .Y(n191) );
  XOR2X1_HVT U156 ( .A1(n113), .A2(in[83]), .Y(n59) );
  XOR2X1_HVT U157 ( .A1(n130), .A2(n37), .Y(n113) );
  XNOR2X1_HVT U158 ( .A1(n190), .A2(n189), .Y(n110) );
  XOR2X1_HVT U159 ( .A1(in[81]), .A2(in[86]), .Y(n189) );
  XOR2X1_HVT U160 ( .A1(in[65]), .A2(n145), .Y(n190) );
  XNOR3X1_HVT U161 ( .A1(n57), .A2(n162), .A3(n117), .Y(n192) );
  XNOR2X1_HVT U162 ( .A1(n160), .A2(in[75]), .Y(n117) );
  XOR2X1_HVT U163 ( .A1(n128), .A2(in[77]), .Y(n160) );
  XOR2X1_HVT U164 ( .A1(in[72]), .A2(in[79]), .Y(n128) );
  XOR2X1_HVT U165 ( .A1(n193), .A2(n153), .Y(n162) );
  XNOR2X1_HVT U166 ( .A1(in[90]), .A2(in[95]), .Y(n57) );
  XNOR3X1_HVT U167 ( .A1(n194), .A2(n118), .A3(n166), .Y(out1[66]) );
  XOR3X1_HVT U168 ( .A1(n64), .A2(in[65]), .A3(n119), .Y(n166) );
  XNOR2X1_HVT U169 ( .A1(n60), .A2(in[90]), .Y(n119) );
  XOR2X1_HVT U170 ( .A1(n177), .A2(in[95]), .Y(n60) );
  XNOR2X1_HVT U171 ( .A1(n121), .A2(in[82]), .Y(n64) );
  XOR2X1_HVT U172 ( .A1(n193), .A2(n130), .Y(n118) );
  XOR2X1_HVT U173 ( .A1(in[80]), .A2(in[87]), .Y(n130) );
  XNOR3X1_HVT U174 ( .A1(in[89]), .A2(n168), .A3(n123), .Y(n194) );
  XNOR2X1_HVT U175 ( .A1(n165), .A2(in[74]), .Y(n123) );
  XOR2X1_HVT U176 ( .A1(in[78]), .A2(in[79]), .Y(n165) );
  XNOR3X1_HVT U177 ( .A1(n195), .A2(n124), .A3(n170), .Y(out1[65]) );
  XOR3X1_HVT U178 ( .A1(n75), .A2(n193), .A3(n125), .Y(n170) );
  XNOR2X1_HVT U179 ( .A1(n70), .A2(in[89]), .Y(n125) );
  XOR2X1_HVT U180 ( .A1(n177), .A2(in[93]), .Y(n70) );
  INVX0_HVT U181 ( .A(in[94]), .Y(n177) );
  XOR2X1_HVT U182 ( .A1(in[64]), .A2(in[71]), .Y(n193) );
  XOR2X1_HVT U183 ( .A1(n127), .A2(in[81]), .Y(n75) );
  XOR2X1_HVT U184 ( .A1(n37), .A2(in[86]), .Y(n127) );
  INVX0_HVT U185 ( .A(in[85]), .Y(n37) );
  XOR2X1_HVT U186 ( .A1(n168), .A2(n121), .Y(n124) );
  XOR2X1_HVT U187 ( .A1(in[87]), .A2(in[86]), .Y(n121) );
  XOR2X1_HVT U188 ( .A1(n196), .A2(n145), .Y(n168) );
  XNOR3X1_HVT U189 ( .A1(n74), .A2(n172), .A3(n131), .Y(n195) );
  XOR2X1_HVT U190 ( .A1(n169), .A2(in[73]), .Y(n131) );
  XOR2X1_HVT U191 ( .A1(in[78]), .A2(n90), .Y(n169) );
  XOR2X1_HVT U192 ( .A1(n153), .A2(n145), .Y(n172) );
  INVX0_HVT U193 ( .A(in[70]), .Y(n145) );
  INVX0_HVT U194 ( .A(in[69]), .Y(n153) );
  XOR2X1_HVT U195 ( .A1(in[88]), .A2(in[95]), .Y(n74) );
  XNOR3X1_HVT U196 ( .A1(n197), .A2(n81), .A3(n174), .Y(out1[64]) );
  XNOR3X1_HVT U197 ( .A1(n80), .A2(n196), .A3(n132), .Y(n174) );
  XNOR2X1_HVT U198 ( .A1(in[88]), .A2(in[93]), .Y(n132) );
  INVX0_HVT U199 ( .A(in[71]), .Y(n196) );
  XOR2X1_HVT U200 ( .A1(in[80]), .A2(in[85]), .Y(n80) );
  XOR2X1_HVT U201 ( .A1(in[69]), .A2(in[86]), .Y(n81) );
  XNOR3X1_HVT U202 ( .A1(in[95]), .A2(in[70]), .A3(n136), .Y(n197) );
  XOR2X1_HVT U203 ( .A1(in[72]), .A2(n90), .Y(n136) );
  INVX0_HVT U204 ( .A(in[77]), .Y(n90) );
  XNOR3X1_HVT U205 ( .A1(n198), .A2(n199), .A3(n200), .Y(out1[63]) );
  XOR3X1_HVT U206 ( .A1(in[54]), .A2(n201), .A3(n202), .Y(n200) );
  XNOR3X1_HVT U207 ( .A1(n203), .A2(n204), .A3(n205), .Y(out1[62]) );
  XNOR3X1_HVT U208 ( .A1(n206), .A2(n199), .A3(n207), .Y(n203) );
  XOR2X1_HVT U209 ( .A1(in[60]), .A2(in[61]), .Y(n199) );
  XNOR3X1_HVT U210 ( .A1(n208), .A2(n209), .A3(n210), .Y(out1[61]) );
  XNOR3X1_HVT U211 ( .A1(in[52]), .A2(n211), .A3(n212), .Y(n208) );
  XOR2X1_HVT U212 ( .A1(n213), .A2(n214), .Y(out1[60]) );
  XNOR3X1_HVT U213 ( .A1(n215), .A2(n216), .A3(n217), .Y(n214) );
  XNOR3X1_HVT U214 ( .A1(n218), .A2(n219), .A3(n209), .Y(n213) );
  XNOR2X1_HVT U215 ( .A1(n220), .A2(n221), .Y(n209) );
  INVX0_HVT U216 ( .A(n222), .Y(n221) );
  XNOR3X1_HVT U217 ( .A1(n223), .A2(n224), .A3(n225), .Y(out1[5]) );
  XNOR3X1_HVT U218 ( .A1(n226), .A2(n227), .A3(n228), .Y(n225) );
  INVX0_HVT U219 ( .A(in[28]), .Y(n226) );
  XNOR3X1_HVT U220 ( .A1(n229), .A2(n230), .A3(n231), .Y(out1[59]) );
  XNOR3X1_HVT U221 ( .A1(n232), .A2(n233), .A3(n234), .Y(n229) );
  XNOR3X1_HVT U222 ( .A1(n235), .A2(n236), .A3(n237), .Y(out1[58]) );
  XNOR3X1_HVT U223 ( .A1(n238), .A2(in[57]), .A3(n239), .Y(n237) );
  XNOR3X1_HVT U224 ( .A1(n240), .A2(n241), .A3(n242), .Y(out1[57]) );
  XNOR3X1_HVT U225 ( .A1(n243), .A2(n244), .A3(n245), .Y(n242) );
  XNOR3X1_HVT U226 ( .A1(n246), .A2(n247), .A3(n248), .Y(out1[56]) );
  XOR2X1_HVT U227 ( .A1(n249), .A2(n250), .Y(n246) );
  INVX0_HVT U228 ( .A(n235), .Y(n249) );
  XNOR3X1_HVT U229 ( .A1(n251), .A2(n252), .A3(n253), .Y(out1[55]) );
  XNOR3X1_HVT U230 ( .A1(in[46]), .A2(n254), .A3(n202), .Y(n253) );
  XOR2X1_HVT U231 ( .A1(n255), .A2(n256), .Y(n202) );
  XNOR3X1_HVT U232 ( .A1(n257), .A2(n258), .A3(n259), .Y(out1[54]) );
  XNOR3X1_HVT U233 ( .A1(n260), .A2(n252), .A3(n205), .Y(n259) );
  XOR2X1_HVT U234 ( .A1(n261), .A2(n262), .Y(n205) );
  XOR2X1_HVT U235 ( .A1(in[52]), .A2(in[53]), .Y(n252) );
  XNOR3X1_HVT U236 ( .A1(n263), .A2(n264), .A3(n265), .Y(out1[53]) );
  XNOR3X1_HVT U237 ( .A1(n266), .A2(n267), .A3(n210), .Y(n265) );
  XNOR2X1_HVT U238 ( .A1(n268), .A2(n269), .Y(n210) );
  INVX0_HVT U239 ( .A(n270), .Y(n267) );
  XOR2X1_HVT U240 ( .A1(n271), .A2(n272), .Y(out1[52]) );
  XNOR3X1_HVT U241 ( .A1(n273), .A2(n264), .A3(n217), .Y(n272) );
  XOR2X1_HVT U242 ( .A1(n274), .A2(n275), .Y(n217) );
  XOR2X1_HVT U243 ( .A1(n276), .A2(n219), .Y(n264) );
  XOR3X1_HVT U244 ( .A1(n277), .A2(n278), .A3(n279), .Y(n271) );
  XNOR3X1_HVT U245 ( .A1(n280), .A2(n281), .A3(n282), .Y(out1[51]) );
  XNOR3X1_HVT U246 ( .A1(n283), .A2(n284), .A3(n231), .Y(n282) );
  XNOR3X1_HVT U247 ( .A1(n285), .A2(n286), .A3(n287), .Y(n231) );
  XNOR3X1_HVT U248 ( .A1(n288), .A2(n289), .A3(n290), .Y(out1[50]) );
  XOR3X1_HVT U249 ( .A1(n291), .A2(in[41]), .A3(n236), .Y(n290) );
  XNOR3X1_HVT U250 ( .A1(n292), .A2(in[49]), .A3(n293), .Y(n236) );
  XOR2X1_HVT U251 ( .A1(n294), .A2(n295), .Y(out1[4]) );
  XNOR3X1_HVT U252 ( .A1(n296), .A2(n297), .A3(n298), .Y(n295) );
  XNOR3X1_HVT U253 ( .A1(n299), .A2(n300), .A3(n224), .Y(n294) );
  XOR2X1_HVT U254 ( .A1(n301), .A2(n302), .Y(n224) );
  XNOR3X1_HVT U255 ( .A1(n303), .A2(n304), .A3(n305), .Y(out1[49]) );
  XNOR3X1_HVT U256 ( .A1(n306), .A2(n307), .A3(n241), .Y(n305) );
  XNOR3X1_HVT U257 ( .A1(n308), .A2(n309), .A3(n310), .Y(n241) );
  XOR3X1_HVT U258 ( .A1(n311), .A2(n312), .A3(n313), .Y(out1[48]) );
  XNOR3X1_HVT U259 ( .A1(in[54]), .A2(in[47]), .A3(n248), .Y(n313) );
  XNOR3X1_HVT U260 ( .A1(n314), .A2(in[55]), .A3(n315), .Y(n248) );
  XNOR3X1_HVT U261 ( .A1(n316), .A2(n317), .A3(n318), .Y(out1[47]) );
  XNOR3X1_HVT U262 ( .A1(n256), .A2(n319), .A3(n247), .Y(n318) );
  XNOR2X1_HVT U263 ( .A1(in[46]), .A2(in[61]), .Y(n247) );
  XOR2X1_HVT U264 ( .A1(in[36]), .A2(in[39]), .Y(n256) );
  XNOR3X1_HVT U265 ( .A1(n317), .A2(n320), .A3(n321), .Y(out1[46]) );
  XNOR3X1_HVT U266 ( .A1(n261), .A2(in[37]), .A3(n211), .Y(n321) );
  XOR2X1_HVT U267 ( .A1(n277), .A2(n322), .Y(n211) );
  INVX0_HVT U268 ( .A(in[60]), .Y(n322) );
  XOR2X1_HVT U269 ( .A1(n323), .A2(n319), .Y(n261) );
  XOR2X1_HVT U270 ( .A1(in[44]), .A2(in[45]), .Y(n317) );
  XNOR3X1_HVT U271 ( .A1(n324), .A2(n325), .A3(n326), .Y(out1[45]) );
  XNOR3X1_HVT U272 ( .A1(in[36]), .A2(n204), .A3(n269), .Y(n324) );
  XNOR2X1_HVT U273 ( .A1(n278), .A2(n327), .Y(n269) );
  XOR2X1_HVT U274 ( .A1(n222), .A2(n266), .Y(n204) );
  XOR2X1_HVT U275 ( .A1(n328), .A2(n329), .Y(out1[44]) );
  XNOR3X1_HVT U276 ( .A1(n275), .A2(n325), .A3(n330), .Y(n329) );
  XNOR2X1_HVT U277 ( .A1(n218), .A2(n277), .Y(n325) );
  XOR2X1_HVT U278 ( .A1(n331), .A2(in[36]), .Y(n275) );
  XNOR3X1_HVT U279 ( .A1(n220), .A2(n323), .A3(n332), .Y(n328) );
  XNOR3X1_HVT U280 ( .A1(n333), .A2(n334), .A3(n335), .Y(out1[43]) );
  XNOR3X1_HVT U281 ( .A1(n284), .A2(n230), .A3(n285), .Y(n333) );
  XOR2X1_HVT U282 ( .A1(n336), .A2(in[35]), .Y(n285) );
  XNOR2X1_HVT U283 ( .A1(n337), .A2(n338), .Y(n230) );
  XOR3X1_HVT U284 ( .A1(n339), .A2(n340), .A3(n341), .Y(out1[42]) );
  XNOR3X1_HVT U285 ( .A1(n238), .A2(in[41]), .A3(n292), .Y(n341) );
  XNOR2X1_HVT U286 ( .A1(n342), .A2(in[34]), .Y(n292) );
  XNOR2X1_HVT U287 ( .A1(n307), .A2(n244), .Y(n238) );
  XNOR3X1_HVT U288 ( .A1(n343), .A2(n344), .A3(n345), .Y(out1[41]) );
  XNOR3X1_HVT U289 ( .A1(n243), .A2(n307), .A3(n308), .Y(n345) );
  XNOR2X1_HVT U290 ( .A1(n346), .A2(in[33]), .Y(n308) );
  XOR2X1_HVT U291 ( .A1(n339), .A2(n235), .Y(n243) );
  XNOR3X1_HVT U292 ( .A1(n347), .A2(n314), .A3(n348), .Y(out1[40]) );
  XOR2X1_HVT U293 ( .A1(in[32]), .A2(in[37]), .Y(n314) );
  XOR2X1_HVT U294 ( .A1(n198), .A2(n339), .Y(n347) );
  XOR2X1_HVT U295 ( .A1(in[62]), .A2(in[45]), .Y(n198) );
  XNOR3X1_HVT U296 ( .A1(n349), .A2(n350), .A3(n351), .Y(out1[3]) );
  XOR3X1_HVT U297 ( .A1(n352), .A2(n353), .A3(n354), .Y(n349) );
  XNOR3X1_HVT U298 ( .A1(n316), .A2(n355), .A3(n356), .Y(out1[39]) );
  XNOR3X1_HVT U299 ( .A1(n255), .A2(n357), .A3(n312), .Y(n356) );
  XNOR2X1_HVT U300 ( .A1(n319), .A2(in[53]), .Y(n312) );
  XOR2X1_HVT U301 ( .A1(n266), .A2(in[47]), .Y(n255) );
  INVX0_HVT U302 ( .A(in[44]), .Y(n266) );
  XNOR2X1_HVT U303 ( .A1(n254), .A2(n201), .Y(n316) );
  XOR2X1_HVT U304 ( .A1(in[52]), .A2(in[55]), .Y(n201) );
  XNOR2X1_HVT U305 ( .A1(in[60]), .A2(in[63]), .Y(n254) );
  XNOR3X1_HVT U306 ( .A1(n320), .A2(n355), .A3(n358), .Y(out1[38]) );
  XNOR3X1_HVT U307 ( .A1(n262), .A2(in[61]), .A3(n263), .Y(n358) );
  XOR2X1_HVT U308 ( .A1(n323), .A2(in[52]), .Y(n263) );
  XOR2X1_HVT U309 ( .A1(n277), .A2(in[46]), .Y(n262) );
  XOR2X1_HVT U310 ( .A1(in[43]), .A2(in[47]), .Y(n277) );
  XNOR2X1_HVT U311 ( .A1(in[36]), .A2(n327), .Y(n355) );
  XOR2X1_HVT U312 ( .A1(n258), .A2(n207), .Y(n320) );
  XNOR2X1_HVT U313 ( .A1(n219), .A2(in[54]), .Y(n207) );
  INVX0_HVT U314 ( .A(n359), .Y(n219) );
  XOR2X1_HVT U315 ( .A1(n222), .A2(n357), .Y(n258) );
  XNOR3X1_HVT U316 ( .A1(n360), .A2(n361), .A3(n326), .Y(out1[37]) );
  XOR2X1_HVT U317 ( .A1(n270), .A2(n212), .Y(n326) );
  XNOR2X1_HVT U318 ( .A1(n276), .A2(in[53]), .Y(n212) );
  XOR2X1_HVT U319 ( .A1(n220), .A2(in[61]), .Y(n270) );
  XOR2X1_HVT U320 ( .A1(n232), .A2(in[62]), .Y(n220) );
  XNOR3X1_HVT U321 ( .A1(n257), .A2(in[60]), .A3(n268), .Y(n360) );
  XOR2X1_HVT U322 ( .A1(n218), .A2(in[45]), .Y(n268) );
  XNOR2X1_HVT U323 ( .A1(n284), .A2(in[46]), .Y(n218) );
  XOR2X1_HVT U324 ( .A1(in[42]), .A2(in[47]), .Y(n284) );
  XOR2X1_HVT U325 ( .A1(n359), .A2(in[36]), .Y(n257) );
  XOR2X1_HVT U326 ( .A1(in[51]), .A2(in[55]), .Y(n359) );
  XOR2X1_HVT U327 ( .A1(n362), .A2(n363), .Y(out1[36]) );
  XOR3X1_HVT U328 ( .A1(n361), .A2(n331), .A3(n330), .Y(n363) );
  XOR2X1_HVT U329 ( .A1(n273), .A2(n215), .Y(n330) );
  XOR2X1_HVT U330 ( .A1(n279), .A2(n364), .Y(n215) );
  INVX0_HVT U331 ( .A(in[52]), .Y(n364) );
  XOR2X1_HVT U332 ( .A1(n365), .A2(n206), .Y(n279) );
  XNOR2X1_HVT U333 ( .A1(n216), .A2(in[60]), .Y(n273) );
  XNOR2X1_HVT U334 ( .A1(n338), .A2(in[61]), .Y(n216) );
  XOR2X1_HVT U335 ( .A1(in[57]), .A2(in[62]), .Y(n338) );
  XNOR2X1_HVT U336 ( .A1(n366), .A2(in[37]), .Y(n331) );
  XNOR2X1_HVT U337 ( .A1(n278), .A2(n323), .Y(n361) );
  XOR2X1_HVT U338 ( .A1(in[35]), .A2(in[39]), .Y(n323) );
  XOR2X1_HVT U339 ( .A1(n367), .A2(n319), .Y(n278) );
  XNOR3X1_HVT U340 ( .A1(n222), .A2(n276), .A3(n274), .Y(n362) );
  XOR2X1_HVT U341 ( .A1(n332), .A2(in[44]), .Y(n274) );
  XOR2X1_HVT U342 ( .A1(n337), .A2(in[45]), .Y(n332) );
  XNOR2X1_HVT U343 ( .A1(in[41]), .A2(in[46]), .Y(n337) );
  XNOR2X1_HVT U344 ( .A1(n286), .A2(in[54]), .Y(n276) );
  XOR2X1_HVT U345 ( .A1(in[50]), .A2(in[55]), .Y(n286) );
  XNOR2X1_HVT U346 ( .A1(in[59]), .A2(in[63]), .Y(n222) );
  XNOR3X1_HVT U347 ( .A1(n368), .A2(n280), .A3(n335), .Y(out1[35]) );
  XOR3X1_HVT U348 ( .A1(n234), .A2(n367), .A3(n281), .Y(n335) );
  XNOR2X1_HVT U349 ( .A1(n233), .A2(in[59]), .Y(n281) );
  XNOR2X1_HVT U350 ( .A1(n244), .A2(in[61]), .Y(n233) );
  XOR2X1_HVT U351 ( .A1(in[34]), .A2(in[39]), .Y(n367) );
  XOR2X1_HVT U352 ( .A1(n283), .A2(in[51]), .Y(n234) );
  XOR2X1_HVT U353 ( .A1(n309), .A2(n206), .Y(n283) );
  XNOR2X1_HVT U354 ( .A1(n366), .A2(n365), .Y(n280) );
  XOR2X1_HVT U355 ( .A1(in[49]), .A2(in[54]), .Y(n365) );
  XOR2X1_HVT U356 ( .A1(in[33]), .A2(n319), .Y(n366) );
  XNOR3X1_HVT U357 ( .A1(n232), .A2(n336), .A3(n287), .Y(n368) );
  XNOR2X1_HVT U358 ( .A1(n334), .A2(in[43]), .Y(n287) );
  XOR2X1_HVT U359 ( .A1(n307), .A2(in[45]), .Y(n334) );
  XOR2X1_HVT U360 ( .A1(in[40]), .A2(in[47]), .Y(n307) );
  XOR2X1_HVT U361 ( .A1(n369), .A2(n327), .Y(n336) );
  XNOR2X1_HVT U362 ( .A1(in[58]), .A2(in[63]), .Y(n232) );
  XNOR3X1_HVT U363 ( .A1(n370), .A2(n288), .A3(n340), .Y(out1[34]) );
  XOR3X1_HVT U364 ( .A1(n239), .A2(in[33]), .A3(n289), .Y(n340) );
  XNOR2X1_HVT U365 ( .A1(n235), .A2(in[58]), .Y(n289) );
  XOR2X1_HVT U366 ( .A1(n357), .A2(in[63]), .Y(n235) );
  XNOR2X1_HVT U367 ( .A1(n291), .A2(in[50]), .Y(n239) );
  XOR2X1_HVT U368 ( .A1(n369), .A2(n309), .Y(n288) );
  XOR2X1_HVT U369 ( .A1(in[48]), .A2(in[55]), .Y(n309) );
  XNOR3X1_HVT U370 ( .A1(in[57]), .A2(n342), .A3(n293), .Y(n370) );
  XNOR2X1_HVT U371 ( .A1(n339), .A2(in[42]), .Y(n293) );
  XOR2X1_HVT U372 ( .A1(in[46]), .A2(in[47]), .Y(n339) );
  XNOR3X1_HVT U373 ( .A1(n371), .A2(n303), .A3(n344), .Y(out1[33]) );
  XOR3X1_HVT U374 ( .A1(n245), .A2(n369), .A3(n304), .Y(n344) );
  XNOR2X1_HVT U375 ( .A1(n240), .A2(in[57]), .Y(n304) );
  XOR2X1_HVT U376 ( .A1(n357), .A2(in[61]), .Y(n240) );
  INVX0_HVT U377 ( .A(in[62]), .Y(n357) );
  XOR2X1_HVT U378 ( .A1(in[32]), .A2(in[39]), .Y(n369) );
  XOR2X1_HVT U379 ( .A1(n306), .A2(in[49]), .Y(n245) );
  XOR2X1_HVT U380 ( .A1(n206), .A2(in[54]), .Y(n306) );
  INVX0_HVT U381 ( .A(in[53]), .Y(n206) );
  XOR2X1_HVT U382 ( .A1(n342), .A2(n291), .Y(n303) );
  XOR2X1_HVT U383 ( .A1(in[55]), .A2(in[54]), .Y(n291) );
  XOR2X1_HVT U384 ( .A1(n372), .A2(n319), .Y(n342) );
  XNOR3X1_HVT U385 ( .A1(n244), .A2(n346), .A3(n310), .Y(n371) );
  XOR2X1_HVT U386 ( .A1(n343), .A2(in[41]), .Y(n310) );
  XOR2X1_HVT U387 ( .A1(in[46]), .A2(n260), .Y(n343) );
  XOR2X1_HVT U388 ( .A1(n327), .A2(n319), .Y(n346) );
  INVX0_HVT U389 ( .A(in[38]), .Y(n319) );
  INVX0_HVT U390 ( .A(in[37]), .Y(n327) );
  XOR2X1_HVT U391 ( .A1(in[56]), .A2(in[63]), .Y(n244) );
  XNOR3X1_HVT U392 ( .A1(n373), .A2(n251), .A3(n348), .Y(out1[32]) );
  XNOR3X1_HVT U393 ( .A1(n250), .A2(n372), .A3(n311), .Y(n348) );
  XNOR2X1_HVT U394 ( .A1(in[56]), .A2(in[61]), .Y(n311) );
  INVX0_HVT U395 ( .A(in[39]), .Y(n372) );
  XOR2X1_HVT U396 ( .A1(in[48]), .A2(in[53]), .Y(n250) );
  XOR2X1_HVT U397 ( .A1(in[37]), .A2(in[54]), .Y(n251) );
  XNOR3X1_HVT U398 ( .A1(in[63]), .A2(in[38]), .A3(n315), .Y(n373) );
  XOR2X1_HVT U399 ( .A1(in[40]), .A2(n260), .Y(n315) );
  INVX0_HVT U400 ( .A(in[45]), .Y(n260) );
  XNOR3X1_HVT U401 ( .A1(n374), .A2(n375), .A3(n376), .Y(out1[31]) );
  XNOR3X1_HVT U402 ( .A1(n69), .A2(n377), .A3(n378), .Y(n376) );
  XOR2X1_HVT U403 ( .A1(in[30]), .A2(in[13]), .Y(n69) );
  XOR3X1_HVT U404 ( .A1(n379), .A2(n380), .A3(n381), .Y(out1[30]) );
  XNOR3X1_HVT U405 ( .A1(n375), .A2(in[21]), .A3(n382), .Y(n379) );
  XOR2X1_HVT U406 ( .A1(in[28]), .A2(in[29]), .Y(n375) );
  XNOR3X1_HVT U407 ( .A1(n383), .A2(n384), .A3(n385), .Y(out1[2]) );
  XNOR3X1_HVT U408 ( .A1(n386), .A2(in[25]), .A3(n387), .Y(n383) );
  XNOR3X1_HVT U409 ( .A1(n388), .A2(n389), .A3(n390), .Y(out1[29]) );
  XNOR3X1_HVT U410 ( .A1(n391), .A2(in[20]), .A3(n392), .Y(n388) );
  XOR2X1_HVT U411 ( .A1(n393), .A2(n394), .Y(out1[28]) );
  XNOR3X1_HVT U412 ( .A1(n395), .A2(n389), .A3(n396), .Y(n394) );
  XNOR2X1_HVT U413 ( .A1(n397), .A2(n299), .Y(n389) );
  XNOR3X1_HVT U414 ( .A1(n398), .A2(n399), .A3(n400), .Y(n393) );
  XNOR3X1_HVT U415 ( .A1(n401), .A2(n402), .A3(n403), .Y(out1[27]) );
  XNOR3X1_HVT U416 ( .A1(n353), .A2(n404), .A3(n405), .Y(n401) );
  XNOR3X1_HVT U417 ( .A1(n406), .A2(n407), .A3(n408), .Y(out1[26]) );
  XNOR3X1_HVT U418 ( .A1(n409), .A2(n410), .A3(n411), .Y(n406) );
  XNOR3X1_HVT U419 ( .A1(n412), .A2(n413), .A3(n414), .Y(out1[25]) );
  XNOR3X1_HVT U420 ( .A1(n415), .A2(n416), .A3(n1), .Y(n412) );
  XOR2X1_HVT U421 ( .A1(n417), .A2(n410), .Y(n1) );
  INVX0_HVT U422 ( .A(n66), .Y(n417) );
  XNOR3X1_HVT U423 ( .A1(n418), .A2(n419), .A3(n420), .Y(out1[24]) );
  XNOR2X1_HVT U424 ( .A1(n410), .A2(n421), .Y(n418) );
  XNOR3X1_HVT U425 ( .A1(n422), .A2(n423), .A3(n424), .Y(out1[23]) );
  XNOR3X1_HVT U426 ( .A1(in[14]), .A2(n425), .A3(n374), .Y(n424) );
  XOR2X1_HVT U427 ( .A1(n426), .A2(n140), .Y(n374) );
  XOR2X1_HVT U428 ( .A1(in[12]), .A2(in[15]), .Y(n140) );
  XNOR3X1_HVT U429 ( .A1(n381), .A2(n423), .A3(n427), .Y(out1[22]) );
  XNOR3X1_HVT U430 ( .A1(n428), .A2(in[13]), .A3(n223), .Y(n427) );
  XOR2X1_HVT U431 ( .A1(n399), .A2(in[4]), .Y(n223) );
  XOR2X1_HVT U432 ( .A1(in[20]), .A2(in[21]), .Y(n423) );
  XOR2X1_HVT U433 ( .A1(n429), .A2(n181), .Y(n381) );
  XOR2X1_HVT U434 ( .A1(n430), .A2(in[14]), .Y(n181) );
  XNOR3X1_HVT U435 ( .A1(n431), .A2(n432), .A3(n390), .Y(out1[21]) );
  XNOR2X1_HVT U436 ( .A1(n433), .A2(n227), .Y(n390) );
  XNOR2X1_HVT U437 ( .A1(n398), .A2(in[13]), .Y(n227) );
  XNOR3X1_HVT U438 ( .A1(in[12]), .A2(n180), .A3(n434), .Y(n431) );
  XNOR2X1_HVT U439 ( .A1(n302), .A2(in[20]), .Y(n180) );
  XOR2X1_HVT U440 ( .A1(n435), .A2(n436), .Y(out1[20]) );
  XOR3X1_HVT U441 ( .A1(n432), .A2(n437), .A3(n396), .Y(n436) );
  XNOR2X1_HVT U442 ( .A1(n297), .A2(n438), .Y(n396) );
  XOR2X1_HVT U443 ( .A1(n439), .A2(in[12]), .Y(n297) );
  XNOR2X1_HVT U444 ( .A1(n300), .A2(n399), .Y(n432) );
  XNOR3X1_HVT U445 ( .A1(n440), .A2(n301), .A3(n441), .Y(n435) );
  XNOR3X1_HVT U446 ( .A1(n442), .A2(n443), .A3(n444), .Y(out1[1]) );
  XOR3X1_HVT U447 ( .A1(n445), .A2(n413), .A3(n6), .Y(n444) );
  XOR3X1_HVT U448 ( .A1(n446), .A2(n447), .A3(n416), .Y(n6) );
  XNOR2X1_HVT U449 ( .A1(n448), .A2(in[17]), .Y(n416) );
  XNOR3X1_HVT U450 ( .A1(n449), .A2(n450), .A3(n403), .Y(out1[19]) );
  XOR3X1_HVT U451 ( .A1(n354), .A2(n451), .A3(n452), .Y(n403) );
  XOR2X1_HVT U452 ( .A1(n453), .A2(in[11]), .Y(n354) );
  XNOR3X1_HVT U453 ( .A1(n454), .A2(n350), .A3(n455), .Y(n449) );
  XNOR2X1_HVT U454 ( .A1(n456), .A2(n457), .Y(n350) );
  XNOR3X1_HVT U455 ( .A1(n458), .A2(n408), .A3(n459), .Y(out1[18]) );
  XNOR3X1_HVT U456 ( .A1(n387), .A2(in[9]), .A3(n460), .Y(n459) );
  XNOR2X1_HVT U457 ( .A1(n461), .A2(n447), .Y(n387) );
  XNOR3X1_HVT U458 ( .A1(n384), .A2(in[17]), .A3(n462), .Y(n408) );
  XNOR2X1_HVT U459 ( .A1(n66), .A2(in[10]), .Y(n384) );
  XNOR3X1_HVT U460 ( .A1(n463), .A2(n443), .A3(n414), .Y(out1[17]) );
  XNOR3X1_HVT U461 ( .A1(n4), .A2(n461), .A3(n442), .Y(n414) );
  XNOR2X1_HVT U462 ( .A1(n2), .A2(in[9]), .Y(n442) );
  XNOR2X1_HVT U463 ( .A1(in[14]), .A2(in[13]), .Y(n2) );
  XNOR2X1_HVT U464 ( .A1(n445), .A2(in[1]), .Y(n4) );
  XOR2X1_HVT U465 ( .A1(n464), .A2(in[6]), .Y(n445) );
  XNOR2X1_HVT U466 ( .A1(n458), .A2(n386), .Y(n443) );
  XNOR3X1_HVT U467 ( .A1(n448), .A2(n5), .A3(n446), .Y(n463) );
  XOR2X1_HVT U468 ( .A1(n415), .A2(in[25]), .Y(n446) );
  XNOR2X1_HVT U469 ( .A1(in[30]), .A2(in[29]), .Y(n415) );
  XOR2X1_HVT U470 ( .A1(in[21]), .A2(in[22]), .Y(n448) );
  XNOR3X1_HVT U471 ( .A1(n465), .A2(n137), .A3(n420), .Y(out1[16]) );
  XNOR3X1_HVT U472 ( .A1(n68), .A2(in[23]), .A3(n466), .Y(n420) );
  XOR2X1_HVT U473 ( .A1(in[0]), .A2(in[5]), .Y(n68) );
  XOR2X1_HVT U474 ( .A1(in[21]), .A2(in[6]), .Y(n137) );
  XNOR3X1_HVT U475 ( .A1(in[22]), .A2(in[15]), .A3(n467), .Y(n465) );
  XNOR3X1_HVT U476 ( .A1(n419), .A2(n468), .A3(n469), .Y(out1[15]) );
  XNOR3X1_HVT U477 ( .A1(n470), .A2(n426), .A3(n141), .Y(n469) );
  XOR2X1_HVT U478 ( .A1(n378), .A2(n425), .Y(n141) );
  XOR2X1_HVT U479 ( .A1(in[28]), .A2(in[31]), .Y(n425) );
  XNOR2X1_HVT U480 ( .A1(in[20]), .A2(in[23]), .Y(n378) );
  XOR2X1_HVT U481 ( .A1(in[4]), .A2(in[7]), .Y(n426) );
  XOR2X1_HVT U482 ( .A1(in[14]), .A2(in[29]), .Y(n419) );
  XNOR3X1_HVT U483 ( .A1(n391), .A2(n468), .A3(n471), .Y(out1[14]) );
  XNOR3X1_HVT U484 ( .A1(in[5]), .A2(n429), .A3(n183), .Y(n471) );
  XNOR2X1_HVT U485 ( .A1(n382), .A2(n428), .Y(n183) );
  XOR2X1_HVT U486 ( .A1(n299), .A2(in[30]), .Y(n428) );
  XOR2X1_HVT U487 ( .A1(n399), .A2(n377), .Y(n382) );
  XOR2X1_HVT U488 ( .A1(in[19]), .A2(in[23]), .Y(n399) );
  XOR2X1_HVT U489 ( .A1(n302), .A2(n470), .Y(n429) );
  XOR2X1_HVT U490 ( .A1(in[12]), .A2(in[13]), .Y(n468) );
  XOR2X1_HVT U491 ( .A1(n430), .A2(in[28]), .Y(n391) );
  INVX0_HVT U492 ( .A(n440), .Y(n430) );
  XNOR3X1_HVT U493 ( .A1(n433), .A2(n472), .A3(n473), .Y(out1[13]) );
  XNOR3X1_HVT U494 ( .A1(n474), .A2(n380), .A3(n228), .Y(n473) );
  XNOR2X1_HVT U495 ( .A1(n434), .A2(n392), .Y(n228) );
  XOR2X1_HVT U496 ( .A1(n300), .A2(in[21]), .Y(n392) );
  XOR2X1_HVT U497 ( .A1(n451), .A2(n377), .Y(n300) );
  XOR2X1_HVT U498 ( .A1(in[18]), .A2(in[23]), .Y(n451) );
  XOR2X1_HVT U499 ( .A1(n397), .A2(in[29]), .Y(n434) );
  XNOR2X1_HVT U500 ( .A1(n299), .A2(n475), .Y(n380) );
  INVX0_HVT U501 ( .A(in[12]), .Y(n475) );
  XOR2X1_HVT U502 ( .A1(in[27]), .A2(in[31]), .Y(n299) );
  XNOR2X1_HVT U503 ( .A1(n301), .A2(in[5]), .Y(n433) );
  XOR2X1_HVT U504 ( .A1(n476), .A2(n470), .Y(n301) );
  XOR2X1_HVT U505 ( .A1(n477), .A2(n478), .Y(out1[12]) );
  XNOR3X1_HVT U506 ( .A1(n472), .A2(n438), .A3(n298), .Y(n478) );
  XOR2X1_HVT U507 ( .A1(n441), .A2(n395), .Y(n298) );
  XOR2X1_HVT U508 ( .A1(n437), .A2(in[20]), .Y(n395) );
  XOR2X1_HVT U509 ( .A1(n457), .A2(in[21]), .Y(n437) );
  XOR2X1_HVT U510 ( .A1(in[17]), .A2(in[22]), .Y(n457) );
  XOR2X1_HVT U511 ( .A1(n400), .A2(in[28]), .Y(n441) );
  XOR2X1_HVT U512 ( .A1(n479), .A2(in[29]), .Y(n400) );
  XOR2X1_HVT U513 ( .A1(n296), .A2(n474), .Y(n438) );
  INVX0_HVT U514 ( .A(in[4]), .Y(n474) );
  XNOR2X1_HVT U515 ( .A1(n456), .A2(n464), .Y(n296) );
  INVX0_HVT U516 ( .A(in[5]), .Y(n464) );
  XOR2X1_HVT U517 ( .A1(in[1]), .A2(n470), .Y(n456) );
  INVX0_HVT U518 ( .A(in[6]), .Y(n470) );
  XOR2X1_HVT U519 ( .A1(n398), .A2(n440), .Y(n472) );
  XNOR2X1_HVT U520 ( .A1(in[11]), .A2(in[15]), .Y(n440) );
  XNOR2X1_HVT U521 ( .A1(n454), .A2(in[14]), .Y(n398) );
  XNOR3X1_HVT U522 ( .A1(n302), .A2(n397), .A3(n439), .Y(n477) );
  XNOR2X1_HVT U523 ( .A1(n480), .A2(in[13]), .Y(n439) );
  XOR2X1_HVT U524 ( .A1(n353), .A2(in[30]), .Y(n397) );
  XNOR2X1_HVT U525 ( .A1(in[26]), .A2(in[31]), .Y(n353) );
  XNOR2X1_HVT U526 ( .A1(in[3]), .A2(in[7]), .Y(n302) );
  XNOR3X1_HVT U527 ( .A1(n481), .A2(n482), .A3(n483), .Y(out1[127]) );
  XNOR3X1_HVT U528 ( .A1(in[118]), .A2(n484), .A3(n485), .Y(n483) );
  XNOR3X1_HVT U529 ( .A1(n486), .A2(n487), .A3(n488), .Y(out1[126]) );
  XNOR3X1_HVT U530 ( .A1(n489), .A2(n482), .A3(n490), .Y(n486) );
  XOR2X1_HVT U531 ( .A1(in[124]), .A2(in[125]), .Y(n482) );
  XNOR3X1_HVT U532 ( .A1(n491), .A2(n492), .A3(n493), .Y(out1[125]) );
  XNOR3X1_HVT U533 ( .A1(in[116]), .A2(n494), .A3(n495), .Y(n491) );
  XOR2X1_HVT U534 ( .A1(n496), .A2(n497), .Y(out1[124]) );
  XNOR3X1_HVT U535 ( .A1(n498), .A2(n499), .A3(n500), .Y(n497) );
  XNOR3X1_HVT U536 ( .A1(n501), .A2(n502), .A3(n492), .Y(n496) );
  XNOR2X1_HVT U537 ( .A1(n503), .A2(n504), .Y(n492) );
  INVX0_HVT U538 ( .A(n505), .Y(n504) );
  XNOR3X1_HVT U539 ( .A1(n506), .A2(n507), .A3(n508), .Y(out1[123]) );
  XOR3X1_HVT U540 ( .A1(n10), .A2(n509), .A3(n510), .Y(n506) );
  XNOR3X1_HVT U541 ( .A1(n511), .A2(n512), .A3(n513), .Y(out1[122]) );
  XOR3X1_HVT U542 ( .A1(in[121]), .A2(n514), .A3(n515), .Y(n511) );
  XNOR3X1_HVT U543 ( .A1(n516), .A2(n517), .A3(n518), .Y(out1[121]) );
  XNOR3X1_HVT U544 ( .A1(n22), .A2(n519), .A3(n520), .Y(n516) );
  XNOR3X1_HVT U545 ( .A1(n521), .A2(n522), .A3(n523), .Y(out1[120]) );
  XNOR2X1_HVT U546 ( .A1(n514), .A2(n524), .Y(n521) );
  XNOR3X1_HVT U547 ( .A1(n402), .A2(n452), .A3(n525), .Y(out1[11]) );
  XNOR3X1_HVT U548 ( .A1(n453), .A2(n454), .A3(n351), .Y(n525) );
  XNOR3X1_HVT U549 ( .A1(n455), .A2(n476), .A3(n405), .Y(n351) );
  XNOR2X1_HVT U550 ( .A1(n450), .A2(in[19]), .Y(n405) );
  XOR2X1_HVT U551 ( .A1(n461), .A2(in[21]), .Y(n450) );
  XOR2X1_HVT U552 ( .A1(in[16]), .A2(in[23]), .Y(n461) );
  XOR2X1_HVT U553 ( .A1(in[2]), .A2(in[7]), .Y(n476) );
  XOR2X1_HVT U554 ( .A1(n404), .A2(in[27]), .Y(n455) );
  XNOR2X1_HVT U555 ( .A1(n413), .A2(in[29]), .Y(n404) );
  XOR2X1_HVT U556 ( .A1(in[10]), .A2(in[15]), .Y(n454) );
  XNOR2X1_HVT U557 ( .A1(n5), .A2(in[13]), .Y(n453) );
  XOR2X1_HVT U558 ( .A1(n352), .A2(in[3]), .Y(n452) );
  XOR2X1_HVT U559 ( .A1(n447), .A2(in[5]), .Y(n352) );
  XOR2X1_HVT U560 ( .A1(in[0]), .A2(in[7]), .Y(n447) );
  XNOR2X1_HVT U561 ( .A1(n479), .A2(n480), .Y(n402) );
  XOR2X1_HVT U562 ( .A1(in[9]), .A2(in[14]), .Y(n480) );
  XOR2X1_HVT U563 ( .A1(n409), .A2(in[30]), .Y(n479) );
  INVX0_HVT U564 ( .A(in[25]), .Y(n409) );
  XNOR3X1_HVT U565 ( .A1(n526), .A2(n527), .A3(n528), .Y(out1[119]) );
  XNOR3X1_HVT U566 ( .A1(in[110]), .A2(n25), .A3(n485), .Y(n528) );
  XNOR2X1_HVT U567 ( .A1(n529), .A2(n530), .Y(n485) );
  XOR2X1_HVT U568 ( .A1(in[101]), .A2(in[118]), .Y(n25) );
  XNOR3X1_HVT U569 ( .A1(n531), .A2(n532), .A3(n533), .Y(out1[118]) );
  XNOR3X1_HVT U570 ( .A1(n534), .A2(n527), .A3(n488), .Y(n533) );
  XOR2X1_HVT U571 ( .A1(n535), .A2(n536), .Y(n488) );
  XOR2X1_HVT U572 ( .A1(in[116]), .A2(in[117]), .Y(n527) );
  XNOR3X1_HVT U573 ( .A1(n537), .A2(n538), .A3(n539), .Y(out1[117]) );
  XNOR3X1_HVT U574 ( .A1(n540), .A2(n541), .A3(n493), .Y(n539) );
  XNOR2X1_HVT U575 ( .A1(n542), .A2(n543), .Y(n493) );
  INVX0_HVT U576 ( .A(n544), .Y(n541) );
  XOR2X1_HVT U577 ( .A1(n545), .A2(n546), .Y(out1[116]) );
  XNOR3X1_HVT U578 ( .A1(n547), .A2(n538), .A3(n500), .Y(n546) );
  XOR2X1_HVT U579 ( .A1(n548), .A2(n549), .Y(n500) );
  XOR2X1_HVT U580 ( .A1(n550), .A2(n502), .Y(n538) );
  XOR3X1_HVT U581 ( .A1(n551), .A2(n552), .A3(n553), .Y(n545) );
  XNOR3X1_HVT U582 ( .A1(n554), .A2(n555), .A3(n508), .Y(out1[115]) );
  XOR3X1_HVT U583 ( .A1(n12), .A2(n556), .A3(n557), .Y(n508) );
  XOR2X1_HVT U584 ( .A1(n558), .A2(in[107]), .Y(n12) );
  XNOR3X1_HVT U585 ( .A1(n559), .A2(n8), .A3(n560), .Y(n554) );
  XNOR2X1_HVT U586 ( .A1(n561), .A2(n562), .Y(n8) );
  XNOR3X1_HVT U587 ( .A1(n563), .A2(n513), .A3(n564), .Y(out1[114]) );
  XNOR3X1_HVT U588 ( .A1(n17), .A2(in[105]), .A3(n565), .Y(n564) );
  XNOR2X1_HVT U589 ( .A1(n566), .A2(n567), .Y(n17) );
  XNOR3X1_HVT U590 ( .A1(n14), .A2(in[113]), .A3(n568), .Y(n513) );
  XOR2X1_HVT U591 ( .A1(n569), .A2(in[106]), .Y(n14) );
  XNOR3X1_HVT U592 ( .A1(n570), .A2(n518), .A3(n571), .Y(out1[113]) );
  XOR3X1_HVT U593 ( .A1(n19), .A2(n572), .A3(n573), .Y(n571) );
  XNOR2X1_HVT U594 ( .A1(n563), .A2(n16), .Y(n19) );
  XOR3X1_HVT U595 ( .A1(n23), .A2(n566), .A3(n574), .Y(n518) );
  XOR2X1_HVT U596 ( .A1(n575), .A2(in[105]), .Y(n23) );
  XNOR3X1_HVT U597 ( .A1(n576), .A2(n577), .A3(n523), .Y(out1[112]) );
  XNOR3X1_HVT U598 ( .A1(n24), .A2(in[119]), .A3(n578), .Y(n523) );
  XOR2X1_HVT U599 ( .A1(in[104]), .A2(in[109]), .Y(n24) );
  XNOR3X1_HVT U600 ( .A1(in[118]), .A2(in[111]), .A3(n579), .Y(n576) );
  XNOR3X1_HVT U601 ( .A1(n580), .A2(n581), .A3(n582), .Y(out1[111]) );
  XNOR3X1_HVT U602 ( .A1(n529), .A2(n27), .A3(n522), .Y(n582) );
  XNOR2X1_HVT U603 ( .A1(n583), .A2(in[125]), .Y(n522) );
  XOR2X1_HVT U604 ( .A1(in[100]), .A2(n584), .Y(n529) );
  XNOR3X1_HVT U605 ( .A1(n581), .A2(n585), .A3(n586), .Y(out1[110]) );
  XNOR3X1_HVT U606 ( .A1(n535), .A2(in[101]), .A3(n494), .Y(n586) );
  XNOR2X1_HVT U607 ( .A1(n551), .A2(in[124]), .Y(n494) );
  XOR2X1_HVT U608 ( .A1(n587), .A2(n27), .Y(n535) );
  XOR2X1_HVT U609 ( .A1(in[108]), .A2(in[109]), .Y(n581) );
  XNOR3X1_HVT U610 ( .A1(n407), .A2(n462), .A3(n588), .Y(out1[10]) );
  XNOR3X1_HVT U611 ( .A1(n66), .A2(in[9]), .A3(n385), .Y(n588) );
  XNOR3X1_HVT U612 ( .A1(n460), .A2(in[1]), .A3(n411), .Y(n385) );
  XOR2X1_HVT U613 ( .A1(n458), .A2(in[18]), .Y(n411) );
  XOR2X1_HVT U614 ( .A1(in[23]), .A2(n377), .Y(n458) );
  INVX0_HVT U615 ( .A(in[22]), .Y(n377) );
  XOR2X1_HVT U616 ( .A1(n410), .A2(in[26]), .Y(n460) );
  XNOR2X1_HVT U617 ( .A1(in[30]), .A2(in[31]), .Y(n410) );
  XNOR2X1_HVT U618 ( .A1(in[14]), .A2(in[15]), .Y(n66) );
  XOR2X1_HVT U619 ( .A1(n386), .A2(in[2]), .Y(n462) );
  XOR2X1_HVT U620 ( .A1(in[7]), .A2(in[6]), .Y(n386) );
  XOR2X1_HVT U621 ( .A1(n413), .A2(n5), .Y(n407) );
  XOR2X1_HVT U622 ( .A1(in[8]), .A2(in[15]), .Y(n5) );
  XOR2X1_HVT U623 ( .A1(in[24]), .A2(in[31]), .Y(n413) );
  XNOR3X1_HVT U624 ( .A1(n589), .A2(n590), .A3(n591), .Y(out1[109]) );
  XNOR3X1_HVT U625 ( .A1(in[100]), .A2(n487), .A3(n543), .Y(n589) );
  XNOR2X1_HVT U626 ( .A1(n552), .A2(n592), .Y(n543) );
  XOR2X1_HVT U627 ( .A1(n505), .A2(n540), .Y(n487) );
  INVX0_HVT U628 ( .A(in[108]), .Y(n540) );
  XOR2X1_HVT U629 ( .A1(n593), .A2(n594), .Y(out1[108]) );
  XNOR3X1_HVT U630 ( .A1(n549), .A2(n590), .A3(n595), .Y(n594) );
  XNOR2X1_HVT U631 ( .A1(n501), .A2(n551), .Y(n590) );
  XOR2X1_HVT U632 ( .A1(n596), .A2(in[100]), .Y(n549) );
  XNOR3X1_HVT U633 ( .A1(n503), .A2(n587), .A3(n597), .Y(n593) );
  XNOR3X1_HVT U634 ( .A1(n507), .A2(n557), .A3(n598), .Y(out1[107]) );
  XNOR3X1_HVT U635 ( .A1(n558), .A2(n555), .A3(n9), .Y(n598) );
  XNOR3X1_HVT U636 ( .A1(n560), .A2(n599), .A3(n510), .Y(n9) );
  XNOR2X1_HVT U637 ( .A1(n559), .A2(in[115]), .Y(n510) );
  XOR2X1_HVT U638 ( .A1(n566), .A2(in[117]), .Y(n559) );
  XOR2X1_HVT U639 ( .A1(in[112]), .A2(in[119]), .Y(n566) );
  XOR2X1_HVT U640 ( .A1(n509), .A2(in[123]), .Y(n560) );
  XNOR2X1_HVT U641 ( .A1(n22), .A2(in[125]), .Y(n509) );
  XOR2X1_HVT U642 ( .A1(n572), .A2(n534), .Y(n558) );
  XOR2X1_HVT U643 ( .A1(n11), .A2(in[99]), .Y(n557) );
  XOR2X1_HVT U644 ( .A1(n567), .A2(in[101]), .Y(n11) );
  XNOR2X1_HVT U645 ( .A1(n600), .A2(n601), .Y(n507) );
  XNOR3X1_HVT U646 ( .A1(n512), .A2(n568), .A3(n602), .Y(out1[106]) );
  XNOR3X1_HVT U647 ( .A1(n569), .A2(n603), .A3(n15), .Y(n602) );
  XNOR3X1_HVT U648 ( .A1(n565), .A2(in[97]), .A3(n515), .Y(n15) );
  XOR2X1_HVT U649 ( .A1(n563), .A2(in[114]), .Y(n515) );
  XOR2X1_HVT U650 ( .A1(n604), .A2(in[118]), .Y(n563) );
  INVX0_HVT U651 ( .A(in[119]), .Y(n604) );
  XOR2X1_HVT U652 ( .A1(n514), .A2(in[122]), .Y(n565) );
  XOR2X1_HVT U653 ( .A1(n16), .A2(in[98]), .Y(n568) );
  XNOR2X1_HVT U654 ( .A1(n584), .A2(in[102]), .Y(n16) );
  XOR2X1_HVT U655 ( .A1(n22), .A2(n572), .Y(n512) );
  XOR2X1_HVT U656 ( .A1(in[120]), .A2(in[127]), .Y(n22) );
  XNOR3X1_HVT U657 ( .A1(n517), .A2(n574), .A3(n605), .Y(out1[105]) );
  XNOR3X1_HVT U658 ( .A1(n575), .A2(n572), .A3(n20), .Y(n605) );
  XNOR3X1_HVT U659 ( .A1(n573), .A2(n567), .A3(n520), .Y(n20) );
  XOR2X1_HVT U660 ( .A1(n570), .A2(in[113]), .Y(n520) );
  XOR2X1_HVT U661 ( .A1(n489), .A2(in[118]), .Y(n570) );
  XOR2X1_HVT U662 ( .A1(in[96]), .A2(in[103]), .Y(n567) );
  XNOR2X1_HVT U663 ( .A1(n519), .A2(in[121]), .Y(n573) );
  XOR2X1_HVT U664 ( .A1(in[126]), .A2(in[125]), .Y(n519) );
  XOR2X1_HVT U665 ( .A1(in[104]), .A2(in[111]), .Y(n572) );
  XOR2X1_HVT U666 ( .A1(n583), .A2(in[109]), .Y(n575) );
  XOR2X1_HVT U667 ( .A1(n21), .A2(in[97]), .Y(n574) );
  XNOR2X1_HVT U668 ( .A1(n592), .A2(in[102]), .Y(n21) );
  XNOR2X1_HVT U669 ( .A1(n514), .A2(n569), .Y(n517) );
  XNOR2X1_HVT U670 ( .A1(in[126]), .A2(in[127]), .Y(n514) );
  XNOR3X1_HVT U671 ( .A1(n606), .A2(n569), .A3(n28), .Y(out1[104]) );
  XNOR3X1_HVT U672 ( .A1(n579), .A2(n584), .A3(n524), .Y(n28) );
  XOR2X1_HVT U673 ( .A1(in[112]), .A2(in[117]), .Y(n524) );
  INVX0_HVT U674 ( .A(in[103]), .Y(n584) );
  XNOR2X1_HVT U675 ( .A1(in[120]), .A2(in[125]), .Y(n579) );
  XNOR2X1_HVT U676 ( .A1(n583), .A2(in[111]), .Y(n569) );
  XOR2X1_HVT U677 ( .A1(n481), .A2(n578), .Y(n606) );
  XOR2X1_HVT U678 ( .A1(in[96]), .A2(in[101]), .Y(n578) );
  XNOR2X1_HVT U679 ( .A1(in[126]), .A2(n534), .Y(n481) );
  INVX0_HVT U680 ( .A(in[109]), .Y(n534) );
  XNOR3X1_HVT U681 ( .A1(n580), .A2(n607), .A3(n608), .Y(out1[103]) );
  XNOR3X1_HVT U682 ( .A1(n530), .A2(in[126]), .A3(n577), .Y(n608) );
  XOR2X1_HVT U683 ( .A1(n27), .A2(n489), .Y(n577) );
  INVX0_HVT U684 ( .A(in[117]), .Y(n489) );
  XOR2X1_HVT U685 ( .A1(in[108]), .A2(in[111]), .Y(n530) );
  XOR2X1_HVT U686 ( .A1(n526), .A2(n484), .Y(n580) );
  XOR2X1_HVT U687 ( .A1(in[116]), .A2(in[119]), .Y(n484) );
  XOR2X1_HVT U688 ( .A1(in[124]), .A2(in[127]), .Y(n526) );
  XNOR3X1_HVT U689 ( .A1(n585), .A2(n607), .A3(n609), .Y(out1[102]) );
  XNOR3X1_HVT U690 ( .A1(n536), .A2(in[125]), .A3(n537), .Y(n609) );
  XOR2X1_HVT U691 ( .A1(n587), .A2(in[116]), .Y(n537) );
  XOR2X1_HVT U692 ( .A1(n551), .A2(in[110]), .Y(n536) );
  XOR2X1_HVT U693 ( .A1(in[107]), .A2(in[111]), .Y(n551) );
  XNOR2X1_HVT U694 ( .A1(in[100]), .A2(n592), .Y(n607) );
  INVX0_HVT U695 ( .A(in[101]), .Y(n592) );
  XOR2X1_HVT U696 ( .A1(n532), .A2(n490), .Y(n585) );
  XNOR2X1_HVT U697 ( .A1(n502), .A2(in[118]), .Y(n490) );
  INVX0_HVT U698 ( .A(n610), .Y(n502) );
  XNOR2X1_HVT U699 ( .A1(n505), .A2(in[126]), .Y(n532) );
  XNOR3X1_HVT U700 ( .A1(n611), .A2(n612), .A3(n591), .Y(out1[101]) );
  XOR2X1_HVT U701 ( .A1(n544), .A2(n495), .Y(n591) );
  XNOR2X1_HVT U702 ( .A1(n550), .A2(in[117]), .Y(n495) );
  XOR2X1_HVT U703 ( .A1(n503), .A2(in[125]), .Y(n544) );
  XNOR2X1_HVT U704 ( .A1(n10), .A2(in[126]), .Y(n503) );
  XOR2X1_HVT U705 ( .A1(in[122]), .A2(in[127]), .Y(n10) );
  XNOR3X1_HVT U706 ( .A1(n531), .A2(in[124]), .A3(n542), .Y(n611) );
  XOR2X1_HVT U707 ( .A1(n501), .A2(in[109]), .Y(n542) );
  XOR2X1_HVT U708 ( .A1(n555), .A2(n583), .Y(n501) );
  INVX0_HVT U709 ( .A(in[110]), .Y(n583) );
  XOR2X1_HVT U710 ( .A1(in[106]), .A2(in[111]), .Y(n555) );
  XOR2X1_HVT U711 ( .A1(n610), .A2(in[100]), .Y(n531) );
  XOR2X1_HVT U712 ( .A1(in[115]), .A2(in[119]), .Y(n610) );
  XOR2X1_HVT U713 ( .A1(n613), .A2(n614), .Y(out1[100]) );
  XOR3X1_HVT U714 ( .A1(n612), .A2(n596), .A3(n595), .Y(n614) );
  XOR2X1_HVT U715 ( .A1(n547), .A2(n498), .Y(n595) );
  XOR2X1_HVT U716 ( .A1(n553), .A2(n615), .Y(n498) );
  INVX0_HVT U717 ( .A(in[116]), .Y(n615) );
  XOR2X1_HVT U718 ( .A1(n561), .A2(in[117]), .Y(n553) );
  XNOR2X1_HVT U719 ( .A1(in[113]), .A2(in[118]), .Y(n561) );
  XNOR2X1_HVT U720 ( .A1(n499), .A2(in[124]), .Y(n547) );
  XNOR2X1_HVT U721 ( .A1(n601), .A2(in[125]), .Y(n499) );
  XOR2X1_HVT U722 ( .A1(in[121]), .A2(in[126]), .Y(n601) );
  XOR2X1_HVT U723 ( .A1(n562), .A2(in[101]), .Y(n596) );
  XOR2X1_HVT U724 ( .A1(in[97]), .A2(in[102]), .Y(n562) );
  XNOR2X1_HVT U725 ( .A1(n552), .A2(n587), .Y(n612) );
  XOR2X1_HVT U726 ( .A1(in[99]), .A2(in[103]), .Y(n587) );
  XOR2X1_HVT U727 ( .A1(n599), .A2(n27), .Y(n552) );
  INVX0_HVT U728 ( .A(in[102]), .Y(n27) );
  XOR2X1_HVT U729 ( .A1(in[98]), .A2(in[103]), .Y(n599) );
  XNOR3X1_HVT U730 ( .A1(n505), .A2(n550), .A3(n548), .Y(n613) );
  XOR2X1_HVT U731 ( .A1(n597), .A2(in[108]), .Y(n548) );
  XOR2X1_HVT U732 ( .A1(n600), .A2(in[109]), .Y(n597) );
  XOR2X1_HVT U733 ( .A1(n603), .A2(in[110]), .Y(n600) );
  INVX0_HVT U734 ( .A(in[105]), .Y(n603) );
  XNOR2X1_HVT U735 ( .A1(n556), .A2(in[118]), .Y(n550) );
  XOR2X1_HVT U736 ( .A1(in[114]), .A2(in[119]), .Y(n556) );
  XNOR2X1_HVT U737 ( .A1(in[123]), .A2(in[127]), .Y(n505) );
  XNOR3X1_HVT U738 ( .A1(n466), .A2(n422), .A3(n616), .Y(out1[0]) );
  XNOR3X1_HVT U739 ( .A1(in[6]), .A2(in[31]), .A3(n67), .Y(n616) );
  XNOR3X1_HVT U740 ( .A1(n467), .A2(in[7]), .A3(n421), .Y(n67) );
  XOR2X1_HVT U741 ( .A1(in[16]), .A2(in[21]), .Y(n421) );
  XNOR2X1_HVT U742 ( .A1(in[24]), .A2(in[29]), .Y(n467) );
  XOR2X1_HVT U743 ( .A1(in[22]), .A2(in[5]), .Y(n422) );
  XOR2X1_HVT U744 ( .A1(in[8]), .A2(in[13]), .Y(n466) );
endmodule

