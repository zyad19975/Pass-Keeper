
module inv_round ( in, last, keyin, out );
  input [127:0] in;
  input [127:0] keyin;
  output [127:0] out;
  input last;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;
  wire   [127:0] sr_out;
  wire   [127:0] sb_out;
  wire   [127:0] oout;
  wire   [127:0] mc_out;

  AO22X1_HVT U2 ( .A1(n68), .A2(n94), .A3(mc_out[9]), .A4(n107), .Y(out[9]) );
  AO22X1_HVT U3 ( .A1(n67), .A2(n95), .A3(mc_out[99]), .A4(n107), .Y(out[99])
         );
  AO22X1_HVT U4 ( .A1(n64), .A2(n95), .A3(mc_out[98]), .A4(n107), .Y(out[98])
         );
  AO22X1_HVT U5 ( .A1(n95), .A2(n24), .A3(mc_out[97]), .A4(n107), .Y(out[97])
         );
  AO22X1_HVT U6 ( .A1(n30), .A2(n96), .A3(mc_out[96]), .A4(n107), .Y(out[96])
         );
  AO22X1_HVT U7 ( .A1(n32), .A2(n96), .A3(mc_out[95]), .A4(n107), .Y(out[95])
         );
  AO22X1_HVT U8 ( .A1(n2), .A2(n96), .A3(mc_out[94]), .A4(n107), .Y(out[94])
         );
  AO22X1_HVT U9 ( .A1(n40), .A2(n96), .A3(mc_out[93]), .A4(n107), .Y(out[93])
         );
  AO22X1_HVT U10 ( .A1(oout[92]), .A2(n96), .A3(mc_out[92]), .A4(n107), .Y(
        out[92]) );
  AO22X1_HVT U11 ( .A1(n33), .A2(n96), .A3(mc_out[91]), .A4(n107), .Y(out[91])
         );
  AO22X1_HVT U12 ( .A1(n28), .A2(n96), .A3(mc_out[90]), .A4(n107), .Y(out[90])
         );
  AO22X1_HVT U13 ( .A1(n96), .A2(n10), .A3(mc_out[8]), .A4(n107), .Y(out[8])
         );
  AO22X1_HVT U14 ( .A1(n22), .A2(n96), .A3(mc_out[89]), .A4(n108), .Y(out[89])
         );
  AO22X1_HVT U15 ( .A1(n31), .A2(n96), .A3(mc_out[88]), .A4(n108), .Y(out[88])
         );
  AO22X1_HVT U16 ( .A1(n88), .A2(n96), .A3(mc_out[87]), .A4(n108), .Y(out[87])
         );
  AO22X1_HVT U17 ( .A1(oout[86]), .A2(n96), .A3(mc_out[86]), .A4(n108), .Y(
        out[86]) );
  AO22X1_HVT U18 ( .A1(n50), .A2(n96), .A3(mc_out[85]), .A4(n108), .Y(out[85])
         );
  AO22X1_HVT U19 ( .A1(oout[84]), .A2(n96), .A3(mc_out[84]), .A4(n108), .Y(
        out[84]) );
  AO22X1_HVT U20 ( .A1(oout[83]), .A2(n96), .A3(mc_out[83]), .A4(n108), .Y(
        out[83]) );
  AO22X1_HVT U21 ( .A1(n42), .A2(n97), .A3(mc_out[82]), .A4(n108), .Y(out[82])
         );
  AO22X1_HVT U22 ( .A1(n97), .A2(n78), .A3(mc_out[81]), .A4(n108), .Y(out[81])
         );
  AO22X1_HVT U23 ( .A1(n46), .A2(n97), .A3(mc_out[80]), .A4(n108), .Y(out[80])
         );
  AO22X1_HVT U24 ( .A1(oout[7]), .A2(n97), .A3(mc_out[7]), .A4(n108), .Y(
        out[7]) );
  AO22X1_HVT U25 ( .A1(n43), .A2(n97), .A3(mc_out[79]), .A4(n108), .Y(out[79])
         );
  AO22X1_HVT U26 ( .A1(n9), .A2(n97), .A3(mc_out[78]), .A4(n109), .Y(out[78])
         );
  AO22X1_HVT U27 ( .A1(n86), .A2(n97), .A3(mc_out[77]), .A4(n109), .Y(out[77])
         );
  AO22X1_HVT U28 ( .A1(oout[76]), .A2(n97), .A3(mc_out[76]), .A4(n109), .Y(
        out[76]) );
  AO22X1_HVT U29 ( .A1(n18), .A2(n97), .A3(mc_out[75]), .A4(n109), .Y(out[75])
         );
  AO22X1_HVT U30 ( .A1(n5), .A2(n97), .A3(mc_out[74]), .A4(n109), .Y(out[74])
         );
  AO22X1_HVT U31 ( .A1(n97), .A2(oout[73]), .A3(mc_out[73]), .A4(n109), .Y(
        out[73]) );
  AO22X1_HVT U32 ( .A1(n41), .A2(n97), .A3(mc_out[72]), .A4(n109), .Y(out[72])
         );
  AO22X1_HVT U33 ( .A1(n44), .A2(n97), .A3(mc_out[71]), .A4(n109), .Y(out[71])
         );
  AO22X1_HVT U34 ( .A1(oout[70]), .A2(n97), .A3(mc_out[70]), .A4(n109), .Y(
        out[70]) );
  AO22X1_HVT U35 ( .A1(n97), .A2(n1), .A3(mc_out[6]), .A4(n109), .Y(out[6]) );
  AO22X1_HVT U36 ( .A1(oout[69]), .A2(n98), .A3(mc_out[69]), .A4(n109), .Y(
        out[69]) );
  AO22X1_HVT U37 ( .A1(oout[68]), .A2(n98), .A3(mc_out[68]), .A4(n109), .Y(
        out[68]) );
  AO22X1_HVT U38 ( .A1(n11), .A2(n98), .A3(mc_out[67]), .A4(n110), .Y(out[67])
         );
  AO22X1_HVT U39 ( .A1(n62), .A2(n98), .A3(mc_out[66]), .A4(n110), .Y(out[66])
         );
  AO22X1_HVT U40 ( .A1(n61), .A2(n98), .A3(mc_out[65]), .A4(n110), .Y(out[65])
         );
  AO22X1_HVT U41 ( .A1(n39), .A2(n98), .A3(n110), .A4(mc_out[64]), .Y(out[64])
         );
  AO22X1_HVT U42 ( .A1(n71), .A2(n98), .A3(mc_out[63]), .A4(n110), .Y(out[63])
         );
  AO22X1_HVT U43 ( .A1(n93), .A2(n98), .A3(mc_out[62]), .A4(n110), .Y(out[62])
         );
  AO22X1_HVT U44 ( .A1(n21), .A2(n98), .A3(mc_out[61]), .A4(n110), .Y(out[61])
         );
  AO22X1_HVT U45 ( .A1(oout[60]), .A2(n98), .A3(mc_out[60]), .A4(n110), .Y(
        out[60]) );
  AO22X1_HVT U46 ( .A1(oout[5]), .A2(n98), .A3(mc_out[5]), .A4(n110), .Y(
        out[5]) );
  AO22X1_HVT U47 ( .A1(n72), .A2(n98), .A3(mc_out[59]), .A4(n110), .Y(out[59])
         );
  AO22X1_HVT U48 ( .A1(oout[58]), .A2(n98), .A3(mc_out[58]), .A4(n110), .Y(
        out[58]) );
  AO22X1_HVT U49 ( .A1(n87), .A2(n98), .A3(mc_out[57]), .A4(n110), .Y(out[57])
         );
  AO22X1_HVT U50 ( .A1(oout[56]), .A2(n98), .A3(mc_out[56]), .A4(n111), .Y(
        out[56]) );
  AO22X1_HVT U51 ( .A1(n90), .A2(n99), .A3(n111), .A4(mc_out[55]), .Y(out[55])
         );
  AO22X1_HVT U52 ( .A1(n99), .A2(n17), .A3(mc_out[54]), .A4(n111), .Y(out[54])
         );
  AO22X1_HVT U53 ( .A1(n63), .A2(n99), .A3(mc_out[53]), .A4(n111), .Y(out[53])
         );
  AO22X1_HVT U54 ( .A1(oout[52]), .A2(n99), .A3(mc_out[52]), .A4(n111), .Y(
        out[52]) );
  AO22X1_HVT U55 ( .A1(n57), .A2(n99), .A3(mc_out[51]), .A4(n111), .Y(out[51])
         );
  AO22X1_HVT U56 ( .A1(n99), .A2(n49), .A3(mc_out[50]), .A4(n111), .Y(out[50])
         );
  AO22X1_HVT U57 ( .A1(n14), .A2(n99), .A3(mc_out[4]), .A4(n111), .Y(out[4])
         );
  AO22X1_HVT U58 ( .A1(n15), .A2(n99), .A3(mc_out[49]), .A4(n111), .Y(out[49])
         );
  AO22X1_HVT U59 ( .A1(n66), .A2(n99), .A3(mc_out[48]), .A4(n111), .Y(out[48])
         );
  AO22X1_HVT U60 ( .A1(n89), .A2(n99), .A3(mc_out[47]), .A4(n111), .Y(out[47])
         );
  AO22X1_HVT U61 ( .A1(oout[46]), .A2(n99), .A3(mc_out[46]), .A4(n111), .Y(
        out[46]) );
  AO22X1_HVT U62 ( .A1(n74), .A2(n99), .A3(mc_out[45]), .A4(n112), .Y(out[45])
         );
  AO22X1_HVT U63 ( .A1(oout[44]), .A2(n99), .A3(mc_out[44]), .A4(n112), .Y(
        out[44]) );
  AO22X1_HVT U64 ( .A1(oout[43]), .A2(n99), .A3(mc_out[43]), .A4(n112), .Y(
        out[43]) );
  AO22X1_HVT U65 ( .A1(n34), .A2(n99), .A3(mc_out[42]), .A4(n112), .Y(out[42])
         );
  AO22X1_HVT U66 ( .A1(oout[41]), .A2(n100), .A3(mc_out[41]), .A4(n112), .Y(
        out[41]) );
  AO22X1_HVT U67 ( .A1(n36), .A2(n100), .A3(mc_out[40]), .A4(n112), .Y(out[40]) );
  AO22X1_HVT U68 ( .A1(oout[3]), .A2(n100), .A3(mc_out[3]), .A4(n112), .Y(
        out[3]) );
  AO22X1_HVT U69 ( .A1(n83), .A2(n100), .A3(mc_out[39]), .A4(n112), .Y(out[39]) );
  AO22X1_HVT U70 ( .A1(n37), .A2(n100), .A3(mc_out[38]), .A4(n112), .Y(out[38]) );
  AO22X1_HVT U71 ( .A1(n77), .A2(n100), .A3(mc_out[37]), .A4(n112), .Y(out[37]) );
  AO22X1_HVT U72 ( .A1(oout[36]), .A2(n100), .A3(mc_out[36]), .A4(n112), .Y(
        out[36]) );
  AO22X1_HVT U73 ( .A1(oout[35]), .A2(n100), .A3(mc_out[35]), .A4(n112), .Y(
        out[35]) );
  AO22X1_HVT U74 ( .A1(n65), .A2(n100), .A3(mc_out[34]), .A4(n113), .Y(out[34]) );
  AO22X1_HVT U75 ( .A1(n100), .A2(n29), .A3(mc_out[33]), .A4(n113), .Y(out[33]) );
  AO22X1_HVT U76 ( .A1(oout[32]), .A2(n100), .A3(mc_out[32]), .A4(n113), .Y(
        out[32]) );
  AO22X1_HVT U77 ( .A1(oout[31]), .A2(n100), .A3(mc_out[31]), .A4(n113), .Y(
        out[31]) );
  AO22X1_HVT U78 ( .A1(n59), .A2(n100), .A3(mc_out[30]), .A4(n113), .Y(out[30]) );
  AO22X1_HVT U79 ( .A1(n12), .A2(n100), .A3(mc_out[2]), .A4(n113), .Y(out[2])
         );
  AO22X1_HVT U80 ( .A1(n16), .A2(n100), .A3(mc_out[29]), .A4(n113), .Y(out[29]) );
  AO22X1_HVT U81 ( .A1(oout[28]), .A2(n101), .A3(mc_out[28]), .A4(n113), .Y(
        out[28]) );
  AO22X1_HVT U82 ( .A1(n19), .A2(n101), .A3(mc_out[27]), .A4(n113), .Y(out[27]) );
  AO22X1_HVT U83 ( .A1(n56), .A2(n101), .A3(mc_out[26]), .A4(n113), .Y(out[26]) );
  AO22X1_HVT U84 ( .A1(n101), .A2(n4), .A3(mc_out[25]), .A4(n113), .Y(out[25])
         );
  AO22X1_HVT U85 ( .A1(n3), .A2(n101), .A3(n113), .A4(mc_out[24]), .Y(out[24])
         );
  AO22X1_HVT U86 ( .A1(n80), .A2(n101), .A3(mc_out[23]), .A4(n114), .Y(out[23]) );
  AO22X1_HVT U87 ( .A1(n101), .A2(n25), .A3(mc_out[22]), .A4(n114), .Y(out[22]) );
  AO22X1_HVT U88 ( .A1(n58), .A2(n101), .A3(mc_out[21]), .A4(n114), .Y(out[21]) );
  AO22X1_HVT U89 ( .A1(oout[20]), .A2(n101), .A3(mc_out[20]), .A4(n114), .Y(
        out[20]) );
  AO22X1_HVT U90 ( .A1(n101), .A2(n45), .A3(mc_out[1]), .A4(n114), .Y(out[1])
         );
  AO22X1_HVT U91 ( .A1(n13), .A2(n101), .A3(mc_out[19]), .A4(n114), .Y(out[19]) );
  AO22X1_HVT U92 ( .A1(n35), .A2(n101), .A3(mc_out[18]), .A4(n114), .Y(out[18]) );
  AO22X1_HVT U93 ( .A1(n55), .A2(n101), .A3(n114), .A4(mc_out[17]), .Y(out[17]) );
  AO22X1_HVT U94 ( .A1(oout[16]), .A2(n101), .A3(mc_out[16]), .A4(n114), .Y(
        out[16]) );
  AO22X1_HVT U95 ( .A1(n92), .A2(n101), .A3(mc_out[15]), .A4(n114), .Y(out[15]) );
  AO22X1_HVT U96 ( .A1(n69), .A2(n102), .A3(mc_out[14]), .A4(n114), .Y(out[14]) );
  AO22X1_HVT U97 ( .A1(n102), .A2(n70), .A3(mc_out[13]), .A4(n114), .Y(out[13]) );
  AO22X1_HVT U98 ( .A1(oout[12]), .A2(n102), .A3(mc_out[12]), .A4(n115), .Y(
        out[12]) );
  AO22X1_HVT U99 ( .A1(n54), .A2(n102), .A3(mc_out[127]), .A4(n115), .Y(
        out[127]) );
  AO22X1_HVT U100 ( .A1(n102), .A2(n60), .A3(mc_out[126]), .A4(n115), .Y(
        out[126]) );
  AO22X1_HVT U101 ( .A1(n51), .A2(n102), .A3(mc_out[125]), .A4(n115), .Y(
        out[125]) );
  AO22X1_HVT U102 ( .A1(oout[124]), .A2(n102), .A3(mc_out[124]), .A4(n115), 
        .Y(out[124]) );
  AO22X1_HVT U103 ( .A1(n53), .A2(n102), .A3(mc_out[123]), .A4(n115), .Y(
        out[123]) );
  AO22X1_HVT U104 ( .A1(n48), .A2(n102), .A3(mc_out[122]), .A4(n115), .Y(
        out[122]) );
  AO22X1_HVT U105 ( .A1(n7), .A2(n102), .A3(mc_out[121]), .A4(n115), .Y(
        out[121]) );
  AO22X1_HVT U106 ( .A1(n6), .A2(n102), .A3(mc_out[120]), .A4(n115), .Y(
        out[120]) );
  AO22X1_HVT U107 ( .A1(oout[11]), .A2(n102), .A3(mc_out[11]), .A4(n115), .Y(
        out[11]) );
  AO22X1_HVT U108 ( .A1(n27), .A2(n102), .A3(mc_out[119]), .A4(n115), .Y(
        out[119]) );
  AO22X1_HVT U109 ( .A1(n73), .A2(n102), .A3(mc_out[118]), .A4(n115), .Y(
        out[118]) );
  AO22X1_HVT U110 ( .A1(n38), .A2(n102), .A3(mc_out[117]), .A4(n116), .Y(
        out[117]) );
  AO22X1_HVT U111 ( .A1(n103), .A2(oout[116]), .A3(mc_out[116]), .A4(n116), 
        .Y(out[116]) );
  AO22X1_HVT U112 ( .A1(oout[115]), .A2(n103), .A3(mc_out[115]), .A4(n116), 
        .Y(out[115]) );
  AO22X1_HVT U113 ( .A1(n76), .A2(n103), .A3(mc_out[114]), .A4(n116), .Y(
        out[114]) );
  AO22X1_HVT U114 ( .A1(oout[113]), .A2(n103), .A3(mc_out[113]), .A4(n116), 
        .Y(out[113]) );
  AO22X1_HVT U115 ( .A1(n103), .A2(oout[112]), .A3(mc_out[112]), .A4(n116), 
        .Y(out[112]) );
  AO22X1_HVT U116 ( .A1(n75), .A2(n103), .A3(mc_out[111]), .A4(n116), .Y(
        out[111]) );
  AO22X1_HVT U117 ( .A1(n8), .A2(n103), .A3(mc_out[110]), .A4(n116), .Y(
        out[110]) );
  AO22X1_HVT U118 ( .A1(n20), .A2(n103), .A3(mc_out[10]), .A4(n116), .Y(
        out[10]) );
  AO22X1_HVT U119 ( .A1(n23), .A2(n103), .A3(mc_out[109]), .A4(n116), .Y(
        out[109]) );
  AO22X1_HVT U120 ( .A1(oout[108]), .A2(n103), .A3(mc_out[108]), .A4(n116), 
        .Y(out[108]) );
  AO22X1_HVT U121 ( .A1(oout[107]), .A2(n103), .A3(mc_out[107]), .A4(n116), 
        .Y(out[107]) );
  AO22X1_HVT U122 ( .A1(n47), .A2(n103), .A3(mc_out[106]), .A4(n117), .Y(
        out[106]) );
  AO22X1_HVT U123 ( .A1(n79), .A2(n103), .A3(mc_out[105]), .A4(n117), .Y(
        out[105]) );
  AO22X1_HVT U124 ( .A1(n52), .A2(n103), .A3(mc_out[104]), .A4(n117), .Y(
        out[104]) );
  AO22X1_HVT U125 ( .A1(n26), .A2(n103), .A3(mc_out[103]), .A4(n117), .Y(
        out[103]) );
  AO22X1_HVT U126 ( .A1(n91), .A2(n104), .A3(mc_out[102]), .A4(n117), .Y(
        out[102]) );
  AO22X1_HVT U127 ( .A1(oout[101]), .A2(n104), .A3(mc_out[101]), .A4(n117), 
        .Y(out[101]) );
  AO22X1_HVT U128 ( .A1(oout[100]), .A2(n104), .A3(mc_out[100]), .A4(n117), 
        .Y(out[100]) );
  AO22X1_HVT U129 ( .A1(oout[0]), .A2(n104), .A3(mc_out[0]), .A4(n117), .Y(
        out[0]) );
  inv_shift_rows sr ( .in({in[127:56], n82, in[54:0]}), .out(sr_out) );
  inv_subbytes sb ( .in({sr_out[127:48], n85, sr_out[46:0]}), .out(sb_out) );
  inv_add_round_keys adk ( .state(sb_out), .subkey(keyin), .out(oout) );
  inv_Mix_Column mc ( .in(oout), .out1(mc_out) );
  DELLN2X2_HVT U1 ( .A(oout[75]), .Y(n18) );
  DELLN1X2_HVT U130 ( .A(oout[40]), .Y(n36) );
  DELLN2X2_HVT U131 ( .A(oout[6]), .Y(n1) );
  DELLN2X2_HVT U132 ( .A(oout[104]), .Y(n52) );
  DELLN2X2_HVT U133 ( .A(oout[94]), .Y(n2) );
  DELLN2X2_HVT U134 ( .A(oout[24]), .Y(n3) );
  DELLN2X2_HVT U135 ( .A(oout[25]), .Y(n4) );
  DELLN2X2_HVT U136 ( .A(oout[74]), .Y(n5) );
  DELLN2X2_HVT U137 ( .A(oout[120]), .Y(n6) );
  DELLN2X2_HVT U138 ( .A(oout[121]), .Y(n7) );
  DELLN1X2_HVT U139 ( .A(oout[42]), .Y(n34) );
  DELLN2X2_HVT U140 ( .A(oout[110]), .Y(n8) );
  DELLN2X2_HVT U141 ( .A(oout[78]), .Y(n9) );
  DELLN2X2_HVT U142 ( .A(oout[62]), .Y(n93) );
  DELLN1X2_HVT U143 ( .A(oout[45]), .Y(n74) );
  DELLN2X2_HVT U144 ( .A(oout[8]), .Y(n10) );
  DELLN2X2_HVT U145 ( .A(oout[67]), .Y(n11) );
  DELLN2X2_HVT U146 ( .A(oout[38]), .Y(n37) );
  DELLN2X2_HVT U147 ( .A(oout[2]), .Y(n12) );
  NBUFFX2_HVT U148 ( .A(oout[53]), .Y(n63) );
  DELLN2X2_HVT U149 ( .A(oout[19]), .Y(n13) );
  DELLN2X2_HVT U150 ( .A(oout[4]), .Y(n14) );
  DELLN2X2_HVT U151 ( .A(oout[49]), .Y(n15) );
  DELLN2X2_HVT U152 ( .A(oout[54]), .Y(n17) );
  DELLN2X2_HVT U153 ( .A(oout[29]), .Y(n16) );
  DELLN2X2_HVT U154 ( .A(oout[27]), .Y(n19) );
  INVX2_HVT U155 ( .A(n84), .Y(n85) );
  DELLN2X2_HVT U156 ( .A(oout[10]), .Y(n20) );
  DELLN2X2_HVT U157 ( .A(oout[61]), .Y(n21) );
  DELLN2X2_HVT U158 ( .A(oout[89]), .Y(n22) );
  DELLN1X2_HVT U159 ( .A(oout[97]), .Y(n24) );
  DELLN2X2_HVT U160 ( .A(oout[109]), .Y(n23) );
  DELLN2X2_HVT U161 ( .A(oout[22]), .Y(n25) );
  DELLN2X2_HVT U162 ( .A(oout[80]), .Y(n46) );
  DELLN2X2_HVT U163 ( .A(oout[103]), .Y(n26) );
  DELLN2X2_HVT U164 ( .A(oout[119]), .Y(n27) );
  DELLN2X2_HVT U165 ( .A(oout[90]), .Y(n28) );
  DELLN2X2_HVT U166 ( .A(oout[33]), .Y(n29) );
  DELLN2X2_HVT U167 ( .A(oout[48]), .Y(n66) );
  DELLN2X2_HVT U168 ( .A(oout[96]), .Y(n30) );
  DELLN2X2_HVT U169 ( .A(oout[88]), .Y(n31) );
  DELLN2X2_HVT U170 ( .A(oout[95]), .Y(n32) );
  DELLN2X2_HVT U171 ( .A(oout[91]), .Y(n33) );
  DELLN2X2_HVT U172 ( .A(oout[18]), .Y(n35) );
  DELLN2X2_HVT U173 ( .A(oout[117]), .Y(n38) );
  DELLN2X2_HVT U174 ( .A(oout[64]), .Y(n39) );
  DELLN2X2_HVT U175 ( .A(oout[93]), .Y(n40) );
  DELLN2X2_HVT U176 ( .A(oout[72]), .Y(n41) );
  DELLN2X2_HVT U177 ( .A(oout[82]), .Y(n42) );
  DELLN2X2_HVT U178 ( .A(oout[79]), .Y(n43) );
  DELLN2X2_HVT U179 ( .A(oout[71]), .Y(n44) );
  DELLN2X2_HVT U180 ( .A(oout[1]), .Y(n45) );
  DELLN2X2_HVT U181 ( .A(oout[106]), .Y(n47) );
  DELLN2X2_HVT U182 ( .A(oout[122]), .Y(n48) );
  DELLN2X2_HVT U183 ( .A(oout[50]), .Y(n49) );
  DELLN2X2_HVT U184 ( .A(oout[85]), .Y(n50) );
  DELLN2X2_HVT U185 ( .A(oout[125]), .Y(n51) );
  DELLN2X2_HVT U186 ( .A(oout[123]), .Y(n53) );
  DELLN2X2_HVT U187 ( .A(oout[127]), .Y(n54) );
  DELLN2X2_HVT U188 ( .A(oout[99]), .Y(n67) );
  DELLN2X2_HVT U189 ( .A(oout[17]), .Y(n55) );
  DELLN2X2_HVT U190 ( .A(oout[26]), .Y(n56) );
  NBUFFX2_HVT U191 ( .A(oout[51]), .Y(n57) );
  DELLN2X2_HVT U192 ( .A(oout[37]), .Y(n77) );
  DELLN2X2_HVT U193 ( .A(oout[21]), .Y(n58) );
  DELLN2X2_HVT U194 ( .A(oout[30]), .Y(n59) );
  DELLN2X2_HVT U195 ( .A(oout[126]), .Y(n60) );
  DELLN2X2_HVT U196 ( .A(oout[65]), .Y(n61) );
  DELLN2X2_HVT U197 ( .A(oout[66]), .Y(n62) );
  DELLN2X2_HVT U198 ( .A(oout[98]), .Y(n64) );
  DELLN2X2_HVT U199 ( .A(oout[34]), .Y(n65) );
  DELLN2X2_HVT U200 ( .A(oout[9]), .Y(n68) );
  DELLN2X2_HVT U201 ( .A(oout[14]), .Y(n69) );
  INVX1_HVT U202 ( .A(n81), .Y(n82) );
  DELLN2X2_HVT U203 ( .A(oout[13]), .Y(n70) );
  DELLN2X2_HVT U204 ( .A(oout[63]), .Y(n71) );
  DELLN2X2_HVT U205 ( .A(oout[59]), .Y(n72) );
  DELLN2X2_HVT U206 ( .A(oout[55]), .Y(n90) );
  DELLN2X2_HVT U207 ( .A(oout[118]), .Y(n73) );
  DELLN2X2_HVT U208 ( .A(oout[111]), .Y(n75) );
  DELLN2X2_HVT U209 ( .A(oout[23]), .Y(n80) );
  DELLN2X2_HVT U210 ( .A(oout[114]), .Y(n76) );
  DELLN2X2_HVT U211 ( .A(oout[81]), .Y(n78) );
  DELLN2X2_HVT U212 ( .A(oout[105]), .Y(n79) );
  INVX0_HVT U213 ( .A(in[55]), .Y(n81) );
  DELLN2X2_HVT U214 ( .A(oout[39]), .Y(n83) );
  INVX0_HVT U215 ( .A(sr_out[47]), .Y(n84) );
  DELLN2X2_HVT U216 ( .A(oout[77]), .Y(n86) );
  DELLN2X2_HVT U217 ( .A(oout[57]), .Y(n87) );
  DELLN2X2_HVT U218 ( .A(oout[87]), .Y(n88) );
  DELLN2X2_HVT U219 ( .A(oout[47]), .Y(n89) );
  DELLN2X2_HVT U220 ( .A(oout[102]), .Y(n91) );
  DELLN2X2_HVT U221 ( .A(oout[15]), .Y(n92) );
  INVX0_HVT U222 ( .A(last), .Y(n105) );
  INVX1_HVT U223 ( .A(n95), .Y(n107) );
  INVX1_HVT U224 ( .A(n95), .Y(n108) );
  INVX1_HVT U225 ( .A(n95), .Y(n111) );
  INVX1_HVT U226 ( .A(n95), .Y(n110) );
  INVX1_HVT U227 ( .A(n95), .Y(n109) );
  INVX1_HVT U228 ( .A(n94), .Y(n113) );
  INVX1_HVT U229 ( .A(n94), .Y(n114) );
  INVX1_HVT U230 ( .A(n94), .Y(n115) );
  INVX1_HVT U231 ( .A(n94), .Y(n116) );
  INVX1_HVT U232 ( .A(n94), .Y(n112) );
  INVX1_HVT U233 ( .A(n94), .Y(n117) );
  INVX1_HVT U234 ( .A(n106), .Y(n96) );
  INVX1_HVT U235 ( .A(n106), .Y(n97) );
  INVX1_HVT U236 ( .A(n105), .Y(n99) );
  INVX1_HVT U237 ( .A(n105), .Y(n101) );
  INVX1_HVT U238 ( .A(n105), .Y(n102) );
  INVX1_HVT U239 ( .A(n105), .Y(n100) );
  INVX1_HVT U240 ( .A(n105), .Y(n103) );
  INVX1_HVT U241 ( .A(n106), .Y(n98) );
  INVX1_HVT U242 ( .A(n106), .Y(n95) );
  INVX1_HVT U243 ( .A(n106), .Y(n94) );
  INVX1_HVT U244 ( .A(n105), .Y(n104) );
  INVX0_HVT U245 ( .A(last), .Y(n106) );
endmodule

