
module keygen_1 ( round_num, keyin, keyout );
  input [0:3] round_num;
  input [0:127] keyin;
  output [0:127] keyout;
  wire   n23, n49, n211, n212, n213, n214, n217, n218, n219, n220, n232, n233,
         n234, n235, n236, n237, n238, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n328, n354, n398, n472, n473, n474,
         n516, n517, n518, n519, n522, n523, n524, n525, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n633, n740, n768, n821, n822, n823, n824,
         n827, n828, n829, n830, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n861, n862, n863, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n938, n963, n965,
         n1083, n1125, n1126, n1127, n1130, n1131, n1132, n1133, n1134, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1169,
         n1170, n1171, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1485, n1486, n1487, n1488, n1489, n1490, n1492, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715;
  wire   [0:31] dummy;

  NAND2X0_HVT U4 ( .A1(n1453), .A2(n1417), .Y(n2712) );
  NAND2X0_HVT U5 ( .A1(n1381), .A2(n217), .Y(n2711) );
  NAND2X0_HVT U6 ( .A1(n1415), .A2(n2712), .Y(n2710) );
  NAND2X0_HVT U15 ( .A1(n2700), .A2(n1421), .Y(n2701) );
  NAND2X0_HVT U17 ( .A1(n2712), .A2(n1684), .Y(n2698) );
  NAND2X0_HVT U21 ( .A1(n1414), .A2(n1458), .Y(n2694) );
  NAND2X0_HVT U25 ( .A1(n1380), .A2(n1458), .Y(n2691) );
  NAND2X0_HVT U33 ( .A1(n1458), .A2(n1689), .Y(n2683) );
  NAND2X0_HVT U34 ( .A1(n1685), .A2(n1458), .Y(n2682) );
  NAND2X0_HVT U39 ( .A1(n214), .A2(n1358), .Y(n2677) );
  MUX41X1_HVT U50 ( .A1(n1671), .A3(n1628), .A2(n2702), .A4(n1648), .S0(n555), 
        .S1(n1246), .Y(n2667) );
  NAND2X0_HVT U52 ( .A1(n2664), .A2(n2674), .Y(n2665) );
  MUX41X1_HVT U55 ( .A1(n1196), .A3(n1647), .A2(n1646), .A4(n1684), .S0(n542), 
        .S1(n1247), .Y(n2661) );
  NAND2X0_HVT U56 ( .A1(n1458), .A2(n1418), .Y(n2660) );
  MUX41X1_HVT U57 ( .A1(n2660), .A3(n1636), .A2(n1666), .A4(n1645), .S0(n542), 
        .S1(n1246), .Y(n2659) );
  NAND2X0_HVT U59 ( .A1(n1415), .A2(n2656), .Y(n2657) );
  MUX41X1_HVT U60 ( .A1(n1672), .A3(n1644), .A2(n2657), .A4(n2705), .S0(n556), 
        .S1(n1247), .Y(n2655) );
  NAND2X0_HVT U61 ( .A1(n1421), .A2(n2712), .Y(n2654) );
  MUX41X1_HVT U62 ( .A1(n1224), .A3(n2654), .A2(n1221), .A4(n1643), .S0(n542), 
        .S1(n1246), .Y(n2653) );
  AO21X1_HVT U65 ( .A1(n1641), .A2(n1252), .A3(n1665), .Y(n2650) );
  MUX41X1_HVT U67 ( .A1(n1639), .A3(n2650), .A2(n2649), .A4(n2651), .S0(n1460), 
        .S1(n1463), .Y(n2648) );
  MUX41X1_HVT U69 ( .A1(n2673), .A3(n1687), .A2(n2691), .A4(n1673), .S0(n1249), 
        .S1(n556), .Y(n2647) );
  NAND2X0_HVT U71 ( .A1(n1419), .A2(n2644), .Y(n2645) );
  MUX41X1_HVT U77 ( .A1(n2671), .A3(n1629), .A2(n2695), .A4(n1420), .S0(n1255), 
        .S1(n1246), .Y(n2637) );
  MUX41X1_HVT U80 ( .A1(n2635), .A3(n1674), .A2(n1675), .A4(n1650), .S0(n1250), 
        .S1(n542), .Y(n2634) );
  MUX41X1_HVT U81 ( .A1(n2706), .A3(n1667), .A2(n1676), .A4(n1688), .S0(n1250), 
        .S1(n1464), .Y(n2633) );
  AND2X1_HVT U82 ( .A1(n1452), .A2(n1384), .Y(n2632) );
  NAND2X0_HVT U83 ( .A1(n1458), .A2(n1687), .Y(n2631) );
  MUX41X1_HVT U84 ( .A1(n2631), .A3(n244), .A2(n1198), .A4(n2632), .S0(n1250), 
        .S1(n542), .Y(n2630) );
  MUX41X1_HVT U85 ( .A1(n1674), .A3(n1649), .A2(n1211), .A4(n2697), .S0(n1249), 
        .S1(n555), .Y(n2629) );
  MUX41X1_HVT U86 ( .A1(n2629), .A3(n2633), .A2(n2630), .A4(n2634), .S0(
        keyin[105]), .S1(n902), .Y(n2628) );
  NAND2X0_HVT U97 ( .A1(n2616), .A2(n2615), .Y(n2617) );
  MUX41X1_HVT U102 ( .A1(n1667), .A3(n1629), .A2(n214), .A4(n1673), .S0(n1249), 
        .S1(n1464), .Y(n2610) );
  MUX41X1_HVT U104 ( .A1(n2669), .A3(n1669), .A2(n1640), .A4(n2683), .S0(n268), 
        .S1(n1248), .Y(n2608) );
  MUX41X1_HVT U106 ( .A1(n1651), .A3(n2712), .A2(n2607), .A4(n1652), .S0(n1250), .S1(n542), .Y(n2606) );
  NAND2X0_HVT U111 ( .A1(n1417), .A2(n2601), .Y(n2602) );
  MUX41X1_HVT U115 ( .A1(n2598), .A3(n2604), .A2(n2600), .A4(n2603), .S0(n1250), .S1(n252), .Y(n2597) );
  NAND2X0_HVT U118 ( .A1(n2593), .A2(n2592), .Y(n2594) );
  MUX41X1_HVT U120 ( .A1(n2694), .A3(n1224), .A2(n1639), .A4(n1678), .S0(n902), 
        .S1(n1464), .Y(n2590) );
  AND2X1_HVT U122 ( .A1(n1453), .A2(n243), .Y(n2588) );
  AO21X1_HVT U125 ( .A1(n1459), .A2(n1419), .A3(n244), .Y(n2585) );
  AND3X1_HVT U129 ( .A1(n1460), .A2(n1458), .A3(n1383), .Y(n2581) );
  MUX41X1_HVT U132 ( .A1(n2579), .A3(n2581), .A2(n2580), .A4(n2582), .S0(n1249), .S1(n251), .Y(n2578) );
  MUX41X1_HVT U133 ( .A1(n2578), .A3(n2583), .A2(n2589), .A4(n2597), .S0(
        keyin[105]), .S1(n1377), .Y(dummy[4]) );
  MUX41X1_HVT U134 ( .A1(n1683), .A3(n2690), .A2(n1678), .A4(n1420), .S0(n556), 
        .S1(n1248), .Y(n2577) );
  MUX41X1_HVT U137 ( .A1(n1684), .A3(n1661), .A2(n1419), .A4(n1656), .S0(n1249), .S1(n542), .Y(n2574) );
  AND2X1_HVT U138 ( .A1(n1420), .A2(n1457), .Y(n2573) );
  MUX41X1_HVT U139 ( .A1(n1649), .A3(n1668), .A2(n2692), .A4(n2573), .S0(n556), 
        .S1(n1245), .Y(n2572) );
  MUX41X1_HVT U140 ( .A1(n2572), .A3(n2574), .A2(n2575), .A4(n2577), .S0(n902), 
        .S1(keyin[105]), .Y(n2571) );
  MUX41X1_HVT U143 ( .A1(n2693), .A3(n1198), .A2(n1660), .A4(n1680), .S0(n1250), .S1(n1464), .Y(n2568) );
  NAND2X0_HVT U144 ( .A1(n1455), .A2(n1421), .Y(n2644) );
  MUX41X1_HVT U148 ( .A1(n1680), .A3(n1667), .A2(n2688), .A4(n1635), .S0(n1464), .S1(n1248), .Y(n2564) );
  MUX41X1_HVT U151 ( .A1(n1196), .A3(n1630), .A2(n1675), .A4(n1683), .S0(n542), 
        .S1(n1248), .Y(n2562) );
  AND2X1_HVT U156 ( .A1(n244), .A2(n2644), .Y(n2556) );
  MUX41X1_HVT U158 ( .A1(n2670), .A3(n2556), .A2(n2555), .A4(n2557), .S0(n1253), .S1(n542), .Y(n2554) );
  MUX41X1_HVT U159 ( .A1(n2694), .A3(n1647), .A2(n1654), .A4(n1213), .S0(n1249), .S1(n542), .Y(n2553) );
  MUX41X1_HVT U160 ( .A1(n2553), .A3(n2554), .A2(n2558), .A4(n2562), .S0(n902), 
        .S1(keyin[105]), .Y(n2552) );
  AND2X1_HVT U161 ( .A1(n251), .A2(n1381), .Y(n2551) );
  NAND2X0_HVT U165 ( .A1(n1453), .A2(n1687), .Y(n2547) );
  MUX41X1_HVT U166 ( .A1(n2701), .A3(n2678), .A2(n2547), .A4(n1676), .S0(n1250), .S1(n1463), .Y(n2546) );
  NAND2X0_HVT U167 ( .A1(n1421), .A2(n2656), .Y(n2545) );
  NAND2X0_HVT U171 ( .A1(n1688), .A2(n1458), .Y(n2541) );
  MUX41X1_HVT U172 ( .A1(n1419), .A3(n1673), .A2(n1672), .A4(n2541), .S0(n555), 
        .S1(n1248), .Y(n2540) );
  NAND2X0_HVT U175 ( .A1(n1452), .A2(n2708), .Y(n2700) );
  NAND2X0_HVT U176 ( .A1(n1454), .A2(n1689), .Y(n2538) );
  MUX41X1_HVT U177 ( .A1(n2538), .A3(n2678), .A2(n1677), .A4(n2700), .S0(n556), 
        .S1(n1245), .Y(n2537) );
  MUX41X1_HVT U179 ( .A1(n2696), .A3(n1689), .A2(n1681), .A4(n2536), .S0(n1251), .S1(n1464), .Y(n2535) );
  MUX41X1_HVT U180 ( .A1(n2631), .A3(n1379), .A2(n1664), .A4(n1632), .S0(n555), 
        .S1(n1245), .Y(n2534) );
  MUX41X1_HVT U184 ( .A1(n2531), .A3(n2535), .A2(n2534), .A4(n2537), .S0(
        keyin[105]), .S1(n1460), .Y(n2530) );
  MUX41X1_HVT U185 ( .A1(n2701), .A3(n1682), .A2(n1197), .A4(n1681), .S0(n1251), .S1(n1463), .Y(n2529) );
  MUX41X1_HVT U186 ( .A1(n1637), .A3(n2689), .A2(n2706), .A4(n1634), .S0(n1251), .S1(n1463), .Y(n2528) );
  MUX41X1_HVT U188 ( .A1(n2527), .A3(n2679), .A2(n1669), .A4(n2670), .S0(n1249), .S1(n270), .Y(n2526) );
  MUX41X1_HVT U190 ( .A1(n2525), .A3(n1204), .A2(n2700), .A4(n2644), .S0(n1251), .S1(n1464), .Y(n2524) );
  MUX41X1_HVT U191 ( .A1(n2524), .A3(n2528), .A2(n2526), .A4(n2529), .S0(
        keyin[105]), .S1(n901), .Y(n2523) );
  MUX41X1_HVT U194 ( .A1(n1679), .A3(n2683), .A2(n1420), .A4(n2522), .S0(n1251), .S1(n1463), .Y(n2521) );
  MUX41X1_HVT U195 ( .A1(n2675), .A3(n2711), .A2(n2690), .A4(n2668), .S0(n1251), .S1(n251), .Y(n2520) );
  MUX41X1_HVT U196 ( .A1(n1663), .A3(n2685), .A2(n2697), .A4(n1197), .S0(n1463), .S1(n1247), .Y(n2519) );
  MUX41X1_HVT U200 ( .A1(n2516), .A3(n2520), .A2(n2519), .A4(n2521), .S0(
        keyin[105]), .S1(n902), .Y(n2515) );
  AO21X1_HVT U202 ( .A1(n1211), .A2(n1255), .A3(n1670), .Y(n2513) );
  MUX41X1_HVT U204 ( .A1(n1638), .A3(n244), .A2(n1681), .A4(n2715), .S0(n1251), 
        .S1(n252), .Y(n2511) );
  MUX41X1_HVT U205 ( .A1(n2712), .A3(n2701), .A2(n1653), .A4(n2693), .S0(n1251), .S1(n1463), .Y(n2510) );
  MUX41X1_HVT U206 ( .A1(n1383), .A3(n2657), .A2(n1682), .A4(n1657), .S0(n1251), .S1(n1464), .Y(n2509) );
  NAND2X0_HVT U211 ( .A1(n1420), .A2(n1455), .Y(n2656) );
  NAND2X0_HVT U212 ( .A1(n1452), .A2(n1414), .Y(n2601) );
  NAND2X0_HVT U215 ( .A1(n244), .A2(n1458), .Y(n2507) );
  NAND2X0_HVT U216 ( .A1(n1419), .A2(n2601), .Y(n2506) );
  NAND2X0_HVT U219 ( .A1(n1455), .A2(n1683), .Y(n2559) );
  NAND2X0_HVT U221 ( .A1(n252), .A2(n2507), .Y(n2639) );
  NAND2X0_HVT U317 ( .A1(n1439), .A2(n1409), .Y(n2491) );
  NAND2X0_HVT U318 ( .A1(n1372), .A2(n1440), .Y(n2490) );
  NAND2X0_HVT U319 ( .A1(n1407), .A2(n2491), .Y(n2489) );
  XOR2X2_HVT U320 ( .A1(n1622), .A2(n1373), .Y(n2487) );
  NAND2X0_HVT U328 ( .A1(n2479), .A2(n1413), .Y(n2480) );
  NAND2X0_HVT U330 ( .A1(n2491), .A2(n1355), .Y(n2477) );
  NAND2X0_HVT U334 ( .A1(n1406), .A2(n1442), .Y(n2473) );
  NAND2X0_HVT U338 ( .A1(n1371), .A2(n1442), .Y(n2470) );
  NAND2X0_HVT U346 ( .A1(n1442), .A2(n1625), .Y(n2462) );
  NAND2X0_HVT U347 ( .A1(n1621), .A2(n1442), .Y(n2461) );
  NAND2X0_HVT U352 ( .A1(n1438), .A2(n599), .Y(n2456) );
  MUX41X1_HVT U363 ( .A1(n1607), .A3(n1565), .A2(n2481), .A4(n1585), .S0(n873), 
        .S1(n1236), .Y(n2446) );
  NAND2X0_HVT U365 ( .A1(n2443), .A2(n2453), .Y(n2444) );
  MUX41X1_HVT U368 ( .A1(n1192), .A3(n1584), .A2(n1583), .A4(n1354), .S0(n873), 
        .S1(n1446), .Y(n2440) );
  NAND2X0_HVT U369 ( .A1(n1442), .A2(n1410), .Y(n2439) );
  MUX41X1_HVT U370 ( .A1(n2439), .A3(n1573), .A2(n1602), .A4(n1582), .S0(n236), 
        .S1(n1236), .Y(n2438) );
  NAND2X0_HVT U372 ( .A1(n1407), .A2(n2435), .Y(n2436) );
  MUX41X1_HVT U373 ( .A1(n1608), .A3(n1581), .A2(n2436), .A4(n2484), .S0(n237), 
        .S1(n1235), .Y(n2434) );
  NAND2X0_HVT U374 ( .A1(n1413), .A2(n2491), .Y(n2433) );
  MUX41X1_HVT U375 ( .A1(n1222), .A3(n2433), .A2(n1218), .A4(n1580), .S0(n237), 
        .S1(n1236), .Y(n2432) );
  AO21X1_HVT U378 ( .A1(n1578), .A2(n1241), .A3(n1601), .Y(n2429) );
  MUX41X1_HVT U380 ( .A1(n1576), .A3(n2429), .A2(n2428), .A4(n2430), .S0(n1443), .S1(n236), .Y(n2427) );
  MUX41X1_HVT U381 ( .A1(n2427), .A3(n2431), .A2(n2437), .A4(n2441), .S0(n1376), .S1(n1369), .Y(dummy[15]) );
  MUX41X1_HVT U382 ( .A1(n2452), .A3(n1623), .A2(n2470), .A4(n1609), .S0(n1238), .S1(n1450), .Y(n2426) );
  NAND2X0_HVT U384 ( .A1(n1412), .A2(n2423), .Y(n2424) );
  AND3X1_HVT U388 ( .A1(n1410), .A2(n2435), .A3(n2418), .Y(n2419) );
  MUX41X1_HVT U390 ( .A1(n2450), .A3(n1566), .A2(n2474), .A4(n1411), .S0(n237), 
        .S1(n1236), .Y(n2416) );
  MUX41X1_HVT U391 ( .A1(n2416), .A3(n2417), .A2(n2421), .A4(n2426), .S0(n247), 
        .S1(n1376), .Y(n2415) );
  MUX41X1_HVT U393 ( .A1(n2414), .A3(n1610), .A2(n1611), .A4(n1587), .S0(n1239), .S1(n236), .Y(n2413) );
  MUX41X1_HVT U394 ( .A1(n2485), .A3(n1603), .A2(n1612), .A4(n1624), .S0(n1239), .S1(n236), .Y(n2412) );
  AND2X1_HVT U395 ( .A1(n1437), .A2(n1375), .Y(n2411) );
  NAND2X0_HVT U396 ( .A1(n1442), .A2(n1623), .Y(n2410) );
  MUX41X1_HVT U397 ( .A1(n2410), .A3(n2487), .A2(n1190), .A4(n2411), .S0(n1239), .S1(n237), .Y(n2409) );
  MUX41X1_HVT U398 ( .A1(n1610), .A3(n1586), .A2(n1207), .A4(n2476), .S0(n1238), .S1(n862), .Y(n2408) );
  MUX41X1_HVT U399 ( .A1(n2408), .A3(n2412), .A2(n2409), .A4(n2413), .S0(
        keyin[113]), .S1(n247), .Y(n2407) );
  AO21X1_HVT U406 ( .A1(n1243), .A2(n2401), .A3(n1606), .Y(n2402) );
  MUX41X1_HVT U407 ( .A1(n2402), .A3(n2404), .A2(n2403), .A4(n2405), .S0(n247), 
        .S1(n1235), .Y(n2400) );
  NAND2X0_HVT U410 ( .A1(n2396), .A2(n2395), .Y(n2397) );
  MUX41X1_HVT U415 ( .A1(n1603), .A3(n1566), .A2(n1437), .A4(n1609), .S0(n1238), .S1(n862), .Y(n2390) );
  MUX41X1_HVT U417 ( .A1(n2448), .A3(n1605), .A2(n1577), .A4(n2462), .S0(n873), 
        .S1(n1237), .Y(n2388) );
  MUX41X1_HVT U419 ( .A1(n1588), .A3(n2491), .A2(n2387), .A4(n1589), .S0(n1239), .S1(n862), .Y(n2386) );
  NAND2X0_HVT U424 ( .A1(n1409), .A2(n2381), .Y(n2382) );
  NAND2X0_HVT U431 ( .A1(n2373), .A2(n2372), .Y(n2374) );
  MUX41X1_HVT U433 ( .A1(n2473), .A3(n1222), .A2(n1576), .A4(n1614), .S0(n1443), .S1(n862), .Y(n2370) );
  AND2X1_HVT U435 ( .A1(n1440), .A2(n1354), .Y(n2368) );
  MUX41X1_HVT U436 ( .A1(n2480), .A3(n2368), .A2(n1587), .A4(n2466), .S0(n1443), .S1(n237), .Y(n2367) );
  AO21X1_HVT U438 ( .A1(n1444), .A2(n1412), .A3(n2487), .Y(n2365) );
  AND3X1_HVT U442 ( .A1(n247), .A2(n1442), .A3(n1374), .Y(n2361) );
  MUX41X1_HVT U445 ( .A1(n2359), .A3(n2361), .A2(n2360), .A4(n2362), .S0(n1238), .S1(n873), .Y(n2358) );
  MUX41X1_HVT U447 ( .A1(n1619), .A3(n2469), .A2(n1614), .A4(n1411), .S0(n236), 
        .S1(n1237), .Y(n2357) );
  MUX41X1_HVT U450 ( .A1(n1354), .A3(n1598), .A2(n1411), .A4(n1593), .S0(n1238), .S1(n237), .Y(n2354) );
  AND2X1_HVT U451 ( .A1(n2493), .A2(n1441), .Y(n2353) );
  MUX41X1_HVT U452 ( .A1(n1586), .A3(n1604), .A2(n2471), .A4(n2353), .S0(n873), 
        .S1(n1235), .Y(n2352) );
  MUX41X1_HVT U453 ( .A1(n2352), .A3(n2354), .A2(n2355), .A4(n2357), .S0(n247), 
        .S1(keyin[113]), .Y(n2351) );
  MUX41X1_HVT U456 ( .A1(n2472), .A3(n1190), .A2(n1597), .A4(n1616), .S0(n1239), .S1(n1450), .Y(n2348) );
  NAND2X0_HVT U457 ( .A1(n1439), .A2(n1413), .Y(n2423) );
  MUX41X1_HVT U461 ( .A1(n1616), .A3(n1603), .A2(n2467), .A4(n1572), .S0(n1243), .S1(n1237), .Y(n2344) );
  MUX41X1_HVT U464 ( .A1(n1192), .A3(n1567), .A2(n1611), .A4(n1619), .S0(n873), 
        .S1(n1237), .Y(n2342) );
  AND2X1_HVT U469 ( .A1(n2487), .A2(n2423), .Y(n2336) );
  MUX41X1_HVT U472 ( .A1(n2473), .A3(n1584), .A2(n1591), .A4(n1209), .S0(n1238), .S1(n862), .Y(n2333) );
  NAND2X0_HVT U478 ( .A1(n1437), .A2(n1623), .Y(n2330) );
  MUX41X1_HVT U479 ( .A1(n2480), .A3(n2457), .A2(n2330), .A4(n1612), .S0(n1239), .S1(n862), .Y(n2329) );
  NAND2X0_HVT U480 ( .A1(n1413), .A2(n2435), .Y(n2328) );
  NAND2X0_HVT U484 ( .A1(n1624), .A2(n1442), .Y(n2324) );
  MUX41X1_HVT U485 ( .A1(n1411), .A3(n1609), .A2(n1608), .A4(n2324), .S0(n873), 
        .S1(n1237), .Y(n2323) );
  NAND2X0_HVT U488 ( .A1(n1439), .A2(n2487), .Y(n2479) );
  NAND2X0_HVT U489 ( .A1(n1437), .A2(n1625), .Y(n2321) );
  MUX41X1_HVT U490 ( .A1(n2321), .A3(n2457), .A2(n1613), .A4(n2479), .S0(n1244), .S1(n1235), .Y(n2320) );
  MUX41X1_HVT U492 ( .A1(n2475), .A3(n1625), .A2(n1617), .A4(n2319), .S0(n1240), .S1(n862), .Y(n2318) );
  MUX41X1_HVT U493 ( .A1(n2410), .A3(n1372), .A2(n1600), .A4(n1569), .S0(n1244), .S1(n1235), .Y(n2317) );
  MUX41X1_HVT U497 ( .A1(n2314), .A3(n2318), .A2(n2317), .A4(n2320), .S0(
        keyin[113]), .S1(n247), .Y(n2313) );
  MUX41X1_HVT U498 ( .A1(n2480), .A3(n1618), .A2(n1194), .A4(n1617), .S0(n1240), .S1(n862), .Y(n2312) );
  MUX41X1_HVT U499 ( .A1(n1574), .A3(n2468), .A2(n2485), .A4(n1571), .S0(n1240), .S1(n862), .Y(n2311) );
  MUX41X1_HVT U501 ( .A1(n2310), .A3(n2458), .A2(n1605), .A4(n2449), .S0(n1238), .S1(n862), .Y(n2309) );
  MUX41X1_HVT U503 ( .A1(n2308), .A3(n1202), .A2(n2479), .A4(n2423), .S0(n1240), .S1(n237), .Y(n2307) );
  MUX41X1_HVT U504 ( .A1(n2307), .A3(n2311), .A2(n2309), .A4(n2312), .S0(n1376), .S1(n247), .Y(n2306) );
  MUX41X1_HVT U507 ( .A1(n1615), .A3(n2462), .A2(n1411), .A4(n2305), .S0(n1240), .S1(n1450), .Y(n2304) );
  MUX41X1_HVT U508 ( .A1(n2454), .A3(n2490), .A2(n2469), .A4(n2447), .S0(n1240), .S1(n236), .Y(n2303) );
  MUX41X1_HVT U509 ( .A1(n1599), .A3(n2464), .A2(n2476), .A4(n1194), .S0(n1450), .S1(n1446), .Y(n2302) );
  AO21X1_HVT U515 ( .A1(n1207), .A2(n873), .A3(n1606), .Y(n2296) );
  MUX41X1_HVT U519 ( .A1(n1374), .A3(n2436), .A2(n1618), .A4(n1594), .S0(n1240), .S1(n1450), .Y(n2292) );
  NAND2X0_HVT U524 ( .A1(n1412), .A2(n1439), .Y(n2435) );
  NAND2X0_HVT U525 ( .A1(n1439), .A2(n1406), .Y(n2381) );
  NAND2X0_HVT U528 ( .A1(n2487), .A2(n1442), .Y(n2290) );
  NAND2X0_HVT U529 ( .A1(n1412), .A2(n2381), .Y(n2289) );
  NAND2X0_HVT U532 ( .A1(n1440), .A2(n1619), .Y(n2339) );
  NAND2X0_HVT U534 ( .A1(n1244), .A2(n2290), .Y(n2418) );
  NAND2X0_HVT U631 ( .A1(n1366), .A2(n1425), .Y(n2273) );
  NAND2X0_HVT U632 ( .A1(n1398), .A2(n2274), .Y(n2272) );
  XOR2X2_HVT U633 ( .A1(n1555), .A2(n1367), .Y(n2270) );
  NAND2X0_HVT U641 ( .A1(n2262), .A2(n1405), .Y(n2263) );
  NAND2X0_HVT U643 ( .A1(n2274), .A2(n1352), .Y(n2260) );
  NAND2X0_HVT U647 ( .A1(n1397), .A2(n1428), .Y(n2256) );
  NAND2X0_HVT U651 ( .A1(n1365), .A2(n1428), .Y(n2253) );
  NAND2X0_HVT U659 ( .A1(n1428), .A2(n1557), .Y(n2245) );
  NAND2X0_HVT U660 ( .A1(n1554), .A2(n1428), .Y(n2244) );
  NAND2X0_HVT U665 ( .A1(n1426), .A2(n1353), .Y(n2239) );
  MUX41X1_HVT U676 ( .A1(n1540), .A3(n1497), .A2(n2264), .A4(n1517), .S0(n283), 
        .S1(n1226), .Y(n2229) );
  NAND2X0_HVT U678 ( .A1(n2226), .A2(n2236), .Y(n2227) );
  MUX41X1_HVT U681 ( .A1(n1193), .A3(n1516), .A2(n1515), .A4(n1351), .S0(n283), 
        .S1(n1226), .Y(n2223) );
  NAND2X0_HVT U682 ( .A1(n1428), .A2(n1401), .Y(n2222) );
  NAND2X0_HVT U685 ( .A1(n1398), .A2(n2218), .Y(n2219) );
  NAND2X0_HVT U687 ( .A1(n1405), .A2(n2274), .Y(n2216) );
  MUX41X1_HVT U688 ( .A1(n1223), .A3(n2216), .A2(n1219), .A4(n1512), .S0(n283), 
        .S1(n1226), .Y(n2215) );
  AO21X1_HVT U691 ( .A1(n1510), .A2(n1231), .A3(n1534), .Y(n2212) );
  NAND2X0_HVT U697 ( .A1(n1403), .A2(n2206), .Y(n2207) );
  AND3X1_HVT U701 ( .A1(n1401), .A2(n2218), .A3(n2201), .Y(n2202) );
  MUX41X1_HVT U706 ( .A1(n2197), .A3(n1543), .A2(n1544), .A4(n1519), .S0(n1229), .S1(n472), .Y(n2196) );
  MUX41X1_HVT U707 ( .A1(n2268), .A3(n1536), .A2(n1545), .A4(n1163), .S0(n1229), .S1(n472), .Y(n2195) );
  AND2X1_HVT U708 ( .A1(n1423), .A2(n1368), .Y(n2194) );
  NAND2X0_HVT U709 ( .A1(n1428), .A2(n1556), .Y(n2193) );
  MUX41X1_HVT U711 ( .A1(n1543), .A3(n1518), .A2(n1208), .A4(n2259), .S0(n1228), .S1(n238), .Y(n2191) );
  AO21X1_HVT U719 ( .A1(n1434), .A2(n2183), .A3(n1539), .Y(n2184) );
  NAND2X0_HVT U723 ( .A1(n2178), .A2(n2177), .Y(n2179) );
  MUX41X1_HVT U728 ( .A1(n1536), .A3(n1498), .A2(n1423), .A4(n1542), .S0(n1228), .S1(n238), .Y(n2172) );
  MUX41X1_HVT U730 ( .A1(n2231), .A3(n1538), .A2(n1509), .A4(n2245), .S0(n283), 
        .S1(n1227), .Y(n2170) );
  MUX41X1_HVT U732 ( .A1(n1520), .A3(n2274), .A2(n2169), .A4(n1521), .S0(n1229), .S1(n238), .Y(n2168) );
  OA21X1_HVT U736 ( .A1(n1528), .A2(n1430), .A3(n1512), .Y(n2165) );
  NAND2X0_HVT U737 ( .A1(n1400), .A2(n2163), .Y(n2164) );
  MUX41X1_HVT U741 ( .A1(n2160), .A3(n2166), .A2(n2162), .A4(n2165), .S0(n1229), .S1(n238), .Y(n2159) );
  NAND2X0_HVT U744 ( .A1(n2155), .A2(n2154), .Y(n2156) );
  MUX41X1_HVT U746 ( .A1(n2256), .A3(n1223), .A2(n1508), .A4(n1547), .S0(n572), 
        .S1(n238), .Y(n2152) );
  AO21X1_HVT U751 ( .A1(n1429), .A2(n1403), .A3(n2270), .Y(n2148) );
  AND3X1_HVT U755 ( .A1(n1429), .A2(n1428), .A3(n1368), .Y(n2144) );
  MUX41X1_HVT U758 ( .A1(n2142), .A3(n2144), .A2(n2143), .A4(n2145), .S0(n1228), .S1(n283), .Y(n2141) );
  MUX41X1_HVT U760 ( .A1(n1552), .A3(n2252), .A2(n1547), .A4(n1402), .S0(n283), 
        .S1(n1227), .Y(n2140) );
  AND2X1_HVT U764 ( .A1(n1404), .A2(n1427), .Y(n2136) );
  MUX41X1_HVT U765 ( .A1(n1518), .A3(n1537), .A2(n2254), .A4(n2136), .S0(n283), 
        .S1(n1431), .Y(n2135) );
  MUX41X1_HVT U769 ( .A1(n2255), .A3(n1191), .A2(n1529), .A4(n1549), .S0(n1229), .S1(n472), .Y(n2131) );
  NAND2X0_HVT U770 ( .A1(n1422), .A2(n1405), .Y(n2206) );
  MUX41X1_HVT U774 ( .A1(n1549), .A3(n1536), .A2(n2250), .A4(n1504), .S0(n283), 
        .S1(n1227), .Y(n2127) );
  MUX41X1_HVT U777 ( .A1(n1193), .A3(n1499), .A2(n1544), .A4(n1552), .S0(n283), 
        .S1(n1227), .Y(n2125) );
  AND2X1_HVT U782 ( .A1(n2270), .A2(n234), .Y(n2120) );
  MUX41X1_HVT U784 ( .A1(n2232), .A3(n2120), .A2(n2119), .A4(n2121), .S0(n1232), .S1(n238), .Y(n2118) );
  MUX41X1_HVT U785 ( .A1(n2256), .A3(n1516), .A2(n1523), .A4(n1210), .S0(n1228), .S1(n238), .Y(n2117) );
  MUX41X1_HVT U786 ( .A1(n2117), .A3(n2118), .A2(n2122), .A4(n2125), .S0(n572), 
        .S1(keyin[121]), .Y(n2116) );
  AND2X1_HVT U787 ( .A1(n1234), .A2(n1366), .Y(n2115) );
  NAND2X0_HVT U791 ( .A1(n1425), .A2(n1556), .Y(n2111) );
  MUX41X1_HVT U792 ( .A1(n2263), .A3(n2240), .A2(n2111), .A4(n1545), .S0(n1229), .S1(n238), .Y(n2110) );
  NAND2X0_HVT U793 ( .A1(n1405), .A2(n2218), .Y(n2109) );
  NAND2X0_HVT U797 ( .A1(n1163), .A2(n1428), .Y(n2105) );
  MUX41X1_HVT U798 ( .A1(n1402), .A3(n1542), .A2(n1541), .A4(n2105), .S0(n283), 
        .S1(n1227), .Y(n2104) );
  MUX41X1_HVT U799 ( .A1(n2104), .A3(n2110), .A2(n2106), .A4(n2112), .S0(
        keyin[121]), .S1(n604), .Y(n2103) );
  NAND2X0_HVT U801 ( .A1(n1423), .A2(n2270), .Y(n2262) );
  NAND2X0_HVT U802 ( .A1(n1423), .A2(n1557), .Y(n2102) );
  MUX41X1_HVT U816 ( .A1(n2089), .A3(n1203), .A2(n2262), .A4(n234), .S0(n1230), 
        .S1(n472), .Y(n2088) );
  MUX41X1_HVT U820 ( .A1(n1548), .A3(n2245), .A2(n1402), .A4(n2086), .S0(n1230), .S1(n472), .Y(n2085) );
  AO21X1_HVT U828 ( .A1(n1208), .A2(n1233), .A3(n1539), .Y(n2077) );
  MUX41X1_HVT U830 ( .A1(n1507), .A3(n2270), .A2(n1550), .A4(n2277), .S0(n1230), .S1(n472), .Y(n2075) );
  MUX41X1_HVT U831 ( .A1(n2274), .A3(n2263), .A2(n1522), .A4(n2255), .S0(n1230), .S1(n472), .Y(n2074) );
  MUX41X1_HVT U832 ( .A1(n1368), .A3(n2219), .A2(n1551), .A4(n1526), .S0(n1230), .S1(n472), .Y(n2073) );
  NAND2X0_HVT U837 ( .A1(n1404), .A2(n1426), .Y(n2218) );
  NAND2X0_HVT U838 ( .A1(n1422), .A2(n1397), .Y(n2163) );
  NAND2X0_HVT U841 ( .A1(n2270), .A2(n1428), .Y(n2071) );
  NAND2X0_HVT U842 ( .A1(n1403), .A2(n2163), .Y(n2070) );
  NAND2X0_HVT U845 ( .A1(n1424), .A2(n1552), .Y(n2123) );
  NAND2X0_HVT U847 ( .A1(n1234), .A2(n2071), .Y(n2201) );
  NAND2X0_HVT U942 ( .A1(n1467), .A2(n1390), .Y(n2056) );
  NAND2X0_HVT U943 ( .A1(n1472), .A2(n1362), .Y(n2054) );
  NAND2X0_HVT U944 ( .A1(n1387), .A2(n1470), .Y(n2053) );
  NAND2X0_HVT U945 ( .A1(n1393), .A2(n2056), .Y(n2052) );
  NAND2X0_HVT U952 ( .A1(n2045), .A2(n1396), .Y(n2046) );
  NAND2X0_HVT U954 ( .A1(n2056), .A2(n1757), .Y(n2043) );
  NAND2X0_HVT U960 ( .A1(n1392), .A2(n1472), .Y(n2037) );
  NAND2X0_HVT U963 ( .A1(n1386), .A2(n1472), .Y(n2035) );
  NAND2X0_HVT U971 ( .A1(n1753), .A2(n1472), .Y(n2026) );
  NAND2X0_HVT U977 ( .A1(n1468), .A2(n1360), .Y(n2020) );
  MUX41X1_HVT U990 ( .A1(n1740), .A3(n1698), .A2(n2039), .A4(n1716), .S0(n1479), .S1(n1345), .Y(n2010) );
  NAND2X0_HVT U992 ( .A1(n2007), .A2(n2017), .Y(n2008) );
  NAND2X0_HVT U995 ( .A1(n1393), .A2(n2003), .Y(n2004) );
  MUX41X1_HVT U996 ( .A1(n1741), .A3(n1715), .A2(n2004), .A4(n2048), .S0(n1348), .S1(n1345), .Y(n2002) );
  NAND2X0_HVT U997 ( .A1(n1396), .A2(n2056), .Y(n2001) );
  MUX41X1_HVT U998 ( .A1(n1225), .A3(n2001), .A2(n1220), .A4(n1714), .S0(n1348), .S1(n1345), .Y(n2000) );
  MUX41X1_HVT U1000 ( .A1(n1201), .A3(n1713), .A2(n1712), .A4(n1361), .S0(
        n1348), .S1(n1345), .Y(n1998) );
  NAND2X0_HVT U1001 ( .A1(n1472), .A2(n1391), .Y(n1997) );
  MUX41X1_HVT U1002 ( .A1(n1997), .A3(n1704), .A2(n1735), .A4(n1711), .S0(
        n1348), .S1(n1344), .Y(n1996) );
  AO21X1_HVT U1005 ( .A1(n1709), .A2(n1347), .A3(n1734), .Y(n1993) );
  MUX41X1_HVT U1007 ( .A1(n1707), .A3(n1993), .A2(n1992), .A4(n1994), .S0(
        n1338), .S1(n240), .Y(n1991) );
  MUX41X1_HVT U1008 ( .A1(n1991), .A3(n1999), .A2(n1995), .A4(n2005), .S0(n573), .S1(n1385), .Y(dummy[31]) );
  NAND2X0_HVT U1012 ( .A1(n2057), .A2(n1986), .Y(n1987) );
  MUX41X1_HVT U1013 ( .A1(n1988), .A3(n2015), .A2(n1987), .A4(n2035), .S0(
        n1338), .S1(n866), .Y(n1985) );
  MUX41X1_HVT U1014 ( .A1(n1738), .A3(n1743), .A2(n1756), .A4(n1718), .S0(
        n1338), .S1(n240), .Y(n1984) );
  MUX41X1_HVT U1016 ( .A1(n2049), .A3(n1745), .A2(n1983), .A4(n1744), .S0(
        n1348), .S1(n1473), .Y(n1982) );
  MUX41X1_HVT U1017 ( .A1(n1982), .A3(n1985), .A2(n1984), .A4(n1989), .S0(
        keyin[103]), .S1(n1345), .Y(n1981) );
  AND3X1_HVT U1019 ( .A1(n2003), .A2(n1390), .A3(n1978), .Y(n1979) );
  MUX41X1_HVT U1021 ( .A1(n2014), .A3(n1716), .A2(n1699), .A4(n2044), .S0(
        n1338), .S1(n1476), .Y(n1976) );
  AND2X1_HVT U1022 ( .A1(n290), .A2(n1389), .Y(n1975) );
  MUX41X1_HVT U1023 ( .A1(n1717), .A3(n254), .A2(n2042), .A4(n1975), .S0(n1338), .S1(n1477), .Y(n1974) );
  NAND2X0_HVT U1024 ( .A1(n1472), .A2(n1755), .Y(n1973) );
  MUX41X1_HVT U1025 ( .A1(n1743), .A3(n1973), .A2(n1206), .A4(n1200), .S0(
        n1339), .S1(n1476), .Y(n1972) );
  MUX41X1_HVT U1026 ( .A1(n1972), .A3(n1976), .A2(n1974), .A4(n1977), .S0(
        n1385), .S1(n1345), .Y(n1971) );
  MUX41X1_HVT U1029 ( .A1(n2013), .A3(n2053), .A2(n1740), .A4(n1970), .S0(
        n1338), .S1(n1476), .Y(n1969) );
  AO21X1_HVT U1032 ( .A1(n1350), .A2(n1965), .A3(n1739), .Y(n1966) );
  MUX41X1_HVT U1036 ( .A1(n1738), .A3(n1212), .A2(n1468), .A4(n2043), .S0(
        n1338), .S1(n240), .Y(n1961) );
  NAND2X0_HVT U1040 ( .A1(n1956), .A2(n1955), .Y(n1957) );
  MUX41X1_HVT U1042 ( .A1(n2056), .A3(n1708), .A2(n1720), .A4(n2054), .S0(
        n1338), .S1(n1477), .Y(n1953) );
  OA21X1_HVT U1048 ( .A1(n1727), .A2(n1475), .A3(n1714), .Y(n1948) );
  NAND2X0_HVT U1049 ( .A1(n1390), .A2(n1946), .Y(n1947) );
  MUX41X1_HVT U1053 ( .A1(n1943), .A3(n1949), .A2(n1945), .A4(n1948), .S0(
        n1347), .S1(n1477), .Y(n1942) );
  AND2X1_HVT U1054 ( .A1(n291), .A2(n1361), .Y(n1941) );
  MUX41X1_HVT U1055 ( .A1(n2046), .A3(n1941), .A2(n1718), .A4(n2028), .S0(
        n1339), .S1(n1477), .Y(n1940) );
  AO21X1_HVT U1057 ( .A1(n1343), .A2(n1394), .A3(n254), .Y(n1938) );
  MUX21X2_HVT U1059 ( .A1(n1937), .A2(n1940), .S0(n1347), .Y(n1936) );
  NAND2X0_HVT U1062 ( .A1(n1932), .A2(n1931), .Y(n1933) );
  MUX41X1_HVT U1064 ( .A1(n2037), .A3(n1225), .A2(n1707), .A4(n1747), .S0(
        n1339), .S1(n1476), .Y(n1929) );
  MUX21X2_HVT U1065 ( .A1(n1929), .A2(n1930), .S0(n1347), .Y(n1928) );
  AND3X1_HVT U1067 ( .A1(n1342), .A2(n1472), .A3(n1388), .Y(n1926) );
  MUX41X1_HVT U1070 ( .A1(n1924), .A3(n1926), .A2(n1925), .A4(n1927), .S0(
        n1347), .S1(n1478), .Y(n1923) );
  MUX41X1_HVT U1071 ( .A1(n1923), .A3(n1936), .A2(n1928), .A4(n1942), .S0(
        keyin[97]), .S1(keyin[103]), .Y(dummy[28]) );
  MUX41X1_HVT U1074 ( .A1(n1748), .A3(n1752), .A2(n2020), .A4(n2032), .S0(
        n1340), .S1(n240), .Y(n1920) );
  MUX41X1_HVT U1075 ( .A1(n1200), .A3(n2026), .A2(n1749), .A4(n2024), .S0(
        n1339), .S1(n1479), .Y(n1919) );
  MUX41X1_HVT U1078 ( .A1(n1917), .A3(n1920), .A2(n1919), .A4(n1921), .S0(
        n1385), .S1(n1344), .Y(n1916) );
  AND2X1_HVT U1079 ( .A1(n1394), .A2(n1471), .Y(n1915) );
  MUX41X1_HVT U1080 ( .A1(n2034), .A3(n1728), .A2(n1915), .A4(n1724), .S0(
        n1340), .S1(n1478), .Y(n1914) );
  MUX41X1_HVT U1081 ( .A1(n1717), .A3(n1361), .A2(n1736), .A4(n1394), .S0(
        n1339), .S1(n1479), .Y(n1913) );
  OA21X1_HVT U1083 ( .A1(n1701), .A2(n1480), .A3(n2028), .Y(n1911) );
  NAND2X0_HVT U1085 ( .A1(n1468), .A2(n1396), .Y(n1986) );
  MUX41X1_HVT U1086 ( .A1(n1749), .A3(n1986), .A2(n1738), .A4(n2013), .S0(
        n1340), .S1(n1479), .Y(n1909) );
  MUX41X1_HVT U1087 ( .A1(n1909), .A3(n1913), .A2(n1910), .A4(n1914), .S0(
        n1385), .S1(n1344), .Y(n1908) );
  OA21X1_HVT U1090 ( .A1(n2019), .A2(n1480), .A3(n1905), .Y(n1906) );
  AND2X1_HVT U1093 ( .A1(n1350), .A2(n1386), .Y(n1902) );
  NAND2X0_HVT U1097 ( .A1(n290), .A2(n1755), .Y(n1898) );
  MUX41X1_HVT U1098 ( .A1(n2046), .A3(n1361), .A2(n1898), .A4(n1730), .S0(
        n1340), .S1(n240), .Y(n1897) );
  NAND2X0_HVT U1105 ( .A1(n1396), .A2(n2003), .Y(n1891) );
  NAND2X0_HVT U1106 ( .A1(n1756), .A2(n1472), .Y(n1890) );
  MUX41X1_HVT U1107 ( .A1(n1741), .A3(n1394), .A2(n1890), .A4(n1891), .S0(
        n1133), .S1(n866), .Y(n1889) );
  OA21X1_HVT U1109 ( .A1(n1220), .A2(n1480), .A3(n2028), .Y(n1887) );
  MUX41X1_HVT U1111 ( .A1(n1886), .A3(n1892), .A2(n1889), .A4(n1894), .S0(
        n1385), .S1(n1346), .Y(n1885) );
  NAND2X0_HVT U1113 ( .A1(n1468), .A2(n2033), .Y(n2045) );
  MUX41X1_HVT U1115 ( .A1(n1363), .A3(n1884), .A2(n1746), .A4(n2045), .S0(
        n1479), .S1(n1473), .Y(n1883) );
  NAND2X0_HVT U1116 ( .A1(n291), .A2(n1363), .Y(n1882) );
  MUX41X1_HVT U1117 ( .A1(n2041), .A3(n1882), .A2(n1750), .A4(n2022), .S0(
        n1133), .S1(n1479), .Y(n1881) );
  MUX41X1_HVT U1118 ( .A1(n2031), .A3(n1751), .A2(n1702), .A4(n1750), .S0(
        n1340), .S1(n1477), .Y(n1880) );
  MUX41X1_HVT U1119 ( .A1(n1705), .A3(n2049), .A2(n2046), .A4(n1199), .S0(
        n1479), .S1(n1473), .Y(n1879) );
  MUX41X1_HVT U1120 ( .A1(n1879), .A3(n1881), .A2(n1880), .A4(n1883), .S0(
        n1385), .S1(n1346), .Y(n1878) );
  MUX41X1_HVT U1121 ( .A1(n1729), .A3(n1393), .A2(n1732), .A4(n1733), .S0(
        n1479), .S1(n1473), .Y(n1877) );
  OA21X1_HVT U1123 ( .A1(n2025), .A2(n1480), .A3(n1717), .Y(n1875) );
  MUX41X1_HVT U1125 ( .A1(n1212), .A3(n2021), .A2(n1986), .A4(n2013), .S0(
        n1133), .S1(n240), .Y(n1873) );
  MUX41X1_HVT U1128 ( .A1(n1871), .A3(n2045), .A2(n1872), .A4(n1737), .S0(
        n1479), .S1(n1473), .Y(n1870) );
  MUX41X1_HVT U1129 ( .A1(n1870), .A3(n1873), .A2(n1874), .A4(n1877), .S0(
        n1346), .S1(n1385), .Y(n1869) );
  MUX21X2_HVT U1130 ( .A1(n1869), .A2(n1878), .S0(keyin[97]), .Y(dummy[25]) );
  MUX41X1_HVT U1132 ( .A1(n2053), .A3(n2054), .A2(n2011), .A4(n1868), .S0(
        n1473), .S1(n1476), .Y(n1867) );
  MUX41X1_HVT U1133 ( .A1(n2018), .A3(n2032), .A2(n1748), .A4(n1394), .S0(
        n1479), .S1(n1473), .Y(n1866) );
  MUX41X1_HVT U1134 ( .A1(n254), .A3(n1742), .A2(n2058), .A4(n2023), .S0(n1133), .S1(n866), .Y(n1865) );
  AO21X1_HVT U1136 ( .A1(n1206), .A2(n1349), .A3(n1739), .Y(n1863) );
  MUX41X1_HVT U1138 ( .A1(n1862), .A3(n1866), .A2(n1865), .A4(n1867), .S0(
        keyin[103]), .S1(n1346), .Y(n1861) );
  OA21X1_HVT U1140 ( .A1(n2050), .A2(n1480), .A3(n1728), .Y(n1859) );
  MUX41X1_HVT U1142 ( .A1(n2024), .A3(n1731), .A2(n2047), .A4(n2027), .S0(
        n1133), .S1(n866), .Y(n1857) );
  MUX41X1_HVT U1143 ( .A1(n2004), .A3(n2046), .A2(n1725), .A4(n2036), .S0(
        n1133), .S1(n1477), .Y(n1856) );
  MUX41X1_HVT U1144 ( .A1(n1389), .A3(n2056), .A2(n1751), .A4(n1723), .S0(
        n1133), .S1(n1476), .Y(n1855) );
  MUX41X1_HVT U1145 ( .A1(n1855), .A3(n1857), .A2(n1856), .A4(n1858), .S0(
        n1385), .S1(n1346), .Y(n1854) );
  MUX21X2_HVT U1146 ( .A1(n1854), .A2(n1861), .S0(keyin[97]), .Y(dummy[24]) );
  NAND2X0_HVT U1147 ( .A1(n1467), .A2(n1392), .Y(n1946) );
  NAND2X0_HVT U1150 ( .A1(n1395), .A2(n290), .Y(n2003) );
  NAND2X0_HVT U1152 ( .A1(n254), .A2(n1472), .Y(n1853) );
  NAND2X0_HVT U1153 ( .A1(n2057), .A2(n1946), .Y(n1852) );
  AO21X1_HVT U1154 ( .A1(n1471), .A2(n1752), .A3(n1480), .Y(n1956) );
  NAND2X0_HVT U1156 ( .A1(n1469), .A2(n1752), .Y(n1905) );
  NAND2X0_HVT U1159 ( .A1(n1349), .A2(n1853), .Y(n1978) );
  XOR2X2_HVT U1256 ( .A1(n867), .A2(n1829), .Y(keyout[94]) );
  XOR2X2_HVT U1257 ( .A1(keyout[29]), .A2(n1828), .Y(keyout[93]) );
  XOR2X2_HVT U1260 ( .A1(keyout[26]), .A2(n1825), .Y(keyout[90]) );
  XOR2X2_HVT U1279 ( .A1(keyin[71]), .A2(keyout[39]), .Y(keyout[71]) );
  XOR3X2_HVT U1281 ( .A1(keyin[67]), .A2(n1839), .A3(n1840), .Y(keyout[67]) );
  XOR2X2_HVT U1296 ( .A1(n1492), .A2(keyin[54]), .Y(keyout[54]) );
  XOR2X2_HVT U1303 ( .A1(keyin[48]), .A2(n1496), .Y(keyout[48]) );
  XOR2X2_HVT U1306 ( .A1(keyin[45]), .A2(n863), .Y(keyout[45]) );
  XOR2X2_HVT U1315 ( .A1(n1803), .A2(n1627), .Y(keyout[36]) );
  XOR2X2_HVT U1317 ( .A1(dummy[3]), .A2(keyin[3]), .Y(n1839) );
  XOR2X2_HVT U1321 ( .A1(keyout[1]), .A2(keyin[33]), .Y(keyout[33]) );
  XOR2X2_HVT U1324 ( .A1(dummy[2]), .A2(keyin[2]), .Y(n1835) );
  XNOR2X2_HVT U1325 ( .A1(n1802), .A2(n1834), .Y(keyout[1]) );
  XOR2X2_HVT U1326 ( .A1(dummy[1]), .A2(keyin[1]), .Y(n1834) );
  XNOR2X2_HVT U1327 ( .A1(keyin[31]), .A2(dummy[31]), .Y(n1787) );
  XNOR2X2_HVT U1331 ( .A1(dummy[29]), .A2(keyin[29]), .Y(n1784) );
  XNOR2X2_HVT U1333 ( .A1(dummy[28]), .A2(keyin[28]), .Y(n1783) );
  XNOR2X2_HVT U1335 ( .A1(dummy[27]), .A2(keyin[27]), .Y(n1782) );
  XNOR2X2_HVT U1337 ( .A1(dummy[26]), .A2(keyin[26]), .Y(n1781) );
  XNOR2X2_HVT U1339 ( .A1(keyin[25]), .A2(dummy[25]), .Y(n1780) );
  XNOR2X2_HVT U1341 ( .A1(keyin[24]), .A2(dummy[24]), .Y(n1779) );
  XNOR2X2_HVT U1343 ( .A1(dummy[23]), .A2(keyin[23]), .Y(n1778) );
  XNOR2X2_HVT U1347 ( .A1(dummy[21]), .A2(keyin[21]), .Y(n1776) );
  XNOR2X2_HVT U1355 ( .A1(dummy[17]), .A2(keyin[17]), .Y(n1772) );
  XNOR2X2_HVT U1359 ( .A1(dummy[15]), .A2(keyin[15]), .Y(n1770) );
  XNOR2X2_HVT U1361 ( .A1(dummy[14]), .A2(keyin[14]), .Y(n1769) );
  XNOR2X2_HVT U1365 ( .A1(dummy[12]), .A2(keyin[12]), .Y(n1767) );
  XNOR2X2_HVT U1367 ( .A1(dummy[11]), .A2(keyin[11]), .Y(n1766) );
  XNOR2X2_HVT U1369 ( .A1(dummy[10]), .A2(keyin[10]), .Y(n1765) );
  XNOR2X2_HVT U1371 ( .A1(dummy[9]), .A2(keyin[9]), .Y(n1797) );
  XNOR2X2_HVT U1373 ( .A1(dummy[8]), .A2(keyin[8]), .Y(n1796) );
  XNOR2X2_HVT U1375 ( .A1(keyout[7]), .A2(keyin[39]), .Y(n1794) );
  XOR3X2_HVT U1376 ( .A1(keyin[7]), .A2(n1764), .A3(dummy[7]), .Y(keyout[7])
         );
  XNOR2X2_HVT U1384 ( .A1(dummy[4]), .A2(keyin[4]), .Y(n1804) );
  XNOR2X2_HVT U1386 ( .A1(n1832), .A2(n1801), .Y(keyout[0]) );
  XOR2X2_HVT U1387 ( .A1(dummy[0]), .A2(keyin[0]), .Y(n1832) );
  XNOR3X1_HVT U1427 ( .A1(keyin[70]), .A2(n1486), .A3(n821), .Y(keyout[70]) );
  XNOR3X1_HVT U1428 ( .A1(keyin[69]), .A2(n1483), .A3(n1626), .Y(keyout[69])
         );
  XNOR3X1_HVT U1430 ( .A1(keyin[32]), .A2(keyin[64]), .A3(n1801), .Y(n1831) );
  NAND3X0_HVT U1431 ( .A1(n1791), .A2(n1790), .A3(n1789), .Y(n1795) );
  NAND4X0_HVT U1432 ( .A1(round_num[1]), .A2(round_num[3]), .A3(n1488), .A4(
        n1490), .Y(n1789) );
  AO21X1_HVT U1433 ( .A1(n1785), .A2(round_num[2]), .A3(n1482), .Y(n1788) );
  NAND4X0_HVT U1434 ( .A1(round_num[1]), .A2(round_num[2]), .A3(round_num[3]), 
        .A4(n1488), .Y(n1802) );
  XNOR3X1_HVT U1435 ( .A1(n1830), .A2(keyin[127]), .A3(n1787), .Y(keyout[127])
         );
  XNOR3X1_HVT U1436 ( .A1(n1829), .A2(n1422), .A3(n1786), .Y(keyout[126]) );
  XNOR3X1_HVT U1437 ( .A1(n1828), .A2(n604), .A3(n1784), .Y(keyout[125]) );
  XNOR3X1_HVT U1438 ( .A1(n1827), .A2(n1366), .A3(n1783), .Y(keyout[124]) );
  XNOR3X1_HVT U1439 ( .A1(n1826), .A2(n1367), .A3(n1782), .Y(keyout[123]) );
  XNOR3X1_HVT U1440 ( .A1(n1825), .A2(n1228), .A3(n1781), .Y(keyout[122]) );
  XNOR3X1_HVT U1441 ( .A1(n1824), .A2(keyin[121]), .A3(n1780), .Y(keyout[121])
         );
  XNOR3X1_HVT U1448 ( .A1(n1817), .A2(n1238), .A3(n869), .Y(keyout[114]) );
  XNOR3X1_HVT U1449 ( .A1(n1816), .A2(n1376), .A3(n865), .Y(keyout[113]) );
  XNOR3X1_HVT U1451 ( .A1(n1814), .A2(n1377), .A3(n1770), .Y(keyout[111]) );
  XNOR3X1_HVT U1452 ( .A1(n1813), .A2(n1456), .A3(n1769), .Y(keyout[110]) );
  XNOR3X1_HVT U1453 ( .A1(n1812), .A2(n901), .A3(n1768), .Y(keyout[109]) );
  XNOR3X1_HVT U1455 ( .A1(n1810), .A2(n1382), .A3(n1766), .Y(keyout[107]) );
  XNOR3X1_HVT U1456 ( .A1(n1809), .A2(n1249), .A3(n1765), .Y(keyout[106]) );
  XNOR3X1_HVT U1457 ( .A1(n1808), .A2(keyin[105]), .A3(n1797), .Y(keyout[105])
         );
  XNOR3X1_HVT U1458 ( .A1(n1807), .A2(n268), .A3(n861), .Y(keyout[104]) );
  XNOR3X1_HVT U1459 ( .A1(keyin[71]), .A2(keyin[103]), .A3(n1794), .Y(
        keyout[103]) );
  AND2X1_HVT U1461 ( .A1(n1790), .A2(n1762), .Y(n1805) );
  NAND3X0_HVT U1462 ( .A1(n1487), .A2(n1489), .A3(round_num[2]), .Y(n1762) );
  AND2X1_HVT U1464 ( .A1(n1791), .A2(n1760), .Y(n1799) );
  NAND4X0_HVT U1465 ( .A1(round_num[2]), .A2(round_num[3]), .A3(n1488), .A4(
        n1487), .Y(n1760) );
  NAND2X0_HVT U1466 ( .A1(round_num[2]), .A2(n1759), .Y(n1791) );
  AO21X1_HVT U1468 ( .A1(n1785), .A2(n1490), .A3(n1485), .Y(n1798) );
  NAND2X0_HVT U1469 ( .A1(round_num[0]), .A2(n1764), .Y(n1790) );
  AND3X1_HVT U1470 ( .A1(n1487), .A2(n1490), .A3(round_num[3]), .Y(n1764) );
  AND3X1_HVT U1471 ( .A1(n1488), .A2(n1489), .A3(round_num[1]), .Y(n1785) );
  NAND2X0_HVT U1472 ( .A1(n1759), .A2(n1490), .Y(n1801) );
  AND3X1_HVT U1473 ( .A1(n1487), .A2(n1489), .A3(round_num[0]), .Y(n1759) );
  MUX21X2_HVT U1 ( .A1(n592), .A2(n591), .S0(n235), .Y(n2192) );
  MUX21X1_HVT U2 ( .A1(n49), .A2(n2456), .S0(n873), .Y(n23) );
  IBUFFX16_HVT U3 ( .A(n1354), .Y(n49) );
  XNOR2X2_HVT U7 ( .A1(keyin[42]), .A2(n1765), .Y(keyout[42]) );
  XOR2X2_HVT U8 ( .A1(dummy[16]), .A2(n211), .Y(n1771) );
  IBUFFX16_HVT U9 ( .A(keyin[16]), .Y(n211) );
  INVX0_HVT U10 ( .A(n1427), .Y(n1423) );
  INVX0_HVT U11 ( .A(n1534), .Y(n234) );
  IBUFFX2_HVT U12 ( .A(n866), .Y(n242) );
  MUX21X2_HVT U13 ( .A1(n1542), .A2(n2242), .S0(n212), .Y(n2078) );
  IBUFFX16_HVT U14 ( .A(n264), .Y(n212) );
  XNOR2X2_HVT U16 ( .A1(n213), .A2(n2252), .Y(n2234) );
  IBUFFX16_HVT U18 ( .A(n1435), .Y(n213) );
  INVX1_HVT U19 ( .A(n1495), .Y(n865) );
  XNOR2X2_HVT U20 ( .A1(keyin[53]), .A2(n1776), .Y(keyout[53]) );
  INVX0_HVT U22 ( .A(n1457), .Y(n214) );
  INVX0_HVT U23 ( .A(n1457), .Y(n217) );
  INVX0_HVT U24 ( .A(n1457), .Y(n1453) );
  NBUFFX2_HVT U26 ( .A(keyin[126]), .Y(n218) );
  IBUFFX2_HVT U27 ( .A(n472), .Y(n235) );
  MUX21X2_HVT U28 ( .A1(n569), .A2(n568), .S0(n219), .Y(n2099) );
  IBUFFX16_HVT U29 ( .A(n238), .Y(n219) );
  MUX21X2_HVT U30 ( .A1(n2202), .A2(n2203), .S0(n220), .Y(n2200) );
  IBUFFX16_HVT U31 ( .A(n1232), .Y(n220) );
  MUX41X1_HVT U32 ( .A1(n2209), .A3(n2204), .A2(n2200), .A4(n2199), .S0(n232), 
        .S1(n233), .Y(n2198) );
  IBUFFX16_HVT U35 ( .A(keyin[125]), .Y(n232) );
  IBUFFX16_HVT U36 ( .A(keyin[121]), .Y(n233) );
  NAND2X2_HVT U37 ( .A1(n1422), .A2(n1400), .Y(n2274) );
  INVX1_HVT U38 ( .A(n1451), .Y(n236) );
  INVX1_HVT U40 ( .A(n1451), .Y(n237) );
  INVX0_HVT U41 ( .A(n1451), .Y(n1449) );
  NBUFFX4_HVT U42 ( .A(keyin[120]), .Y(n238) );
  XOR2X2_HVT U43 ( .A1(dummy[21]), .A2(keyin[21]), .Y(keyout[21]) );
  INVX1_HVT U44 ( .A(keyin[120]), .Y(n1435) );
  IBUFFX2_HVT U45 ( .A(n1480), .Y(n240) );
  MUX41X1_HVT U46 ( .A1(n1737), .A3(n1952), .A2(n2012), .A4(n1719), .S0(n241), 
        .S1(n242), .Y(n1951) );
  IBUFFX16_HVT U47 ( .A(n1338), .Y(n241) );
  INVX0_HVT U48 ( .A(n2708), .Y(n243) );
  INVX2_HVT U49 ( .A(n243), .Y(n244) );
  INVX1_HVT U51 ( .A(n2708), .Y(n1684) );
  MUX21X1_HVT U53 ( .A1(n1380), .A2(n1684), .S0(n245), .Y(n2693) );
  IBUFFX16_HVT U54 ( .A(n1454), .Y(n245) );
  INVX1_HVT U58 ( .A(n2693), .Y(n1649) );
  NBUFFX4_HVT U63 ( .A(keyin[112]), .Y(n862) );
  NBUFFX2_HVT U64 ( .A(n1451), .Y(n280) );
  INVX1_HVT U66 ( .A(n1451), .Y(n1450) );
  INVX2_HVT U68 ( .A(n1427), .Y(n1422) );
  MUX41X1_HVT U70 ( .A1(n2093), .A3(n2092), .A2(n2090), .A4(n2088), .S0(n246), 
        .S1(n516), .Y(n2087) );
  IBUFFX16_HVT U72 ( .A(n474), .Y(n246) );
  IBUFFX2_HVT U73 ( .A(n1445), .Y(n247) );
  MUX21X1_HVT U74 ( .A1(n2532), .A2(n2533), .S0(n1253), .Y(n2531) );
  OA21X1_HVT U75 ( .A1(n2684), .A2(n1466), .A3(n1649), .Y(n2532) );
  MUX41X1_HVT U76 ( .A1(n2358), .A3(n2363), .A2(n2369), .A4(n2377), .S0(n1376), 
        .S1(n248), .Y(n852) );
  IBUFFX16_HVT U78 ( .A(n892), .Y(n248) );
  XOR3X1_HVT U79 ( .A1(n249), .A2(n250), .A3(n875), .Y(keyout[108]) );
  IBUFFX16_HVT U87 ( .A(n1811), .Y(n249) );
  IBUFFX16_HVT U88 ( .A(n255), .Y(n250) );
  INVX0_HVT U89 ( .A(n1466), .Y(n251) );
  INVX0_HVT U90 ( .A(n1466), .Y(n252) );
  INVX0_HVT U91 ( .A(n1466), .Y(n1465) );
  INVX1_HVT U92 ( .A(n875), .Y(keyout[12]) );
  INVX1_HVT U93 ( .A(n2033), .Y(n253) );
  INVX2_HVT U94 ( .A(n253), .Y(n254) );
  IBUFFX16_HVT U95 ( .A(n1379), .Y(n255) );
  MUX21X2_HVT U96 ( .A1(n1387), .A2(n1361), .S0(n256), .Y(n2036) );
  IBUFFX16_HVT U98 ( .A(n1470), .Y(n256) );
  INVX1_HVT U99 ( .A(n1427), .Y(n1425) );
  INVX1_HVT U100 ( .A(n1427), .Y(n1424) );
  MUX41X1_HVT U101 ( .A1(n2188), .A3(n2185), .A2(n2186), .A4(n2184), .S0(n257), 
        .S1(n258), .Y(n2182) );
  IBUFFX16_HVT U103 ( .A(n572), .Y(n257) );
  IBUFFX16_HVT U105 ( .A(n1226), .Y(n258) );
  MUX41X1_HVT U107 ( .A1(n2358), .A3(n2363), .A2(n2369), .A4(n2377), .S0(n1376), .S1(n259), .Y(dummy[12]) );
  IBUFFX16_HVT U108 ( .A(n892), .Y(n259) );
  MUX21X1_HVT U109 ( .A1(n2370), .A2(n2371), .S0(n1236), .Y(n2369) );
  MUX21X2_HVT U110 ( .A1(n2266), .A2(n2243), .S0(n260), .Y(n2082) );
  IBUFFX16_HVT U112 ( .A(n1234), .Y(n260) );
  MUX21X1_HVT U113 ( .A1(n1363), .A2(n1361), .S0(n261), .Y(n1955) );
  IBUFFX16_HVT U114 ( .A(n1468), .Y(n261) );
  MUX21X2_HVT U116 ( .A1(n1722), .A2(n1957), .S0(n262), .Y(n1954) );
  IBUFFX16_HVT U117 ( .A(n1342), .Y(n262) );
  MUX41X1_HVT U119 ( .A1(n2167), .A3(n2176), .A2(n2171), .A4(n2182), .S0(
        keyin[127]), .S1(n263), .Y(dummy[21]) );
  IBUFFX16_HVT U121 ( .A(n594), .Y(n263) );
  IBUFFX16_HVT U123 ( .A(n1233), .Y(n264) );
  MUX41X1_HVT U124 ( .A1(n2076), .A3(n2074), .A2(n2075), .A4(n2073), .S0(n265), 
        .S1(n266), .Y(n2072) );
  IBUFFX16_HVT U126 ( .A(keyin[121]), .Y(n265) );
  IBUFFX16_HVT U127 ( .A(n572), .Y(n266) );
  MUX21X2_HVT U128 ( .A1(n2081), .A2(n2082), .S0(n267), .Y(n2080) );
  IBUFFX16_HVT U130 ( .A(n1232), .Y(n267) );
  OA21X1_HVT U131 ( .A1(n2269), .A2(n1435), .A3(n1530), .Y(n2081) );
  INVX1_HVT U135 ( .A(n285), .Y(n268) );
  INVX0_HVT U136 ( .A(n555), .Y(n285) );
  INVX1_HVT U141 ( .A(n2498), .Y(n1679) );
  IBUFFX2_HVT U142 ( .A(n1445), .Y(n1443) );
  INVX4_HVT U145 ( .A(keyin[117]), .Y(n1445) );
  MUX21X2_HVT U146 ( .A1(n1193), .A2(n2261), .S0(n269), .Y(n2181) );
  IBUFFX16_HVT U147 ( .A(n1234), .Y(n269) );
  XOR2X2_HVT U149 ( .A1(n1357), .A2(n1382), .Y(n2708) );
  NBUFFX4_HVT U150 ( .A(n1686), .Y(n1357) );
  INVX2_HVT U152 ( .A(n279), .Y(n270) );
  INVX1_HVT U153 ( .A(n554), .Y(n279) );
  XOR3X2_HVT U154 ( .A1(n1834), .A2(n271), .A3(n1833), .Y(keyout[97]) );
  IBUFFX16_HVT U155 ( .A(n573), .Y(n271) );
  MUX21X2_HVT U157 ( .A1(n1753), .A2(n1361), .S0(n272), .Y(n1963) );
  IBUFFX16_HVT U162 ( .A(n1469), .Y(n272) );
  MUX41X1_HVT U163 ( .A1(n1212), .A3(n1699), .A2(n1963), .A4(n1742), .S0(n273), 
        .S1(n866), .Y(n1962) );
  IBUFFX16_HVT U164 ( .A(n1340), .Y(n273) );
  MUX21X2_HVT U168 ( .A1(n2672), .A2(n2643), .S0(n274), .Y(n2642) );
  IBUFFX16_HVT U169 ( .A(n1252), .Y(n274) );
  MUX41X1_HVT U170 ( .A1(n2642), .A3(n2647), .A2(n2637), .A4(n2638), .S0(n901), 
        .S1(n275), .Y(n2636) );
  IBUFFX16_HVT U173 ( .A(keyin[105]), .Y(n275) );
  IBUFFX2_HVT U174 ( .A(n1480), .Y(n866) );
  IBUFFX2_HVT U178 ( .A(n1480), .Y(n1476) );
  IBUFFX2_HVT U181 ( .A(n1480), .Y(n1477) );
  INVX1_HVT U182 ( .A(n1457), .Y(n1456) );
  INVX1_HVT U183 ( .A(n1457), .Y(n1455) );
  XNOR2X2_HVT U187 ( .A1(keyout[0]), .A2(n276), .Y(keyout[32]) );
  IBUFFX16_HVT U189 ( .A(keyin[32]), .Y(n276) );
  NBUFFX2_HVT U192 ( .A(n214), .Y(n277) );
  MUX41X1_HVT U193 ( .A1(n2687), .A3(n1650), .A2(n2588), .A4(n2701), .S0(n278), 
        .S1(n279), .Y(n2587) );
  IBUFFX16_HVT U197 ( .A(n1460), .Y(n278) );
  INVX1_HVT U198 ( .A(keyin[112]), .Y(n1451) );
  INVX0_HVT U199 ( .A(n873), .Y(n293) );
  INVX0_HVT U201 ( .A(n289), .Y(n281) );
  MUX21X2_HVT U203 ( .A1(n2513), .A2(n2514), .S0(n1252), .Y(n2512) );
  XOR2X2_HVT U207 ( .A1(n1831), .A2(n1832), .Y(keyout[64]) );
  OA21X1_HVT U208 ( .A1(n1570), .A2(n280), .A3(n2466), .Y(n2346) );
  IBUFFX16_HVT U209 ( .A(n1466), .Y(n1464) );
  INVX2_HVT U210 ( .A(keyin[126]), .Y(n1427) );
  MUX41X1_HVT U213 ( .A1(n2179), .A3(n1524), .A2(n2180), .A4(n2181), .S0(n572), 
        .S1(n1431), .Y(n2176) );
  MUX41X1_HVT U214 ( .A1(n2652), .A3(n2648), .A2(n2662), .A4(n2658), .S0(n595), 
        .S1(n282), .Y(dummy[7]) );
  IBUFFX16_HVT U217 ( .A(n596), .Y(n282) );
  MUX21X1_HVT U218 ( .A1(n2661), .A2(n2659), .S0(n549), .Y(n2658) );
  INVX1_HVT U220 ( .A(n1441), .Y(n1438) );
  INVX0_HVT U222 ( .A(n1441), .Y(n1439) );
  INVX1_HVT U223 ( .A(n1441), .Y(n1436) );
  NBUFFX2_HVT U224 ( .A(keyin[120]), .Y(n283) );
  MUX41X1_HVT U225 ( .A1(n2259), .A3(n1195), .A2(n1532), .A4(n2247), .S0(n283), 
        .S1(n284), .Y(n2083) );
  IBUFFX16_HVT U226 ( .A(n1226), .Y(n284) );
  INVX2_HVT U227 ( .A(n1441), .Y(n1437) );
  INVX1_HVT U228 ( .A(n2283), .Y(n1592) );
  MUX21X2_HVT U229 ( .A1(n2594), .A2(n2595), .S0(n285), .Y(n2591) );
  MUX21X1_HVT U230 ( .A1(n2587), .A2(n2584), .S0(n844), .Y(n2583) );
  INVX1_HVT U231 ( .A(n1769), .Y(keyout[14]) );
  MUX21X2_HVT U232 ( .A1(n2612), .A2(n1204), .S0(n288), .Y(n2611) );
  IBUFFX2_HVT U233 ( .A(n1255), .Y(n288) );
  MUX21X2_HVT U234 ( .A1(n2698), .A2(n2613), .S0(n1253), .Y(n2612) );
  MUX41X1_HVT U235 ( .A1(n2348), .A3(n2344), .A2(n2349), .A4(n2345), .S0(n286), 
        .S1(n1443), .Y(n2343) );
  IBUFFX16_HVT U236 ( .A(keyin[113]), .Y(n286) );
  MUX21X2_HVT U237 ( .A1(n2313), .A2(n2306), .S0(n287), .Y(dummy[9]) );
  IBUFFX16_HVT U238 ( .A(n1370), .Y(n287) );
  NAND2X0_HVT U239 ( .A1(n588), .A2(n589), .Y(n289) );
  INVX0_HVT U240 ( .A(n1471), .Y(n290) );
  INVX1_HVT U241 ( .A(n1471), .Y(n291) );
  MUX21X1_HVT U242 ( .A1(n1757), .A2(n1395), .S0(n292), .Y(n1952) );
  IBUFFX16_HVT U243 ( .A(n1469), .Y(n292) );
  INVX0_HVT U244 ( .A(n1471), .Y(n1468) );
  NAND2X0_HVT U245 ( .A1(n2552), .A2(n1175), .Y(n1176) );
  INVX2_HVT U246 ( .A(n1457), .Y(n1454) );
  INVX2_HVT U247 ( .A(keyin[110]), .Y(n1457) );
  MUX21X2_HVT U248 ( .A1(n2392), .A2(n1202), .S0(n293), .Y(n2391) );
  MUX21X2_HVT U249 ( .A1(n2343), .A2(n2351), .S0(n294), .Y(dummy[11]) );
  IBUFFX16_HVT U250 ( .A(n1184), .Y(n294) );
  MUX21X1_HVT U251 ( .A1(n296), .A2(n1371), .S0(n543), .Y(n295) );
  IBUFFX16_HVT U252 ( .A(n1375), .Y(n296) );
  INVX1_HVT U253 ( .A(n1244), .Y(n543) );
  MUX41X1_HVT U254 ( .A1(n2569), .A3(n2565), .A2(n2568), .A4(n2564), .S0(n297), 
        .S1(n298), .Y(n2563) );
  IBUFFX16_HVT U255 ( .A(keyin[105]), .Y(n297) );
  IBUFFX16_HVT U256 ( .A(n1460), .Y(n298) );
  XOR3X2_HVT U257 ( .A1(n299), .A2(n1839), .A3(n1838), .Y(keyout[99]) );
  IBUFFX16_HVT U258 ( .A(n1840), .Y(n299) );
  MUX41X1_HVT U259 ( .A1(n2546), .A3(n2540), .A2(n2548), .A4(n2542), .S0(n300), 
        .S1(n301), .Y(n2539) );
  IBUFFX16_HVT U260 ( .A(keyin[105]), .Y(n300) );
  IBUFFX16_HVT U261 ( .A(n843), .Y(n301) );
  NAND2X0_HVT U262 ( .A1(n2523), .A2(n609), .Y(n610) );
  XOR3X1_HVT U263 ( .A1(n302), .A2(keyin[66]), .A3(n1837), .Y(keyout[98]) );
  IBUFFX16_HVT U264 ( .A(n1346), .Y(n302) );
  XNOR2X2_HVT U265 ( .A1(n1836), .A2(n1835), .Y(n1837) );
  INVX2_HVT U266 ( .A(n1471), .Y(n1467) );
  INVX2_HVT U267 ( .A(keyin[102]), .Y(n1471) );
  INVX1_HVT U268 ( .A(n1967), .Y(n522) );
  XOR3X1_HVT U269 ( .A1(n303), .A2(n304), .A3(n305), .Y(keyout[100]) );
  IBUFFX16_HVT U270 ( .A(keyin[68]), .Y(n303) );
  IBUFFX16_HVT U271 ( .A(n1387), .Y(n304) );
  XNOR2X2_HVT U272 ( .A1(n1803), .A2(n1804), .Y(n305) );
  INVX2_HVT U273 ( .A(keyin[96]), .Y(n1481) );
  XOR3X2_HVT U274 ( .A1(keyin[68]), .A2(n328), .A3(n1804), .Y(keyout[68]) );
  IBUFFX16_HVT U275 ( .A(n1803), .Y(n328) );
  XOR2X2_HVT U276 ( .A1(n1798), .A2(n1627), .Y(keyout[4]) );
  MUX21X2_HVT U277 ( .A1(n2407), .A2(n2415), .S0(n354), .Y(dummy[14]) );
  IBUFFX16_HVT U278 ( .A(n903), .Y(n354) );
  MUX21X2_HVT U279 ( .A1(n2611), .A2(n2610), .S0(n398), .Y(n2609) );
  IBUFFX16_HVT U280 ( .A(n1460), .Y(n398) );
  NBUFFX4_HVT U281 ( .A(keyin[120]), .Y(n472) );
  XOR2X2_HVT U282 ( .A1(dummy[22]), .A2(n473), .Y(n1777) );
  IBUFFX16_HVT U283 ( .A(keyin[22]), .Y(n473) );
  IBUFFX16_HVT U284 ( .A(n582), .Y(n474) );
  IBUFFX16_HVT U285 ( .A(keyin[121]), .Y(n516) );
  XNOR2X2_HVT U286 ( .A1(n1765), .A2(n1809), .Y(keyout[74]) );
  INVX1_HVT U287 ( .A(n1765), .Y(keyout[10]) );
  XOR3X2_HVT U288 ( .A1(n1792), .A2(n1761), .A3(n1626), .Y(keyout[101]) );
  XNOR2X2_HVT U289 ( .A1(n1799), .A2(keyin[37]), .Y(n1792) );
  INVX1_HVT U290 ( .A(n2286), .Y(n1609) );
  MUX41X1_HVT U291 ( .A1(n2334), .A3(n2333), .A2(n2342), .A4(n2338), .S0(n1445), .S1(n517), .Y(n2332) );
  IBUFFX16_HVT U292 ( .A(n524), .Y(n517) );
  XOR2X2_HVT U293 ( .A1(n1792), .A2(n281), .Y(keyout[37]) );
  MUX21X1_HVT U294 ( .A1(n1396), .A2(n1393), .S0(n1471), .Y(n1965) );
  MUX21X1_HVT U295 ( .A1(n522), .A2(n519), .S0(n523), .Y(n518) );
  IBUFFX16_HVT U296 ( .A(n518), .Y(n1964) );
  IBUFFX16_HVT U297 ( .A(n1966), .Y(n519) );
  IBUFFX16_HVT U298 ( .A(n1342), .Y(n523) );
  MUX21X2_HVT U299 ( .A1(n1585), .A2(n2478), .S0(n1243), .Y(n2420) );
  IBUFFX16_HVT U300 ( .A(keyin[113]), .Y(n524) );
  INVX0_HVT U301 ( .A(n861), .Y(n525) );
  NBUFFX4_HVT U302 ( .A(n1796), .Y(n861) );
  INVX2_HVT U303 ( .A(n1796), .Y(keyout[8]) );
  MUX21X2_HVT U304 ( .A1(n2300), .A2(n2301), .S0(n537), .Y(n2299) );
  IBUFFX16_HVT U305 ( .A(n1242), .Y(n537) );
  INVX0_HVT U306 ( .A(n543), .Y(n538) );
  MUX41X1_HVT U307 ( .A1(n2480), .A3(n2491), .A2(n2472), .A4(n1590), .S0(n539), 
        .S1(n1450), .Y(n2293) );
  IBUFFX16_HVT U308 ( .A(n1240), .Y(n539) );
  MUX21X1_HVT U309 ( .A1(n2296), .A2(n2297), .S0(n1241), .Y(n2295) );
  MUX41X1_HVT U310 ( .A1(n2294), .A3(n2292), .A2(n2295), .A4(n2293), .S0(n540), 
        .S1(n1443), .Y(n2291) );
  IBUFFX16_HVT U311 ( .A(n1376), .Y(n540) );
  MUX21X1_HVT U312 ( .A1(n2326), .A2(n2327), .S0(n1241), .Y(n2325) );
  INVX4_HVT U313 ( .A(n1784), .Y(keyout[29]) );
  MUX41X1_HVT U314 ( .A1(n1550), .A3(n1195), .A2(n1551), .A4(n2263), .S0(n541), 
        .S1(n1162), .Y(n2093) );
  IBUFFX16_HVT U315 ( .A(n1230), .Y(n541) );
  NBUFFX2_HVT U316 ( .A(keyin[104]), .Y(n542) );
  INVX2_HVT U321 ( .A(keyin[104]), .Y(n1466) );
  MUX21X2_HVT U322 ( .A1(n1609), .A2(n2459), .S0(n873), .Y(n2297) );
  NAND2X0_HVT U323 ( .A1(n2460), .A2(n543), .Y(n544) );
  NAND2X0_HVT U324 ( .A1(n2483), .A2(n1244), .Y(n545) );
  NAND2X0_HVT U325 ( .A1(n544), .A2(n545), .Y(n2301) );
  MUX41X1_HVT U326 ( .A1(n2085), .A3(n2083), .A2(n2084), .A4(n2080), .S0(n594), 
        .S1(n1430), .Y(n2079) );
  MUX21X1_HVT U327 ( .A1(n2273), .A2(n2237), .S0(n548), .Y(n546) );
  MUX21X1_HVT U329 ( .A1(n2230), .A2(n2252), .S0(n548), .Y(n547) );
  MUX21X1_HVT U331 ( .A1(n546), .A2(n547), .S0(n472), .Y(n2084) );
  INVX0_HVT U332 ( .A(keyin[121]), .Y(n594) );
  IBUFFX2_HVT U333 ( .A(n1230), .Y(n548) );
  IBUFFX2_HVT U335 ( .A(keyin[118]), .Y(n1442) );
  XOR2X2_HVT U336 ( .A1(keyout[21]), .A2(n1820), .Y(keyout[85]) );
  IBUFFX2_HVT U337 ( .A(n2483), .Y(n1579) );
  MUX21X2_HVT U339 ( .A1(n2518), .A2(n2517), .S0(n1253), .Y(n2516) );
  IBUFFX16_HVT U340 ( .A(n902), .Y(n549) );
  NAND2X0_HVT U341 ( .A1(n1655), .A2(n550), .Y(n551) );
  NAND2X0_HVT U342 ( .A1(n2576), .A2(n844), .Y(n552) );
  NAND2X0_HVT U343 ( .A1(n551), .A2(n552), .Y(n2575) );
  IBUFFX2_HVT U344 ( .A(n844), .Y(n550) );
  MUX21X2_HVT U345 ( .A1(n2591), .A2(n2590), .S0(n553), .Y(n2589) );
  IBUFFX16_HVT U348 ( .A(n1252), .Y(n553) );
  NBUFFX2_HVT U349 ( .A(n1465), .Y(n554) );
  NBUFFX2_HVT U350 ( .A(n1465), .Y(n555) );
  NBUFFX2_HVT U351 ( .A(n1465), .Y(n556) );
  IBUFFX2_HVT U353 ( .A(n1466), .Y(n1463) );
  NBUFFX2_HVT U354 ( .A(n1467), .Y(n557) );
  NBUFFX2_HVT U355 ( .A(n1467), .Y(n558) );
  NBUFFX2_HVT U356 ( .A(n1467), .Y(n559) );
  IBUFFX2_HVT U357 ( .A(n1471), .Y(n1469) );
  NBUFFX2_HVT U358 ( .A(n1439), .Y(n560) );
  NBUFFX2_HVT U359 ( .A(n1439), .Y(n561) );
  NBUFFX2_HVT U360 ( .A(n1439), .Y(n562) );
  AND3X1_HVT U361 ( .A1(n1418), .A2(n2656), .A3(n2639), .Y(n2640) );
  INVX1_HVT U362 ( .A(n1435), .Y(n1434) );
  INVX0_HVT U364 ( .A(n1380), .Y(n823) );
  INVX0_HVT U366 ( .A(n1440), .Y(n580) );
  INVX1_HVT U367 ( .A(n579), .Y(n1187) );
  MUX21X1_HVT U371 ( .A1(n1196), .A2(n1653), .S0(n1255), .Y(n2618) );
  OA21X1_HVT U376 ( .A1(n280), .A2(n2486), .A3(n1598), .Y(n2300) );
  INVX0_HVT U377 ( .A(n1228), .Y(n583) );
  OA21X1_HVT U379 ( .A1(n1218), .A2(n280), .A3(n2466), .Y(n2326) );
  OA21X1_HVT U383 ( .A1(n2455), .A2(n280), .A3(n2339), .Y(n2340) );
  MUX21X1_HVT U385 ( .A1(n1660), .A2(n1414), .S0(n1254), .Y(n2533) );
  MUX21X1_HVT U386 ( .A1(n2058), .A2(n1395), .S0(n557), .Y(n2028) );
  XOR2X1_HVT U387 ( .A1(n1480), .A2(n2032), .Y(n2016) );
  INVX1_HVT U389 ( .A(n1475), .Y(n1474) );
  MUX21X1_HVT U392 ( .A1(n1673), .A2(n2680), .S0(n270), .Y(n2514) );
  INVX1_HVT U400 ( .A(keyin[101]), .Y(n1475) );
  INVX1_HVT U401 ( .A(n1377), .Y(n596) );
  INVX1_HVT U402 ( .A(n830), .Y(n824) );
  NAND2X0_HVT U403 ( .A1(n912), .A2(n911), .Y(n2138) );
  NAND2X0_HVT U404 ( .A1(n2628), .A2(n601), .Y(n602) );
  INVX1_HVT U405 ( .A(n893), .Y(n600) );
  INVX1_HVT U408 ( .A(keyin[20]), .Y(n571) );
  INVX1_HVT U409 ( .A(n1794), .Y(keyout[39]) );
  INVX2_HVT U411 ( .A(n1481), .Y(n1478) );
  INVX0_HVT U412 ( .A(n1836), .Y(n563) );
  INVX0_HVT U413 ( .A(n1242), .Y(n581) );
  INVX0_HVT U414 ( .A(n2033), .Y(n1757) );
  INVX1_HVT U416 ( .A(n1245), .Y(n590) );
  XNOR3X1_HVT U418 ( .A1(n1823), .A2(n283), .A3(n1779), .Y(keyout[120]) );
  INVX1_HVT U420 ( .A(n1214), .Y(n577) );
  INVX1_HVT U421 ( .A(n1344), .Y(n564) );
  INVX1_HVT U422 ( .A(n901), .Y(n843) );
  INVX0_HVT U423 ( .A(keyin[125]), .Y(n582) );
  INVX0_HVT U425 ( .A(n1430), .Y(n572) );
  INVX1_HVT U426 ( .A(n582), .Y(n604) );
  INVX1_HVT U427 ( .A(n1371), .Y(n599) );
  INVX1_HVT U428 ( .A(keyin[105]), .Y(n595) );
  INVX0_HVT U429 ( .A(n1473), .Y(n584) );
  INVX1_HVT U430 ( .A(n1247), .Y(n844) );
  INVX1_HVT U432 ( .A(n1364), .Y(n856) );
  INVX0_HVT U434 ( .A(keyin[127]), .Y(n1148) );
  INVX0_HVT U437 ( .A(keyin[97]), .Y(n593) );
  MUX21X2_HVT U439 ( .A1(n1938), .A2(n1939), .S0(n1349), .Y(n1937) );
  MUX41X1_HVT U440 ( .A1(n2620), .A3(n2609), .A2(n2614), .A4(n2605), .S0(n1178), .S1(n595), .Y(dummy[5]) );
  XNOR2X2_HVT U441 ( .A1(n563), .A2(n1835), .Y(keyout[34]) );
  MUX41X1_HVT U443 ( .A1(n1969), .A3(n1962), .A2(n1964), .A4(n1961), .S0(n884), 
        .S1(n564), .Y(n1960) );
  MUX41X1_HVT U444 ( .A1(n1402), .A3(n2257), .A2(n1498), .A4(n2233), .S0(n1162), .S1(n907), .Y(n2199) );
  XNOR2X2_HVT U446 ( .A1(keyin[52]), .A2(n1775), .Y(keyout[52]) );
  INVX1_HVT U448 ( .A(n1775), .Y(keyout[20]) );
  XOR2X1_HVT U449 ( .A1(dummy[20]), .A2(n571), .Y(n1775) );
  NAND2X0_HVT U454 ( .A1(n1885), .A2(n565), .Y(n566) );
  NAND2X0_HVT U455 ( .A1(n1896), .A2(n573), .Y(n567) );
  NAND2X0_HVT U458 ( .A1(n566), .A2(n567), .Y(dummy[26]) );
  INVX1_HVT U459 ( .A(n573), .Y(n565) );
  INVX1_HVT U460 ( .A(n593), .Y(n573) );
  MUX41X1_HVT U462 ( .A1(n2151), .A3(n2159), .A2(n2141), .A4(n2146), .S0(
        keyin[121]), .S1(n965), .Y(dummy[20]) );
  MUX21X2_HVT U463 ( .A1(n2147), .A2(n2150), .S0(n1231), .Y(n2146) );
  MUX21X2_HVT U465 ( .A1(n2560), .A2(n2561), .S0(n844), .Y(n2558) );
  MUX21X1_HVT U466 ( .A1(n1557), .A2(n2258), .S0(n570), .Y(n568) );
  MUX21X1_HVT U467 ( .A1(n2100), .A2(n1550), .S0(n570), .Y(n569) );
  INVX1_HVT U468 ( .A(n2060), .Y(n1550) );
  IBUFFX2_HVT U470 ( .A(n1230), .Y(n570) );
  XOR3X2_HVT U471 ( .A1(n1819), .A2(n599), .A3(n871), .Y(keyout[116]) );
  MUX41X1_HVT U473 ( .A1(n2099), .A3(n2095), .A2(n2101), .A4(n2098), .S0(n594), 
        .S1(n572), .Y(n2094) );
  MUX41X1_HVT U474 ( .A1(n2325), .A3(n2323), .A2(n2331), .A4(n2329), .S0(n1445), .S1(keyin[113]), .Y(n2322) );
  MUX41X1_HVT U475 ( .A1(n2235), .A3(n2253), .A2(n1556), .A4(n1542), .S0(n472), 
        .S1(n1228), .Y(n2209) );
  INVX1_HVT U476 ( .A(n2067), .Y(n1542) );
  MUX41X1_HVT U477 ( .A1(n2195), .A3(n2196), .A2(n2191), .A4(n2192), .S0(n572), 
        .S1(n594), .Y(n2190) );
  MUX41X1_HVT U481 ( .A1(n1508), .A3(n2212), .A2(n2211), .A4(n2213), .S0(n572), 
        .S1(n472), .Y(n2210) );
  INVX1_HVT U482 ( .A(keyin[125]), .Y(n1430) );
  MUX41X1_HVT U483 ( .A1(n2224), .A3(n2220), .A2(n2214), .A4(n2210), .S0(n594), 
        .S1(n856), .Y(dummy[23]) );
  NAND2X0_HVT U486 ( .A1(n2225), .A2(n582), .Y(n574) );
  NAND2X0_HVT U487 ( .A1(n2229), .A2(n1429), .Y(n575) );
  NAND2X0_HVT U491 ( .A1(n574), .A2(n575), .Y(n2224) );
  INVX1_HVT U494 ( .A(n1430), .Y(n1429) );
  XNOR2X1_HVT U495 ( .A1(dummy[20]), .A2(keyin[20]), .Y(n871) );
  MUX21X1_HVT U496 ( .A1(n1624), .A2(n578), .S0(n577), .Y(n576) );
  NAND2X0_HVT U500 ( .A1(n1244), .A2(n1372), .Y(n578) );
  MUX21X1_HVT U502 ( .A1(n23), .A2(n576), .S0(n1239), .Y(n1179) );
  XOR2X1_HVT U505 ( .A1(n1445), .A2(n580), .Y(n579) );
  MUX41X1_HVT U506 ( .A1(n2383), .A3(n2380), .A2(n2384), .A4(n2378), .S0(n581), 
        .S1(n543), .Y(n2377) );
  MUX41X1_HVT U510 ( .A1(n2337), .A3(n2335), .A2(n2336), .A4(n2449), .S0(n581), 
        .S1(n543), .Y(n2334) );
  XNOR2X2_HVT U511 ( .A1(keyin[49]), .A2(n865), .Y(keyout[49]) );
  MUX41X1_HVT U512 ( .A1(n2241), .A3(n2091), .A2(n2232), .A4(n1538), .S0(n583), 
        .S1(n238), .Y(n2090) );
  AO21X1_HVT U513 ( .A1(n1255), .A2(n2621), .A3(n1670), .Y(n2622) );
  MUX21X1_HVT U514 ( .A1(n2699), .A2(n1196), .S0(n554), .Y(n2619) );
  MUX41X1_HVT U516 ( .A1(n1893), .A3(n2013), .A2(n1721), .A4(n2037), .S0(n1480), .S1(n584), .Y(n1892) );
  INVX2_HVT U517 ( .A(keyin[96]), .Y(n1480) );
  IBUFFX2_HVT U518 ( .A(n1768), .Y(keyout[13]) );
  XNOR2X2_HVT U520 ( .A1(dummy[13]), .A2(keyin[13]), .Y(n1768) );
  XOR2X1_HVT U521 ( .A1(dummy[13]), .A2(keyin[13]), .Y(n863) );
  NAND2X0_HVT U522 ( .A1(dummy[5]), .A2(keyin[5]), .Y(n588) );
  NAND2X0_HVT U523 ( .A1(n586), .A2(n587), .Y(n589) );
  NAND2X0_HVT U526 ( .A1(n588), .A2(n589), .Y(n1800) );
  INVX1_HVT U527 ( .A(dummy[5]), .Y(n586) );
  INVX0_HVT U530 ( .A(keyin[5]), .Y(n587) );
  INVX1_HVT U531 ( .A(n1800), .Y(n1626) );
  MUX41X1_HVT U533 ( .A1(n2618), .A3(n2619), .A2(n2617), .A4(n1655), .S0(n1460), .S1(n590), .Y(n2614) );
  XOR3X2_HVT U535 ( .A1(n1793), .A2(n821), .A3(n1763), .Y(keyout[102]) );
  INVX1_HVT U536 ( .A(n1793), .Y(n1486) );
  XNOR2X2_HVT U537 ( .A1(n1805), .A2(keyin[38]), .Y(n1793) );
  IBUFFX2_HVT U538 ( .A(n1461), .Y(n901) );
  MUX21X1_HVT U539 ( .A1(n2193), .A2(n2270), .S0(n1229), .Y(n591) );
  MUX21X1_HVT U540 ( .A1(n1191), .A2(n2194), .S0(n1229), .Y(n592) );
  NAND2X0_HVT U541 ( .A1(n2332), .A2(n896), .Y(n897) );
  NAND2X0_HVT U542 ( .A1(n2543), .A2(n590), .Y(n597) );
  NAND2X0_HVT U543 ( .A1(n2544), .A2(n1252), .Y(n598) );
  NAND2X0_HVT U544 ( .A1(n597), .A2(n598), .Y(n2542) );
  XOR2X1_HVT U545 ( .A1(n1788), .A2(n1835), .Y(keyout[2]) );
  MUX21X1_HVT U546 ( .A1(n1420), .A2(n2545), .S0(n554), .Y(n2544) );
  MUX41X1_HVT U547 ( .A1(n2512), .A3(n2510), .A2(n2511), .A4(n2509), .S0(n595), 
        .S1(n843), .Y(n2508) );
  MUX41X1_HVT U548 ( .A1(n1506), .A3(n2268), .A2(n2251), .A4(n1503), .S0(n238), 
        .S1(n1230), .Y(n2092) );
  MUX41X1_HVT U549 ( .A1(n2389), .A3(n2400), .A2(n2385), .A4(n2394), .S0(n600), 
        .S1(n894), .Y(dummy[13]) );
  NAND2X0_HVT U550 ( .A1(n2636), .A2(n1378), .Y(n603) );
  NAND2X0_HVT U551 ( .A1(n602), .A2(n603), .Y(dummy[6]) );
  IBUFFX2_HVT U552 ( .A(n1378), .Y(n601) );
  XOR2X2_HVT U553 ( .A1(n821), .A2(n1793), .Y(keyout[38]) );
  IBUFFX2_HVT U554 ( .A(n1481), .Y(n1479) );
  XNOR2X1_HVT U555 ( .A1(dummy[6]), .A2(keyin[6]), .Y(n1806) );
  NAND2X0_HVT U556 ( .A1(n2173), .A2(n604), .Y(n605) );
  NAND2X0_HVT U557 ( .A1(n2172), .A2(n582), .Y(n606) );
  NAND2X0_HVT U558 ( .A1(n605), .A2(n606), .Y(n2171) );
  INVX2_HVT U559 ( .A(keyin[118]), .Y(n1441) );
  NAND2X0_HVT U560 ( .A1(n2710), .A2(n590), .Y(n607) );
  NAND2X0_HVT U561 ( .A1(n2570), .A2(n1253), .Y(n608) );
  NAND2X0_HVT U562 ( .A1(n607), .A2(n608), .Y(n2569) );
  NAND2X0_HVT U563 ( .A1(n2530), .A2(n1378), .Y(n633) );
  NAND2X0_HVT U564 ( .A1(n633), .A2(n610), .Y(dummy[1]) );
  IBUFFX2_HVT U565 ( .A(n1378), .Y(n609) );
  MUX41X1_HVT U566 ( .A1(n2137), .A3(n2135), .A2(n2140), .A4(n2138), .S0(n1430), .S1(keyin[121]), .Y(n2134) );
  MUX41X1_HVT U567 ( .A1(n1351), .A3(n1402), .A2(n1530), .A4(n1525), .S0(n283), 
        .S1(n1228), .Y(n2137) );
  INVX2_HVT U568 ( .A(n1783), .Y(keyout[28]) );
  INVX2_HVT U569 ( .A(n1786), .Y(keyout[30]) );
  NAND2X0_HVT U570 ( .A1(n1981), .A2(n573), .Y(n740) );
  NAND2X0_HVT U571 ( .A1(n1971), .A2(n565), .Y(n768) );
  NAND2X0_HVT U572 ( .A1(n740), .A2(n768), .Y(dummy[30]) );
  XOR2X2_HVT U573 ( .A1(dummy[6]), .A2(keyin[6]), .Y(n821) );
  INVX1_HVT U574 ( .A(n822), .Y(n2625) );
  MUX21X1_HVT U575 ( .A1(n823), .A2(n1384), .S0(n1463), .Y(n822) );
  NAND2X0_HVT U576 ( .A1(n830), .A2(n827), .Y(n828) );
  NAND2X0_HVT U577 ( .A1(n824), .A2(n842), .Y(n829) );
  NAND2X0_HVT U578 ( .A1(n828), .A2(n829), .Y(n1155) );
  INVX0_HVT U579 ( .A(n842), .Y(n827) );
  INVX1_HVT U580 ( .A(keyin[19]), .Y(n830) );
  AND2X1_HVT U581 ( .A1(n1156), .A2(n1157), .Y(n842) );
  XNOR2X2_HVT U582 ( .A1(dummy[19]), .A2(keyin[19]), .Y(n1774) );
  MUX21X2_HVT U583 ( .A1(n2640), .A2(n2641), .S0(n844), .Y(n2638) );
  MUX21X1_HVT U584 ( .A1(n1648), .A2(n2699), .S0(n1465), .Y(n2641) );
  IBUFFX2_HVT U585 ( .A(n1778), .Y(keyout[23]) );
  MUX21X1_HVT U586 ( .A1(n2682), .A2(n2681), .S0(n270), .Y(n2570) );
  MUX41X1_HVT U587 ( .A1(n2626), .A3(n2623), .A2(n2624), .A4(n2622), .S0(n843), 
        .S1(n844), .Y(n2620) );
  XOR2X2_HVT U588 ( .A1(n1806), .A2(n1805), .Y(keyout[6]) );
  NAND2X0_HVT U589 ( .A1(n2217), .A2(n572), .Y(n845) );
  NAND2X0_HVT U590 ( .A1(n2215), .A2(n582), .Y(n846) );
  NAND2X0_HVT U591 ( .A1(n845), .A2(n846), .Y(n2214) );
  XOR2X2_HVT U592 ( .A1(n1840), .A2(n1839), .Y(keyout[35]) );
  NAND2X0_HVT U593 ( .A1(n1400), .A2(n847), .Y(n848) );
  NAND2X0_HVT U594 ( .A1(n2161), .A2(n1188), .Y(n849) );
  NAND2X0_HVT U595 ( .A1(n848), .A2(n849), .Y(n2160) );
  INVX0_HVT U596 ( .A(n1188), .Y(n847) );
  MUX21X1_HVT U597 ( .A1(n2376), .A2(n1568), .S0(n1445), .Y(n2375) );
  MUX21X1_HVT U598 ( .A1(n2375), .A2(n2374), .S0(n538), .Y(n2371) );
  NAND2X0_HVT U599 ( .A1(n2072), .A2(n1148), .Y(n850) );
  NAND2X0_HVT U600 ( .A1(n2079), .A2(n1364), .Y(n851) );
  NAND2X0_HVT U601 ( .A1(n850), .A2(n851), .Y(dummy[16]) );
  NAND2X0_HVT U602 ( .A1(n2515), .A2(n853), .Y(n854) );
  NAND2X0_HVT U603 ( .A1(n2508), .A2(n859), .Y(n855) );
  NAND2X0_HVT U604 ( .A1(n854), .A2(n855), .Y(dummy[0]) );
  INVX1_HVT U605 ( .A(n859), .Y(n853) );
  IBUFFX2_HVT U606 ( .A(n1378), .Y(n859) );
  NAND2X0_HVT U607 ( .A1(n2190), .A2(n856), .Y(n857) );
  NAND2X0_HVT U608 ( .A1(n2198), .A2(n1364), .Y(n858) );
  NAND2X0_HVT U609 ( .A1(n857), .A2(n858), .Y(dummy[22]) );
  MUX21X2_HVT U610 ( .A1(n2016), .A2(n1990), .S0(n1341), .Y(n1989) );
  MUX41X1_HVT U611 ( .A1(n2494), .A3(n1617), .A2(n2487), .A4(n1575), .S0(n581), 
        .S1(n543), .Y(n2294) );
  AO21X2_HVT U612 ( .A1(n1458), .A2(n1683), .A3(n1466), .Y(n2616) );
  OA21X2_HVT U613 ( .A1(n1221), .A2(n1466), .A3(n2687), .Y(n2543) );
  OA21X2_HVT U614 ( .A1(n2676), .A2(n1466), .A3(n2559), .Y(n2560) );
  OA21X2_HVT U615 ( .A1(n1633), .A2(n1466), .A3(n2687), .Y(n2566) );
  OA21X2_HVT U616 ( .A1(n2707), .A2(n1466), .A3(n1661), .Y(n2517) );
  XNOR2X1_HVT U617 ( .A1(dummy[30]), .A2(keyin[30]), .Y(n1786) );
  MUX21X1_HVT U618 ( .A1(n2232), .A2(n234), .S0(n1435), .Y(n2130) );
  MUX41X1_HVT U619 ( .A1(n2127), .A3(n2131), .A2(n2128), .A4(n2132), .S0(
        keyin[121]), .S1(keyin[125]), .Y(n2126) );
  IBUFFX2_HVT U620 ( .A(n1155), .Y(n1153) );
  MUX21X1_HVT U621 ( .A1(n2239), .A2(n1548), .S0(n1435), .Y(n2139) );
  INVX1_HVT U622 ( .A(n1445), .Y(n1444) );
  INVX1_HVT U623 ( .A(n2124), .Y(n882) );
  INVX1_HVT U624 ( .A(n1369), .Y(n892) );
  INVX1_HVT U625 ( .A(n1895), .Y(n879) );
  INVX0_HVT U626 ( .A(n1713), .Y(n877) );
  INVX0_HVT U627 ( .A(n881), .Y(n2122) );
  INVX1_HVT U628 ( .A(keyin[109]), .Y(n1461) );
  INVX0_HVT U629 ( .A(n1373), .Y(n872) );
  INVX0_HVT U630 ( .A(n1130), .Y(n895) );
  INVX0_HVT U634 ( .A(n1811), .Y(n1130) );
  INVX0_HVT U635 ( .A(n1461), .Y(n1459) );
  INVX0_HVT U636 ( .A(n1179), .Y(n2331) );
  NAND2X0_HVT U637 ( .A1(n2549), .A2(n590), .Y(n1173) );
  INVX0_HVT U638 ( .A(n1151), .Y(n2150) );
  INVX0_HVT U639 ( .A(n876), .Y(n1894) );
  INVX0_HVT U640 ( .A(n1205), .Y(n878) );
  INVX0_HVT U642 ( .A(n1178), .Y(n1175) );
  NAND2X0_HVT U644 ( .A1(n2103), .A2(n965), .Y(n1083) );
  INVX1_HVT U645 ( .A(keyin[18]), .Y(n870) );
  INVX0_HVT U646 ( .A(n1369), .Y(n893) );
  INVX1_HVT U648 ( .A(n1804), .Y(n1627) );
  NAND2X0_HVT U649 ( .A1(n1960), .A2(keyin[97]), .Y(n890) );
  NAND2X0_HVT U650 ( .A1(n2087), .A2(n1148), .Y(n1126) );
  INVX1_HVT U652 ( .A(n1822), .Y(n868) );
  INVX1_HVT U653 ( .A(n1153), .Y(keyout[19]) );
  INVX1_HVT U654 ( .A(n1431), .Y(n907) );
  INVX0_HVT U655 ( .A(n1231), .Y(n1150) );
  INVX1_HVT U656 ( .A(n1149), .Y(n965) );
  INVX1_HVT U657 ( .A(n1376), .Y(n894) );
  INVX0_HVT U658 ( .A(n1370), .Y(n903) );
  INVX0_HVT U661 ( .A(n1370), .Y(n1184) );
  INVX1_HVT U662 ( .A(n1378), .Y(n1178) );
  INVX1_HVT U663 ( .A(n1771), .Y(n1496) );
  INVX1_HVT U664 ( .A(n1777), .Y(n1492) );
  XNOR2X2_HVT U666 ( .A1(n1768), .A2(n1812), .Y(keyout[77]) );
  INVX1_HVT U667 ( .A(n1399), .Y(n1163) );
  INVX1_HVT U668 ( .A(keyin[103]), .Y(n884) );
  XNOR2X1_HVT U669 ( .A1(keyin[40]), .A2(n861), .Y(keyout[40]) );
  IBUFFX2_HVT U670 ( .A(n1772), .Y(keyout[17]) );
  INVX1_HVT U671 ( .A(n1772), .Y(n1495) );
  XOR2X2_HVT U672 ( .A1(dummy[30]), .A2(keyin[30]), .Y(n867) );
  INVX0_HVT U673 ( .A(n1773), .Y(keyout[18]) );
  XOR2X1_HVT U674 ( .A1(dummy[18]), .A2(n870), .Y(n1773) );
  XOR3X2_HVT U675 ( .A1(n1821), .A2(n1441), .A3(n1777), .Y(keyout[118]) );
  XOR3X2_HVT U677 ( .A1(n1815), .A2(n543), .A3(n1771), .Y(keyout[112]) );
  XNOR2X2_HVT U679 ( .A1(keyin[50]), .A2(n869), .Y(keyout[50]) );
  XOR3X2_HVT U680 ( .A1(n868), .A2(n896), .A3(n1778), .Y(keyout[119]) );
  XOR2X1_HVT U683 ( .A1(dummy[18]), .A2(n870), .Y(n869) );
  MUX41X1_HVT U684 ( .A1(n1697), .A3(n2055), .A2(n1201), .A4(n1947), .S0(n584), 
        .S1(n1481), .Y(n1903) );
  MUX41X1_HVT U686 ( .A1(n1904), .A3(n1899), .A2(n1903), .A4(n1897), .S0(n884), 
        .S1(n564), .Y(n1896) );
  INVX2_HVT U689 ( .A(n1781), .Y(keyout[26]) );
  XNOR2X2_HVT U690 ( .A1(keyin[55]), .A2(n1778), .Y(keyout[55]) );
  INVX0_HVT U692 ( .A(n1777), .Y(keyout[22]) );
  INVX0_HVT U693 ( .A(n1771), .Y(keyout[16]) );
  XOR2X1_HVT U694 ( .A1(keyin[62]), .A2(n867), .Y(keyout[62]) );
  XOR3X1_HVT U695 ( .A1(n1818), .A2(n872), .A3(n1774), .Y(keyout[115]) );
  NBUFFX2_HVT U696 ( .A(keyin[112]), .Y(n873) );
  MUX21X1_HVT U698 ( .A1(n2388), .A2(n2386), .S0(n1445), .Y(n2385) );
  XNOR2X2_HVT U699 ( .A1(n871), .A2(n1819), .Y(keyout[84]) );
  XNOR3X1_HVT U700 ( .A1(n1820), .A2(n1443), .A3(n1776), .Y(keyout[117]) );
  XOR2X2_HVT U702 ( .A1(n1492), .A2(n1821), .Y(keyout[86]) );
  XOR2X2_HVT U703 ( .A1(n1496), .A2(n1815), .Y(keyout[80]) );
  MUX41X1_HVT U704 ( .A1(n2304), .A3(n2302), .A2(n2303), .A4(n2299), .S0(n894), 
        .S1(n1445), .Y(n2298) );
  XNOR2X2_HVT U705 ( .A1(n852), .A2(keyin[12]), .Y(n875) );
  MUX41X1_HVT U710 ( .A1(n879), .A3(n878), .A2(n880), .A4(n877), .S0(n584), 
        .S1(n1481), .Y(n876) );
  NAND2X0_HVT U712 ( .A1(n254), .A2(n1986), .Y(n880) );
  XNOR2X2_HVT U713 ( .A1(n1779), .A2(n1823), .Y(keyout[88]) );
  IBUFFX2_HVT U714 ( .A(n1779), .Y(keyout[24]) );
  XNOR2X2_HVT U715 ( .A1(n1787), .A2(n1830), .Y(keyout[95]) );
  IBUFFX2_HVT U716 ( .A(n1787), .Y(keyout[31]) );
  MUX21X1_HVT U717 ( .A1(n1401), .A2(n2164), .S0(n1162), .Y(n2124) );
  MUX21X1_HVT U718 ( .A1(n883), .A2(n882), .S0(n1150), .Y(n881) );
  OAI21X1_HVT U720 ( .A1(n2238), .A2(n1435), .A3(n2123), .Y(n883) );
  MUX41X1_HVT U721 ( .A1(n2399), .A3(n2398), .A2(n1592), .A4(n2397), .S0(n1445), .S1(n581), .Y(n2394) );
  XNOR2X1_HVT U722 ( .A1(n1475), .A2(n1481), .Y(n1185) );
  XNOR2X1_HVT U724 ( .A1(keyin[61]), .A2(n1784), .Y(keyout[61]) );
  XNOR2X2_HVT U725 ( .A1(n1783), .A2(n1827), .Y(keyout[92]) );
  MUX41X1_HVT U726 ( .A1(n1958), .A3(n1954), .A2(n1953), .A4(n1951), .S0(n564), 
        .S1(n884), .Y(n1950) );
  XOR3X2_HVT U727 ( .A1(n1479), .A2(n1831), .A3(n1832), .Y(keyout[96]) );
  XNOR2X2_HVT U729 ( .A1(keyin[56]), .A2(n1779), .Y(keyout[56]) );
  XNOR2X2_HVT U731 ( .A1(n1780), .A2(n1824), .Y(keyout[89]) );
  IBUFFX2_HVT U733 ( .A(n1780), .Y(keyout[25]) );
  XNOR2X2_HVT U734 ( .A1(keyin[63]), .A2(n1787), .Y(keyout[63]) );
  XNOR2X2_HVT U735 ( .A1(n1782), .A2(n1826), .Y(keyout[91]) );
  IBUFFX2_HVT U738 ( .A(n1782), .Y(keyout[27]) );
  MUX21X2_HVT U739 ( .A1(n1916), .A2(n1908), .S0(n565), .Y(dummy[27]) );
  XNOR2X2_HVT U740 ( .A1(keyin[57]), .A2(n1780), .Y(keyout[57]) );
  MUX41X1_HVT U742 ( .A1(n2262), .A3(n1546), .A2(n2240), .A4(n2102), .S0(n1162), .S1(n907), .Y(n2101) );
  INVX1_HVT U743 ( .A(n1434), .Y(n1162) );
  XNOR2X2_HVT U745 ( .A1(keyin[59]), .A2(n1782), .Y(keyout[59]) );
  XNOR2X1_HVT U747 ( .A1(keyin[58]), .A2(n1781), .Y(keyout[58]) );
  NAND2X0_HVT U748 ( .A1(n2152), .A2(n1150), .Y(n885) );
  NAND2X0_HVT U749 ( .A1(n2153), .A2(n1231), .Y(n886) );
  NAND2X0_HVT U750 ( .A1(n886), .A2(n885), .Y(n2151) );
  NAND2X0_HVT U752 ( .A1(n1959), .A2(n887), .Y(n888) );
  NAND2X0_HVT U753 ( .A1(n1201), .A2(n1185), .Y(n889) );
  NAND2X0_HVT U754 ( .A1(n888), .A2(n889), .Y(n1958) );
  INVX0_HVT U756 ( .A(n1185), .Y(n887) );
  NAND2X0_HVT U757 ( .A1(n1950), .A2(n593), .Y(n891) );
  NAND2X0_HVT U759 ( .A1(n890), .A2(n891), .Y(dummy[29]) );
  MUX21X1_HVT U761 ( .A1(n1375), .A2(n1372), .S0(n1445), .Y(n2379) );
  XNOR2X1_HVT U762 ( .A1(keyin[47]), .A2(n1770), .Y(keyout[47]) );
  IBUFFX2_HVT U763 ( .A(n1770), .Y(keyout[15]) );
  OA21X2_HVT U766 ( .A1(n1596), .A2(n1445), .A3(n1580), .Y(n2383) );
  MUX21X1_HVT U767 ( .A1(n2438), .A2(n2440), .S0(n1443), .Y(n2437) );
  XNOR2X2_HVT U768 ( .A1(n1767), .A2(n895), .Y(keyout[76]) );
  XNOR2X2_HVT U771 ( .A1(keyin[44]), .A2(n875), .Y(keyout[44]) );
  NAND2X0_HVT U772 ( .A1(n2322), .A2(n1184), .Y(n898) );
  NAND2X0_HVT U773 ( .A1(n897), .A2(n898), .Y(dummy[10]) );
  INVX1_HVT U775 ( .A(n1184), .Y(n896) );
  XNOR2X2_HVT U776 ( .A1(n1766), .A2(n1810), .Y(keyout[75]) );
  IBUFFX2_HVT U778 ( .A(n1766), .Y(keyout[11]) );
  XNOR2X2_HVT U779 ( .A1(n1769), .A2(n1813), .Y(keyout[78]) );
  NAND2X0_HVT U780 ( .A1(n2291), .A2(n903), .Y(n899) );
  NAND2X0_HVT U781 ( .A1(n2298), .A2(n1370), .Y(n900) );
  NAND2X0_HVT U783 ( .A1(n899), .A2(n900), .Y(dummy[8]) );
  XNOR2X2_HVT U788 ( .A1(n1797), .A2(n1808), .Y(keyout[73]) );
  IBUFFX2_HVT U789 ( .A(n1797), .Y(keyout[9]) );
  XNOR2X2_HVT U790 ( .A1(n1770), .A2(n1814), .Y(keyout[79]) );
  IBUFFX2_HVT U794 ( .A(n1461), .Y(n902) );
  OA21X2_HVT U795 ( .A1(n1659), .A2(n1461), .A3(n1643), .Y(n2603) );
  IBUFFX2_HVT U796 ( .A(n1461), .Y(n1460) );
  XNOR2X2_HVT U800 ( .A1(keyin[43]), .A2(n1766), .Y(keyout[43]) );
  XNOR2X2_HVT U803 ( .A1(keyin[46]), .A2(n1769), .Y(keyout[46]) );
  XNOR2X2_HVT U804 ( .A1(keyin[41]), .A2(n1797), .Y(keyout[41]) );
  NAND2X0_HVT U805 ( .A1(n1417), .A2(n904), .Y(n905) );
  NAND2X0_HVT U806 ( .A1(n2599), .A2(n1189), .Y(n906) );
  NAND2X0_HVT U807 ( .A1(n906), .A2(n905), .Y(n2598) );
  INVX0_HVT U808 ( .A(n1189), .Y(n904) );
  MUX41X1_HVT U809 ( .A1(n1501), .A3(n1533), .A2(n1366), .A4(n2193), .S0(n1162), .S1(n907), .Y(n2098) );
  NAND2X0_HVT U810 ( .A1(n2129), .A2(n908), .Y(n909) );
  NAND2X0_HVT U811 ( .A1(n2130), .A2(n907), .Y(n910) );
  NAND2X0_HVT U812 ( .A1(n909), .A2(n910), .Y(n2128) );
  INVX0_HVT U813 ( .A(n1150), .Y(n908) );
  XOR2X2_HVT U814 ( .A1(n525), .A2(n1807), .Y(keyout[72]) );
  NAND2X0_HVT U815 ( .A1(n1524), .A2(n908), .Y(n911) );
  NAND2X0_HVT U817 ( .A1(n2139), .A2(n1150), .Y(n912) );
  NAND2X0_HVT U818 ( .A1(n2168), .A2(n582), .Y(n913) );
  NAND2X0_HVT U819 ( .A1(n2170), .A2(n1429), .Y(n914) );
  NAND2X0_HVT U821 ( .A1(n913), .A2(n914), .Y(n2167) );
  XNOR2X2_HVT U822 ( .A1(n1774), .A2(n1818), .Y(keyout[83]) );
  XNOR2X1_HVT U823 ( .A1(n1778), .A2(n1822), .Y(keyout[87]) );
  MUX41X1_HVT U824 ( .A1(n2219), .A3(n2267), .A2(n1541), .A4(n1513), .S0(n283), 
        .S1(n907), .Y(n2217) );
  NAND2X0_HVT U825 ( .A1(n2221), .A2(n582), .Y(n938) );
  NAND2X0_HVT U826 ( .A1(n2223), .A2(n1429), .Y(n963) );
  NAND2X0_HVT U827 ( .A1(n938), .A2(n963), .Y(n2220) );
  NAND2X0_HVT U829 ( .A1(n2116), .A2(n1149), .Y(n1125) );
  NAND2X0_HVT U833 ( .A1(n1083), .A2(n1125), .Y(dummy[18]) );
  INVX1_HVT U834 ( .A(n1148), .Y(n1149) );
  NAND2X0_HVT U835 ( .A1(n2094), .A2(n1364), .Y(n1127) );
  NAND2X0_HVT U836 ( .A1(n1127), .A2(n1126), .Y(dummy[17]) );
  XOR2X2_HVT U839 ( .A1(n1495), .A2(n1816), .Y(keyout[81]) );
  NAND2X0_HVT U840 ( .A1(n1409), .A2(n579), .Y(n1131) );
  NAND2X0_HVT U843 ( .A1(n2379), .A2(n1187), .Y(n1132) );
  NAND2X0_HVT U844 ( .A1(n1132), .A2(n1131), .Y(n2378) );
  IBUFFX2_HVT U846 ( .A(n1475), .Y(n1133) );
  INVX2_HVT U848 ( .A(n1475), .Y(n1473) );
  NAND2X0_HVT U849 ( .A1(n1391), .A2(n1134), .Y(n1146) );
  NAND2X0_HVT U850 ( .A1(n1944), .A2(n1186), .Y(n1147) );
  NAND2X0_HVT U851 ( .A1(n1146), .A2(n1147), .Y(n1943) );
  INVX0_HVT U852 ( .A(n1186), .Y(n1134) );
  MUX41X1_HVT U853 ( .A1(n1514), .A3(n1535), .A2(n1505), .A4(n2222), .S0(n1162), .S1(n1150), .Y(n2221) );
  OA21X2_HVT U854 ( .A1(n1502), .A2(n1435), .A3(n2249), .Y(n2129) );
  OA21X2_HVT U855 ( .A1(n1219), .A2(n1435), .A3(n2249), .Y(n2107) );
  AO21X2_HVT U856 ( .A1(n1428), .A2(n1552), .A3(n1435), .Y(n2178) );
  MUX41X1_HVT U857 ( .A1(n1522), .A3(n2254), .A2(n1152), .A4(n1535), .S0(n1430), .S1(n1162), .Y(n1151) );
  NAND2X0_HVT U858 ( .A1(n1424), .A2(n1351), .Y(n1152) );
  INVX1_HVT U859 ( .A(n2249), .Y(n1522) );
  OA21X2_HVT U860 ( .A1(n2246), .A2(n1435), .A3(n1518), .Y(n2096) );
  MUX21X1_HVT U861 ( .A1(n2157), .A2(n2156), .S0(n283), .Y(n2153) );
  NAND2X0_HVT U862 ( .A1(n2126), .A2(n1148), .Y(n1156) );
  NAND2X0_HVT U863 ( .A1(n2134), .A2(n1364), .Y(n1157) );
  NAND2X0_HVT U864 ( .A1(n1156), .A2(n1157), .Y(dummy[19]) );
  XOR2X2_HVT U865 ( .A1(n1155), .A2(keyin[51]), .Y(keyout[51]) );
  XOR2X2_HVT U866 ( .A1(n1835), .A2(n1164), .Y(keyout[66]) );
  NAND2X0_HVT U867 ( .A1(n2663), .A2(n1461), .Y(n1158) );
  NAND2X0_HVT U868 ( .A1(n2667), .A2(n901), .Y(n1159) );
  NAND2X0_HVT U869 ( .A1(n1158), .A2(n1159), .Y(n2662) );
  MUX21X1_HVT U870 ( .A1(n2665), .A2(n2666), .S0(n1255), .Y(n2663) );
  NAND2X0_HVT U871 ( .A1(n2563), .A2(n1178), .Y(n1160) );
  NAND2X0_HVT U872 ( .A1(n2571), .A2(n1378), .Y(n1161) );
  NAND2X0_HVT U873 ( .A1(n1160), .A2(n1161), .Y(dummy[3]) );
  MUX21X2_HVT U874 ( .A1(n2566), .A2(n2567), .S0(n590), .Y(n2565) );
  INVX0_HVT U875 ( .A(n1216), .Y(n1169) );
  XOR2X2_HVT U876 ( .A1(n289), .A2(n1799), .Y(keyout[5]) );
  OR2X1_HVT U877 ( .A1(n1163), .A2(n1215), .Y(n1182) );
  XOR2X1_HVT U878 ( .A1(n1836), .A2(keyin[66]), .Y(n1164) );
  NAND2X0_HVT U879 ( .A1(n2551), .A2(n1169), .Y(n1165) );
  NAND2X0_HVT U880 ( .A1(n1417), .A2(n1216), .Y(n1166) );
  NAND2X0_HVT U881 ( .A1(n1165), .A2(n1166), .Y(n2550) );
  NAND2X0_HVT U882 ( .A1(n1416), .A2(n1169), .Y(n1170) );
  NAND2X0_HVT U883 ( .A1(n1216), .A2(n2625), .Y(n1171) );
  NAND2X0_HVT U884 ( .A1(n1170), .A2(n1171), .Y(n2624) );
  XNOR2X2_HVT U885 ( .A1(n1773), .A2(n1817), .Y(keyout[82]) );
  NAND2X0_HVT U886 ( .A1(n2550), .A2(n1253), .Y(n1174) );
  NAND2X0_HVT U887 ( .A1(n1173), .A2(n1174), .Y(n2548) );
  NAND2X0_HVT U888 ( .A1(n2539), .A2(n1178), .Y(n1177) );
  NAND2X0_HVT U889 ( .A1(n1176), .A2(n1177), .Y(dummy[2]) );
  XNOR2X2_HVT U890 ( .A1(n218), .A2(n1162), .Y(n1215) );
  MUX21X2_HVT U891 ( .A1(n2115), .A2(n1400), .S0(n1215), .Y(n2114) );
  AO21X2_HVT U892 ( .A1(n1442), .A2(n1619), .A3(n280), .Y(n2396) );
  OA21X2_HVT U893 ( .A1(n2463), .A2(n280), .A3(n1586), .Y(n2315) );
  NAND2X0_HVT U894 ( .A1(n1408), .A2(n577), .Y(n1180) );
  NAND2X0_HVT U895 ( .A1(n295), .A2(n1214), .Y(n1181) );
  NAND2X0_HVT U896 ( .A1(n1180), .A2(n1181), .Y(n2404) );
  NAND2X0_HVT U897 ( .A1(n2187), .A2(n1215), .Y(n1183) );
  NAND2X0_HVT U898 ( .A1(n1183), .A2(n1182), .Y(n2186) );
  MUX21X2_HVT U899 ( .A1(n2113), .A2(n2114), .S0(n1232), .Y(n2112) );
  MUX21X1_HVT U900 ( .A1(n1859), .A2(n1860), .S0(n1342), .Y(n1858) );
  MUX21X1_HVT U901 ( .A1(n2442), .A2(n2446), .S0(n1443), .Y(n2441) );
  MUX21X1_HVT U902 ( .A1(n1588), .A2(n2465), .S0(n1444), .Y(n2362) );
  MUX21X1_HVT U903 ( .A1(n1520), .A2(n2248), .S0(n1429), .Y(n2145) );
  MUX21X1_HVT U904 ( .A1(n1567), .A2(n1594), .S0(n1444), .Y(n2366) );
  MUX21X1_HVT U905 ( .A1(n1209), .A2(n1583), .S0(n1444), .Y(n2360) );
  MUX21X1_HVT U906 ( .A1(n1210), .A2(n1515), .S0(n1429), .Y(n2143) );
  MUX21X2_HVT U907 ( .A1(n2653), .A2(n2655), .S0(n901), .Y(n2652) );
  MUX21X2_HVT U908 ( .A1(n2606), .A2(n2608), .S0(n901), .Y(n2605) );
  MUX21X2_HVT U909 ( .A1(n2006), .A2(n2010), .S0(n1341), .Y(n2005) );
  MUX21X2_HVT U910 ( .A1(n2008), .A2(n2009), .S0(n1348), .Y(n2006) );
  XOR2X2_HVT U911 ( .A1(n1758), .A2(keyin[100]), .Y(n2033) );
  INVX0_HVT U912 ( .A(n1471), .Y(n1470) );
  XOR2X1_HVT U913 ( .A1(n1798), .A2(keyin[36]), .Y(n1803) );
  XOR2X1_HVT U914 ( .A1(keyin[40]), .A2(keyin[72]), .Y(n1807) );
  XOR2X1_HVT U915 ( .A1(keyin[41]), .A2(keyin[73]), .Y(n1808) );
  XOR2X1_HVT U916 ( .A1(keyin[42]), .A2(keyin[74]), .Y(n1809) );
  XOR2X1_HVT U917 ( .A1(keyin[43]), .A2(keyin[75]), .Y(n1810) );
  XOR2X1_HVT U918 ( .A1(keyin[44]), .A2(keyin[76]), .Y(n1811) );
  XOR2X1_HVT U919 ( .A1(keyin[45]), .A2(keyin[77]), .Y(n1812) );
  XOR2X1_HVT U920 ( .A1(keyin[46]), .A2(keyin[78]), .Y(n1813) );
  XOR2X1_HVT U921 ( .A1(keyin[47]), .A2(keyin[79]), .Y(n1814) );
  XOR2X1_HVT U922 ( .A1(keyin[48]), .A2(keyin[80]), .Y(n1815) );
  XOR2X1_HVT U923 ( .A1(keyin[49]), .A2(keyin[81]), .Y(n1816) );
  XOR2X1_HVT U924 ( .A1(keyin[50]), .A2(keyin[82]), .Y(n1817) );
  XOR2X1_HVT U925 ( .A1(keyin[51]), .A2(keyin[83]), .Y(n1818) );
  XOR2X1_HVT U926 ( .A1(keyin[52]), .A2(keyin[84]), .Y(n1819) );
  XOR2X1_HVT U927 ( .A1(keyin[53]), .A2(keyin[85]), .Y(n1820) );
  XOR2X1_HVT U928 ( .A1(keyin[54]), .A2(keyin[86]), .Y(n1821) );
  XOR2X1_HVT U929 ( .A1(keyin[55]), .A2(keyin[87]), .Y(n1822) );
  XOR2X1_HVT U930 ( .A1(keyin[56]), .A2(keyin[88]), .Y(n1823) );
  XOR2X1_HVT U931 ( .A1(keyin[57]), .A2(keyin[89]), .Y(n1824) );
  XOR2X1_HVT U932 ( .A1(keyin[58]), .A2(keyin[90]), .Y(n1825) );
  XOR2X1_HVT U933 ( .A1(keyin[62]), .A2(keyin[94]), .Y(n1829) );
  XNOR2X1_HVT U934 ( .A1(n1473), .A2(n291), .Y(n1186) );
  XNOR2X1_HVT U935 ( .A1(n604), .A2(n1424), .Y(n1188) );
  XNOR2X1_HVT U936 ( .A1(n1459), .A2(n1453), .Y(n1189) );
  XOR2X2_HVT U937 ( .A1(keyin[60]), .A2(keyout[28]), .Y(keyout[60]) );
  XOR2X2_HVT U938 ( .A1(n1788), .A2(keyin[34]), .Y(n1836) );
  XOR3X2_HVT U939 ( .A1(keyin[65]), .A2(keyin[33]), .A3(n1802), .Y(n1833) );
  XOR2X2_HVT U940 ( .A1(keyin[60]), .A2(keyin[92]), .Y(n1827) );
  XOR2X2_HVT U941 ( .A1(keyin[61]), .A2(keyin[93]), .Y(n1828) );
  XOR2X2_HVT U946 ( .A1(keyin[63]), .A2(keyin[95]), .Y(n1830) );
  XOR2X2_HVT U947 ( .A1(keyin[59]), .A2(keyin[91]), .Y(n1826) );
  INVX1_HVT U948 ( .A(n2051), .Y(n1753) );
  INVX1_HVT U949 ( .A(n2488), .Y(n1621) );
  INVX1_HVT U950 ( .A(n2271), .Y(n1554) );
  INVX1_HVT U951 ( .A(n2709), .Y(n1685) );
  NBUFFX2_HVT U953 ( .A(n2051), .Y(n1392) );
  NBUFFX2_HVT U955 ( .A(n2051), .Y(n1393) );
  AND2X1_HVT U956 ( .A1(n1409), .A2(n2423), .Y(n1190) );
  AND2X1_HVT U957 ( .A1(n1400), .A2(n2206), .Y(n1191) );
  MUX21X1_HVT U958 ( .A1(n1192), .A2(n1590), .S0(n873), .Y(n2398) );
  MUX21X1_HVT U959 ( .A1(n1193), .A2(n1522), .S0(n1233), .Y(n2180) );
  MUX21X1_HVT U961 ( .A1(n2478), .A2(n1192), .S0(n1244), .Y(n2399) );
  AND2X1_HVT U962 ( .A1(n1413), .A2(n2381), .Y(n1192) );
  AND2X1_HVT U964 ( .A1(n1405), .A2(n2163), .Y(n1193) );
  AND2X1_HVT U965 ( .A1(n1356), .A2(n2435), .Y(n1194) );
  AND2X1_HVT U966 ( .A1(n1553), .A2(n2218), .Y(n1195) );
  AND2X1_HVT U967 ( .A1(n1421), .A2(n2601), .Y(n1196) );
  MUX21X1_HVT U968 ( .A1(n1722), .A2(n1922), .S0(n1339), .Y(n1921) );
  MUX21X1_HVT U969 ( .A1(n1747), .A2(n1395), .S0(n1349), .Y(n1922) );
  AND2X1_HVT U970 ( .A1(n1684), .A2(n2656), .Y(n1197) );
  AND2X1_HVT U972 ( .A1(n1417), .A2(n2644), .Y(n1198) );
  MUX21X1_HVT U973 ( .A1(n1708), .A2(n1752), .S0(n1347), .Y(n1992) );
  AND2X1_HVT U974 ( .A1(n2003), .A2(n1757), .Y(n1199) );
  AND2X1_HVT U975 ( .A1(n1390), .A2(n1986), .Y(n1200) );
  AND2X1_HVT U976 ( .A1(n1396), .A2(n1946), .Y(n1201) );
  NBUFFX2_HVT U978 ( .A(n2488), .Y(n1406) );
  NBUFFX2_HVT U979 ( .A(n2271), .Y(n1397) );
  NBUFFX2_HVT U980 ( .A(n253), .Y(n1361) );
  NBUFFX2_HVT U981 ( .A(n1620), .Y(n1354) );
  NBUFFX2_HVT U982 ( .A(n1553), .Y(n1351) );
  NBUFFX2_HVT U983 ( .A(n1620), .Y(n1355) );
  NBUFFX2_HVT U984 ( .A(n1553), .Y(n1352) );
  NBUFFX2_HVT U985 ( .A(n1620), .Y(n1356) );
  INVX1_HVT U986 ( .A(n1411), .Y(n1619) );
  INVX1_HVT U987 ( .A(n1402), .Y(n1552) );
  NBUFFX2_HVT U988 ( .A(n2709), .Y(n1414) );
  INVX1_HVT U989 ( .A(n1394), .Y(n1752) );
  INVX1_HVT U991 ( .A(n2494), .Y(n1623) );
  INVX1_HVT U993 ( .A(n2277), .Y(n1556) );
  NAND2X0_HVT U994 ( .A1(n1362), .A2(n1754), .Y(n2051) );
  NBUFFX2_HVT U999 ( .A(n2488), .Y(n1407) );
  NBUFFX2_HVT U1003 ( .A(n2271), .Y(n1398) );
  INVX1_HVT U1004 ( .A(n2058), .Y(n1755) );
  NBUFFX2_HVT U1006 ( .A(n2709), .Y(n1415) );
  INVX1_HVT U1009 ( .A(n2714), .Y(n1683) );
  INVX1_HVT U1010 ( .A(n2715), .Y(n1687) );
  MUX21X1_HVT U1011 ( .A1(n1351), .A2(n1531), .S0(n1233), .Y(n2113) );
  MUX21X1_HVT U1015 ( .A1(n2449), .A2(n1607), .S0(n1244), .Y(n2403) );
  MUX21X1_HVT U1018 ( .A1(n2490), .A2(n2406), .S0(n873), .Y(n2405) );
  MUX21X1_HVT U1020 ( .A1(n2232), .A2(n1540), .S0(n1234), .Y(n2185) );
  MUX21X1_HVT U1027 ( .A1(n2273), .A2(n2189), .S0(n1233), .Y(n2188) );
  MUX21X1_HVT U1028 ( .A1(n2356), .A2(n1592), .S0(n1242), .Y(n2355) );
  MUX21X1_HVT U1030 ( .A1(n1615), .A2(n2456), .S0(n1244), .Y(n2356) );
  MUX21X1_HVT U1031 ( .A1(n2364), .A2(n2367), .S0(n1241), .Y(n2363) );
  MUX21X1_HVT U1033 ( .A1(n2365), .A2(n2366), .S0(n1243), .Y(n2364) );
  MUX21X1_HVT U1034 ( .A1(n2148), .A2(n2149), .S0(n1434), .Y(n2147) );
  MUX21X1_HVT U1035 ( .A1(n243), .A2(n1662), .S0(n270), .Y(n2549) );
  MUX21X1_HVT U1037 ( .A1(n2444), .A2(n2445), .S0(n1243), .Y(n2442) );
  MUX21X1_HVT U1038 ( .A1(n2227), .A2(n2228), .S0(n1434), .Y(n2225) );
  MUX21X1_HVT U1039 ( .A1(n2432), .A2(n2434), .S0(n247), .Y(n2431) );
  MUX21X1_HVT U1041 ( .A1(n2670), .A2(n1671), .S0(n1463), .Y(n2623) );
  MUX21X1_HVT U1043 ( .A1(n2711), .A2(n2627), .S0(n1255), .Y(n2626) );
  XOR2X1_HVT U1044 ( .A1(n1437), .A2(n1619), .Y(n2450) );
  XOR2X1_HVT U1045 ( .A1(n1425), .A2(n1552), .Y(n2233) );
  MUX21X1_HVT U1046 ( .A1(n1679), .A2(n2677), .S0(n542), .Y(n2576) );
  MUX21X1_HVT U1047 ( .A1(n2585), .A2(n2586), .S0(n1255), .Y(n2584) );
  XOR2X1_HVT U1050 ( .A1(n217), .A2(n1683), .Y(n2671) );
  MUX21X1_HVT U1051 ( .A1(n1723), .A2(n2044), .S0(n1342), .Y(n1959) );
  MUX21X1_HVT U1052 ( .A1(n1625), .A2(n599), .S0(n1437), .Y(n2376) );
  MUX21X1_HVT U1056 ( .A1(n1500), .A2(n2158), .S0(n604), .Y(n2157) );
  MUX21X1_HVT U1058 ( .A1(n1557), .A2(n1353), .S0(n1426), .Y(n2158) );
  MUX21X1_HVT U1060 ( .A1(n1752), .A2(n1756), .S0(n1470), .Y(n1893) );
  MUX21X1_HVT U1061 ( .A1(n1753), .A2(n1756), .S0(n1468), .Y(n1884) );
  MUX21X1_HVT U1063 ( .A1(n1360), .A2(n1396), .S0(n1470), .Y(n1871) );
  MUX21X1_HVT U1066 ( .A1(n2058), .A2(n1390), .S0(n290), .Y(n1872) );
  MUX21X1_HVT U1068 ( .A1(n254), .A2(n1363), .S0(n558), .Y(n1983) );
  MUX21X1_HVT U1069 ( .A1(n1755), .A2(n1757), .S0(n1469), .Y(n1895) );
  XOR2X1_HVT U1072 ( .A1(n1391), .A2(n1469), .Y(n2011) );
  MUX21X1_HVT U1073 ( .A1(n1360), .A2(n1363), .S0(n291), .Y(n1868) );
  MUX21X1_HVT U1076 ( .A1(n1631), .A2(n2596), .S0(n1459), .Y(n2595) );
  MUX21X1_HVT U1077 ( .A1(n1689), .A2(n1358), .S0(n1456), .Y(n2596) );
  MUX21X1_HVT U1082 ( .A1(n1619), .A2(n1624), .S0(n1437), .Y(n2335) );
  MUX21X1_HVT U1084 ( .A1(n1623), .A2(n1355), .S0(n1440), .Y(n2337) );
  MUX21X1_HVT U1088 ( .A1(n1552), .A2(n1163), .S0(n1423), .Y(n2119) );
  MUX21X1_HVT U1089 ( .A1(n1556), .A2(n1352), .S0(n1423), .Y(n2121) );
  MUX21X1_HVT U1091 ( .A1(n2494), .A2(n1410), .S0(n1436), .Y(n2310) );
  MUX21X1_HVT U1092 ( .A1(n2277), .A2(n1401), .S0(n1424), .Y(n2091) );
  MUX21X1_HVT U1094 ( .A1(n2465), .A2(n2289), .S0(n873), .Y(n2283) );
  MUX21X1_HVT U1095 ( .A1(n2248), .A2(n2070), .S0(n1233), .Y(n2064) );
  MUX21X1_HVT U1096 ( .A1(n1595), .A2(n2491), .S0(n1444), .Y(n2384) );
  MUX21X1_HVT U1099 ( .A1(n1527), .A2(n2274), .S0(n1429), .Y(n2166) );
  MUX21X1_HVT U1100 ( .A1(n2420), .A2(n2419), .S0(n1242), .Y(n2417) );
  MUX21X1_HVT U1101 ( .A1(n1517), .A2(n2261), .S0(n1233), .Y(n2203) );
  MUX21X1_HVT U1102 ( .A1(n2477), .A2(n2393), .S0(n1242), .Y(n2392) );
  MUX21X1_HVT U1103 ( .A1(n1355), .A2(n1621), .S0(n1438), .Y(n2393) );
  MUX21X1_HVT U1104 ( .A1(n1203), .A2(n2174), .S0(n1233), .Y(n2173) );
  MUX21X1_HVT U1108 ( .A1(n2260), .A2(n2175), .S0(n1232), .Y(n2174) );
  MUX21X1_HVT U1110 ( .A1(n1352), .A2(n1554), .S0(n1422), .Y(n2175) );
  XOR2X1_HVT U1112 ( .A1(n1408), .A2(n1440), .Y(n2447) );
  XOR2X1_HVT U1114 ( .A1(n1399), .A2(n1426), .Y(n2230) );
  MUX21X1_HVT U1122 ( .A1(n599), .A2(n1413), .S0(n1436), .Y(n2308) );
  MUX21X1_HVT U1124 ( .A1(n1353), .A2(n1405), .S0(n1422), .Y(n2089) );
  AND2X1_HVT U1126 ( .A1(n1440), .A2(n1624), .Y(n1202) );
  AND2X1_HVT U1127 ( .A1(n1426), .A2(n1163), .Y(n1203) );
  MUX21X1_HVT U1131 ( .A1(n1756), .A2(n1755), .S0(n559), .Y(n2032) );
  MUX21X1_HVT U1135 ( .A1(n1391), .A2(n1395), .S0(n559), .Y(n2044) );
  MUX21X1_HVT U1137 ( .A1(n1757), .A2(n1360), .S0(n291), .Y(n2042) );
  MUX21X1_HVT U1139 ( .A1(n2077), .A2(n2078), .S0(n1231), .Y(n2076) );
  MUX21X1_HVT U1141 ( .A1(n1980), .A2(n1979), .S0(n1343), .Y(n1977) );
  MUX21X1_HVT U1148 ( .A1(n2038), .A2(n1395), .S0(n1349), .Y(n1980) );
  MUX21X1_HVT U1149 ( .A1(n2466), .A2(n2382), .S0(n1444), .Y(n2380) );
  MUX21X1_HVT U1151 ( .A1(n2249), .A2(n2164), .S0(n1429), .Y(n2162) );
  MUX21X1_HVT U1155 ( .A1(n1413), .A2(n1412), .S0(n562), .Y(n2466) );
  MUX21X1_HVT U1157 ( .A1(n2277), .A2(n1403), .S0(n1424), .Y(n2249) );
  MUX21X1_HVT U1158 ( .A1(n1755), .A2(n1753), .S0(n291), .Y(n2022) );
  MUX21X1_HVT U1160 ( .A1(n1755), .A2(n1360), .S0(n557), .Y(n2025) );
  MUX21X1_HVT U1161 ( .A1(n254), .A2(n1756), .S0(n558), .Y(n2034) );
  MUX21X1_HVT U1162 ( .A1(n1390), .A2(n1360), .S0(n558), .Y(n2039) );
  MUX21X1_HVT U1163 ( .A1(n1392), .A2(n1360), .S0(n559), .Y(n2047) );
  MUX21X1_HVT U1164 ( .A1(n1393), .A2(n254), .S0(n558), .Y(n2023) );
  MUX21X1_HVT U1165 ( .A1(n1360), .A2(n1756), .S0(n557), .Y(n2019) );
  MUX21X1_HVT U1166 ( .A1(n1363), .A2(n1753), .S0(n558), .Y(n2030) );
  MUX21X1_HVT U1167 ( .A1(n1406), .A2(n2487), .S0(n560), .Y(n2459) );
  MUX21X1_HVT U1168 ( .A1(n1397), .A2(n2270), .S0(n1422), .Y(n2242) );
  MUX21X1_HVT U1169 ( .A1(n1719), .A2(n2029), .S0(n1339), .Y(n1927) );
  MUX21X1_HVT U1170 ( .A1(n2000), .A2(n2002), .S0(n1341), .Y(n1999) );
  MUX21X1_HVT U1171 ( .A1(n2489), .A2(n2350), .S0(n1242), .Y(n2349) );
  MUX21X1_HVT U1172 ( .A1(n2461), .A2(n2460), .S0(n1243), .Y(n2350) );
  MUX21X1_HVT U1173 ( .A1(n2272), .A2(n2133), .S0(n1232), .Y(n2132) );
  MUX21X1_HVT U1174 ( .A1(n2244), .A2(n2243), .S0(n1234), .Y(n2133) );
  MUX21X1_HVT U1175 ( .A1(n1918), .A2(n2052), .S0(n1340), .Y(n1917) );
  MUX21X1_HVT U1176 ( .A1(n2036), .A2(n1729), .S0(n1350), .Y(n1918) );
  MUX21X1_HVT U1177 ( .A1(n1864), .A2(n1863), .S0(n1341), .Y(n1862) );
  MUX21X1_HVT U1178 ( .A1(n1706), .A2(n1750), .S0(n1349), .Y(n1864) );
  MUX21X1_HVT U1179 ( .A1(n1697), .A2(n1725), .S0(n1339), .Y(n1939) );
  MUX21X1_HVT U1180 ( .A1(n1934), .A2(n1933), .S0(n1350), .Y(n1930) );
  MUX21X1_HVT U1181 ( .A1(n1700), .A2(n1935), .S0(n1343), .Y(n1934) );
  MUX21X1_HVT U1182 ( .A1(n1395), .A2(n1396), .S0(n1341), .Y(n1932) );
  MUX21X1_HVT U1183 ( .A1(n1362), .A2(n1360), .S0(n1467), .Y(n1935) );
  XOR2X1_HVT U1184 ( .A1(n290), .A2(n1752), .Y(n2014) );
  MUX21X1_HVT U1185 ( .A1(n1395), .A2(n1362), .S0(n1470), .Y(n1988) );
  MUX21X1_HVT U1186 ( .A1(n1392), .A2(n1395), .S0(n1470), .Y(n1970) );
  MUX21X1_HVT U1187 ( .A1(n1412), .A2(n599), .S0(n1436), .Y(n2286) );
  MUX21X1_HVT U1188 ( .A1(n1403), .A2(n1353), .S0(n1425), .Y(n2067) );
  MUX21X1_HVT U1189 ( .A1(n1395), .A2(n1360), .S0(n1468), .Y(n1849) );
  MUX21X1_HVT U1190 ( .A1(n1753), .A2(n1362), .S0(n291), .Y(n1845) );
  MUX21X1_HVT U1191 ( .A1(n1360), .A2(n254), .S0(n290), .Y(n1847) );
  MUX21X1_HVT U1192 ( .A1(n2029), .A2(n1852), .S0(n1348), .Y(n1846) );
  MUX21X1_HVT U1193 ( .A1(n1752), .A2(n1753), .S0(n559), .Y(n2040) );
  MUX21X1_HVT U1194 ( .A1(n1624), .A2(n1623), .S0(n562), .Y(n2469) );
  MUX21X1_HVT U1195 ( .A1(n1163), .A2(n1556), .S0(n218), .Y(n2252) );
  MUX21X1_HVT U1196 ( .A1(n1623), .A2(n1621), .S0(n560), .Y(n2457) );
  MUX21X1_HVT U1197 ( .A1(n1556), .A2(n1554), .S0(n1425), .Y(n2240) );
  MUX21X1_HVT U1198 ( .A1(n1355), .A2(n599), .S0(n1438), .Y(n2476) );
  MUX21X1_HVT U1199 ( .A1(n1352), .A2(n1353), .S0(n1425), .Y(n2259) );
  MUX21X1_HVT U1200 ( .A1(n1410), .A2(n1412), .S0(n1439), .Y(n2478) );
  MUX21X1_HVT U1201 ( .A1(n1401), .A2(n1403), .S0(n1422), .Y(n2261) );
  MUX21X1_HVT U1202 ( .A1(n1623), .A2(n599), .S0(n562), .Y(n2463) );
  MUX21X1_HVT U1203 ( .A1(n1556), .A2(n1353), .S0(n218), .Y(n2246) );
  MUX21X1_HVT U1204 ( .A1(n2487), .A2(n1624), .S0(n1438), .Y(n2471) );
  MUX21X1_HVT U1205 ( .A1(n2270), .A2(n1163), .S0(n1422), .Y(n2254) );
  MUX21X1_HVT U1206 ( .A1(n1408), .A2(n1355), .S0(n562), .Y(n2454) );
  MUX21X1_HVT U1207 ( .A1(n1399), .A2(n1352), .S0(n1424), .Y(n2237) );
  MUX21X1_HVT U1208 ( .A1(n599), .A2(n1623), .S0(n1440), .Y(n2484) );
  MUX21X1_HVT U1209 ( .A1(n1353), .A2(n1556), .S0(n1424), .Y(n2267) );
  MUX21X1_HVT U1210 ( .A1(n1391), .A2(n1757), .S0(n557), .Y(n2018) );
  MUX21X1_HVT U1211 ( .A1(n1409), .A2(n599), .S0(n561), .Y(n2481) );
  MUX21X1_HVT U1212 ( .A1(n1400), .A2(n1353), .S0(n1422), .Y(n2264) );
  MUX21X1_HVT U1213 ( .A1(n599), .A2(n1624), .S0(n561), .Y(n2455) );
  MUX21X1_HVT U1214 ( .A1(n1353), .A2(n1163), .S0(n1424), .Y(n2238) );
  MUX21X1_HVT U1215 ( .A1(n1356), .A2(n1623), .S0(n1437), .Y(n2486) );
  MUX21X1_HVT U1216 ( .A1(n1553), .A2(n1556), .S0(n1426), .Y(n2269) );
  MUX21X1_HVT U1217 ( .A1(n1407), .A2(n599), .S0(n1440), .Y(n2483) );
  MUX21X1_HVT U1218 ( .A1(n1398), .A2(n1353), .S0(n218), .Y(n2266) );
  MUX21X1_HVT U1219 ( .A1(n1354), .A2(n1625), .S0(n1440), .Y(n2395) );
  MUX21X1_HVT U1220 ( .A1(n1351), .A2(n1557), .S0(n1424), .Y(n2177) );
  MUX21X1_HVT U1221 ( .A1(n1407), .A2(n1412), .S0(n562), .Y(n2406) );
  MUX21X1_HVT U1222 ( .A1(n1398), .A2(n1404), .S0(n218), .Y(n2189) );
  MUX21X1_HVT U1223 ( .A1(n1412), .A2(n1356), .S0(n561), .Y(n2387) );
  MUX21X1_HVT U1224 ( .A1(n1403), .A2(n1351), .S0(n1426), .Y(n2169) );
  MUX21X1_HVT U1225 ( .A1(n1499), .A2(n1526), .S0(n1429), .Y(n2149) );
  XOR2X1_HVT U1226 ( .A1(n1416), .A2(n1454), .Y(n2668) );
  MUX21X1_HVT U1227 ( .A1(n1621), .A2(n1624), .S0(n562), .Y(n2319) );
  MUX21X1_HVT U1228 ( .A1(n1554), .A2(n1163), .S0(n218), .Y(n2100) );
  MUX21X1_HVT U1229 ( .A1(n2715), .A2(n1418), .S0(n1456), .Y(n2527) );
  MUX21X1_HVT U1230 ( .A1(n599), .A2(n1625), .S0(n561), .Y(n2305) );
  MUX21X1_HVT U1231 ( .A1(n1555), .A2(n1557), .S0(n1423), .Y(n2086) );
  MUX21X1_HVT U1232 ( .A1(n2487), .A2(n1625), .S0(n1438), .Y(n2414) );
  MUX21X1_HVT U1233 ( .A1(n2270), .A2(n1557), .S0(n1424), .Y(n2197) );
  MUX21X1_HVT U1234 ( .A1(n254), .A2(n1752), .S0(n1470), .Y(n1844) );
  MUX21X1_HVT U1235 ( .A1(n1391), .A2(n1362), .S0(n1469), .Y(n1851) );
  MUX21X1_HVT U1236 ( .A1(n599), .A2(n2487), .S0(n1438), .Y(n2284) );
  MUX21X1_HVT U1237 ( .A1(n1555), .A2(n2270), .S0(n1425), .Y(n2065) );
  MUX21X1_HVT U1238 ( .A1(n2686), .A2(n2506), .S0(n270), .Y(n2500) );
  MUX21X1_HVT U1239 ( .A1(n2487), .A2(n1619), .S0(n1436), .Y(n2281) );
  MUX21X1_HVT U1240 ( .A1(n2270), .A2(n1552), .S0(n1426), .Y(n2062) );
  MUX21X1_HVT U1241 ( .A1(n1408), .A2(n1625), .S0(n1438), .Y(n2288) );
  MUX21X1_HVT U1242 ( .A1(n1399), .A2(n1557), .S0(n1426), .Y(n2069) );
  AND2X1_HVT U1243 ( .A1(n1455), .A2(n1688), .Y(n1204) );
  MUX21X1_HVT U1244 ( .A1(n1625), .A2(n1621), .S0(n1437), .Y(n2467) );
  MUX21X1_HVT U1245 ( .A1(n1557), .A2(n1554), .S0(n1425), .Y(n2250) );
  MUX21X1_HVT U1246 ( .A1(n1577), .A2(n1619), .S0(n1241), .Y(n2428) );
  MUX21X1_HVT U1247 ( .A1(n1509), .A2(n1552), .S0(n1231), .Y(n2211) );
  MUX21X1_HVT U1248 ( .A1(n2475), .A2(n1593), .S0(n1444), .Y(n2359) );
  MUX21X1_HVT U1249 ( .A1(n2258), .A2(n1525), .S0(n1429), .Y(n2142) );
  MUX21X1_HVT U1250 ( .A1(n1621), .A2(n1623), .S0(n1241), .Y(n2443) );
  MUX21X1_HVT U1251 ( .A1(n1554), .A2(n1556), .S0(n1231), .Y(n2226) );
  MUX21X1_HVT U1252 ( .A1(n1683), .A2(n1688), .S0(n1453), .Y(n2555) );
  MUX21X1_HVT U1253 ( .A1(n1687), .A2(n1684), .S0(n1456), .Y(n2557) );
  MUX21X1_HVT U1254 ( .A1(n1359), .A2(n1421), .S0(n1454), .Y(n2525) );
  XOR2X1_HVT U1255 ( .A1(n2033), .A2(n1469), .Y(n2013) );
  MUX21X1_HVT U1258 ( .A1(n1619), .A2(n1621), .S0(n1436), .Y(n2482) );
  MUX21X1_HVT U1259 ( .A1(n1552), .A2(n1554), .S0(n1425), .Y(n2265) );
  MUX21X1_HVT U1261 ( .A1(n1358), .A2(n1687), .S0(n1455), .Y(n2705) );
  MUX21X1_HVT U1262 ( .A1(n1417), .A2(n1359), .S0(n277), .Y(n2702) );
  MUX21X1_HVT U1263 ( .A1(n1683), .A2(n1685), .S0(n214), .Y(n2703) );
  MUX21X1_HVT U1264 ( .A1(n1658), .A2(n2712), .S0(n1459), .Y(n2604) );
  MUX21X1_HVT U1265 ( .A1(n1684), .A2(n1685), .S0(n1452), .Y(n2613) );
  XOR2X1_HVT U1266 ( .A1(n2487), .A2(n1439), .Y(n2449) );
  XOR2X1_HVT U1267 ( .A1(n2270), .A2(n1425), .Y(n2232) );
  XOR2X1_HVT U1268 ( .A1(n1363), .A2(n1469), .Y(n2015) );
  XNOR2X1_HVT U1269 ( .A1(n1392), .A2(n1468), .Y(n1205) );
  MUX21X1_HVT U1270 ( .A1(n1416), .A2(n1689), .S0(n1456), .Y(n2505) );
  XNOR2X1_HVT U1271 ( .A1(n1396), .A2(n291), .Y(n1206) );
  MUX21X1_HVT U1272 ( .A1(n1688), .A2(n1687), .S0(n1455), .Y(n2690) );
  MUX21X1_HVT U1273 ( .A1(n1687), .A2(n1685), .S0(n214), .Y(n2678) );
  MUX21X1_HVT U1274 ( .A1(n1684), .A2(n1358), .S0(n217), .Y(n2697) );
  MUX21X1_HVT U1275 ( .A1(n1418), .A2(n1419), .S0(n1452), .Y(n2699) );
  MUX21X1_HVT U1276 ( .A1(n1687), .A2(n1359), .S0(n1452), .Y(n2684) );
  MUX21X1_HVT U1277 ( .A1(n1407), .A2(n1413), .S0(n1438), .Y(n2401) );
  MUX21X1_HVT U1278 ( .A1(n1398), .A2(n1405), .S0(n1424), .Y(n2183) );
  MUX21X1_HVT U1280 ( .A1(n1757), .A2(n1755), .S0(n1470), .Y(n2050) );
  MUX21X1_HVT U1282 ( .A1(n1414), .A2(n244), .S0(n1453), .Y(n2680) );
  MUX21X1_HVT U1283 ( .A1(n1415), .A2(n1358), .S0(n1456), .Y(n2704) );
  MUX21X1_HVT U1284 ( .A1(n1621), .A2(n1625), .S0(n1438), .Y(n2282) );
  MUX21X1_HVT U1285 ( .A1(n1554), .A2(n1557), .S0(n1426), .Y(n2063) );
  MUX21X1_HVT U1286 ( .A1(n1640), .A2(n1683), .S0(n1252), .Y(n2649) );
  MUX21X1_HVT U1287 ( .A1(n2687), .A2(n2602), .S0(n1459), .Y(n2600) );
  MUX21X1_HVT U1288 ( .A1(n1408), .A2(n1407), .S0(n1438), .Y(n2280) );
  MUX21X1_HVT U1289 ( .A1(n1399), .A2(n1398), .S0(n1422), .Y(n2061) );
  MUX21X1_HVT U1290 ( .A1(n1685), .A2(n1687), .S0(n1252), .Y(n2664) );
  MUX21X1_HVT U1291 ( .A1(n1685), .A2(n1688), .S0(n277), .Y(n2536) );
  MUX21X1_HVT U1292 ( .A1(n1357), .A2(n1689), .S0(n1453), .Y(n2522) );
  XNOR2X1_HVT U1293 ( .A1(n2494), .A2(n1436), .Y(n1207) );
  XNOR2X1_HVT U1294 ( .A1(n2277), .A2(n1424), .Y(n1208) );
  XOR2X1_HVT U1295 ( .A1(n1237), .A2(n1436), .Y(n2453) );
  XOR2X1_HVT U1297 ( .A1(n1227), .A2(n1422), .Y(n2236) );
  MUX21X1_HVT U1298 ( .A1(n1419), .A2(n1359), .S0(n1456), .Y(n2503) );
  MUX21X1_HVT U1299 ( .A1(n1753), .A2(n1755), .S0(n1347), .Y(n2007) );
  XOR2X1_HVT U1300 ( .A1(n291), .A2(n1346), .Y(n2017) );
  MUX21X1_HVT U1301 ( .A1(n1391), .A2(n1392), .S0(n1468), .Y(n1843) );
  XNOR2X1_HVT U1302 ( .A1(n1406), .A2(n1439), .Y(n1209) );
  XNOR2X1_HVT U1304 ( .A1(n1398), .A2(n1426), .Y(n1210) );
  MUX21X1_HVT U1305 ( .A1(n2715), .A2(n1419), .S0(n1455), .Y(n2687) );
  MUX21X1_HVT U1307 ( .A1(n1416), .A2(n1684), .S0(n277), .Y(n2675) );
  MUX21X1_HVT U1308 ( .A1(n1360), .A2(n1755), .S0(n290), .Y(n2048) );
  MUX21X1_HVT U1309 ( .A1(n1358), .A2(n1688), .S0(n1456), .Y(n2676) );
  MUX21X1_HVT U1310 ( .A1(n1684), .A2(n1687), .S0(n1452), .Y(n2707) );
  MUX21X1_HVT U1311 ( .A1(n243), .A2(n1689), .S0(n1453), .Y(n2615) );
  MUX21X1_HVT U1312 ( .A1(n244), .A2(n1683), .S0(n1454), .Y(n2498) );
  MUX21X1_HVT U1313 ( .A1(n1414), .A2(n1420), .S0(n277), .Y(n2627) );
  MUX21X1_HVT U1314 ( .A1(n1630), .A2(n1657), .S0(n1459), .Y(n2586) );
  MUX21X1_HVT U1316 ( .A1(n244), .A2(n1689), .S0(n1455), .Y(n2635) );
  MUX21X1_HVT U1318 ( .A1(n1689), .A2(n1685), .S0(n1454), .Y(n2688) );
  MUX21X1_HVT U1319 ( .A1(n244), .A2(n1688), .S0(n214), .Y(n2692) );
  MUX21X1_HVT U1320 ( .A1(n1651), .A2(n2686), .S0(n901), .Y(n2582) );
  MUX21X1_HVT U1322 ( .A1(n1357), .A2(n244), .S0(n1454), .Y(n2501) );
  MUX21X1_HVT U1323 ( .A1(n1419), .A2(n1684), .S0(n277), .Y(n2607) );
  NBUFFX2_HVT U1328 ( .A(n2492), .Y(n1409) );
  NBUFFX2_HVT U1329 ( .A(n2275), .Y(n1400) );
  XOR2X1_HVT U1330 ( .A1(n1248), .A2(n1452), .Y(n2674) );
  NBUFFX2_HVT U1332 ( .A(n2492), .Y(n1408) );
  NBUFFX2_HVT U1334 ( .A(n2275), .Y(n1399) );
  NAND2X0_HVT U1336 ( .A1(n1622), .A2(n1625), .Y(n2488) );
  NAND2X0_HVT U1338 ( .A1(n1353), .A2(n1557), .Y(n2271) );
  INVX0_HVT U1340 ( .A(n2487), .Y(n1620) );
  INVX0_HVT U1342 ( .A(n2270), .Y(n1553) );
  MUX21X1_HVT U1344 ( .A1(n1213), .A2(n1646), .S0(n1460), .Y(n2580) );
  MUX21X1_HVT U1345 ( .A1(n2696), .A2(n1656), .S0(n902), .Y(n2579) );
  NBUFFX2_HVT U1346 ( .A(n2713), .Y(n1417) );
  NBUFFX2_HVT U1348 ( .A(n2492), .Y(n1410) );
  NBUFFX2_HVT U1349 ( .A(n2275), .Y(n1401) );
  XOR2X1_HVT U1350 ( .A1(n2708), .A2(n217), .Y(n2670) );
  XNOR2X1_HVT U1351 ( .A1(n1421), .A2(n1452), .Y(n1211) );
  AND2X1_HVT U1352 ( .A1(n1756), .A2(n290), .Y(n1212) );
  NBUFFX2_HVT U1353 ( .A(n2493), .Y(n1411) );
  NBUFFX2_HVT U1354 ( .A(n2276), .Y(n1402) );
  MUX21X1_HVT U1356 ( .A1(n1414), .A2(n1421), .S0(n1453), .Y(n2621) );
  MUX21X1_HVT U1357 ( .A1(n2493), .A2(n1413), .S0(n1444), .Y(n2373) );
  MUX21X1_HVT U1358 ( .A1(n1404), .A2(n1405), .S0(n1429), .Y(n2155) );
  NAND2X0_HVT U1360 ( .A1(n1357), .A2(n1689), .Y(n2709) );
  MUX21X1_HVT U1362 ( .A1(n1416), .A2(n1415), .S0(n214), .Y(n2497) );
  NBUFFX2_HVT U1363 ( .A(n2057), .Y(n1394) );
  XNOR2X1_HVT U1364 ( .A1(n1415), .A2(n217), .Y(n1213) );
  MUX21X1_HVT U1366 ( .A1(n1685), .A2(n1689), .S0(n1456), .Y(n2499) );
  NBUFFX2_HVT U1368 ( .A(n1758), .Y(n1363) );
  NBUFFX2_HVT U1370 ( .A(n2055), .Y(n1390) );
  NBUFFX2_HVT U1372 ( .A(n2713), .Y(n1418) );
  NBUFFX2_HVT U1374 ( .A(n2057), .Y(n1395) );
  NBUFFX2_HVT U1377 ( .A(n2713), .Y(n1416) );
  NBUFFX2_HVT U1378 ( .A(n2055), .Y(n1391) );
  NBUFFX2_HVT U1379 ( .A(n2493), .Y(n1412) );
  NBUFFX2_HVT U1380 ( .A(n2276), .Y(n1403) );
  NBUFFX2_HVT U1381 ( .A(n2276), .Y(n1404) );
  NBUFFX2_HVT U1382 ( .A(keyin[112]), .Y(n1244) );
  NBUFFX2_HVT U1383 ( .A(n1434), .Y(n1234) );
  NBUFFX2_HVT U1385 ( .A(n2494), .Y(n1413) );
  NBUFFX2_HVT U1388 ( .A(n2277), .Y(n1405) );
  NBUFFX2_HVT U1389 ( .A(n2058), .Y(n1396) );
  NBUFFX2_HVT U1390 ( .A(keyin[112]), .Y(n1243) );
  NBUFFX2_HVT U1391 ( .A(n1434), .Y(n1233) );
  NBUFFX2_HVT U1392 ( .A(keyin[98]), .Y(n1347) );
  NBUFFX2_HVT U1393 ( .A(n1478), .Y(n1350) );
  NBUFFX2_HVT U1394 ( .A(n1478), .Y(n1349) );
  MUX21X1_HVT U1395 ( .A1(n1420), .A2(n1421), .S0(n1459), .Y(n2593) );
  NBUFFX2_HVT U1396 ( .A(keyin[98]), .Y(n1346) );
  NBUFFX2_HVT U1397 ( .A(n1478), .Y(n1348) );
  NBUFFX2_HVT U1398 ( .A(n1474), .Y(n1339) );
  NBUFFX2_HVT U1399 ( .A(n1754), .Y(n1360) );
  NBUFFX2_HVT U1400 ( .A(n2714), .Y(n1419) );
  NBUFFX2_HVT U1401 ( .A(n2714), .Y(n1420) );
  NBUFFX2_HVT U1402 ( .A(n1474), .Y(n1343) );
  NBUFFX2_HVT U1403 ( .A(n1555), .Y(n1353) );
  NBUFFX2_HVT U1404 ( .A(n1758), .Y(n1362) );
  NBUFFX2_HVT U1405 ( .A(n2715), .Y(n1421) );
  NBUFFX2_HVT U1406 ( .A(n1465), .Y(n1255) );
  NBUFFX2_HVT U1407 ( .A(n1474), .Y(n1342) );
  NBUFFX2_HVT U1408 ( .A(n1474), .Y(n1340) );
  NBUFFX2_HVT U1409 ( .A(keyin[98]), .Y(n1344) );
  NBUFFX2_HVT U1410 ( .A(keyin[98]), .Y(n1345) );
  NBUFFX2_HVT U1411 ( .A(n1465), .Y(n1254) );
  NBUFFX2_HVT U1412 ( .A(n1474), .Y(n1341) );
  NBUFFX2_HVT U1413 ( .A(n1343), .Y(n1338) );
  NBUFFX2_HVT U1414 ( .A(n1686), .Y(n1358) );
  NBUFFX2_HVT U1415 ( .A(n1686), .Y(n1359) );
  MUX21X1_HVT U1416 ( .A1(n1365), .A2(n1557), .S0(n1234), .Y(n2187) );
  XNOR2X1_HVT U1417 ( .A1(n1441), .A2(n1449), .Y(n1214) );
  MUX21X1_HVT U1418 ( .A1(n2347), .A2(n2346), .S0(n1242), .Y(n2345) );
  MUX21X1_HVT U1419 ( .A1(n2423), .A2(n2449), .S0(n1449), .Y(n2347) );
  MUX21X1_HVT U1420 ( .A1(n2341), .A2(n2340), .S0(n1241), .Y(n2338) );
  MUX21X1_HVT U1421 ( .A1(n2382), .A2(n1410), .S0(n1243), .Y(n2341) );
  XNOR2X1_HVT U1422 ( .A1(n1457), .A2(n554), .Y(n1216) );
  MUX21X1_HVT U1423 ( .A1(n2644), .A2(n2670), .S0(n555), .Y(n2567) );
  MUX21X1_HVT U1424 ( .A1(n2602), .A2(n1418), .S0(n554), .Y(n2561) );
  XOR2X1_HVT U1425 ( .A1(n1795), .A2(n1839), .Y(keyout[3]) );
  XNOR2X1_HVT U1426 ( .A1(n1833), .A2(n1834), .Y(keyout[65]) );
  MUX21X1_HVT U1429 ( .A1(n1386), .A2(n1389), .S0(n1343), .Y(n1944) );
  MUX21X1_HVT U1442 ( .A1(n1726), .A2(n2056), .S0(n1343), .Y(n1949) );
  MUX21X1_HVT U1443 ( .A1(n2028), .A2(n1947), .S0(n1339), .Y(n1945) );
  MUX21X1_HVT U1444 ( .A1(n1366), .A2(n1368), .S0(n604), .Y(n2161) );
  MUX21X1_HVT U1445 ( .A1(n1381), .A2(n1384), .S0(n1459), .Y(n2599) );
  MUX21X1_HVT U1446 ( .A1(n1386), .A2(n2054), .S0(n1347), .Y(n2009) );
  MUX21X1_HVT U1447 ( .A1(n1205), .A2(n1712), .S0(n1342), .Y(n1925) );
  MUX21X1_HVT U1450 ( .A1(n2041), .A2(n1724), .S0(n1340), .Y(n1924) );
  INVX1_HVT U1454 ( .A(n1441), .Y(n1440) );
  INVX1_HVT U1460 ( .A(n1427), .Y(n1426) );
  MUX21X1_HVT U1463 ( .A1(n1412), .A2(n2328), .S0(n1244), .Y(n2327) );
  MUX21X1_HVT U1467 ( .A1(n2107), .A2(n2108), .S0(n1231), .Y(n2106) );
  MUX21X1_HVT U1474 ( .A1(n1404), .A2(n2109), .S0(n1234), .Y(n2108) );
  MUX21X1_HVT U1475 ( .A1(n1389), .A2(n1391), .S0(n558), .Y(n2038) );
  MUX21X1_HVT U1476 ( .A1(n2042), .A2(n1199), .S0(n1348), .Y(n1860) );
  MUX21X1_HVT U1477 ( .A1(n1755), .A2(n1742), .S0(n1350), .Y(n1990) );
  MUX21X1_HVT U1478 ( .A1(n2422), .A2(n2451), .S0(n1241), .Y(n2421) );
  XOR2X1_HVT U1479 ( .A1(n280), .A2(n2469), .Y(n2451) );
  MUX21X1_HVT U1480 ( .A1(n2425), .A2(n2424), .S0(n1243), .Y(n2422) );
  MUX21X1_HVT U1481 ( .A1(n1412), .A2(n1625), .S0(n561), .Y(n2425) );
  MUX21X1_HVT U1482 ( .A1(n2205), .A2(n2234), .S0(n1231), .Y(n2204) );
  MUX21X1_HVT U1483 ( .A1(n2208), .A2(n2207), .S0(n1233), .Y(n2205) );
  MUX21X1_HVT U1484 ( .A1(n1404), .A2(n1557), .S0(n1424), .Y(n2208) );
  MUX21X1_HVT U1485 ( .A1(n2491), .A2(n1442), .S0(n1444), .Y(n2372) );
  MUX21X1_HVT U1486 ( .A1(n2274), .A2(n1428), .S0(n1429), .Y(n2154) );
  MUX21X1_HVT U1487 ( .A1(n1388), .A2(n1755), .S0(n557), .Y(n2024) );
  MUX21X1_HVT U1488 ( .A1(n1393), .A2(n1386), .S0(n558), .Y(n2049) );
  MUX21X1_HVT U1489 ( .A1(n1388), .A2(n1752), .S0(n559), .Y(n2041) );
  MUX21X1_HVT U1490 ( .A1(n1374), .A2(n1623), .S0(n560), .Y(n2460) );
  MUX21X1_HVT U1491 ( .A1(n1368), .A2(n1556), .S0(n1426), .Y(n2243) );
  MUX21X1_HVT U1492 ( .A1(n1360), .A2(n1389), .S0(n557), .Y(n2029) );
  MUX21X1_HVT U1493 ( .A1(n1387), .A2(n1753), .S0(n559), .Y(n2021) );
  MUX21X1_HVT U1494 ( .A1(n1753), .A2(n1388), .S0(n559), .Y(n2027) );
  MUX21X1_HVT U1495 ( .A1(n1391), .A2(n1968), .S0(n1217), .Y(n1967) );
  MUX21X1_HVT U1496 ( .A1(n1387), .A2(n1362), .S0(n1350), .Y(n1968) );
  MUX21X1_HVT U1497 ( .A1(n1906), .A2(n1907), .S0(n1342), .Y(n1904) );
  MUX21X1_HVT U1498 ( .A1(n1744), .A2(n1752), .S0(n1350), .Y(n1907) );
  MUX21X1_HVT U1499 ( .A1(n1875), .A2(n1876), .S0(n1343), .Y(n1874) );
  MUX21X1_HVT U1500 ( .A1(n1973), .A2(n1386), .S0(n1349), .Y(n1876) );
  MUX21X1_HVT U1501 ( .A1(n1888), .A2(n1887), .S0(n1342), .Y(n1886) );
  MUX21X1_HVT U1502 ( .A1(n1395), .A2(n1742), .S0(n1350), .Y(n1888) );
  MUX21X1_HVT U1503 ( .A1(n1900), .A2(n1901), .S0(n1343), .Y(n1899) );
  MUX21X1_HVT U1504 ( .A1(n1902), .A2(n1391), .S0(n1217), .Y(n1901) );
  MUX21X1_HVT U1505 ( .A1(n2022), .A2(n1745), .S0(n1349), .Y(n1900) );
  MUX21X1_HVT U1506 ( .A1(n1912), .A2(n1911), .S0(n1340), .Y(n1910) );
  MUX21X1_HVT U1507 ( .A1(n2030), .A2(n1703), .S0(n1349), .Y(n1912) );
  MUX21X1_HVT U1508 ( .A1(n1388), .A2(n2057), .S0(n1469), .Y(n1842) );
  MUX21X1_HVT U1509 ( .A1(n1356), .A2(n1371), .S0(n1437), .Y(n2472) );
  MUX21X1_HVT U1510 ( .A1(n1553), .A2(n1365), .S0(n1426), .Y(n2255) );
  MUX21X1_HVT U1511 ( .A1(n1406), .A2(n1372), .S0(n1436), .Y(n2485) );
  MUX21X1_HVT U1512 ( .A1(n1397), .A2(n1366), .S0(n1425), .Y(n2268) );
  MUX21X1_HVT U1513 ( .A1(n1375), .A2(n1410), .S0(n1438), .Y(n2474) );
  MUX21X1_HVT U1514 ( .A1(n1368), .A2(n1401), .S0(n1424), .Y(n2257) );
  MUX21X1_HVT U1515 ( .A1(n1371), .A2(n1621), .S0(n561), .Y(n2458) );
  MUX21X1_HVT U1516 ( .A1(n1365), .A2(n1554), .S0(n218), .Y(n2241) );
  MUX21X1_HVT U1517 ( .A1(n1413), .A2(n1374), .S0(n1438), .Y(n2468) );
  MUX21X1_HVT U1518 ( .A1(n1405), .A2(n1368), .S0(n1422), .Y(n2251) );
  MUX21X1_HVT U1519 ( .A1(n1396), .A2(n1388), .S0(n558), .Y(n2031) );
  MUX21X1_HVT U1520 ( .A1(n2315), .A2(n2316), .S0(n1242), .Y(n2314) );
  MUX21X1_HVT U1521 ( .A1(n1597), .A2(n1406), .S0(n1243), .Y(n2316) );
  MUX21X1_HVT U1522 ( .A1(n2096), .A2(n2097), .S0(n1232), .Y(n2095) );
  MUX21X1_HVT U1523 ( .A1(n1529), .A2(n1397), .S0(n1234), .Y(n2097) );
  MUX21X1_HVT U1524 ( .A1(n1710), .A2(n1471), .S0(n1347), .Y(n1994) );
  MUX21X1_HVT U1525 ( .A1(n1371), .A2(n1619), .S0(n1436), .Y(n2285) );
  MUX21X1_HVT U1526 ( .A1(n1365), .A2(n1552), .S0(n1425), .Y(n2066) );
  MUX21X1_HVT U1527 ( .A1(n1372), .A2(n2462), .S0(n1242), .Y(n2445) );
  MUX21X1_HVT U1528 ( .A1(n1366), .A2(n2245), .S0(n1232), .Y(n2228) );
  XOR2X1_HVT U1529 ( .A1(n1386), .A2(n290), .Y(n2012) );
  MUX21X1_HVT U1530 ( .A1(n1374), .A2(n1412), .S0(n1436), .Y(n2279) );
  MUX21X1_HVT U1531 ( .A1(n1368), .A2(n1404), .S0(n1426), .Y(n2060) );
  MUX21X1_HVT U1532 ( .A1(n1387), .A2(n1752), .S0(n291), .Y(n1848) );
  MUX21X1_HVT U1533 ( .A1(n1389), .A2(n254), .S0(n290), .Y(n1850) );
  NBUFFX2_HVT U1534 ( .A(n1448), .Y(n1242) );
  NBUFFX2_HVT U1535 ( .A(n1433), .Y(n1232) );
  MUX21X1_HVT U1536 ( .A1(n1374), .A2(n1619), .S0(n1440), .Y(n2475) );
  MUX21X1_HVT U1537 ( .A1(n1368), .A2(n1552), .S0(n1422), .Y(n2258) );
  MUX21X1_HVT U1538 ( .A1(n599), .A2(n1375), .S0(n1440), .Y(n2465) );
  MUX21X1_HVT U1539 ( .A1(n1353), .A2(n1368), .S0(n1425), .Y(n2248) );
  MUX21X1_HVT U1540 ( .A1(n1621), .A2(n1374), .S0(n1437), .Y(n2464) );
  MUX21X1_HVT U1541 ( .A1(n1554), .A2(n1368), .S0(n1423), .Y(n2247) );
  MUX21X1_HVT U1542 ( .A1(n1579), .A2(n1442), .S0(n1241), .Y(n2430) );
  MUX21X1_HVT U1543 ( .A1(n1511), .A2(n1428), .S0(n1231), .Y(n2213) );
  XNOR2X1_HVT U1544 ( .A1(n1480), .A2(n1467), .Y(n1217) );
  MUX21X1_HVT U1545 ( .A1(n1375), .A2(n2487), .S0(n1436), .Y(n2287) );
  MUX21X1_HVT U1546 ( .A1(n1368), .A2(n2270), .S0(n1423), .Y(n2068) );
  NBUFFX2_HVT U1547 ( .A(n1448), .Y(n1241) );
  NBUFFX2_HVT U1548 ( .A(n1433), .Y(n1231) );
  MUX21X1_HVT U1549 ( .A1(n1384), .A2(n1418), .S0(n1454), .Y(n2695) );
  MUX21X1_HVT U1550 ( .A1(n1381), .A2(n2683), .S0(n1253), .Y(n2666) );
  MUX21X1_HVT U1551 ( .A1(n2712), .A2(n1458), .S0(n1459), .Y(n2592) );
  MUX21X1_HVT U1552 ( .A1(n1389), .A2(n1396), .S0(n1470), .Y(n1841) );
  MUX21X1_HVT U1553 ( .A1(n1384), .A2(n244), .S0(n214), .Y(n2504) );
  NBUFFX2_HVT U1554 ( .A(n1462), .Y(n1253) );
  MUX21X1_HVT U1555 ( .A1(n1414), .A2(n1381), .S0(n214), .Y(n2706) );
  MUX21X1_HVT U1556 ( .A1(n1383), .A2(n1683), .S0(n1456), .Y(n2696) );
  MUX21X1_HVT U1557 ( .A1(n1383), .A2(n1687), .S0(n217), .Y(n2681) );
  MUX21X1_HVT U1558 ( .A1(n1380), .A2(n1685), .S0(n277), .Y(n2679) );
  MUX21X1_HVT U1559 ( .A1(n1642), .A2(n1458), .S0(n1252), .Y(n2651) );
  MUX21X1_HVT U1560 ( .A1(n2681), .A2(n2704), .S0(n556), .Y(n2518) );
  XOR2X1_HVT U1561 ( .A1(n1466), .A2(n2690), .Y(n2672) );
  MUX21X1_HVT U1562 ( .A1(n2646), .A2(n2645), .S0(n270), .Y(n2643) );
  MUX21X1_HVT U1563 ( .A1(n1420), .A2(n1689), .S0(n217), .Y(n2646) );
  MUX21X1_HVT U1564 ( .A1(n1383), .A2(n1420), .S0(n1452), .Y(n2496) );
  XOR2X1_HVT U1565 ( .A1(n1372), .A2(n1437), .Y(n2448) );
  XOR2X1_HVT U1566 ( .A1(n1366), .A2(n1425), .Y(n2231) );
  MUX21X1_HVT U1567 ( .A1(n1375), .A2(n1413), .S0(n1440), .Y(n2278) );
  MUX21X1_HVT U1568 ( .A1(n1368), .A2(n1405), .S0(n1422), .Y(n2059) );
  NBUFFX2_HVT U1569 ( .A(n1462), .Y(n1252) );
  MUX21X1_HVT U1570 ( .A1(n1685), .A2(n1383), .S0(n214), .Y(n2685) );
  MUX21X1_HVT U1571 ( .A1(n1421), .A2(n1383), .S0(n1454), .Y(n2689) );
  MUX21X1_HVT U1572 ( .A1(n2056), .A2(n1472), .S0(n1341), .Y(n1931) );
  INVX1_HVT U1573 ( .A(keyin[99]), .Y(n1758) );
  NBUFFX2_HVT U1574 ( .A(n1448), .Y(n1240) );
  NBUFFX2_HVT U1575 ( .A(n1433), .Y(n1230) );
  MUX21X1_HVT U1576 ( .A1(n1359), .A2(n1384), .S0(n1455), .Y(n2686) );
  MUX21X1_HVT U1577 ( .A1(n1380), .A2(n1683), .S0(n1455), .Y(n2502) );
  NAND2X0_HVT U1578 ( .A1(n1625), .A2(n1372), .Y(n2492) );
  NAND2X0_HVT U1579 ( .A1(n1557), .A2(n1366), .Y(n2275) );
  INVX1_HVT U1580 ( .A(n1375), .Y(n1625) );
  INVX1_HVT U1581 ( .A(keyin[123]), .Y(n1557) );
  INVX1_HVT U1582 ( .A(n1457), .Y(n1452) );
  INVX1_HVT U1583 ( .A(keyin[116]), .Y(n1622) );
  INVX1_HVT U1584 ( .A(keyin[124]), .Y(n1555) );
  NAND2X0_HVT U1585 ( .A1(n1689), .A2(n1381), .Y(n2713) );
  NAND2X0_HVT U1586 ( .A1(n1373), .A2(n1622), .Y(n2493) );
  NAND2X0_HVT U1587 ( .A1(n1367), .A2(n1555), .Y(n2276) );
  MUX21X1_HVT U1588 ( .A1(n1384), .A2(n1421), .S0(n217), .Y(n2495) );
  INVX1_HVT U1589 ( .A(n1384), .Y(n1689) );
  NAND2X0_HVT U1590 ( .A1(n1373), .A2(n1371), .Y(n2494) );
  NAND2X0_HVT U1591 ( .A1(n1367), .A2(n1365), .Y(n2277) );
  NAND2X0_HVT U1592 ( .A1(n1754), .A2(n1389), .Y(n2057) );
  AND2X1_HVT U1593 ( .A1(n1356), .A2(n1442), .Y(n1218) );
  AND2X1_HVT U1594 ( .A1(n1351), .A2(n1428), .Y(n1219) );
  AND2X1_HVT U1595 ( .A1(n1757), .A2(n1472), .Y(n1220) );
  INVX1_HVT U1596 ( .A(n1379), .Y(n1686) );
  INVX1_HVT U1597 ( .A(n1387), .Y(n1754) );
  NBUFFX2_HVT U1598 ( .A(n1462), .Y(n1251) );
  XOR2X1_HVT U1599 ( .A1(n1379), .A2(n217), .Y(n2669) );
  NAND2X0_HVT U1600 ( .A1(n1386), .A2(n1388), .Y(n2058) );
  NAND2X0_HVT U1601 ( .A1(n1387), .A2(n1363), .Y(n2055) );
  NAND2X0_HVT U1602 ( .A1(n1382), .A2(n1357), .Y(n2714) );
  AND2X1_HVT U1603 ( .A1(n243), .A2(n1458), .Y(n1221) );
  XOR2X1_HVT U1604 ( .A1(n1442), .A2(n1373), .Y(n2452) );
  XOR2X1_HVT U1605 ( .A1(n1428), .A2(n1367), .Y(n2235) );
  NAND2X0_HVT U1606 ( .A1(n1382), .A2(n1380), .Y(n2715) );
  AND2X1_HVT U1607 ( .A1(n1442), .A2(n599), .Y(n1222) );
  AND2X1_HVT U1608 ( .A1(n1428), .A2(n1353), .Y(n1223) );
  AND2X1_HVT U1609 ( .A1(n1458), .A2(n1359), .Y(n1224) );
  NBUFFX2_HVT U1610 ( .A(n1447), .Y(n1237) );
  NBUFFX2_HVT U1611 ( .A(n1432), .Y(n1227) );
  XOR2X1_HVT U1612 ( .A1(n1458), .A2(n1382), .Y(n2673) );
  NBUFFX2_HVT U1613 ( .A(n1447), .Y(n1238) );
  NBUFFX2_HVT U1614 ( .A(n1432), .Y(n1228) );
  AND2X1_HVT U1615 ( .A1(n1754), .A2(n1472), .Y(n1225) );
  NBUFFX2_HVT U1616 ( .A(keyin[106]), .Y(n1248) );
  NBUFFX2_HVT U1617 ( .A(n1447), .Y(n1239) );
  NBUFFX2_HVT U1618 ( .A(n1432), .Y(n1229) );
  NBUFFX2_HVT U1619 ( .A(n1446), .Y(n1235) );
  NBUFFX2_HVT U1620 ( .A(n1431), .Y(n1226) );
  NBUFFX2_HVT U1621 ( .A(n1446), .Y(n1236) );
  NBUFFX2_HVT U1622 ( .A(keyin[106]), .Y(n1247) );
  NBUFFX2_HVT U1623 ( .A(n1462), .Y(n1246) );
  NBUFFX2_HVT U1624 ( .A(n1247), .Y(n1249) );
  NBUFFX2_HVT U1625 ( .A(keyin[106]), .Y(n1245) );
  NBUFFX2_HVT U1626 ( .A(n1245), .Y(n1250) );
  MUX21X1_HVT U1627 ( .A1(n2390), .A2(n2391), .S0(n1443), .Y(n2389) );
  XOR2X1_HVT U1628 ( .A1(keyin[69]), .A2(n1133), .Y(n1761) );
  XNOR2X1_HVT U1629 ( .A1(keyin[67]), .A2(n1388), .Y(n1838) );
  XOR2X1_HVT U1630 ( .A1(keyin[70]), .A2(n1468), .Y(n1763) );
  MUX21X1_HVT U1631 ( .A1(n1996), .A2(n1998), .S0(n1341), .Y(n1995) );
  NBUFFX2_HVT U1632 ( .A(keyin[114]), .Y(n1448) );
  NBUFFX2_HVT U1633 ( .A(keyin[122]), .Y(n1433) );
  NBUFFX2_HVT U1634 ( .A(keyin[106]), .Y(n1462) );
  NBUFFX2_HVT U1635 ( .A(keyin[115]), .Y(n1375) );
  NBUFFX2_HVT U1636 ( .A(keyin[115]), .Y(n1373) );
  NBUFFX2_HVT U1637 ( .A(keyin[123]), .Y(n1367) );
  NBUFFX2_HVT U1638 ( .A(keyin[107]), .Y(n1384) );
  NBUFFX2_HVT U1639 ( .A(keyin[116]), .Y(n1371) );
  NBUFFX2_HVT U1640 ( .A(keyin[124]), .Y(n1365) );
  NBUFFX2_HVT U1641 ( .A(keyin[108]), .Y(n1379) );
  NBUFFX2_HVT U1642 ( .A(keyin[100]), .Y(n1387) );
  NBUFFX2_HVT U1643 ( .A(keyin[107]), .Y(n1382) );
  NBUFFX2_HVT U1644 ( .A(keyin[116]), .Y(n1372) );
  NBUFFX2_HVT U1645 ( .A(keyin[124]), .Y(n1366) );
  INVX0_HVT U1646 ( .A(keyin[126]), .Y(n1428) );
  NBUFFX2_HVT U1647 ( .A(keyin[108]), .Y(n1380) );
  NBUFFX2_HVT U1648 ( .A(keyin[108]), .Y(n1381) );
  INVX0_HVT U1649 ( .A(keyin[110]), .Y(n1458) );
  INVX0_HVT U1650 ( .A(keyin[102]), .Y(n1472) );
  NBUFFX2_HVT U1651 ( .A(keyin[99]), .Y(n1388) );
  NBUFFX2_HVT U1652 ( .A(keyin[99]), .Y(n1389) );
  NBUFFX2_HVT U1653 ( .A(keyin[115]), .Y(n1374) );
  NBUFFX2_HVT U1654 ( .A(keyin[123]), .Y(n1368) );
  NBUFFX2_HVT U1655 ( .A(keyin[114]), .Y(n1447) );
  NBUFFX2_HVT U1656 ( .A(keyin[122]), .Y(n1432) );
  NBUFFX2_HVT U1657 ( .A(keyin[100]), .Y(n1386) );
  NBUFFX2_HVT U1658 ( .A(keyin[107]), .Y(n1383) );
  NBUFFX2_HVT U1659 ( .A(keyin[114]), .Y(n1446) );
  NBUFFX2_HVT U1660 ( .A(keyin[122]), .Y(n1431) );
  NBUFFX2_HVT U1661 ( .A(keyin[103]), .Y(n1385) );
  NBUFFX2_HVT U1662 ( .A(keyin[113]), .Y(n1376) );
  NBUFFX2_HVT U1663 ( .A(keyin[119]), .Y(n1370) );
  NBUFFX2_HVT U1664 ( .A(keyin[127]), .Y(n1364) );
  NBUFFX2_HVT U1665 ( .A(keyin[119]), .Y(n1369) );
  NBUFFX2_HVT U1666 ( .A(keyin[111]), .Y(n1377) );
  NBUFFX2_HVT U1667 ( .A(keyin[111]), .Y(n1378) );
  XOR2X1_HVT U1668 ( .A1(n1795), .A2(keyin[35]), .Y(n1840) );
  INVX0_HVT U1669 ( .A(n1791), .Y(n1482) );
  INVX0_HVT U1670 ( .A(n1792), .Y(n1483) );
  INVX0_HVT U1671 ( .A(n1790), .Y(n1485) );
  INVX0_HVT U1672 ( .A(round_num[1]), .Y(n1487) );
  INVX0_HVT U1673 ( .A(round_num[0]), .Y(n1488) );
  INVX0_HVT U1674 ( .A(round_num[3]), .Y(n1489) );
  INVX0_HVT U1675 ( .A(round_num[2]), .Y(n1490) );
  INVX0_HVT U1676 ( .A(n2256), .Y(n1497) );
  INVX0_HVT U1677 ( .A(n2253), .Y(n1498) );
  INVX0_HVT U1678 ( .A(n2245), .Y(n1499) );
  INVX0_HVT U1679 ( .A(n2244), .Y(n1500) );
  INVX0_HVT U1680 ( .A(n2235), .Y(n1501) );
  INVX0_HVT U1681 ( .A(n2105), .Y(n1502) );
  INVX0_HVT U1682 ( .A(n2071), .Y(n1503) );
  INVX0_HVT U1683 ( .A(n2274), .Y(n1504) );
  INVX0_HVT U1684 ( .A(n2260), .Y(n1505) );
  INVX0_HVT U1685 ( .A(n2272), .Y(n1506) );
  INVX0_HVT U1686 ( .A(n2273), .Y(n1507) );
  INVX0_HVT U1687 ( .A(n2269), .Y(n1508) );
  INVX0_HVT U1688 ( .A(n2268), .Y(n1509) );
  INVX0_HVT U1689 ( .A(n2267), .Y(n1510) );
  INVX0_HVT U1690 ( .A(n2266), .Y(n1511) );
  INVX0_HVT U1691 ( .A(n2265), .Y(n1512) );
  INVX0_HVT U1692 ( .A(n2264), .Y(n1513) );
  INVX0_HVT U1693 ( .A(n2261), .Y(n1514) );
  INVX0_HVT U1694 ( .A(n2259), .Y(n1515) );
  INVX0_HVT U1695 ( .A(n2258), .Y(n1516) );
  INVX0_HVT U1696 ( .A(n2257), .Y(n1517) );
  INVX0_HVT U1697 ( .A(n2255), .Y(n1518) );
  INVX0_HVT U1698 ( .A(n2254), .Y(n1519) );
  INVX0_HVT U1699 ( .A(n2251), .Y(n1520) );
  INVX0_HVT U1700 ( .A(n2250), .Y(n1521) );
  INVX0_HVT U1701 ( .A(n2248), .Y(n1523) );
  INVX0_HVT U1702 ( .A(n2064), .Y(n1524) );
  INVX0_HVT U1703 ( .A(n2247), .Y(n1525) );
  INVX0_HVT U1704 ( .A(n2246), .Y(n1526) );
  INVX0_HVT U1705 ( .A(n2243), .Y(n1527) );
  INVX0_HVT U1706 ( .A(n2242), .Y(n1528) );
  INVX0_HVT U1707 ( .A(n2241), .Y(n1529) );
  INVX0_HVT U1708 ( .A(n2240), .Y(n1530) );
  INVX0_HVT U1709 ( .A(n2239), .Y(n1531) );
  INVX0_HVT U1710 ( .A(n2238), .Y(n1532) );
  INVX0_HVT U1711 ( .A(n2237), .Y(n1533) );
  INVX0_HVT U1712 ( .A(n2206), .Y(n1534) );
  INVX0_HVT U1713 ( .A(n2263), .Y(n1535) );
  INVX0_HVT U1714 ( .A(n2218), .Y(n1536) );
  INVX0_HVT U1715 ( .A(n2163), .Y(n1537) );
  INVX0_HVT U1716 ( .A(n2070), .Y(n1538) );
  INVX0_HVT U1717 ( .A(n2123), .Y(n1539) );
  INVX0_HVT U1718 ( .A(n2069), .Y(n1540) );
  INVX0_HVT U1719 ( .A(n2068), .Y(n1541) );
  INVX0_HVT U1720 ( .A(n2066), .Y(n1543) );
  INVX0_HVT U1721 ( .A(n2065), .Y(n1544) );
  INVX0_HVT U1722 ( .A(n2183), .Y(n1545) );
  INVX0_HVT U1723 ( .A(n2177), .Y(n1546) );
  INVX0_HVT U1724 ( .A(n2063), .Y(n1547) );
  INVX0_HVT U1725 ( .A(n2062), .Y(n1548) );
  INVX0_HVT U1726 ( .A(n2061), .Y(n1549) );
  INVX0_HVT U1727 ( .A(n2059), .Y(n1551) );
  INVX0_HVT U1728 ( .A(n2473), .Y(n1565) );
  INVX0_HVT U1729 ( .A(n2470), .Y(n1566) );
  INVX0_HVT U1730 ( .A(n2462), .Y(n1567) );
  INVX0_HVT U1731 ( .A(n2461), .Y(n1568) );
  INVX0_HVT U1732 ( .A(n2452), .Y(n1569) );
  INVX0_HVT U1733 ( .A(n2324), .Y(n1570) );
  INVX0_HVT U1734 ( .A(n2290), .Y(n1571) );
  INVX0_HVT U1735 ( .A(n2491), .Y(n1572) );
  INVX0_HVT U1736 ( .A(n2477), .Y(n1573) );
  INVX0_HVT U1737 ( .A(n2489), .Y(n1574) );
  INVX0_HVT U1738 ( .A(n2490), .Y(n1575) );
  INVX0_HVT U1739 ( .A(n2486), .Y(n1576) );
  INVX0_HVT U1740 ( .A(n2485), .Y(n1577) );
  INVX0_HVT U1741 ( .A(n2484), .Y(n1578) );
  INVX0_HVT U1742 ( .A(n2482), .Y(n1580) );
  INVX0_HVT U1743 ( .A(n2481), .Y(n1581) );
  INVX0_HVT U1744 ( .A(n2478), .Y(n1582) );
  INVX0_HVT U1745 ( .A(n2476), .Y(n1583) );
  INVX0_HVT U1746 ( .A(n2475), .Y(n1584) );
  INVX0_HVT U1747 ( .A(n2474), .Y(n1585) );
  INVX0_HVT U1748 ( .A(n2472), .Y(n1586) );
  INVX0_HVT U1749 ( .A(n2471), .Y(n1587) );
  INVX0_HVT U1750 ( .A(n2468), .Y(n1588) );
  INVX0_HVT U1751 ( .A(n2467), .Y(n1589) );
  INVX0_HVT U1752 ( .A(n2466), .Y(n1590) );
  INVX0_HVT U1753 ( .A(n2465), .Y(n1591) );
  INVX0_HVT U1754 ( .A(n2464), .Y(n1593) );
  INVX0_HVT U1755 ( .A(n2463), .Y(n1594) );
  INVX0_HVT U1756 ( .A(n2460), .Y(n1595) );
  INVX0_HVT U1757 ( .A(n2459), .Y(n1596) );
  INVX0_HVT U1758 ( .A(n2458), .Y(n1597) );
  INVX0_HVT U1759 ( .A(n2457), .Y(n1598) );
  INVX0_HVT U1760 ( .A(n2455), .Y(n1599) );
  INVX0_HVT U1761 ( .A(n2454), .Y(n1600) );
  INVX0_HVT U1762 ( .A(n2423), .Y(n1601) );
  INVX0_HVT U1763 ( .A(n2480), .Y(n1602) );
  INVX0_HVT U1764 ( .A(n2435), .Y(n1603) );
  INVX0_HVT U1765 ( .A(n2381), .Y(n1604) );
  INVX0_HVT U1766 ( .A(n2289), .Y(n1605) );
  INVX0_HVT U1767 ( .A(n2339), .Y(n1606) );
  INVX0_HVT U1768 ( .A(n2288), .Y(n1607) );
  INVX0_HVT U1769 ( .A(n2287), .Y(n1608) );
  INVX0_HVT U1770 ( .A(n2285), .Y(n1610) );
  INVX0_HVT U1771 ( .A(n2284), .Y(n1611) );
  INVX0_HVT U1772 ( .A(n2401), .Y(n1612) );
  INVX0_HVT U1773 ( .A(n2395), .Y(n1613) );
  INVX0_HVT U1774 ( .A(n2282), .Y(n1614) );
  INVX0_HVT U1775 ( .A(n2281), .Y(n1615) );
  INVX0_HVT U1776 ( .A(n2280), .Y(n1616) );
  INVX0_HVT U1777 ( .A(n2279), .Y(n1617) );
  INVX0_HVT U1778 ( .A(n2278), .Y(n1618) );
  INVX0_HVT U1779 ( .A(n1408), .Y(n1624) );
  INVX0_HVT U1780 ( .A(n2694), .Y(n1628) );
  INVX0_HVT U1781 ( .A(n2691), .Y(n1629) );
  INVX0_HVT U1782 ( .A(n2683), .Y(n1630) );
  INVX0_HVT U1783 ( .A(n2682), .Y(n1631) );
  INVX0_HVT U1784 ( .A(n2673), .Y(n1632) );
  INVX0_HVT U1785 ( .A(n2541), .Y(n1633) );
  INVX0_HVT U1786 ( .A(n2507), .Y(n1634) );
  INVX0_HVT U1787 ( .A(n2712), .Y(n1635) );
  INVX0_HVT U1788 ( .A(n2698), .Y(n1636) );
  INVX0_HVT U1789 ( .A(n2710), .Y(n1637) );
  INVX0_HVT U1790 ( .A(n2711), .Y(n1638) );
  INVX0_HVT U1791 ( .A(n2707), .Y(n1639) );
  INVX0_HVT U1792 ( .A(n2706), .Y(n1640) );
  INVX0_HVT U1793 ( .A(n2705), .Y(n1641) );
  INVX0_HVT U1794 ( .A(n2704), .Y(n1642) );
  INVX0_HVT U1795 ( .A(n2703), .Y(n1643) );
  INVX0_HVT U1796 ( .A(n2702), .Y(n1644) );
  INVX0_HVT U1797 ( .A(n2699), .Y(n1645) );
  INVX0_HVT U1798 ( .A(n2697), .Y(n1646) );
  INVX0_HVT U1799 ( .A(n2696), .Y(n1647) );
  INVX0_HVT U1800 ( .A(n2695), .Y(n1648) );
  INVX0_HVT U1801 ( .A(n2692), .Y(n1650) );
  INVX0_HVT U1802 ( .A(n2689), .Y(n1651) );
  INVX0_HVT U1803 ( .A(n2688), .Y(n1652) );
  INVX0_HVT U1804 ( .A(n2687), .Y(n1653) );
  INVX0_HVT U1805 ( .A(n2686), .Y(n1654) );
  INVX0_HVT U1806 ( .A(n2500), .Y(n1655) );
  INVX0_HVT U1807 ( .A(n2685), .Y(n1656) );
  INVX0_HVT U1808 ( .A(n2684), .Y(n1657) );
  INVX0_HVT U1809 ( .A(n2681), .Y(n1658) );
  INVX0_HVT U1810 ( .A(n2680), .Y(n1659) );
  INVX0_HVT U1811 ( .A(n2679), .Y(n1660) );
  INVX0_HVT U1812 ( .A(n2678), .Y(n1661) );
  INVX0_HVT U1813 ( .A(n2677), .Y(n1662) );
  INVX0_HVT U1814 ( .A(n2676), .Y(n1663) );
  INVX0_HVT U1815 ( .A(n2675), .Y(n1664) );
  INVX0_HVT U1816 ( .A(n2644), .Y(n1665) );
  INVX0_HVT U1817 ( .A(n2701), .Y(n1666) );
  INVX0_HVT U1818 ( .A(n2656), .Y(n1667) );
  INVX0_HVT U1819 ( .A(n2601), .Y(n1668) );
  INVX0_HVT U1820 ( .A(n2506), .Y(n1669) );
  INVX0_HVT U1821 ( .A(n2559), .Y(n1670) );
  INVX0_HVT U1822 ( .A(n2505), .Y(n1671) );
  INVX0_HVT U1823 ( .A(n2504), .Y(n1672) );
  INVX0_HVT U1824 ( .A(n2503), .Y(n1673) );
  INVX0_HVT U1825 ( .A(n2502), .Y(n1674) );
  INVX0_HVT U1826 ( .A(n2501), .Y(n1675) );
  INVX0_HVT U1827 ( .A(n2621), .Y(n1676) );
  INVX0_HVT U1828 ( .A(n2615), .Y(n1677) );
  INVX0_HVT U1829 ( .A(n2499), .Y(n1678) );
  INVX0_HVT U1830 ( .A(n2497), .Y(n1680) );
  INVX0_HVT U1831 ( .A(n2496), .Y(n1681) );
  INVX0_HVT U1832 ( .A(n2495), .Y(n1682) );
  INVX0_HVT U1833 ( .A(n1416), .Y(n1688) );
  INVX0_HVT U1834 ( .A(n2054), .Y(n1697) );
  INVX0_HVT U1835 ( .A(n2037), .Y(n1698) );
  INVX0_HVT U1836 ( .A(n2035), .Y(n1699) );
  INVX0_HVT U1837 ( .A(n2026), .Y(n1700) );
  INVX0_HVT U1838 ( .A(n1890), .Y(n1701) );
  INVX0_HVT U1839 ( .A(n1853), .Y(n1702) );
  INVX0_HVT U1840 ( .A(n2056), .Y(n1703) );
  INVX0_HVT U1841 ( .A(n2043), .Y(n1704) );
  INVX0_HVT U1842 ( .A(n2052), .Y(n1705) );
  INVX0_HVT U1843 ( .A(n2053), .Y(n1706) );
  INVX0_HVT U1844 ( .A(n2050), .Y(n1707) );
  INVX0_HVT U1845 ( .A(n2049), .Y(n1708) );
  INVX0_HVT U1846 ( .A(n2048), .Y(n1709) );
  INVX0_HVT U1847 ( .A(n2047), .Y(n1710) );
  INVX0_HVT U1848 ( .A(n2044), .Y(n1711) );
  INVX0_HVT U1849 ( .A(n2042), .Y(n1712) );
  INVX0_HVT U1850 ( .A(n2041), .Y(n1713) );
  INVX0_HVT U1851 ( .A(n2040), .Y(n1714) );
  INVX0_HVT U1852 ( .A(n2039), .Y(n1715) );
  INVX0_HVT U1853 ( .A(n2038), .Y(n1716) );
  INVX0_HVT U1854 ( .A(n2036), .Y(n1717) );
  INVX0_HVT U1855 ( .A(n2034), .Y(n1718) );
  INVX0_HVT U1856 ( .A(n2031), .Y(n1719) );
  INVX0_HVT U1857 ( .A(n2030), .Y(n1720) );
  INVX0_HVT U1858 ( .A(n2029), .Y(n1721) );
  INVX0_HVT U1859 ( .A(n1846), .Y(n1722) );
  INVX0_HVT U1860 ( .A(n2028), .Y(n1723) );
  INVX0_HVT U1861 ( .A(n2027), .Y(n1724) );
  INVX0_HVT U1862 ( .A(n2025), .Y(n1725) );
  INVX0_HVT U1863 ( .A(n2024), .Y(n1726) );
  INVX0_HVT U1864 ( .A(n2023), .Y(n1727) );
  INVX0_HVT U1865 ( .A(n2022), .Y(n1728) );
  INVX0_HVT U1866 ( .A(n2021), .Y(n1729) );
  INVX0_HVT U1867 ( .A(n2020), .Y(n1730) );
  INVX0_HVT U1868 ( .A(n2019), .Y(n1731) );
  INVX0_HVT U1869 ( .A(n2018), .Y(n1732) );
  INVX0_HVT U1870 ( .A(n2015), .Y(n1733) );
  INVX0_HVT U1871 ( .A(n1986), .Y(n1734) );
  INVX0_HVT U1872 ( .A(n2046), .Y(n1735) );
  INVX0_HVT U1873 ( .A(n1946), .Y(n1736) );
  INVX0_HVT U1874 ( .A(n1852), .Y(n1737) );
  INVX0_HVT U1875 ( .A(n2003), .Y(n1738) );
  INVX0_HVT U1876 ( .A(n1905), .Y(n1739) );
  INVX0_HVT U1877 ( .A(n1851), .Y(n1740) );
  INVX0_HVT U1878 ( .A(n1850), .Y(n1741) );
  INVX0_HVT U1879 ( .A(n1849), .Y(n1742) );
  INVX0_HVT U1880 ( .A(n1848), .Y(n1743) );
  INVX0_HVT U1881 ( .A(n1847), .Y(n1744) );
  INVX0_HVT U1882 ( .A(n1965), .Y(n1745) );
  INVX0_HVT U1883 ( .A(n1955), .Y(n1746) );
  INVX0_HVT U1884 ( .A(n1845), .Y(n1747) );
  INVX0_HVT U1885 ( .A(n1844), .Y(n1748) );
  INVX0_HVT U1886 ( .A(n1843), .Y(n1749) );
  INVX0_HVT U1887 ( .A(n1842), .Y(n1750) );
  INVX0_HVT U1888 ( .A(n1841), .Y(n1751) );
  INVX0_HVT U1889 ( .A(n2055), .Y(n1756) );
endmodule

