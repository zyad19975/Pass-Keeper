
module aes ( plaintext, key, clk, reset, start, cipher_text, ready );
  input [127:0] plaintext;
  input [127:0] key;
  output [127:0] cipher_text;
  input clk, reset, start;
  output ready;
  wire   n4, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316;
  wire   [127:0] adk_out0;
  wire   [127:0] adk_in;
  wire   [3:0] round_number;
  wire   [127:0] key_round;
  wire   [127:0] keyout;

  add_round_keys_0 adk_0 ( .state(plaintext), .subkey(key), .out(adk_out0) );
  round r1 ( .in(adk_in), .round_num(round_number), .keyin(key_round), 
        .keyout(keyout), .out(cipher_text) );
  DFFX1_HVT \round_number_reg[0]  ( .D(n291), .CLK(clk), .Q(round_number[0]), 
        .QN(n292) );
  DFFX1_HVT d_reg ( .D(n289), .CLK(clk), .Q(n294), .QN(n4) );
  DFFX1_HVT \round_number_reg[3]  ( .D(n290), .CLK(clk), .Q(round_number[3])
         );
  DFFX1_HVT \round_number_reg[1]  ( .D(n288), .CLK(clk), .Q(round_number[1]), 
        .QN(n293) );
  DFFX1_HVT \round_number_reg[2]  ( .D(n287), .CLK(clk), .Q(round_number[2]), 
        .QN(n295) );
  DFFX1_HVT ready_reg ( .D(n30), .CLK(clk), .Q(ready) );
  DFFX1_HVT \adk_in_reg[0]  ( .D(n286), .CLK(clk), .Q(adk_in[0]) );
  DFFX1_HVT \adk_in_reg[1]  ( .D(n285), .CLK(clk), .Q(adk_in[1]) );
  DFFX1_HVT \adk_in_reg[2]  ( .D(n284), .CLK(clk), .Q(adk_in[2]) );
  DFFX1_HVT \adk_in_reg[3]  ( .D(n283), .CLK(clk), .Q(adk_in[3]) );
  DFFX1_HVT \adk_in_reg[4]  ( .D(n282), .CLK(clk), .Q(adk_in[4]) );
  DFFX1_HVT \adk_in_reg[5]  ( .D(n281), .CLK(clk), .Q(adk_in[5]) );
  DFFX1_HVT \adk_in_reg[6]  ( .D(n280), .CLK(clk), .Q(adk_in[6]) );
  DFFX1_HVT \adk_in_reg[7]  ( .D(n279), .CLK(clk), .Q(adk_in[7]) );
  DFFX1_HVT \adk_in_reg[8]  ( .D(n278), .CLK(clk), .Q(adk_in[8]) );
  DFFX1_HVT \adk_in_reg[9]  ( .D(n277), .CLK(clk), .Q(adk_in[9]) );
  DFFX1_HVT \adk_in_reg[10]  ( .D(n276), .CLK(clk), .Q(adk_in[10]) );
  DFFX1_HVT \adk_in_reg[11]  ( .D(n275), .CLK(clk), .Q(adk_in[11]) );
  DFFX1_HVT \adk_in_reg[12]  ( .D(n274), .CLK(clk), .Q(adk_in[12]) );
  DFFX1_HVT \adk_in_reg[13]  ( .D(n273), .CLK(clk), .Q(adk_in[13]) );
  DFFX1_HVT \adk_in_reg[14]  ( .D(n272), .CLK(clk), .Q(adk_in[14]) );
  DFFX1_HVT \adk_in_reg[15]  ( .D(n271), .CLK(clk), .Q(adk_in[15]) );
  DFFX1_HVT \adk_in_reg[16]  ( .D(n270), .CLK(clk), .Q(adk_in[16]) );
  DFFX1_HVT \adk_in_reg[17]  ( .D(n269), .CLK(clk), .Q(adk_in[17]) );
  DFFX1_HVT \adk_in_reg[18]  ( .D(n268), .CLK(clk), .Q(adk_in[18]) );
  DFFX1_HVT \adk_in_reg[19]  ( .D(n267), .CLK(clk), .Q(adk_in[19]) );
  DFFX1_HVT \adk_in_reg[20]  ( .D(n266), .CLK(clk), .Q(adk_in[20]) );
  DFFX1_HVT \adk_in_reg[21]  ( .D(n265), .CLK(clk), .Q(adk_in[21]) );
  DFFX1_HVT \adk_in_reg[22]  ( .D(n264), .CLK(clk), .Q(adk_in[22]) );
  DFFX1_HVT \adk_in_reg[23]  ( .D(n263), .CLK(clk), .Q(adk_in[23]) );
  DFFX1_HVT \adk_in_reg[24]  ( .D(n262), .CLK(clk), .Q(adk_in[24]) );
  DFFX1_HVT \adk_in_reg[25]  ( .D(n261), .CLK(clk), .Q(adk_in[25]) );
  DFFX1_HVT \adk_in_reg[26]  ( .D(n260), .CLK(clk), .Q(adk_in[26]) );
  DFFX1_HVT \adk_in_reg[27]  ( .D(n259), .CLK(clk), .Q(adk_in[27]) );
  DFFX1_HVT \adk_in_reg[28]  ( .D(n258), .CLK(clk), .Q(adk_in[28]) );
  DFFX1_HVT \adk_in_reg[29]  ( .D(n257), .CLK(clk), .Q(adk_in[29]) );
  DFFX1_HVT \adk_in_reg[30]  ( .D(n256), .CLK(clk), .Q(adk_in[30]) );
  DFFX1_HVT \adk_in_reg[31]  ( .D(n255), .CLK(clk), .Q(adk_in[31]) );
  DFFX1_HVT \adk_in_reg[32]  ( .D(n254), .CLK(clk), .Q(adk_in[32]) );
  DFFX1_HVT \adk_in_reg[33]  ( .D(n253), .CLK(clk), .Q(adk_in[33]) );
  DFFX1_HVT \adk_in_reg[34]  ( .D(n252), .CLK(clk), .Q(adk_in[34]) );
  DFFX1_HVT \adk_in_reg[35]  ( .D(n251), .CLK(clk), .Q(adk_in[35]) );
  DFFX1_HVT \adk_in_reg[36]  ( .D(n250), .CLK(clk), .Q(adk_in[36]) );
  DFFX1_HVT \adk_in_reg[37]  ( .D(n249), .CLK(clk), .Q(adk_in[37]) );
  DFFX1_HVT \adk_in_reg[38]  ( .D(n248), .CLK(clk), .Q(adk_in[38]) );
  DFFX1_HVT \adk_in_reg[39]  ( .D(n247), .CLK(clk), .Q(adk_in[39]) );
  DFFX1_HVT \adk_in_reg[40]  ( .D(n246), .CLK(clk), .Q(adk_in[40]) );
  DFFX1_HVT \adk_in_reg[41]  ( .D(n245), .CLK(clk), .Q(adk_in[41]) );
  DFFX1_HVT \adk_in_reg[42]  ( .D(n244), .CLK(clk), .Q(adk_in[42]) );
  DFFX1_HVT \adk_in_reg[43]  ( .D(n243), .CLK(clk), .Q(adk_in[43]) );
  DFFX1_HVT \adk_in_reg[44]  ( .D(n242), .CLK(clk), .Q(adk_in[44]) );
  DFFX1_HVT \adk_in_reg[45]  ( .D(n241), .CLK(clk), .Q(adk_in[45]) );
  DFFX1_HVT \adk_in_reg[46]  ( .D(n240), .CLK(clk), .Q(adk_in[46]) );
  DFFX1_HVT \adk_in_reg[47]  ( .D(n239), .CLK(clk), .Q(adk_in[47]) );
  DFFX1_HVT \adk_in_reg[48]  ( .D(n238), .CLK(clk), .Q(adk_in[48]) );
  DFFX1_HVT \adk_in_reg[49]  ( .D(n237), .CLK(clk), .Q(adk_in[49]) );
  DFFX1_HVT \adk_in_reg[50]  ( .D(n236), .CLK(clk), .Q(adk_in[50]) );
  DFFX1_HVT \adk_in_reg[51]  ( .D(n235), .CLK(clk), .Q(adk_in[51]) );
  DFFX1_HVT \adk_in_reg[52]  ( .D(n234), .CLK(clk), .Q(adk_in[52]) );
  DFFX1_HVT \adk_in_reg[53]  ( .D(n233), .CLK(clk), .Q(adk_in[53]) );
  DFFX1_HVT \adk_in_reg[54]  ( .D(n232), .CLK(clk), .Q(adk_in[54]) );
  DFFX1_HVT \adk_in_reg[55]  ( .D(n231), .CLK(clk), .Q(adk_in[55]) );
  DFFX1_HVT \adk_in_reg[56]  ( .D(n230), .CLK(clk), .Q(adk_in[56]) );
  DFFX1_HVT \adk_in_reg[57]  ( .D(n229), .CLK(clk), .Q(adk_in[57]) );
  DFFX1_HVT \adk_in_reg[58]  ( .D(n228), .CLK(clk), .Q(adk_in[58]) );
  DFFX1_HVT \adk_in_reg[59]  ( .D(n227), .CLK(clk), .Q(adk_in[59]) );
  DFFX1_HVT \adk_in_reg[60]  ( .D(n226), .CLK(clk), .Q(adk_in[60]) );
  DFFX1_HVT \adk_in_reg[61]  ( .D(n225), .CLK(clk), .Q(adk_in[61]) );
  DFFX1_HVT \adk_in_reg[62]  ( .D(n224), .CLK(clk), .Q(adk_in[62]) );
  DFFX1_HVT \adk_in_reg[63]  ( .D(n223), .CLK(clk), .Q(adk_in[63]) );
  DFFX1_HVT \adk_in_reg[64]  ( .D(n222), .CLK(clk), .Q(adk_in[64]) );
  DFFX1_HVT \adk_in_reg[65]  ( .D(n221), .CLK(clk), .Q(adk_in[65]) );
  DFFX1_HVT \adk_in_reg[66]  ( .D(n220), .CLK(clk), .Q(adk_in[66]) );
  DFFX1_HVT \adk_in_reg[67]  ( .D(n219), .CLK(clk), .Q(adk_in[67]) );
  DFFX1_HVT \adk_in_reg[68]  ( .D(n218), .CLK(clk), .Q(adk_in[68]) );
  DFFX1_HVT \adk_in_reg[69]  ( .D(n217), .CLK(clk), .Q(adk_in[69]) );
  DFFX1_HVT \adk_in_reg[70]  ( .D(n216), .CLK(clk), .Q(adk_in[70]) );
  DFFX1_HVT \adk_in_reg[71]  ( .D(n215), .CLK(clk), .Q(adk_in[71]) );
  DFFX1_HVT \adk_in_reg[72]  ( .D(n214), .CLK(clk), .Q(adk_in[72]) );
  DFFX1_HVT \adk_in_reg[73]  ( .D(n213), .CLK(clk), .Q(adk_in[73]) );
  DFFX1_HVT \adk_in_reg[74]  ( .D(n212), .CLK(clk), .Q(adk_in[74]) );
  DFFX1_HVT \adk_in_reg[75]  ( .D(n211), .CLK(clk), .Q(adk_in[75]) );
  DFFX1_HVT \adk_in_reg[76]  ( .D(n210), .CLK(clk), .Q(adk_in[76]) );
  DFFX1_HVT \adk_in_reg[77]  ( .D(n209), .CLK(clk), .Q(adk_in[77]) );
  DFFX1_HVT \adk_in_reg[78]  ( .D(n208), .CLK(clk), .Q(adk_in[78]) );
  DFFX1_HVT \adk_in_reg[79]  ( .D(n207), .CLK(clk), .Q(adk_in[79]) );
  DFFX1_HVT \adk_in_reg[80]  ( .D(n206), .CLK(clk), .Q(adk_in[80]) );
  DFFX1_HVT \adk_in_reg[81]  ( .D(n205), .CLK(clk), .Q(adk_in[81]) );
  DFFX1_HVT \adk_in_reg[82]  ( .D(n204), .CLK(clk), .Q(adk_in[82]) );
  DFFX1_HVT \adk_in_reg[83]  ( .D(n203), .CLK(clk), .Q(adk_in[83]) );
  DFFX1_HVT \adk_in_reg[84]  ( .D(n202), .CLK(clk), .Q(adk_in[84]) );
  DFFX1_HVT \adk_in_reg[85]  ( .D(n201), .CLK(clk), .Q(adk_in[85]) );
  DFFX1_HVT \adk_in_reg[86]  ( .D(n200), .CLK(clk), .Q(adk_in[86]) );
  DFFX1_HVT \adk_in_reg[87]  ( .D(n199), .CLK(clk), .Q(adk_in[87]) );
  DFFX1_HVT \adk_in_reg[88]  ( .D(n198), .CLK(clk), .Q(adk_in[88]) );
  DFFX1_HVT \adk_in_reg[89]  ( .D(n197), .CLK(clk), .Q(adk_in[89]) );
  DFFX1_HVT \adk_in_reg[90]  ( .D(n196), .CLK(clk), .Q(adk_in[90]) );
  DFFX1_HVT \adk_in_reg[91]  ( .D(n195), .CLK(clk), .Q(adk_in[91]) );
  DFFX1_HVT \adk_in_reg[92]  ( .D(n194), .CLK(clk), .Q(adk_in[92]) );
  DFFX1_HVT \adk_in_reg[93]  ( .D(n193), .CLK(clk), .Q(adk_in[93]) );
  DFFX1_HVT \adk_in_reg[94]  ( .D(n192), .CLK(clk), .Q(adk_in[94]) );
  DFFX1_HVT \adk_in_reg[95]  ( .D(n191), .CLK(clk), .Q(adk_in[95]) );
  DFFX1_HVT \adk_in_reg[96]  ( .D(n190), .CLK(clk), .Q(adk_in[96]) );
  DFFX1_HVT \adk_in_reg[97]  ( .D(n189), .CLK(clk), .Q(adk_in[97]) );
  DFFX1_HVT \adk_in_reg[98]  ( .D(n188), .CLK(clk), .Q(adk_in[98]) );
  DFFX1_HVT \adk_in_reg[99]  ( .D(n187), .CLK(clk), .Q(adk_in[99]) );
  DFFX1_HVT \adk_in_reg[100]  ( .D(n186), .CLK(clk), .Q(adk_in[100]) );
  DFFX1_HVT \adk_in_reg[101]  ( .D(n185), .CLK(clk), .Q(adk_in[101]) );
  DFFX1_HVT \adk_in_reg[102]  ( .D(n184), .CLK(clk), .Q(adk_in[102]) );
  DFFX1_HVT \adk_in_reg[103]  ( .D(n183), .CLK(clk), .Q(adk_in[103]) );
  DFFX1_HVT \adk_in_reg[104]  ( .D(n182), .CLK(clk), .Q(adk_in[104]) );
  DFFX1_HVT \adk_in_reg[105]  ( .D(n181), .CLK(clk), .Q(adk_in[105]) );
  DFFX1_HVT \adk_in_reg[106]  ( .D(n180), .CLK(clk), .Q(adk_in[106]) );
  DFFX1_HVT \adk_in_reg[107]  ( .D(n179), .CLK(clk), .Q(adk_in[107]) );
  DFFX1_HVT \adk_in_reg[108]  ( .D(n178), .CLK(clk), .Q(adk_in[108]) );
  DFFX1_HVT \adk_in_reg[109]  ( .D(n177), .CLK(clk), .Q(adk_in[109]) );
  DFFX1_HVT \adk_in_reg[110]  ( .D(n176), .CLK(clk), .Q(adk_in[110]) );
  DFFX1_HVT \adk_in_reg[111]  ( .D(n175), .CLK(clk), .Q(adk_in[111]) );
  DFFX1_HVT \adk_in_reg[112]  ( .D(n174), .CLK(clk), .Q(adk_in[112]) );
  DFFX1_HVT \adk_in_reg[113]  ( .D(n173), .CLK(clk), .Q(adk_in[113]) );
  DFFX1_HVT \adk_in_reg[114]  ( .D(n172), .CLK(clk), .Q(adk_in[114]) );
  DFFX1_HVT \adk_in_reg[115]  ( .D(n171), .CLK(clk), .Q(adk_in[115]) );
  DFFX1_HVT \adk_in_reg[116]  ( .D(n170), .CLK(clk), .Q(adk_in[116]) );
  DFFX1_HVT \adk_in_reg[117]  ( .D(n169), .CLK(clk), .Q(adk_in[117]) );
  DFFX1_HVT \adk_in_reg[118]  ( .D(n168), .CLK(clk), .Q(adk_in[118]) );
  DFFX1_HVT \adk_in_reg[119]  ( .D(n167), .CLK(clk), .Q(adk_in[119]) );
  DFFX1_HVT \adk_in_reg[120]  ( .D(n166), .CLK(clk), .Q(adk_in[120]) );
  DFFX1_HVT \adk_in_reg[121]  ( .D(n165), .CLK(clk), .Q(adk_in[121]) );
  DFFX1_HVT \adk_in_reg[122]  ( .D(n164), .CLK(clk), .Q(adk_in[122]) );
  DFFX1_HVT \adk_in_reg[123]  ( .D(n163), .CLK(clk), .Q(adk_in[123]) );
  DFFX1_HVT \adk_in_reg[124]  ( .D(n162), .CLK(clk), .Q(adk_in[124]) );
  DFFX1_HVT \adk_in_reg[125]  ( .D(n161), .CLK(clk), .Q(adk_in[125]) );
  DFFX1_HVT \adk_in_reg[126]  ( .D(n160), .CLK(clk), .Q(adk_in[126]) );
  DFFX1_HVT \adk_in_reg[127]  ( .D(n159), .CLK(clk), .Q(adk_in[127]) );
  DFFX1_HVT \key_round_reg[0]  ( .D(n158), .CLK(clk), .Q(key_round[0]) );
  DFFX1_HVT \key_round_reg[1]  ( .D(n157), .CLK(clk), .Q(key_round[1]) );
  DFFX1_HVT \key_round_reg[2]  ( .D(n156), .CLK(clk), .Q(key_round[2]) );
  DFFX1_HVT \key_round_reg[3]  ( .D(n155), .CLK(clk), .Q(key_round[3]) );
  DFFX1_HVT \key_round_reg[4]  ( .D(n154), .CLK(clk), .Q(key_round[4]) );
  DFFX1_HVT \key_round_reg[5]  ( .D(n153), .CLK(clk), .Q(key_round[5]) );
  DFFX1_HVT \key_round_reg[6]  ( .D(n152), .CLK(clk), .Q(key_round[6]) );
  DFFX1_HVT \key_round_reg[7]  ( .D(n151), .CLK(clk), .Q(key_round[7]) );
  DFFX1_HVT \key_round_reg[8]  ( .D(n150), .CLK(clk), .Q(key_round[8]) );
  DFFX1_HVT \key_round_reg[9]  ( .D(n149), .CLK(clk), .Q(key_round[9]) );
  DFFX1_HVT \key_round_reg[10]  ( .D(n148), .CLK(clk), .Q(key_round[10]) );
  DFFX1_HVT \key_round_reg[11]  ( .D(n147), .CLK(clk), .Q(key_round[11]) );
  DFFX1_HVT \key_round_reg[12]  ( .D(n146), .CLK(clk), .Q(key_round[12]) );
  DFFX1_HVT \key_round_reg[13]  ( .D(n145), .CLK(clk), .Q(key_round[13]) );
  DFFX1_HVT \key_round_reg[14]  ( .D(n144), .CLK(clk), .Q(key_round[14]) );
  DFFX1_HVT \key_round_reg[15]  ( .D(n143), .CLK(clk), .Q(key_round[15]) );
  DFFX1_HVT \key_round_reg[16]  ( .D(n142), .CLK(clk), .Q(key_round[16]) );
  DFFX1_HVT \key_round_reg[17]  ( .D(n141), .CLK(clk), .Q(key_round[17]) );
  DFFX1_HVT \key_round_reg[18]  ( .D(n140), .CLK(clk), .Q(key_round[18]) );
  DFFX1_HVT \key_round_reg[19]  ( .D(n139), .CLK(clk), .Q(key_round[19]) );
  DFFX1_HVT \key_round_reg[20]  ( .D(n138), .CLK(clk), .Q(key_round[20]) );
  DFFX1_HVT \key_round_reg[21]  ( .D(n137), .CLK(clk), .Q(key_round[21]) );
  DFFX1_HVT \key_round_reg[22]  ( .D(n136), .CLK(clk), .Q(key_round[22]) );
  DFFX1_HVT \key_round_reg[23]  ( .D(n135), .CLK(clk), .Q(key_round[23]) );
  DFFX1_HVT \key_round_reg[24]  ( .D(n134), .CLK(clk), .Q(key_round[24]) );
  DFFX1_HVT \key_round_reg[25]  ( .D(n133), .CLK(clk), .Q(key_round[25]) );
  DFFX1_HVT \key_round_reg[26]  ( .D(n132), .CLK(clk), .Q(key_round[26]) );
  DFFX1_HVT \key_round_reg[27]  ( .D(n131), .CLK(clk), .Q(key_round[27]) );
  DFFX1_HVT \key_round_reg[28]  ( .D(n130), .CLK(clk), .Q(key_round[28]) );
  DFFX1_HVT \key_round_reg[29]  ( .D(n129), .CLK(clk), .Q(key_round[29]) );
  DFFX1_HVT \key_round_reg[30]  ( .D(n128), .CLK(clk), .Q(key_round[30]) );
  DFFX1_HVT \key_round_reg[31]  ( .D(n127), .CLK(clk), .Q(key_round[31]) );
  DFFX1_HVT \key_round_reg[32]  ( .D(n126), .CLK(clk), .Q(key_round[32]) );
  DFFX1_HVT \key_round_reg[33]  ( .D(n125), .CLK(clk), .Q(key_round[33]) );
  DFFX1_HVT \key_round_reg[34]  ( .D(n124), .CLK(clk), .Q(key_round[34]) );
  DFFX1_HVT \key_round_reg[35]  ( .D(n123), .CLK(clk), .Q(key_round[35]) );
  DFFX1_HVT \key_round_reg[36]  ( .D(n122), .CLK(clk), .Q(key_round[36]) );
  DFFX1_HVT \key_round_reg[37]  ( .D(n121), .CLK(clk), .Q(key_round[37]) );
  DFFX1_HVT \key_round_reg[38]  ( .D(n120), .CLK(clk), .Q(key_round[38]) );
  DFFX1_HVT \key_round_reg[39]  ( .D(n119), .CLK(clk), .Q(key_round[39]) );
  DFFX1_HVT \key_round_reg[40]  ( .D(n118), .CLK(clk), .Q(key_round[40]) );
  DFFX1_HVT \key_round_reg[41]  ( .D(n117), .CLK(clk), .Q(key_round[41]) );
  DFFX1_HVT \key_round_reg[42]  ( .D(n116), .CLK(clk), .Q(key_round[42]) );
  DFFX1_HVT \key_round_reg[43]  ( .D(n115), .CLK(clk), .Q(key_round[43]) );
  DFFX1_HVT \key_round_reg[44]  ( .D(n114), .CLK(clk), .Q(key_round[44]) );
  DFFX1_HVT \key_round_reg[45]  ( .D(n113), .CLK(clk), .Q(key_round[45]) );
  DFFX1_HVT \key_round_reg[46]  ( .D(n112), .CLK(clk), .Q(key_round[46]) );
  DFFX1_HVT \key_round_reg[47]  ( .D(n111), .CLK(clk), .Q(key_round[47]) );
  DFFX1_HVT \key_round_reg[48]  ( .D(n110), .CLK(clk), .Q(key_round[48]) );
  DFFX1_HVT \key_round_reg[49]  ( .D(n109), .CLK(clk), .Q(key_round[49]) );
  DFFX1_HVT \key_round_reg[50]  ( .D(n108), .CLK(clk), .Q(key_round[50]) );
  DFFX1_HVT \key_round_reg[51]  ( .D(n107), .CLK(clk), .Q(key_round[51]) );
  DFFX1_HVT \key_round_reg[52]  ( .D(n106), .CLK(clk), .Q(key_round[52]) );
  DFFX1_HVT \key_round_reg[53]  ( .D(n105), .CLK(clk), .Q(key_round[53]) );
  DFFX1_HVT \key_round_reg[54]  ( .D(n104), .CLK(clk), .Q(key_round[54]) );
  DFFX1_HVT \key_round_reg[55]  ( .D(n103), .CLK(clk), .Q(key_round[55]) );
  DFFX1_HVT \key_round_reg[56]  ( .D(n102), .CLK(clk), .Q(key_round[56]) );
  DFFX1_HVT \key_round_reg[57]  ( .D(n101), .CLK(clk), .Q(key_round[57]) );
  DFFX1_HVT \key_round_reg[58]  ( .D(n100), .CLK(clk), .Q(key_round[58]) );
  DFFX1_HVT \key_round_reg[59]  ( .D(n99), .CLK(clk), .Q(key_round[59]) );
  DFFX1_HVT \key_round_reg[60]  ( .D(n98), .CLK(clk), .Q(key_round[60]) );
  DFFX1_HVT \key_round_reg[61]  ( .D(n97), .CLK(clk), .Q(key_round[61]) );
  DFFX1_HVT \key_round_reg[62]  ( .D(n96), .CLK(clk), .Q(key_round[62]) );
  DFFX1_HVT \key_round_reg[63]  ( .D(n95), .CLK(clk), .Q(key_round[63]) );
  DFFX1_HVT \key_round_reg[64]  ( .D(n94), .CLK(clk), .Q(key_round[64]) );
  DFFX1_HVT \key_round_reg[65]  ( .D(n93), .CLK(clk), .Q(key_round[65]) );
  DFFX1_HVT \key_round_reg[66]  ( .D(n92), .CLK(clk), .Q(key_round[66]) );
  DFFX1_HVT \key_round_reg[67]  ( .D(n91), .CLK(clk), .Q(key_round[67]) );
  DFFX1_HVT \key_round_reg[68]  ( .D(n90), .CLK(clk), .Q(key_round[68]) );
  DFFX1_HVT \key_round_reg[69]  ( .D(n89), .CLK(clk), .Q(key_round[69]) );
  DFFX1_HVT \key_round_reg[70]  ( .D(n88), .CLK(clk), .Q(key_round[70]) );
  DFFX1_HVT \key_round_reg[71]  ( .D(n87), .CLK(clk), .Q(key_round[71]) );
  DFFX1_HVT \key_round_reg[72]  ( .D(n86), .CLK(clk), .Q(key_round[72]) );
  DFFX1_HVT \key_round_reg[73]  ( .D(n85), .CLK(clk), .Q(key_round[73]) );
  DFFX1_HVT \key_round_reg[74]  ( .D(n84), .CLK(clk), .Q(key_round[74]) );
  DFFX1_HVT \key_round_reg[75]  ( .D(n83), .CLK(clk), .Q(key_round[75]) );
  DFFX1_HVT \key_round_reg[76]  ( .D(n82), .CLK(clk), .Q(key_round[76]) );
  DFFX1_HVT \key_round_reg[77]  ( .D(n81), .CLK(clk), .Q(key_round[77]) );
  DFFX1_HVT \key_round_reg[78]  ( .D(n80), .CLK(clk), .Q(key_round[78]) );
  DFFX1_HVT \key_round_reg[79]  ( .D(n79), .CLK(clk), .Q(key_round[79]) );
  DFFX1_HVT \key_round_reg[80]  ( .D(n78), .CLK(clk), .Q(key_round[80]) );
  DFFX1_HVT \key_round_reg[81]  ( .D(n77), .CLK(clk), .Q(key_round[81]) );
  DFFX1_HVT \key_round_reg[82]  ( .D(n76), .CLK(clk), .Q(key_round[82]) );
  DFFX1_HVT \key_round_reg[83]  ( .D(n75), .CLK(clk), .Q(key_round[83]) );
  DFFX1_HVT \key_round_reg[84]  ( .D(n74), .CLK(clk), .Q(key_round[84]) );
  DFFX1_HVT \key_round_reg[85]  ( .D(n73), .CLK(clk), .Q(key_round[85]) );
  DFFX1_HVT \key_round_reg[86]  ( .D(n72), .CLK(clk), .Q(key_round[86]) );
  DFFX1_HVT \key_round_reg[87]  ( .D(n71), .CLK(clk), .Q(key_round[87]) );
  DFFX1_HVT \key_round_reg[88]  ( .D(n70), .CLK(clk), .Q(key_round[88]) );
  DFFX1_HVT \key_round_reg[89]  ( .D(n69), .CLK(clk), .Q(key_round[89]) );
  DFFX1_HVT \key_round_reg[90]  ( .D(n68), .CLK(clk), .Q(key_round[90]) );
  DFFX1_HVT \key_round_reg[91]  ( .D(n67), .CLK(clk), .Q(key_round[91]) );
  DFFX1_HVT \key_round_reg[92]  ( .D(n66), .CLK(clk), .Q(key_round[92]) );
  DFFX1_HVT \key_round_reg[93]  ( .D(n65), .CLK(clk), .Q(key_round[93]) );
  DFFX1_HVT \key_round_reg[94]  ( .D(n64), .CLK(clk), .Q(key_round[94]) );
  DFFX1_HVT \key_round_reg[95]  ( .D(n63), .CLK(clk), .Q(key_round[95]) );
  DFFX1_HVT \key_round_reg[96]  ( .D(n62), .CLK(clk), .Q(key_round[96]) );
  DFFX1_HVT \key_round_reg[97]  ( .D(n61), .CLK(clk), .Q(key_round[97]) );
  DFFX1_HVT \key_round_reg[98]  ( .D(n60), .CLK(clk), .Q(key_round[98]) );
  DFFX1_HVT \key_round_reg[99]  ( .D(n59), .CLK(clk), .Q(key_round[99]) );
  DFFX1_HVT \key_round_reg[100]  ( .D(n58), .CLK(clk), .Q(key_round[100]) );
  DFFX1_HVT \key_round_reg[101]  ( .D(n57), .CLK(clk), .Q(key_round[101]) );
  DFFX1_HVT \key_round_reg[102]  ( .D(n56), .CLK(clk), .Q(key_round[102]) );
  DFFX1_HVT \key_round_reg[103]  ( .D(n55), .CLK(clk), .Q(key_round[103]) );
  DFFX1_HVT \key_round_reg[104]  ( .D(n54), .CLK(clk), .Q(key_round[104]) );
  DFFX1_HVT \key_round_reg[105]  ( .D(n53), .CLK(clk), .Q(key_round[105]) );
  DFFX1_HVT \key_round_reg[106]  ( .D(n52), .CLK(clk), .Q(key_round[106]) );
  DFFX1_HVT \key_round_reg[107]  ( .D(n51), .CLK(clk), .Q(key_round[107]) );
  DFFX1_HVT \key_round_reg[108]  ( .D(n50), .CLK(clk), .Q(key_round[108]) );
  DFFX1_HVT \key_round_reg[109]  ( .D(n49), .CLK(clk), .Q(key_round[109]) );
  DFFX1_HVT \key_round_reg[110]  ( .D(n48), .CLK(clk), .Q(key_round[110]) );
  DFFX1_HVT \key_round_reg[111]  ( .D(n47), .CLK(clk), .Q(key_round[111]) );
  DFFX1_HVT \key_round_reg[112]  ( .D(n46), .CLK(clk), .Q(key_round[112]) );
  DFFX1_HVT \key_round_reg[113]  ( .D(n45), .CLK(clk), .Q(key_round[113]) );
  DFFX1_HVT \key_round_reg[114]  ( .D(n44), .CLK(clk), .Q(key_round[114]) );
  DFFX1_HVT \key_round_reg[115]  ( .D(n43), .CLK(clk), .Q(key_round[115]) );
  DFFX1_HVT \key_round_reg[116]  ( .D(n42), .CLK(clk), .Q(key_round[116]) );
  DFFX1_HVT \key_round_reg[117]  ( .D(n41), .CLK(clk), .Q(key_round[117]) );
  DFFX1_HVT \key_round_reg[118]  ( .D(n40), .CLK(clk), .Q(key_round[118]) );
  DFFX1_HVT \key_round_reg[119]  ( .D(n39), .CLK(clk), .Q(key_round[119]) );
  DFFX1_HVT \key_round_reg[120]  ( .D(n38), .CLK(clk), .Q(key_round[120]) );
  DFFX1_HVT \key_round_reg[121]  ( .D(n37), .CLK(clk), .Q(key_round[121]) );
  DFFX1_HVT \key_round_reg[122]  ( .D(n36), .CLK(clk), .Q(key_round[122]) );
  DFFX1_HVT \key_round_reg[123]  ( .D(n35), .CLK(clk), .Q(key_round[123]) );
  DFFX1_HVT \key_round_reg[124]  ( .D(n34), .CLK(clk), .Q(key_round[124]) );
  DFFX1_HVT \key_round_reg[125]  ( .D(n33), .CLK(clk), .Q(key_round[125]) );
  DFFX1_HVT \key_round_reg[126]  ( .D(n32), .CLK(clk), .Q(key_round[126]) );
  DFFX1_HVT \key_round_reg[127]  ( .D(n31), .CLK(clk), .Q(key_round[127]) );
  AO222X1_HVT U288 ( .A1(key[59]), .A2(n296), .A3(n297), .A4(key_round[59]), 
        .A5(keyout[59]), .A6(n298), .Y(n99) );
  AO222X1_HVT U289 ( .A1(key[60]), .A2(n296), .A3(n297), .A4(key_round[60]), 
        .A5(keyout[60]), .A6(n298), .Y(n98) );
  AO222X1_HVT U290 ( .A1(key[61]), .A2(n296), .A3(n297), .A4(key_round[61]), 
        .A5(keyout[61]), .A6(n298), .Y(n97) );
  AO222X1_HVT U291 ( .A1(key[62]), .A2(n296), .A3(n297), .A4(key_round[62]), 
        .A5(keyout[62]), .A6(n298), .Y(n96) );
  AO222X1_HVT U292 ( .A1(key[63]), .A2(n296), .A3(n297), .A4(key_round[63]), 
        .A5(keyout[63]), .A6(n298), .Y(n95) );
  AO222X1_HVT U293 ( .A1(key[64]), .A2(n296), .A3(n297), .A4(key_round[64]), 
        .A5(keyout[64]), .A6(n298), .Y(n94) );
  AO222X1_HVT U294 ( .A1(key[65]), .A2(n296), .A3(n297), .A4(key_round[65]), 
        .A5(keyout[65]), .A6(n298), .Y(n93) );
  AO222X1_HVT U295 ( .A1(key[66]), .A2(n296), .A3(n297), .A4(key_round[66]), 
        .A5(keyout[66]), .A6(n298), .Y(n92) );
  AO222X1_HVT U296 ( .A1(key[67]), .A2(n296), .A3(n297), .A4(key_round[67]), 
        .A5(keyout[67]), .A6(n298), .Y(n91) );
  AO222X1_HVT U297 ( .A1(key[68]), .A2(n296), .A3(n297), .A4(key_round[68]), 
        .A5(keyout[68]), .A6(n298), .Y(n90) );
  AO222X1_HVT U298 ( .A1(key[69]), .A2(n296), .A3(n297), .A4(key_round[69]), 
        .A5(keyout[69]), .A6(n298), .Y(n89) );
  AO222X1_HVT U299 ( .A1(key[70]), .A2(n296), .A3(n297), .A4(key_round[70]), 
        .A5(keyout[70]), .A6(n298), .Y(n88) );
  AO222X1_HVT U300 ( .A1(key[71]), .A2(n296), .A3(n297), .A4(key_round[71]), 
        .A5(keyout[71]), .A6(n298), .Y(n87) );
  AO222X1_HVT U301 ( .A1(key[72]), .A2(n296), .A3(n297), .A4(key_round[72]), 
        .A5(keyout[72]), .A6(n298), .Y(n86) );
  AO222X1_HVT U302 ( .A1(key[73]), .A2(n296), .A3(n297), .A4(key_round[73]), 
        .A5(keyout[73]), .A6(n298), .Y(n85) );
  AO222X1_HVT U303 ( .A1(key[74]), .A2(n296), .A3(n297), .A4(key_round[74]), 
        .A5(keyout[74]), .A6(n298), .Y(n84) );
  AO222X1_HVT U304 ( .A1(key[75]), .A2(n296), .A3(n297), .A4(key_round[75]), 
        .A5(keyout[75]), .A6(n298), .Y(n83) );
  AO222X1_HVT U305 ( .A1(key[76]), .A2(n296), .A3(n297), .A4(key_round[76]), 
        .A5(keyout[76]), .A6(n298), .Y(n82) );
  AO222X1_HVT U306 ( .A1(key[77]), .A2(n296), .A3(n297), .A4(key_round[77]), 
        .A5(keyout[77]), .A6(n298), .Y(n81) );
  AO222X1_HVT U307 ( .A1(key[78]), .A2(n296), .A3(n297), .A4(key_round[78]), 
        .A5(keyout[78]), .A6(n298), .Y(n80) );
  AO222X1_HVT U308 ( .A1(key[79]), .A2(n296), .A3(n297), .A4(key_round[79]), 
        .A5(keyout[79]), .A6(n298), .Y(n79) );
  AO222X1_HVT U309 ( .A1(key[80]), .A2(n296), .A3(n297), .A4(key_round[80]), 
        .A5(keyout[80]), .A6(n298), .Y(n78) );
  AO222X1_HVT U310 ( .A1(key[81]), .A2(n296), .A3(n297), .A4(key_round[81]), 
        .A5(keyout[81]), .A6(n298), .Y(n77) );
  AO222X1_HVT U311 ( .A1(key[82]), .A2(n296), .A3(n297), .A4(key_round[82]), 
        .A5(keyout[82]), .A6(n298), .Y(n76) );
  AO222X1_HVT U312 ( .A1(key[83]), .A2(n296), .A3(n297), .A4(key_round[83]), 
        .A5(keyout[83]), .A6(n298), .Y(n75) );
  AO222X1_HVT U313 ( .A1(key[84]), .A2(n296), .A3(n297), .A4(key_round[84]), 
        .A5(keyout[84]), .A6(n298), .Y(n74) );
  AO222X1_HVT U314 ( .A1(key[85]), .A2(n296), .A3(n297), .A4(key_round[85]), 
        .A5(keyout[85]), .A6(n298), .Y(n73) );
  AO222X1_HVT U315 ( .A1(key[86]), .A2(n296), .A3(n297), .A4(key_round[86]), 
        .A5(keyout[86]), .A6(n298), .Y(n72) );
  AO222X1_HVT U316 ( .A1(key[87]), .A2(n296), .A3(n297), .A4(key_round[87]), 
        .A5(keyout[87]), .A6(n298), .Y(n71) );
  AO222X1_HVT U317 ( .A1(key[88]), .A2(n296), .A3(n297), .A4(key_round[88]), 
        .A5(keyout[88]), .A6(n298), .Y(n70) );
  AO222X1_HVT U318 ( .A1(key[89]), .A2(n296), .A3(n297), .A4(key_round[89]), 
        .A5(keyout[89]), .A6(n298), .Y(n69) );
  AO222X1_HVT U319 ( .A1(key[90]), .A2(n296), .A3(n297), .A4(key_round[90]), 
        .A5(keyout[90]), .A6(n298), .Y(n68) );
  AO222X1_HVT U320 ( .A1(key[91]), .A2(n296), .A3(n297), .A4(key_round[91]), 
        .A5(keyout[91]), .A6(n298), .Y(n67) );
  AO222X1_HVT U321 ( .A1(key[92]), .A2(n296), .A3(n297), .A4(key_round[92]), 
        .A5(keyout[92]), .A6(n298), .Y(n66) );
  AO222X1_HVT U322 ( .A1(key[93]), .A2(n296), .A3(n297), .A4(key_round[93]), 
        .A5(keyout[93]), .A6(n298), .Y(n65) );
  AO222X1_HVT U323 ( .A1(key[94]), .A2(n296), .A3(n297), .A4(key_round[94]), 
        .A5(keyout[94]), .A6(n298), .Y(n64) );
  AO222X1_HVT U324 ( .A1(key[95]), .A2(n296), .A3(n297), .A4(key_round[95]), 
        .A5(keyout[95]), .A6(n298), .Y(n63) );
  AO222X1_HVT U325 ( .A1(key[96]), .A2(n296), .A3(n297), .A4(key_round[96]), 
        .A5(keyout[96]), .A6(n298), .Y(n62) );
  AO222X1_HVT U326 ( .A1(key[97]), .A2(n296), .A3(n297), .A4(key_round[97]), 
        .A5(keyout[97]), .A6(n298), .Y(n61) );
  AO222X1_HVT U327 ( .A1(key[98]), .A2(n296), .A3(n297), .A4(key_round[98]), 
        .A5(keyout[98]), .A6(n298), .Y(n60) );
  AO222X1_HVT U328 ( .A1(key[99]), .A2(n296), .A3(n297), .A4(key_round[99]), 
        .A5(keyout[99]), .A6(n298), .Y(n59) );
  AO222X1_HVT U329 ( .A1(key[100]), .A2(n296), .A3(n297), .A4(key_round[100]), 
        .A5(keyout[100]), .A6(n298), .Y(n58) );
  AO222X1_HVT U330 ( .A1(key[101]), .A2(n296), .A3(n297), .A4(key_round[101]), 
        .A5(keyout[101]), .A6(n298), .Y(n57) );
  AO222X1_HVT U331 ( .A1(key[102]), .A2(n296), .A3(n297), .A4(key_round[102]), 
        .A5(keyout[102]), .A6(n298), .Y(n56) );
  AO222X1_HVT U332 ( .A1(key[103]), .A2(n296), .A3(n297), .A4(key_round[103]), 
        .A5(keyout[103]), .A6(n298), .Y(n55) );
  AO222X1_HVT U333 ( .A1(key[104]), .A2(n296), .A3(n297), .A4(key_round[104]), 
        .A5(keyout[104]), .A6(n298), .Y(n54) );
  AO222X1_HVT U334 ( .A1(key[105]), .A2(n296), .A3(n297), .A4(key_round[105]), 
        .A5(keyout[105]), .A6(n298), .Y(n53) );
  AO222X1_HVT U335 ( .A1(key[106]), .A2(n296), .A3(n297), .A4(key_round[106]), 
        .A5(keyout[106]), .A6(n298), .Y(n52) );
  AO222X1_HVT U336 ( .A1(key[107]), .A2(n296), .A3(n297), .A4(key_round[107]), 
        .A5(keyout[107]), .A6(n298), .Y(n51) );
  AO222X1_HVT U337 ( .A1(key[108]), .A2(n296), .A3(n297), .A4(key_round[108]), 
        .A5(keyout[108]), .A6(n298), .Y(n50) );
  AO222X1_HVT U338 ( .A1(key[109]), .A2(n296), .A3(n297), .A4(key_round[109]), 
        .A5(keyout[109]), .A6(n298), .Y(n49) );
  AO222X1_HVT U339 ( .A1(key[110]), .A2(n296), .A3(n297), .A4(key_round[110]), 
        .A5(keyout[110]), .A6(n298), .Y(n48) );
  AO222X1_HVT U340 ( .A1(key[111]), .A2(n296), .A3(n297), .A4(key_round[111]), 
        .A5(keyout[111]), .A6(n298), .Y(n47) );
  AO222X1_HVT U341 ( .A1(key[112]), .A2(n296), .A3(n297), .A4(key_round[112]), 
        .A5(keyout[112]), .A6(n298), .Y(n46) );
  AO222X1_HVT U342 ( .A1(key[113]), .A2(n296), .A3(n297), .A4(key_round[113]), 
        .A5(keyout[113]), .A6(n298), .Y(n45) );
  AO222X1_HVT U343 ( .A1(key[114]), .A2(n296), .A3(n297), .A4(key_round[114]), 
        .A5(keyout[114]), .A6(n298), .Y(n44) );
  AO222X1_HVT U344 ( .A1(key[115]), .A2(n296), .A3(n297), .A4(key_round[115]), 
        .A5(keyout[115]), .A6(n298), .Y(n43) );
  AO222X1_HVT U345 ( .A1(key[116]), .A2(n296), .A3(n297), .A4(key_round[116]), 
        .A5(keyout[116]), .A6(n298), .Y(n42) );
  AO222X1_HVT U346 ( .A1(key[117]), .A2(n296), .A3(n297), .A4(key_round[117]), 
        .A5(keyout[117]), .A6(n298), .Y(n41) );
  AO222X1_HVT U347 ( .A1(key[118]), .A2(n296), .A3(n297), .A4(key_round[118]), 
        .A5(keyout[118]), .A6(n298), .Y(n40) );
  AO222X1_HVT U348 ( .A1(key[119]), .A2(n296), .A3(n297), .A4(key_round[119]), 
        .A5(keyout[119]), .A6(n298), .Y(n39) );
  AO222X1_HVT U349 ( .A1(key[120]), .A2(n296), .A3(n297), .A4(key_round[120]), 
        .A5(keyout[120]), .A6(n298), .Y(n38) );
  AO222X1_HVT U350 ( .A1(key[121]), .A2(n296), .A3(n297), .A4(key_round[121]), 
        .A5(keyout[121]), .A6(n298), .Y(n37) );
  AO222X1_HVT U351 ( .A1(key[122]), .A2(n296), .A3(n297), .A4(key_round[122]), 
        .A5(keyout[122]), .A6(n298), .Y(n36) );
  AO222X1_HVT U352 ( .A1(key[123]), .A2(n296), .A3(n297), .A4(key_round[123]), 
        .A5(keyout[123]), .A6(n298), .Y(n35) );
  AO222X1_HVT U353 ( .A1(key[124]), .A2(n296), .A3(n297), .A4(key_round[124]), 
        .A5(keyout[124]), .A6(n298), .Y(n34) );
  AO222X1_HVT U354 ( .A1(key[125]), .A2(n296), .A3(n297), .A4(key_round[125]), 
        .A5(keyout[125]), .A6(n298), .Y(n33) );
  AO222X1_HVT U355 ( .A1(key[126]), .A2(n296), .A3(n297), .A4(key_round[126]), 
        .A5(keyout[126]), .A6(n298), .Y(n32) );
  AO222X1_HVT U356 ( .A1(key[127]), .A2(n296), .A3(n297), .A4(key_round[127]), 
        .A5(keyout[127]), .A6(n298), .Y(n31) );
  OA21X1_HVT U357 ( .A1(n299), .A2(n300), .A3(n301), .Y(n30) );
  INVX0_HVT U358 ( .A(n302), .Y(n300) );
  AND2X1_HVT U359 ( .A1(ready), .A2(n303), .Y(n299) );
  MUX21X1_HVT U360 ( .A1(n304), .A2(n305), .S0(round_number[0]), .Y(n291) );
  AND2X1_HVT U361 ( .A1(n297), .A2(n306), .Y(n305) );
  AO22X1_HVT U362 ( .A1(round_number[3]), .A2(n307), .A3(round_number[2]), 
        .A4(n308), .Y(n290) );
  NAND3X0_HVT U363 ( .A1(n302), .A2(n301), .A3(n309), .Y(n289) );
  NAND2X0_HVT U364 ( .A1(n306), .A2(n294), .Y(n309) );
  NAND4X0_HVT U365 ( .A1(n292), .A2(n295), .A3(round_number[3]), .A4(n310), 
        .Y(n302) );
  AND2X1_HVT U366 ( .A1(round_number[1]), .A2(n4), .Y(n310) );
  MUX21X1_HVT U367 ( .A1(n311), .A2(n312), .S0(round_number[1]), .Y(n288) );
  AND2X1_HVT U368 ( .A1(round_number[0]), .A2(n304), .Y(n311) );
  MUX21X1_HVT U369 ( .A1(n308), .A2(n307), .S0(round_number[2]), .Y(n287) );
  AO21X1_HVT U370 ( .A1(n304), .A2(n293), .A3(n312), .Y(n307) );
  AO22X1_HVT U371 ( .A1(n304), .A2(n292), .A3(n297), .A4(n306), .Y(n312) );
  NAND2X0_HVT U372 ( .A1(start), .A2(n313), .Y(n306) );
  INVX0_HVT U373 ( .A(n303), .Y(n313) );
  NAND3X0_HVT U374 ( .A1(n314), .A2(n294), .A3(round_number[3]), .Y(n303) );
  AND3X1_HVT U375 ( .A1(round_number[1]), .A2(n304), .A3(round_number[0]), .Y(
        n308) );
  AO222X1_HVT U376 ( .A1(adk_out0[0]), .A2(n296), .A3(n297), .A4(adk_in[0]), 
        .A5(cipher_text[0]), .A6(n298), .Y(n286) );
  AO222X1_HVT U377 ( .A1(adk_out0[1]), .A2(n296), .A3(n297), .A4(adk_in[1]), 
        .A5(cipher_text[1]), .A6(n298), .Y(n285) );
  AO222X1_HVT U378 ( .A1(adk_out0[2]), .A2(n296), .A3(n297), .A4(adk_in[2]), 
        .A5(cipher_text[2]), .A6(n298), .Y(n284) );
  AO222X1_HVT U379 ( .A1(adk_out0[3]), .A2(n296), .A3(n297), .A4(adk_in[3]), 
        .A5(cipher_text[3]), .A6(n298), .Y(n283) );
  AO222X1_HVT U380 ( .A1(adk_out0[4]), .A2(n296), .A3(n297), .A4(adk_in[4]), 
        .A5(cipher_text[4]), .A6(n298), .Y(n282) );
  AO222X1_HVT U381 ( .A1(adk_out0[5]), .A2(n296), .A3(n297), .A4(adk_in[5]), 
        .A5(cipher_text[5]), .A6(n298), .Y(n281) );
  AO222X1_HVT U382 ( .A1(adk_out0[6]), .A2(n296), .A3(n297), .A4(adk_in[6]), 
        .A5(cipher_text[6]), .A6(n298), .Y(n280) );
  AO222X1_HVT U383 ( .A1(adk_out0[7]), .A2(n296), .A3(n297), .A4(adk_in[7]), 
        .A5(cipher_text[7]), .A6(n298), .Y(n279) );
  AO222X1_HVT U384 ( .A1(adk_out0[8]), .A2(n296), .A3(n297), .A4(adk_in[8]), 
        .A5(cipher_text[8]), .A6(n298), .Y(n278) );
  AO222X1_HVT U385 ( .A1(adk_out0[9]), .A2(n296), .A3(n297), .A4(adk_in[9]), 
        .A5(cipher_text[9]), .A6(n298), .Y(n277) );
  AO222X1_HVT U386 ( .A1(adk_out0[10]), .A2(n296), .A3(n297), .A4(adk_in[10]), 
        .A5(cipher_text[10]), .A6(n298), .Y(n276) );
  AO222X1_HVT U387 ( .A1(adk_out0[11]), .A2(n296), .A3(n297), .A4(adk_in[11]), 
        .A5(cipher_text[11]), .A6(n298), .Y(n275) );
  AO222X1_HVT U388 ( .A1(adk_out0[12]), .A2(n296), .A3(n297), .A4(adk_in[12]), 
        .A5(cipher_text[12]), .A6(n298), .Y(n274) );
  AO222X1_HVT U389 ( .A1(adk_out0[13]), .A2(n296), .A3(n297), .A4(adk_in[13]), 
        .A5(cipher_text[13]), .A6(n298), .Y(n273) );
  AO222X1_HVT U390 ( .A1(adk_out0[14]), .A2(n296), .A3(n297), .A4(adk_in[14]), 
        .A5(cipher_text[14]), .A6(n298), .Y(n272) );
  AO222X1_HVT U391 ( .A1(adk_out0[15]), .A2(n296), .A3(n297), .A4(adk_in[15]), 
        .A5(cipher_text[15]), .A6(n298), .Y(n271) );
  AO222X1_HVT U392 ( .A1(adk_out0[16]), .A2(n296), .A3(n297), .A4(adk_in[16]), 
        .A5(cipher_text[16]), .A6(n298), .Y(n270) );
  AO222X1_HVT U393 ( .A1(adk_out0[17]), .A2(n296), .A3(n297), .A4(adk_in[17]), 
        .A5(cipher_text[17]), .A6(n298), .Y(n269) );
  AO222X1_HVT U394 ( .A1(adk_out0[18]), .A2(n296), .A3(n297), .A4(adk_in[18]), 
        .A5(cipher_text[18]), .A6(n298), .Y(n268) );
  AO222X1_HVT U395 ( .A1(adk_out0[19]), .A2(n296), .A3(n297), .A4(adk_in[19]), 
        .A5(cipher_text[19]), .A6(n298), .Y(n267) );
  AO222X1_HVT U396 ( .A1(adk_out0[20]), .A2(n296), .A3(n297), .A4(adk_in[20]), 
        .A5(cipher_text[20]), .A6(n298), .Y(n266) );
  AO222X1_HVT U397 ( .A1(adk_out0[21]), .A2(n296), .A3(n297), .A4(adk_in[21]), 
        .A5(cipher_text[21]), .A6(n298), .Y(n265) );
  AO222X1_HVT U398 ( .A1(adk_out0[22]), .A2(n296), .A3(n297), .A4(adk_in[22]), 
        .A5(cipher_text[22]), .A6(n298), .Y(n264) );
  AO222X1_HVT U399 ( .A1(adk_out0[23]), .A2(n296), .A3(n297), .A4(adk_in[23]), 
        .A5(cipher_text[23]), .A6(n298), .Y(n263) );
  AO222X1_HVT U400 ( .A1(adk_out0[24]), .A2(n296), .A3(n297), .A4(adk_in[24]), 
        .A5(cipher_text[24]), .A6(n298), .Y(n262) );
  AO222X1_HVT U401 ( .A1(adk_out0[25]), .A2(n296), .A3(n297), .A4(adk_in[25]), 
        .A5(cipher_text[25]), .A6(n298), .Y(n261) );
  AO222X1_HVT U402 ( .A1(adk_out0[26]), .A2(n296), .A3(n297), .A4(adk_in[26]), 
        .A5(cipher_text[26]), .A6(n298), .Y(n260) );
  AO222X1_HVT U403 ( .A1(adk_out0[27]), .A2(n296), .A3(n297), .A4(adk_in[27]), 
        .A5(cipher_text[27]), .A6(n298), .Y(n259) );
  AO222X1_HVT U404 ( .A1(adk_out0[28]), .A2(n296), .A3(n297), .A4(adk_in[28]), 
        .A5(cipher_text[28]), .A6(n298), .Y(n258) );
  AO222X1_HVT U405 ( .A1(adk_out0[29]), .A2(n296), .A3(n297), .A4(adk_in[29]), 
        .A5(cipher_text[29]), .A6(n298), .Y(n257) );
  AO222X1_HVT U406 ( .A1(adk_out0[30]), .A2(n296), .A3(n297), .A4(adk_in[30]), 
        .A5(cipher_text[30]), .A6(n298), .Y(n256) );
  AO222X1_HVT U407 ( .A1(adk_out0[31]), .A2(n296), .A3(n297), .A4(adk_in[31]), 
        .A5(cipher_text[31]), .A6(n298), .Y(n255) );
  AO222X1_HVT U408 ( .A1(adk_out0[32]), .A2(n296), .A3(n297), .A4(adk_in[32]), 
        .A5(cipher_text[32]), .A6(n298), .Y(n254) );
  AO222X1_HVT U409 ( .A1(adk_out0[33]), .A2(n296), .A3(n297), .A4(adk_in[33]), 
        .A5(cipher_text[33]), .A6(n298), .Y(n253) );
  AO222X1_HVT U410 ( .A1(adk_out0[34]), .A2(n296), .A3(n297), .A4(adk_in[34]), 
        .A5(cipher_text[34]), .A6(n298), .Y(n252) );
  AO222X1_HVT U411 ( .A1(adk_out0[35]), .A2(n296), .A3(n297), .A4(adk_in[35]), 
        .A5(cipher_text[35]), .A6(n298), .Y(n251) );
  AO222X1_HVT U412 ( .A1(adk_out0[36]), .A2(n296), .A3(n297), .A4(adk_in[36]), 
        .A5(cipher_text[36]), .A6(n298), .Y(n250) );
  AO222X1_HVT U413 ( .A1(adk_out0[37]), .A2(n296), .A3(n297), .A4(adk_in[37]), 
        .A5(cipher_text[37]), .A6(n298), .Y(n249) );
  AO222X1_HVT U414 ( .A1(adk_out0[38]), .A2(n296), .A3(n297), .A4(adk_in[38]), 
        .A5(cipher_text[38]), .A6(n298), .Y(n248) );
  AO222X1_HVT U415 ( .A1(adk_out0[39]), .A2(n296), .A3(n297), .A4(adk_in[39]), 
        .A5(cipher_text[39]), .A6(n298), .Y(n247) );
  AO222X1_HVT U416 ( .A1(adk_out0[40]), .A2(n296), .A3(n297), .A4(adk_in[40]), 
        .A5(cipher_text[40]), .A6(n298), .Y(n246) );
  AO222X1_HVT U417 ( .A1(adk_out0[41]), .A2(n296), .A3(n297), .A4(adk_in[41]), 
        .A5(cipher_text[41]), .A6(n298), .Y(n245) );
  AO222X1_HVT U418 ( .A1(adk_out0[42]), .A2(n296), .A3(n297), .A4(adk_in[42]), 
        .A5(cipher_text[42]), .A6(n298), .Y(n244) );
  AO222X1_HVT U419 ( .A1(adk_out0[43]), .A2(n296), .A3(n297), .A4(adk_in[43]), 
        .A5(cipher_text[43]), .A6(n298), .Y(n243) );
  AO222X1_HVT U420 ( .A1(adk_out0[44]), .A2(n296), .A3(n297), .A4(adk_in[44]), 
        .A5(cipher_text[44]), .A6(n298), .Y(n242) );
  AO222X1_HVT U421 ( .A1(adk_out0[45]), .A2(n296), .A3(n297), .A4(adk_in[45]), 
        .A5(cipher_text[45]), .A6(n298), .Y(n241) );
  AO222X1_HVT U422 ( .A1(adk_out0[46]), .A2(n296), .A3(n297), .A4(adk_in[46]), 
        .A5(cipher_text[46]), .A6(n298), .Y(n240) );
  AO222X1_HVT U423 ( .A1(adk_out0[47]), .A2(n296), .A3(n297), .A4(adk_in[47]), 
        .A5(cipher_text[47]), .A6(n298), .Y(n239) );
  AO222X1_HVT U424 ( .A1(adk_out0[48]), .A2(n296), .A3(n297), .A4(adk_in[48]), 
        .A5(cipher_text[48]), .A6(n298), .Y(n238) );
  AO222X1_HVT U425 ( .A1(adk_out0[49]), .A2(n296), .A3(n297), .A4(adk_in[49]), 
        .A5(cipher_text[49]), .A6(n298), .Y(n237) );
  AO222X1_HVT U426 ( .A1(adk_out0[50]), .A2(n296), .A3(n297), .A4(adk_in[50]), 
        .A5(cipher_text[50]), .A6(n298), .Y(n236) );
  AO222X1_HVT U427 ( .A1(adk_out0[51]), .A2(n296), .A3(n297), .A4(adk_in[51]), 
        .A5(cipher_text[51]), .A6(n298), .Y(n235) );
  AO222X1_HVT U428 ( .A1(adk_out0[52]), .A2(n296), .A3(n297), .A4(adk_in[52]), 
        .A5(cipher_text[52]), .A6(n298), .Y(n234) );
  AO222X1_HVT U429 ( .A1(adk_out0[53]), .A2(n296), .A3(n297), .A4(adk_in[53]), 
        .A5(cipher_text[53]), .A6(n298), .Y(n233) );
  AO222X1_HVT U430 ( .A1(adk_out0[54]), .A2(n296), .A3(n297), .A4(adk_in[54]), 
        .A5(cipher_text[54]), .A6(n298), .Y(n232) );
  AO222X1_HVT U431 ( .A1(adk_out0[55]), .A2(n296), .A3(n297), .A4(adk_in[55]), 
        .A5(cipher_text[55]), .A6(n298), .Y(n231) );
  AO222X1_HVT U432 ( .A1(adk_out0[56]), .A2(n296), .A3(n297), .A4(adk_in[56]), 
        .A5(cipher_text[56]), .A6(n298), .Y(n230) );
  AO222X1_HVT U433 ( .A1(adk_out0[57]), .A2(n296), .A3(n297), .A4(adk_in[57]), 
        .A5(cipher_text[57]), .A6(n298), .Y(n229) );
  AO222X1_HVT U434 ( .A1(adk_out0[58]), .A2(n296), .A3(n297), .A4(adk_in[58]), 
        .A5(cipher_text[58]), .A6(n298), .Y(n228) );
  AO222X1_HVT U435 ( .A1(adk_out0[59]), .A2(n296), .A3(n297), .A4(adk_in[59]), 
        .A5(cipher_text[59]), .A6(n298), .Y(n227) );
  AO222X1_HVT U436 ( .A1(adk_out0[60]), .A2(n296), .A3(n297), .A4(adk_in[60]), 
        .A5(cipher_text[60]), .A6(n298), .Y(n226) );
  AO222X1_HVT U437 ( .A1(adk_out0[61]), .A2(n296), .A3(n297), .A4(adk_in[61]), 
        .A5(cipher_text[61]), .A6(n298), .Y(n225) );
  AO222X1_HVT U438 ( .A1(adk_out0[62]), .A2(n296), .A3(n297), .A4(adk_in[62]), 
        .A5(cipher_text[62]), .A6(n298), .Y(n224) );
  AO222X1_HVT U439 ( .A1(adk_out0[63]), .A2(n296), .A3(n297), .A4(adk_in[63]), 
        .A5(cipher_text[63]), .A6(n298), .Y(n223) );
  AO222X1_HVT U440 ( .A1(adk_out0[64]), .A2(n296), .A3(n297), .A4(adk_in[64]), 
        .A5(cipher_text[64]), .A6(n298), .Y(n222) );
  AO222X1_HVT U441 ( .A1(adk_out0[65]), .A2(n296), .A3(n297), .A4(adk_in[65]), 
        .A5(cipher_text[65]), .A6(n298), .Y(n221) );
  AO222X1_HVT U442 ( .A1(adk_out0[66]), .A2(n296), .A3(n297), .A4(adk_in[66]), 
        .A5(cipher_text[66]), .A6(n298), .Y(n220) );
  AO222X1_HVT U443 ( .A1(adk_out0[67]), .A2(n296), .A3(n297), .A4(adk_in[67]), 
        .A5(cipher_text[67]), .A6(n298), .Y(n219) );
  AO222X1_HVT U444 ( .A1(adk_out0[68]), .A2(n296), .A3(n297), .A4(adk_in[68]), 
        .A5(cipher_text[68]), .A6(n298), .Y(n218) );
  AO222X1_HVT U445 ( .A1(adk_out0[69]), .A2(n296), .A3(n297), .A4(adk_in[69]), 
        .A5(cipher_text[69]), .A6(n298), .Y(n217) );
  AO222X1_HVT U446 ( .A1(adk_out0[70]), .A2(n296), .A3(n297), .A4(adk_in[70]), 
        .A5(cipher_text[70]), .A6(n298), .Y(n216) );
  AO222X1_HVT U447 ( .A1(adk_out0[71]), .A2(n296), .A3(n297), .A4(adk_in[71]), 
        .A5(cipher_text[71]), .A6(n298), .Y(n215) );
  AO222X1_HVT U448 ( .A1(adk_out0[72]), .A2(n296), .A3(n297), .A4(adk_in[72]), 
        .A5(cipher_text[72]), .A6(n298), .Y(n214) );
  AO222X1_HVT U449 ( .A1(adk_out0[73]), .A2(n296), .A3(n297), .A4(adk_in[73]), 
        .A5(cipher_text[73]), .A6(n298), .Y(n213) );
  AO222X1_HVT U450 ( .A1(adk_out0[74]), .A2(n296), .A3(n297), .A4(adk_in[74]), 
        .A5(cipher_text[74]), .A6(n298), .Y(n212) );
  AO222X1_HVT U451 ( .A1(adk_out0[75]), .A2(n296), .A3(n297), .A4(adk_in[75]), 
        .A5(cipher_text[75]), .A6(n298), .Y(n211) );
  AO222X1_HVT U452 ( .A1(adk_out0[76]), .A2(n296), .A3(n297), .A4(adk_in[76]), 
        .A5(cipher_text[76]), .A6(n298), .Y(n210) );
  AO222X1_HVT U453 ( .A1(adk_out0[77]), .A2(n296), .A3(n297), .A4(adk_in[77]), 
        .A5(cipher_text[77]), .A6(n298), .Y(n209) );
  AO222X1_HVT U454 ( .A1(adk_out0[78]), .A2(n296), .A3(n297), .A4(adk_in[78]), 
        .A5(cipher_text[78]), .A6(n298), .Y(n208) );
  AO222X1_HVT U455 ( .A1(adk_out0[79]), .A2(n296), .A3(n297), .A4(adk_in[79]), 
        .A5(cipher_text[79]), .A6(n298), .Y(n207) );
  AO222X1_HVT U456 ( .A1(adk_out0[80]), .A2(n296), .A3(n297), .A4(adk_in[80]), 
        .A5(cipher_text[80]), .A6(n298), .Y(n206) );
  AO222X1_HVT U457 ( .A1(adk_out0[81]), .A2(n296), .A3(n297), .A4(adk_in[81]), 
        .A5(cipher_text[81]), .A6(n298), .Y(n205) );
  AO222X1_HVT U458 ( .A1(adk_out0[82]), .A2(n296), .A3(n297), .A4(adk_in[82]), 
        .A5(cipher_text[82]), .A6(n298), .Y(n204) );
  AO222X1_HVT U459 ( .A1(adk_out0[83]), .A2(n296), .A3(n297), .A4(adk_in[83]), 
        .A5(cipher_text[83]), .A6(n298), .Y(n203) );
  AO222X1_HVT U460 ( .A1(adk_out0[84]), .A2(n296), .A3(n297), .A4(adk_in[84]), 
        .A5(cipher_text[84]), .A6(n298), .Y(n202) );
  AO222X1_HVT U461 ( .A1(adk_out0[85]), .A2(n296), .A3(n297), .A4(adk_in[85]), 
        .A5(cipher_text[85]), .A6(n298), .Y(n201) );
  AO222X1_HVT U462 ( .A1(adk_out0[86]), .A2(n296), .A3(n297), .A4(adk_in[86]), 
        .A5(cipher_text[86]), .A6(n298), .Y(n200) );
  AO222X1_HVT U463 ( .A1(adk_out0[87]), .A2(n296), .A3(n297), .A4(adk_in[87]), 
        .A5(cipher_text[87]), .A6(n298), .Y(n199) );
  AO222X1_HVT U464 ( .A1(adk_out0[88]), .A2(n296), .A3(n297), .A4(adk_in[88]), 
        .A5(cipher_text[88]), .A6(n298), .Y(n198) );
  AO222X1_HVT U465 ( .A1(adk_out0[89]), .A2(n296), .A3(n297), .A4(adk_in[89]), 
        .A5(cipher_text[89]), .A6(n298), .Y(n197) );
  AO222X1_HVT U466 ( .A1(adk_out0[90]), .A2(n296), .A3(n297), .A4(adk_in[90]), 
        .A5(cipher_text[90]), .A6(n298), .Y(n196) );
  AO222X1_HVT U467 ( .A1(adk_out0[91]), .A2(n296), .A3(n297), .A4(adk_in[91]), 
        .A5(cipher_text[91]), .A6(n298), .Y(n195) );
  AO222X1_HVT U468 ( .A1(adk_out0[92]), .A2(n296), .A3(n297), .A4(adk_in[92]), 
        .A5(cipher_text[92]), .A6(n298), .Y(n194) );
  AO222X1_HVT U469 ( .A1(adk_out0[93]), .A2(n296), .A3(n297), .A4(adk_in[93]), 
        .A5(cipher_text[93]), .A6(n298), .Y(n193) );
  AO222X1_HVT U470 ( .A1(adk_out0[94]), .A2(n296), .A3(n297), .A4(adk_in[94]), 
        .A5(cipher_text[94]), .A6(n298), .Y(n192) );
  AO222X1_HVT U471 ( .A1(adk_out0[95]), .A2(n296), .A3(n297), .A4(adk_in[95]), 
        .A5(cipher_text[95]), .A6(n298), .Y(n191) );
  AO222X1_HVT U472 ( .A1(adk_out0[96]), .A2(n296), .A3(n297), .A4(adk_in[96]), 
        .A5(cipher_text[96]), .A6(n298), .Y(n190) );
  AO222X1_HVT U473 ( .A1(adk_out0[97]), .A2(n296), .A3(n297), .A4(adk_in[97]), 
        .A5(cipher_text[97]), .A6(n298), .Y(n189) );
  AO222X1_HVT U474 ( .A1(adk_out0[98]), .A2(n296), .A3(n297), .A4(adk_in[98]), 
        .A5(cipher_text[98]), .A6(n298), .Y(n188) );
  AO222X1_HVT U475 ( .A1(adk_out0[99]), .A2(n296), .A3(n297), .A4(adk_in[99]), 
        .A5(cipher_text[99]), .A6(n298), .Y(n187) );
  AO222X1_HVT U476 ( .A1(adk_out0[100]), .A2(n296), .A3(n297), .A4(adk_in[100]), .A5(cipher_text[100]), .A6(n298), .Y(n186) );
  AO222X1_HVT U477 ( .A1(adk_out0[101]), .A2(n296), .A3(n297), .A4(adk_in[101]), .A5(cipher_text[101]), .A6(n298), .Y(n185) );
  AO222X1_HVT U478 ( .A1(adk_out0[102]), .A2(n296), .A3(n297), .A4(adk_in[102]), .A5(cipher_text[102]), .A6(n298), .Y(n184) );
  AO222X1_HVT U479 ( .A1(adk_out0[103]), .A2(n296), .A3(n297), .A4(adk_in[103]), .A5(cipher_text[103]), .A6(n298), .Y(n183) );
  AO222X1_HVT U480 ( .A1(adk_out0[104]), .A2(n296), .A3(n297), .A4(adk_in[104]), .A5(cipher_text[104]), .A6(n298), .Y(n182) );
  AO222X1_HVT U481 ( .A1(adk_out0[105]), .A2(n296), .A3(n297), .A4(adk_in[105]), .A5(cipher_text[105]), .A6(n298), .Y(n181) );
  AO222X1_HVT U482 ( .A1(adk_out0[106]), .A2(n296), .A3(n297), .A4(adk_in[106]), .A5(cipher_text[106]), .A6(n298), .Y(n180) );
  AO222X1_HVT U483 ( .A1(adk_out0[107]), .A2(n296), .A3(n297), .A4(adk_in[107]), .A5(cipher_text[107]), .A6(n298), .Y(n179) );
  AO222X1_HVT U484 ( .A1(adk_out0[108]), .A2(n296), .A3(n297), .A4(adk_in[108]), .A5(cipher_text[108]), .A6(n298), .Y(n178) );
  AO222X1_HVT U485 ( .A1(adk_out0[109]), .A2(n296), .A3(n297), .A4(adk_in[109]), .A5(cipher_text[109]), .A6(n298), .Y(n177) );
  AO222X1_HVT U486 ( .A1(adk_out0[110]), .A2(n296), .A3(n297), .A4(adk_in[110]), .A5(cipher_text[110]), .A6(n298), .Y(n176) );
  AO222X1_HVT U487 ( .A1(adk_out0[111]), .A2(n296), .A3(n297), .A4(adk_in[111]), .A5(cipher_text[111]), .A6(n298), .Y(n175) );
  AO222X1_HVT U488 ( .A1(adk_out0[112]), .A2(n296), .A3(n297), .A4(adk_in[112]), .A5(cipher_text[112]), .A6(n298), .Y(n174) );
  AO222X1_HVT U489 ( .A1(adk_out0[113]), .A2(n296), .A3(n297), .A4(adk_in[113]), .A5(cipher_text[113]), .A6(n298), .Y(n173) );
  AO222X1_HVT U490 ( .A1(adk_out0[114]), .A2(n296), .A3(n297), .A4(adk_in[114]), .A5(cipher_text[114]), .A6(n298), .Y(n172) );
  AO222X1_HVT U491 ( .A1(adk_out0[115]), .A2(n296), .A3(n297), .A4(adk_in[115]), .A5(cipher_text[115]), .A6(n298), .Y(n171) );
  AO222X1_HVT U492 ( .A1(adk_out0[116]), .A2(n296), .A3(n297), .A4(adk_in[116]), .A5(cipher_text[116]), .A6(n298), .Y(n170) );
  AO222X1_HVT U493 ( .A1(adk_out0[117]), .A2(n296), .A3(n297), .A4(adk_in[117]), .A5(cipher_text[117]), .A6(n298), .Y(n169) );
  AO222X1_HVT U494 ( .A1(adk_out0[118]), .A2(n296), .A3(n297), .A4(adk_in[118]), .A5(cipher_text[118]), .A6(n298), .Y(n168) );
  AO222X1_HVT U495 ( .A1(adk_out0[119]), .A2(n296), .A3(n297), .A4(adk_in[119]), .A5(cipher_text[119]), .A6(n298), .Y(n167) );
  AO222X1_HVT U496 ( .A1(adk_out0[120]), .A2(n296), .A3(n297), .A4(adk_in[120]), .A5(cipher_text[120]), .A6(n298), .Y(n166) );
  AO222X1_HVT U497 ( .A1(adk_out0[121]), .A2(n296), .A3(n297), .A4(adk_in[121]), .A5(cipher_text[121]), .A6(n298), .Y(n165) );
  AO222X1_HVT U498 ( .A1(adk_out0[122]), .A2(n296), .A3(n297), .A4(adk_in[122]), .A5(cipher_text[122]), .A6(n298), .Y(n164) );
  AO222X1_HVT U499 ( .A1(adk_out0[123]), .A2(n296), .A3(n297), .A4(adk_in[123]), .A5(cipher_text[123]), .A6(n298), .Y(n163) );
  AO222X1_HVT U500 ( .A1(adk_out0[124]), .A2(n296), .A3(n297), .A4(adk_in[124]), .A5(cipher_text[124]), .A6(n298), .Y(n162) );
  AO222X1_HVT U501 ( .A1(adk_out0[125]), .A2(n296), .A3(n297), .A4(adk_in[125]), .A5(cipher_text[125]), .A6(n298), .Y(n161) );
  AO222X1_HVT U502 ( .A1(adk_out0[126]), .A2(n296), .A3(n297), .A4(adk_in[126]), .A5(cipher_text[126]), .A6(n298), .Y(n160) );
  AO222X1_HVT U503 ( .A1(adk_out0[127]), .A2(n296), .A3(n297), .A4(adk_in[127]), .A5(cipher_text[127]), .A6(n298), .Y(n159) );
  AO222X1_HVT U504 ( .A1(key[0]), .A2(n296), .A3(n297), .A4(key_round[0]), 
        .A5(keyout[0]), .A6(n298), .Y(n158) );
  AO222X1_HVT U505 ( .A1(key[1]), .A2(n296), .A3(n297), .A4(key_round[1]), 
        .A5(keyout[1]), .A6(n298), .Y(n157) );
  AO222X1_HVT U506 ( .A1(key[2]), .A2(n296), .A3(n297), .A4(key_round[2]), 
        .A5(keyout[2]), .A6(n298), .Y(n156) );
  AO222X1_HVT U507 ( .A1(key[3]), .A2(n296), .A3(n297), .A4(key_round[3]), 
        .A5(keyout[3]), .A6(n298), .Y(n155) );
  AO222X1_HVT U508 ( .A1(key[4]), .A2(n296), .A3(n297), .A4(key_round[4]), 
        .A5(keyout[4]), .A6(n298), .Y(n154) );
  AO222X1_HVT U509 ( .A1(key[5]), .A2(n296), .A3(n297), .A4(key_round[5]), 
        .A5(keyout[5]), .A6(n298), .Y(n153) );
  AO222X1_HVT U510 ( .A1(key[6]), .A2(n296), .A3(n297), .A4(key_round[6]), 
        .A5(keyout[6]), .A6(n298), .Y(n152) );
  AO222X1_HVT U511 ( .A1(key[7]), .A2(n296), .A3(n297), .A4(key_round[7]), 
        .A5(keyout[7]), .A6(n298), .Y(n151) );
  AO222X1_HVT U512 ( .A1(key[8]), .A2(n296), .A3(n297), .A4(key_round[8]), 
        .A5(keyout[8]), .A6(n298), .Y(n150) );
  AO222X1_HVT U513 ( .A1(key[9]), .A2(n296), .A3(n297), .A4(key_round[9]), 
        .A5(keyout[9]), .A6(n298), .Y(n149) );
  AO222X1_HVT U514 ( .A1(key[10]), .A2(n296), .A3(n297), .A4(key_round[10]), 
        .A5(keyout[10]), .A6(n298), .Y(n148) );
  AO222X1_HVT U515 ( .A1(key[11]), .A2(n296), .A3(n297), .A4(key_round[11]), 
        .A5(keyout[11]), .A6(n298), .Y(n147) );
  AO222X1_HVT U516 ( .A1(key[12]), .A2(n296), .A3(n297), .A4(key_round[12]), 
        .A5(keyout[12]), .A6(n298), .Y(n146) );
  AO222X1_HVT U517 ( .A1(key[13]), .A2(n296), .A3(n297), .A4(key_round[13]), 
        .A5(keyout[13]), .A6(n298), .Y(n145) );
  AO222X1_HVT U518 ( .A1(key[14]), .A2(n296), .A3(n297), .A4(key_round[14]), 
        .A5(keyout[14]), .A6(n298), .Y(n144) );
  AO222X1_HVT U519 ( .A1(key[15]), .A2(n296), .A3(n297), .A4(key_round[15]), 
        .A5(keyout[15]), .A6(n298), .Y(n143) );
  AO222X1_HVT U520 ( .A1(key[16]), .A2(n296), .A3(n297), .A4(key_round[16]), 
        .A5(keyout[16]), .A6(n298), .Y(n142) );
  AO222X1_HVT U521 ( .A1(key[17]), .A2(n296), .A3(n297), .A4(key_round[17]), 
        .A5(keyout[17]), .A6(n298), .Y(n141) );
  AO222X1_HVT U522 ( .A1(key[18]), .A2(n296), .A3(n297), .A4(key_round[18]), 
        .A5(keyout[18]), .A6(n298), .Y(n140) );
  AO222X1_HVT U523 ( .A1(key[19]), .A2(n296), .A3(n297), .A4(key_round[19]), 
        .A5(keyout[19]), .A6(n298), .Y(n139) );
  AO222X1_HVT U524 ( .A1(key[20]), .A2(n296), .A3(n297), .A4(key_round[20]), 
        .A5(keyout[20]), .A6(n298), .Y(n138) );
  AO222X1_HVT U525 ( .A1(key[21]), .A2(n296), .A3(n297), .A4(key_round[21]), 
        .A5(keyout[21]), .A6(n298), .Y(n137) );
  AO222X1_HVT U526 ( .A1(key[22]), .A2(n296), .A3(n297), .A4(key_round[22]), 
        .A5(keyout[22]), .A6(n298), .Y(n136) );
  AO222X1_HVT U527 ( .A1(key[23]), .A2(n296), .A3(n297), .A4(key_round[23]), 
        .A5(keyout[23]), .A6(n298), .Y(n135) );
  AO222X1_HVT U528 ( .A1(key[24]), .A2(n296), .A3(n297), .A4(key_round[24]), 
        .A5(keyout[24]), .A6(n298), .Y(n134) );
  AO222X1_HVT U529 ( .A1(key[25]), .A2(n296), .A3(n297), .A4(key_round[25]), 
        .A5(keyout[25]), .A6(n298), .Y(n133) );
  AO222X1_HVT U530 ( .A1(key[26]), .A2(n296), .A3(n297), .A4(key_round[26]), 
        .A5(keyout[26]), .A6(n298), .Y(n132) );
  AO222X1_HVT U531 ( .A1(key[27]), .A2(n296), .A3(n297), .A4(key_round[27]), 
        .A5(keyout[27]), .A6(n298), .Y(n131) );
  AO222X1_HVT U532 ( .A1(key[28]), .A2(n296), .A3(n297), .A4(key_round[28]), 
        .A5(keyout[28]), .A6(n298), .Y(n130) );
  AO222X1_HVT U533 ( .A1(key[29]), .A2(n296), .A3(n297), .A4(key_round[29]), 
        .A5(keyout[29]), .A6(n298), .Y(n129) );
  AO222X1_HVT U534 ( .A1(key[30]), .A2(n296), .A3(n297), .A4(key_round[30]), 
        .A5(keyout[30]), .A6(n298), .Y(n128) );
  AO222X1_HVT U535 ( .A1(key[31]), .A2(n296), .A3(n297), .A4(key_round[31]), 
        .A5(keyout[31]), .A6(n298), .Y(n127) );
  AO222X1_HVT U536 ( .A1(key[32]), .A2(n296), .A3(n297), .A4(key_round[32]), 
        .A5(keyout[32]), .A6(n298), .Y(n126) );
  AO222X1_HVT U537 ( .A1(key[33]), .A2(n296), .A3(n297), .A4(key_round[33]), 
        .A5(keyout[33]), .A6(n298), .Y(n125) );
  AO222X1_HVT U538 ( .A1(key[34]), .A2(n296), .A3(n297), .A4(key_round[34]), 
        .A5(keyout[34]), .A6(n298), .Y(n124) );
  AO222X1_HVT U539 ( .A1(key[35]), .A2(n296), .A3(n297), .A4(key_round[35]), 
        .A5(keyout[35]), .A6(n298), .Y(n123) );
  AO222X1_HVT U540 ( .A1(key[36]), .A2(n296), .A3(n297), .A4(key_round[36]), 
        .A5(keyout[36]), .A6(n298), .Y(n122) );
  AO222X1_HVT U541 ( .A1(key[37]), .A2(n296), .A3(n297), .A4(key_round[37]), 
        .A5(keyout[37]), .A6(n298), .Y(n121) );
  AO222X1_HVT U542 ( .A1(key[38]), .A2(n296), .A3(n297), .A4(key_round[38]), 
        .A5(keyout[38]), .A6(n298), .Y(n120) );
  AO222X1_HVT U543 ( .A1(key[39]), .A2(n296), .A3(n297), .A4(key_round[39]), 
        .A5(keyout[39]), .A6(n298), .Y(n119) );
  AO222X1_HVT U544 ( .A1(key[40]), .A2(n296), .A3(n297), .A4(key_round[40]), 
        .A5(keyout[40]), .A6(n298), .Y(n118) );
  AO222X1_HVT U545 ( .A1(key[41]), .A2(n296), .A3(n297), .A4(key_round[41]), 
        .A5(keyout[41]), .A6(n298), .Y(n117) );
  AO222X1_HVT U546 ( .A1(key[42]), .A2(n296), .A3(n297), .A4(key_round[42]), 
        .A5(keyout[42]), .A6(n298), .Y(n116) );
  AO222X1_HVT U547 ( .A1(key[43]), .A2(n296), .A3(n297), .A4(key_round[43]), 
        .A5(keyout[43]), .A6(n298), .Y(n115) );
  AO222X1_HVT U548 ( .A1(key[44]), .A2(n296), .A3(n297), .A4(key_round[44]), 
        .A5(keyout[44]), .A6(n298), .Y(n114) );
  AO222X1_HVT U549 ( .A1(key[45]), .A2(n296), .A3(n297), .A4(key_round[45]), 
        .A5(keyout[45]), .A6(n298), .Y(n113) );
  AO222X1_HVT U550 ( .A1(key[46]), .A2(n296), .A3(n297), .A4(key_round[46]), 
        .A5(keyout[46]), .A6(n298), .Y(n112) );
  AO222X1_HVT U551 ( .A1(key[47]), .A2(n296), .A3(n297), .A4(key_round[47]), 
        .A5(keyout[47]), .A6(n298), .Y(n111) );
  AO222X1_HVT U552 ( .A1(key[48]), .A2(n296), .A3(n297), .A4(key_round[48]), 
        .A5(keyout[48]), .A6(n298), .Y(n110) );
  AO222X1_HVT U553 ( .A1(key[49]), .A2(n296), .A3(n297), .A4(key_round[49]), 
        .A5(keyout[49]), .A6(n298), .Y(n109) );
  AO222X1_HVT U554 ( .A1(key[50]), .A2(n296), .A3(n297), .A4(key_round[50]), 
        .A5(keyout[50]), .A6(n298), .Y(n108) );
  AO222X1_HVT U555 ( .A1(key[51]), .A2(n296), .A3(n297), .A4(key_round[51]), 
        .A5(keyout[51]), .A6(n298), .Y(n107) );
  AO222X1_HVT U556 ( .A1(key[52]), .A2(n296), .A3(n297), .A4(key_round[52]), 
        .A5(keyout[52]), .A6(n298), .Y(n106) );
  AO222X1_HVT U557 ( .A1(key[53]), .A2(n296), .A3(n297), .A4(key_round[53]), 
        .A5(keyout[53]), .A6(n298), .Y(n105) );
  AO222X1_HVT U558 ( .A1(key[54]), .A2(n296), .A3(n297), .A4(key_round[54]), 
        .A5(keyout[54]), .A6(n298), .Y(n104) );
  AO222X1_HVT U559 ( .A1(key[55]), .A2(n296), .A3(n297), .A4(key_round[55]), 
        .A5(keyout[55]), .A6(n298), .Y(n103) );
  AO222X1_HVT U560 ( .A1(key[56]), .A2(n296), .A3(n297), .A4(key_round[56]), 
        .A5(keyout[56]), .A6(n298), .Y(n102) );
  AO222X1_HVT U561 ( .A1(key[57]), .A2(n296), .A3(n297), .A4(key_round[57]), 
        .A5(keyout[57]), .A6(n298), .Y(n101) );
  AO222X1_HVT U562 ( .A1(key[58]), .A2(n296), .A3(n297), .A4(key_round[58]), 
        .A5(keyout[58]), .A6(n298), .Y(n100) );
  AND2X1_HVT U563 ( .A1(n304), .A2(n315), .Y(n298) );
  INVX0_HVT U564 ( .A(n316), .Y(n304) );
  AND2X1_HVT U565 ( .A1(n301), .A2(n316), .Y(n297) );
  INVX0_HVT U566 ( .A(reset), .Y(n301) );
  NOR2X0_HVT U567 ( .A1(n316), .A2(n315), .Y(n296) );
  OR3X1_HVT U568 ( .A1(round_number[0]), .A2(round_number[3]), .A3(n314), .Y(
        n315) );
  AO21X1_HVT U569 ( .A1(round_number[3]), .A2(n314), .A3(reset), .Y(n316) );
  NAND2X0_HVT U570 ( .A1(n295), .A2(n293), .Y(n314) );
endmodule

