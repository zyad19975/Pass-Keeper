
module sbox_13 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n2, n10, n23, n38, n50, n51, n95, n96, n113, n114, n117, n119, n210,
         n211, n212, n213, n216, n217, n218, n219, n231, n232, n234, n236,
         n238, n240, n242, n246, n255, n256, n258, n259, n261, n264, n272,
         n274, n275, n282, n283, n285, n286, n293, n297, n300, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774;

  NAND2X0_HVT U4 ( .A1(n432), .A2(n437), .Y(n772) );
  NAND2X0_HVT U5 ( .A1(n96), .A2(n500), .Y(n770) );
  NAND2X0_HVT U15 ( .A1(n773), .A2(n454), .Y(n761) );
  NAND2X0_HVT U21 ( .A1(n436), .A2(n507), .Y(n755) );
  NAND2X0_HVT U24 ( .A1(n119), .A2(n348), .Y(n753) );
  NAND2X0_HVT U33 ( .A1(n293), .A2(n348), .Y(n744) );
  NAND2X0_HVT U42 ( .A1(n383), .A2(n388), .Y(n736) );
  NAND2X0_HVT U53 ( .A1(n726), .A2(n735), .Y(n727) );
  NAND2X0_HVT U56 ( .A1(n432), .A2(n722), .Y(n723) );
  NAND2X0_HVT U58 ( .A1(n415), .A2(n773), .Y(n720) );
  NAND2X0_HVT U62 ( .A1(n348), .A2(n339), .Y(n716) );
  MUX41X1_HVT U63 ( .A1(n716), .A3(n528), .A2(n217), .A4(n526), .S0(n470), 
        .S1(n491), .Y(n715) );
  MUX41X1_HVT U68 ( .A1(n407), .A3(n712), .A2(n711), .A4(n713), .S0(n307), 
        .S1(n513), .Y(n710) );
  NAND2X0_HVT U73 ( .A1(n431), .A2(n705), .Y(n706) );
  AND2X1_HVT U83 ( .A1(n333), .A2(n399), .Y(n694) );
  NAND2X0_HVT U85 ( .A1(n507), .A2(n417), .Y(n692) );
  MUX41X1_HVT U86 ( .A1(n556), .A3(n692), .A2(n474), .A4(n472), .S0(n307), 
        .S1(n470), .Y(n691) );
  MUX41X1_HVT U97 ( .A1(n558), .A3(n475), .A2(n383), .A4(n761), .S0(n307), 
        .S1(n391), .Y(n682) );
  NAND2X0_HVT U101 ( .A1(n677), .A2(n676), .Y(n678) );
  MUX41X1_HVT U103 ( .A1(n437), .A3(n95), .A2(n357), .A4(n742), .S0(n308), 
        .S1(n512), .Y(n674) );
  MUX41X1_HVT U105 ( .A1(n553), .A3(n730), .A2(n673), .A4(n546), .S0(n489), 
        .S1(n391), .Y(n672) );
  NAND2X0_HVT U110 ( .A1(n339), .A2(n669), .Y(n670) );
  AND2X1_HVT U115 ( .A1(n96), .A2(n455), .Y(n666) );
  MUX41X1_HVT U116 ( .A1(n764), .A3(n666), .A2(n354), .A4(n746), .S0(n487), 
        .S1(n468), .Y(n665) );
  NAND2X0_HVT U123 ( .A1(n657), .A2(n656), .Y(n658) );
  MUX41X1_HVT U125 ( .A1(n755), .A3(n479), .A2(n407), .A4(n542), .S0(n308), 
        .S1(n468), .Y(n654) );
  MUX41X1_HVT U136 ( .A1(n472), .A3(n744), .A2(n522), .A4(n741), .S0(n486), 
        .S1(n470), .Y(n644) );
  AND2X1_HVT U140 ( .A1(n431), .A2(n507), .Y(n640) );
  MUX41X1_HVT U142 ( .A1(n530), .A3(n454), .A2(n545), .A4(n431), .S0(n489), 
        .S1(n469), .Y(n638) );
  OA21X1_HVT U151 ( .A1(n738), .A2(n389), .A3(n630), .Y(n631) );
  MUX41X1_HVT U153 ( .A1(n670), .A3(n476), .A2(n339), .A4(n363), .S0(n488), 
        .S1(n513), .Y(n628) );
  AND2X1_HVT U154 ( .A1(n495), .A2(n388), .Y(n627) );
  NAND2X0_HVT U158 ( .A1(n505), .A2(n417), .Y(n623) );
  MUX41X1_HVT U159 ( .A1(n764), .A3(n453), .A2(n623), .A4(n562), .S0(n508), 
        .S1(n458), .Y(n622) );
  AND2X1_HVT U162 ( .A1(n451), .A2(n286), .Y(n619) );
  NAND2X0_HVT U166 ( .A1(n418), .A2(n722), .Y(n615) );
  NAND2X0_HVT U167 ( .A1(n411), .A2(n507), .Y(n614) );
  MUX41X1_HVT U168 ( .A1(n535), .A3(n51), .A2(n614), .A4(n615), .S0(n314), 
        .S1(n513), .Y(n613) );
  MUX41X1_HVT U176 ( .A1(n497), .A3(n608), .A2(n531), .A4(n327), .S0(n470), 
        .S1(n508), .Y(n607) );
  NAND2X0_HVT U177 ( .A1(n503), .A2(n212), .Y(n606) );
  MUX41X1_HVT U179 ( .A1(n749), .A3(n549), .A2(n536), .A4(n550), .S0(n314), 
        .S1(n512), .Y(n604) );
  MUX41X1_HVT U180 ( .A1(n529), .A3(n767), .A2(n352), .A4(n471), .S0(n493), 
        .S1(n508), .Y(n603) );
  MUX41X1_HVT U182 ( .A1(n541), .A3(n436), .A2(n524), .A4(n548), .S0(n470), 
        .S1(n486), .Y(n601) );
  MUX41X1_HVT U189 ( .A1(n595), .A3(n327), .A2(n596), .A4(n546), .S0(n493), 
        .S1(n307), .Y(n594) );
  MUX41X1_HVT U194 ( .A1(n737), .A3(n750), .A2(n533), .A4(n350), .S0(n493), 
        .S1(n307), .Y(n590) );
  AO21X1_HVT U197 ( .A1(n474), .A2(n494), .A3(n555), .Y(n587) );
  MUX41X1_HVT U203 ( .A1(n741), .A3(n519), .A2(n765), .A4(n745), .S0(n486), 
        .S1(n458), .Y(n581) );
  NAND2X0_HVT U208 ( .A1(n504), .A2(n433), .Y(n669) );
  NAND2X0_HVT U212 ( .A1(n333), .A2(n381), .Y(n722) );
  NAND2X0_HVT U214 ( .A1(n451), .A2(n507), .Y(n577) );
  NAND2X0_HVT U215 ( .A1(n669), .A2(n51), .Y(n576) );
  NAND2X0_HVT U218 ( .A1(n349), .A2(n413), .Y(n630) );
  NAND2X0_HVT U220 ( .A1(n494), .A2(n577), .Y(n697) );
  INVX0_HVT U241 ( .A(n753), .Y(n564) );
  INVX0_HVT U245 ( .A(n770), .Y(n562) );
  INVX0_HVT U251 ( .A(n746), .Y(n559) );
  INVX0_HVT U256 ( .A(n630), .Y(n555) );
  INVX0_HVT U265 ( .A(n751), .Y(n548) );
  INVX0_HVT U268 ( .A(n755), .Y(n547) );
  INVX0_HVT U270 ( .A(n576), .Y(n546) );
  INVX0_HVT U278 ( .A(n744), .Y(n539) );
  INVX0_HVT U284 ( .A(n577), .Y(n536) );
  INVX0_HVT U285 ( .A(n574), .Y(n535) );
  INVX0_HVT U289 ( .A(n676), .Y(n531) );
  INVX0_HVT U295 ( .A(n772), .Y(n529) );
  INVX0_HVT U296 ( .A(n761), .Y(n528) );
  INVX0_HVT U300 ( .A(n737), .Y(n524) );
  INVX0_HVT U306 ( .A(n614), .Y(n520) );
  INVX0_HVT U309 ( .A(n757), .Y(n518) );
  INVX1_HVT U1 ( .A(n498), .Y(n399) );
  INVX1_HVT U2 ( .A(n438), .Y(n382) );
  INVX1_HVT U3 ( .A(n359), .Y(n507) );
  MUX21X1_HVT U6 ( .A1(n381), .A2(n453), .S0(n219), .Y(n673) );
  MUX21X1_HVT U7 ( .A1(n663), .A2(n664), .S0(n494), .Y(n662) );
  AO21X1_HVT U8 ( .A1(n487), .A2(n51), .A3(n451), .Y(n663) );
  NOR3X0_HVT U9 ( .A1(n242), .A2(n219), .A3(n212), .Y(n651) );
  INVX1_HVT U10 ( .A(n443), .Y(n96) );
  INVX1_HVT U11 ( .A(n486), .Y(n353) );
  AND2X1_HVT U12 ( .A1(n231), .A2(n232), .Y(n2) );
  AND2X1_HVT U13 ( .A1(n439), .A2(n467), .Y(n10) );
  INVX1_HVT U14 ( .A(n349), .Y(n350) );
  INVX1_HVT U16 ( .A(n495), .Y(n445) );
  INVX1_HVT U17 ( .A(in[7]), .Y(n516) );
  INVX1_HVT U18 ( .A(n317), .Y(n521) );
  INVX0_HVT U19 ( .A(n399), .Y(n212) );
  MUX21X1_HVT U20 ( .A1(n560), .A2(n363), .S0(n510), .Y(n664) );
  NAND2X0_HVT U22 ( .A1(n417), .A2(n342), .Y(n23) );
  NAND2X0_HVT U23 ( .A1(n453), .A2(n414), .Y(n38) );
  NAND2X0_HVT U25 ( .A1(n23), .A2(n38), .Y(n620) );
  NBUFFX2_HVT U26 ( .A(n359), .Y(n414) );
  AND3X1_HVT U27 ( .A1(n339), .A2(n117), .A3(n697), .Y(n698) );
  INVX1_HVT U28 ( .A(n722), .Y(n558) );
  AO21X1_HVT U29 ( .A1(n507), .A2(n325), .A3(n389), .Y(n677) );
  INVX1_HVT U30 ( .A(n516), .Y(n514) );
  MUX21X1_HVT U31 ( .A1(n747), .A2(n576), .S0(n493), .Y(n570) );
  INVX1_HVT U32 ( .A(n669), .Y(n545) );
  MUX21X1_HVT U34 ( .A1(n527), .A2(n748), .S0(n445), .Y(n637) );
  INVX1_HVT U35 ( .A(n516), .Y(n513) );
  INVX1_HVT U36 ( .A(n317), .Y(n411) );
  INVX1_HVT U37 ( .A(n510), .Y(n508) );
  INVX1_HVT U38 ( .A(n275), .Y(n503) );
  MUX21X1_HVT U39 ( .A1(n415), .A2(n339), .S0(n503), .Y(n596) );
  INVX1_HVT U40 ( .A(n510), .Y(n509) );
  MUX21X1_HVT U41 ( .A1(n95), .A2(n325), .S0(n490), .Y(n711) );
  XNOR2X1_HVT U43 ( .A1(n463), .A2(n508), .Y(n483) );
  INVX1_HVT U44 ( .A(n282), .Y(n275) );
  INVX1_HVT U45 ( .A(n308), .Y(n242) );
  INVX1_HVT U46 ( .A(n468), .Y(n389) );
  INVX1_HVT U47 ( .A(n308), .Y(n394) );
  MUX21X1_HVT U48 ( .A1(n325), .A2(n573), .S0(n495), .Y(n338) );
  INVX1_HVT U49 ( .A(n442), .Y(n617) );
  INVX1_HVT U50 ( .A(n747), .Y(n552) );
  INVX1_HVT U51 ( .A(n488), .Y(n365) );
  MUX21X1_HVT U52 ( .A1(n431), .A2(n756), .S0(n445), .Y(n699) );
  INVX1_HVT U54 ( .A(n488), .Y(n351) );
  XNOR2X1_HVT U55 ( .A1(n246), .A2(n430), .Y(n733) );
  MUX21X1_HVT U57 ( .A1(n454), .A2(n434), .S0(n383), .Y(n684) );
  MUX21X1_HVT U59 ( .A1(n431), .A2(n436), .S0(n342), .Y(n689) );
  MUX21X1_HVT U60 ( .A1(n476), .A2(n680), .S0(n731), .Y(n679) );
  MUX21X1_HVT U61 ( .A1(n636), .A2(n637), .S0(n365), .Y(n635) );
  MUX21X1_HVT U64 ( .A1(n631), .A2(n632), .S0(n488), .Y(n629) );
  INVX1_HVT U65 ( .A(n494), .Y(n345) );
  MUX21X1_HVT U66 ( .A1(n293), .A2(n411), .S0(n504), .Y(n608) );
  MUX21X1_HVT U67 ( .A1(n599), .A2(n600), .S0(n487), .Y(n598) );
  INVX1_HVT U69 ( .A(n738), .Y(n519) );
  MUX21X1_HVT U70 ( .A1(n729), .A2(n725), .S0(n365), .Y(n724) );
  INVX1_HVT U71 ( .A(n470), .Y(n218) );
  INVX1_HVT U72 ( .A(n489), .Y(n444) );
  INVX1_HVT U74 ( .A(n491), .Y(n309) );
  INVX1_HVT U75 ( .A(n345), .Y(n512) );
  INVX1_HVT U76 ( .A(n429), .Y(n408) );
  NBUFFX2_HVT U77 ( .A(n509), .Y(n307) );
  INVX1_HVT U78 ( .A(n490), .Y(n429) );
  NBUFFX2_HVT U79 ( .A(n515), .Y(n493) );
  INVX1_HVT U80 ( .A(n493), .Y(n421) );
  INVX0_HVT U81 ( .A(n332), .Y(n219) );
  INVX1_HVT U82 ( .A(n440), .Y(n358) );
  INVX0_HVT U84 ( .A(n358), .Y(n359) );
  NBUFFX2_HVT U87 ( .A(n509), .Y(n308) );
  INVX0_HVT U88 ( .A(n543), .Y(n432) );
  INVX1_HVT U89 ( .A(n432), .Y(n434) );
  INVX0_HVT U90 ( .A(n381), .Y(n325) );
  INVX0_HVT U91 ( .A(n321), .Y(n119) );
  NBUFFX2_HVT U92 ( .A(n326), .Y(n499) );
  INVX0_HVT U93 ( .A(n499), .Y(n467) );
  INVX1_HVT U94 ( .A(n499), .Y(n274) );
  INVX1_HVT U95 ( .A(n543), .Y(n433) );
  NBUFFX2_HVT U96 ( .A(in[0]), .Y(n496) );
  INVX1_HVT U98 ( .A(n742), .Y(n363) );
  INVX1_HVT U99 ( .A(n561), .Y(n286) );
  XNOR2X1_HVT U100 ( .A1(n420), .A2(n414), .Y(n474) );
  AND2X1_HVT U102 ( .A1(n334), .A2(n335), .Y(n50) );
  INVX0_HVT U104 ( .A(n360), .Y(n760) );
  MUX21X1_HVT U106 ( .A1(n318), .A2(n119), .S0(n383), .Y(n360) );
  INVX0_HVT U107 ( .A(n354), .Y(n752) );
  INVX1_HVT U108 ( .A(n275), .Y(n464) );
  INVX1_HVT U109 ( .A(in[0]), .Y(n297) );
  INVX1_HVT U111 ( .A(n743), .Y(n560) );
  INVX0_HVT U112 ( .A(n433), .Y(n293) );
  MUX41X1_HVT U113 ( .A1(n736), .A3(n732), .A2(n689), .A4(n523), .S0(n351), 
        .S1(n513), .Y(n688) );
  INVX1_HVT U114 ( .A(n745), .Y(n538) );
  INVX1_HVT U117 ( .A(n445), .Y(n458) );
  NBUFFX2_HVT U118 ( .A(n359), .Y(n383) );
  XOR2X1_HVT U119 ( .A1(n750), .A2(n389), .Y(n734) );
  INVX0_HVT U120 ( .A(n358), .Y(n504) );
  INVX1_HVT U121 ( .A(in[4]), .Y(n326) );
  MUX21X1_HVT U122 ( .A1(n356), .A2(n559), .S0(n394), .Y(n355) );
  INVX1_HVT U124 ( .A(n10), .Y(n418) );
  INVX0_HVT U126 ( .A(n449), .Y(n451) );
  INVX0_HVT U127 ( .A(n440), .Y(n441) );
  INVX1_HVT U128 ( .A(n736), .Y(n362) );
  MUX41X1_HVT U129 ( .A1(n672), .A3(n675), .A2(n674), .A4(n679), .S0(n496), 
        .S1(n408), .Y(n671) );
  MUX21X1_HVT U130 ( .A1(n501), .A2(n521), .S0(n503), .Y(n738) );
  MUX41X1_HVT U131 ( .A1(n475), .A3(n564), .A2(n684), .A4(n557), .S0(n444), 
        .S1(n512), .Y(n683) );
  INVX1_HVT U132 ( .A(n319), .Y(n452) );
  MUX21X1_HVT U133 ( .A1(n612), .A2(n611), .S0(n508), .Y(n610) );
  MUX41X1_HVT U134 ( .A1(n649), .A3(n651), .A2(n650), .A4(n652), .S0(n492), 
        .S1(n469), .Y(n648) );
  INVX0_HVT U135 ( .A(n325), .Y(n51) );
  INVX1_HVT U137 ( .A(n765), .Y(n261) );
  AND2X1_HVT U138 ( .A1(n312), .A2(n313), .Y(n95) );
  MUX41X1_HVT U139 ( .A1(n606), .A3(n759), .A2(n740), .A4(n550), .S0(n426), 
        .S1(n512), .Y(n605) );
  NBUFFX2_HVT U141 ( .A(n498), .Y(n497) );
  MUX41X1_HVT U143 ( .A1(n620), .A3(n473), .A2(n619), .A4(n554), .S0(n242), 
        .S1(n421), .Y(n618) );
  MUX21X1_HVT U144 ( .A1(n320), .A2(n349), .S0(n413), .Y(n568) );
  MUX21X1_HVT U145 ( .A1(n430), .A2(n434), .S0(n503), .Y(n758) );
  INVX1_HVT U146 ( .A(n451), .Y(n453) );
  NAND2X0_HVT U147 ( .A1(n420), .A2(n96), .Y(n113) );
  NAND2X0_HVT U148 ( .A1(n320), .A2(n443), .Y(n114) );
  NAND2X0_HVT U149 ( .A1(n113), .A2(n114), .Y(n407) );
  INVX0_HVT U150 ( .A(n319), .Y(n320) );
  INVX0_HVT U152 ( .A(n504), .Y(n443) );
  INVX0_HVT U155 ( .A(n407), .Y(n768) );
  INVX0_HVT U156 ( .A(n558), .Y(n117) );
  INVX1_HVT U157 ( .A(n484), .Y(n667) );
  NAND2X0_HVT U160 ( .A1(n119), .A2(n96), .Y(n210) );
  NAND2X0_HVT U161 ( .A1(n532), .A2(n332), .Y(n211) );
  NAND2X0_HVT U163 ( .A1(n210), .A2(n211), .Y(n754) );
  INVX1_HVT U164 ( .A(n382), .Y(n321) );
  INVX0_HVT U165 ( .A(n504), .Y(n332) );
  OR2X1_HVT U169 ( .A1(n275), .A2(n532), .Y(n763) );
  INVX1_HVT U170 ( .A(n275), .Y(n505) );
  MUX41X1_HVT U171 ( .A1(n701), .A3(n704), .A2(n703), .A4(n708), .S0(n496), 
        .S1(n408), .Y(n700) );
  MUX41X1_HVT U172 ( .A1(n760), .A3(n694), .A2(n530), .A4(n451), .S0(n487), 
        .S1(n390), .Y(n693) );
  MUX21X1_HVT U173 ( .A1(n532), .A2(n306), .S0(n333), .Y(n354) );
  NBUFFX2_HVT U174 ( .A(n326), .Y(n498) );
  INVX1_HVT U175 ( .A(n338), .Y(n612) );
  MUX21X1_HVT U178 ( .A1(n626), .A2(n625), .S0(n351), .Y(n624) );
  INVX0_HVT U181 ( .A(n769), .Y(n532) );
  MUX21X1_HVT U183 ( .A1(n325), .A2(n534), .S0(n345), .Y(n632) );
  MUX21X2_HVT U184 ( .A1(n759), .A2(n538), .S0(n486), .Y(n649) );
  MUX21X1_HVT U185 ( .A1(n261), .A2(n348), .S0(n490), .Y(n713) );
  MUX41X1_HVT U186 ( .A1(n557), .A3(n2), .A2(n451), .A4(n418), .S0(n512), .S1(
        n353), .Y(n589) );
  NAND2X0_HVT U187 ( .A1(n715), .A2(n365), .Y(n213) );
  NAND2X0_HVT U188 ( .A1(n717), .A2(n314), .Y(n216) );
  NAND2X0_HVT U190 ( .A1(n213), .A2(n216), .Y(n714) );
  INVX0_HVT U191 ( .A(n764), .Y(n217) );
  INVX1_HVT U192 ( .A(n272), .Y(n764) );
  INVX0_HVT U193 ( .A(n739), .Y(n541) );
  INVX0_HVT U195 ( .A(n771), .Y(n543) );
  MUX41X1_HVT U196 ( .A1(n616), .A3(n610), .A2(n618), .A4(n613), .S0(n297), 
        .S1(n408), .Y(n609) );
  MUX41X1_HVT U198 ( .A1(n648), .A3(n653), .A2(n661), .A4(n667), .S0(n496), 
        .S1(in[6]), .Y(out[3]) );
  MUX41X1_HVT U199 ( .A1(n635), .A3(n634), .A2(n639), .A4(n638), .S0(n429), 
        .S1(n496), .Y(n633) );
  MUX41X1_HVT U200 ( .A1(n538), .A3(n540), .A2(n640), .A4(n752), .S0(n218), 
        .S1(n353), .Y(n639) );
  NAND2X0_HVT U201 ( .A1(n532), .A2(n219), .Y(n231) );
  NAND2X0_HVT U202 ( .A1(n434), .A2(n332), .Y(n232) );
  MUX21X2_HVT U204 ( .A1(n274), .A2(n430), .S0(n414), .Y(n759) );
  MUX41X1_HVT U205 ( .A1(n559), .A3(n549), .A2(n437), .A4(n378), .S0(n242), 
        .S1(n390), .Y(n579) );
  NAND2X0_HVT U206 ( .A1(n747), .A2(n489), .Y(n234) );
  NAND2X0_HVT U207 ( .A1(n553), .A2(n365), .Y(n236) );
  NAND2X0_HVT U209 ( .A1(n234), .A2(n236), .Y(n652) );
  MUX41X1_HVT U210 ( .A1(n688), .A3(n683), .A2(n685), .A4(n682), .S0(n297), 
        .S1(n309), .Y(n681) );
  NBUFFX2_HVT U211 ( .A(n384), .Y(n306) );
  NAND2X0_HVT U213 ( .A1(n473), .A2(n444), .Y(n238) );
  NAND2X0_HVT U216 ( .A1(n360), .A2(n489), .Y(n240) );
  NAND2X0_HVT U217 ( .A1(n238), .A2(n240), .Y(n650) );
  INVX1_HVT U219 ( .A(n375), .Y(n430) );
  MUX21X2_HVT U221 ( .A1(n584), .A2(n583), .S0(n353), .Y(n582) );
  INVX1_HVT U222 ( .A(n449), .Y(n318) );
  INVX1_HVT U223 ( .A(n318), .Y(n319) );
  MUX21X1_HVT U224 ( .A1(n497), .A2(n320), .S0(n332), .Y(n702) );
  INVX1_HVT U225 ( .A(n272), .Y(n352) );
  MUX41X1_HVT U226 ( .A1(n642), .A3(n644), .A2(n645), .A4(n646), .S0(n408), 
        .S1(n496), .Y(n641) );
  INVX1_HVT U227 ( .A(n483), .Y(n446) );
  NAND2X0_HVT U228 ( .A1(n433), .A2(n246), .Y(n255) );
  NAND2X0_HVT U229 ( .A1(n501), .A2(n406), .Y(n256) );
  NAND2X0_HVT U230 ( .A1(n255), .A2(n256), .Y(n765) );
  INVX1_HVT U231 ( .A(n406), .Y(n246) );
  INVX0_HVT U232 ( .A(n441), .Y(n406) );
  MUX41X1_HVT U233 ( .A1(n607), .A3(n604), .A2(n605), .A4(n603), .S0(n297), 
        .S1(n429), .Y(n602) );
  NAND2X0_HVT U234 ( .A1(n436), .A2(n505), .Y(n258) );
  NAND2X0_HVT U235 ( .A1(n293), .A2(n246), .Y(n259) );
  NAND2X0_HVT U236 ( .A1(n258), .A2(n259), .Y(n473) );
  XOR2X1_HVT U237 ( .A1(n508), .A2(n468), .Y(n731) );
  INVX0_HVT U238 ( .A(n771), .Y(n435) );
  INVX0_HVT U239 ( .A(n740), .Y(n540) );
  INVX0_HVT U240 ( .A(n317), .Y(n482) );
  INVX1_HVT U242 ( .A(in[2]), .Y(n510) );
  NAND2X0_HVT U243 ( .A1(n489), .A2(n2), .Y(n264) );
  NAND2X0_HVT U244 ( .A1(n264), .A2(n537), .Y(n485) );
  MUX21X1_HVT U246 ( .A1(n419), .A2(n435), .S0(n503), .Y(n740) );
  INVX0_HVT U247 ( .A(n416), .Y(n417) );
  INVX1_HVT U248 ( .A(n321), .Y(n439) );
  INVX1_HVT U249 ( .A(n419), .Y(n420) );
  MUX41X1_HVT U250 ( .A1(n533), .A3(n325), .A2(n770), .A4(n750), .S0(n487), 
        .S1(n470), .Y(n645) );
  AND2X1_HVT U252 ( .A1(n763), .A2(n415), .Y(n272) );
  INVX1_HVT U253 ( .A(n741), .Y(n551) );
  INVX1_HVT U254 ( .A(n769), .Y(n449) );
  INVX1_HVT U255 ( .A(n506), .Y(n282) );
  MUX41X1_HVT U257 ( .A1(n598), .A3(n601), .A2(n594), .A4(n597), .S0(n492), 
        .S1(n297), .Y(n593) );
  MUX21X1_HVT U258 ( .A1(n432), .A2(n418), .S0(n414), .Y(n686) );
  INVX1_HVT U259 ( .A(in[3]), .Y(n438) );
  INVX0_HVT U260 ( .A(n413), .Y(n283) );
  INVX0_HVT U261 ( .A(n441), .Y(n413) );
  INVX0_HVT U262 ( .A(n10), .Y(n415) );
  NAND2X0_HVT U263 ( .A1(n387), .A2(n490), .Y(n285) );
  NAND2X0_HVT U264 ( .A1(n285), .A2(n286), .Y(n712) );
  MUX21X1_HVT U266 ( .A1(n388), .A2(n415), .S0(n503), .Y(n387) );
  INVX0_HVT U267 ( .A(n705), .Y(n561) );
  INVX0_HVT U269 ( .A(n387), .Y(n766) );
  MUX21X2_HVT U271 ( .A1(n274), .A2(n419), .S0(n463), .Y(n741) );
  INVX1_HVT U272 ( .A(n438), .Y(n322) );
  MUX21X1_HVT U273 ( .A1(n119), .A2(n430), .S0(n96), .Y(n572) );
  INVX1_HVT U274 ( .A(n565), .Y(n549) );
  INVX1_HVT U275 ( .A(in[1]), .Y(n506) );
  INVX0_HVT U276 ( .A(n441), .Y(n463) );
  INVX0_HVT U277 ( .A(n435), .Y(n436) );
  MUX41X1_HVT U279 ( .A1(n589), .A3(n591), .A2(n586), .A4(n590), .S0(n496), 
        .S1(n429), .Y(n585) );
  INVX0_HVT U280 ( .A(n749), .Y(n553) );
  MUX21X1_HVT U281 ( .A1(n500), .A2(n274), .S0(n282), .Y(n747) );
  OA21X1_HVT U282 ( .A1(n445), .A2(n743), .A3(n530), .Y(n599) );
  MUX41X1_HVT U283 ( .A1(n558), .A3(n522), .A2(n732), .A4(n286), .S0(n445), 
        .S1(n489), .Y(n634) );
  MUX41X1_HVT U286 ( .A1(n714), .A3(n724), .A2(n710), .A4(n718), .S0(n323), 
        .S1(n297), .Y(out[0]) );
  NAND2X0_HVT U287 ( .A1(n719), .A2(n444), .Y(n300) );
  NAND2X0_HVT U288 ( .A1(n721), .A2(n487), .Y(n303) );
  NAND2X0_HVT U290 ( .A1(n300), .A2(n303), .Y(n718) );
  INVX1_HVT U291 ( .A(n532), .Y(n450) );
  INVX0_HVT U292 ( .A(n419), .Y(n416) );
  MUX41X1_HVT U293 ( .A1(n762), .A3(n525), .A2(n564), .A4(n733), .S0(n218), 
        .S1(n351), .Y(n695) );
  NAND2X0_HVT U294 ( .A1(n350), .A2(n219), .Y(n304) );
  NAND2X0_HVT U297 ( .A1(n339), .A2(n283), .Y(n305) );
  NAND2X0_HVT U298 ( .A1(n304), .A2(n305), .Y(n762) );
  INVX1_HVT U299 ( .A(n567), .Y(n522) );
  MUX41X1_HVT U301 ( .A1(n360), .A3(n455), .A2(n476), .A4(n554), .S0(n469), 
        .S1(n309), .Y(n717) );
  INVX0_HVT U302 ( .A(n756), .Y(n525) );
  NAND2X0_HVT U303 ( .A1(n772), .A2(n314), .Y(n310) );
  NAND2X0_HVT U304 ( .A1(n643), .A2(n242), .Y(n311) );
  NAND2X0_HVT U305 ( .A1(n310), .A2(n311), .Y(n642) );
  NBUFFX2_HVT U307 ( .A(n509), .Y(n489) );
  NBUFFX2_HVT U308 ( .A(n509), .Y(n488) );
  NAND2X0_HVT U310 ( .A1(n436), .A2(n283), .Y(n312) );
  NAND2X0_HVT U311 ( .A1(n388), .A2(n219), .Y(n313) );
  NAND2X0_HVT U312 ( .A1(n312), .A2(n313), .Y(n767) );
  INVX1_HVT U313 ( .A(n324), .Y(n707) );
  NAND2X0_HVT U314 ( .A1(n587), .A2(n314), .Y(n315) );
  NAND2X0_HVT U315 ( .A1(n588), .A2(n242), .Y(n316) );
  NAND2X0_HVT U316 ( .A1(n315), .A2(n316), .Y(n586) );
  INVX0_HVT U317 ( .A(n353), .Y(n314) );
  MUX21X1_HVT U318 ( .A1(n550), .A2(n362), .S0(n390), .Y(n588) );
  NAND2X0_HVT U319 ( .A1(n439), .A2(n498), .Y(n317) );
  INVX1_HVT U320 ( .A(n773), .Y(n527) );
  INVX1_HVT U321 ( .A(n573), .Y(n557) );
  NAND2X0_HVT U322 ( .A1(n367), .A2(n368), .Y(out[1]) );
  INVX1_HVT U323 ( .A(n774), .Y(n419) );
  INVX1_HVT U324 ( .A(n412), .Y(n323) );
  INVX1_HVT U325 ( .A(in[6]), .Y(n412) );
  MUX21X1_HVT U326 ( .A1(n399), .A2(n349), .S0(n441), .Y(n324) );
  MUX41X1_HVT U327 ( .A1(n720), .A3(n479), .A2(n537), .A4(n477), .S0(n445), 
        .S1(n491), .Y(n719) );
  NBUFFX2_HVT U328 ( .A(n763), .Y(n327) );
  NAND2X0_HVT U329 ( .A1(n406), .A2(n416), .Y(n705) );
  OA21X1_HVT U330 ( .A1(n768), .A2(n389), .A3(n540), .Y(n583) );
  NAND2X0_HVT U331 ( .A1(n10), .A2(n414), .Y(n328) );
  NAND2X0_HVT U332 ( .A1(n342), .A2(n521), .Y(n329) );
  NAND2X0_HVT U333 ( .A1(n328), .A2(n329), .Y(n750) );
  INVX0_HVT U334 ( .A(n413), .Y(n342) );
  MUX21X1_HVT U335 ( .A1(n119), .A2(n521), .S0(n441), .Y(n757) );
  MUX41X1_HVT U336 ( .A1(n354), .A3(n556), .A2(n411), .A4(n558), .S0(n390), 
        .S1(n394), .Y(n703) );
  INVX1_HVT U337 ( .A(n494), .Y(n390) );
  OR2X1_HVT U338 ( .A1(n332), .A2(n482), .Y(n773) );
  NAND2X0_HVT U339 ( .A1(n293), .A2(n283), .Y(n330) );
  NAND2X0_HVT U340 ( .A1(n274), .A2(n464), .Y(n331) );
  NAND2X0_HVT U341 ( .A1(n330), .A2(n331), .Y(n745) );
  NAND2X0_HVT U342 ( .A1(n337), .A2(n336), .Y(out[2]) );
  NBUFFX2_HVT U343 ( .A(n504), .Y(n333) );
  MUX41X1_HVT U344 ( .A1(n547), .A3(n523), .A2(n525), .A4(n518), .S0(n218), 
        .S1(n491), .Y(n729) );
  MUX41X1_HVT U345 ( .A1(n757), .A3(n535), .A2(n766), .A4(n723), .S0(n421), 
        .S1(n491), .Y(n721) );
  NAND2X0_HVT U346 ( .A1(n773), .A2(n487), .Y(n334) );
  NAND2X0_HVT U347 ( .A1(n551), .A2(n394), .Y(n335) );
  INVX1_HVT U348 ( .A(n345), .Y(n391) );
  INVX1_HVT U349 ( .A(n322), .Y(n563) );
  MUX41X1_HVT U350 ( .A1(n702), .A3(n534), .A2(n767), .A4(n544), .S0(n493), 
        .S1(n351), .Y(n701) );
  INVX0_HVT U351 ( .A(n686), .Y(n544) );
  INVX0_HVT U352 ( .A(n754), .Y(n530) );
  NAND2X0_HVT U353 ( .A1(n681), .A2(n323), .Y(n336) );
  NAND2X0_HVT U354 ( .A1(n671), .A2(n412), .Y(n337) );
  INVX0_HVT U355 ( .A(n425), .Y(n685) );
  INVX0_HVT U356 ( .A(n430), .Y(n431) );
  INVX1_HVT U357 ( .A(n482), .Y(n339) );
  NAND2X0_HVT U358 ( .A1(n502), .A2(n283), .Y(n340) );
  NAND2X0_HVT U359 ( .A1(n454), .A2(n464), .Y(n341) );
  NAND2X0_HVT U360 ( .A1(n340), .A2(n341), .Y(n737) );
  MUX21X1_HVT U361 ( .A1(n274), .A2(n420), .S0(n342), .Y(n749) );
  NAND2X0_HVT U362 ( .A1(n699), .A2(n242), .Y(n343) );
  NAND2X0_HVT U363 ( .A1(n698), .A2(n488), .Y(n344) );
  NAND2X0_HVT U364 ( .A1(n343), .A2(n344), .Y(n696) );
  MUX21X1_HVT U365 ( .A1(n399), .A2(n502), .S0(n505), .Y(n756) );
  NAND2X0_HVT U366 ( .A1(n394), .A2(n559), .Y(n395) );
  INVX0_HVT U367 ( .A(n357), .Y(n748) );
  MUX41X1_HVT U368 ( .A1(n739), .A3(n475), .A2(n732), .A4(n286), .S0(n365), 
        .S1(n514), .Y(n597) );
  INVX1_HVT U369 ( .A(n450), .Y(n454) );
  NAND2X0_HVT U370 ( .A1(n381), .A2(n464), .Y(n346) );
  NAND2X0_HVT U371 ( .A1(n774), .A2(n443), .Y(n347) );
  NAND2X0_HVT U372 ( .A1(n347), .A2(n346), .Y(n746) );
  INVX0_HVT U373 ( .A(n361), .Y(n591) );
  NBUFFX2_HVT U374 ( .A(n507), .Y(n348) );
  INVX0_HVT U375 ( .A(n762), .Y(n526) );
  INVX0_HVT U376 ( .A(n375), .Y(n349) );
  MUX41X1_HVT U377 ( .A1(n751), .A3(n707), .A2(n753), .A4(n706), .S0(n426), 
        .S1(n469), .Y(n704) );
  MUX41X1_HVT U378 ( .A1(n352), .A3(n723), .A2(n754), .A4(n560), .S0(n242), 
        .S1(n468), .Y(n580) );
  INVX1_HVT U379 ( .A(n571), .Y(n534) );
  INVX1_HVT U380 ( .A(n572), .Y(n556) );
  INVX1_HVT U381 ( .A(n592), .Y(n364) );
  INVX0_HVT U382 ( .A(n670), .Y(n356) );
  NAND2X0_HVT U383 ( .A1(n404), .A2(n405), .Y(out[4]) );
  MUX21X1_HVT U384 ( .A1(n399), .A2(n433), .S0(n464), .Y(n357) );
  INVX1_HVT U385 ( .A(n506), .Y(n440) );
  INVX0_HVT U386 ( .A(n308), .Y(n426) );
  OR2X1_HVT U387 ( .A1(n399), .A2(n333), .Y(n742) );
  INVX0_HVT U388 ( .A(n759), .Y(n554) );
  INVX1_HVT U389 ( .A(n575), .Y(n523) );
  XOR2X2_HVT U390 ( .A1(n452), .A2(n463), .Y(n732) );
  INVX1_HVT U391 ( .A(n501), .Y(n388) );
  MUX41X1_HVT U392 ( .A1(n363), .A3(n362), .A2(n364), .A4(n366), .S0(n365), 
        .S1(n513), .Y(n361) );
  XNOR2X1_HVT U393 ( .A1(n306), .A2(n464), .Y(n366) );
  NAND2X0_HVT U394 ( .A1(n700), .A2(n323), .Y(n367) );
  NAND2X0_HVT U395 ( .A1(n690), .A2(n412), .Y(n368) );
  NAND2X0_HVT U396 ( .A1(n517), .A2(n394), .Y(n369) );
  NAND2X0_HVT U397 ( .A1(n647), .A2(n489), .Y(n370) );
  NAND2X0_HVT U398 ( .A1(n369), .A2(n370), .Y(n646) );
  MUX21X1_HVT U399 ( .A1(n428), .A2(n427), .S0(n314), .Y(n425) );
  NAND2X0_HVT U400 ( .A1(n602), .A2(n323), .Y(n397) );
  NAND2X0_HVT U401 ( .A1(n541), .A2(n469), .Y(n371) );
  NAND2X0_HVT U402 ( .A1(n754), .A2(n421), .Y(n372) );
  NAND2X0_HVT U403 ( .A1(n371), .A2(n372), .Y(n643) );
  NAND2X0_HVT U404 ( .A1(n544), .A2(n469), .Y(n373) );
  NAND2X0_HVT U405 ( .A1(n740), .A2(n421), .Y(n374) );
  NAND2X0_HVT U406 ( .A1(n373), .A2(n374), .Y(n625) );
  NAND2X0_HVT U407 ( .A1(n467), .A2(n563), .Y(n375) );
  OA21X1_HVT U408 ( .A1(n520), .A2(n389), .A3(n746), .Y(n636) );
  XOR2X2_HVT U409 ( .A1(n326), .A2(n382), .Y(n769) );
  NBUFFX2_HVT U410 ( .A(n509), .Y(n487) );
  INVX0_HVT U411 ( .A(n668), .Y(n481) );
  NAND2X0_HVT U412 ( .A1(n709), .A2(n314), .Y(n376) );
  NAND2X0_HVT U413 ( .A1(n734), .A2(n444), .Y(n377) );
  NAND2X0_HVT U414 ( .A1(n376), .A2(n377), .Y(n708) );
  NBUFFX2_HVT U415 ( .A(n399), .Y(n378) );
  NAND2X0_HVT U416 ( .A1(n379), .A2(n469), .Y(n380) );
  AND2X1_HVT U417 ( .A1(n380), .A2(n746), .Y(n611) );
  INVX0_HVT U418 ( .A(n477), .Y(n379) );
  NAND2X0_HVT U419 ( .A1(n467), .A2(n321), .Y(n381) );
  NAND2X0_HVT U420 ( .A1(n439), .A2(n498), .Y(n384) );
  NAND2X0_HVT U421 ( .A1(n350), .A2(n494), .Y(n385) );
  NAND2X0_HVT U422 ( .A1(n542), .A2(n390), .Y(n386) );
  NAND2X0_HVT U423 ( .A1(n385), .A2(n386), .Y(n647) );
  NAND2X0_HVT U424 ( .A1(n658), .A2(n391), .Y(n392) );
  NAND2X0_HVT U425 ( .A1(n659), .A2(n421), .Y(n393) );
  NAND2X0_HVT U426 ( .A1(n392), .A2(n393), .Y(n655) );
  MUX21X1_HVT U427 ( .A1(n539), .A2(n660), .S0(n308), .Y(n659) );
  NAND2X0_HVT U428 ( .A1(n487), .A2(n762), .Y(n396) );
  NAND2X0_HVT U429 ( .A1(n396), .A2(n395), .Y(n680) );
  NAND2X0_HVT U430 ( .A1(n593), .A2(n412), .Y(n398) );
  NAND2X0_HVT U431 ( .A1(n397), .A2(n398), .Y(out[6]) );
  MUX41X1_HVT U432 ( .A1(n624), .A3(n622), .A2(n629), .A4(n628), .S0(n309), 
        .S1(n496), .Y(n621) );
  NAND2X0_HVT U433 ( .A1(n578), .A2(n412), .Y(n400) );
  NAND2X0_HVT U434 ( .A1(n585), .A2(n323), .Y(n401) );
  NAND2X0_HVT U435 ( .A1(n400), .A2(n401), .Y(out[7]) );
  NAND2X0_HVT U436 ( .A1(n727), .A2(n218), .Y(n402) );
  NAND2X0_HVT U437 ( .A1(n728), .A2(n493), .Y(n403) );
  NAND2X0_HVT U438 ( .A1(n403), .A2(n402), .Y(n725) );
  MUX21X1_HVT U439 ( .A1(n388), .A2(n742), .S0(n492), .Y(n728) );
  NAND2X0_HVT U440 ( .A1(n633), .A2(n412), .Y(n404) );
  NAND2X0_HVT U441 ( .A1(n641), .A2(n323), .Y(n405) );
  MUX21X1_HVT U442 ( .A1(n381), .A2(n274), .S0(n246), .Y(n566) );
  NAND2X0_HVT U443 ( .A1(n665), .A2(n408), .Y(n409) );
  NAND2X0_HVT U444 ( .A1(n662), .A2(n429), .Y(n410) );
  NAND2X0_HVT U445 ( .A1(n409), .A2(n410), .Y(n661) );
  MUX41X1_HVT U446 ( .A1(n695), .A3(n691), .A2(n696), .A4(n693), .S0(n297), 
        .S1(n490), .Y(n690) );
  MUX41X1_HVT U447 ( .A1(n582), .A3(n580), .A2(n581), .A4(n579), .S0(n297), 
        .S1(n429), .Y(n578) );
  INVX1_HVT U448 ( .A(n566), .Y(n550) );
  NAND2X0_HVT U449 ( .A1(n502), .A2(n422), .Y(n423) );
  NAND2X0_HVT U450 ( .A1(n687), .A2(n478), .Y(n424) );
  INVX0_HVT U451 ( .A(n478), .Y(n422) );
  AND2X1_HVT U452 ( .A1(n423), .A2(n424), .Y(n427) );
  AOI21X1_HVT U453 ( .A1(n686), .A2(n495), .A3(n555), .Y(n428) );
  INVX1_HVT U454 ( .A(n758), .Y(n537) );
  INVX1_HVT U455 ( .A(n527), .Y(n437) );
  INVX1_HVT U456 ( .A(n570), .Y(n517) );
  INVX1_HVT U457 ( .A(n569), .Y(n542) );
  MUX21X1_HVT U458 ( .A1(n10), .A2(n500), .S0(n383), .Y(n743) );
  INVX1_HVT U459 ( .A(n568), .Y(n533) );
  MUX21X1_HVT U460 ( .A1(n502), .A2(n431), .S0(n283), .Y(n442) );
  MUX41X1_HVT U461 ( .A1(n617), .A3(n732), .A2(n552), .A4(n755), .S0(n421), 
        .S1(n444), .Y(n616) );
  MUX21X1_HVT U462 ( .A1(n417), .A2(n557), .S0(n495), .Y(n709) );
  NAND2X0_HVT U463 ( .A1(n482), .A2(n446), .Y(n447) );
  NAND2X0_HVT U464 ( .A1(n481), .A2(n483), .Y(n448) );
  NAND2X0_HVT U465 ( .A1(n447), .A2(n448), .Y(n480) );
  INVX1_HVT U466 ( .A(n450), .Y(n455) );
  NAND2X0_HVT U467 ( .A1(n654), .A2(n309), .Y(n456) );
  NAND2X0_HVT U468 ( .A1(n655), .A2(n490), .Y(n457) );
  NAND2X0_HVT U469 ( .A1(n456), .A2(n457), .Y(n653) );
  NAND2X0_HVT U470 ( .A1(n471), .A2(n458), .Y(n459) );
  NAND2X0_HVT U471 ( .A1(n760), .A2(n345), .Y(n460) );
  NAND2X0_HVT U472 ( .A1(n459), .A2(n460), .Y(n584) );
  NAND2X0_HVT U473 ( .A1(n466), .A2(n465), .Y(out[5]) );
  NAND2X0_HVT U474 ( .A1(n627), .A2(n422), .Y(n461) );
  NAND2X0_HVT U475 ( .A1(n384), .A2(n478), .Y(n462) );
  NAND2X0_HVT U476 ( .A1(n461), .A2(n462), .Y(n626) );
  NAND2X0_HVT U477 ( .A1(n609), .A2(n412), .Y(n465) );
  NAND2X0_HVT U478 ( .A1(n621), .A2(n323), .Y(n466) );
  NBUFFX2_HVT U479 ( .A(n514), .Y(n468) );
  NBUFFX2_HVT U480 ( .A(n514), .Y(n469) );
  NBUFFX2_HVT U481 ( .A(n514), .Y(n470) );
  AND2X1_HVT U482 ( .A1(n453), .A2(n722), .Y(n471) );
  MUX21X1_HVT U483 ( .A1(n434), .A2(n417), .S0(n492), .Y(n726) );
  AND2X1_HVT U484 ( .A1(n339), .A2(n705), .Y(n472) );
  MUX21X1_HVT U485 ( .A1(n455), .A2(n212), .S0(n464), .Y(n676) );
  MUX21X1_HVT U486 ( .A1(n500), .A2(n450), .S0(n333), .Y(n571) );
  NAND2X0_HVT U487 ( .A1(n498), .A2(n563), .Y(n771) );
  MUX21X1_HVT U488 ( .A1(n434), .A2(n497), .S0(n505), .Y(n569) );
  NBUFFX2_HVT U489 ( .A(n384), .Y(n502) );
  MUX21X1_HVT U490 ( .A1(n497), .A2(n501), .S0(n383), .Y(n660) );
  MUX21X1_HVT U491 ( .A1(n500), .A2(n212), .S0(n413), .Y(n592) );
  MUX21X1_HVT U492 ( .A1(n502), .A2(n436), .S0(n463), .Y(n567) );
  MUX21X1_HVT U493 ( .A1(n306), .A2(n497), .S0(n333), .Y(n575) );
  AND2X1_HVT U494 ( .A1(n383), .A2(n411), .Y(n475) );
  MUX21X1_HVT U495 ( .A1(n350), .A2(n500), .S0(n414), .Y(n573) );
  AND2X1_HVT U496 ( .A1(n415), .A2(n669), .Y(n476) );
  MUX21X1_HVT U497 ( .A1(n350), .A2(n415), .S0(n307), .Y(n657) );
  XOR2X1_HVT U498 ( .A1(n497), .A2(n464), .Y(n751) );
  NBUFFX2_HVT U499 ( .A(n509), .Y(n486) );
  NBUFFX2_HVT U500 ( .A(n563), .Y(n500) );
  NBUFFX2_HVT U501 ( .A(n563), .Y(n501) );
  NBUFFX2_HVT U502 ( .A(n515), .Y(n494) );
  NBUFFX2_HVT U503 ( .A(n515), .Y(n495) );
  NBUFFX2_HVT U504 ( .A(n511), .Y(n492) );
  NBUFFX2_HVT U505 ( .A(n511), .Y(n491) );
  NBUFFX2_HVT U506 ( .A(n511), .Y(n490) );
  MUX21X1_HVT U507 ( .A1(n692), .A2(n119), .S0(n494), .Y(n600) );
  MUX21X1_HVT U508 ( .A1(n678), .A2(n517), .S0(n488), .Y(n675) );
  XOR2X1_HVT U509 ( .A1(n406), .A2(n119), .Y(n730) );
  AND2X1_HVT U510 ( .A1(n455), .A2(n507), .Y(n477) );
  MUX21X1_HVT U511 ( .A1(n388), .A2(n293), .S0(n505), .Y(n739) );
  XOR2X1_HVT U512 ( .A1(n406), .A2(n492), .Y(n735) );
  MUX21X1_HVT U513 ( .A1(n437), .A2(n348), .S0(n488), .Y(n656) );
  MUX21X1_HVT U514 ( .A1(n388), .A2(n212), .S0(n495), .Y(n687) );
  XNOR2X1_HVT U515 ( .A1(n516), .A2(n505), .Y(n478) );
  AND2X1_HVT U516 ( .A1(n501), .A2(n348), .Y(n479) );
  INVX1_HVT U517 ( .A(n516), .Y(n515) );
  NBUFFX2_HVT U518 ( .A(in[5]), .Y(n511) );
  NAND2X0_HVT U519 ( .A1(n439), .A2(n467), .Y(n774) );
  MUX21X1_HVT U520 ( .A1(n563), .A2(n420), .S0(n505), .Y(n595) );
  MUX21X1_HVT U521 ( .A1(n274), .A2(n451), .S0(n503), .Y(n574) );
  MUX21X1_HVT U522 ( .A1(n274), .A2(n418), .S0(n96), .Y(n565) );
  MUX21X1_HVT U523 ( .A1(n388), .A2(n378), .S0(n509), .Y(n668) );
  MUX41X1_HVT U524 ( .A1(n355), .A3(n485), .A2(n480), .A4(n50), .S0(n492), 
        .S1(n421), .Y(n484) );
endmodule

