
module inv_sbox_12 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n103, n196, n197, n198, n199, n200, n201, n202, n206, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623;

  NAND2X0_HVT U1 ( .A1(in[3]), .A2(n330), .Y(n623) );
  NAND2X0_HVT U4 ( .A1(n349), .A2(n201), .Y(n620) );
  NAND2X0_HVT U5 ( .A1(n620), .A2(n340), .Y(n619) );
  NAND2X0_HVT U8 ( .A1(n282), .A2(n339), .Y(n615) );
  NAND2X0_HVT U9 ( .A1(n345), .A2(n615), .Y(n614) );
  NAND2X0_HVT U10 ( .A1(n345), .A2(n612), .Y(n613) );
  NAND2X0_HVT U11 ( .A1(n351), .A2(n344), .Y(n611) );
  NAND2X0_HVT U12 ( .A1(n292), .A2(n329), .Y(n610) );
  NAND2X0_HVT U13 ( .A1(n343), .A2(n223), .Y(n609) );
  NAND2X0_HVT U15 ( .A1(n338), .A2(n291), .Y(n607) );
  NAND2X0_HVT U19 ( .A1(n284), .A2(n413), .Y(n602) );
  NAND2X0_HVT U25 ( .A1(n264), .A2(n329), .Y(n618) );
  NAND2X0_HVT U38 ( .A1(n329), .A2(n271), .Y(n584) );
  OA21X1_HVT U53 ( .A1(n358), .A2(n572), .A3(n380), .Y(n570) );
  NAND2X0_HVT U55 ( .A1(n343), .A2(n620), .Y(n568) );
  MUX41X1_HVT U56 ( .A1(n394), .A3(n337), .A2(n378), .A4(n568), .S0(n321), 
        .S1(n354), .Y(n567) );
  MUX41X1_HVT U62 ( .A1(n561), .A3(n567), .A2(n565), .A4(n569), .S0(in[5]), 
        .S1(n333), .Y(n560) );
  MUX41X1_HVT U65 ( .A1(n268), .A3(n374), .A2(n373), .A4(n584), .S0(n321), 
        .S1(n356), .Y(n557) );
  NAND2X0_HVT U66 ( .A1(n290), .A2(n316), .Y(n556) );
  MUX41X1_HVT U67 ( .A1(n303), .A3(n395), .A2(n372), .A4(n556), .S0(n327), 
        .S1(n317), .Y(n555) );
  MUX41X1_HVT U68 ( .A1(n303), .A3(n308), .A2(n371), .A4(n345), .S0(n320), 
        .S1(n356), .Y(n554) );
  MUX41X1_HVT U69 ( .A1(n554), .A3(n557), .A2(n555), .A4(n558), .S0(n336), 
        .S1(n333), .Y(n553) );
  NAND2X0_HVT U72 ( .A1(n337), .A2(n616), .Y(n551) );
  MUX41X1_HVT U73 ( .A1(n231), .A3(n551), .A2(n396), .A4(n328), .S0(n326), 
        .S1(n318), .Y(n550) );
  MUX41X1_HVT U74 ( .A1(n613), .A3(n385), .A2(n384), .A4(n375), .S0(n321), 
        .S1(n300), .Y(n549) );
  MUX41X1_HVT U78 ( .A1(n546), .A3(n550), .A2(n549), .A4(n552), .S0(n336), 
        .S1(n333), .Y(n545) );
  MUX41X1_HVT U79 ( .A1(n381), .A3(n604), .A2(n383), .A4(n605), .S0(n321), 
        .S1(n300), .Y(n544) );
  MUX41X1_HVT U80 ( .A1(n397), .A3(n394), .A2(n614), .A4(n619), .S0(n320), 
        .S1(n355), .Y(n543) );
  NAND2X0_HVT U81 ( .A1(n258), .A2(n616), .Y(n542) );
  AND2X1_HVT U82 ( .A1(n617), .A2(n341), .Y(n541) );
  MUX41X1_HVT U84 ( .A1(n314), .A3(n381), .A2(n399), .A4(n597), .S0(n321), 
        .S1(n356), .Y(n539) );
  MUX41X1_HVT U87 ( .A1(n363), .A3(n314), .A2(n400), .A4(n378), .S0(n319), 
        .S1(n301), .Y(n537) );
  MUX41X1_HVT U88 ( .A1(n372), .A3(n360), .A2(n592), .A4(n576), .S0(n320), 
        .S1(n293), .Y(n536) );
  NAND2X0_HVT U89 ( .A1(n271), .A2(n257), .Y(n535) );
  MUX41X1_HVT U96 ( .A1(n395), .A3(n609), .A2(n379), .A4(n401), .S0(n321), 
        .S1(n354), .Y(n528) );
  MUX41X1_HVT U98 ( .A1(n527), .A3(n402), .A2(n387), .A4(n594), .S0(n321), 
        .S1(n300), .Y(n526) );
  MUX41X1_HVT U99 ( .A1(n590), .A3(n373), .A2(n574), .A4(n337), .S0(n356), 
        .S1(n317), .Y(n525) );
  NAND2X0_HVT U100 ( .A1(n351), .A2(n409), .Y(n524) );
  MUX41X1_HVT U101 ( .A1(n403), .A3(n610), .A2(n386), .A4(n524), .S0(n356), 
        .S1(n317), .Y(n523) );
  MUX41X1_HVT U107 ( .A1(n403), .A3(n341), .A2(n520), .A4(n365), .S0(n320), 
        .S1(n301), .Y(n519) );
  MUX41X1_HVT U108 ( .A1(n259), .A3(n337), .A2(n378), .A4(n258), .S0(n321), 
        .S1(n354), .Y(n518) );
  MUX41X1_HVT U109 ( .A1(n402), .A3(n360), .A2(n399), .A4(n392), .S0(n320), 
        .S1(n300), .Y(n517) );
  AO21X1_HVT U112 ( .A1(n389), .A2(n326), .A3(n598), .Y(n514) );
  NAND2X0_HVT U114 ( .A1(n345), .A2(n616), .Y(n512) );
  MUX41X1_HVT U115 ( .A1(n512), .A3(n611), .A2(n389), .A4(n341), .S0(n356), 
        .S1(n318), .Y(n511) );
  MUX41X1_HVT U116 ( .A1(n388), .A3(n381), .A2(n360), .A4(n200), .S0(n319), 
        .S1(n301), .Y(n510) );
  NAND2X0_HVT U118 ( .A1(n271), .A2(n308), .Y(n508) );
  MUX41X1_HVT U119 ( .A1(n405), .A3(n509), .A2(n585), .A4(n508), .S0(n319), 
        .S1(n354), .Y(n507) );
  MUX41X1_HVT U122 ( .A1(n393), .A3(n310), .A2(n576), .A4(n265), .S0(n319), 
        .S1(n293), .Y(n505) );
  MUX41X1_HVT U124 ( .A1(n312), .A3(n504), .A2(n599), .A4(n376), .S0(n325), 
        .S1(n319), .Y(n503) );
  AOI21X1_HVT U127 ( .A1(n324), .A2(n499), .A3(n366), .Y(n500) );
  NAND2X0_HVT U129 ( .A1(n323), .A2(n345), .Y(n497) );
  MUX41X1_HVT U130 ( .A1(n497), .A3(n498), .A2(n501), .A4(n500), .S0(n327), 
        .S1(n334), .Y(n496) );
  AND2X1_HVT U131 ( .A1(n316), .A2(n227), .Y(n495) );
  MUX41X1_HVT U132 ( .A1(n364), .A3(n495), .A2(n407), .A4(n303), .S0(n326), 
        .S1(n318), .Y(n494) );
  MUX41X1_HVT U133 ( .A1(n408), .A3(n365), .A2(n568), .A4(n294), .S0(n325), 
        .S1(n317), .Y(n493) );
  MUX41X1_HVT U136 ( .A1(n573), .A3(n524), .A2(n491), .A4(n369), .S0(n323), 
        .S1(n293), .Y(n490) );
  MUX41X1_HVT U137 ( .A1(n223), .A3(n593), .A2(n597), .A4(n401), .S0(n327), 
        .S1(n317), .Y(n489) );
  MUX41X1_HVT U139 ( .A1(n488), .A3(n492), .A2(n496), .A4(n502), .S0(n336), 
        .S1(n307), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n384), .A3(n311), .A2(n236), .A4(n611), .S0(n326), 
        .S1(n318), .Y(n487) );
  NAND2X0_HVT U141 ( .A1(n337), .A2(n351), .Y(n486) );
  MUX41X1_HVT U142 ( .A1(n486), .A3(n583), .A2(n406), .A4(n236), .S0(n324), 
        .S1(n356), .Y(n485) );
  MUX41X1_HVT U143 ( .A1(n257), .A3(n390), .A2(n602), .A4(n599), .S0(n322), 
        .S1(n300), .Y(n484) );
  MUX41X1_HVT U145 ( .A1(n591), .A3(n404), .A2(n483), .A4(n542), .S0(n324), 
        .S1(n300), .Y(n482) );
  MUX41X1_HVT U146 ( .A1(n482), .A3(n484), .A2(n485), .A4(n487), .S0(n334), 
        .S1(n336), .Y(n481) );
  MUX41X1_HVT U151 ( .A1(n398), .A3(n387), .A2(n252), .A4(n477), .S0(n325), 
        .S1(n317), .Y(n476) );
  MUX41X1_HVT U155 ( .A1(n236), .A3(n611), .A2(n603), .A4(n379), .S0(n322), 
        .S1(n301), .Y(n472) );
  MUX41X1_HVT U156 ( .A1(n472), .A3(n476), .A2(n473), .A4(n478), .S0(n336), 
        .S1(n334), .Y(n471) );
  NAND2X0_HVT U159 ( .A1(n468), .A2(n467), .Y(n469) );
  MUX41X1_HVT U162 ( .A1(n286), .A3(n374), .A2(n587), .A4(n465), .S0(n322), 
        .S1(n300), .Y(n464) );
  NAND2X0_HVT U163 ( .A1(n292), .A2(n257), .Y(n463) );
  MUX41X1_HVT U164 ( .A1(n614), .A3(n463), .A2(n585), .A4(n259), .S0(n319), 
        .S1(n354), .Y(n462) );
  NAND2X0_HVT U166 ( .A1(n612), .A2(n459), .Y(n460) );
  MUX41X1_HVT U170 ( .A1(n313), .A3(n309), .A2(n312), .A4(n456), .S0(n322), 
        .S1(n301), .Y(n455) );
  MUX41X1_HVT U172 ( .A1(n535), .A3(n454), .A2(n309), .A4(n600), .S0(n322), 
        .S1(n301), .Y(n453) );
  MUX41X1_HVT U173 ( .A1(n345), .A3(n412), .A2(n258), .A4(n586), .S0(n322), 
        .S1(n356), .Y(n452) );
  MUX41X1_HVT U174 ( .A1(n400), .A3(n568), .A2(n408), .A4(n414), .S0(n322), 
        .S1(n300), .Y(n451) );
  NAND2X0_HVT U177 ( .A1(n284), .A2(n308), .Y(n449) );
  MUX41X1_HVT U178 ( .A1(n313), .A3(n449), .A2(n412), .A4(n578), .S0(n322), 
        .S1(n354), .Y(n448) );
  AND2X1_HVT U179 ( .A1(n617), .A2(n340), .Y(n447) );
  MUX41X1_HVT U180 ( .A1(n590), .A3(n359), .A2(n447), .A4(n577), .S0(n322), 
        .S1(n354), .Y(n446) );
  AND2X1_HVT U185 ( .A1(n414), .A2(n350), .Y(n441) );
  NAND2X0_HVT U191 ( .A1(n358), .A2(n370), .Y(n435) );
  AND2X1_HVT U192 ( .A1(n385), .A2(n433), .Y(n434) );
  NAND2X0_HVT U194 ( .A1(n580), .A2(n433), .Y(n431) );
  MUX41X1_HVT U195 ( .A1(n432), .A3(n431), .A2(n434), .A4(n435), .S0(n320), 
        .S1(n334), .Y(n430) );
  NAND2X0_HVT U198 ( .A1(n284), .A2(n414), .Y(n612) );
  NAND2X0_HVT U200 ( .A1(n340), .A2(n271), .Y(n499) );
  NAND2X0_HVT U207 ( .A1(n271), .A2(n412), .Y(n562) );
  INVX1_HVT U2 ( .A(n350), .Y(n291) );
  NBUFFX2_HVT U3 ( .A(n411), .Y(n329) );
  XNOR2X1_HVT U6 ( .A1(n415), .A2(n411), .Y(n606) );
  NBUFFX2_HVT U7 ( .A(n411), .Y(n328) );
  MUX21X1_HVT U14 ( .A1(n265), .A2(n579), .S0(n287), .Y(n470) );
  INVX1_HVT U16 ( .A(n417), .Y(n407) );
  XNOR2X1_HVT U17 ( .A1(n410), .A2(n349), .Y(n574) );
  INVX1_HVT U18 ( .A(n579), .Y(n390) );
  INVX1_HVT U20 ( .A(n618), .Y(n257) );
  IBUFFX2_HVT U21 ( .A(n605), .Y(n372) );
  MUX21X2_HVT U22 ( .A1(n314), .A2(n574), .S0(n327), .Y(n439) );
  OA21X2_HVT U23 ( .A1(n362), .A2(n358), .A3(n601), .Y(n547) );
  MUX21X1_HVT U24 ( .A1(n413), .A2(n316), .S0(n227), .Y(n581) );
  IBUFFX2_HVT U26 ( .A(n350), .Y(n348) );
  NAND2X0_HVT U27 ( .A1(n308), .A2(n103), .Y(n196) );
  NAND2X0_HVT U28 ( .A1(n409), .A2(n260), .Y(n197) );
  NAND2X0_HVT U29 ( .A1(n196), .A2(n197), .Y(n599) );
  INVX0_HVT U30 ( .A(n260), .Y(n103) );
  NBUFFX2_HVT U31 ( .A(n415), .Y(n330) );
  INVX0_HVT U32 ( .A(n415), .Y(n316) );
  MUX21X2_HVT U33 ( .A1(n329), .A2(n338), .S0(n227), .Y(n601) );
  MUX21X1_HVT U34 ( .A1(n375), .A2(n559), .S0(n315), .Y(n558) );
  AO21X2_HVT U35 ( .A1(n562), .A2(n325), .A3(n601), .Y(n563) );
  MUX21X1_HVT U36 ( .A1(n308), .A2(n331), .S0(n256), .Y(n595) );
  IBUFFX2_HVT U37 ( .A(n350), .Y(n347) );
  INVX0_HVT U39 ( .A(n285), .Y(n256) );
  NAND2X0_HVT U40 ( .A1(n348), .A2(n342), .Y(n616) );
  IBUFFX2_HVT U41 ( .A(n263), .Y(n248) );
  INVX1_HVT U42 ( .A(n580), .Y(n365) );
  MUX41X1_HVT U43 ( .A1(n528), .A3(n525), .A2(n526), .A4(n523), .S0(n198), 
        .S1(n199), .Y(n522) );
  IBUFFX16_HVT U44 ( .A(n336), .Y(n198) );
  IBUFFX16_HVT U45 ( .A(n333), .Y(n199) );
  MUX21X2_HVT U46 ( .A1(n460), .A2(n461), .S0(n323), .Y(n458) );
  INVX1_HVT U47 ( .A(in[4]), .Y(n357) );
  INVX0_HVT U48 ( .A(n618), .Y(n410) );
  NOR2X0_HVT U49 ( .A1(n350), .A2(n295), .Y(n294) );
  MUX41X1_HVT U50 ( .A1(n580), .A3(n394), .A2(n375), .A4(n390), .S0(n305), 
        .S1(n298), .Y(n443) );
  INVX2_HVT U51 ( .A(n357), .Y(n300) );
  INVX0_HVT U52 ( .A(n371), .Y(n200) );
  INVX0_HVT U54 ( .A(n607), .Y(n371) );
  INVX0_HVT U57 ( .A(n601), .Y(n259) );
  MUX21X1_HVT U58 ( .A1(n568), .A2(n376), .S0(n222), .Y(n564) );
  INVX0_HVT U59 ( .A(n326), .Y(n222) );
  INVX1_HVT U60 ( .A(n270), .Y(n201) );
  INVX2_HVT U61 ( .A(n622), .Y(n270) );
  NAND2X0_HVT U63 ( .A1(n328), .A2(n415), .Y(n622) );
  MUX41X1_HVT U64 ( .A1(n440), .A3(n439), .A2(n437), .A4(n438), .S0(n202), 
        .S1(n206), .Y(n436) );
  IBUFFX16_HVT U70 ( .A(n318), .Y(n202) );
  IBUFFX16_HVT U71 ( .A(n334), .Y(n206) );
  INVX0_HVT U75 ( .A(n599), .Y(n376) );
  INVX0_HVT U76 ( .A(n327), .Y(n232) );
  INVX0_HVT U77 ( .A(n285), .Y(n227) );
  INVX1_HVT U83 ( .A(n277), .Y(n218) );
  INVX0_HVT U85 ( .A(n330), .Y(n277) );
  NBUFFX2_HVT U86 ( .A(n415), .Y(n331) );
  MUX21X1_HVT U90 ( .A1(n295), .A2(n410), .S0(n291), .Y(n594) );
  MUX21X1_HVT U91 ( .A1(n329), .A2(n330), .S0(n291), .Y(n577) );
  INVX0_HVT U92 ( .A(n595), .Y(n379) );
  MUX21X1_HVT U93 ( .A1(n595), .A2(n607), .S0(n327), .Y(n219) );
  IBUFFX16_HVT U94 ( .A(n219), .Y(n571) );
  IBUFFX2_HVT U95 ( .A(n594), .Y(n380) );
  INVX0_HVT U97 ( .A(n302), .Y(n521) );
  INVX0_HVT U102 ( .A(n268), .Y(n604) );
  INVX0_HVT U103 ( .A(n285), .Y(n260) );
  MUX21X1_HVT U104 ( .A1(n441), .A2(n397), .S0(n325), .Y(n440) );
  INVX1_HVT U105 ( .A(n276), .Y(n590) );
  MUX21X2_HVT U106 ( .A1(n346), .A2(n316), .S0(n271), .Y(n605) );
  IBUFFX2_HVT U110 ( .A(n577), .Y(n391) );
  INVX1_HVT U111 ( .A(n220), .Y(n265) );
  MUX21X1_HVT U113 ( .A1(n265), .A2(n276), .S0(n327), .Y(n548) );
  INVX1_HVT U117 ( .A(n299), .Y(n238) );
  MUX21X2_HVT U120 ( .A1(n269), .A2(n270), .S0(n291), .Y(n268) );
  MUX21X1_HVT U121 ( .A1(n221), .A2(n329), .S0(n290), .Y(n220) );
  IBUFFX16_HVT U123 ( .A(n341), .Y(n221) );
  MUX21X1_HVT U125 ( .A1(n344), .A2(n329), .S0(n260), .Y(n426) );
  IBUFFX2_HVT U126 ( .A(n350), .Y(n292) );
  NOR2X4_HVT U128 ( .A1(n277), .A2(n292), .Y(n276) );
  AO21X2_HVT U134 ( .A1(n337), .A2(n620), .A3(n358), .Y(n459) );
  MUX21X2_HVT U135 ( .A1(n339), .A2(n316), .S0(n282), .Y(n593) );
  INVX0_HVT U138 ( .A(n290), .Y(n243) );
  INVX0_HVT U144 ( .A(n611), .Y(n359) );
  AO21X2_HVT U147 ( .A1(n327), .A2(n367), .A3(n409), .Y(n479) );
  INVX1_HVT U148 ( .A(n367), .Y(n223) );
  INVX0_HVT U149 ( .A(n615), .Y(n367) );
  OR2X1_HVT U150 ( .A1(n294), .A2(n338), .Y(n580) );
  INVX1_HVT U152 ( .A(n294), .Y(n617) );
  NAND2X0_HVT U153 ( .A1(n342), .A2(n224), .Y(n225) );
  NAND2X0_HVT U154 ( .A1(n533), .A2(n275), .Y(n226) );
  NAND2X0_HVT U157 ( .A1(n226), .A2(n225), .Y(n532) );
  INVX0_HVT U158 ( .A(n275), .Y(n224) );
  NBUFFX4_HVT U160 ( .A(n621), .Y(n342) );
  MUX21X1_HVT U161 ( .A1(n338), .A2(n218), .S0(n326), .Y(n533) );
  MUX21X2_HVT U165 ( .A1(n564), .A2(n563), .S0(n323), .Y(n561) );
  NBUFFX16_HVT U167 ( .A(n355), .Y(n326) );
  NAND2X0_HVT U168 ( .A1(n391), .A2(n228), .Y(n229) );
  NAND2X0_HVT U169 ( .A1(n312), .A2(n325), .Y(n230) );
  NAND2X0_HVT U171 ( .A1(n229), .A2(n230), .Y(n432) );
  IBUFFX2_HVT U175 ( .A(n325), .Y(n228) );
  INVX1_HVT U176 ( .A(n601), .Y(n375) );
  NBUFFX2_HVT U181 ( .A(n595), .Y(n231) );
  IBUFFX2_HVT U182 ( .A(n326), .Y(n287) );
  IBUFFX4_HVT U183 ( .A(n326), .Y(n251) );
  MUX21X1_HVT U184 ( .A1(n337), .A2(n237), .S0(n232), .Y(n531) );
  IBUFFX2_HVT U186 ( .A(n237), .Y(n587) );
  NAND2X0_HVT U187 ( .A1(n377), .A2(n233), .Y(n234) );
  NAND2X0_HVT U188 ( .A1(n566), .A2(n315), .Y(n235) );
  NAND2X0_HVT U189 ( .A1(n234), .A2(n235), .Y(n565) );
  INVX0_HVT U190 ( .A(n315), .Y(n233) );
  AND2X1_HVT U193 ( .A1(n249), .A2(n250), .Y(n236) );
  INVX0_HVT U196 ( .A(n598), .Y(n377) );
  MUX21X1_HVT U197 ( .A1(n236), .A2(n619), .S0(n324), .Y(n566) );
  AND2X1_HVT U199 ( .A1(n615), .A2(n414), .Y(n237) );
  MUX41X1_HVT U201 ( .A1(n436), .A3(n430), .A2(n445), .A4(n442), .S0(n335), 
        .S1(n238), .Y(out[7]) );
  MUX21X1_HVT U202 ( .A1(n596), .A2(n599), .S0(n325), .Y(n461) );
  MUX21X2_HVT U203 ( .A1(n516), .A2(n506), .S0(n239), .Y(out[3]) );
  IBUFFX16_HVT U204 ( .A(n307), .Y(n239) );
  NAND2X0_HVT U205 ( .A1(n396), .A2(n240), .Y(n241) );
  NAND2X0_HVT U206 ( .A1(n581), .A2(n326), .Y(n242) );
  NAND2X0_HVT U208 ( .A1(n241), .A2(n242), .Y(n438) );
  IBUFFX2_HVT U209 ( .A(n326), .Y(n240) );
  MUX21X1_HVT U210 ( .A1(n330), .A2(n409), .S0(n243), .Y(n427) );
  NAND2X0_HVT U211 ( .A1(n515), .A2(n244), .Y(n245) );
  NAND2X0_HVT U212 ( .A1(n514), .A2(n281), .Y(n246) );
  NAND2X0_HVT U213 ( .A1(n245), .A2(n246), .Y(n513) );
  INVX0_HVT U214 ( .A(n281), .Y(n244) );
  IBUFFX2_HVT U215 ( .A(n324), .Y(n281) );
  MUX21X2_HVT U216 ( .A1(n316), .A2(n412), .S0(n284), .Y(n598) );
  INVX0_HVT U217 ( .A(n292), .Y(n351) );
  MUX21X2_HVT U218 ( .A1(n532), .A2(n531), .S0(n247), .Y(n530) );
  IBUFFX16_HVT U219 ( .A(n323), .Y(n247) );
  MUX21X2_HVT U220 ( .A1(n480), .A2(n479), .S0(n323), .Y(n478) );
  MUX21X2_HVT U221 ( .A1(n407), .A2(n364), .S0(n325), .Y(n480) );
  NAND2X0_HVT U222 ( .A1(n218), .A2(n248), .Y(n249) );
  NAND2X0_HVT U223 ( .A1(n337), .A2(n263), .Y(n250) );
  NAND2X0_HVT U224 ( .A1(n249), .A2(n250), .Y(n597) );
  IBUFFX2_HVT U225 ( .A(n349), .Y(n263) );
  MUX21X1_HVT U226 ( .A1(n314), .A2(n597), .S0(n251), .Y(n475) );
  NBUFFX2_HVT U227 ( .A(n355), .Y(n327) );
  OA21X2_HVT U228 ( .A1(n361), .A2(n358), .A3(n368), .Y(n474) );
  MUX21X1_HVT U229 ( .A1(n338), .A2(n201), .S0(n285), .Y(n252) );
  IBUFFX16_HVT U230 ( .A(n252), .Y(n600) );
  INVX1_HVT U231 ( .A(n338), .Y(n414) );
  INVX1_HVT U232 ( .A(n427), .Y(n396) );
  NAND2X0_HVT U233 ( .A1(n444), .A2(n253), .Y(n254) );
  NAND2X0_HVT U234 ( .A1(n443), .A2(n289), .Y(n255) );
  NAND2X0_HVT U235 ( .A1(n254), .A2(n255), .Y(n442) );
  IBUFFX2_HVT U236 ( .A(n289), .Y(n253) );
  MUX21X1_HVT U237 ( .A1(n257), .A2(n316), .S0(n256), .Y(n429) );
  INVX0_HVT U238 ( .A(n333), .Y(n289) );
  INVX1_HVT U239 ( .A(n270), .Y(n258) );
  MUX21X2_HVT U240 ( .A1(n474), .A2(n475), .S0(n324), .Y(n473) );
  INVX1_HVT U241 ( .A(n426), .Y(n397) );
  MUX41X1_HVT U242 ( .A1(n398), .A3(n363), .A2(n620), .A4(n365), .S0(n261), 
        .S1(n358), .Y(n444) );
  IBUFFX16_HVT U243 ( .A(n319), .Y(n261) );
  INVX1_HVT U244 ( .A(n425), .Y(n398) );
  MUX21X2_HVT U245 ( .A1(n620), .A2(n252), .S0(n262), .Y(n559) );
  IBUFFX16_HVT U246 ( .A(n323), .Y(n262) );
  OR2X1_HVT U247 ( .A1(n328), .A2(n330), .Y(n621) );
  IBUFFX2_HVT U248 ( .A(n411), .Y(n308) );
  INVX1_HVT U249 ( .A(n429), .Y(n394) );
  IBUFFX2_HVT U250 ( .A(n614), .Y(n369) );
  MUX21X2_HVT U251 ( .A1(n553), .A2(n560), .S0(n307), .Y(out[0]) );
  INVX1_HVT U252 ( .A(in[3]), .Y(n411) );
  INVX0_HVT U253 ( .A(n331), .Y(n264) );
  MUX21X2_HVT U254 ( .A1(n471), .A2(n481), .S0(n307), .Y(out[5]) );
  MUX21X2_HVT U255 ( .A1(n548), .A2(n547), .S0(n266), .Y(n546) );
  IBUFFX16_HVT U256 ( .A(n267), .Y(n266) );
  INVX1_HVT U257 ( .A(n341), .Y(n413) );
  MUX21X1_HVT U258 ( .A1(n331), .A2(n414), .S0(n282), .Y(n586) );
  IBUFFX16_HVT U259 ( .A(n324), .Y(n267) );
  IBUFFX2_HVT U260 ( .A(n290), .Y(n275) );
  IBUFFX16_HVT U261 ( .A(n343), .Y(n269) );
  IBUFFX2_HVT U262 ( .A(in[4]), .Y(n358) );
  INVX1_HVT U263 ( .A(n349), .Y(n271) );
  IBUFFX2_HVT U264 ( .A(n355), .Y(n280) );
  NAND2X0_HVT U265 ( .A1(n450), .A2(n272), .Y(n273) );
  NAND2X0_HVT U266 ( .A1(n457), .A2(in[7]), .Y(n274) );
  NAND2X0_HVT U267 ( .A1(n273), .A2(n274), .Y(out[6]) );
  IBUFFX2_HVT U268 ( .A(in[7]), .Y(n272) );
  MUX41X1_HVT U269 ( .A1(n540), .A3(n544), .A2(n539), .A4(n543), .S0(n336), 
        .S1(n278), .Y(n538) );
  IBUFFX16_HVT U270 ( .A(n333), .Y(n278) );
  INVX1_HVT U271 ( .A(n593), .Y(n381) );
  MUX41X1_HVT U272 ( .A1(n464), .A3(n458), .A2(n466), .A4(n462), .S0(n335), 
        .S1(n288), .Y(n457) );
  MUX41X1_HVT U273 ( .A1(n237), .A3(n611), .A2(n412), .A4(n617), .S0(n279), 
        .S1(n280), .Y(n552) );
  IBUFFX16_HVT U274 ( .A(n320), .Y(n279) );
  INVX2_HVT U275 ( .A(n332), .Y(n334) );
  MUX21X2_HVT U276 ( .A1(n469), .A2(n470), .S0(n324), .Y(n466) );
  IBUFFX16_HVT U277 ( .A(n357), .Y(n354) );
  INVX1_HVT U278 ( .A(n350), .Y(n349) );
  INVX1_HVT U279 ( .A(n350), .Y(n290) );
  MUX41X1_HVT U280 ( .A1(n513), .A3(n510), .A2(n511), .A4(n507), .S0(n335), 
        .S1(n332), .Y(n506) );
  INVX2_HVT U281 ( .A(n335), .Y(n336) );
  INVX0_HVT U282 ( .A(n345), .Y(n412) );
  INVX1_HVT U283 ( .A(n346), .Y(n295) );
  NBUFFX2_HVT U284 ( .A(n349), .Y(n282) );
  NBUFFX2_HVT U285 ( .A(n349), .Y(n283) );
  NBUFFX2_HVT U286 ( .A(n291), .Y(n284) );
  AO21X1_HVT U287 ( .A1(n290), .A2(n409), .A3(n358), .Y(n433) );
  INVX1_HVT U288 ( .A(n286), .Y(n578) );
  NBUFFX2_HVT U289 ( .A(in[0]), .Y(n285) );
  INVX2_HVT U290 ( .A(n357), .Y(n355) );
  MUX21X1_HVT U291 ( .A1(n340), .A2(n345), .S0(n348), .Y(n286) );
  IBUFFX2_HVT U292 ( .A(n357), .Y(n301) );
  INVX0_HVT U293 ( .A(n325), .Y(n298) );
  MUX41X1_HVT U294 ( .A1(n412), .A3(n616), .A2(n575), .A4(n535), .S0(n320), 
        .S1(n301), .Y(n534) );
  INVX1_HVT U295 ( .A(n307), .Y(n299) );
  INVX1_HVT U296 ( .A(n357), .Y(n356) );
  NBUFFX2_HVT U297 ( .A(n355), .Y(n293) );
  INVX0_HVT U298 ( .A(n321), .Y(n305) );
  MUX41X1_HVT U299 ( .A1(n530), .A3(n534), .A2(n536), .A4(n537), .S0(n288), 
        .S1(in[5]), .Y(n529) );
  INVX1_HVT U300 ( .A(n289), .Y(n288) );
  MUX41X1_HVT U301 ( .A1(n517), .A3(n519), .A2(n518), .A4(n521), .S0(n336), 
        .S1(n288), .Y(n516) );
  OA21X1_HVT U302 ( .A1(n381), .A2(n358), .A3(n562), .Y(n437) );
  MUX41X1_HVT U303 ( .A1(n455), .A3(n452), .A2(n453), .A4(n451), .S0(n335), 
        .S1(n332), .Y(n450) );
  INVX1_HVT U304 ( .A(in[1]), .Y(n332) );
  NAND2X0_HVT U305 ( .A1(n448), .A2(n334), .Y(n296) );
  NAND2X0_HVT U306 ( .A1(n446), .A2(n289), .Y(n297) );
  NAND2X0_HVT U307 ( .A1(n297), .A2(n296), .Y(n445) );
  NBUFFX2_HVT U308 ( .A(n201), .Y(n344) );
  INVX0_HVT U309 ( .A(n542), .Y(n304) );
  INVX1_HVT U310 ( .A(n608), .Y(n303) );
  MUX41X1_HVT U311 ( .A1(n306), .A3(n304), .A2(n419), .A4(n303), .S0(n305), 
        .S1(n358), .Y(n302) );
  NAND2X0_HVT U312 ( .A1(n616), .A2(n339), .Y(n306) );
  INVX1_HVT U313 ( .A(in[0]), .Y(n350) );
  MUX41X1_HVT U314 ( .A1(n542), .A3(n398), .A2(n382), .A4(n541), .S0(n305), 
        .S1(n358), .Y(n540) );
  AO21X2_HVT U315 ( .A1(n350), .A2(n345), .A3(n358), .Y(n467) );
  NBUFFX2_HVT U316 ( .A(in[7]), .Y(n307) );
  INVX1_HVT U317 ( .A(n622), .Y(n409) );
  MUX21X2_HVT U318 ( .A1(n571), .A2(n570), .S0(n323), .Y(n569) );
  MUX21X2_HVT U319 ( .A1(n538), .A2(n545), .S0(n307), .Y(out[1]) );
  MUX21X2_HVT U320 ( .A1(n522), .A2(n529), .S0(n307), .Y(out[2]) );
  MUX21X2_HVT U321 ( .A1(n489), .A2(n490), .S0(n288), .Y(n488) );
  MUX21X2_HVT U322 ( .A1(n493), .A2(n494), .S0(n334), .Y(n492) );
  INVX0_HVT U323 ( .A(in[5]), .Y(n335) );
  NBUFFX2_HVT U324 ( .A(n618), .Y(n339) );
  AND2X1_HVT U325 ( .A1(n617), .A2(n201), .Y(n309) );
  NBUFFX2_HVT U326 ( .A(n618), .Y(n340) );
  AND2X1_HVT U327 ( .A1(n201), .A2(n200), .Y(n310) );
  MUX21X1_HVT U328 ( .A1(n330), .A2(n409), .S0(n349), .Y(n596) );
  MUX21X1_HVT U329 ( .A1(n295), .A2(n218), .S0(n347), .Y(n454) );
  MUX21X1_HVT U330 ( .A1(n295), .A2(n413), .S0(n348), .Y(n456) );
  MUX21X1_HVT U331 ( .A1(n409), .A2(n414), .S0(n347), .Y(n589) );
  MUX21X1_HVT U332 ( .A1(n339), .A2(n342), .S0(n290), .Y(n465) );
  MUX21X1_HVT U333 ( .A1(n218), .A2(n257), .S0(n285), .Y(n477) );
  MUX21X1_HVT U334 ( .A1(n328), .A2(n414), .S0(n282), .Y(n425) );
  MUX21X1_HVT U335 ( .A1(n295), .A2(n337), .S0(n348), .Y(n423) );
  MUX21X1_HVT U336 ( .A1(n329), .A2(n409), .S0(n291), .Y(n592) );
  MUX21X1_HVT U337 ( .A1(n329), .A2(n413), .S0(n348), .Y(n579) );
  MUX21X1_HVT U338 ( .A1(n337), .A2(n257), .S0(n283), .Y(n588) );
  MUX21X1_HVT U339 ( .A1(n414), .A2(n329), .S0(n347), .Y(n583) );
  MUX21X1_HVT U340 ( .A1(n337), .A2(n295), .S0(n283), .Y(n591) );
  MUX21X1_HVT U341 ( .A1(n366), .A2(n581), .S0(n327), .Y(n515) );
  MUX21X1_HVT U342 ( .A1(n409), .A2(n413), .S0(n292), .Y(n572) );
  MUX21X1_HVT U343 ( .A1(n258), .A2(n339), .S0(n348), .Y(n483) );
  MUX21X1_HVT U344 ( .A1(n414), .A2(n218), .S0(n283), .Y(n418) );
  MUX21X1_HVT U345 ( .A1(n340), .A2(n344), .S0(n283), .Y(n417) );
  MUX21X1_HVT U346 ( .A1(n218), .A2(n344), .S0(n285), .Y(n520) );
  XOR2X1_HVT U347 ( .A1(n341), .A2(n291), .Y(n575) );
  XNOR2X1_HVT U348 ( .A1(n344), .A2(n285), .Y(n311) );
  MUX21X1_HVT U349 ( .A1(n346), .A2(n344), .S0(n348), .Y(n608) );
  MUX21X1_HVT U350 ( .A1(n589), .A2(n310), .S0(n324), .Y(n498) );
  MUX21X1_HVT U351 ( .A1(n406), .A2(n311), .S0(n323), .Y(n501) );
  XOR2X1_HVT U352 ( .A1(n338), .A2(n290), .Y(n576) );
  XOR2X1_HVT U353 ( .A1(n346), .A2(n347), .Y(n585) );
  MUX21X1_HVT U354 ( .A1(n218), .A2(n337), .S0(n284), .Y(n582) );
  MUX21X1_HVT U355 ( .A1(n342), .A2(n329), .S0(n292), .Y(n603) );
  MUX21X1_HVT U356 ( .A1(n328), .A2(n342), .S0(n285), .Y(n420) );
  MUX21X1_HVT U357 ( .A1(n343), .A2(n330), .S0(n285), .Y(n504) );
  AND2X1_HVT U358 ( .A1(n284), .A2(n218), .Y(n312) );
  NBUFFX2_HVT U359 ( .A(n355), .Y(n325) );
  NBUFFX2_HVT U360 ( .A(n606), .Y(n337) );
  NBUFFX2_HVT U361 ( .A(n606), .Y(n338) );
  AND2X1_HVT U362 ( .A1(n413), .A2(n271), .Y(n313) );
  NBUFFX2_HVT U363 ( .A(n621), .Y(n341) );
  AND2X1_HVT U364 ( .A1(n343), .A2(n351), .Y(n314) );
  NBUFFX2_HVT U365 ( .A(n621), .Y(n343) );
  MUX21X1_HVT U366 ( .A1(n503), .A2(n505), .S0(n288), .Y(n502) );
  NBUFFX2_HVT U367 ( .A(n352), .Y(n322) );
  NBUFFX2_HVT U368 ( .A(n352), .Y(n324) );
  NBUFFX2_HVT U369 ( .A(n353), .Y(n323) );
  XNOR2X1_HVT U370 ( .A1(n357), .A2(n319), .Y(n315) );
  NBUFFX2_HVT U371 ( .A(n352), .Y(n318) );
  NBUFFX2_HVT U372 ( .A(n353), .Y(n319) );
  NBUFFX2_HVT U373 ( .A(n353), .Y(n320) );
  NBUFFX2_HVT U374 ( .A(n353), .Y(n321) );
  NBUFFX2_HVT U375 ( .A(n352), .Y(n317) );
  INVX1_HVT U376 ( .A(n332), .Y(n333) );
  MUX21X1_HVT U377 ( .A1(n295), .A2(n308), .S0(n290), .Y(n416) );
  MUX21X1_HVT U378 ( .A1(n339), .A2(n308), .S0(n347), .Y(n527) );
  MUX21X1_HVT U379 ( .A1(n413), .A2(n257), .S0(n347), .Y(n509) );
  MUX21X1_HVT U380 ( .A1(n345), .A2(n308), .S0(n292), .Y(n468) );
  MUX21X1_HVT U381 ( .A1(n308), .A2(n340), .S0(n290), .Y(n421) );
  MUX21X1_HVT U382 ( .A1(n308), .A2(n345), .S0(n283), .Y(n422) );
  NBUFFX2_HVT U383 ( .A(in[2]), .Y(n353) );
  NBUFFX2_HVT U384 ( .A(in[2]), .Y(n352) );
  INVX1_HVT U385 ( .A(in[6]), .Y(n415) );
  MUX21X1_HVT U386 ( .A1(n409), .A2(n316), .S0(n347), .Y(n491) );
  XOR2X1_HVT U387 ( .A1(n285), .A2(n316), .Y(n573) );
  MUX21X1_HVT U388 ( .A1(n316), .A2(n343), .S0(n282), .Y(n428) );
  MUX21X1_HVT U389 ( .A1(n342), .A2(n316), .S0(n291), .Y(n424) );
  MUX21X1_HVT U390 ( .A1(n328), .A2(n316), .S0(n292), .Y(n419) );
  NBUFFX2_HVT U391 ( .A(n623), .Y(n345) );
  NBUFFX2_HVT U392 ( .A(n623), .Y(n346) );
  INVX0_HVT U393 ( .A(n584), .Y(n360) );
  INVX0_HVT U394 ( .A(n524), .Y(n361) );
  INVX0_HVT U395 ( .A(n486), .Y(n362) );
  INVX0_HVT U396 ( .A(n620), .Y(n363) );
  INVX0_HVT U397 ( .A(n619), .Y(n364) );
  INVX0_HVT U398 ( .A(n616), .Y(n366) );
  INVX0_HVT U399 ( .A(n609), .Y(n368) );
  INVX0_HVT U400 ( .A(n610), .Y(n370) );
  INVX0_HVT U401 ( .A(n603), .Y(n373) );
  INVX0_HVT U402 ( .A(n602), .Y(n374) );
  INVX0_HVT U403 ( .A(n596), .Y(n378) );
  INVX0_HVT U404 ( .A(n592), .Y(n382) );
  INVX0_HVT U405 ( .A(n591), .Y(n383) );
  INVX0_HVT U406 ( .A(n589), .Y(n384) );
  INVX0_HVT U407 ( .A(n588), .Y(n385) );
  INVX0_HVT U408 ( .A(n586), .Y(n386) );
  INVX0_HVT U409 ( .A(n585), .Y(n387) );
  INVX0_HVT U410 ( .A(n583), .Y(n388) );
  INVX0_HVT U411 ( .A(n582), .Y(n389) );
  INVX0_HVT U412 ( .A(n576), .Y(n392) );
  INVX0_HVT U413 ( .A(n613), .Y(n393) );
  INVX0_HVT U414 ( .A(n428), .Y(n395) );
  INVX0_HVT U415 ( .A(n424), .Y(n399) );
  INVX0_HVT U416 ( .A(n423), .Y(n400) );
  INVX0_HVT U417 ( .A(n422), .Y(n401) );
  INVX0_HVT U418 ( .A(n421), .Y(n402) );
  INVX0_HVT U419 ( .A(n420), .Y(n403) );
  INVX0_HVT U420 ( .A(n419), .Y(n404) );
  INVX0_HVT U421 ( .A(n468), .Y(n405) );
  INVX0_HVT U422 ( .A(n418), .Y(n406) );
  INVX0_HVT U423 ( .A(n416), .Y(n408) );
endmodule

