
module inv_sbox_3 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n5, n196, n197, n198, n199, n200, n201, n202, n208, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597;

  NAND2X0_HVT U1 ( .A1(n265), .A2(n303), .Y(n597) );
  NAND2X0_HVT U4 ( .A1(n252), .A2(n200), .Y(n594) );
  NAND2X0_HVT U8 ( .A1(n247), .A2(n311), .Y(n590) );
  NAND2X0_HVT U9 ( .A1(n288), .A2(n254), .Y(n589) );
  NAND2X0_HVT U10 ( .A1(n287), .A2(n587), .Y(n588) );
  NAND2X0_HVT U11 ( .A1(n322), .A2(n201), .Y(n586) );
  NAND2X0_HVT U12 ( .A1(n252), .A2(n301), .Y(n585) );
  NAND2X0_HVT U13 ( .A1(n590), .A2(n314), .Y(n584) );
  NAND2X0_HVT U15 ( .A1(n309), .A2(n320), .Y(n582) );
  NAND2X0_HVT U19 ( .A1(n319), .A2(n387), .Y(n577) );
  NAND2X0_HVT U25 ( .A1(in[6]), .A2(n264), .Y(n593) );
  NAND2X0_HVT U32 ( .A1(n238), .A2(n322), .Y(n565) );
  NAND2X0_HVT U35 ( .A1(n590), .A2(n388), .Y(n562) );
  NAND2X0_HVT U38 ( .A1(n301), .A2(n322), .Y(n559) );
  NAND2X0_HVT U42 ( .A1(n592), .A2(n388), .Y(n555) );
  OA21X1_HVT U53 ( .A1(n328), .A2(n547), .A3(n356), .Y(n545) );
  NAND2X0_HVT U55 ( .A1(n314), .A2(n594), .Y(n543) );
  AO21X1_HVT U60 ( .A1(n537), .A2(n298), .A3(n576), .Y(n538) );
  MUX41X1_HVT U62 ( .A1(n536), .A3(n542), .A2(n540), .A4(n544), .S0(in[5]), 
        .S1(n305), .Y(n535) );
  MUX41X1_HVT U65 ( .A1(n346), .A3(n348), .A2(n347), .A4(n559), .S0(n294), 
        .S1(n249), .Y(n532) );
  NAND2X0_HVT U66 ( .A1(n316), .A2(n263), .Y(n531) );
  MUX41X1_HVT U67 ( .A1(n343), .A3(n371), .A2(n345), .A4(n531), .S0(n300), 
        .S1(n291), .Y(n530) );
  MUX41X1_HVT U71 ( .A1(n592), .A3(n284), .A2(n586), .A4(n339), .S0(n293), 
        .S1(n324), .Y(n527) );
  NAND2X0_HVT U72 ( .A1(n310), .A2(n591), .Y(n526) );
  MUX41X1_HVT U73 ( .A1(n570), .A3(n526), .A2(n372), .A4(n301), .S0(n299), 
        .S1(n290), .Y(n525) );
  MUX41X1_HVT U74 ( .A1(n588), .A3(n361), .A2(n360), .A4(n349), .S0(n294), 
        .S1(n249), .Y(n524) );
  NAND2X0_HVT U81 ( .A1(n201), .A2(n591), .Y(n517) );
  AND2X1_HVT U82 ( .A1(n592), .A2(n240), .Y(n516) );
  MUX41X1_HVT U84 ( .A1(n279), .A3(n357), .A2(n375), .A4(n572), .S0(n294), 
        .S1(n250), .Y(n514) );
  MUX41X1_HVT U87 ( .A1(n334), .A3(n279), .A2(n376), .A4(n354), .S0(n292), 
        .S1(n250), .Y(n512) );
  MUX41X1_HVT U88 ( .A1(n345), .A3(n331), .A2(n567), .A4(n551), .S0(n293), 
        .S1(n324), .Y(n511) );
  NAND2X0_HVT U89 ( .A1(n322), .A2(n386), .Y(n510) );
  MUX41X1_HVT U90 ( .A1(n282), .A3(n591), .A2(n550), .A4(n510), .S0(n293), 
        .S1(n326), .Y(n509) );
  MUX41X1_HVT U96 ( .A1(n371), .A3(n584), .A2(n355), .A4(n377), .S0(n294), 
        .S1(n324), .Y(n503) );
  MUX41X1_HVT U98 ( .A1(n502), .A3(n378), .A2(n362), .A4(n569), .S0(n294), 
        .S1(n250), .Y(n501) );
  MUX41X1_HVT U99 ( .A1(n565), .A3(n347), .A2(n549), .A4(n202), .S0(n249), 
        .S1(n291), .Y(n500) );
  MUX41X1_HVT U101 ( .A1(n379), .A3(n585), .A2(n272), .A4(n499), .S0(n324), 
        .S1(n289), .Y(n498) );
  AND2X1_HVT U104 ( .A1(n591), .A2(n593), .Y(n496) );
  MUX41X1_HVT U105 ( .A1(n583), .A3(n380), .A2(n517), .A4(n496), .S0(n294), 
        .S1(n249), .Y(n495) );
  MUX41X1_HVT U107 ( .A1(n379), .A3(n240), .A2(n494), .A4(n336), .S0(n293), 
        .S1(n326), .Y(n493) );
  MUX41X1_HVT U108 ( .A1(n349), .A3(n202), .A2(n354), .A4(n201), .S0(n294), 
        .S1(n324), .Y(n492) );
  MUX41X1_HVT U109 ( .A1(n378), .A3(n331), .A2(n375), .A4(n368), .S0(n293), 
        .S1(n250), .Y(n491) );
  MUX41X1_HVT U110 ( .A1(n491), .A3(n493), .A2(n492), .A4(n495), .S0(n308), 
        .S1(n305), .Y(n490) );
  NAND2X0_HVT U114 ( .A1(n288), .A2(n591), .Y(n486) );
  MUX41X1_HVT U115 ( .A1(n486), .A3(n586), .A2(n364), .A4(n240), .S0(n324), 
        .S1(n291), .Y(n485) );
  MUX41X1_HVT U116 ( .A1(n363), .A3(n357), .A2(n331), .A4(n582), .S0(n292), 
        .S1(n250), .Y(n484) );
  NAND2X0_HVT U118 ( .A1(n322), .A2(n265), .Y(n482) );
  MUX41X1_HVT U119 ( .A1(n381), .A3(n483), .A2(n560), .A4(n482), .S0(n292), 
        .S1(n249), .Y(n481) );
  MUX41X1_HVT U120 ( .A1(n481), .A3(n485), .A2(n484), .A4(n487), .S0(n308), 
        .S1(n306), .Y(n480) );
  MUX41X1_HVT U122 ( .A1(n369), .A3(n276), .A2(n551), .A4(n373), .S0(n292), 
        .S1(n326), .Y(n479) );
  MUX41X1_HVT U124 ( .A1(n278), .A3(n478), .A2(n574), .A4(n351), .S0(n298), 
        .S1(n292), .Y(n477) );
  AOI21X1_HVT U127 ( .A1(n297), .A2(n473), .A3(n337), .Y(n474) );
  NAND2X0_HVT U129 ( .A1(n296), .A2(n286), .Y(n471) );
  MUX41X1_HVT U130 ( .A1(n471), .A3(n472), .A2(n475), .A4(n474), .S0(n300), 
        .S1(n305), .Y(n470) );
  AND2X1_HVT U131 ( .A1(n263), .A2(n241), .Y(n469) );
  MUX41X1_HVT U132 ( .A1(n245), .A3(n469), .A2(n383), .A4(n343), .S0(n299), 
        .S1(n290), .Y(n468) );
  MUX41X1_HVT U133 ( .A1(n384), .A3(n336), .A2(n543), .A4(n335), .S0(n298), 
        .S1(n289), .Y(n467) );
  MUX41X1_HVT U136 ( .A1(n548), .A3(n499), .A2(n465), .A4(n341), .S0(n296), 
        .S1(n326), .Y(n464) );
  MUX41X1_HVT U137 ( .A1(n254), .A3(n568), .A2(n572), .A4(n377), .S0(n300), 
        .S1(n289), .Y(n463) );
  MUX41X1_HVT U139 ( .A1(n462), .A3(n466), .A2(n470), .A4(n476), .S0(n308), 
        .S1(n260), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n360), .A3(n277), .A2(n353), .A4(n586), .S0(n299), 
        .S1(n291), .Y(n461) );
  NAND2X0_HVT U141 ( .A1(n309), .A2(n322), .Y(n460) );
  MUX41X1_HVT U143 ( .A1(n386), .A3(n365), .A2(n577), .A4(n574), .S0(n295), 
        .S1(n326), .Y(n458) );
  MUX41X1_HVT U145 ( .A1(n566), .A3(n380), .A2(n457), .A4(n517), .S0(n297), 
        .S1(n325), .Y(n456) );
  AO21X1_HVT U148 ( .A1(n300), .A2(n338), .A3(n197), .Y(n453) );
  NAND2X0_HVT U159 ( .A1(n442), .A2(n441), .Y(n443) );
  MUX41X1_HVT U162 ( .A1(n366), .A3(n348), .A2(n562), .A4(n439), .S0(n295), 
        .S1(n325), .Y(n438) );
  NAND2X0_HVT U163 ( .A1(n320), .A2(n386), .Y(n437) );
  MUX41X1_HVT U164 ( .A1(n589), .A3(n437), .A2(n560), .A4(n349), .S0(n292), 
        .S1(n325), .Y(n436) );
  MUX41X1_HVT U170 ( .A1(n280), .A3(n275), .A2(n278), .A4(n430), .S0(n295), 
        .S1(n325), .Y(n429) );
  MUX41X1_HVT U173 ( .A1(n287), .A3(n284), .A2(n200), .A4(n561), .S0(n295), 
        .S1(n325), .Y(n426) );
  MUX41X1_HVT U174 ( .A1(n376), .A3(n543), .A2(n384), .A4(n388), .S0(n295), 
        .S1(n249), .Y(n425) );
  MUX41X1_HVT U175 ( .A1(n425), .A3(n426), .A2(n427), .A4(n429), .S0(n306), 
        .S1(n308), .Y(n424) );
  NAND2X0_HVT U177 ( .A1(n319), .A2(n265), .Y(n423) );
  MUX41X1_HVT U178 ( .A1(n280), .A3(n423), .A2(n282), .A4(n553), .S0(n295), 
        .S1(n325), .Y(n422) );
  AND2X1_HVT U179 ( .A1(n592), .A2(n593), .Y(n421) );
  MUX41X1_HVT U182 ( .A1(n336), .A3(n594), .A2(n334), .A4(n239), .S0(n292), 
        .S1(n326), .Y(n418) );
  MUX41X1_HVT U183 ( .A1(n365), .A3(n370), .A2(n349), .A4(n555), .S0(n298), 
        .S1(n290), .Y(n417) );
  AND2X1_HVT U185 ( .A1(n388), .A2(n241), .Y(n415) );
  MUX41X1_HVT U190 ( .A1(n412), .A3(n413), .A2(n411), .A4(n414), .S0(n306), 
        .S1(n290), .Y(n410) );
  NAND2X0_HVT U191 ( .A1(n328), .A2(n342), .Y(n409) );
  AND2X1_HVT U192 ( .A1(n361), .A2(n407), .Y(n408) );
  NAND2X0_HVT U194 ( .A1(n555), .A2(n407), .Y(n405) );
  NAND2X0_HVT U198 ( .A1(n316), .A2(n388), .Y(n587) );
  NAND2X0_HVT U200 ( .A1(n311), .A2(n322), .Y(n473) );
  NAND2X0_HVT U207 ( .A1(n322), .A2(n283), .Y(n537) );
  MUX21X2_HVT U2 ( .A1(n358), .A2(n516), .S0(n242), .Y(n258) );
  INVX2_HVT U3 ( .A(n327), .Y(n250) );
  INVX1_HVT U5 ( .A(n321), .Y(n248) );
  MUX21X2_HVT U6 ( .A1(n386), .A2(n282), .S0(n320), .Y(n553) );
  IBUFFX2_HVT U7 ( .A(n321), .Y(n320) );
  MUX21X2_HVT U14 ( .A1(n594), .A2(n350), .S0(n242), .Y(n534) );
  IBUFFX2_HVT U16 ( .A(n327), .Y(n249) );
  IBUFFX2_HVT U17 ( .A(n327), .Y(n325) );
  INVX1_HVT U18 ( .A(n385), .Y(n5) );
  INVX1_HVT U20 ( .A(n385), .Y(n196) );
  INVX1_HVT U21 ( .A(n5), .Y(n197) );
  INVX1_HVT U22 ( .A(n196), .Y(n198) );
  IBUFFX2_HVT U23 ( .A(n596), .Y(n199) );
  INVX1_HVT U24 ( .A(n199), .Y(n200) );
  INVX1_HVT U26 ( .A(n199), .Y(n201) );
  IBUFFX2_HVT U27 ( .A(n596), .Y(n385) );
  IBUFFX2_HVT U28 ( .A(n274), .Y(n236) );
  MUX21X1_HVT U29 ( .A1(n255), .A2(n256), .S0(n324), .Y(n420) );
  IBUFFX16_HVT U30 ( .A(n327), .Y(n324) );
  IBUFFX2_HVT U31 ( .A(n388), .Y(n202) );
  MUX21X2_HVT U33 ( .A1(n449), .A2(n448), .S0(n208), .Y(n447) );
  IBUFFX16_HVT U34 ( .A(n297), .Y(n208) );
  NAND2X0_HVT U36 ( .A1(n445), .A2(n218), .Y(n219) );
  NAND2X0_HVT U37 ( .A1(n455), .A2(n260), .Y(n220) );
  NAND2X0_HVT U39 ( .A1(n219), .A2(n220), .Y(out[5]) );
  IBUFFX2_HVT U40 ( .A(n260), .Y(n218) );
  MUX21X1_HVT U41 ( .A1(n310), .A2(n303), .S0(n317), .Y(n572) );
  INVX2_HVT U43 ( .A(n581), .Y(n388) );
  INVX1_HVT U44 ( .A(n317), .Y(n241) );
  MUX21X2_HVT U45 ( .A1(n517), .A2(n239), .S0(n242), .Y(n259) );
  NAND2X0_HVT U46 ( .A1(n552), .A2(n221), .Y(n222) );
  NAND2X0_HVT U47 ( .A1(n421), .A2(n225), .Y(n223) );
  NAND2X0_HVT U48 ( .A1(n222), .A2(n223), .Y(n256) );
  INVX0_HVT U49 ( .A(n225), .Y(n221) );
  IBUFFX2_HVT U50 ( .A(n294), .Y(n225) );
  OA21X1_HVT U51 ( .A1(n333), .A2(n328), .A3(n576), .Y(n522) );
  INVX1_HVT U52 ( .A(n576), .Y(n349) );
  INVX2_HVT U54 ( .A(in[3]), .Y(n264) );
  MUX21X2_HVT U56 ( .A1(n279), .A2(n572), .S0(n224), .Y(n449) );
  IBUFFX16_HVT U57 ( .A(n299), .Y(n224) );
  INVX1_HVT U58 ( .A(in[4]), .Y(n327) );
  INVX0_HVT U59 ( .A(n552), .Y(n367) );
  MUX41X1_HVT U61 ( .A1(n406), .A3(n405), .A2(n408), .A4(n409), .S0(n293), 
        .S1(n306), .Y(n404) );
  MUX21X1_HVT U63 ( .A1(n367), .A2(n278), .S0(n298), .Y(n406) );
  OA21X1_HVT U64 ( .A1(n332), .A2(n328), .A3(n340), .Y(n448) );
  MUX41X1_HVT U68 ( .A1(n362), .A3(n239), .A2(n451), .A4(n350), .S0(n226), 
        .S1(n289), .Y(n450) );
  IBUFFX16_HVT U69 ( .A(n298), .Y(n226) );
  MUX41X1_HVT U70 ( .A1(n519), .A3(n518), .A2(n515), .A4(n514), .S0(n227), 
        .S1(n228), .Y(n513) );
  IBUFFX16_HVT U75 ( .A(n305), .Y(n227) );
  IBUFFX16_HVT U76 ( .A(in[5]), .Y(n228) );
  NAND2X1_HVT U77 ( .A1(n248), .A2(n313), .Y(n591) );
  MUX41X1_HVT U78 ( .A1(n428), .A3(n510), .A2(n575), .A4(n275), .S0(n229), 
        .S1(n250), .Y(n427) );
  IBUFFX16_HVT U79 ( .A(n295), .Y(n229) );
  NAND2X2_HVT U80 ( .A1(n316), .A2(n315), .Y(n592) );
  MUX21X2_HVT U83 ( .A1(n372), .A2(n556), .S0(n299), .Y(n412) );
  MUX21X1_HVT U85 ( .A1(n263), .A2(n387), .S0(n318), .Y(n556) );
  NAND2X0_HVT U86 ( .A1(n313), .A2(n230), .Y(n231) );
  NAND2X0_HVT U91 ( .A1(n508), .A2(n237), .Y(n232) );
  NAND2X0_HVT U92 ( .A1(n231), .A2(n232), .Y(n507) );
  INVX0_HVT U93 ( .A(n237), .Y(n230) );
  NAND2X0_HVT U94 ( .A1(n497), .A2(n233), .Y(n234) );
  NAND2X0_HVT U95 ( .A1(n504), .A2(n260), .Y(n235) );
  NAND2X0_HVT U97 ( .A1(n234), .A2(n235), .Y(out[2]) );
  IBUFFX2_HVT U100 ( .A(n260), .Y(n233) );
  NBUFFX4_HVT U102 ( .A(n595), .Y(n313) );
  MUX21X1_HVT U103 ( .A1(n309), .A2(n303), .S0(n299), .Y(n508) );
  IBUFFX2_HVT U106 ( .A(n248), .Y(n237) );
  MUX21X2_HVT U111 ( .A1(n258), .A2(n259), .S0(n324), .Y(n515) );
  IBUFFX2_HVT U112 ( .A(n321), .Y(n247) );
  MUX41X1_HVT U113 ( .A1(n432), .A3(n438), .A2(n436), .A4(n440), .S0(n308), 
        .S1(n236), .Y(n431) );
  AO21X2_HVT U117 ( .A1(n364), .A2(n299), .A3(n573), .Y(n488) );
  MUX41X1_HVT U121 ( .A1(n419), .A3(n416), .A2(n410), .A4(n404), .S0(n307), 
        .S1(n266), .Y(out[7]) );
  INVX0_HVT U123 ( .A(in[7]), .Y(n266) );
  INVX1_HVT U125 ( .A(n321), .Y(n252) );
  NBUFFX4_HVT U126 ( .A(n389), .Y(n302) );
  MUX21X2_HVT U128 ( .A1(n571), .A2(n574), .S0(n298), .Y(n435) );
  INVX0_HVT U134 ( .A(n574), .Y(n351) );
  MUX21X2_HVT U135 ( .A1(n198), .A2(n265), .S0(n318), .Y(n574) );
  INVX1_HVT U138 ( .A(n264), .Y(n265) );
  INVX2_HVT U142 ( .A(n241), .Y(n318) );
  MUX21X2_HVT U144 ( .A1(n422), .A2(n420), .S0(n304), .Y(n419) );
  MUX21X1_HVT U146 ( .A1(n383), .A2(n245), .S0(n298), .Y(n454) );
  MUX21X1_HVT U147 ( .A1(n454), .A2(n453), .S0(n296), .Y(n452) );
  INVX0_HVT U149 ( .A(n321), .Y(n316) );
  INVX1_HVT U150 ( .A(n317), .Y(n322) );
  AO21X1_HVT U151 ( .A1(n241), .A2(n288), .A3(n328), .Y(n441) );
  INVX0_HVT U152 ( .A(n285), .Y(n286) );
  INVX1_HVT U153 ( .A(n241), .Y(n319) );
  INVX1_HVT U154 ( .A(n273), .Y(n238) );
  INVX0_HVT U155 ( .A(n302), .Y(n273) );
  OR2X1_HVT U156 ( .A1(n264), .A2(n389), .Y(n595) );
  IBUFFX2_HVT U157 ( .A(n389), .Y(n263) );
  MUX21X2_HVT U158 ( .A1(n373), .A2(n330), .S0(n300), .Y(n523) );
  OA21X1_HVT U160 ( .A1(n357), .A2(n328), .A3(n537), .Y(n411) );
  MUX21X1_HVT U161 ( .A1(n279), .A2(n549), .S0(n300), .Y(n413) );
  INVX1_HVT U165 ( .A(in[0]), .Y(n321) );
  NBUFFX2_HVT U166 ( .A(n246), .Y(n299) );
  AO21X1_HVT U167 ( .A1(n316), .A2(n198), .A3(n328), .Y(n407) );
  NAND2X0_HVT U168 ( .A1(n587), .A2(n433), .Y(n434) );
  AND2X1_HVT U169 ( .A1(n559), .A2(n271), .Y(n239) );
  INVX1_HVT U171 ( .A(n266), .Y(n260) );
  INVX1_HVT U172 ( .A(n297), .Y(n242) );
  NBUFFX2_HVT U176 ( .A(n323), .Y(n293) );
  INVX0_HVT U180 ( .A(n295), .Y(n257) );
  INVX1_HVT U181 ( .A(in[5]), .Y(n307) );
  INVX1_HVT U184 ( .A(n307), .Y(n308) );
  MUX21X2_HVT U186 ( .A1(n523), .A2(n522), .S0(n297), .Y(n521) );
  MUX21X2_HVT U187 ( .A1(n337), .A2(n556), .S0(n300), .Y(n489) );
  INVX1_HVT U188 ( .A(n400), .Y(n373) );
  MUX21X2_HVT U189 ( .A1(n488), .A2(n489), .S0(n297), .Y(n487) );
  INVX2_HVT U193 ( .A(n312), .Y(n387) );
  NBUFFX2_HVT U195 ( .A(n312), .Y(n240) );
  INVX1_HVT U196 ( .A(n321), .Y(n317) );
  NAND2X0_HVT U197 ( .A1(n443), .A2(n242), .Y(n243) );
  NAND2X0_HVT U199 ( .A1(n444), .A2(n297), .Y(n244) );
  NAND2X0_HVT U201 ( .A1(n243), .A2(n244), .Y(n440) );
  MUX21X1_HVT U202 ( .A1(n373), .A2(n554), .S0(n251), .Y(n444) );
  AND2X1_HVT U203 ( .A1(n594), .A2(n311), .Y(n245) );
  AO21X1_HVT U204 ( .A1(n310), .A2(n594), .A3(n328), .Y(n433) );
  INVX0_HVT U205 ( .A(n586), .Y(n329) );
  MUX21X2_HVT U206 ( .A1(n329), .A2(n565), .S0(n257), .Y(n255) );
  NBUFFX2_HVT U208 ( .A(in[4]), .Y(n246) );
  INVX1_HVT U209 ( .A(in[4]), .Y(n328) );
  MUX21X1_HVT U210 ( .A1(n352), .A2(n541), .S0(n281), .Y(n540) );
  IBUFFX2_HVT U211 ( .A(n299), .Y(n251) );
  XNOR2X2_HVT U212 ( .A1(n302), .A2(n264), .Y(n581) );
  MUX21X1_HVT U213 ( .A1(n351), .A2(n543), .S0(n299), .Y(n539) );
  MUX21X1_HVT U214 ( .A1(n339), .A2(n309), .S0(n300), .Y(n506) );
  MUX21X2_HVT U215 ( .A1(n539), .A2(n538), .S0(n296), .Y(n536) );
  MUX21X2_HVT U216 ( .A1(n480), .A2(n490), .S0(n260), .Y(out[3]) );
  MUX21X1_HVT U217 ( .A1(n415), .A2(n374), .S0(n298), .Y(n414) );
  IBUFFX2_HVT U218 ( .A(n594), .Y(n334) );
  INVX0_HVT U219 ( .A(n245), .Y(n253) );
  INVX0_HVT U220 ( .A(n338), .Y(n254) );
  MUX21X2_HVT U221 ( .A1(n506), .A2(n507), .S0(n296), .Y(n505) );
  MUX41X1_HVT U222 ( .A1(n543), .A3(n354), .A2(n202), .A4(n370), .S0(n242), 
        .S1(n327), .Y(n542) );
  IBUFFX2_HVT U223 ( .A(n327), .Y(n326) );
  INVX0_HVT U224 ( .A(n272), .Y(n561) );
  INVX0_HVT U225 ( .A(n572), .Y(n353) );
  MUX41X1_HVT U226 ( .A1(n580), .A3(n359), .A2(n579), .A4(n357), .S0(n257), 
        .S1(n328), .Y(n519) );
  INVX1_HVT U227 ( .A(n305), .Y(n274) );
  INVX1_HVT U228 ( .A(n304), .Y(n306) );
  MUX41X1_HVT U229 ( .A1(n353), .A3(n382), .A2(n558), .A4(n460), .S0(n242), 
        .S1(n327), .Y(n459) );
  MUX41X1_HVT U230 ( .A1(n461), .A3(n459), .A2(n458), .A4(n456), .S0(n274), 
        .S1(n307), .Y(n455) );
  IBUFFX2_HVT U231 ( .A(n554), .Y(n365) );
  MUX41X1_HVT U232 ( .A1(n501), .A3(n498), .A2(n503), .A4(n500), .S0(n307), 
        .S1(n305), .Y(n497) );
  MUX41X1_HVT U233 ( .A1(n512), .A3(n509), .A2(n511), .A4(n505), .S0(n307), 
        .S1(n274), .Y(n504) );
  MUX21X2_HVT U234 ( .A1(n513), .A2(n520), .S0(in[7]), .Y(out[1]) );
  MUX21X2_HVT U235 ( .A1(n477), .A2(n479), .S0(n306), .Y(n476) );
  MUX41X1_HVT U236 ( .A1(n374), .A3(n589), .A2(n370), .A4(n253), .S0(n249), 
        .S1(n293), .Y(n518) );
  INVX1_HVT U237 ( .A(n304), .Y(n305) );
  INVX1_HVT U238 ( .A(n403), .Y(n370) );
  MUX41X1_HVT U239 ( .A1(n527), .A3(n524), .A2(n525), .A4(n521), .S0(n307), 
        .S1(n304), .Y(n520) );
  MUX41X1_HVT U240 ( .A1(n343), .A3(n344), .A2(n265), .A4(n286), .S0(n250), 
        .S1(n293), .Y(n529) );
  NAND2X0_HVT U241 ( .A1(n535), .A2(n260), .Y(n261) );
  NAND2X0_HVT U242 ( .A1(n528), .A2(n266), .Y(n262) );
  NAND2X0_HVT U243 ( .A1(n261), .A2(n262), .Y(out[0]) );
  MUX41X1_HVT U244 ( .A1(n355), .A3(n578), .A2(n586), .A4(n353), .S0(n242), 
        .S1(n328), .Y(n446) );
  MUX21X1_HVT U245 ( .A1(n546), .A2(n545), .S0(n296), .Y(n544) );
  NAND2X0_HVT U246 ( .A1(n424), .A2(n266), .Y(n267) );
  INVX1_HVT U247 ( .A(in[6]), .Y(n389) );
  NBUFFX2_HVT U248 ( .A(n389), .Y(n303) );
  MUX21X1_HVT U249 ( .A1(n467), .A2(n468), .S0(n306), .Y(n466) );
  MUX21X1_HVT U250 ( .A1(n463), .A2(n464), .S0(n306), .Y(n462) );
  MUX21X1_HVT U251 ( .A1(n284), .A2(n238), .S0(n316), .Y(n428) );
  INVX1_HVT U252 ( .A(n401), .Y(n372) );
  NAND2X0_HVT U253 ( .A1(n431), .A2(in[7]), .Y(n268) );
  NAND2X0_HVT U254 ( .A1(n267), .A2(n268), .Y(out[6]) );
  MUX41X1_HVT U255 ( .A1(n533), .A3(n530), .A2(n532), .A4(n529), .S0(n307), 
        .S1(n274), .Y(n528) );
  MUX21X2_HVT U256 ( .A1(n349), .A2(n534), .S0(n281), .Y(n533) );
  NAND2X0_HVT U257 ( .A1(n417), .A2(n304), .Y(n269) );
  NAND2X0_HVT U258 ( .A1(n418), .A2(n306), .Y(n270) );
  NAND2X0_HVT U259 ( .A1(n269), .A2(n270), .Y(n416) );
  NAND2X0_HVT U260 ( .A1(n388), .A2(n318), .Y(n271) );
  MUX21X2_HVT U261 ( .A1(n434), .A2(n435), .S0(n296), .Y(n432) );
  MUX21X1_HVT U262 ( .A1(n309), .A2(n273), .S0(n322), .Y(n272) );
  MUX41X1_HVT U263 ( .A1(n452), .A3(n447), .A2(n450), .A4(n446), .S0(n307), 
        .S1(n274), .Y(n445) );
  MUX21X2_HVT U264 ( .A1(n355), .A2(n344), .S0(n300), .Y(n546) );
  INVX0_HVT U265 ( .A(n597), .Y(n285) );
  AND2X1_HVT U266 ( .A1(n592), .A2(n200), .Y(n275) );
  AND2X1_HVT U267 ( .A1(n201), .A2(n582), .Y(n276) );
  MUX21X1_HVT U268 ( .A1(n302), .A2(n386), .S0(n318), .Y(n451) );
  MUX21X1_HVT U269 ( .A1(n388), .A2(n301), .S0(n318), .Y(n558) );
  MUX21X1_HVT U270 ( .A1(n197), .A2(n238), .S0(n319), .Y(n401) );
  MUX21X1_HVT U271 ( .A1(n593), .A2(n313), .S0(n318), .Y(n439) );
  NAND2X0_HVT U272 ( .A1(n264), .A2(n302), .Y(n596) );
  MUX21X1_HVT U273 ( .A1(n388), .A2(n238), .S0(n320), .Y(n392) );
  MUX21X1_HVT U274 ( .A1(n303), .A2(n197), .S0(n252), .Y(n571) );
  MUX21X1_HVT U275 ( .A1(n309), .A2(n301), .S0(n252), .Y(n576) );
  MUX21X1_HVT U276 ( .A1(n309), .A2(n284), .S0(n248), .Y(n566) );
  MUX21X1_HVT U277 ( .A1(n301), .A2(n197), .S0(n318), .Y(n567) );
  MUX21X1_HVT U278 ( .A1(n382), .A2(n277), .S0(n296), .Y(n475) );
  MUX21X1_HVT U279 ( .A1(n282), .A2(n310), .S0(n247), .Y(n397) );
  MUX21X1_HVT U280 ( .A1(n198), .A2(n387), .S0(n252), .Y(n547) );
  XOR2X1_HVT U281 ( .A1(n287), .A2(n248), .Y(n560) );
  XNOR2X1_HVT U282 ( .A1(n201), .A2(n247), .Y(n277) );
  MUX21X1_HVT U283 ( .A1(n283), .A2(n387), .S0(n318), .Y(n430) );
  MUX21X1_HVT U284 ( .A1(n302), .A2(n200), .S0(n319), .Y(n494) );
  XOR2X1_HVT U285 ( .A1(n309), .A2(n252), .Y(n551) );
  MUX21X1_HVT U286 ( .A1(n310), .A2(n386), .S0(n319), .Y(n563) );
  MUX21X1_HVT U287 ( .A1(n593), .A2(n201), .S0(n248), .Y(n391) );
  MUX21X1_HVT U288 ( .A1(n301), .A2(n200), .S0(n319), .Y(n399) );
  INVX1_HVT U289 ( .A(n593), .Y(n386) );
  MUX21X1_HVT U290 ( .A1(n314), .A2(n200), .S0(n316), .Y(n579) );
  MUX21X1_HVT U291 ( .A1(n283), .A2(n386), .S0(n316), .Y(n569) );
  MUX21X1_HVT U292 ( .A1(n301), .A2(n387), .S0(n248), .Y(n554) );
  MUX21X1_HVT U293 ( .A1(n387), .A2(n301), .S0(n247), .Y(n400) );
  MUX21X1_HVT U294 ( .A1(n286), .A2(n200), .S0(n248), .Y(n583) );
  MUX21X1_HVT U295 ( .A1(n301), .A2(n303), .S0(n252), .Y(n552) );
  XOR2X1_HVT U296 ( .A1(n593), .A2(n316), .Y(n549) );
  MUX21X1_HVT U297 ( .A1(n302), .A2(n310), .S0(n319), .Y(n557) );
  MUX21X1_HVT U298 ( .A1(n313), .A2(n301), .S0(n247), .Y(n578) );
  XOR2X1_HVT U299 ( .A1(n240), .A2(n248), .Y(n550) );
  AND2X1_HVT U300 ( .A1(n319), .A2(n238), .Y(n278) );
  MUX21X1_HVT U301 ( .A1(n301), .A2(n313), .S0(n247), .Y(n394) );
  MUX21X1_HVT U302 ( .A1(n314), .A2(n238), .S0(n316), .Y(n478) );
  NBUFFX2_HVT U303 ( .A(n246), .Y(n298) );
  NBUFFX2_HVT U304 ( .A(n246), .Y(n300) );
  NAND2X0_HVT U305 ( .A1(n322), .A2(n197), .Y(n499) );
  MUX21X1_HVT U306 ( .A1(n201), .A2(n311), .S0(n252), .Y(n457) );
  MUX21X1_HVT U307 ( .A1(n353), .A2(n253), .S0(n297), .Y(n541) );
  AND2X1_HVT U308 ( .A1(n314), .A2(n322), .Y(n279) );
  AND2X1_HVT U309 ( .A1(n387), .A2(n322), .Y(n280) );
  NBUFFX2_HVT U310 ( .A(n593), .Y(n311) );
  NBUFFX2_HVT U311 ( .A(n264), .Y(n301) );
  XNOR2X1_HVT U312 ( .A1(n328), .A2(n292), .Y(n281) );
  NBUFFX2_HVT U313 ( .A(n323), .Y(n292) );
  NBUFFX2_HVT U314 ( .A(n296), .Y(n291) );
  NBUFFX2_HVT U315 ( .A(n294), .Y(n289) );
  NBUFFX2_HVT U316 ( .A(n296), .Y(n290) );
  NBUFFX2_HVT U317 ( .A(n323), .Y(n294) );
  MUX21X1_HVT U318 ( .A1(n387), .A2(n386), .S0(n247), .Y(n483) );
  MUX21X1_HVT U319 ( .A1(n198), .A2(n263), .S0(n319), .Y(n465) );
  XOR2X1_HVT U320 ( .A1(n248), .A2(n263), .Y(n548) );
  MUX21X1_HVT U321 ( .A1(n263), .A2(n284), .S0(n252), .Y(n573) );
  MUX21X1_HVT U322 ( .A1(n313), .A2(n263), .S0(n247), .Y(n398) );
  MUX21X1_HVT U323 ( .A1(n263), .A2(n314), .S0(n320), .Y(n402) );
  MUX21X1_HVT U324 ( .A1(n263), .A2(n287), .S0(n320), .Y(n580) );
  MUX21X1_HVT U325 ( .A1(n301), .A2(n263), .S0(n319), .Y(n393) );
  MUX21X1_HVT U326 ( .A1(n311), .A2(n263), .S0(n248), .Y(n568) );
  MUX21X1_HVT U327 ( .A1(n263), .A2(n386), .S0(n252), .Y(n403) );
  NBUFFX2_HVT U328 ( .A(n581), .Y(n309) );
  INVX1_HVT U329 ( .A(n575), .Y(n350) );
  MUX21X1_HVT U330 ( .A1(n564), .A2(n276), .S0(n297), .Y(n472) );
  MUX21X1_HVT U331 ( .A1(n197), .A2(n388), .S0(n247), .Y(n564) );
  MUX21X1_HVT U332 ( .A1(n388), .A2(n198), .S0(n316), .Y(n575) );
  INVX1_HVT U333 ( .A(n315), .Y(n282) );
  INVX1_HVT U334 ( .A(n315), .Y(n283) );
  INVX1_HVT U335 ( .A(n288), .Y(n284) );
  INVX0_HVT U336 ( .A(n285), .Y(n287) );
  INVX0_HVT U337 ( .A(n285), .Y(n288) );
  NBUFFX2_HVT U338 ( .A(n597), .Y(n315) );
  INVX1_HVT U339 ( .A(in[1]), .Y(n304) );
  NBUFFX2_HVT U340 ( .A(in[2]), .Y(n323) );
  NBUFFX2_HVT U341 ( .A(n323), .Y(n295) );
  NBUFFX2_HVT U342 ( .A(n323), .Y(n296) );
  NBUFFX2_HVT U343 ( .A(n323), .Y(n297) );
  MUX21X1_HVT U344 ( .A1(n283), .A2(n265), .S0(n247), .Y(n390) );
  MUX21X1_HVT U345 ( .A1(n286), .A2(n265), .S0(n320), .Y(n442) );
  MUX21X1_HVT U346 ( .A1(n265), .A2(n311), .S0(n320), .Y(n395) );
  MUX21X1_HVT U347 ( .A1(n265), .A2(n288), .S0(n320), .Y(n396) );
  MUX21X1_HVT U348 ( .A1(n311), .A2(n265), .S0(n320), .Y(n502) );
  MUX21X1_HVT U349 ( .A1(n303), .A2(n265), .S0(n318), .Y(n570) );
  NBUFFX2_HVT U350 ( .A(n581), .Y(n310) );
  NBUFFX2_HVT U351 ( .A(n595), .Y(n312) );
  NBUFFX2_HVT U352 ( .A(n595), .Y(n314) );
  INVX0_HVT U353 ( .A(n565), .Y(n330) );
  INVX0_HVT U354 ( .A(n559), .Y(n331) );
  INVX0_HVT U355 ( .A(n499), .Y(n332) );
  INVX0_HVT U356 ( .A(n460), .Y(n333) );
  INVX0_HVT U357 ( .A(n592), .Y(n335) );
  INVX0_HVT U358 ( .A(n555), .Y(n336) );
  INVX0_HVT U359 ( .A(n591), .Y(n337) );
  INVX0_HVT U360 ( .A(n590), .Y(n338) );
  INVX0_HVT U361 ( .A(n562), .Y(n339) );
  INVX0_HVT U362 ( .A(n584), .Y(n340) );
  INVX0_HVT U363 ( .A(n589), .Y(n341) );
  INVX0_HVT U364 ( .A(n585), .Y(n342) );
  INVX0_HVT U365 ( .A(n583), .Y(n343) );
  INVX0_HVT U366 ( .A(n582), .Y(n344) );
  INVX0_HVT U367 ( .A(n580), .Y(n345) );
  INVX0_HVT U368 ( .A(n579), .Y(n346) );
  INVX0_HVT U369 ( .A(n578), .Y(n347) );
  INVX0_HVT U370 ( .A(n577), .Y(n348) );
  INVX0_HVT U371 ( .A(n573), .Y(n352) );
  INVX0_HVT U372 ( .A(n571), .Y(n354) );
  INVX0_HVT U373 ( .A(n570), .Y(n355) );
  INVX0_HVT U374 ( .A(n569), .Y(n356) );
  INVX0_HVT U375 ( .A(n568), .Y(n357) );
  INVX0_HVT U376 ( .A(n567), .Y(n358) );
  INVX0_HVT U377 ( .A(n566), .Y(n359) );
  INVX0_HVT U378 ( .A(n564), .Y(n360) );
  INVX0_HVT U379 ( .A(n563), .Y(n361) );
  INVX0_HVT U380 ( .A(n560), .Y(n362) );
  INVX0_HVT U381 ( .A(n558), .Y(n363) );
  INVX0_HVT U382 ( .A(n557), .Y(n364) );
  INVX0_HVT U383 ( .A(n553), .Y(n366) );
  INVX0_HVT U384 ( .A(n551), .Y(n368) );
  INVX0_HVT U385 ( .A(n588), .Y(n369) );
  INVX0_HVT U386 ( .A(n402), .Y(n371) );
  INVX0_HVT U387 ( .A(n399), .Y(n374) );
  INVX0_HVT U388 ( .A(n398), .Y(n375) );
  INVX0_HVT U389 ( .A(n397), .Y(n376) );
  INVX0_HVT U390 ( .A(n396), .Y(n377) );
  INVX0_HVT U391 ( .A(n395), .Y(n378) );
  INVX0_HVT U392 ( .A(n394), .Y(n379) );
  INVX0_HVT U393 ( .A(n393), .Y(n380) );
  INVX0_HVT U394 ( .A(n442), .Y(n381) );
  INVX0_HVT U395 ( .A(n392), .Y(n382) );
  INVX0_HVT U396 ( .A(n391), .Y(n383) );
  INVX0_HVT U397 ( .A(n390), .Y(n384) );
endmodule

