
module add_round_keys_1 ( state, subkey, out );
  input [127:0] state;
  input [127:0] subkey;
  output [127:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233;

  XOR2X2_HVT U2 ( .A1(state[99]), .A2(subkey[99]), .Y(out[99]) );
  XOR2X2_HVT U3 ( .A1(subkey[98]), .A2(state[98]), .Y(out[98]) );
  XOR2X2_HVT U4 ( .A1(subkey[97]), .A2(state[97]), .Y(out[97]) );
  XOR2X2_HVT U5 ( .A1(subkey[96]), .A2(state[96]), .Y(out[96]) );
  XOR2X2_HVT U7 ( .A1(subkey[94]), .A2(state[94]), .Y(out[94]) );
  XOR2X2_HVT U11 ( .A1(subkey[90]), .A2(state[90]), .Y(out[90]) );
  XOR2X2_HVT U12 ( .A1(subkey[8]), .A2(state[8]), .Y(out[8]) );
  XOR2X2_HVT U14 ( .A1(state[88]), .A2(subkey[88]), .Y(out[88]) );
  XOR2X2_HVT U16 ( .A1(state[86]), .A2(subkey[86]), .Y(out[86]) );
  XOR2X2_HVT U20 ( .A1(subkey[82]), .A2(state[82]), .Y(out[82]) );
  XOR2X2_HVT U23 ( .A1(subkey[7]), .A2(state[7]), .Y(out[7]) );
  XOR2X2_HVT U24 ( .A1(subkey[79]), .A2(state[79]), .Y(out[79]) );
  XOR2X2_HVT U25 ( .A1(subkey[78]), .A2(state[78]), .Y(out[78]) );
  XOR2X2_HVT U26 ( .A1(state[77]), .A2(subkey[77]), .Y(out[77]) );
  XOR2X2_HVT U29 ( .A1(subkey[74]), .A2(state[74]), .Y(out[74]) );
  XOR2X2_HVT U32 ( .A1(subkey[71]), .A2(state[71]), .Y(out[71]) );
  XOR2X2_HVT U33 ( .A1(subkey[70]), .A2(state[70]), .Y(out[70]) );
  XOR2X2_HVT U34 ( .A1(subkey[6]), .A2(state[6]), .Y(out[6]) );
  XOR2X2_HVT U38 ( .A1(subkey[66]), .A2(state[66]), .Y(out[66]) );
  XOR2X2_HVT U40 ( .A1(subkey[64]), .A2(state[64]), .Y(out[64]) );
  XOR2X2_HVT U42 ( .A1(subkey[62]), .A2(state[62]), .Y(out[62]) );
  XOR2X2_HVT U47 ( .A1(subkey[58]), .A2(state[58]), .Y(out[58]) );
  XOR2X2_HVT U49 ( .A1(subkey[56]), .A2(state[56]), .Y(out[56]) );
  XOR2X2_HVT U50 ( .A1(state[55]), .A2(subkey[55]), .Y(out[55]) );
  XOR2X2_HVT U58 ( .A1(subkey[48]), .A2(state[48]), .Y(out[48]) );
  XOR2X2_HVT U59 ( .A1(subkey[47]), .A2(state[47]), .Y(out[47]) );
  XOR2X2_HVT U66 ( .A1(subkey[40]), .A2(state[40]), .Y(out[40]) );
  XOR2X2_HVT U75 ( .A1(state[32]), .A2(subkey[32]), .Y(out[32]) );
  XOR2X2_HVT U76 ( .A1(subkey[31]), .A2(state[31]), .Y(out[31]) );
  XOR2X2_HVT U77 ( .A1(subkey[30]), .A2(state[30]), .Y(out[30]) );
  XOR2X2_HVT U78 ( .A1(subkey[2]), .A2(state[2]), .Y(out[2]) );
  XOR2X2_HVT U83 ( .A1(subkey[25]), .A2(state[25]), .Y(out[25]) );
  XOR2X2_HVT U84 ( .A1(state[24]), .A2(subkey[24]), .Y(out[24]) );
  XOR2X2_HVT U85 ( .A1(subkey[23]), .A2(state[23]), .Y(out[23]) );
  XOR2X2_HVT U86 ( .A1(state[22]), .A2(subkey[22]), .Y(out[22]) );
  XOR2X2_HVT U87 ( .A1(subkey[21]), .A2(state[21]), .Y(out[21]) );
  XOR2X2_HVT U89 ( .A1(subkey[1]), .A2(state[1]), .Y(out[1]) );
  XOR2X2_HVT U91 ( .A1(subkey[18]), .A2(state[18]), .Y(out[18]) );
  XOR2X2_HVT U93 ( .A1(subkey[16]), .A2(state[16]), .Y(out[16]) );
  XOR2X2_HVT U94 ( .A1(state[15]), .A2(subkey[15]), .Y(out[15]) );
  XOR2X2_HVT U95 ( .A1(subkey[14]), .A2(state[14]), .Y(out[14]) );
  XOR2X2_HVT U96 ( .A1(subkey[13]), .A2(state[13]), .Y(out[13]) );
  XOR2X2_HVT U101 ( .A1(subkey[124]), .A2(state[124]), .Y(out[124]) );
  XOR2X2_HVT U103 ( .A1(subkey[122]), .A2(state[122]), .Y(out[122]) );
  XOR2X2_HVT U104 ( .A1(subkey[121]), .A2(state[121]), .Y(out[121]) );
  XOR2X2_HVT U105 ( .A1(state[120]), .A2(subkey[120]), .Y(out[120]) );
  XOR2X2_HVT U109 ( .A1(subkey[117]), .A2(state[117]), .Y(out[117]) );
  XOR2X2_HVT U113 ( .A1(state[113]), .A2(subkey[113]), .Y(out[113]) );
  XOR2X2_HVT U116 ( .A1(subkey[110]), .A2(state[110]), .Y(out[110]) );
  XOR2X2_HVT U117 ( .A1(state[10]), .A2(subkey[10]), .Y(out[10]) );
  XOR2X2_HVT U118 ( .A1(subkey[109]), .A2(state[109]), .Y(out[109]) );
  XOR2X2_HVT U121 ( .A1(subkey[106]), .A2(state[106]), .Y(out[106]) );
  XOR2X2_HVT U122 ( .A1(subkey[105]), .A2(state[105]), .Y(out[105]) );
  XOR2X2_HVT U124 ( .A1(subkey[103]), .A2(state[103]), .Y(out[103]) );
  XOR2X2_HVT U126 ( .A1(subkey[101]), .A2(state[101]), .Y(out[101]) );
  XOR2X2_HVT U128 ( .A1(state[0]), .A2(subkey[0]), .Y(out[0]) );
  XOR2X1_HVT U1 ( .A1(state[112]), .A2(subkey[112]), .Y(out[112]) );
  INVX2_HVT U6 ( .A(subkey[19]), .Y(n62) );
  NAND2X0_HVT U8 ( .A1(state[37]), .A2(n2), .Y(n3) );
  NAND2X0_HVT U9 ( .A1(n1), .A2(subkey[37]), .Y(n4) );
  NAND2X0_HVT U10 ( .A1(n3), .A2(n4), .Y(out[37]) );
  INVX0_HVT U13 ( .A(state[37]), .Y(n1) );
  INVX0_HVT U15 ( .A(subkey[37]), .Y(n2) );
  NAND2X0_HVT U17 ( .A1(subkey[104]), .A2(n6), .Y(n7) );
  NAND2X0_HVT U18 ( .A1(n5), .A2(state[104]), .Y(n8) );
  NAND2X0_HVT U19 ( .A1(n7), .A2(n8), .Y(out[104]) );
  IBUFFX2_HVT U21 ( .A(subkey[104]), .Y(n5) );
  INVX0_HVT U22 ( .A(state[104]), .Y(n6) );
  NAND2X0_HVT U27 ( .A1(subkey[50]), .A2(n10), .Y(n11) );
  NAND2X0_HVT U28 ( .A1(n9), .A2(state[50]), .Y(n12) );
  NAND2X0_HVT U30 ( .A1(n11), .A2(n12), .Y(out[50]) );
  IBUFFX2_HVT U31 ( .A(subkey[50]), .Y(n9) );
  INVX0_HVT U35 ( .A(state[50]), .Y(n10) );
  NAND2X0_HVT U36 ( .A1(state[4]), .A2(n14), .Y(n15) );
  NAND2X0_HVT U37 ( .A1(n13), .A2(subkey[4]), .Y(n16) );
  NAND2X0_HVT U39 ( .A1(n15), .A2(n16), .Y(out[4]) );
  INVX0_HVT U41 ( .A(state[4]), .Y(n13) );
  IBUFFX2_HVT U43 ( .A(subkey[4]), .Y(n14) );
  XNOR2X2_HVT U44 ( .A1(state[93]), .A2(n17), .Y(out[93]) );
  IBUFFX16_HVT U45 ( .A(subkey[93]), .Y(n17) );
  NAND2X0_HVT U46 ( .A1(subkey[45]), .A2(n19), .Y(n20) );
  NAND2X0_HVT U48 ( .A1(n18), .A2(state[45]), .Y(n21) );
  NAND2X0_HVT U51 ( .A1(n20), .A2(n21), .Y(out[45]) );
  INVX0_HVT U52 ( .A(subkey[45]), .Y(n18) );
  INVX0_HVT U53 ( .A(state[45]), .Y(n19) );
  XNOR2X2_HVT U54 ( .A1(n22), .A2(state[100]), .Y(out[100]) );
  IBUFFX16_HVT U55 ( .A(subkey[100]), .Y(n22) );
  NAND2X0_HVT U56 ( .A1(state[28]), .A2(n27), .Y(n25) );
  NAND2X0_HVT U57 ( .A1(n23), .A2(n24), .Y(n26) );
  NAND2X0_HVT U60 ( .A1(n25), .A2(n26), .Y(out[28]) );
  INVX0_HVT U61 ( .A(state[28]), .Y(n23) );
  INVX16_HVT U62 ( .A(n27), .Y(n24) );
  IBUFFX16_HVT U63 ( .A(subkey[28]), .Y(n27) );
  XNOR2X2_HVT U64 ( .A1(state[115]), .A2(n28), .Y(out[115]) );
  IBUFFX16_HVT U65 ( .A(subkey[115]), .Y(n28) );
  NAND2X0_HVT U67 ( .A1(state[19]), .A2(n62), .Y(n31) );
  NAND2X0_HVT U68 ( .A1(n29), .A2(n30), .Y(n32) );
  NAND2X0_HVT U69 ( .A1(n31), .A2(n32), .Y(out[19]) );
  INVX0_HVT U70 ( .A(state[19]), .Y(n29) );
  INVX0_HVT U71 ( .A(n62), .Y(n30) );
  NAND2X0_HVT U72 ( .A1(state[89]), .A2(n61), .Y(n35) );
  NAND2X0_HVT U73 ( .A1(n33), .A2(n34), .Y(n36) );
  NAND2X0_HVT U74 ( .A1(n35), .A2(n36), .Y(out[89]) );
  INVX0_HVT U79 ( .A(state[89]), .Y(n33) );
  INVX0_HVT U80 ( .A(n61), .Y(n34) );
  IBUFFX2_HVT U81 ( .A(subkey[89]), .Y(n61) );
  NAND2X0_HVT U82 ( .A1(subkey[53]), .A2(n38), .Y(n39) );
  NAND2X0_HVT U88 ( .A1(n37), .A2(state[53]), .Y(n40) );
  NAND2X0_HVT U90 ( .A1(n39), .A2(n40), .Y(out[53]) );
  IBUFFX2_HVT U92 ( .A(subkey[53]), .Y(n37) );
  INVX0_HVT U97 ( .A(state[53]), .Y(n38) );
  NAND2X0_HVT U98 ( .A1(subkey[11]), .A2(n42), .Y(n43) );
  NAND2X0_HVT U99 ( .A1(n41), .A2(state[11]), .Y(n44) );
  NAND2X0_HVT U100 ( .A1(n43), .A2(n44), .Y(out[11]) );
  IBUFFX2_HVT U102 ( .A(subkey[11]), .Y(n41) );
  INVX0_HVT U106 ( .A(state[11]), .Y(n42) );
  INVX1_HVT U107 ( .A(subkey[76]), .Y(n123) );
  NAND2X0_HVT U108 ( .A1(subkey[20]), .A2(n46), .Y(n47) );
  NAND2X0_HVT U110 ( .A1(n45), .A2(state[20]), .Y(n48) );
  NAND2X0_HVT U111 ( .A1(n47), .A2(n48), .Y(out[20]) );
  IBUFFX2_HVT U112 ( .A(subkey[20]), .Y(n45) );
  INVX0_HVT U114 ( .A(state[20]), .Y(n46) );
  NAND2X0_HVT U115 ( .A1(state[34]), .A2(n50), .Y(n51) );
  NAND2X0_HVT U119 ( .A1(n49), .A2(subkey[34]), .Y(n52) );
  NAND2X0_HVT U120 ( .A1(n51), .A2(n52), .Y(out[34]) );
  INVX0_HVT U123 ( .A(state[34]), .Y(n49) );
  INVX0_HVT U125 ( .A(subkey[34]), .Y(n50) );
  NAND2X0_HVT U127 ( .A1(subkey[72]), .A2(n54), .Y(n55) );
  NAND2X0_HVT U129 ( .A1(n53), .A2(state[72]), .Y(n56) );
  NAND2X0_HVT U130 ( .A1(n55), .A2(n56), .Y(out[72]) );
  INVX0_HVT U131 ( .A(subkey[72]), .Y(n53) );
  INVX0_HVT U132 ( .A(state[72]), .Y(n54) );
  XOR2X2_HVT U133 ( .A1(state[42]), .A2(subkey[42]), .Y(out[42]) );
  NAND2X0_HVT U134 ( .A1(state[12]), .A2(n58), .Y(n59) );
  NAND2X0_HVT U135 ( .A1(n57), .A2(subkey[12]), .Y(n60) );
  NAND2X0_HVT U136 ( .A1(n59), .A2(n60), .Y(out[12]) );
  INVX0_HVT U137 ( .A(state[12]), .Y(n57) );
  INVX0_HVT U138 ( .A(subkey[12]), .Y(n58) );
  INVX0_HVT U139 ( .A(subkey[108]), .Y(n91) );
  OR2X1_HVT U140 ( .A1(n198), .A2(state[35]), .Y(n192) );
  INVX0_HVT U141 ( .A(subkey[69]), .Y(n71) );
  XOR2X2_HVT U142 ( .A1(subkey[102]), .A2(state[102]), .Y(out[102]) );
  XOR2X2_HVT U143 ( .A1(subkey[118]), .A2(state[118]), .Y(out[118]) );
  NAND2X0_HVT U144 ( .A1(subkey[87]), .A2(n64), .Y(n65) );
  NAND2X0_HVT U145 ( .A1(n63), .A2(state[87]), .Y(n66) );
  NAND2X0_HVT U146 ( .A1(n65), .A2(n66), .Y(out[87]) );
  IBUFFX2_HVT U147 ( .A(subkey[87]), .Y(n63) );
  INVX0_HVT U148 ( .A(state[87]), .Y(n64) );
  NAND2X0_HVT U149 ( .A1(subkey[80]), .A2(n68), .Y(n69) );
  NAND2X0_HVT U150 ( .A1(n67), .A2(state[80]), .Y(n70) );
  NAND2X0_HVT U151 ( .A1(n69), .A2(n70), .Y(out[80]) );
  INVX0_HVT U152 ( .A(subkey[80]), .Y(n67) );
  INVX0_HVT U153 ( .A(state[80]), .Y(n68) );
  NAND2X0_HVT U154 ( .A1(subkey[69]), .A2(n72), .Y(n73) );
  NAND2X0_HVT U155 ( .A1(n71), .A2(state[69]), .Y(n74) );
  NAND2X0_HVT U156 ( .A1(n73), .A2(n74), .Y(out[69]) );
  INVX0_HVT U157 ( .A(state[69]), .Y(n72) );
  NAND2X0_HVT U158 ( .A1(state[26]), .A2(n76), .Y(n77) );
  NAND2X0_HVT U159 ( .A1(n75), .A2(subkey[26]), .Y(n78) );
  NAND2X0_HVT U160 ( .A1(n77), .A2(n78), .Y(out[26]) );
  INVX0_HVT U161 ( .A(state[26]), .Y(n75) );
  IBUFFX2_HVT U162 ( .A(subkey[26]), .Y(n76) );
  NAND2X0_HVT U163 ( .A1(subkey[9]), .A2(n80), .Y(n81) );
  NAND2X0_HVT U164 ( .A1(n79), .A2(state[9]), .Y(n82) );
  NAND2X0_HVT U165 ( .A1(n81), .A2(n82), .Y(out[9]) );
  INVX0_HVT U166 ( .A(subkey[9]), .Y(n79) );
  INVX0_HVT U167 ( .A(state[9]), .Y(n80) );
  NAND2X0_HVT U168 ( .A1(subkey[95]), .A2(n84), .Y(n85) );
  NAND2X0_HVT U169 ( .A1(n83), .A2(state[95]), .Y(n86) );
  NAND2X0_HVT U170 ( .A1(n85), .A2(n86), .Y(out[95]) );
  INVX0_HVT U171 ( .A(subkey[95]), .Y(n83) );
  INVX0_HVT U172 ( .A(state[95]), .Y(n84) );
  NAND2X0_HVT U173 ( .A1(state[59]), .A2(n193), .Y(n89) );
  NAND2X0_HVT U174 ( .A1(n87), .A2(n88), .Y(n90) );
  NAND2X0_HVT U175 ( .A1(n89), .A2(n90), .Y(out[59]) );
  INVX0_HVT U176 ( .A(state[59]), .Y(n87) );
  INVX0_HVT U177 ( .A(n193), .Y(n88) );
  INVX0_HVT U178 ( .A(subkey[59]), .Y(n193) );
  NAND2X0_HVT U179 ( .A1(subkey[108]), .A2(n92), .Y(n93) );
  NAND2X0_HVT U180 ( .A1(n91), .A2(state[108]), .Y(n94) );
  NAND2X0_HVT U181 ( .A1(n93), .A2(n94), .Y(out[108]) );
  INVX0_HVT U182 ( .A(state[108]), .Y(n92) );
  XOR2X2_HVT U183 ( .A1(subkey[114]), .A2(state[114]), .Y(out[114]) );
  INVX0_HVT U184 ( .A(subkey[92]), .Y(n119) );
  INVX0_HVT U185 ( .A(subkey[91]), .Y(n159) );
  INVX0_HVT U186 ( .A(subkey[61]), .Y(n95) );
  INVX0_HVT U187 ( .A(subkey[38]), .Y(n204) );
  INVX0_HVT U188 ( .A(subkey[33]), .Y(n209) );
  INVX0_HVT U189 ( .A(subkey[111]), .Y(n199) );
  NAND2X0_HVT U190 ( .A1(subkey[61]), .A2(n96), .Y(n97) );
  NAND2X0_HVT U191 ( .A1(n95), .A2(state[61]), .Y(n98) );
  NAND2X0_HVT U192 ( .A1(n97), .A2(n98), .Y(out[61]) );
  INVX0_HVT U193 ( .A(state[61]), .Y(n96) );
  NAND2X0_HVT U194 ( .A1(subkey[65]), .A2(n100), .Y(n101) );
  NAND2X0_HVT U195 ( .A1(state[65]), .A2(n99), .Y(n102) );
  NAND2X0_HVT U196 ( .A1(n101), .A2(n102), .Y(out[65]) );
  INVX0_HVT U197 ( .A(subkey[65]), .Y(n99) );
  INVX0_HVT U198 ( .A(state[65]), .Y(n100) );
  NAND2X0_HVT U199 ( .A1(state[83]), .A2(n104), .Y(n105) );
  NAND2X0_HVT U200 ( .A1(n103), .A2(subkey[83]), .Y(n106) );
  NAND2X0_HVT U201 ( .A1(n105), .A2(n106), .Y(out[83]) );
  INVX0_HVT U202 ( .A(state[83]), .Y(n103) );
  INVX0_HVT U203 ( .A(subkey[83]), .Y(n104) );
  NAND2X0_HVT U204 ( .A1(subkey[85]), .A2(n108), .Y(n109) );
  NAND2X0_HVT U205 ( .A1(n107), .A2(state[85]), .Y(n110) );
  NAND2X0_HVT U206 ( .A1(n109), .A2(n110), .Y(out[85]) );
  INVX0_HVT U207 ( .A(subkey[85]), .Y(n107) );
  INVX0_HVT U208 ( .A(state[85]), .Y(n108) );
  NAND2X0_HVT U209 ( .A1(subkey[17]), .A2(n112), .Y(n113) );
  NAND2X0_HVT U210 ( .A1(n111), .A2(state[17]), .Y(n114) );
  NAND2X0_HVT U211 ( .A1(n113), .A2(n114), .Y(out[17]) );
  INVX0_HVT U212 ( .A(subkey[17]), .Y(n111) );
  INVX0_HVT U213 ( .A(state[17]), .Y(n112) );
  NAND2X0_HVT U214 ( .A1(subkey[46]), .A2(n116), .Y(n117) );
  NAND2X0_HVT U215 ( .A1(n115), .A2(state[46]), .Y(n118) );
  NAND2X0_HVT U216 ( .A1(n117), .A2(n118), .Y(out[46]) );
  INVX0_HVT U217 ( .A(subkey[46]), .Y(n115) );
  INVX0_HVT U218 ( .A(state[46]), .Y(n116) );
  NAND2X0_HVT U219 ( .A1(subkey[92]), .A2(n120), .Y(n121) );
  NAND2X0_HVT U220 ( .A1(n119), .A2(state[92]), .Y(n122) );
  NAND2X0_HVT U221 ( .A1(n121), .A2(n122), .Y(out[92]) );
  INVX0_HVT U222 ( .A(state[92]), .Y(n120) );
  NAND2X0_HVT U223 ( .A1(subkey[76]), .A2(n124), .Y(n125) );
  NAND2X0_HVT U224 ( .A1(state[76]), .A2(n123), .Y(n126) );
  NAND2X0_HVT U225 ( .A1(n125), .A2(n126), .Y(out[76]) );
  INVX0_HVT U226 ( .A(state[76]), .Y(n124) );
  XOR2X2_HVT U227 ( .A1(subkey[119]), .A2(state[119]), .Y(out[119]) );
  NAND2X0_HVT U228 ( .A1(subkey[68]), .A2(n128), .Y(n129) );
  NAND2X0_HVT U229 ( .A1(n127), .A2(state[68]), .Y(n130) );
  NAND2X0_HVT U230 ( .A1(n129), .A2(n130), .Y(out[68]) );
  INVX0_HVT U231 ( .A(subkey[68]), .Y(n127) );
  INVX0_HVT U232 ( .A(state[68]), .Y(n128) );
  XOR2X2_HVT U233 ( .A1(subkey[126]), .A2(state[126]), .Y(out[126]) );
  NAND2X0_HVT U234 ( .A1(subkey[52]), .A2(n132), .Y(n133) );
  NAND2X0_HVT U235 ( .A1(n131), .A2(state[52]), .Y(n134) );
  NAND2X0_HVT U236 ( .A1(n133), .A2(n134), .Y(out[52]) );
  INVX0_HVT U237 ( .A(subkey[52]), .Y(n131) );
  INVX0_HVT U238 ( .A(state[52]), .Y(n132) );
  NAND2X0_HVT U239 ( .A1(subkey[44]), .A2(n136), .Y(n137) );
  NAND2X0_HVT U240 ( .A1(n135), .A2(state[44]), .Y(n138) );
  NAND2X0_HVT U241 ( .A1(n137), .A2(n138), .Y(out[44]) );
  INVX0_HVT U242 ( .A(subkey[44]), .Y(n135) );
  INVX0_HVT U243 ( .A(state[44]), .Y(n136) );
  NAND2X0_HVT U244 ( .A1(subkey[125]), .A2(n140), .Y(n141) );
  NAND2X0_HVT U245 ( .A1(n139), .A2(state[125]), .Y(n142) );
  NAND2X0_HVT U246 ( .A1(n141), .A2(n142), .Y(out[125]) );
  INVX0_HVT U247 ( .A(subkey[125]), .Y(n139) );
  INVX0_HVT U248 ( .A(state[125]), .Y(n140) );
  NAND2X0_HVT U249 ( .A1(n144), .A2(state[75]), .Y(n145) );
  NAND2X0_HVT U250 ( .A1(n143), .A2(subkey[75]), .Y(n146) );
  NAND2X0_HVT U251 ( .A1(n146), .A2(n145), .Y(out[75]) );
  INVX0_HVT U252 ( .A(state[75]), .Y(n143) );
  INVX0_HVT U253 ( .A(subkey[75]), .Y(n144) );
  NAND2X0_HVT U254 ( .A1(state[3]), .A2(n148), .Y(n149) );
  NAND2X0_HVT U255 ( .A1(n147), .A2(subkey[3]), .Y(n150) );
  NAND2X0_HVT U256 ( .A1(n149), .A2(n150), .Y(out[3]) );
  INVX0_HVT U257 ( .A(state[3]), .Y(n147) );
  INVX0_HVT U258 ( .A(subkey[3]), .Y(n148) );
  NAND2X0_HVT U259 ( .A1(state[41]), .A2(n152), .Y(n153) );
  NAND2X0_HVT U260 ( .A1(n151), .A2(subkey[41]), .Y(n154) );
  NAND2X0_HVT U261 ( .A1(n153), .A2(n154), .Y(out[41]) );
  INVX0_HVT U262 ( .A(state[41]), .Y(n151) );
  INVX0_HVT U263 ( .A(subkey[41]), .Y(n152) );
  INVX1_HVT U264 ( .A(subkey[60]), .Y(n208) );
  NAND2X0_HVT U265 ( .A1(n156), .A2(state[51]), .Y(n157) );
  NAND2X0_HVT U266 ( .A1(n155), .A2(subkey[51]), .Y(n158) );
  NAND2X0_HVT U267 ( .A1(n157), .A2(n158), .Y(out[51]) );
  INVX0_HVT U268 ( .A(state[51]), .Y(n155) );
  INVX0_HVT U269 ( .A(subkey[51]), .Y(n156) );
  NAND2X0_HVT U270 ( .A1(subkey[91]), .A2(n160), .Y(n161) );
  NAND2X0_HVT U271 ( .A1(state[91]), .A2(n159), .Y(n162) );
  NAND2X0_HVT U272 ( .A1(n161), .A2(n162), .Y(out[91]) );
  INVX0_HVT U273 ( .A(state[91]), .Y(n160) );
  INVX1_HVT U274 ( .A(subkey[35]), .Y(n198) );
  NAND2X0_HVT U275 ( .A1(subkey[54]), .A2(n164), .Y(n165) );
  NAND2X0_HVT U276 ( .A1(n163), .A2(state[54]), .Y(n166) );
  NAND2X0_HVT U277 ( .A1(n165), .A2(n166), .Y(out[54]) );
  INVX0_HVT U278 ( .A(subkey[54]), .Y(n163) );
  INVX0_HVT U279 ( .A(state[54]), .Y(n164) );
  NAND2X0_HVT U280 ( .A1(state[84]), .A2(n168), .Y(n169) );
  NAND2X0_HVT U281 ( .A1(n167), .A2(subkey[84]), .Y(n170) );
  NAND2X0_HVT U282 ( .A1(n169), .A2(n170), .Y(out[84]) );
  INVX0_HVT U283 ( .A(state[84]), .Y(n167) );
  INVX0_HVT U284 ( .A(subkey[84]), .Y(n168) );
  NAND2X0_HVT U285 ( .A1(subkey[73]), .A2(n172), .Y(n173) );
  NAND2X0_HVT U286 ( .A1(n171), .A2(state[73]), .Y(n174) );
  NAND2X0_HVT U287 ( .A1(n173), .A2(n174), .Y(out[73]) );
  INVX0_HVT U288 ( .A(subkey[73]), .Y(n171) );
  INVX0_HVT U289 ( .A(state[73]), .Y(n172) );
  NAND2X0_HVT U290 ( .A1(subkey[107]), .A2(n176), .Y(n177) );
  NAND2X0_HVT U291 ( .A1(n175), .A2(state[107]), .Y(n178) );
  NAND2X0_HVT U292 ( .A1(n177), .A2(n178), .Y(out[107]) );
  IBUFFX2_HVT U293 ( .A(subkey[107]), .Y(n175) );
  INVX0_HVT U294 ( .A(state[107]), .Y(n176) );
  NAND2X0_HVT U295 ( .A1(subkey[57]), .A2(n180), .Y(n181) );
  NAND2X0_HVT U296 ( .A1(state[57]), .A2(n179), .Y(n182) );
  NAND2X0_HVT U297 ( .A1(n181), .A2(n182), .Y(out[57]) );
  INVX0_HVT U298 ( .A(subkey[57]), .Y(n179) );
  INVX0_HVT U299 ( .A(state[57]), .Y(n180) );
  NAND2X0_HVT U300 ( .A1(subkey[63]), .A2(n184), .Y(n185) );
  NAND2X0_HVT U301 ( .A1(state[63]), .A2(n183), .Y(n186) );
  NAND2X0_HVT U302 ( .A1(n185), .A2(n186), .Y(out[63]) );
  INVX0_HVT U303 ( .A(subkey[63]), .Y(n183) );
  INVX0_HVT U304 ( .A(state[63]), .Y(n184) );
  NAND2X0_HVT U305 ( .A1(subkey[81]), .A2(n188), .Y(n189) );
  NAND2X0_HVT U306 ( .A1(state[81]), .A2(n187), .Y(n190) );
  NAND2X0_HVT U307 ( .A1(n190), .A2(n189), .Y(out[81]) );
  INVX0_HVT U308 ( .A(subkey[81]), .Y(n187) );
  INVX0_HVT U309 ( .A(state[81]), .Y(n188) );
  NAND2X0_HVT U310 ( .A1(n198), .A2(state[35]), .Y(n191) );
  NAND2X0_HVT U311 ( .A1(n191), .A2(n192), .Y(out[35]) );
  NAND2X0_HVT U312 ( .A1(subkey[49]), .A2(n195), .Y(n196) );
  NAND2X0_HVT U313 ( .A1(state[49]), .A2(n194), .Y(n197) );
  NAND2X0_HVT U314 ( .A1(n196), .A2(n197), .Y(out[49]) );
  INVX0_HVT U315 ( .A(subkey[49]), .Y(n194) );
  INVX0_HVT U316 ( .A(state[49]), .Y(n195) );
  XNOR2X2_HVT U317 ( .A1(state[111]), .A2(n199), .Y(out[111]) );
  NAND2X0_HVT U318 ( .A1(subkey[39]), .A2(n201), .Y(n202) );
  NAND2X0_HVT U319 ( .A1(state[39]), .A2(n200), .Y(n203) );
  NAND2X0_HVT U320 ( .A1(n202), .A2(n203), .Y(out[39]) );
  INVX0_HVT U321 ( .A(subkey[39]), .Y(n200) );
  INVX0_HVT U322 ( .A(state[39]), .Y(n201) );
  NAND2X0_HVT U323 ( .A1(subkey[38]), .A2(n205), .Y(n206) );
  NAND2X0_HVT U324 ( .A1(n204), .A2(state[38]), .Y(n207) );
  NAND2X0_HVT U325 ( .A1(n206), .A2(n207), .Y(out[38]) );
  INVX0_HVT U326 ( .A(state[38]), .Y(n205) );
  XNOR2X2_HVT U327 ( .A1(state[60]), .A2(n208), .Y(out[60]) );
  XOR2X2_HVT U328 ( .A1(subkey[127]), .A2(state[127]), .Y(out[127]) );
  NAND2X0_HVT U329 ( .A1(subkey[33]), .A2(n210), .Y(n211) );
  NAND2X0_HVT U330 ( .A1(n209), .A2(state[33]), .Y(n212) );
  NAND2X0_HVT U331 ( .A1(n211), .A2(n212), .Y(out[33]) );
  INVX0_HVT U332 ( .A(state[33]), .Y(n210) );
  INVX0_HVT U333 ( .A(subkey[116]), .Y(n213) );
  INVX0_HVT U334 ( .A(subkey[67]), .Y(n214) );
  INVX0_HVT U335 ( .A(subkey[36]), .Y(n218) );
  XOR2X2_HVT U336 ( .A1(subkey[29]), .A2(state[29]), .Y(out[29]) );
  XNOR2X2_HVT U337 ( .A1(state[116]), .A2(n213), .Y(out[116]) );
  NAND2X0_HVT U338 ( .A1(subkey[67]), .A2(n215), .Y(n216) );
  NAND2X0_HVT U339 ( .A1(n214), .A2(state[67]), .Y(n217) );
  NAND2X0_HVT U340 ( .A1(n216), .A2(n217), .Y(out[67]) );
  INVX0_HVT U341 ( .A(state[67]), .Y(n215) );
  XOR2X2_HVT U342 ( .A1(subkey[5]), .A2(state[5]), .Y(out[5]) );
  INVX0_HVT U343 ( .A(subkey[43]), .Y(n222) );
  NAND2X0_HVT U344 ( .A1(subkey[36]), .A2(n219), .Y(n220) );
  NAND2X0_HVT U345 ( .A1(n218), .A2(state[36]), .Y(n221) );
  NAND2X0_HVT U346 ( .A1(n221), .A2(n220), .Y(out[36]) );
  INVX0_HVT U347 ( .A(state[36]), .Y(n219) );
  NAND2X0_HVT U348 ( .A1(subkey[43]), .A2(n223), .Y(n224) );
  NAND2X0_HVT U349 ( .A1(state[43]), .A2(n222), .Y(n225) );
  NAND2X0_HVT U350 ( .A1(n224), .A2(n225), .Y(out[43]) );
  INVX0_HVT U351 ( .A(state[43]), .Y(n223) );
  NAND2X0_HVT U352 ( .A1(subkey[27]), .A2(n227), .Y(n228) );
  NAND2X0_HVT U353 ( .A1(n226), .A2(state[27]), .Y(n229) );
  NAND2X0_HVT U354 ( .A1(n228), .A2(n229), .Y(out[27]) );
  INVX0_HVT U355 ( .A(subkey[27]), .Y(n226) );
  INVX0_HVT U356 ( .A(state[27]), .Y(n227) );
  NAND2X0_HVT U357 ( .A1(subkey[123]), .A2(n231), .Y(n232) );
  NAND2X0_HVT U358 ( .A1(n230), .A2(state[123]), .Y(n233) );
  NAND2X0_HVT U359 ( .A1(n232), .A2(n233), .Y(out[123]) );
  INVX0_HVT U360 ( .A(subkey[123]), .Y(n230) );
  INVX0_HVT U361 ( .A(state[123]), .Y(n231) );
endmodule

