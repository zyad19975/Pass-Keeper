
module sbox_1 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n19, n23, n48, n50, n210, n211, n212, n213, n216, n217, n218, n219,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626;

  NAND2X0_HVT U3 ( .A1(n337), .A2(n331), .Y(n624) );
  NAND2X0_HVT U4 ( .A1(n245), .A2(n624), .Y(n623) );
  NAND2X0_HVT U5 ( .A1(n339), .A2(n405), .Y(n621) );
  NAND2X0_HVT U13 ( .A1(n613), .A2(n333), .Y(n614) );
  NAND2X0_HVT U15 ( .A1(n624), .A2(n322), .Y(n611) );
  NAND2X0_HVT U21 ( .A1(n246), .A2(n341), .Y(n606) );
  NAND2X0_HVT U24 ( .A1(n326), .A2(n341), .Y(n604) );
  NAND2X0_HVT U33 ( .A1(n242), .A2(n341), .Y(n595) );
  NAND2X0_HVT U35 ( .A1(n324), .A2(n341), .Y(n593) );
  NAND2X0_HVT U42 ( .A1(n335), .A2(n326), .Y(n586) );
  MUX41X1_HVT U51 ( .A1(n391), .A3(n352), .A2(n367), .A4(n368), .S0(n263), 
        .S1(n319), .Y(n579) );
  NAND2X0_HVT U53 ( .A1(n576), .A2(n585), .Y(n577) );
  NAND2X0_HVT U56 ( .A1(n246), .A2(n572), .Y(n573) );
  MUX41X1_HVT U57 ( .A1(n392), .A3(n608), .A2(n573), .A4(n616), .S0(n262), 
        .S1(n319), .Y(n571) );
  NAND2X0_HVT U58 ( .A1(n333), .A2(n624), .Y(n570) );
  MUX41X1_HVT U61 ( .A1(n309), .A3(n267), .A2(n366), .A4(n322), .S0(n262), 
        .S1(n319), .Y(n567) );
  NAND2X0_HVT U62 ( .A1(n341), .A2(n332), .Y(n566) );
  MUX41X1_HVT U63 ( .A1(n566), .A3(n359), .A2(n386), .A4(n365), .S0(n350), 
        .S1(n319), .Y(n565) );
  AO21X1_HVT U66 ( .A1(n19), .A2(n346), .A3(n385), .Y(n562) );
  MUX41X1_HVT U68 ( .A1(n362), .A3(n562), .A2(n561), .A4(n563), .S0(n298), 
        .S1(n349), .Y(n560) );
  MUX41X1_HVT U69 ( .A1(n560), .A3(n568), .A2(n564), .A4(n574), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n328), .A2(n555), .Y(n556) );
  MUX41X1_HVT U74 ( .A1(n557), .A3(n602), .A2(n556), .A4(n604), .S0(n315), 
        .S1(n261), .Y(n554) );
  MUX41X1_HVT U75 ( .A1(n389), .A3(n394), .A2(n407), .A4(n272), .S0(n298), 
        .S1(n263), .Y(n553) );
  MUX41X1_HVT U77 ( .A1(n618), .A3(n396), .A2(n552), .A4(n395), .S0(n321), 
        .S1(n343), .Y(n551) );
  AND3X1_HVT U80 ( .A1(n331), .A2(n572), .A3(n547), .Y(n548) );
  MUX41X1_HVT U82 ( .A1(n583), .A3(n368), .A2(n353), .A4(n612), .S0(n316), 
        .S1(n261), .Y(n545) );
  AND2X1_HVT U83 ( .A1(n336), .A2(n270), .Y(n544) );
  MUX41X1_HVT U84 ( .A1(n369), .A3(n620), .A2(n610), .A4(n544), .S0(n316), 
        .S1(n263), .Y(n543) );
  NAND2X0_HVT U85 ( .A1(n341), .A2(n406), .Y(n542) );
  MUX41X1_HVT U86 ( .A1(n394), .A3(n542), .A2(n307), .A4(n306), .S0(n298), 
        .S1(n350), .Y(n541) );
  MUX41X1_HVT U90 ( .A1(n582), .A3(n586), .A2(n391), .A4(n539), .S0(n314), 
        .S1(n349), .Y(n538) );
  AO21X1_HVT U93 ( .A1(n321), .A2(n534), .A3(n390), .Y(n535) );
  MUX41X1_HVT U96 ( .A1(n353), .A3(n308), .A2(n393), .A4(n532), .S0(n298), 
        .S1(n262), .Y(n531) );
  MUX41X1_HVT U97 ( .A1(n389), .A3(n308), .A2(n335), .A4(n611), .S0(n298), 
        .S1(n349), .Y(n530) );
  MUX41X1_HVT U98 ( .A1(n530), .A3(n533), .A2(n531), .A4(n538), .S0(n325), 
        .S1(n346), .Y(n529) );
  NAND2X0_HVT U101 ( .A1(n525), .A2(n524), .Y(n526) );
  MUX41X1_HVT U103 ( .A1(n624), .A3(n363), .A2(n372), .A4(n593), .S0(n298), 
        .S1(n262), .Y(n522) );
  MUX41X1_HVT U105 ( .A1(n371), .A3(n581), .A2(n521), .A4(n388), .S0(n317), 
        .S1(n349), .Y(n520) );
  MUX41X1_HVT U106 ( .A1(n520), .A3(n523), .A2(n522), .A4(n527), .S0(in[0]), 
        .S1(in[5]), .Y(n519) );
  NAND2X0_HVT U110 ( .A1(n331), .A2(n515), .Y(n516) );
  AND2X1_HVT U115 ( .A1(n335), .A2(n322), .Y(n510) );
  NAND2X0_HVT U123 ( .A1(n501), .A2(n500), .Y(n502) );
  MUX41X1_HVT U125 ( .A1(n606), .A3(n313), .A2(n362), .A4(n398), .S0(n314), 
        .S1(n261), .Y(n498) );
  MUX41X1_HVT U131 ( .A1(n493), .A3(n495), .A2(n494), .A4(n496), .S0(in[5]), 
        .S1(n262), .Y(n492) );
  MUX41X1_HVT U136 ( .A1(n306), .A3(n595), .A2(n400), .A4(n592), .S0(n314), 
        .S1(n348), .Y(n488) );
  MUX41X1_HVT U139 ( .A1(n486), .A3(n489), .A2(n488), .A4(n490), .S0(n325), 
        .S1(n346), .Y(n485) );
  AND2X1_HVT U140 ( .A1(n327), .A2(n340), .Y(n484) );
  MUX41X1_HVT U141 ( .A1(n603), .A3(n380), .A2(n484), .A4(n376), .S0(n315), 
        .S1(n348), .Y(n483) );
  MUX41X1_HVT U142 ( .A1(n369), .A3(n323), .A2(n387), .A4(n327), .S0(n314), 
        .S1(n348), .Y(n482) );
  NAND2X0_HVT U146 ( .A1(n339), .A2(n334), .Y(n555) );
  OA21X1_HVT U151 ( .A1(n588), .A2(n294), .A3(n474), .Y(n475) );
  MUX41X1_HVT U153 ( .A1(n516), .A3(n309), .A2(n330), .A4(n355), .S0(n314), 
        .S1(n350), .Y(n472) );
  AND2X1_HVT U154 ( .A1(n321), .A2(n326), .Y(n471) );
  NAND2X0_HVT U158 ( .A1(n335), .A2(n406), .Y(n467) );
  MUX41X1_HVT U159 ( .A1(n614), .A3(n322), .A2(n467), .A4(n361), .S0(n343), 
        .S1(n263), .Y(n466) );
  MUX41X1_HVT U160 ( .A1(n466), .A3(n472), .A2(n468), .A4(n473), .S0(n325), 
        .S1(n345), .Y(n465) );
  AND2X1_HVT U162 ( .A1(n620), .A2(n555), .Y(n463) );
  MUX41X1_HVT U163 ( .A1(n267), .A3(n463), .A2(n310), .A4(n464), .S0(n314), 
        .S1(n348), .Y(n462) );
  MUX41X1_HVT U165 ( .A1(n606), .A3(n373), .A2(n582), .A4(n461), .S0(n262), 
        .S1(n317), .Y(n460) );
  NAND2X0_HVT U166 ( .A1(n333), .A2(n572), .Y(n459) );
  NAND2X0_HVT U167 ( .A1(n407), .A2(n341), .Y(n458) );
  MUX41X1_HVT U168 ( .A1(n392), .A3(n327), .A2(n458), .A4(n459), .S0(n343), 
        .S1(n349), .Y(n457) );
  MUX41X1_HVT U172 ( .A1(n454), .A3(n460), .A2(n457), .A4(n462), .S0(in[0]), 
        .S1(in[5]), .Y(n453) );
  MUX41X1_HVT U176 ( .A1(n324), .A3(n452), .A2(n397), .A4(n613), .S0(n263), 
        .S1(n343), .Y(n451) );
  NAND2X0_HVT U177 ( .A1(n335), .A2(n324), .Y(n450) );
  MUX41X1_HVT U178 ( .A1(n609), .A3(n450), .A2(n401), .A4(n590), .S0(n315), 
        .S1(n263), .Y(n449) );
  MUX41X1_HVT U179 ( .A1(n600), .A3(n402), .A2(n357), .A4(n401), .S0(n342), 
        .S1(n350), .Y(n448) );
  MUX41X1_HVT U180 ( .A1(n360), .A3(n618), .A2(n614), .A4(n305), .S0(n321), 
        .S1(n343), .Y(n447) );
  MUX41X1_HVT U181 ( .A1(n447), .A3(n449), .A2(n448), .A4(n451), .S0(n325), 
        .S1(n345), .Y(n446) );
  MUX41X1_HVT U182 ( .A1(n381), .A3(n245), .A2(n383), .A4(n370), .S0(n350), 
        .S1(n343), .Y(n445) );
  OA21X1_HVT U184 ( .A1(n294), .A2(n594), .A3(n369), .Y(n443) );
  MUX41X1_HVT U186 ( .A1(n308), .A3(n589), .A2(n555), .A4(n582), .S0(n342), 
        .S1(n350), .Y(n441) );
  MUX41X1_HVT U189 ( .A1(n439), .A3(n613), .A2(n440), .A4(n388), .S0(n349), 
        .S1(n316), .Y(n438) );
  MUX41X1_HVT U190 ( .A1(n438), .A3(n441), .A2(n442), .A4(n445), .S0(n346), 
        .S1(in[0]), .Y(n437) );
  MUX41X1_HVT U193 ( .A1(n586), .A3(n593), .A2(n580), .A4(n436), .S0(n342), 
        .S1(n261), .Y(n435) );
  MUX41X1_HVT U195 ( .A1(n620), .A3(n393), .A2(n333), .A4(n591), .S0(n343), 
        .S1(n348), .Y(n433) );
  AO21X1_HVT U197 ( .A1(n307), .A2(n320), .A3(n390), .Y(n431) );
  MUX41X1_HVT U199 ( .A1(n430), .A3(n434), .A2(n433), .A4(n435), .S0(n325), 
        .S1(in[5]), .Y(n429) );
  OA21X1_HVT U201 ( .A1(n619), .A2(n294), .A3(n380), .Y(n427) );
  MUX41X1_HVT U203 ( .A1(n592), .A3(n382), .A2(n615), .A4(n596), .S0(n343), 
        .S1(n261), .Y(n425) );
  MUX41X1_HVT U204 ( .A1(n573), .A3(n614), .A2(n377), .A4(n605), .S0(n318), 
        .S1(n262), .Y(n424) );
  MUX41X1_HVT U205 ( .A1(n270), .A3(n624), .A2(n402), .A4(n375), .S0(n342), 
        .S1(n349), .Y(n423) );
  MUX41X1_HVT U206 ( .A1(n423), .A3(n425), .A2(n424), .A4(n426), .S0(n325), 
        .S1(in[5]), .Y(n422) );
  NAND2X0_HVT U208 ( .A1(n339), .A2(n245), .Y(n515) );
  NAND2X0_HVT U212 ( .A1(n339), .A2(n328), .Y(n572) );
  NAND2X0_HVT U214 ( .A1(n620), .A2(n341), .Y(n421) );
  NAND2X0_HVT U215 ( .A1(n515), .A2(n329), .Y(n420) );
  NAND2X0_HVT U218 ( .A1(n404), .A2(n338), .Y(n474) );
  NAND2X0_HVT U220 ( .A1(n320), .A2(n421), .Y(n547) );
  MUX21X1_HVT U1 ( .A1(n23), .A2(n626), .S0(n336), .Y(n19) );
  INVX8_HVT U2 ( .A(n19), .Y(n616) );
  IBUFFX16_HVT U6 ( .A(n405), .Y(n23) );
  INVX1_HVT U7 ( .A(n231), .Y(n601) );
  MUX21X2_HVT U8 ( .A1(n476), .A2(n475), .S0(n48), .Y(n473) );
  IBUFFX16_HVT U9 ( .A(n318), .Y(n48) );
  INVX0_HVT U10 ( .A(n272), .Y(n603) );
  MUX21X1_HVT U11 ( .A1(n330), .A2(n295), .S0(n273), .Y(n272) );
  MUX21X1_HVT U12 ( .A1(n371), .A2(n598), .S0(n315), .Y(n496) );
  INVX0_HVT U14 ( .A(n598), .Y(n373) );
  MUX41X1_HVT U16 ( .A1(n570), .A3(n313), .A2(n258), .A4(n311), .S0(n50), .S1(
        n319), .Y(n569) );
  IBUFFX16_HVT U17 ( .A(n263), .Y(n50) );
  OA21X2_HVT U18 ( .A1(n379), .A2(n344), .A3(n258), .Y(n517) );
  MUX21X2_HVT U19 ( .A1(n569), .A2(n571), .S0(n210), .Y(n568) );
  IBUFFX16_HVT U20 ( .A(n259), .Y(n210) );
  MUX21X2_HVT U22 ( .A1(n529), .A2(n519), .S0(n211), .Y(out[2]) );
  IBUFFX16_HVT U23 ( .A(in[6]), .Y(n211) );
  NAND2X0_HVT U25 ( .A1(n565), .A2(n212), .Y(n213) );
  NAND2X0_HVT U26 ( .A1(n567), .A2(n298), .Y(n216) );
  NAND2X0_HVT U27 ( .A1(n213), .A2(n216), .Y(n564) );
  IBUFFX2_HVT U28 ( .A(n298), .Y(n212) );
  NAND2X0_HVT U29 ( .A1(n327), .A2(n217), .Y(n218) );
  NAND2X0_HVT U30 ( .A1(n408), .A2(n268), .Y(n219) );
  NAND2X0_HVT U31 ( .A1(n218), .A2(n219), .Y(n267) );
  INVX0_HVT U32 ( .A(n268), .Y(n217) );
  INVX1_HVT U34 ( .A(in[4]), .Y(n408) );
  MUX21X1_HVT U36 ( .A1(n626), .A2(n330), .S0(n232), .Y(n231) );
  IBUFFX16_HVT U37 ( .A(n337), .Y(n232) );
  MUX41X1_HVT U38 ( .A1(n234), .A3(n412), .A2(n231), .A4(n235), .S0(n236), 
        .S1(n348), .Y(n233) );
  IBUFFX16_HVT U39 ( .A(n233), .Y(n489) );
  IBUFFX16_HVT U40 ( .A(n265), .Y(n234) );
  IBUFFX16_HVT U41 ( .A(n621), .Y(n235) );
  IBUFFX16_HVT U43 ( .A(n315), .Y(n236) );
  INVX0_HVT U44 ( .A(n412), .Y(n399) );
  INVX0_HVT U45 ( .A(n315), .Y(n269) );
  INVX1_HVT U46 ( .A(n344), .Y(n342) );
  INVX2_HVT U47 ( .A(in[2]), .Y(n344) );
  AO21X2_HVT U48 ( .A1(n340), .A2(n265), .A3(n294), .Y(n525) );
  INVX1_HVT U49 ( .A(n338), .Y(n256) );
  NBUFFX2_HVT U50 ( .A(n337), .Y(n280) );
  NAND2X0_HVT U52 ( .A1(n374), .A2(n237), .Y(n238) );
  NAND2X0_HVT U54 ( .A1(n491), .A2(n317), .Y(n239) );
  NAND2X0_HVT U55 ( .A1(n238), .A2(n239), .Y(n490) );
  IBUFFX2_HVT U59 ( .A(n317), .Y(n237) );
  INVX1_HVT U60 ( .A(n403), .Y(n240) );
  INVX1_HVT U64 ( .A(n403), .Y(n241) );
  INVX1_HVT U65 ( .A(n240), .Y(n242) );
  INVX1_HVT U67 ( .A(n241), .Y(n243) );
  IBUFFX2_HVT U70 ( .A(n622), .Y(n244) );
  INVX1_HVT U71 ( .A(n244), .Y(n245) );
  INVX1_HVT U72 ( .A(n244), .Y(n246) );
  INVX1_HVT U76 ( .A(n414), .Y(n374) );
  MUX21X1_HVT U78 ( .A1(n398), .A2(n329), .S0(n320), .Y(n491) );
  INVX0_HVT U79 ( .A(n622), .Y(n403) );
  INVX2_HVT U81 ( .A(n340), .Y(n336) );
  IBUFFX2_HVT U87 ( .A(n612), .Y(n365) );
  NAND2X0_HVT U88 ( .A1(n577), .A2(n247), .Y(n248) );
  NAND2X0_HVT U89 ( .A1(n578), .A2(n321), .Y(n249) );
  NAND2X0_HVT U91 ( .A1(n248), .A2(n249), .Y(n575) );
  IBUFFX2_HVT U92 ( .A(n321), .Y(n247) );
  NAND2X0_HVT U94 ( .A1(n579), .A2(n250), .Y(n251) );
  NAND2X0_HVT U95 ( .A1(n575), .A2(n260), .Y(n252) );
  NAND2X0_HVT U99 ( .A1(n251), .A2(n252), .Y(n574) );
  INVX0_HVT U100 ( .A(n260), .Y(n250) );
  NBUFFX4_HVT U102 ( .A(n347), .Y(n321) );
  IBUFFX2_HVT U104 ( .A(n317), .Y(n260) );
  MUX41X1_HVT U107 ( .A1(n558), .A3(n553), .A2(n554), .A4(n551), .S0(n253), 
        .S1(n254), .Y(n550) );
  IBUFFX16_HVT U108 ( .A(n325), .Y(n253) );
  IBUFFX16_HVT U109 ( .A(n319), .Y(n254) );
  INVX1_HVT U111 ( .A(n340), .Y(n335) );
  INVX1_HVT U112 ( .A(in[3]), .Y(n405) );
  NAND2X2_HVT U113 ( .A1(n284), .A2(n285), .Y(out[1]) );
  MUX21X1_HVT U114 ( .A1(n584), .A2(n559), .S0(n316), .Y(n558) );
  XOR2X2_HVT U116 ( .A1(n294), .A2(n601), .Y(n584) );
  OR2X1_HVT U117 ( .A1(n255), .A2(in[3]), .Y(n617) );
  IBUFFX16_HVT U118 ( .A(in[4]), .Y(n255) );
  XNOR2X1_HVT U119 ( .A1(n256), .A2(n404), .Y(n583) );
  MUX41X1_HVT U120 ( .A1(n545), .A3(n541), .A2(n546), .A4(n543), .S0(n257), 
        .S1(in[5]), .Y(n540) );
  IBUFFX16_HVT U121 ( .A(in[0]), .Y(n257) );
  MUX21X1_HVT U122 ( .A1(n327), .A2(n245), .S0(n335), .Y(n258) );
  IBUFFX16_HVT U124 ( .A(n316), .Y(n259) );
  INVX1_HVT U126 ( .A(n327), .Y(n404) );
  INVX0_HVT U127 ( .A(n267), .Y(n609) );
  INVX0_HVT U128 ( .A(n338), .Y(n268) );
  INVX0_HVT U129 ( .A(n335), .Y(n273) );
  INVX1_HVT U130 ( .A(n351), .Y(n261) );
  INVX1_HVT U132 ( .A(n351), .Y(n347) );
  INVX2_HVT U133 ( .A(in[7]), .Y(n351) );
  INVX1_HVT U134 ( .A(n266), .Y(n262) );
  INVX1_HVT U135 ( .A(n266), .Y(n263) );
  INVX1_HVT U137 ( .A(n266), .Y(n348) );
  XNOR2X1_HVT U138 ( .A1(n408), .A2(in[3]), .Y(n295) );
  AO21X1_HVT U143 ( .A1(n318), .A2(n327), .A3(n620), .Y(n507) );
  INVX1_HVT U144 ( .A(in[7]), .Y(n266) );
  INVX2_HVT U145 ( .A(n266), .Y(n350) );
  INVX2_HVT U147 ( .A(n266), .Y(n349) );
  MUX21X1_HVT U148 ( .A1(n406), .A2(n393), .S0(n321), .Y(n559) );
  INVX0_HVT U149 ( .A(n404), .Y(n264) );
  INVX1_HVT U150 ( .A(n264), .Y(n265) );
  OA21X1_HVT U152 ( .A1(n356), .A2(n294), .A3(n597), .Y(n480) );
  OA21X1_HVT U155 ( .A1(n311), .A2(n294), .A3(n597), .Y(n455) );
  MUX21X1_HVT U156 ( .A1(n470), .A2(n469), .S0(n344), .Y(n468) );
  MUX21X2_HVT U157 ( .A1(n376), .A2(n609), .S0(n269), .Y(n493) );
  INVX1_HVT U161 ( .A(n408), .Y(n270) );
  MUX21X2_HVT U164 ( .A1(n453), .A2(n465), .S0(n271), .Y(out[5]) );
  IBUFFX16_HVT U169 ( .A(n299), .Y(n271) );
  MUX41X1_HVT U170 ( .A1(n483), .A3(n479), .A2(n482), .A4(n478), .S0(n274), 
        .S1(n275), .Y(n477) );
  IBUFFX16_HVT U171 ( .A(in[0]), .Y(n274) );
  IBUFFX16_HVT U173 ( .A(n345), .Y(n275) );
  IBUFFX2_HVT U174 ( .A(n588), .Y(n382) );
  MUX21X2_HVT U175 ( .A1(n355), .A2(n377), .S0(n314), .Y(n508) );
  INVX1_HVT U183 ( .A(n594), .Y(n377) );
  NAND2X0_HVT U185 ( .A1(n481), .A2(n276), .Y(n277) );
  NAND2X0_HVT U187 ( .A1(n480), .A2(n317), .Y(n278) );
  NAND2X0_HVT U188 ( .A1(n277), .A2(n278), .Y(n479) );
  IBUFFX2_HVT U191 ( .A(n317), .Y(n276) );
  NBUFFX2_HVT U192 ( .A(n337), .Y(n279) );
  NAND2X0_HVT U194 ( .A1(n502), .A2(n320), .Y(n288) );
  NAND2X0_HVT U196 ( .A1(n427), .A2(n344), .Y(n296) );
  INVX0_HVT U198 ( .A(n346), .Y(n290) );
  INVX1_HVT U200 ( .A(n347), .Y(n294) );
  INVX0_HVT U202 ( .A(in[6]), .Y(n299) );
  NBUFFX2_HVT U207 ( .A(n342), .Y(n314) );
  INVX1_HVT U209 ( .A(n315), .Y(n293) );
  MUX21X2_HVT U210 ( .A1(n506), .A2(n509), .S0(n346), .Y(n505) );
  INVX2_HVT U211 ( .A(n291), .Y(n341) );
  IBUFFX2_HVT U213 ( .A(n340), .Y(n339) );
  NAND2X0_HVT U216 ( .A1(n516), .A2(n298), .Y(n281) );
  NAND2X0_HVT U217 ( .A1(n597), .A2(n293), .Y(n282) );
  NAND2X0_HVT U219 ( .A1(n281), .A2(n282), .Y(n514) );
  MUX21X2_HVT U221 ( .A1(n309), .A2(n528), .S0(n283), .Y(n527) );
  XOR2X1_HVT U222 ( .A1(n318), .A2(n261), .Y(n283) );
  MUX21X1_HVT U223 ( .A1(n332), .A2(n537), .S0(n312), .Y(n536) );
  NAND2X0_HVT U224 ( .A1(n540), .A2(n299), .Y(n284) );
  NAND2X0_HVT U225 ( .A1(n550), .A2(in[6]), .Y(n285) );
  INVX1_HVT U226 ( .A(n596), .Y(n376) );
  MUX21X2_HVT U227 ( .A1(n535), .A2(n536), .S0(n318), .Y(n533) );
  XOR2X1_HVT U228 ( .A1(n295), .A2(n292), .Y(n582) );
  INVX1_HVT U229 ( .A(n295), .Y(n620) );
  MUX21X2_HVT U230 ( .A1(n612), .A2(n375), .S0(n293), .Y(n528) );
  MUX21X2_HVT U231 ( .A1(n507), .A2(n508), .S0(n320), .Y(n506) );
  INVX1_HVT U232 ( .A(n415), .Y(n395) );
  MUX21X2_HVT U233 ( .A1(n590), .A2(n396), .S0(n320), .Y(n469) );
  NAND2X0_HVT U234 ( .A1(n422), .A2(n299), .Y(n286) );
  NAND2X0_HVT U235 ( .A1(n429), .A2(in[6]), .Y(n287) );
  NAND2X0_HVT U236 ( .A1(n286), .A2(n287), .Y(out[7]) );
  NAND2X0_HVT U237 ( .A1(n503), .A2(n294), .Y(n289) );
  NAND2X0_HVT U238 ( .A1(n288), .A2(n289), .Y(n499) );
  MUX21X2_HVT U239 ( .A1(n499), .A2(n498), .S0(n290), .Y(n497) );
  INVX1_HVT U240 ( .A(n417), .Y(n393) );
  INVX2_HVT U241 ( .A(n340), .Y(n337) );
  MUX21X2_HVT U242 ( .A1(n354), .A2(n504), .S0(n315), .Y(n503) );
  MUX41X1_HVT U243 ( .A1(n597), .A3(n272), .A2(n510), .A4(n614), .S0(n293), 
        .S1(n266), .Y(n509) );
  INVX0_HVT U244 ( .A(n292), .Y(n291) );
  INVX0_HVT U245 ( .A(n337), .Y(n292) );
  INVX2_HVT U246 ( .A(in[1]), .Y(n340) );
  OR2X1_HVT U247 ( .A1(n292), .A2(n295), .Y(n613) );
  MUX41X1_HVT U248 ( .A1(n582), .A3(n389), .A2(n555), .A4(n400), .S0(n293), 
        .S1(n294), .Y(n478) );
  INVX0_HVT U249 ( .A(n614), .Y(n386) );
  AND3X2_HVT U250 ( .A1(n317), .A2(n341), .A3(n270), .Y(n495) );
  NAND2X0_HVT U251 ( .A1(n428), .A2(n316), .Y(n297) );
  NAND2X0_HVT U252 ( .A1(n296), .A2(n297), .Y(n426) );
  MUX21X2_HVT U253 ( .A1(n610), .A2(n305), .S0(n320), .Y(n428) );
  INVX1_HVT U254 ( .A(in[0]), .Y(n300) );
  INVX1_HVT U255 ( .A(n344), .Y(n298) );
  MUX21X2_HVT U256 ( .A1(n437), .A2(n446), .S0(in[6]), .Y(out[6]) );
  MUX21X1_HVT U257 ( .A1(n326), .A2(n323), .S0(n340), .Y(n605) );
  MUX21X2_HVT U258 ( .A1(n623), .A2(n487), .S0(n344), .Y(n486) );
  IBUFFX2_HVT U259 ( .A(n340), .Y(n338) );
  MUX21X2_HVT U260 ( .A1(n477), .A2(n485), .S0(in[6]), .Y(out[4]) );
  MUX41X1_HVT U261 ( .A1(n511), .A3(n497), .A2(n505), .A4(n492), .S0(n299), 
        .S1(n300), .Y(out[3]) );
  MUX41X1_HVT U262 ( .A1(n327), .A3(n399), .A2(n601), .A4(n587), .S0(n294), 
        .S1(n344), .Y(n434) );
  MUX41X1_HVT U263 ( .A1(n512), .A3(n514), .A2(n518), .A4(n517), .S0(n350), 
        .S1(n345), .Y(n511) );
  NAND2X0_HVT U264 ( .A1(n332), .A2(n301), .Y(n302) );
  NAND2X0_HVT U265 ( .A1(n513), .A2(n304), .Y(n303) );
  NAND2X0_HVT U266 ( .A1(n302), .A2(n303), .Y(n512) );
  INVX0_HVT U267 ( .A(n304), .Y(n301) );
  INVX0_HVT U268 ( .A(n344), .Y(n343) );
  XNOR2X1_HVT U269 ( .A1(n336), .A2(n343), .Y(n304) );
  NBUFFX2_HVT U270 ( .A(n295), .Y(n322) );
  NBUFFX2_HVT U271 ( .A(n295), .Y(n323) );
  AND2X1_HVT U272 ( .A1(n323), .A2(n572), .Y(n305) );
  MUX21X1_HVT U273 ( .A1(n310), .A2(n366), .S0(n314), .Y(n494) );
  INVX1_HVT U274 ( .A(n330), .Y(n407) );
  MUX21X1_HVT U275 ( .A1(n242), .A2(n406), .S0(n346), .Y(n576) );
  MUX21X1_HVT U276 ( .A1(n363), .A2(n404), .S0(n346), .Y(n561) );
  AND2X1_HVT U277 ( .A1(n331), .A2(n555), .Y(n306) );
  MUX21X1_HVT U278 ( .A1(n322), .A2(n405), .S0(n339), .Y(n610) );
  MUX21X1_HVT U279 ( .A1(n323), .A2(n406), .S0(n338), .Y(n619) );
  MUX21X1_HVT U280 ( .A1(n331), .A2(n322), .S0(n338), .Y(n587) );
  MUX21X1_HVT U281 ( .A1(n245), .A2(n620), .S0(n339), .Y(n591) );
  MUX21X1_HVT U282 ( .A1(n322), .A2(n408), .S0(n280), .Y(n524) );
  MUX21X1_HVT U283 ( .A1(n605), .A2(n381), .S0(n320), .Y(n487) );
  MUX21X1_HVT U284 ( .A1(n620), .A2(n404), .S0(n280), .Y(n412) );
  MUX21X1_HVT U285 ( .A1(n406), .A2(n243), .S0(n336), .Y(n590) );
  MUX21X1_HVT U286 ( .A1(n405), .A2(n407), .S0(n338), .Y(n588) );
  MUX21X1_HVT U287 ( .A1(n243), .A2(n407), .S0(n339), .Y(n452) );
  MUX21X1_HVT U288 ( .A1(n406), .A2(n322), .S0(n280), .Y(n464) );
  MUX21X1_HVT U289 ( .A1(n322), .A2(n243), .S0(n280), .Y(n532) );
  NAND2X0_HVT U290 ( .A1(n408), .A2(n405), .Y(n622) );
  NBUFFX2_HVT U291 ( .A(n625), .Y(n330) );
  MUX21X1_HVT U292 ( .A1(n245), .A2(n329), .S0(n336), .Y(n539) );
  MUX21X1_HVT U293 ( .A1(n405), .A2(n620), .S0(n279), .Y(n415) );
  INVX1_HVT U294 ( .A(n626), .Y(n406) );
  MUX21X1_HVT U295 ( .A1(n406), .A2(n405), .S0(n339), .Y(n594) );
  MUX21X1_HVT U296 ( .A1(n324), .A2(n243), .S0(n336), .Y(n599) );
  NBUFFX2_HVT U297 ( .A(n625), .Y(n331) );
  MUX21X1_HVT U298 ( .A1(n405), .A2(n324), .S0(n279), .Y(n436) );
  XOR2X1_HVT U299 ( .A1(n330), .A2(n339), .Y(n580) );
  MUX21X1_HVT U300 ( .A1(n620), .A2(n324), .S0(n338), .Y(n552) );
  MUX21X1_HVT U301 ( .A1(n242), .A2(n324), .S0(n337), .Y(n413) );
  MUX21X1_HVT U302 ( .A1(n334), .A2(n328), .S0(n338), .Y(n597) );
  MUX21X1_HVT U303 ( .A1(n246), .A2(n405), .S0(n336), .Y(n615) );
  MUX21X1_HVT U304 ( .A1(n324), .A2(n405), .S0(n279), .Y(n504) );
  MUX21X1_HVT U305 ( .A1(n332), .A2(n328), .S0(n336), .Y(n612) );
  MUX21X1_HVT U306 ( .A1(n246), .A2(n334), .S0(n335), .Y(n534) );
  NBUFFX2_HVT U307 ( .A(n625), .Y(n332) );
  MUX21X1_HVT U308 ( .A1(n405), .A2(n334), .S0(n280), .Y(n439) );
  MUX21X1_HVT U309 ( .A1(n333), .A2(n331), .S0(n280), .Y(n440) );
  MUX21X1_HVT U310 ( .A1(n328), .A2(n405), .S0(n279), .Y(n417) );
  MUX21X1_HVT U311 ( .A1(n330), .A2(n324), .S0(n279), .Y(n419) );
  XNOR2X1_HVT U312 ( .A1(n333), .A2(n336), .Y(n307) );
  AND2X1_HVT U313 ( .A1(n335), .A2(n407), .Y(n308) );
  MUX21X1_HVT U314 ( .A1(n330), .A2(n246), .S0(n338), .Y(n411) );
  AND2X1_HVT U315 ( .A1(n333), .A2(n515), .Y(n309) );
  XNOR2X1_HVT U316 ( .A1(n246), .A2(n337), .Y(n310) );
  MUX21X1_HVT U317 ( .A1(n329), .A2(n324), .S0(n336), .Y(n557) );
  MUX21X1_HVT U318 ( .A1(n329), .A2(n334), .S0(n317), .Y(n501) );
  XOR2X1_HVT U319 ( .A1(n324), .A2(n338), .Y(n602) );
  NBUFFX2_HVT U320 ( .A(n347), .Y(n320) );
  NBUFFX2_HVT U321 ( .A(n342), .Y(n316) );
  NBUFFX2_HVT U322 ( .A(n342), .Y(n315) );
  NBUFFX2_HVT U323 ( .A(n342), .Y(n318) );
  NBUFFX2_HVT U324 ( .A(n345), .Y(n319) );
  NBUFFX2_HVT U325 ( .A(n342), .Y(n317) );
  MUX21X1_HVT U326 ( .A1(n526), .A2(n374), .S0(n317), .Y(n523) );
  MUX21X1_HVT U327 ( .A1(n443), .A2(n444), .S0(n316), .Y(n442) );
  MUX21X1_HVT U328 ( .A1(n542), .A2(n326), .S0(n320), .Y(n444) );
  XOR2X1_HVT U329 ( .A1(n335), .A2(in[3]), .Y(n581) );
  MUX21X1_HVT U330 ( .A1(n328), .A2(n323), .S0(n339), .Y(n521) );
  NAND2X0_HVT U331 ( .A1(n326), .A2(n408), .Y(n625) );
  MUX21X1_HVT U332 ( .A1(n395), .A2(n404), .S0(n320), .Y(n476) );
  MUX21X1_HVT U333 ( .A1(n549), .A2(n548), .S0(n318), .Y(n546) );
  MUX21X1_HVT U334 ( .A1(n607), .A2(n329), .S0(n321), .Y(n549) );
  MUX21X1_HVT U335 ( .A1(n456), .A2(n455), .S0(n317), .Y(n454) );
  MUX21X1_HVT U336 ( .A1(n329), .A2(n393), .S0(n321), .Y(n456) );
  AND2X1_HVT U337 ( .A1(n323), .A2(n341), .Y(n311) );
  NBUFFX2_HVT U338 ( .A(n617), .Y(n327) );
  MUX21X1_HVT U339 ( .A1(n326), .A2(n242), .S0(n338), .Y(n589) );
  MUX21X1_HVT U340 ( .A1(n599), .A2(n358), .S0(n321), .Y(n481) );
  MUX21X1_HVT U341 ( .A1(n404), .A2(n407), .S0(n280), .Y(n461) );
  MUX21X1_HVT U342 ( .A1(n407), .A2(n326), .S0(n339), .Y(n608) );
  MUX21X1_HVT U343 ( .A1(n378), .A2(n624), .S0(n315), .Y(n518) );
  MUX21X1_HVT U344 ( .A1(n471), .A2(n332), .S0(n312), .Y(n470) );
  MUX21X1_HVT U345 ( .A1(n326), .A2(n593), .S0(n346), .Y(n578) );
  XOR2X1_HVT U346 ( .A1(n335), .A2(n345), .Y(n585) );
  NBUFFX2_HVT U347 ( .A(n617), .Y(n328) );
  MUX21X1_HVT U348 ( .A1(n384), .A2(n401), .S0(n320), .Y(n432) );
  MUX21X1_HVT U349 ( .A1(n624), .A2(n340), .S0(n316), .Y(n500) );
  MUX21X1_HVT U350 ( .A1(n326), .A2(n404), .S0(n280), .Y(n416) );
  MUX21X1_HVT U351 ( .A1(n364), .A2(n341), .S0(n346), .Y(n563) );
  NBUFFX2_HVT U352 ( .A(n626), .Y(n333) );
  MUX21X1_HVT U353 ( .A1(n598), .A2(n420), .S0(n321), .Y(n414) );
  MUX21X1_HVT U354 ( .A1(n245), .A2(n326), .S0(n335), .Y(n618) );
  MUX21X1_HVT U355 ( .A1(n326), .A2(n324), .S0(n321), .Y(n537) );
  NBUFFX2_HVT U356 ( .A(n617), .Y(n329) );
  NBUFFX2_HVT U357 ( .A(n626), .Y(n334) );
  NBUFFX2_HVT U358 ( .A(n408), .Y(n324) );
  XNOR2X1_HVT U359 ( .A1(n294), .A2(n337), .Y(n312) );
  AND2X1_HVT U360 ( .A1(n405), .A2(n341), .Y(n313) );
  NBUFFX2_HVT U361 ( .A(in[5]), .Y(n346) );
  NBUFFX2_HVT U362 ( .A(in[5]), .Y(n345) );
  MUX21X1_HVT U363 ( .A1(n432), .A2(n431), .S0(n316), .Y(n430) );
  MUX21X1_HVT U364 ( .A1(n242), .A2(n270), .S0(n336), .Y(n596) );
  MUX21X1_HVT U365 ( .A1(n270), .A2(n406), .S0(n336), .Y(n592) );
  NAND2X0_HVT U366 ( .A1(in[3]), .A2(in[4]), .Y(n626) );
  MUX21X1_HVT U367 ( .A1(n270), .A2(n620), .S0(n279), .Y(n418) );
  MUX21X1_HVT U368 ( .A1(n270), .A2(n332), .S0(n337), .Y(n607) );
  MUX21X1_HVT U369 ( .A1(n270), .A2(n328), .S0(n279), .Y(n410) );
  MUX21X1_HVT U370 ( .A1(n270), .A2(n333), .S0(n338), .Y(n409) );
  MUX21X1_HVT U371 ( .A1(n326), .A2(n270), .S0(n314), .Y(n513) );
  MUX21X1_HVT U372 ( .A1(n334), .A2(n270), .S0(n339), .Y(n600) );
  MUX21X1_HVT U373 ( .A1(n405), .A2(n270), .S0(n335), .Y(n598) );
  NBUFFX2_HVT U374 ( .A(in[3]), .Y(n326) );
  NBUFFX2_HVT U375 ( .A(in[0]), .Y(n325) );
  INVX0_HVT U376 ( .A(n606), .Y(n352) );
  INVX0_HVT U377 ( .A(n604), .Y(n353) );
  INVX0_HVT U378 ( .A(n595), .Y(n354) );
  INVX0_HVT U379 ( .A(n593), .Y(n355) );
  INVX0_HVT U380 ( .A(n458), .Y(n356) );
  INVX0_HVT U381 ( .A(n421), .Y(n357) );
  INVX0_HVT U382 ( .A(n624), .Y(n358) );
  INVX0_HVT U383 ( .A(n611), .Y(n359) );
  INVX0_HVT U384 ( .A(n623), .Y(n360) );
  INVX0_HVT U385 ( .A(n621), .Y(n361) );
  INVX0_HVT U386 ( .A(n619), .Y(n362) );
  INVX0_HVT U387 ( .A(n618), .Y(n363) );
  INVX0_HVT U388 ( .A(n615), .Y(n364) );
  INVX0_HVT U389 ( .A(n610), .Y(n366) );
  INVX0_HVT U390 ( .A(n608), .Y(n367) );
  INVX0_HVT U391 ( .A(n607), .Y(n368) );
  INVX0_HVT U392 ( .A(n605), .Y(n369) );
  INVX0_HVT U393 ( .A(n602), .Y(n370) );
  INVX0_HVT U394 ( .A(n600), .Y(n371) );
  INVX0_HVT U395 ( .A(n599), .Y(n372) );
  INVX0_HVT U396 ( .A(n597), .Y(n375) );
  INVX0_HVT U397 ( .A(n592), .Y(n378) );
  INVX0_HVT U398 ( .A(n591), .Y(n379) );
  INVX0_HVT U399 ( .A(n590), .Y(n380) );
  INVX0_HVT U400 ( .A(n589), .Y(n381) );
  INVX0_HVT U401 ( .A(n587), .Y(n383) );
  INVX0_HVT U402 ( .A(n586), .Y(n384) );
  INVX0_HVT U403 ( .A(n555), .Y(n385) );
  INVX0_HVT U404 ( .A(n515), .Y(n387) );
  INVX0_HVT U405 ( .A(n420), .Y(n388) );
  INVX0_HVT U406 ( .A(n572), .Y(n389) );
  INVX0_HVT U407 ( .A(n474), .Y(n390) );
  INVX0_HVT U408 ( .A(n419), .Y(n391) );
  INVX0_HVT U409 ( .A(n418), .Y(n392) );
  INVX0_HVT U410 ( .A(n416), .Y(n394) );
  INVX0_HVT U411 ( .A(n534), .Y(n396) );
  INVX0_HVT U412 ( .A(n524), .Y(n397) );
  INVX0_HVT U413 ( .A(n413), .Y(n398) );
  INVX0_HVT U414 ( .A(n411), .Y(n400) );
  INVX0_HVT U415 ( .A(n410), .Y(n401) );
  INVX0_HVT U416 ( .A(n409), .Y(n402) );
endmodule

