
module Mix_Column ( in, out );
  input [127:0] in;
  output [127:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203;

  XNOR3X1_HVT U1 ( .A1(n1), .A2(n2), .A3(n3), .Y(out[9]) );
  XOR2X1_HVT U2 ( .A1(n4), .A2(in[1]), .Y(n3) );
  XOR2X1_HVT U3 ( .A1(n5), .A2(n6), .Y(out[99]) );
  XNOR3X1_HVT U4 ( .A1(in[122]), .A2(in[103]), .A3(n7), .Y(n6) );
  XNOR3X1_HVT U5 ( .A1(in[98]), .A2(in[127]), .A3(in[123]), .Y(n5) );
  XNOR3X1_HVT U6 ( .A1(n8), .A2(in[106]), .A3(n9), .Y(out[98]) );
  INVX0_HVT U7 ( .A(n10), .Y(n8) );
  XNOR3X1_HVT U8 ( .A1(n11), .A2(n12), .A3(n13), .Y(out[97]) );
  XOR2X1_HVT U9 ( .A1(n14), .A2(in[121]), .Y(n13) );
  XNOR3X1_HVT U10 ( .A1(n15), .A2(in[103]), .A3(n11), .Y(out[96]) );
  XOR2X1_HVT U11 ( .A1(in[112]), .A2(in[104]), .Y(n15) );
  XNOR3X1_HVT U12 ( .A1(n16), .A2(in[87]), .A3(n17), .Y(out[95]) );
  XNOR3X1_HVT U13 ( .A1(n18), .A2(in[86]), .A3(n19), .Y(out[94]) );
  XNOR3X1_HVT U14 ( .A1(n20), .A2(in[85]), .A3(n21), .Y(out[93]) );
  XNOR3X1_HVT U15 ( .A1(n22), .A2(n23), .A3(n24), .Y(out[92]) );
  XNOR3X1_HVT U16 ( .A1(in[95]), .A2(in[84]), .A3(in[83]), .Y(n24) );
  XNOR3X1_HVT U17 ( .A1(n25), .A2(n26), .A3(n27), .Y(out[91]) );
  XNOR3X1_HVT U18 ( .A1(in[95]), .A2(in[90]), .A3(in[82]), .Y(n27) );
  XOR3X1_HVT U19 ( .A1(n28), .A2(in[82]), .A3(n29), .Y(out[90]) );
  XNOR3X1_HVT U20 ( .A1(n30), .A2(n31), .A3(n1), .Y(out[8]) );
  XOR2X1_HVT U21 ( .A1(in[24]), .A2(in[16]), .Y(n30) );
  XOR3X1_HVT U22 ( .A1(n32), .A2(n33), .A3(n34), .Y(out[89]) );
  XOR2X1_HVT U23 ( .A1(n35), .A2(in[81]), .Y(n34) );
  XOR3X1_HVT U24 ( .A1(n36), .A2(in[64]), .A3(n32), .Y(out[88]) );
  XOR2X1_HVT U25 ( .A1(in[95]), .A2(in[72]), .Y(n36) );
  XNOR3X1_HVT U26 ( .A1(n37), .A2(in[78]), .A3(n38), .Y(out[87]) );
  XOR2X1_HVT U27 ( .A1(in[95]), .A2(in[86]), .Y(n37) );
  XOR3X1_HVT U28 ( .A1(n39), .A2(in[77]), .A3(n18), .Y(out[86]) );
  XOR2X1_HVT U29 ( .A1(in[94]), .A2(in[85]), .Y(n39) );
  XNOR3X1_HVT U30 ( .A1(n40), .A2(in[93]), .A3(n20), .Y(out[85]) );
  XNOR3X1_HVT U31 ( .A1(n26), .A2(n41), .A3(n42), .Y(out[84]) );
  XNOR3X1_HVT U32 ( .A1(in[79]), .A2(in[76]), .A3(in[75]), .Y(n42) );
  XNOR2X1_HVT U33 ( .A1(in[83]), .A2(n43), .Y(n26) );
  INVX0_HVT U34 ( .A(in[87]), .Y(n43) );
  XNOR3X1_HVT U35 ( .A1(n23), .A2(n25), .A3(n44), .Y(out[83]) );
  XNOR3X1_HVT U36 ( .A1(in[82]), .A2(in[79]), .A3(in[74]), .Y(n44) );
  XOR2X1_HVT U37 ( .A1(in[67]), .A2(in[75]), .Y(n25) );
  XOR2X1_HVT U38 ( .A1(in[91]), .A2(in[87]), .Y(n23) );
  XNOR3X1_HVT U39 ( .A1(n45), .A2(in[90]), .A3(n28), .Y(out[82]) );
  XNOR2X1_HVT U40 ( .A1(in[66]), .A2(in[74]), .Y(n28) );
  XNOR3X1_HVT U41 ( .A1(n46), .A2(n47), .A3(n48), .Y(out[81]) );
  XOR2X1_HVT U42 ( .A1(n32), .A2(n49), .Y(n48) );
  XOR2X1_HVT U43 ( .A1(in[80]), .A2(in[87]), .Y(n32) );
  XNOR3X1_HVT U44 ( .A1(n50), .A2(in[64]), .A3(n47), .Y(out[80]) );
  XOR2X1_HVT U45 ( .A1(in[88]), .A2(in[87]), .Y(n50) );
  XNOR3X1_HVT U46 ( .A1(n51), .A2(n31), .A3(n52), .Y(out[7]) );
  XOR2X1_HVT U47 ( .A1(in[6]), .A2(in[30]), .Y(n51) );
  XNOR3X1_HVT U48 ( .A1(n53), .A2(in[71]), .A3(n18), .Y(out[79]) );
  XOR2X1_HVT U49 ( .A1(in[70]), .A2(in[78]), .Y(n18) );
  XOR3X1_HVT U50 ( .A1(n20), .A2(in[70]), .A3(n17), .Y(out[78]) );
  XNOR2X1_HVT U51 ( .A1(in[69]), .A2(in[77]), .Y(n20) );
  XNOR3X1_HVT U52 ( .A1(n22), .A2(in[69]), .A3(n19), .Y(out[77]) );
  XOR2X1_HVT U53 ( .A1(in[68]), .A2(in[76]), .Y(n22) );
  XNOR3X1_HVT U54 ( .A1(n16), .A2(n21), .A3(n54), .Y(out[76]) );
  XNOR3X1_HVT U55 ( .A1(in[75]), .A2(in[68]), .A3(in[67]), .Y(n54) );
  XOR2X1_HVT U56 ( .A1(in[84]), .A2(in[92]), .Y(n21) );
  INVX0_HVT U57 ( .A(n38), .Y(n16) );
  XNOR2X1_HVT U58 ( .A1(in[71]), .A2(in[79]), .Y(n38) );
  XOR2X1_HVT U59 ( .A1(n55), .A2(n56), .Y(out[75]) );
  XNOR3X1_HVT U60 ( .A1(in[74]), .A2(in[67]), .A3(n57), .Y(n56) );
  XNOR3X1_HVT U61 ( .A1(in[91]), .A2(in[83]), .A3(in[79]), .Y(n55) );
  XNOR3X1_HVT U62 ( .A1(n58), .A2(in[66]), .A3(n33), .Y(out[74]) );
  XOR2X1_HVT U63 ( .A1(in[65]), .A2(n49), .Y(n33) );
  INVX0_HVT U64 ( .A(in[73]), .Y(n49) );
  XNOR3X1_HVT U65 ( .A1(n47), .A2(n59), .A3(n60), .Y(out[73]) );
  XOR2X1_HVT U66 ( .A1(n29), .A2(in[65]), .Y(n60) );
  XNOR2X1_HVT U67 ( .A1(in[81]), .A2(in[89]), .Y(n29) );
  XOR2X1_HVT U68 ( .A1(n61), .A2(in[79]), .Y(n47) );
  INVX0_HVT U69 ( .A(in[72]), .Y(n61) );
  XNOR3X1_HVT U70 ( .A1(n62), .A2(in[79]), .A3(n59), .Y(out[72]) );
  XOR2X1_HVT U71 ( .A1(in[88]), .A2(in[80]), .Y(n62) );
  XNOR3X1_HVT U72 ( .A1(n63), .A2(in[70]), .A3(n53), .Y(out[71]) );
  XNOR2X1_HVT U73 ( .A1(in[87]), .A2(in[95]), .Y(n53) );
  XOR2X1_HVT U74 ( .A1(in[94]), .A2(in[79]), .Y(n63) );
  XNOR3X1_HVT U75 ( .A1(n64), .A2(in[69]), .A3(n17), .Y(out[70]) );
  XNOR2X1_HVT U76 ( .A1(in[86]), .A2(in[94]), .Y(n17) );
  XOR2X1_HVT U77 ( .A1(in[93]), .A2(in[78]), .Y(n64) );
  XNOR3X1_HVT U78 ( .A1(n65), .A2(in[14]), .A3(n66), .Y(out[6]) );
  XOR2X1_HVT U79 ( .A1(in[5]), .A2(in[29]), .Y(n65) );
  XNOR3X1_HVT U80 ( .A1(n41), .A2(in[77]), .A3(n19), .Y(out[69]) );
  XNOR2X1_HVT U81 ( .A1(in[85]), .A2(in[93]), .Y(n19) );
  XOR2X1_HVT U82 ( .A1(in[68]), .A2(in[92]), .Y(n41) );
  XNOR3X1_HVT U83 ( .A1(n40), .A2(n67), .A3(n68), .Y(out[68]) );
  XNOR3X1_HVT U84 ( .A1(in[92]), .A2(in[71]), .A3(in[67]), .Y(n68) );
  XOR2X1_HVT U85 ( .A1(in[76]), .A2(in[84]), .Y(n40) );
  XNOR3X1_HVT U86 ( .A1(n57), .A2(n67), .A3(n69), .Y(out[67]) );
  XNOR3X1_HVT U87 ( .A1(in[90]), .A2(in[83]), .A3(in[75]), .Y(n69) );
  XOR2X1_HVT U88 ( .A1(in[91]), .A2(in[95]), .Y(n67) );
  XOR2X1_HVT U89 ( .A1(in[66]), .A2(in[71]), .Y(n57) );
  XNOR3X1_HVT U90 ( .A1(n58), .A2(in[74]), .A3(n46), .Y(out[66]) );
  XNOR2X1_HVT U91 ( .A1(in[65]), .A2(in[89]), .Y(n46) );
  XOR2X1_HVT U92 ( .A1(in[82]), .A2(in[90]), .Y(n58) );
  XOR3X1_HVT U93 ( .A1(n45), .A2(n59), .A3(n70), .Y(out[65]) );
  XOR2X1_HVT U94 ( .A1(n35), .A2(in[89]), .Y(n70) );
  XNOR2X1_HVT U95 ( .A1(in[64]), .A2(in[71]), .Y(n59) );
  XOR2X1_HVT U96 ( .A1(in[73]), .A2(in[81]), .Y(n45) );
  XNOR3X1_HVT U97 ( .A1(n71), .A2(in[71]), .A3(n35), .Y(out[64]) );
  XNOR2X1_HVT U98 ( .A1(in[88]), .A2(in[95]), .Y(n35) );
  XOR2X1_HVT U99 ( .A1(in[80]), .A2(in[72]), .Y(n71) );
  XNOR3X1_HVT U100 ( .A1(n72), .A2(in[55]), .A3(n73), .Y(out[63]) );
  XNOR3X1_HVT U101 ( .A1(n74), .A2(in[54]), .A3(n75), .Y(out[62]) );
  XNOR3X1_HVT U102 ( .A1(n76), .A2(in[53]), .A3(n77), .Y(out[61]) );
  XNOR3X1_HVT U103 ( .A1(n78), .A2(n79), .A3(n80), .Y(out[60]) );
  XNOR3X1_HVT U104 ( .A1(in[63]), .A2(in[52]), .A3(in[51]), .Y(n80) );
  XNOR3X1_HVT U105 ( .A1(n81), .A2(in[13]), .A3(n82), .Y(out[5]) );
  XNOR3X1_HVT U106 ( .A1(n83), .A2(n84), .A3(n85), .Y(out[59]) );
  XNOR3X1_HVT U107 ( .A1(in[63]), .A2(in[58]), .A3(in[50]), .Y(n85) );
  XOR3X1_HVT U108 ( .A1(n86), .A2(in[50]), .A3(n87), .Y(out[58]) );
  XOR3X1_HVT U109 ( .A1(n88), .A2(n89), .A3(n90), .Y(out[57]) );
  XOR2X1_HVT U110 ( .A1(n91), .A2(in[49]), .Y(n90) );
  XOR3X1_HVT U111 ( .A1(n92), .A2(in[32]), .A3(n88), .Y(out[56]) );
  XOR2X1_HVT U112 ( .A1(in[63]), .A2(in[40]), .Y(n92) );
  XNOR3X1_HVT U113 ( .A1(n93), .A2(in[46]), .A3(n94), .Y(out[55]) );
  XOR2X1_HVT U114 ( .A1(in[63]), .A2(in[54]), .Y(n93) );
  XOR3X1_HVT U115 ( .A1(n95), .A2(in[45]), .A3(n74), .Y(out[54]) );
  XOR2X1_HVT U116 ( .A1(in[62]), .A2(in[53]), .Y(n95) );
  XNOR3X1_HVT U117 ( .A1(n96), .A2(in[61]), .A3(n76), .Y(out[53]) );
  XNOR3X1_HVT U118 ( .A1(n84), .A2(n97), .A3(n98), .Y(out[52]) );
  XNOR3X1_HVT U119 ( .A1(in[47]), .A2(in[44]), .A3(in[43]), .Y(n98) );
  XNOR2X1_HVT U120 ( .A1(in[51]), .A2(n99), .Y(n84) );
  INVX0_HVT U121 ( .A(in[55]), .Y(n99) );
  XNOR3X1_HVT U122 ( .A1(n79), .A2(n83), .A3(n100), .Y(out[51]) );
  XNOR3X1_HVT U123 ( .A1(in[50]), .A2(in[47]), .A3(in[42]), .Y(n100) );
  XOR2X1_HVT U124 ( .A1(in[35]), .A2(in[43]), .Y(n83) );
  XOR2X1_HVT U125 ( .A1(in[59]), .A2(in[55]), .Y(n79) );
  XNOR3X1_HVT U126 ( .A1(n101), .A2(in[58]), .A3(n86), .Y(out[50]) );
  XNOR2X1_HVT U127 ( .A1(in[34]), .A2(in[42]), .Y(n86) );
  XNOR3X1_HVT U128 ( .A1(n102), .A2(n103), .A3(n104), .Y(out[4]) );
  XNOR3X1_HVT U129 ( .A1(in[3]), .A2(in[28]), .A3(in[27]), .Y(n104) );
  XNOR3X1_HVT U130 ( .A1(n105), .A2(n106), .A3(n107), .Y(out[49]) );
  XOR2X1_HVT U131 ( .A1(n88), .A2(n108), .Y(n107) );
  XOR2X1_HVT U132 ( .A1(in[48]), .A2(in[55]), .Y(n88) );
  XNOR3X1_HVT U133 ( .A1(n109), .A2(in[32]), .A3(n106), .Y(out[48]) );
  XOR2X1_HVT U134 ( .A1(in[56]), .A2(in[55]), .Y(n109) );
  XNOR3X1_HVT U135 ( .A1(n110), .A2(in[39]), .A3(n74), .Y(out[47]) );
  XOR2X1_HVT U136 ( .A1(in[38]), .A2(in[46]), .Y(n74) );
  XOR3X1_HVT U137 ( .A1(n76), .A2(in[38]), .A3(n73), .Y(out[46]) );
  XNOR2X1_HVT U138 ( .A1(in[37]), .A2(in[45]), .Y(n76) );
  XNOR3X1_HVT U139 ( .A1(n78), .A2(in[37]), .A3(n75), .Y(out[45]) );
  XOR2X1_HVT U140 ( .A1(in[36]), .A2(in[44]), .Y(n78) );
  XNOR3X1_HVT U141 ( .A1(n72), .A2(n77), .A3(n111), .Y(out[44]) );
  XNOR3X1_HVT U142 ( .A1(in[43]), .A2(in[36]), .A3(in[35]), .Y(n111) );
  XOR2X1_HVT U143 ( .A1(in[52]), .A2(in[60]), .Y(n77) );
  INVX0_HVT U144 ( .A(n94), .Y(n72) );
  XNOR2X1_HVT U145 ( .A1(in[39]), .A2(in[47]), .Y(n94) );
  XOR2X1_HVT U146 ( .A1(n112), .A2(n113), .Y(out[43]) );
  XNOR3X1_HVT U147 ( .A1(in[42]), .A2(in[35]), .A3(n114), .Y(n113) );
  XNOR3X1_HVT U148 ( .A1(in[59]), .A2(in[51]), .A3(in[47]), .Y(n112) );
  XNOR3X1_HVT U149 ( .A1(n115), .A2(in[34]), .A3(n89), .Y(out[42]) );
  XOR2X1_HVT U150 ( .A1(in[33]), .A2(n108), .Y(n89) );
  INVX0_HVT U151 ( .A(in[41]), .Y(n108) );
  XNOR3X1_HVT U152 ( .A1(n106), .A2(n116), .A3(n117), .Y(out[41]) );
  XOR2X1_HVT U153 ( .A1(n87), .A2(in[33]), .Y(n117) );
  XNOR2X1_HVT U154 ( .A1(in[49]), .A2(in[57]), .Y(n87) );
  XOR2X1_HVT U155 ( .A1(n118), .A2(in[47]), .Y(n106) );
  INVX0_HVT U156 ( .A(in[40]), .Y(n118) );
  XNOR3X1_HVT U157 ( .A1(n119), .A2(in[47]), .A3(n116), .Y(out[40]) );
  XOR2X1_HVT U158 ( .A1(in[56]), .A2(in[48]), .Y(n119) );
  XNOR3X1_HVT U159 ( .A1(n120), .A2(n121), .A3(n122), .Y(out[3]) );
  XOR2X1_HVT U160 ( .A1(n103), .A2(in[26]), .Y(n122) );
  XOR2X1_HVT U161 ( .A1(n123), .A2(in[7]), .Y(n103) );
  XNOR3X1_HVT U162 ( .A1(n124), .A2(in[38]), .A3(n110), .Y(out[39]) );
  XNOR2X1_HVT U163 ( .A1(in[55]), .A2(in[63]), .Y(n110) );
  XOR2X1_HVT U164 ( .A1(in[62]), .A2(in[47]), .Y(n124) );
  XNOR3X1_HVT U165 ( .A1(n125), .A2(in[37]), .A3(n73), .Y(out[38]) );
  XNOR2X1_HVT U166 ( .A1(in[54]), .A2(in[62]), .Y(n73) );
  XOR2X1_HVT U167 ( .A1(in[61]), .A2(in[46]), .Y(n125) );
  XNOR3X1_HVT U168 ( .A1(n97), .A2(in[45]), .A3(n75), .Y(out[37]) );
  XNOR2X1_HVT U169 ( .A1(in[53]), .A2(in[61]), .Y(n75) );
  XOR2X1_HVT U170 ( .A1(in[36]), .A2(in[60]), .Y(n97) );
  XNOR3X1_HVT U171 ( .A1(n96), .A2(n126), .A3(n127), .Y(out[36]) );
  XNOR3X1_HVT U172 ( .A1(in[60]), .A2(in[39]), .A3(in[35]), .Y(n127) );
  XOR2X1_HVT U173 ( .A1(in[44]), .A2(in[52]), .Y(n96) );
  XNOR3X1_HVT U174 ( .A1(n114), .A2(n126), .A3(n128), .Y(out[35]) );
  XNOR3X1_HVT U175 ( .A1(in[58]), .A2(in[51]), .A3(in[43]), .Y(n128) );
  XOR2X1_HVT U176 ( .A1(in[59]), .A2(in[63]), .Y(n126) );
  XOR2X1_HVT U177 ( .A1(in[34]), .A2(in[39]), .Y(n114) );
  XNOR3X1_HVT U178 ( .A1(n115), .A2(in[42]), .A3(n105), .Y(out[34]) );
  XNOR2X1_HVT U179 ( .A1(in[33]), .A2(in[57]), .Y(n105) );
  XOR2X1_HVT U180 ( .A1(in[50]), .A2(in[58]), .Y(n115) );
  XOR3X1_HVT U181 ( .A1(n101), .A2(n116), .A3(n129), .Y(out[33]) );
  XOR2X1_HVT U182 ( .A1(n91), .A2(in[57]), .Y(n129) );
  XNOR2X1_HVT U183 ( .A1(in[32]), .A2(in[39]), .Y(n116) );
  XOR2X1_HVT U184 ( .A1(in[41]), .A2(in[49]), .Y(n101) );
  XNOR3X1_HVT U185 ( .A1(n130), .A2(in[39]), .A3(n91), .Y(out[32]) );
  XNOR2X1_HVT U186 ( .A1(in[56]), .A2(in[63]), .Y(n91) );
  XOR2X1_HVT U187 ( .A1(in[48]), .A2(in[40]), .Y(n130) );
  XNOR3X1_HVT U188 ( .A1(n131), .A2(in[23]), .A3(n66), .Y(out[31]) );
  XNOR3X1_HVT U189 ( .A1(n132), .A2(in[22]), .A3(n82), .Y(out[30]) );
  XNOR3X1_HVT U190 ( .A1(n133), .A2(in[10]), .A3(n134), .Y(out[2]) );
  XOR3X1_HVT U191 ( .A1(n135), .A2(in[21]), .A3(n136), .Y(out[29]) );
  XNOR3X1_HVT U192 ( .A1(n52), .A2(n137), .A3(n138), .Y(out[28]) );
  XNOR3X1_HVT U193 ( .A1(in[27]), .A2(in[20]), .A3(in[19]), .Y(n138) );
  XOR2X1_HVT U194 ( .A1(n139), .A2(n140), .Y(out[27]) );
  XNOR3X1_HVT U195 ( .A1(in[23]), .A2(in[18]), .A3(n120), .Y(n140) );
  XOR2X1_HVT U196 ( .A1(in[11]), .A2(in[19]), .Y(n120) );
  XNOR3X1_HVT U197 ( .A1(in[3]), .A2(in[31]), .A3(in[26]), .Y(n139) );
  XNOR3X1_HVT U198 ( .A1(n141), .A2(in[18]), .A3(n2), .Y(out[26]) );
  XOR2X1_HVT U199 ( .A1(in[17]), .A2(in[25]), .Y(n2) );
  XNOR3X1_HVT U200 ( .A1(n142), .A2(n143), .A3(n144), .Y(out[25]) );
  XNOR2X1_HVT U201 ( .A1(n145), .A2(in[17]), .Y(n144) );
  XOR3X1_HVT U202 ( .A1(n146), .A2(in[0]), .A3(n142), .Y(out[24]) );
  XOR2X1_HVT U203 ( .A1(in[8]), .A2(in[31]), .Y(n146) );
  XOR3X1_HVT U204 ( .A1(n147), .A2(in[14]), .A3(n131), .Y(out[23]) );
  XNOR2X1_HVT U205 ( .A1(n31), .A2(in[7]), .Y(n131) );
  XOR2X1_HVT U206 ( .A1(in[31]), .A2(in[22]), .Y(n147) );
  XOR3X1_HVT U207 ( .A1(n148), .A2(in[13]), .A3(n132), .Y(out[22]) );
  XOR2X1_HVT U208 ( .A1(in[30]), .A2(in[21]), .Y(n148) );
  XNOR3X1_HVT U209 ( .A1(n136), .A2(in[29]), .A3(n102), .Y(out[21]) );
  XNOR2X1_HVT U210 ( .A1(in[12]), .A2(in[20]), .Y(n102) );
  XOR2X1_HVT U211 ( .A1(n149), .A2(n150), .Y(out[20]) );
  XNOR3X1_HVT U212 ( .A1(in[12]), .A2(in[11]), .A3(n81), .Y(n150) );
  XOR2X1_HVT U213 ( .A1(in[28]), .A2(in[4]), .Y(n81) );
  XNOR3X1_HVT U214 ( .A1(in[23]), .A2(in[19]), .A3(in[15]), .Y(n149) );
  XNOR3X1_HVT U215 ( .A1(n145), .A2(n151), .A3(n152), .Y(out[1]) );
  XNOR2X1_HVT U216 ( .A1(n1), .A2(in[25]), .Y(n152) );
  XOR2X1_HVT U217 ( .A1(in[0]), .A2(in[7]), .Y(n1) );
  XOR2X1_HVT U218 ( .A1(n153), .A2(n154), .Y(out[19]) );
  XNOR3X1_HVT U219 ( .A1(in[18]), .A2(in[11]), .A3(n155), .Y(n154) );
  XNOR3X1_HVT U220 ( .A1(in[3]), .A2(in[27]), .A3(in[23]), .Y(n153) );
  XNOR3X1_HVT U221 ( .A1(n151), .A2(in[26]), .A3(n141), .Y(out[18]) );
  XNOR2X1_HVT U222 ( .A1(in[10]), .A2(in[2]), .Y(n141) );
  XOR2X1_HVT U223 ( .A1(in[17]), .A2(in[9]), .Y(n151) );
  XNOR3X1_HVT U224 ( .A1(n133), .A2(n142), .A3(n156), .Y(out[17]) );
  XOR2X1_HVT U225 ( .A1(n4), .A2(in[9]), .Y(n156) );
  XOR2X1_HVT U226 ( .A1(in[16]), .A2(in[23]), .Y(n142) );
  XOR2X1_HVT U227 ( .A1(in[1]), .A2(in[25]), .Y(n133) );
  XNOR3X1_HVT U228 ( .A1(n157), .A2(in[0]), .A3(n4), .Y(out[16]) );
  XOR2X1_HVT U229 ( .A1(in[8]), .A2(n31), .Y(n4) );
  XOR2X1_HVT U230 ( .A1(in[24]), .A2(in[23]), .Y(n157) );
  XOR3X1_HVT U231 ( .A1(n132), .A2(in[7]), .A3(n52), .Y(out[15]) );
  XOR2X1_HVT U232 ( .A1(in[23]), .A2(in[31]), .Y(n52) );
  XOR2X1_HVT U233 ( .A1(in[14]), .A2(in[6]), .Y(n132) );
  XNOR3X1_HVT U234 ( .A1(n136), .A2(in[6]), .A3(n66), .Y(out[14]) );
  XNOR2X1_HVT U235 ( .A1(in[22]), .A2(in[30]), .Y(n66) );
  XOR2X1_HVT U236 ( .A1(in[13]), .A2(in[5]), .Y(n136) );
  XNOR3X1_HVT U237 ( .A1(n137), .A2(in[5]), .A3(n82), .Y(out[13]) );
  XNOR2X1_HVT U238 ( .A1(in[21]), .A2(in[29]), .Y(n82) );
  XOR2X1_HVT U239 ( .A1(in[12]), .A2(in[4]), .Y(n137) );
  XNOR3X1_HVT U240 ( .A1(n135), .A2(n158), .A3(n159), .Y(out[12]) );
  XNOR3X1_HVT U241 ( .A1(in[4]), .A2(in[15]), .A3(in[11]), .Y(n159) );
  XOR2X1_HVT U242 ( .A1(in[20]), .A2(in[28]), .Y(n135) );
  XNOR3X1_HVT U243 ( .A1(n160), .A2(n161), .A3(n162), .Y(out[127]) );
  XOR3X1_HVT U244 ( .A1(n163), .A2(in[118]), .A3(n164), .Y(out[126]) );
  XNOR3X1_HVT U245 ( .A1(n165), .A2(in[117]), .A3(n166), .Y(out[125]) );
  XOR3X1_HVT U246 ( .A1(n167), .A2(n168), .A3(n169), .Y(out[124]) );
  XNOR3X1_HVT U247 ( .A1(in[123]), .A2(in[116]), .A3(in[115]), .Y(n169) );
  XNOR3X1_HVT U248 ( .A1(n7), .A2(n170), .A3(n171), .Y(out[123]) );
  XNOR3X1_HVT U249 ( .A1(in[122]), .A2(in[119]), .A3(in[114]), .Y(n171) );
  XOR2X1_HVT U250 ( .A1(in[107]), .A2(in[115]), .Y(n7) );
  XOR3X1_HVT U251 ( .A1(n172), .A2(in[114]), .A3(n173), .Y(out[122]) );
  XNOR3X1_HVT U252 ( .A1(n174), .A2(n175), .A3(n176), .Y(out[121]) );
  XOR2X1_HVT U253 ( .A1(n11), .A2(in[113]), .Y(n176) );
  XNOR2X1_HVT U254 ( .A1(in[120]), .A2(in[127]), .Y(n11) );
  XOR3X1_HVT U255 ( .A1(n177), .A2(in[104]), .A3(n175), .Y(out[120]) );
  XOR2X1_HVT U256 ( .A1(in[96]), .A2(in[127]), .Y(n177) );
  XNOR3X1_HVT U257 ( .A1(n155), .A2(n158), .A3(n178), .Y(out[11]) );
  XNOR2X1_HVT U258 ( .A1(n121), .A2(in[19]), .Y(n178) );
  XOR2X1_HVT U259 ( .A1(in[2]), .A2(in[27]), .Y(n121) );
  XOR2X1_HVT U260 ( .A1(in[3]), .A2(in[7]), .Y(n158) );
  XNOR2X1_HVT U261 ( .A1(in[10]), .A2(n31), .Y(n155) );
  INVX0_HVT U262 ( .A(in[15]), .Y(n31) );
  XNOR3X1_HVT U263 ( .A1(n179), .A2(in[110]), .A3(n160), .Y(out[119]) );
  XOR2X1_HVT U264 ( .A1(in[127]), .A2(in[118]), .Y(n179) );
  XNOR3X1_HVT U265 ( .A1(n180), .A2(in[109]), .A3(n164), .Y(out[118]) );
  XOR2X1_HVT U266 ( .A1(in[126]), .A2(in[117]), .Y(n180) );
  XNOR3X1_HVT U267 ( .A1(n181), .A2(in[125]), .A3(n165), .Y(out[117]) );
  XOR2X1_HVT U268 ( .A1(n182), .A2(n183), .Y(out[116]) );
  XNOR3X1_HVT U269 ( .A1(in[108]), .A2(in[107]), .A3(n184), .Y(n183) );
  XNOR3X1_HVT U270 ( .A1(in[119]), .A2(in[115]), .A3(in[111]), .Y(n182) );
  XOR2X1_HVT U271 ( .A1(n185), .A2(n186), .Y(out[115]) );
  XNOR3X1_HVT U272 ( .A1(in[114]), .A2(in[106]), .A3(n187), .Y(n186) );
  XNOR3X1_HVT U273 ( .A1(in[99]), .A2(in[123]), .A3(in[119]), .Y(n185) );
  XNOR3X1_HVT U274 ( .A1(n173), .A2(in[122]), .A3(n12), .Y(out[114]) );
  XNOR2X1_HVT U275 ( .A1(in[105]), .A2(in[113]), .Y(n12) );
  XNOR2X1_HVT U276 ( .A1(n188), .A2(in[98]), .Y(n173) );
  XNOR3X1_HVT U277 ( .A1(n175), .A2(n189), .A3(n190), .Y(out[113]) );
  XOR2X1_HVT U278 ( .A1(n10), .A2(in[105]), .Y(n190) );
  XNOR2X1_HVT U279 ( .A1(in[121]), .A2(in[97]), .Y(n10) );
  XOR2X1_HVT U280 ( .A1(n191), .A2(n161), .Y(n175) );
  INVX0_HVT U281 ( .A(in[112]), .Y(n191) );
  XNOR3X1_HVT U282 ( .A1(n192), .A2(n161), .A3(n189), .Y(out[112]) );
  XOR2X1_HVT U283 ( .A1(in[96]), .A2(in[120]), .Y(n192) );
  XNOR3X1_HVT U284 ( .A1(n168), .A2(n193), .A3(n164), .Y(out[111]) );
  XNOR2X1_HVT U285 ( .A1(in[102]), .A2(in[110]), .Y(n164) );
  XOR3X1_HVT U286 ( .A1(n165), .A2(in[102]), .A3(n162), .Y(out[110]) );
  XNOR2X1_HVT U287 ( .A1(in[101]), .A2(in[109]), .Y(n165) );
  XNOR3X1_HVT U288 ( .A1(n143), .A2(in[2]), .A3(n134), .Y(out[10]) );
  XNOR2X1_HVT U289 ( .A1(in[18]), .A2(in[26]), .Y(n134) );
  XOR2X1_HVT U290 ( .A1(in[1]), .A2(in[9]), .Y(n143) );
  XNOR3X1_HVT U291 ( .A1(n167), .A2(in[101]), .A3(n163), .Y(out[109]) );
  XOR2X1_HVT U292 ( .A1(in[100]), .A2(in[108]), .Y(n167) );
  XNOR3X1_HVT U293 ( .A1(n166), .A2(n187), .A3(n194), .Y(out[108]) );
  XNOR3X1_HVT U294 ( .A1(in[99]), .A2(in[103]), .A3(in[100]), .Y(n194) );
  XOR2X1_HVT U295 ( .A1(in[107]), .A2(in[111]), .Y(n187) );
  XOR2X1_HVT U296 ( .A1(in[116]), .A2(in[124]), .Y(n166) );
  XOR2X1_HVT U297 ( .A1(n195), .A2(n196), .Y(out[107]) );
  XNOR3X1_HVT U298 ( .A1(in[115]), .A2(n188), .A3(n160), .Y(n196) );
  XNOR2X1_HVT U299 ( .A1(in[103]), .A2(in[111]), .Y(n160) );
  INVX0_HVT U300 ( .A(in[106]), .Y(n188) );
  XNOR3X1_HVT U301 ( .A1(in[99]), .A2(in[98]), .A3(in[123]), .Y(n195) );
  XNOR3X1_HVT U302 ( .A1(n174), .A2(in[98]), .A3(n9), .Y(out[106]) );
  XNOR2X1_HVT U303 ( .A1(in[114]), .A2(in[122]), .Y(n9) );
  XOR2X1_HVT U304 ( .A1(in[105]), .A2(in[97]), .Y(n174) );
  XNOR3X1_HVT U305 ( .A1(n172), .A2(n189), .A3(n197), .Y(out[105]) );
  XOR2X1_HVT U306 ( .A1(n14), .A2(in[97]), .Y(n197) );
  XOR2X1_HVT U307 ( .A1(in[104]), .A2(in[111]), .Y(n189) );
  XOR2X1_HVT U308 ( .A1(in[113]), .A2(in[121]), .Y(n172) );
  XNOR3X1_HVT U309 ( .A1(n198), .A2(in[111]), .A3(n14), .Y(out[104]) );
  XOR2X1_HVT U310 ( .A1(in[96]), .A2(n193), .Y(n14) );
  INVX0_HVT U311 ( .A(in[103]), .Y(n193) );
  XOR2X1_HVT U312 ( .A1(in[120]), .A2(in[112]), .Y(n198) );
  XNOR3X1_HVT U313 ( .A1(n199), .A2(in[102]), .A3(n168), .Y(out[103]) );
  XOR2X1_HVT U314 ( .A1(n161), .A2(in[127]), .Y(n168) );
  INVX0_HVT U315 ( .A(in[119]), .Y(n161) );
  XOR2X1_HVT U316 ( .A1(in[126]), .A2(in[111]), .Y(n199) );
  XNOR3X1_HVT U317 ( .A1(n200), .A2(in[101]), .A3(n162), .Y(out[102]) );
  XNOR2X1_HVT U318 ( .A1(in[118]), .A2(in[126]), .Y(n162) );
  XOR2X1_HVT U319 ( .A1(in[125]), .A2(in[110]), .Y(n200) );
  XNOR3X1_HVT U320 ( .A1(n184), .A2(in[109]), .A3(n163), .Y(out[101]) );
  XNOR2X1_HVT U321 ( .A1(in[117]), .A2(in[125]), .Y(n163) );
  XOR2X1_HVT U322 ( .A1(in[100]), .A2(in[124]), .Y(n184) );
  XNOR3X1_HVT U323 ( .A1(n170), .A2(n181), .A3(n201), .Y(out[100]) );
  XNOR3X1_HVT U324 ( .A1(in[124]), .A2(in[123]), .A3(in[103]), .Y(n201) );
  XOR2X1_HVT U325 ( .A1(in[108]), .A2(in[116]), .Y(n181) );
  XOR2X1_HVT U326 ( .A1(in[99]), .A2(in[127]), .Y(n170) );
  XOR3X1_HVT U327 ( .A1(n202), .A2(in[16]), .A3(n145), .Y(out[0]) );
  XOR2X1_HVT U328 ( .A1(n203), .A2(n123), .Y(n145) );
  INVX0_HVT U329 ( .A(in[31]), .Y(n123) );
  INVX0_HVT U330 ( .A(in[24]), .Y(n203) );
  XOR2X1_HVT U331 ( .A1(in[8]), .A2(in[7]), .Y(n202) );
endmodule

