
module sbox_13 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n50, n121, n210, n211, n212, n213, n216, n217, n218, n219,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575;

  NAND2X0_HVT U3 ( .A1(n284), .A2(n277), .Y(n573) );
  NAND2X0_HVT U4 ( .A1(n275), .A2(n573), .Y(n572) );
  NAND2X0_HVT U5 ( .A1(n282), .A2(n267), .Y(n570) );
  NAND2X0_HVT U13 ( .A1(n562), .A2(n279), .Y(n563) );
  NAND2X0_HVT U15 ( .A1(n573), .A2(n356), .Y(n560) );
  NAND2X0_HVT U21 ( .A1(n274), .A2(n286), .Y(n554) );
  NAND2X0_HVT U24 ( .A1(n271), .A2(n286), .Y(n552) );
  NAND2X0_HVT U33 ( .A1(n351), .A2(n286), .Y(n543) );
  NAND2X0_HVT U35 ( .A1(n269), .A2(n286), .Y(n541) );
  NAND2X0_HVT U42 ( .A1(n280), .A2(n271), .Y(n534) );
  MUX41X1_HVT U51 ( .A1(n339), .A3(n299), .A2(n317), .A4(n318), .S0(n296), 
        .S1(n291), .Y(n527) );
  NAND2X0_HVT U53 ( .A1(n524), .A2(n533), .Y(n525) );
  NAND2X0_HVT U56 ( .A1(n275), .A2(n520), .Y(n521) );
  MUX41X1_HVT U57 ( .A1(n340), .A3(n556), .A2(n521), .A4(n565), .S0(n296), 
        .S1(n291), .Y(n519) );
  NAND2X0_HVT U58 ( .A1(n279), .A2(n573), .Y(n518) );
  MUX41X1_HVT U59 ( .A1(n256), .A3(n518), .A2(n254), .A4(n316), .S0(n296), 
        .S1(n291), .Y(n517) );
  MUX41X1_HVT U61 ( .A1(n253), .A3(n315), .A2(n314), .A4(n268), .S0(n296), 
        .S1(in[5]), .Y(n515) );
  NAND2X0_HVT U62 ( .A1(n286), .A2(n278), .Y(n514) );
  MUX41X1_HVT U63 ( .A1(n514), .A3(n306), .A2(n241), .A4(n313), .S0(n296), 
        .S1(n291), .Y(n513) );
  AO21X1_HVT U66 ( .A1(n311), .A2(n263), .A3(n334), .Y(n510) );
  MUX41X1_HVT U68 ( .A1(n309), .A3(n510), .A2(n509), .A4(n511), .S0(n257), 
        .S1(n235), .Y(n508) );
  MUX41X1_HVT U69 ( .A1(n508), .A3(n516), .A2(n512), .A4(n522), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n272), .A2(n503), .Y(n504) );
  MUX41X1_HVT U74 ( .A1(n505), .A3(n550), .A2(n504), .A4(n552), .S0(n259), 
        .S1(n293), .Y(n502) );
  MUX41X1_HVT U75 ( .A1(n337), .A3(n342), .A2(n355), .A4(n320), .S0(n257), 
        .S1(n235), .Y(n501) );
  MUX41X1_HVT U77 ( .A1(n567), .A3(n344), .A2(n500), .A4(n343), .S0(n264), 
        .S1(n289), .Y(n499) );
  MUX41X1_HVT U78 ( .A1(n499), .A3(n502), .A2(n501), .A4(n506), .S0(in[0]), 
        .S1(n292), .Y(n498) );
  AND3X1_HVT U80 ( .A1(n277), .A2(n520), .A3(n495), .Y(n496) );
  AND2X1_HVT U83 ( .A1(n281), .A2(n219), .Y(n492) );
  MUX41X1_HVT U84 ( .A1(n319), .A3(n237), .A2(n559), .A4(n492), .S0(n257), 
        .S1(n235), .Y(n491) );
  NAND2X0_HVT U85 ( .A1(n286), .A2(n354), .Y(n490) );
  MUX41X1_HVT U86 ( .A1(n342), .A3(n490), .A2(n251), .A4(n249), .S0(n257), 
        .S1(n294), .Y(n489) );
  MUX41X1_HVT U87 ( .A1(n489), .A3(n493), .A2(n491), .A4(n494), .S0(in[0]), 
        .S1(n291), .Y(n488) );
  MUX41X1_HVT U90 ( .A1(n530), .A3(n534), .A2(n339), .A4(n487), .S0(n258), 
        .S1(n235), .Y(n486) );
  AO21X1_HVT U93 ( .A1(n266), .A2(n482), .A3(n338), .Y(n483) );
  MUX41X1_HVT U96 ( .A1(n300), .A3(n252), .A2(n341), .A4(n480), .S0(n257), 
        .S1(n294), .Y(n479) );
  MUX41X1_HVT U97 ( .A1(n337), .A3(n252), .A2(n280), .A4(n560), .S0(n257), 
        .S1(n293), .Y(n478) );
  MUX41X1_HVT U98 ( .A1(n478), .A3(n481), .A2(n479), .A4(n486), .S0(n270), 
        .S1(n292), .Y(n477) );
  NAND2X0_HVT U101 ( .A1(n473), .A2(n472), .Y(n474) );
  MUX41X1_HVT U103 ( .A1(n573), .A3(n310), .A2(n323), .A4(n541), .S0(n257), 
        .S1(n293), .Y(n470) );
  MUX21X2_HVT U107 ( .A1(n467), .A2(n477), .S0(in[6]), .Y(out[2]) );
  NAND2X0_HVT U110 ( .A1(n277), .A2(n463), .Y(n464) );
  AO21X1_HVT U118 ( .A1(n260), .A2(n566), .A3(n237), .Y(n456) );
  NAND2X0_HVT U123 ( .A1(n450), .A2(n449), .Y(n451) );
  MUX41X1_HVT U131 ( .A1(n442), .A3(n444), .A2(n443), .A4(n445), .S0(n263), 
        .S1(n296), .Y(n441) );
  MUX41X1_HVT U132 ( .A1(n441), .A3(n454), .A2(n446), .A4(n459), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  MUX41X1_HVT U135 ( .A1(n347), .A3(n352), .A2(n570), .A4(n549), .S0(n259), 
        .S1(n295), .Y(n438) );
  MUX41X1_HVT U136 ( .A1(n249), .A3(n543), .A2(n348), .A4(n540), .S0(n258), 
        .S1(n296), .Y(n437) );
  MUX41X1_HVT U139 ( .A1(n435), .A3(n438), .A2(n437), .A4(n439), .S0(n270), 
        .S1(n291), .Y(n434) );
  AND2X1_HVT U140 ( .A1(n566), .A2(n285), .Y(n433) );
  MUX41X1_HVT U141 ( .A1(n551), .A3(n329), .A2(n433), .A4(n326), .S0(n259), 
        .S1(n295), .Y(n432) );
  MUX41X1_HVT U142 ( .A1(n319), .A3(n268), .A2(n335), .A4(n566), .S0(n258), 
        .S1(n295), .Y(n431) );
  NAND2X0_HVT U146 ( .A1(n284), .A2(n279), .Y(n503) );
  MUX41X1_HVT U147 ( .A1(n348), .A3(n503), .A2(n337), .A4(n530), .S0(n259), 
        .S1(n296), .Y(n427) );
  MUX41X1_HVT U148 ( .A1(n427), .A3(n431), .A2(n428), .A4(n432), .S0(n270), 
        .S1(n291), .Y(n426) );
  OA21X1_HVT U151 ( .A1(n536), .A2(n297), .A3(n423), .Y(n424) );
  MUX41X1_HVT U153 ( .A1(n464), .A3(n253), .A2(n276), .A4(n302), .S0(n258), 
        .S1(n235), .Y(n421) );
  AND2X1_HVT U154 ( .A1(n266), .A2(n271), .Y(n420) );
  NAND2X0_HVT U158 ( .A1(n283), .A2(n354), .Y(n416) );
  MUX41X1_HVT U159 ( .A1(n563), .A3(n268), .A2(n416), .A4(n308), .S0(n289), 
        .S1(n294), .Y(n415) );
  MUX41X1_HVT U160 ( .A1(n415), .A3(n421), .A2(n417), .A4(n422), .S0(n270), 
        .S1(n262), .Y(n414) );
  AND2X1_HVT U162 ( .A1(n237), .A2(n503), .Y(n412) );
  MUX41X1_HVT U163 ( .A1(n315), .A3(n412), .A2(n250), .A4(n413), .S0(n289), 
        .S1(n293), .Y(n411) );
  MUX41X1_HVT U165 ( .A1(n554), .A3(n324), .A2(n530), .A4(n410), .S0(n296), 
        .S1(n289), .Y(n409) );
  NAND2X0_HVT U166 ( .A1(n279), .A2(n520), .Y(n408) );
  NAND2X0_HVT U167 ( .A1(n355), .A2(n286), .Y(n407) );
  MUX41X1_HVT U168 ( .A1(n340), .A3(n566), .A2(n407), .A4(n408), .S0(n289), 
        .S1(n294), .Y(n406) );
  MUX41X1_HVT U172 ( .A1(n403), .A3(n409), .A2(n406), .A4(n411), .S0(in[0]), 
        .S1(n262), .Y(n402) );
  MUX21X2_HVT U173 ( .A1(n402), .A2(n414), .S0(in[6]), .Y(out[5]) );
  NAND2X0_HVT U174 ( .A1(n280), .A2(n569), .Y(n562) );
  MUX41X1_HVT U176 ( .A1(n269), .A3(n401), .A2(n345), .A4(n562), .S0(n296), 
        .S1(n288), .Y(n400) );
  NAND2X0_HVT U177 ( .A1(n50), .A2(n269), .Y(n399) );
  MUX41X1_HVT U178 ( .A1(n558), .A3(n399), .A2(n349), .A4(n538), .S0(n259), 
        .S1(n294), .Y(n398) );
  MUX41X1_HVT U179 ( .A1(n548), .A3(n350), .A2(n304), .A4(n349), .S0(n288), 
        .S1(n235), .Y(n397) );
  MUX41X1_HVT U180 ( .A1(n307), .A3(n567), .A2(n563), .A4(n248), .S0(n264), 
        .S1(n288), .Y(n396) );
  MUX41X1_HVT U181 ( .A1(n396), .A3(n398), .A2(n397), .A4(n400), .S0(n270), 
        .S1(n262), .Y(n395) );
  MUX41X1_HVT U182 ( .A1(n330), .A3(n273), .A2(n332), .A4(n321), .S0(n296), 
        .S1(n288), .Y(n394) );
  OA21X1_HVT U184 ( .A1(n542), .A2(n297), .A3(n319), .Y(n392) );
  MUX41X1_HVT U186 ( .A1(n252), .A3(n537), .A2(n503), .A4(n530), .S0(n288), 
        .S1(n293), .Y(n390) );
  MUX41X1_HVT U189 ( .A1(n388), .A3(n562), .A2(n389), .A4(n336), .S0(n264), 
        .S1(n288), .Y(n387) );
  MUX41X1_HVT U190 ( .A1(n387), .A3(n390), .A2(n391), .A4(n394), .S0(n262), 
        .S1(in[0]), .Y(n386) );
  MUX41X1_HVT U194 ( .A1(n535), .A3(n549), .A2(n347), .A4(n566), .S0(n264), 
        .S1(n289), .Y(n383) );
  MUX41X1_HVT U195 ( .A1(n237), .A3(n341), .A2(n575), .A4(n539), .S0(n288), 
        .S1(n235), .Y(n382) );
  AO21X1_HVT U197 ( .A1(n251), .A2(n265), .A3(n338), .Y(n380) );
  MUX41X1_HVT U199 ( .A1(n379), .A3(n383), .A2(n382), .A4(n384), .S0(in[0]), 
        .S1(n262), .Y(n378) );
  OA21X1_HVT U201 ( .A1(n568), .A2(n297), .A3(n329), .Y(n376) );
  MUX41X1_HVT U203 ( .A1(n540), .A3(n331), .A2(n564), .A4(n544), .S0(n288), 
        .S1(n294), .Y(n374) );
  MUX41X1_HVT U204 ( .A1(n521), .A3(n563), .A2(n327), .A4(n553), .S0(n288), 
        .S1(n293), .Y(n373) );
  MUX41X1_HVT U205 ( .A1(n219), .A3(n573), .A2(n350), .A4(n242), .S0(n289), 
        .S1(n294), .Y(n372) );
  NAND2X0_HVT U208 ( .A1(n121), .A2(n274), .Y(n463) );
  NAND2X0_HVT U212 ( .A1(n50), .A2(n272), .Y(n520) );
  NAND2X0_HVT U214 ( .A1(n237), .A2(n286), .Y(n370) );
  NAND2X0_HVT U215 ( .A1(n463), .A2(n272), .Y(n369) );
  AO21X1_HVT U216 ( .A1(n285), .A2(n352), .A3(n297), .Y(n473) );
  NAND2X0_HVT U218 ( .A1(n352), .A2(n121), .Y(n423) );
  NAND2X0_HVT U220 ( .A1(n265), .A2(n370), .Y(n495) );
  IBUFFX16_HVT U1 ( .A(n297), .Y(n294) );
  INVX2_HVT U2 ( .A(in[7]), .Y(n297) );
  MUX21X1_HVT U6 ( .A1(n559), .A2(n248), .S0(n264), .Y(n377) );
  NAND2X2_HVT U7 ( .A1(in[4]), .A2(n353), .Y(n566) );
  MUX41X1_HVT U8 ( .A1(n336), .A3(n469), .A2(n529), .A4(n322), .S0(n23), .S1(
        n231), .Y(n468) );
  IBUFFX16_HVT U9 ( .A(n257), .Y(n23) );
  INVX1_HVT U10 ( .A(n297), .Y(n235) );
  INVX2_HVT U11 ( .A(n266), .Y(n231) );
  MUX41X1_HVT U12 ( .A1(n561), .A3(n300), .A2(n318), .A4(n531), .S0(n48), .S1(
        n231), .Y(n493) );
  IBUFFX16_HVT U14 ( .A(n257), .Y(n48) );
  IBUFFX2_HVT U16 ( .A(n285), .Y(n50) );
  IBUFFX2_HVT U17 ( .A(n285), .Y(n121) );
  MUX21X1_HVT U18 ( .A1(n507), .A2(n532), .S0(n243), .Y(n506) );
  MUX21X2_HVT U19 ( .A1(n498), .A2(n488), .S0(n239), .Y(out[1]) );
  INVX1_HVT U20 ( .A(n285), .Y(n284) );
  IBUFFX2_HVT U22 ( .A(n285), .Y(n280) );
  OA21X2_HVT U23 ( .A1(n303), .A2(n297), .A3(n545), .Y(n429) );
  OA21X2_HVT U25 ( .A1(n254), .A2(n297), .A3(n545), .Y(n404) );
  MUX21X2_HVT U26 ( .A1(n354), .A2(n341), .S0(n266), .Y(n507) );
  IBUFFX2_HVT U27 ( .A(n285), .Y(n281) );
  MUX21X2_HVT U28 ( .A1(n419), .A2(n418), .S0(n210), .Y(n417) );
  IBUFFX16_HVT U29 ( .A(n261), .Y(n210) );
  NAND2X0_HVT U30 ( .A1(n464), .A2(n211), .Y(n212) );
  NAND2X0_HVT U31 ( .A1(n545), .A2(n243), .Y(n213) );
  NAND2X0_HVT U32 ( .A1(n212), .A2(n213), .Y(n462) );
  IBUFFX2_HVT U34 ( .A(n243), .Y(n211) );
  IBUFFX2_HVT U36 ( .A(n285), .Y(n282) );
  INVX1_HVT U37 ( .A(n276), .Y(n355) );
  INVX1_HVT U38 ( .A(n357), .Y(n219) );
  INVX1_HVT U39 ( .A(n273), .Y(n351) );
  MUX21X1_HVT U40 ( .A1(n234), .A2(n236), .S0(n121), .Y(n233) );
  INVX0_HVT U41 ( .A(n275), .Y(n234) );
  INVX0_HVT U43 ( .A(n233), .Y(n539) );
  MUX21X1_HVT U44 ( .A1(n377), .A2(n376), .S0(n243), .Y(n375) );
  INVX0_HVT U45 ( .A(in[6]), .Y(n239) );
  INVX1_HVT U46 ( .A(n569), .Y(n356) );
  INVX1_HVT U47 ( .A(in[3]), .Y(n353) );
  INVX0_HVT U48 ( .A(n258), .Y(n243) );
  NAND2X0_HVT U49 ( .A1(n378), .A2(n216), .Y(n217) );
  NAND2X0_HVT U50 ( .A1(n371), .A2(n239), .Y(n218) );
  NAND2X0_HVT U52 ( .A1(n217), .A2(n218), .Y(out[7]) );
  INVX0_HVT U54 ( .A(n239), .Y(n216) );
  INVX1_HVT U55 ( .A(n359), .Y(n349) );
  MUX21X2_HVT U60 ( .A1(n381), .A2(n380), .S0(n260), .Y(n379) );
  MUX21X2_HVT U64 ( .A1(n333), .A2(n349), .S0(n265), .Y(n381) );
  INVX1_HVT U65 ( .A(n361), .Y(n347) );
  MUX21X1_HVT U67 ( .A1(n354), .A2(n355), .S0(n232), .Y(n549) );
  INVX0_HVT U70 ( .A(n284), .Y(n232) );
  INVX1_HVT U71 ( .A(in[4]), .Y(n357) );
  INVX0_HVT U72 ( .A(n569), .Y(n236) );
  MUX21X2_HVT U76 ( .A1(n424), .A2(n425), .S0(n257), .Y(n422) );
  MUX41X1_HVT U79 ( .A1(n385), .A3(n528), .A2(n541), .A4(n534), .S0(n290), 
        .S1(n231), .Y(n384) );
  INVX1_HVT U81 ( .A(n545), .Y(n242) );
  INVX0_HVT U82 ( .A(n240), .Y(n458) );
  MUX21X2_HVT U88 ( .A1(n302), .A2(n327), .S0(n258), .Y(n457) );
  MUX21X2_HVT U89 ( .A1(n451), .A2(n452), .S0(n231), .Y(n448) );
  XOR2X1_HVT U91 ( .A1(n297), .A2(n549), .Y(n532) );
  MUX41X1_HVT U92 ( .A1(n554), .A3(n256), .A2(n309), .A4(n346), .S0(n258), 
        .S1(n295), .Y(n447) );
  INVX1_HVT U94 ( .A(n362), .Y(n346) );
  MUX21X2_HVT U95 ( .A1(n305), .A2(n547), .S0(n231), .Y(n430) );
  MUX21X2_HVT U99 ( .A1(n455), .A2(n458), .S0(n263), .Y(n454) );
  IBUFFX2_HVT U100 ( .A(n538), .Y(n329) );
  MUX21X2_HVT U102 ( .A1(n538), .A2(n344), .S0(n264), .Y(n418) );
  MUX21X2_HVT U104 ( .A1(n456), .A2(n457), .S0(n265), .Y(n455) );
  MUX21X2_HVT U105 ( .A1(n301), .A2(n453), .S0(n259), .Y(n452) );
  INVX1_HVT U106 ( .A(n542), .Y(n327) );
  MUX41X1_HVT U108 ( .A1(n462), .A3(n465), .A2(n460), .A4(n466), .S0(n263), 
        .S1(n297), .Y(n459) );
  IBUFFX2_HVT U109 ( .A(n297), .Y(n293) );
  MUX21X2_HVT U111 ( .A1(n447), .A2(n448), .S0(n263), .Y(n446) );
  INVX2_HVT U112 ( .A(in[1]), .Y(n285) );
  AND3X2_HVT U113 ( .A1(n261), .A2(n286), .A3(n219), .Y(n444) );
  INVX1_HVT U114 ( .A(in[2]), .Y(n290) );
  INVX1_HVT U115 ( .A(in[7]), .Y(n298) );
  INVX2_HVT U116 ( .A(n298), .Y(n295) );
  OA21X1_HVT U117 ( .A1(n233), .A2(n290), .A3(n316), .Y(n465) );
  MUX21X1_HVT U119 ( .A1(n278), .A2(n461), .S0(n247), .Y(n460) );
  INVX1_HVT U120 ( .A(n236), .Y(n237) );
  INVX0_HVT U121 ( .A(n563), .Y(n241) );
  INVX1_HVT U122 ( .A(n291), .Y(n245) );
  INVX1_HVT U124 ( .A(n270), .Y(n238) );
  MUX41X1_HVT U125 ( .A1(n375), .A3(n373), .A2(n374), .A4(n372), .S0(n238), 
        .S1(n245), .Y(n371) );
  MUX21X1_HVT U126 ( .A1(n267), .A2(n356), .S0(n285), .Y(n559) );
  IBUFFX2_HVT U127 ( .A(n285), .Y(n283) );
  XOR2X2_HVT U128 ( .A1(n357), .A2(in[3]), .Y(n569) );
  MUX41X1_HVT U129 ( .A1(n242), .A3(n551), .A2(n244), .A4(n241), .S0(n243), 
        .S1(n298), .Y(n240) );
  NAND2X0_HVT U130 ( .A1(n284), .A2(n268), .Y(n244) );
  MUX41X1_HVT U133 ( .A1(n475), .A3(n470), .A2(n471), .A4(n468), .S0(n238), 
        .S1(n245), .Y(n467) );
  MUX21X2_HVT U134 ( .A1(n426), .A2(n434), .S0(in[6]), .Y(out[4]) );
  INVX1_HVT U137 ( .A(n290), .Y(n287) );
  IBUFFX2_HVT U138 ( .A(n290), .Y(n288) );
  MUX21X2_HVT U143 ( .A1(n476), .A2(n253), .S0(n246), .Y(n475) );
  XNOR2X1_HVT U144 ( .A1(n286), .A2(n290), .Y(n247) );
  IBUFFX2_HVT U145 ( .A(in[1]), .Y(n286) );
  IBUFFX2_HVT U149 ( .A(n290), .Y(n289) );
  NBUFFX4_HVT U150 ( .A(n287), .Y(n258) );
  INVX0_HVT U152 ( .A(n298), .Y(n296) );
  MUX21X2_HVT U155 ( .A1(n386), .A2(n395), .S0(in[6]), .Y(out[6]) );
  XNOR2X1_HVT U156 ( .A1(n289), .A2(n295), .Y(n246) );
  MUX21X1_HVT U157 ( .A1(n250), .A2(n314), .S0(n258), .Y(n443) );
  NBUFFX2_HVT U161 ( .A(n356), .Y(n268) );
  AND2X1_HVT U164 ( .A1(n356), .A2(n520), .Y(n248) );
  NBUFFX2_HVT U169 ( .A(n571), .Y(n273) );
  MUX21X1_HVT U170 ( .A1(n351), .A2(n354), .S0(n263), .Y(n524) );
  NBUFFX2_HVT U171 ( .A(n571), .Y(n274) );
  NBUFFX2_HVT U175 ( .A(n571), .Y(n275) );
  MUX21X1_HVT U183 ( .A1(n310), .A2(n352), .S0(n263), .Y(n509) );
  AND2X1_HVT U185 ( .A1(n277), .A2(n503), .Y(n249) );
  MUX21X1_HVT U187 ( .A1(n356), .A2(n354), .S0(n283), .Y(n568) );
  MUX21X1_HVT U188 ( .A1(n277), .A2(n268), .S0(n283), .Y(n535) );
  MUX21X1_HVT U191 ( .A1(n268), .A2(n269), .S0(n283), .Y(n472) );
  MUX21X1_HVT U192 ( .A1(n436), .A2(n572), .S0(n260), .Y(n435) );
  MUX21X1_HVT U193 ( .A1(n553), .A2(n330), .S0(n265), .Y(n436) );
  MUX21X1_HVT U196 ( .A1(n351), .A2(n355), .S0(n282), .Y(n401) );
  MUX21X1_HVT U198 ( .A1(n354), .A2(n356), .S0(n121), .Y(n413) );
  MUX21X1_HVT U200 ( .A1(n356), .A2(n351), .S0(n50), .Y(n480) );
  MUX21X1_HVT U202 ( .A1(n237), .A2(n352), .S0(n121), .Y(n361) );
  MUX21X1_HVT U206 ( .A1(n569), .A2(n355), .S0(n283), .Y(n551) );
  MUX21X1_HVT U207 ( .A1(n237), .A2(n269), .S0(n282), .Y(n500) );
  XOR2X1_HVT U209 ( .A1(n569), .A2(n121), .Y(n530) );
  MUX21X1_HVT U210 ( .A1(n267), .A2(n237), .S0(n283), .Y(n364) );
  MUX21X1_HVT U211 ( .A1(n354), .A2(n351), .S0(n50), .Y(n538) );
  MUX21X1_HVT U213 ( .A1(n267), .A2(n355), .S0(n282), .Y(n536) );
  MUX21X1_HVT U217 ( .A1(n269), .A2(n351), .S0(n50), .Y(n547) );
  MUX21X1_HVT U219 ( .A1(n325), .A2(n440), .S0(n261), .Y(n439) );
  MUX21X1_HVT U221 ( .A1(n346), .A2(n272), .S0(n265), .Y(n440) );
  MUX21X1_HVT U222 ( .A1(n274), .A2(n272), .S0(n284), .Y(n487) );
  NAND2X0_HVT U223 ( .A1(n357), .A2(n353), .Y(n571) );
  MUX21X1_HVT U224 ( .A1(n351), .A2(n269), .S0(n121), .Y(n362) );
  NBUFFX2_HVT U225 ( .A(n574), .Y(n276) );
  INVX1_HVT U226 ( .A(n575), .Y(n354) );
  MUX21X1_HVT U227 ( .A1(n354), .A2(n267), .S0(n280), .Y(n542) );
  MUX21X1_HVT U228 ( .A1(n269), .A2(n267), .S0(n283), .Y(n453) );
  NBUFFX2_HVT U229 ( .A(n574), .Y(n277) );
  MUX21X1_HVT U230 ( .A1(n267), .A2(n279), .S0(n121), .Y(n388) );
  MUX21X1_HVT U231 ( .A1(n575), .A2(n277), .S0(n282), .Y(n389) );
  MUX21X1_HVT U232 ( .A1(n352), .A2(n351), .S0(n281), .Y(n557) );
  INVX1_HVT U233 ( .A(n566), .Y(n352) );
  MUX21X1_HVT U234 ( .A1(n278), .A2(n272), .S0(n282), .Y(n561) );
  MUX21X1_HVT U235 ( .A1(n273), .A2(n279), .S0(n280), .Y(n482) );
  MUX21X1_HVT U236 ( .A1(n267), .A2(n354), .S0(n281), .Y(n565) );
  MUX21X1_HVT U237 ( .A1(n274), .A2(n267), .S0(n121), .Y(n564) );
  MUX21X1_HVT U238 ( .A1(n242), .A2(n561), .S0(n261), .Y(n476) );
  NBUFFX2_HVT U239 ( .A(n574), .Y(n278) );
  XOR2X1_HVT U240 ( .A1(n284), .A2(n352), .Y(n531) );
  MUX21X1_HVT U241 ( .A1(n267), .A2(n269), .S0(n282), .Y(n385) );
  XOR2X1_HVT U242 ( .A1(n276), .A2(n284), .Y(n528) );
  XNOR2X1_HVT U243 ( .A1(n273), .A2(n284), .Y(n250) );
  MUX21X1_HVT U244 ( .A1(n279), .A2(n272), .S0(n282), .Y(n545) );
  MUX21X1_HVT U245 ( .A1(n276), .A2(n269), .S0(n282), .Y(n368) );
  MUX21X1_HVT U246 ( .A1(n276), .A2(n274), .S0(n284), .Y(n360) );
  XNOR2X1_HVT U247 ( .A1(n575), .A2(n284), .Y(n251) );
  AND2X1_HVT U248 ( .A1(n280), .A2(n355), .Y(n252) );
  MUX21X1_HVT U249 ( .A1(n272), .A2(n267), .S0(n281), .Y(n366) );
  AND2X1_HVT U250 ( .A1(n279), .A2(n463), .Y(n253) );
  MUX21X1_HVT U251 ( .A1(n272), .A2(n269), .S0(n281), .Y(n505) );
  MUX21X1_HVT U252 ( .A1(n566), .A2(n279), .S0(n261), .Y(n450) );
  XOR2X1_HVT U253 ( .A1(n269), .A2(n50), .Y(n550) );
  NBUFFX2_HVT U254 ( .A(n295), .Y(n266) );
  NBUFFX2_HVT U255 ( .A(n295), .Y(n264) );
  NBUFFX2_HVT U256 ( .A(n295), .Y(n265) );
  NBUFFX2_HVT U257 ( .A(n353), .Y(n267) );
  NBUFFX2_HVT U258 ( .A(n292), .Y(n263) );
  NBUFFX2_HVT U259 ( .A(n287), .Y(n259) );
  NBUFFX2_HVT U260 ( .A(n287), .Y(n261) );
  NBUFFX2_HVT U261 ( .A(n287), .Y(n260) );
  NBUFFX2_HVT U262 ( .A(n292), .Y(n262) );
  NBUFFX2_HVT U263 ( .A(n287), .Y(n257) );
  MUX21X1_HVT U264 ( .A1(n356), .A2(n271), .S0(n281), .Y(n553) );
  MUX21X1_HVT U265 ( .A1(n392), .A2(n393), .S0(n260), .Y(n391) );
  MUX21X1_HVT U266 ( .A1(n490), .A2(n271), .S0(n265), .Y(n393) );
  MUX21X1_HVT U267 ( .A1(n474), .A2(n325), .S0(n261), .Y(n471) );
  MUX21X1_HVT U268 ( .A1(n513), .A2(n515), .S0(n260), .Y(n512) );
  XOR2X1_HVT U269 ( .A1(n283), .A2(n271), .Y(n529) );
  MUX21X1_HVT U270 ( .A1(n272), .A2(n268), .S0(n50), .Y(n469) );
  MUX21X1_HVT U271 ( .A1(n497), .A2(n496), .S0(n260), .Y(n494) );
  MUX21X1_HVT U272 ( .A1(n555), .A2(n272), .S0(n266), .Y(n497) );
  MUX21X1_HVT U273 ( .A1(n405), .A2(n404), .S0(n261), .Y(n403) );
  MUX21X1_HVT U274 ( .A1(n566), .A2(n341), .S0(n266), .Y(n405) );
  MUX21X1_HVT U275 ( .A1(n343), .A2(n352), .S0(n265), .Y(n425) );
  AND2X1_HVT U276 ( .A1(n236), .A2(n286), .Y(n254) );
  MUX21X1_HVT U277 ( .A1(n430), .A2(n429), .S0(n261), .Y(n428) );
  MUX21X1_HVT U278 ( .A1(n352), .A2(n355), .S0(n283), .Y(n410) );
  NAND2X0_HVT U279 ( .A1(in[3]), .A2(n357), .Y(n574) );
  MUX21X1_HVT U280 ( .A1(n355), .A2(n271), .S0(n280), .Y(n556) );
  MUX21X1_HVT U281 ( .A1(n271), .A2(n351), .S0(n281), .Y(n537) );
  MUX21X1_HVT U282 ( .A1(n328), .A2(n573), .S0(n259), .Y(n466) );
  MUX21X1_HVT U283 ( .A1(n420), .A2(n278), .S0(n255), .Y(n419) );
  MUX21X1_HVT U284 ( .A1(n558), .A2(n326), .S0(n259), .Y(n442) );
  MUX21X1_HVT U285 ( .A1(n573), .A2(n285), .S0(n260), .Y(n449) );
  MUX21X1_HVT U286 ( .A1(n525), .A2(n526), .S0(n264), .Y(n523) );
  MUX21X1_HVT U287 ( .A1(n271), .A2(n541), .S0(n263), .Y(n526) );
  XOR2X1_HVT U288 ( .A1(n281), .A2(n262), .Y(n533) );
  MUX21X1_HVT U289 ( .A1(n271), .A2(n352), .S0(n50), .Y(n365) );
  NBUFFX2_HVT U290 ( .A(n566), .Y(n272) );
  MUX21X1_HVT U291 ( .A1(n546), .A2(n369), .S0(n264), .Y(n363) );
  MUX21X1_HVT U292 ( .A1(n275), .A2(n271), .S0(n280), .Y(n567) );
  MUX21X1_HVT U293 ( .A1(n322), .A2(n546), .S0(n259), .Y(n445) );
  MUX21X1_HVT U294 ( .A1(n312), .A2(n286), .S0(n263), .Y(n511) );
  MUX21X1_HVT U295 ( .A1(n278), .A2(n485), .S0(n255), .Y(n484) );
  MUX21X1_HVT U296 ( .A1(n271), .A2(n269), .S0(n266), .Y(n485) );
  NBUFFX2_HVT U297 ( .A(n575), .Y(n279) );
  NBUFFX2_HVT U298 ( .A(n357), .Y(n269) );
  XNOR2X1_HVT U299 ( .A1(n297), .A2(n282), .Y(n255) );
  AND2X1_HVT U300 ( .A1(n267), .A2(n286), .Y(n256) );
  NBUFFX2_HVT U301 ( .A(in[5]), .Y(n292) );
  NBUFFX2_HVT U302 ( .A(in[5]), .Y(n291) );
  MUX21X1_HVT U303 ( .A1(n483), .A2(n484), .S0(n261), .Y(n481) );
  MUX21X1_HVT U304 ( .A1(n523), .A2(n527), .S0(n261), .Y(n522) );
  MUX21X1_HVT U305 ( .A1(n517), .A2(n519), .S0(n260), .Y(n516) );
  MUX21X1_HVT U306 ( .A1(n351), .A2(n219), .S0(n50), .Y(n544) );
  NAND2X0_HVT U307 ( .A1(in[3]), .A2(in[4]), .Y(n575) );
  MUX21X1_HVT U308 ( .A1(n219), .A2(n354), .S0(n280), .Y(n540) );
  MUX21X1_HVT U309 ( .A1(n219), .A2(n352), .S0(n280), .Y(n558) );
  MUX21X1_HVT U310 ( .A1(n219), .A2(n237), .S0(n283), .Y(n367) );
  MUX21X1_HVT U311 ( .A1(n219), .A2(n278), .S0(n50), .Y(n555) );
  MUX21X1_HVT U312 ( .A1(n219), .A2(n272), .S0(n281), .Y(n359) );
  MUX21X1_HVT U313 ( .A1(n279), .A2(n219), .S0(n281), .Y(n548) );
  MUX21X1_HVT U314 ( .A1(n271), .A2(n219), .S0(n258), .Y(n461) );
  MUX21X1_HVT U315 ( .A1(n219), .A2(n279), .S0(n280), .Y(n358) );
  MUX21X1_HVT U316 ( .A1(n267), .A2(n219), .S0(n121), .Y(n546) );
  NBUFFX2_HVT U317 ( .A(in[3]), .Y(n271) );
  NBUFFX2_HVT U318 ( .A(in[0]), .Y(n270) );
  INVX0_HVT U319 ( .A(n554), .Y(n299) );
  INVX0_HVT U320 ( .A(n552), .Y(n300) );
  INVX0_HVT U321 ( .A(n543), .Y(n301) );
  INVX0_HVT U322 ( .A(n541), .Y(n302) );
  INVX0_HVT U323 ( .A(n407), .Y(n303) );
  INVX0_HVT U324 ( .A(n370), .Y(n304) );
  INVX0_HVT U325 ( .A(n573), .Y(n305) );
  INVX0_HVT U326 ( .A(n560), .Y(n306) );
  INVX0_HVT U327 ( .A(n572), .Y(n307) );
  INVX0_HVT U328 ( .A(n570), .Y(n308) );
  INVX0_HVT U329 ( .A(n568), .Y(n309) );
  INVX0_HVT U330 ( .A(n567), .Y(n310) );
  INVX0_HVT U331 ( .A(n565), .Y(n311) );
  INVX0_HVT U332 ( .A(n564), .Y(n312) );
  INVX0_HVT U333 ( .A(n561), .Y(n313) );
  INVX0_HVT U334 ( .A(n559), .Y(n314) );
  INVX0_HVT U335 ( .A(n558), .Y(n315) );
  INVX0_HVT U336 ( .A(n557), .Y(n316) );
  INVX0_HVT U337 ( .A(n556), .Y(n317) );
  INVX0_HVT U338 ( .A(n555), .Y(n318) );
  INVX0_HVT U339 ( .A(n553), .Y(n319) );
  INVX0_HVT U340 ( .A(n551), .Y(n320) );
  INVX0_HVT U341 ( .A(n550), .Y(n321) );
  INVX0_HVT U342 ( .A(n548), .Y(n322) );
  INVX0_HVT U343 ( .A(n547), .Y(n323) );
  INVX0_HVT U344 ( .A(n546), .Y(n324) );
  INVX0_HVT U345 ( .A(n363), .Y(n325) );
  INVX0_HVT U346 ( .A(n544), .Y(n326) );
  INVX0_HVT U347 ( .A(n540), .Y(n328) );
  INVX0_HVT U348 ( .A(n537), .Y(n330) );
  INVX0_HVT U349 ( .A(n536), .Y(n331) );
  INVX0_HVT U350 ( .A(n535), .Y(n332) );
  INVX0_HVT U351 ( .A(n534), .Y(n333) );
  INVX0_HVT U352 ( .A(n503), .Y(n334) );
  INVX0_HVT U353 ( .A(n463), .Y(n335) );
  INVX0_HVT U354 ( .A(n369), .Y(n336) );
  INVX0_HVT U355 ( .A(n520), .Y(n337) );
  INVX0_HVT U356 ( .A(n423), .Y(n338) );
  INVX0_HVT U357 ( .A(n368), .Y(n339) );
  INVX0_HVT U358 ( .A(n367), .Y(n340) );
  INVX0_HVT U359 ( .A(n366), .Y(n341) );
  INVX0_HVT U360 ( .A(n365), .Y(n342) );
  INVX0_HVT U361 ( .A(n364), .Y(n343) );
  INVX0_HVT U362 ( .A(n482), .Y(n344) );
  INVX0_HVT U363 ( .A(n472), .Y(n345) );
  INVX0_HVT U364 ( .A(n360), .Y(n348) );
  INVX0_HVT U365 ( .A(n358), .Y(n350) );
endmodule

