
module sbox_2 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n28, n48, n50, n114, n119, n168, n210, n211, n212, n213, n216,
         n217, n218, n219, n224, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599;

  NAND2X0_HVT U4 ( .A1(n312), .A2(n597), .Y(n596) );
  NAND2X0_HVT U5 ( .A1(n318), .A2(n300), .Y(n594) );
  NAND2X0_HVT U15 ( .A1(n597), .A2(n302), .Y(n584) );
  NAND2X0_HVT U21 ( .A1(n312), .A2(n23), .Y(n578) );
  NAND2X0_HVT U24 ( .A1(n308), .A2(n23), .Y(n576) );
  NAND2X0_HVT U33 ( .A1(n381), .A2(n23), .Y(n568) );
  NAND2X0_HVT U35 ( .A1(n304), .A2(n23), .Y(n566) );
  NAND2X0_HVT U42 ( .A1(n239), .A2(n307), .Y(n559) );
  MUX41X1_HVT U51 ( .A1(n370), .A3(n329), .A2(n347), .A4(n348), .S0(n326), 
        .S1(n321), .Y(n552) );
  NAND2X0_HVT U53 ( .A1(n549), .A2(n558), .Y(n550) );
  NAND2X0_HVT U56 ( .A1(n312), .A2(n545), .Y(n546) );
  MUX41X1_HVT U57 ( .A1(n371), .A3(n580), .A2(n546), .A4(n589), .S0(n326), 
        .S1(n321), .Y(n544) );
  NAND2X0_HVT U58 ( .A1(n315), .A2(n597), .Y(n543) );
  MUX41X1_HVT U59 ( .A1(n291), .A3(n543), .A2(n289), .A4(n346), .S0(n326), 
        .S1(n321), .Y(n542) );
  MUX41X1_HVT U61 ( .A1(n287), .A3(n345), .A2(n344), .A4(n301), .S0(n326), 
        .S1(n321), .Y(n540) );
  NAND2X0_HVT U62 ( .A1(n23), .A2(n314), .Y(n539) );
  MUX41X1_HVT U63 ( .A1(n539), .A3(n336), .A2(n365), .A4(n343), .S0(n326), 
        .S1(n321), .Y(n538) );
  AO21X1_HVT U66 ( .A1(n341), .A2(n297), .A3(n364), .Y(n535) );
  MUX41X1_HVT U68 ( .A1(n339), .A3(n535), .A2(n534), .A4(n536), .S0(n293), 
        .S1(n324), .Y(n533) );
  NAND2X0_HVT U73 ( .A1(n310), .A2(n528), .Y(n529) );
  MUX41X1_HVT U74 ( .A1(n530), .A3(n574), .A2(n529), .A4(n576), .S0(n293), 
        .S1(n324), .Y(n527) );
  MUX41X1_HVT U75 ( .A1(n368), .A3(n373), .A2(n384), .A4(n350), .S0(n295), 
        .S1(n324), .Y(n526) );
  MUX41X1_HVT U77 ( .A1(n591), .A3(n374), .A2(n525), .A4(n255), .S0(n243), 
        .S1(n294), .Y(n524) );
  AND3X1_HVT U80 ( .A1(n314), .A2(n545), .A3(n520), .Y(n521) );
  MUX41X1_HVT U82 ( .A1(n556), .A3(n348), .A2(n330), .A4(n585), .S0(n295), 
        .S1(n323), .Y(n518) );
  AND2X1_HVT U83 ( .A1(n318), .A2(n247), .Y(n517) );
  MUX41X1_HVT U84 ( .A1(n349), .A3(n593), .A2(n583), .A4(n517), .S0(n295), 
        .S1(n323), .Y(n516) );
  NAND2X0_HVT U85 ( .A1(n23), .A2(n236), .Y(n515) );
  AO21X1_HVT U93 ( .A1(n299), .A2(n507), .A3(n369), .Y(n508) );
  MUX41X1_HVT U96 ( .A1(n330), .A3(n286), .A2(n372), .A4(n505), .S0(n296), 
        .S1(n324), .Y(n504) );
  MUX41X1_HVT U97 ( .A1(n368), .A3(n286), .A2(n217), .A4(n584), .S0(n295), 
        .S1(n324), .Y(n503) );
  MUX41X1_HVT U98 ( .A1(n503), .A3(n506), .A2(n504), .A4(n511), .S0(n306), 
        .S1(n321), .Y(n502) );
  NAND2X0_HVT U101 ( .A1(n498), .A2(n497), .Y(n499) );
  MUX41X1_HVT U103 ( .A1(n212), .A3(n340), .A2(n257), .A4(n213), .S0(n296), 
        .S1(n324), .Y(n495) );
  MUX41X1_HVT U105 ( .A1(n352), .A3(n554), .A2(n494), .A4(n367), .S0(n295), 
        .S1(n324), .Y(n493) );
  NAND2X0_HVT U110 ( .A1(n314), .A2(n489), .Y(n490) );
  AND2X1_HVT U115 ( .A1(n218), .A2(n301), .Y(n485) );
  NAND2X0_HVT U123 ( .A1(n476), .A2(n475), .Y(n477) );
  MUX41X1_HVT U125 ( .A1(n578), .A3(n291), .A2(n339), .A4(n376), .S0(n292), 
        .S1(n325), .Y(n473) );
  MUX41X1_HVT U131 ( .A1(n468), .A3(n470), .A2(n469), .A4(n471), .S0(n297), 
        .S1(n326), .Y(n467) );
  MUX41X1_HVT U135 ( .A1(n377), .A3(n382), .A2(n594), .A4(n234), .S0(n293), 
        .S1(n325), .Y(n464) );
  MUX41X1_HVT U136 ( .A1(n284), .A3(n568), .A2(n378), .A4(n565), .S0(n292), 
        .S1(n326), .Y(n463) );
  AND2X1_HVT U140 ( .A1(n309), .A2(n320), .Y(n459) );
  MUX41X1_HVT U141 ( .A1(n575), .A3(n248), .A2(n459), .A4(n356), .S0(n293), 
        .S1(n325), .Y(n458) );
  MUX41X1_HVT U142 ( .A1(n349), .A3(n301), .A2(n366), .A4(n309), .S0(n292), 
        .S1(n325), .Y(n457) );
  NAND2X0_HVT U146 ( .A1(n317), .A2(n315), .Y(n528) );
  MUX41X1_HVT U148 ( .A1(n453), .A3(n457), .A2(n454), .A4(n458), .S0(n306), 
        .S1(n321), .Y(n452) );
  OA21X1_HVT U151 ( .A1(n561), .A2(n281), .A3(n449), .Y(n450) );
  MUX41X1_HVT U153 ( .A1(n490), .A3(n287), .A2(n313), .A4(n332), .S0(n292), 
        .S1(n323), .Y(n447) );
  AND2X1_HVT U154 ( .A1(n299), .A2(n308), .Y(n446) );
  NAND2X0_HVT U158 ( .A1(n318), .A2(n236), .Y(n442) );
  MUX41X1_HVT U159 ( .A1(n259), .A3(n301), .A2(n442), .A4(n338), .S0(n292), 
        .S1(n323), .Y(n441) );
  NAND2X0_HVT U166 ( .A1(n315), .A2(n545), .Y(n435) );
  NAND2X0_HVT U167 ( .A1(n384), .A2(n23), .Y(n434) );
  NAND2X0_HVT U174 ( .A1(n317), .A2(n593), .Y(n586) );
  NAND2X0_HVT U177 ( .A1(n318), .A2(n303), .Y(n426) );
  MUX41X1_HVT U178 ( .A1(n582), .A3(n426), .A2(n379), .A4(n563), .S0(n293), 
        .S1(n324), .Y(n425) );
  MUX41X1_HVT U179 ( .A1(n573), .A3(n380), .A2(n334), .A4(n379), .S0(n293), 
        .S1(n324), .Y(n424) );
  MUX41X1_HVT U180 ( .A1(n337), .A3(n591), .A2(n259), .A4(n283), .S0(n243), 
        .S1(n294), .Y(n423) );
  MUX41X1_HVT U181 ( .A1(n423), .A3(n425), .A2(n424), .A4(n427), .S0(n306), 
        .S1(in[5]), .Y(n422) );
  OA21X1_HVT U184 ( .A1(n567), .A2(n281), .A3(n349), .Y(n419) );
  MUX41X1_HVT U189 ( .A1(n415), .A3(n586), .A2(n416), .A4(n367), .S0(n243), 
        .S1(n294), .Y(n414) );
  MUX41X1_HVT U190 ( .A1(n414), .A3(n417), .A2(n418), .A4(n421), .S0(in[5]), 
        .S1(n305), .Y(n413) );
  MUX41X1_HVT U193 ( .A1(n559), .A3(n213), .A2(n553), .A4(n412), .S0(n293), 
        .S1(n323), .Y(n411) );
  MUX41X1_HVT U195 ( .A1(n593), .A3(n372), .A2(n599), .A4(n564), .S0(n294), 
        .S1(n323), .Y(n409) );
  AO21X1_HVT U197 ( .A1(n288), .A2(n298), .A3(n369), .Y(n407) );
  MUX41X1_HVT U199 ( .A1(n406), .A3(n410), .A2(n409), .A4(n411), .S0(n306), 
        .S1(n322), .Y(n405) );
  OA21X1_HVT U201 ( .A1(n592), .A2(n281), .A3(n248), .Y(n403) );
  MUX41X1_HVT U204 ( .A1(n546), .A3(n587), .A2(n357), .A4(n577), .S0(n293), 
        .S1(n323), .Y(n400) );
  MUX41X1_HVT U205 ( .A1(n247), .A3(n597), .A2(n380), .A4(n355), .S0(n294), 
        .S1(n323), .Y(n399) );
  NAND2X0_HVT U208 ( .A1(n317), .A2(n312), .Y(n489) );
  NAND2X0_HVT U212 ( .A1(n239), .A2(n310), .Y(n545) );
  NAND2X0_HVT U214 ( .A1(n593), .A2(n23), .Y(n397) );
  NAND2X0_HVT U215 ( .A1(n489), .A2(n311), .Y(n396) );
  AO21X1_HVT U216 ( .A1(n320), .A2(n382), .A3(n281), .Y(n498) );
  NAND2X0_HVT U218 ( .A1(n382), .A2(n318), .Y(n449) );
  NAND2X0_HVT U220 ( .A1(n298), .A2(n397), .Y(n520) );
  INVX2_HVT U1 ( .A(n327), .Y(n324) );
  NBUFFX2_HVT U2 ( .A(n238), .Y(n23) );
  INVX0_HVT U3 ( .A(in[1]), .Y(n238) );
  INVX1_HVT U6 ( .A(n238), .Y(n239) );
  MUX41X1_HVT U7 ( .A1(n486), .A3(n472), .A2(n480), .A4(n467), .S0(n246), .S1(
        n249), .Y(out[3]) );
  INVX2_HVT U8 ( .A(n305), .Y(n249) );
  MUX21X2_HVT U9 ( .A1(n550), .A2(n551), .S0(n243), .Y(n548) );
  INVX1_HVT U10 ( .A(in[6]), .Y(n48) );
  MUX21X2_HVT U11 ( .A1(n484), .A2(n481), .S0(n28), .Y(n480) );
  IBUFFX16_HVT U12 ( .A(n297), .Y(n28) );
  INVX2_HVT U13 ( .A(in[1]), .Y(n320) );
  INVX1_HVT U14 ( .A(n320), .Y(n316) );
  MUX21X2_HVT U16 ( .A1(n422), .A2(n413), .S0(n48), .Y(out[6]) );
  IBUFFX2_HVT U17 ( .A(n592), .Y(n339) );
  MUX21X2_HVT U18 ( .A1(n477), .A2(n478), .S0(n50), .Y(n474) );
  IBUFFX16_HVT U19 ( .A(n299), .Y(n50) );
  MUX21X2_HVT U20 ( .A1(n482), .A2(n483), .S0(n298), .Y(n481) );
  OR2X1_HVT U22 ( .A1(n320), .A2(n114), .Y(n597) );
  IBUFFX16_HVT U23 ( .A(n598), .Y(n114) );
  IBUFFX2_HVT U25 ( .A(n320), .Y(n319) );
  MUX21X2_HVT U26 ( .A1(n450), .A2(n451), .S0(n119), .Y(n448) );
  IBUFFX16_HVT U27 ( .A(n219), .Y(n119) );
  MUX41X1_HVT U28 ( .A1(n447), .A3(n441), .A2(n448), .A4(n443), .S0(n168), 
        .S1(n210), .Y(n440) );
  IBUFFX16_HVT U29 ( .A(n306), .Y(n168) );
  IBUFFX16_HVT U30 ( .A(n256), .Y(n210) );
  MUX41X1_HVT U31 ( .A1(n284), .A3(n288), .A2(n515), .A4(n373), .S0(n211), 
        .S1(n327), .Y(n514) );
  IBUFFX16_HVT U32 ( .A(n295), .Y(n211) );
  MUX41X1_HVT U34 ( .A1(n518), .A3(n514), .A2(n519), .A4(n516), .S0(n237), 
        .S1(n322), .Y(n513) );
  INVX0_HVT U36 ( .A(n335), .Y(n212) );
  INVX0_HVT U37 ( .A(n332), .Y(n213) );
  INVX4_HVT U38 ( .A(n327), .Y(n323) );
  NBUFFX2_HVT U39 ( .A(n316), .Y(n216) );
  NBUFFX2_HVT U40 ( .A(n316), .Y(n217) );
  NBUFFX2_HVT U41 ( .A(n316), .Y(n218) );
  IBUFFX2_HVT U43 ( .A(n320), .Y(n317) );
  INVX0_HVT U44 ( .A(n298), .Y(n254) );
  MUX21X1_HVT U45 ( .A1(n311), .A2(n579), .S0(n328), .Y(n522) );
  INVX1_HVT U46 ( .A(n306), .Y(n237) );
  MUX21X1_HVT U47 ( .A1(n255), .A2(n382), .S0(n298), .Y(n451) );
  NAND2X0_HVT U48 ( .A1(n444), .A2(n219), .Y(n224) );
  INVX1_HVT U49 ( .A(n328), .Y(n326) );
  MUX21X1_HVT U50 ( .A1(n354), .A2(n466), .S0(n295), .Y(n465) );
  MUX21X1_HVT U52 ( .A1(n253), .A2(n390), .S0(n254), .Y(n252) );
  INVX0_HVT U54 ( .A(n311), .Y(n253) );
  MUX21X1_HVT U55 ( .A1(n462), .A2(n596), .S0(n296), .Y(n461) );
  MUX21X1_HVT U60 ( .A1(n532), .A2(n557), .S0(n265), .Y(n531) );
  INVX1_HVT U64 ( .A(n326), .Y(n260) );
  INVX1_HVT U65 ( .A(in[6]), .Y(n246) );
  INVX1_HVT U67 ( .A(n320), .Y(n318) );
  INVX0_HVT U69 ( .A(n294), .Y(n265) );
  NBUFFX2_HVT U70 ( .A(in[2]), .Y(n292) );
  NBUFFX2_HVT U71 ( .A(n239), .Y(n240) );
  INVX1_HVT U72 ( .A(n313), .Y(n235) );
  NBUFFX2_HVT U76 ( .A(n385), .Y(n303) );
  INVX1_HVT U78 ( .A(n599), .Y(n236) );
  INVX0_HVT U79 ( .A(n281), .Y(n243) );
  INVX1_HVT U81 ( .A(n322), .Y(n256) );
  NBUFFX2_HVT U86 ( .A(in[2]), .Y(n293) );
  INVX1_HVT U87 ( .A(n296), .Y(n219) );
  NBUFFX2_HVT U88 ( .A(in[2]), .Y(n296) );
  INVX1_HVT U89 ( .A(n293), .Y(n258) );
  NAND2X0_HVT U90 ( .A1(n445), .A2(n296), .Y(n231) );
  NAND2X0_HVT U91 ( .A1(n224), .A2(n231), .Y(n443) );
  NAND2X0_HVT U92 ( .A1(n429), .A2(n246), .Y(n232) );
  NAND2X0_HVT U94 ( .A1(n440), .A2(in[6]), .Y(n233) );
  NAND2X0_HVT U95 ( .A1(n232), .A2(n233), .Y(out[5]) );
  MUX21X1_HVT U99 ( .A1(n374), .A2(n563), .S0(n260), .Y(n444) );
  MUX21X1_HVT U100 ( .A1(n446), .A2(n314), .S0(n290), .Y(n445) );
  MUX41X1_HVT U102 ( .A1(n547), .A3(n537), .A2(n541), .A4(n533), .S0(n246), 
        .S1(n249), .Y(out[0]) );
  MUX21X1_HVT U104 ( .A1(n235), .A2(n236), .S0(n239), .Y(n234) );
  MUX21X2_HVT U106 ( .A1(n473), .A2(n474), .S0(n297), .Y(n472) );
  MUX41X1_HVT U107 ( .A1(n555), .A3(n528), .A2(n562), .A4(n286), .S0(n219), 
        .S1(n327), .Y(n417) );
  IBUFFX2_HVT U108 ( .A(n589), .Y(n341) );
  MUX21X2_HVT U109 ( .A1(n452), .A2(n460), .S0(in[6]), .Y(out[4]) );
  MUX41X1_HVT U111 ( .A1(n570), .A3(n350), .A2(n485), .A4(n259), .S0(n219), 
        .S1(n260), .Y(n484) );
  MUX21X2_HVT U112 ( .A1(n521), .A2(n522), .S0(n265), .Y(n519) );
  IBUFFX2_HVT U113 ( .A(n579), .Y(n348) );
  INVX0_HVT U114 ( .A(n390), .Y(n376) );
  INVX0_HVT U116 ( .A(n257), .Y(n572) );
  OA21X1_HVT U117 ( .A1(n289), .A2(n328), .A3(n570), .Y(n431) );
  OA21X1_HVT U118 ( .A1(n333), .A2(n281), .A3(n570), .Y(n455) );
  MUX41X1_HVT U119 ( .A1(n370), .A3(n512), .A2(n555), .A4(n559), .S0(n292), 
        .S1(n327), .Y(n511) );
  NAND2X0_HVT U120 ( .A1(n502), .A2(n261), .Y(n241) );
  NAND2X0_HVT U121 ( .A1(n492), .A2(n246), .Y(n242) );
  NAND2X0_HVT U122 ( .A1(n241), .A2(n242), .Y(out[2]) );
  MUX21X1_HVT U124 ( .A1(n355), .A2(n585), .S0(n296), .Y(n501) );
  INVX0_HVT U126 ( .A(n570), .Y(n355) );
  MUX21X1_HVT U127 ( .A1(n599), .A2(n310), .S0(n216), .Y(n570) );
  XNOR2X2_HVT U128 ( .A1(n243), .A2(n234), .Y(n557) );
  XOR2X2_HVT U129 ( .A1(n262), .A2(n238), .Y(n555) );
  NAND2X0_HVT U130 ( .A1(n508), .A2(n258), .Y(n244) );
  NAND2X0_HVT U132 ( .A1(n509), .A2(n296), .Y(n245) );
  NAND2X0_HVT U133 ( .A1(n244), .A2(n245), .Y(n506) );
  MUX21X1_HVT U134 ( .A1(n314), .A2(n510), .S0(n290), .Y(n509) );
  INVX1_HVT U137 ( .A(n252), .Y(n466) );
  MUX21X1_HVT U138 ( .A1(n384), .A2(n307), .S0(n318), .Y(n580) );
  INVX2_HVT U139 ( .A(in[7]), .Y(n327) );
  MUX21X1_HVT U143 ( .A1(n300), .A2(n384), .S0(n239), .Y(n561) );
  INVX1_HVT U144 ( .A(n248), .Y(n563) );
  NBUFFX2_HVT U145 ( .A(in[4]), .Y(n247) );
  MUX21X1_HVT U147 ( .A1(n595), .A2(n599), .S0(n238), .Y(n248) );
  INVX1_HVT U149 ( .A(n595), .Y(n381) );
  MUX41X1_HVT U150 ( .A1(n531), .A3(n526), .A2(n527), .A4(n524), .S0(n249), 
        .S1(n256), .Y(n523) );
  INVX1_HVT U152 ( .A(n313), .Y(n384) );
  MUX21X2_HVT U155 ( .A1(n542), .A2(n544), .S0(n294), .Y(n541) );
  NAND2X0_HVT U156 ( .A1(n398), .A2(n246), .Y(n250) );
  NAND2X0_HVT U157 ( .A1(n405), .A2(n261), .Y(n251) );
  NAND2X0_HVT U160 ( .A1(n250), .A2(n251), .Y(out[7]) );
  INVX0_HVT U161 ( .A(n246), .Y(n261) );
  IBUFFX2_HVT U162 ( .A(n561), .Y(n361) );
  MUX41X1_HVT U163 ( .A1(n463), .A3(n465), .A2(n461), .A4(n464), .S0(n306), 
        .S1(n256), .Y(n460) );
  MUX21X1_HVT U164 ( .A1(n303), .A2(n381), .S0(n238), .Y(n390) );
  INVX0_HVT U165 ( .A(n569), .Y(n356) );
  MUX21X1_HVT U168 ( .A1(n308), .A2(n262), .S0(n316), .Y(n255) );
  INVX1_HVT U169 ( .A(n262), .Y(n593) );
  MUX21X1_HVT U170 ( .A1(n247), .A2(n595), .S0(n216), .Y(n257) );
  MUX41X1_HVT U171 ( .A1(n569), .A3(n588), .A2(n361), .A4(n565), .S0(n258), 
        .S1(n327), .Y(n401) );
  INVX0_HVT U172 ( .A(n365), .Y(n259) );
  NAND2X0_HVT U173 ( .A1(n586), .A2(n315), .Y(n587) );
  MUX21X2_HVT U175 ( .A1(n572), .A2(n335), .S0(n299), .Y(n456) );
  MUX21X2_HVT U176 ( .A1(n456), .A2(n455), .S0(n295), .Y(n454) );
  MUX21X1_HVT U182 ( .A1(n577), .A2(n360), .S0(n298), .Y(n462) );
  INVX1_HVT U183 ( .A(n562), .Y(n360) );
  MUX41X1_HVT U185 ( .A1(n555), .A3(n368), .A2(n528), .A4(n378), .S0(n219), 
        .S1(n260), .Y(n453) );
  INVX1_HVT U186 ( .A(in[4]), .Y(n385) );
  MUX41X1_HVT U187 ( .A1(n586), .A3(n375), .A2(n428), .A4(n304), .S0(n260), 
        .S1(n265), .Y(n427) );
  MUX21X2_HVT U188 ( .A1(n432), .A2(n431), .S0(n295), .Y(n430) );
  MUX21X2_HVT U191 ( .A1(n538), .A2(n540), .S0(n294), .Y(n537) );
  INVX1_HVT U192 ( .A(n393), .Y(n372) );
  MUX21X2_HVT U194 ( .A1(n331), .A2(n479), .S0(n293), .Y(n478) );
  MUX21X1_HVT U196 ( .A1(n308), .A2(n302), .S0(n320), .Y(n577) );
  XNOR2X2_HVT U198 ( .A1(n385), .A2(in[3]), .Y(n262) );
  IBUFFX2_HVT U200 ( .A(n560), .Y(n362) );
  MUX41X1_HVT U202 ( .A1(n351), .A3(n362), .A2(n595), .A4(n360), .S0(n328), 
        .S1(n219), .Y(n421) );
  INVX1_HVT U203 ( .A(n281), .Y(n325) );
  NBUFFX2_HVT U206 ( .A(n385), .Y(n304) );
  INVX1_HVT U207 ( .A(n501), .Y(n273) );
  INVX0_HVT U209 ( .A(n285), .Y(n268) );
  INVX0_HVT U210 ( .A(n491), .Y(n279) );
  INVX1_HVT U211 ( .A(n266), .Y(n274) );
  INVX0_HVT U213 ( .A(n287), .Y(n272) );
  INVX1_HVT U217 ( .A(n487), .Y(n276) );
  INVX1_HVT U219 ( .A(n488), .Y(n280) );
  MUX21X1_HVT U221 ( .A1(n285), .A2(n344), .S0(n292), .Y(n469) );
  INVX1_HVT U222 ( .A(n267), .Y(n438) );
  MUX21X1_HVT U223 ( .A1(n302), .A2(n300), .S0(n240), .Y(n583) );
  INVX1_HVT U224 ( .A(n577), .Y(n349) );
  INVX1_HVT U225 ( .A(in[7]), .Y(n328) );
  INVX1_HVT U226 ( .A(in[7]), .Y(n281) );
  MUX41X1_HVT U227 ( .A1(n435), .A3(n434), .A2(n309), .A4(n371), .S0(n258), 
        .S1(n328), .Y(n433) );
  MUX41X1_HVT U228 ( .A1(n438), .A3(n433), .A2(n436), .A4(n430), .S0(n249), 
        .S1(n256), .Y(n429) );
  NBUFFX2_HVT U229 ( .A(n262), .Y(n302) );
  NAND2X0_HVT U230 ( .A1(n283), .A2(n243), .Y(n263) );
  NAND2X0_HVT U231 ( .A1(n583), .A2(n260), .Y(n264) );
  NAND2X0_HVT U232 ( .A1(n263), .A2(n264), .Y(n404) );
  MUX21X2_HVT U233 ( .A1(n404), .A2(n403), .S0(n265), .Y(n402) );
  MUX41X1_HVT U234 ( .A1(n402), .A3(n400), .A2(n401), .A4(n399), .S0(n249), 
        .S1(n256), .Y(n398) );
  AND3X2_HVT U235 ( .A1(n295), .A2(n23), .A3(n247), .Y(n470) );
  AO21X2_HVT U236 ( .A1(n296), .A2(n309), .A3(n593), .Y(n482) );
  XOR2X1_HVT U237 ( .A1(n219), .A2(n328), .Y(n266) );
  MUX41X1_HVT U238 ( .A1(n500), .A3(n495), .A2(n496), .A4(n493), .S0(n249), 
        .S1(n256), .Y(n492) );
  INVX1_HVT U239 ( .A(n439), .Y(n269) );
  MUX41X1_HVT U240 ( .A1(n270), .A3(n582), .A2(n269), .A4(n268), .S0(n258), 
        .S1(n323), .Y(n267) );
  NAND2X0_HVT U241 ( .A1(n593), .A2(n528), .Y(n270) );
  INVX0_HVT U242 ( .A(n271), .Y(n500) );
  MUX21X2_HVT U243 ( .A1(n513), .A2(n523), .S0(in[6]), .Y(out[1]) );
  MUX41X1_HVT U244 ( .A1(n309), .A3(n377), .A2(n234), .A4(n560), .S0(n260), 
        .S1(n265), .Y(n410) );
  MUX41X1_HVT U245 ( .A1(n437), .A3(n555), .A2(n353), .A4(n578), .S0(n281), 
        .S1(n219), .Y(n436) );
  MUX21X1_HVT U246 ( .A1(n273), .A2(n272), .S0(n274), .Y(n271) );
  XNOR2X1_HVT U247 ( .A1(n23), .A2(n219), .Y(n277) );
  INVX1_HVT U248 ( .A(n278), .Y(n486) );
  MUX21X2_HVT U249 ( .A1(n235), .A2(n276), .S0(n277), .Y(n275) );
  MUX41X1_HVT U250 ( .A1(n280), .A3(n282), .A2(n275), .A4(n279), .S0(in[5]), 
        .S1(n328), .Y(n278) );
  OAI21X1_HVT U251 ( .A1(n359), .A2(n219), .A3(n346), .Y(n282) );
  INVX0_HVT U252 ( .A(in[3]), .Y(n383) );
  NBUFFX2_HVT U253 ( .A(n262), .Y(n301) );
  AND2X1_HVT U254 ( .A1(n301), .A2(n545), .Y(n283) );
  MUX21X1_HVT U255 ( .A1(n381), .A2(n236), .S0(n297), .Y(n549) );
  NBUFFX2_HVT U256 ( .A(n595), .Y(n312) );
  MUX21X1_HVT U257 ( .A1(n340), .A2(n382), .S0(n297), .Y(n534) );
  MUX21X1_HVT U258 ( .A1(n570), .A2(n490), .S0(n292), .Y(n488) );
  AND2X1_HVT U259 ( .A1(n314), .A2(n528), .Y(n284) );
  MUX21X1_HVT U260 ( .A1(n301), .A2(n236), .S0(n319), .Y(n592) );
  MUX21X1_HVT U261 ( .A1(n314), .A2(n302), .S0(n316), .Y(n560) );
  MUX21X1_HVT U262 ( .A1(n301), .A2(n303), .S0(n319), .Y(n497) );
  MUX21X1_HVT U263 ( .A1(n381), .A2(n384), .S0(n318), .Y(n428) );
  MUX21X1_HVT U264 ( .A1(n236), .A2(n302), .S0(n317), .Y(n439) );
  MUX21X1_HVT U265 ( .A1(n302), .A2(n381), .S0(n319), .Y(n505) );
  MUX21X1_HVT U266 ( .A1(n312), .A2(n593), .S0(n317), .Y(n564) );
  MUX21X1_HVT U267 ( .A1(n593), .A2(n382), .S0(n318), .Y(n389) );
  MUX21X1_HVT U268 ( .A1(n593), .A2(n384), .S0(n217), .Y(n575) );
  MUX21X1_HVT U269 ( .A1(n312), .A2(n311), .S0(n317), .Y(n512) );
  MUX21X1_HVT U270 ( .A1(n593), .A2(n304), .S0(n217), .Y(n525) );
  MUX21X1_HVT U271 ( .A1(n236), .A2(n300), .S0(n316), .Y(n567) );
  MUX21X1_HVT U272 ( .A1(n332), .A2(n357), .S0(n292), .Y(n483) );
  NAND2X0_HVT U273 ( .A1(n304), .A2(n383), .Y(n595) );
  NBUFFX2_HVT U274 ( .A(n598), .Y(n313) );
  MUX21X1_HVT U275 ( .A1(n314), .A2(n310), .S0(n216), .Y(n585) );
  MUX21X1_HVT U276 ( .A1(n595), .A2(n315), .S0(n319), .Y(n507) );
  MUX21X1_HVT U277 ( .A1(n382), .A2(n381), .S0(n240), .Y(n581) );
  MUX21X1_HVT U278 ( .A1(n303), .A2(n300), .S0(n316), .Y(n479) );
  NBUFFX2_HVT U279 ( .A(n598), .Y(n314) );
  XOR2X1_HVT U280 ( .A1(n218), .A2(n382), .Y(n556) );
  MUX21X1_HVT U281 ( .A1(n300), .A2(n315), .S0(n218), .Y(n415) );
  MUX21X1_HVT U282 ( .A1(n599), .A2(n314), .S0(n319), .Y(n416) );
  INVX1_HVT U283 ( .A(n309), .Y(n382) );
  MUX21X1_HVT U284 ( .A1(n300), .A2(n236), .S0(n318), .Y(n589) );
  MUX21X1_HVT U285 ( .A1(n312), .A2(n300), .S0(n319), .Y(n588) );
  MUX21X1_HVT U286 ( .A1(n300), .A2(n304), .S0(n216), .Y(n412) );
  XOR2X1_HVT U287 ( .A1(n313), .A2(n317), .Y(n553) );
  MUX21X1_HVT U288 ( .A1(n313), .A2(n303), .S0(n317), .Y(n395) );
  XNOR2X1_HVT U289 ( .A1(n595), .A2(n317), .Y(n285) );
  AND2X1_HVT U290 ( .A1(n239), .A2(n384), .Y(n286) );
  MUX21X1_HVT U291 ( .A1(n313), .A2(n312), .S0(n239), .Y(n388) );
  AND2X1_HVT U292 ( .A1(n315), .A2(n489), .Y(n287) );
  XNOR2X1_HVT U293 ( .A1(n599), .A2(n319), .Y(n288) );
  MUX21X1_HVT U294 ( .A1(n310), .A2(n300), .S0(n239), .Y(n393) );
  MUX21X1_HVT U295 ( .A1(n311), .A2(n304), .S0(n217), .Y(n530) );
  MUX21X1_HVT U296 ( .A1(n311), .A2(n315), .S0(n295), .Y(n476) );
  XOR2X1_HVT U297 ( .A1(n304), .A2(n217), .Y(n574) );
  NBUFFX2_HVT U298 ( .A(n325), .Y(n299) );
  NBUFFX2_HVT U299 ( .A(n325), .Y(n298) );
  NBUFFX2_HVT U300 ( .A(n383), .Y(n300) );
  NBUFFX2_HVT U301 ( .A(n322), .Y(n297) );
  NBUFFX2_HVT U302 ( .A(in[2]), .Y(n295) );
  NBUFFX2_HVT U303 ( .A(in[2]), .Y(n294) );
  MUX21X1_HVT U304 ( .A1(n499), .A2(n354), .S0(n295), .Y(n496) );
  MUX21X1_HVT U305 ( .A1(n419), .A2(n420), .S0(n294), .Y(n418) );
  MUX21X1_HVT U306 ( .A1(n515), .A2(n307), .S0(n298), .Y(n420) );
  XOR2X1_HVT U307 ( .A1(n240), .A2(n308), .Y(n554) );
  MUX21X1_HVT U308 ( .A1(n310), .A2(n301), .S0(n239), .Y(n494) );
  MUX21X1_HVT U309 ( .A1(n311), .A2(n372), .S0(n299), .Y(n432) );
  MUX21X1_HVT U310 ( .A1(n382), .A2(n384), .S0(n319), .Y(n437) );
  AND2X1_HVT U311 ( .A1(n301), .A2(n23), .Y(n289) );
  MUX21X1_HVT U312 ( .A1(n307), .A2(n381), .S0(n316), .Y(n562) );
  MUX21X1_HVT U313 ( .A1(n236), .A2(n372), .S0(n299), .Y(n532) );
  MUX21X1_HVT U314 ( .A1(n582), .A2(n356), .S0(n293), .Y(n468) );
  NAND2X0_HVT U315 ( .A1(n308), .A2(n303), .Y(n598) );
  MUX21X1_HVT U316 ( .A1(n358), .A2(n597), .S0(n293), .Y(n491) );
  MUX21X1_HVT U317 ( .A1(n308), .A2(n566), .S0(n297), .Y(n551) );
  XOR2X1_HVT U318 ( .A1(n318), .A2(n322), .Y(n558) );
  MUX21X1_HVT U319 ( .A1(n597), .A2(n320), .S0(n294), .Y(n475) );
  NBUFFX2_HVT U320 ( .A(n590), .Y(n309) );
  MUX21X1_HVT U321 ( .A1(n307), .A2(n382), .S0(n317), .Y(n392) );
  MUX21X1_HVT U322 ( .A1(n571), .A2(n396), .S0(n243), .Y(n391) );
  MUX21X1_HVT U323 ( .A1(n312), .A2(n308), .S0(n316), .Y(n591) );
  MUX21X1_HVT U324 ( .A1(n342), .A2(n23), .S0(n297), .Y(n536) );
  MUX21X1_HVT U325 ( .A1(n363), .A2(n379), .S0(n298), .Y(n408) );
  MUX21X1_HVT U326 ( .A1(n307), .A2(n303), .S0(n299), .Y(n510) );
  NBUFFX2_HVT U327 ( .A(n590), .Y(n310) );
  MUX21X1_HVT U328 ( .A1(n352), .A2(n571), .S0(n293), .Y(n471) );
  NBUFFX2_HVT U329 ( .A(n590), .Y(n311) );
  NBUFFX2_HVT U330 ( .A(n599), .Y(n315) );
  XNOR2X1_HVT U331 ( .A1(n328), .A2(n319), .Y(n290) );
  AND2X1_HVT U332 ( .A1(n300), .A2(n23), .Y(n291) );
  NBUFFX2_HVT U333 ( .A(in[5]), .Y(n322) );
  NBUFFX2_HVT U334 ( .A(in[5]), .Y(n321) );
  MUX21X1_HVT U335 ( .A1(n408), .A2(n407), .S0(n294), .Y(n406) );
  MUX21X1_HVT U336 ( .A1(n548), .A2(n552), .S0(n295), .Y(n547) );
  MUX21X1_HVT U337 ( .A1(n381), .A2(n247), .S0(n318), .Y(n569) );
  NAND2X0_HVT U338 ( .A1(n307), .A2(in[4]), .Y(n599) );
  MUX21X1_HVT U339 ( .A1(n247), .A2(n593), .S0(n319), .Y(n394) );
  MUX21X1_HVT U340 ( .A1(n247), .A2(n236), .S0(n218), .Y(n565) );
  MUX21X1_HVT U341 ( .A1(n247), .A2(n382), .S0(n240), .Y(n582) );
  NAND2X0_HVT U342 ( .A1(in[4]), .A2(n383), .Y(n590) );
  MUX21X1_HVT U343 ( .A1(n247), .A2(n314), .S0(n239), .Y(n579) );
  MUX21X1_HVT U344 ( .A1(n247), .A2(n310), .S0(n239), .Y(n387) );
  MUX21X1_HVT U345 ( .A1(n315), .A2(n247), .S0(n218), .Y(n573) );
  MUX21X1_HVT U346 ( .A1(n308), .A2(n247), .S0(n292), .Y(n487) );
  MUX21X1_HVT U347 ( .A1(n247), .A2(n315), .S0(n317), .Y(n386) );
  MUX21X1_HVT U348 ( .A1(n300), .A2(n247), .S0(n316), .Y(n571) );
  NBUFFX2_HVT U349 ( .A(in[3]), .Y(n307) );
  NBUFFX2_HVT U350 ( .A(in[3]), .Y(n308) );
  NBUFFX2_HVT U351 ( .A(in[0]), .Y(n306) );
  NBUFFX2_HVT U352 ( .A(in[0]), .Y(n305) );
  INVX0_HVT U353 ( .A(n578), .Y(n329) );
  INVX0_HVT U354 ( .A(n576), .Y(n330) );
  INVX0_HVT U355 ( .A(n568), .Y(n331) );
  INVX0_HVT U356 ( .A(n566), .Y(n332) );
  INVX0_HVT U357 ( .A(n434), .Y(n333) );
  INVX0_HVT U358 ( .A(n397), .Y(n334) );
  INVX0_HVT U359 ( .A(n597), .Y(n335) );
  INVX0_HVT U360 ( .A(n584), .Y(n336) );
  INVX0_HVT U361 ( .A(n596), .Y(n337) );
  INVX0_HVT U362 ( .A(n594), .Y(n338) );
  INVX0_HVT U363 ( .A(n591), .Y(n340) );
  INVX0_HVT U364 ( .A(n588), .Y(n342) );
  INVX0_HVT U365 ( .A(n585), .Y(n343) );
  INVX0_HVT U366 ( .A(n583), .Y(n344) );
  INVX0_HVT U367 ( .A(n582), .Y(n345) );
  INVX0_HVT U368 ( .A(n581), .Y(n346) );
  INVX0_HVT U369 ( .A(n580), .Y(n347) );
  INVX0_HVT U370 ( .A(n575), .Y(n350) );
  INVX0_HVT U371 ( .A(n574), .Y(n351) );
  INVX0_HVT U372 ( .A(n573), .Y(n352) );
  INVX0_HVT U373 ( .A(n571), .Y(n353) );
  INVX0_HVT U374 ( .A(n391), .Y(n354) );
  INVX0_HVT U375 ( .A(n567), .Y(n357) );
  INVX0_HVT U376 ( .A(n565), .Y(n358) );
  INVX0_HVT U377 ( .A(n564), .Y(n359) );
  INVX0_HVT U378 ( .A(n559), .Y(n363) );
  INVX0_HVT U379 ( .A(n528), .Y(n364) );
  INVX0_HVT U380 ( .A(n587), .Y(n365) );
  INVX0_HVT U381 ( .A(n489), .Y(n366) );
  INVX0_HVT U382 ( .A(n396), .Y(n367) );
  INVX0_HVT U383 ( .A(n545), .Y(n368) );
  INVX0_HVT U384 ( .A(n449), .Y(n369) );
  INVX0_HVT U385 ( .A(n395), .Y(n370) );
  INVX0_HVT U386 ( .A(n394), .Y(n371) );
  INVX0_HVT U387 ( .A(n392), .Y(n373) );
  INVX0_HVT U388 ( .A(n507), .Y(n374) );
  INVX0_HVT U389 ( .A(n497), .Y(n375) );
  INVX0_HVT U390 ( .A(n389), .Y(n377) );
  INVX0_HVT U391 ( .A(n388), .Y(n378) );
  INVX0_HVT U392 ( .A(n387), .Y(n379) );
  INVX0_HVT U393 ( .A(n386), .Y(n380) );
endmodule

