
module sbox_2 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n26, n45, n48, n50, n87, n121, n210, n211, n212, n213, n216,
         n217, n218, n219, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600;

  NAND2X0_HVT U4 ( .A1(n310), .A2(n598), .Y(n597) );
  NAND2X0_HVT U5 ( .A1(n319), .A2(n382), .Y(n595) );
  NAND2X0_HVT U13 ( .A1(n587), .A2(n314), .Y(n588) );
  NAND2X0_HVT U15 ( .A1(n598), .A2(n301), .Y(n585) );
  NAND2X0_HVT U21 ( .A1(n309), .A2(n322), .Y(n579) );
  NAND2X0_HVT U24 ( .A1(n212), .A2(n210), .Y(n577) );
  NAND2X0_HVT U33 ( .A1(n380), .A2(n322), .Y(n569) );
  NAND2X0_HVT U35 ( .A1(n302), .A2(n322), .Y(n567) );
  NAND2X0_HVT U42 ( .A1(n87), .A2(n23), .Y(n560) );
  MUX41X1_HVT U51 ( .A1(n368), .A3(n329), .A2(n346), .A4(n347), .S0(n325), 
        .S1(n294), .Y(n554) );
  NAND2X0_HVT U53 ( .A1(n551), .A2(n559), .Y(n552) );
  NAND2X0_HVT U56 ( .A1(n310), .A2(n547), .Y(n548) );
  MUX41X1_HVT U57 ( .A1(n369), .A3(n581), .A2(n548), .A4(n590), .S0(n325), 
        .S1(n294), .Y(n546) );
  NAND2X0_HVT U58 ( .A1(n314), .A2(n598), .Y(n545) );
  MUX41X1_HVT U59 ( .A1(n287), .A3(n545), .A2(n285), .A4(n345), .S0(n325), 
        .S1(n294), .Y(n544) );
  MUX41X1_HVT U61 ( .A1(n283), .A3(n344), .A2(n250), .A4(n300), .S0(n325), 
        .S1(n294), .Y(n542) );
  NAND2X0_HVT U62 ( .A1(n322), .A2(n313), .Y(n541) );
  MUX41X1_HVT U63 ( .A1(n541), .A3(n336), .A2(n273), .A4(n343), .S0(n325), 
        .S1(n294), .Y(n540) );
  AO21X1_HVT U66 ( .A1(n341), .A2(n296), .A3(n363), .Y(n537) );
  MUX41X1_HVT U68 ( .A1(n339), .A3(n537), .A2(n536), .A4(n538), .S0(n288), 
        .S1(n264), .Y(n535) );
  NAND2X0_HVT U73 ( .A1(n307), .A2(n530), .Y(n531) );
  MUX41X1_HVT U74 ( .A1(n532), .A3(n576), .A2(n531), .A4(n577), .S0(n290), 
        .S1(n264), .Y(n529) );
  MUX41X1_HVT U75 ( .A1(n366), .A3(n371), .A2(n384), .A4(n241), .S0(n288), 
        .S1(n264), .Y(n528) );
  MUX41X1_HVT U77 ( .A1(n592), .A3(n373), .A2(n527), .A4(n372), .S0(n297), 
        .S1(n323), .Y(n526) );
  MUX41X1_HVT U78 ( .A1(n526), .A3(n529), .A2(n528), .A4(n533), .S0(n304), 
        .S1(n294), .Y(n525) );
  AND3X1_HVT U80 ( .A1(n312), .A2(n547), .A3(n522), .Y(n523) );
  NAND2X0_HVT U85 ( .A1(n322), .A2(n383), .Y(n518) );
  MUX41X1_HVT U86 ( .A1(n371), .A3(n518), .A2(n284), .A4(n280), .S0(n288), 
        .S1(n216), .Y(n517) );
  MUX41X1_HVT U87 ( .A1(n517), .A3(n520), .A2(n519), .A4(n521), .S0(n304), 
        .S1(in[5]), .Y(n516) );
  AO21X1_HVT U93 ( .A1(n326), .A2(n510), .A3(n367), .Y(n511) );
  MUX41X1_HVT U96 ( .A1(n330), .A3(n282), .A2(n370), .A4(n508), .S0(n288), 
        .S1(n216), .Y(n507) );
  MUX41X1_HVT U97 ( .A1(n366), .A3(n282), .A2(n121), .A4(n585), .S0(n288), 
        .S1(n216), .Y(n506) );
  NAND2X0_HVT U101 ( .A1(n501), .A2(n500), .Y(n502) );
  MUX41X1_HVT U105 ( .A1(n350), .A3(n556), .A2(n497), .A4(n365), .S0(n288), 
        .S1(n216), .Y(n496) );
  MUX41X1_HVT U106 ( .A1(n496), .A3(n499), .A2(n498), .A4(n503), .S0(in[0]), 
        .S1(in[5]), .Y(n495) );
  OA21X1_HVT U109 ( .A1(n357), .A2(n238), .A3(n345), .Y(n493) );
  NAND2X0_HVT U110 ( .A1(n312), .A2(n491), .Y(n492) );
  MUX41X1_HVT U114 ( .A1(n488), .A3(n494), .A2(n490), .A4(n493), .S0(n296), 
        .S1(n216), .Y(n487) );
  NAND2X0_HVT U123 ( .A1(n478), .A2(n477), .Y(n479) );
  MUX41X1_HVT U125 ( .A1(n579), .A3(n287), .A2(n339), .A4(n375), .S0(n289), 
        .S1(n325), .Y(n475) );
  MUX41X1_HVT U131 ( .A1(n470), .A3(n472), .A2(n471), .A4(n473), .S0(n296), 
        .S1(n325), .Y(n469) );
  MUX41X1_HVT U132 ( .A1(n469), .A3(n482), .A2(n474), .A4(n487), .S0(in[6]), 
        .S1(n304), .Y(out[3]) );
  MUX41X1_HVT U135 ( .A1(n376), .A3(n381), .A2(n595), .A4(n575), .S0(n290), 
        .S1(n325), .Y(n466) );
  AND2X1_HVT U140 ( .A1(n308), .A2(n210), .Y(n461) );
  OA21X1_HVT U144 ( .A1(n333), .A2(n327), .A3(n571), .Y(n457) );
  NAND2X0_HVT U146 ( .A1(n320), .A2(n315), .Y(n530) );
  MUX41X1_HVT U147 ( .A1(n377), .A3(n530), .A2(n366), .A4(n557), .S0(n290), 
        .S1(n325), .Y(n455) );
  MUX41X1_HVT U148 ( .A1(n455), .A3(n459), .A2(n456), .A4(n460), .S0(n304), 
        .S1(n295), .Y(n454) );
  OA21X1_HVT U151 ( .A1(n562), .A2(n327), .A3(n451), .Y(n452) );
  MUX41X1_HVT U153 ( .A1(n492), .A3(n283), .A2(n311), .A4(n332), .S0(n289), 
        .S1(n216), .Y(n449) );
  AND2X1_HVT U154 ( .A1(n326), .A2(n306), .Y(n448) );
  NAND2X0_HVT U158 ( .A1(n320), .A2(n383), .Y(n444) );
  MUX41X1_HVT U159 ( .A1(n245), .A3(n300), .A2(n444), .A4(n338), .S0(n290), 
        .S1(n216), .Y(n443) );
  MUX41X1_HVT U160 ( .A1(n443), .A3(n449), .A2(n445), .A4(n450), .S0(n305), 
        .S1(n295), .Y(n442) );
  AND2X1_HVT U162 ( .A1(n594), .A2(n530), .Y(n440) );
  MUX41X1_HVT U163 ( .A1(n344), .A3(n440), .A2(n281), .A4(n441), .S0(n323), 
        .S1(n216), .Y(n439) );
  MUX41X1_HVT U165 ( .A1(n579), .A3(n352), .A2(n557), .A4(n438), .S0(n325), 
        .S1(n323), .Y(n437) );
  NAND2X0_HVT U166 ( .A1(n314), .A2(n547), .Y(n436) );
  NAND2X0_HVT U167 ( .A1(n384), .A2(n210), .Y(n435) );
  MUX41X1_HVT U168 ( .A1(n369), .A3(n308), .A2(n435), .A4(n436), .S0(n323), 
        .S1(n264), .Y(n434) );
  OA21X1_HVT U170 ( .A1(n285), .A2(n327), .A3(n571), .Y(n432) );
  NAND2X0_HVT U174 ( .A1(n316), .A2(n594), .Y(n587) );
  MUX41X1_HVT U176 ( .A1(n303), .A3(n429), .A2(n374), .A4(n587), .S0(n325), 
        .S1(n253), .Y(n428) );
  NAND2X0_HVT U177 ( .A1(n319), .A2(n303), .Y(n427) );
  MUX41X1_HVT U178 ( .A1(n583), .A3(n427), .A2(n378), .A4(n564), .S0(n290), 
        .S1(n324), .Y(n426) );
  MUX41X1_HVT U179 ( .A1(n574), .A3(n379), .A2(n334), .A4(n378), .S0(n291), 
        .S1(n324), .Y(n425) );
  MUX41X1_HVT U180 ( .A1(n337), .A3(n592), .A2(n588), .A4(n279), .S0(n297), 
        .S1(n323), .Y(n424) );
  MUX41X1_HVT U181 ( .A1(n424), .A3(n426), .A2(n425), .A4(n428), .S0(n305), 
        .S1(n295), .Y(n423) );
  MUX41X1_HVT U186 ( .A1(n282), .A3(n563), .A2(n530), .A4(n557), .S0(n291), 
        .S1(n324), .Y(n418) );
  MUX41X1_HVT U189 ( .A1(n416), .A3(n587), .A2(n417), .A4(n365), .S0(n297), 
        .S1(n253), .Y(n415) );
  MUX41X1_HVT U195 ( .A1(n594), .A3(n370), .A2(n314), .A4(n565), .S0(n253), 
        .S1(n264), .Y(n410) );
  AO21X1_HVT U197 ( .A1(n284), .A2(n298), .A3(n367), .Y(n408) );
  MUX41X1_HVT U199 ( .A1(n407), .A3(n411), .A2(n410), .A4(n412), .S0(n304), 
        .S1(n295), .Y(n406) );
  OA21X1_HVT U201 ( .A1(n593), .A2(n327), .A3(n358), .Y(n404) );
  MUX41X1_HVT U203 ( .A1(n566), .A3(n360), .A2(n589), .A4(n570), .S0(n323), 
        .S1(n324), .Y(n402) );
  MUX41X1_HVT U204 ( .A1(n548), .A3(n588), .A2(n355), .A4(n578), .S0(n323), 
        .S1(n324), .Y(n401) );
  MUX41X1_HVT U205 ( .A1(n211), .A3(n598), .A2(n379), .A4(n275), .S0(n290), 
        .S1(n324), .Y(n400) );
  NAND2X0_HVT U208 ( .A1(n319), .A2(n309), .Y(n491) );
  NAND2X0_HVT U212 ( .A1(n317), .A2(n307), .Y(n547) );
  NAND2X0_HVT U214 ( .A1(n594), .A2(n322), .Y(n398) );
  NAND2X0_HVT U215 ( .A1(n491), .A2(n308), .Y(n397) );
  AO21X1_HVT U216 ( .A1(n210), .A2(n381), .A3(n327), .Y(n501) );
  NAND2X0_HVT U218 ( .A1(n381), .A2(n320), .Y(n451) );
  NAND2X0_HVT U220 ( .A1(n298), .A2(n398), .Y(n522) );
  INVX2_HVT U1 ( .A(n256), .Y(n323) );
  INVX0_HVT U2 ( .A(n299), .Y(n23) );
  MUX21X2_HVT U3 ( .A1(n372), .A2(n381), .S0(n298), .Y(n453) );
  NAND2X0_HVT U6 ( .A1(n279), .A2(n26), .Y(n45) );
  NAND2X0_HVT U7 ( .A1(n584), .A2(n270), .Y(n48) );
  NAND2X0_HVT U8 ( .A1(n45), .A2(n48), .Y(n405) );
  IBUFFX2_HVT U9 ( .A(n270), .Y(n26) );
  INVX0_HVT U10 ( .A(n297), .Y(n270) );
  MUX21X1_HVT U11 ( .A1(n404), .A2(n405), .S0(n291), .Y(n403) );
  INVX1_HVT U12 ( .A(n588), .Y(n273) );
  MUX41X1_HVT U14 ( .A1(n566), .A3(n377), .A2(n569), .A4(n280), .S0(n50), .S1(
        n328), .Y(n465) );
  IBUFFX16_HVT U16 ( .A(n289), .Y(n50) );
  IBUFFX2_HVT U17 ( .A(n328), .Y(n325) );
  INVX1_HVT U18 ( .A(n272), .Y(n486) );
  INVX1_HVT U19 ( .A(n321), .Y(n87) );
  INVX1_HVT U20 ( .A(n321), .Y(n121) );
  INVX1_HVT U22 ( .A(n321), .Y(n317) );
  INVX0_HVT U23 ( .A(n321), .Y(n319) );
  INVX1_HVT U25 ( .A(n321), .Y(n316) );
  INVX1_HVT U26 ( .A(in[1]), .Y(n321) );
  INVX1_HVT U27 ( .A(in[1]), .Y(n210) );
  MUX41X1_HVT U28 ( .A1(n467), .A3(n465), .A2(n466), .A4(n463), .S0(n259), 
        .S1(n240), .Y(n462) );
  INVX1_HVT U29 ( .A(n385), .Y(n211) );
  INVX2_HVT U30 ( .A(in[4]), .Y(n385) );
  MUX21X1_HVT U31 ( .A1(n23), .A2(n384), .S0(n210), .Y(n581) );
  INVX0_HVT U32 ( .A(n382), .Y(n212) );
  INVX0_HVT U34 ( .A(in[3]), .Y(n213) );
  NBUFFX4_HVT U36 ( .A(in[7]), .Y(n216) );
  INVX1_HVT U37 ( .A(in[7]), .Y(n327) );
  MUX21X1_HVT U38 ( .A1(n302), .A2(n299), .S0(n322), .Y(n413) );
  MUX41X1_HVT U39 ( .A1(n413), .A3(n555), .A2(n567), .A4(n560), .S0(n217), 
        .S1(n218), .Y(n412) );
  IBUFFX16_HVT U40 ( .A(n290), .Y(n217) );
  IBUFFX16_HVT U41 ( .A(n324), .Y(n218) );
  MUX41X1_HVT U43 ( .A1(n308), .A3(n364), .A2(n300), .A4(n348), .S0(n219), 
        .S1(n327), .Y(n459) );
  IBUFFX16_HVT U44 ( .A(n289), .Y(n219) );
  NBUFFX2_HVT U45 ( .A(n318), .Y(n231) );
  NBUFFX2_HVT U46 ( .A(n318), .Y(n232) );
  IBUFFX2_HVT U47 ( .A(n322), .Y(n318) );
  NAND2X0_HVT U48 ( .A1(n542), .A2(n253), .Y(n254) );
  INVX0_HVT U49 ( .A(n319), .Y(n242) );
  INVX0_HVT U50 ( .A(n249), .Y(n519) );
  XNOR2X1_HVT U52 ( .A1(n327), .A2(n575), .Y(n267) );
  INVX0_HVT U54 ( .A(n317), .Y(n252) );
  NBUFFX2_HVT U55 ( .A(n385), .Y(n303) );
  INVX0_HVT U60 ( .A(n578), .Y(n348) );
  INVX1_HVT U64 ( .A(n304), .Y(n259) );
  INVX1_HVT U65 ( .A(n306), .Y(n382) );
  XNOR2X1_HVT U67 ( .A1(n276), .A2(n328), .Y(n233) );
  MUX21X1_HVT U69 ( .A1(n382), .A2(n300), .S0(n210), .Y(n584) );
  INVX1_HVT U70 ( .A(n584), .Y(n250) );
  NBUFFX2_HVT U71 ( .A(n269), .Y(n301) );
  NBUFFX2_HVT U72 ( .A(in[5]), .Y(n296) );
  INVX1_HVT U76 ( .A(n295), .Y(n240) );
  INVX1_HVT U79 ( .A(in[6]), .Y(n271) );
  INVX1_HVT U81 ( .A(n271), .Y(n268) );
  INVX1_HVT U82 ( .A(n289), .Y(n276) );
  INVX1_HVT U83 ( .A(n289), .Y(n238) );
  NBUFFX2_HVT U84 ( .A(in[2]), .Y(n289) );
  INVX1_HVT U88 ( .A(n291), .Y(n256) );
  INVX0_HVT U89 ( .A(n268), .Y(n246) );
  IBUFFX2_HVT U90 ( .A(n568), .Y(n355) );
  MUX21X1_HVT U91 ( .A1(n340), .A2(n598), .S0(n239), .Y(n234) );
  MUX21X1_HVT U92 ( .A1(n567), .A2(n351), .S0(n239), .Y(n235) );
  MUX21X1_HVT U94 ( .A1(n234), .A2(n235), .S0(n216), .Y(n498) );
  NAND2X0_HVT U95 ( .A1(n495), .A2(n246), .Y(n236) );
  NAND2X0_HVT U98 ( .A1(n505), .A2(in[6]), .Y(n237) );
  NAND2X0_HVT U99 ( .A1(n236), .A2(n237), .Y(out[2]) );
  NAND2X0_HVT U100 ( .A1(n317), .A2(n312), .Y(n598) );
  IBUFFX2_HVT U102 ( .A(n288), .Y(n239) );
  MUX21X2_HVT U103 ( .A1(n492), .A2(n571), .S0(n238), .Y(n490) );
  NAND2X0_HVT U104 ( .A1(n483), .A2(n240), .Y(n257) );
  INVX1_HVT U107 ( .A(n269), .Y(n594) );
  INVX1_HVT U108 ( .A(n392), .Y(n372) );
  MUX41X1_HVT U111 ( .A1(n439), .A3(n434), .A2(n437), .A4(n431), .S0(n259), 
        .S1(n240), .Y(n430) );
  MUX21X2_HVT U112 ( .A1(n516), .A2(n525), .S0(n268), .Y(out[1]) );
  MUX21X2_HVT U113 ( .A1(n586), .A2(n275), .S0(n238), .Y(n504) );
  MUX21X2_HVT U115 ( .A1(n353), .A2(n468), .S0(n292), .Y(n467) );
  MUX21X2_HVT U116 ( .A1(n452), .A2(n453), .S0(n293), .Y(n450) );
  MUX21X1_HVT U117 ( .A1(n359), .A2(n578), .S0(n270), .Y(n464) );
  OA21X1_HVT U118 ( .A1(n568), .A2(n328), .A3(n348), .Y(n420) );
  NBUFFX2_HVT U119 ( .A(n385), .Y(n302) );
  MUX21X1_HVT U120 ( .A1(n311), .A2(n269), .S0(n242), .Y(n241) );
  MUX21X1_HVT U121 ( .A1(n560), .A2(n557), .S0(n238), .Y(n243) );
  MUX21X1_HVT U122 ( .A1(n515), .A2(n368), .S0(n238), .Y(n244) );
  MUX21X1_HVT U124 ( .A1(n243), .A2(n244), .S0(n216), .Y(n514) );
  MUX21X2_HVT U126 ( .A1(n430), .A2(n442), .S0(in[6]), .Y(out[5]) );
  INVX1_HVT U127 ( .A(n534), .Y(n266) );
  INVX1_HVT U128 ( .A(n394), .Y(n370) );
  INVX0_HVT U129 ( .A(n273), .Y(n245) );
  NAND2X0_HVT U130 ( .A1(n399), .A2(n246), .Y(n247) );
  NAND2X0_HVT U133 ( .A1(n406), .A2(n268), .Y(n248) );
  NAND2X0_HVT U134 ( .A1(n247), .A2(n248), .Y(out[7]) );
  MUX41X1_HVT U136 ( .A1(n251), .A3(n250), .A2(n269), .A4(n578), .S0(n276), 
        .S1(n327), .Y(n249) );
  NAND2X0_HVT U137 ( .A1(n316), .A2(n211), .Y(n251) );
  XOR2X1_HVT U138 ( .A1(n269), .A2(n252), .Y(n557) );
  NAND2X0_HVT U139 ( .A1(n540), .A2(n256), .Y(n255) );
  NAND2X0_HVT U141 ( .A1(n254), .A2(n255), .Y(n539) );
  INVX1_HVT U142 ( .A(n256), .Y(n253) );
  NAND2X0_HVT U143 ( .A1(n486), .A2(n296), .Y(n258) );
  NAND2X0_HVT U145 ( .A1(n257), .A2(n258), .Y(n482) );
  INVX1_HVT U149 ( .A(n311), .Y(n384) );
  INVX0_HVT U150 ( .A(n265), .Y(n533) );
  MUX21X2_HVT U152 ( .A1(n384), .A2(n383), .S0(n316), .Y(n575) );
  MUX41X1_HVT U155 ( .A1(n549), .A3(n539), .A2(n543), .A4(n535), .S0(n271), 
        .S1(n259), .Y(out[0]) );
  MUX21X2_HVT U156 ( .A1(n544), .A2(n546), .S0(n291), .Y(n543) );
  NAND2X0_HVT U157 ( .A1(n550), .A2(n256), .Y(n260) );
  NAND2X0_HVT U161 ( .A1(n554), .A2(n292), .Y(n261) );
  NAND2X0_HVT U164 ( .A1(n260), .A2(n261), .Y(n549) );
  MUX41X1_HVT U169 ( .A1(n354), .A3(n461), .A2(n358), .A4(n274), .S0(n238), 
        .S1(n327), .Y(n460) );
  MUX41X1_HVT U171 ( .A1(n586), .A3(n330), .A2(n347), .A4(n558), .S0(n276), 
        .S1(n327), .Y(n520) );
  NAND2X0_HVT U172 ( .A1(n476), .A2(in[5]), .Y(n262) );
  NAND2X0_HVT U173 ( .A1(n475), .A2(n240), .Y(n263) );
  NAND2X0_HVT U175 ( .A1(n262), .A2(n263), .Y(n474) );
  MUX41X1_HVT U182 ( .A1(n507), .A3(n514), .A2(n506), .A4(n509), .S0(n305), 
        .S1(n240), .Y(n505) );
  INVX2_HVT U183 ( .A(in[7]), .Y(n328) );
  NBUFFX2_HVT U184 ( .A(n324), .Y(n264) );
  MUX41X1_HVT U185 ( .A1(n400), .A3(n401), .A2(n402), .A4(n403), .S0(in[5]), 
        .S1(n305), .Y(n399) );
  IBUFFX2_HVT U187 ( .A(n328), .Y(n324) );
  MUX21X1_HVT U188 ( .A1(n266), .A2(n267), .S0(n238), .Y(n265) );
  MUX41X1_HVT U190 ( .A1(n418), .A3(n415), .A2(n422), .A4(n419), .S0(n240), 
        .S1(in[0]), .Y(n414) );
  MUX21X2_HVT U191 ( .A1(n414), .A2(n423), .S0(in[6]), .Y(out[6]) );
  XNOR2X2_HVT U192 ( .A1(n385), .A2(n306), .Y(n269) );
  AND3X2_HVT U193 ( .A1(n292), .A2(n210), .A3(n211), .Y(n472) );
  AO21X2_HVT U194 ( .A1(n293), .A2(n308), .A3(n594), .Y(n484) );
  MUX21X1_HVT U196 ( .A1(n313), .A2(n489), .S0(n278), .Y(n488) );
  INVX1_HVT U198 ( .A(n571), .Y(n275) );
  INVX1_HVT U200 ( .A(in[1]), .Y(n322) );
  MUX21X1_HVT U202 ( .A1(n23), .A2(n301), .S0(n322), .Y(n578) );
  MUX21X2_HVT U206 ( .A1(n597), .A2(n464), .S0(n276), .Y(n463) );
  MUX21X2_HVT U207 ( .A1(n421), .A2(n420), .S0(n276), .Y(n419) );
  INVX0_HVT U209 ( .A(n241), .Y(n274) );
  MUX21X2_HVT U210 ( .A1(n454), .A2(n462), .S0(in[6]), .Y(out[4]) );
  MUX41X1_HVT U211 ( .A1(n349), .A3(n361), .A2(n309), .A4(n359), .S0(n327), 
        .S1(n238), .Y(n422) );
  MUX41X1_HVT U213 ( .A1(n275), .A3(n274), .A2(n277), .A4(n273), .S0(n276), 
        .S1(n327), .Y(n272) );
  NAND2X0_HVT U217 ( .A1(n87), .A2(n300), .Y(n277) );
  MUX41X1_HVT U219 ( .A1(n307), .A3(n376), .A2(n575), .A4(n561), .S0(n270), 
        .S1(n238), .Y(n411) );
  MUX21X2_HVT U221 ( .A1(n504), .A2(n283), .S0(n233), .Y(n503) );
  XNOR2X1_HVT U222 ( .A1(n210), .A2(n276), .Y(n278) );
  INVX0_HVT U223 ( .A(n321), .Y(n320) );
  INVX0_HVT U224 ( .A(n328), .Y(n326) );
  INVX1_HVT U225 ( .A(n596), .Y(n380) );
  MUX21X1_HVT U226 ( .A1(n281), .A2(n250), .S0(n289), .Y(n471) );
  NBUFFX2_HVT U227 ( .A(n269), .Y(n300) );
  AND2X1_HVT U228 ( .A1(n301), .A2(n547), .Y(n279) );
  MUX21X1_HVT U229 ( .A1(n380), .A2(n383), .S0(n296), .Y(n551) );
  NBUFFX2_HVT U230 ( .A(n596), .Y(n309) );
  NBUFFX2_HVT U231 ( .A(n596), .Y(n310) );
  MUX21X1_HVT U232 ( .A1(n340), .A2(n381), .S0(n296), .Y(n536) );
  AND2X1_HVT U233 ( .A1(n312), .A2(n530), .Y(n280) );
  MUX21X1_HVT U234 ( .A1(n301), .A2(n383), .S0(n320), .Y(n593) );
  MUX21X1_HVT U235 ( .A1(n480), .A2(n479), .S0(n326), .Y(n476) );
  MUX21X1_HVT U236 ( .A1(n312), .A2(n300), .S0(n231), .Y(n561) );
  MUX21X1_HVT U237 ( .A1(n300), .A2(n303), .S0(n320), .Y(n500) );
  MUX21X1_HVT U238 ( .A1(n380), .A2(n384), .S0(n232), .Y(n429) );
  MUX21X1_HVT U239 ( .A1(n383), .A2(n269), .S0(n316), .Y(n441) );
  MUX21X1_HVT U240 ( .A1(n269), .A2(n380), .S0(n121), .Y(n508) );
  MUX21X1_HVT U241 ( .A1(n310), .A2(n594), .S0(n231), .Y(n565) );
  MUX21X1_HVT U242 ( .A1(n594), .A2(n381), .S0(n87), .Y(n389) );
  MUX21X1_HVT U243 ( .A1(n309), .A2(n308), .S0(n231), .Y(n515) );
  MUX21X1_HVT U244 ( .A1(n594), .A2(n303), .S0(n232), .Y(n527) );
  MUX21X1_HVT U245 ( .A1(n299), .A2(n594), .S0(n121), .Y(n392) );
  MUX21X1_HVT U246 ( .A1(n383), .A2(n380), .S0(n231), .Y(n564) );
  MUX21X1_HVT U247 ( .A1(n383), .A2(n382), .S0(n231), .Y(n568) );
  MUX21X1_HVT U248 ( .A1(n382), .A2(n384), .S0(n232), .Y(n562) );
  MUX21X1_HVT U249 ( .A1(n302), .A2(n380), .S0(n317), .Y(n573) );
  MUX21X1_HVT U250 ( .A1(n375), .A2(n308), .S0(n298), .Y(n468) );
  MUX21X1_HVT U251 ( .A1(n484), .A2(n485), .S0(n298), .Y(n483) );
  MUX21X1_HVT U252 ( .A1(n332), .A2(n355), .S0(n289), .Y(n485) );
  NAND2X0_HVT U253 ( .A1(n302), .A2(n299), .Y(n596) );
  MUX21X1_HVT U254 ( .A1(n380), .A2(n303), .S0(n121), .Y(n390) );
  NBUFFX2_HVT U255 ( .A(n599), .Y(n311) );
  INVX1_HVT U256 ( .A(n600), .Y(n383) );
  MUX21X1_HVT U257 ( .A1(n313), .A2(n307), .S0(n317), .Y(n586) );
  MUX21X1_HVT U258 ( .A1(n310), .A2(n315), .S0(n320), .Y(n510) );
  MUX21X1_HVT U259 ( .A1(n381), .A2(n380), .S0(n121), .Y(n582) );
  MUX21X1_HVT U260 ( .A1(n331), .A2(n481), .S0(n290), .Y(n480) );
  MUX21X1_HVT U261 ( .A1(n302), .A2(n382), .S0(n319), .Y(n481) );
  NBUFFX2_HVT U262 ( .A(n599), .Y(n312) );
  NBUFFX2_HVT U263 ( .A(n599), .Y(n313) );
  MUX21X1_HVT U264 ( .A1(n299), .A2(n315), .S0(n319), .Y(n416) );
  MUX21X1_HVT U265 ( .A1(n314), .A2(n312), .S0(n316), .Y(n417) );
  INVX1_HVT U266 ( .A(n591), .Y(n381) );
  MUX21X1_HVT U267 ( .A1(n382), .A2(n383), .S0(n317), .Y(n590) );
  XOR2X1_HVT U268 ( .A1(n311), .A2(n87), .Y(n555) );
  XOR2X1_HVT U269 ( .A1(n319), .A2(n381), .Y(n558) );
  MUX21X1_HVT U270 ( .A1(n311), .A2(n303), .S0(n316), .Y(n396) );
  XNOR2X1_HVT U271 ( .A1(n310), .A2(n320), .Y(n281) );
  AND2X1_HVT U272 ( .A1(n121), .A2(n384), .Y(n282) );
  MUX21X1_HVT U273 ( .A1(n315), .A2(n307), .S0(n231), .Y(n571) );
  MUX21X1_HVT U274 ( .A1(n309), .A2(n382), .S0(n317), .Y(n589) );
  MUX21X1_HVT U275 ( .A1(n311), .A2(n309), .S0(n121), .Y(n388) );
  AND2X1_HVT U276 ( .A1(n314), .A2(n491), .Y(n283) );
  XNOR2X1_HVT U277 ( .A1(n314), .A2(n121), .Y(n284) );
  MUX21X1_HVT U278 ( .A1(n307), .A2(n382), .S0(n320), .Y(n394) );
  MUX21X1_HVT U279 ( .A1(n308), .A2(n303), .S0(n232), .Y(n532) );
  MUX21X1_HVT U280 ( .A1(n308), .A2(n315), .S0(n292), .Y(n478) );
  XOR2X1_HVT U281 ( .A1(n303), .A2(n87), .Y(n576) );
  NBUFFX2_HVT U282 ( .A(n213), .Y(n299) );
  NBUFFX2_HVT U283 ( .A(n326), .Y(n297) );
  NBUFFX2_HVT U284 ( .A(n326), .Y(n298) );
  NBUFFX2_HVT U285 ( .A(in[2]), .Y(n290) );
  NBUFFX2_HVT U286 ( .A(in[5]), .Y(n295) );
  NBUFFX2_HVT U287 ( .A(n253), .Y(n292) );
  NBUFFX2_HVT U288 ( .A(n291), .Y(n293) );
  NBUFFX2_HVT U289 ( .A(in[2]), .Y(n291) );
  NBUFFX2_HVT U290 ( .A(in[5]), .Y(n294) );
  NBUFFX2_HVT U291 ( .A(n323), .Y(n288) );
  MUX21X1_HVT U292 ( .A1(n502), .A2(n353), .S0(n292), .Y(n499) );
  MUX21X1_HVT U293 ( .A1(n518), .A2(n23), .S0(n298), .Y(n421) );
  XOR2X1_HVT U294 ( .A1(n320), .A2(n306), .Y(n556) );
  MUX21X1_HVT U295 ( .A1(n307), .A2(n301), .S0(n232), .Y(n497) );
  MUX21X1_HVT U296 ( .A1(n524), .A2(n523), .S0(n293), .Y(n521) );
  MUX21X1_HVT U297 ( .A1(n580), .A2(n308), .S0(n298), .Y(n524) );
  MUX21X1_HVT U298 ( .A1(n381), .A2(n384), .S0(n87), .Y(n438) );
  MUX21X1_HVT U299 ( .A1(n433), .A2(n432), .S0(n292), .Y(n431) );
  MUX21X1_HVT U300 ( .A1(n308), .A2(n370), .S0(n326), .Y(n433) );
  AND2X1_HVT U301 ( .A1(n301), .A2(n210), .Y(n285) );
  MUX21X1_HVT U302 ( .A1(n306), .A2(n380), .S0(n232), .Y(n563) );
  MUX21X1_HVT U303 ( .A1(n383), .A2(n370), .S0(n326), .Y(n534) );
  MUX21X1_HVT U304 ( .A1(n458), .A2(n457), .S0(n292), .Y(n456) );
  MUX21X1_HVT U305 ( .A1(n573), .A2(n335), .S0(n326), .Y(n458) );
  NAND2X0_HVT U306 ( .A1(n306), .A2(n302), .Y(n599) );
  MUX21X1_HVT U307 ( .A1(n356), .A2(n598), .S0(n290), .Y(n494) );
  MUX21X1_HVT U308 ( .A1(n446), .A2(n447), .S0(n293), .Y(n445) );
  MUX21X1_HVT U309 ( .A1(n448), .A2(n313), .S0(n286), .Y(n447) );
  MUX21X1_HVT U310 ( .A1(n564), .A2(n373), .S0(n297), .Y(n446) );
  MUX21X1_HVT U311 ( .A1(n583), .A2(n354), .S0(n290), .Y(n470) );
  MUX21X1_HVT U312 ( .A1(n552), .A2(n553), .S0(n297), .Y(n550) );
  MUX21X1_HVT U313 ( .A1(n212), .A2(n567), .S0(n296), .Y(n553) );
  XOR2X1_HVT U314 ( .A1(n87), .A2(n295), .Y(n559) );
  MUX21X1_HVT U315 ( .A1(n598), .A2(n322), .S0(n291), .Y(n477) );
  MUX21X1_HVT U316 ( .A1(n23), .A2(n381), .S0(n316), .Y(n393) );
  MUX21X1_HVT U317 ( .A1(n572), .A2(n397), .S0(n297), .Y(n391) );
  MUX21X1_HVT U318 ( .A1(n310), .A2(n23), .S0(n121), .Y(n592) );
  MUX21X1_HVT U319 ( .A1(n342), .A2(n322), .S0(n296), .Y(n538) );
  NBUFFX2_HVT U320 ( .A(n591), .Y(n307) );
  MUX21X1_HVT U321 ( .A1(n350), .A2(n572), .S0(n290), .Y(n473) );
  MUX21X1_HVT U322 ( .A1(n362), .A2(n378), .S0(n298), .Y(n409) );
  MUX21X1_HVT U323 ( .A1(n313), .A2(n513), .S0(n286), .Y(n512) );
  MUX21X1_HVT U324 ( .A1(n23), .A2(n302), .S0(n326), .Y(n513) );
  NBUFFX2_HVT U325 ( .A(n600), .Y(n315) );
  NBUFFX2_HVT U326 ( .A(n591), .Y(n308) );
  NBUFFX2_HVT U327 ( .A(n600), .Y(n314) );
  XNOR2X1_HVT U328 ( .A1(n328), .A2(n316), .Y(n286) );
  AND2X1_HVT U329 ( .A1(n382), .A2(n210), .Y(n287) );
  MUX21X1_HVT U330 ( .A1(n409), .A2(n408), .S0(n291), .Y(n407) );
  MUX21X1_HVT U331 ( .A1(n511), .A2(n512), .S0(n293), .Y(n509) );
  MUX21X1_HVT U332 ( .A1(n380), .A2(n211), .S0(n232), .Y(n570) );
  NAND2X0_HVT U333 ( .A1(n306), .A2(in[4]), .Y(n600) );
  MUX21X1_HVT U334 ( .A1(n211), .A2(n594), .S0(n319), .Y(n395) );
  MUX21X1_HVT U335 ( .A1(n211), .A2(n383), .S0(n231), .Y(n566) );
  MUX21X1_HVT U336 ( .A1(n211), .A2(n381), .S0(n319), .Y(n583) );
  NAND2X0_HVT U337 ( .A1(in[4]), .A2(n299), .Y(n591) );
  MUX21X1_HVT U338 ( .A1(n211), .A2(n313), .S0(n317), .Y(n580) );
  MUX21X1_HVT U339 ( .A1(n315), .A2(n211), .S0(n316), .Y(n574) );
  MUX21X1_HVT U340 ( .A1(n23), .A2(n211), .S0(n289), .Y(n489) );
  MUX21X1_HVT U341 ( .A1(n211), .A2(n307), .S0(n87), .Y(n387) );
  MUX21X1_HVT U342 ( .A1(n211), .A2(n314), .S0(n232), .Y(n386) );
  MUX21X1_HVT U343 ( .A1(n382), .A2(n211), .S0(n87), .Y(n572) );
  NBUFFX2_HVT U344 ( .A(in[3]), .Y(n306) );
  NBUFFX2_HVT U345 ( .A(in[0]), .Y(n305) );
  NBUFFX2_HVT U346 ( .A(in[0]), .Y(n304) );
  INVX0_HVT U347 ( .A(n579), .Y(n329) );
  INVX0_HVT U348 ( .A(n577), .Y(n330) );
  INVX0_HVT U349 ( .A(n569), .Y(n331) );
  INVX0_HVT U350 ( .A(n567), .Y(n332) );
  INVX0_HVT U351 ( .A(n435), .Y(n333) );
  INVX0_HVT U352 ( .A(n398), .Y(n334) );
  INVX0_HVT U353 ( .A(n598), .Y(n335) );
  INVX0_HVT U354 ( .A(n585), .Y(n336) );
  INVX0_HVT U355 ( .A(n597), .Y(n337) );
  INVX0_HVT U356 ( .A(n595), .Y(n338) );
  INVX0_HVT U357 ( .A(n593), .Y(n339) );
  INVX0_HVT U358 ( .A(n592), .Y(n340) );
  INVX0_HVT U359 ( .A(n590), .Y(n341) );
  INVX0_HVT U360 ( .A(n589), .Y(n342) );
  INVX0_HVT U361 ( .A(n586), .Y(n343) );
  INVX0_HVT U362 ( .A(n583), .Y(n344) );
  INVX0_HVT U363 ( .A(n582), .Y(n345) );
  INVX0_HVT U364 ( .A(n581), .Y(n346) );
  INVX0_HVT U365 ( .A(n580), .Y(n347) );
  INVX0_HVT U366 ( .A(n576), .Y(n349) );
  INVX0_HVT U367 ( .A(n574), .Y(n350) );
  INVX0_HVT U368 ( .A(n573), .Y(n351) );
  INVX0_HVT U369 ( .A(n572), .Y(n352) );
  INVX0_HVT U370 ( .A(n391), .Y(n353) );
  INVX0_HVT U371 ( .A(n570), .Y(n354) );
  INVX0_HVT U372 ( .A(n566), .Y(n356) );
  INVX0_HVT U373 ( .A(n565), .Y(n357) );
  INVX0_HVT U374 ( .A(n564), .Y(n358) );
  INVX0_HVT U375 ( .A(n563), .Y(n359) );
  INVX0_HVT U376 ( .A(n562), .Y(n360) );
  INVX0_HVT U377 ( .A(n561), .Y(n361) );
  INVX0_HVT U378 ( .A(n560), .Y(n362) );
  INVX0_HVT U379 ( .A(n530), .Y(n363) );
  INVX0_HVT U380 ( .A(n491), .Y(n364) );
  INVX0_HVT U381 ( .A(n397), .Y(n365) );
  INVX0_HVT U382 ( .A(n547), .Y(n366) );
  INVX0_HVT U383 ( .A(n451), .Y(n367) );
  INVX0_HVT U384 ( .A(n396), .Y(n368) );
  INVX0_HVT U385 ( .A(n395), .Y(n369) );
  INVX0_HVT U386 ( .A(n393), .Y(n371) );
  INVX0_HVT U387 ( .A(n510), .Y(n373) );
  INVX0_HVT U388 ( .A(n500), .Y(n374) );
  INVX0_HVT U389 ( .A(n390), .Y(n375) );
  INVX0_HVT U390 ( .A(n389), .Y(n376) );
  INVX0_HVT U391 ( .A(n388), .Y(n377) );
  INVX0_HVT U392 ( .A(n387), .Y(n378) );
  INVX0_HVT U393 ( .A(n386), .Y(n379) );
endmodule

