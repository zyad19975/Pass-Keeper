
module Get_key ( clk, rest, local_key, rount_no, key_round, done );
  input [127:0] local_key;
  input [3:0] rount_no;
  output [127:0] key_round;
  input clk, rest;
  output done;
  wire   \keys[0][127] , \keys[0][126] , \keys[0][125] , \keys[0][124] ,
         \keys[0][123] , \keys[0][122] , \keys[0][121] , \keys[0][120] ,
         \keys[0][119] , \keys[0][118] , \keys[0][117] , \keys[0][116] ,
         \keys[0][115] , \keys[0][114] , \keys[0][113] , \keys[0][112] ,
         \keys[0][111] , \keys[0][110] , \keys[0][109] , \keys[0][108] ,
         \keys[0][107] , \keys[0][106] , \keys[0][105] , \keys[0][104] ,
         \keys[0][103] , \keys[0][102] , \keys[0][101] , \keys[0][100] ,
         \keys[0][99] , \keys[0][98] , \keys[0][97] , \keys[0][96] ,
         \keys[0][95] , \keys[0][94] , \keys[0][93] , \keys[0][92] ,
         \keys[0][91] , \keys[0][90] , \keys[0][89] , \keys[0][88] ,
         \keys[0][87] , \keys[0][86] , \keys[0][85] , \keys[0][84] ,
         \keys[0][83] , \keys[0][82] , \keys[0][81] , \keys[0][80] ,
         \keys[0][79] , \keys[0][78] , \keys[0][77] , \keys[0][76] ,
         \keys[0][75] , \keys[0][74] , \keys[0][73] , \keys[0][72] ,
         \keys[0][71] , \keys[0][70] , \keys[0][69] , \keys[0][68] ,
         \keys[0][67] , \keys[0][66] , \keys[0][65] , \keys[0][64] ,
         \keys[0][63] , \keys[0][62] , \keys[0][61] , \keys[0][60] ,
         \keys[0][59] , \keys[0][58] , \keys[0][57] , \keys[0][56] ,
         \keys[0][55] , \keys[0][54] , \keys[0][53] , \keys[0][52] ,
         \keys[0][51] , \keys[0][50] , \keys[0][49] , \keys[0][48] ,
         \keys[0][47] , \keys[0][46] , \keys[0][45] , \keys[0][44] ,
         \keys[0][43] , \keys[0][42] , \keys[0][41] , \keys[0][40] ,
         \keys[0][39] , \keys[0][38] , \keys[0][37] , \keys[0][36] ,
         \keys[0][35] , \keys[0][34] , \keys[0][33] , \keys[0][32] ,
         \keys[0][31] , \keys[0][30] , \keys[0][29] , \keys[0][28] ,
         \keys[0][27] , \keys[0][26] , \keys[0][25] , \keys[0][24] ,
         \keys[0][23] , \keys[0][22] , \keys[0][21] , \keys[0][20] ,
         \keys[0][19] , \keys[0][18] , \keys[0][17] , \keys[0][16] ,
         \keys[0][15] , \keys[0][14] , \keys[0][13] , \keys[0][12] ,
         \keys[0][11] , \keys[0][10] , \keys[0][9] , \keys[0][8] ,
         \keys[0][7] , \keys[0][6] , \keys[0][5] , \keys[0][4] , \keys[0][3] ,
         \keys[0][2] , \keys[0][1] , \keys[0][0] , \keys[1][127] ,
         \keys[1][126] , \keys[1][125] , \keys[1][124] , \keys[1][123] ,
         \keys[1][122] , \keys[1][121] , \keys[1][120] , \keys[1][119] ,
         \keys[1][118] , \keys[1][117] , \keys[1][116] , \keys[1][115] ,
         \keys[1][114] , \keys[1][113] , \keys[1][112] , \keys[1][111] ,
         \keys[1][110] , \keys[1][109] , \keys[1][108] , \keys[1][107] ,
         \keys[1][106] , \keys[1][105] , \keys[1][104] , \keys[1][103] ,
         \keys[1][102] , \keys[1][101] , \keys[1][100] , \keys[1][99] ,
         \keys[1][98] , \keys[1][97] , \keys[1][96] , \keys[1][95] ,
         \keys[1][94] , \keys[1][93] , \keys[1][92] , \keys[1][91] ,
         \keys[1][90] , \keys[1][89] , \keys[1][88] , \keys[1][87] ,
         \keys[1][86] , \keys[1][85] , \keys[1][84] , \keys[1][83] ,
         \keys[1][82] , \keys[1][81] , \keys[1][80] , \keys[1][79] ,
         \keys[1][78] , \keys[1][77] , \keys[1][76] , \keys[1][75] ,
         \keys[1][74] , \keys[1][73] , \keys[1][72] , \keys[1][71] ,
         \keys[1][70] , \keys[1][69] , \keys[1][68] , \keys[1][67] ,
         \keys[1][66] , \keys[1][65] , \keys[1][64] , \keys[1][63] ,
         \keys[1][62] , \keys[1][61] , \keys[1][60] , \keys[1][59] ,
         \keys[1][58] , \keys[1][57] , \keys[1][56] , \keys[1][55] ,
         \keys[1][54] , \keys[1][53] , \keys[1][52] , \keys[1][51] ,
         \keys[1][50] , \keys[1][49] , \keys[1][48] , \keys[1][47] ,
         \keys[1][46] , \keys[1][45] , \keys[1][44] , \keys[1][42] ,
         \keys[1][41] , \keys[1][40] , \keys[1][39] , \keys[1][38] ,
         \keys[1][37] , \keys[1][36] , \keys[1][35] , \keys[1][34] ,
         \keys[1][33] , \keys[1][32] , \keys[1][31] , \keys[1][30] ,
         \keys[1][29] , \keys[1][28] , \keys[1][27] , \keys[1][26] ,
         \keys[1][25] , \keys[1][24] , \keys[1][23] , \keys[1][22] ,
         \keys[1][21] , \keys[1][20] , \keys[1][19] , \keys[1][18] ,
         \keys[1][17] , \keys[1][16] , \keys[1][15] , \keys[1][14] ,
         \keys[1][13] , \keys[1][12] , \keys[1][11] , \keys[1][10] ,
         \keys[1][9] , \keys[1][8] , \keys[1][7] , \keys[1][6] , \keys[1][5] ,
         \keys[1][4] , \keys[1][3] , \keys[1][2] , \keys[1][1] , \keys[1][0] ,
         \keys[2][127] , \keys[2][126] , \keys[2][125] , \keys[2][124] ,
         \keys[2][123] , \keys[2][122] , \keys[2][121] , \keys[2][120] ,
         \keys[2][119] , \keys[2][118] , \keys[2][117] , \keys[2][116] ,
         \keys[2][115] , \keys[2][114] , \keys[2][113] , \keys[2][112] ,
         \keys[2][111] , \keys[2][110] , \keys[2][109] , \keys[2][108] ,
         \keys[2][107] , \keys[2][106] , \keys[2][105] , \keys[2][104] ,
         \keys[2][103] , \keys[2][102] , \keys[2][101] , \keys[2][100] ,
         \keys[2][99] , \keys[2][98] , \keys[2][97] , \keys[2][96] ,
         \keys[2][95] , \keys[2][94] , \keys[2][93] , \keys[2][92] ,
         \keys[2][91] , \keys[2][90] , \keys[2][89] , \keys[2][88] ,
         \keys[2][87] , \keys[2][86] , \keys[2][85] , \keys[2][84] ,
         \keys[2][83] , \keys[2][82] , \keys[2][81] , \keys[2][80] ,
         \keys[2][79] , \keys[2][78] , \keys[2][77] , \keys[2][76] ,
         \keys[2][75] , \keys[2][74] , \keys[2][73] , \keys[2][72] ,
         \keys[2][71] , \keys[2][70] , \keys[2][69] , \keys[2][68] ,
         \keys[2][67] , \keys[2][66] , \keys[2][65] , \keys[2][64] ,
         \keys[2][63] , \keys[2][62] , \keys[2][61] , \keys[2][60] ,
         \keys[2][59] , \keys[2][58] , \keys[2][57] , \keys[2][56] ,
         \keys[2][55] , \keys[2][54] , \keys[2][53] , \keys[2][52] ,
         \keys[2][51] , \keys[2][50] , \keys[2][49] , \keys[2][48] ,
         \keys[2][46] , \keys[2][44] , \keys[2][43] , \keys[2][42] ,
         \keys[2][40] , \keys[2][39] , \keys[2][38] , \keys[2][37] ,
         \keys[2][36] , \keys[2][35] , \keys[2][34] , \keys[2][33] ,
         \keys[2][32] , \keys[2][31] , \keys[2][30] , \keys[2][29] ,
         \keys[2][28] , \keys[2][27] , \keys[2][26] , \keys[2][25] ,
         \keys[2][24] , \keys[2][23] , \keys[2][22] , \keys[2][21] ,
         \keys[2][20] , \keys[2][19] , \keys[2][18] , \keys[2][17] ,
         \keys[2][16] , \keys[2][15] , \keys[2][14] , \keys[2][13] ,
         \keys[2][12] , \keys[2][11] , \keys[2][10] , \keys[2][9] ,
         \keys[2][8] , \keys[2][7] , \keys[2][6] , \keys[2][5] , \keys[2][4] ,
         \keys[2][3] , \keys[2][2] , \keys[2][1] , \keys[2][0] ,
         \keys[3][127] , \keys[3][126] , \keys[3][125] , \keys[3][124] ,
         \keys[3][123] , \keys[3][122] , \keys[3][121] , \keys[3][120] ,
         \keys[3][119] , \keys[3][118] , \keys[3][117] , \keys[3][116] ,
         \keys[3][115] , \keys[3][114] , \keys[3][113] , \keys[3][112] ,
         \keys[3][111] , \keys[3][110] , \keys[3][109] , \keys[3][108] ,
         \keys[3][107] , \keys[3][106] , \keys[3][105] , \keys[3][104] ,
         \keys[3][103] , \keys[3][102] , \keys[3][101] , \keys[3][100] ,
         \keys[3][99] , \keys[3][98] , \keys[3][97] , \keys[3][96] ,
         \keys[3][95] , \keys[3][94] , \keys[3][93] , \keys[3][92] ,
         \keys[3][89] , \keys[3][88] , \keys[3][87] , \keys[3][86] ,
         \keys[3][85] , \keys[3][84] , \keys[3][83] , \keys[3][82] ,
         \keys[3][81] , \keys[3][80] , \keys[3][79] , \keys[3][78] ,
         \keys[3][77] , \keys[3][76] , \keys[3][75] , \keys[3][74] ,
         \keys[3][73] , \keys[3][72] , \keys[3][71] , \keys[3][70] ,
         \keys[3][69] , \keys[3][68] , \keys[3][67] , \keys[3][66] ,
         \keys[3][65] , \keys[3][64] , \keys[3][63] , \keys[3][62] ,
         \keys[3][61] , \keys[3][60] , \keys[3][59] , \keys[3][58] ,
         \keys[3][57] , \keys[3][56] , \keys[3][55] , \keys[3][54] ,
         \keys[3][53] , \keys[3][52] , \keys[3][51] , \keys[3][50] ,
         \keys[3][49] , \keys[3][48] , \keys[3][47] , \keys[3][46] ,
         \keys[3][45] , \keys[3][44] , \keys[3][43] , \keys[3][42] ,
         \keys[3][41] , \keys[3][40] , \keys[3][39] , \keys[3][38] ,
         \keys[3][37] , \keys[3][36] , \keys[3][35] , \keys[3][34] ,
         \keys[3][33] , \keys[3][32] , \keys[3][31] , \keys[3][30] ,
         \keys[3][29] , \keys[3][28] , \keys[3][27] , \keys[3][26] ,
         \keys[3][25] , \keys[3][24] , \keys[3][23] , \keys[3][22] ,
         \keys[3][21] , \keys[3][20] , \keys[3][19] , \keys[3][18] ,
         \keys[3][17] , \keys[3][16] , \keys[3][15] , \keys[3][14] ,
         \keys[3][13] , \keys[3][12] , \keys[3][11] , \keys[3][10] ,
         \keys[3][9] , \keys[3][8] , \keys[3][7] , \keys[3][6] , \keys[3][5] ,
         \keys[3][4] , \keys[3][3] , \keys[3][2] , \keys[3][1] , \keys[3][0] ,
         \keys[4][127] , \keys[4][126] , \keys[4][125] , \keys[4][124] ,
         \keys[4][123] , \keys[4][122] , \keys[4][121] , \keys[4][120] ,
         \keys[4][119] , \keys[4][118] , \keys[4][117] , \keys[4][116] ,
         \keys[4][115] , \keys[4][114] , \keys[4][113] , \keys[4][112] ,
         \keys[4][111] , \keys[4][110] , \keys[4][109] , \keys[4][108] ,
         \keys[4][107] , \keys[4][106] , \keys[4][105] , \keys[4][104] ,
         \keys[4][103] , \keys[4][102] , \keys[4][101] , \keys[4][100] ,
         \keys[4][99] , \keys[4][98] , \keys[4][97] , \keys[4][96] ,
         \keys[4][95] , \keys[4][94] , \keys[4][93] , \keys[4][92] ,
         \keys[4][91] , \keys[4][90] , \keys[4][89] , \keys[4][88] ,
         \keys[4][87] , \keys[4][86] , \keys[4][85] , \keys[4][84] ,
         \keys[4][83] , \keys[4][82] , \keys[4][81] , \keys[4][80] ,
         \keys[4][79] , \keys[4][78] , \keys[4][77] , \keys[4][76] ,
         \keys[4][73] , \keys[4][72] , \keys[4][71] , \keys[4][70] ,
         \keys[4][69] , \keys[4][68] , \keys[4][67] , \keys[4][66] ,
         \keys[4][65] , \keys[4][64] , \keys[4][63] , \keys[4][62] ,
         \keys[4][61] , \keys[4][60] , \keys[4][59] , \keys[4][58] ,
         \keys[4][57] , \keys[4][56] , \keys[4][55] , \keys[4][54] ,
         \keys[4][53] , \keys[4][52] , \keys[4][51] , \keys[4][50] ,
         \keys[4][49] , \keys[4][48] , \keys[4][47] , \keys[4][46] ,
         \keys[4][45] , \keys[4][43] , \keys[4][42] , \keys[4][41] ,
         \keys[4][40] , \keys[4][39] , \keys[4][38] , \keys[4][37] ,
         \keys[4][36] , \keys[4][35] , \keys[4][34] , \keys[4][33] ,
         \keys[4][32] , \keys[4][31] , \keys[4][30] , \keys[4][29] ,
         \keys[4][28] , \keys[4][27] , \keys[4][26] , \keys[4][25] ,
         \keys[4][24] , \keys[4][23] , \keys[4][22] , \keys[4][21] ,
         \keys[4][20] , \keys[4][19] , \keys[4][18] , \keys[4][17] ,
         \keys[4][16] , \keys[4][15] , \keys[4][14] , \keys[4][13] ,
         \keys[4][12] , \keys[4][11] , \keys[4][10] , \keys[4][9] ,
         \keys[4][8] , \keys[4][7] , \keys[4][6] , \keys[4][5] , \keys[4][4] ,
         \keys[4][3] , \keys[4][2] , \keys[4][1] , \keys[4][0] ,
         \keys[5][127] , \keys[5][126] , \keys[5][125] , \keys[5][124] ,
         \keys[5][123] , \keys[5][122] , \keys[5][121] , \keys[5][120] ,
         \keys[5][119] , \keys[5][118] , \keys[5][117] , \keys[5][116] ,
         \keys[5][115] , \keys[5][114] , \keys[5][113] , \keys[5][112] ,
         \keys[5][111] , \keys[5][110] , \keys[5][109] , \keys[5][108] ,
         \keys[5][107] , \keys[5][106] , \keys[5][105] , \keys[5][104] ,
         \keys[5][103] , \keys[5][102] , \keys[5][101] , \keys[5][100] ,
         \keys[5][99] , \keys[5][98] , \keys[5][97] , \keys[5][96] ,
         \keys[5][95] , \keys[5][94] , \keys[5][93] , \keys[5][92] ,
         \keys[5][91] , \keys[5][90] , \keys[5][89] , \keys[5][88] ,
         \keys[5][87] , \keys[5][86] , \keys[5][85] , \keys[5][84] ,
         \keys[5][83] , \keys[5][82] , \keys[5][81] , \keys[5][80] ,
         \keys[5][79] , \keys[5][78] , \keys[5][77] , \keys[5][76] ,
         \keys[5][75] , \keys[5][74] , \keys[5][73] , \keys[5][72] ,
         \keys[5][71] , \keys[5][70] , \keys[5][69] , \keys[5][68] ,
         \keys[5][67] , \keys[5][66] , \keys[5][65] , \keys[5][64] ,
         \keys[5][63] , \keys[5][62] , \keys[5][61] , \keys[5][60] ,
         \keys[5][59] , \keys[5][58] , \keys[5][57] , \keys[5][56] ,
         \keys[5][54] , \keys[5][53] , \keys[5][52] , \keys[5][51] ,
         \keys[5][50] , \keys[5][49] , \keys[5][48] , \keys[5][47] ,
         \keys[5][46] , \keys[5][45] , \keys[5][44] , \keys[5][43] ,
         \keys[5][42] , \keys[5][41] , \keys[5][40] , \keys[5][39] ,
         \keys[5][38] , \keys[5][37] , \keys[5][36] , \keys[5][35] ,
         \keys[5][34] , \keys[5][33] , \keys[5][32] , \keys[5][31] ,
         \keys[5][30] , \keys[5][29] , \keys[5][28] , \keys[5][27] ,
         \keys[5][26] , \keys[5][25] , \keys[5][24] , \keys[5][23] ,
         \keys[5][22] , \keys[5][21] , \keys[5][20] , \keys[5][19] ,
         \keys[5][18] , \keys[5][17] , \keys[5][16] , \keys[5][15] ,
         \keys[5][14] , \keys[5][13] , \keys[5][12] , \keys[5][11] ,
         \keys[5][10] , \keys[5][9] , \keys[5][8] , \keys[5][7] , \keys[5][6] ,
         \keys[5][5] , \keys[5][4] , \keys[5][3] , \keys[5][2] , \keys[5][1] ,
         \keys[5][0] , \keys[6][127] , \keys[6][126] , \keys[6][125] ,
         \keys[6][124] , \keys[6][123] , \keys[6][122] , \keys[6][121] ,
         \keys[6][120] , \keys[6][119] , \keys[6][118] , \keys[6][117] ,
         \keys[6][116] , \keys[6][115] , \keys[6][114] , \keys[6][113] ,
         \keys[6][112] , \keys[6][111] , \keys[6][110] , \keys[6][109] ,
         \keys[6][107] , \keys[6][106] , \keys[6][105] , \keys[6][104] ,
         \keys[6][103] , \keys[6][102] , \keys[6][101] , \keys[6][100] ,
         \keys[6][99] , \keys[6][98] , \keys[6][97] , \keys[6][96] ,
         \keys[6][95] , \keys[6][94] , \keys[6][93] , \keys[6][92] ,
         \keys[6][91] , \keys[6][90] , \keys[6][89] , \keys[6][88] ,
         \keys[6][87] , \keys[6][86] , \keys[6][85] , \keys[6][84] ,
         \keys[6][83] , \keys[6][82] , \keys[6][81] , \keys[6][80] ,
         \keys[6][79] , \keys[6][78] , \keys[6][77] , \keys[6][76] ,
         \keys[6][75] , \keys[6][74] , \keys[6][73] , \keys[6][72] ,
         \keys[6][71] , \keys[6][70] , \keys[6][69] , \keys[6][68] ,
         \keys[6][67] , \keys[6][66] , \keys[6][65] , \keys[6][64] ,
         \keys[6][63] , \keys[6][62] , \keys[6][61] , \keys[6][60] ,
         \keys[6][59] , \keys[6][58] , \keys[6][57] , \keys[6][56] ,
         \keys[6][55] , \keys[6][54] , \keys[6][53] , \keys[6][52] ,
         \keys[6][51] , \keys[6][50] , \keys[6][49] , \keys[6][48] ,
         \keys[6][47] , \keys[6][46] , \keys[6][45] , \keys[6][44] ,
         \keys[6][43] , \keys[6][42] , \keys[6][41] , \keys[6][40] ,
         \keys[6][39] , \keys[6][38] , \keys[6][37] , \keys[6][36] ,
         \keys[6][35] , \keys[6][34] , \keys[6][33] , \keys[6][32] ,
         \keys[6][31] , \keys[6][30] , \keys[6][29] , \keys[6][28] ,
         \keys[6][27] , \keys[6][26] , \keys[6][25] , \keys[6][24] ,
         \keys[6][23] , \keys[6][22] , \keys[6][21] , \keys[6][20] ,
         \keys[6][19] , \keys[6][18] , \keys[6][17] , \keys[6][16] ,
         \keys[6][15] , \keys[6][14] , \keys[6][13] , \keys[6][12] ,
         \keys[6][11] , \keys[6][10] , \keys[6][9] , \keys[6][8] ,
         \keys[6][7] , \keys[6][6] , \keys[6][5] , \keys[6][4] , \keys[6][3] ,
         \keys[6][2] , \keys[6][1] , \keys[6][0] , \keys[7][127] ,
         \keys[7][126] , \keys[7][125] , \keys[7][124] , \keys[7][123] ,
         \keys[7][122] , \keys[7][121] , \keys[7][120] , \keys[7][119] ,
         \keys[7][118] , \keys[7][117] , \keys[7][116] , \keys[7][115] ,
         \keys[7][114] , \keys[7][113] , \keys[7][112] , \keys[7][111] ,
         \keys[7][110] , \keys[7][109] , \keys[7][108] , \keys[7][107] ,
         \keys[7][106] , \keys[7][105] , \keys[7][104] , \keys[7][103] ,
         \keys[7][102] , \keys[7][101] , \keys[7][100] , \keys[7][99] ,
         \keys[7][98] , \keys[7][97] , \keys[7][96] , \keys[7][95] ,
         \keys[7][94] , \keys[7][93] , \keys[7][92] , \keys[7][91] ,
         \keys[7][90] , \keys[7][89] , \keys[7][88] , \keys[7][87] ,
         \keys[7][86] , \keys[7][85] , \keys[7][84] , \keys[7][83] ,
         \keys[7][82] , \keys[7][81] , \keys[7][80] , \keys[7][78] ,
         \keys[7][77] , \keys[7][76] , \keys[7][75] , \keys[7][72] ,
         \keys[7][71] , \keys[7][70] , \keys[7][69] , \keys[7][68] ,
         \keys[7][67] , \keys[7][66] , \keys[7][65] , \keys[7][64] ,
         \keys[7][63] , \keys[7][62] , \keys[7][61] , \keys[7][60] ,
         \keys[7][59] , \keys[7][58] , \keys[7][57] , \keys[7][56] ,
         \keys[7][55] , \keys[7][54] , \keys[7][53] , \keys[7][52] ,
         \keys[7][51] , \keys[7][50] , \keys[7][49] , \keys[7][48] ,
         \keys[7][47] , \keys[7][46] , \keys[7][45] , \keys[7][44] ,
         \keys[7][43] , \keys[7][42] , \keys[7][41] , \keys[7][40] ,
         \keys[7][39] , \keys[7][38] , \keys[7][37] , \keys[7][36] ,
         \keys[7][35] , \keys[7][34] , \keys[7][33] , \keys[7][32] ,
         \keys[7][31] , \keys[7][30] , \keys[7][29] , \keys[7][28] ,
         \keys[7][27] , \keys[7][26] , \keys[7][25] , \keys[7][24] ,
         \keys[7][23] , \keys[7][22] , \keys[7][21] , \keys[7][20] ,
         \keys[7][19] , \keys[7][18] , \keys[7][17] , \keys[7][16] ,
         \keys[7][15] , \keys[7][14] , \keys[7][13] , \keys[7][12] ,
         \keys[7][11] , \keys[7][10] , \keys[7][9] , \keys[7][8] ,
         \keys[7][7] , \keys[7][6] , \keys[7][5] , \keys[7][4] , \keys[7][3] ,
         \keys[7][2] , \keys[7][1] , \keys[7][0] , \keys[8][127] ,
         \keys[8][126] , \keys[8][125] , \keys[8][124] , \keys[8][123] ,
         \keys[8][122] , \keys[8][121] , \keys[8][120] , \keys[8][119] ,
         \keys[8][118] , \keys[8][117] , \keys[8][116] , \keys[8][115] ,
         \keys[8][114] , \keys[8][113] , \keys[8][112] , \keys[8][111] ,
         \keys[8][110] , \keys[8][109] , \keys[8][108] , \keys[8][107] ,
         \keys[8][106] , \keys[8][105] , \keys[8][104] , \keys[8][103] ,
         \keys[8][102] , \keys[8][101] , \keys[8][100] , \keys[8][99] ,
         \keys[8][98] , \keys[8][97] , \keys[8][96] , \keys[8][95] ,
         \keys[8][94] , \keys[8][93] , \keys[8][92] , \keys[8][91] ,
         \keys[8][90] , \keys[8][89] , \keys[8][88] , \keys[8][87] ,
         \keys[8][86] , \keys[8][85] , \keys[8][84] , \keys[8][83] ,
         \keys[8][82] , \keys[8][81] , \keys[8][80] , \keys[8][79] ,
         \keys[8][78] , \keys[8][77] , \keys[8][76] , \keys[8][75] ,
         \keys[8][74] , \keys[8][73] , \keys[8][72] , \keys[8][71] ,
         \keys[8][70] , \keys[8][69] , \keys[8][68] , \keys[8][67] ,
         \keys[8][66] , \keys[8][65] , \keys[8][64] , \keys[8][63] ,
         \keys[8][62] , \keys[8][61] , \keys[8][60] , \keys[8][59] ,
         \keys[8][58] , \keys[8][57] , \keys[8][56] , \keys[8][55] ,
         \keys[8][54] , \keys[8][53] , \keys[8][52] , \keys[8][51] ,
         \keys[8][50] , \keys[8][49] , \keys[8][48] , \keys[8][47] ,
         \keys[8][46] , \keys[8][45] , \keys[8][44] , \keys[8][43] ,
         \keys[8][42] , \keys[8][41] , \keys[8][40] , \keys[8][39] ,
         \keys[8][38] , \keys[8][37] , \keys[8][36] , \keys[8][35] ,
         \keys[8][34] , \keys[8][33] , \keys[8][32] , \keys[8][31] ,
         \keys[8][30] , \keys[8][29] , \keys[8][28] , \keys[8][27] ,
         \keys[8][26] , \keys[8][25] , \keys[8][24] , \keys[8][23] ,
         \keys[8][22] , \keys[8][21] , \keys[8][20] , \keys[8][19] ,
         \keys[8][18] , \keys[8][17] , \keys[8][16] , \keys[8][15] ,
         \keys[8][14] , \keys[8][13] , \keys[8][12] , \keys[8][11] ,
         \keys[8][10] , \keys[8][9] , \keys[8][8] , \keys[8][7] , \keys[8][6] ,
         \keys[8][5] , \keys[8][4] , \keys[8][3] , \keys[8][2] , \keys[8][1] ,
         \keys[8][0] , \keys[9][127] , \keys[9][126] , \keys[9][125] ,
         \keys[9][124] , \keys[9][123] , \keys[9][122] , \keys[9][121] ,
         \keys[9][120] , \keys[9][119] , \keys[9][118] , \keys[9][117] ,
         \keys[9][116] , \keys[9][115] , \keys[9][114] , \keys[9][113] ,
         \keys[9][112] , \keys[9][111] , \keys[9][110] , \keys[9][109] ,
         \keys[9][108] , \keys[9][107] , \keys[9][106] , \keys[9][105] ,
         \keys[9][104] , \keys[9][103] , \keys[9][102] , \keys[9][101] ,
         \keys[9][100] , \keys[9][99] , \keys[9][98] , \keys[9][97] ,
         \keys[9][96] , \keys[9][95] , \keys[9][94] , \keys[9][93] ,
         \keys[9][92] , \keys[9][91] , \keys[9][90] , \keys[9][89] ,
         \keys[9][88] , \keys[9][87] , \keys[9][86] , \keys[9][85] ,
         \keys[9][84] , \keys[9][83] , \keys[9][82] , \keys[9][81] ,
         \keys[9][80] , \keys[9][79] , \keys[9][78] , \keys[9][77] ,
         \keys[9][76] , \keys[9][75] , \keys[9][74] , \keys[9][73] ,
         \keys[9][72] , \keys[9][71] , \keys[9][70] , \keys[9][69] ,
         \keys[9][68] , \keys[9][67] , \keys[9][66] , \keys[9][65] ,
         \keys[9][64] , \keys[9][63] , \keys[9][62] , \keys[9][61] ,
         \keys[9][60] , \keys[9][59] , \keys[9][58] , \keys[9][57] ,
         \keys[9][56] , \keys[9][55] , \keys[9][54] , \keys[9][53] ,
         \keys[9][52] , \keys[9][51] , \keys[9][50] , \keys[9][49] ,
         \keys[9][48] , \keys[9][47] , \keys[9][46] , \keys[9][45] ,
         \keys[9][44] , \keys[9][43] , \keys[9][42] , \keys[9][41] ,
         \keys[9][40] , \keys[9][39] , \keys[9][38] , \keys[9][37] ,
         \keys[9][36] , \keys[9][35] , \keys[9][34] , \keys[9][33] ,
         \keys[9][32] , \keys[9][31] , \keys[9][30] , \keys[9][29] ,
         \keys[9][28] , \keys[9][27] , \keys[9][26] , \keys[9][25] ,
         \keys[9][24] , \keys[9][23] , \keys[9][22] , \keys[9][21] ,
         \keys[9][20] , \keys[9][19] , \keys[9][18] , \keys[9][17] ,
         \keys[9][16] , \keys[9][15] , \keys[9][14] , \keys[9][13] ,
         \keys[9][12] , \keys[9][11] , \keys[9][10] , \keys[9][9] ,
         \keys[9][8] , \keys[9][7] , \keys[9][6] , \keys[9][5] , \keys[9][4] ,
         \keys[9][3] , \keys[9][2] , \keys[9][1] , \keys[9][0] ,
         \keys[10][127] , \keys[10][126] , \keys[10][125] , \keys[10][124] ,
         \keys[10][123] , \keys[10][122] , \keys[10][121] , \keys[10][120] ,
         \keys[10][119] , \keys[10][118] , \keys[10][117] , \keys[10][116] ,
         \keys[10][115] , \keys[10][114] , \keys[10][113] , \keys[10][112] ,
         \keys[10][111] , \keys[10][110] , \keys[10][109] , \keys[10][108] ,
         \keys[10][107] , \keys[10][106] , \keys[10][105] , \keys[10][104] ,
         \keys[10][103] , \keys[10][102] , \keys[10][101] , \keys[10][100] ,
         \keys[10][99] , \keys[10][98] , \keys[10][97] , \keys[10][96] ,
         \keys[10][95] , \keys[10][94] , \keys[10][93] , \keys[10][92] ,
         \keys[10][91] , \keys[10][89] , \keys[10][88] , \keys[10][87] ,
         \keys[10][86] , \keys[10][85] , \keys[10][84] , \keys[10][83] ,
         \keys[10][82] , \keys[10][81] , \keys[10][80] , \keys[10][79] ,
         \keys[10][78] , \keys[10][77] , \keys[10][76] , \keys[10][75] ,
         \keys[10][74] , \keys[10][73] , \keys[10][72] , \keys[10][71] ,
         \keys[10][70] , \keys[10][69] , \keys[10][68] , \keys[10][67] ,
         \keys[10][66] , \keys[10][65] , \keys[10][64] , \keys[10][63] ,
         \keys[10][62] , \keys[10][61] , \keys[10][60] , \keys[10][59] ,
         \keys[10][58] , \keys[10][57] , \keys[10][56] , \keys[10][55] ,
         \keys[10][54] , \keys[10][53] , \keys[10][52] , \keys[10][51] ,
         \keys[10][50] , \keys[10][49] , \keys[10][48] , \keys[10][47] ,
         \keys[10][46] , \keys[10][45] , \keys[10][44] , \keys[10][43] ,
         \keys[10][42] , \keys[10][41] , \keys[10][40] , \keys[10][39] ,
         \keys[10][38] , \keys[10][37] , \keys[10][36] , \keys[10][35] ,
         \keys[10][34] , \keys[10][33] , \keys[10][32] , \keys[10][31] ,
         \keys[10][30] , \keys[10][29] , \keys[10][28] , \keys[10][27] ,
         \keys[10][26] , \keys[10][25] , \keys[10][24] , \keys[10][23] ,
         \keys[10][22] , \keys[10][21] , \keys[10][20] , \keys[10][19] ,
         \keys[10][18] , \keys[10][17] , \keys[10][16] , \keys[10][15] ,
         \keys[10][14] , \keys[10][13] , \keys[10][12] , \keys[10][11] ,
         \keys[10][10] , \keys[10][9] , \keys[10][8] , \keys[10][7] ,
         \keys[10][6] , \keys[10][5] , \keys[10][4] , \keys[10][3] ,
         \keys[10][2] , \keys[10][1] , \keys[10][0] , n11, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1430, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n1427,
         n1428, n1429, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559;
  wire   [3:0] round_number;
  wire   [127:0] prev_key;
  wire   [127:0] keyout;
  wire   [3:0] state;
  tri   clk;
  tri   rest;

  DFFX1_HVT \state_reg[0]  ( .D(n3797), .CLK(clk), .Q(state[0]), .QN(n18) );
  DFFX1_HVT \state_reg[3]  ( .D(n3796), .CLK(clk), .Q(state[3]), .QN(n11) );
  DFFX1_HVT \state_reg[2]  ( .D(n3794), .CLK(clk), .Q(state[2]), .QN(n16) );
  DFFX1_HVT \state_reg[1]  ( .D(n3795), .CLK(clk), .Q(state[1]), .QN(n17) );
  DFFX1_HVT done_reg ( .D(n3793), .CLK(clk), .Q(done) );
  DFFX1_HVT \round_number_reg[2]  ( .D(n3790), .CLK(clk), .Q(round_number[2])
         );
  DFFX1_HVT \round_number_reg[3]  ( .D(n3789), .CLK(clk), .Q(round_number[3])
         );
  DFFX1_HVT \round_number_reg[0]  ( .D(n3792), .CLK(clk), .Q(round_number[0])
         );
  DFFX1_HVT \round_number_reg[1]  ( .D(n3791), .CLK(clk), .Q(round_number[1])
         );
  DFFX1_HVT \prev_key_reg[0]  ( .D(n3788), .CLK(clk), .Q(prev_key[0]) );
  DFFX1_HVT \prev_key_reg[1]  ( .D(n3787), .CLK(clk), .Q(prev_key[1]) );
  DFFX1_HVT \prev_key_reg[2]  ( .D(n3786), .CLK(clk), .Q(prev_key[2]), .QN(
        n3847) );
  DFFX1_HVT \prev_key_reg[3]  ( .D(n3785), .CLK(clk), .Q(prev_key[3]) );
  DFFX1_HVT \prev_key_reg[4]  ( .D(n3784), .CLK(clk), .Q(prev_key[4]) );
  DFFX1_HVT \prev_key_reg[5]  ( .D(n3783), .CLK(clk), .Q(prev_key[5]) );
  DFFX1_HVT \prev_key_reg[6]  ( .D(n3782), .CLK(clk), .Q(prev_key[6]) );
  DFFX1_HVT \prev_key_reg[7]  ( .D(n3781), .CLK(clk), .Q(prev_key[7]), .QN(
        n3899) );
  DFFX1_HVT \prev_key_reg[8]  ( .D(n3780), .CLK(clk), .Q(prev_key[8]) );
  DFFX1_HVT \prev_key_reg[9]  ( .D(n3779), .CLK(clk), .Q(prev_key[9]) );
  DFFX1_HVT \prev_key_reg[10]  ( .D(n3778), .CLK(clk), .Q(prev_key[10]), .QN(
        n3917) );
  DFFX1_HVT \prev_key_reg[11]  ( .D(n3777), .CLK(clk), .Q(prev_key[11]) );
  DFFX1_HVT \prev_key_reg[12]  ( .D(n3776), .CLK(clk), .Q(prev_key[12]) );
  DFFX1_HVT \prev_key_reg[13]  ( .D(n3775), .CLK(clk), .Q(prev_key[13]) );
  DFFX1_HVT \prev_key_reg[14]  ( .D(n3774), .CLK(clk), .Q(prev_key[14]) );
  DFFX1_HVT \prev_key_reg[15]  ( .D(n3773), .CLK(clk), .Q(n3975), .QN(n6) );
  DFFX1_HVT \prev_key_reg[16]  ( .D(n3772), .CLK(clk), .Q(prev_key[16]) );
  DFFX1_HVT \prev_key_reg[17]  ( .D(n3771), .CLK(clk), .Q(prev_key[17]), .QN(
        n8) );
  DFFX1_HVT \prev_key_reg[18]  ( .D(n3770), .CLK(clk), .Q(prev_key[18]), .QN(
        n3932) );
  DFFX1_HVT \prev_key_reg[19]  ( .D(n3769), .CLK(clk), .Q(prev_key[19]) );
  DFFX1_HVT \prev_key_reg[20]  ( .D(n3768), .CLK(clk), .Q(prev_key[20]) );
  DFFX1_HVT \prev_key_reg[21]  ( .D(n3767), .CLK(clk), .Q(prev_key[21]) );
  DFFX1_HVT \prev_key_reg[22]  ( .D(n3766), .CLK(clk), .Q(prev_key[22]) );
  DFFX1_HVT \prev_key_reg[23]  ( .D(n3765), .CLK(clk), .Q(n3954), .QN(n3821)
         );
  DFFX1_HVT \prev_key_reg[24]  ( .D(n3764), .CLK(clk), .Q(prev_key[24]) );
  DFFX1_HVT \prev_key_reg[25]  ( .D(n3763), .CLK(clk), .Q(prev_key[25]) );
  DFFX1_HVT \prev_key_reg[26]  ( .D(n3762), .CLK(clk), .Q(prev_key[26]) );
  DFFX1_HVT \prev_key_reg[27]  ( .D(n3761), .CLK(clk), .Q(prev_key[27]) );
  DFFX1_HVT \prev_key_reg[28]  ( .D(n3760), .CLK(clk), .Q(prev_key[28]) );
  DFFX1_HVT \prev_key_reg[29]  ( .D(n3759), .CLK(clk), .Q(prev_key[29]) );
  DFFX1_HVT \prev_key_reg[30]  ( .D(n3758), .CLK(clk), .Q(prev_key[30]) );
  DFFX1_HVT \prev_key_reg[31]  ( .D(n3757), .CLK(clk), .Q(prev_key[31]) );
  DFFX1_HVT \prev_key_reg[32]  ( .D(n3756), .CLK(clk), .Q(prev_key[32]) );
  DFFX1_HVT \prev_key_reg[33]  ( .D(n3755), .CLK(clk), .Q(prev_key[33]) );
  DFFX1_HVT \prev_key_reg[34]  ( .D(n3754), .CLK(clk), .Q(prev_key[34]) );
  DFFX1_HVT \prev_key_reg[35]  ( .D(n3753), .CLK(clk), .Q(prev_key[35]) );
  DFFX1_HVT \prev_key_reg[36]  ( .D(n3752), .CLK(clk), .Q(prev_key[36]) );
  DFFX1_HVT \prev_key_reg[37]  ( .D(n3751), .CLK(clk), .Q(prev_key[37]) );
  DFFX1_HVT \prev_key_reg[38]  ( .D(n3750), .CLK(clk), .Q(prev_key[38]) );
  DFFX1_HVT \prev_key_reg[39]  ( .D(n3749), .CLK(clk), .Q(prev_key[39]) );
  DFFX1_HVT \prev_key_reg[40]  ( .D(n3748), .CLK(clk), .Q(prev_key[40]) );
  DFFX1_HVT \prev_key_reg[41]  ( .D(n3747), .CLK(clk), .Q(prev_key[41]) );
  DFFX1_HVT \prev_key_reg[42]  ( .D(n3746), .CLK(clk), .Q(prev_key[42]) );
  DFFX1_HVT \prev_key_reg[43]  ( .D(n3745), .CLK(clk), .Q(prev_key[43]) );
  DFFX1_HVT \prev_key_reg[44]  ( .D(n3744), .CLK(clk), .Q(prev_key[44]) );
  DFFX1_HVT \prev_key_reg[45]  ( .D(n3743), .CLK(clk), .Q(prev_key[45]) );
  DFFX1_HVT \prev_key_reg[46]  ( .D(n3742), .CLK(clk), .Q(prev_key[46]) );
  DFFX1_HVT \prev_key_reg[47]  ( .D(n3741), .CLK(clk), .Q(prev_key[47]) );
  DFFX1_HVT \prev_key_reg[48]  ( .D(n3740), .CLK(clk), .Q(prev_key[48]) );
  DFFX1_HVT \prev_key_reg[49]  ( .D(n3739), .CLK(clk), .Q(prev_key[49]) );
  DFFX1_HVT \prev_key_reg[50]  ( .D(n3738), .CLK(clk), .Q(prev_key[50]) );
  DFFX1_HVT \prev_key_reg[51]  ( .D(n3737), .CLK(clk), .Q(prev_key[51]) );
  DFFX1_HVT \prev_key_reg[52]  ( .D(n3736), .CLK(clk), .Q(prev_key[52]) );
  DFFX1_HVT \prev_key_reg[53]  ( .D(n3735), .CLK(clk), .Q(prev_key[53]) );
  DFFX1_HVT \prev_key_reg[54]  ( .D(n3734), .CLK(clk), .Q(prev_key[54]) );
  DFFX1_HVT \prev_key_reg[55]  ( .D(n3733), .CLK(clk), .Q(prev_key[55]) );
  DFFX1_HVT \prev_key_reg[56]  ( .D(n3732), .CLK(clk), .Q(prev_key[56]) );
  DFFX1_HVT \prev_key_reg[57]  ( .D(n3731), .CLK(clk), .Q(prev_key[57]) );
  DFFX1_HVT \prev_key_reg[58]  ( .D(n3730), .CLK(clk), .Q(prev_key[58]) );
  DFFX1_HVT \prev_key_reg[59]  ( .D(n3729), .CLK(clk), .Q(prev_key[59]) );
  DFFX1_HVT \prev_key_reg[60]  ( .D(n3728), .CLK(clk), .Q(prev_key[60]) );
  DFFX1_HVT \prev_key_reg[61]  ( .D(n3727), .CLK(clk), .Q(prev_key[61]), .QN(
        n3807) );
  DFFX1_HVT \prev_key_reg[62]  ( .D(n3726), .CLK(clk), .Q(prev_key[62]) );
  DFFX1_HVT \prev_key_reg[63]  ( .D(n3725), .CLK(clk), .Q(prev_key[63]) );
  DFFX1_HVT \prev_key_reg[64]  ( .D(n3724), .CLK(clk), .Q(prev_key[64]) );
  DFFX1_HVT \prev_key_reg[65]  ( .D(n3723), .CLK(clk), .Q(prev_key[65]) );
  DFFX1_HVT \prev_key_reg[66]  ( .D(n3722), .CLK(clk), .Q(prev_key[66]) );
  DFFX1_HVT \prev_key_reg[67]  ( .D(n3721), .CLK(clk), .Q(prev_key[67]) );
  DFFX1_HVT \prev_key_reg[68]  ( .D(n3720), .CLK(clk), .Q(prev_key[68]) );
  DFFX1_HVT \prev_key_reg[69]  ( .D(n3719), .CLK(clk), .Q(prev_key[69]) );
  DFFX1_HVT \prev_key_reg[70]  ( .D(n3718), .CLK(clk), .Q(prev_key[70]) );
  DFFX1_HVT \prev_key_reg[71]  ( .D(n3717), .CLK(clk), .Q(prev_key[71]) );
  DFFX1_HVT \prev_key_reg[72]  ( .D(n3716), .CLK(clk), .Q(prev_key[72]) );
  DFFX1_HVT \prev_key_reg[73]  ( .D(n3715), .CLK(clk), .Q(prev_key[73]) );
  DFFX1_HVT \prev_key_reg[74]  ( .D(n3714), .CLK(clk), .Q(prev_key[74]) );
  DFFX1_HVT \prev_key_reg[75]  ( .D(n3713), .CLK(clk), .Q(prev_key[75]) );
  DFFX1_HVT \prev_key_reg[76]  ( .D(n3712), .CLK(clk), .Q(prev_key[76]) );
  DFFX1_HVT \prev_key_reg[77]  ( .D(n3711), .CLK(clk), .Q(prev_key[77]) );
  DFFX1_HVT \prev_key_reg[78]  ( .D(n3710), .CLK(clk), .Q(prev_key[78]) );
  DFFX1_HVT \prev_key_reg[79]  ( .D(n3709), .CLK(clk), .Q(prev_key[79]) );
  DFFX1_HVT \prev_key_reg[80]  ( .D(n3708), .CLK(clk), .Q(prev_key[80]) );
  DFFX1_HVT \prev_key_reg[81]  ( .D(n3707), .CLK(clk), .Q(prev_key[81]) );
  DFFX1_HVT \prev_key_reg[82]  ( .D(n3706), .CLK(clk), .Q(prev_key[82]) );
  DFFX1_HVT \prev_key_reg[83]  ( .D(n3705), .CLK(clk), .Q(prev_key[83]) );
  DFFX1_HVT \prev_key_reg[84]  ( .D(n3704), .CLK(clk), .Q(prev_key[84]) );
  DFFX1_HVT \prev_key_reg[85]  ( .D(n3703), .CLK(clk), .Q(prev_key[85]) );
  DFFX1_HVT \prev_key_reg[86]  ( .D(n3702), .CLK(clk), .Q(prev_key[86]) );
  DFFX1_HVT \prev_key_reg[87]  ( .D(n3701), .CLK(clk), .Q(prev_key[87]), .QN(
        n3801) );
  DFFX1_HVT \prev_key_reg[88]  ( .D(n3700), .CLK(clk), .Q(prev_key[88]) );
  DFFX1_HVT \prev_key_reg[89]  ( .D(n3699), .CLK(clk), .Q(prev_key[89]) );
  DFFX1_HVT \prev_key_reg[90]  ( .D(n3698), .CLK(clk), .Q(prev_key[90]) );
  DFFX1_HVT \prev_key_reg[91]  ( .D(n3697), .CLK(clk), .Q(prev_key[91]) );
  DFFX1_HVT \prev_key_reg[92]  ( .D(n3696), .CLK(clk), .Q(prev_key[92]) );
  DFFX1_HVT \prev_key_reg[93]  ( .D(n3695), .CLK(clk), .Q(prev_key[93]) );
  DFFX1_HVT \prev_key_reg[94]  ( .D(n3694), .CLK(clk), .Q(prev_key[94]) );
  DFFX1_HVT \prev_key_reg[95]  ( .D(n3693), .CLK(clk), .Q(prev_key[95]) );
  DFFX1_HVT \prev_key_reg[96]  ( .D(n3692), .CLK(clk), .Q(prev_key[96]) );
  DFFX1_HVT \prev_key_reg[97]  ( .D(n3691), .CLK(clk), .Q(prev_key[97]) );
  DFFX1_HVT \prev_key_reg[98]  ( .D(n3690), .CLK(clk), .Q(prev_key[98]) );
  DFFX1_HVT \prev_key_reg[99]  ( .D(n3689), .CLK(clk), .Q(prev_key[99]) );
  DFFX1_HVT \prev_key_reg[100]  ( .D(n3688), .CLK(clk), .Q(prev_key[100]) );
  DFFX1_HVT \prev_key_reg[101]  ( .D(n3687), .CLK(clk), .Q(prev_key[101]) );
  DFFX1_HVT \prev_key_reg[102]  ( .D(n3686), .CLK(clk), .Q(prev_key[102]) );
  DFFX1_HVT \prev_key_reg[103]  ( .D(n3685), .CLK(clk), .Q(prev_key[103]) );
  DFFX1_HVT \prev_key_reg[104]  ( .D(n3684), .CLK(clk), .Q(prev_key[104]) );
  DFFX1_HVT \prev_key_reg[105]  ( .D(n3683), .CLK(clk), .Q(prev_key[105]) );
  DFFX1_HVT \prev_key_reg[106]  ( .D(n3682), .CLK(clk), .Q(prev_key[106]) );
  DFFX1_HVT \prev_key_reg[107]  ( .D(n3681), .CLK(clk), .Q(prev_key[107]) );
  DFFX1_HVT \prev_key_reg[108]  ( .D(n3680), .CLK(clk), .Q(prev_key[108]) );
  DFFX1_HVT \prev_key_reg[109]  ( .D(n3679), .CLK(clk), .Q(prev_key[109]) );
  DFFX1_HVT \prev_key_reg[110]  ( .D(n3678), .CLK(clk), .Q(prev_key[110]) );
  DFFX1_HVT \prev_key_reg[111]  ( .D(n3677), .CLK(clk), .Q(prev_key[111]) );
  DFFX1_HVT \prev_key_reg[112]  ( .D(n3676), .CLK(clk), .Q(prev_key[112]) );
  DFFX1_HVT \prev_key_reg[113]  ( .D(n3675), .CLK(clk), .Q(prev_key[113]) );
  DFFX1_HVT \prev_key_reg[114]  ( .D(n3674), .CLK(clk), .Q(prev_key[114]) );
  DFFX1_HVT \prev_key_reg[115]  ( .D(n3673), .CLK(clk), .Q(prev_key[115]) );
  DFFX1_HVT \prev_key_reg[116]  ( .D(n3672), .CLK(clk), .Q(prev_key[116]) );
  DFFX1_HVT \prev_key_reg[117]  ( .D(n3671), .CLK(clk), .Q(prev_key[117]) );
  DFFX1_HVT \prev_key_reg[118]  ( .D(n3670), .CLK(clk), .Q(prev_key[118]) );
  DFFX1_HVT \prev_key_reg[119]  ( .D(n3669), .CLK(clk), .Q(prev_key[119]) );
  DFFX1_HVT \prev_key_reg[120]  ( .D(n3668), .CLK(clk), .Q(prev_key[120]) );
  DFFX1_HVT \prev_key_reg[121]  ( .D(n3667), .CLK(clk), .Q(prev_key[121]) );
  DFFX1_HVT \prev_key_reg[122]  ( .D(n3666), .CLK(clk), .Q(prev_key[122]) );
  DFFX1_HVT \prev_key_reg[123]  ( .D(n3665), .CLK(clk), .Q(prev_key[123]) );
  DFFX1_HVT \prev_key_reg[124]  ( .D(n3664), .CLK(clk), .Q(prev_key[124]) );
  DFFX1_HVT \prev_key_reg[125]  ( .D(n3663), .CLK(clk), .Q(prev_key[125]) );
  DFFX1_HVT \prev_key_reg[126]  ( .D(n3662), .CLK(clk), .Q(prev_key[126]) );
  DFFX1_HVT \prev_key_reg[127]  ( .D(n3661), .CLK(clk), .Q(prev_key[127]) );
  DFFX1_HVT \keys_reg[0][127]  ( .D(n3660), .CLK(clk), .Q(\keys[0][127] ), 
        .QN(n19) );
  DFFX1_HVT \keys_reg[0][126]  ( .D(n3659), .CLK(clk), .Q(\keys[0][126] ), 
        .QN(n20) );
  DFFX1_HVT \keys_reg[0][125]  ( .D(n3658), .CLK(clk), .Q(\keys[0][125] ), 
        .QN(n21) );
  DFFX1_HVT \keys_reg[0][124]  ( .D(n3657), .CLK(clk), .Q(\keys[0][124] ), 
        .QN(n22) );
  DFFX1_HVT \keys_reg[0][123]  ( .D(n3656), .CLK(clk), .Q(\keys[0][123] ), 
        .QN(n23) );
  DFFX1_HVT \keys_reg[0][122]  ( .D(n3655), .CLK(clk), .Q(\keys[0][122] ), 
        .QN(n24) );
  DFFX1_HVT \keys_reg[0][121]  ( .D(n3654), .CLK(clk), .Q(\keys[0][121] ), 
        .QN(n25) );
  DFFX1_HVT \keys_reg[0][120]  ( .D(n3653), .CLK(clk), .Q(\keys[0][120] ), 
        .QN(n26) );
  DFFX1_HVT \keys_reg[0][119]  ( .D(n3652), .CLK(clk), .Q(\keys[0][119] ), 
        .QN(n27) );
  DFFX1_HVT \keys_reg[0][118]  ( .D(n3651), .CLK(clk), .Q(\keys[0][118] ), 
        .QN(n28) );
  DFFX1_HVT \keys_reg[0][117]  ( .D(n3650), .CLK(clk), .Q(\keys[0][117] ), 
        .QN(n29) );
  DFFX1_HVT \keys_reg[0][116]  ( .D(n3649), .CLK(clk), .Q(\keys[0][116] ), 
        .QN(n30) );
  DFFX1_HVT \keys_reg[0][115]  ( .D(n3648), .CLK(clk), .Q(\keys[0][115] ), 
        .QN(n31) );
  DFFX1_HVT \keys_reg[0][114]  ( .D(n3647), .CLK(clk), .Q(\keys[0][114] ), 
        .QN(n32) );
  DFFX1_HVT \keys_reg[0][113]  ( .D(n3646), .CLK(clk), .Q(\keys[0][113] ), 
        .QN(n33) );
  DFFX1_HVT \keys_reg[0][112]  ( .D(n3645), .CLK(clk), .Q(\keys[0][112] ), 
        .QN(n34) );
  DFFX1_HVT \keys_reg[0][111]  ( .D(n3644), .CLK(clk), .Q(\keys[0][111] ), 
        .QN(n35) );
  DFFX1_HVT \keys_reg[0][110]  ( .D(n3643), .CLK(clk), .Q(\keys[0][110] ), 
        .QN(n36) );
  DFFX1_HVT \keys_reg[0][109]  ( .D(n3642), .CLK(clk), .Q(\keys[0][109] ), 
        .QN(n37) );
  DFFX1_HVT \keys_reg[0][108]  ( .D(n3641), .CLK(clk), .Q(\keys[0][108] ), 
        .QN(n38) );
  DFFX1_HVT \keys_reg[0][107]  ( .D(n3640), .CLK(clk), .Q(\keys[0][107] ), 
        .QN(n39) );
  DFFX1_HVT \keys_reg[0][106]  ( .D(n3639), .CLK(clk), .Q(\keys[0][106] ), 
        .QN(n40) );
  DFFX1_HVT \keys_reg[0][105]  ( .D(n3638), .CLK(clk), .Q(\keys[0][105] ), 
        .QN(n41) );
  DFFX1_HVT \keys_reg[0][104]  ( .D(n3637), .CLK(clk), .Q(\keys[0][104] ), 
        .QN(n42) );
  DFFX1_HVT \keys_reg[0][103]  ( .D(n3636), .CLK(clk), .Q(\keys[0][103] ), 
        .QN(n43) );
  DFFX1_HVT \keys_reg[0][102]  ( .D(n3635), .CLK(clk), .Q(\keys[0][102] ), 
        .QN(n44) );
  DFFX1_HVT \keys_reg[0][101]  ( .D(n3634), .CLK(clk), .Q(\keys[0][101] ), 
        .QN(n45) );
  DFFX1_HVT \keys_reg[0][100]  ( .D(n3633), .CLK(clk), .Q(\keys[0][100] ), 
        .QN(n46) );
  DFFX1_HVT \keys_reg[0][99]  ( .D(n3632), .CLK(clk), .Q(\keys[0][99] ), .QN(
        n47) );
  DFFX1_HVT \keys_reg[0][98]  ( .D(n3631), .CLK(clk), .Q(\keys[0][98] ), .QN(
        n48) );
  DFFX1_HVT \keys_reg[0][97]  ( .D(n3630), .CLK(clk), .Q(\keys[0][97] ), .QN(
        n49) );
  DFFX1_HVT \keys_reg[0][96]  ( .D(n3629), .CLK(clk), .Q(\keys[0][96] ), .QN(
        n50) );
  DFFX1_HVT \keys_reg[0][95]  ( .D(n3628), .CLK(clk), .Q(\keys[0][95] ), .QN(
        n51) );
  DFFX1_HVT \keys_reg[0][94]  ( .D(n3627), .CLK(clk), .Q(\keys[0][94] ), .QN(
        n52) );
  DFFX1_HVT \keys_reg[0][93]  ( .D(n3626), .CLK(clk), .Q(\keys[0][93] ), .QN(
        n53) );
  DFFX1_HVT \keys_reg[0][92]  ( .D(n3625), .CLK(clk), .Q(\keys[0][92] ), .QN(
        n54) );
  DFFX1_HVT \keys_reg[0][91]  ( .D(n3624), .CLK(clk), .Q(\keys[0][91] ), .QN(
        n55) );
  DFFX1_HVT \keys_reg[0][90]  ( .D(n3623), .CLK(clk), .Q(\keys[0][90] ), .QN(
        n56) );
  DFFX1_HVT \keys_reg[0][89]  ( .D(n3622), .CLK(clk), .Q(\keys[0][89] ), .QN(
        n57) );
  DFFX1_HVT \keys_reg[0][88]  ( .D(n3621), .CLK(clk), .Q(\keys[0][88] ), .QN(
        n58) );
  DFFX1_HVT \keys_reg[0][87]  ( .D(n3620), .CLK(clk), .Q(\keys[0][87] ), .QN(
        n59) );
  DFFX1_HVT \keys_reg[0][86]  ( .D(n3619), .CLK(clk), .Q(\keys[0][86] ), .QN(
        n60) );
  DFFX1_HVT \keys_reg[0][85]  ( .D(n3618), .CLK(clk), .Q(\keys[0][85] ), .QN(
        n61) );
  DFFX1_HVT \keys_reg[0][84]  ( .D(n3617), .CLK(clk), .Q(\keys[0][84] ), .QN(
        n62) );
  DFFX1_HVT \keys_reg[0][83]  ( .D(n3616), .CLK(clk), .Q(\keys[0][83] ), .QN(
        n63) );
  DFFX1_HVT \keys_reg[0][82]  ( .D(n3615), .CLK(clk), .Q(\keys[0][82] ), .QN(
        n64) );
  DFFX1_HVT \keys_reg[0][81]  ( .D(n3614), .CLK(clk), .Q(\keys[0][81] ), .QN(
        n65) );
  DFFX1_HVT \keys_reg[0][80]  ( .D(n3613), .CLK(clk), .Q(\keys[0][80] ), .QN(
        n66) );
  DFFX1_HVT \keys_reg[0][79]  ( .D(n3612), .CLK(clk), .Q(\keys[0][79] ), .QN(
        n67) );
  DFFX1_HVT \keys_reg[0][78]  ( .D(n3611), .CLK(clk), .Q(\keys[0][78] ), .QN(
        n68) );
  DFFX1_HVT \keys_reg[0][77]  ( .D(n3610), .CLK(clk), .Q(\keys[0][77] ), .QN(
        n69) );
  DFFX1_HVT \keys_reg[0][76]  ( .D(n3609), .CLK(clk), .Q(\keys[0][76] ), .QN(
        n70) );
  DFFX1_HVT \keys_reg[0][75]  ( .D(n3608), .CLK(clk), .Q(\keys[0][75] ), .QN(
        n71) );
  DFFX1_HVT \keys_reg[0][74]  ( .D(n3607), .CLK(clk), .Q(\keys[0][74] ), .QN(
        n72) );
  DFFX1_HVT \keys_reg[0][73]  ( .D(n3606), .CLK(clk), .Q(\keys[0][73] ), .QN(
        n73) );
  DFFX1_HVT \keys_reg[0][72]  ( .D(n3605), .CLK(clk), .Q(\keys[0][72] ), .QN(
        n74) );
  DFFX1_HVT \keys_reg[0][71]  ( .D(n3604), .CLK(clk), .Q(\keys[0][71] ), .QN(
        n75) );
  DFFX1_HVT \keys_reg[0][70]  ( .D(n3603), .CLK(clk), .Q(\keys[0][70] ), .QN(
        n76) );
  DFFX1_HVT \keys_reg[0][69]  ( .D(n3602), .CLK(clk), .Q(\keys[0][69] ), .QN(
        n77) );
  DFFX1_HVT \keys_reg[0][68]  ( .D(n3601), .CLK(clk), .Q(\keys[0][68] ), .QN(
        n78) );
  DFFX1_HVT \keys_reg[0][67]  ( .D(n3600), .CLK(clk), .Q(\keys[0][67] ), .QN(
        n79) );
  DFFX1_HVT \keys_reg[0][66]  ( .D(n3599), .CLK(clk), .Q(\keys[0][66] ), .QN(
        n80) );
  DFFX1_HVT \keys_reg[0][65]  ( .D(n3598), .CLK(clk), .Q(\keys[0][65] ), .QN(
        n81) );
  DFFX1_HVT \keys_reg[0][64]  ( .D(n3597), .CLK(clk), .Q(\keys[0][64] ), .QN(
        n82) );
  DFFX1_HVT \keys_reg[0][63]  ( .D(n3596), .CLK(clk), .Q(\keys[0][63] ), .QN(
        n83) );
  DFFX1_HVT \keys_reg[0][62]  ( .D(n3595), .CLK(clk), .Q(\keys[0][62] ), .QN(
        n84) );
  DFFX1_HVT \keys_reg[0][61]  ( .D(n3594), .CLK(clk), .Q(\keys[0][61] ), .QN(
        n85) );
  DFFX1_HVT \keys_reg[0][60]  ( .D(n3593), .CLK(clk), .Q(\keys[0][60] ), .QN(
        n86) );
  DFFX1_HVT \keys_reg[0][59]  ( .D(n3592), .CLK(clk), .Q(\keys[0][59] ), .QN(
        n87) );
  DFFX1_HVT \keys_reg[0][58]  ( .D(n3591), .CLK(clk), .Q(\keys[0][58] ), .QN(
        n88) );
  DFFX1_HVT \keys_reg[0][57]  ( .D(n3590), .CLK(clk), .Q(\keys[0][57] ), .QN(
        n89) );
  DFFX1_HVT \keys_reg[0][56]  ( .D(n3589), .CLK(clk), .Q(\keys[0][56] ), .QN(
        n90) );
  DFFX1_HVT \keys_reg[0][55]  ( .D(n3588), .CLK(clk), .Q(\keys[0][55] ), .QN(
        n91) );
  DFFX1_HVT \keys_reg[0][54]  ( .D(n3587), .CLK(clk), .Q(\keys[0][54] ), .QN(
        n92) );
  DFFX1_HVT \keys_reg[0][53]  ( .D(n3586), .CLK(clk), .Q(\keys[0][53] ), .QN(
        n93) );
  DFFX1_HVT \keys_reg[0][52]  ( .D(n3585), .CLK(clk), .Q(\keys[0][52] ), .QN(
        n94) );
  DFFX1_HVT \keys_reg[0][51]  ( .D(n3584), .CLK(clk), .Q(\keys[0][51] ), .QN(
        n95) );
  DFFX1_HVT \keys_reg[0][50]  ( .D(n3583), .CLK(clk), .Q(\keys[0][50] ), .QN(
        n96) );
  DFFX1_HVT \keys_reg[0][49]  ( .D(n3582), .CLK(clk), .Q(\keys[0][49] ), .QN(
        n97) );
  DFFX1_HVT \keys_reg[0][48]  ( .D(n3581), .CLK(clk), .Q(\keys[0][48] ), .QN(
        n98) );
  DFFX1_HVT \keys_reg[0][47]  ( .D(n3580), .CLK(clk), .Q(\keys[0][47] ), .QN(
        n99) );
  DFFX1_HVT \keys_reg[0][46]  ( .D(n3579), .CLK(clk), .Q(\keys[0][46] ), .QN(
        n100) );
  DFFX1_HVT \keys_reg[0][45]  ( .D(n3578), .CLK(clk), .Q(\keys[0][45] ), .QN(
        n101) );
  DFFX1_HVT \keys_reg[0][44]  ( .D(n3577), .CLK(clk), .Q(\keys[0][44] ), .QN(
        n102) );
  DFFX1_HVT \keys_reg[0][43]  ( .D(n3576), .CLK(clk), .Q(\keys[0][43] ), .QN(
        n103) );
  DFFX1_HVT \keys_reg[0][42]  ( .D(n3575), .CLK(clk), .Q(\keys[0][42] ), .QN(
        n104) );
  DFFX1_HVT \keys_reg[0][41]  ( .D(n3574), .CLK(clk), .Q(\keys[0][41] ), .QN(
        n105) );
  DFFX1_HVT \keys_reg[0][40]  ( .D(n3573), .CLK(clk), .Q(\keys[0][40] ), .QN(
        n106) );
  DFFX1_HVT \keys_reg[0][39]  ( .D(n3572), .CLK(clk), .Q(\keys[0][39] ), .QN(
        n107) );
  DFFX1_HVT \keys_reg[0][38]  ( .D(n3571), .CLK(clk), .Q(\keys[0][38] ), .QN(
        n108) );
  DFFX1_HVT \keys_reg[0][37]  ( .D(n3570), .CLK(clk), .Q(\keys[0][37] ), .QN(
        n109) );
  DFFX1_HVT \keys_reg[0][36]  ( .D(n3569), .CLK(clk), .Q(\keys[0][36] ), .QN(
        n110) );
  DFFX1_HVT \keys_reg[0][35]  ( .D(n3568), .CLK(clk), .Q(\keys[0][35] ), .QN(
        n111) );
  DFFX1_HVT \keys_reg[0][34]  ( .D(n3567), .CLK(clk), .Q(\keys[0][34] ), .QN(
        n112) );
  DFFX1_HVT \keys_reg[0][33]  ( .D(n3566), .CLK(clk), .Q(\keys[0][33] ), .QN(
        n113) );
  DFFX1_HVT \keys_reg[0][32]  ( .D(n3565), .CLK(clk), .Q(\keys[0][32] ), .QN(
        n114) );
  DFFX1_HVT \keys_reg[0][31]  ( .D(n3564), .CLK(clk), .Q(\keys[0][31] ), .QN(
        n115) );
  DFFX1_HVT \keys_reg[0][30]  ( .D(n3563), .CLK(clk), .Q(\keys[0][30] ), .QN(
        n116) );
  DFFX1_HVT \keys_reg[0][29]  ( .D(n3562), .CLK(clk), .Q(\keys[0][29] ), .QN(
        n117) );
  DFFX1_HVT \keys_reg[0][28]  ( .D(n3561), .CLK(clk), .Q(\keys[0][28] ), .QN(
        n118) );
  DFFX1_HVT \keys_reg[0][27]  ( .D(n3560), .CLK(clk), .Q(\keys[0][27] ), .QN(
        n119) );
  DFFX1_HVT \keys_reg[0][26]  ( .D(n3559), .CLK(clk), .Q(\keys[0][26] ), .QN(
        n120) );
  DFFX1_HVT \keys_reg[0][25]  ( .D(n3558), .CLK(clk), .Q(\keys[0][25] ), .QN(
        n121) );
  DFFX1_HVT \keys_reg[0][24]  ( .D(n3557), .CLK(clk), .Q(\keys[0][24] ), .QN(
        n122) );
  DFFX1_HVT \keys_reg[0][23]  ( .D(n3556), .CLK(clk), .Q(\keys[0][23] ), .QN(
        n123) );
  DFFX1_HVT \keys_reg[0][22]  ( .D(n3555), .CLK(clk), .Q(\keys[0][22] ), .QN(
        n124) );
  DFFX1_HVT \keys_reg[0][21]  ( .D(n3554), .CLK(clk), .Q(\keys[0][21] ), .QN(
        n125) );
  DFFX1_HVT \keys_reg[0][20]  ( .D(n3553), .CLK(clk), .Q(\keys[0][20] ), .QN(
        n126) );
  DFFX1_HVT \keys_reg[0][19]  ( .D(n3552), .CLK(clk), .Q(\keys[0][19] ), .QN(
        n127) );
  DFFX1_HVT \keys_reg[0][18]  ( .D(n3551), .CLK(clk), .Q(\keys[0][18] ), .QN(
        n128) );
  DFFX1_HVT \keys_reg[0][17]  ( .D(n3550), .CLK(clk), .Q(\keys[0][17] ), .QN(
        n129) );
  DFFX1_HVT \keys_reg[0][16]  ( .D(n3549), .CLK(clk), .Q(\keys[0][16] ), .QN(
        n130) );
  DFFX1_HVT \keys_reg[0][15]  ( .D(n3548), .CLK(clk), .Q(\keys[0][15] ), .QN(
        n131) );
  DFFX1_HVT \keys_reg[0][14]  ( .D(n3547), .CLK(clk), .Q(\keys[0][14] ), .QN(
        n132) );
  DFFX1_HVT \keys_reg[0][13]  ( .D(n3546), .CLK(clk), .Q(\keys[0][13] ), .QN(
        n133) );
  DFFX1_HVT \keys_reg[0][12]  ( .D(n3545), .CLK(clk), .Q(\keys[0][12] ), .QN(
        n134) );
  DFFX1_HVT \keys_reg[0][11]  ( .D(n3544), .CLK(clk), .Q(\keys[0][11] ), .QN(
        n135) );
  DFFX1_HVT \keys_reg[0][10]  ( .D(n3543), .CLK(clk), .Q(\keys[0][10] ), .QN(
        n136) );
  DFFX1_HVT \keys_reg[0][9]  ( .D(n3542), .CLK(clk), .Q(\keys[0][9] ), .QN(
        n137) );
  DFFX1_HVT \keys_reg[0][8]  ( .D(n3541), .CLK(clk), .Q(\keys[0][8] ), .QN(
        n138) );
  DFFX1_HVT \keys_reg[0][7]  ( .D(n3540), .CLK(clk), .Q(\keys[0][7] ), .QN(
        n139) );
  DFFX1_HVT \keys_reg[0][6]  ( .D(n3539), .CLK(clk), .Q(\keys[0][6] ), .QN(
        n140) );
  DFFX1_HVT \keys_reg[0][5]  ( .D(n3538), .CLK(clk), .Q(\keys[0][5] ), .QN(
        n141) );
  DFFX1_HVT \keys_reg[0][4]  ( .D(n3537), .CLK(clk), .Q(\keys[0][4] ), .QN(
        n142) );
  DFFX1_HVT \keys_reg[0][3]  ( .D(n3536), .CLK(clk), .Q(\keys[0][3] ), .QN(
        n143) );
  DFFX1_HVT \keys_reg[0][2]  ( .D(n3535), .CLK(clk), .Q(\keys[0][2] ), .QN(
        n144) );
  DFFX1_HVT \keys_reg[0][1]  ( .D(n3534), .CLK(clk), .Q(\keys[0][1] ), .QN(
        n145) );
  DFFX1_HVT \keys_reg[0][0]  ( .D(n3533), .CLK(clk), .Q(\keys[0][0] ), .QN(
        n146) );
  DFFX1_HVT \keys_reg[1][127]  ( .D(n3532), .CLK(clk), .Q(\keys[1][127] ), 
        .QN(n147) );
  DFFX1_HVT \keys_reg[1][126]  ( .D(n3531), .CLK(clk), .Q(\keys[1][126] ), 
        .QN(n148) );
  DFFX1_HVT \keys_reg[1][125]  ( .D(n3530), .CLK(clk), .Q(\keys[1][125] ), 
        .QN(n149) );
  DFFX1_HVT \keys_reg[1][124]  ( .D(n3529), .CLK(clk), .Q(\keys[1][124] ), 
        .QN(n150) );
  DFFX1_HVT \keys_reg[1][123]  ( .D(n3528), .CLK(clk), .Q(\keys[1][123] ), 
        .QN(n151) );
  DFFX1_HVT \keys_reg[1][122]  ( .D(n3527), .CLK(clk), .Q(\keys[1][122] ), 
        .QN(n152) );
  DFFX1_HVT \keys_reg[1][121]  ( .D(n3526), .CLK(clk), .Q(\keys[1][121] ), 
        .QN(n153) );
  DFFX1_HVT \keys_reg[1][120]  ( .D(n3525), .CLK(clk), .Q(\keys[1][120] ), 
        .QN(n154) );
  DFFX1_HVT \keys_reg[1][119]  ( .D(n3524), .CLK(clk), .Q(\keys[1][119] ), 
        .QN(n155) );
  DFFX1_HVT \keys_reg[1][118]  ( .D(n3523), .CLK(clk), .Q(\keys[1][118] ), 
        .QN(n156) );
  DFFX1_HVT \keys_reg[1][117]  ( .D(n3522), .CLK(clk), .Q(\keys[1][117] ), 
        .QN(n157) );
  DFFX1_HVT \keys_reg[1][116]  ( .D(n3521), .CLK(clk), .Q(\keys[1][116] ), 
        .QN(n158) );
  DFFX1_HVT \keys_reg[1][115]  ( .D(n3520), .CLK(clk), .Q(\keys[1][115] ), 
        .QN(n159) );
  DFFX1_HVT \keys_reg[1][114]  ( .D(n3519), .CLK(clk), .Q(\keys[1][114] ), 
        .QN(n160) );
  DFFX1_HVT \keys_reg[1][113]  ( .D(n3518), .CLK(clk), .Q(\keys[1][113] ), 
        .QN(n161) );
  DFFX1_HVT \keys_reg[1][112]  ( .D(n3517), .CLK(clk), .Q(\keys[1][112] ), 
        .QN(n162) );
  DFFX1_HVT \keys_reg[1][111]  ( .D(n3516), .CLK(clk), .Q(\keys[1][111] ), 
        .QN(n163) );
  DFFX1_HVT \keys_reg[1][110]  ( .D(n3515), .CLK(clk), .Q(\keys[1][110] ), 
        .QN(n164) );
  DFFX1_HVT \keys_reg[1][109]  ( .D(n3514), .CLK(clk), .Q(\keys[1][109] ), 
        .QN(n165) );
  DFFX1_HVT \keys_reg[1][108]  ( .D(n3513), .CLK(clk), .Q(\keys[1][108] ), 
        .QN(n166) );
  DFFX1_HVT \keys_reg[1][107]  ( .D(n3512), .CLK(clk), .Q(\keys[1][107] ), 
        .QN(n167) );
  DFFX1_HVT \keys_reg[1][106]  ( .D(n3511), .CLK(clk), .Q(\keys[1][106] ), 
        .QN(n168) );
  DFFX1_HVT \keys_reg[1][105]  ( .D(n3510), .CLK(clk), .Q(\keys[1][105] ), 
        .QN(n169) );
  DFFX1_HVT \keys_reg[1][104]  ( .D(n3509), .CLK(clk), .Q(\keys[1][104] ), 
        .QN(n170) );
  DFFX1_HVT \keys_reg[1][103]  ( .D(n3508), .CLK(clk), .Q(\keys[1][103] ), 
        .QN(n171) );
  DFFX1_HVT \keys_reg[1][102]  ( .D(n3507), .CLK(clk), .Q(\keys[1][102] ), 
        .QN(n172) );
  DFFX1_HVT \keys_reg[1][101]  ( .D(n3506), .CLK(clk), .Q(\keys[1][101] ), 
        .QN(n173) );
  DFFX1_HVT \keys_reg[1][100]  ( .D(n3505), .CLK(clk), .Q(\keys[1][100] ), 
        .QN(n174) );
  DFFX1_HVT \keys_reg[1][99]  ( .D(n3504), .CLK(clk), .Q(\keys[1][99] ), .QN(
        n175) );
  DFFX1_HVT \keys_reg[1][98]  ( .D(n3503), .CLK(clk), .Q(\keys[1][98] ), .QN(
        n176) );
  DFFX1_HVT \keys_reg[1][97]  ( .D(n3502), .CLK(clk), .Q(\keys[1][97] ), .QN(
        n177) );
  DFFX1_HVT \keys_reg[1][96]  ( .D(n3501), .CLK(clk), .Q(\keys[1][96] ), .QN(
        n178) );
  DFFX1_HVT \keys_reg[1][95]  ( .D(n3500), .CLK(clk), .Q(\keys[1][95] ), .QN(
        n179) );
  DFFX1_HVT \keys_reg[1][94]  ( .D(n3499), .CLK(clk), .Q(\keys[1][94] ), .QN(
        n180) );
  DFFX1_HVT \keys_reg[1][93]  ( .D(n3498), .CLK(clk), .Q(\keys[1][93] ), .QN(
        n181) );
  DFFX1_HVT \keys_reg[1][92]  ( .D(n3497), .CLK(clk), .Q(\keys[1][92] ), .QN(
        n182) );
  DFFX1_HVT \keys_reg[1][91]  ( .D(n3496), .CLK(clk), .Q(\keys[1][91] ), .QN(
        n183) );
  DFFX1_HVT \keys_reg[1][90]  ( .D(n3495), .CLK(clk), .Q(\keys[1][90] ), .QN(
        n184) );
  DFFX1_HVT \keys_reg[1][89]  ( .D(n3494), .CLK(clk), .Q(\keys[1][89] ), .QN(
        n185) );
  DFFX1_HVT \keys_reg[1][88]  ( .D(n3493), .CLK(clk), .Q(\keys[1][88] ), .QN(
        n186) );
  DFFX1_HVT \keys_reg[1][87]  ( .D(n3492), .CLK(clk), .Q(\keys[1][87] ), .QN(
        n187) );
  DFFX1_HVT \keys_reg[1][86]  ( .D(n3491), .CLK(clk), .Q(\keys[1][86] ), .QN(
        n188) );
  DFFX1_HVT \keys_reg[1][85]  ( .D(n3490), .CLK(clk), .Q(\keys[1][85] ), .QN(
        n189) );
  DFFX1_HVT \keys_reg[1][84]  ( .D(n3489), .CLK(clk), .Q(\keys[1][84] ), .QN(
        n190) );
  DFFX1_HVT \keys_reg[1][83]  ( .D(n3488), .CLK(clk), .Q(\keys[1][83] ), .QN(
        n191) );
  DFFX1_HVT \keys_reg[1][82]  ( .D(n3487), .CLK(clk), .Q(\keys[1][82] ), .QN(
        n192) );
  DFFX1_HVT \keys_reg[1][81]  ( .D(n3486), .CLK(clk), .Q(\keys[1][81] ), .QN(
        n193) );
  DFFX1_HVT \keys_reg[1][80]  ( .D(n3485), .CLK(clk), .Q(\keys[1][80] ), .QN(
        n194) );
  DFFX1_HVT \keys_reg[1][79]  ( .D(n3484), .CLK(clk), .Q(\keys[1][79] ), .QN(
        n195) );
  DFFX1_HVT \keys_reg[1][78]  ( .D(n3483), .CLK(clk), .Q(\keys[1][78] ), .QN(
        n196) );
  DFFX1_HVT \keys_reg[1][77]  ( .D(n3482), .CLK(clk), .Q(\keys[1][77] ), .QN(
        n197) );
  DFFX1_HVT \keys_reg[1][76]  ( .D(n3481), .CLK(clk), .Q(\keys[1][76] ), .QN(
        n198) );
  DFFX1_HVT \keys_reg[1][75]  ( .D(n3480), .CLK(clk), .Q(\keys[1][75] ), .QN(
        n199) );
  DFFX1_HVT \keys_reg[1][74]  ( .D(n3479), .CLK(clk), .Q(\keys[1][74] ), .QN(
        n200) );
  DFFX1_HVT \keys_reg[1][73]  ( .D(n3478), .CLK(clk), .Q(\keys[1][73] ), .QN(
        n201) );
  DFFX1_HVT \keys_reg[1][72]  ( .D(n3477), .CLK(clk), .Q(\keys[1][72] ), .QN(
        n202) );
  DFFX1_HVT \keys_reg[1][71]  ( .D(n3476), .CLK(clk), .Q(\keys[1][71] ), .QN(
        n203) );
  DFFX1_HVT \keys_reg[1][70]  ( .D(n3475), .CLK(clk), .Q(\keys[1][70] ), .QN(
        n204) );
  DFFX1_HVT \keys_reg[1][69]  ( .D(n3474), .CLK(clk), .Q(\keys[1][69] ), .QN(
        n205) );
  DFFX1_HVT \keys_reg[1][68]  ( .D(n3473), .CLK(clk), .Q(\keys[1][68] ), .QN(
        n206) );
  DFFX1_HVT \keys_reg[1][67]  ( .D(n3472), .CLK(clk), .Q(\keys[1][67] ), .QN(
        n207) );
  DFFX1_HVT \keys_reg[1][66]  ( .D(n3471), .CLK(clk), .Q(\keys[1][66] ), .QN(
        n208) );
  DFFX1_HVT \keys_reg[1][65]  ( .D(n3470), .CLK(clk), .Q(\keys[1][65] ), .QN(
        n209) );
  DFFX1_HVT \keys_reg[1][64]  ( .D(n3469), .CLK(clk), .Q(\keys[1][64] ), .QN(
        n210) );
  DFFX1_HVT \keys_reg[1][63]  ( .D(n3468), .CLK(clk), .Q(\keys[1][63] ), .QN(
        n211) );
  DFFX1_HVT \keys_reg[1][62]  ( .D(n3467), .CLK(clk), .Q(\keys[1][62] ), .QN(
        n212) );
  DFFX1_HVT \keys_reg[1][61]  ( .D(n3466), .CLK(clk), .Q(\keys[1][61] ), .QN(
        n213) );
  DFFX1_HVT \keys_reg[1][60]  ( .D(n3465), .CLK(clk), .Q(\keys[1][60] ), .QN(
        n214) );
  DFFX1_HVT \keys_reg[1][59]  ( .D(n3464), .CLK(clk), .Q(\keys[1][59] ), .QN(
        n215) );
  DFFX1_HVT \keys_reg[1][58]  ( .D(n3463), .CLK(clk), .Q(\keys[1][58] ), .QN(
        n216) );
  DFFX1_HVT \keys_reg[1][57]  ( .D(n3462), .CLK(clk), .Q(\keys[1][57] ), .QN(
        n217) );
  DFFX1_HVT \keys_reg[1][56]  ( .D(n3461), .CLK(clk), .Q(\keys[1][56] ), .QN(
        n218) );
  DFFX1_HVT \keys_reg[1][55]  ( .D(n3460), .CLK(clk), .Q(\keys[1][55] ), .QN(
        n219) );
  DFFX1_HVT \keys_reg[1][54]  ( .D(n3459), .CLK(clk), .Q(\keys[1][54] ), .QN(
        n220) );
  DFFX1_HVT \keys_reg[1][53]  ( .D(n3458), .CLK(clk), .Q(\keys[1][53] ), .QN(
        n221) );
  DFFX1_HVT \keys_reg[1][52]  ( .D(n3457), .CLK(clk), .Q(\keys[1][52] ), .QN(
        n222) );
  DFFX1_HVT \keys_reg[1][51]  ( .D(n3456), .CLK(clk), .Q(\keys[1][51] ), .QN(
        n223) );
  DFFX1_HVT \keys_reg[1][50]  ( .D(n3455), .CLK(clk), .Q(\keys[1][50] ), .QN(
        n224) );
  DFFX1_HVT \keys_reg[1][49]  ( .D(n3454), .CLK(clk), .Q(\keys[1][49] ), .QN(
        n225) );
  DFFX1_HVT \keys_reg[1][48]  ( .D(n3453), .CLK(clk), .Q(\keys[1][48] ), .QN(
        n226) );
  DFFX1_HVT \keys_reg[1][47]  ( .D(n3452), .CLK(clk), .Q(\keys[1][47] ), .QN(
        n227) );
  DFFX1_HVT \keys_reg[1][46]  ( .D(n3451), .CLK(clk), .Q(\keys[1][46] ), .QN(
        n228) );
  DFFX1_HVT \keys_reg[1][45]  ( .D(n3450), .CLK(clk), .Q(\keys[1][45] ), .QN(
        n229) );
  DFFX1_HVT \keys_reg[1][44]  ( .D(n3449), .CLK(clk), .Q(\keys[1][44] ), .QN(
        n230) );
  DFFX1_HVT \keys_reg[1][43]  ( .D(n3448), .CLK(clk), .QN(n231) );
  DFFX1_HVT \keys_reg[1][42]  ( .D(n3447), .CLK(clk), .Q(\keys[1][42] ), .QN(
        n232) );
  DFFX1_HVT \keys_reg[1][41]  ( .D(n3446), .CLK(clk), .Q(\keys[1][41] ), .QN(
        n233) );
  DFFX1_HVT \keys_reg[1][40]  ( .D(n3445), .CLK(clk), .Q(\keys[1][40] ), .QN(
        n234) );
  DFFX1_HVT \keys_reg[1][39]  ( .D(n3444), .CLK(clk), .Q(\keys[1][39] ), .QN(
        n235) );
  DFFX1_HVT \keys_reg[1][38]  ( .D(n3443), .CLK(clk), .Q(\keys[1][38] ), .QN(
        n236) );
  DFFX1_HVT \keys_reg[1][37]  ( .D(n3442), .CLK(clk), .Q(\keys[1][37] ), .QN(
        n237) );
  DFFX1_HVT \keys_reg[1][36]  ( .D(n3441), .CLK(clk), .Q(\keys[1][36] ), .QN(
        n238) );
  DFFX1_HVT \keys_reg[1][35]  ( .D(n3440), .CLK(clk), .Q(\keys[1][35] ), .QN(
        n239) );
  DFFX1_HVT \keys_reg[1][34]  ( .D(n3439), .CLK(clk), .Q(\keys[1][34] ), .QN(
        n240) );
  DFFX1_HVT \keys_reg[1][33]  ( .D(n3438), .CLK(clk), .Q(\keys[1][33] ), .QN(
        n241) );
  DFFX1_HVT \keys_reg[1][32]  ( .D(n3437), .CLK(clk), .Q(\keys[1][32] ), .QN(
        n242) );
  DFFX1_HVT \keys_reg[1][31]  ( .D(n3436), .CLK(clk), .Q(\keys[1][31] ), .QN(
        n243) );
  DFFX1_HVT \keys_reg[1][30]  ( .D(n3435), .CLK(clk), .Q(\keys[1][30] ), .QN(
        n244) );
  DFFX1_HVT \keys_reg[1][29]  ( .D(n3434), .CLK(clk), .Q(\keys[1][29] ), .QN(
        n245) );
  DFFX1_HVT \keys_reg[1][28]  ( .D(n3433), .CLK(clk), .Q(\keys[1][28] ), .QN(
        n246) );
  DFFX1_HVT \keys_reg[1][27]  ( .D(n3432), .CLK(clk), .Q(\keys[1][27] ), .QN(
        n247) );
  DFFX1_HVT \keys_reg[1][26]  ( .D(n3431), .CLK(clk), .Q(\keys[1][26] ), .QN(
        n248) );
  DFFX1_HVT \keys_reg[1][25]  ( .D(n3430), .CLK(clk), .Q(\keys[1][25] ), .QN(
        n249) );
  DFFX1_HVT \keys_reg[1][24]  ( .D(n3429), .CLK(clk), .Q(\keys[1][24] ), .QN(
        n250) );
  DFFX1_HVT \keys_reg[1][23]  ( .D(n3428), .CLK(clk), .Q(\keys[1][23] ), .QN(
        n251) );
  DFFX1_HVT \keys_reg[1][22]  ( .D(n3427), .CLK(clk), .Q(\keys[1][22] ), .QN(
        n252) );
  DFFX1_HVT \keys_reg[1][21]  ( .D(n3426), .CLK(clk), .Q(\keys[1][21] ), .QN(
        n253) );
  DFFX1_HVT \keys_reg[1][20]  ( .D(n3425), .CLK(clk), .Q(\keys[1][20] ), .QN(
        n254) );
  DFFX1_HVT \keys_reg[1][19]  ( .D(n3424), .CLK(clk), .Q(\keys[1][19] ), .QN(
        n255) );
  DFFX1_HVT \keys_reg[1][18]  ( .D(n3423), .CLK(clk), .Q(\keys[1][18] ), .QN(
        n256) );
  DFFX1_HVT \keys_reg[1][17]  ( .D(n3422), .CLK(clk), .Q(\keys[1][17] ), .QN(
        n257) );
  DFFX1_HVT \keys_reg[1][16]  ( .D(n3421), .CLK(clk), .Q(\keys[1][16] ), .QN(
        n258) );
  DFFX1_HVT \keys_reg[1][15]  ( .D(n3420), .CLK(clk), .Q(\keys[1][15] ), .QN(
        n259) );
  DFFX1_HVT \keys_reg[1][14]  ( .D(n3419), .CLK(clk), .Q(\keys[1][14] ), .QN(
        n260) );
  DFFX1_HVT \keys_reg[1][13]  ( .D(n3418), .CLK(clk), .Q(\keys[1][13] ), .QN(
        n261) );
  DFFX1_HVT \keys_reg[1][12]  ( .D(n3417), .CLK(clk), .Q(\keys[1][12] ), .QN(
        n262) );
  DFFX1_HVT \keys_reg[1][11]  ( .D(n3416), .CLK(clk), .Q(\keys[1][11] ), .QN(
        n263) );
  DFFX1_HVT \keys_reg[1][10]  ( .D(n3415), .CLK(clk), .Q(\keys[1][10] ), .QN(
        n264) );
  DFFX1_HVT \keys_reg[1][9]  ( .D(n3414), .CLK(clk), .Q(\keys[1][9] ), .QN(
        n265) );
  DFFX1_HVT \keys_reg[1][8]  ( .D(n3413), .CLK(clk), .Q(\keys[1][8] ), .QN(
        n266) );
  DFFX1_HVT \keys_reg[1][7]  ( .D(n3412), .CLK(clk), .Q(\keys[1][7] ), .QN(
        n267) );
  DFFX1_HVT \keys_reg[1][6]  ( .D(n3411), .CLK(clk), .Q(\keys[1][6] ), .QN(
        n268) );
  DFFX1_HVT \keys_reg[1][5]  ( .D(n3410), .CLK(clk), .Q(\keys[1][5] ), .QN(
        n269) );
  DFFX1_HVT \keys_reg[1][4]  ( .D(n3409), .CLK(clk), .Q(\keys[1][4] ), .QN(
        n270) );
  DFFX1_HVT \keys_reg[1][3]  ( .D(n3408), .CLK(clk), .Q(\keys[1][3] ), .QN(
        n271) );
  DFFX1_HVT \keys_reg[1][2]  ( .D(n3407), .CLK(clk), .Q(\keys[1][2] ), .QN(
        n272) );
  DFFX1_HVT \keys_reg[1][1]  ( .D(n3406), .CLK(clk), .Q(\keys[1][1] ), .QN(
        n273) );
  DFFX1_HVT \keys_reg[1][0]  ( .D(n3405), .CLK(clk), .Q(\keys[1][0] ), .QN(
        n274) );
  DFFX1_HVT \keys_reg[2][127]  ( .D(n3404), .CLK(clk), .Q(\keys[2][127] ), 
        .QN(n275) );
  DFFX1_HVT \keys_reg[2][126]  ( .D(n3403), .CLK(clk), .Q(\keys[2][126] ), 
        .QN(n276) );
  DFFX1_HVT \keys_reg[2][125]  ( .D(n3402), .CLK(clk), .Q(\keys[2][125] ), 
        .QN(n277) );
  DFFX1_HVT \keys_reg[2][124]  ( .D(n3401), .CLK(clk), .Q(\keys[2][124] ), 
        .QN(n278) );
  DFFX1_HVT \keys_reg[2][123]  ( .D(n3400), .CLK(clk), .Q(\keys[2][123] ), 
        .QN(n279) );
  DFFX1_HVT \keys_reg[2][122]  ( .D(n3399), .CLK(clk), .Q(\keys[2][122] ), 
        .QN(n280) );
  DFFX1_HVT \keys_reg[2][121]  ( .D(n3398), .CLK(clk), .Q(\keys[2][121] ), 
        .QN(n281) );
  DFFX1_HVT \keys_reg[2][120]  ( .D(n3397), .CLK(clk), .Q(\keys[2][120] ), 
        .QN(n282) );
  DFFX1_HVT \keys_reg[2][119]  ( .D(n3396), .CLK(clk), .Q(\keys[2][119] ), 
        .QN(n283) );
  DFFX1_HVT \keys_reg[2][118]  ( .D(n3395), .CLK(clk), .Q(\keys[2][118] ), 
        .QN(n284) );
  DFFX1_HVT \keys_reg[2][117]  ( .D(n3394), .CLK(clk), .Q(\keys[2][117] ), 
        .QN(n285) );
  DFFX1_HVT \keys_reg[2][116]  ( .D(n3393), .CLK(clk), .Q(\keys[2][116] ), 
        .QN(n286) );
  DFFX1_HVT \keys_reg[2][115]  ( .D(n3392), .CLK(clk), .Q(\keys[2][115] ), 
        .QN(n287) );
  DFFX1_HVT \keys_reg[2][114]  ( .D(n3391), .CLK(clk), .Q(\keys[2][114] ), 
        .QN(n288) );
  DFFX1_HVT \keys_reg[2][113]  ( .D(n3390), .CLK(clk), .Q(\keys[2][113] ), 
        .QN(n289) );
  DFFX1_HVT \keys_reg[2][112]  ( .D(n3389), .CLK(clk), .Q(\keys[2][112] ), 
        .QN(n290) );
  DFFX1_HVT \keys_reg[2][111]  ( .D(n3388), .CLK(clk), .Q(\keys[2][111] ), 
        .QN(n291) );
  DFFX1_HVT \keys_reg[2][110]  ( .D(n3387), .CLK(clk), .Q(\keys[2][110] ), 
        .QN(n292) );
  DFFX1_HVT \keys_reg[2][109]  ( .D(n3386), .CLK(clk), .Q(\keys[2][109] ), 
        .QN(n293) );
  DFFX1_HVT \keys_reg[2][108]  ( .D(n3385), .CLK(clk), .Q(\keys[2][108] ), 
        .QN(n294) );
  DFFX1_HVT \keys_reg[2][107]  ( .D(n3384), .CLK(clk), .Q(\keys[2][107] ), 
        .QN(n295) );
  DFFX1_HVT \keys_reg[2][106]  ( .D(n3383), .CLK(clk), .Q(\keys[2][106] ), 
        .QN(n296) );
  DFFX1_HVT \keys_reg[2][105]  ( .D(n3382), .CLK(clk), .Q(\keys[2][105] ), 
        .QN(n297) );
  DFFX1_HVT \keys_reg[2][104]  ( .D(n3381), .CLK(clk), .Q(\keys[2][104] ), 
        .QN(n298) );
  DFFX1_HVT \keys_reg[2][103]  ( .D(n3380), .CLK(clk), .Q(\keys[2][103] ), 
        .QN(n299) );
  DFFX1_HVT \keys_reg[2][102]  ( .D(n3379), .CLK(clk), .Q(\keys[2][102] ), 
        .QN(n300) );
  DFFX1_HVT \keys_reg[2][101]  ( .D(n3378), .CLK(clk), .Q(\keys[2][101] ), 
        .QN(n301) );
  DFFX1_HVT \keys_reg[2][100]  ( .D(n3377), .CLK(clk), .Q(\keys[2][100] ), 
        .QN(n302) );
  DFFX1_HVT \keys_reg[2][99]  ( .D(n3376), .CLK(clk), .Q(\keys[2][99] ), .QN(
        n303) );
  DFFX1_HVT \keys_reg[2][98]  ( .D(n3375), .CLK(clk), .Q(\keys[2][98] ), .QN(
        n304) );
  DFFX1_HVT \keys_reg[2][97]  ( .D(n3374), .CLK(clk), .Q(\keys[2][97] ), .QN(
        n305) );
  DFFX1_HVT \keys_reg[2][96]  ( .D(n3373), .CLK(clk), .Q(\keys[2][96] ), .QN(
        n306) );
  DFFX1_HVT \keys_reg[2][95]  ( .D(n3372), .CLK(clk), .Q(\keys[2][95] ), .QN(
        n307) );
  DFFX1_HVT \keys_reg[2][94]  ( .D(n3371), .CLK(clk), .Q(\keys[2][94] ), .QN(
        n308) );
  DFFX1_HVT \keys_reg[2][93]  ( .D(n3370), .CLK(clk), .Q(\keys[2][93] ), .QN(
        n309) );
  DFFX1_HVT \keys_reg[2][92]  ( .D(n3369), .CLK(clk), .Q(\keys[2][92] ), .QN(
        n310) );
  DFFX1_HVT \keys_reg[2][91]  ( .D(n3368), .CLK(clk), .Q(\keys[2][91] ), .QN(
        n311) );
  DFFX1_HVT \keys_reg[2][90]  ( .D(n3367), .CLK(clk), .Q(\keys[2][90] ), .QN(
        n312) );
  DFFX1_HVT \keys_reg[2][89]  ( .D(n3366), .CLK(clk), .Q(\keys[2][89] ), .QN(
        n313) );
  DFFX1_HVT \keys_reg[2][88]  ( .D(n3365), .CLK(clk), .Q(\keys[2][88] ), .QN(
        n314) );
  DFFX1_HVT \keys_reg[2][87]  ( .D(n3364), .CLK(clk), .Q(\keys[2][87] ), .QN(
        n315) );
  DFFX1_HVT \keys_reg[2][86]  ( .D(n3363), .CLK(clk), .Q(\keys[2][86] ), .QN(
        n316) );
  DFFX1_HVT \keys_reg[2][85]  ( .D(n3362), .CLK(clk), .Q(\keys[2][85] ), .QN(
        n317) );
  DFFX1_HVT \keys_reg[2][84]  ( .D(n3361), .CLK(clk), .Q(\keys[2][84] ), .QN(
        n318) );
  DFFX1_HVT \keys_reg[2][83]  ( .D(n3360), .CLK(clk), .Q(\keys[2][83] ), .QN(
        n319) );
  DFFX1_HVT \keys_reg[2][82]  ( .D(n3359), .CLK(clk), .Q(\keys[2][82] ), .QN(
        n320) );
  DFFX1_HVT \keys_reg[2][81]  ( .D(n3358), .CLK(clk), .Q(\keys[2][81] ), .QN(
        n321) );
  DFFX1_HVT \keys_reg[2][80]  ( .D(n3357), .CLK(clk), .Q(\keys[2][80] ), .QN(
        n322) );
  DFFX1_HVT \keys_reg[2][79]  ( .D(n3356), .CLK(clk), .Q(\keys[2][79] ), .QN(
        n323) );
  DFFX1_HVT \keys_reg[2][78]  ( .D(n3355), .CLK(clk), .Q(\keys[2][78] ), .QN(
        n324) );
  DFFX1_HVT \keys_reg[2][77]  ( .D(n3354), .CLK(clk), .Q(\keys[2][77] ), .QN(
        n325) );
  DFFX1_HVT \keys_reg[2][76]  ( .D(n3353), .CLK(clk), .Q(\keys[2][76] ), .QN(
        n326) );
  DFFX1_HVT \keys_reg[2][75]  ( .D(n3352), .CLK(clk), .Q(\keys[2][75] ), .QN(
        n327) );
  DFFX1_HVT \keys_reg[2][74]  ( .D(n3351), .CLK(clk), .Q(\keys[2][74] ), .QN(
        n328) );
  DFFX1_HVT \keys_reg[2][73]  ( .D(n3350), .CLK(clk), .Q(\keys[2][73] ), .QN(
        n329) );
  DFFX1_HVT \keys_reg[2][72]  ( .D(n3349), .CLK(clk), .Q(\keys[2][72] ), .QN(
        n330) );
  DFFX1_HVT \keys_reg[2][71]  ( .D(n3348), .CLK(clk), .Q(\keys[2][71] ), .QN(
        n331) );
  DFFX1_HVT \keys_reg[2][70]  ( .D(n3347), .CLK(clk), .Q(\keys[2][70] ), .QN(
        n332) );
  DFFX1_HVT \keys_reg[2][69]  ( .D(n3346), .CLK(clk), .Q(\keys[2][69] ), .QN(
        n333) );
  DFFX1_HVT \keys_reg[2][68]  ( .D(n3345), .CLK(clk), .Q(\keys[2][68] ), .QN(
        n334) );
  DFFX1_HVT \keys_reg[2][67]  ( .D(n3344), .CLK(clk), .Q(\keys[2][67] ), .QN(
        n335) );
  DFFX1_HVT \keys_reg[2][66]  ( .D(n3343), .CLK(clk), .Q(\keys[2][66] ), .QN(
        n336) );
  DFFX1_HVT \keys_reg[2][65]  ( .D(n3342), .CLK(clk), .Q(\keys[2][65] ), .QN(
        n337) );
  DFFX1_HVT \keys_reg[2][64]  ( .D(n3341), .CLK(clk), .Q(\keys[2][64] ), .QN(
        n338) );
  DFFX1_HVT \keys_reg[2][63]  ( .D(n3340), .CLK(clk), .Q(\keys[2][63] ), .QN(
        n339) );
  DFFX1_HVT \keys_reg[2][62]  ( .D(n3339), .CLK(clk), .Q(\keys[2][62] ), .QN(
        n340) );
  DFFX1_HVT \keys_reg[2][61]  ( .D(n3338), .CLK(clk), .Q(\keys[2][61] ), .QN(
        n341) );
  DFFX1_HVT \keys_reg[2][60]  ( .D(n3337), .CLK(clk), .Q(\keys[2][60] ), .QN(
        n342) );
  DFFX1_HVT \keys_reg[2][59]  ( .D(n3336), .CLK(clk), .Q(\keys[2][59] ), .QN(
        n343) );
  DFFX1_HVT \keys_reg[2][58]  ( .D(n3335), .CLK(clk), .Q(\keys[2][58] ), .QN(
        n344) );
  DFFX1_HVT \keys_reg[2][57]  ( .D(n3334), .CLK(clk), .Q(\keys[2][57] ), .QN(
        n345) );
  DFFX1_HVT \keys_reg[2][56]  ( .D(n3333), .CLK(clk), .Q(\keys[2][56] ), .QN(
        n346) );
  DFFX1_HVT \keys_reg[2][55]  ( .D(n3332), .CLK(clk), .Q(\keys[2][55] ), .QN(
        n347) );
  DFFX1_HVT \keys_reg[2][54]  ( .D(n3331), .CLK(clk), .Q(\keys[2][54] ), .QN(
        n348) );
  DFFX1_HVT \keys_reg[2][53]  ( .D(n3330), .CLK(clk), .Q(\keys[2][53] ), .QN(
        n349) );
  DFFX1_HVT \keys_reg[2][52]  ( .D(n3329), .CLK(clk), .Q(\keys[2][52] ), .QN(
        n350) );
  DFFX1_HVT \keys_reg[2][51]  ( .D(n3328), .CLK(clk), .Q(\keys[2][51] ), .QN(
        n351) );
  DFFX1_HVT \keys_reg[2][50]  ( .D(n3327), .CLK(clk), .Q(\keys[2][50] ), .QN(
        n352) );
  DFFX1_HVT \keys_reg[2][49]  ( .D(n3326), .CLK(clk), .Q(\keys[2][49] ), .QN(
        n353) );
  DFFX1_HVT \keys_reg[2][48]  ( .D(n3325), .CLK(clk), .Q(\keys[2][48] ), .QN(
        n354) );
  DFFX1_HVT \keys_reg[2][47]  ( .D(n3324), .CLK(clk), .QN(n355) );
  DFFX1_HVT \keys_reg[2][46]  ( .D(n3323), .CLK(clk), .Q(\keys[2][46] ), .QN(
        n356) );
  DFFX1_HVT \keys_reg[2][45]  ( .D(n3322), .CLK(clk), .QN(n357) );
  DFFX1_HVT \keys_reg[2][44]  ( .D(n3321), .CLK(clk), .Q(\keys[2][44] ), .QN(
        n358) );
  DFFX1_HVT \keys_reg[2][43]  ( .D(n3320), .CLK(clk), .Q(\keys[2][43] ), .QN(
        n359) );
  DFFX1_HVT \keys_reg[2][42]  ( .D(n3319), .CLK(clk), .Q(\keys[2][42] ), .QN(
        n360) );
  DFFX1_HVT \keys_reg[2][41]  ( .D(n3318), .CLK(clk), .QN(n361) );
  DFFX1_HVT \keys_reg[2][40]  ( .D(n3317), .CLK(clk), .Q(\keys[2][40] ), .QN(
        n362) );
  DFFX1_HVT \keys_reg[2][39]  ( .D(n3316), .CLK(clk), .Q(\keys[2][39] ), .QN(
        n363) );
  DFFX1_HVT \keys_reg[2][38]  ( .D(n3315), .CLK(clk), .Q(\keys[2][38] ), .QN(
        n364) );
  DFFX1_HVT \keys_reg[2][37]  ( .D(n3314), .CLK(clk), .Q(\keys[2][37] ), .QN(
        n365) );
  DFFX1_HVT \keys_reg[2][36]  ( .D(n3313), .CLK(clk), .Q(\keys[2][36] ), .QN(
        n366) );
  DFFX1_HVT \keys_reg[2][35]  ( .D(n3312), .CLK(clk), .Q(\keys[2][35] ), .QN(
        n367) );
  DFFX1_HVT \keys_reg[2][34]  ( .D(n3311), .CLK(clk), .Q(\keys[2][34] ), .QN(
        n368) );
  DFFX1_HVT \keys_reg[2][33]  ( .D(n3310), .CLK(clk), .Q(\keys[2][33] ), .QN(
        n369) );
  DFFX1_HVT \keys_reg[2][32]  ( .D(n3309), .CLK(clk), .Q(\keys[2][32] ), .QN(
        n370) );
  DFFX1_HVT \keys_reg[2][31]  ( .D(n3308), .CLK(clk), .Q(\keys[2][31] ), .QN(
        n371) );
  DFFX1_HVT \keys_reg[2][30]  ( .D(n3307), .CLK(clk), .Q(\keys[2][30] ), .QN(
        n372) );
  DFFX1_HVT \keys_reg[2][29]  ( .D(n3306), .CLK(clk), .Q(\keys[2][29] ), .QN(
        n373) );
  DFFX1_HVT \keys_reg[2][28]  ( .D(n3305), .CLK(clk), .Q(\keys[2][28] ), .QN(
        n374) );
  DFFX1_HVT \keys_reg[2][27]  ( .D(n3304), .CLK(clk), .Q(\keys[2][27] ), .QN(
        n375) );
  DFFX1_HVT \keys_reg[2][26]  ( .D(n3303), .CLK(clk), .Q(\keys[2][26] ), .QN(
        n376) );
  DFFX1_HVT \keys_reg[2][25]  ( .D(n3302), .CLK(clk), .Q(\keys[2][25] ), .QN(
        n377) );
  DFFX1_HVT \keys_reg[2][24]  ( .D(n3301), .CLK(clk), .Q(\keys[2][24] ), .QN(
        n378) );
  DFFX1_HVT \keys_reg[2][23]  ( .D(n3300), .CLK(clk), .Q(\keys[2][23] ), .QN(
        n379) );
  DFFX1_HVT \keys_reg[2][22]  ( .D(n3299), .CLK(clk), .Q(\keys[2][22] ), .QN(
        n380) );
  DFFX1_HVT \keys_reg[2][21]  ( .D(n3298), .CLK(clk), .Q(\keys[2][21] ), .QN(
        n381) );
  DFFX1_HVT \keys_reg[2][20]  ( .D(n3297), .CLK(clk), .Q(\keys[2][20] ), .QN(
        n382) );
  DFFX1_HVT \keys_reg[2][19]  ( .D(n3296), .CLK(clk), .Q(\keys[2][19] ), .QN(
        n383) );
  DFFX1_HVT \keys_reg[2][18]  ( .D(n3295), .CLK(clk), .Q(\keys[2][18] ), .QN(
        n384) );
  DFFX1_HVT \keys_reg[2][17]  ( .D(n3294), .CLK(clk), .Q(\keys[2][17] ), .QN(
        n385) );
  DFFX1_HVT \keys_reg[2][16]  ( .D(n3293), .CLK(clk), .Q(\keys[2][16] ), .QN(
        n386) );
  DFFX1_HVT \keys_reg[2][15]  ( .D(n3292), .CLK(clk), .Q(\keys[2][15] ), .QN(
        n387) );
  DFFX1_HVT \keys_reg[2][14]  ( .D(n3291), .CLK(clk), .Q(\keys[2][14] ), .QN(
        n388) );
  DFFX1_HVT \keys_reg[2][13]  ( .D(n3290), .CLK(clk), .Q(\keys[2][13] ), .QN(
        n389) );
  DFFX1_HVT \keys_reg[2][12]  ( .D(n3289), .CLK(clk), .Q(\keys[2][12] ), .QN(
        n390) );
  DFFX1_HVT \keys_reg[2][11]  ( .D(n3288), .CLK(clk), .Q(\keys[2][11] ), .QN(
        n391) );
  DFFX1_HVT \keys_reg[2][10]  ( .D(n3287), .CLK(clk), .Q(\keys[2][10] ), .QN(
        n392) );
  DFFX1_HVT \keys_reg[2][9]  ( .D(n3286), .CLK(clk), .Q(\keys[2][9] ), .QN(
        n393) );
  DFFX1_HVT \keys_reg[2][8]  ( .D(n3285), .CLK(clk), .Q(\keys[2][8] ), .QN(
        n394) );
  DFFX1_HVT \keys_reg[2][7]  ( .D(n3284), .CLK(clk), .Q(\keys[2][7] ), .QN(
        n395) );
  DFFX1_HVT \keys_reg[2][6]  ( .D(n3283), .CLK(clk), .Q(\keys[2][6] ), .QN(
        n396) );
  DFFX1_HVT \keys_reg[2][5]  ( .D(n3282), .CLK(clk), .Q(\keys[2][5] ), .QN(
        n397) );
  DFFX1_HVT \keys_reg[2][4]  ( .D(n3281), .CLK(clk), .Q(\keys[2][4] ), .QN(
        n398) );
  DFFX1_HVT \keys_reg[2][3]  ( .D(n3280), .CLK(clk), .Q(\keys[2][3] ), .QN(
        n399) );
  DFFX1_HVT \keys_reg[2][2]  ( .D(n3279), .CLK(clk), .Q(\keys[2][2] ), .QN(
        n400) );
  DFFX1_HVT \keys_reg[2][1]  ( .D(n3278), .CLK(clk), .Q(\keys[2][1] ), .QN(
        n401) );
  DFFX1_HVT \keys_reg[2][0]  ( .D(n3277), .CLK(clk), .Q(\keys[2][0] ), .QN(
        n402) );
  DFFX1_HVT \keys_reg[3][127]  ( .D(n3276), .CLK(clk), .Q(\keys[3][127] ), 
        .QN(n403) );
  DFFX1_HVT \keys_reg[3][126]  ( .D(n3275), .CLK(clk), .Q(\keys[3][126] ), 
        .QN(n404) );
  DFFX1_HVT \keys_reg[3][125]  ( .D(n3274), .CLK(clk), .Q(\keys[3][125] ), 
        .QN(n405) );
  DFFX1_HVT \keys_reg[3][124]  ( .D(n3273), .CLK(clk), .Q(\keys[3][124] ), 
        .QN(n406) );
  DFFX1_HVT \keys_reg[3][123]  ( .D(n3272), .CLK(clk), .Q(\keys[3][123] ), 
        .QN(n407) );
  DFFX1_HVT \keys_reg[3][122]  ( .D(n3271), .CLK(clk), .Q(\keys[3][122] ), 
        .QN(n408) );
  DFFX1_HVT \keys_reg[3][121]  ( .D(n3270), .CLK(clk), .Q(\keys[3][121] ), 
        .QN(n409) );
  DFFX1_HVT \keys_reg[3][120]  ( .D(n3269), .CLK(clk), .Q(\keys[3][120] ), 
        .QN(n410) );
  DFFX1_HVT \keys_reg[3][119]  ( .D(n3268), .CLK(clk), .Q(\keys[3][119] ), 
        .QN(n411) );
  DFFX1_HVT \keys_reg[3][118]  ( .D(n3267), .CLK(clk), .Q(\keys[3][118] ), 
        .QN(n412) );
  DFFX1_HVT \keys_reg[3][117]  ( .D(n3266), .CLK(clk), .Q(\keys[3][117] ), 
        .QN(n413) );
  DFFX1_HVT \keys_reg[3][116]  ( .D(n3265), .CLK(clk), .Q(\keys[3][116] ), 
        .QN(n414) );
  DFFX1_HVT \keys_reg[3][115]  ( .D(n3264), .CLK(clk), .Q(\keys[3][115] ), 
        .QN(n415) );
  DFFX1_HVT \keys_reg[3][114]  ( .D(n3263), .CLK(clk), .Q(\keys[3][114] ), 
        .QN(n416) );
  DFFX1_HVT \keys_reg[3][113]  ( .D(n3262), .CLK(clk), .Q(\keys[3][113] ), 
        .QN(n417) );
  DFFX1_HVT \keys_reg[3][112]  ( .D(n3261), .CLK(clk), .Q(\keys[3][112] ), 
        .QN(n418) );
  DFFX1_HVT \keys_reg[3][111]  ( .D(n3260), .CLK(clk), .Q(\keys[3][111] ), 
        .QN(n419) );
  DFFX1_HVT \keys_reg[3][110]  ( .D(n3259), .CLK(clk), .Q(\keys[3][110] ), 
        .QN(n420) );
  DFFX1_HVT \keys_reg[3][109]  ( .D(n3258), .CLK(clk), .Q(\keys[3][109] ), 
        .QN(n421) );
  DFFX1_HVT \keys_reg[3][108]  ( .D(n3257), .CLK(clk), .Q(\keys[3][108] ), 
        .QN(n422) );
  DFFX1_HVT \keys_reg[3][107]  ( .D(n3256), .CLK(clk), .Q(\keys[3][107] ), 
        .QN(n423) );
  DFFX1_HVT \keys_reg[3][106]  ( .D(n3255), .CLK(clk), .Q(\keys[3][106] ), 
        .QN(n424) );
  DFFX1_HVT \keys_reg[3][105]  ( .D(n3254), .CLK(clk), .Q(\keys[3][105] ), 
        .QN(n425) );
  DFFX1_HVT \keys_reg[3][104]  ( .D(n3253), .CLK(clk), .Q(\keys[3][104] ), 
        .QN(n426) );
  DFFX1_HVT \keys_reg[3][103]  ( .D(n3252), .CLK(clk), .Q(\keys[3][103] ), 
        .QN(n427) );
  DFFX1_HVT \keys_reg[3][102]  ( .D(n3251), .CLK(clk), .Q(\keys[3][102] ), 
        .QN(n428) );
  DFFX1_HVT \keys_reg[3][101]  ( .D(n3250), .CLK(clk), .Q(\keys[3][101] ), 
        .QN(n429) );
  DFFX1_HVT \keys_reg[3][100]  ( .D(n3249), .CLK(clk), .Q(\keys[3][100] ), 
        .QN(n430) );
  DFFX1_HVT \keys_reg[3][99]  ( .D(n3248), .CLK(clk), .Q(\keys[3][99] ), .QN(
        n431) );
  DFFX1_HVT \keys_reg[3][98]  ( .D(n3247), .CLK(clk), .Q(\keys[3][98] ), .QN(
        n432) );
  DFFX1_HVT \keys_reg[3][97]  ( .D(n3246), .CLK(clk), .Q(\keys[3][97] ), .QN(
        n433) );
  DFFX1_HVT \keys_reg[3][96]  ( .D(n3245), .CLK(clk), .Q(\keys[3][96] ), .QN(
        n434) );
  DFFX1_HVT \keys_reg[3][95]  ( .D(n3244), .CLK(clk), .Q(\keys[3][95] ), .QN(
        n435) );
  DFFX1_HVT \keys_reg[3][94]  ( .D(n3243), .CLK(clk), .Q(\keys[3][94] ), .QN(
        n436) );
  DFFX1_HVT \keys_reg[3][93]  ( .D(n3242), .CLK(clk), .Q(\keys[3][93] ), .QN(
        n437) );
  DFFX1_HVT \keys_reg[3][92]  ( .D(n3241), .CLK(clk), .Q(\keys[3][92] ), .QN(
        n438) );
  DFFX1_HVT \keys_reg[3][91]  ( .D(n3240), .CLK(clk), .QN(n439) );
  DFFX1_HVT \keys_reg[3][90]  ( .D(n3239), .CLK(clk), .QN(n440) );
  DFFX1_HVT \keys_reg[3][89]  ( .D(n3238), .CLK(clk), .Q(\keys[3][89] ), .QN(
        n441) );
  DFFX1_HVT \keys_reg[3][88]  ( .D(n3237), .CLK(clk), .Q(\keys[3][88] ), .QN(
        n442) );
  DFFX1_HVT \keys_reg[3][87]  ( .D(n3236), .CLK(clk), .Q(\keys[3][87] ), .QN(
        n443) );
  DFFX1_HVT \keys_reg[3][86]  ( .D(n3235), .CLK(clk), .Q(\keys[3][86] ), .QN(
        n444) );
  DFFX1_HVT \keys_reg[3][85]  ( .D(n3234), .CLK(clk), .Q(\keys[3][85] ), .QN(
        n445) );
  DFFX1_HVT \keys_reg[3][84]  ( .D(n3233), .CLK(clk), .Q(\keys[3][84] ), .QN(
        n446) );
  DFFX1_HVT \keys_reg[3][83]  ( .D(n3232), .CLK(clk), .Q(\keys[3][83] ), .QN(
        n447) );
  DFFX1_HVT \keys_reg[3][82]  ( .D(n3231), .CLK(clk), .Q(\keys[3][82] ), .QN(
        n448) );
  DFFX1_HVT \keys_reg[3][81]  ( .D(n3230), .CLK(clk), .Q(\keys[3][81] ), .QN(
        n449) );
  DFFX1_HVT \keys_reg[3][80]  ( .D(n3229), .CLK(clk), .Q(\keys[3][80] ), .QN(
        n450) );
  DFFX1_HVT \keys_reg[3][79]  ( .D(n3228), .CLK(clk), .Q(\keys[3][79] ), .QN(
        n451) );
  DFFX1_HVT \keys_reg[3][78]  ( .D(n3227), .CLK(clk), .Q(\keys[3][78] ), .QN(
        n452) );
  DFFX1_HVT \keys_reg[3][77]  ( .D(n3226), .CLK(clk), .Q(\keys[3][77] ), .QN(
        n453) );
  DFFX1_HVT \keys_reg[3][76]  ( .D(n3225), .CLK(clk), .Q(\keys[3][76] ), .QN(
        n454) );
  DFFX1_HVT \keys_reg[3][75]  ( .D(n3224), .CLK(clk), .Q(\keys[3][75] ), .QN(
        n455) );
  DFFX1_HVT \keys_reg[3][74]  ( .D(n3223), .CLK(clk), .Q(\keys[3][74] ), .QN(
        n456) );
  DFFX1_HVT \keys_reg[3][73]  ( .D(n3222), .CLK(clk), .Q(\keys[3][73] ), .QN(
        n457) );
  DFFX1_HVT \keys_reg[3][72]  ( .D(n3221), .CLK(clk), .Q(\keys[3][72] ), .QN(
        n458) );
  DFFX1_HVT \keys_reg[3][71]  ( .D(n3220), .CLK(clk), .Q(\keys[3][71] ), .QN(
        n459) );
  DFFX1_HVT \keys_reg[3][70]  ( .D(n3219), .CLK(clk), .Q(\keys[3][70] ), .QN(
        n460) );
  DFFX1_HVT \keys_reg[3][69]  ( .D(n3218), .CLK(clk), .Q(\keys[3][69] ), .QN(
        n461) );
  DFFX1_HVT \keys_reg[3][68]  ( .D(n3217), .CLK(clk), .Q(\keys[3][68] ), .QN(
        n462) );
  DFFX1_HVT \keys_reg[3][67]  ( .D(n3216), .CLK(clk), .Q(\keys[3][67] ), .QN(
        n463) );
  DFFX1_HVT \keys_reg[3][66]  ( .D(n3215), .CLK(clk), .Q(\keys[3][66] ), .QN(
        n464) );
  DFFX1_HVT \keys_reg[3][65]  ( .D(n3214), .CLK(clk), .Q(\keys[3][65] ), .QN(
        n465) );
  DFFX1_HVT \keys_reg[3][64]  ( .D(n3213), .CLK(clk), .Q(\keys[3][64] ), .QN(
        n466) );
  DFFX1_HVT \keys_reg[3][63]  ( .D(n3212), .CLK(clk), .Q(\keys[3][63] ), .QN(
        n467) );
  DFFX1_HVT \keys_reg[3][62]  ( .D(n3211), .CLK(clk), .Q(\keys[3][62] ), .QN(
        n468) );
  DFFX1_HVT \keys_reg[3][61]  ( .D(n3210), .CLK(clk), .Q(\keys[3][61] ), .QN(
        n469) );
  DFFX1_HVT \keys_reg[3][60]  ( .D(n3209), .CLK(clk), .Q(\keys[3][60] ), .QN(
        n470) );
  DFFX1_HVT \keys_reg[3][59]  ( .D(n3208), .CLK(clk), .Q(\keys[3][59] ), .QN(
        n471) );
  DFFX1_HVT \keys_reg[3][58]  ( .D(n3207), .CLK(clk), .Q(\keys[3][58] ), .QN(
        n472) );
  DFFX1_HVT \keys_reg[3][57]  ( .D(n3206), .CLK(clk), .Q(\keys[3][57] ), .QN(
        n473) );
  DFFX1_HVT \keys_reg[3][56]  ( .D(n3205), .CLK(clk), .Q(\keys[3][56] ), .QN(
        n474) );
  DFFX1_HVT \keys_reg[3][55]  ( .D(n3204), .CLK(clk), .Q(\keys[3][55] ), .QN(
        n475) );
  DFFX1_HVT \keys_reg[3][54]  ( .D(n3203), .CLK(clk), .Q(\keys[3][54] ), .QN(
        n476) );
  DFFX1_HVT \keys_reg[3][53]  ( .D(n3202), .CLK(clk), .Q(\keys[3][53] ), .QN(
        n477) );
  DFFX1_HVT \keys_reg[3][52]  ( .D(n3201), .CLK(clk), .Q(\keys[3][52] ), .QN(
        n478) );
  DFFX1_HVT \keys_reg[3][51]  ( .D(n3200), .CLK(clk), .Q(\keys[3][51] ), .QN(
        n479) );
  DFFX1_HVT \keys_reg[3][50]  ( .D(n3199), .CLK(clk), .Q(\keys[3][50] ), .QN(
        n480) );
  DFFX1_HVT \keys_reg[3][49]  ( .D(n3198), .CLK(clk), .Q(\keys[3][49] ), .QN(
        n481) );
  DFFX1_HVT \keys_reg[3][48]  ( .D(n3197), .CLK(clk), .Q(\keys[3][48] ), .QN(
        n482) );
  DFFX1_HVT \keys_reg[3][47]  ( .D(n3196), .CLK(clk), .Q(\keys[3][47] ), .QN(
        n483) );
  DFFX1_HVT \keys_reg[3][46]  ( .D(n3195), .CLK(clk), .Q(\keys[3][46] ), .QN(
        n484) );
  DFFX1_HVT \keys_reg[3][45]  ( .D(n3194), .CLK(clk), .Q(\keys[3][45] ), .QN(
        n485) );
  DFFX1_HVT \keys_reg[3][44]  ( .D(n3193), .CLK(clk), .Q(\keys[3][44] ), .QN(
        n486) );
  DFFX1_HVT \keys_reg[3][43]  ( .D(n3192), .CLK(clk), .Q(\keys[3][43] ), .QN(
        n487) );
  DFFX1_HVT \keys_reg[3][42]  ( .D(n3191), .CLK(clk), .Q(\keys[3][42] ), .QN(
        n488) );
  DFFX1_HVT \keys_reg[3][41]  ( .D(n3190), .CLK(clk), .Q(\keys[3][41] ), .QN(
        n489) );
  DFFX1_HVT \keys_reg[3][40]  ( .D(n3189), .CLK(clk), .Q(\keys[3][40] ), .QN(
        n490) );
  DFFX1_HVT \keys_reg[3][39]  ( .D(n3188), .CLK(clk), .Q(\keys[3][39] ), .QN(
        n491) );
  DFFX1_HVT \keys_reg[3][38]  ( .D(n3187), .CLK(clk), .Q(\keys[3][38] ), .QN(
        n492) );
  DFFX1_HVT \keys_reg[3][37]  ( .D(n3186), .CLK(clk), .Q(\keys[3][37] ), .QN(
        n493) );
  DFFX1_HVT \keys_reg[3][36]  ( .D(n3185), .CLK(clk), .Q(\keys[3][36] ), .QN(
        n494) );
  DFFX1_HVT \keys_reg[3][35]  ( .D(n3184), .CLK(clk), .Q(\keys[3][35] ), .QN(
        n495) );
  DFFX1_HVT \keys_reg[3][34]  ( .D(n3183), .CLK(clk), .Q(\keys[3][34] ), .QN(
        n496) );
  DFFX1_HVT \keys_reg[3][33]  ( .D(n3182), .CLK(clk), .Q(\keys[3][33] ), .QN(
        n497) );
  DFFX1_HVT \keys_reg[3][32]  ( .D(n3181), .CLK(clk), .Q(\keys[3][32] ), .QN(
        n498) );
  DFFX1_HVT \keys_reg[3][31]  ( .D(n3180), .CLK(clk), .Q(\keys[3][31] ), .QN(
        n499) );
  DFFX1_HVT \keys_reg[3][30]  ( .D(n3179), .CLK(clk), .Q(\keys[3][30] ), .QN(
        n500) );
  DFFX1_HVT \keys_reg[3][29]  ( .D(n3178), .CLK(clk), .Q(\keys[3][29] ), .QN(
        n501) );
  DFFX1_HVT \keys_reg[3][28]  ( .D(n3177), .CLK(clk), .Q(\keys[3][28] ), .QN(
        n502) );
  DFFX1_HVT \keys_reg[3][27]  ( .D(n3176), .CLK(clk), .Q(\keys[3][27] ), .QN(
        n503) );
  DFFX1_HVT \keys_reg[3][26]  ( .D(n3175), .CLK(clk), .Q(\keys[3][26] ), .QN(
        n504) );
  DFFX1_HVT \keys_reg[3][25]  ( .D(n3174), .CLK(clk), .Q(\keys[3][25] ), .QN(
        n505) );
  DFFX1_HVT \keys_reg[3][24]  ( .D(n3173), .CLK(clk), .Q(\keys[3][24] ), .QN(
        n506) );
  DFFX1_HVT \keys_reg[3][23]  ( .D(n3172), .CLK(clk), .Q(\keys[3][23] ), .QN(
        n507) );
  DFFX1_HVT \keys_reg[3][22]  ( .D(n3171), .CLK(clk), .Q(\keys[3][22] ), .QN(
        n508) );
  DFFX1_HVT \keys_reg[3][21]  ( .D(n3170), .CLK(clk), .Q(\keys[3][21] ), .QN(
        n509) );
  DFFX1_HVT \keys_reg[3][20]  ( .D(n3169), .CLK(clk), .Q(\keys[3][20] ), .QN(
        n510) );
  DFFX1_HVT \keys_reg[3][19]  ( .D(n3168), .CLK(clk), .Q(\keys[3][19] ), .QN(
        n511) );
  DFFX1_HVT \keys_reg[3][18]  ( .D(n3167), .CLK(clk), .Q(\keys[3][18] ), .QN(
        n512) );
  DFFX1_HVT \keys_reg[3][17]  ( .D(n3166), .CLK(clk), .Q(\keys[3][17] ), .QN(
        n513) );
  DFFX1_HVT \keys_reg[3][16]  ( .D(n3165), .CLK(clk), .Q(\keys[3][16] ), .QN(
        n514) );
  DFFX1_HVT \keys_reg[3][15]  ( .D(n3164), .CLK(clk), .Q(\keys[3][15] ), .QN(
        n515) );
  DFFX1_HVT \keys_reg[3][14]  ( .D(n3163), .CLK(clk), .Q(\keys[3][14] ), .QN(
        n516) );
  DFFX1_HVT \keys_reg[3][13]  ( .D(n3162), .CLK(clk), .Q(\keys[3][13] ), .QN(
        n517) );
  DFFX1_HVT \keys_reg[3][12]  ( .D(n3161), .CLK(clk), .Q(\keys[3][12] ), .QN(
        n518) );
  DFFX1_HVT \keys_reg[3][11]  ( .D(n3160), .CLK(clk), .Q(\keys[3][11] ), .QN(
        n519) );
  DFFX1_HVT \keys_reg[3][10]  ( .D(n3159), .CLK(clk), .Q(\keys[3][10] ), .QN(
        n520) );
  DFFX1_HVT \keys_reg[3][9]  ( .D(n3158), .CLK(clk), .Q(\keys[3][9] ), .QN(
        n521) );
  DFFX1_HVT \keys_reg[3][8]  ( .D(n3157), .CLK(clk), .Q(\keys[3][8] ), .QN(
        n522) );
  DFFX1_HVT \keys_reg[3][7]  ( .D(n3156), .CLK(clk), .Q(\keys[3][7] ), .QN(
        n523) );
  DFFX1_HVT \keys_reg[3][6]  ( .D(n3155), .CLK(clk), .Q(\keys[3][6] ), .QN(
        n524) );
  DFFX1_HVT \keys_reg[3][5]  ( .D(n3154), .CLK(clk), .Q(\keys[3][5] ), .QN(
        n525) );
  DFFX1_HVT \keys_reg[3][4]  ( .D(n3153), .CLK(clk), .Q(\keys[3][4] ), .QN(
        n526) );
  DFFX1_HVT \keys_reg[3][3]  ( .D(n3152), .CLK(clk), .Q(\keys[3][3] ), .QN(
        n527) );
  DFFX1_HVT \keys_reg[3][2]  ( .D(n3151), .CLK(clk), .Q(\keys[3][2] ), .QN(
        n528) );
  DFFX1_HVT \keys_reg[3][1]  ( .D(n3150), .CLK(clk), .Q(\keys[3][1] ), .QN(
        n529) );
  DFFX1_HVT \keys_reg[3][0]  ( .D(n3149), .CLK(clk), .Q(\keys[3][0] ), .QN(
        n530) );
  DFFX1_HVT \keys_reg[4][127]  ( .D(n3148), .CLK(clk), .Q(\keys[4][127] ), 
        .QN(n531) );
  DFFX1_HVT \keys_reg[4][126]  ( .D(n3147), .CLK(clk), .Q(\keys[4][126] ), 
        .QN(n532) );
  DFFX1_HVT \keys_reg[4][125]  ( .D(n3146), .CLK(clk), .Q(\keys[4][125] ), 
        .QN(n533) );
  DFFX1_HVT \keys_reg[4][124]  ( .D(n3145), .CLK(clk), .Q(\keys[4][124] ), 
        .QN(n534) );
  DFFX1_HVT \keys_reg[4][123]  ( .D(n3144), .CLK(clk), .Q(\keys[4][123] ), 
        .QN(n535) );
  DFFX1_HVT \keys_reg[4][122]  ( .D(n3143), .CLK(clk), .Q(\keys[4][122] ), 
        .QN(n536) );
  DFFX1_HVT \keys_reg[4][121]  ( .D(n3142), .CLK(clk), .Q(\keys[4][121] ), 
        .QN(n537) );
  DFFX1_HVT \keys_reg[4][120]  ( .D(n3141), .CLK(clk), .Q(\keys[4][120] ), 
        .QN(n538) );
  DFFX1_HVT \keys_reg[4][119]  ( .D(n3140), .CLK(clk), .Q(\keys[4][119] ), 
        .QN(n539) );
  DFFX1_HVT \keys_reg[4][118]  ( .D(n3139), .CLK(clk), .Q(\keys[4][118] ), 
        .QN(n540) );
  DFFX1_HVT \keys_reg[4][117]  ( .D(n3138), .CLK(clk), .Q(\keys[4][117] ), 
        .QN(n541) );
  DFFX1_HVT \keys_reg[4][116]  ( .D(n3137), .CLK(clk), .Q(\keys[4][116] ), 
        .QN(n542) );
  DFFX1_HVT \keys_reg[4][115]  ( .D(n3136), .CLK(clk), .Q(\keys[4][115] ), 
        .QN(n543) );
  DFFX1_HVT \keys_reg[4][114]  ( .D(n3135), .CLK(clk), .Q(\keys[4][114] ), 
        .QN(n544) );
  DFFX1_HVT \keys_reg[4][113]  ( .D(n3134), .CLK(clk), .Q(\keys[4][113] ), 
        .QN(n545) );
  DFFX1_HVT \keys_reg[4][112]  ( .D(n3133), .CLK(clk), .Q(\keys[4][112] ), 
        .QN(n546) );
  DFFX1_HVT \keys_reg[4][111]  ( .D(n3132), .CLK(clk), .Q(\keys[4][111] ), 
        .QN(n547) );
  DFFX1_HVT \keys_reg[4][110]  ( .D(n3131), .CLK(clk), .Q(\keys[4][110] ), 
        .QN(n548) );
  DFFX1_HVT \keys_reg[4][109]  ( .D(n3130), .CLK(clk), .Q(\keys[4][109] ), 
        .QN(n549) );
  DFFX1_HVT \keys_reg[4][108]  ( .D(n3129), .CLK(clk), .Q(\keys[4][108] ), 
        .QN(n550) );
  DFFX1_HVT \keys_reg[4][107]  ( .D(n3128), .CLK(clk), .Q(\keys[4][107] ), 
        .QN(n551) );
  DFFX1_HVT \keys_reg[4][106]  ( .D(n3127), .CLK(clk), .Q(\keys[4][106] ), 
        .QN(n552) );
  DFFX1_HVT \keys_reg[4][105]  ( .D(n3126), .CLK(clk), .Q(\keys[4][105] ), 
        .QN(n553) );
  DFFX1_HVT \keys_reg[4][104]  ( .D(n3125), .CLK(clk), .Q(\keys[4][104] ), 
        .QN(n554) );
  DFFX1_HVT \keys_reg[4][103]  ( .D(n3124), .CLK(clk), .Q(\keys[4][103] ), 
        .QN(n555) );
  DFFX1_HVT \keys_reg[4][102]  ( .D(n3123), .CLK(clk), .Q(\keys[4][102] ), 
        .QN(n556) );
  DFFX1_HVT \keys_reg[4][101]  ( .D(n3122), .CLK(clk), .Q(\keys[4][101] ), 
        .QN(n557) );
  DFFX1_HVT \keys_reg[4][100]  ( .D(n3121), .CLK(clk), .Q(\keys[4][100] ), 
        .QN(n558) );
  DFFX1_HVT \keys_reg[4][99]  ( .D(n3120), .CLK(clk), .Q(\keys[4][99] ), .QN(
        n559) );
  DFFX1_HVT \keys_reg[4][98]  ( .D(n3119), .CLK(clk), .Q(\keys[4][98] ), .QN(
        n560) );
  DFFX1_HVT \keys_reg[4][97]  ( .D(n3118), .CLK(clk), .Q(\keys[4][97] ), .QN(
        n561) );
  DFFX1_HVT \keys_reg[4][96]  ( .D(n3117), .CLK(clk), .Q(\keys[4][96] ), .QN(
        n562) );
  DFFX1_HVT \keys_reg[4][95]  ( .D(n3116), .CLK(clk), .Q(\keys[4][95] ), .QN(
        n563) );
  DFFX1_HVT \keys_reg[4][94]  ( .D(n3115), .CLK(clk), .Q(\keys[4][94] ), .QN(
        n564) );
  DFFX1_HVT \keys_reg[4][93]  ( .D(n3114), .CLK(clk), .Q(\keys[4][93] ), .QN(
        n565) );
  DFFX1_HVT \keys_reg[4][92]  ( .D(n3113), .CLK(clk), .Q(\keys[4][92] ), .QN(
        n566) );
  DFFX1_HVT \keys_reg[4][91]  ( .D(n3112), .CLK(clk), .Q(\keys[4][91] ), .QN(
        n567) );
  DFFX1_HVT \keys_reg[4][90]  ( .D(n3111), .CLK(clk), .Q(\keys[4][90] ), .QN(
        n568) );
  DFFX1_HVT \keys_reg[4][89]  ( .D(n3110), .CLK(clk), .Q(\keys[4][89] ), .QN(
        n569) );
  DFFX1_HVT \keys_reg[4][88]  ( .D(n3109), .CLK(clk), .Q(\keys[4][88] ), .QN(
        n570) );
  DFFX1_HVT \keys_reg[4][87]  ( .D(n3108), .CLK(clk), .Q(\keys[4][87] ), .QN(
        n571) );
  DFFX1_HVT \keys_reg[4][86]  ( .D(n3107), .CLK(clk), .Q(\keys[4][86] ), .QN(
        n572) );
  DFFX1_HVT \keys_reg[4][85]  ( .D(n3106), .CLK(clk), .Q(\keys[4][85] ), .QN(
        n573) );
  DFFX1_HVT \keys_reg[4][84]  ( .D(n3105), .CLK(clk), .Q(\keys[4][84] ), .QN(
        n574) );
  DFFX1_HVT \keys_reg[4][83]  ( .D(n3104), .CLK(clk), .Q(\keys[4][83] ), .QN(
        n575) );
  DFFX1_HVT \keys_reg[4][82]  ( .D(n3103), .CLK(clk), .Q(\keys[4][82] ), .QN(
        n576) );
  DFFX1_HVT \keys_reg[4][81]  ( .D(n3102), .CLK(clk), .Q(\keys[4][81] ), .QN(
        n577) );
  DFFX1_HVT \keys_reg[4][80]  ( .D(n3101), .CLK(clk), .Q(\keys[4][80] ), .QN(
        n578) );
  DFFX1_HVT \keys_reg[4][79]  ( .D(n3100), .CLK(clk), .Q(\keys[4][79] ), .QN(
        n579) );
  DFFX1_HVT \keys_reg[4][78]  ( .D(n3099), .CLK(clk), .Q(\keys[4][78] ), .QN(
        n580) );
  DFFX1_HVT \keys_reg[4][77]  ( .D(n3098), .CLK(clk), .Q(\keys[4][77] ), .QN(
        n581) );
  DFFX1_HVT \keys_reg[4][76]  ( .D(n3097), .CLK(clk), .Q(\keys[4][76] ), .QN(
        n582) );
  DFFX1_HVT \keys_reg[4][75]  ( .D(n3096), .CLK(clk), .QN(n583) );
  DFFX1_HVT \keys_reg[4][74]  ( .D(n3095), .CLK(clk), .QN(n584) );
  DFFX1_HVT \keys_reg[4][73]  ( .D(n3094), .CLK(clk), .Q(\keys[4][73] ), .QN(
        n585) );
  DFFX1_HVT \keys_reg[4][72]  ( .D(n3093), .CLK(clk), .Q(\keys[4][72] ), .QN(
        n586) );
  DFFX1_HVT \keys_reg[4][71]  ( .D(n3092), .CLK(clk), .Q(\keys[4][71] ), .QN(
        n587) );
  DFFX1_HVT \keys_reg[4][70]  ( .D(n3091), .CLK(clk), .Q(\keys[4][70] ), .QN(
        n588) );
  DFFX1_HVT \keys_reg[4][69]  ( .D(n3090), .CLK(clk), .Q(\keys[4][69] ), .QN(
        n589) );
  DFFX1_HVT \keys_reg[4][68]  ( .D(n3089), .CLK(clk), .Q(\keys[4][68] ), .QN(
        n590) );
  DFFX1_HVT \keys_reg[4][67]  ( .D(n3088), .CLK(clk), .Q(\keys[4][67] ), .QN(
        n591) );
  DFFX1_HVT \keys_reg[4][66]  ( .D(n3087), .CLK(clk), .Q(\keys[4][66] ), .QN(
        n592) );
  DFFX1_HVT \keys_reg[4][65]  ( .D(n3086), .CLK(clk), .Q(\keys[4][65] ), .QN(
        n593) );
  DFFX1_HVT \keys_reg[4][64]  ( .D(n3085), .CLK(clk), .Q(\keys[4][64] ), .QN(
        n594) );
  DFFX1_HVT \keys_reg[4][63]  ( .D(n3084), .CLK(clk), .Q(\keys[4][63] ), .QN(
        n595) );
  DFFX1_HVT \keys_reg[4][62]  ( .D(n3083), .CLK(clk), .Q(\keys[4][62] ), .QN(
        n596) );
  DFFX1_HVT \keys_reg[4][61]  ( .D(n3082), .CLK(clk), .Q(\keys[4][61] ), .QN(
        n597) );
  DFFX1_HVT \keys_reg[4][60]  ( .D(n3081), .CLK(clk), .Q(\keys[4][60] ), .QN(
        n598) );
  DFFX1_HVT \keys_reg[4][59]  ( .D(n3080), .CLK(clk), .Q(\keys[4][59] ), .QN(
        n599) );
  DFFX1_HVT \keys_reg[4][58]  ( .D(n3079), .CLK(clk), .Q(\keys[4][58] ), .QN(
        n600) );
  DFFX1_HVT \keys_reg[4][57]  ( .D(n3078), .CLK(clk), .Q(\keys[4][57] ), .QN(
        n601) );
  DFFX1_HVT \keys_reg[4][56]  ( .D(n3077), .CLK(clk), .Q(\keys[4][56] ), .QN(
        n602) );
  DFFX1_HVT \keys_reg[4][55]  ( .D(n3076), .CLK(clk), .Q(\keys[4][55] ), .QN(
        n603) );
  DFFX1_HVT \keys_reg[4][54]  ( .D(n3075), .CLK(clk), .Q(\keys[4][54] ), .QN(
        n604) );
  DFFX1_HVT \keys_reg[4][53]  ( .D(n3074), .CLK(clk), .Q(\keys[4][53] ), .QN(
        n605) );
  DFFX1_HVT \keys_reg[4][52]  ( .D(n3073), .CLK(clk), .Q(\keys[4][52] ), .QN(
        n606) );
  DFFX1_HVT \keys_reg[4][51]  ( .D(n3072), .CLK(clk), .Q(\keys[4][51] ), .QN(
        n607) );
  DFFX1_HVT \keys_reg[4][50]  ( .D(n3071), .CLK(clk), .Q(\keys[4][50] ), .QN(
        n608) );
  DFFX1_HVT \keys_reg[4][49]  ( .D(n3070), .CLK(clk), .Q(\keys[4][49] ), .QN(
        n609) );
  DFFX1_HVT \keys_reg[4][48]  ( .D(n3069), .CLK(clk), .Q(\keys[4][48] ), .QN(
        n610) );
  DFFX1_HVT \keys_reg[4][47]  ( .D(n3068), .CLK(clk), .Q(\keys[4][47] ), .QN(
        n611) );
  DFFX1_HVT \keys_reg[4][46]  ( .D(n3067), .CLK(clk), .Q(\keys[4][46] ), .QN(
        n612) );
  DFFX1_HVT \keys_reg[4][45]  ( .D(n3066), .CLK(clk), .Q(\keys[4][45] ), .QN(
        n613) );
  DFFX1_HVT \keys_reg[4][44]  ( .D(n3065), .CLK(clk), .Q(n3877), .QN(n614) );
  DFFX1_HVT \keys_reg[4][43]  ( .D(n3064), .CLK(clk), .Q(\keys[4][43] ), .QN(
        n615) );
  DFFX1_HVT \keys_reg[4][42]  ( .D(n3063), .CLK(clk), .Q(\keys[4][42] ), .QN(
        n616) );
  DFFX1_HVT \keys_reg[4][41]  ( .D(n3062), .CLK(clk), .Q(\keys[4][41] ), .QN(
        n617) );
  DFFX1_HVT \keys_reg[4][40]  ( .D(n3061), .CLK(clk), .Q(\keys[4][40] ), .QN(
        n618) );
  DFFX1_HVT \keys_reg[4][39]  ( .D(n3060), .CLK(clk), .Q(\keys[4][39] ), .QN(
        n619) );
  DFFX1_HVT \keys_reg[4][38]  ( .D(n3059), .CLK(clk), .Q(\keys[4][38] ), .QN(
        n620) );
  DFFX1_HVT \keys_reg[4][37]  ( .D(n3058), .CLK(clk), .Q(\keys[4][37] ), .QN(
        n621) );
  DFFX1_HVT \keys_reg[4][36]  ( .D(n3057), .CLK(clk), .Q(\keys[4][36] ), .QN(
        n622) );
  DFFX1_HVT \keys_reg[4][35]  ( .D(n3056), .CLK(clk), .Q(\keys[4][35] ), .QN(
        n623) );
  DFFX1_HVT \keys_reg[4][34]  ( .D(n3055), .CLK(clk), .Q(\keys[4][34] ), .QN(
        n624) );
  DFFX1_HVT \keys_reg[4][33]  ( .D(n3054), .CLK(clk), .Q(\keys[4][33] ), .QN(
        n625) );
  DFFX1_HVT \keys_reg[4][32]  ( .D(n3053), .CLK(clk), .Q(\keys[4][32] ), .QN(
        n626) );
  DFFX1_HVT \keys_reg[4][31]  ( .D(n3052), .CLK(clk), .Q(\keys[4][31] ), .QN(
        n627) );
  DFFX1_HVT \keys_reg[4][30]  ( .D(n3051), .CLK(clk), .Q(\keys[4][30] ), .QN(
        n628) );
  DFFX1_HVT \keys_reg[4][29]  ( .D(n3050), .CLK(clk), .Q(\keys[4][29] ), .QN(
        n629) );
  DFFX1_HVT \keys_reg[4][28]  ( .D(n3049), .CLK(clk), .Q(\keys[4][28] ), .QN(
        n630) );
  DFFX1_HVT \keys_reg[4][27]  ( .D(n3048), .CLK(clk), .Q(\keys[4][27] ), .QN(
        n631) );
  DFFX1_HVT \keys_reg[4][26]  ( .D(n3047), .CLK(clk), .Q(\keys[4][26] ), .QN(
        n632) );
  DFFX1_HVT \keys_reg[4][25]  ( .D(n3046), .CLK(clk), .Q(\keys[4][25] ), .QN(
        n633) );
  DFFX1_HVT \keys_reg[4][24]  ( .D(n3045), .CLK(clk), .Q(\keys[4][24] ), .QN(
        n634) );
  DFFX1_HVT \keys_reg[4][23]  ( .D(n3044), .CLK(clk), .Q(\keys[4][23] ), .QN(
        n635) );
  DFFX1_HVT \keys_reg[4][22]  ( .D(n3043), .CLK(clk), .Q(\keys[4][22] ), .QN(
        n636) );
  DFFX1_HVT \keys_reg[4][21]  ( .D(n3042), .CLK(clk), .Q(\keys[4][21] ), .QN(
        n637) );
  DFFX1_HVT \keys_reg[4][20]  ( .D(n3041), .CLK(clk), .Q(\keys[4][20] ), .QN(
        n638) );
  DFFX1_HVT \keys_reg[4][19]  ( .D(n3040), .CLK(clk), .Q(\keys[4][19] ), .QN(
        n639) );
  DFFX1_HVT \keys_reg[4][18]  ( .D(n3039), .CLK(clk), .Q(\keys[4][18] ), .QN(
        n640) );
  DFFX1_HVT \keys_reg[4][17]  ( .D(n3038), .CLK(clk), .Q(\keys[4][17] ), .QN(
        n641) );
  DFFX1_HVT \keys_reg[4][16]  ( .D(n3037), .CLK(clk), .Q(\keys[4][16] ), .QN(
        n642) );
  DFFX1_HVT \keys_reg[4][15]  ( .D(n3036), .CLK(clk), .Q(\keys[4][15] ), .QN(
        n643) );
  DFFX1_HVT \keys_reg[4][14]  ( .D(n3035), .CLK(clk), .Q(\keys[4][14] ), .QN(
        n644) );
  DFFX1_HVT \keys_reg[4][13]  ( .D(n3034), .CLK(clk), .Q(\keys[4][13] ), .QN(
        n645) );
  DFFX1_HVT \keys_reg[4][12]  ( .D(n3033), .CLK(clk), .Q(\keys[4][12] ), .QN(
        n646) );
  DFFX1_HVT \keys_reg[4][11]  ( .D(n3032), .CLK(clk), .Q(\keys[4][11] ), .QN(
        n647) );
  DFFX1_HVT \keys_reg[4][10]  ( .D(n3031), .CLK(clk), .Q(\keys[4][10] ), .QN(
        n648) );
  DFFX1_HVT \keys_reg[4][9]  ( .D(n3030), .CLK(clk), .Q(\keys[4][9] ), .QN(
        n649) );
  DFFX1_HVT \keys_reg[4][8]  ( .D(n3029), .CLK(clk), .Q(\keys[4][8] ), .QN(
        n650) );
  DFFX1_HVT \keys_reg[4][7]  ( .D(n3028), .CLK(clk), .Q(\keys[4][7] ), .QN(
        n651) );
  DFFX1_HVT \keys_reg[4][6]  ( .D(n3027), .CLK(clk), .Q(\keys[4][6] ), .QN(
        n652) );
  DFFX1_HVT \keys_reg[4][5]  ( .D(n3026), .CLK(clk), .Q(\keys[4][5] ), .QN(
        n653) );
  DFFX1_HVT \keys_reg[4][4]  ( .D(n3025), .CLK(clk), .Q(\keys[4][4] ), .QN(
        n654) );
  DFFX1_HVT \keys_reg[4][3]  ( .D(n3024), .CLK(clk), .Q(\keys[4][3] ), .QN(
        n655) );
  DFFX1_HVT \keys_reg[4][2]  ( .D(n3023), .CLK(clk), .Q(\keys[4][2] ), .QN(
        n656) );
  DFFX1_HVT \keys_reg[4][1]  ( .D(n3022), .CLK(clk), .Q(\keys[4][1] ), .QN(
        n657) );
  DFFX1_HVT \keys_reg[4][0]  ( .D(n3021), .CLK(clk), .Q(\keys[4][0] ), .QN(
        n658) );
  DFFX1_HVT \keys_reg[5][127]  ( .D(n3020), .CLK(clk), .Q(\keys[5][127] ), 
        .QN(n659) );
  DFFX1_HVT \keys_reg[5][126]  ( .D(n3019), .CLK(clk), .Q(\keys[5][126] ), 
        .QN(n660) );
  DFFX1_HVT \keys_reg[5][125]  ( .D(n3018), .CLK(clk), .Q(\keys[5][125] ), 
        .QN(n661) );
  DFFX1_HVT \keys_reg[5][124]  ( .D(n3017), .CLK(clk), .Q(\keys[5][124] ), 
        .QN(n662) );
  DFFX1_HVT \keys_reg[5][123]  ( .D(n3016), .CLK(clk), .Q(\keys[5][123] ), 
        .QN(n663) );
  DFFX1_HVT \keys_reg[5][122]  ( .D(n3015), .CLK(clk), .Q(\keys[5][122] ), 
        .QN(n664) );
  DFFX1_HVT \keys_reg[5][121]  ( .D(n3014), .CLK(clk), .Q(\keys[5][121] ), 
        .QN(n665) );
  DFFX1_HVT \keys_reg[5][120]  ( .D(n3013), .CLK(clk), .Q(\keys[5][120] ), 
        .QN(n666) );
  DFFX1_HVT \keys_reg[5][119]  ( .D(n3012), .CLK(clk), .Q(\keys[5][119] ), 
        .QN(n667) );
  DFFX1_HVT \keys_reg[5][118]  ( .D(n3011), .CLK(clk), .Q(\keys[5][118] ), 
        .QN(n668) );
  DFFX1_HVT \keys_reg[5][117]  ( .D(n3010), .CLK(clk), .Q(\keys[5][117] ), 
        .QN(n669) );
  DFFX1_HVT \keys_reg[5][116]  ( .D(n3009), .CLK(clk), .Q(\keys[5][116] ), 
        .QN(n670) );
  DFFX1_HVT \keys_reg[5][115]  ( .D(n3008), .CLK(clk), .Q(\keys[5][115] ), 
        .QN(n671) );
  DFFX1_HVT \keys_reg[5][114]  ( .D(n3007), .CLK(clk), .Q(\keys[5][114] ), 
        .QN(n672) );
  DFFX1_HVT \keys_reg[5][113]  ( .D(n3006), .CLK(clk), .Q(\keys[5][113] ), 
        .QN(n673) );
  DFFX1_HVT \keys_reg[5][112]  ( .D(n3005), .CLK(clk), .Q(\keys[5][112] ), 
        .QN(n674) );
  DFFX1_HVT \keys_reg[5][111]  ( .D(n3004), .CLK(clk), .Q(\keys[5][111] ), 
        .QN(n675) );
  DFFX1_HVT \keys_reg[5][110]  ( .D(n3003), .CLK(clk), .Q(\keys[5][110] ), 
        .QN(n676) );
  DFFX1_HVT \keys_reg[5][109]  ( .D(n3002), .CLK(clk), .Q(\keys[5][109] ), 
        .QN(n677) );
  DFFX1_HVT \keys_reg[5][108]  ( .D(n3001), .CLK(clk), .Q(\keys[5][108] ), 
        .QN(n678) );
  DFFX1_HVT \keys_reg[5][107]  ( .D(n3000), .CLK(clk), .Q(\keys[5][107] ), 
        .QN(n679) );
  DFFX1_HVT \keys_reg[5][106]  ( .D(n2999), .CLK(clk), .Q(\keys[5][106] ), 
        .QN(n680) );
  DFFX1_HVT \keys_reg[5][105]  ( .D(n2998), .CLK(clk), .Q(\keys[5][105] ), 
        .QN(n681) );
  DFFX1_HVT \keys_reg[5][104]  ( .D(n2997), .CLK(clk), .Q(\keys[5][104] ), 
        .QN(n682) );
  DFFX1_HVT \keys_reg[5][103]  ( .D(n2996), .CLK(clk), .Q(\keys[5][103] ), 
        .QN(n683) );
  DFFX1_HVT \keys_reg[5][102]  ( .D(n2995), .CLK(clk), .Q(\keys[5][102] ), 
        .QN(n684) );
  DFFX1_HVT \keys_reg[5][101]  ( .D(n2994), .CLK(clk), .Q(\keys[5][101] ), 
        .QN(n685) );
  DFFX1_HVT \keys_reg[5][100]  ( .D(n2993), .CLK(clk), .Q(\keys[5][100] ), 
        .QN(n686) );
  DFFX1_HVT \keys_reg[5][99]  ( .D(n2992), .CLK(clk), .Q(\keys[5][99] ), .QN(
        n687) );
  DFFX1_HVT \keys_reg[5][98]  ( .D(n2991), .CLK(clk), .Q(\keys[5][98] ), .QN(
        n688) );
  DFFX1_HVT \keys_reg[5][97]  ( .D(n2990), .CLK(clk), .Q(\keys[5][97] ), .QN(
        n689) );
  DFFX1_HVT \keys_reg[5][96]  ( .D(n2989), .CLK(clk), .Q(\keys[5][96] ), .QN(
        n690) );
  DFFX1_HVT \keys_reg[5][95]  ( .D(n2988), .CLK(clk), .Q(\keys[5][95] ), .QN(
        n691) );
  DFFX1_HVT \keys_reg[5][94]  ( .D(n2987), .CLK(clk), .Q(\keys[5][94] ), .QN(
        n692) );
  DFFX1_HVT \keys_reg[5][93]  ( .D(n2986), .CLK(clk), .Q(\keys[5][93] ), .QN(
        n693) );
  DFFX1_HVT \keys_reg[5][92]  ( .D(n2985), .CLK(clk), .Q(\keys[5][92] ), .QN(
        n694) );
  DFFX1_HVT \keys_reg[5][91]  ( .D(n2984), .CLK(clk), .Q(\keys[5][91] ), .QN(
        n695) );
  DFFX1_HVT \keys_reg[5][90]  ( .D(n2983), .CLK(clk), .Q(\keys[5][90] ), .QN(
        n696) );
  DFFX1_HVT \keys_reg[5][89]  ( .D(n2982), .CLK(clk), .Q(\keys[5][89] ), .QN(
        n697) );
  DFFX1_HVT \keys_reg[5][88]  ( .D(n2981), .CLK(clk), .Q(\keys[5][88] ), .QN(
        n698) );
  DFFX1_HVT \keys_reg[5][87]  ( .D(n2980), .CLK(clk), .Q(\keys[5][87] ), .QN(
        n699) );
  DFFX1_HVT \keys_reg[5][86]  ( .D(n2979), .CLK(clk), .Q(\keys[5][86] ), .QN(
        n700) );
  DFFX1_HVT \keys_reg[5][85]  ( .D(n2978), .CLK(clk), .Q(\keys[5][85] ), .QN(
        n701) );
  DFFX1_HVT \keys_reg[5][84]  ( .D(n2977), .CLK(clk), .Q(\keys[5][84] ), .QN(
        n702) );
  DFFX1_HVT \keys_reg[5][83]  ( .D(n2976), .CLK(clk), .Q(\keys[5][83] ), .QN(
        n703) );
  DFFX1_HVT \keys_reg[5][82]  ( .D(n2975), .CLK(clk), .Q(\keys[5][82] ), .QN(
        n704) );
  DFFX1_HVT \keys_reg[5][81]  ( .D(n2974), .CLK(clk), .Q(\keys[5][81] ), .QN(
        n705) );
  DFFX1_HVT \keys_reg[5][80]  ( .D(n2973), .CLK(clk), .Q(\keys[5][80] ), .QN(
        n706) );
  DFFX1_HVT \keys_reg[5][79]  ( .D(n2972), .CLK(clk), .Q(\keys[5][79] ), .QN(
        n707) );
  DFFX1_HVT \keys_reg[5][78]  ( .D(n2971), .CLK(clk), .Q(\keys[5][78] ), .QN(
        n708) );
  DFFX1_HVT \keys_reg[5][77]  ( .D(n2970), .CLK(clk), .Q(\keys[5][77] ), .QN(
        n709) );
  DFFX1_HVT \keys_reg[5][76]  ( .D(n2969), .CLK(clk), .Q(\keys[5][76] ), .QN(
        n710) );
  DFFX1_HVT \keys_reg[5][75]  ( .D(n2968), .CLK(clk), .Q(\keys[5][75] ), .QN(
        n711) );
  DFFX1_HVT \keys_reg[5][74]  ( .D(n2967), .CLK(clk), .Q(\keys[5][74] ), .QN(
        n712) );
  DFFX1_HVT \keys_reg[5][73]  ( .D(n2966), .CLK(clk), .Q(\keys[5][73] ), .QN(
        n713) );
  DFFX1_HVT \keys_reg[5][72]  ( .D(n2965), .CLK(clk), .Q(\keys[5][72] ), .QN(
        n714) );
  DFFX1_HVT \keys_reg[5][71]  ( .D(n2964), .CLK(clk), .Q(\keys[5][71] ), .QN(
        n715) );
  DFFX1_HVT \keys_reg[5][70]  ( .D(n2963), .CLK(clk), .Q(\keys[5][70] ), .QN(
        n716) );
  DFFX1_HVT \keys_reg[5][69]  ( .D(n2962), .CLK(clk), .Q(\keys[5][69] ), .QN(
        n717) );
  DFFX1_HVT \keys_reg[5][68]  ( .D(n2961), .CLK(clk), .Q(\keys[5][68] ), .QN(
        n718) );
  DFFX1_HVT \keys_reg[5][67]  ( .D(n2960), .CLK(clk), .Q(\keys[5][67] ), .QN(
        n719) );
  DFFX1_HVT \keys_reg[5][66]  ( .D(n2959), .CLK(clk), .Q(\keys[5][66] ), .QN(
        n720) );
  DFFX1_HVT \keys_reg[5][65]  ( .D(n2958), .CLK(clk), .Q(\keys[5][65] ), .QN(
        n721) );
  DFFX1_HVT \keys_reg[5][64]  ( .D(n2957), .CLK(clk), .Q(\keys[5][64] ), .QN(
        n722) );
  DFFX1_HVT \keys_reg[5][63]  ( .D(n2956), .CLK(clk), .Q(\keys[5][63] ), .QN(
        n723) );
  DFFX1_HVT \keys_reg[5][62]  ( .D(n2955), .CLK(clk), .Q(\keys[5][62] ), .QN(
        n724) );
  DFFX1_HVT \keys_reg[5][61]  ( .D(n2954), .CLK(clk), .Q(\keys[5][61] ), .QN(
        n725) );
  DFFX1_HVT \keys_reg[5][60]  ( .D(n2953), .CLK(clk), .Q(\keys[5][60] ), .QN(
        n726) );
  DFFX1_HVT \keys_reg[5][59]  ( .D(n2952), .CLK(clk), .Q(\keys[5][59] ), .QN(
        n727) );
  DFFX1_HVT \keys_reg[5][58]  ( .D(n2951), .CLK(clk), .Q(\keys[5][58] ), .QN(
        n728) );
  DFFX1_HVT \keys_reg[5][57]  ( .D(n2950), .CLK(clk), .Q(\keys[5][57] ), .QN(
        n729) );
  DFFX1_HVT \keys_reg[5][56]  ( .D(n2949), .CLK(clk), .Q(\keys[5][56] ), .QN(
        n730) );
  DFFX1_HVT \keys_reg[5][55]  ( .D(n2948), .CLK(clk), .QN(n731) );
  DFFX1_HVT \keys_reg[5][54]  ( .D(n2947), .CLK(clk), .Q(\keys[5][54] ), .QN(
        n732) );
  DFFX1_HVT \keys_reg[5][53]  ( .D(n2946), .CLK(clk), .Q(\keys[5][53] ), .QN(
        n733) );
  DFFX1_HVT \keys_reg[5][52]  ( .D(n2945), .CLK(clk), .Q(\keys[5][52] ), .QN(
        n734) );
  DFFX1_HVT \keys_reg[5][51]  ( .D(n2944), .CLK(clk), .Q(\keys[5][51] ), .QN(
        n735) );
  DFFX1_HVT \keys_reg[5][50]  ( .D(n2943), .CLK(clk), .Q(\keys[5][50] ), .QN(
        n736) );
  DFFX1_HVT \keys_reg[5][49]  ( .D(n2942), .CLK(clk), .Q(\keys[5][49] ), .QN(
        n737) );
  DFFX1_HVT \keys_reg[5][48]  ( .D(n2941), .CLK(clk), .Q(\keys[5][48] ), .QN(
        n738) );
  DFFX1_HVT \keys_reg[5][47]  ( .D(n2940), .CLK(clk), .Q(\keys[5][47] ), .QN(
        n739) );
  DFFX1_HVT \keys_reg[5][46]  ( .D(n2939), .CLK(clk), .Q(\keys[5][46] ), .QN(
        n740) );
  DFFX1_HVT \keys_reg[5][45]  ( .D(n2938), .CLK(clk), .Q(\keys[5][45] ), .QN(
        n741) );
  DFFX1_HVT \keys_reg[5][44]  ( .D(n2937), .CLK(clk), .Q(\keys[5][44] ), .QN(
        n742) );
  DFFX1_HVT \keys_reg[5][43]  ( .D(n2936), .CLK(clk), .Q(\keys[5][43] ), .QN(
        n743) );
  DFFX1_HVT \keys_reg[5][42]  ( .D(n2935), .CLK(clk), .Q(\keys[5][42] ), .QN(
        n744) );
  DFFX1_HVT \keys_reg[5][41]  ( .D(n2934), .CLK(clk), .Q(\keys[5][41] ), .QN(
        n745) );
  DFFX1_HVT \keys_reg[5][40]  ( .D(n2933), .CLK(clk), .Q(\keys[5][40] ), .QN(
        n746) );
  DFFX1_HVT \keys_reg[5][39]  ( .D(n2932), .CLK(clk), .Q(\keys[5][39] ), .QN(
        n747) );
  DFFX1_HVT \keys_reg[5][38]  ( .D(n2931), .CLK(clk), .Q(\keys[5][38] ), .QN(
        n748) );
  DFFX1_HVT \keys_reg[5][37]  ( .D(n2930), .CLK(clk), .Q(\keys[5][37] ), .QN(
        n749) );
  DFFX1_HVT \keys_reg[5][36]  ( .D(n2929), .CLK(clk), .Q(\keys[5][36] ), .QN(
        n750) );
  DFFX1_HVT \keys_reg[5][35]  ( .D(n2928), .CLK(clk), .Q(\keys[5][35] ), .QN(
        n751) );
  DFFX1_HVT \keys_reg[5][34]  ( .D(n2927), .CLK(clk), .Q(\keys[5][34] ), .QN(
        n752) );
  DFFX1_HVT \keys_reg[5][33]  ( .D(n2926), .CLK(clk), .Q(\keys[5][33] ), .QN(
        n753) );
  DFFX1_HVT \keys_reg[5][32]  ( .D(n2925), .CLK(clk), .Q(\keys[5][32] ), .QN(
        n754) );
  DFFX1_HVT \keys_reg[5][31]  ( .D(n2924), .CLK(clk), .Q(\keys[5][31] ), .QN(
        n755) );
  DFFX1_HVT \keys_reg[5][30]  ( .D(n2923), .CLK(clk), .Q(\keys[5][30] ), .QN(
        n756) );
  DFFX1_HVT \keys_reg[5][29]  ( .D(n2922), .CLK(clk), .Q(\keys[5][29] ), .QN(
        n757) );
  DFFX1_HVT \keys_reg[5][28]  ( .D(n2921), .CLK(clk), .Q(\keys[5][28] ), .QN(
        n758) );
  DFFX1_HVT \keys_reg[5][27]  ( .D(n2920), .CLK(clk), .Q(\keys[5][27] ), .QN(
        n759) );
  DFFX1_HVT \keys_reg[5][26]  ( .D(n2919), .CLK(clk), .Q(\keys[5][26] ), .QN(
        n760) );
  DFFX1_HVT \keys_reg[5][25]  ( .D(n2918), .CLK(clk), .Q(\keys[5][25] ), .QN(
        n761) );
  DFFX1_HVT \keys_reg[5][24]  ( .D(n2917), .CLK(clk), .Q(\keys[5][24] ), .QN(
        n762) );
  DFFX1_HVT \keys_reg[5][23]  ( .D(n2916), .CLK(clk), .Q(\keys[5][23] ), .QN(
        n763) );
  DFFX1_HVT \keys_reg[5][22]  ( .D(n2915), .CLK(clk), .Q(\keys[5][22] ), .QN(
        n764) );
  DFFX1_HVT \keys_reg[5][21]  ( .D(n2914), .CLK(clk), .Q(\keys[5][21] ), .QN(
        n765) );
  DFFX1_HVT \keys_reg[5][20]  ( .D(n2913), .CLK(clk), .Q(\keys[5][20] ), .QN(
        n766) );
  DFFX1_HVT \keys_reg[5][19]  ( .D(n2912), .CLK(clk), .Q(\keys[5][19] ), .QN(
        n767) );
  DFFX1_HVT \keys_reg[5][18]  ( .D(n2911), .CLK(clk), .Q(\keys[5][18] ), .QN(
        n768) );
  DFFX1_HVT \keys_reg[5][17]  ( .D(n2910), .CLK(clk), .Q(\keys[5][17] ), .QN(
        n769) );
  DFFX1_HVT \keys_reg[5][16]  ( .D(n2909), .CLK(clk), .Q(\keys[5][16] ), .QN(
        n770) );
  DFFX1_HVT \keys_reg[5][15]  ( .D(n2908), .CLK(clk), .Q(\keys[5][15] ), .QN(
        n771) );
  DFFX1_HVT \keys_reg[5][14]  ( .D(n2907), .CLK(clk), .Q(\keys[5][14] ), .QN(
        n772) );
  DFFX1_HVT \keys_reg[5][13]  ( .D(n2906), .CLK(clk), .Q(\keys[5][13] ), .QN(
        n773) );
  DFFX1_HVT \keys_reg[5][12]  ( .D(n2905), .CLK(clk), .Q(\keys[5][12] ), .QN(
        n774) );
  DFFX1_HVT \keys_reg[5][11]  ( .D(n2904), .CLK(clk), .Q(\keys[5][11] ), .QN(
        n775) );
  DFFX1_HVT \keys_reg[5][10]  ( .D(n2903), .CLK(clk), .Q(\keys[5][10] ), .QN(
        n776) );
  DFFX1_HVT \keys_reg[5][9]  ( .D(n2902), .CLK(clk), .Q(\keys[5][9] ), .QN(
        n777) );
  DFFX1_HVT \keys_reg[5][8]  ( .D(n2901), .CLK(clk), .Q(\keys[5][8] ), .QN(
        n778) );
  DFFX1_HVT \keys_reg[5][7]  ( .D(n2900), .CLK(clk), .Q(\keys[5][7] ), .QN(
        n779) );
  DFFX1_HVT \keys_reg[5][6]  ( .D(n2899), .CLK(clk), .Q(\keys[5][6] ), .QN(
        n780) );
  DFFX1_HVT \keys_reg[5][5]  ( .D(n2898), .CLK(clk), .Q(\keys[5][5] ), .QN(
        n781) );
  DFFX1_HVT \keys_reg[5][4]  ( .D(n2897), .CLK(clk), .Q(\keys[5][4] ), .QN(
        n782) );
  DFFX1_HVT \keys_reg[5][3]  ( .D(n2896), .CLK(clk), .Q(\keys[5][3] ), .QN(
        n783) );
  DFFX1_HVT \keys_reg[5][2]  ( .D(n2895), .CLK(clk), .Q(\keys[5][2] ), .QN(
        n784) );
  DFFX1_HVT \keys_reg[5][1]  ( .D(n2894), .CLK(clk), .Q(\keys[5][1] ), .QN(
        n785) );
  DFFX1_HVT \keys_reg[5][0]  ( .D(n2893), .CLK(clk), .Q(\keys[5][0] ), .QN(
        n786) );
  DFFX1_HVT \keys_reg[6][127]  ( .D(n2892), .CLK(clk), .Q(\keys[6][127] ), 
        .QN(n787) );
  DFFX1_HVT \keys_reg[6][126]  ( .D(n2891), .CLK(clk), .Q(\keys[6][126] ), 
        .QN(n788) );
  DFFX1_HVT \keys_reg[6][125]  ( .D(n2890), .CLK(clk), .Q(\keys[6][125] ), 
        .QN(n789) );
  DFFX1_HVT \keys_reg[6][124]  ( .D(n2889), .CLK(clk), .Q(\keys[6][124] ), 
        .QN(n790) );
  DFFX1_HVT \keys_reg[6][123]  ( .D(n2888), .CLK(clk), .Q(\keys[6][123] ), 
        .QN(n791) );
  DFFX1_HVT \keys_reg[6][122]  ( .D(n2887), .CLK(clk), .Q(\keys[6][122] ), 
        .QN(n792) );
  DFFX1_HVT \keys_reg[6][121]  ( .D(n2886), .CLK(clk), .Q(\keys[6][121] ), 
        .QN(n793) );
  DFFX1_HVT \keys_reg[6][120]  ( .D(n2885), .CLK(clk), .Q(\keys[6][120] ), 
        .QN(n794) );
  DFFX1_HVT \keys_reg[6][119]  ( .D(n2884), .CLK(clk), .Q(\keys[6][119] ), 
        .QN(n795) );
  DFFX1_HVT \keys_reg[6][118]  ( .D(n2883), .CLK(clk), .Q(\keys[6][118] ), 
        .QN(n796) );
  DFFX1_HVT \keys_reg[6][117]  ( .D(n2882), .CLK(clk), .Q(\keys[6][117] ), 
        .QN(n797) );
  DFFX1_HVT \keys_reg[6][116]  ( .D(n2881), .CLK(clk), .Q(\keys[6][116] ), 
        .QN(n798) );
  DFFX1_HVT \keys_reg[6][115]  ( .D(n2880), .CLK(clk), .Q(\keys[6][115] ), 
        .QN(n799) );
  DFFX1_HVT \keys_reg[6][114]  ( .D(n2879), .CLK(clk), .Q(\keys[6][114] ), 
        .QN(n800) );
  DFFX1_HVT \keys_reg[6][113]  ( .D(n2878), .CLK(clk), .Q(\keys[6][113] ), 
        .QN(n801) );
  DFFX1_HVT \keys_reg[6][112]  ( .D(n2877), .CLK(clk), .Q(\keys[6][112] ), 
        .QN(n802) );
  DFFX1_HVT \keys_reg[6][111]  ( .D(n2876), .CLK(clk), .Q(\keys[6][111] ), 
        .QN(n803) );
  DFFX1_HVT \keys_reg[6][110]  ( .D(n2875), .CLK(clk), .Q(\keys[6][110] ), 
        .QN(n804) );
  DFFX1_HVT \keys_reg[6][109]  ( .D(n2874), .CLK(clk), .Q(\keys[6][109] ), 
        .QN(n805) );
  DFFX1_HVT \keys_reg[6][108]  ( .D(n2873), .CLK(clk), .QN(n806) );
  DFFX1_HVT \keys_reg[6][107]  ( .D(n2872), .CLK(clk), .Q(\keys[6][107] ), 
        .QN(n807) );
  DFFX1_HVT \keys_reg[6][106]  ( .D(n2871), .CLK(clk), .Q(\keys[6][106] ), 
        .QN(n808) );
  DFFX1_HVT \keys_reg[6][105]  ( .D(n2870), .CLK(clk), .Q(\keys[6][105] ), 
        .QN(n809) );
  DFFX1_HVT \keys_reg[6][104]  ( .D(n2869), .CLK(clk), .Q(\keys[6][104] ), 
        .QN(n810) );
  DFFX1_HVT \keys_reg[6][103]  ( .D(n2868), .CLK(clk), .Q(\keys[6][103] ), 
        .QN(n811) );
  DFFX1_HVT \keys_reg[6][102]  ( .D(n2867), .CLK(clk), .Q(\keys[6][102] ), 
        .QN(n812) );
  DFFX1_HVT \keys_reg[6][101]  ( .D(n2866), .CLK(clk), .Q(\keys[6][101] ), 
        .QN(n813) );
  DFFX1_HVT \keys_reg[6][100]  ( .D(n2865), .CLK(clk), .Q(\keys[6][100] ), 
        .QN(n814) );
  DFFX1_HVT \keys_reg[6][99]  ( .D(n2864), .CLK(clk), .Q(\keys[6][99] ), .QN(
        n815) );
  DFFX1_HVT \keys_reg[6][98]  ( .D(n2863), .CLK(clk), .Q(\keys[6][98] ), .QN(
        n816) );
  DFFX1_HVT \keys_reg[6][97]  ( .D(n2862), .CLK(clk), .Q(\keys[6][97] ), .QN(
        n817) );
  DFFX1_HVT \keys_reg[6][96]  ( .D(n2861), .CLK(clk), .Q(\keys[6][96] ), .QN(
        n818) );
  DFFX1_HVT \keys_reg[6][95]  ( .D(n2860), .CLK(clk), .Q(\keys[6][95] ), .QN(
        n819) );
  DFFX1_HVT \keys_reg[6][94]  ( .D(n2859), .CLK(clk), .Q(\keys[6][94] ), .QN(
        n820) );
  DFFX1_HVT \keys_reg[6][93]  ( .D(n2858), .CLK(clk), .Q(\keys[6][93] ), .QN(
        n821) );
  DFFX1_HVT \keys_reg[6][92]  ( .D(n2857), .CLK(clk), .Q(\keys[6][92] ), .QN(
        n822) );
  DFFX1_HVT \keys_reg[6][91]  ( .D(n2856), .CLK(clk), .Q(\keys[6][91] ), .QN(
        n823) );
  DFFX1_HVT \keys_reg[6][90]  ( .D(n2855), .CLK(clk), .Q(\keys[6][90] ), .QN(
        n824) );
  DFFX1_HVT \keys_reg[6][89]  ( .D(n2854), .CLK(clk), .Q(\keys[6][89] ), .QN(
        n825) );
  DFFX1_HVT \keys_reg[6][88]  ( .D(n2853), .CLK(clk), .Q(\keys[6][88] ), .QN(
        n826) );
  DFFX1_HVT \keys_reg[6][87]  ( .D(n2852), .CLK(clk), .Q(\keys[6][87] ), .QN(
        n827) );
  DFFX1_HVT \keys_reg[6][86]  ( .D(n2851), .CLK(clk), .Q(\keys[6][86] ), .QN(
        n828) );
  DFFX1_HVT \keys_reg[6][85]  ( .D(n2850), .CLK(clk), .Q(\keys[6][85] ), .QN(
        n829) );
  DFFX1_HVT \keys_reg[6][84]  ( .D(n2849), .CLK(clk), .Q(\keys[6][84] ), .QN(
        n830) );
  DFFX1_HVT \keys_reg[6][83]  ( .D(n2848), .CLK(clk), .Q(\keys[6][83] ), .QN(
        n831) );
  DFFX1_HVT \keys_reg[6][82]  ( .D(n2847), .CLK(clk), .Q(\keys[6][82] ), .QN(
        n832) );
  DFFX1_HVT \keys_reg[6][81]  ( .D(n2846), .CLK(clk), .Q(\keys[6][81] ), .QN(
        n833) );
  DFFX1_HVT \keys_reg[6][80]  ( .D(n2845), .CLK(clk), .Q(\keys[6][80] ), .QN(
        n834) );
  DFFX1_HVT \keys_reg[6][79]  ( .D(n2844), .CLK(clk), .Q(\keys[6][79] ), .QN(
        n835) );
  DFFX1_HVT \keys_reg[6][78]  ( .D(n2843), .CLK(clk), .Q(\keys[6][78] ), .QN(
        n836) );
  DFFX1_HVT \keys_reg[6][77]  ( .D(n2842), .CLK(clk), .Q(\keys[6][77] ), .QN(
        n837) );
  DFFX1_HVT \keys_reg[6][76]  ( .D(n2841), .CLK(clk), .Q(\keys[6][76] ), .QN(
        n838) );
  DFFX1_HVT \keys_reg[6][75]  ( .D(n2840), .CLK(clk), .Q(\keys[6][75] ), .QN(
        n839) );
  DFFX1_HVT \keys_reg[6][74]  ( .D(n2839), .CLK(clk), .Q(\keys[6][74] ), .QN(
        n840) );
  DFFX1_HVT \keys_reg[6][73]  ( .D(n2838), .CLK(clk), .Q(\keys[6][73] ), .QN(
        n841) );
  DFFX1_HVT \keys_reg[6][72]  ( .D(n2837), .CLK(clk), .Q(\keys[6][72] ), .QN(
        n842) );
  DFFX1_HVT \keys_reg[6][71]  ( .D(n2836), .CLK(clk), .Q(\keys[6][71] ), .QN(
        n843) );
  DFFX1_HVT \keys_reg[6][70]  ( .D(n2835), .CLK(clk), .Q(\keys[6][70] ), .QN(
        n844) );
  DFFX1_HVT \keys_reg[6][69]  ( .D(n2834), .CLK(clk), .Q(\keys[6][69] ), .QN(
        n845) );
  DFFX1_HVT \keys_reg[6][68]  ( .D(n2833), .CLK(clk), .Q(\keys[6][68] ), .QN(
        n846) );
  DFFX1_HVT \keys_reg[6][67]  ( .D(n2832), .CLK(clk), .Q(\keys[6][67] ), .QN(
        n847) );
  DFFX1_HVT \keys_reg[6][66]  ( .D(n2831), .CLK(clk), .Q(\keys[6][66] ), .QN(
        n848) );
  DFFX1_HVT \keys_reg[6][65]  ( .D(n2830), .CLK(clk), .Q(\keys[6][65] ), .QN(
        n849) );
  DFFX1_HVT \keys_reg[6][64]  ( .D(n2829), .CLK(clk), .Q(\keys[6][64] ), .QN(
        n850) );
  DFFX1_HVT \keys_reg[6][63]  ( .D(n2828), .CLK(clk), .Q(\keys[6][63] ), .QN(
        n851) );
  DFFX1_HVT \keys_reg[6][62]  ( .D(n2827), .CLK(clk), .Q(\keys[6][62] ), .QN(
        n852) );
  DFFX1_HVT \keys_reg[6][61]  ( .D(n2826), .CLK(clk), .Q(\keys[6][61] ), .QN(
        n853) );
  DFFX1_HVT \keys_reg[6][60]  ( .D(n2825), .CLK(clk), .Q(\keys[6][60] ), .QN(
        n854) );
  DFFX1_HVT \keys_reg[6][59]  ( .D(n2824), .CLK(clk), .Q(\keys[6][59] ), .QN(
        n855) );
  DFFX1_HVT \keys_reg[6][58]  ( .D(n2823), .CLK(clk), .Q(\keys[6][58] ), .QN(
        n856) );
  DFFX1_HVT \keys_reg[6][57]  ( .D(n2822), .CLK(clk), .Q(\keys[6][57] ), .QN(
        n857) );
  DFFX1_HVT \keys_reg[6][56]  ( .D(n2821), .CLK(clk), .Q(\keys[6][56] ), .QN(
        n858) );
  DFFX1_HVT \keys_reg[6][55]  ( .D(n2820), .CLK(clk), .Q(\keys[6][55] ), .QN(
        n859) );
  DFFX1_HVT \keys_reg[6][54]  ( .D(n2819), .CLK(clk), .Q(\keys[6][54] ), .QN(
        n860) );
  DFFX1_HVT \keys_reg[6][53]  ( .D(n2818), .CLK(clk), .Q(\keys[6][53] ), .QN(
        n861) );
  DFFX1_HVT \keys_reg[6][52]  ( .D(n2817), .CLK(clk), .Q(\keys[6][52] ), .QN(
        n862) );
  DFFX1_HVT \keys_reg[6][51]  ( .D(n2816), .CLK(clk), .Q(\keys[6][51] ), .QN(
        n863) );
  DFFX1_HVT \keys_reg[6][50]  ( .D(n2815), .CLK(clk), .Q(\keys[6][50] ), .QN(
        n864) );
  DFFX1_HVT \keys_reg[6][49]  ( .D(n2814), .CLK(clk), .Q(\keys[6][49] ), .QN(
        n865) );
  DFFX1_HVT \keys_reg[6][48]  ( .D(n2813), .CLK(clk), .Q(\keys[6][48] ), .QN(
        n866) );
  DFFX1_HVT \keys_reg[6][47]  ( .D(n2812), .CLK(clk), .Q(\keys[6][47] ), .QN(
        n867) );
  DFFX1_HVT \keys_reg[6][46]  ( .D(n2811), .CLK(clk), .Q(\keys[6][46] ), .QN(
        n868) );
  DFFX1_HVT \keys_reg[6][45]  ( .D(n2810), .CLK(clk), .Q(\keys[6][45] ), .QN(
        n869) );
  DFFX1_HVT \keys_reg[6][44]  ( .D(n2809), .CLK(clk), .Q(\keys[6][44] ), .QN(
        n870) );
  DFFX1_HVT \keys_reg[6][43]  ( .D(n2808), .CLK(clk), .Q(\keys[6][43] ), .QN(
        n871) );
  DFFX1_HVT \keys_reg[6][42]  ( .D(n2807), .CLK(clk), .Q(\keys[6][42] ), .QN(
        n872) );
  DFFX1_HVT \keys_reg[6][41]  ( .D(n2806), .CLK(clk), .Q(\keys[6][41] ), .QN(
        n873) );
  DFFX1_HVT \keys_reg[6][40]  ( .D(n2805), .CLK(clk), .Q(\keys[6][40] ), .QN(
        n874) );
  DFFX1_HVT \keys_reg[6][39]  ( .D(n2804), .CLK(clk), .Q(\keys[6][39] ), .QN(
        n875) );
  DFFX1_HVT \keys_reg[6][38]  ( .D(n2803), .CLK(clk), .Q(\keys[6][38] ), .QN(
        n876) );
  DFFX1_HVT \keys_reg[6][37]  ( .D(n2802), .CLK(clk), .Q(\keys[6][37] ), .QN(
        n877) );
  DFFX1_HVT \keys_reg[6][36]  ( .D(n2801), .CLK(clk), .Q(\keys[6][36] ), .QN(
        n878) );
  DFFX1_HVT \keys_reg[6][35]  ( .D(n2800), .CLK(clk), .Q(\keys[6][35] ), .QN(
        n879) );
  DFFX1_HVT \keys_reg[6][34]  ( .D(n2799), .CLK(clk), .Q(\keys[6][34] ), .QN(
        n880) );
  DFFX1_HVT \keys_reg[6][33]  ( .D(n2798), .CLK(clk), .Q(\keys[6][33] ), .QN(
        n881) );
  DFFX1_HVT \keys_reg[6][32]  ( .D(n2797), .CLK(clk), .Q(\keys[6][32] ), .QN(
        n882) );
  DFFX1_HVT \keys_reg[6][31]  ( .D(n2796), .CLK(clk), .Q(\keys[6][31] ), .QN(
        n883) );
  DFFX1_HVT \keys_reg[6][30]  ( .D(n2795), .CLK(clk), .Q(\keys[6][30] ), .QN(
        n884) );
  DFFX1_HVT \keys_reg[6][29]  ( .D(n2794), .CLK(clk), .Q(\keys[6][29] ), .QN(
        n885) );
  DFFX1_HVT \keys_reg[6][28]  ( .D(n2793), .CLK(clk), .Q(\keys[6][28] ), .QN(
        n886) );
  DFFX1_HVT \keys_reg[6][27]  ( .D(n2792), .CLK(clk), .Q(\keys[6][27] ), .QN(
        n887) );
  DFFX1_HVT \keys_reg[6][26]  ( .D(n2791), .CLK(clk), .Q(\keys[6][26] ), .QN(
        n888) );
  DFFX1_HVT \keys_reg[6][25]  ( .D(n2790), .CLK(clk), .Q(\keys[6][25] ), .QN(
        n889) );
  DFFX1_HVT \keys_reg[6][24]  ( .D(n2789), .CLK(clk), .Q(\keys[6][24] ), .QN(
        n890) );
  DFFX1_HVT \keys_reg[6][23]  ( .D(n2788), .CLK(clk), .Q(\keys[6][23] ), .QN(
        n891) );
  DFFX1_HVT \keys_reg[6][22]  ( .D(n2787), .CLK(clk), .Q(\keys[6][22] ), .QN(
        n892) );
  DFFX1_HVT \keys_reg[6][21]  ( .D(n2786), .CLK(clk), .Q(\keys[6][21] ), .QN(
        n893) );
  DFFX1_HVT \keys_reg[6][20]  ( .D(n2785), .CLK(clk), .Q(\keys[6][20] ), .QN(
        n894) );
  DFFX1_HVT \keys_reg[6][19]  ( .D(n2784), .CLK(clk), .Q(\keys[6][19] ), .QN(
        n895) );
  DFFX1_HVT \keys_reg[6][18]  ( .D(n2783), .CLK(clk), .Q(\keys[6][18] ), .QN(
        n896) );
  DFFX1_HVT \keys_reg[6][17]  ( .D(n2782), .CLK(clk), .Q(\keys[6][17] ), .QN(
        n897) );
  DFFX1_HVT \keys_reg[6][16]  ( .D(n2781), .CLK(clk), .Q(\keys[6][16] ), .QN(
        n898) );
  DFFX1_HVT \keys_reg[6][15]  ( .D(n2780), .CLK(clk), .Q(\keys[6][15] ), .QN(
        n899) );
  DFFX1_HVT \keys_reg[6][14]  ( .D(n2779), .CLK(clk), .Q(\keys[6][14] ), .QN(
        n900) );
  DFFX1_HVT \keys_reg[6][13]  ( .D(n2778), .CLK(clk), .Q(\keys[6][13] ), .QN(
        n901) );
  DFFX1_HVT \keys_reg[6][12]  ( .D(n2777), .CLK(clk), .Q(\keys[6][12] ), .QN(
        n902) );
  DFFX1_HVT \keys_reg[6][11]  ( .D(n2776), .CLK(clk), .Q(\keys[6][11] ), .QN(
        n903) );
  DFFX1_HVT \keys_reg[6][10]  ( .D(n2775), .CLK(clk), .Q(\keys[6][10] ), .QN(
        n904) );
  DFFX1_HVT \keys_reg[6][9]  ( .D(n2774), .CLK(clk), .Q(\keys[6][9] ), .QN(
        n905) );
  DFFX1_HVT \keys_reg[6][8]  ( .D(n2773), .CLK(clk), .Q(\keys[6][8] ), .QN(
        n906) );
  DFFX1_HVT \keys_reg[6][7]  ( .D(n2772), .CLK(clk), .Q(\keys[6][7] ), .QN(
        n907) );
  DFFX1_HVT \keys_reg[6][6]  ( .D(n2771), .CLK(clk), .Q(\keys[6][6] ), .QN(
        n908) );
  DFFX1_HVT \keys_reg[6][5]  ( .D(n2770), .CLK(clk), .Q(\keys[6][5] ), .QN(
        n909) );
  DFFX1_HVT \keys_reg[6][4]  ( .D(n2769), .CLK(clk), .Q(\keys[6][4] ), .QN(
        n910) );
  DFFX1_HVT \keys_reg[6][3]  ( .D(n2768), .CLK(clk), .Q(\keys[6][3] ), .QN(
        n911) );
  DFFX1_HVT \keys_reg[6][2]  ( .D(n2767), .CLK(clk), .Q(\keys[6][2] ), .QN(
        n912) );
  DFFX1_HVT \keys_reg[6][1]  ( .D(n2766), .CLK(clk), .Q(\keys[6][1] ), .QN(
        n913) );
  DFFX1_HVT \keys_reg[6][0]  ( .D(n2765), .CLK(clk), .Q(\keys[6][0] ), .QN(
        n914) );
  DFFX1_HVT \keys_reg[7][127]  ( .D(n2764), .CLK(clk), .Q(\keys[7][127] ), 
        .QN(n915) );
  DFFX1_HVT \keys_reg[7][126]  ( .D(n2763), .CLK(clk), .Q(\keys[7][126] ), 
        .QN(n916) );
  DFFX1_HVT \keys_reg[7][125]  ( .D(n2762), .CLK(clk), .Q(\keys[7][125] ), 
        .QN(n917) );
  DFFX1_HVT \keys_reg[7][124]  ( .D(n2761), .CLK(clk), .Q(\keys[7][124] ), 
        .QN(n918) );
  DFFX1_HVT \keys_reg[7][123]  ( .D(n2760), .CLK(clk), .Q(\keys[7][123] ), 
        .QN(n919) );
  DFFX1_HVT \keys_reg[7][122]  ( .D(n2759), .CLK(clk), .Q(\keys[7][122] ), 
        .QN(n920) );
  DFFX1_HVT \keys_reg[7][121]  ( .D(n2758), .CLK(clk), .Q(\keys[7][121] ), 
        .QN(n921) );
  DFFX1_HVT \keys_reg[7][120]  ( .D(n2757), .CLK(clk), .Q(\keys[7][120] ), 
        .QN(n922) );
  DFFX1_HVT \keys_reg[7][119]  ( .D(n2756), .CLK(clk), .Q(\keys[7][119] ), 
        .QN(n923) );
  DFFX1_HVT \keys_reg[7][118]  ( .D(n2755), .CLK(clk), .Q(\keys[7][118] ), 
        .QN(n924) );
  DFFX1_HVT \keys_reg[7][117]  ( .D(n2754), .CLK(clk), .Q(\keys[7][117] ), 
        .QN(n925) );
  DFFX1_HVT \keys_reg[7][116]  ( .D(n2753), .CLK(clk), .Q(\keys[7][116] ), 
        .QN(n926) );
  DFFX1_HVT \keys_reg[7][115]  ( .D(n2752), .CLK(clk), .Q(\keys[7][115] ), 
        .QN(n927) );
  DFFX1_HVT \keys_reg[7][114]  ( .D(n2751), .CLK(clk), .Q(\keys[7][114] ), 
        .QN(n928) );
  DFFX1_HVT \keys_reg[7][113]  ( .D(n2750), .CLK(clk), .Q(\keys[7][113] ), 
        .QN(n929) );
  DFFX1_HVT \keys_reg[7][112]  ( .D(n2749), .CLK(clk), .Q(\keys[7][112] ), 
        .QN(n930) );
  DFFX1_HVT \keys_reg[7][111]  ( .D(n2748), .CLK(clk), .Q(\keys[7][111] ), 
        .QN(n931) );
  DFFX1_HVT \keys_reg[7][110]  ( .D(n2747), .CLK(clk), .Q(\keys[7][110] ), 
        .QN(n932) );
  DFFX1_HVT \keys_reg[7][109]  ( .D(n2746), .CLK(clk), .Q(\keys[7][109] ), 
        .QN(n933) );
  DFFX1_HVT \keys_reg[7][108]  ( .D(n2745), .CLK(clk), .Q(\keys[7][108] ), 
        .QN(n934) );
  DFFX1_HVT \keys_reg[7][107]  ( .D(n2744), .CLK(clk), .Q(\keys[7][107] ), 
        .QN(n935) );
  DFFX1_HVT \keys_reg[7][106]  ( .D(n2743), .CLK(clk), .Q(\keys[7][106] ), 
        .QN(n936) );
  DFFX1_HVT \keys_reg[7][105]  ( .D(n2742), .CLK(clk), .Q(\keys[7][105] ), 
        .QN(n937) );
  DFFX1_HVT \keys_reg[7][104]  ( .D(n2741), .CLK(clk), .Q(\keys[7][104] ), 
        .QN(n938) );
  DFFX1_HVT \keys_reg[7][103]  ( .D(n2740), .CLK(clk), .Q(\keys[7][103] ), 
        .QN(n939) );
  DFFX1_HVT \keys_reg[7][102]  ( .D(n2739), .CLK(clk), .Q(\keys[7][102] ), 
        .QN(n940) );
  DFFX1_HVT \keys_reg[7][101]  ( .D(n2738), .CLK(clk), .Q(\keys[7][101] ), 
        .QN(n941) );
  DFFX1_HVT \keys_reg[7][100]  ( .D(n2737), .CLK(clk), .Q(\keys[7][100] ), 
        .QN(n942) );
  DFFX1_HVT \keys_reg[7][99]  ( .D(n2736), .CLK(clk), .Q(\keys[7][99] ), .QN(
        n943) );
  DFFX1_HVT \keys_reg[7][98]  ( .D(n2735), .CLK(clk), .Q(\keys[7][98] ), .QN(
        n944) );
  DFFX1_HVT \keys_reg[7][97]  ( .D(n2734), .CLK(clk), .Q(\keys[7][97] ), .QN(
        n945) );
  DFFX1_HVT \keys_reg[7][96]  ( .D(n2733), .CLK(clk), .Q(\keys[7][96] ), .QN(
        n946) );
  DFFX1_HVT \keys_reg[7][95]  ( .D(n2732), .CLK(clk), .Q(\keys[7][95] ), .QN(
        n947) );
  DFFX1_HVT \keys_reg[7][94]  ( .D(n2731), .CLK(clk), .Q(\keys[7][94] ), .QN(
        n948) );
  DFFX1_HVT \keys_reg[7][93]  ( .D(n2730), .CLK(clk), .Q(\keys[7][93] ), .QN(
        n949) );
  DFFX1_HVT \keys_reg[7][92]  ( .D(n2729), .CLK(clk), .Q(\keys[7][92] ), .QN(
        n950) );
  DFFX1_HVT \keys_reg[7][91]  ( .D(n2728), .CLK(clk), .Q(\keys[7][91] ), .QN(
        n951) );
  DFFX1_HVT \keys_reg[7][90]  ( .D(n2727), .CLK(clk), .Q(\keys[7][90] ), .QN(
        n952) );
  DFFX1_HVT \keys_reg[7][89]  ( .D(n2726), .CLK(clk), .Q(\keys[7][89] ), .QN(
        n953) );
  DFFX1_HVT \keys_reg[7][88]  ( .D(n2725), .CLK(clk), .Q(\keys[7][88] ), .QN(
        n954) );
  DFFX1_HVT \keys_reg[7][87]  ( .D(n2724), .CLK(clk), .Q(\keys[7][87] ), .QN(
        n955) );
  DFFX1_HVT \keys_reg[7][86]  ( .D(n2723), .CLK(clk), .Q(\keys[7][86] ), .QN(
        n956) );
  DFFX1_HVT \keys_reg[7][85]  ( .D(n2722), .CLK(clk), .Q(\keys[7][85] ), .QN(
        n957) );
  DFFX1_HVT \keys_reg[7][84]  ( .D(n2721), .CLK(clk), .Q(\keys[7][84] ), .QN(
        n958) );
  DFFX1_HVT \keys_reg[7][83]  ( .D(n2720), .CLK(clk), .Q(\keys[7][83] ), .QN(
        n959) );
  DFFX1_HVT \keys_reg[7][82]  ( .D(n2719), .CLK(clk), .Q(\keys[7][82] ), .QN(
        n960) );
  DFFX1_HVT \keys_reg[7][81]  ( .D(n2718), .CLK(clk), .Q(\keys[7][81] ), .QN(
        n961) );
  DFFX1_HVT \keys_reg[7][80]  ( .D(n2717), .CLK(clk), .Q(\keys[7][80] ), .QN(
        n962) );
  DFFX1_HVT \keys_reg[7][79]  ( .D(n2716), .CLK(clk), .QN(n963) );
  DFFX1_HVT \keys_reg[7][78]  ( .D(n2715), .CLK(clk), .Q(\keys[7][78] ), .QN(
        n964) );
  DFFX1_HVT \keys_reg[7][77]  ( .D(n2714), .CLK(clk), .Q(\keys[7][77] ), .QN(
        n965) );
  DFFX1_HVT \keys_reg[7][76]  ( .D(n2713), .CLK(clk), .Q(\keys[7][76] ), .QN(
        n966) );
  DFFX1_HVT \keys_reg[7][75]  ( .D(n2712), .CLK(clk), .Q(\keys[7][75] ), .QN(
        n967) );
  DFFX1_HVT \keys_reg[7][74]  ( .D(n2711), .CLK(clk), .QN(n968) );
  DFFX1_HVT \keys_reg[7][73]  ( .D(n2710), .CLK(clk), .QN(n969) );
  DFFX1_HVT \keys_reg[7][72]  ( .D(n2709), .CLK(clk), .Q(\keys[7][72] ), .QN(
        n970) );
  DFFX1_HVT \keys_reg[7][71]  ( .D(n2708), .CLK(clk), .Q(\keys[7][71] ), .QN(
        n971) );
  DFFX1_HVT \keys_reg[7][70]  ( .D(n2707), .CLK(clk), .Q(\keys[7][70] ), .QN(
        n972) );
  DFFX1_HVT \keys_reg[7][69]  ( .D(n2706), .CLK(clk), .Q(\keys[7][69] ), .QN(
        n973) );
  DFFX1_HVT \keys_reg[7][68]  ( .D(n2705), .CLK(clk), .Q(\keys[7][68] ), .QN(
        n974) );
  DFFX1_HVT \keys_reg[7][67]  ( .D(n2704), .CLK(clk), .Q(\keys[7][67] ), .QN(
        n975) );
  DFFX1_HVT \keys_reg[7][66]  ( .D(n2703), .CLK(clk), .Q(\keys[7][66] ), .QN(
        n976) );
  DFFX1_HVT \keys_reg[7][65]  ( .D(n2702), .CLK(clk), .Q(\keys[7][65] ), .QN(
        n977) );
  DFFX1_HVT \keys_reg[7][64]  ( .D(n2701), .CLK(clk), .Q(\keys[7][64] ), .QN(
        n978) );
  DFFX1_HVT \keys_reg[7][63]  ( .D(n2700), .CLK(clk), .Q(\keys[7][63] ), .QN(
        n979) );
  DFFX1_HVT \keys_reg[7][62]  ( .D(n2699), .CLK(clk), .Q(\keys[7][62] ), .QN(
        n980) );
  DFFX1_HVT \keys_reg[7][61]  ( .D(n2698), .CLK(clk), .Q(\keys[7][61] ), .QN(
        n981) );
  DFFX1_HVT \keys_reg[7][60]  ( .D(n2697), .CLK(clk), .Q(\keys[7][60] ), .QN(
        n982) );
  DFFX1_HVT \keys_reg[7][59]  ( .D(n2696), .CLK(clk), .Q(\keys[7][59] ), .QN(
        n983) );
  DFFX1_HVT \keys_reg[7][58]  ( .D(n2695), .CLK(clk), .Q(\keys[7][58] ), .QN(
        n984) );
  DFFX1_HVT \keys_reg[7][57]  ( .D(n2694), .CLK(clk), .Q(\keys[7][57] ), .QN(
        n985) );
  DFFX1_HVT \keys_reg[7][56]  ( .D(n2693), .CLK(clk), .Q(\keys[7][56] ), .QN(
        n986) );
  DFFX1_HVT \keys_reg[7][55]  ( .D(n2692), .CLK(clk), .Q(\keys[7][55] ), .QN(
        n987) );
  DFFX1_HVT \keys_reg[7][54]  ( .D(n2691), .CLK(clk), .Q(\keys[7][54] ), .QN(
        n988) );
  DFFX1_HVT \keys_reg[7][53]  ( .D(n2690), .CLK(clk), .Q(\keys[7][53] ), .QN(
        n989) );
  DFFX1_HVT \keys_reg[7][52]  ( .D(n2689), .CLK(clk), .Q(\keys[7][52] ), .QN(
        n990) );
  DFFX1_HVT \keys_reg[7][51]  ( .D(n2688), .CLK(clk), .Q(\keys[7][51] ), .QN(
        n991) );
  DFFX1_HVT \keys_reg[7][50]  ( .D(n2687), .CLK(clk), .Q(\keys[7][50] ), .QN(
        n992) );
  DFFX1_HVT \keys_reg[7][49]  ( .D(n2686), .CLK(clk), .Q(\keys[7][49] ), .QN(
        n993) );
  DFFX1_HVT \keys_reg[7][48]  ( .D(n2685), .CLK(clk), .Q(\keys[7][48] ), .QN(
        n994) );
  DFFX1_HVT \keys_reg[7][47]  ( .D(n2684), .CLK(clk), .Q(\keys[7][47] ), .QN(
        n995) );
  DFFX1_HVT \keys_reg[7][46]  ( .D(n2683), .CLK(clk), .Q(\keys[7][46] ), .QN(
        n996) );
  DFFX1_HVT \keys_reg[7][45]  ( .D(n2682), .CLK(clk), .Q(\keys[7][45] ), .QN(
        n997) );
  DFFX1_HVT \keys_reg[7][44]  ( .D(n2681), .CLK(clk), .Q(\keys[7][44] ), .QN(
        n998) );
  DFFX1_HVT \keys_reg[7][43]  ( .D(n2680), .CLK(clk), .Q(\keys[7][43] ), .QN(
        n999) );
  DFFX1_HVT \keys_reg[7][42]  ( .D(n2679), .CLK(clk), .Q(\keys[7][42] ), .QN(
        n1000) );
  DFFX1_HVT \keys_reg[7][41]  ( .D(n2678), .CLK(clk), .Q(\keys[7][41] ), .QN(
        n1001) );
  DFFX1_HVT \keys_reg[7][40]  ( .D(n2677), .CLK(clk), .Q(\keys[7][40] ), .QN(
        n1002) );
  DFFX1_HVT \keys_reg[7][39]  ( .D(n2676), .CLK(clk), .Q(\keys[7][39] ), .QN(
        n1003) );
  DFFX1_HVT \keys_reg[7][38]  ( .D(n2675), .CLK(clk), .Q(\keys[7][38] ), .QN(
        n1004) );
  DFFX1_HVT \keys_reg[7][37]  ( .D(n2674), .CLK(clk), .Q(\keys[7][37] ), .QN(
        n1005) );
  DFFX1_HVT \keys_reg[7][36]  ( .D(n2673), .CLK(clk), .Q(\keys[7][36] ), .QN(
        n1006) );
  DFFX1_HVT \keys_reg[7][35]  ( .D(n2672), .CLK(clk), .Q(\keys[7][35] ), .QN(
        n1007) );
  DFFX1_HVT \keys_reg[7][34]  ( .D(n2671), .CLK(clk), .Q(\keys[7][34] ), .QN(
        n1008) );
  DFFX1_HVT \keys_reg[7][33]  ( .D(n2670), .CLK(clk), .Q(\keys[7][33] ), .QN(
        n1009) );
  DFFX1_HVT \keys_reg[7][32]  ( .D(n2669), .CLK(clk), .Q(\keys[7][32] ), .QN(
        n1010) );
  DFFX1_HVT \keys_reg[7][31]  ( .D(n2668), .CLK(clk), .Q(\keys[7][31] ), .QN(
        n1011) );
  DFFX1_HVT \keys_reg[7][30]  ( .D(n2667), .CLK(clk), .Q(\keys[7][30] ), .QN(
        n1012) );
  DFFX1_HVT \keys_reg[7][29]  ( .D(n2666), .CLK(clk), .Q(\keys[7][29] ), .QN(
        n1013) );
  DFFX1_HVT \keys_reg[7][28]  ( .D(n2665), .CLK(clk), .Q(\keys[7][28] ), .QN(
        n1014) );
  DFFX1_HVT \keys_reg[7][27]  ( .D(n2664), .CLK(clk), .Q(\keys[7][27] ), .QN(
        n1015) );
  DFFX1_HVT \keys_reg[7][26]  ( .D(n2663), .CLK(clk), .Q(\keys[7][26] ), .QN(
        n1016) );
  DFFX1_HVT \keys_reg[7][25]  ( .D(n2662), .CLK(clk), .Q(\keys[7][25] ), .QN(
        n1017) );
  DFFX1_HVT \keys_reg[7][24]  ( .D(n2661), .CLK(clk), .Q(\keys[7][24] ), .QN(
        n1018) );
  DFFX1_HVT \keys_reg[7][23]  ( .D(n2660), .CLK(clk), .Q(\keys[7][23] ), .QN(
        n1019) );
  DFFX1_HVT \keys_reg[7][22]  ( .D(n2659), .CLK(clk), .Q(\keys[7][22] ), .QN(
        n1020) );
  DFFX1_HVT \keys_reg[7][21]  ( .D(n2658), .CLK(clk), .Q(\keys[7][21] ), .QN(
        n1021) );
  DFFX1_HVT \keys_reg[7][20]  ( .D(n2657), .CLK(clk), .Q(\keys[7][20] ), .QN(
        n1022) );
  DFFX1_HVT \keys_reg[7][19]  ( .D(n2656), .CLK(clk), .Q(\keys[7][19] ), .QN(
        n1023) );
  DFFX1_HVT \keys_reg[7][18]  ( .D(n2655), .CLK(clk), .Q(\keys[7][18] ), .QN(
        n1024) );
  DFFX1_HVT \keys_reg[7][17]  ( .D(n2654), .CLK(clk), .Q(\keys[7][17] ), .QN(
        n1025) );
  DFFX1_HVT \keys_reg[7][16]  ( .D(n2653), .CLK(clk), .Q(\keys[7][16] ), .QN(
        n1026) );
  DFFX1_HVT \keys_reg[7][15]  ( .D(n2652), .CLK(clk), .Q(\keys[7][15] ), .QN(
        n1027) );
  DFFX1_HVT \keys_reg[7][14]  ( .D(n2651), .CLK(clk), .Q(\keys[7][14] ), .QN(
        n1028) );
  DFFX1_HVT \keys_reg[7][13]  ( .D(n2650), .CLK(clk), .Q(\keys[7][13] ), .QN(
        n1029) );
  DFFX1_HVT \keys_reg[7][12]  ( .D(n2649), .CLK(clk), .Q(\keys[7][12] ), .QN(
        n1030) );
  DFFX1_HVT \keys_reg[7][11]  ( .D(n2648), .CLK(clk), .Q(\keys[7][11] ), .QN(
        n1031) );
  DFFX1_HVT \keys_reg[7][10]  ( .D(n2647), .CLK(clk), .Q(\keys[7][10] ), .QN(
        n1032) );
  DFFX1_HVT \keys_reg[7][9]  ( .D(n2646), .CLK(clk), .Q(\keys[7][9] ), .QN(
        n1033) );
  DFFX1_HVT \keys_reg[7][8]  ( .D(n2645), .CLK(clk), .Q(\keys[7][8] ), .QN(
        n1034) );
  DFFX1_HVT \keys_reg[7][7]  ( .D(n2644), .CLK(clk), .Q(\keys[7][7] ), .QN(
        n1035) );
  DFFX1_HVT \keys_reg[7][6]  ( .D(n2643), .CLK(clk), .Q(\keys[7][6] ), .QN(
        n1036) );
  DFFX1_HVT \keys_reg[7][5]  ( .D(n2642), .CLK(clk), .Q(\keys[7][5] ), .QN(
        n1037) );
  DFFX1_HVT \keys_reg[7][4]  ( .D(n2641), .CLK(clk), .Q(\keys[7][4] ), .QN(
        n1038) );
  DFFX1_HVT \keys_reg[7][3]  ( .D(n2640), .CLK(clk), .Q(\keys[7][3] ), .QN(
        n1039) );
  DFFX1_HVT \keys_reg[7][2]  ( .D(n2639), .CLK(clk), .Q(\keys[7][2] ), .QN(
        n1040) );
  DFFX1_HVT \keys_reg[7][1]  ( .D(n2638), .CLK(clk), .Q(\keys[7][1] ), .QN(
        n1041) );
  DFFX1_HVT \keys_reg[7][0]  ( .D(n2637), .CLK(clk), .Q(\keys[7][0] ), .QN(
        n1042) );
  DFFX1_HVT \keys_reg[8][127]  ( .D(n2636), .CLK(clk), .Q(\keys[8][127] ), 
        .QN(n1043) );
  DFFX1_HVT \keys_reg[8][126]  ( .D(n2635), .CLK(clk), .Q(\keys[8][126] ), 
        .QN(n1044) );
  DFFX1_HVT \keys_reg[8][125]  ( .D(n2634), .CLK(clk), .Q(\keys[8][125] ), 
        .QN(n1045) );
  DFFX1_HVT \keys_reg[8][124]  ( .D(n2633), .CLK(clk), .Q(\keys[8][124] ), 
        .QN(n1046) );
  DFFX1_HVT \keys_reg[8][123]  ( .D(n2632), .CLK(clk), .Q(\keys[8][123] ), 
        .QN(n1047) );
  DFFX1_HVT \keys_reg[8][122]  ( .D(n2631), .CLK(clk), .Q(\keys[8][122] ), 
        .QN(n1048) );
  DFFX1_HVT \keys_reg[8][121]  ( .D(n2630), .CLK(clk), .Q(\keys[8][121] ), 
        .QN(n1049) );
  DFFX1_HVT \keys_reg[8][120]  ( .D(n2629), .CLK(clk), .Q(\keys[8][120] ), 
        .QN(n1050) );
  DFFX1_HVT \keys_reg[8][119]  ( .D(n2628), .CLK(clk), .Q(\keys[8][119] ), 
        .QN(n1051) );
  DFFX1_HVT \keys_reg[8][118]  ( .D(n2627), .CLK(clk), .Q(\keys[8][118] ), 
        .QN(n1052) );
  DFFX1_HVT \keys_reg[8][117]  ( .D(n2626), .CLK(clk), .Q(\keys[8][117] ), 
        .QN(n1053) );
  DFFX1_HVT \keys_reg[8][116]  ( .D(n2625), .CLK(clk), .Q(\keys[8][116] ), 
        .QN(n1054) );
  DFFX1_HVT \keys_reg[8][115]  ( .D(n2624), .CLK(clk), .Q(\keys[8][115] ), 
        .QN(n1055) );
  DFFX1_HVT \keys_reg[8][114]  ( .D(n2623), .CLK(clk), .Q(\keys[8][114] ), 
        .QN(n1056) );
  DFFX1_HVT \keys_reg[8][113]  ( .D(n2622), .CLK(clk), .Q(\keys[8][113] ), 
        .QN(n1057) );
  DFFX1_HVT \keys_reg[8][112]  ( .D(n2621), .CLK(clk), .Q(\keys[8][112] ), 
        .QN(n1058) );
  DFFX1_HVT \keys_reg[8][111]  ( .D(n2620), .CLK(clk), .Q(\keys[8][111] ), 
        .QN(n1059) );
  DFFX1_HVT \keys_reg[8][110]  ( .D(n2619), .CLK(clk), .Q(\keys[8][110] ), 
        .QN(n1060) );
  DFFX1_HVT \keys_reg[8][109]  ( .D(n2618), .CLK(clk), .Q(\keys[8][109] ), 
        .QN(n1061) );
  DFFX1_HVT \keys_reg[8][108]  ( .D(n2617), .CLK(clk), .Q(\keys[8][108] ), 
        .QN(n1062) );
  DFFX1_HVT \keys_reg[8][107]  ( .D(n2616), .CLK(clk), .Q(\keys[8][107] ), 
        .QN(n1063) );
  DFFX1_HVT \keys_reg[8][106]  ( .D(n2615), .CLK(clk), .Q(\keys[8][106] ), 
        .QN(n1064) );
  DFFX1_HVT \keys_reg[8][105]  ( .D(n2614), .CLK(clk), .Q(\keys[8][105] ), 
        .QN(n1065) );
  DFFX1_HVT \keys_reg[8][104]  ( .D(n2613), .CLK(clk), .Q(\keys[8][104] ), 
        .QN(n1066) );
  DFFX1_HVT \keys_reg[8][103]  ( .D(n2612), .CLK(clk), .Q(\keys[8][103] ), 
        .QN(n1067) );
  DFFX1_HVT \keys_reg[8][102]  ( .D(n2611), .CLK(clk), .Q(\keys[8][102] ), 
        .QN(n1068) );
  DFFX1_HVT \keys_reg[8][101]  ( .D(n2610), .CLK(clk), .Q(\keys[8][101] ), 
        .QN(n1069) );
  DFFX1_HVT \keys_reg[8][100]  ( .D(n2609), .CLK(clk), .Q(\keys[8][100] ), 
        .QN(n1070) );
  DFFX1_HVT \keys_reg[8][99]  ( .D(n2608), .CLK(clk), .Q(\keys[8][99] ), .QN(
        n1071) );
  DFFX1_HVT \keys_reg[8][98]  ( .D(n2607), .CLK(clk), .Q(\keys[8][98] ), .QN(
        n1072) );
  DFFX1_HVT \keys_reg[8][97]  ( .D(n2606), .CLK(clk), .Q(\keys[8][97] ), .QN(
        n1073) );
  DFFX1_HVT \keys_reg[8][96]  ( .D(n2605), .CLK(clk), .Q(\keys[8][96] ), .QN(
        n1074) );
  DFFX1_HVT \keys_reg[8][95]  ( .D(n2604), .CLK(clk), .Q(\keys[8][95] ), .QN(
        n1075) );
  DFFX1_HVT \keys_reg[8][94]  ( .D(n2603), .CLK(clk), .Q(\keys[8][94] ), .QN(
        n1076) );
  DFFX1_HVT \keys_reg[8][93]  ( .D(n2602), .CLK(clk), .Q(\keys[8][93] ), .QN(
        n1077) );
  DFFX1_HVT \keys_reg[8][92]  ( .D(n2601), .CLK(clk), .Q(\keys[8][92] ), .QN(
        n1078) );
  DFFX1_HVT \keys_reg[8][91]  ( .D(n2600), .CLK(clk), .Q(\keys[8][91] ), .QN(
        n1079) );
  DFFX1_HVT \keys_reg[8][90]  ( .D(n2599), .CLK(clk), .Q(\keys[8][90] ), .QN(
        n1080) );
  DFFX1_HVT \keys_reg[8][89]  ( .D(n2598), .CLK(clk), .Q(\keys[8][89] ), .QN(
        n1081) );
  DFFX1_HVT \keys_reg[8][88]  ( .D(n2597), .CLK(clk), .Q(\keys[8][88] ), .QN(
        n1082) );
  DFFX1_HVT \keys_reg[8][87]  ( .D(n2596), .CLK(clk), .Q(\keys[8][87] ), .QN(
        n1083) );
  DFFX1_HVT \keys_reg[8][86]  ( .D(n2595), .CLK(clk), .Q(\keys[8][86] ), .QN(
        n1084) );
  DFFX1_HVT \keys_reg[8][85]  ( .D(n2594), .CLK(clk), .Q(\keys[8][85] ), .QN(
        n1085) );
  DFFX1_HVT \keys_reg[8][84]  ( .D(n2593), .CLK(clk), .Q(\keys[8][84] ), .QN(
        n1086) );
  DFFX1_HVT \keys_reg[8][83]  ( .D(n2592), .CLK(clk), .Q(\keys[8][83] ), .QN(
        n1087) );
  DFFX1_HVT \keys_reg[8][82]  ( .D(n2591), .CLK(clk), .Q(\keys[8][82] ), .QN(
        n1088) );
  DFFX1_HVT \keys_reg[8][81]  ( .D(n2590), .CLK(clk), .Q(\keys[8][81] ), .QN(
        n1089) );
  DFFX1_HVT \keys_reg[8][80]  ( .D(n2589), .CLK(clk), .Q(\keys[8][80] ), .QN(
        n1090) );
  DFFX1_HVT \keys_reg[8][79]  ( .D(n2588), .CLK(clk), .Q(\keys[8][79] ), .QN(
        n1091) );
  DFFX1_HVT \keys_reg[8][78]  ( .D(n2587), .CLK(clk), .Q(\keys[8][78] ), .QN(
        n1092) );
  DFFX1_HVT \keys_reg[8][77]  ( .D(n2586), .CLK(clk), .Q(\keys[8][77] ), .QN(
        n1093) );
  DFFX1_HVT \keys_reg[8][76]  ( .D(n2585), .CLK(clk), .Q(\keys[8][76] ), .QN(
        n1094) );
  DFFX1_HVT \keys_reg[8][75]  ( .D(n2584), .CLK(clk), .Q(\keys[8][75] ), .QN(
        n1095) );
  DFFX1_HVT \keys_reg[8][74]  ( .D(n2583), .CLK(clk), .Q(\keys[8][74] ), .QN(
        n1096) );
  DFFX1_HVT \keys_reg[8][73]  ( .D(n2582), .CLK(clk), .Q(\keys[8][73] ), .QN(
        n1097) );
  DFFX1_HVT \keys_reg[8][72]  ( .D(n2581), .CLK(clk), .Q(\keys[8][72] ), .QN(
        n1098) );
  DFFX1_HVT \keys_reg[8][71]  ( .D(n2580), .CLK(clk), .Q(\keys[8][71] ), .QN(
        n1099) );
  DFFX1_HVT \keys_reg[8][70]  ( .D(n2579), .CLK(clk), .Q(\keys[8][70] ), .QN(
        n1100) );
  DFFX1_HVT \keys_reg[8][69]  ( .D(n2578), .CLK(clk), .Q(\keys[8][69] ), .QN(
        n1101) );
  DFFX1_HVT \keys_reg[8][68]  ( .D(n2577), .CLK(clk), .Q(\keys[8][68] ), .QN(
        n1102) );
  DFFX1_HVT \keys_reg[8][67]  ( .D(n2576), .CLK(clk), .Q(\keys[8][67] ), .QN(
        n1103) );
  DFFX1_HVT \keys_reg[8][66]  ( .D(n2575), .CLK(clk), .Q(\keys[8][66] ), .QN(
        n1104) );
  DFFX1_HVT \keys_reg[8][65]  ( .D(n2574), .CLK(clk), .Q(\keys[8][65] ), .QN(
        n1105) );
  DFFX1_HVT \keys_reg[8][64]  ( .D(n2573), .CLK(clk), .Q(\keys[8][64] ), .QN(
        n1106) );
  DFFX1_HVT \keys_reg[8][63]  ( .D(n2572), .CLK(clk), .Q(\keys[8][63] ), .QN(
        n1107) );
  DFFX1_HVT \keys_reg[8][62]  ( .D(n2571), .CLK(clk), .Q(\keys[8][62] ), .QN(
        n1108) );
  DFFX1_HVT \keys_reg[8][61]  ( .D(n2570), .CLK(clk), .Q(\keys[8][61] ), .QN(
        n1109) );
  DFFX1_HVT \keys_reg[8][60]  ( .D(n2569), .CLK(clk), .Q(\keys[8][60] ), .QN(
        n1110) );
  DFFX1_HVT \keys_reg[8][59]  ( .D(n2568), .CLK(clk), .Q(\keys[8][59] ), .QN(
        n1111) );
  DFFX1_HVT \keys_reg[8][58]  ( .D(n2567), .CLK(clk), .Q(\keys[8][58] ), .QN(
        n1112) );
  DFFX1_HVT \keys_reg[8][57]  ( .D(n2566), .CLK(clk), .Q(\keys[8][57] ), .QN(
        n1113) );
  DFFX1_HVT \keys_reg[8][56]  ( .D(n2565), .CLK(clk), .Q(\keys[8][56] ), .QN(
        n1114) );
  DFFX1_HVT \keys_reg[8][55]  ( .D(n2564), .CLK(clk), .Q(\keys[8][55] ), .QN(
        n1115) );
  DFFX1_HVT \keys_reg[8][54]  ( .D(n2563), .CLK(clk), .Q(\keys[8][54] ), .QN(
        n1116) );
  DFFX1_HVT \keys_reg[8][53]  ( .D(n2562), .CLK(clk), .Q(\keys[8][53] ), .QN(
        n1117) );
  DFFX1_HVT \keys_reg[8][52]  ( .D(n2561), .CLK(clk), .Q(\keys[8][52] ), .QN(
        n1118) );
  DFFX1_HVT \keys_reg[8][51]  ( .D(n2560), .CLK(clk), .Q(\keys[8][51] ), .QN(
        n1119) );
  DFFX1_HVT \keys_reg[8][50]  ( .D(n2559), .CLK(clk), .Q(\keys[8][50] ), .QN(
        n1120) );
  DFFX1_HVT \keys_reg[8][49]  ( .D(n2558), .CLK(clk), .Q(\keys[8][49] ), .QN(
        n1121) );
  DFFX1_HVT \keys_reg[8][48]  ( .D(n2557), .CLK(clk), .Q(\keys[8][48] ), .QN(
        n1122) );
  DFFX1_HVT \keys_reg[8][47]  ( .D(n2556), .CLK(clk), .Q(\keys[8][47] ), .QN(
        n1123) );
  DFFX1_HVT \keys_reg[8][46]  ( .D(n2555), .CLK(clk), .Q(\keys[8][46] ), .QN(
        n1124) );
  DFFX1_HVT \keys_reg[8][45]  ( .D(n2554), .CLK(clk), .Q(\keys[8][45] ), .QN(
        n1125) );
  DFFX1_HVT \keys_reg[8][44]  ( .D(n2553), .CLK(clk), .Q(\keys[8][44] ), .QN(
        n1126) );
  DFFX1_HVT \keys_reg[8][43]  ( .D(n2552), .CLK(clk), .Q(\keys[8][43] ), .QN(
        n1127) );
  DFFX1_HVT \keys_reg[8][42]  ( .D(n2551), .CLK(clk), .Q(\keys[8][42] ), .QN(
        n1128) );
  DFFX1_HVT \keys_reg[8][41]  ( .D(n2550), .CLK(clk), .Q(\keys[8][41] ), .QN(
        n1129) );
  DFFX1_HVT \keys_reg[8][40]  ( .D(n2549), .CLK(clk), .Q(\keys[8][40] ), .QN(
        n1130) );
  DFFX1_HVT \keys_reg[8][39]  ( .D(n2548), .CLK(clk), .Q(\keys[8][39] ), .QN(
        n1131) );
  DFFX1_HVT \keys_reg[8][38]  ( .D(n2547), .CLK(clk), .Q(\keys[8][38] ), .QN(
        n1132) );
  DFFX1_HVT \keys_reg[8][37]  ( .D(n2546), .CLK(clk), .Q(\keys[8][37] ), .QN(
        n1133) );
  DFFX1_HVT \keys_reg[8][36]  ( .D(n2545), .CLK(clk), .Q(\keys[8][36] ), .QN(
        n1134) );
  DFFX1_HVT \keys_reg[8][35]  ( .D(n2544), .CLK(clk), .Q(\keys[8][35] ), .QN(
        n1135) );
  DFFX1_HVT \keys_reg[8][34]  ( .D(n2543), .CLK(clk), .Q(\keys[8][34] ), .QN(
        n1136) );
  DFFX1_HVT \keys_reg[8][33]  ( .D(n2542), .CLK(clk), .Q(\keys[8][33] ), .QN(
        n1137) );
  DFFX1_HVT \keys_reg[8][32]  ( .D(n2541), .CLK(clk), .Q(\keys[8][32] ), .QN(
        n1138) );
  DFFX1_HVT \keys_reg[8][31]  ( .D(n2540), .CLK(clk), .Q(\keys[8][31] ), .QN(
        n1139) );
  DFFX1_HVT \keys_reg[8][30]  ( .D(n2539), .CLK(clk), .Q(\keys[8][30] ), .QN(
        n1140) );
  DFFX1_HVT \keys_reg[8][29]  ( .D(n2538), .CLK(clk), .Q(\keys[8][29] ), .QN(
        n1141) );
  DFFX1_HVT \keys_reg[8][28]  ( .D(n2537), .CLK(clk), .Q(\keys[8][28] ), .QN(
        n1142) );
  DFFX1_HVT \keys_reg[8][27]  ( .D(n2536), .CLK(clk), .Q(\keys[8][27] ), .QN(
        n1143) );
  DFFX1_HVT \keys_reg[8][26]  ( .D(n2535), .CLK(clk), .Q(\keys[8][26] ), .QN(
        n1144) );
  DFFX1_HVT \keys_reg[8][25]  ( .D(n2534), .CLK(clk), .Q(\keys[8][25] ), .QN(
        n1145) );
  DFFX1_HVT \keys_reg[8][24]  ( .D(n2533), .CLK(clk), .Q(\keys[8][24] ), .QN(
        n1146) );
  DFFX1_HVT \keys_reg[8][23]  ( .D(n2532), .CLK(clk), .Q(\keys[8][23] ), .QN(
        n1147) );
  DFFX1_HVT \keys_reg[8][22]  ( .D(n2531), .CLK(clk), .Q(\keys[8][22] ), .QN(
        n1148) );
  DFFX1_HVT \keys_reg[8][21]  ( .D(n2530), .CLK(clk), .Q(\keys[8][21] ), .QN(
        n1149) );
  DFFX1_HVT \keys_reg[8][20]  ( .D(n2529), .CLK(clk), .Q(\keys[8][20] ), .QN(
        n1150) );
  DFFX1_HVT \keys_reg[8][19]  ( .D(n2528), .CLK(clk), .Q(\keys[8][19] ), .QN(
        n1151) );
  DFFX1_HVT \keys_reg[8][18]  ( .D(n2527), .CLK(clk), .Q(\keys[8][18] ), .QN(
        n1152) );
  DFFX1_HVT \keys_reg[8][17]  ( .D(n2526), .CLK(clk), .Q(\keys[8][17] ), .QN(
        n1153) );
  DFFX1_HVT \keys_reg[8][16]  ( .D(n2525), .CLK(clk), .Q(\keys[8][16] ), .QN(
        n1154) );
  DFFX1_HVT \keys_reg[8][15]  ( .D(n2524), .CLK(clk), .Q(\keys[8][15] ), .QN(
        n1155) );
  DFFX1_HVT \keys_reg[8][14]  ( .D(n2523), .CLK(clk), .Q(\keys[8][14] ), .QN(
        n1156) );
  DFFX1_HVT \keys_reg[8][13]  ( .D(n2522), .CLK(clk), .Q(\keys[8][13] ), .QN(
        n1157) );
  DFFX1_HVT \keys_reg[8][12]  ( .D(n2521), .CLK(clk), .Q(\keys[8][12] ), .QN(
        n1158) );
  DFFX1_HVT \keys_reg[8][11]  ( .D(n2520), .CLK(clk), .Q(\keys[8][11] ), .QN(
        n1159) );
  DFFX1_HVT \keys_reg[8][10]  ( .D(n2519), .CLK(clk), .Q(\keys[8][10] ), .QN(
        n1160) );
  DFFX1_HVT \keys_reg[8][9]  ( .D(n2518), .CLK(clk), .Q(\keys[8][9] ), .QN(
        n1161) );
  DFFX1_HVT \keys_reg[8][8]  ( .D(n2517), .CLK(clk), .Q(\keys[8][8] ), .QN(
        n1162) );
  DFFX1_HVT \keys_reg[8][7]  ( .D(n2516), .CLK(clk), .Q(\keys[8][7] ), .QN(
        n1163) );
  DFFX1_HVT \keys_reg[8][6]  ( .D(n2515), .CLK(clk), .Q(\keys[8][6] ), .QN(
        n1164) );
  DFFX1_HVT \keys_reg[8][5]  ( .D(n2514), .CLK(clk), .Q(\keys[8][5] ), .QN(
        n1165) );
  DFFX1_HVT \keys_reg[8][4]  ( .D(n2513), .CLK(clk), .Q(\keys[8][4] ), .QN(
        n1166) );
  DFFX1_HVT \keys_reg[8][3]  ( .D(n2512), .CLK(clk), .Q(\keys[8][3] ), .QN(
        n1167) );
  DFFX1_HVT \keys_reg[8][2]  ( .D(n2511), .CLK(clk), .Q(\keys[8][2] ), .QN(
        n1168) );
  DFFX1_HVT \keys_reg[8][1]  ( .D(n2510), .CLK(clk), .Q(\keys[8][1] ), .QN(
        n1169) );
  DFFX1_HVT \keys_reg[8][0]  ( .D(n2509), .CLK(clk), .Q(\keys[8][0] ), .QN(
        n1170) );
  DFFX1_HVT \keys_reg[9][127]  ( .D(n2508), .CLK(clk), .Q(\keys[9][127] ), 
        .QN(n1171) );
  DFFX1_HVT \keys_reg[9][126]  ( .D(n2507), .CLK(clk), .Q(\keys[9][126] ), 
        .QN(n1172) );
  DFFX1_HVT \keys_reg[9][125]  ( .D(n2506), .CLK(clk), .Q(\keys[9][125] ), 
        .QN(n1173) );
  DFFX1_HVT \keys_reg[9][124]  ( .D(n2505), .CLK(clk), .Q(\keys[9][124] ), 
        .QN(n1174) );
  DFFX1_HVT \keys_reg[9][123]  ( .D(n2504), .CLK(clk), .Q(\keys[9][123] ), 
        .QN(n1175) );
  DFFX1_HVT \keys_reg[9][122]  ( .D(n2503), .CLK(clk), .Q(\keys[9][122] ), 
        .QN(n1176) );
  DFFX1_HVT \keys_reg[9][121]  ( .D(n2502), .CLK(clk), .Q(\keys[9][121] ), 
        .QN(n1177) );
  DFFX1_HVT \keys_reg[9][120]  ( .D(n2501), .CLK(clk), .Q(\keys[9][120] ), 
        .QN(n1178) );
  DFFX1_HVT \keys_reg[9][119]  ( .D(n2500), .CLK(clk), .Q(\keys[9][119] ), 
        .QN(n1179) );
  DFFX1_HVT \keys_reg[9][118]  ( .D(n2499), .CLK(clk), .Q(\keys[9][118] ), 
        .QN(n1180) );
  DFFX1_HVT \keys_reg[9][117]  ( .D(n2498), .CLK(clk), .Q(\keys[9][117] ), 
        .QN(n1181) );
  DFFX1_HVT \keys_reg[9][116]  ( .D(n2497), .CLK(clk), .Q(\keys[9][116] ), 
        .QN(n1182) );
  DFFX1_HVT \keys_reg[9][115]  ( .D(n2496), .CLK(clk), .Q(\keys[9][115] ), 
        .QN(n1183) );
  DFFX1_HVT \keys_reg[9][114]  ( .D(n2495), .CLK(clk), .Q(\keys[9][114] ), 
        .QN(n1184) );
  DFFX1_HVT \keys_reg[9][113]  ( .D(n2494), .CLK(clk), .Q(\keys[9][113] ), 
        .QN(n1185) );
  DFFX1_HVT \keys_reg[9][112]  ( .D(n2493), .CLK(clk), .Q(\keys[9][112] ), 
        .QN(n1186) );
  DFFX1_HVT \keys_reg[9][111]  ( .D(n2492), .CLK(clk), .Q(\keys[9][111] ), 
        .QN(n1187) );
  DFFX1_HVT \keys_reg[9][110]  ( .D(n2491), .CLK(clk), .Q(\keys[9][110] ), 
        .QN(n1188) );
  DFFX1_HVT \keys_reg[9][109]  ( .D(n2490), .CLK(clk), .Q(\keys[9][109] ), 
        .QN(n1189) );
  DFFX1_HVT \keys_reg[9][108]  ( .D(n2489), .CLK(clk), .Q(\keys[9][108] ), 
        .QN(n1190) );
  DFFX1_HVT \keys_reg[9][107]  ( .D(n2488), .CLK(clk), .Q(\keys[9][107] ), 
        .QN(n1191) );
  DFFX1_HVT \keys_reg[9][106]  ( .D(n2487), .CLK(clk), .Q(\keys[9][106] ), 
        .QN(n1192) );
  DFFX1_HVT \keys_reg[9][105]  ( .D(n2486), .CLK(clk), .Q(\keys[9][105] ), 
        .QN(n1193) );
  DFFX1_HVT \keys_reg[9][104]  ( .D(n2485), .CLK(clk), .Q(\keys[9][104] ), 
        .QN(n1194) );
  DFFX1_HVT \keys_reg[9][103]  ( .D(n2484), .CLK(clk), .Q(\keys[9][103] ), 
        .QN(n1195) );
  DFFX1_HVT \keys_reg[9][102]  ( .D(n2483), .CLK(clk), .Q(\keys[9][102] ), 
        .QN(n1196) );
  DFFX1_HVT \keys_reg[9][101]  ( .D(n2482), .CLK(clk), .Q(\keys[9][101] ), 
        .QN(n1197) );
  DFFX1_HVT \keys_reg[9][100]  ( .D(n2481), .CLK(clk), .Q(\keys[9][100] ), 
        .QN(n1198) );
  DFFX1_HVT \keys_reg[9][99]  ( .D(n2480), .CLK(clk), .Q(\keys[9][99] ), .QN(
        n1199) );
  DFFX1_HVT \keys_reg[9][98]  ( .D(n2479), .CLK(clk), .Q(\keys[9][98] ), .QN(
        n1200) );
  DFFX1_HVT \keys_reg[9][97]  ( .D(n2478), .CLK(clk), .Q(\keys[9][97] ), .QN(
        n1201) );
  DFFX1_HVT \keys_reg[9][96]  ( .D(n2477), .CLK(clk), .Q(\keys[9][96] ), .QN(
        n1202) );
  DFFX1_HVT \keys_reg[9][95]  ( .D(n2476), .CLK(clk), .Q(\keys[9][95] ), .QN(
        n1203) );
  DFFX1_HVT \keys_reg[9][94]  ( .D(n2475), .CLK(clk), .Q(\keys[9][94] ), .QN(
        n1204) );
  DFFX1_HVT \keys_reg[9][93]  ( .D(n2474), .CLK(clk), .Q(\keys[9][93] ), .QN(
        n1205) );
  DFFX1_HVT \keys_reg[9][92]  ( .D(n2473), .CLK(clk), .Q(\keys[9][92] ), .QN(
        n1206) );
  DFFX1_HVT \keys_reg[9][91]  ( .D(n2472), .CLK(clk), .Q(\keys[9][91] ), .QN(
        n1207) );
  DFFX1_HVT \keys_reg[9][90]  ( .D(n2471), .CLK(clk), .Q(\keys[9][90] ), .QN(
        n1208) );
  DFFX1_HVT \keys_reg[9][89]  ( .D(n2470), .CLK(clk), .Q(\keys[9][89] ), .QN(
        n1209) );
  DFFX1_HVT \keys_reg[9][88]  ( .D(n2469), .CLK(clk), .Q(\keys[9][88] ), .QN(
        n1210) );
  DFFX1_HVT \keys_reg[9][87]  ( .D(n2468), .CLK(clk), .Q(\keys[9][87] ), .QN(
        n1211) );
  DFFX1_HVT \keys_reg[9][86]  ( .D(n2467), .CLK(clk), .Q(\keys[9][86] ), .QN(
        n1212) );
  DFFX1_HVT \keys_reg[9][85]  ( .D(n2466), .CLK(clk), .Q(\keys[9][85] ), .QN(
        n1213) );
  DFFX1_HVT \keys_reg[9][84]  ( .D(n2465), .CLK(clk), .Q(\keys[9][84] ), .QN(
        n1214) );
  DFFX1_HVT \keys_reg[9][83]  ( .D(n2464), .CLK(clk), .Q(\keys[9][83] ), .QN(
        n1215) );
  DFFX1_HVT \keys_reg[9][82]  ( .D(n2463), .CLK(clk), .Q(\keys[9][82] ), .QN(
        n1216) );
  DFFX1_HVT \keys_reg[9][81]  ( .D(n2462), .CLK(clk), .Q(\keys[9][81] ), .QN(
        n1217) );
  DFFX1_HVT \keys_reg[9][80]  ( .D(n2461), .CLK(clk), .Q(\keys[9][80] ), .QN(
        n1218) );
  DFFX1_HVT \keys_reg[9][79]  ( .D(n2460), .CLK(clk), .Q(\keys[9][79] ), .QN(
        n1219) );
  DFFX1_HVT \keys_reg[9][78]  ( .D(n2459), .CLK(clk), .Q(\keys[9][78] ), .QN(
        n1220) );
  DFFX1_HVT \keys_reg[9][77]  ( .D(n2458), .CLK(clk), .Q(\keys[9][77] ), .QN(
        n1221) );
  DFFX1_HVT \keys_reg[9][76]  ( .D(n2457), .CLK(clk), .Q(\keys[9][76] ), .QN(
        n1222) );
  DFFX1_HVT \keys_reg[9][75]  ( .D(n2456), .CLK(clk), .Q(\keys[9][75] ), .QN(
        n1223) );
  DFFX1_HVT \keys_reg[9][74]  ( .D(n2455), .CLK(clk), .Q(\keys[9][74] ), .QN(
        n1224) );
  DFFX1_HVT \keys_reg[9][73]  ( .D(n2454), .CLK(clk), .Q(\keys[9][73] ), .QN(
        n1225) );
  DFFX1_HVT \keys_reg[9][72]  ( .D(n2453), .CLK(clk), .Q(\keys[9][72] ), .QN(
        n1226) );
  DFFX1_HVT \keys_reg[9][71]  ( .D(n2452), .CLK(clk), .Q(\keys[9][71] ), .QN(
        n1227) );
  DFFX1_HVT \keys_reg[9][70]  ( .D(n2451), .CLK(clk), .Q(\keys[9][70] ), .QN(
        n1228) );
  DFFX1_HVT \keys_reg[9][69]  ( .D(n2450), .CLK(clk), .Q(\keys[9][69] ), .QN(
        n1229) );
  DFFX1_HVT \keys_reg[9][68]  ( .D(n2449), .CLK(clk), .Q(\keys[9][68] ), .QN(
        n1230) );
  DFFX1_HVT \keys_reg[9][67]  ( .D(n2448), .CLK(clk), .Q(\keys[9][67] ), .QN(
        n1231) );
  DFFX1_HVT \keys_reg[9][66]  ( .D(n2447), .CLK(clk), .Q(\keys[9][66] ), .QN(
        n1232) );
  DFFX1_HVT \keys_reg[9][65]  ( .D(n2446), .CLK(clk), .Q(\keys[9][65] ), .QN(
        n1233) );
  DFFX1_HVT \keys_reg[9][64]  ( .D(n2445), .CLK(clk), .Q(\keys[9][64] ), .QN(
        n1234) );
  DFFX1_HVT \keys_reg[9][63]  ( .D(n2444), .CLK(clk), .Q(\keys[9][63] ), .QN(
        n1235) );
  DFFX1_HVT \keys_reg[9][62]  ( .D(n2443), .CLK(clk), .Q(\keys[9][62] ), .QN(
        n1236) );
  DFFX1_HVT \keys_reg[9][61]  ( .D(n2442), .CLK(clk), .Q(\keys[9][61] ), .QN(
        n1237) );
  DFFX1_HVT \keys_reg[9][60]  ( .D(n2441), .CLK(clk), .Q(\keys[9][60] ), .QN(
        n1238) );
  DFFX1_HVT \keys_reg[9][59]  ( .D(n2440), .CLK(clk), .Q(\keys[9][59] ), .QN(
        n1239) );
  DFFX1_HVT \keys_reg[9][58]  ( .D(n2439), .CLK(clk), .Q(\keys[9][58] ), .QN(
        n1240) );
  DFFX1_HVT \keys_reg[9][57]  ( .D(n2438), .CLK(clk), .Q(\keys[9][57] ), .QN(
        n1241) );
  DFFX1_HVT \keys_reg[9][56]  ( .D(n2437), .CLK(clk), .Q(\keys[9][56] ), .QN(
        n1242) );
  DFFX1_HVT \keys_reg[9][55]  ( .D(n2436), .CLK(clk), .Q(\keys[9][55] ), .QN(
        n1243) );
  DFFX1_HVT \keys_reg[9][54]  ( .D(n2435), .CLK(clk), .Q(\keys[9][54] ), .QN(
        n1244) );
  DFFX1_HVT \keys_reg[9][53]  ( .D(n2434), .CLK(clk), .Q(\keys[9][53] ), .QN(
        n1245) );
  DFFX1_HVT \keys_reg[9][52]  ( .D(n2433), .CLK(clk), .Q(\keys[9][52] ), .QN(
        n1246) );
  DFFX1_HVT \keys_reg[9][51]  ( .D(n2432), .CLK(clk), .Q(\keys[9][51] ), .QN(
        n1247) );
  DFFX1_HVT \keys_reg[9][50]  ( .D(n2431), .CLK(clk), .Q(\keys[9][50] ), .QN(
        n1248) );
  DFFX1_HVT \keys_reg[9][49]  ( .D(n2430), .CLK(clk), .Q(\keys[9][49] ), .QN(
        n1249) );
  DFFX1_HVT \keys_reg[9][48]  ( .D(n2429), .CLK(clk), .Q(\keys[9][48] ), .QN(
        n1250) );
  DFFX1_HVT \keys_reg[9][47]  ( .D(n2428), .CLK(clk), .Q(\keys[9][47] ), .QN(
        n1251) );
  DFFX1_HVT \keys_reg[9][46]  ( .D(n2427), .CLK(clk), .Q(\keys[9][46] ), .QN(
        n1252) );
  DFFX1_HVT \keys_reg[9][45]  ( .D(n2426), .CLK(clk), .Q(\keys[9][45] ), .QN(
        n1253) );
  DFFX1_HVT \keys_reg[9][44]  ( .D(n2425), .CLK(clk), .Q(\keys[9][44] ), .QN(
        n1254) );
  DFFX1_HVT \keys_reg[9][43]  ( .D(n2424), .CLK(clk), .Q(\keys[9][43] ), .QN(
        n1255) );
  DFFX1_HVT \keys_reg[9][42]  ( .D(n2423), .CLK(clk), .Q(\keys[9][42] ), .QN(
        n1256) );
  DFFX1_HVT \keys_reg[9][41]  ( .D(n2422), .CLK(clk), .Q(\keys[9][41] ), .QN(
        n1257) );
  DFFX1_HVT \keys_reg[9][40]  ( .D(n2421), .CLK(clk), .Q(\keys[9][40] ), .QN(
        n1258) );
  DFFX1_HVT \keys_reg[9][39]  ( .D(n2420), .CLK(clk), .Q(\keys[9][39] ), .QN(
        n1259) );
  DFFX1_HVT \keys_reg[9][38]  ( .D(n2419), .CLK(clk), .Q(\keys[9][38] ), .QN(
        n1260) );
  DFFX1_HVT \keys_reg[9][37]  ( .D(n2418), .CLK(clk), .Q(\keys[9][37] ), .QN(
        n1261) );
  DFFX1_HVT \keys_reg[9][36]  ( .D(n2417), .CLK(clk), .Q(\keys[9][36] ), .QN(
        n1262) );
  DFFX1_HVT \keys_reg[9][35]  ( .D(n2416), .CLK(clk), .Q(\keys[9][35] ), .QN(
        n1263) );
  DFFX1_HVT \keys_reg[9][34]  ( .D(n2415), .CLK(clk), .Q(\keys[9][34] ), .QN(
        n1264) );
  DFFX1_HVT \keys_reg[9][33]  ( .D(n2414), .CLK(clk), .Q(\keys[9][33] ), .QN(
        n1265) );
  DFFX1_HVT \keys_reg[9][32]  ( .D(n2413), .CLK(clk), .Q(\keys[9][32] ), .QN(
        n1266) );
  DFFX1_HVT \keys_reg[9][31]  ( .D(n2412), .CLK(clk), .Q(\keys[9][31] ), .QN(
        n1267) );
  DFFX1_HVT \keys_reg[9][30]  ( .D(n2411), .CLK(clk), .Q(\keys[9][30] ), .QN(
        n1268) );
  DFFX1_HVT \keys_reg[9][29]  ( .D(n2410), .CLK(clk), .Q(\keys[9][29] ), .QN(
        n1269) );
  DFFX1_HVT \keys_reg[9][28]  ( .D(n2409), .CLK(clk), .Q(\keys[9][28] ), .QN(
        n1270) );
  DFFX1_HVT \keys_reg[9][27]  ( .D(n2408), .CLK(clk), .Q(\keys[9][27] ), .QN(
        n1271) );
  DFFX1_HVT \keys_reg[9][26]  ( .D(n2407), .CLK(clk), .Q(\keys[9][26] ), .QN(
        n1272) );
  DFFX1_HVT \keys_reg[9][25]  ( .D(n2406), .CLK(clk), .Q(\keys[9][25] ), .QN(
        n1273) );
  DFFX1_HVT \keys_reg[9][24]  ( .D(n2405), .CLK(clk), .Q(\keys[9][24] ), .QN(
        n1274) );
  DFFX1_HVT \keys_reg[9][23]  ( .D(n2404), .CLK(clk), .Q(\keys[9][23] ), .QN(
        n1275) );
  DFFX1_HVT \keys_reg[9][22]  ( .D(n2403), .CLK(clk), .Q(\keys[9][22] ), .QN(
        n1276) );
  DFFX1_HVT \keys_reg[9][21]  ( .D(n2402), .CLK(clk), .Q(\keys[9][21] ), .QN(
        n1277) );
  DFFX1_HVT \keys_reg[9][20]  ( .D(n2401), .CLK(clk), .Q(\keys[9][20] ), .QN(
        n1278) );
  DFFX1_HVT \keys_reg[9][19]  ( .D(n2400), .CLK(clk), .Q(\keys[9][19] ), .QN(
        n1279) );
  DFFX1_HVT \keys_reg[9][18]  ( .D(n2399), .CLK(clk), .Q(\keys[9][18] ), .QN(
        n1280) );
  DFFX1_HVT \keys_reg[9][17]  ( .D(n2398), .CLK(clk), .Q(\keys[9][17] ), .QN(
        n1281) );
  DFFX1_HVT \keys_reg[9][16]  ( .D(n2397), .CLK(clk), .Q(\keys[9][16] ), .QN(
        n1282) );
  DFFX1_HVT \keys_reg[9][15]  ( .D(n2396), .CLK(clk), .Q(\keys[9][15] ), .QN(
        n1283) );
  DFFX1_HVT \keys_reg[9][14]  ( .D(n2395), .CLK(clk), .Q(\keys[9][14] ), .QN(
        n1284) );
  DFFX1_HVT \keys_reg[9][13]  ( .D(n2394), .CLK(clk), .Q(\keys[9][13] ), .QN(
        n1285) );
  DFFX1_HVT \keys_reg[9][12]  ( .D(n2393), .CLK(clk), .Q(\keys[9][12] ), .QN(
        n1286) );
  DFFX1_HVT \keys_reg[9][11]  ( .D(n2392), .CLK(clk), .Q(\keys[9][11] ), .QN(
        n1287) );
  DFFX1_HVT \keys_reg[9][10]  ( .D(n2391), .CLK(clk), .Q(\keys[9][10] ), .QN(
        n1288) );
  DFFX1_HVT \keys_reg[9][9]  ( .D(n2390), .CLK(clk), .Q(\keys[9][9] ), .QN(
        n1289) );
  DFFX1_HVT \keys_reg[9][8]  ( .D(n2389), .CLK(clk), .Q(\keys[9][8] ), .QN(
        n1290) );
  DFFX1_HVT \keys_reg[9][7]  ( .D(n2388), .CLK(clk), .Q(\keys[9][7] ), .QN(
        n1291) );
  DFFX1_HVT \keys_reg[9][6]  ( .D(n2387), .CLK(clk), .Q(\keys[9][6] ), .QN(
        n1292) );
  DFFX1_HVT \keys_reg[9][5]  ( .D(n2386), .CLK(clk), .Q(\keys[9][5] ), .QN(
        n1293) );
  DFFX1_HVT \keys_reg[9][4]  ( .D(n2385), .CLK(clk), .Q(\keys[9][4] ), .QN(
        n1294) );
  DFFX1_HVT \keys_reg[9][3]  ( .D(n2384), .CLK(clk), .Q(\keys[9][3] ), .QN(
        n1295) );
  DFFX1_HVT \keys_reg[9][2]  ( .D(n2383), .CLK(clk), .Q(\keys[9][2] ), .QN(
        n1296) );
  DFFX1_HVT \keys_reg[9][1]  ( .D(n2382), .CLK(clk), .Q(\keys[9][1] ), .QN(
        n1297) );
  DFFX1_HVT \keys_reg[9][0]  ( .D(n2381), .CLK(clk), .Q(\keys[9][0] ), .QN(
        n1298) );
  DFFX1_HVT \keys_reg[10][127]  ( .D(n2380), .CLK(clk), .Q(\keys[10][127] ), 
        .QN(n1299) );
  DFFX1_HVT \keys_reg[10][126]  ( .D(n2379), .CLK(clk), .Q(\keys[10][126] ), 
        .QN(n1300) );
  DFFX1_HVT \keys_reg[10][125]  ( .D(n2378), .CLK(clk), .Q(\keys[10][125] ), 
        .QN(n1301) );
  DFFX1_HVT \keys_reg[10][124]  ( .D(n2377), .CLK(clk), .Q(\keys[10][124] ), 
        .QN(n1302) );
  DFFX1_HVT \keys_reg[10][123]  ( .D(n2376), .CLK(clk), .Q(\keys[10][123] ), 
        .QN(n1303) );
  DFFX1_HVT \keys_reg[10][122]  ( .D(n2375), .CLK(clk), .Q(\keys[10][122] ), 
        .QN(n1304) );
  DFFX1_HVT \keys_reg[10][121]  ( .D(n2374), .CLK(clk), .Q(\keys[10][121] ), 
        .QN(n1305) );
  DFFX1_HVT \keys_reg[10][120]  ( .D(n2373), .CLK(clk), .Q(\keys[10][120] ), 
        .QN(n1306) );
  DFFX1_HVT \keys_reg[10][119]  ( .D(n2372), .CLK(clk), .Q(\keys[10][119] ), 
        .QN(n1307) );
  DFFX1_HVT \keys_reg[10][118]  ( .D(n2371), .CLK(clk), .Q(\keys[10][118] ), 
        .QN(n1308) );
  DFFX1_HVT \keys_reg[10][117]  ( .D(n2370), .CLK(clk), .Q(\keys[10][117] ), 
        .QN(n1309) );
  DFFX1_HVT \keys_reg[10][116]  ( .D(n2369), .CLK(clk), .Q(\keys[10][116] ), 
        .QN(n1310) );
  DFFX1_HVT \keys_reg[10][115]  ( .D(n2368), .CLK(clk), .Q(\keys[10][115] ), 
        .QN(n1311) );
  DFFX1_HVT \keys_reg[10][114]  ( .D(n2367), .CLK(clk), .Q(\keys[10][114] ), 
        .QN(n1312) );
  DFFX1_HVT \keys_reg[10][113]  ( .D(n2366), .CLK(clk), .Q(\keys[10][113] ), 
        .QN(n1313) );
  DFFX1_HVT \keys_reg[10][112]  ( .D(n2365), .CLK(clk), .Q(\keys[10][112] ), 
        .QN(n1314) );
  DFFX1_HVT \keys_reg[10][111]  ( .D(n2364), .CLK(clk), .Q(\keys[10][111] ), 
        .QN(n1315) );
  DFFX1_HVT \keys_reg[10][110]  ( .D(n2363), .CLK(clk), .Q(\keys[10][110] ), 
        .QN(n1316) );
  DFFX1_HVT \keys_reg[10][109]  ( .D(n2362), .CLK(clk), .Q(\keys[10][109] ), 
        .QN(n1317) );
  DFFX1_HVT \keys_reg[10][108]  ( .D(n2361), .CLK(clk), .Q(\keys[10][108] ), 
        .QN(n1318) );
  DFFX1_HVT \keys_reg[10][107]  ( .D(n2360), .CLK(clk), .Q(\keys[10][107] ), 
        .QN(n1319) );
  DFFX1_HVT \keys_reg[10][106]  ( .D(n2359), .CLK(clk), .Q(\keys[10][106] ), 
        .QN(n1320) );
  DFFX1_HVT \keys_reg[10][105]  ( .D(n2358), .CLK(clk), .Q(\keys[10][105] ), 
        .QN(n1321) );
  DFFX1_HVT \keys_reg[10][104]  ( .D(n2357), .CLK(clk), .Q(\keys[10][104] ), 
        .QN(n1322) );
  DFFX1_HVT \keys_reg[10][103]  ( .D(n2356), .CLK(clk), .Q(\keys[10][103] ), 
        .QN(n1323) );
  DFFX1_HVT \keys_reg[10][102]  ( .D(n2355), .CLK(clk), .Q(\keys[10][102] ), 
        .QN(n1324) );
  DFFX1_HVT \keys_reg[10][101]  ( .D(n2354), .CLK(clk), .Q(\keys[10][101] ), 
        .QN(n1325) );
  DFFX1_HVT \keys_reg[10][100]  ( .D(n2353), .CLK(clk), .Q(\keys[10][100] ), 
        .QN(n1326) );
  DFFX1_HVT \keys_reg[10][99]  ( .D(n2352), .CLK(clk), .Q(\keys[10][99] ), 
        .QN(n1327) );
  DFFX1_HVT \keys_reg[10][98]  ( .D(n2351), .CLK(clk), .Q(\keys[10][98] ), 
        .QN(n1328) );
  DFFX1_HVT \keys_reg[10][97]  ( .D(n2350), .CLK(clk), .Q(\keys[10][97] ), 
        .QN(n1329) );
  DFFX1_HVT \keys_reg[10][96]  ( .D(n2349), .CLK(clk), .Q(\keys[10][96] ), 
        .QN(n1330) );
  DFFX1_HVT \keys_reg[10][95]  ( .D(n2348), .CLK(clk), .Q(\keys[10][95] ), 
        .QN(n1331) );
  DFFX1_HVT \keys_reg[10][94]  ( .D(n2347), .CLK(clk), .Q(\keys[10][94] ), 
        .QN(n1332) );
  DFFX1_HVT \keys_reg[10][93]  ( .D(n2346), .CLK(clk), .Q(\keys[10][93] ), 
        .QN(n1333) );
  DFFX1_HVT \keys_reg[10][92]  ( .D(n2345), .CLK(clk), .Q(\keys[10][92] ), 
        .QN(n1334) );
  DFFX1_HVT \keys_reg[10][91]  ( .D(n2344), .CLK(clk), .Q(\keys[10][91] ), 
        .QN(n1335) );
  DFFX1_HVT \keys_reg[10][90]  ( .D(n2343), .CLK(clk), .QN(n1336) );
  DFFX1_HVT \keys_reg[10][89]  ( .D(n2342), .CLK(clk), .Q(\keys[10][89] ), 
        .QN(n1337) );
  DFFX1_HVT \keys_reg[10][88]  ( .D(n2341), .CLK(clk), .Q(\keys[10][88] ), 
        .QN(n1338) );
  DFFX1_HVT \keys_reg[10][87]  ( .D(n2340), .CLK(clk), .Q(\keys[10][87] ), 
        .QN(n1339) );
  DFFX1_HVT \keys_reg[10][86]  ( .D(n2339), .CLK(clk), .Q(\keys[10][86] ), 
        .QN(n1340) );
  DFFX1_HVT \keys_reg[10][85]  ( .D(n2338), .CLK(clk), .Q(\keys[10][85] ), 
        .QN(n1341) );
  DFFX1_HVT \keys_reg[10][84]  ( .D(n2337), .CLK(clk), .Q(\keys[10][84] ), 
        .QN(n1342) );
  DFFX1_HVT \keys_reg[10][83]  ( .D(n2336), .CLK(clk), .Q(\keys[10][83] ), 
        .QN(n1343) );
  DFFX1_HVT \keys_reg[10][82]  ( .D(n2335), .CLK(clk), .Q(\keys[10][82] ), 
        .QN(n1344) );
  DFFX1_HVT \keys_reg[10][81]  ( .D(n2334), .CLK(clk), .Q(\keys[10][81] ), 
        .QN(n1345) );
  DFFX1_HVT \keys_reg[10][80]  ( .D(n2333), .CLK(clk), .Q(\keys[10][80] ), 
        .QN(n1346) );
  DFFX1_HVT \keys_reg[10][79]  ( .D(n2332), .CLK(clk), .Q(\keys[10][79] ), 
        .QN(n1347) );
  DFFX1_HVT \keys_reg[10][78]  ( .D(n2331), .CLK(clk), .Q(\keys[10][78] ), 
        .QN(n1348) );
  DFFX1_HVT \keys_reg[10][77]  ( .D(n2330), .CLK(clk), .Q(\keys[10][77] ), 
        .QN(n1349) );
  DFFX1_HVT \keys_reg[10][76]  ( .D(n2329), .CLK(clk), .Q(\keys[10][76] ), 
        .QN(n1350) );
  DFFX1_HVT \keys_reg[10][75]  ( .D(n2328), .CLK(clk), .Q(\keys[10][75] ), 
        .QN(n1351) );
  DFFX1_HVT \keys_reg[10][74]  ( .D(n2327), .CLK(clk), .Q(\keys[10][74] ), 
        .QN(n1352) );
  DFFX1_HVT \keys_reg[10][73]  ( .D(n2326), .CLK(clk), .Q(\keys[10][73] ), 
        .QN(n1353) );
  DFFX1_HVT \keys_reg[10][72]  ( .D(n2325), .CLK(clk), .Q(\keys[10][72] ), 
        .QN(n1354) );
  DFFX1_HVT \keys_reg[10][71]  ( .D(n2324), .CLK(clk), .Q(\keys[10][71] ), 
        .QN(n1355) );
  DFFX1_HVT \keys_reg[10][70]  ( .D(n2323), .CLK(clk), .Q(\keys[10][70] ), 
        .QN(n1356) );
  DFFX1_HVT \keys_reg[10][69]  ( .D(n2322), .CLK(clk), .Q(\keys[10][69] ), 
        .QN(n1357) );
  DFFX1_HVT \keys_reg[10][68]  ( .D(n2321), .CLK(clk), .Q(\keys[10][68] ), 
        .QN(n1358) );
  DFFX1_HVT \keys_reg[10][67]  ( .D(n2320), .CLK(clk), .Q(\keys[10][67] ), 
        .QN(n1359) );
  DFFX1_HVT \keys_reg[10][66]  ( .D(n2319), .CLK(clk), .Q(\keys[10][66] ), 
        .QN(n1360) );
  DFFX1_HVT \keys_reg[10][65]  ( .D(n2318), .CLK(clk), .Q(\keys[10][65] ), 
        .QN(n1361) );
  DFFX1_HVT \keys_reg[10][64]  ( .D(n2317), .CLK(clk), .Q(\keys[10][64] ), 
        .QN(n1362) );
  DFFX1_HVT \keys_reg[10][63]  ( .D(n2316), .CLK(clk), .Q(\keys[10][63] ), 
        .QN(n1363) );
  DFFX1_HVT \keys_reg[10][62]  ( .D(n2315), .CLK(clk), .Q(\keys[10][62] ), 
        .QN(n1364) );
  DFFX1_HVT \keys_reg[10][61]  ( .D(n2314), .CLK(clk), .Q(\keys[10][61] ), 
        .QN(n1365) );
  DFFX1_HVT \keys_reg[10][60]  ( .D(n2313), .CLK(clk), .Q(\keys[10][60] ), 
        .QN(n1366) );
  DFFX1_HVT \keys_reg[10][59]  ( .D(n2312), .CLK(clk), .Q(\keys[10][59] ), 
        .QN(n1367) );
  DFFX1_HVT \keys_reg[10][58]  ( .D(n2311), .CLK(clk), .Q(\keys[10][58] ), 
        .QN(n1368) );
  DFFX1_HVT \keys_reg[10][57]  ( .D(n2310), .CLK(clk), .Q(\keys[10][57] ), 
        .QN(n1369) );
  DFFX1_HVT \keys_reg[10][56]  ( .D(n2309), .CLK(clk), .Q(\keys[10][56] ), 
        .QN(n1370) );
  DFFX1_HVT \keys_reg[10][55]  ( .D(n2308), .CLK(clk), .Q(\keys[10][55] ), 
        .QN(n1371) );
  DFFX1_HVT \keys_reg[10][54]  ( .D(n2307), .CLK(clk), .Q(\keys[10][54] ), 
        .QN(n1372) );
  DFFX1_HVT \keys_reg[10][53]  ( .D(n2306), .CLK(clk), .Q(\keys[10][53] ), 
        .QN(n1373) );
  DFFX1_HVT \keys_reg[10][52]  ( .D(n2305), .CLK(clk), .Q(\keys[10][52] ), 
        .QN(n1374) );
  DFFX1_HVT \keys_reg[10][51]  ( .D(n2304), .CLK(clk), .Q(\keys[10][51] ), 
        .QN(n1375) );
  DFFX1_HVT \keys_reg[10][50]  ( .D(n2303), .CLK(clk), .Q(\keys[10][50] ), 
        .QN(n1376) );
  DFFX1_HVT \keys_reg[10][49]  ( .D(n2302), .CLK(clk), .Q(\keys[10][49] ), 
        .QN(n1377) );
  DFFX1_HVT \keys_reg[10][48]  ( .D(n2301), .CLK(clk), .Q(\keys[10][48] ), 
        .QN(n1378) );
  DFFX1_HVT \keys_reg[10][47]  ( .D(n2300), .CLK(clk), .Q(\keys[10][47] ), 
        .QN(n1379) );
  DFFX1_HVT \keys_reg[10][46]  ( .D(n2299), .CLK(clk), .Q(\keys[10][46] ), 
        .QN(n1380) );
  DFFX1_HVT \keys_reg[10][45]  ( .D(n2298), .CLK(clk), .Q(\keys[10][45] ), 
        .QN(n1381) );
  DFFX1_HVT \keys_reg[10][44]  ( .D(n2297), .CLK(clk), .Q(\keys[10][44] ), 
        .QN(n1382) );
  DFFX1_HVT \keys_reg[10][43]  ( .D(n2296), .CLK(clk), .Q(\keys[10][43] ), 
        .QN(n1383) );
  DFFX1_HVT \keys_reg[10][42]  ( .D(n2295), .CLK(clk), .Q(\keys[10][42] ), 
        .QN(n1384) );
  DFFX1_HVT \keys_reg[10][41]  ( .D(n2294), .CLK(clk), .Q(\keys[10][41] ), 
        .QN(n1385) );
  DFFX1_HVT \keys_reg[10][40]  ( .D(n2293), .CLK(clk), .Q(\keys[10][40] ), 
        .QN(n1386) );
  DFFX1_HVT \keys_reg[10][39]  ( .D(n2292), .CLK(clk), .Q(\keys[10][39] ), 
        .QN(n1387) );
  DFFX1_HVT \keys_reg[10][38]  ( .D(n2291), .CLK(clk), .Q(\keys[10][38] ), 
        .QN(n1388) );
  DFFX1_HVT \keys_reg[10][37]  ( .D(n2290), .CLK(clk), .Q(\keys[10][37] ), 
        .QN(n1389) );
  DFFX1_HVT \keys_reg[10][36]  ( .D(n2289), .CLK(clk), .Q(\keys[10][36] ), 
        .QN(n1390) );
  DFFX1_HVT \keys_reg[10][35]  ( .D(n2288), .CLK(clk), .Q(\keys[10][35] ), 
        .QN(n1391) );
  DFFX1_HVT \keys_reg[10][34]  ( .D(n2287), .CLK(clk), .Q(\keys[10][34] ), 
        .QN(n1392) );
  DFFX1_HVT \keys_reg[10][33]  ( .D(n2286), .CLK(clk), .Q(\keys[10][33] ), 
        .QN(n1393) );
  DFFX1_HVT \keys_reg[10][32]  ( .D(n2285), .CLK(clk), .Q(\keys[10][32] ), 
        .QN(n1394) );
  DFFX1_HVT \keys_reg[10][31]  ( .D(n2284), .CLK(clk), .Q(\keys[10][31] ), 
        .QN(n1395) );
  DFFX1_HVT \keys_reg[10][30]  ( .D(n2283), .CLK(clk), .Q(\keys[10][30] ), 
        .QN(n1396) );
  DFFX1_HVT \keys_reg[10][29]  ( .D(n2282), .CLK(clk), .Q(\keys[10][29] ), 
        .QN(n1397) );
  DFFX1_HVT \keys_reg[10][28]  ( .D(n2281), .CLK(clk), .Q(\keys[10][28] ), 
        .QN(n1398) );
  DFFX1_HVT \keys_reg[10][27]  ( .D(n2280), .CLK(clk), .Q(\keys[10][27] ), 
        .QN(n1399) );
  DFFX1_HVT \keys_reg[10][26]  ( .D(n2279), .CLK(clk), .Q(\keys[10][26] ), 
        .QN(n1400) );
  DFFX1_HVT \keys_reg[10][25]  ( .D(n2278), .CLK(clk), .Q(\keys[10][25] ), 
        .QN(n1401) );
  DFFX1_HVT \keys_reg[10][24]  ( .D(n2277), .CLK(clk), .Q(\keys[10][24] ), 
        .QN(n1402) );
  DFFX1_HVT \keys_reg[10][23]  ( .D(n2276), .CLK(clk), .Q(\keys[10][23] ), 
        .QN(n1403) );
  DFFX1_HVT \keys_reg[10][22]  ( .D(n2275), .CLK(clk), .Q(\keys[10][22] ), 
        .QN(n1404) );
  DFFX1_HVT \keys_reg[10][21]  ( .D(n2274), .CLK(clk), .Q(\keys[10][21] ), 
        .QN(n1405) );
  DFFX1_HVT \keys_reg[10][20]  ( .D(n2273), .CLK(clk), .Q(\keys[10][20] ), 
        .QN(n1406) );
  DFFX1_HVT \keys_reg[10][19]  ( .D(n2272), .CLK(clk), .Q(\keys[10][19] ), 
        .QN(n1407) );
  DFFX1_HVT \keys_reg[10][18]  ( .D(n2271), .CLK(clk), .Q(\keys[10][18] ), 
        .QN(n1408) );
  DFFX1_HVT \keys_reg[10][17]  ( .D(n2270), .CLK(clk), .Q(\keys[10][17] ), 
        .QN(n1409) );
  DFFX1_HVT \keys_reg[10][16]  ( .D(n2269), .CLK(clk), .Q(\keys[10][16] ), 
        .QN(n1410) );
  DFFX1_HVT \keys_reg[10][15]  ( .D(n2268), .CLK(clk), .Q(\keys[10][15] ), 
        .QN(n1411) );
  DFFX1_HVT \keys_reg[10][14]  ( .D(n2267), .CLK(clk), .Q(\keys[10][14] ), 
        .QN(n1412) );
  DFFX1_HVT \keys_reg[10][13]  ( .D(n2266), .CLK(clk), .Q(\keys[10][13] ), 
        .QN(n1413) );
  DFFX1_HVT \keys_reg[10][12]  ( .D(n2265), .CLK(clk), .Q(\keys[10][12] ), 
        .QN(n1414) );
  DFFX1_HVT \keys_reg[10][11]  ( .D(n2264), .CLK(clk), .Q(\keys[10][11] ), 
        .QN(n1415) );
  DFFX1_HVT \keys_reg[10][10]  ( .D(n2263), .CLK(clk), .Q(\keys[10][10] ), 
        .QN(n1416) );
  DFFX1_HVT \keys_reg[10][9]  ( .D(n2262), .CLK(clk), .Q(\keys[10][9] ), .QN(
        n1417) );
  DFFX1_HVT \keys_reg[10][8]  ( .D(n2261), .CLK(clk), .Q(\keys[10][8] ), .QN(
        n1418) );
  DFFX1_HVT \keys_reg[10][7]  ( .D(n2260), .CLK(clk), .Q(\keys[10][7] ), .QN(
        n1419) );
  DFFX1_HVT \keys_reg[10][6]  ( .D(n2259), .CLK(clk), .Q(\keys[10][6] ), .QN(
        n1420) );
  DFFX1_HVT \keys_reg[10][5]  ( .D(n2258), .CLK(clk), .Q(\keys[10][5] ), .QN(
        n1421) );
  DFFX1_HVT \keys_reg[10][4]  ( .D(n2257), .CLK(clk), .Q(\keys[10][4] ), .QN(
        n1422) );
  DFFX1_HVT \keys_reg[10][3]  ( .D(n2256), .CLK(clk), .Q(\keys[10][3] ), .QN(
        n1423) );
  DFFX1_HVT \keys_reg[10][2]  ( .D(n2255), .CLK(clk), .Q(\keys[10][2] ), .QN(
        n1424) );
  DFFX1_HVT \keys_reg[10][1]  ( .D(n2254), .CLK(clk), .Q(\keys[10][1] ), .QN(
        n1425) );
  DFFX1_HVT \keys_reg[10][0]  ( .D(n2253), .CLK(clk), .Q(\keys[10][0] ), .QN(
        n1426) );
  DFFX1_HVT \key_round_reg[127]  ( .D(n2252), .CLK(clk), .Q(key_round[127]) );
  DFFX1_HVT \key_round_reg[126]  ( .D(n2251), .CLK(clk), .Q(key_round[126]) );
  DFFX1_HVT \key_round_reg[125]  ( .D(n2250), .CLK(clk), .Q(key_round[125]) );
  DFFX1_HVT \key_round_reg[124]  ( .D(n2249), .CLK(clk), .Q(key_round[124]) );
  DFFX1_HVT \key_round_reg[123]  ( .D(n2248), .CLK(clk), .Q(key_round[123]) );
  DFFX1_HVT \key_round_reg[122]  ( .D(n2247), .CLK(clk), .Q(key_round[122]) );
  DFFX1_HVT \key_round_reg[121]  ( .D(n2246), .CLK(clk), .Q(key_round[121]) );
  DFFX1_HVT \key_round_reg[120]  ( .D(n2245), .CLK(clk), .Q(key_round[120]) );
  DFFX1_HVT \key_round_reg[119]  ( .D(n2244), .CLK(clk), .Q(key_round[119]) );
  DFFX1_HVT \key_round_reg[118]  ( .D(n2243), .CLK(clk), .Q(key_round[118]) );
  DFFX1_HVT \key_round_reg[117]  ( .D(n2242), .CLK(clk), .Q(key_round[117]) );
  DFFX1_HVT \key_round_reg[116]  ( .D(n2241), .CLK(clk), .Q(key_round[116]) );
  DFFX1_HVT \key_round_reg[115]  ( .D(n2240), .CLK(clk), .Q(key_round[115]) );
  DFFX1_HVT \key_round_reg[114]  ( .D(n2239), .CLK(clk), .Q(key_round[114]) );
  DFFX1_HVT \key_round_reg[113]  ( .D(n2238), .CLK(clk), .Q(key_round[113]) );
  DFFX1_HVT \key_round_reg[112]  ( .D(n2237), .CLK(clk), .Q(key_round[112]) );
  DFFX1_HVT \key_round_reg[111]  ( .D(n2236), .CLK(clk), .Q(key_round[111]) );
  DFFX1_HVT \key_round_reg[110]  ( .D(n2235), .CLK(clk), .Q(key_round[110]) );
  DFFX1_HVT \key_round_reg[109]  ( .D(n2234), .CLK(clk), .Q(key_round[109]) );
  DFFX1_HVT \key_round_reg[108]  ( .D(n2233), .CLK(clk), .Q(key_round[108]) );
  DFFX1_HVT \key_round_reg[107]  ( .D(n2232), .CLK(clk), .Q(key_round[107]) );
  DFFX1_HVT \key_round_reg[106]  ( .D(n2231), .CLK(clk), .Q(key_round[106]) );
  DFFX1_HVT \key_round_reg[105]  ( .D(n2230), .CLK(clk), .Q(key_round[105]) );
  DFFX1_HVT \key_round_reg[104]  ( .D(n2229), .CLK(clk), .Q(key_round[104]) );
  DFFX1_HVT \key_round_reg[103]  ( .D(n2228), .CLK(clk), .Q(key_round[103]) );
  DFFX1_HVT \key_round_reg[102]  ( .D(n2227), .CLK(clk), .Q(key_round[102]) );
  DFFX1_HVT \key_round_reg[101]  ( .D(n2226), .CLK(clk), .Q(key_round[101]) );
  DFFX1_HVT \key_round_reg[100]  ( .D(n2225), .CLK(clk), .Q(key_round[100]) );
  DFFX1_HVT \key_round_reg[99]  ( .D(n2224), .CLK(clk), .Q(key_round[99]) );
  DFFX1_HVT \key_round_reg[98]  ( .D(n2223), .CLK(clk), .Q(key_round[98]) );
  DFFX1_HVT \key_round_reg[97]  ( .D(n2222), .CLK(clk), .Q(key_round[97]) );
  DFFX1_HVT \key_round_reg[96]  ( .D(n2221), .CLK(clk), .Q(key_round[96]) );
  DFFX1_HVT \key_round_reg[95]  ( .D(n2220), .CLK(clk), .Q(key_round[95]) );
  DFFX1_HVT \key_round_reg[94]  ( .D(n2219), .CLK(clk), .Q(key_round[94]) );
  DFFX1_HVT \key_round_reg[93]  ( .D(n2218), .CLK(clk), .Q(key_round[93]) );
  DFFX1_HVT \key_round_reg[92]  ( .D(n2217), .CLK(clk), .Q(key_round[92]) );
  DFFX1_HVT \key_round_reg[91]  ( .D(n2216), .CLK(clk), .Q(key_round[91]) );
  DFFX1_HVT \key_round_reg[90]  ( .D(n2215), .CLK(clk), .Q(key_round[90]) );
  DFFX1_HVT \key_round_reg[89]  ( .D(n2214), .CLK(clk), .Q(key_round[89]) );
  DFFX1_HVT \key_round_reg[88]  ( .D(n2213), .CLK(clk), .Q(key_round[88]) );
  DFFX1_HVT \key_round_reg[87]  ( .D(n2212), .CLK(clk), .Q(key_round[87]) );
  DFFX1_HVT \key_round_reg[86]  ( .D(n2211), .CLK(clk), .Q(key_round[86]) );
  DFFX1_HVT \key_round_reg[85]  ( .D(n2210), .CLK(clk), .Q(key_round[85]) );
  DFFX1_HVT \key_round_reg[84]  ( .D(n2209), .CLK(clk), .Q(key_round[84]) );
  DFFX1_HVT \key_round_reg[83]  ( .D(n2208), .CLK(clk), .Q(key_round[83]) );
  DFFX1_HVT \key_round_reg[82]  ( .D(n2207), .CLK(clk), .Q(key_round[82]) );
  DFFX1_HVT \key_round_reg[81]  ( .D(n2206), .CLK(clk), .Q(key_round[81]) );
  DFFX1_HVT \key_round_reg[80]  ( .D(n2205), .CLK(clk), .Q(key_round[80]) );
  DFFX1_HVT \key_round_reg[79]  ( .D(n2204), .CLK(clk), .Q(key_round[79]) );
  DFFX1_HVT \key_round_reg[78]  ( .D(n2203), .CLK(clk), .Q(key_round[78]) );
  DFFX1_HVT \key_round_reg[77]  ( .D(n2202), .CLK(clk), .Q(key_round[77]) );
  DFFX1_HVT \key_round_reg[76]  ( .D(n2201), .CLK(clk), .Q(key_round[76]) );
  DFFX1_HVT \key_round_reg[75]  ( .D(n2200), .CLK(clk), .Q(key_round[75]) );
  DFFX1_HVT \key_round_reg[74]  ( .D(n2199), .CLK(clk), .Q(key_round[74]) );
  DFFX1_HVT \key_round_reg[73]  ( .D(n2198), .CLK(clk), .Q(key_round[73]) );
  DFFX1_HVT \key_round_reg[72]  ( .D(n2197), .CLK(clk), .Q(key_round[72]) );
  DFFX1_HVT \key_round_reg[71]  ( .D(n2196), .CLK(clk), .Q(key_round[71]) );
  DFFX1_HVT \key_round_reg[70]  ( .D(n2195), .CLK(clk), .Q(key_round[70]) );
  DFFX1_HVT \key_round_reg[69]  ( .D(n2194), .CLK(clk), .Q(key_round[69]) );
  DFFX1_HVT \key_round_reg[68]  ( .D(n2193), .CLK(clk), .Q(key_round[68]) );
  DFFX1_HVT \key_round_reg[67]  ( .D(n2192), .CLK(clk), .Q(key_round[67]) );
  DFFX1_HVT \key_round_reg[66]  ( .D(n2191), .CLK(clk), .Q(key_round[66]) );
  DFFX1_HVT \key_round_reg[65]  ( .D(n2190), .CLK(clk), .Q(key_round[65]) );
  DFFX1_HVT \key_round_reg[64]  ( .D(n2189), .CLK(clk), .Q(key_round[64]) );
  DFFX1_HVT \key_round_reg[63]  ( .D(n2188), .CLK(clk), .Q(key_round[63]) );
  DFFX1_HVT \key_round_reg[62]  ( .D(n2187), .CLK(clk), .Q(key_round[62]) );
  DFFX1_HVT \key_round_reg[61]  ( .D(n2186), .CLK(clk), .Q(key_round[61]) );
  DFFX1_HVT \key_round_reg[60]  ( .D(n2185), .CLK(clk), .Q(key_round[60]) );
  DFFX1_HVT \key_round_reg[59]  ( .D(n2184), .CLK(clk), .Q(key_round[59]) );
  DFFX1_HVT \key_round_reg[58]  ( .D(n2183), .CLK(clk), .Q(key_round[58]) );
  DFFX1_HVT \key_round_reg[57]  ( .D(n2182), .CLK(clk), .Q(key_round[57]) );
  DFFX1_HVT \key_round_reg[56]  ( .D(n2181), .CLK(clk), .Q(key_round[56]) );
  DFFX1_HVT \key_round_reg[55]  ( .D(n2180), .CLK(clk), .Q(key_round[55]) );
  DFFX1_HVT \key_round_reg[54]  ( .D(n2179), .CLK(clk), .Q(key_round[54]) );
  DFFX1_HVT \key_round_reg[53]  ( .D(n2178), .CLK(clk), .Q(key_round[53]) );
  DFFX1_HVT \key_round_reg[52]  ( .D(n2177), .CLK(clk), .Q(key_round[52]) );
  DFFX1_HVT \key_round_reg[51]  ( .D(n2176), .CLK(clk), .Q(key_round[51]) );
  DFFX1_HVT \key_round_reg[50]  ( .D(n2175), .CLK(clk), .Q(key_round[50]) );
  DFFX1_HVT \key_round_reg[49]  ( .D(n2174), .CLK(clk), .Q(key_round[49]) );
  DFFX1_HVT \key_round_reg[48]  ( .D(n2173), .CLK(clk), .Q(key_round[48]) );
  DFFX1_HVT \key_round_reg[47]  ( .D(n2172), .CLK(clk), .Q(key_round[47]) );
  DFFX1_HVT \key_round_reg[46]  ( .D(n2171), .CLK(clk), .Q(key_round[46]) );
  DFFX1_HVT \key_round_reg[45]  ( .D(n2170), .CLK(clk), .Q(key_round[45]) );
  DFFX1_HVT \key_round_reg[44]  ( .D(n2169), .CLK(clk), .Q(key_round[44]) );
  DFFX1_HVT \key_round_reg[43]  ( .D(n2168), .CLK(clk), .Q(key_round[43]) );
  DFFX1_HVT \key_round_reg[42]  ( .D(n2167), .CLK(clk), .Q(key_round[42]) );
  DFFX1_HVT \key_round_reg[41]  ( .D(n2166), .CLK(clk), .Q(key_round[41]) );
  DFFX1_HVT \key_round_reg[40]  ( .D(n2165), .CLK(clk), .Q(key_round[40]) );
  DFFX1_HVT \key_round_reg[39]  ( .D(n2164), .CLK(clk), .Q(key_round[39]) );
  DFFX1_HVT \key_round_reg[38]  ( .D(n2163), .CLK(clk), .Q(key_round[38]) );
  DFFX1_HVT \key_round_reg[37]  ( .D(n2162), .CLK(clk), .Q(key_round[37]) );
  DFFX1_HVT \key_round_reg[36]  ( .D(n2161), .CLK(clk), .Q(key_round[36]) );
  DFFX1_HVT \key_round_reg[35]  ( .D(n2160), .CLK(clk), .Q(key_round[35]) );
  DFFX1_HVT \key_round_reg[34]  ( .D(n2159), .CLK(clk), .Q(key_round[34]) );
  DFFX1_HVT \key_round_reg[33]  ( .D(n2158), .CLK(clk), .Q(key_round[33]) );
  DFFX1_HVT \key_round_reg[32]  ( .D(n2157), .CLK(clk), .Q(key_round[32]) );
  DFFX1_HVT \key_round_reg[31]  ( .D(n2156), .CLK(clk), .Q(key_round[31]) );
  DFFX1_HVT \key_round_reg[30]  ( .D(n2155), .CLK(clk), .Q(key_round[30]) );
  DFFX1_HVT \key_round_reg[29]  ( .D(n2154), .CLK(clk), .Q(key_round[29]) );
  DFFX1_HVT \key_round_reg[28]  ( .D(n2153), .CLK(clk), .Q(key_round[28]) );
  DFFX1_HVT \key_round_reg[27]  ( .D(n2152), .CLK(clk), .Q(key_round[27]) );
  DFFX1_HVT \key_round_reg[26]  ( .D(n2151), .CLK(clk), .Q(key_round[26]) );
  DFFX1_HVT \key_round_reg[25]  ( .D(n2150), .CLK(clk), .Q(key_round[25]) );
  DFFX1_HVT \key_round_reg[24]  ( .D(n2149), .CLK(clk), .Q(key_round[24]) );
  DFFX1_HVT \key_round_reg[23]  ( .D(n2148), .CLK(clk), .Q(key_round[23]) );
  DFFX1_HVT \key_round_reg[22]  ( .D(n2147), .CLK(clk), .Q(key_round[22]) );
  DFFX1_HVT \key_round_reg[21]  ( .D(n2146), .CLK(clk), .Q(key_round[21]) );
  DFFX1_HVT \key_round_reg[20]  ( .D(n2145), .CLK(clk), .Q(key_round[20]) );
  DFFX1_HVT \key_round_reg[19]  ( .D(n2144), .CLK(clk), .Q(key_round[19]) );
  DFFX1_HVT \key_round_reg[18]  ( .D(n2143), .CLK(clk), .Q(key_round[18]) );
  DFFX1_HVT \key_round_reg[17]  ( .D(n2142), .CLK(clk), .Q(key_round[17]) );
  DFFX1_HVT \key_round_reg[16]  ( .D(n2141), .CLK(clk), .Q(key_round[16]) );
  DFFX1_HVT \key_round_reg[15]  ( .D(n2140), .CLK(clk), .Q(key_round[15]) );
  DFFX1_HVT \key_round_reg[14]  ( .D(n2139), .CLK(clk), .Q(key_round[14]) );
  DFFX1_HVT \key_round_reg[13]  ( .D(n2138), .CLK(clk), .Q(key_round[13]) );
  DFFX1_HVT \key_round_reg[12]  ( .D(n2137), .CLK(clk), .Q(key_round[12]) );
  DFFX1_HVT \key_round_reg[11]  ( .D(n2136), .CLK(clk), .Q(key_round[11]) );
  DFFX1_HVT \key_round_reg[10]  ( .D(n2135), .CLK(clk), .Q(key_round[10]) );
  DFFX1_HVT \key_round_reg[9]  ( .D(n2134), .CLK(clk), .Q(key_round[9]) );
  DFFX1_HVT \key_round_reg[8]  ( .D(n2133), .CLK(clk), .Q(key_round[8]) );
  DFFX1_HVT \key_round_reg[7]  ( .D(n2132), .CLK(clk), .Q(key_round[7]) );
  DFFX1_HVT \key_round_reg[6]  ( .D(n2131), .CLK(clk), .Q(key_round[6]) );
  DFFX1_HVT \key_round_reg[5]  ( .D(n2130), .CLK(clk), .Q(key_round[5]) );
  DFFX1_HVT \key_round_reg[4]  ( .D(n2129), .CLK(clk), .Q(key_round[4]) );
  DFFX1_HVT \key_round_reg[3]  ( .D(n2128), .CLK(clk), .Q(key_round[3]) );
  DFFX1_HVT \key_round_reg[2]  ( .D(n2127), .CLK(clk), .Q(key_round[2]) );
  DFFX1_HVT \key_round_reg[1]  ( .D(n2126), .CLK(clk), .Q(key_round[1]) );
  DFFX1_HVT \key_round_reg[0]  ( .D(n2125), .CLK(clk), .Q(key_round[0]) );
  AO22X1_HVT U20 ( .A1(n1427), .A2(n4534), .A3(\keys[10][48] ), .A4(n4518), 
        .Y(n2301) );
  AO22X1_HVT U21 ( .A1(n1429), .A2(n4542), .A3(\keys[10][49] ), .A4(n4512), 
        .Y(n2302) );
  AO22X1_HVT U22 ( .A1(n1432), .A2(n4544), .A3(\keys[10][50] ), .A4(n4512), 
        .Y(n2303) );
  AO22X1_HVT U23 ( .A1(n3937), .A2(n4544), .A3(\keys[10][51] ), .A4(n4512), 
        .Y(n2304) );
  AO22X1_HVT U24 ( .A1(n1434), .A2(n4544), .A3(\keys[10][52] ), .A4(n4512), 
        .Y(n2305) );
  AO22X1_HVT U25 ( .A1(n3920), .A2(n4544), .A3(\keys[10][53] ), .A4(n4512), 
        .Y(n2306) );
  AO22X1_HVT U26 ( .A1(n13), .A2(n4544), .A3(\keys[10][54] ), .A4(n4512), .Y(
        n2307) );
  AO22X1_HVT U27 ( .A1(n3922), .A2(n4544), .A3(\keys[10][55] ), .A4(n4512), 
        .Y(n2308) );
  AO22X1_HVT U28 ( .A1(n3941), .A2(n4544), .A3(\keys[10][56] ), .A4(n4512), 
        .Y(n2309) );
  AO22X1_HVT U29 ( .A1(n4084), .A2(n4544), .A3(\keys[10][57] ), .A4(n4512), 
        .Y(n2310) );
  AO22X1_HVT U30 ( .A1(n4086), .A2(n4544), .A3(\keys[10][58] ), .A4(n4512), 
        .Y(n2311) );
  AO22X1_HVT U31 ( .A1(n4089), .A2(n4544), .A3(\keys[10][59] ), .A4(n4512), 
        .Y(n2312) );
  AO22X1_HVT U32 ( .A1(n3943), .A2(n4544), .A3(\keys[10][60] ), .A4(n4513), 
        .Y(n2313) );
  AO22X1_HVT U33 ( .A1(n3805), .A2(n4544), .A3(\keys[10][61] ), .A4(n4513), 
        .Y(n2314) );
  AO22X1_HVT U34 ( .A1(n3832), .A2(n4544), .A3(\keys[10][62] ), .A4(n4513), 
        .Y(n2315) );
  AO22X1_HVT U35 ( .A1(n3860), .A2(n4544), .A3(\keys[10][63] ), .A4(n4513), 
        .Y(n2316) );
  AO22X1_HVT U36 ( .A1(keyout[64]), .A2(n4544), .A3(\keys[10][64] ), .A4(n4513), .Y(n2317) );
  AO22X1_HVT U37 ( .A1(n3883), .A2(n4543), .A3(\keys[10][65] ), .A4(n4513), 
        .Y(n2318) );
  AO22X1_HVT U38 ( .A1(n3914), .A2(n4543), .A3(\keys[10][66] ), .A4(n4513), 
        .Y(n2319) );
  AO22X1_HVT U39 ( .A1(n3825), .A2(n4543), .A3(\keys[10][67] ), .A4(n4513), 
        .Y(n2320) );
  AO22X1_HVT U40 ( .A1(keyout[68]), .A2(n4543), .A3(\keys[10][68] ), .A4(n4513), .Y(n2321) );
  AO22X1_HVT U41 ( .A1(keyout[69]), .A2(n4543), .A3(\keys[10][69] ), .A4(n4513), .Y(n2322) );
  AO22X1_HVT U42 ( .A1(keyout[70]), .A2(n4543), .A3(\keys[10][70] ), .A4(n4513), .Y(n2323) );
  AO22X1_HVT U43 ( .A1(keyout[71]), .A2(n4543), .A3(\keys[10][71] ), .A4(n4513), .Y(n2324) );
  AO22X1_HVT U44 ( .A1(n3951), .A2(n4543), .A3(\keys[10][72] ), .A4(n4514), 
        .Y(n2325) );
  AO22X1_HVT U45 ( .A1(n3896), .A2(n4543), .A3(\keys[10][73] ), .A4(n4514), 
        .Y(n2326) );
  AO22X1_HVT U46 ( .A1(n3979), .A2(n4543), .A3(\keys[10][74] ), .A4(n4514), 
        .Y(n2327) );
  AO22X1_HVT U47 ( .A1(n3959), .A2(n4543), .A3(\keys[10][75] ), .A4(n4514), 
        .Y(n2328) );
  AO22X1_HVT U48 ( .A1(n3966), .A2(n4543), .A3(\keys[10][76] ), .A4(n4514), 
        .Y(n2329) );
  AO22X1_HVT U49 ( .A1(n3985), .A2(n4543), .A3(\keys[10][77] ), .A4(n4514), 
        .Y(n2330) );
  AO22X1_HVT U50 ( .A1(n3946), .A2(n4543), .A3(\keys[10][78] ), .A4(n4514), 
        .Y(n2331) );
  AO22X1_HVT U51 ( .A1(n3898), .A2(n4542), .A3(\keys[10][79] ), .A4(n4514), 
        .Y(n2332) );
  AO22X1_HVT U52 ( .A1(n3931), .A2(n4542), .A3(\keys[10][80] ), .A4(n4514), 
        .Y(n2333) );
  AO22X1_HVT U53 ( .A1(n3811), .A2(n4542), .A3(\keys[10][81] ), .A4(n4514), 
        .Y(n2334) );
  AO22X1_HVT U54 ( .A1(n3977), .A2(n4542), .A3(\keys[10][82] ), .A4(n4514), 
        .Y(n2335) );
  AO22X1_HVT U55 ( .A1(n3916), .A2(n4542), .A3(\keys[10][83] ), .A4(n4514), 
        .Y(n2336) );
  AO22X1_HVT U56 ( .A1(n1438), .A2(n4542), .A3(\keys[10][84] ), .A4(n4515), 
        .Y(n2337) );
  AO22X1_HVT U57 ( .A1(n2), .A2(n4542), .A3(\keys[10][85] ), .A4(n4515), .Y(
        n2338) );
  AO22X1_HVT U58 ( .A1(n1436), .A2(n4542), .A3(\keys[10][86] ), .A4(n4515), 
        .Y(n2339) );
  AO22X1_HVT U59 ( .A1(n1439), .A2(n4542), .A3(\keys[10][87] ), .A4(n4515), 
        .Y(n2340) );
  AO22X1_HVT U60 ( .A1(n4093), .A2(n4542), .A3(\keys[10][88] ), .A4(n4515), 
        .Y(n2341) );
  AO22X1_HVT U61 ( .A1(n3863), .A2(n4542), .A3(\keys[10][89] ), .A4(n4515), 
        .Y(n2342) );
  AO22X1_HVT U63 ( .A1(n3816), .A2(n4542), .A3(\keys[10][91] ), .A4(n4515), 
        .Y(n2344) );
  AO22X1_HVT U64 ( .A1(n3831), .A2(n4542), .A3(\keys[10][92] ), .A4(n4515), 
        .Y(n2345) );
  AO22X1_HVT U65 ( .A1(keyout[93]), .A2(n4541), .A3(\keys[10][93] ), .A4(n4515), .Y(n2346) );
  AO22X1_HVT U66 ( .A1(n3835), .A2(n4541), .A3(\keys[10][94] ), .A4(n4515), 
        .Y(n2347) );
  AO22X1_HVT U67 ( .A1(n3869), .A2(n4541), .A3(\keys[10][95] ), .A4(n4515), 
        .Y(n2348) );
  AO22X1_HVT U68 ( .A1(keyout[96]), .A2(n4541), .A3(\keys[10][96] ), .A4(n4516), .Y(n2349) );
  AO22X1_HVT U69 ( .A1(keyout[97]), .A2(n4545), .A3(\keys[10][97] ), .A4(n4516), .Y(n2350) );
  AO22X1_HVT U70 ( .A1(keyout[98]), .A2(n4545), .A3(\keys[10][98] ), .A4(n4516), .Y(n2351) );
  AO22X1_HVT U71 ( .A1(keyout[99]), .A2(n4545), .A3(\keys[10][99] ), .A4(n4516), .Y(n2352) );
  AO22X1_HVT U72 ( .A1(keyout[100]), .A2(n4545), .A3(\keys[10][100] ), .A4(
        n4516), .Y(n2353) );
  AO22X1_HVT U73 ( .A1(keyout[101]), .A2(n4545), .A3(\keys[10][101] ), .A4(
        n4516), .Y(n2354) );
  AO22X1_HVT U74 ( .A1(keyout[102]), .A2(n4545), .A3(\keys[10][102] ), .A4(
        n4516), .Y(n2355) );
  AO22X1_HVT U75 ( .A1(keyout[103]), .A2(n4545), .A3(\keys[10][103] ), .A4(
        n4516), .Y(n2356) );
  AO22X1_HVT U76 ( .A1(n3839), .A2(n4545), .A3(\keys[10][104] ), .A4(n4516), 
        .Y(n2357) );
  AO22X1_HVT U77 ( .A1(keyout[105]), .A2(n4545), .A3(\keys[10][105] ), .A4(
        n4516), .Y(n2358) );
  AO22X1_HVT U78 ( .A1(n3880), .A2(n4545), .A3(\keys[10][106] ), .A4(n4516), 
        .Y(n2359) );
  AO22X1_HVT U79 ( .A1(n3820), .A2(n4545), .A3(\keys[10][107] ), .A4(n4516), 
        .Y(n2360) );
  AO22X1_HVT U80 ( .A1(n3892), .A2(n4545), .A3(\keys[10][108] ), .A4(n4517), 
        .Y(n2361) );
  AO22X1_HVT U81 ( .A1(n3873), .A2(n4545), .A3(\keys[10][109] ), .A4(n4517), 
        .Y(n2362) );
  AO22X1_HVT U82 ( .A1(keyout[110]), .A2(n4545), .A3(\keys[10][110] ), .A4(
        n4517), .Y(n2363) );
  AO22X1_HVT U83 ( .A1(keyout[111]), .A2(n4545), .A3(\keys[10][111] ), .A4(
        n4517), .Y(n2364) );
  AO22X1_HVT U84 ( .A1(keyout[112]), .A2(n4541), .A3(\keys[10][112] ), .A4(
        n4517), .Y(n2365) );
  AO22X1_HVT U85 ( .A1(keyout[113]), .A2(n4541), .A3(\keys[10][113] ), .A4(
        n4517), .Y(n2366) );
  AO22X1_HVT U86 ( .A1(keyout[114]), .A2(n4541), .A3(\keys[10][114] ), .A4(
        n4517), .Y(n2367) );
  AO22X1_HVT U87 ( .A1(n3915), .A2(n4541), .A3(\keys[10][115] ), .A4(n4517), 
        .Y(n2368) );
  AO22X1_HVT U88 ( .A1(keyout[116]), .A2(n4541), .A3(\keys[10][116] ), .A4(
        n4517), .Y(n2369) );
  AO22X1_HVT U89 ( .A1(keyout[117]), .A2(n4541), .A3(\keys[10][117] ), .A4(
        n4517), .Y(n2370) );
  AO22X1_HVT U90 ( .A1(keyout[118]), .A2(n4541), .A3(\keys[10][118] ), .A4(
        n4517), .Y(n2371) );
  AO22X1_HVT U91 ( .A1(keyout[119]), .A2(n4541), .A3(\keys[10][119] ), .A4(
        n4517), .Y(n2372) );
  AO22X1_HVT U92 ( .A1(n4096), .A2(n4541), .A3(\keys[10][120] ), .A4(n4518), 
        .Y(n2373) );
  AO22X1_HVT U93 ( .A1(n3829), .A2(n4541), .A3(\keys[10][121] ), .A4(n4518), 
        .Y(n2374) );
  AO22X1_HVT U94 ( .A1(n3803), .A2(n4541), .A3(\keys[10][122] ), .A4(n4518), 
        .Y(n2375) );
  AO22X1_HVT U95 ( .A1(n3817), .A2(n4540), .A3(\keys[10][123] ), .A4(n4518), 
        .Y(n2376) );
  AO22X1_HVT U96 ( .A1(n3845), .A2(n4540), .A3(\keys[10][124] ), .A4(n4518), 
        .Y(n2377) );
  AO22X1_HVT U97 ( .A1(n3823), .A2(n4540), .A3(\keys[10][125] ), .A4(n4518), 
        .Y(n2378) );
  AO22X1_HVT U98 ( .A1(n4099), .A2(n4540), .A3(\keys[10][126] ), .A4(n4518), 
        .Y(n2379) );
  AO22X1_HVT U99 ( .A1(n4102), .A2(n4540), .A3(\keys[10][127] ), .A4(n4518), 
        .Y(n2380) );
  AO22X1_HVT U100 ( .A1(n3999), .A2(n4497), .A3(\keys[9][0] ), .A4(n4491), .Y(
        n2381) );
  AO22X1_HVT U101 ( .A1(n4002), .A2(n4498), .A3(\keys[9][1] ), .A4(n4486), .Y(
        n2382) );
  AO22X1_HVT U102 ( .A1(n4003), .A2(n4498), .A3(\keys[9][2] ), .A4(n4486), .Y(
        n2383) );
  AO22X1_HVT U103 ( .A1(n4006), .A2(n4498), .A3(\keys[9][3] ), .A4(n4486), .Y(
        n2384) );
  AO22X1_HVT U104 ( .A1(n4009), .A2(n4499), .A3(\keys[9][4] ), .A4(n4486), .Y(
        n2385) );
  AO22X1_HVT U105 ( .A1(n4012), .A2(n4499), .A3(\keys[9][5] ), .A4(n4486), .Y(
        n2386) );
  AO22X1_HVT U106 ( .A1(n4015), .A2(n4499), .A3(\keys[9][6] ), .A4(n4486), .Y(
        n2387) );
  AO22X1_HVT U107 ( .A1(n4016), .A2(n4499), .A3(\keys[9][7] ), .A4(n4486), .Y(
        n2388) );
  AO22X1_HVT U108 ( .A1(n4019), .A2(n4499), .A3(\keys[9][8] ), .A4(n4486), .Y(
        n2389) );
  AO22X1_HVT U109 ( .A1(n4499), .A2(n4022), .A3(\keys[9][9] ), .A4(n4486), .Y(
        n2390) );
  AO22X1_HVT U110 ( .A1(n4025), .A2(n4499), .A3(\keys[9][10] ), .A4(n4486), 
        .Y(n2391) );
  AO22X1_HVT U111 ( .A1(n4499), .A2(n4028), .A3(\keys[9][11] ), .A4(n4486), 
        .Y(n2392) );
  AO22X1_HVT U112 ( .A1(n4031), .A2(n4499), .A3(\keys[9][12] ), .A4(n4486), 
        .Y(n2393) );
  AO22X1_HVT U113 ( .A1(n4034), .A2(n4499), .A3(\keys[9][13] ), .A4(n4487), 
        .Y(n2394) );
  AO22X1_HVT U114 ( .A1(n4037), .A2(n4499), .A3(\keys[9][14] ), .A4(n4487), 
        .Y(n2395) );
  AO22X1_HVT U115 ( .A1(n4040), .A2(n4499), .A3(\keys[9][15] ), .A4(n4487), 
        .Y(n2396) );
  AO22X1_HVT U116 ( .A1(n4043), .A2(n4499), .A3(\keys[9][16] ), .A4(n4487), 
        .Y(n2397) );
  AO22X1_HVT U117 ( .A1(n4046), .A2(n4499), .A3(\keys[9][17] ), .A4(n4487), 
        .Y(n2398) );
  AO22X1_HVT U118 ( .A1(n4049), .A2(n4499), .A3(\keys[9][18] ), .A4(n4487), 
        .Y(n2399) );
  AO22X1_HVT U119 ( .A1(n4052), .A2(n4500), .A3(\keys[9][19] ), .A4(n4487), 
        .Y(n2400) );
  AO22X1_HVT U120 ( .A1(n4055), .A2(n4500), .A3(\keys[9][20] ), .A4(n4487), 
        .Y(n2401) );
  AO22X1_HVT U121 ( .A1(n4058), .A2(n4500), .A3(\keys[9][21] ), .A4(n4487), 
        .Y(n2402) );
  AO22X1_HVT U122 ( .A1(n4061), .A2(n4500), .A3(\keys[9][22] ), .A4(n4487), 
        .Y(n2403) );
  AO22X1_HVT U123 ( .A1(n4064), .A2(n4500), .A3(\keys[9][23] ), .A4(n4487), 
        .Y(n2404) );
  AO22X1_HVT U124 ( .A1(n4067), .A2(n4500), .A3(\keys[9][24] ), .A4(n4487), 
        .Y(n2405) );
  AO22X1_HVT U125 ( .A1(n4069), .A2(n4500), .A3(\keys[9][25] ), .A4(n4488), 
        .Y(n2406) );
  AO22X1_HVT U126 ( .A1(n4072), .A2(n4500), .A3(\keys[9][26] ), .A4(n4488), 
        .Y(n2407) );
  AO22X1_HVT U127 ( .A1(n4075), .A2(n4500), .A3(\keys[9][27] ), .A4(n4488), 
        .Y(n2408) );
  AO22X1_HVT U128 ( .A1(n4078), .A2(n4500), .A3(\keys[9][28] ), .A4(n4488), 
        .Y(n2409) );
  AO22X1_HVT U129 ( .A1(n4081), .A2(n4500), .A3(\keys[9][29] ), .A4(n4488), 
        .Y(n2410) );
  AO22X1_HVT U130 ( .A1(n4083), .A2(n4500), .A3(\keys[9][30] ), .A4(n4488), 
        .Y(n2411) );
  AO22X1_HVT U131 ( .A1(n3852), .A2(n4500), .A3(\keys[9][31] ), .A4(n4488), 
        .Y(n2412) );
  AO22X1_HVT U132 ( .A1(keyout[32]), .A2(n4500), .A3(\keys[9][32] ), .A4(n4488), .Y(n2413) );
  AO22X1_HVT U133 ( .A1(n3876), .A2(n4500), .A3(\keys[9][33] ), .A4(n4488), 
        .Y(n2414) );
  AO22X1_HVT U134 ( .A1(n3913), .A2(n4501), .A3(\keys[9][34] ), .A4(n4488), 
        .Y(n2415) );
  AO22X1_HVT U135 ( .A1(keyout[35]), .A2(n4501), .A3(\keys[9][35] ), .A4(n4488), .Y(n2416) );
  AO22X1_HVT U136 ( .A1(keyout[36]), .A2(n4501), .A3(\keys[9][36] ), .A4(n4488), .Y(n2417) );
  AO22X1_HVT U137 ( .A1(n3911), .A2(n4501), .A3(\keys[9][37] ), .A4(n4489), 
        .Y(n2418) );
  AO22X1_HVT U138 ( .A1(keyout[38]), .A2(n4501), .A3(\keys[9][38] ), .A4(n4489), .Y(n2419) );
  AO22X1_HVT U139 ( .A1(keyout[39]), .A2(n4501), .A3(\keys[9][39] ), .A4(n4489), .Y(n2420) );
  AO22X1_HVT U140 ( .A1(n3953), .A2(n4501), .A3(\keys[9][40] ), .A4(n4489), 
        .Y(n2421) );
  AO22X1_HVT U141 ( .A1(n3854), .A2(n4501), .A3(\keys[9][41] ), .A4(n4489), 
        .Y(n2422) );
  AO22X1_HVT U142 ( .A1(n3973), .A2(n4501), .A3(\keys[9][42] ), .A4(n4489), 
        .Y(n2423) );
  AO22X1_HVT U143 ( .A1(n3890), .A2(n4501), .A3(\keys[9][43] ), .A4(n4489), 
        .Y(n2424) );
  AO22X1_HVT U144 ( .A1(n3902), .A2(n4501), .A3(\keys[9][44] ), .A4(n4489), 
        .Y(n2425) );
  AO22X1_HVT U145 ( .A1(n3935), .A2(n4501), .A3(\keys[9][45] ), .A4(n4489), 
        .Y(n2426) );
  AO22X1_HVT U146 ( .A1(n3945), .A2(n4501), .A3(\keys[9][46] ), .A4(n4489), 
        .Y(n2427) );
  AO22X1_HVT U147 ( .A1(n3885), .A2(n4501), .A3(\keys[9][47] ), .A4(n4489), 
        .Y(n2428) );
  AO22X1_HVT U148 ( .A1(n4501), .A2(keyout[48]), .A3(\keys[9][48] ), .A4(n4489), .Y(n2429) );
  AO22X1_HVT U149 ( .A1(n4502), .A2(n14), .A3(\keys[9][49] ), .A4(n4490), .Y(
        n2430) );
  AO22X1_HVT U150 ( .A1(n4502), .A2(keyout[50]), .A3(\keys[9][50] ), .A4(n4490), .Y(n2431) );
  AO22X1_HVT U151 ( .A1(n4502), .A2(keyout[51]), .A3(\keys[9][51] ), .A4(n4490), .Y(n2432) );
  AO22X1_HVT U152 ( .A1(n4502), .A2(keyout[52]), .A3(\keys[9][52] ), .A4(n4490), .Y(n2433) );
  AO22X1_HVT U153 ( .A1(n4502), .A2(n3874), .A3(\keys[9][53] ), .A4(n4490), 
        .Y(n2434) );
  AO22X1_HVT U154 ( .A1(n4502), .A2(keyout[54]), .A3(\keys[9][54] ), .A4(n4490), .Y(n2435) );
  AO22X1_HVT U155 ( .A1(n4502), .A2(n3866), .A3(\keys[9][55] ), .A4(n4490), 
        .Y(n2436) );
  AO22X1_HVT U156 ( .A1(n4502), .A2(keyout[56]), .A3(\keys[9][56] ), .A4(n4490), .Y(n2437) );
  AO22X1_HVT U157 ( .A1(n4502), .A2(n4084), .A3(\keys[9][57] ), .A4(n4490), 
        .Y(n2438) );
  AO22X1_HVT U158 ( .A1(n4502), .A2(n4086), .A3(\keys[9][58] ), .A4(n4490), 
        .Y(n2439) );
  AO22X1_HVT U159 ( .A1(n4502), .A2(n4088), .A3(\keys[9][59] ), .A4(n4490), 
        .Y(n2440) );
  AO22X1_HVT U160 ( .A1(n4502), .A2(keyout[60]), .A3(\keys[9][60] ), .A4(n4490), .Y(n2441) );
  AO22X1_HVT U161 ( .A1(n4502), .A2(keyout[61]), .A3(\keys[9][61] ), .A4(n4491), .Y(n2442) );
  AO22X1_HVT U162 ( .A1(n4502), .A2(n3833), .A3(\keys[9][62] ), .A4(n4491), 
        .Y(n2443) );
  AO22X1_HVT U163 ( .A1(n4502), .A2(n3859), .A3(\keys[9][63] ), .A4(n4491), 
        .Y(n2444) );
  AO22X1_HVT U164 ( .A1(n4502), .A2(keyout[64]), .A3(\keys[9][64] ), .A4(n4491), .Y(n2445) );
  AO22X1_HVT U165 ( .A1(n4503), .A2(n3870), .A3(\keys[9][65] ), .A4(n4491), 
        .Y(n2446) );
  AO22X1_HVT U166 ( .A1(n4503), .A2(keyout[66]), .A3(\keys[9][66] ), .A4(n4491), .Y(n2447) );
  AO22X1_HVT U167 ( .A1(n4503), .A2(n3938), .A3(\keys[9][67] ), .A4(n4491), 
        .Y(n2448) );
  AO22X1_HVT U168 ( .A1(n4503), .A2(keyout[68]), .A3(\keys[9][68] ), .A4(n4491), .Y(n2449) );
  AO22X1_HVT U169 ( .A1(n4503), .A2(keyout[69]), .A3(\keys[9][69] ), .A4(n4491), .Y(n2450) );
  AO22X1_HVT U170 ( .A1(n4503), .A2(keyout[70]), .A3(\keys[9][70] ), .A4(n4491), .Y(n2451) );
  AO22X1_HVT U171 ( .A1(n4503), .A2(keyout[71]), .A3(\keys[9][71] ), .A4(n4491), .Y(n2452) );
  AO22X1_HVT U172 ( .A1(n4503), .A2(n3939), .A3(\keys[9][72] ), .A4(n4492), 
        .Y(n2453) );
  AO22X1_HVT U173 ( .A1(n4503), .A2(n3886), .A3(\keys[9][73] ), .A4(n4492), 
        .Y(n2454) );
  AO22X1_HVT U174 ( .A1(n4503), .A2(n3872), .A3(\keys[9][74] ), .A4(n4492), 
        .Y(n2455) );
  AO22X1_HVT U175 ( .A1(n4503), .A2(n3960), .A3(\keys[9][75] ), .A4(n4492), 
        .Y(n2456) );
  AO22X1_HVT U176 ( .A1(n4503), .A2(n3965), .A3(\keys[9][76] ), .A4(n4492), 
        .Y(n2457) );
  AO22X1_HVT U177 ( .A1(n4503), .A2(n3984), .A3(\keys[9][77] ), .A4(n4492), 
        .Y(n2458) );
  AO22X1_HVT U178 ( .A1(n4503), .A2(n3947), .A3(\keys[9][78] ), .A4(n4492), 
        .Y(n2459) );
  AO22X1_HVT U179 ( .A1(n4503), .A2(n3887), .A3(\keys[9][79] ), .A4(n4492), 
        .Y(n2460) );
  AO22X1_HVT U180 ( .A1(n4503), .A2(keyout[80]), .A3(\keys[9][80] ), .A4(n4492), .Y(n2461) );
  AO22X1_HVT U181 ( .A1(n4504), .A2(keyout[81]), .A3(\keys[9][81] ), .A4(n4492), .Y(n2462) );
  AO22X1_HVT U182 ( .A1(n4504), .A2(keyout[82]), .A3(\keys[9][82] ), .A4(n4492), .Y(n2463) );
  AO22X1_HVT U183 ( .A1(n4504), .A2(n3904), .A3(\keys[9][83] ), .A4(n4492), 
        .Y(n2464) );
  AO22X1_HVT U184 ( .A1(n4504), .A2(keyout[84]), .A3(\keys[9][84] ), .A4(n4493), .Y(n2465) );
  AO22X1_HVT U185 ( .A1(n4504), .A2(n1), .A3(\keys[9][85] ), .A4(n4493), .Y(
        n2466) );
  AO22X1_HVT U186 ( .A1(n4504), .A2(keyout[86]), .A3(\keys[9][86] ), .A4(n4493), .Y(n2467) );
  AO22X1_HVT U187 ( .A1(n4504), .A2(n1440), .A3(\keys[9][87] ), .A4(n4493), 
        .Y(n2468) );
  AO22X1_HVT U188 ( .A1(n4504), .A2(n4092), .A3(\keys[9][88] ), .A4(n4493), 
        .Y(n2469) );
  AO22X1_HVT U189 ( .A1(n4504), .A2(n3827), .A3(\keys[9][89] ), .A4(n4493), 
        .Y(n2470) );
  AO22X1_HVT U190 ( .A1(n4504), .A2(keyout[90]), .A3(\keys[9][90] ), .A4(n4493), .Y(n2471) );
  AO22X1_HVT U191 ( .A1(n4504), .A2(keyout[91]), .A3(\keys[9][91] ), .A4(n4493), .Y(n2472) );
  AO22X1_HVT U192 ( .A1(n4504), .A2(keyout[92]), .A3(\keys[9][92] ), .A4(n4493), .Y(n2473) );
  AO22X1_HVT U193 ( .A1(n4504), .A2(keyout[93]), .A3(\keys[9][93] ), .A4(n4493), .Y(n2474) );
  AO22X1_HVT U194 ( .A1(n4504), .A2(n3865), .A3(\keys[9][94] ), .A4(n4493), 
        .Y(n2475) );
  AO22X1_HVT U195 ( .A1(n4504), .A2(keyout[95]), .A3(\keys[9][95] ), .A4(n4493), .Y(n2476) );
  AO22X1_HVT U196 ( .A1(n4504), .A2(keyout[96]), .A3(\keys[9][96] ), .A4(n4494), .Y(n2477) );
  AO22X1_HVT U197 ( .A1(n4505), .A2(keyout[97]), .A3(\keys[9][97] ), .A4(n4494), .Y(n2478) );
  AO22X1_HVT U198 ( .A1(n4505), .A2(keyout[98]), .A3(\keys[9][98] ), .A4(n4494), .Y(n2479) );
  AO22X1_HVT U199 ( .A1(n4505), .A2(keyout[99]), .A3(\keys[9][99] ), .A4(n4494), .Y(n2480) );
  AO22X1_HVT U200 ( .A1(n4505), .A2(keyout[100]), .A3(\keys[9][100] ), .A4(
        n4494), .Y(n2481) );
  AO22X1_HVT U201 ( .A1(n4505), .A2(keyout[101]), .A3(\keys[9][101] ), .A4(
        n4494), .Y(n2482) );
  AO22X1_HVT U202 ( .A1(n4505), .A2(keyout[102]), .A3(\keys[9][102] ), .A4(
        n4494), .Y(n2483) );
  AO22X1_HVT U203 ( .A1(n4505), .A2(keyout[103]), .A3(\keys[9][103] ), .A4(
        n4494), .Y(n2484) );
  AO22X1_HVT U204 ( .A1(n4505), .A2(keyout[104]), .A3(\keys[9][104] ), .A4(
        n4494), .Y(n2485) );
  AO22X1_HVT U205 ( .A1(n4505), .A2(keyout[105]), .A3(\keys[9][105] ), .A4(
        n4494), .Y(n2486) );
  AO22X1_HVT U206 ( .A1(n4505), .A2(keyout[106]), .A3(\keys[9][106] ), .A4(
        n4494), .Y(n2487) );
  AO22X1_HVT U207 ( .A1(n4505), .A2(keyout[107]), .A3(\keys[9][107] ), .A4(
        n4494), .Y(n2488) );
  AO22X1_HVT U208 ( .A1(n4505), .A2(n3881), .A3(\keys[9][108] ), .A4(n4495), 
        .Y(n2489) );
  AO22X1_HVT U209 ( .A1(n4505), .A2(keyout[109]), .A3(\keys[9][109] ), .A4(
        n4495), .Y(n2490) );
  AO22X1_HVT U210 ( .A1(n4505), .A2(keyout[110]), .A3(\keys[9][110] ), .A4(
        n4495), .Y(n2491) );
  AO22X1_HVT U211 ( .A1(n4505), .A2(keyout[111]), .A3(\keys[9][111] ), .A4(
        n4495), .Y(n2492) );
  AO22X1_HVT U212 ( .A1(n4505), .A2(keyout[112]), .A3(\keys[9][112] ), .A4(
        n4495), .Y(n2493) );
  AO22X1_HVT U213 ( .A1(n4506), .A2(keyout[113]), .A3(\keys[9][113] ), .A4(
        n4495), .Y(n2494) );
  AO22X1_HVT U214 ( .A1(n4506), .A2(keyout[114]), .A3(\keys[9][114] ), .A4(
        n4495), .Y(n2495) );
  AO22X1_HVT U215 ( .A1(n4506), .A2(keyout[115]), .A3(\keys[9][115] ), .A4(
        n4495), .Y(n2496) );
  AO22X1_HVT U216 ( .A1(n4506), .A2(keyout[116]), .A3(\keys[9][116] ), .A4(
        n4495), .Y(n2497) );
  AO22X1_HVT U217 ( .A1(n4506), .A2(keyout[117]), .A3(\keys[9][117] ), .A4(
        n4495), .Y(n2498) );
  AO22X1_HVT U218 ( .A1(n4506), .A2(keyout[118]), .A3(\keys[9][118] ), .A4(
        n4495), .Y(n2499) );
  AO22X1_HVT U219 ( .A1(n4506), .A2(keyout[119]), .A3(\keys[9][119] ), .A4(
        n4495), .Y(n2500) );
  AO22X1_HVT U220 ( .A1(n4506), .A2(n4095), .A3(\keys[9][120] ), .A4(n4496), 
        .Y(n2501) );
  AO22X1_HVT U221 ( .A1(n4506), .A2(n3829), .A3(\keys[9][121] ), .A4(n4496), 
        .Y(n2502) );
  AO22X1_HVT U222 ( .A1(n4506), .A2(n3803), .A3(\keys[9][122] ), .A4(n4496), 
        .Y(n2503) );
  AO22X1_HVT U223 ( .A1(n4506), .A2(n3817), .A3(\keys[9][123] ), .A4(n4496), 
        .Y(n2504) );
  AO22X1_HVT U224 ( .A1(n4506), .A2(n3846), .A3(\keys[9][124] ), .A4(n4496), 
        .Y(n2505) );
  AO22X1_HVT U225 ( .A1(n4506), .A2(n3823), .A3(\keys[9][125] ), .A4(n4496), 
        .Y(n2506) );
  AO22X1_HVT U226 ( .A1(n4506), .A2(n4098), .A3(\keys[9][126] ), .A4(n4496), 
        .Y(n2507) );
  AO22X1_HVT U227 ( .A1(n4506), .A2(n4101), .A3(\keys[9][127] ), .A4(n4496), 
        .Y(n2508) );
  AO22X1_HVT U228 ( .A1(n4474), .A2(n3997), .A3(\keys[8][0] ), .A4(n4473), .Y(
        n2509) );
  AO22X1_HVT U229 ( .A1(n4475), .A2(n4000), .A3(\keys[8][1] ), .A4(n4473), .Y(
        n2510) );
  AO22X1_HVT U230 ( .A1(n4475), .A2(keyout[2]), .A3(\keys[8][2] ), .A4(n4473), 
        .Y(n2511) );
  AO22X1_HVT U231 ( .A1(n4475), .A2(n4004), .A3(\keys[8][3] ), .A4(n4473), .Y(
        n2512) );
  AO22X1_HVT U232 ( .A1(n4475), .A2(n4007), .A3(\keys[8][4] ), .A4(n4473), .Y(
        n2513) );
  AO22X1_HVT U233 ( .A1(n4475), .A2(n4010), .A3(\keys[8][5] ), .A4(n4473), .Y(
        n2514) );
  AO22X1_HVT U234 ( .A1(n4475), .A2(n4013), .A3(\keys[8][6] ), .A4(n4473), .Y(
        n2515) );
  AO22X1_HVT U235 ( .A1(n4476), .A2(keyout[7]), .A3(\keys[8][7] ), .A4(n4473), 
        .Y(n2516) );
  AO22X1_HVT U236 ( .A1(n4476), .A2(n4017), .A3(\keys[8][8] ), .A4(n4473), .Y(
        n2517) );
  AO22X1_HVT U237 ( .A1(n4476), .A2(n4020), .A3(\keys[8][9] ), .A4(n4473), .Y(
        n2518) );
  AO22X1_HVT U238 ( .A1(n4476), .A2(n4023), .A3(\keys[8][10] ), .A4(n4473), 
        .Y(n2519) );
  AO22X1_HVT U239 ( .A1(n4476), .A2(n4026), .A3(\keys[8][11] ), .A4(n4473), 
        .Y(n2520) );
  AO22X1_HVT U240 ( .A1(n4476), .A2(n4029), .A3(\keys[8][12] ), .A4(n4473), 
        .Y(n2521) );
  AO22X1_HVT U241 ( .A1(n4476), .A2(n4032), .A3(\keys[8][13] ), .A4(n4472), 
        .Y(n2522) );
  AO22X1_HVT U242 ( .A1(n4476), .A2(n4035), .A3(\keys[8][14] ), .A4(n4472), 
        .Y(n2523) );
  AO22X1_HVT U243 ( .A1(n4476), .A2(n4038), .A3(\keys[8][15] ), .A4(n4472), 
        .Y(n2524) );
  AO22X1_HVT U244 ( .A1(n4476), .A2(n4041), .A3(\keys[8][16] ), .A4(n4472), 
        .Y(n2525) );
  AO22X1_HVT U245 ( .A1(n4476), .A2(n4044), .A3(\keys[8][17] ), .A4(n4472), 
        .Y(n2526) );
  AO22X1_HVT U246 ( .A1(n4476), .A2(n4047), .A3(\keys[8][18] ), .A4(n4472), 
        .Y(n2527) );
  AO22X1_HVT U247 ( .A1(n4476), .A2(n4050), .A3(\keys[8][19] ), .A4(n4472), 
        .Y(n2528) );
  AO22X1_HVT U248 ( .A1(n4476), .A2(n4053), .A3(\keys[8][20] ), .A4(n4472), 
        .Y(n2529) );
  AO22X1_HVT U249 ( .A1(n4476), .A2(n4056), .A3(\keys[8][21] ), .A4(n4472), 
        .Y(n2530) );
  AO22X1_HVT U250 ( .A1(n4476), .A2(n4059), .A3(\keys[8][22] ), .A4(n4472), 
        .Y(n2531) );
  AO22X1_HVT U251 ( .A1(n4477), .A2(n4062), .A3(\keys[8][23] ), .A4(n4472), 
        .Y(n2532) );
  AO22X1_HVT U252 ( .A1(n4477), .A2(n4065), .A3(\keys[8][24] ), .A4(n4472), 
        .Y(n2533) );
  AO22X1_HVT U253 ( .A1(n4477), .A2(keyout[25]), .A3(\keys[8][25] ), .A4(n4472), .Y(n2534) );
  AO22X1_HVT U254 ( .A1(n4477), .A2(n4070), .A3(\keys[8][26] ), .A4(n4471), 
        .Y(n2535) );
  AO22X1_HVT U255 ( .A1(n4477), .A2(n4073), .A3(\keys[8][27] ), .A4(n4471), 
        .Y(n2536) );
  AO22X1_HVT U256 ( .A1(n4477), .A2(n4076), .A3(\keys[8][28] ), .A4(n4471), 
        .Y(n2537) );
  AO22X1_HVT U257 ( .A1(n4477), .A2(n4079), .A3(\keys[8][29] ), .A4(n4471), 
        .Y(n2538) );
  AO22X1_HVT U258 ( .A1(n4477), .A2(n4082), .A3(\keys[8][30] ), .A4(n4471), 
        .Y(n2539) );
  AO22X1_HVT U259 ( .A1(n4477), .A2(keyout[31]), .A3(\keys[8][31] ), .A4(n4471), .Y(n2540) );
  AO22X1_HVT U260 ( .A1(n4477), .A2(keyout[32]), .A3(\keys[8][32] ), .A4(n4471), .Y(n2541) );
  AO22X1_HVT U261 ( .A1(n4477), .A2(keyout[33]), .A3(\keys[8][33] ), .A4(n4471), .Y(n2542) );
  AO22X1_HVT U262 ( .A1(n4477), .A2(keyout[34]), .A3(\keys[8][34] ), .A4(n4471), .Y(n2543) );
  AO22X1_HVT U263 ( .A1(n4477), .A2(keyout[35]), .A3(\keys[8][35] ), .A4(n4471), .Y(n2544) );
  AO22X1_HVT U264 ( .A1(n4477), .A2(keyout[36]), .A3(\keys[8][36] ), .A4(n4471), .Y(n2545) );
  AO22X1_HVT U265 ( .A1(n4477), .A2(n3910), .A3(\keys[8][37] ), .A4(n4471), 
        .Y(n2546) );
  AO22X1_HVT U266 ( .A1(n4477), .A2(keyout[38]), .A3(\keys[8][38] ), .A4(n4471), .Y(n2547) );
  AO22X1_HVT U267 ( .A1(n4478), .A2(keyout[39]), .A3(\keys[8][39] ), .A4(n4470), .Y(n2548) );
  AO22X1_HVT U268 ( .A1(n4478), .A2(n3953), .A3(\keys[8][40] ), .A4(n4470), 
        .Y(n2549) );
  AO22X1_HVT U269 ( .A1(n4478), .A2(n3884), .A3(\keys[8][41] ), .A4(n4470), 
        .Y(n2550) );
  AO22X1_HVT U270 ( .A1(n4478), .A2(n3972), .A3(\keys[8][42] ), .A4(n4470), 
        .Y(n2551) );
  AO22X1_HVT U271 ( .A1(n4478), .A2(n3878), .A3(\keys[8][43] ), .A4(n4470), 
        .Y(n2552) );
  AO22X1_HVT U272 ( .A1(n4478), .A2(keyout[44]), .A3(\keys[8][44] ), .A4(n4470), .Y(n2553) );
  AO22X1_HVT U273 ( .A1(n4478), .A2(n3871), .A3(\keys[8][45] ), .A4(n4470), 
        .Y(n2554) );
  AO22X1_HVT U274 ( .A1(n4478), .A2(n3945), .A3(\keys[8][46] ), .A4(n4470), 
        .Y(n2555) );
  AO22X1_HVT U275 ( .A1(n4478), .A2(n3885), .A3(\keys[8][47] ), .A4(n4470), 
        .Y(n2556) );
  AO22X1_HVT U276 ( .A1(n4478), .A2(n1427), .A3(\keys[8][48] ), .A4(n4470), 
        .Y(n2557) );
  AO22X1_HVT U277 ( .A1(n4478), .A2(n14), .A3(\keys[8][49] ), .A4(n4470), .Y(
        n2558) );
  AO22X1_HVT U278 ( .A1(n4478), .A2(n1432), .A3(\keys[8][50] ), .A4(n4470), 
        .Y(n2559) );
  AO22X1_HVT U279 ( .A1(n4478), .A2(n3), .A3(\keys[8][51] ), .A4(n4470), .Y(
        n2560) );
  AO22X1_HVT U280 ( .A1(n4478), .A2(keyout[52]), .A3(\keys[8][52] ), .A4(n4469), .Y(n2561) );
  AO22X1_HVT U281 ( .A1(n4478), .A2(n3874), .A3(\keys[8][53] ), .A4(n4469), 
        .Y(n2562) );
  AO22X1_HVT U282 ( .A1(n4478), .A2(keyout[54]), .A3(\keys[8][54] ), .A4(n4469), .Y(n2563) );
  AO22X1_HVT U283 ( .A1(n4479), .A2(n3866), .A3(\keys[8][55] ), .A4(n4469), 
        .Y(n2564) );
  AO22X1_HVT U284 ( .A1(n4479), .A2(n10), .A3(\keys[8][56] ), .A4(n4469), .Y(
        n2565) );
  AO22X1_HVT U285 ( .A1(n4479), .A2(n4084), .A3(\keys[8][57] ), .A4(n4469), 
        .Y(n2566) );
  AO22X1_HVT U286 ( .A1(n4479), .A2(n4086), .A3(\keys[8][58] ), .A4(n4469), 
        .Y(n2567) );
  AO22X1_HVT U287 ( .A1(n4479), .A2(n4088), .A3(\keys[8][59] ), .A4(n4469), 
        .Y(n2568) );
  AO22X1_HVT U288 ( .A1(n4479), .A2(keyout[60]), .A3(\keys[8][60] ), .A4(n4469), .Y(n2569) );
  AO22X1_HVT U289 ( .A1(n4479), .A2(keyout[61]), .A3(\keys[8][61] ), .A4(n4469), .Y(n2570) );
  AO22X1_HVT U290 ( .A1(n4479), .A2(n3832), .A3(\keys[8][62] ), .A4(n4469), 
        .Y(n2571) );
  AO22X1_HVT U291 ( .A1(n4479), .A2(n3860), .A3(\keys[8][63] ), .A4(n4469), 
        .Y(n2572) );
  AO22X1_HVT U292 ( .A1(n4479), .A2(keyout[64]), .A3(\keys[8][64] ), .A4(n4469), .Y(n2573) );
  AO22X1_HVT U293 ( .A1(n4479), .A2(n3870), .A3(\keys[8][65] ), .A4(n4468), 
        .Y(n2574) );
  AO22X1_HVT U294 ( .A1(n4479), .A2(keyout[66]), .A3(\keys[8][66] ), .A4(n4468), .Y(n2575) );
  AO22X1_HVT U295 ( .A1(n4479), .A2(n3938), .A3(\keys[8][67] ), .A4(n4468), 
        .Y(n2576) );
  AO22X1_HVT U296 ( .A1(n4479), .A2(keyout[68]), .A3(\keys[8][68] ), .A4(n4468), .Y(n2577) );
  AO22X1_HVT U297 ( .A1(n4479), .A2(keyout[69]), .A3(\keys[8][69] ), .A4(n4468), .Y(n2578) );
  AO22X1_HVT U298 ( .A1(n4479), .A2(keyout[70]), .A3(\keys[8][70] ), .A4(n4468), .Y(n2579) );
  AO22X1_HVT U299 ( .A1(n4480), .A2(keyout[71]), .A3(\keys[8][71] ), .A4(n4468), .Y(n2580) );
  AO22X1_HVT U300 ( .A1(n4480), .A2(n3939), .A3(\keys[8][72] ), .A4(n4468), 
        .Y(n2581) );
  AO22X1_HVT U301 ( .A1(n4480), .A2(n3886), .A3(\keys[8][73] ), .A4(n4468), 
        .Y(n2582) );
  AO22X1_HVT U302 ( .A1(n4480), .A2(n3872), .A3(\keys[8][74] ), .A4(n4468), 
        .Y(n2583) );
  AO22X1_HVT U303 ( .A1(n4480), .A2(n3959), .A3(\keys[8][75] ), .A4(n4468), 
        .Y(n2584) );
  AO22X1_HVT U304 ( .A1(n4480), .A2(n3966), .A3(\keys[8][76] ), .A4(n4468), 
        .Y(n2585) );
  AO22X1_HVT U305 ( .A1(n4480), .A2(n3985), .A3(\keys[8][77] ), .A4(n4468), 
        .Y(n2586) );
  AO22X1_HVT U306 ( .A1(n4480), .A2(n3946), .A3(\keys[8][78] ), .A4(n4467), 
        .Y(n2587) );
  AO22X1_HVT U307 ( .A1(n4480), .A2(n3887), .A3(\keys[8][79] ), .A4(n4467), 
        .Y(n2588) );
  AO22X1_HVT U308 ( .A1(n4480), .A2(keyout[80]), .A3(\keys[8][80] ), .A4(n4467), .Y(n2589) );
  AO22X1_HVT U309 ( .A1(n4480), .A2(n3811), .A3(\keys[8][81] ), .A4(n4467), 
        .Y(n2590) );
  AO22X1_HVT U310 ( .A1(n4480), .A2(n3905), .A3(\keys[8][82] ), .A4(n4467), 
        .Y(n2591) );
  AO22X1_HVT U311 ( .A1(n4480), .A2(n3904), .A3(\keys[8][83] ), .A4(n4467), 
        .Y(n2592) );
  AO22X1_HVT U312 ( .A1(n4480), .A2(n1438), .A3(\keys[8][84] ), .A4(n4467), 
        .Y(n2593) );
  AO22X1_HVT U313 ( .A1(n4480), .A2(n2), .A3(\keys[8][85] ), .A4(n4467), .Y(
        n2594) );
  AO22X1_HVT U314 ( .A1(n4480), .A2(n1436), .A3(\keys[8][86] ), .A4(n4467), 
        .Y(n2595) );
  AO22X1_HVT U315 ( .A1(n4481), .A2(n1439), .A3(\keys[8][87] ), .A4(n4467), 
        .Y(n2596) );
  AO22X1_HVT U316 ( .A1(n4481), .A2(n4092), .A3(\keys[8][88] ), .A4(n4467), 
        .Y(n2597) );
  AO22X1_HVT U317 ( .A1(n4481), .A2(n3863), .A3(\keys[8][89] ), .A4(n4467), 
        .Y(n2598) );
  AO22X1_HVT U318 ( .A1(n4481), .A2(keyout[90]), .A3(\keys[8][90] ), .A4(n4467), .Y(n2599) );
  AO22X1_HVT U319 ( .A1(n4481), .A2(n3816), .A3(\keys[8][91] ), .A4(n4466), 
        .Y(n2600) );
  AO22X1_HVT U320 ( .A1(n4481), .A2(n3831), .A3(\keys[8][92] ), .A4(n4466), 
        .Y(n2601) );
  AO22X1_HVT U321 ( .A1(n4481), .A2(keyout[93]), .A3(\keys[8][93] ), .A4(n4466), .Y(n2602) );
  AO22X1_HVT U322 ( .A1(n4481), .A2(n3865), .A3(\keys[8][94] ), .A4(n4466), 
        .Y(n2603) );
  AO22X1_HVT U323 ( .A1(n4481), .A2(n3869), .A3(\keys[8][95] ), .A4(n4466), 
        .Y(n2604) );
  AO22X1_HVT U324 ( .A1(n4481), .A2(keyout[96]), .A3(\keys[8][96] ), .A4(n4466), .Y(n2605) );
  AO22X1_HVT U325 ( .A1(n4481), .A2(keyout[97]), .A3(\keys[8][97] ), .A4(n4466), .Y(n2606) );
  AO22X1_HVT U326 ( .A1(n4481), .A2(keyout[98]), .A3(\keys[8][98] ), .A4(n4466), .Y(n2607) );
  AO22X1_HVT U327 ( .A1(n4481), .A2(keyout[99]), .A3(\keys[8][99] ), .A4(n4466), .Y(n2608) );
  AO22X1_HVT U328 ( .A1(n4481), .A2(keyout[100]), .A3(\keys[8][100] ), .A4(
        n4466), .Y(n2609) );
  AO22X1_HVT U329 ( .A1(n4481), .A2(keyout[101]), .A3(\keys[8][101] ), .A4(
        n4466), .Y(n2610) );
  AO22X1_HVT U330 ( .A1(n4481), .A2(keyout[102]), .A3(\keys[8][102] ), .A4(
        n4466), .Y(n2611) );
  AO22X1_HVT U331 ( .A1(n4482), .A2(keyout[103]), .A3(\keys[8][103] ), .A4(
        n4466), .Y(n2612) );
  AO22X1_HVT U332 ( .A1(n4482), .A2(keyout[104]), .A3(\keys[8][104] ), .A4(
        n4465), .Y(n2613) );
  AO22X1_HVT U333 ( .A1(n4482), .A2(keyout[105]), .A3(\keys[8][105] ), .A4(
        n4465), .Y(n2614) );
  AO22X1_HVT U334 ( .A1(n4482), .A2(n3880), .A3(\keys[8][106] ), .A4(n4465), 
        .Y(n2615) );
  AO22X1_HVT U335 ( .A1(n4482), .A2(n3820), .A3(\keys[8][107] ), .A4(n4465), 
        .Y(n2616) );
  AO22X1_HVT U336 ( .A1(n4482), .A2(n3881), .A3(\keys[8][108] ), .A4(n4465), 
        .Y(n2617) );
  AO22X1_HVT U337 ( .A1(n4482), .A2(n3873), .A3(\keys[8][109] ), .A4(n4465), 
        .Y(n2618) );
  AO22X1_HVT U338 ( .A1(n4482), .A2(keyout[110]), .A3(\keys[8][110] ), .A4(
        n4465), .Y(n2619) );
  AO22X1_HVT U339 ( .A1(n4482), .A2(keyout[111]), .A3(\keys[8][111] ), .A4(
        n4465), .Y(n2620) );
  AO22X1_HVT U340 ( .A1(n4482), .A2(keyout[112]), .A3(\keys[8][112] ), .A4(
        n4465), .Y(n2621) );
  AO22X1_HVT U341 ( .A1(n4482), .A2(keyout[113]), .A3(\keys[8][113] ), .A4(
        n4465), .Y(n2622) );
  AO22X1_HVT U342 ( .A1(n4482), .A2(keyout[114]), .A3(\keys[8][114] ), .A4(
        n4465), .Y(n2623) );
  AO22X1_HVT U343 ( .A1(n4482), .A2(keyout[115]), .A3(\keys[8][115] ), .A4(
        n4465), .Y(n2624) );
  AO22X1_HVT U344 ( .A1(n4482), .A2(keyout[116]), .A3(\keys[8][116] ), .A4(
        n4465), .Y(n2625) );
  AO22X1_HVT U345 ( .A1(n4482), .A2(keyout[117]), .A3(\keys[8][117] ), .A4(
        n4464), .Y(n2626) );
  AO22X1_HVT U346 ( .A1(n4482), .A2(keyout[118]), .A3(\keys[8][118] ), .A4(
        n4464), .Y(n2627) );
  AO22X1_HVT U347 ( .A1(n4483), .A2(keyout[119]), .A3(\keys[8][119] ), .A4(
        n4464), .Y(n2628) );
  AO22X1_HVT U348 ( .A1(n4483), .A2(n4095), .A3(\keys[8][120] ), .A4(n4464), 
        .Y(n2629) );
  AO22X1_HVT U349 ( .A1(n4483), .A2(keyout[121]), .A3(\keys[8][121] ), .A4(
        n4464), .Y(n2630) );
  AO22X1_HVT U350 ( .A1(n4483), .A2(keyout[122]), .A3(\keys[8][122] ), .A4(
        n4464), .Y(n2631) );
  AO22X1_HVT U351 ( .A1(n4483), .A2(n3809), .A3(\keys[8][123] ), .A4(n4464), 
        .Y(n2632) );
  AO22X1_HVT U352 ( .A1(n4483), .A2(n3844), .A3(\keys[8][124] ), .A4(n4464), 
        .Y(n2633) );
  AO22X1_HVT U353 ( .A1(n4483), .A2(keyout[125]), .A3(\keys[8][125] ), .A4(
        n4464), .Y(n2634) );
  AO22X1_HVT U354 ( .A1(n4483), .A2(n4098), .A3(\keys[8][126] ), .A4(n4464), 
        .Y(n2635) );
  AO22X1_HVT U355 ( .A1(n4483), .A2(n4101), .A3(\keys[8][127] ), .A4(n4464), 
        .Y(n2636) );
  AO22X1_HVT U356 ( .A1(n4452), .A2(n3997), .A3(\keys[7][0] ), .A4(n4447), .Y(
        n2637) );
  AO22X1_HVT U357 ( .A1(n4453), .A2(n4000), .A3(\keys[7][1] ), .A4(n4442), .Y(
        n2638) );
  AO22X1_HVT U358 ( .A1(n4453), .A2(keyout[2]), .A3(\keys[7][2] ), .A4(n4442), 
        .Y(n2639) );
  AO22X1_HVT U359 ( .A1(n4453), .A2(n4004), .A3(\keys[7][3] ), .A4(n4442), .Y(
        n2640) );
  AO22X1_HVT U360 ( .A1(n4453), .A2(n4007), .A3(\keys[7][4] ), .A4(n4442), .Y(
        n2641) );
  AO22X1_HVT U361 ( .A1(n4453), .A2(n4010), .A3(\keys[7][5] ), .A4(n4442), .Y(
        n2642) );
  AO22X1_HVT U362 ( .A1(n4453), .A2(n4013), .A3(\keys[7][6] ), .A4(n4442), .Y(
        n2643) );
  AO22X1_HVT U363 ( .A1(n4454), .A2(keyout[7]), .A3(\keys[7][7] ), .A4(n4442), 
        .Y(n2644) );
  AO22X1_HVT U364 ( .A1(n4454), .A2(n4017), .A3(\keys[7][8] ), .A4(n4442), .Y(
        n2645) );
  AO22X1_HVT U365 ( .A1(n4454), .A2(n4020), .A3(\keys[7][9] ), .A4(n4442), .Y(
        n2646) );
  AO22X1_HVT U366 ( .A1(n4454), .A2(n4023), .A3(\keys[7][10] ), .A4(n4442), 
        .Y(n2647) );
  AO22X1_HVT U367 ( .A1(n4454), .A2(n4026), .A3(\keys[7][11] ), .A4(n4443), 
        .Y(n2648) );
  AO22X1_HVT U368 ( .A1(n4454), .A2(n4029), .A3(\keys[7][12] ), .A4(n4443), 
        .Y(n2649) );
  AO22X1_HVT U369 ( .A1(n4454), .A2(n4032), .A3(\keys[7][13] ), .A4(n4443), 
        .Y(n2650) );
  AO22X1_HVT U370 ( .A1(n4454), .A2(n4035), .A3(\keys[7][14] ), .A4(n4443), 
        .Y(n2651) );
  AO22X1_HVT U371 ( .A1(n4454), .A2(n4038), .A3(\keys[7][15] ), .A4(n4443), 
        .Y(n2652) );
  AO22X1_HVT U372 ( .A1(n4454), .A2(n4041), .A3(\keys[7][16] ), .A4(n4443), 
        .Y(n2653) );
  AO22X1_HVT U373 ( .A1(n4454), .A2(n4044), .A3(\keys[7][17] ), .A4(n4443), 
        .Y(n2654) );
  AO22X1_HVT U374 ( .A1(n4454), .A2(n4047), .A3(\keys[7][18] ), .A4(n4443), 
        .Y(n2655) );
  AO22X1_HVT U375 ( .A1(n4454), .A2(n4050), .A3(\keys[7][19] ), .A4(n4443), 
        .Y(n2656) );
  AO22X1_HVT U376 ( .A1(n4454), .A2(n4053), .A3(\keys[7][20] ), .A4(n4443), 
        .Y(n2657) );
  AO22X1_HVT U377 ( .A1(n4454), .A2(n4056), .A3(\keys[7][21] ), .A4(n4443), 
        .Y(n2658) );
  AO22X1_HVT U378 ( .A1(n4454), .A2(n4059), .A3(\keys[7][22] ), .A4(n4443), 
        .Y(n2659) );
  AO22X1_HVT U379 ( .A1(n4455), .A2(n4062), .A3(\keys[7][23] ), .A4(n4443), 
        .Y(n2660) );
  AO22X1_HVT U380 ( .A1(n4455), .A2(n4065), .A3(\keys[7][24] ), .A4(n4444), 
        .Y(n2661) );
  AO22X1_HVT U381 ( .A1(n4455), .A2(keyout[25]), .A3(\keys[7][25] ), .A4(n4444), .Y(n2662) );
  AO22X1_HVT U382 ( .A1(n4455), .A2(n4070), .A3(\keys[7][26] ), .A4(n4444), 
        .Y(n2663) );
  AO22X1_HVT U383 ( .A1(n4455), .A2(n4073), .A3(\keys[7][27] ), .A4(n4444), 
        .Y(n2664) );
  AO22X1_HVT U384 ( .A1(n4455), .A2(n4076), .A3(\keys[7][28] ), .A4(n4444), 
        .Y(n2665) );
  AO22X1_HVT U385 ( .A1(n4455), .A2(n4079), .A3(\keys[7][29] ), .A4(n4444), 
        .Y(n2666) );
  AO22X1_HVT U386 ( .A1(n4455), .A2(n4082), .A3(\keys[7][30] ), .A4(n4444), 
        .Y(n2667) );
  AO22X1_HVT U387 ( .A1(n4455), .A2(keyout[31]), .A3(\keys[7][31] ), .A4(n4444), .Y(n2668) );
  AO22X1_HVT U388 ( .A1(n4455), .A2(keyout[32]), .A3(\keys[7][32] ), .A4(n4444), .Y(n2669) );
  AO22X1_HVT U389 ( .A1(n4455), .A2(keyout[33]), .A3(\keys[7][33] ), .A4(n4444), .Y(n2670) );
  AO22X1_HVT U390 ( .A1(n4455), .A2(keyout[34]), .A3(\keys[7][34] ), .A4(n4444), .Y(n2671) );
  AO22X1_HVT U391 ( .A1(n4455), .A2(keyout[35]), .A3(\keys[7][35] ), .A4(n4444), .Y(n2672) );
  AO22X1_HVT U392 ( .A1(n4455), .A2(keyout[36]), .A3(\keys[7][36] ), .A4(n4444), .Y(n2673) );
  AO22X1_HVT U393 ( .A1(n4455), .A2(n3910), .A3(\keys[7][37] ), .A4(n4445), 
        .Y(n2674) );
  AO22X1_HVT U394 ( .A1(n4455), .A2(keyout[38]), .A3(\keys[7][38] ), .A4(n4445), .Y(n2675) );
  AO22X1_HVT U395 ( .A1(n4456), .A2(keyout[39]), .A3(\keys[7][39] ), .A4(n4445), .Y(n2676) );
  AO22X1_HVT U396 ( .A1(n4456), .A2(n3952), .A3(\keys[7][40] ), .A4(n4445), 
        .Y(n2677) );
  AO22X1_HVT U397 ( .A1(n4456), .A2(n3884), .A3(\keys[7][41] ), .A4(n4445), 
        .Y(n2678) );
  AO22X1_HVT U398 ( .A1(n4456), .A2(n3972), .A3(\keys[7][42] ), .A4(n4445), 
        .Y(n2679) );
  AO22X1_HVT U399 ( .A1(n4456), .A2(n3878), .A3(\keys[7][43] ), .A4(n4445), 
        .Y(n2680) );
  AO22X1_HVT U400 ( .A1(n4456), .A2(n3888), .A3(\keys[7][44] ), .A4(n4445), 
        .Y(n2681) );
  AO22X1_HVT U401 ( .A1(n4456), .A2(n3871), .A3(\keys[7][45] ), .A4(n4445), 
        .Y(n2682) );
  AO22X1_HVT U402 ( .A1(n4456), .A2(n3813), .A3(\keys[7][46] ), .A4(n4445), 
        .Y(n2683) );
  AO22X1_HVT U403 ( .A1(n4456), .A2(n3885), .A3(\keys[7][47] ), .A4(n4445), 
        .Y(n2684) );
  AO22X1_HVT U404 ( .A1(n4456), .A2(n1427), .A3(\keys[7][48] ), .A4(n4445), 
        .Y(n2685) );
  AO22X1_HVT U405 ( .A1(n4456), .A2(n14), .A3(\keys[7][49] ), .A4(n4445), .Y(
        n2686) );
  AO22X1_HVT U406 ( .A1(n4456), .A2(n1432), .A3(\keys[7][50] ), .A4(n4446), 
        .Y(n2687) );
  AO22X1_HVT U407 ( .A1(n4456), .A2(n3), .A3(\keys[7][51] ), .A4(n4446), .Y(
        n2688) );
  AO22X1_HVT U408 ( .A1(n4456), .A2(keyout[52]), .A3(\keys[7][52] ), .A4(n4446), .Y(n2689) );
  AO22X1_HVT U409 ( .A1(n4456), .A2(n3874), .A3(\keys[7][53] ), .A4(n4446), 
        .Y(n2690) );
  AO22X1_HVT U410 ( .A1(n4456), .A2(keyout[54]), .A3(\keys[7][54] ), .A4(n4446), .Y(n2691) );
  AO22X1_HVT U411 ( .A1(n4457), .A2(n3866), .A3(\keys[7][55] ), .A4(n4446), 
        .Y(n2692) );
  AO22X1_HVT U412 ( .A1(n4457), .A2(n10), .A3(\keys[7][56] ), .A4(n4446), .Y(
        n2693) );
  AO22X1_HVT U413 ( .A1(n4457), .A2(n4085), .A3(\keys[7][57] ), .A4(n4446), 
        .Y(n2694) );
  AO22X1_HVT U414 ( .A1(n4457), .A2(n4087), .A3(\keys[7][58] ), .A4(n4446), 
        .Y(n2695) );
  AO22X1_HVT U415 ( .A1(n4457), .A2(n4090), .A3(\keys[7][59] ), .A4(n4446), 
        .Y(n2696) );
  AO22X1_HVT U416 ( .A1(n4457), .A2(keyout[60]), .A3(\keys[7][60] ), .A4(n4446), .Y(n2697) );
  AO22X1_HVT U417 ( .A1(n4457), .A2(n3805), .A3(\keys[7][61] ), .A4(n4446), 
        .Y(n2698) );
  AO22X1_HVT U418 ( .A1(n4457), .A2(n3833), .A3(\keys[7][62] ), .A4(n4446), 
        .Y(n2699) );
  AO22X1_HVT U419 ( .A1(n4457), .A2(n3861), .A3(\keys[7][63] ), .A4(n4447), 
        .Y(n2700) );
  AO22X1_HVT U420 ( .A1(n4457), .A2(keyout[64]), .A3(\keys[7][64] ), .A4(n4447), .Y(n2701) );
  AO22X1_HVT U421 ( .A1(n4457), .A2(n3870), .A3(\keys[7][65] ), .A4(n4447), 
        .Y(n2702) );
  AO22X1_HVT U422 ( .A1(n4457), .A2(keyout[66]), .A3(\keys[7][66] ), .A4(n4447), .Y(n2703) );
  AO22X1_HVT U423 ( .A1(n4457), .A2(n3825), .A3(\keys[7][67] ), .A4(n4447), 
        .Y(n2704) );
  AO22X1_HVT U424 ( .A1(n4457), .A2(keyout[68]), .A3(\keys[7][68] ), .A4(n4447), .Y(n2705) );
  AO22X1_HVT U425 ( .A1(n4457), .A2(keyout[69]), .A3(\keys[7][69] ), .A4(n4447), .Y(n2706) );
  AO22X1_HVT U426 ( .A1(n4457), .A2(keyout[70]), .A3(\keys[7][70] ), .A4(n4447), .Y(n2707) );
  AO22X1_HVT U427 ( .A1(n4458), .A2(keyout[71]), .A3(\keys[7][71] ), .A4(n4447), .Y(n2708) );
  AO22X1_HVT U428 ( .A1(n4458), .A2(n3951), .A3(\keys[7][72] ), .A4(n4447), 
        .Y(n2709) );
  AO22X1_HVT U431 ( .A1(n4458), .A2(n3960), .A3(\keys[7][75] ), .A4(n4448), 
        .Y(n2712) );
  AO22X1_HVT U432 ( .A1(n4458), .A2(n3967), .A3(\keys[7][76] ), .A4(n4448), 
        .Y(n2713) );
  AO22X1_HVT U433 ( .A1(n4458), .A2(n3986), .A3(\keys[7][77] ), .A4(n4448), 
        .Y(n2714) );
  AO22X1_HVT U434 ( .A1(n4458), .A2(n3947), .A3(\keys[7][78] ), .A4(n4448), 
        .Y(n2715) );
  AO22X1_HVT U436 ( .A1(n4458), .A2(n3931), .A3(\keys[7][80] ), .A4(n4448), 
        .Y(n2717) );
  AO22X1_HVT U437 ( .A1(n4458), .A2(keyout[81]), .A3(\keys[7][81] ), .A4(n4448), .Y(n2718) );
  AO22X1_HVT U438 ( .A1(n4458), .A2(n3977), .A3(\keys[7][82] ), .A4(n4448), 
        .Y(n2719) );
  AO22X1_HVT U439 ( .A1(n4458), .A2(n3927), .A3(\keys[7][83] ), .A4(n4448), 
        .Y(n2720) );
  AO22X1_HVT U440 ( .A1(n4458), .A2(keyout[84]), .A3(\keys[7][84] ), .A4(n4448), .Y(n2721) );
  AO22X1_HVT U441 ( .A1(n4458), .A2(n1), .A3(\keys[7][85] ), .A4(n4448), .Y(
        n2722) );
  AO22X1_HVT U442 ( .A1(n4458), .A2(keyout[86]), .A3(\keys[7][86] ), .A4(n4448), .Y(n2723) );
  AO22X1_HVT U443 ( .A1(n4459), .A2(n1440), .A3(\keys[7][87] ), .A4(n4448), 
        .Y(n2724) );
  AO22X1_HVT U444 ( .A1(n4459), .A2(n4092), .A3(\keys[7][88] ), .A4(n4449), 
        .Y(n2725) );
  AO22X1_HVT U445 ( .A1(n4459), .A2(n3863), .A3(\keys[7][89] ), .A4(n4449), 
        .Y(n2726) );
  AO22X1_HVT U446 ( .A1(n4459), .A2(n3949), .A3(\keys[7][90] ), .A4(n4449), 
        .Y(n2727) );
  AO22X1_HVT U447 ( .A1(n4459), .A2(n3816), .A3(\keys[7][91] ), .A4(n4449), 
        .Y(n2728) );
  AO22X1_HVT U448 ( .A1(n4459), .A2(n3831), .A3(\keys[7][92] ), .A4(n4449), 
        .Y(n2729) );
  AO22X1_HVT U449 ( .A1(n4459), .A2(keyout[93]), .A3(\keys[7][93] ), .A4(n4449), .Y(n2730) );
  AO22X1_HVT U450 ( .A1(n4459), .A2(n3865), .A3(\keys[7][94] ), .A4(n4449), 
        .Y(n2731) );
  AO22X1_HVT U451 ( .A1(n4459), .A2(n3869), .A3(\keys[7][95] ), .A4(n4449), 
        .Y(n2732) );
  AO22X1_HVT U452 ( .A1(n4459), .A2(keyout[96]), .A3(\keys[7][96] ), .A4(n4449), .Y(n2733) );
  AO22X1_HVT U453 ( .A1(n4459), .A2(keyout[97]), .A3(\keys[7][97] ), .A4(n4449), .Y(n2734) );
  AO22X1_HVT U454 ( .A1(n4459), .A2(keyout[98]), .A3(\keys[7][98] ), .A4(n4449), .Y(n2735) );
  AO22X1_HVT U455 ( .A1(n4459), .A2(keyout[99]), .A3(\keys[7][99] ), .A4(n4449), .Y(n2736) );
  AO22X1_HVT U456 ( .A1(n4459), .A2(keyout[100]), .A3(\keys[7][100] ), .A4(
        n4449), .Y(n2737) );
  AO22X1_HVT U457 ( .A1(n4459), .A2(keyout[101]), .A3(\keys[7][101] ), .A4(
        n4450), .Y(n2738) );
  AO22X1_HVT U458 ( .A1(n4459), .A2(keyout[102]), .A3(\keys[7][102] ), .A4(
        n4450), .Y(n2739) );
  AO22X1_HVT U459 ( .A1(n4460), .A2(keyout[103]), .A3(\keys[7][103] ), .A4(
        n4450), .Y(n2740) );
  AO22X1_HVT U460 ( .A1(n4460), .A2(n3839), .A3(\keys[7][104] ), .A4(n4450), 
        .Y(n2741) );
  AO22X1_HVT U461 ( .A1(n4460), .A2(keyout[105]), .A3(\keys[7][105] ), .A4(
        n4450), .Y(n2742) );
  AO22X1_HVT U462 ( .A1(n4460), .A2(n3880), .A3(\keys[7][106] ), .A4(n4450), 
        .Y(n2743) );
  AO22X1_HVT U463 ( .A1(n4460), .A2(n3820), .A3(\keys[7][107] ), .A4(n4450), 
        .Y(n2744) );
  AO22X1_HVT U464 ( .A1(n4460), .A2(n3892), .A3(\keys[7][108] ), .A4(n4450), 
        .Y(n2745) );
  AO22X1_HVT U465 ( .A1(n4460), .A2(n3873), .A3(\keys[7][109] ), .A4(n4450), 
        .Y(n2746) );
  AO22X1_HVT U466 ( .A1(n4460), .A2(keyout[110]), .A3(\keys[7][110] ), .A4(
        n4450), .Y(n2747) );
  AO22X1_HVT U467 ( .A1(n4460), .A2(keyout[111]), .A3(\keys[7][111] ), .A4(
        n4450), .Y(n2748) );
  AO22X1_HVT U468 ( .A1(n4460), .A2(keyout[112]), .A3(\keys[7][112] ), .A4(
        n4450), .Y(n2749) );
  AO22X1_HVT U469 ( .A1(n4460), .A2(keyout[113]), .A3(\keys[7][113] ), .A4(
        n4450), .Y(n2750) );
  AO22X1_HVT U470 ( .A1(n4460), .A2(keyout[114]), .A3(\keys[7][114] ), .A4(
        n4451), .Y(n2751) );
  AO22X1_HVT U471 ( .A1(n4460), .A2(n3915), .A3(\keys[7][115] ), .A4(n4451), 
        .Y(n2752) );
  AO22X1_HVT U472 ( .A1(n4460), .A2(keyout[116]), .A3(\keys[7][116] ), .A4(
        n4451), .Y(n2753) );
  AO22X1_HVT U473 ( .A1(n4460), .A2(keyout[117]), .A3(\keys[7][117] ), .A4(
        n4451), .Y(n2754) );
  AO22X1_HVT U474 ( .A1(n4460), .A2(keyout[118]), .A3(\keys[7][118] ), .A4(
        n4451), .Y(n2755) );
  AO22X1_HVT U475 ( .A1(n4461), .A2(keyout[119]), .A3(\keys[7][119] ), .A4(
        n4451), .Y(n2756) );
  AO22X1_HVT U476 ( .A1(n4461), .A2(n4095), .A3(\keys[7][120] ), .A4(n4451), 
        .Y(n2757) );
  AO22X1_HVT U477 ( .A1(n4461), .A2(n3829), .A3(\keys[7][121] ), .A4(n4451), 
        .Y(n2758) );
  AO22X1_HVT U478 ( .A1(n4461), .A2(n3803), .A3(\keys[7][122] ), .A4(n4451), 
        .Y(n2759) );
  AO22X1_HVT U479 ( .A1(n4461), .A2(n3817), .A3(\keys[7][123] ), .A4(n4451), 
        .Y(n2760) );
  AO22X1_HVT U480 ( .A1(n4461), .A2(n3845), .A3(\keys[7][124] ), .A4(n4451), 
        .Y(n2761) );
  AO22X1_HVT U481 ( .A1(n4461), .A2(n3823), .A3(\keys[7][125] ), .A4(n4451), 
        .Y(n2762) );
  AO22X1_HVT U482 ( .A1(n4461), .A2(n4098), .A3(\keys[7][126] ), .A4(n4451), 
        .Y(n2763) );
  AO22X1_HVT U483 ( .A1(n4461), .A2(n4101), .A3(\keys[7][127] ), .A4(n4442), 
        .Y(n2764) );
  AO22X1_HVT U484 ( .A1(n4430), .A2(n3999), .A3(\keys[6][0] ), .A4(n4429), .Y(
        n2765) );
  AO22X1_HVT U485 ( .A1(n4431), .A2(n4002), .A3(\keys[6][1] ), .A4(n4429), .Y(
        n2766) );
  AO22X1_HVT U486 ( .A1(n4431), .A2(n4003), .A3(\keys[6][2] ), .A4(n4429), .Y(
        n2767) );
  AO22X1_HVT U487 ( .A1(n4431), .A2(n4006), .A3(\keys[6][3] ), .A4(n4429), .Y(
        n2768) );
  AO22X1_HVT U488 ( .A1(n4431), .A2(n4009), .A3(\keys[6][4] ), .A4(n4429), .Y(
        n2769) );
  AO22X1_HVT U489 ( .A1(n4431), .A2(n4012), .A3(\keys[6][5] ), .A4(n4429), .Y(
        n2770) );
  AO22X1_HVT U490 ( .A1(n4431), .A2(n4015), .A3(\keys[6][6] ), .A4(n4429), .Y(
        n2771) );
  AO22X1_HVT U491 ( .A1(n4432), .A2(n4016), .A3(\keys[6][7] ), .A4(n4429), .Y(
        n2772) );
  AO22X1_HVT U492 ( .A1(n4432), .A2(n4019), .A3(\keys[6][8] ), .A4(n4429), .Y(
        n2773) );
  AO22X1_HVT U493 ( .A1(n4432), .A2(n4022), .A3(\keys[6][9] ), .A4(n4429), .Y(
        n2774) );
  AO22X1_HVT U494 ( .A1(n4432), .A2(n4025), .A3(\keys[6][10] ), .A4(n4429), 
        .Y(n2775) );
  AO22X1_HVT U495 ( .A1(n4432), .A2(n4028), .A3(\keys[6][11] ), .A4(n4429), 
        .Y(n2776) );
  AO22X1_HVT U496 ( .A1(n4432), .A2(n4031), .A3(\keys[6][12] ), .A4(n4428), 
        .Y(n2777) );
  AO22X1_HVT U497 ( .A1(n4432), .A2(n4034), .A3(\keys[6][13] ), .A4(n4428), 
        .Y(n2778) );
  AO22X1_HVT U498 ( .A1(n4432), .A2(n4037), .A3(\keys[6][14] ), .A4(n4428), 
        .Y(n2779) );
  AO22X1_HVT U499 ( .A1(n4432), .A2(n4040), .A3(\keys[6][15] ), .A4(n4428), 
        .Y(n2780) );
  AO22X1_HVT U500 ( .A1(n4432), .A2(n4043), .A3(\keys[6][16] ), .A4(n4428), 
        .Y(n2781) );
  AO22X1_HVT U501 ( .A1(n4432), .A2(n4046), .A3(\keys[6][17] ), .A4(n4428), 
        .Y(n2782) );
  AO22X1_HVT U502 ( .A1(n4432), .A2(n4049), .A3(\keys[6][18] ), .A4(n4428), 
        .Y(n2783) );
  AO22X1_HVT U503 ( .A1(n4432), .A2(n4052), .A3(\keys[6][19] ), .A4(n4428), 
        .Y(n2784) );
  AO22X1_HVT U504 ( .A1(n4432), .A2(n4055), .A3(\keys[6][20] ), .A4(n4428), 
        .Y(n2785) );
  AO22X1_HVT U505 ( .A1(n4432), .A2(n4058), .A3(\keys[6][21] ), .A4(n4428), 
        .Y(n2786) );
  AO22X1_HVT U506 ( .A1(n4432), .A2(n4061), .A3(\keys[6][22] ), .A4(n4428), 
        .Y(n2787) );
  AO22X1_HVT U507 ( .A1(n4433), .A2(n4064), .A3(\keys[6][23] ), .A4(n4428), 
        .Y(n2788) );
  AO22X1_HVT U508 ( .A1(n4433), .A2(n4067), .A3(\keys[6][24] ), .A4(n4428), 
        .Y(n2789) );
  AO22X1_HVT U509 ( .A1(n4433), .A2(n4069), .A3(\keys[6][25] ), .A4(n4427), 
        .Y(n2790) );
  AO22X1_HVT U510 ( .A1(n4433), .A2(n4072), .A3(\keys[6][26] ), .A4(n4427), 
        .Y(n2791) );
  AO22X1_HVT U511 ( .A1(n4433), .A2(n4075), .A3(\keys[6][27] ), .A4(n4427), 
        .Y(n2792) );
  AO22X1_HVT U512 ( .A1(n4433), .A2(n4078), .A3(\keys[6][28] ), .A4(n4427), 
        .Y(n2793) );
  AO22X1_HVT U513 ( .A1(n4433), .A2(n4081), .A3(\keys[6][29] ), .A4(n4427), 
        .Y(n2794) );
  AO22X1_HVT U514 ( .A1(n4433), .A2(n4083), .A3(\keys[6][30] ), .A4(n4427), 
        .Y(n2795) );
  AO22X1_HVT U515 ( .A1(n4433), .A2(keyout[31]), .A3(\keys[6][31] ), .A4(n4427), .Y(n2796) );
  AO22X1_HVT U516 ( .A1(n4433), .A2(keyout[32]), .A3(\keys[6][32] ), .A4(n4427), .Y(n2797) );
  AO22X1_HVT U517 ( .A1(n4433), .A2(keyout[33]), .A3(\keys[6][33] ), .A4(n4427), .Y(n2798) );
  AO22X1_HVT U518 ( .A1(n4433), .A2(keyout[34]), .A3(\keys[6][34] ), .A4(n4427), .Y(n2799) );
  AO22X1_HVT U519 ( .A1(n4433), .A2(keyout[35]), .A3(\keys[6][35] ), .A4(n4427), .Y(n2800) );
  AO22X1_HVT U520 ( .A1(n4433), .A2(keyout[36]), .A3(\keys[6][36] ), .A4(n4427), .Y(n2801) );
  AO22X1_HVT U521 ( .A1(n4433), .A2(n3910), .A3(\keys[6][37] ), .A4(n4427), 
        .Y(n2802) );
  AO22X1_HVT U522 ( .A1(n4433), .A2(keyout[38]), .A3(\keys[6][38] ), .A4(n4426), .Y(n2803) );
  AO22X1_HVT U523 ( .A1(n4434), .A2(keyout[39]), .A3(\keys[6][39] ), .A4(n4426), .Y(n2804) );
  AO22X1_HVT U524 ( .A1(n4434), .A2(n3953), .A3(\keys[6][40] ), .A4(n4426), 
        .Y(n2805) );
  AO22X1_HVT U525 ( .A1(n4434), .A2(n3854), .A3(\keys[6][41] ), .A4(n4426), 
        .Y(n2806) );
  AO22X1_HVT U526 ( .A1(n3972), .A2(n4434), .A3(\keys[6][42] ), .A4(n4426), 
        .Y(n2807) );
  AO22X1_HVT U527 ( .A1(n4434), .A2(n3890), .A3(\keys[6][43] ), .A4(n4426), 
        .Y(n2808) );
  AO22X1_HVT U528 ( .A1(n4434), .A2(n3888), .A3(\keys[6][44] ), .A4(n4426), 
        .Y(n2809) );
  AO22X1_HVT U529 ( .A1(n4434), .A2(n3871), .A3(\keys[6][45] ), .A4(n4426), 
        .Y(n2810) );
  AO22X1_HVT U530 ( .A1(n4434), .A2(n3945), .A3(\keys[6][46] ), .A4(n4426), 
        .Y(n2811) );
  AO22X1_HVT U531 ( .A1(n4434), .A2(n3850), .A3(\keys[6][47] ), .A4(n4426), 
        .Y(n2812) );
  AO22X1_HVT U532 ( .A1(n4434), .A2(n1427), .A3(\keys[6][48] ), .A4(n4426), 
        .Y(n2813) );
  AO22X1_HVT U533 ( .A1(n4434), .A2(n14), .A3(\keys[6][49] ), .A4(n4426), .Y(
        n2814) );
  AO22X1_HVT U534 ( .A1(n4434), .A2(n1432), .A3(\keys[6][50] ), .A4(n4426), 
        .Y(n2815) );
  AO22X1_HVT U535 ( .A1(n4434), .A2(n3), .A3(\keys[6][51] ), .A4(n4425), .Y(
        n2816) );
  AO22X1_HVT U536 ( .A1(n4434), .A2(keyout[52]), .A3(\keys[6][52] ), .A4(n4425), .Y(n2817) );
  AO22X1_HVT U537 ( .A1(n4434), .A2(keyout[53]), .A3(\keys[6][53] ), .A4(n4425), .Y(n2818) );
  AO22X1_HVT U538 ( .A1(n4434), .A2(keyout[54]), .A3(\keys[6][54] ), .A4(n4425), .Y(n2819) );
  AO22X1_HVT U539 ( .A1(n4435), .A2(n3866), .A3(\keys[6][55] ), .A4(n4425), 
        .Y(n2820) );
  AO22X1_HVT U540 ( .A1(n4435), .A2(n10), .A3(\keys[6][56] ), .A4(n4425), .Y(
        n2821) );
  AO22X1_HVT U541 ( .A1(n4435), .A2(n4085), .A3(\keys[6][57] ), .A4(n4425), 
        .Y(n2822) );
  AO22X1_HVT U542 ( .A1(n4435), .A2(n4087), .A3(\keys[6][58] ), .A4(n4425), 
        .Y(n2823) );
  AO22X1_HVT U543 ( .A1(n4435), .A2(n4089), .A3(\keys[6][59] ), .A4(n4425), 
        .Y(n2824) );
  AO22X1_HVT U544 ( .A1(n4435), .A2(keyout[60]), .A3(\keys[6][60] ), .A4(n4425), .Y(n2825) );
  AO22X1_HVT U545 ( .A1(n4435), .A2(n3805), .A3(\keys[6][61] ), .A4(n4425), 
        .Y(n2826) );
  AO22X1_HVT U546 ( .A1(n4435), .A2(n3832), .A3(\keys[6][62] ), .A4(n4425), 
        .Y(n2827) );
  AO22X1_HVT U547 ( .A1(n4435), .A2(n3860), .A3(\keys[6][63] ), .A4(n4425), 
        .Y(n2828) );
  AO22X1_HVT U548 ( .A1(n4435), .A2(keyout[64]), .A3(\keys[6][64] ), .A4(n4424), .Y(n2829) );
  AO22X1_HVT U549 ( .A1(n4435), .A2(n3870), .A3(\keys[6][65] ), .A4(n4424), 
        .Y(n2830) );
  AO22X1_HVT U550 ( .A1(n4435), .A2(keyout[66]), .A3(\keys[6][66] ), .A4(n4424), .Y(n2831) );
  AO22X1_HVT U551 ( .A1(n4435), .A2(n3825), .A3(\keys[6][67] ), .A4(n4424), 
        .Y(n2832) );
  AO22X1_HVT U552 ( .A1(n4435), .A2(keyout[68]), .A3(\keys[6][68] ), .A4(n4424), .Y(n2833) );
  AO22X1_HVT U553 ( .A1(n4435), .A2(keyout[69]), .A3(\keys[6][69] ), .A4(n4424), .Y(n2834) );
  AO22X1_HVT U554 ( .A1(n4435), .A2(keyout[70]), .A3(\keys[6][70] ), .A4(n4424), .Y(n2835) );
  AO22X1_HVT U555 ( .A1(n4436), .A2(keyout[71]), .A3(\keys[6][71] ), .A4(n4424), .Y(n2836) );
  AO22X1_HVT U556 ( .A1(n4436), .A2(n3951), .A3(\keys[6][72] ), .A4(n4424), 
        .Y(n2837) );
  AO22X1_HVT U557 ( .A1(n4436), .A2(n3896), .A3(\keys[6][73] ), .A4(n4424), 
        .Y(n2838) );
  AO22X1_HVT U558 ( .A1(n4436), .A2(n3979), .A3(\keys[6][74] ), .A4(n4424), 
        .Y(n2839) );
  AO22X1_HVT U559 ( .A1(n4436), .A2(n3959), .A3(\keys[6][75] ), .A4(n4424), 
        .Y(n2840) );
  AO22X1_HVT U560 ( .A1(n4436), .A2(n3966), .A3(\keys[6][76] ), .A4(n4424), 
        .Y(n2841) );
  AO22X1_HVT U561 ( .A1(n4436), .A2(n3985), .A3(\keys[6][77] ), .A4(n4423), 
        .Y(n2842) );
  AO22X1_HVT U562 ( .A1(n4436), .A2(n3946), .A3(\keys[6][78] ), .A4(n4423), 
        .Y(n2843) );
  AO22X1_HVT U563 ( .A1(n4436), .A2(n3898), .A3(\keys[6][79] ), .A4(n4423), 
        .Y(n2844) );
  AO22X1_HVT U564 ( .A1(n4436), .A2(n3931), .A3(\keys[6][80] ), .A4(n4423), 
        .Y(n2845) );
  AO22X1_HVT U565 ( .A1(n4436), .A2(n3811), .A3(\keys[6][81] ), .A4(n4423), 
        .Y(n2846) );
  AO22X1_HVT U566 ( .A1(n4436), .A2(n3977), .A3(\keys[6][82] ), .A4(n4423), 
        .Y(n2847) );
  AO22X1_HVT U567 ( .A1(n4436), .A2(n3927), .A3(\keys[6][83] ), .A4(n4423), 
        .Y(n2848) );
  AO22X1_HVT U568 ( .A1(n4436), .A2(n1438), .A3(\keys[6][84] ), .A4(n4423), 
        .Y(n2849) );
  AO22X1_HVT U569 ( .A1(n4436), .A2(n2), .A3(\keys[6][85] ), .A4(n4423), .Y(
        n2850) );
  AO22X1_HVT U570 ( .A1(n4436), .A2(n1436), .A3(\keys[6][86] ), .A4(n4423), 
        .Y(n2851) );
  AO22X1_HVT U571 ( .A1(n4437), .A2(n1440), .A3(\keys[6][87] ), .A4(n4423), 
        .Y(n2852) );
  AO22X1_HVT U572 ( .A1(n4437), .A2(n4092), .A3(\keys[6][88] ), .A4(n4423), 
        .Y(n2853) );
  AO22X1_HVT U573 ( .A1(n4437), .A2(n3863), .A3(\keys[6][89] ), .A4(n4423), 
        .Y(n2854) );
  AO22X1_HVT U574 ( .A1(n4437), .A2(n3949), .A3(\keys[6][90] ), .A4(n4422), 
        .Y(n2855) );
  AO22X1_HVT U575 ( .A1(n4437), .A2(n4), .A3(\keys[6][91] ), .A4(n4422), .Y(
        n2856) );
  AO22X1_HVT U576 ( .A1(n4437), .A2(keyout[92]), .A3(\keys[6][92] ), .A4(n4422), .Y(n2857) );
  AO22X1_HVT U577 ( .A1(n4437), .A2(keyout[93]), .A3(\keys[6][93] ), .A4(n4422), .Y(n2858) );
  AO22X1_HVT U578 ( .A1(n4437), .A2(n3835), .A3(\keys[6][94] ), .A4(n4422), 
        .Y(n2859) );
  AO22X1_HVT U579 ( .A1(n4437), .A2(n3869), .A3(\keys[6][95] ), .A4(n4422), 
        .Y(n2860) );
  AO22X1_HVT U580 ( .A1(n4437), .A2(keyout[96]), .A3(\keys[6][96] ), .A4(n4422), .Y(n2861) );
  AO22X1_HVT U581 ( .A1(n4437), .A2(keyout[97]), .A3(\keys[6][97] ), .A4(n4422), .Y(n2862) );
  AO22X1_HVT U582 ( .A1(n4437), .A2(keyout[98]), .A3(\keys[6][98] ), .A4(n4422), .Y(n2863) );
  AO22X1_HVT U583 ( .A1(n4437), .A2(keyout[99]), .A3(\keys[6][99] ), .A4(n4422), .Y(n2864) );
  AO22X1_HVT U584 ( .A1(n4437), .A2(keyout[100]), .A3(\keys[6][100] ), .A4(
        n4422), .Y(n2865) );
  AO22X1_HVT U585 ( .A1(n4437), .A2(keyout[101]), .A3(\keys[6][101] ), .A4(
        n4422), .Y(n2866) );
  AO22X1_HVT U586 ( .A1(n4437), .A2(keyout[102]), .A3(\keys[6][102] ), .A4(
        n4422), .Y(n2867) );
  AO22X1_HVT U587 ( .A1(n4438), .A2(keyout[103]), .A3(\keys[6][103] ), .A4(
        n4421), .Y(n2868) );
  AO22X1_HVT U588 ( .A1(n4438), .A2(keyout[104]), .A3(\keys[6][104] ), .A4(
        n4421), .Y(n2869) );
  AO22X1_HVT U589 ( .A1(n4438), .A2(keyout[105]), .A3(\keys[6][105] ), .A4(
        n4421), .Y(n2870) );
  AO22X1_HVT U590 ( .A1(n4438), .A2(keyout[106]), .A3(\keys[6][106] ), .A4(
        n4421), .Y(n2871) );
  AO22X1_HVT U591 ( .A1(n4438), .A2(keyout[107]), .A3(\keys[6][107] ), .A4(
        n4421), .Y(n2872) );
  AO22X1_HVT U593 ( .A1(n4438), .A2(keyout[109]), .A3(\keys[6][109] ), .A4(
        n4421), .Y(n2874) );
  AO22X1_HVT U594 ( .A1(n4438), .A2(keyout[110]), .A3(\keys[6][110] ), .A4(
        n4421), .Y(n2875) );
  AO22X1_HVT U595 ( .A1(n4438), .A2(keyout[111]), .A3(\keys[6][111] ), .A4(
        n4421), .Y(n2876) );
  AO22X1_HVT U596 ( .A1(n4438), .A2(keyout[112]), .A3(\keys[6][112] ), .A4(
        n4421), .Y(n2877) );
  AO22X1_HVT U597 ( .A1(n4438), .A2(keyout[113]), .A3(\keys[6][113] ), .A4(
        n4421), .Y(n2878) );
  AO22X1_HVT U598 ( .A1(n4438), .A2(keyout[114]), .A3(\keys[6][114] ), .A4(
        n4421), .Y(n2879) );
  AO22X1_HVT U599 ( .A1(n4438), .A2(n3915), .A3(\keys[6][115] ), .A4(n4421), 
        .Y(n2880) );
  AO22X1_HVT U600 ( .A1(n4438), .A2(keyout[116]), .A3(\keys[6][116] ), .A4(
        n4420), .Y(n2881) );
  AO22X1_HVT U601 ( .A1(n4438), .A2(keyout[117]), .A3(\keys[6][117] ), .A4(
        n4420), .Y(n2882) );
  AO22X1_HVT U602 ( .A1(n4438), .A2(keyout[118]), .A3(\keys[6][118] ), .A4(
        n4420), .Y(n2883) );
  AO22X1_HVT U603 ( .A1(n4439), .A2(keyout[119]), .A3(\keys[6][119] ), .A4(
        n4420), .Y(n2884) );
  AO22X1_HVT U604 ( .A1(n4439), .A2(n4095), .A3(\keys[6][120] ), .A4(n4420), 
        .Y(n2885) );
  AO22X1_HVT U605 ( .A1(n4439), .A2(keyout[121]), .A3(\keys[6][121] ), .A4(
        n4420), .Y(n2886) );
  AO22X1_HVT U606 ( .A1(n4439), .A2(keyout[122]), .A3(\keys[6][122] ), .A4(
        n4420), .Y(n2887) );
  AO22X1_HVT U607 ( .A1(n4439), .A2(n3809), .A3(\keys[6][123] ), .A4(n4420), 
        .Y(n2888) );
  AO22X1_HVT U608 ( .A1(n4439), .A2(n3844), .A3(\keys[6][124] ), .A4(n4420), 
        .Y(n2889) );
  AO22X1_HVT U609 ( .A1(n4439), .A2(keyout[125]), .A3(\keys[6][125] ), .A4(
        n4420), .Y(n2890) );
  AO22X1_HVT U610 ( .A1(n4439), .A2(n4098), .A3(\keys[6][126] ), .A4(n4420), 
        .Y(n2891) );
  AO22X1_HVT U611 ( .A1(n4439), .A2(n4101), .A3(\keys[6][127] ), .A4(n4420), 
        .Y(n2892) );
  AO22X1_HVT U612 ( .A1(n4408), .A2(n3998), .A3(\keys[5][0] ), .A4(n4402), .Y(
        n2893) );
  AO22X1_HVT U613 ( .A1(n4409), .A2(n4001), .A3(\keys[5][1] ), .A4(n4397), .Y(
        n2894) );
  AO22X1_HVT U614 ( .A1(n4409), .A2(n4003), .A3(\keys[5][2] ), .A4(n4397), .Y(
        n2895) );
  AO22X1_HVT U615 ( .A1(n4409), .A2(n4005), .A3(\keys[5][3] ), .A4(n4397), .Y(
        n2896) );
  AO22X1_HVT U616 ( .A1(n4410), .A2(n4008), .A3(\keys[5][4] ), .A4(n4397), .Y(
        n2897) );
  AO22X1_HVT U617 ( .A1(n4410), .A2(n4011), .A3(\keys[5][5] ), .A4(n4397), .Y(
        n2898) );
  AO22X1_HVT U618 ( .A1(n4410), .A2(n4014), .A3(\keys[5][6] ), .A4(n4397), .Y(
        n2899) );
  AO22X1_HVT U619 ( .A1(n4410), .A2(n4016), .A3(\keys[5][7] ), .A4(n4397), .Y(
        n2900) );
  AO22X1_HVT U620 ( .A1(n4410), .A2(n4018), .A3(\keys[5][8] ), .A4(n4397), .Y(
        n2901) );
  AO22X1_HVT U621 ( .A1(n4410), .A2(n4021), .A3(\keys[5][9] ), .A4(n4397), .Y(
        n2902) );
  AO22X1_HVT U622 ( .A1(n4410), .A2(n4024), .A3(\keys[5][10] ), .A4(n4397), 
        .Y(n2903) );
  AO22X1_HVT U623 ( .A1(n4410), .A2(n4027), .A3(\keys[5][11] ), .A4(n4397), 
        .Y(n2904) );
  AO22X1_HVT U624 ( .A1(n4410), .A2(n4030), .A3(\keys[5][12] ), .A4(n4397), 
        .Y(n2905) );
  AO22X1_HVT U625 ( .A1(n4410), .A2(n4033), .A3(\keys[5][13] ), .A4(n4398), 
        .Y(n2906) );
  AO22X1_HVT U626 ( .A1(n4410), .A2(n4036), .A3(\keys[5][14] ), .A4(n4398), 
        .Y(n2907) );
  AO22X1_HVT U627 ( .A1(n4410), .A2(n4039), .A3(\keys[5][15] ), .A4(n4398), 
        .Y(n2908) );
  AO22X1_HVT U628 ( .A1(n4410), .A2(n4042), .A3(\keys[5][16] ), .A4(n4398), 
        .Y(n2909) );
  AO22X1_HVT U629 ( .A1(n4410), .A2(n4045), .A3(\keys[5][17] ), .A4(n4398), 
        .Y(n2910) );
  AO22X1_HVT U630 ( .A1(n4410), .A2(n4048), .A3(\keys[5][18] ), .A4(n4398), 
        .Y(n2911) );
  AO22X1_HVT U631 ( .A1(n4410), .A2(n4051), .A3(\keys[5][19] ), .A4(n4398), 
        .Y(n2912) );
  AO22X1_HVT U632 ( .A1(n4411), .A2(n4054), .A3(\keys[5][20] ), .A4(n4398), 
        .Y(n2913) );
  AO22X1_HVT U633 ( .A1(n4411), .A2(n4057), .A3(\keys[5][21] ), .A4(n4398), 
        .Y(n2914) );
  AO22X1_HVT U634 ( .A1(n4411), .A2(n4060), .A3(\keys[5][22] ), .A4(n4398), 
        .Y(n2915) );
  AO22X1_HVT U635 ( .A1(n4411), .A2(n4063), .A3(\keys[5][23] ), .A4(n4398), 
        .Y(n2916) );
  AO22X1_HVT U636 ( .A1(n4411), .A2(n4066), .A3(\keys[5][24] ), .A4(n4398), 
        .Y(n2917) );
  AO22X1_HVT U637 ( .A1(n4411), .A2(n4068), .A3(\keys[5][25] ), .A4(n4399), 
        .Y(n2918) );
  AO22X1_HVT U638 ( .A1(n4411), .A2(n4071), .A3(\keys[5][26] ), .A4(n4399), 
        .Y(n2919) );
  AO22X1_HVT U639 ( .A1(n4411), .A2(n4074), .A3(\keys[5][27] ), .A4(n4399), 
        .Y(n2920) );
  AO22X1_HVT U640 ( .A1(n4411), .A2(n4077), .A3(\keys[5][28] ), .A4(n4399), 
        .Y(n2921) );
  AO22X1_HVT U641 ( .A1(n4411), .A2(n4080), .A3(\keys[5][29] ), .A4(n4399), 
        .Y(n2922) );
  AO22X1_HVT U642 ( .A1(n4411), .A2(n4083), .A3(\keys[5][30] ), .A4(n4399), 
        .Y(n2923) );
  AO22X1_HVT U643 ( .A1(n4411), .A2(n3852), .A3(\keys[5][31] ), .A4(n4399), 
        .Y(n2924) );
  AO22X1_HVT U644 ( .A1(n4411), .A2(keyout[32]), .A3(\keys[5][32] ), .A4(n4399), .Y(n2925) );
  AO22X1_HVT U645 ( .A1(n4411), .A2(keyout[33]), .A3(\keys[5][33] ), .A4(n4399), .Y(n2926) );
  AO22X1_HVT U646 ( .A1(n4411), .A2(keyout[34]), .A3(\keys[5][34] ), .A4(n4399), .Y(n2927) );
  AO22X1_HVT U647 ( .A1(n4411), .A2(keyout[35]), .A3(\keys[5][35] ), .A4(n4399), .Y(n2928) );
  AO22X1_HVT U648 ( .A1(n4412), .A2(keyout[36]), .A3(\keys[5][36] ), .A4(n4399), .Y(n2929) );
  AO22X1_HVT U649 ( .A1(n4412), .A2(n3911), .A3(\keys[5][37] ), .A4(n4400), 
        .Y(n2930) );
  AO22X1_HVT U650 ( .A1(n4412), .A2(keyout[38]), .A3(\keys[5][38] ), .A4(n4400), .Y(n2931) );
  AO22X1_HVT U651 ( .A1(n4412), .A2(keyout[39]), .A3(\keys[5][39] ), .A4(n4400), .Y(n2932) );
  AO22X1_HVT U652 ( .A1(n4412), .A2(n3952), .A3(\keys[5][40] ), .A4(n4400), 
        .Y(n2933) );
  AO22X1_HVT U653 ( .A1(n4412), .A2(n3884), .A3(\keys[5][41] ), .A4(n4400), 
        .Y(n2934) );
  AO22X1_HVT U654 ( .A1(n4412), .A2(n3973), .A3(\keys[5][42] ), .A4(n4400), 
        .Y(n2935) );
  AO22X1_HVT U655 ( .A1(n4412), .A2(n3878), .A3(\keys[5][43] ), .A4(n4400), 
        .Y(n2936) );
  AO22X1_HVT U656 ( .A1(n4412), .A2(n3888), .A3(\keys[5][44] ), .A4(n4400), 
        .Y(n2937) );
  AO22X1_HVT U657 ( .A1(n4412), .A2(n3871), .A3(\keys[5][45] ), .A4(n4400), 
        .Y(n2938) );
  AO22X1_HVT U658 ( .A1(n4412), .A2(n3813), .A3(\keys[5][46] ), .A4(n4400), 
        .Y(n2939) );
  AO22X1_HVT U659 ( .A1(n4412), .A2(n3885), .A3(\keys[5][47] ), .A4(n4400), 
        .Y(n2940) );
  AO22X1_HVT U660 ( .A1(n4412), .A2(n1427), .A3(\keys[5][48] ), .A4(n4400), 
        .Y(n2941) );
  AO22X1_HVT U661 ( .A1(n4412), .A2(n1429), .A3(\keys[5][49] ), .A4(n4401), 
        .Y(n2942) );
  AO22X1_HVT U662 ( .A1(n4412), .A2(n1432), .A3(\keys[5][50] ), .A4(n4401), 
        .Y(n2943) );
  AO22X1_HVT U663 ( .A1(n4412), .A2(n3937), .A3(\keys[5][51] ), .A4(n4401), 
        .Y(n2944) );
  AO22X1_HVT U664 ( .A1(n4413), .A2(keyout[52]), .A3(\keys[5][52] ), .A4(n4401), .Y(n2945) );
  AO22X1_HVT U665 ( .A1(n4413), .A2(n3920), .A3(\keys[5][53] ), .A4(n4401), 
        .Y(n2946) );
  AO22X1_HVT U666 ( .A1(n4413), .A2(keyout[54]), .A3(\keys[5][54] ), .A4(n4401), .Y(n2947) );
  AO22X1_HVT U668 ( .A1(n4413), .A2(n3941), .A3(\keys[5][56] ), .A4(n4401), 
        .Y(n2949) );
  AO22X1_HVT U669 ( .A1(n4413), .A2(keyout[57]), .A3(\keys[5][57] ), .A4(n4401), .Y(n2950) );
  AO22X1_HVT U670 ( .A1(n4413), .A2(keyout[58]), .A3(\keys[5][58] ), .A4(n4401), .Y(n2951) );
  AO22X1_HVT U671 ( .A1(n4413), .A2(n4089), .A3(\keys[5][59] ), .A4(n4401), 
        .Y(n2952) );
  AO22X1_HVT U672 ( .A1(n4413), .A2(n3943), .A3(\keys[5][60] ), .A4(n4401), 
        .Y(n2953) );
  AO22X1_HVT U673 ( .A1(n4413), .A2(keyout[61]), .A3(\keys[5][61] ), .A4(n4402), .Y(n2954) );
  AO22X1_HVT U674 ( .A1(n4413), .A2(n3833), .A3(\keys[5][62] ), .A4(n4402), 
        .Y(n2955) );
  AO22X1_HVT U675 ( .A1(n4413), .A2(n3859), .A3(\keys[5][63] ), .A4(n4402), 
        .Y(n2956) );
  AO22X1_HVT U676 ( .A1(n4413), .A2(keyout[64]), .A3(\keys[5][64] ), .A4(n4402), .Y(n2957) );
  AO22X1_HVT U677 ( .A1(n4413), .A2(n3883), .A3(\keys[5][65] ), .A4(n4402), 
        .Y(n2958) );
  AO22X1_HVT U678 ( .A1(n4413), .A2(n3914), .A3(\keys[5][66] ), .A4(n4402), 
        .Y(n2959) );
  AO22X1_HVT U679 ( .A1(n4413), .A2(n3938), .A3(\keys[5][67] ), .A4(n4402), 
        .Y(n2960) );
  AO22X1_HVT U680 ( .A1(n4414), .A2(keyout[68]), .A3(\keys[5][68] ), .A4(n4402), .Y(n2961) );
  AO22X1_HVT U681 ( .A1(n4414), .A2(keyout[69]), .A3(\keys[5][69] ), .A4(n4402), .Y(n2962) );
  AO22X1_HVT U682 ( .A1(n4414), .A2(keyout[70]), .A3(\keys[5][70] ), .A4(n4402), .Y(n2963) );
  AO22X1_HVT U683 ( .A1(n4414), .A2(keyout[71]), .A3(\keys[5][71] ), .A4(n4402), .Y(n2964) );
  AO22X1_HVT U684 ( .A1(n4414), .A2(n3939), .A3(\keys[5][72] ), .A4(n4403), 
        .Y(n2965) );
  AO22X1_HVT U685 ( .A1(n4414), .A2(n3886), .A3(\keys[5][73] ), .A4(n4403), 
        .Y(n2966) );
  AO22X1_HVT U686 ( .A1(n4414), .A2(n3872), .A3(\keys[5][74] ), .A4(n4403), 
        .Y(n2967) );
  AO22X1_HVT U687 ( .A1(n4414), .A2(n3960), .A3(\keys[5][75] ), .A4(n4403), 
        .Y(n2968) );
  AO22X1_HVT U688 ( .A1(n4414), .A2(n3965), .A3(\keys[5][76] ), .A4(n4403), 
        .Y(n2969) );
  AO22X1_HVT U689 ( .A1(n4414), .A2(n3984), .A3(\keys[5][77] ), .A4(n4403), 
        .Y(n2970) );
  AO22X1_HVT U690 ( .A1(n4414), .A2(n3946), .A3(\keys[5][78] ), .A4(n4403), 
        .Y(n2971) );
  AO22X1_HVT U691 ( .A1(n4414), .A2(n3887), .A3(\keys[5][79] ), .A4(n4403), 
        .Y(n2972) );
  AO22X1_HVT U692 ( .A1(n4414), .A2(keyout[80]), .A3(\keys[5][80] ), .A4(n4403), .Y(n2973) );
  AO22X1_HVT U693 ( .A1(n4414), .A2(keyout[81]), .A3(\keys[5][81] ), .A4(n4403), .Y(n2974) );
  AO22X1_HVT U694 ( .A1(n4414), .A2(n3905), .A3(\keys[5][82] ), .A4(n4403), 
        .Y(n2975) );
  AO22X1_HVT U695 ( .A1(n4414), .A2(n3904), .A3(\keys[5][83] ), .A4(n4403), 
        .Y(n2976) );
  AO22X1_HVT U696 ( .A1(n4415), .A2(keyout[84]), .A3(\keys[5][84] ), .A4(n4404), .Y(n2977) );
  AO22X1_HVT U697 ( .A1(n4415), .A2(n1), .A3(\keys[5][85] ), .A4(n4404), .Y(
        n2978) );
  AO22X1_HVT U698 ( .A1(n4415), .A2(keyout[86]), .A3(\keys[5][86] ), .A4(n4404), .Y(n2979) );
  AO22X1_HVT U699 ( .A1(n4415), .A2(n1439), .A3(\keys[5][87] ), .A4(n4404), 
        .Y(n2980) );
  AO22X1_HVT U700 ( .A1(n4415), .A2(n4092), .A3(\keys[5][88] ), .A4(n4404), 
        .Y(n2981) );
  AO22X1_HVT U701 ( .A1(n4415), .A2(n3827), .A3(\keys[5][89] ), .A4(n4404), 
        .Y(n2982) );
  AO22X1_HVT U702 ( .A1(n4415), .A2(keyout[90]), .A3(\keys[5][90] ), .A4(n4404), .Y(n2983) );
  AO22X1_HVT U703 ( .A1(n4415), .A2(n4), .A3(\keys[5][91] ), .A4(n4404), .Y(
        n2984) );
  AO22X1_HVT U704 ( .A1(n4415), .A2(keyout[92]), .A3(\keys[5][92] ), .A4(n4404), .Y(n2985) );
  AO22X1_HVT U705 ( .A1(n4415), .A2(keyout[93]), .A3(\keys[5][93] ), .A4(n4404), .Y(n2986) );
  AO22X1_HVT U706 ( .A1(n4415), .A2(n3835), .A3(\keys[5][94] ), .A4(n4404), 
        .Y(n2987) );
  AO22X1_HVT U707 ( .A1(n4415), .A2(n3834), .A3(\keys[5][95] ), .A4(n4404), 
        .Y(n2988) );
  AO22X1_HVT U708 ( .A1(n4415), .A2(keyout[96]), .A3(\keys[5][96] ), .A4(n4405), .Y(n2989) );
  AO22X1_HVT U709 ( .A1(n4415), .A2(keyout[97]), .A3(\keys[5][97] ), .A4(n4405), .Y(n2990) );
  AO22X1_HVT U710 ( .A1(n4415), .A2(keyout[98]), .A3(\keys[5][98] ), .A4(n4405), .Y(n2991) );
  AO22X1_HVT U711 ( .A1(n4415), .A2(keyout[99]), .A3(\keys[5][99] ), .A4(n4405), .Y(n2992) );
  AO22X1_HVT U712 ( .A1(n4416), .A2(keyout[100]), .A3(\keys[5][100] ), .A4(
        n4405), .Y(n2993) );
  AO22X1_HVT U713 ( .A1(n4416), .A2(keyout[101]), .A3(\keys[5][101] ), .A4(
        n4405), .Y(n2994) );
  AO22X1_HVT U714 ( .A1(n4416), .A2(keyout[102]), .A3(\keys[5][102] ), .A4(
        n4405), .Y(n2995) );
  AO22X1_HVT U715 ( .A1(n4416), .A2(keyout[103]), .A3(\keys[5][103] ), .A4(
        n4405), .Y(n2996) );
  AO22X1_HVT U716 ( .A1(n4416), .A2(keyout[104]), .A3(\keys[5][104] ), .A4(
        n4405), .Y(n2997) );
  AO22X1_HVT U717 ( .A1(n4416), .A2(keyout[105]), .A3(\keys[5][105] ), .A4(
        n4405), .Y(n2998) );
  AO22X1_HVT U718 ( .A1(n4416), .A2(n3880), .A3(\keys[5][106] ), .A4(n4405), 
        .Y(n2999) );
  AO22X1_HVT U719 ( .A1(n4416), .A2(keyout[107]), .A3(\keys[5][107] ), .A4(
        n4405), .Y(n3000) );
  AO22X1_HVT U720 ( .A1(n4416), .A2(n3881), .A3(\keys[5][108] ), .A4(n4406), 
        .Y(n3001) );
  AO22X1_HVT U721 ( .A1(n4416), .A2(keyout[109]), .A3(\keys[5][109] ), .A4(
        n4406), .Y(n3002) );
  AO22X1_HVT U722 ( .A1(n4416), .A2(keyout[110]), .A3(\keys[5][110] ), .A4(
        n4406), .Y(n3003) );
  AO22X1_HVT U723 ( .A1(n4416), .A2(keyout[111]), .A3(\keys[5][111] ), .A4(
        n4406), .Y(n3004) );
  AO22X1_HVT U724 ( .A1(n4416), .A2(keyout[112]), .A3(\keys[5][112] ), .A4(
        n4406), .Y(n3005) );
  AO22X1_HVT U725 ( .A1(n4416), .A2(keyout[113]), .A3(\keys[5][113] ), .A4(
        n4406), .Y(n3006) );
  AO22X1_HVT U726 ( .A1(n4416), .A2(keyout[114]), .A3(\keys[5][114] ), .A4(
        n4406), .Y(n3007) );
  AO22X1_HVT U727 ( .A1(n4416), .A2(keyout[115]), .A3(\keys[5][115] ), .A4(
        n4406), .Y(n3008) );
  AO22X1_HVT U728 ( .A1(n4417), .A2(keyout[116]), .A3(\keys[5][116] ), .A4(
        n4406), .Y(n3009) );
  AO22X1_HVT U729 ( .A1(n4417), .A2(keyout[117]), .A3(\keys[5][117] ), .A4(
        n4406), .Y(n3010) );
  AO22X1_HVT U730 ( .A1(n4417), .A2(keyout[118]), .A3(\keys[5][118] ), .A4(
        n4406), .Y(n3011) );
  AO22X1_HVT U731 ( .A1(n4417), .A2(keyout[119]), .A3(\keys[5][119] ), .A4(
        n4406), .Y(n3012) );
  AO22X1_HVT U732 ( .A1(n4417), .A2(n4095), .A3(\keys[5][120] ), .A4(n4407), 
        .Y(n3013) );
  AO22X1_HVT U733 ( .A1(n4417), .A2(n3829), .A3(\keys[5][121] ), .A4(n4407), 
        .Y(n3014) );
  AO22X1_HVT U734 ( .A1(n4417), .A2(n3803), .A3(\keys[5][122] ), .A4(n4407), 
        .Y(n3015) );
  AO22X1_HVT U735 ( .A1(n4417), .A2(n3817), .A3(\keys[5][123] ), .A4(n4407), 
        .Y(n3016) );
  AO22X1_HVT U736 ( .A1(n4417), .A2(n3846), .A3(\keys[5][124] ), .A4(n4407), 
        .Y(n3017) );
  AO22X1_HVT U737 ( .A1(n4417), .A2(n3823), .A3(\keys[5][125] ), .A4(n4407), 
        .Y(n3018) );
  AO22X1_HVT U738 ( .A1(n4417), .A2(n4098), .A3(\keys[5][126] ), .A4(n4407), 
        .Y(n3019) );
  AO22X1_HVT U739 ( .A1(n4417), .A2(n4101), .A3(\keys[5][127] ), .A4(n4407), 
        .Y(n3020) );
  AO22X1_HVT U740 ( .A1(n4385), .A2(n3999), .A3(\keys[4][0] ), .A4(n4384), .Y(
        n3021) );
  AO22X1_HVT U741 ( .A1(n4386), .A2(n4002), .A3(\keys[4][1] ), .A4(n4384), .Y(
        n3022) );
  AO22X1_HVT U742 ( .A1(n4386), .A2(n4003), .A3(\keys[4][2] ), .A4(n4384), .Y(
        n3023) );
  AO22X1_HVT U743 ( .A1(n4386), .A2(n4006), .A3(\keys[4][3] ), .A4(n4384), .Y(
        n3024) );
  AO22X1_HVT U744 ( .A1(n4386), .A2(n4009), .A3(\keys[4][4] ), .A4(n4384), .Y(
        n3025) );
  AO22X1_HVT U745 ( .A1(n4386), .A2(n4012), .A3(\keys[4][5] ), .A4(n4384), .Y(
        n3026) );
  AO22X1_HVT U746 ( .A1(n4386), .A2(n4015), .A3(\keys[4][6] ), .A4(n4384), .Y(
        n3027) );
  AO22X1_HVT U747 ( .A1(n4387), .A2(n4016), .A3(\keys[4][7] ), .A4(n4384), .Y(
        n3028) );
  AO22X1_HVT U748 ( .A1(n4387), .A2(n4019), .A3(\keys[4][8] ), .A4(n4384), .Y(
        n3029) );
  AO22X1_HVT U749 ( .A1(n4387), .A2(n4022), .A3(\keys[4][9] ), .A4(n4384), .Y(
        n3030) );
  AO22X1_HVT U750 ( .A1(n4387), .A2(n4025), .A3(\keys[4][10] ), .A4(n4384), 
        .Y(n3031) );
  AO22X1_HVT U751 ( .A1(n4387), .A2(n4028), .A3(\keys[4][11] ), .A4(n4384), 
        .Y(n3032) );
  AO22X1_HVT U752 ( .A1(n4387), .A2(n4031), .A3(\keys[4][12] ), .A4(n4384), 
        .Y(n3033) );
  AO22X1_HVT U753 ( .A1(n4387), .A2(n4034), .A3(\keys[4][13] ), .A4(n4383), 
        .Y(n3034) );
  AO22X1_HVT U754 ( .A1(n4387), .A2(n4037), .A3(\keys[4][14] ), .A4(n4383), 
        .Y(n3035) );
  AO22X1_HVT U755 ( .A1(n4387), .A2(n4040), .A3(\keys[4][15] ), .A4(n4383), 
        .Y(n3036) );
  AO22X1_HVT U756 ( .A1(n4387), .A2(n4043), .A3(\keys[4][16] ), .A4(n4383), 
        .Y(n3037) );
  AO22X1_HVT U757 ( .A1(n4387), .A2(n4046), .A3(\keys[4][17] ), .A4(n4383), 
        .Y(n3038) );
  AO22X1_HVT U758 ( .A1(n4387), .A2(n4049), .A3(\keys[4][18] ), .A4(n4383), 
        .Y(n3039) );
  AO22X1_HVT U759 ( .A1(n4387), .A2(n4052), .A3(\keys[4][19] ), .A4(n4383), 
        .Y(n3040) );
  AO22X1_HVT U760 ( .A1(n4387), .A2(n4055), .A3(\keys[4][20] ), .A4(n4383), 
        .Y(n3041) );
  AO22X1_HVT U761 ( .A1(n4387), .A2(n4058), .A3(\keys[4][21] ), .A4(n4383), 
        .Y(n3042) );
  AO22X1_HVT U762 ( .A1(n4387), .A2(n4061), .A3(\keys[4][22] ), .A4(n4383), 
        .Y(n3043) );
  AO22X1_HVT U763 ( .A1(n4388), .A2(n4064), .A3(\keys[4][23] ), .A4(n4383), 
        .Y(n3044) );
  AO22X1_HVT U764 ( .A1(n4388), .A2(n4067), .A3(\keys[4][24] ), .A4(n4383), 
        .Y(n3045) );
  AO22X1_HVT U765 ( .A1(n4388), .A2(n4069), .A3(\keys[4][25] ), .A4(n4383), 
        .Y(n3046) );
  AO22X1_HVT U766 ( .A1(n4388), .A2(n4072), .A3(\keys[4][26] ), .A4(n4382), 
        .Y(n3047) );
  AO22X1_HVT U767 ( .A1(n4388), .A2(n4075), .A3(\keys[4][27] ), .A4(n4382), 
        .Y(n3048) );
  AO22X1_HVT U768 ( .A1(n4388), .A2(n4078), .A3(\keys[4][28] ), .A4(n4382), 
        .Y(n3049) );
  AO22X1_HVT U769 ( .A1(n4388), .A2(n4081), .A3(\keys[4][29] ), .A4(n4382), 
        .Y(n3050) );
  AO22X1_HVT U770 ( .A1(n4388), .A2(n4083), .A3(\keys[4][30] ), .A4(n4382), 
        .Y(n3051) );
  AO22X1_HVT U771 ( .A1(n4388), .A2(keyout[31]), .A3(\keys[4][31] ), .A4(n4382), .Y(n3052) );
  AO22X1_HVT U772 ( .A1(n4388), .A2(keyout[32]), .A3(\keys[4][32] ), .A4(n4382), .Y(n3053) );
  AO22X1_HVT U773 ( .A1(n4388), .A2(n3876), .A3(\keys[4][33] ), .A4(n4382), 
        .Y(n3054) );
  AO22X1_HVT U774 ( .A1(n4388), .A2(n3913), .A3(\keys[4][34] ), .A4(n4382), 
        .Y(n3055) );
  AO22X1_HVT U775 ( .A1(n4388), .A2(keyout[35]), .A3(\keys[4][35] ), .A4(n4382), .Y(n3056) );
  AO22X1_HVT U776 ( .A1(n4388), .A2(keyout[36]), .A3(\keys[4][36] ), .A4(n4382), .Y(n3057) );
  AO22X1_HVT U777 ( .A1(n4388), .A2(n3819), .A3(\keys[4][37] ), .A4(n4382), 
        .Y(n3058) );
  AO22X1_HVT U778 ( .A1(n4388), .A2(keyout[38]), .A3(\keys[4][38] ), .A4(n4382), .Y(n3059) );
  AO22X1_HVT U779 ( .A1(n4389), .A2(keyout[39]), .A3(\keys[4][39] ), .A4(n4381), .Y(n3060) );
  AO22X1_HVT U780 ( .A1(n4389), .A2(n3953), .A3(\keys[4][40] ), .A4(n4381), 
        .Y(n3061) );
  AO22X1_HVT U781 ( .A1(n4389), .A2(n3884), .A3(\keys[4][41] ), .A4(n4381), 
        .Y(n3062) );
  AO22X1_HVT U782 ( .A1(n4389), .A2(n3974), .A3(\keys[4][42] ), .A4(n4381), 
        .Y(n3063) );
  AO22X1_HVT U783 ( .A1(n4389), .A2(keyout[43]), .A3(\keys[4][43] ), .A4(n4381), .Y(n3064) );
  AO22X1_HVT U785 ( .A1(n4389), .A2(n3935), .A3(\keys[4][45] ), .A4(n4381), 
        .Y(n3066) );
  AO22X1_HVT U786 ( .A1(n4389), .A2(n3945), .A3(\keys[4][46] ), .A4(n4381), 
        .Y(n3067) );
  AO22X1_HVT U787 ( .A1(n4389), .A2(n3885), .A3(\keys[4][47] ), .A4(n4381), 
        .Y(n3068) );
  AO22X1_HVT U788 ( .A1(n4389), .A2(keyout[48]), .A3(\keys[4][48] ), .A4(n4381), .Y(n3069) );
  AO22X1_HVT U789 ( .A1(n4389), .A2(keyout[49]), .A3(\keys[4][49] ), .A4(n4381), .Y(n3070) );
  AO22X1_HVT U790 ( .A1(n4389), .A2(keyout[50]), .A3(\keys[4][50] ), .A4(n4381), .Y(n3071) );
  AO22X1_HVT U791 ( .A1(n4389), .A2(n3937), .A3(\keys[4][51] ), .A4(n4381), 
        .Y(n3072) );
  AO22X1_HVT U792 ( .A1(n4389), .A2(keyout[52]), .A3(\keys[4][52] ), .A4(n4380), .Y(n3073) );
  AO22X1_HVT U793 ( .A1(n4389), .A2(n3920), .A3(\keys[4][53] ), .A4(n4380), 
        .Y(n3074) );
  AO22X1_HVT U794 ( .A1(n4389), .A2(keyout[54]), .A3(\keys[4][54] ), .A4(n4380), .Y(n3075) );
  AO22X1_HVT U795 ( .A1(n4390), .A2(n3922), .A3(\keys[4][55] ), .A4(n4380), 
        .Y(n3076) );
  AO22X1_HVT U796 ( .A1(n4390), .A2(n3941), .A3(\keys[4][56] ), .A4(n4380), 
        .Y(n3077) );
  AO22X1_HVT U797 ( .A1(n4390), .A2(keyout[57]), .A3(\keys[4][57] ), .A4(n4380), .Y(n3078) );
  AO22X1_HVT U798 ( .A1(n4390), .A2(keyout[58]), .A3(\keys[4][58] ), .A4(n4380), .Y(n3079) );
  AO22X1_HVT U799 ( .A1(n4390), .A2(n4089), .A3(\keys[4][59] ), .A4(n4380), 
        .Y(n3080) );
  AO22X1_HVT U800 ( .A1(n4390), .A2(n3943), .A3(\keys[4][60] ), .A4(n4380), 
        .Y(n3081) );
  AO22X1_HVT U801 ( .A1(n4390), .A2(keyout[61]), .A3(\keys[4][61] ), .A4(n4380), .Y(n3082) );
  AO22X1_HVT U802 ( .A1(n4390), .A2(n3832), .A3(\keys[4][62] ), .A4(n4380), 
        .Y(n3083) );
  AO22X1_HVT U803 ( .A1(n4390), .A2(n3859), .A3(\keys[4][63] ), .A4(n4380), 
        .Y(n3084) );
  AO22X1_HVT U804 ( .A1(n4390), .A2(keyout[64]), .A3(\keys[4][64] ), .A4(n4380), .Y(n3085) );
  AO22X1_HVT U805 ( .A1(n4390), .A2(n3883), .A3(\keys[4][65] ), .A4(n4379), 
        .Y(n3086) );
  AO22X1_HVT U806 ( .A1(n4390), .A2(n3914), .A3(\keys[4][66] ), .A4(n4379), 
        .Y(n3087) );
  AO22X1_HVT U807 ( .A1(n4390), .A2(n3825), .A3(\keys[4][67] ), .A4(n4379), 
        .Y(n3088) );
  AO22X1_HVT U808 ( .A1(n4390), .A2(keyout[68]), .A3(\keys[4][68] ), .A4(n4379), .Y(n3089) );
  AO22X1_HVT U809 ( .A1(n4390), .A2(keyout[69]), .A3(\keys[4][69] ), .A4(n4379), .Y(n3090) );
  AO22X1_HVT U810 ( .A1(n4390), .A2(keyout[70]), .A3(\keys[4][70] ), .A4(n4379), .Y(n3091) );
  AO22X1_HVT U811 ( .A1(n4391), .A2(keyout[71]), .A3(\keys[4][71] ), .A4(n4379), .Y(n3092) );
  AO22X1_HVT U812 ( .A1(n4391), .A2(n3951), .A3(\keys[4][72] ), .A4(n4379), 
        .Y(n3093) );
  AO22X1_HVT U813 ( .A1(n4391), .A2(n3896), .A3(\keys[4][73] ), .A4(n4379), 
        .Y(n3094) );
  AO22X1_HVT U816 ( .A1(n4391), .A2(n3967), .A3(\keys[4][76] ), .A4(n4379), 
        .Y(n3097) );
  AO22X1_HVT U817 ( .A1(n4391), .A2(n3986), .A3(\keys[4][77] ), .A4(n4379), 
        .Y(n3098) );
  AO22X1_HVT U818 ( .A1(n4391), .A2(n3947), .A3(\keys[4][78] ), .A4(n4378), 
        .Y(n3099) );
  AO22X1_HVT U819 ( .A1(n4391), .A2(n3898), .A3(\keys[4][79] ), .A4(n4378), 
        .Y(n3100) );
  AO22X1_HVT U820 ( .A1(n4391), .A2(n3931), .A3(\keys[4][80] ), .A4(n4378), 
        .Y(n3101) );
  AO22X1_HVT U821 ( .A1(n4391), .A2(n3811), .A3(\keys[4][81] ), .A4(n4378), 
        .Y(n3102) );
  AO22X1_HVT U822 ( .A1(n4391), .A2(n3977), .A3(\keys[4][82] ), .A4(n4378), 
        .Y(n3103) );
  AO22X1_HVT U823 ( .A1(n4391), .A2(n3927), .A3(\keys[4][83] ), .A4(n4378), 
        .Y(n3104) );
  AO22X1_HVT U824 ( .A1(n4391), .A2(n1438), .A3(\keys[4][84] ), .A4(n4378), 
        .Y(n3105) );
  AO22X1_HVT U825 ( .A1(n4391), .A2(n1), .A3(\keys[4][85] ), .A4(n4378), .Y(
        n3106) );
  AO22X1_HVT U826 ( .A1(n4391), .A2(n1436), .A3(\keys[4][86] ), .A4(n4378), 
        .Y(n3107) );
  AO22X1_HVT U827 ( .A1(n4392), .A2(n1439), .A3(\keys[4][87] ), .A4(n4378), 
        .Y(n3108) );
  AO22X1_HVT U828 ( .A1(n4392), .A2(n4093), .A3(\keys[4][88] ), .A4(n4378), 
        .Y(n3109) );
  AO22X1_HVT U829 ( .A1(n4392), .A2(n3827), .A3(\keys[4][89] ), .A4(n4378), 
        .Y(n3110) );
  AO22X1_HVT U830 ( .A1(n4392), .A2(n3949), .A3(\keys[4][90] ), .A4(n4378), 
        .Y(n3111) );
  AO22X1_HVT U831 ( .A1(n4392), .A2(n3816), .A3(\keys[4][91] ), .A4(n4377), 
        .Y(n3112) );
  AO22X1_HVT U832 ( .A1(n4392), .A2(n3831), .A3(\keys[4][92] ), .A4(n4377), 
        .Y(n3113) );
  AO22X1_HVT U833 ( .A1(n4392), .A2(keyout[93]), .A3(\keys[4][93] ), .A4(n4377), .Y(n3114) );
  AO22X1_HVT U834 ( .A1(n4392), .A2(n3835), .A3(\keys[4][94] ), .A4(n4377), 
        .Y(n3115) );
  AO22X1_HVT U835 ( .A1(n4392), .A2(n3834), .A3(\keys[4][95] ), .A4(n4377), 
        .Y(n3116) );
  AO22X1_HVT U836 ( .A1(n4392), .A2(keyout[96]), .A3(\keys[4][96] ), .A4(n4377), .Y(n3117) );
  AO22X1_HVT U837 ( .A1(n4392), .A2(keyout[97]), .A3(\keys[4][97] ), .A4(n4377), .Y(n3118) );
  AO22X1_HVT U838 ( .A1(n4392), .A2(keyout[98]), .A3(\keys[4][98] ), .A4(n4377), .Y(n3119) );
  AO22X1_HVT U839 ( .A1(n4392), .A2(keyout[99]), .A3(\keys[4][99] ), .A4(n4377), .Y(n3120) );
  AO22X1_HVT U840 ( .A1(n4392), .A2(keyout[100]), .A3(\keys[4][100] ), .A4(
        n4377), .Y(n3121) );
  AO22X1_HVT U841 ( .A1(n4392), .A2(keyout[101]), .A3(\keys[4][101] ), .A4(
        n4377), .Y(n3122) );
  AO22X1_HVT U842 ( .A1(n4392), .A2(keyout[102]), .A3(\keys[4][102] ), .A4(
        n4377), .Y(n3123) );
  AO22X1_HVT U843 ( .A1(n4393), .A2(keyout[103]), .A3(\keys[4][103] ), .A4(
        n4377), .Y(n3124) );
  AO22X1_HVT U844 ( .A1(n4393), .A2(n3839), .A3(\keys[4][104] ), .A4(n4376), 
        .Y(n3125) );
  AO22X1_HVT U845 ( .A1(n4393), .A2(keyout[105]), .A3(\keys[4][105] ), .A4(
        n4376), .Y(n3126) );
  AO22X1_HVT U846 ( .A1(n4393), .A2(n3880), .A3(\keys[4][106] ), .A4(n4376), 
        .Y(n3127) );
  AO22X1_HVT U847 ( .A1(n4393), .A2(n3820), .A3(\keys[4][107] ), .A4(n4376), 
        .Y(n3128) );
  AO22X1_HVT U848 ( .A1(n4393), .A2(n3892), .A3(\keys[4][108] ), .A4(n4376), 
        .Y(n3129) );
  AO22X1_HVT U849 ( .A1(n4393), .A2(n3873), .A3(\keys[4][109] ), .A4(n4376), 
        .Y(n3130) );
  AO22X1_HVT U850 ( .A1(n4393), .A2(keyout[110]), .A3(\keys[4][110] ), .A4(
        n4376), .Y(n3131) );
  AO22X1_HVT U851 ( .A1(n4393), .A2(keyout[111]), .A3(\keys[4][111] ), .A4(
        n4376), .Y(n3132) );
  AO22X1_HVT U852 ( .A1(n4393), .A2(keyout[112]), .A3(\keys[4][112] ), .A4(
        n4376), .Y(n3133) );
  AO22X1_HVT U853 ( .A1(n4393), .A2(keyout[113]), .A3(\keys[4][113] ), .A4(
        n4376), .Y(n3134) );
  AO22X1_HVT U854 ( .A1(n4393), .A2(keyout[114]), .A3(\keys[4][114] ), .A4(
        n4376), .Y(n3135) );
  AO22X1_HVT U855 ( .A1(n4393), .A2(n3915), .A3(\keys[4][115] ), .A4(n4376), 
        .Y(n3136) );
  AO22X1_HVT U856 ( .A1(n4393), .A2(keyout[116]), .A3(\keys[4][116] ), .A4(
        n4376), .Y(n3137) );
  AO22X1_HVT U857 ( .A1(n4393), .A2(keyout[117]), .A3(\keys[4][117] ), .A4(
        n4375), .Y(n3138) );
  AO22X1_HVT U858 ( .A1(n4393), .A2(keyout[118]), .A3(\keys[4][118] ), .A4(
        n4375), .Y(n3139) );
  AO22X1_HVT U859 ( .A1(n4394), .A2(keyout[119]), .A3(\keys[4][119] ), .A4(
        n4375), .Y(n3140) );
  AO22X1_HVT U860 ( .A1(n4394), .A2(n4096), .A3(\keys[4][120] ), .A4(n4375), 
        .Y(n3141) );
  AO22X1_HVT U861 ( .A1(n4394), .A2(n3829), .A3(\keys[4][121] ), .A4(n4375), 
        .Y(n3142) );
  AO22X1_HVT U862 ( .A1(n4394), .A2(n3803), .A3(\keys[4][122] ), .A4(n4375), 
        .Y(n3143) );
  AO22X1_HVT U863 ( .A1(n4394), .A2(n3817), .A3(\keys[4][123] ), .A4(n4375), 
        .Y(n3144) );
  AO22X1_HVT U864 ( .A1(n4394), .A2(n3846), .A3(\keys[4][124] ), .A4(n4375), 
        .Y(n3145) );
  AO22X1_HVT U865 ( .A1(n4394), .A2(n3823), .A3(\keys[4][125] ), .A4(n4375), 
        .Y(n3146) );
  AO22X1_HVT U866 ( .A1(n4394), .A2(n4099), .A3(\keys[4][126] ), .A4(n4375), 
        .Y(n3147) );
  AO22X1_HVT U867 ( .A1(n4394), .A2(n4102), .A3(\keys[4][127] ), .A4(n4375), 
        .Y(n3148) );
  AO22X1_HVT U868 ( .A1(n4363), .A2(n3999), .A3(\keys[3][0] ), .A4(n4362), .Y(
        n3149) );
  AO22X1_HVT U869 ( .A1(n4364), .A2(n4002), .A3(\keys[3][1] ), .A4(n4362), .Y(
        n3150) );
  AO22X1_HVT U870 ( .A1(n4364), .A2(n4003), .A3(\keys[3][2] ), .A4(n4362), .Y(
        n3151) );
  AO22X1_HVT U871 ( .A1(n4364), .A2(n4006), .A3(\keys[3][3] ), .A4(n4362), .Y(
        n3152) );
  AO22X1_HVT U872 ( .A1(n4364), .A2(n4009), .A3(\keys[3][4] ), .A4(n4362), .Y(
        n3153) );
  AO22X1_HVT U873 ( .A1(n4364), .A2(n4012), .A3(\keys[3][5] ), .A4(n4362), .Y(
        n3154) );
  AO22X1_HVT U874 ( .A1(n4364), .A2(n4015), .A3(\keys[3][6] ), .A4(n4362), .Y(
        n3155) );
  AO22X1_HVT U875 ( .A1(n4365), .A2(n4016), .A3(\keys[3][7] ), .A4(n4362), .Y(
        n3156) );
  AO22X1_HVT U876 ( .A1(n4365), .A2(n4019), .A3(\keys[3][8] ), .A4(n4362), .Y(
        n3157) );
  AO22X1_HVT U877 ( .A1(n4365), .A2(n4022), .A3(\keys[3][9] ), .A4(n4362), .Y(
        n3158) );
  AO22X1_HVT U878 ( .A1(n4365), .A2(n4025), .A3(\keys[3][10] ), .A4(n4362), 
        .Y(n3159) );
  AO22X1_HVT U879 ( .A1(n4365), .A2(n4028), .A3(\keys[3][11] ), .A4(n4362), 
        .Y(n3160) );
  AO22X1_HVT U880 ( .A1(n4365), .A2(n4031), .A3(\keys[3][12] ), .A4(n4362), 
        .Y(n3161) );
  AO22X1_HVT U881 ( .A1(n4365), .A2(n4034), .A3(\keys[3][13] ), .A4(n4361), 
        .Y(n3162) );
  AO22X1_HVT U882 ( .A1(n4365), .A2(n4037), .A3(\keys[3][14] ), .A4(n4361), 
        .Y(n3163) );
  AO22X1_HVT U883 ( .A1(n4365), .A2(n4040), .A3(\keys[3][15] ), .A4(n4361), 
        .Y(n3164) );
  AO22X1_HVT U884 ( .A1(n4365), .A2(n4043), .A3(\keys[3][16] ), .A4(n4361), 
        .Y(n3165) );
  AO22X1_HVT U885 ( .A1(n4365), .A2(n4046), .A3(\keys[3][17] ), .A4(n4361), 
        .Y(n3166) );
  AO22X1_HVT U886 ( .A1(n4365), .A2(n4049), .A3(\keys[3][18] ), .A4(n4361), 
        .Y(n3167) );
  AO22X1_HVT U887 ( .A1(n4365), .A2(n4052), .A3(\keys[3][19] ), .A4(n4361), 
        .Y(n3168) );
  AO22X1_HVT U888 ( .A1(n4365), .A2(n4055), .A3(\keys[3][20] ), .A4(n4361), 
        .Y(n3169) );
  AO22X1_HVT U889 ( .A1(n4365), .A2(n4058), .A3(\keys[3][21] ), .A4(n4361), 
        .Y(n3170) );
  AO22X1_HVT U890 ( .A1(n4365), .A2(n4061), .A3(\keys[3][22] ), .A4(n4361), 
        .Y(n3171) );
  AO22X1_HVT U891 ( .A1(n4366), .A2(n4064), .A3(\keys[3][23] ), .A4(n4361), 
        .Y(n3172) );
  AO22X1_HVT U892 ( .A1(n4366), .A2(n4067), .A3(\keys[3][24] ), .A4(n4361), 
        .Y(n3173) );
  AO22X1_HVT U893 ( .A1(n4366), .A2(n4069), .A3(\keys[3][25] ), .A4(n4361), 
        .Y(n3174) );
  AO22X1_HVT U894 ( .A1(n4366), .A2(n4072), .A3(\keys[3][26] ), .A4(n4360), 
        .Y(n3175) );
  AO22X1_HVT U895 ( .A1(n4366), .A2(n4075), .A3(\keys[3][27] ), .A4(n4360), 
        .Y(n3176) );
  AO22X1_HVT U896 ( .A1(n4366), .A2(n4078), .A3(\keys[3][28] ), .A4(n4360), 
        .Y(n3177) );
  AO22X1_HVT U897 ( .A1(n4366), .A2(n4081), .A3(\keys[3][29] ), .A4(n4360), 
        .Y(n3178) );
  AO22X1_HVT U898 ( .A1(n4366), .A2(n4083), .A3(\keys[3][30] ), .A4(n4360), 
        .Y(n3179) );
  AO22X1_HVT U899 ( .A1(n4366), .A2(n3852), .A3(\keys[3][31] ), .A4(n4360), 
        .Y(n3180) );
  AO22X1_HVT U900 ( .A1(n4366), .A2(keyout[32]), .A3(\keys[3][32] ), .A4(n4360), .Y(n3181) );
  AO22X1_HVT U901 ( .A1(n4366), .A2(n3876), .A3(\keys[3][33] ), .A4(n4360), 
        .Y(n3182) );
  AO22X1_HVT U902 ( .A1(n4366), .A2(n3913), .A3(\keys[3][34] ), .A4(n4360), 
        .Y(n3183) );
  AO22X1_HVT U903 ( .A1(n4366), .A2(keyout[35]), .A3(\keys[3][35] ), .A4(n4360), .Y(n3184) );
  AO22X1_HVT U904 ( .A1(n4366), .A2(keyout[36]), .A3(\keys[3][36] ), .A4(n4360), .Y(n3185) );
  AO22X1_HVT U905 ( .A1(n4366), .A2(n3819), .A3(\keys[3][37] ), .A4(n4360), 
        .Y(n3186) );
  AO22X1_HVT U906 ( .A1(n4366), .A2(keyout[38]), .A3(\keys[3][38] ), .A4(n4360), .Y(n3187) );
  AO22X1_HVT U907 ( .A1(n4367), .A2(keyout[39]), .A3(\keys[3][39] ), .A4(n4359), .Y(n3188) );
  AO22X1_HVT U908 ( .A1(n4367), .A2(n3952), .A3(\keys[3][40] ), .A4(n4359), 
        .Y(n3189) );
  AO22X1_HVT U909 ( .A1(n4367), .A2(n3854), .A3(\keys[3][41] ), .A4(n4359), 
        .Y(n3190) );
  AO22X1_HVT U910 ( .A1(n4367), .A2(n3974), .A3(\keys[3][42] ), .A4(n4359), 
        .Y(n3191) );
  AO22X1_HVT U911 ( .A1(n4367), .A2(n3890), .A3(\keys[3][43] ), .A4(n4359), 
        .Y(n3192) );
  AO22X1_HVT U912 ( .A1(n4367), .A2(n3902), .A3(\keys[3][44] ), .A4(n4359), 
        .Y(n3193) );
  AO22X1_HVT U913 ( .A1(n4367), .A2(n3935), .A3(\keys[3][45] ), .A4(n4359), 
        .Y(n3194) );
  AO22X1_HVT U914 ( .A1(n4367), .A2(n3944), .A3(\keys[3][46] ), .A4(n4359), 
        .Y(n3195) );
  AO22X1_HVT U915 ( .A1(n4367), .A2(n3850), .A3(\keys[3][47] ), .A4(n4359), 
        .Y(n3196) );
  AO22X1_HVT U916 ( .A1(n4367), .A2(n1427), .A3(\keys[3][48] ), .A4(n4359), 
        .Y(n3197) );
  AO22X1_HVT U917 ( .A1(n4367), .A2(n14), .A3(\keys[3][49] ), .A4(n4359), .Y(
        n3198) );
  AO22X1_HVT U918 ( .A1(n4367), .A2(n1432), .A3(\keys[3][50] ), .A4(n4359), 
        .Y(n3199) );
  AO22X1_HVT U919 ( .A1(n4367), .A2(n3937), .A3(\keys[3][51] ), .A4(n4359), 
        .Y(n3200) );
  AO22X1_HVT U920 ( .A1(n4367), .A2(keyout[52]), .A3(\keys[3][52] ), .A4(n4358), .Y(n3201) );
  AO22X1_HVT U921 ( .A1(n4367), .A2(n3920), .A3(\keys[3][53] ), .A4(n4358), 
        .Y(n3202) );
  AO22X1_HVT U922 ( .A1(n4367), .A2(keyout[54]), .A3(\keys[3][54] ), .A4(n4358), .Y(n3203) );
  AO22X1_HVT U923 ( .A1(n4368), .A2(n3922), .A3(\keys[3][55] ), .A4(n4358), 
        .Y(n3204) );
  AO22X1_HVT U924 ( .A1(n4368), .A2(n3941), .A3(\keys[3][56] ), .A4(n4358), 
        .Y(n3205) );
  AO22X1_HVT U925 ( .A1(n4368), .A2(n4085), .A3(\keys[3][57] ), .A4(n4358), 
        .Y(n3206) );
  AO22X1_HVT U926 ( .A1(n4368), .A2(n4087), .A3(\keys[3][58] ), .A4(n4358), 
        .Y(n3207) );
  AO22X1_HVT U927 ( .A1(n4368), .A2(n4090), .A3(\keys[3][59] ), .A4(n4358), 
        .Y(n3208) );
  AO22X1_HVT U928 ( .A1(n4368), .A2(n3943), .A3(\keys[3][60] ), .A4(n4358), 
        .Y(n3209) );
  AO22X1_HVT U929 ( .A1(n4368), .A2(n3805), .A3(\keys[3][61] ), .A4(n4358), 
        .Y(n3210) );
  AO22X1_HVT U930 ( .A1(n4368), .A2(n3833), .A3(\keys[3][62] ), .A4(n4358), 
        .Y(n3211) );
  AO22X1_HVT U931 ( .A1(n4368), .A2(n3861), .A3(\keys[3][63] ), .A4(n4358), 
        .Y(n3212) );
  AO22X1_HVT U932 ( .A1(n4368), .A2(keyout[64]), .A3(\keys[3][64] ), .A4(n4358), .Y(n3213) );
  AO22X1_HVT U933 ( .A1(n4368), .A2(n3883), .A3(\keys[3][65] ), .A4(n4357), 
        .Y(n3214) );
  AO22X1_HVT U934 ( .A1(n4368), .A2(n3914), .A3(\keys[3][66] ), .A4(n4357), 
        .Y(n3215) );
  AO22X1_HVT U935 ( .A1(n4368), .A2(n3938), .A3(\keys[3][67] ), .A4(n4357), 
        .Y(n3216) );
  AO22X1_HVT U936 ( .A1(n4368), .A2(keyout[68]), .A3(\keys[3][68] ), .A4(n4357), .Y(n3217) );
  AO22X1_HVT U937 ( .A1(n4368), .A2(keyout[69]), .A3(\keys[3][69] ), .A4(n4357), .Y(n3218) );
  AO22X1_HVT U938 ( .A1(n4368), .A2(keyout[70]), .A3(\keys[3][70] ), .A4(n4357), .Y(n3219) );
  AO22X1_HVT U939 ( .A1(n4369), .A2(keyout[71]), .A3(\keys[3][71] ), .A4(n4357), .Y(n3220) );
  AO22X1_HVT U940 ( .A1(n4369), .A2(n3951), .A3(\keys[3][72] ), .A4(n4357), 
        .Y(n3221) );
  AO22X1_HVT U941 ( .A1(n4369), .A2(n3896), .A3(\keys[3][73] ), .A4(n4357), 
        .Y(n3222) );
  AO22X1_HVT U942 ( .A1(n4369), .A2(n3979), .A3(\keys[3][74] ), .A4(n4357), 
        .Y(n3223) );
  AO22X1_HVT U943 ( .A1(n4369), .A2(n3959), .A3(\keys[3][75] ), .A4(n4357), 
        .Y(n3224) );
  AO22X1_HVT U944 ( .A1(n4369), .A2(n3966), .A3(\keys[3][76] ), .A4(n4357), 
        .Y(n3225) );
  AO22X1_HVT U945 ( .A1(n4369), .A2(n3985), .A3(\keys[3][77] ), .A4(n4357), 
        .Y(n3226) );
  AO22X1_HVT U946 ( .A1(n4369), .A2(n3946), .A3(\keys[3][78] ), .A4(n4356), 
        .Y(n3227) );
  AO22X1_HVT U947 ( .A1(n4369), .A2(n3898), .A3(\keys[3][79] ), .A4(n4356), 
        .Y(n3228) );
  AO22X1_HVT U948 ( .A1(n4369), .A2(n3931), .A3(\keys[3][80] ), .A4(n4356), 
        .Y(n3229) );
  AO22X1_HVT U949 ( .A1(n4369), .A2(n3811), .A3(\keys[3][81] ), .A4(n4356), 
        .Y(n3230) );
  AO22X1_HVT U950 ( .A1(n4369), .A2(n3977), .A3(\keys[3][82] ), .A4(n4356), 
        .Y(n3231) );
  AO22X1_HVT U951 ( .A1(n4369), .A2(n3916), .A3(\keys[3][83] ), .A4(n4356), 
        .Y(n3232) );
  AO22X1_HVT U952 ( .A1(n4369), .A2(n1438), .A3(\keys[3][84] ), .A4(n4356), 
        .Y(n3233) );
  AO22X1_HVT U953 ( .A1(n4369), .A2(n2), .A3(\keys[3][85] ), .A4(n4356), .Y(
        n3234) );
  AO22X1_HVT U954 ( .A1(n4369), .A2(n1436), .A3(\keys[3][86] ), .A4(n4356), 
        .Y(n3235) );
  AO22X1_HVT U955 ( .A1(n4370), .A2(n1439), .A3(\keys[3][87] ), .A4(n4356), 
        .Y(n3236) );
  AO22X1_HVT U956 ( .A1(n4370), .A2(n4093), .A3(\keys[3][88] ), .A4(n4356), 
        .Y(n3237) );
  AO22X1_HVT U957 ( .A1(n4370), .A2(n3863), .A3(\keys[3][89] ), .A4(n4356), 
        .Y(n3238) );
  AO22X1_HVT U960 ( .A1(n4370), .A2(n3831), .A3(\keys[3][92] ), .A4(n4355), 
        .Y(n3241) );
  AO22X1_HVT U961 ( .A1(n4370), .A2(keyout[93]), .A3(\keys[3][93] ), .A4(n4355), .Y(n3242) );
  AO22X1_HVT U962 ( .A1(n4370), .A2(n3865), .A3(\keys[3][94] ), .A4(n4355), 
        .Y(n3243) );
  AO22X1_HVT U963 ( .A1(n4370), .A2(n3869), .A3(\keys[3][95] ), .A4(n4355), 
        .Y(n3244) );
  AO22X1_HVT U964 ( .A1(n4370), .A2(keyout[96]), .A3(\keys[3][96] ), .A4(n4355), .Y(n3245) );
  AO22X1_HVT U965 ( .A1(n4370), .A2(keyout[97]), .A3(\keys[3][97] ), .A4(n4355), .Y(n3246) );
  AO22X1_HVT U966 ( .A1(n4370), .A2(keyout[98]), .A3(\keys[3][98] ), .A4(n4355), .Y(n3247) );
  AO22X1_HVT U967 ( .A1(n4370), .A2(keyout[99]), .A3(\keys[3][99] ), .A4(n4355), .Y(n3248) );
  AO22X1_HVT U968 ( .A1(n4370), .A2(keyout[100]), .A3(\keys[3][100] ), .A4(
        n4355), .Y(n3249) );
  AO22X1_HVT U969 ( .A1(n4370), .A2(keyout[101]), .A3(\keys[3][101] ), .A4(
        n4355), .Y(n3250) );
  AO22X1_HVT U970 ( .A1(n4370), .A2(keyout[102]), .A3(\keys[3][102] ), .A4(
        n4355), .Y(n3251) );
  AO22X1_HVT U971 ( .A1(n4371), .A2(keyout[103]), .A3(\keys[3][103] ), .A4(
        n4355), .Y(n3252) );
  AO22X1_HVT U972 ( .A1(n4371), .A2(keyout[104]), .A3(\keys[3][104] ), .A4(
        n4354), .Y(n3253) );
  AO22X1_HVT U973 ( .A1(n4371), .A2(keyout[105]), .A3(\keys[3][105] ), .A4(
        n4354), .Y(n3254) );
  AO22X1_HVT U974 ( .A1(n4371), .A2(n3880), .A3(\keys[3][106] ), .A4(n4354), 
        .Y(n3255) );
  AO22X1_HVT U975 ( .A1(n4371), .A2(n3820), .A3(\keys[3][107] ), .A4(n4354), 
        .Y(n3256) );
  AO22X1_HVT U976 ( .A1(n4371), .A2(n3892), .A3(\keys[3][108] ), .A4(n4354), 
        .Y(n3257) );
  AO22X1_HVT U977 ( .A1(n4371), .A2(n3873), .A3(\keys[3][109] ), .A4(n4354), 
        .Y(n3258) );
  AO22X1_HVT U978 ( .A1(n4371), .A2(keyout[110]), .A3(\keys[3][110] ), .A4(
        n4354), .Y(n3259) );
  AO22X1_HVT U979 ( .A1(n4371), .A2(keyout[111]), .A3(\keys[3][111] ), .A4(
        n4354), .Y(n3260) );
  AO22X1_HVT U980 ( .A1(n4371), .A2(keyout[112]), .A3(\keys[3][112] ), .A4(
        n4354), .Y(n3261) );
  AO22X1_HVT U981 ( .A1(n4371), .A2(keyout[113]), .A3(\keys[3][113] ), .A4(
        n4354), .Y(n3262) );
  AO22X1_HVT U982 ( .A1(n4371), .A2(keyout[114]), .A3(\keys[3][114] ), .A4(
        n4354), .Y(n3263) );
  AO22X1_HVT U983 ( .A1(n4371), .A2(n3915), .A3(\keys[3][115] ), .A4(n4354), 
        .Y(n3264) );
  AO22X1_HVT U984 ( .A1(n4371), .A2(keyout[116]), .A3(\keys[3][116] ), .A4(
        n4354), .Y(n3265) );
  AO22X1_HVT U985 ( .A1(n4371), .A2(keyout[117]), .A3(\keys[3][117] ), .A4(
        n4353), .Y(n3266) );
  AO22X1_HVT U986 ( .A1(n4371), .A2(keyout[118]), .A3(\keys[3][118] ), .A4(
        n4353), .Y(n3267) );
  AO22X1_HVT U987 ( .A1(n4372), .A2(keyout[119]), .A3(\keys[3][119] ), .A4(
        n4353), .Y(n3268) );
  AO22X1_HVT U988 ( .A1(n4372), .A2(n4096), .A3(\keys[3][120] ), .A4(n4353), 
        .Y(n3269) );
  AO22X1_HVT U989 ( .A1(n4372), .A2(keyout[121]), .A3(\keys[3][121] ), .A4(
        n4353), .Y(n3270) );
  AO22X1_HVT U990 ( .A1(n4372), .A2(keyout[122]), .A3(\keys[3][122] ), .A4(
        n4353), .Y(n3271) );
  AO22X1_HVT U991 ( .A1(n4372), .A2(n3809), .A3(\keys[3][123] ), .A4(n4353), 
        .Y(n3272) );
  AO22X1_HVT U992 ( .A1(n4372), .A2(n3844), .A3(\keys[3][124] ), .A4(n4353), 
        .Y(n3273) );
  AO22X1_HVT U993 ( .A1(n4372), .A2(keyout[125]), .A3(\keys[3][125] ), .A4(
        n4353), .Y(n3274) );
  AO22X1_HVT U994 ( .A1(n4372), .A2(n4099), .A3(\keys[3][126] ), .A4(n4353), 
        .Y(n3275) );
  AO22X1_HVT U995 ( .A1(n4372), .A2(n4102), .A3(\keys[3][127] ), .A4(n4353), 
        .Y(n3276) );
  AO22X1_HVT U996 ( .A1(n4341), .A2(n3998), .A3(\keys[2][0] ), .A4(n4340), .Y(
        n3277) );
  AO22X1_HVT U997 ( .A1(n4342), .A2(n4001), .A3(\keys[2][1] ), .A4(n4340), .Y(
        n3278) );
  AO22X1_HVT U998 ( .A1(n4342), .A2(keyout[2]), .A3(\keys[2][2] ), .A4(n4340), 
        .Y(n3279) );
  AO22X1_HVT U999 ( .A1(n4342), .A2(n4005), .A3(\keys[2][3] ), .A4(n4340), .Y(
        n3280) );
  AO22X1_HVT U1000 ( .A1(n4342), .A2(n4008), .A3(\keys[2][4] ), .A4(n4340), 
        .Y(n3281) );
  AO22X1_HVT U1001 ( .A1(n4342), .A2(n4011), .A3(\keys[2][5] ), .A4(n4340), 
        .Y(n3282) );
  AO22X1_HVT U1002 ( .A1(n4342), .A2(n4014), .A3(\keys[2][6] ), .A4(n4340), 
        .Y(n3283) );
  AO22X1_HVT U1003 ( .A1(n4343), .A2(n4016), .A3(\keys[2][7] ), .A4(n4340), 
        .Y(n3284) );
  AO22X1_HVT U1004 ( .A1(n4343), .A2(n4018), .A3(\keys[2][8] ), .A4(n4340), 
        .Y(n3285) );
  AO22X1_HVT U1005 ( .A1(n4343), .A2(n4021), .A3(\keys[2][9] ), .A4(n4340), 
        .Y(n3286) );
  AO22X1_HVT U1006 ( .A1(n4343), .A2(n4024), .A3(\keys[2][10] ), .A4(n4340), 
        .Y(n3287) );
  AO22X1_HVT U1007 ( .A1(n4343), .A2(n4027), .A3(\keys[2][11] ), .A4(n4340), 
        .Y(n3288) );
  AO22X1_HVT U1008 ( .A1(n4343), .A2(n4030), .A3(\keys[2][12] ), .A4(n4339), 
        .Y(n3289) );
  AO22X1_HVT U1009 ( .A1(n4343), .A2(n4033), .A3(\keys[2][13] ), .A4(n4339), 
        .Y(n3290) );
  AO22X1_HVT U1010 ( .A1(n4343), .A2(n4036), .A3(\keys[2][14] ), .A4(n4339), 
        .Y(n3291) );
  AO22X1_HVT U1011 ( .A1(n4343), .A2(n4039), .A3(\keys[2][15] ), .A4(n4339), 
        .Y(n3292) );
  AO22X1_HVT U1012 ( .A1(n4343), .A2(n4042), .A3(\keys[2][16] ), .A4(n4339), 
        .Y(n3293) );
  AO22X1_HVT U1013 ( .A1(n4343), .A2(n4045), .A3(\keys[2][17] ), .A4(n4339), 
        .Y(n3294) );
  AO22X1_HVT U1014 ( .A1(n4343), .A2(n4048), .A3(\keys[2][18] ), .A4(n4339), 
        .Y(n3295) );
  AO22X1_HVT U1015 ( .A1(n4343), .A2(n4051), .A3(\keys[2][19] ), .A4(n4339), 
        .Y(n3296) );
  AO22X1_HVT U1016 ( .A1(n4343), .A2(n4054), .A3(\keys[2][20] ), .A4(n4339), 
        .Y(n3297) );
  AO22X1_HVT U1017 ( .A1(n4343), .A2(n4057), .A3(\keys[2][21] ), .A4(n4339), 
        .Y(n3298) );
  AO22X1_HVT U1018 ( .A1(n4343), .A2(n4060), .A3(\keys[2][22] ), .A4(n4339), 
        .Y(n3299) );
  AO22X1_HVT U1019 ( .A1(n4344), .A2(n4063), .A3(\keys[2][23] ), .A4(n4339), 
        .Y(n3300) );
  AO22X1_HVT U1020 ( .A1(n4344), .A2(n4066), .A3(\keys[2][24] ), .A4(n4339), 
        .Y(n3301) );
  AO22X1_HVT U1021 ( .A1(n4344), .A2(n4068), .A3(\keys[2][25] ), .A4(n4338), 
        .Y(n3302) );
  AO22X1_HVT U1022 ( .A1(n4344), .A2(n4071), .A3(\keys[2][26] ), .A4(n4338), 
        .Y(n3303) );
  AO22X1_HVT U1023 ( .A1(n4344), .A2(n4074), .A3(\keys[2][27] ), .A4(n4338), 
        .Y(n3304) );
  AO22X1_HVT U1024 ( .A1(n4344), .A2(n4077), .A3(\keys[2][28] ), .A4(n4338), 
        .Y(n3305) );
  AO22X1_HVT U1025 ( .A1(n4344), .A2(n4080), .A3(\keys[2][29] ), .A4(n4338), 
        .Y(n3306) );
  AO22X1_HVT U1026 ( .A1(n4344), .A2(n4082), .A3(\keys[2][30] ), .A4(n4338), 
        .Y(n3307) );
  AO22X1_HVT U1027 ( .A1(n4344), .A2(n3852), .A3(\keys[2][31] ), .A4(n4338), 
        .Y(n3308) );
  AO22X1_HVT U1028 ( .A1(n4344), .A2(keyout[32]), .A3(\keys[2][32] ), .A4(
        n4338), .Y(n3309) );
  AO22X1_HVT U1029 ( .A1(n4344), .A2(n3876), .A3(\keys[2][33] ), .A4(n4338), 
        .Y(n3310) );
  AO22X1_HVT U1030 ( .A1(n4344), .A2(n3913), .A3(\keys[2][34] ), .A4(n4338), 
        .Y(n3311) );
  AO22X1_HVT U1031 ( .A1(n4344), .A2(keyout[35]), .A3(\keys[2][35] ), .A4(
        n4338), .Y(n3312) );
  AO22X1_HVT U1032 ( .A1(n4344), .A2(keyout[36]), .A3(\keys[2][36] ), .A4(
        n4338), .Y(n3313) );
  AO22X1_HVT U1033 ( .A1(n4344), .A2(n3819), .A3(\keys[2][37] ), .A4(n4338), 
        .Y(n3314) );
  AO22X1_HVT U1034 ( .A1(n4344), .A2(keyout[38]), .A3(\keys[2][38] ), .A4(
        n4337), .Y(n3315) );
  AO22X1_HVT U1035 ( .A1(n4345), .A2(keyout[39]), .A3(\keys[2][39] ), .A4(
        n4337), .Y(n3316) );
  AO22X1_HVT U1036 ( .A1(n4345), .A2(n3953), .A3(\keys[2][40] ), .A4(n4337), 
        .Y(n3317) );
  AO22X1_HVT U1038 ( .A1(n4345), .A2(n3974), .A3(\keys[2][42] ), .A4(n4337), 
        .Y(n3319) );
  AO22X1_HVT U1039 ( .A1(n4345), .A2(n3890), .A3(\keys[2][43] ), .A4(n4337), 
        .Y(n3320) );
  AO22X1_HVT U1040 ( .A1(n4345), .A2(n3902), .A3(\keys[2][44] ), .A4(n4337), 
        .Y(n3321) );
  AO22X1_HVT U1042 ( .A1(n4345), .A2(n3945), .A3(\keys[2][46] ), .A4(n4337), 
        .Y(n3323) );
  AO22X1_HVT U1044 ( .A1(n4345), .A2(keyout[48]), .A3(\keys[2][48] ), .A4(
        n4337), .Y(n3325) );
  AO22X1_HVT U1045 ( .A1(n4345), .A2(keyout[49]), .A3(\keys[2][49] ), .A4(
        n4337), .Y(n3326) );
  AO22X1_HVT U1046 ( .A1(n4345), .A2(keyout[50]), .A3(\keys[2][50] ), .A4(
        n4337), .Y(n3327) );
  AO22X1_HVT U1047 ( .A1(n4345), .A2(n3937), .A3(\keys[2][51] ), .A4(n4336), 
        .Y(n3328) );
  AO22X1_HVT U1048 ( .A1(n4345), .A2(keyout[52]), .A3(\keys[2][52] ), .A4(
        n4336), .Y(n3329) );
  AO22X1_HVT U1049 ( .A1(n4345), .A2(n3920), .A3(\keys[2][53] ), .A4(n4336), 
        .Y(n3330) );
  AO22X1_HVT U1050 ( .A1(n4345), .A2(keyout[54]), .A3(\keys[2][54] ), .A4(
        n4336), .Y(n3331) );
  AO22X1_HVT U1051 ( .A1(n4346), .A2(n3922), .A3(\keys[2][55] ), .A4(n4336), 
        .Y(n3332) );
  AO22X1_HVT U1052 ( .A1(n4346), .A2(n3941), .A3(\keys[2][56] ), .A4(n4336), 
        .Y(n3333) );
  AO22X1_HVT U1053 ( .A1(n4346), .A2(n4085), .A3(\keys[2][57] ), .A4(n4336), 
        .Y(n3334) );
  AO22X1_HVT U1054 ( .A1(n4346), .A2(n4087), .A3(\keys[2][58] ), .A4(n4336), 
        .Y(n3335) );
  AO22X1_HVT U1055 ( .A1(n4346), .A2(n4090), .A3(\keys[2][59] ), .A4(n4336), 
        .Y(n3336) );
  AO22X1_HVT U1056 ( .A1(n4346), .A2(n3943), .A3(\keys[2][60] ), .A4(n4336), 
        .Y(n3337) );
  AO22X1_HVT U1057 ( .A1(n4346), .A2(n3805), .A3(\keys[2][61] ), .A4(n4336), 
        .Y(n3338) );
  AO22X1_HVT U1058 ( .A1(n4346), .A2(n3833), .A3(\keys[2][62] ), .A4(n4336), 
        .Y(n3339) );
  AO22X1_HVT U1059 ( .A1(n4346), .A2(n3861), .A3(\keys[2][63] ), .A4(n4336), 
        .Y(n3340) );
  AO22X1_HVT U1060 ( .A1(n4346), .A2(keyout[64]), .A3(\keys[2][64] ), .A4(
        n4335), .Y(n3341) );
  AO22X1_HVT U1061 ( .A1(n4346), .A2(n3883), .A3(\keys[2][65] ), .A4(n4335), 
        .Y(n3342) );
  AO22X1_HVT U1062 ( .A1(n4346), .A2(n3914), .A3(\keys[2][66] ), .A4(n4335), 
        .Y(n3343) );
  AO22X1_HVT U1063 ( .A1(n4346), .A2(n3938), .A3(\keys[2][67] ), .A4(n4335), 
        .Y(n3344) );
  AO22X1_HVT U1064 ( .A1(n4346), .A2(keyout[68]), .A3(\keys[2][68] ), .A4(
        n4335), .Y(n3345) );
  AO22X1_HVT U1065 ( .A1(n4346), .A2(keyout[69]), .A3(\keys[2][69] ), .A4(
        n4335), .Y(n3346) );
  AO22X1_HVT U1066 ( .A1(n4346), .A2(keyout[70]), .A3(\keys[2][70] ), .A4(
        n4335), .Y(n3347) );
  AO22X1_HVT U1067 ( .A1(n4347), .A2(keyout[71]), .A3(\keys[2][71] ), .A4(
        n4335), .Y(n3348) );
  AO22X1_HVT U1068 ( .A1(n4347), .A2(n3951), .A3(\keys[2][72] ), .A4(n4335), 
        .Y(n3349) );
  AO22X1_HVT U1069 ( .A1(n4347), .A2(n3896), .A3(\keys[2][73] ), .A4(n4335), 
        .Y(n3350) );
  AO22X1_HVT U1070 ( .A1(n4347), .A2(n3979), .A3(\keys[2][74] ), .A4(n4335), 
        .Y(n3351) );
  AO22X1_HVT U1071 ( .A1(n4347), .A2(n3960), .A3(\keys[2][75] ), .A4(n4335), 
        .Y(n3352) );
  AO22X1_HVT U1072 ( .A1(n4347), .A2(n3967), .A3(\keys[2][76] ), .A4(n4335), 
        .Y(n3353) );
  AO22X1_HVT U1073 ( .A1(n4347), .A2(n3986), .A3(\keys[2][77] ), .A4(n4334), 
        .Y(n3354) );
  AO22X1_HVT U1074 ( .A1(n4347), .A2(n3947), .A3(\keys[2][78] ), .A4(n4334), 
        .Y(n3355) );
  AO22X1_HVT U1075 ( .A1(n4347), .A2(n3898), .A3(\keys[2][79] ), .A4(n4334), 
        .Y(n3356) );
  AO22X1_HVT U1076 ( .A1(n4347), .A2(n3931), .A3(\keys[2][80] ), .A4(n4334), 
        .Y(n3357) );
  AO22X1_HVT U1077 ( .A1(n4347), .A2(n3811), .A3(\keys[2][81] ), .A4(n4334), 
        .Y(n3358) );
  AO22X1_HVT U1078 ( .A1(n4347), .A2(n3977), .A3(\keys[2][82] ), .A4(n4334), 
        .Y(n3359) );
  AO22X1_HVT U1079 ( .A1(n4347), .A2(n3916), .A3(\keys[2][83] ), .A4(n4334), 
        .Y(n3360) );
  AO22X1_HVT U1080 ( .A1(n4347), .A2(n1438), .A3(\keys[2][84] ), .A4(n4334), 
        .Y(n3361) );
  AO22X1_HVT U1081 ( .A1(n4347), .A2(n2), .A3(\keys[2][85] ), .A4(n4334), .Y(
        n3362) );
  AO22X1_HVT U1082 ( .A1(n4347), .A2(n1436), .A3(\keys[2][86] ), .A4(n4334), 
        .Y(n3363) );
  AO22X1_HVT U1083 ( .A1(n4348), .A2(n1440), .A3(\keys[2][87] ), .A4(n4334), 
        .Y(n3364) );
  AO22X1_HVT U1084 ( .A1(n4348), .A2(n4093), .A3(\keys[2][88] ), .A4(n4334), 
        .Y(n3365) );
  AO22X1_HVT U1085 ( .A1(n4348), .A2(n3863), .A3(\keys[2][89] ), .A4(n4334), 
        .Y(n3366) );
  AO22X1_HVT U1086 ( .A1(n4348), .A2(n3949), .A3(\keys[2][90] ), .A4(n4333), 
        .Y(n3367) );
  AO22X1_HVT U1087 ( .A1(n4348), .A2(n3816), .A3(\keys[2][91] ), .A4(n4333), 
        .Y(n3368) );
  AO22X1_HVT U1088 ( .A1(n4348), .A2(n3831), .A3(\keys[2][92] ), .A4(n4333), 
        .Y(n3369) );
  AO22X1_HVT U1089 ( .A1(n4348), .A2(keyout[93]), .A3(\keys[2][93] ), .A4(
        n4333), .Y(n3370) );
  AO22X1_HVT U1090 ( .A1(n4348), .A2(n3835), .A3(\keys[2][94] ), .A4(n4333), 
        .Y(n3371) );
  AO22X1_HVT U1091 ( .A1(n4348), .A2(n3869), .A3(\keys[2][95] ), .A4(n4333), 
        .Y(n3372) );
  AO22X1_HVT U1092 ( .A1(n4348), .A2(keyout[96]), .A3(\keys[2][96] ), .A4(
        n4333), .Y(n3373) );
  AO22X1_HVT U1093 ( .A1(n4348), .A2(keyout[97]), .A3(\keys[2][97] ), .A4(
        n4333), .Y(n3374) );
  AO22X1_HVT U1094 ( .A1(n4348), .A2(keyout[98]), .A3(\keys[2][98] ), .A4(
        n4333), .Y(n3375) );
  AO22X1_HVT U1095 ( .A1(n4348), .A2(keyout[99]), .A3(\keys[2][99] ), .A4(
        n4333), .Y(n3376) );
  AO22X1_HVT U1096 ( .A1(n4348), .A2(keyout[100]), .A3(\keys[2][100] ), .A4(
        n4333), .Y(n3377) );
  AO22X1_HVT U1097 ( .A1(n4348), .A2(keyout[101]), .A3(\keys[2][101] ), .A4(
        n4333), .Y(n3378) );
  AO22X1_HVT U1098 ( .A1(n4348), .A2(keyout[102]), .A3(\keys[2][102] ), .A4(
        n4333), .Y(n3379) );
  AO22X1_HVT U1099 ( .A1(n4349), .A2(keyout[103]), .A3(\keys[2][103] ), .A4(
        n4332), .Y(n3380) );
  AO22X1_HVT U1100 ( .A1(n4349), .A2(keyout[104]), .A3(\keys[2][104] ), .A4(
        n4332), .Y(n3381) );
  AO22X1_HVT U1101 ( .A1(n4349), .A2(keyout[105]), .A3(\keys[2][105] ), .A4(
        n4332), .Y(n3382) );
  AO22X1_HVT U1102 ( .A1(n4349), .A2(n3880), .A3(\keys[2][106] ), .A4(n4332), 
        .Y(n3383) );
  AO22X1_HVT U1103 ( .A1(n4349), .A2(n3820), .A3(\keys[2][107] ), .A4(n4332), 
        .Y(n3384) );
  AO22X1_HVT U1104 ( .A1(n4349), .A2(n3892), .A3(\keys[2][108] ), .A4(n4332), 
        .Y(n3385) );
  AO22X1_HVT U1105 ( .A1(n4349), .A2(n3873), .A3(\keys[2][109] ), .A4(n4332), 
        .Y(n3386) );
  AO22X1_HVT U1106 ( .A1(n4349), .A2(keyout[110]), .A3(\keys[2][110] ), .A4(
        n4332), .Y(n3387) );
  AO22X1_HVT U1107 ( .A1(n4349), .A2(keyout[111]), .A3(\keys[2][111] ), .A4(
        n4332), .Y(n3388) );
  AO22X1_HVT U1108 ( .A1(n4349), .A2(keyout[112]), .A3(\keys[2][112] ), .A4(
        n4332), .Y(n3389) );
  AO22X1_HVT U1109 ( .A1(n4349), .A2(keyout[113]), .A3(\keys[2][113] ), .A4(
        n4332), .Y(n3390) );
  AO22X1_HVT U1110 ( .A1(n4349), .A2(keyout[114]), .A3(\keys[2][114] ), .A4(
        n4332), .Y(n3391) );
  AO22X1_HVT U1111 ( .A1(n4349), .A2(n3915), .A3(\keys[2][115] ), .A4(n4332), 
        .Y(n3392) );
  AO22X1_HVT U1112 ( .A1(n4349), .A2(keyout[116]), .A3(\keys[2][116] ), .A4(
        n4331), .Y(n3393) );
  AO22X1_HVT U1113 ( .A1(n4349), .A2(keyout[117]), .A3(\keys[2][117] ), .A4(
        n4331), .Y(n3394) );
  AO22X1_HVT U1114 ( .A1(n4349), .A2(keyout[118]), .A3(\keys[2][118] ), .A4(
        n4331), .Y(n3395) );
  AO22X1_HVT U1115 ( .A1(n4350), .A2(keyout[119]), .A3(\keys[2][119] ), .A4(
        n4331), .Y(n3396) );
  AO22X1_HVT U1116 ( .A1(n4350), .A2(n4096), .A3(\keys[2][120] ), .A4(n4331), 
        .Y(n3397) );
  AO22X1_HVT U1117 ( .A1(n4350), .A2(keyout[121]), .A3(\keys[2][121] ), .A4(
        n4331), .Y(n3398) );
  AO22X1_HVT U1118 ( .A1(n4350), .A2(keyout[122]), .A3(\keys[2][122] ), .A4(
        n4331), .Y(n3399) );
  AO22X1_HVT U1119 ( .A1(n4350), .A2(n3809), .A3(\keys[2][123] ), .A4(n4331), 
        .Y(n3400) );
  AO22X1_HVT U1120 ( .A1(n4350), .A2(n3845), .A3(\keys[2][124] ), .A4(n4331), 
        .Y(n3401) );
  AO22X1_HVT U1121 ( .A1(n4350), .A2(keyout[125]), .A3(\keys[2][125] ), .A4(
        n4331), .Y(n3402) );
  AO22X1_HVT U1122 ( .A1(n4350), .A2(n4099), .A3(\keys[2][126] ), .A4(n4331), 
        .Y(n3403) );
  AO22X1_HVT U1123 ( .A1(n4350), .A2(n4102), .A3(\keys[2][127] ), .A4(n4331), 
        .Y(n3404) );
  AO22X1_HVT U1124 ( .A1(n4319), .A2(n3998), .A3(\keys[1][0] ), .A4(n4308), 
        .Y(n3405) );
  AO22X1_HVT U1125 ( .A1(n4320), .A2(n4001), .A3(\keys[1][1] ), .A4(n4308), 
        .Y(n3406) );
  AO22X1_HVT U1126 ( .A1(n4320), .A2(keyout[2]), .A3(\keys[1][2] ), .A4(n4308), 
        .Y(n3407) );
  AO22X1_HVT U1127 ( .A1(n4320), .A2(n4005), .A3(\keys[1][3] ), .A4(n4308), 
        .Y(n3408) );
  AO22X1_HVT U1128 ( .A1(n4321), .A2(n4008), .A3(\keys[1][4] ), .A4(n4308), 
        .Y(n3409) );
  AO22X1_HVT U1129 ( .A1(n4321), .A2(n4011), .A3(\keys[1][5] ), .A4(n4308), 
        .Y(n3410) );
  AO22X1_HVT U1130 ( .A1(n4321), .A2(n4014), .A3(\keys[1][6] ), .A4(n4308), 
        .Y(n3411) );
  AO22X1_HVT U1131 ( .A1(n4321), .A2(keyout[7]), .A3(\keys[1][7] ), .A4(n4308), 
        .Y(n3412) );
  AO22X1_HVT U1132 ( .A1(n4321), .A2(n4018), .A3(\keys[1][8] ), .A4(n4308), 
        .Y(n3413) );
  AO22X1_HVT U1133 ( .A1(n4321), .A2(n4021), .A3(\keys[1][9] ), .A4(n4308), 
        .Y(n3414) );
  AO22X1_HVT U1134 ( .A1(n4321), .A2(n4024), .A3(\keys[1][10] ), .A4(n4308), 
        .Y(n3415) );
  AO22X1_HVT U1135 ( .A1(n4321), .A2(n4027), .A3(\keys[1][11] ), .A4(n4308), 
        .Y(n3416) );
  AO22X1_HVT U1136 ( .A1(n4321), .A2(n4030), .A3(\keys[1][12] ), .A4(n4309), 
        .Y(n3417) );
  AO22X1_HVT U1137 ( .A1(n4321), .A2(n4033), .A3(\keys[1][13] ), .A4(n4309), 
        .Y(n3418) );
  AO22X1_HVT U1138 ( .A1(n4321), .A2(n4036), .A3(\keys[1][14] ), .A4(n4309), 
        .Y(n3419) );
  AO22X1_HVT U1139 ( .A1(n4321), .A2(n4039), .A3(\keys[1][15] ), .A4(n4309), 
        .Y(n3420) );
  AO22X1_HVT U1140 ( .A1(n4321), .A2(n4042), .A3(\keys[1][16] ), .A4(n4309), 
        .Y(n3421) );
  AO22X1_HVT U1141 ( .A1(n4321), .A2(n4045), .A3(\keys[1][17] ), .A4(n4309), 
        .Y(n3422) );
  AO22X1_HVT U1142 ( .A1(n4321), .A2(n4048), .A3(\keys[1][18] ), .A4(n4309), 
        .Y(n3423) );
  AO22X1_HVT U1143 ( .A1(n4321), .A2(n4051), .A3(\keys[1][19] ), .A4(n4309), 
        .Y(n3424) );
  AO22X1_HVT U1144 ( .A1(n4322), .A2(n4054), .A3(\keys[1][20] ), .A4(n4309), 
        .Y(n3425) );
  AO22X1_HVT U1145 ( .A1(n4322), .A2(n4057), .A3(\keys[1][21] ), .A4(n4309), 
        .Y(n3426) );
  AO22X1_HVT U1146 ( .A1(n4322), .A2(n4060), .A3(\keys[1][22] ), .A4(n4309), 
        .Y(n3427) );
  AO22X1_HVT U1147 ( .A1(n4322), .A2(n4063), .A3(\keys[1][23] ), .A4(n4309), 
        .Y(n3428) );
  AO22X1_HVT U1148 ( .A1(n4322), .A2(n4066), .A3(\keys[1][24] ), .A4(n4310), 
        .Y(n3429) );
  AO22X1_HVT U1149 ( .A1(n4322), .A2(n4068), .A3(\keys[1][25] ), .A4(n4310), 
        .Y(n3430) );
  AO22X1_HVT U1150 ( .A1(n4322), .A2(n4071), .A3(\keys[1][26] ), .A4(n4310), 
        .Y(n3431) );
  AO22X1_HVT U1151 ( .A1(n4322), .A2(n4074), .A3(\keys[1][27] ), .A4(n4310), 
        .Y(n3432) );
  AO22X1_HVT U1152 ( .A1(n4322), .A2(n4077), .A3(\keys[1][28] ), .A4(n4310), 
        .Y(n3433) );
  AO22X1_HVT U1153 ( .A1(n4322), .A2(n4080), .A3(\keys[1][29] ), .A4(n4310), 
        .Y(n3434) );
  AO22X1_HVT U1154 ( .A1(n4322), .A2(keyout[30]), .A3(\keys[1][30] ), .A4(
        n4310), .Y(n3435) );
  AO22X1_HVT U1155 ( .A1(n4322), .A2(n3852), .A3(\keys[1][31] ), .A4(n4310), 
        .Y(n3436) );
  AO22X1_HVT U1156 ( .A1(n4322), .A2(keyout[32]), .A3(\keys[1][32] ), .A4(
        n4310), .Y(n3437) );
  AO22X1_HVT U1157 ( .A1(n4322), .A2(n3876), .A3(\keys[1][33] ), .A4(n4310), 
        .Y(n3438) );
  AO22X1_HVT U1158 ( .A1(n4322), .A2(n3913), .A3(\keys[1][34] ), .A4(n4310), 
        .Y(n3439) );
  AO22X1_HVT U1159 ( .A1(n4322), .A2(keyout[35]), .A3(\keys[1][35] ), .A4(
        n4310), .Y(n3440) );
  AO22X1_HVT U1160 ( .A1(n4323), .A2(keyout[36]), .A3(\keys[1][36] ), .A4(
        n4311), .Y(n3441) );
  AO22X1_HVT U1161 ( .A1(n4323), .A2(n3911), .A3(\keys[1][37] ), .A4(n4311), 
        .Y(n3442) );
  AO22X1_HVT U1162 ( .A1(n4323), .A2(keyout[38]), .A3(\keys[1][38] ), .A4(
        n4311), .Y(n3443) );
  AO22X1_HVT U1163 ( .A1(n4323), .A2(keyout[39]), .A3(\keys[1][39] ), .A4(
        n4311), .Y(n3444) );
  AO22X1_HVT U1164 ( .A1(n4323), .A2(n3952), .A3(\keys[1][40] ), .A4(n4311), 
        .Y(n3445) );
  AO22X1_HVT U1165 ( .A1(n4323), .A2(n3854), .A3(\keys[1][41] ), .A4(n4311), 
        .Y(n3446) );
  AO22X1_HVT U1168 ( .A1(n4323), .A2(n3902), .A3(\keys[1][44] ), .A4(n4311), 
        .Y(n3449) );
  AO22X1_HVT U1169 ( .A1(n4323), .A2(n3935), .A3(\keys[1][45] ), .A4(n4311), 
        .Y(n3450) );
  AO22X1_HVT U1170 ( .A1(n4323), .A2(n3944), .A3(\keys[1][46] ), .A4(n4311), 
        .Y(n3451) );
  AO22X1_HVT U1171 ( .A1(n4323), .A2(n3850), .A3(\keys[1][47] ), .A4(n4311), 
        .Y(n3452) );
  AO22X1_HVT U1172 ( .A1(n4323), .A2(keyout[48]), .A3(\keys[1][48] ), .A4(
        n4312), .Y(n3453) );
  AO22X1_HVT U1173 ( .A1(n4323), .A2(keyout[49]), .A3(\keys[1][49] ), .A4(
        n4312), .Y(n3454) );
  AO22X1_HVT U1174 ( .A1(n4323), .A2(keyout[50]), .A3(\keys[1][50] ), .A4(
        n4312), .Y(n3455) );
  AO22X1_HVT U1175 ( .A1(n4323), .A2(n3937), .A3(\keys[1][51] ), .A4(n4312), 
        .Y(n3456) );
  AO22X1_HVT U1176 ( .A1(n4324), .A2(n1434), .A3(\keys[1][52] ), .A4(n4312), 
        .Y(n3457) );
  AO22X1_HVT U1177 ( .A1(n4324), .A2(n3920), .A3(\keys[1][53] ), .A4(n4312), 
        .Y(n3458) );
  AO22X1_HVT U1178 ( .A1(n4324), .A2(n13), .A3(\keys[1][54] ), .A4(n4312), .Y(
        n3459) );
  AO22X1_HVT U1179 ( .A1(n4324), .A2(n3922), .A3(\keys[1][55] ), .A4(n4312), 
        .Y(n3460) );
  AO22X1_HVT U1180 ( .A1(n4324), .A2(n3941), .A3(\keys[1][56] ), .A4(n4312), 
        .Y(n3461) );
  AO22X1_HVT U1181 ( .A1(n4324), .A2(n4085), .A3(\keys[1][57] ), .A4(n4312), 
        .Y(n3462) );
  AO22X1_HVT U1182 ( .A1(n4324), .A2(n4087), .A3(\keys[1][58] ), .A4(n4312), 
        .Y(n3463) );
  AO22X1_HVT U1183 ( .A1(n4324), .A2(n4090), .A3(\keys[1][59] ), .A4(n4312), 
        .Y(n3464) );
  AO22X1_HVT U1184 ( .A1(n4324), .A2(n3943), .A3(\keys[1][60] ), .A4(n4313), 
        .Y(n3465) );
  AO22X1_HVT U1185 ( .A1(n4324), .A2(n3805), .A3(\keys[1][61] ), .A4(n4313), 
        .Y(n3466) );
  AO22X1_HVT U1186 ( .A1(n4324), .A2(n3832), .A3(\keys[1][62] ), .A4(n4313), 
        .Y(n3467) );
  AO22X1_HVT U1187 ( .A1(n4324), .A2(n3860), .A3(\keys[1][63] ), .A4(n4313), 
        .Y(n3468) );
  AO22X1_HVT U1188 ( .A1(n4324), .A2(keyout[64]), .A3(\keys[1][64] ), .A4(
        n4313), .Y(n3469) );
  AO22X1_HVT U1189 ( .A1(n4324), .A2(n3883), .A3(\keys[1][65] ), .A4(n4313), 
        .Y(n3470) );
  AO22X1_HVT U1190 ( .A1(n4324), .A2(n3914), .A3(\keys[1][66] ), .A4(n4313), 
        .Y(n3471) );
  AO22X1_HVT U1191 ( .A1(n4324), .A2(n3825), .A3(\keys[1][67] ), .A4(n4313), 
        .Y(n3472) );
  AO22X1_HVT U1192 ( .A1(n4325), .A2(keyout[68]), .A3(\keys[1][68] ), .A4(
        n4313), .Y(n3473) );
  AO22X1_HVT U1193 ( .A1(n4325), .A2(keyout[69]), .A3(\keys[1][69] ), .A4(
        n4313), .Y(n3474) );
  AO22X1_HVT U1194 ( .A1(n4325), .A2(keyout[70]), .A3(\keys[1][70] ), .A4(
        n4313), .Y(n3475) );
  AO22X1_HVT U1195 ( .A1(n4325), .A2(keyout[71]), .A3(\keys[1][71] ), .A4(
        n4313), .Y(n3476) );
  AO22X1_HVT U1196 ( .A1(n4325), .A2(n3939), .A3(\keys[1][72] ), .A4(n4314), 
        .Y(n3477) );
  AO22X1_HVT U1197 ( .A1(n4325), .A2(n3886), .A3(\keys[1][73] ), .A4(n4314), 
        .Y(n3478) );
  AO22X1_HVT U1198 ( .A1(n4325), .A2(n3872), .A3(\keys[1][74] ), .A4(n4314), 
        .Y(n3479) );
  AO22X1_HVT U1199 ( .A1(n4325), .A2(keyout[75]), .A3(\keys[1][75] ), .A4(
        n4314), .Y(n3480) );
  AO22X1_HVT U1200 ( .A1(n4325), .A2(n3965), .A3(\keys[1][76] ), .A4(n4314), 
        .Y(n3481) );
  AO22X1_HVT U1201 ( .A1(n4325), .A2(n3984), .A3(\keys[1][77] ), .A4(n4314), 
        .Y(n3482) );
  AO22X1_HVT U1202 ( .A1(n4325), .A2(n3947), .A3(\keys[1][78] ), .A4(n4314), 
        .Y(n3483) );
  AO22X1_HVT U1203 ( .A1(n4325), .A2(n3887), .A3(\keys[1][79] ), .A4(n4314), 
        .Y(n3484) );
  AO22X1_HVT U1204 ( .A1(n4325), .A2(keyout[80]), .A3(\keys[1][80] ), .A4(
        n4314), .Y(n3485) );
  AO22X1_HVT U1205 ( .A1(n4325), .A2(keyout[81]), .A3(\keys[1][81] ), .A4(
        n4314), .Y(n3486) );
  AO22X1_HVT U1206 ( .A1(n4325), .A2(n3905), .A3(\keys[1][82] ), .A4(n4314), 
        .Y(n3487) );
  AO22X1_HVT U1207 ( .A1(n4325), .A2(n3904), .A3(\keys[1][83] ), .A4(n4314), 
        .Y(n3488) );
  AO22X1_HVT U1208 ( .A1(n4326), .A2(keyout[84]), .A3(\keys[1][84] ), .A4(
        n4315), .Y(n3489) );
  AO22X1_HVT U1209 ( .A1(n4326), .A2(n2), .A3(\keys[1][85] ), .A4(n4315), .Y(
        n3490) );
  AO22X1_HVT U1210 ( .A1(n4326), .A2(keyout[86]), .A3(\keys[1][86] ), .A4(
        n4315), .Y(n3491) );
  AO22X1_HVT U1211 ( .A1(n4326), .A2(n1440), .A3(\keys[1][87] ), .A4(n4315), 
        .Y(n3492) );
  AO22X1_HVT U1212 ( .A1(n4326), .A2(n4093), .A3(\keys[1][88] ), .A4(n4315), 
        .Y(n3493) );
  AO22X1_HVT U1213 ( .A1(n4326), .A2(n3827), .A3(\keys[1][89] ), .A4(n4315), 
        .Y(n3494) );
  AO22X1_HVT U1214 ( .A1(n4326), .A2(keyout[90]), .A3(\keys[1][90] ), .A4(
        n4315), .Y(n3495) );
  AO22X1_HVT U1215 ( .A1(n4326), .A2(n4), .A3(\keys[1][91] ), .A4(n4315), .Y(
        n3496) );
  AO22X1_HVT U1216 ( .A1(n4326), .A2(keyout[92]), .A3(\keys[1][92] ), .A4(
        n4315), .Y(n3497) );
  AO22X1_HVT U1217 ( .A1(n4326), .A2(keyout[93]), .A3(\keys[1][93] ), .A4(
        n4315), .Y(n3498) );
  AO22X1_HVT U1218 ( .A1(n4326), .A2(n3865), .A3(\keys[1][94] ), .A4(n4315), 
        .Y(n3499) );
  AO22X1_HVT U1219 ( .A1(n4326), .A2(n3834), .A3(\keys[1][95] ), .A4(n4315), 
        .Y(n3500) );
  AO22X1_HVT U1220 ( .A1(n4326), .A2(keyout[96]), .A3(\keys[1][96] ), .A4(
        n4316), .Y(n3501) );
  AO22X1_HVT U1221 ( .A1(n4326), .A2(keyout[97]), .A3(\keys[1][97] ), .A4(
        n4316), .Y(n3502) );
  AO22X1_HVT U1222 ( .A1(n4326), .A2(keyout[98]), .A3(\keys[1][98] ), .A4(
        n4316), .Y(n3503) );
  AO22X1_HVT U1223 ( .A1(n4326), .A2(keyout[99]), .A3(\keys[1][99] ), .A4(
        n4316), .Y(n3504) );
  AO22X1_HVT U1224 ( .A1(n4327), .A2(keyout[100]), .A3(\keys[1][100] ), .A4(
        n4316), .Y(n3505) );
  AO22X1_HVT U1225 ( .A1(n4327), .A2(keyout[101]), .A3(\keys[1][101] ), .A4(
        n4316), .Y(n3506) );
  AO22X1_HVT U1226 ( .A1(n4327), .A2(keyout[102]), .A3(\keys[1][102] ), .A4(
        n4316), .Y(n3507) );
  AO22X1_HVT U1227 ( .A1(n4327), .A2(keyout[103]), .A3(\keys[1][103] ), .A4(
        n4316), .Y(n3508) );
  AO22X1_HVT U1228 ( .A1(n4327), .A2(keyout[104]), .A3(\keys[1][104] ), .A4(
        n4316), .Y(n3509) );
  AO22X1_HVT U1229 ( .A1(n4327), .A2(keyout[105]), .A3(\keys[1][105] ), .A4(
        n4316), .Y(n3510) );
  AO22X1_HVT U1230 ( .A1(n4327), .A2(n3880), .A3(\keys[1][106] ), .A4(n4316), 
        .Y(n3511) );
  AO22X1_HVT U1231 ( .A1(n4327), .A2(keyout[107]), .A3(\keys[1][107] ), .A4(
        n4316), .Y(n3512) );
  AO22X1_HVT U1232 ( .A1(n4327), .A2(n3881), .A3(\keys[1][108] ), .A4(n4317), 
        .Y(n3513) );
  AO22X1_HVT U1233 ( .A1(n4327), .A2(keyout[109]), .A3(\keys[1][109] ), .A4(
        n4317), .Y(n3514) );
  AO22X1_HVT U1234 ( .A1(n4327), .A2(keyout[110]), .A3(\keys[1][110] ), .A4(
        n4317), .Y(n3515) );
  AO22X1_HVT U1235 ( .A1(n4327), .A2(keyout[111]), .A3(\keys[1][111] ), .A4(
        n4317), .Y(n3516) );
  AO22X1_HVT U1236 ( .A1(n4327), .A2(keyout[112]), .A3(\keys[1][112] ), .A4(
        n4317), .Y(n3517) );
  AO22X1_HVT U1237 ( .A1(n4327), .A2(keyout[113]), .A3(\keys[1][113] ), .A4(
        n4317), .Y(n3518) );
  AO22X1_HVT U1238 ( .A1(n4327), .A2(keyout[114]), .A3(\keys[1][114] ), .A4(
        n4317), .Y(n3519) );
  AO22X1_HVT U1239 ( .A1(n4327), .A2(keyout[115]), .A3(\keys[1][115] ), .A4(
        n4317), .Y(n3520) );
  AO22X1_HVT U1240 ( .A1(n4328), .A2(keyout[116]), .A3(\keys[1][116] ), .A4(
        n4317), .Y(n3521) );
  AO22X1_HVT U1241 ( .A1(n4328), .A2(keyout[117]), .A3(\keys[1][117] ), .A4(
        n4317), .Y(n3522) );
  AO22X1_HVT U1242 ( .A1(n4328), .A2(keyout[118]), .A3(\keys[1][118] ), .A4(
        n4317), .Y(n3523) );
  AO22X1_HVT U1243 ( .A1(n4328), .A2(keyout[119]), .A3(\keys[1][119] ), .A4(
        n4317), .Y(n3524) );
  AO22X1_HVT U1244 ( .A1(n4328), .A2(n4096), .A3(\keys[1][120] ), .A4(n4318), 
        .Y(n3525) );
  AO22X1_HVT U1245 ( .A1(n4328), .A2(n3829), .A3(\keys[1][121] ), .A4(n4318), 
        .Y(n3526) );
  AO22X1_HVT U1246 ( .A1(n4328), .A2(n3803), .A3(\keys[1][122] ), .A4(n4318), 
        .Y(n3527) );
  AO22X1_HVT U1247 ( .A1(n4328), .A2(n3817), .A3(\keys[1][123] ), .A4(n4318), 
        .Y(n3528) );
  AO22X1_HVT U1248 ( .A1(n4328), .A2(n3845), .A3(\keys[1][124] ), .A4(n4318), 
        .Y(n3529) );
  AO22X1_HVT U1249 ( .A1(n4328), .A2(n3823), .A3(\keys[1][125] ), .A4(n4318), 
        .Y(n3530) );
  AO22X1_HVT U1250 ( .A1(n4328), .A2(n4099), .A3(\keys[1][126] ), .A4(n4318), 
        .Y(n3531) );
  AO22X1_HVT U1251 ( .A1(n4328), .A2(n4102), .A3(\keys[1][127] ), .A4(n4318), 
        .Y(n3532) );
  AO22X1_HVT U1252 ( .A1(local_key[0]), .A2(n4295), .A3(\keys[0][0] ), .A4(
        n4294), .Y(n3533) );
  AO22X1_HVT U1253 ( .A1(local_key[1]), .A2(n4296), .A3(\keys[0][1] ), .A4(
        n4294), .Y(n3534) );
  AO22X1_HVT U1254 ( .A1(local_key[2]), .A2(n4296), .A3(\keys[0][2] ), .A4(
        n4294), .Y(n3535) );
  AO22X1_HVT U1255 ( .A1(local_key[3]), .A2(n4296), .A3(\keys[0][3] ), .A4(
        n4294), .Y(n3536) );
  AO22X1_HVT U1256 ( .A1(local_key[4]), .A2(n4296), .A3(\keys[0][4] ), .A4(
        n4294), .Y(n3537) );
  AO22X1_HVT U1257 ( .A1(local_key[5]), .A2(n4296), .A3(\keys[0][5] ), .A4(
        n4294), .Y(n3538) );
  AO22X1_HVT U1258 ( .A1(local_key[6]), .A2(n4297), .A3(\keys[0][6] ), .A4(
        n4294), .Y(n3539) );
  AO22X1_HVT U1259 ( .A1(local_key[7]), .A2(n4297), .A3(\keys[0][7] ), .A4(
        n4294), .Y(n3540) );
  AO22X1_HVT U1260 ( .A1(local_key[8]), .A2(n4297), .A3(\keys[0][8] ), .A4(
        n4294), .Y(n3541) );
  AO22X1_HVT U1261 ( .A1(local_key[9]), .A2(n4297), .A3(\keys[0][9] ), .A4(
        n4294), .Y(n3542) );
  AO22X1_HVT U1262 ( .A1(local_key[10]), .A2(n4297), .A3(\keys[0][10] ), .A4(
        n4294), .Y(n3543) );
  AO22X1_HVT U1263 ( .A1(local_key[11]), .A2(n4297), .A3(\keys[0][11] ), .A4(
        n4294), .Y(n3544) );
  AO22X1_HVT U1264 ( .A1(local_key[12]), .A2(n4297), .A3(\keys[0][12] ), .A4(
        n4293), .Y(n3545) );
  AO22X1_HVT U1265 ( .A1(local_key[13]), .A2(n4297), .A3(\keys[0][13] ), .A4(
        n4293), .Y(n3546) );
  AO22X1_HVT U1266 ( .A1(local_key[14]), .A2(n4297), .A3(\keys[0][14] ), .A4(
        n4293), .Y(n3547) );
  AO22X1_HVT U1267 ( .A1(local_key[15]), .A2(n4297), .A3(\keys[0][15] ), .A4(
        n4293), .Y(n3548) );
  AO22X1_HVT U1268 ( .A1(local_key[16]), .A2(n4297), .A3(\keys[0][16] ), .A4(
        n4293), .Y(n3549) );
  AO22X1_HVT U1269 ( .A1(local_key[17]), .A2(n4297), .A3(\keys[0][17] ), .A4(
        n4293), .Y(n3550) );
  AO22X1_HVT U1270 ( .A1(local_key[18]), .A2(n4297), .A3(\keys[0][18] ), .A4(
        n4293), .Y(n3551) );
  AO22X1_HVT U1271 ( .A1(local_key[19]), .A2(n4297), .A3(\keys[0][19] ), .A4(
        n4293), .Y(n3552) );
  AO22X1_HVT U1272 ( .A1(local_key[20]), .A2(n4297), .A3(\keys[0][20] ), .A4(
        n4293), .Y(n3553) );
  AO22X1_HVT U1273 ( .A1(local_key[21]), .A2(n4298), .A3(\keys[0][21] ), .A4(
        n4293), .Y(n3554) );
  AO22X1_HVT U1274 ( .A1(local_key[22]), .A2(n4298), .A3(\keys[0][22] ), .A4(
        n4293), .Y(n3555) );
  AO22X1_HVT U1275 ( .A1(local_key[23]), .A2(n4298), .A3(\keys[0][23] ), .A4(
        n4293), .Y(n3556) );
  AO22X1_HVT U1276 ( .A1(local_key[24]), .A2(n4298), .A3(\keys[0][24] ), .A4(
        n4293), .Y(n3557) );
  AO22X1_HVT U1277 ( .A1(local_key[25]), .A2(n4298), .A3(\keys[0][25] ), .A4(
        n4292), .Y(n3558) );
  AO22X1_HVT U1278 ( .A1(local_key[26]), .A2(n4298), .A3(\keys[0][26] ), .A4(
        n4292), .Y(n3559) );
  AO22X1_HVT U1279 ( .A1(local_key[27]), .A2(n4298), .A3(\keys[0][27] ), .A4(
        n4292), .Y(n3560) );
  AO22X1_HVT U1280 ( .A1(local_key[28]), .A2(n4298), .A3(\keys[0][28] ), .A4(
        n4292), .Y(n3561) );
  AO22X1_HVT U1281 ( .A1(local_key[29]), .A2(n4298), .A3(\keys[0][29] ), .A4(
        n4292), .Y(n3562) );
  AO22X1_HVT U1282 ( .A1(local_key[30]), .A2(n4298), .A3(\keys[0][30] ), .A4(
        n4292), .Y(n3563) );
  AO22X1_HVT U1283 ( .A1(local_key[31]), .A2(n4298), .A3(\keys[0][31] ), .A4(
        n4292), .Y(n3564) );
  AO22X1_HVT U1284 ( .A1(local_key[32]), .A2(n4298), .A3(\keys[0][32] ), .A4(
        n4292), .Y(n3565) );
  AO22X1_HVT U1285 ( .A1(local_key[33]), .A2(n4298), .A3(\keys[0][33] ), .A4(
        n4292), .Y(n3566) );
  AO22X1_HVT U1286 ( .A1(local_key[34]), .A2(n4298), .A3(\keys[0][34] ), .A4(
        n4292), .Y(n3567) );
  AO22X1_HVT U1287 ( .A1(local_key[35]), .A2(n4298), .A3(\keys[0][35] ), .A4(
        n4292), .Y(n3568) );
  AO22X1_HVT U1288 ( .A1(local_key[36]), .A2(n4299), .A3(\keys[0][36] ), .A4(
        n4292), .Y(n3569) );
  AO22X1_HVT U1289 ( .A1(local_key[37]), .A2(n4299), .A3(\keys[0][37] ), .A4(
        n4292), .Y(n3570) );
  AO22X1_HVT U1290 ( .A1(local_key[38]), .A2(n4299), .A3(\keys[0][38] ), .A4(
        n4291), .Y(n3571) );
  AO22X1_HVT U1291 ( .A1(local_key[39]), .A2(n4299), .A3(\keys[0][39] ), .A4(
        n4291), .Y(n3572) );
  AO22X1_HVT U1292 ( .A1(local_key[40]), .A2(n4299), .A3(\keys[0][40] ), .A4(
        n4291), .Y(n3573) );
  AO22X1_HVT U1293 ( .A1(local_key[41]), .A2(n4299), .A3(\keys[0][41] ), .A4(
        n4291), .Y(n3574) );
  AO22X1_HVT U1294 ( .A1(local_key[42]), .A2(n4299), .A3(\keys[0][42] ), .A4(
        n4291), .Y(n3575) );
  AO22X1_HVT U1295 ( .A1(local_key[43]), .A2(n4299), .A3(\keys[0][43] ), .A4(
        n4291), .Y(n3576) );
  AO22X1_HVT U1296 ( .A1(local_key[44]), .A2(n4299), .A3(\keys[0][44] ), .A4(
        n4291), .Y(n3577) );
  AO22X1_HVT U1297 ( .A1(local_key[45]), .A2(n4299), .A3(\keys[0][45] ), .A4(
        n4291), .Y(n3578) );
  AO22X1_HVT U1298 ( .A1(local_key[46]), .A2(n4299), .A3(\keys[0][46] ), .A4(
        n4291), .Y(n3579) );
  AO22X1_HVT U1299 ( .A1(local_key[47]), .A2(n4299), .A3(\keys[0][47] ), .A4(
        n4291), .Y(n3580) );
  AO22X1_HVT U1300 ( .A1(local_key[48]), .A2(n4299), .A3(\keys[0][48] ), .A4(
        n4291), .Y(n3581) );
  AO22X1_HVT U1301 ( .A1(local_key[49]), .A2(n4299), .A3(\keys[0][49] ), .A4(
        n4291), .Y(n3582) );
  AO22X1_HVT U1302 ( .A1(local_key[50]), .A2(n4299), .A3(\keys[0][50] ), .A4(
        n4291), .Y(n3583) );
  AO22X1_HVT U1303 ( .A1(local_key[51]), .A2(n4300), .A3(\keys[0][51] ), .A4(
        n4290), .Y(n3584) );
  AO22X1_HVT U1304 ( .A1(local_key[52]), .A2(n4300), .A3(\keys[0][52] ), .A4(
        n4290), .Y(n3585) );
  AO22X1_HVT U1305 ( .A1(local_key[53]), .A2(n4300), .A3(\keys[0][53] ), .A4(
        n4290), .Y(n3586) );
  AO22X1_HVT U1306 ( .A1(local_key[54]), .A2(n4300), .A3(\keys[0][54] ), .A4(
        n4290), .Y(n3587) );
  AO22X1_HVT U1307 ( .A1(local_key[55]), .A2(n4300), .A3(\keys[0][55] ), .A4(
        n4290), .Y(n3588) );
  AO22X1_HVT U1308 ( .A1(local_key[56]), .A2(n4300), .A3(\keys[0][56] ), .A4(
        n4290), .Y(n3589) );
  AO22X1_HVT U1309 ( .A1(local_key[57]), .A2(n4300), .A3(\keys[0][57] ), .A4(
        n4290), .Y(n3590) );
  AO22X1_HVT U1310 ( .A1(local_key[58]), .A2(n4300), .A3(\keys[0][58] ), .A4(
        n4290), .Y(n3591) );
  AO22X1_HVT U1311 ( .A1(local_key[59]), .A2(n4300), .A3(\keys[0][59] ), .A4(
        n4290), .Y(n3592) );
  AO22X1_HVT U1312 ( .A1(local_key[60]), .A2(n4300), .A3(\keys[0][60] ), .A4(
        n4290), .Y(n3593) );
  AO22X1_HVT U1313 ( .A1(local_key[61]), .A2(n4300), .A3(\keys[0][61] ), .A4(
        n4290), .Y(n3594) );
  AO22X1_HVT U1314 ( .A1(local_key[62]), .A2(n4300), .A3(\keys[0][62] ), .A4(
        n4290), .Y(n3595) );
  AO22X1_HVT U1315 ( .A1(local_key[63]), .A2(n4300), .A3(\keys[0][63] ), .A4(
        n4290), .Y(n3596) );
  AO22X1_HVT U1316 ( .A1(local_key[64]), .A2(n4300), .A3(\keys[0][64] ), .A4(
        n4289), .Y(n3597) );
  AO22X1_HVT U1317 ( .A1(local_key[65]), .A2(n4300), .A3(\keys[0][65] ), .A4(
        n4289), .Y(n3598) );
  AO22X1_HVT U1318 ( .A1(local_key[66]), .A2(n4301), .A3(\keys[0][66] ), .A4(
        n4289), .Y(n3599) );
  AO22X1_HVT U1319 ( .A1(local_key[67]), .A2(n4301), .A3(\keys[0][67] ), .A4(
        n4289), .Y(n3600) );
  AO22X1_HVT U1320 ( .A1(local_key[68]), .A2(n4301), .A3(\keys[0][68] ), .A4(
        n4289), .Y(n3601) );
  AO22X1_HVT U1321 ( .A1(local_key[69]), .A2(n4301), .A3(\keys[0][69] ), .A4(
        n4289), .Y(n3602) );
  AO22X1_HVT U1322 ( .A1(local_key[70]), .A2(n4301), .A3(\keys[0][70] ), .A4(
        n4289), .Y(n3603) );
  AO22X1_HVT U1323 ( .A1(local_key[71]), .A2(n4301), .A3(\keys[0][71] ), .A4(
        n4289), .Y(n3604) );
  AO22X1_HVT U1324 ( .A1(local_key[72]), .A2(n4301), .A3(\keys[0][72] ), .A4(
        n4289), .Y(n3605) );
  AO22X1_HVT U1325 ( .A1(local_key[73]), .A2(n4301), .A3(\keys[0][73] ), .A4(
        n4289), .Y(n3606) );
  AO22X1_HVT U1326 ( .A1(local_key[74]), .A2(n4301), .A3(\keys[0][74] ), .A4(
        n4289), .Y(n3607) );
  AO22X1_HVT U1327 ( .A1(local_key[75]), .A2(n4301), .A3(\keys[0][75] ), .A4(
        n4289), .Y(n3608) );
  AO22X1_HVT U1328 ( .A1(local_key[76]), .A2(n4301), .A3(\keys[0][76] ), .A4(
        n4289), .Y(n3609) );
  AO22X1_HVT U1329 ( .A1(local_key[77]), .A2(n4301), .A3(\keys[0][77] ), .A4(
        n4288), .Y(n3610) );
  AO22X1_HVT U1330 ( .A1(local_key[78]), .A2(n4301), .A3(\keys[0][78] ), .A4(
        n4288), .Y(n3611) );
  AO22X1_HVT U1331 ( .A1(local_key[79]), .A2(n4301), .A3(\keys[0][79] ), .A4(
        n4288), .Y(n3612) );
  AO22X1_HVT U1332 ( .A1(local_key[80]), .A2(n4301), .A3(\keys[0][80] ), .A4(
        n4288), .Y(n3613) );
  AO22X1_HVT U1333 ( .A1(local_key[81]), .A2(n4302), .A3(\keys[0][81] ), .A4(
        n4288), .Y(n3614) );
  AO22X1_HVT U1334 ( .A1(local_key[82]), .A2(n4302), .A3(\keys[0][82] ), .A4(
        n4288), .Y(n3615) );
  AO22X1_HVT U1335 ( .A1(local_key[83]), .A2(n4302), .A3(\keys[0][83] ), .A4(
        n4288), .Y(n3616) );
  AO22X1_HVT U1336 ( .A1(local_key[84]), .A2(n4302), .A3(\keys[0][84] ), .A4(
        n4288), .Y(n3617) );
  AO22X1_HVT U1337 ( .A1(local_key[85]), .A2(n4302), .A3(\keys[0][85] ), .A4(
        n4288), .Y(n3618) );
  AO22X1_HVT U1338 ( .A1(local_key[86]), .A2(n4302), .A3(\keys[0][86] ), .A4(
        n4288), .Y(n3619) );
  AO22X1_HVT U1339 ( .A1(local_key[87]), .A2(n4302), .A3(\keys[0][87] ), .A4(
        n4288), .Y(n3620) );
  AO22X1_HVT U1340 ( .A1(local_key[88]), .A2(n4302), .A3(\keys[0][88] ), .A4(
        n4288), .Y(n3621) );
  AO22X1_HVT U1341 ( .A1(local_key[89]), .A2(n4302), .A3(\keys[0][89] ), .A4(
        n4288), .Y(n3622) );
  AO22X1_HVT U1342 ( .A1(local_key[90]), .A2(n4302), .A3(\keys[0][90] ), .A4(
        n4287), .Y(n3623) );
  AO22X1_HVT U1343 ( .A1(local_key[91]), .A2(n4302), .A3(\keys[0][91] ), .A4(
        n4287), .Y(n3624) );
  AO22X1_HVT U1344 ( .A1(local_key[92]), .A2(n4302), .A3(\keys[0][92] ), .A4(
        n4287), .Y(n3625) );
  AO22X1_HVT U1345 ( .A1(local_key[93]), .A2(n4302), .A3(\keys[0][93] ), .A4(
        n4287), .Y(n3626) );
  AO22X1_HVT U1346 ( .A1(local_key[94]), .A2(n4302), .A3(\keys[0][94] ), .A4(
        n4287), .Y(n3627) );
  AO22X1_HVT U1347 ( .A1(local_key[95]), .A2(n4302), .A3(\keys[0][95] ), .A4(
        n4287), .Y(n3628) );
  AO22X1_HVT U1348 ( .A1(local_key[96]), .A2(n4303), .A3(\keys[0][96] ), .A4(
        n4287), .Y(n3629) );
  AO22X1_HVT U1349 ( .A1(local_key[97]), .A2(n4303), .A3(\keys[0][97] ), .A4(
        n4287), .Y(n3630) );
  AO22X1_HVT U1350 ( .A1(local_key[98]), .A2(n4303), .A3(\keys[0][98] ), .A4(
        n4287), .Y(n3631) );
  AO22X1_HVT U1351 ( .A1(local_key[99]), .A2(n4303), .A3(\keys[0][99] ), .A4(
        n4287), .Y(n3632) );
  AO22X1_HVT U1352 ( .A1(local_key[100]), .A2(n4303), .A3(\keys[0][100] ), 
        .A4(n4287), .Y(n3633) );
  AO22X1_HVT U1353 ( .A1(local_key[101]), .A2(n4303), .A3(\keys[0][101] ), 
        .A4(n4287), .Y(n3634) );
  AO22X1_HVT U1354 ( .A1(local_key[102]), .A2(n4303), .A3(\keys[0][102] ), 
        .A4(n4287), .Y(n3635) );
  AO22X1_HVT U1355 ( .A1(local_key[103]), .A2(n4303), .A3(\keys[0][103] ), 
        .A4(n4286), .Y(n3636) );
  AO22X1_HVT U1356 ( .A1(local_key[104]), .A2(n4303), .A3(\keys[0][104] ), 
        .A4(n4286), .Y(n3637) );
  AO22X1_HVT U1357 ( .A1(local_key[105]), .A2(n4303), .A3(\keys[0][105] ), 
        .A4(n4286), .Y(n3638) );
  AO22X1_HVT U1358 ( .A1(local_key[106]), .A2(n4303), .A3(\keys[0][106] ), 
        .A4(n4286), .Y(n3639) );
  AO22X1_HVT U1359 ( .A1(local_key[107]), .A2(n4303), .A3(\keys[0][107] ), 
        .A4(n4286), .Y(n3640) );
  AO22X1_HVT U1360 ( .A1(local_key[108]), .A2(n4303), .A3(\keys[0][108] ), 
        .A4(n4286), .Y(n3641) );
  AO22X1_HVT U1361 ( .A1(local_key[109]), .A2(n4303), .A3(\keys[0][109] ), 
        .A4(n4286), .Y(n3642) );
  AO22X1_HVT U1362 ( .A1(local_key[110]), .A2(n4303), .A3(\keys[0][110] ), 
        .A4(n4286), .Y(n3643) );
  AO22X1_HVT U1363 ( .A1(local_key[111]), .A2(n4304), .A3(\keys[0][111] ), 
        .A4(n4286), .Y(n3644) );
  AO22X1_HVT U1364 ( .A1(local_key[112]), .A2(n4304), .A3(\keys[0][112] ), 
        .A4(n4286), .Y(n3645) );
  AO22X1_HVT U1365 ( .A1(local_key[113]), .A2(n4304), .A3(\keys[0][113] ), 
        .A4(n4286), .Y(n3646) );
  AO22X1_HVT U1366 ( .A1(local_key[114]), .A2(n4304), .A3(\keys[0][114] ), 
        .A4(n4286), .Y(n3647) );
  AO22X1_HVT U1367 ( .A1(local_key[115]), .A2(n4304), .A3(\keys[0][115] ), 
        .A4(n4286), .Y(n3648) );
  AO22X1_HVT U1368 ( .A1(local_key[116]), .A2(n4304), .A3(\keys[0][116] ), 
        .A4(n4285), .Y(n3649) );
  AO22X1_HVT U1369 ( .A1(local_key[117]), .A2(n4304), .A3(\keys[0][117] ), 
        .A4(n4285), .Y(n3650) );
  AO22X1_HVT U1370 ( .A1(local_key[118]), .A2(n4304), .A3(\keys[0][118] ), 
        .A4(n4285), .Y(n3651) );
  AO22X1_HVT U1371 ( .A1(local_key[119]), .A2(n4304), .A3(\keys[0][119] ), 
        .A4(n4285), .Y(n3652) );
  AO22X1_HVT U1372 ( .A1(local_key[120]), .A2(n4304), .A3(\keys[0][120] ), 
        .A4(n4285), .Y(n3653) );
  AO22X1_HVT U1373 ( .A1(local_key[121]), .A2(n4304), .A3(\keys[0][121] ), 
        .A4(n4285), .Y(n3654) );
  AO22X1_HVT U1374 ( .A1(local_key[122]), .A2(n4304), .A3(\keys[0][122] ), 
        .A4(n4285), .Y(n3655) );
  AO22X1_HVT U1375 ( .A1(local_key[123]), .A2(n4304), .A3(\keys[0][123] ), 
        .A4(n4285), .Y(n3656) );
  AO22X1_HVT U1376 ( .A1(local_key[124]), .A2(n4304), .A3(\keys[0][124] ), 
        .A4(n4285), .Y(n3657) );
  AO22X1_HVT U1377 ( .A1(local_key[125]), .A2(n4304), .A3(\keys[0][125] ), 
        .A4(n4285), .Y(n3658) );
  AO22X1_HVT U1378 ( .A1(local_key[126]), .A2(n4305), .A3(\keys[0][126] ), 
        .A4(n4285), .Y(n3659) );
  AO22X1_HVT U1379 ( .A1(local_key[127]), .A2(n4305), .A3(\keys[0][127] ), 
        .A4(n4285), .Y(n3660) );
  AO222X1_HVT U1380 ( .A1(n4272), .A2(local_key[127]), .A3(n4259), .A4(n4101), 
        .A5(prev_key[127]), .A6(n4250), .Y(n3661) );
  AO222X1_HVT U1381 ( .A1(n4272), .A2(local_key[126]), .A3(n4259), .A4(n4098), 
        .A5(prev_key[126]), .A6(n4245), .Y(n3662) );
  AO222X1_HVT U1382 ( .A1(n4272), .A2(local_key[125]), .A3(n4259), .A4(
        keyout[125]), .A5(prev_key[125]), .A6(n4245), .Y(n3663) );
  AO222X1_HVT U1384 ( .A1(n4272), .A2(local_key[123]), .A3(n4259), .A4(
        keyout[123]), .A5(prev_key[123]), .A6(n4245), .Y(n3665) );
  AO222X1_HVT U1385 ( .A1(n4272), .A2(local_key[122]), .A3(n4259), .A4(
        keyout[122]), .A5(prev_key[122]), .A6(n4245), .Y(n3666) );
  AO222X1_HVT U1386 ( .A1(n4272), .A2(local_key[121]), .A3(n4259), .A4(
        keyout[121]), .A5(prev_key[121]), .A6(n4245), .Y(n3667) );
  AO222X1_HVT U1387 ( .A1(n4272), .A2(local_key[120]), .A3(n4259), .A4(n4095), 
        .A5(prev_key[120]), .A6(n4245), .Y(n3668) );
  AO222X1_HVT U1388 ( .A1(n4272), .A2(local_key[119]), .A3(n4259), .A4(
        keyout[119]), .A5(prev_key[119]), .A6(n4245), .Y(n3669) );
  AO222X1_HVT U1389 ( .A1(n4272), .A2(local_key[118]), .A3(n4259), .A4(
        keyout[118]), .A5(prev_key[118]), .A6(n4245), .Y(n3670) );
  AO222X1_HVT U1390 ( .A1(n4272), .A2(local_key[117]), .A3(n4259), .A4(
        keyout[117]), .A5(prev_key[117]), .A6(n4245), .Y(n3671) );
  AO222X1_HVT U1391 ( .A1(n4272), .A2(local_key[116]), .A3(n4259), .A4(
        keyout[116]), .A5(prev_key[116]), .A6(n4245), .Y(n3672) );
  AO222X1_HVT U1392 ( .A1(n4273), .A2(local_key[115]), .A3(n4260), .A4(
        keyout[115]), .A5(prev_key[115]), .A6(n4245), .Y(n3673) );
  AO222X1_HVT U1393 ( .A1(n4273), .A2(local_key[114]), .A3(n4260), .A4(
        keyout[114]), .A5(prev_key[114]), .A6(n4246), .Y(n3674) );
  AO222X1_HVT U1394 ( .A1(n4273), .A2(local_key[113]), .A3(n4260), .A4(
        keyout[113]), .A5(prev_key[113]), .A6(n4246), .Y(n3675) );
  AO222X1_HVT U1395 ( .A1(n4273), .A2(local_key[112]), .A3(n4260), .A4(
        keyout[112]), .A5(prev_key[112]), .A6(n4246), .Y(n3676) );
  AO222X1_HVT U1396 ( .A1(n4273), .A2(local_key[111]), .A3(n4260), .A4(
        keyout[111]), .A5(prev_key[111]), .A6(n4246), .Y(n3677) );
  AO222X1_HVT U1397 ( .A1(n4273), .A2(local_key[110]), .A3(n4260), .A4(
        keyout[110]), .A5(prev_key[110]), .A6(n4246), .Y(n3678) );
  AO222X1_HVT U1398 ( .A1(n4273), .A2(local_key[109]), .A3(n4260), .A4(
        keyout[109]), .A5(prev_key[109]), .A6(n4246), .Y(n3679) );
  AO222X1_HVT U1399 ( .A1(n4273), .A2(local_key[108]), .A3(n4260), .A4(
        keyout[108]), .A5(prev_key[108]), .A6(n4246), .Y(n3680) );
  AO222X1_HVT U1400 ( .A1(n4273), .A2(local_key[107]), .A3(n4260), .A4(
        keyout[107]), .A5(prev_key[107]), .A6(n4246), .Y(n3681) );
  AO222X1_HVT U1401 ( .A1(n4273), .A2(local_key[106]), .A3(n4260), .A4(
        keyout[106]), .A5(prev_key[106]), .A6(n4246), .Y(n3682) );
  AO222X1_HVT U1402 ( .A1(n4273), .A2(local_key[105]), .A3(n4260), .A4(
        keyout[105]), .A5(prev_key[105]), .A6(n4246), .Y(n3683) );
  AO222X1_HVT U1403 ( .A1(n4273), .A2(local_key[104]), .A3(n4260), .A4(
        keyout[104]), .A5(prev_key[104]), .A6(n4246), .Y(n3684) );
  AO222X1_HVT U1404 ( .A1(n4274), .A2(local_key[103]), .A3(n4261), .A4(
        keyout[103]), .A5(prev_key[103]), .A6(n4246), .Y(n3685) );
  AO222X1_HVT U1405 ( .A1(n4274), .A2(local_key[102]), .A3(n4261), .A4(
        keyout[102]), .A5(prev_key[102]), .A6(n4247), .Y(n3686) );
  AO222X1_HVT U1406 ( .A1(n4274), .A2(local_key[101]), .A3(n4261), .A4(
        keyout[101]), .A5(prev_key[101]), .A6(n4247), .Y(n3687) );
  AO222X1_HVT U1407 ( .A1(n4274), .A2(local_key[100]), .A3(n4261), .A4(
        keyout[100]), .A5(prev_key[100]), .A6(n4247), .Y(n3688) );
  AO222X1_HVT U1408 ( .A1(n4274), .A2(local_key[99]), .A3(n4261), .A4(
        keyout[99]), .A5(prev_key[99]), .A6(n4247), .Y(n3689) );
  AO222X1_HVT U1409 ( .A1(n4274), .A2(local_key[98]), .A3(n4261), .A4(
        keyout[98]), .A5(prev_key[98]), .A6(n4247), .Y(n3690) );
  AO222X1_HVT U1410 ( .A1(n4274), .A2(local_key[97]), .A3(n4261), .A4(
        keyout[97]), .A5(prev_key[97]), .A6(n4247), .Y(n3691) );
  AO222X1_HVT U1411 ( .A1(n4274), .A2(local_key[96]), .A3(n4261), .A4(
        keyout[96]), .A5(prev_key[96]), .A6(n4247), .Y(n3692) );
  AO222X1_HVT U1412 ( .A1(n4274), .A2(local_key[95]), .A3(n4261), .A4(
        keyout[95]), .A5(prev_key[95]), .A6(n4247), .Y(n3693) );
  AO222X1_HVT U1413 ( .A1(n4274), .A2(local_key[94]), .A3(n4261), .A4(
        keyout[94]), .A5(prev_key[94]), .A6(n4247), .Y(n3694) );
  AO222X1_HVT U1414 ( .A1(n4274), .A2(local_key[93]), .A3(n4261), .A4(
        keyout[93]), .A5(prev_key[93]), .A6(n4247), .Y(n3695) );
  AO222X1_HVT U1415 ( .A1(n4274), .A2(local_key[92]), .A3(n4261), .A4(
        keyout[92]), .A5(prev_key[92]), .A6(n4247), .Y(n3696) );
  AO222X1_HVT U1416 ( .A1(n4275), .A2(local_key[91]), .A3(n4262), .A4(
        keyout[91]), .A5(prev_key[91]), .A6(n4247), .Y(n3697) );
  AO222X1_HVT U1417 ( .A1(n4275), .A2(local_key[90]), .A3(n4262), .A4(
        keyout[90]), .A5(prev_key[90]), .A6(n4248), .Y(n3698) );
  AO222X1_HVT U1418 ( .A1(n4275), .A2(local_key[89]), .A3(n4262), .A4(
        keyout[89]), .A5(prev_key[89]), .A6(n4248), .Y(n3699) );
  AO222X1_HVT U1419 ( .A1(n4275), .A2(local_key[88]), .A3(n4262), .A4(n4092), 
        .A5(prev_key[88]), .A6(n4248), .Y(n3700) );
  AO222X1_HVT U1421 ( .A1(n4275), .A2(local_key[86]), .A3(n4262), .A4(
        keyout[86]), .A5(prev_key[86]), .A6(n4248), .Y(n3702) );
  AO222X1_HVT U1422 ( .A1(n4275), .A2(local_key[85]), .A3(n4262), .A4(n1), 
        .A5(prev_key[85]), .A6(n4248), .Y(n3703) );
  AO222X1_HVT U1423 ( .A1(n4275), .A2(local_key[84]), .A3(n4262), .A4(
        keyout[84]), .A5(prev_key[84]), .A6(n4248), .Y(n3704) );
  AO222X1_HVT U1425 ( .A1(n4275), .A2(local_key[82]), .A3(n4262), .A4(
        keyout[82]), .A5(prev_key[82]), .A6(n4248), .Y(n3706) );
  AO222X1_HVT U1426 ( .A1(n4275), .A2(local_key[81]), .A3(n4262), .A4(
        keyout[81]), .A5(prev_key[81]), .A6(n4248), .Y(n3707) );
  AO222X1_HVT U1428 ( .A1(n4276), .A2(local_key[79]), .A3(keyout[79]), .A4(
        n4263), .A5(prev_key[79]), .A6(n4248), .Y(n3709) );
  AO222X1_HVT U1429 ( .A1(n4276), .A2(local_key[78]), .A3(n4263), .A4(
        keyout[78]), .A5(prev_key[78]), .A6(n4249), .Y(n3710) );
  AO222X1_HVT U1433 ( .A1(n4276), .A2(local_key[74]), .A3(n4263), .A4(
        keyout[74]), .A5(prev_key[74]), .A6(n4249), .Y(n3714) );
  AO222X1_HVT U1434 ( .A1(n4276), .A2(local_key[73]), .A3(n4263), .A4(
        keyout[73]), .A5(prev_key[73]), .A6(n4249), .Y(n3715) );
  AO222X1_HVT U1435 ( .A1(n4276), .A2(local_key[72]), .A3(n4263), .A4(
        keyout[72]), .A5(prev_key[72]), .A6(n4249), .Y(n3716) );
  AO222X1_HVT U1436 ( .A1(n4276), .A2(local_key[71]), .A3(n4263), .A4(
        keyout[71]), .A5(prev_key[71]), .A6(n4249), .Y(n3717) );
  AO222X1_HVT U1437 ( .A1(n4276), .A2(local_key[70]), .A3(n4263), .A4(
        keyout[70]), .A5(prev_key[70]), .A6(n4249), .Y(n3718) );
  AO222X1_HVT U1438 ( .A1(n4276), .A2(local_key[69]), .A3(n4263), .A4(
        keyout[69]), .A5(prev_key[69]), .A6(n4249), .Y(n3719) );
  AO222X1_HVT U1439 ( .A1(n4276), .A2(local_key[68]), .A3(n4263), .A4(
        keyout[68]), .A5(prev_key[68]), .A6(n4249), .Y(n3720) );
  AO222X1_HVT U1440 ( .A1(n4277), .A2(local_key[67]), .A3(n4264), .A4(
        keyout[67]), .A5(prev_key[67]), .A6(n4249), .Y(n3721) );
  AO222X1_HVT U1441 ( .A1(n4277), .A2(local_key[66]), .A3(n4264), .A4(
        keyout[66]), .A5(prev_key[66]), .A6(n4250), .Y(n3722) );
  AO222X1_HVT U1442 ( .A1(n4277), .A2(local_key[65]), .A3(n4264), .A4(n3870), 
        .A5(prev_key[65]), .A6(n4250), .Y(n3723) );
  AO222X1_HVT U1443 ( .A1(n4277), .A2(local_key[64]), .A3(n4264), .A4(
        keyout[64]), .A5(prev_key[64]), .A6(n4250), .Y(n3724) );
  AO222X1_HVT U1445 ( .A1(n4277), .A2(local_key[62]), .A3(n4264), .A4(
        keyout[62]), .A5(prev_key[62]), .A6(n4250), .Y(n3726) );
  AO222X1_HVT U1447 ( .A1(n4277), .A2(local_key[60]), .A3(n4264), .A4(
        keyout[60]), .A5(prev_key[60]), .A6(n4250), .Y(n3728) );
  AO222X1_HVT U1448 ( .A1(n4277), .A2(local_key[59]), .A3(n4264), .A4(n4088), 
        .A5(prev_key[59]), .A6(n4250), .Y(n3729) );
  AO222X1_HVT U1449 ( .A1(n4277), .A2(local_key[58]), .A3(n4264), .A4(n4086), 
        .A5(prev_key[58]), .A6(n4250), .Y(n3730) );
  AO222X1_HVT U1450 ( .A1(n4277), .A2(local_key[57]), .A3(n4264), .A4(n4084), 
        .A5(prev_key[57]), .A6(n4250), .Y(n3731) );
  AO222X1_HVT U1451 ( .A1(n4277), .A2(local_key[56]), .A3(n4264), .A4(
        keyout[56]), .A5(prev_key[56]), .A6(n4250), .Y(n3732) );
  AO222X1_HVT U1452 ( .A1(n4278), .A2(local_key[55]), .A3(keyout[55]), .A4(
        n4265), .A5(prev_key[55]), .A6(n4251), .Y(n3733) );
  AO222X1_HVT U1453 ( .A1(n4278), .A2(local_key[54]), .A3(n4265), .A4(
        keyout[54]), .A5(prev_key[54]), .A6(n4251), .Y(n3734) );
  AO222X1_HVT U1454 ( .A1(n4278), .A2(local_key[53]), .A3(n4265), .A4(n3874), 
        .A5(prev_key[53]), .A6(n4251), .Y(n3735) );
  AO222X1_HVT U1455 ( .A1(n4278), .A2(local_key[52]), .A3(n4265), .A4(
        keyout[52]), .A5(prev_key[52]), .A6(n4251), .Y(n3736) );
  AO222X1_HVT U1456 ( .A1(n4278), .A2(local_key[51]), .A3(n4265), .A4(
        keyout[51]), .A5(prev_key[51]), .A6(n4251), .Y(n3737) );
  AO222X1_HVT U1457 ( .A1(n4278), .A2(local_key[50]), .A3(n4265), .A4(
        keyout[50]), .A5(prev_key[50]), .A6(n4251), .Y(n3738) );
  AO222X1_HVT U1458 ( .A1(n4278), .A2(local_key[49]), .A3(n4265), .A4(
        keyout[49]), .A5(prev_key[49]), .A6(n4251), .Y(n3739) );
  AO222X1_HVT U1459 ( .A1(n4278), .A2(local_key[48]), .A3(n4265), .A4(
        keyout[48]), .A5(prev_key[48]), .A6(n4251), .Y(n3740) );
  AO222X1_HVT U1460 ( .A1(n4278), .A2(local_key[47]), .A3(n4265), .A4(
        keyout[47]), .A5(prev_key[47]), .A6(n4251), .Y(n3741) );
  AO222X1_HVT U1461 ( .A1(n4278), .A2(local_key[46]), .A3(n4265), .A4(n3944), 
        .A5(prev_key[46]), .A6(n4251), .Y(n3742) );
  AO222X1_HVT U1462 ( .A1(n4278), .A2(local_key[45]), .A3(n4265), .A4(
        keyout[45]), .A5(prev_key[45]), .A6(n4251), .Y(n3743) );
  AO222X1_HVT U1463 ( .A1(n4278), .A2(local_key[44]), .A3(n4265), .A4(
        keyout[44]), .A5(prev_key[44]), .A6(n4251), .Y(n3744) );
  AO222X1_HVT U1464 ( .A1(n4279), .A2(local_key[43]), .A3(n4266), .A4(
        keyout[43]), .A5(prev_key[43]), .A6(n4252), .Y(n3745) );
  AO222X1_HVT U1466 ( .A1(n4279), .A2(local_key[41]), .A3(n4266), .A4(
        keyout[41]), .A5(prev_key[41]), .A6(n4252), .Y(n3747) );
  AO222X1_HVT U1467 ( .A1(n4279), .A2(local_key[40]), .A3(n4266), .A4(
        keyout[40]), .A5(prev_key[40]), .A6(n4252), .Y(n3748) );
  AO222X1_HVT U1468 ( .A1(n4279), .A2(local_key[39]), .A3(n4266), .A4(
        keyout[39]), .A5(prev_key[39]), .A6(n4252), .Y(n3749) );
  AO222X1_HVT U1469 ( .A1(n4279), .A2(local_key[38]), .A3(n4266), .A4(
        keyout[38]), .A5(prev_key[38]), .A6(n4252), .Y(n3750) );
  AO222X1_HVT U1471 ( .A1(n4279), .A2(local_key[36]), .A3(n4266), .A4(
        keyout[36]), .A5(prev_key[36]), .A6(n4252), .Y(n3752) );
  AO222X1_HVT U1472 ( .A1(n4279), .A2(local_key[35]), .A3(n4266), .A4(
        keyout[35]), .A5(prev_key[35]), .A6(n4252), .Y(n3753) );
  AO222X1_HVT U1473 ( .A1(n4279), .A2(local_key[34]), .A3(n4266), .A4(
        keyout[34]), .A5(prev_key[34]), .A6(n4252), .Y(n3754) );
  AO222X1_HVT U1474 ( .A1(n4279), .A2(local_key[33]), .A3(n4266), .A4(
        keyout[33]), .A5(prev_key[33]), .A6(n4252), .Y(n3755) );
  AO222X1_HVT U1475 ( .A1(n4279), .A2(local_key[32]), .A3(n4266), .A4(
        keyout[32]), .A5(prev_key[32]), .A6(n4252), .Y(n3756) );
  AO222X1_HVT U1476 ( .A1(n4280), .A2(local_key[31]), .A3(n4267), .A4(
        keyout[31]), .A5(prev_key[31]), .A6(n4253), .Y(n3757) );
  AO222X1_HVT U1477 ( .A1(n4280), .A2(local_key[30]), .A3(n4267), .A4(n4082), 
        .A5(prev_key[30]), .A6(n4253), .Y(n3758) );
  AO222X1_HVT U1478 ( .A1(n4280), .A2(local_key[29]), .A3(n4267), .A4(n4079), 
        .A5(prev_key[29]), .A6(n4253), .Y(n3759) );
  AO222X1_HVT U1479 ( .A1(n4280), .A2(local_key[28]), .A3(n4267), .A4(n4076), 
        .A5(prev_key[28]), .A6(n4253), .Y(n3760) );
  AO222X1_HVT U1480 ( .A1(n4280), .A2(local_key[27]), .A3(n4267), .A4(n4073), 
        .A5(prev_key[27]), .A6(n4253), .Y(n3761) );
  AO222X1_HVT U1481 ( .A1(n4280), .A2(local_key[26]), .A3(n4267), .A4(n4070), 
        .A5(prev_key[26]), .A6(n4253), .Y(n3762) );
  AO222X1_HVT U1482 ( .A1(n4280), .A2(local_key[25]), .A3(n4267), .A4(
        keyout[25]), .A5(prev_key[25]), .A6(n4253), .Y(n3763) );
  AO222X1_HVT U1483 ( .A1(n4280), .A2(local_key[24]), .A3(n4267), .A4(n4065), 
        .A5(prev_key[24]), .A6(n4253), .Y(n3764) );
  AO222X1_HVT U1484 ( .A1(n4280), .A2(local_key[23]), .A3(n4267), .A4(n4062), 
        .A5(n3954), .A6(n4253), .Y(n3765) );
  AO222X1_HVT U1485 ( .A1(n4280), .A2(local_key[22]), .A3(n4267), .A4(n4059), 
        .A5(prev_key[22]), .A6(n4253), .Y(n3766) );
  AO222X1_HVT U1486 ( .A1(n4280), .A2(local_key[21]), .A3(n4267), .A4(n4056), 
        .A5(prev_key[21]), .A6(n4253), .Y(n3767) );
  AO222X1_HVT U1487 ( .A1(n4280), .A2(local_key[20]), .A3(n4267), .A4(n4053), 
        .A5(prev_key[20]), .A6(n4253), .Y(n3768) );
  AO222X1_HVT U1488 ( .A1(n4281), .A2(local_key[19]), .A3(n4268), .A4(n4050), 
        .A5(prev_key[19]), .A6(n4254), .Y(n3769) );
  AO222X1_HVT U1489 ( .A1(n4281), .A2(local_key[18]), .A3(n4268), .A4(n4047), 
        .A5(prev_key[18]), .A6(n4254), .Y(n3770) );
  AO222X1_HVT U1490 ( .A1(n4281), .A2(local_key[17]), .A3(n4268), .A4(n4044), 
        .A5(prev_key[17]), .A6(n4254), .Y(n3771) );
  AO222X1_HVT U1491 ( .A1(n4281), .A2(local_key[16]), .A3(n4268), .A4(n4041), 
        .A5(prev_key[16]), .A6(n4254), .Y(n3772) );
  AO222X1_HVT U1492 ( .A1(n4281), .A2(local_key[15]), .A3(n4268), .A4(n4038), 
        .A5(n3975), .A6(n4254), .Y(n3773) );
  AO222X1_HVT U1493 ( .A1(n4281), .A2(local_key[14]), .A3(n4268), .A4(n4035), 
        .A5(prev_key[14]), .A6(n4254), .Y(n3774) );
  AO222X1_HVT U1494 ( .A1(n4281), .A2(local_key[13]), .A3(n4268), .A4(n4032), 
        .A5(prev_key[13]), .A6(n4254), .Y(n3775) );
  AO222X1_HVT U1495 ( .A1(n4281), .A2(local_key[12]), .A3(n4268), .A4(n4029), 
        .A5(prev_key[12]), .A6(n4254), .Y(n3776) );
  AO222X1_HVT U1496 ( .A1(n4281), .A2(local_key[11]), .A3(n4268), .A4(n4026), 
        .A5(prev_key[11]), .A6(n4254), .Y(n3777) );
  AO222X1_HVT U1497 ( .A1(n4281), .A2(local_key[10]), .A3(n4268), .A4(n4023), 
        .A5(prev_key[10]), .A6(n4254), .Y(n3778) );
  AO222X1_HVT U1498 ( .A1(n4281), .A2(local_key[9]), .A3(n4268), .A4(n4020), 
        .A5(prev_key[9]), .A6(n4254), .Y(n3779) );
  AO222X1_HVT U1499 ( .A1(n4281), .A2(local_key[8]), .A3(n4268), .A4(n4017), 
        .A5(prev_key[8]), .A6(n4254), .Y(n3780) );
  AO222X1_HVT U1500 ( .A1(n1441), .A2(local_key[7]), .A3(n4269), .A4(keyout[7]), .A5(prev_key[7]), .A6(n4255), .Y(n3781) );
  AO222X1_HVT U1501 ( .A1(n1441), .A2(local_key[6]), .A3(n4269), .A4(n4013), 
        .A5(prev_key[6]), .A6(n4255), .Y(n3782) );
  AO222X1_HVT U1502 ( .A1(n1441), .A2(local_key[5]), .A3(n4269), .A4(n4010), 
        .A5(prev_key[5]), .A6(n4255), .Y(n3783) );
  AO222X1_HVT U1503 ( .A1(n1441), .A2(local_key[4]), .A3(n4269), .A4(n4007), 
        .A5(prev_key[4]), .A6(n4255), .Y(n3784) );
  AO222X1_HVT U1504 ( .A1(n1441), .A2(local_key[3]), .A3(n4269), .A4(n4004), 
        .A5(prev_key[3]), .A6(n4255), .Y(n3785) );
  AO222X1_HVT U1505 ( .A1(n1441), .A2(local_key[2]), .A3(n4269), .A4(keyout[2]), .A5(prev_key[2]), .A6(n4255), .Y(n3786) );
  AO222X1_HVT U1506 ( .A1(n1441), .A2(local_key[1]), .A3(n4269), .A4(n4000), 
        .A5(prev_key[1]), .A6(n4255), .Y(n3787) );
  AO222X1_HVT U1507 ( .A1(n1441), .A2(local_key[0]), .A3(n4269), .A4(n3997), 
        .A5(prev_key[0]), .A6(n4255), .Y(n3788) );
  AND2X1_HVT U1508 ( .A1(n4256), .A2(n1444), .Y(n1442) );
  AO22X1_HVT U1509 ( .A1(round_number[3]), .A2(n4255), .A3(n4257), .A4(n1445), 
        .Y(n3789) );
  NAND2X0_HVT U1510 ( .A1(n1446), .A2(n1447), .Y(n1445) );
  AO22X1_HVT U1511 ( .A1(round_number[2]), .A2(n4255), .A3(n4257), .A4(n1448), 
        .Y(n3790) );
  NAND3X0_HVT U1512 ( .A1(n1449), .A2(n1450), .A3(n1451), .Y(n1448) );
  AO22X1_HVT U1513 ( .A1(round_number[1]), .A2(n4255), .A3(n4258), .A4(n1452), 
        .Y(n3791) );
  AO221X1_HVT U1514 ( .A1(n4258), .A2(n1453), .A3(round_number[0]), .A4(n4255), 
        .A5(n1441), .Y(n3792) );
  AND2X1_HVT U1515 ( .A1(n4257), .A2(n1454), .Y(n1441) );
  NAND3X0_HVT U1516 ( .A1(n1455), .A2(n1456), .A3(n1451), .Y(n1453) );
  AND2X1_HVT U1517 ( .A1(n1457), .A2(n1458), .Y(n1451) );
  NAND2X0_HVT U1518 ( .A1(n1459), .A2(n4559), .Y(n1443) );
  AO21X1_HVT U1519 ( .A1(done), .A2(n4559), .A3(n4546), .Y(n3793) );
  NAND4X0_HVT U1520 ( .A1(n4353), .A2(n4331), .A3(n4375), .A4(n1460), .Y(n3794) );
  OA21X1_HVT U1521 ( .A1(n16), .A2(n1461), .A3(n4407), .Y(n1460) );
  NAND4X0_HVT U1523 ( .A1(n4375), .A2(n4285), .A3(n4464), .A4(n1462), .Y(n3795) );
  OA21X1_HVT U1524 ( .A1(n17), .A2(n1461), .A3(n1463), .Y(n1462) );
  NAND4X0_HVT U1527 ( .A1(n4442), .A2(n4420), .A3(n4464), .A4(n1464), .Y(n3796) );
  OA21X1_HVT U1528 ( .A1(n11), .A2(n1461), .A3(n4496), .Y(n1464) );
  NAND4X0_HVT U1531 ( .A1(n1463), .A2(n1465), .A3(n4442), .A4(n4353), .Y(n3797) );
  OR2X1_HVT U1534 ( .A1(n1461), .A2(n18), .Y(n1465) );
  OR2X1_HVT U1535 ( .A1(n1459), .A2(rest), .Y(n1461) );
  OR2X1_HVT U1536 ( .A1(n1444), .A2(n1454), .Y(n1459) );
  AND4X1_HVT U1537 ( .A1(n18), .A2(n17), .A3(n16), .A4(n11), .Y(n1454) );
  NAND4X0_HVT U1538 ( .A1(n4555), .A2(n1446), .A3(n1449), .A4(n1457), .Y(n1444) );
  NAND2X0_HVT U1539 ( .A1(n1467), .A2(state[0]), .Y(n1457) );
  NAND2X0_HVT U1540 ( .A1(n1467), .A2(n18), .Y(n1449) );
  AND3X1_HVT U1541 ( .A1(n17), .A2(n11), .A3(state[2]), .Y(n1467) );
  AND2X1_HVT U1542 ( .A1(n1466), .A2(n1456), .Y(n1446) );
  NAND3X0_HVT U1543 ( .A1(n1468), .A2(n17), .A3(state[0]), .Y(n1456) );
  NAND3X0_HVT U1544 ( .A1(n18), .A2(n17), .A3(n1468), .Y(n1466) );
  OR3X1_HVT U1545 ( .A1(n4556), .A2(n1469), .A3(n1470), .Y(n1452) );
  NAND3X0_HVT U1546 ( .A1(n1458), .A2(n1447), .A3(n1450), .Y(n1470) );
  NAND3X0_HVT U1547 ( .A1(n1471), .A2(state[0]), .A3(state[2]), .Y(n1458) );
  NAND3X0_HVT U1548 ( .A1(state[0]), .A2(n16), .A3(n1471), .Y(n1455) );
  AND3X1_HVT U1549 ( .A1(n4407), .A2(n4318), .A3(n4496), .Y(n1463) );
  NAND3X0_HVT U1551 ( .A1(n1468), .A2(n18), .A3(state[1]), .Y(n1447) );
  AND3X1_HVT U1553 ( .A1(n18), .A2(n16), .A3(n1471), .Y(n1469) );
  NAND3X0_HVT U1555 ( .A1(n1471), .A2(n18), .A3(state[2]), .Y(n1450) );
  AND2X1_HVT U1556 ( .A1(state[1]), .A2(n11), .Y(n1471) );
  AO22X1_HVT U1557 ( .A1(key_round[0]), .A2(n4525), .A3(n4546), .A4(n1472), 
        .Y(n2125) );
  NAND4X0_HVT U1558 ( .A1(n1473), .A2(n1474), .A3(n1475), .A4(n1476), .Y(n1472) );
  OA222X1_HVT U1559 ( .A1(n1170), .A2(n4232), .A3(n4220), .A4(n1426), .A5(
        n1298), .A6(n4207), .Y(n1476) );
  OA222X1_HVT U1560 ( .A1(n786), .A2(n4194), .A3(n1042), .A4(n4181), .A5(n914), 
        .A6(n4168), .Y(n1475) );
  OA222X1_HVT U1561 ( .A1(n402), .A2(n4155), .A3(n658), .A4(n4142), .A5(n530), 
        .A6(n4129), .Y(n1474) );
  OA22X1_HVT U1562 ( .A1(n274), .A2(n4116), .A3(n146), .A4(n4103), .Y(n1473)
         );
  AO22X1_HVT U1563 ( .A1(key_round[1]), .A2(n4525), .A3(n4554), .A4(n1488), 
        .Y(n2126) );
  NAND4X0_HVT U1564 ( .A1(n1489), .A2(n1490), .A3(n1491), .A4(n1492), .Y(n1488) );
  OA222X1_HVT U1565 ( .A1(n1169), .A2(n4232), .A3(n4220), .A4(n1425), .A5(
        n1297), .A6(n4207), .Y(n1492) );
  OA222X1_HVT U1566 ( .A1(n785), .A2(n4194), .A3(n1041), .A4(n4181), .A5(n913), 
        .A6(n4168), .Y(n1491) );
  OA222X1_HVT U1567 ( .A1(n401), .A2(n4155), .A3(n657), .A4(n4142), .A5(n529), 
        .A6(n4129), .Y(n1490) );
  OA22X1_HVT U1568 ( .A1(n273), .A2(n4116), .A3(n145), .A4(n4103), .Y(n1489)
         );
  AO22X1_HVT U1569 ( .A1(key_round[2]), .A2(n4525), .A3(n4554), .A4(n1493), 
        .Y(n2127) );
  NAND4X0_HVT U1570 ( .A1(n1494), .A2(n1495), .A3(n1496), .A4(n1497), .Y(n1493) );
  OA222X1_HVT U1571 ( .A1(n1168), .A2(n4232), .A3(n4220), .A4(n1424), .A5(
        n1296), .A6(n4207), .Y(n1497) );
  OA222X1_HVT U1572 ( .A1(n784), .A2(n4194), .A3(n1040), .A4(n4181), .A5(n912), 
        .A6(n4168), .Y(n1496) );
  OA222X1_HVT U1573 ( .A1(n400), .A2(n4155), .A3(n656), .A4(n4142), .A5(n528), 
        .A6(n4129), .Y(n1495) );
  OA22X1_HVT U1574 ( .A1(n272), .A2(n4116), .A3(n144), .A4(n4103), .Y(n1494)
         );
  AO22X1_HVT U1575 ( .A1(key_round[3]), .A2(n4525), .A3(n4554), .A4(n1498), 
        .Y(n2128) );
  NAND4X0_HVT U1576 ( .A1(n1499), .A2(n1500), .A3(n1501), .A4(n1502), .Y(n1498) );
  OA222X1_HVT U1577 ( .A1(n1167), .A2(n4232), .A3(n4220), .A4(n1423), .A5(
        n1295), .A6(n4207), .Y(n1502) );
  OA222X1_HVT U1578 ( .A1(n783), .A2(n4194), .A3(n1039), .A4(n4181), .A5(n911), 
        .A6(n4168), .Y(n1501) );
  OA222X1_HVT U1579 ( .A1(n399), .A2(n4155), .A3(n655), .A4(n4142), .A5(n527), 
        .A6(n4129), .Y(n1500) );
  OA22X1_HVT U1580 ( .A1(n271), .A2(n4116), .A3(n143), .A4(n4103), .Y(n1499)
         );
  AO22X1_HVT U1581 ( .A1(key_round[4]), .A2(n4525), .A3(n4554), .A4(n1503), 
        .Y(n2129) );
  NAND4X0_HVT U1582 ( .A1(n1504), .A2(n1505), .A3(n1506), .A4(n1507), .Y(n1503) );
  OA222X1_HVT U1583 ( .A1(n1166), .A2(n4232), .A3(n4220), .A4(n1422), .A5(
        n1294), .A6(n4207), .Y(n1507) );
  OA222X1_HVT U1584 ( .A1(n782), .A2(n4194), .A3(n1038), .A4(n4181), .A5(n910), 
        .A6(n4168), .Y(n1506) );
  OA222X1_HVT U1585 ( .A1(n398), .A2(n4155), .A3(n654), .A4(n4142), .A5(n526), 
        .A6(n4129), .Y(n1505) );
  OA22X1_HVT U1586 ( .A1(n270), .A2(n4116), .A3(n142), .A4(n4103), .Y(n1504)
         );
  AO22X1_HVT U1587 ( .A1(key_round[5]), .A2(n4525), .A3(n4554), .A4(n1508), 
        .Y(n2130) );
  NAND4X0_HVT U1588 ( .A1(n1509), .A2(n1510), .A3(n1511), .A4(n1512), .Y(n1508) );
  OA222X1_HVT U1589 ( .A1(n1165), .A2(n4232), .A3(n4220), .A4(n1421), .A5(
        n1293), .A6(n4207), .Y(n1512) );
  OA222X1_HVT U1590 ( .A1(n781), .A2(n4194), .A3(n1037), .A4(n4181), .A5(n909), 
        .A6(n4168), .Y(n1511) );
  OA222X1_HVT U1591 ( .A1(n397), .A2(n4155), .A3(n653), .A4(n4142), .A5(n525), 
        .A6(n4129), .Y(n1510) );
  OA22X1_HVT U1592 ( .A1(n269), .A2(n4116), .A3(n141), .A4(n4103), .Y(n1509)
         );
  AO22X1_HVT U1593 ( .A1(key_round[6]), .A2(n4526), .A3(n4554), .A4(n1513), 
        .Y(n2131) );
  NAND4X0_HVT U1594 ( .A1(n1514), .A2(n1515), .A3(n1516), .A4(n1517), .Y(n1513) );
  OA222X1_HVT U1595 ( .A1(n1164), .A2(n4232), .A3(n4220), .A4(n1420), .A5(
        n1292), .A6(n4207), .Y(n1517) );
  OA222X1_HVT U1596 ( .A1(n780), .A2(n4194), .A3(n1036), .A4(n4181), .A5(n908), 
        .A6(n4168), .Y(n1516) );
  OA222X1_HVT U1597 ( .A1(n396), .A2(n4155), .A3(n652), .A4(n4142), .A5(n524), 
        .A6(n4129), .Y(n1515) );
  OA22X1_HVT U1598 ( .A1(n268), .A2(n4116), .A3(n140), .A4(n4103), .Y(n1514)
         );
  AO22X1_HVT U1599 ( .A1(key_round[7]), .A2(n4526), .A3(n4554), .A4(n1518), 
        .Y(n2132) );
  NAND4X0_HVT U1600 ( .A1(n1519), .A2(n1520), .A3(n1521), .A4(n1522), .Y(n1518) );
  OA222X1_HVT U1601 ( .A1(n1163), .A2(n4232), .A3(n4220), .A4(n1419), .A5(
        n1291), .A6(n4207), .Y(n1522) );
  OA222X1_HVT U1602 ( .A1(n779), .A2(n4194), .A3(n1035), .A4(n4181), .A5(n907), 
        .A6(n4168), .Y(n1521) );
  OA222X1_HVT U1603 ( .A1(n395), .A2(n4155), .A3(n651), .A4(n4142), .A5(n523), 
        .A6(n4129), .Y(n1520) );
  OA22X1_HVT U1604 ( .A1(n267), .A2(n4116), .A3(n139), .A4(n4103), .Y(n1519)
         );
  AO22X1_HVT U1605 ( .A1(key_round[8]), .A2(n4526), .A3(n4554), .A4(n1523), 
        .Y(n2133) );
  NAND4X0_HVT U1606 ( .A1(n1524), .A2(n1525), .A3(n1526), .A4(n1527), .Y(n1523) );
  OA222X1_HVT U1607 ( .A1(n1162), .A2(n4232), .A3(n4220), .A4(n1418), .A5(
        n1290), .A6(n4207), .Y(n1527) );
  OA222X1_HVT U1608 ( .A1(n778), .A2(n4194), .A3(n1034), .A4(n4181), .A5(n906), 
        .A6(n4168), .Y(n1526) );
  OA222X1_HVT U1609 ( .A1(n394), .A2(n4155), .A3(n650), .A4(n4142), .A5(n522), 
        .A6(n4129), .Y(n1525) );
  OA22X1_HVT U1610 ( .A1(n266), .A2(n4116), .A3(n138), .A4(n4103), .Y(n1524)
         );
  AO22X1_HVT U1611 ( .A1(key_round[9]), .A2(n4526), .A3(n4554), .A4(n1528), 
        .Y(n2134) );
  NAND4X0_HVT U1612 ( .A1(n1529), .A2(n1530), .A3(n1531), .A4(n1532), .Y(n1528) );
  OA222X1_HVT U1613 ( .A1(n1161), .A2(n4232), .A3(n4220), .A4(n1417), .A5(
        n1289), .A6(n4207), .Y(n1532) );
  OA222X1_HVT U1614 ( .A1(n777), .A2(n4194), .A3(n1033), .A4(n4181), .A5(n905), 
        .A6(n4168), .Y(n1531) );
  OA222X1_HVT U1615 ( .A1(n393), .A2(n4155), .A3(n649), .A4(n4142), .A5(n521), 
        .A6(n4129), .Y(n1530) );
  OA22X1_HVT U1616 ( .A1(n265), .A2(n4116), .A3(n137), .A4(n4103), .Y(n1529)
         );
  AO22X1_HVT U1617 ( .A1(key_round[10]), .A2(n4526), .A3(n4553), .A4(n1533), 
        .Y(n2135) );
  NAND4X0_HVT U1618 ( .A1(n1534), .A2(n1535), .A3(n1536), .A4(n1537), .Y(n1533) );
  OA222X1_HVT U1619 ( .A1(n1160), .A2(n4232), .A3(n4220), .A4(n1416), .A5(
        n1288), .A6(n4207), .Y(n1537) );
  OA222X1_HVT U1620 ( .A1(n776), .A2(n4194), .A3(n1032), .A4(n4181), .A5(n904), 
        .A6(n4168), .Y(n1536) );
  OA222X1_HVT U1621 ( .A1(n392), .A2(n4155), .A3(n648), .A4(n4142), .A5(n520), 
        .A6(n4129), .Y(n1535) );
  OA22X1_HVT U1622 ( .A1(n264), .A2(n4116), .A3(n136), .A4(n4103), .Y(n1534)
         );
  AO22X1_HVT U1623 ( .A1(key_round[11]), .A2(n4526), .A3(n4553), .A4(n1538), 
        .Y(n2136) );
  NAND4X0_HVT U1624 ( .A1(n1539), .A2(n1540), .A3(n1541), .A4(n1542), .Y(n1538) );
  OA222X1_HVT U1625 ( .A1(n1159), .A2(n4232), .A3(n4220), .A4(n1415), .A5(
        n1287), .A6(n4207), .Y(n1542) );
  OA222X1_HVT U1626 ( .A1(n775), .A2(n4194), .A3(n1031), .A4(n4181), .A5(n903), 
        .A6(n4168), .Y(n1541) );
  OA222X1_HVT U1627 ( .A1(n391), .A2(n4155), .A3(n647), .A4(n4142), .A5(n519), 
        .A6(n4129), .Y(n1540) );
  OA22X1_HVT U1628 ( .A1(n263), .A2(n4116), .A3(n135), .A4(n4103), .Y(n1539)
         );
  AO22X1_HVT U1629 ( .A1(key_round[12]), .A2(n4526), .A3(n4553), .A4(n1543), 
        .Y(n2137) );
  NAND4X0_HVT U1630 ( .A1(n1544), .A2(n1545), .A3(n1546), .A4(n1547), .Y(n1543) );
  OA222X1_HVT U1631 ( .A1(n1158), .A2(n4233), .A3(n4221), .A4(n1414), .A5(
        n1286), .A6(n4208), .Y(n1547) );
  OA222X1_HVT U1632 ( .A1(n774), .A2(n4195), .A3(n1030), .A4(n4182), .A5(n902), 
        .A6(n4169), .Y(n1546) );
  OA222X1_HVT U1633 ( .A1(n390), .A2(n4156), .A3(n646), .A4(n4143), .A5(n518), 
        .A6(n4130), .Y(n1545) );
  OA22X1_HVT U1634 ( .A1(n262), .A2(n4117), .A3(n134), .A4(n4104), .Y(n1544)
         );
  AO22X1_HVT U1635 ( .A1(key_round[13]), .A2(n4526), .A3(n4553), .A4(n1548), 
        .Y(n2138) );
  NAND4X0_HVT U1636 ( .A1(n1549), .A2(n1550), .A3(n1551), .A4(n1552), .Y(n1548) );
  OA222X1_HVT U1637 ( .A1(n1157), .A2(n4233), .A3(n4221), .A4(n1413), .A5(
        n1285), .A6(n4208), .Y(n1552) );
  OA222X1_HVT U1638 ( .A1(n773), .A2(n4195), .A3(n1029), .A4(n4182), .A5(n901), 
        .A6(n4169), .Y(n1551) );
  OA222X1_HVT U1639 ( .A1(n389), .A2(n4156), .A3(n645), .A4(n4143), .A5(n517), 
        .A6(n4130), .Y(n1550) );
  OA22X1_HVT U1640 ( .A1(n261), .A2(n4117), .A3(n133), .A4(n4104), .Y(n1549)
         );
  AO22X1_HVT U1641 ( .A1(key_round[14]), .A2(n4526), .A3(n4553), .A4(n1553), 
        .Y(n2139) );
  NAND4X0_HVT U1642 ( .A1(n1554), .A2(n1555), .A3(n1556), .A4(n1557), .Y(n1553) );
  OA222X1_HVT U1643 ( .A1(n1156), .A2(n4233), .A3(n4221), .A4(n1412), .A5(
        n1284), .A6(n4208), .Y(n1557) );
  OA222X1_HVT U1644 ( .A1(n772), .A2(n4195), .A3(n1028), .A4(n4182), .A5(n900), 
        .A6(n4169), .Y(n1556) );
  OA222X1_HVT U1645 ( .A1(n388), .A2(n4156), .A3(n644), .A4(n4143), .A5(n516), 
        .A6(n4130), .Y(n1555) );
  OA22X1_HVT U1646 ( .A1(n260), .A2(n4117), .A3(n132), .A4(n4104), .Y(n1554)
         );
  AO22X1_HVT U1647 ( .A1(key_round[15]), .A2(n4526), .A3(n4553), .A4(n1558), 
        .Y(n2140) );
  NAND4X0_HVT U1648 ( .A1(n1559), .A2(n1560), .A3(n1561), .A4(n1562), .Y(n1558) );
  OA222X1_HVT U1649 ( .A1(n1155), .A2(n4233), .A3(n4221), .A4(n1411), .A5(
        n1283), .A6(n4208), .Y(n1562) );
  OA222X1_HVT U1650 ( .A1(n771), .A2(n4195), .A3(n1027), .A4(n4182), .A5(n899), 
        .A6(n4169), .Y(n1561) );
  OA222X1_HVT U1651 ( .A1(n387), .A2(n4156), .A3(n643), .A4(n4143), .A5(n515), 
        .A6(n4130), .Y(n1560) );
  OA22X1_HVT U1652 ( .A1(n259), .A2(n4117), .A3(n131), .A4(n4104), .Y(n1559)
         );
  AO22X1_HVT U1653 ( .A1(key_round[16]), .A2(n4526), .A3(n4553), .A4(n1563), 
        .Y(n2141) );
  NAND4X0_HVT U1654 ( .A1(n1564), .A2(n1565), .A3(n1566), .A4(n1567), .Y(n1563) );
  OA222X1_HVT U1655 ( .A1(n1154), .A2(n4233), .A3(n4221), .A4(n1410), .A5(
        n1282), .A6(n4208), .Y(n1567) );
  OA222X1_HVT U1656 ( .A1(n770), .A2(n4195), .A3(n1026), .A4(n4182), .A5(n898), 
        .A6(n4169), .Y(n1566) );
  OA222X1_HVT U1657 ( .A1(n386), .A2(n4156), .A3(n642), .A4(n4143), .A5(n514), 
        .A6(n4130), .Y(n1565) );
  OA22X1_HVT U1658 ( .A1(n258), .A2(n4117), .A3(n130), .A4(n4104), .Y(n1564)
         );
  AO22X1_HVT U1659 ( .A1(key_round[17]), .A2(n4527), .A3(n4553), .A4(n1568), 
        .Y(n2142) );
  NAND4X0_HVT U1660 ( .A1(n1569), .A2(n1570), .A3(n1571), .A4(n1572), .Y(n1568) );
  OA222X1_HVT U1661 ( .A1(n1153), .A2(n4233), .A3(n4221), .A4(n1409), .A5(
        n1281), .A6(n4208), .Y(n1572) );
  OA222X1_HVT U1662 ( .A1(n769), .A2(n4195), .A3(n1025), .A4(n4182), .A5(n897), 
        .A6(n4169), .Y(n1571) );
  OA222X1_HVT U1663 ( .A1(n385), .A2(n4156), .A3(n641), .A4(n4143), .A5(n513), 
        .A6(n4130), .Y(n1570) );
  OA22X1_HVT U1664 ( .A1(n257), .A2(n4117), .A3(n129), .A4(n4104), .Y(n1569)
         );
  AO22X1_HVT U1665 ( .A1(key_round[18]), .A2(n4527), .A3(n4553), .A4(n1573), 
        .Y(n2143) );
  NAND4X0_HVT U1666 ( .A1(n1574), .A2(n1575), .A3(n1576), .A4(n1577), .Y(n1573) );
  OA222X1_HVT U1667 ( .A1(n1152), .A2(n4233), .A3(n4221), .A4(n1408), .A5(
        n1280), .A6(n4208), .Y(n1577) );
  OA222X1_HVT U1668 ( .A1(n768), .A2(n4195), .A3(n1024), .A4(n4182), .A5(n896), 
        .A6(n4169), .Y(n1576) );
  OA222X1_HVT U1669 ( .A1(n384), .A2(n4156), .A3(n640), .A4(n4143), .A5(n512), 
        .A6(n4130), .Y(n1575) );
  OA22X1_HVT U1670 ( .A1(n256), .A2(n4117), .A3(n128), .A4(n4104), .Y(n1574)
         );
  AO22X1_HVT U1671 ( .A1(key_round[19]), .A2(n4527), .A3(n4553), .A4(n1578), 
        .Y(n2144) );
  NAND4X0_HVT U1672 ( .A1(n1579), .A2(n1580), .A3(n1581), .A4(n1582), .Y(n1578) );
  OA222X1_HVT U1673 ( .A1(n1151), .A2(n4233), .A3(n4221), .A4(n1407), .A5(
        n1279), .A6(n4208), .Y(n1582) );
  OA222X1_HVT U1674 ( .A1(n767), .A2(n4195), .A3(n1023), .A4(n4182), .A5(n895), 
        .A6(n4169), .Y(n1581) );
  OA222X1_HVT U1675 ( .A1(n383), .A2(n4156), .A3(n639), .A4(n4143), .A5(n511), 
        .A6(n4130), .Y(n1580) );
  OA22X1_HVT U1676 ( .A1(n255), .A2(n4117), .A3(n127), .A4(n4104), .Y(n1579)
         );
  AO22X1_HVT U1677 ( .A1(key_round[20]), .A2(n4527), .A3(n4553), .A4(n1583), 
        .Y(n2145) );
  NAND4X0_HVT U1678 ( .A1(n1584), .A2(n1585), .A3(n1586), .A4(n1587), .Y(n1583) );
  OA222X1_HVT U1679 ( .A1(n1150), .A2(n4233), .A3(n4221), .A4(n1406), .A5(
        n1278), .A6(n4208), .Y(n1587) );
  OA222X1_HVT U1680 ( .A1(n766), .A2(n4195), .A3(n1022), .A4(n4182), .A5(n894), 
        .A6(n4169), .Y(n1586) );
  OA222X1_HVT U1681 ( .A1(n382), .A2(n4156), .A3(n638), .A4(n4143), .A5(n510), 
        .A6(n4130), .Y(n1585) );
  OA22X1_HVT U1682 ( .A1(n254), .A2(n4117), .A3(n126), .A4(n4104), .Y(n1584)
         );
  AO22X1_HVT U1683 ( .A1(key_round[21]), .A2(n4527), .A3(n4553), .A4(n1588), 
        .Y(n2146) );
  NAND4X0_HVT U1684 ( .A1(n1589), .A2(n1590), .A3(n1591), .A4(n1592), .Y(n1588) );
  OA222X1_HVT U1685 ( .A1(n1149), .A2(n4233), .A3(n4221), .A4(n1405), .A5(
        n1277), .A6(n4208), .Y(n1592) );
  OA222X1_HVT U1686 ( .A1(n765), .A2(n4195), .A3(n1021), .A4(n4182), .A5(n893), 
        .A6(n4169), .Y(n1591) );
  OA222X1_HVT U1687 ( .A1(n381), .A2(n4156), .A3(n637), .A4(n4143), .A5(n509), 
        .A6(n4130), .Y(n1590) );
  OA22X1_HVT U1688 ( .A1(n253), .A2(n4117), .A3(n125), .A4(n4104), .Y(n1589)
         );
  AO22X1_HVT U1689 ( .A1(key_round[22]), .A2(n4527), .A3(n4553), .A4(n1593), 
        .Y(n2147) );
  NAND4X0_HVT U1690 ( .A1(n1594), .A2(n1595), .A3(n1596), .A4(n1597), .Y(n1593) );
  OA222X1_HVT U1691 ( .A1(n1148), .A2(n4233), .A3(n4221), .A4(n1404), .A5(
        n1276), .A6(n4208), .Y(n1597) );
  OA222X1_HVT U1692 ( .A1(n764), .A2(n4195), .A3(n1020), .A4(n4182), .A5(n892), 
        .A6(n4169), .Y(n1596) );
  OA222X1_HVT U1693 ( .A1(n380), .A2(n4156), .A3(n636), .A4(n4143), .A5(n508), 
        .A6(n4130), .Y(n1595) );
  OA22X1_HVT U1694 ( .A1(n252), .A2(n4117), .A3(n124), .A4(n4104), .Y(n1594)
         );
  AO22X1_HVT U1695 ( .A1(key_round[23]), .A2(n4527), .A3(n4553), .A4(n1598), 
        .Y(n2148) );
  NAND4X0_HVT U1696 ( .A1(n1599), .A2(n1600), .A3(n1601), .A4(n1602), .Y(n1598) );
  OA222X1_HVT U1697 ( .A1(n1147), .A2(n4233), .A3(n4221), .A4(n1403), .A5(
        n1275), .A6(n4208), .Y(n1602) );
  OA222X1_HVT U1698 ( .A1(n763), .A2(n4195), .A3(n1019), .A4(n4182), .A5(n891), 
        .A6(n4169), .Y(n1601) );
  OA222X1_HVT U1699 ( .A1(n379), .A2(n4156), .A3(n635), .A4(n4143), .A5(n507), 
        .A6(n4130), .Y(n1600) );
  OA22X1_HVT U1700 ( .A1(n251), .A2(n4117), .A3(n123), .A4(n4104), .Y(n1599)
         );
  AO22X1_HVT U1701 ( .A1(key_round[24]), .A2(n4527), .A3(n4553), .A4(n1603), 
        .Y(n2149) );
  NAND4X0_HVT U1702 ( .A1(n1604), .A2(n1605), .A3(n1606), .A4(n1607), .Y(n1603) );
  OA222X1_HVT U1703 ( .A1(n1146), .A2(n4234), .A3(n4221), .A4(n1402), .A5(
        n1274), .A6(n4209), .Y(n1607) );
  OA222X1_HVT U1704 ( .A1(n762), .A2(n4196), .A3(n1018), .A4(n4183), .A5(n890), 
        .A6(n4170), .Y(n1606) );
  OA222X1_HVT U1705 ( .A1(n378), .A2(n4157), .A3(n634), .A4(n4144), .A5(n506), 
        .A6(n4131), .Y(n1605) );
  OA22X1_HVT U1706 ( .A1(n250), .A2(n4118), .A3(n122), .A4(n4105), .Y(n1604)
         );
  AO22X1_HVT U1707 ( .A1(key_round[25]), .A2(n4527), .A3(n4552), .A4(n1608), 
        .Y(n2150) );
  NAND4X0_HVT U1708 ( .A1(n1609), .A2(n1610), .A3(n1611), .A4(n1612), .Y(n1608) );
  OA222X1_HVT U1709 ( .A1(n1145), .A2(n4234), .A3(n4220), .A4(n1401), .A5(
        n1273), .A6(n4209), .Y(n1612) );
  OA222X1_HVT U1710 ( .A1(n761), .A2(n4196), .A3(n1017), .A4(n4183), .A5(n889), 
        .A6(n4170), .Y(n1611) );
  OA222X1_HVT U1711 ( .A1(n377), .A2(n4157), .A3(n633), .A4(n4144), .A5(n505), 
        .A6(n4131), .Y(n1610) );
  OA22X1_HVT U1712 ( .A1(n249), .A2(n4118), .A3(n121), .A4(n4105), .Y(n1609)
         );
  AO22X1_HVT U1713 ( .A1(key_round[26]), .A2(n4527), .A3(n4552), .A4(n1613), 
        .Y(n2151) );
  NAND4X0_HVT U1714 ( .A1(n1614), .A2(n1615), .A3(n1616), .A4(n1617), .Y(n1613) );
  OA222X1_HVT U1715 ( .A1(n1144), .A2(n4234), .A3(n4229), .A4(n1400), .A5(
        n1272), .A6(n4209), .Y(n1617) );
  OA222X1_HVT U1716 ( .A1(n760), .A2(n4196), .A3(n1016), .A4(n4183), .A5(n888), 
        .A6(n4170), .Y(n1616) );
  OA222X1_HVT U1717 ( .A1(n376), .A2(n4157), .A3(n632), .A4(n4144), .A5(n504), 
        .A6(n4131), .Y(n1615) );
  OA22X1_HVT U1718 ( .A1(n248), .A2(n4118), .A3(n120), .A4(n4105), .Y(n1614)
         );
  AO22X1_HVT U1719 ( .A1(key_round[27]), .A2(n4527), .A3(n4552), .A4(n1618), 
        .Y(n2152) );
  NAND4X0_HVT U1720 ( .A1(n1619), .A2(n1620), .A3(n1621), .A4(n1622), .Y(n1618) );
  OA222X1_HVT U1721 ( .A1(n1143), .A2(n4234), .A3(n4229), .A4(n1399), .A5(
        n1271), .A6(n4209), .Y(n1622) );
  OA222X1_HVT U1722 ( .A1(n759), .A2(n4196), .A3(n1015), .A4(n4183), .A5(n887), 
        .A6(n4170), .Y(n1621) );
  OA222X1_HVT U1723 ( .A1(n375), .A2(n4157), .A3(n631), .A4(n4144), .A5(n503), 
        .A6(n4131), .Y(n1620) );
  OA22X1_HVT U1724 ( .A1(n247), .A2(n4118), .A3(n119), .A4(n4105), .Y(n1619)
         );
  AO22X1_HVT U1725 ( .A1(key_round[28]), .A2(n4527), .A3(n4552), .A4(n1623), 
        .Y(n2153) );
  NAND4X0_HVT U1726 ( .A1(n1624), .A2(n1625), .A3(n1626), .A4(n1627), .Y(n1623) );
  OA222X1_HVT U1727 ( .A1(n1142), .A2(n4234), .A3(n4229), .A4(n1398), .A5(
        n1270), .A6(n4209), .Y(n1627) );
  OA222X1_HVT U1728 ( .A1(n758), .A2(n4196), .A3(n1014), .A4(n4183), .A5(n886), 
        .A6(n4170), .Y(n1626) );
  OA222X1_HVT U1729 ( .A1(n374), .A2(n4157), .A3(n630), .A4(n4144), .A5(n502), 
        .A6(n4131), .Y(n1625) );
  OA22X1_HVT U1730 ( .A1(n246), .A2(n4118), .A3(n118), .A4(n4105), .Y(n1624)
         );
  AO22X1_HVT U1731 ( .A1(key_round[29]), .A2(n4528), .A3(n4552), .A4(n1628), 
        .Y(n2154) );
  NAND4X0_HVT U1732 ( .A1(n1629), .A2(n1630), .A3(n1631), .A4(n1632), .Y(n1628) );
  OA222X1_HVT U1733 ( .A1(n1141), .A2(n4234), .A3(n4229), .A4(n1397), .A5(
        n1269), .A6(n4209), .Y(n1632) );
  OA222X1_HVT U1734 ( .A1(n757), .A2(n4196), .A3(n1013), .A4(n4183), .A5(n885), 
        .A6(n4170), .Y(n1631) );
  OA222X1_HVT U1735 ( .A1(n373), .A2(n4157), .A3(n629), .A4(n4144), .A5(n501), 
        .A6(n4131), .Y(n1630) );
  OA22X1_HVT U1736 ( .A1(n245), .A2(n4118), .A3(n117), .A4(n4105), .Y(n1629)
         );
  AO22X1_HVT U1737 ( .A1(key_round[30]), .A2(n4528), .A3(n4552), .A4(n1633), 
        .Y(n2155) );
  NAND4X0_HVT U1738 ( .A1(n1634), .A2(n1635), .A3(n1636), .A4(n1637), .Y(n1633) );
  OA222X1_HVT U1739 ( .A1(n1140), .A2(n4234), .A3(n4229), .A4(n1396), .A5(
        n1268), .A6(n4209), .Y(n1637) );
  OA222X1_HVT U1740 ( .A1(n756), .A2(n4196), .A3(n1012), .A4(n4183), .A5(n884), 
        .A6(n4170), .Y(n1636) );
  OA222X1_HVT U1741 ( .A1(n372), .A2(n4157), .A3(n628), .A4(n4144), .A5(n500), 
        .A6(n4131), .Y(n1635) );
  OA22X1_HVT U1742 ( .A1(n244), .A2(n4118), .A3(n116), .A4(n4105), .Y(n1634)
         );
  AO22X1_HVT U1743 ( .A1(key_round[31]), .A2(n4528), .A3(n4548), .A4(n1638), 
        .Y(n2156) );
  NAND4X0_HVT U1744 ( .A1(n1639), .A2(n1640), .A3(n1641), .A4(n1642), .Y(n1638) );
  OA222X1_HVT U1745 ( .A1(n1139), .A2(n4234), .A3(n4229), .A4(n1395), .A5(
        n1267), .A6(n4209), .Y(n1642) );
  OA222X1_HVT U1746 ( .A1(n755), .A2(n4196), .A3(n1011), .A4(n4183), .A5(n883), 
        .A6(n4170), .Y(n1641) );
  OA222X1_HVT U1747 ( .A1(n371), .A2(n4157), .A3(n627), .A4(n4144), .A5(n499), 
        .A6(n4131), .Y(n1640) );
  OA22X1_HVT U1748 ( .A1(n243), .A2(n4118), .A3(n115), .A4(n4105), .Y(n1639)
         );
  AO22X1_HVT U1749 ( .A1(key_round[32]), .A2(n4528), .A3(n4552), .A4(n1643), 
        .Y(n2157) );
  NAND4X0_HVT U1750 ( .A1(n1644), .A2(n1645), .A3(n1646), .A4(n1647), .Y(n1643) );
  OA222X1_HVT U1751 ( .A1(n1138), .A2(n4234), .A3(n4229), .A4(n1394), .A5(
        n1266), .A6(n4209), .Y(n1647) );
  OA222X1_HVT U1752 ( .A1(n754), .A2(n4196), .A3(n1010), .A4(n4183), .A5(n882), 
        .A6(n4170), .Y(n1646) );
  OA222X1_HVT U1753 ( .A1(n370), .A2(n4157), .A3(n626), .A4(n4144), .A5(n498), 
        .A6(n4131), .Y(n1645) );
  OA22X1_HVT U1754 ( .A1(n242), .A2(n4118), .A3(n114), .A4(n4105), .Y(n1644)
         );
  AO22X1_HVT U1755 ( .A1(key_round[33]), .A2(n4528), .A3(n4552), .A4(n1648), 
        .Y(n2158) );
  NAND4X0_HVT U1756 ( .A1(n1649), .A2(n1650), .A3(n1651), .A4(n1652), .Y(n1648) );
  OA222X1_HVT U1757 ( .A1(n1137), .A2(n4234), .A3(n4229), .A4(n1393), .A5(
        n1265), .A6(n4209), .Y(n1652) );
  OA222X1_HVT U1758 ( .A1(n753), .A2(n4196), .A3(n1009), .A4(n4183), .A5(n881), 
        .A6(n4170), .Y(n1651) );
  OA222X1_HVT U1759 ( .A1(n369), .A2(n4157), .A3(n625), .A4(n4144), .A5(n497), 
        .A6(n4131), .Y(n1650) );
  OA22X1_HVT U1760 ( .A1(n241), .A2(n4118), .A3(n113), .A4(n4105), .Y(n1649)
         );
  AO22X1_HVT U1761 ( .A1(key_round[34]), .A2(n4528), .A3(n4552), .A4(n1653), 
        .Y(n2159) );
  NAND4X0_HVT U1762 ( .A1(n1654), .A2(n1655), .A3(n1656), .A4(n1657), .Y(n1653) );
  OA222X1_HVT U1763 ( .A1(n1136), .A2(n4234), .A3(n4229), .A4(n1392), .A5(
        n1264), .A6(n4209), .Y(n1657) );
  OA222X1_HVT U1764 ( .A1(n752), .A2(n4196), .A3(n1008), .A4(n4183), .A5(n880), 
        .A6(n4170), .Y(n1656) );
  OA222X1_HVT U1765 ( .A1(n368), .A2(n4157), .A3(n624), .A4(n4144), .A5(n496), 
        .A6(n4131), .Y(n1655) );
  OA22X1_HVT U1766 ( .A1(n240), .A2(n4118), .A3(n112), .A4(n4105), .Y(n1654)
         );
  AO22X1_HVT U1767 ( .A1(key_round[35]), .A2(n4528), .A3(n4552), .A4(n1658), 
        .Y(n2160) );
  NAND4X0_HVT U1768 ( .A1(n1659), .A2(n1660), .A3(n1661), .A4(n1662), .Y(n1658) );
  OA222X1_HVT U1769 ( .A1(n1135), .A2(n4234), .A3(n4229), .A4(n1391), .A5(
        n1263), .A6(n4209), .Y(n1662) );
  OA222X1_HVT U1770 ( .A1(n751), .A2(n4196), .A3(n1007), .A4(n4183), .A5(n879), 
        .A6(n4170), .Y(n1661) );
  OA222X1_HVT U1771 ( .A1(n367), .A2(n4157), .A3(n623), .A4(n4144), .A5(n495), 
        .A6(n4131), .Y(n1660) );
  OA22X1_HVT U1772 ( .A1(n239), .A2(n4118), .A3(n111), .A4(n4105), .Y(n1659)
         );
  AO22X1_HVT U1773 ( .A1(key_round[36]), .A2(n4528), .A3(n4552), .A4(n1663), 
        .Y(n2161) );
  NAND4X0_HVT U1774 ( .A1(n1664), .A2(n1665), .A3(n1666), .A4(n1667), .Y(n1663) );
  OA222X1_HVT U1775 ( .A1(n1134), .A2(n4235), .A3(n4222), .A4(n1390), .A5(
        n1262), .A6(n4210), .Y(n1667) );
  OA222X1_HVT U1776 ( .A1(n750), .A2(n4197), .A3(n1006), .A4(n4184), .A5(n878), 
        .A6(n4171), .Y(n1666) );
  OA222X1_HVT U1777 ( .A1(n366), .A2(n4158), .A3(n622), .A4(n4145), .A5(n494), 
        .A6(n4132), .Y(n1665) );
  OA22X1_HVT U1778 ( .A1(n238), .A2(n4119), .A3(n110), .A4(n4106), .Y(n1664)
         );
  AO22X1_HVT U1779 ( .A1(key_round[37]), .A2(n4528), .A3(n4552), .A4(n1668), 
        .Y(n2162) );
  NAND4X0_HVT U1780 ( .A1(n1669), .A2(n1670), .A3(n1671), .A4(n1672), .Y(n1668) );
  OA222X1_HVT U1781 ( .A1(n1133), .A2(n4235), .A3(n4222), .A4(n1389), .A5(
        n1261), .A6(n4210), .Y(n1672) );
  OA222X1_HVT U1782 ( .A1(n749), .A2(n4197), .A3(n1005), .A4(n4184), .A5(n877), 
        .A6(n4171), .Y(n1671) );
  OA222X1_HVT U1783 ( .A1(n365), .A2(n4158), .A3(n621), .A4(n4145), .A5(n493), 
        .A6(n4132), .Y(n1670) );
  OA22X1_HVT U1784 ( .A1(n237), .A2(n4119), .A3(n109), .A4(n4106), .Y(n1669)
         );
  AO22X1_HVT U1785 ( .A1(key_round[38]), .A2(n4528), .A3(n4552), .A4(n1673), 
        .Y(n2163) );
  NAND4X0_HVT U1786 ( .A1(n1674), .A2(n1675), .A3(n1676), .A4(n1677), .Y(n1673) );
  OA222X1_HVT U1787 ( .A1(n1132), .A2(n4235), .A3(n4222), .A4(n1388), .A5(
        n1260), .A6(n4210), .Y(n1677) );
  OA222X1_HVT U1788 ( .A1(n748), .A2(n4197), .A3(n1004), .A4(n4184), .A5(n876), 
        .A6(n4171), .Y(n1676) );
  OA222X1_HVT U1789 ( .A1(n364), .A2(n4158), .A3(n620), .A4(n4145), .A5(n492), 
        .A6(n4132), .Y(n1675) );
  OA22X1_HVT U1790 ( .A1(n236), .A2(n4119), .A3(n108), .A4(n4106), .Y(n1674)
         );
  AO22X1_HVT U1791 ( .A1(key_round[39]), .A2(n4528), .A3(n4552), .A4(n1678), 
        .Y(n2164) );
  NAND4X0_HVT U1792 ( .A1(n1679), .A2(n1680), .A3(n1681), .A4(n1682), .Y(n1678) );
  OA222X1_HVT U1793 ( .A1(n1131), .A2(n4235), .A3(n4222), .A4(n1387), .A5(
        n1259), .A6(n4210), .Y(n1682) );
  OA222X1_HVT U1794 ( .A1(n747), .A2(n4197), .A3(n1003), .A4(n4184), .A5(n875), 
        .A6(n4171), .Y(n1681) );
  OA222X1_HVT U1795 ( .A1(n363), .A2(n4158), .A3(n619), .A4(n4145), .A5(n491), 
        .A6(n4132), .Y(n1680) );
  OA22X1_HVT U1796 ( .A1(n235), .A2(n4119), .A3(n107), .A4(n4106), .Y(n1679)
         );
  AO22X1_HVT U1797 ( .A1(key_round[40]), .A2(n4528), .A3(n4552), .A4(n1683), 
        .Y(n2165) );
  NAND4X0_HVT U1798 ( .A1(n1684), .A2(n1685), .A3(n1686), .A4(n1687), .Y(n1683) );
  OA222X1_HVT U1799 ( .A1(n1130), .A2(n4235), .A3(n4222), .A4(n1386), .A5(
        n1258), .A6(n4210), .Y(n1687) );
  OA222X1_HVT U1800 ( .A1(n746), .A2(n4197), .A3(n1002), .A4(n4184), .A5(n874), 
        .A6(n4171), .Y(n1686) );
  OA222X1_HVT U1801 ( .A1(n362), .A2(n4158), .A3(n618), .A4(n4145), .A5(n490), 
        .A6(n4132), .Y(n1685) );
  OA22X1_HVT U1802 ( .A1(n234), .A2(n4119), .A3(n106), .A4(n4106), .Y(n1684)
         );
  AO22X1_HVT U1803 ( .A1(key_round[41]), .A2(n4529), .A3(n4551), .A4(n1688), 
        .Y(n2166) );
  NAND4X0_HVT U1804 ( .A1(n1689), .A2(n1690), .A3(n1691), .A4(n1692), .Y(n1688) );
  OA222X1_HVT U1805 ( .A1(n1129), .A2(n4235), .A3(n4222), .A4(n1385), .A5(
        n1257), .A6(n4210), .Y(n1692) );
  OA222X1_HVT U1806 ( .A1(n745), .A2(n4197), .A3(n1001), .A4(n4184), .A5(n873), 
        .A6(n4171), .Y(n1691) );
  OA222X1_HVT U1807 ( .A1(n361), .A2(n4158), .A3(n617), .A4(n4145), .A5(n489), 
        .A6(n4132), .Y(n1690) );
  OA22X1_HVT U1808 ( .A1(n233), .A2(n4119), .A3(n105), .A4(n4106), .Y(n1689)
         );
  AO22X1_HVT U1809 ( .A1(key_round[42]), .A2(n4529), .A3(n4551), .A4(n1693), 
        .Y(n2167) );
  NAND4X0_HVT U1810 ( .A1(n1694), .A2(n1695), .A3(n1696), .A4(n1697), .Y(n1693) );
  OA222X1_HVT U1811 ( .A1(n1128), .A2(n4235), .A3(n4222), .A4(n1384), .A5(
        n1256), .A6(n4210), .Y(n1697) );
  OA222X1_HVT U1812 ( .A1(n744), .A2(n4197), .A3(n1000), .A4(n4184), .A5(n872), 
        .A6(n4171), .Y(n1696) );
  OA222X1_HVT U1813 ( .A1(n360), .A2(n4158), .A3(n616), .A4(n4145), .A5(n488), 
        .A6(n4132), .Y(n1695) );
  OA22X1_HVT U1814 ( .A1(n232), .A2(n4119), .A3(n104), .A4(n4106), .Y(n1694)
         );
  AO22X1_HVT U1815 ( .A1(key_round[43]), .A2(n4529), .A3(n4551), .A4(n1698), 
        .Y(n2168) );
  NAND4X0_HVT U1816 ( .A1(n1699), .A2(n1700), .A3(n1701), .A4(n1702), .Y(n1698) );
  OA222X1_HVT U1817 ( .A1(n1127), .A2(n4235), .A3(n4222), .A4(n1383), .A5(
        n1255), .A6(n4210), .Y(n1702) );
  OA222X1_HVT U1818 ( .A1(n743), .A2(n4197), .A3(n999), .A4(n4184), .A5(n871), 
        .A6(n4171), .Y(n1701) );
  OA222X1_HVT U1819 ( .A1(n359), .A2(n4158), .A3(n615), .A4(n4145), .A5(n487), 
        .A6(n4132), .Y(n1700) );
  OA22X1_HVT U1820 ( .A1(n231), .A2(n4119), .A3(n103), .A4(n4106), .Y(n1699)
         );
  AO22X1_HVT U1821 ( .A1(key_round[44]), .A2(n4529), .A3(n4551), .A4(n1703), 
        .Y(n2169) );
  NAND4X0_HVT U1822 ( .A1(n1704), .A2(n1705), .A3(n1706), .A4(n1707), .Y(n1703) );
  OA222X1_HVT U1823 ( .A1(n1126), .A2(n4235), .A3(n4222), .A4(n1382), .A5(
        n1254), .A6(n4210), .Y(n1707) );
  OA222X1_HVT U1824 ( .A1(n742), .A2(n4197), .A3(n998), .A4(n4184), .A5(n870), 
        .A6(n4171), .Y(n1706) );
  OA222X1_HVT U1825 ( .A1(n358), .A2(n4158), .A3(n614), .A4(n4145), .A5(n486), 
        .A6(n4132), .Y(n1705) );
  OA22X1_HVT U1826 ( .A1(n230), .A2(n4119), .A3(n102), .A4(n4106), .Y(n1704)
         );
  AO22X1_HVT U1827 ( .A1(key_round[45]), .A2(n4529), .A3(n4551), .A4(n1708), 
        .Y(n2170) );
  NAND4X0_HVT U1828 ( .A1(n1709), .A2(n1710), .A3(n1711), .A4(n1712), .Y(n1708) );
  OA222X1_HVT U1829 ( .A1(n1125), .A2(n4235), .A3(n4222), .A4(n1381), .A5(
        n1253), .A6(n4210), .Y(n1712) );
  OA222X1_HVT U1830 ( .A1(n741), .A2(n4197), .A3(n997), .A4(n4184), .A5(n869), 
        .A6(n4171), .Y(n1711) );
  OA222X1_HVT U1831 ( .A1(n357), .A2(n4158), .A3(n613), .A4(n4145), .A5(n485), 
        .A6(n4132), .Y(n1710) );
  OA22X1_HVT U1832 ( .A1(n229), .A2(n4119), .A3(n101), .A4(n4106), .Y(n1709)
         );
  AO22X1_HVT U1833 ( .A1(key_round[46]), .A2(n4529), .A3(n4551), .A4(n1713), 
        .Y(n2171) );
  NAND4X0_HVT U1834 ( .A1(n1714), .A2(n1715), .A3(n1716), .A4(n1717), .Y(n1713) );
  OA222X1_HVT U1835 ( .A1(n1124), .A2(n4235), .A3(n4222), .A4(n1380), .A5(
        n1252), .A6(n4210), .Y(n1717) );
  OA222X1_HVT U1836 ( .A1(n740), .A2(n4197), .A3(n996), .A4(n4184), .A5(n868), 
        .A6(n4171), .Y(n1716) );
  OA222X1_HVT U1837 ( .A1(n356), .A2(n4158), .A3(n612), .A4(n4145), .A5(n484), 
        .A6(n4132), .Y(n1715) );
  OA22X1_HVT U1838 ( .A1(n228), .A2(n4119), .A3(n100), .A4(n4106), .Y(n1714)
         );
  AO22X1_HVT U1839 ( .A1(key_round[47]), .A2(n4529), .A3(n4551), .A4(n1718), 
        .Y(n2172) );
  NAND4X0_HVT U1840 ( .A1(n1719), .A2(n1720), .A3(n1721), .A4(n1722), .Y(n1718) );
  OA222X1_HVT U1841 ( .A1(n1123), .A2(n4235), .A3(n4222), .A4(n1379), .A5(
        n1251), .A6(n4210), .Y(n1722) );
  OA222X1_HVT U1842 ( .A1(n739), .A2(n4197), .A3(n995), .A4(n4184), .A5(n867), 
        .A6(n4171), .Y(n1721) );
  OA222X1_HVT U1843 ( .A1(n355), .A2(n4158), .A3(n611), .A4(n4145), .A5(n483), 
        .A6(n4132), .Y(n1720) );
  OA22X1_HVT U1844 ( .A1(n227), .A2(n4119), .A3(n99), .A4(n4106), .Y(n1719) );
  AO22X1_HVT U1845 ( .A1(key_round[48]), .A2(n4529), .A3(n4551), .A4(n1723), 
        .Y(n2173) );
  NAND4X0_HVT U1846 ( .A1(n1724), .A2(n1725), .A3(n1726), .A4(n1727), .Y(n1723) );
  OA222X1_HVT U1847 ( .A1(n1122), .A2(n4236), .A3(n1378), .A4(n4223), .A5(
        n1250), .A6(n4211), .Y(n1727) );
  OA222X1_HVT U1848 ( .A1(n738), .A2(n4198), .A3(n994), .A4(n4185), .A5(n866), 
        .A6(n4172), .Y(n1726) );
  OA222X1_HVT U1849 ( .A1(n354), .A2(n4159), .A3(n610), .A4(n4146), .A5(n482), 
        .A6(n4133), .Y(n1725) );
  OA22X1_HVT U1850 ( .A1(n226), .A2(n4120), .A3(n98), .A4(n4107), .Y(n1724) );
  AO22X1_HVT U1851 ( .A1(key_round[49]), .A2(n4529), .A3(n4551), .A4(n1728), 
        .Y(n2174) );
  NAND4X0_HVT U1852 ( .A1(n1729), .A2(n1730), .A3(n1731), .A4(n1732), .Y(n1728) );
  OA222X1_HVT U1853 ( .A1(n1121), .A2(n4236), .A3(n1377), .A4(n4223), .A5(
        n1249), .A6(n4211), .Y(n1732) );
  OA222X1_HVT U1854 ( .A1(n737), .A2(n4198), .A3(n993), .A4(n4185), .A5(n865), 
        .A6(n4172), .Y(n1731) );
  OA222X1_HVT U1855 ( .A1(n353), .A2(n4159), .A3(n609), .A4(n4146), .A5(n481), 
        .A6(n4133), .Y(n1730) );
  OA22X1_HVT U1856 ( .A1(n225), .A2(n4120), .A3(n97), .A4(n4107), .Y(n1729) );
  AO22X1_HVT U1857 ( .A1(key_round[50]), .A2(n4529), .A3(n4551), .A4(n1733), 
        .Y(n2175) );
  NAND4X0_HVT U1858 ( .A1(n1734), .A2(n1735), .A3(n1736), .A4(n1737), .Y(n1733) );
  OA222X1_HVT U1859 ( .A1(n1120), .A2(n4236), .A3(n1376), .A4(n4223), .A5(
        n1248), .A6(n4211), .Y(n1737) );
  OA222X1_HVT U1860 ( .A1(n736), .A2(n4198), .A3(n992), .A4(n4185), .A5(n864), 
        .A6(n4172), .Y(n1736) );
  OA222X1_HVT U1861 ( .A1(n352), .A2(n4159), .A3(n608), .A4(n4146), .A5(n480), 
        .A6(n4133), .Y(n1735) );
  OA22X1_HVT U1862 ( .A1(n224), .A2(n4120), .A3(n96), .A4(n4107), .Y(n1734) );
  AO22X1_HVT U1863 ( .A1(key_round[51]), .A2(n4526), .A3(n4551), .A4(n1738), 
        .Y(n2176) );
  NAND4X0_HVT U1864 ( .A1(n1739), .A2(n1740), .A3(n1741), .A4(n1742), .Y(n1738) );
  OA222X1_HVT U1865 ( .A1(n1119), .A2(n4236), .A3(n1375), .A4(n4223), .A5(
        n1247), .A6(n4211), .Y(n1742) );
  OA222X1_HVT U1866 ( .A1(n735), .A2(n4198), .A3(n991), .A4(n4185), .A5(n863), 
        .A6(n4172), .Y(n1741) );
  OA222X1_HVT U1867 ( .A1(n351), .A2(n4159), .A3(n607), .A4(n4146), .A5(n479), 
        .A6(n4133), .Y(n1740) );
  OA22X1_HVT U1868 ( .A1(n223), .A2(n4120), .A3(n95), .A4(n4107), .Y(n1739) );
  AO22X1_HVT U1869 ( .A1(key_round[52]), .A2(n4529), .A3(n4551), .A4(n1743), 
        .Y(n2177) );
  NAND4X0_HVT U1870 ( .A1(n1744), .A2(n1745), .A3(n1746), .A4(n1747), .Y(n1743) );
  OA222X1_HVT U1871 ( .A1(n1118), .A2(n4236), .A3(n1374), .A4(n4223), .A5(
        n1246), .A6(n4211), .Y(n1747) );
  OA222X1_HVT U1872 ( .A1(n734), .A2(n4198), .A3(n990), .A4(n4185), .A5(n862), 
        .A6(n4172), .Y(n1746) );
  OA222X1_HVT U1873 ( .A1(n350), .A2(n4159), .A3(n606), .A4(n4146), .A5(n478), 
        .A6(n4133), .Y(n1745) );
  OA22X1_HVT U1874 ( .A1(n222), .A2(n4120), .A3(n94), .A4(n4107), .Y(n1744) );
  AO22X1_HVT U1875 ( .A1(key_round[53]), .A2(n4529), .A3(n4551), .A4(n1748), 
        .Y(n2178) );
  NAND4X0_HVT U1876 ( .A1(n1749), .A2(n1750), .A3(n1751), .A4(n1752), .Y(n1748) );
  OA222X1_HVT U1877 ( .A1(n1117), .A2(n4236), .A3(n1373), .A4(n4223), .A5(
        n1245), .A6(n4211), .Y(n1752) );
  OA222X1_HVT U1878 ( .A1(n733), .A2(n4198), .A3(n989), .A4(n4185), .A5(n861), 
        .A6(n4172), .Y(n1751) );
  OA222X1_HVT U1879 ( .A1(n349), .A2(n4159), .A3(n605), .A4(n4146), .A5(n477), 
        .A6(n4133), .Y(n1750) );
  OA22X1_HVT U1880 ( .A1(n221), .A2(n4120), .A3(n93), .A4(n4107), .Y(n1749) );
  AO22X1_HVT U1881 ( .A1(key_round[54]), .A2(n4530), .A3(n4551), .A4(n1753), 
        .Y(n2179) );
  NAND4X0_HVT U1882 ( .A1(n1754), .A2(n1755), .A3(n1756), .A4(n1757), .Y(n1753) );
  OA222X1_HVT U1883 ( .A1(n1116), .A2(n4236), .A3(n1372), .A4(n4223), .A5(
        n1244), .A6(n4211), .Y(n1757) );
  OA222X1_HVT U1884 ( .A1(n732), .A2(n4198), .A3(n988), .A4(n4185), .A5(n860), 
        .A6(n4172), .Y(n1756) );
  OA222X1_HVT U1885 ( .A1(n348), .A2(n4159), .A3(n604), .A4(n4146), .A5(n476), 
        .A6(n4133), .Y(n1755) );
  OA22X1_HVT U1886 ( .A1(n220), .A2(n4120), .A3(n92), .A4(n4107), .Y(n1754) );
  AO22X1_HVT U1887 ( .A1(key_round[55]), .A2(n4530), .A3(n4551), .A4(n1758), 
        .Y(n2180) );
  NAND4X0_HVT U1888 ( .A1(n1759), .A2(n1760), .A3(n1761), .A4(n1762), .Y(n1758) );
  OA222X1_HVT U1889 ( .A1(n1115), .A2(n4236), .A3(n1371), .A4(n4223), .A5(
        n1243), .A6(n4211), .Y(n1762) );
  OA222X1_HVT U1890 ( .A1(n731), .A2(n4198), .A3(n987), .A4(n4185), .A5(n859), 
        .A6(n4172), .Y(n1761) );
  OA222X1_HVT U1891 ( .A1(n347), .A2(n4159), .A3(n603), .A4(n4146), .A5(n475), 
        .A6(n4133), .Y(n1760) );
  OA22X1_HVT U1892 ( .A1(n219), .A2(n4120), .A3(n91), .A4(n4107), .Y(n1759) );
  AO22X1_HVT U1893 ( .A1(key_round[56]), .A2(n4530), .A3(n4550), .A4(n1763), 
        .Y(n2181) );
  NAND4X0_HVT U1894 ( .A1(n1764), .A2(n1765), .A3(n1766), .A4(n1767), .Y(n1763) );
  OA222X1_HVT U1895 ( .A1(n1114), .A2(n4236), .A3(n1370), .A4(n4223), .A5(
        n1242), .A6(n4211), .Y(n1767) );
  OA222X1_HVT U1896 ( .A1(n730), .A2(n4198), .A3(n986), .A4(n4185), .A5(n858), 
        .A6(n4172), .Y(n1766) );
  OA222X1_HVT U1897 ( .A1(n346), .A2(n4159), .A3(n602), .A4(n4146), .A5(n474), 
        .A6(n4133), .Y(n1765) );
  OA22X1_HVT U1898 ( .A1(n218), .A2(n4120), .A3(n90), .A4(n4107), .Y(n1764) );
  AO22X1_HVT U1899 ( .A1(key_round[57]), .A2(n4530), .A3(n4550), .A4(n1768), 
        .Y(n2182) );
  NAND4X0_HVT U1900 ( .A1(n1769), .A2(n1770), .A3(n1771), .A4(n1772), .Y(n1768) );
  OA222X1_HVT U1901 ( .A1(n1113), .A2(n4236), .A3(n1369), .A4(n4223), .A5(
        n1241), .A6(n4211), .Y(n1772) );
  OA222X1_HVT U1902 ( .A1(n729), .A2(n4198), .A3(n985), .A4(n4185), .A5(n857), 
        .A6(n4172), .Y(n1771) );
  OA222X1_HVT U1903 ( .A1(n345), .A2(n4159), .A3(n601), .A4(n4146), .A5(n473), 
        .A6(n4133), .Y(n1770) );
  OA22X1_HVT U1904 ( .A1(n217), .A2(n4120), .A3(n89), .A4(n4107), .Y(n1769) );
  AO22X1_HVT U1905 ( .A1(key_round[58]), .A2(n4530), .A3(n4550), .A4(n1773), 
        .Y(n2183) );
  NAND4X0_HVT U1906 ( .A1(n1774), .A2(n1775), .A3(n1776), .A4(n1777), .Y(n1773) );
  OA222X1_HVT U1907 ( .A1(n1112), .A2(n4236), .A3(n1368), .A4(n4223), .A5(
        n1240), .A6(n4211), .Y(n1777) );
  OA222X1_HVT U1908 ( .A1(n728), .A2(n4198), .A3(n984), .A4(n4185), .A5(n856), 
        .A6(n4172), .Y(n1776) );
  OA222X1_HVT U1909 ( .A1(n344), .A2(n4159), .A3(n600), .A4(n4146), .A5(n472), 
        .A6(n4133), .Y(n1775) );
  OA22X1_HVT U1910 ( .A1(n216), .A2(n4120), .A3(n88), .A4(n4107), .Y(n1774) );
  AO22X1_HVT U1911 ( .A1(key_round[59]), .A2(n4530), .A3(n4550), .A4(n1778), 
        .Y(n2184) );
  NAND4X0_HVT U1912 ( .A1(n1779), .A2(n1780), .A3(n1781), .A4(n1782), .Y(n1778) );
  OA222X1_HVT U1913 ( .A1(n1111), .A2(n4236), .A3(n1367), .A4(n4223), .A5(
        n1239), .A6(n4211), .Y(n1782) );
  OA222X1_HVT U1914 ( .A1(n727), .A2(n4198), .A3(n983), .A4(n4185), .A5(n855), 
        .A6(n4172), .Y(n1781) );
  OA222X1_HVT U1915 ( .A1(n343), .A2(n4159), .A3(n599), .A4(n4146), .A5(n471), 
        .A6(n4133), .Y(n1780) );
  OA22X1_HVT U1916 ( .A1(n215), .A2(n4120), .A3(n87), .A4(n4107), .Y(n1779) );
  AO22X1_HVT U1917 ( .A1(key_round[60]), .A2(n4530), .A3(n4550), .A4(n1783), 
        .Y(n2185) );
  NAND4X0_HVT U1918 ( .A1(n1784), .A2(n1785), .A3(n1786), .A4(n1787), .Y(n1783) );
  OA222X1_HVT U1919 ( .A1(n1110), .A2(n4237), .A3(n1366), .A4(n4223), .A5(
        n1238), .A6(n4212), .Y(n1787) );
  OA222X1_HVT U1920 ( .A1(n726), .A2(n4199), .A3(n982), .A4(n4186), .A5(n854), 
        .A6(n4173), .Y(n1786) );
  OA222X1_HVT U1921 ( .A1(n342), .A2(n4160), .A3(n598), .A4(n4147), .A5(n470), 
        .A6(n4134), .Y(n1785) );
  OA22X1_HVT U1922 ( .A1(n214), .A2(n4121), .A3(n86), .A4(n4108), .Y(n1784) );
  AO22X1_HVT U1923 ( .A1(key_round[61]), .A2(n4530), .A3(n4550), .A4(n1788), 
        .Y(n2186) );
  NAND4X0_HVT U1924 ( .A1(n1789), .A2(n1790), .A3(n1791), .A4(n1792), .Y(n1788) );
  OA222X1_HVT U1925 ( .A1(n1109), .A2(n4237), .A3(n1365), .A4(n4224), .A5(
        n1237), .A6(n4212), .Y(n1792) );
  OA222X1_HVT U1926 ( .A1(n725), .A2(n4199), .A3(n981), .A4(n4186), .A5(n853), 
        .A6(n4173), .Y(n1791) );
  OA222X1_HVT U1927 ( .A1(n341), .A2(n4160), .A3(n597), .A4(n4147), .A5(n469), 
        .A6(n4134), .Y(n1790) );
  OA22X1_HVT U1928 ( .A1(n213), .A2(n4121), .A3(n85), .A4(n4108), .Y(n1789) );
  AO22X1_HVT U1929 ( .A1(key_round[62]), .A2(n4530), .A3(n4550), .A4(n1793), 
        .Y(n2187) );
  NAND4X0_HVT U1930 ( .A1(n1794), .A2(n1795), .A3(n1796), .A4(n1797), .Y(n1793) );
  OA222X1_HVT U1931 ( .A1(n1108), .A2(n4237), .A3(n1364), .A4(n4224), .A5(
        n1236), .A6(n4212), .Y(n1797) );
  OA222X1_HVT U1932 ( .A1(n724), .A2(n4199), .A3(n980), .A4(n4186), .A5(n852), 
        .A6(n4173), .Y(n1796) );
  OA222X1_HVT U1933 ( .A1(n340), .A2(n4160), .A3(n596), .A4(n4147), .A5(n468), 
        .A6(n4134), .Y(n1795) );
  OA22X1_HVT U1934 ( .A1(n212), .A2(n4121), .A3(n84), .A4(n4108), .Y(n1794) );
  AO22X1_HVT U1935 ( .A1(key_round[63]), .A2(n4530), .A3(n4550), .A4(n1798), 
        .Y(n2188) );
  NAND4X0_HVT U1936 ( .A1(n1799), .A2(n1800), .A3(n1801), .A4(n1802), .Y(n1798) );
  OA222X1_HVT U1937 ( .A1(n1107), .A2(n4237), .A3(n1363), .A4(n4224), .A5(
        n1235), .A6(n4212), .Y(n1802) );
  OA222X1_HVT U1938 ( .A1(n723), .A2(n4199), .A3(n979), .A4(n4186), .A5(n851), 
        .A6(n4173), .Y(n1801) );
  OA222X1_HVT U1939 ( .A1(n339), .A2(n4160), .A3(n595), .A4(n4147), .A5(n467), 
        .A6(n4134), .Y(n1800) );
  OA22X1_HVT U1940 ( .A1(n211), .A2(n4121), .A3(n83), .A4(n4108), .Y(n1799) );
  AO22X1_HVT U1941 ( .A1(key_round[64]), .A2(n4530), .A3(n4550), .A4(n1803), 
        .Y(n2189) );
  NAND4X0_HVT U1942 ( .A1(n1804), .A2(n1805), .A3(n1806), .A4(n1807), .Y(n1803) );
  OA222X1_HVT U1943 ( .A1(n1106), .A2(n4237), .A3(n1362), .A4(n4224), .A5(
        n1234), .A6(n4212), .Y(n1807) );
  OA222X1_HVT U1944 ( .A1(n722), .A2(n4199), .A3(n978), .A4(n4186), .A5(n850), 
        .A6(n4173), .Y(n1806) );
  OA222X1_HVT U1945 ( .A1(n338), .A2(n4160), .A3(n594), .A4(n4147), .A5(n466), 
        .A6(n4134), .Y(n1805) );
  OA22X1_HVT U1946 ( .A1(n210), .A2(n4121), .A3(n82), .A4(n4108), .Y(n1804) );
  AO22X1_HVT U1947 ( .A1(key_round[65]), .A2(n4530), .A3(n4550), .A4(n1808), 
        .Y(n2190) );
  NAND4X0_HVT U1948 ( .A1(n1809), .A2(n1810), .A3(n1811), .A4(n1812), .Y(n1808) );
  OA222X1_HVT U1949 ( .A1(n1105), .A2(n4237), .A3(n1361), .A4(n4224), .A5(
        n1233), .A6(n4212), .Y(n1812) );
  OA222X1_HVT U1950 ( .A1(n721), .A2(n4199), .A3(n977), .A4(n4186), .A5(n849), 
        .A6(n4173), .Y(n1811) );
  OA222X1_HVT U1951 ( .A1(n337), .A2(n4160), .A3(n593), .A4(n4147), .A5(n465), 
        .A6(n4134), .Y(n1810) );
  OA22X1_HVT U1952 ( .A1(n209), .A2(n4121), .A3(n81), .A4(n4108), .Y(n1809) );
  AO22X1_HVT U1953 ( .A1(key_round[66]), .A2(n4531), .A3(n4550), .A4(n1813), 
        .Y(n2191) );
  NAND4X0_HVT U1954 ( .A1(n1814), .A2(n1815), .A3(n1816), .A4(n1817), .Y(n1813) );
  OA222X1_HVT U1955 ( .A1(n1104), .A2(n4237), .A3(n1360), .A4(n4224), .A5(
        n1232), .A6(n4212), .Y(n1817) );
  OA222X1_HVT U1956 ( .A1(n720), .A2(n4199), .A3(n976), .A4(n4186), .A5(n848), 
        .A6(n4173), .Y(n1816) );
  OA222X1_HVT U1957 ( .A1(n336), .A2(n4160), .A3(n592), .A4(n4147), .A5(n464), 
        .A6(n4134), .Y(n1815) );
  OA22X1_HVT U1958 ( .A1(n208), .A2(n4121), .A3(n80), .A4(n4108), .Y(n1814) );
  AO22X1_HVT U1959 ( .A1(key_round[67]), .A2(n4531), .A3(n4550), .A4(n1818), 
        .Y(n2192) );
  NAND4X0_HVT U1960 ( .A1(n1819), .A2(n1820), .A3(n1821), .A4(n1822), .Y(n1818) );
  OA222X1_HVT U1961 ( .A1(n1103), .A2(n4237), .A3(n1359), .A4(n4224), .A5(
        n1231), .A6(n4212), .Y(n1822) );
  OA222X1_HVT U1962 ( .A1(n719), .A2(n4199), .A3(n975), .A4(n4186), .A5(n847), 
        .A6(n4173), .Y(n1821) );
  OA222X1_HVT U1963 ( .A1(n335), .A2(n4160), .A3(n591), .A4(n4147), .A5(n463), 
        .A6(n4134), .Y(n1820) );
  OA22X1_HVT U1964 ( .A1(n207), .A2(n4121), .A3(n79), .A4(n4108), .Y(n1819) );
  AO22X1_HVT U1965 ( .A1(key_round[68]), .A2(n4531), .A3(n4550), .A4(n1823), 
        .Y(n2193) );
  NAND4X0_HVT U1966 ( .A1(n1824), .A2(n1825), .A3(n1826), .A4(n1827), .Y(n1823) );
  OA222X1_HVT U1967 ( .A1(n1102), .A2(n4237), .A3(n1358), .A4(n4224), .A5(
        n1230), .A6(n4212), .Y(n1827) );
  OA222X1_HVT U1968 ( .A1(n718), .A2(n4199), .A3(n974), .A4(n4186), .A5(n846), 
        .A6(n4173), .Y(n1826) );
  OA222X1_HVT U1969 ( .A1(n334), .A2(n4160), .A3(n590), .A4(n4147), .A5(n462), 
        .A6(n4134), .Y(n1825) );
  OA22X1_HVT U1970 ( .A1(n206), .A2(n4121), .A3(n78), .A4(n4108), .Y(n1824) );
  AO22X1_HVT U1971 ( .A1(key_round[69]), .A2(n4531), .A3(n4550), .A4(n1828), 
        .Y(n2194) );
  NAND4X0_HVT U1972 ( .A1(n1829), .A2(n1830), .A3(n1831), .A4(n1832), .Y(n1828) );
  OA222X1_HVT U1973 ( .A1(n1101), .A2(n4237), .A3(n1357), .A4(n4224), .A5(
        n1229), .A6(n4212), .Y(n1832) );
  OA222X1_HVT U1974 ( .A1(n717), .A2(n4199), .A3(n973), .A4(n4186), .A5(n845), 
        .A6(n4173), .Y(n1831) );
  OA222X1_HVT U1975 ( .A1(n333), .A2(n4160), .A3(n589), .A4(n4147), .A5(n461), 
        .A6(n4134), .Y(n1830) );
  OA22X1_HVT U1976 ( .A1(n205), .A2(n4121), .A3(n77), .A4(n4108), .Y(n1829) );
  AO22X1_HVT U1977 ( .A1(key_round[70]), .A2(n4531), .A3(n4550), .A4(n1833), 
        .Y(n2195) );
  NAND4X0_HVT U1978 ( .A1(n1834), .A2(n1835), .A3(n1836), .A4(n1837), .Y(n1833) );
  OA222X1_HVT U1979 ( .A1(n1100), .A2(n4237), .A3(n1356), .A4(n4224), .A5(
        n1228), .A6(n4212), .Y(n1837) );
  OA222X1_HVT U1980 ( .A1(n716), .A2(n4199), .A3(n972), .A4(n4186), .A5(n844), 
        .A6(n4173), .Y(n1836) );
  OA222X1_HVT U1981 ( .A1(n332), .A2(n4160), .A3(n588), .A4(n4147), .A5(n460), 
        .A6(n4134), .Y(n1835) );
  OA22X1_HVT U1982 ( .A1(n204), .A2(n4121), .A3(n76), .A4(n4108), .Y(n1834) );
  AO22X1_HVT U1983 ( .A1(key_round[71]), .A2(n4531), .A3(n4549), .A4(n1838), 
        .Y(n2196) );
  NAND4X0_HVT U1984 ( .A1(n1839), .A2(n1840), .A3(n1841), .A4(n1842), .Y(n1838) );
  OA222X1_HVT U1985 ( .A1(n1099), .A2(n4237), .A3(n1355), .A4(n4224), .A5(
        n1227), .A6(n4212), .Y(n1842) );
  OA222X1_HVT U1986 ( .A1(n715), .A2(n4199), .A3(n971), .A4(n4186), .A5(n843), 
        .A6(n4173), .Y(n1841) );
  OA222X1_HVT U1987 ( .A1(n331), .A2(n4160), .A3(n587), .A4(n4147), .A5(n459), 
        .A6(n4134), .Y(n1840) );
  OA22X1_HVT U1988 ( .A1(n203), .A2(n4121), .A3(n75), .A4(n4108), .Y(n1839) );
  AO22X1_HVT U1989 ( .A1(key_round[72]), .A2(n4531), .A3(n4549), .A4(n1843), 
        .Y(n2197) );
  NAND4X0_HVT U1990 ( .A1(n1844), .A2(n1845), .A3(n1846), .A4(n1847), .Y(n1843) );
  OA222X1_HVT U1991 ( .A1(n1098), .A2(n4238), .A3(n1354), .A4(n4224), .A5(
        n1226), .A6(n4213), .Y(n1847) );
  OA222X1_HVT U1992 ( .A1(n714), .A2(n4200), .A3(n970), .A4(n4187), .A5(n842), 
        .A6(n4174), .Y(n1846) );
  OA222X1_HVT U1993 ( .A1(n330), .A2(n4161), .A3(n586), .A4(n4148), .A5(n458), 
        .A6(n4135), .Y(n1845) );
  OA22X1_HVT U1994 ( .A1(n202), .A2(n4122), .A3(n74), .A4(n4109), .Y(n1844) );
  AO22X1_HVT U1995 ( .A1(key_round[73]), .A2(n4531), .A3(n4549), .A4(n1848), 
        .Y(n2198) );
  NAND4X0_HVT U1996 ( .A1(n1849), .A2(n1850), .A3(n1851), .A4(n1852), .Y(n1848) );
  OA222X1_HVT U1997 ( .A1(n1097), .A2(n4238), .A3(n1353), .A4(n4224), .A5(
        n1225), .A6(n4213), .Y(n1852) );
  OA222X1_HVT U1998 ( .A1(n713), .A2(n4200), .A3(n969), .A4(n4187), .A5(n841), 
        .A6(n4174), .Y(n1851) );
  OA222X1_HVT U1999 ( .A1(n329), .A2(n4161), .A3(n585), .A4(n4148), .A5(n457), 
        .A6(n4135), .Y(n1850) );
  OA22X1_HVT U2000 ( .A1(n201), .A2(n4122), .A3(n73), .A4(n4109), .Y(n1849) );
  AO22X1_HVT U2001 ( .A1(key_round[74]), .A2(n4531), .A3(n4549), .A4(n1853), 
        .Y(n2199) );
  NAND4X0_HVT U2002 ( .A1(n1854), .A2(n1855), .A3(n1856), .A4(n1857), .Y(n1853) );
  OA222X1_HVT U2003 ( .A1(n1096), .A2(n4238), .A3(n1352), .A4(n4225), .A5(
        n1224), .A6(n4213), .Y(n1857) );
  OA222X1_HVT U2004 ( .A1(n712), .A2(n4200), .A3(n968), .A4(n4187), .A5(n840), 
        .A6(n4174), .Y(n1856) );
  OA222X1_HVT U2005 ( .A1(n328), .A2(n4161), .A3(n584), .A4(n4148), .A5(n456), 
        .A6(n4135), .Y(n1855) );
  OA22X1_HVT U2006 ( .A1(n200), .A2(n4122), .A3(n72), .A4(n4109), .Y(n1854) );
  AO22X1_HVT U2007 ( .A1(key_round[75]), .A2(n4531), .A3(n4549), .A4(n1858), 
        .Y(n2200) );
  NAND4X0_HVT U2008 ( .A1(n1859), .A2(n1860), .A3(n1861), .A4(n1862), .Y(n1858) );
  OA222X1_HVT U2009 ( .A1(n1095), .A2(n4238), .A3(n1351), .A4(n4225), .A5(
        n1223), .A6(n4213), .Y(n1862) );
  OA222X1_HVT U2010 ( .A1(n711), .A2(n4200), .A3(n967), .A4(n4187), .A5(n839), 
        .A6(n4174), .Y(n1861) );
  OA222X1_HVT U2011 ( .A1(n327), .A2(n4161), .A3(n583), .A4(n4148), .A5(n455), 
        .A6(n4135), .Y(n1860) );
  OA22X1_HVT U2012 ( .A1(n199), .A2(n4122), .A3(n71), .A4(n4109), .Y(n1859) );
  AO22X1_HVT U2013 ( .A1(key_round[76]), .A2(n4531), .A3(n4549), .A4(n1863), 
        .Y(n2201) );
  NAND4X0_HVT U2014 ( .A1(n1864), .A2(n1865), .A3(n1866), .A4(n1867), .Y(n1863) );
  OA222X1_HVT U2015 ( .A1(n1094), .A2(n4238), .A3(n1350), .A4(n4225), .A5(
        n1222), .A6(n4213), .Y(n1867) );
  OA222X1_HVT U2016 ( .A1(n710), .A2(n4200), .A3(n966), .A4(n4187), .A5(n838), 
        .A6(n4174), .Y(n1866) );
  OA222X1_HVT U2017 ( .A1(n326), .A2(n4161), .A3(n582), .A4(n4148), .A5(n454), 
        .A6(n4135), .Y(n1865) );
  OA22X1_HVT U2018 ( .A1(n198), .A2(n4122), .A3(n70), .A4(n4109), .Y(n1864) );
  AO22X1_HVT U2019 ( .A1(key_round[77]), .A2(n4531), .A3(n4549), .A4(n1868), 
        .Y(n2202) );
  NAND4X0_HVT U2020 ( .A1(n1869), .A2(n1870), .A3(n1871), .A4(n1872), .Y(n1868) );
  OA222X1_HVT U2021 ( .A1(n1093), .A2(n4238), .A3(n1349), .A4(n4225), .A5(
        n1221), .A6(n4213), .Y(n1872) );
  OA222X1_HVT U2022 ( .A1(n709), .A2(n4200), .A3(n965), .A4(n4187), .A5(n837), 
        .A6(n4174), .Y(n1871) );
  OA222X1_HVT U2023 ( .A1(n325), .A2(n4161), .A3(n581), .A4(n4148), .A5(n453), 
        .A6(n4135), .Y(n1870) );
  OA22X1_HVT U2024 ( .A1(n197), .A2(n4122), .A3(n69), .A4(n4109), .Y(n1869) );
  AO22X1_HVT U2025 ( .A1(key_round[78]), .A2(n4532), .A3(n4549), .A4(n1873), 
        .Y(n2203) );
  NAND4X0_HVT U2026 ( .A1(n1874), .A2(n1875), .A3(n1876), .A4(n1877), .Y(n1873) );
  OA222X1_HVT U2027 ( .A1(n1092), .A2(n4238), .A3(n1348), .A4(n4225), .A5(
        n1220), .A6(n4213), .Y(n1877) );
  OA222X1_HVT U2028 ( .A1(n708), .A2(n4200), .A3(n964), .A4(n4187), .A5(n836), 
        .A6(n4174), .Y(n1876) );
  OA222X1_HVT U2029 ( .A1(n324), .A2(n4161), .A3(n580), .A4(n4148), .A5(n452), 
        .A6(n4135), .Y(n1875) );
  OA22X1_HVT U2030 ( .A1(n196), .A2(n4122), .A3(n68), .A4(n4109), .Y(n1874) );
  AO22X1_HVT U2031 ( .A1(key_round[79]), .A2(n4532), .A3(n4549), .A4(n1878), 
        .Y(n2204) );
  NAND4X0_HVT U2032 ( .A1(n1879), .A2(n1880), .A3(n1881), .A4(n1882), .Y(n1878) );
  OA222X1_HVT U2033 ( .A1(n1091), .A2(n4238), .A3(n1347), .A4(n4225), .A5(
        n1219), .A6(n4213), .Y(n1882) );
  OA222X1_HVT U2034 ( .A1(n707), .A2(n4200), .A3(n963), .A4(n4187), .A5(n835), 
        .A6(n4174), .Y(n1881) );
  OA222X1_HVT U2035 ( .A1(n323), .A2(n4161), .A3(n579), .A4(n4148), .A5(n451), 
        .A6(n4135), .Y(n1880) );
  OA22X1_HVT U2036 ( .A1(n195), .A2(n4122), .A3(n67), .A4(n4109), .Y(n1879) );
  AO22X1_HVT U2037 ( .A1(key_round[80]), .A2(n4532), .A3(n4549), .A4(n1883), 
        .Y(n2205) );
  NAND4X0_HVT U2038 ( .A1(n1884), .A2(n1885), .A3(n1886), .A4(n1887), .Y(n1883) );
  OA222X1_HVT U2039 ( .A1(n1090), .A2(n4238), .A3(n1346), .A4(n4225), .A5(
        n1218), .A6(n4213), .Y(n1887) );
  OA222X1_HVT U2040 ( .A1(n706), .A2(n4200), .A3(n962), .A4(n4187), .A5(n834), 
        .A6(n4174), .Y(n1886) );
  OA222X1_HVT U2041 ( .A1(n322), .A2(n4161), .A3(n578), .A4(n4148), .A5(n450), 
        .A6(n4135), .Y(n1885) );
  OA22X1_HVT U2042 ( .A1(n194), .A2(n4122), .A3(n66), .A4(n4109), .Y(n1884) );
  AO22X1_HVT U2043 ( .A1(key_round[81]), .A2(n4532), .A3(n4549), .A4(n1888), 
        .Y(n2206) );
  NAND4X0_HVT U2044 ( .A1(n1889), .A2(n1890), .A3(n1891), .A4(n1892), .Y(n1888) );
  OA222X1_HVT U2045 ( .A1(n1089), .A2(n4238), .A3(n1345), .A4(n4225), .A5(
        n1217), .A6(n4213), .Y(n1892) );
  OA222X1_HVT U2046 ( .A1(n705), .A2(n4200), .A3(n961), .A4(n4187), .A5(n833), 
        .A6(n4174), .Y(n1891) );
  OA222X1_HVT U2047 ( .A1(n321), .A2(n4161), .A3(n577), .A4(n4148), .A5(n449), 
        .A6(n4135), .Y(n1890) );
  OA22X1_HVT U2048 ( .A1(n193), .A2(n4122), .A3(n65), .A4(n4109), .Y(n1889) );
  AO22X1_HVT U2049 ( .A1(key_round[82]), .A2(n4532), .A3(n4549), .A4(n1893), 
        .Y(n2207) );
  NAND4X0_HVT U2050 ( .A1(n1894), .A2(n1895), .A3(n1896), .A4(n1897), .Y(n1893) );
  OA222X1_HVT U2051 ( .A1(n1088), .A2(n4238), .A3(n1344), .A4(n4225), .A5(
        n1216), .A6(n4213), .Y(n1897) );
  OA222X1_HVT U2052 ( .A1(n704), .A2(n4200), .A3(n960), .A4(n4187), .A5(n832), 
        .A6(n4174), .Y(n1896) );
  OA222X1_HVT U2053 ( .A1(n320), .A2(n4161), .A3(n576), .A4(n4148), .A5(n448), 
        .A6(n4135), .Y(n1895) );
  OA22X1_HVT U2054 ( .A1(n192), .A2(n4122), .A3(n64), .A4(n4109), .Y(n1894) );
  AO22X1_HVT U2055 ( .A1(key_round[83]), .A2(n4532), .A3(n4549), .A4(n1898), 
        .Y(n2208) );
  NAND4X0_HVT U2056 ( .A1(n1899), .A2(n1900), .A3(n1901), .A4(n1902), .Y(n1898) );
  OA222X1_HVT U2057 ( .A1(n1087), .A2(n4238), .A3(n1343), .A4(n4225), .A5(
        n1215), .A6(n4213), .Y(n1902) );
  OA222X1_HVT U2058 ( .A1(n703), .A2(n4200), .A3(n959), .A4(n4187), .A5(n831), 
        .A6(n4174), .Y(n1901) );
  OA222X1_HVT U2059 ( .A1(n319), .A2(n4161), .A3(n575), .A4(n4148), .A5(n447), 
        .A6(n4135), .Y(n1900) );
  OA22X1_HVT U2060 ( .A1(n191), .A2(n4122), .A3(n63), .A4(n4109), .Y(n1899) );
  AO22X1_HVT U2061 ( .A1(key_round[84]), .A2(n4532), .A3(n4549), .A4(n1903), 
        .Y(n2209) );
  NAND4X0_HVT U2062 ( .A1(n1904), .A2(n1905), .A3(n1906), .A4(n1907), .Y(n1903) );
  OA222X1_HVT U2063 ( .A1(n1086), .A2(n4239), .A3(n1342), .A4(n4225), .A5(
        n1214), .A6(n4214), .Y(n1907) );
  OA222X1_HVT U2064 ( .A1(n702), .A2(n4201), .A3(n958), .A4(n4188), .A5(n830), 
        .A6(n4175), .Y(n1906) );
  OA222X1_HVT U2065 ( .A1(n318), .A2(n4162), .A3(n574), .A4(n4149), .A5(n446), 
        .A6(n4136), .Y(n1905) );
  OA22X1_HVT U2066 ( .A1(n190), .A2(n4123), .A3(n62), .A4(n4110), .Y(n1904) );
  AO22X1_HVT U2067 ( .A1(key_round[85]), .A2(n4532), .A3(n4549), .A4(n1908), 
        .Y(n2210) );
  NAND4X0_HVT U2068 ( .A1(n1909), .A2(n1910), .A3(n1911), .A4(n1912), .Y(n1908) );
  OA222X1_HVT U2069 ( .A1(n1085), .A2(n4239), .A3(n1341), .A4(n4225), .A5(
        n1213), .A6(n4214), .Y(n1912) );
  OA222X1_HVT U2070 ( .A1(n701), .A2(n4201), .A3(n957), .A4(n4188), .A5(n829), 
        .A6(n4175), .Y(n1911) );
  OA222X1_HVT U2071 ( .A1(n317), .A2(n4162), .A3(n573), .A4(n4149), .A5(n445), 
        .A6(n4136), .Y(n1910) );
  OA22X1_HVT U2072 ( .A1(n189), .A2(n4123), .A3(n61), .A4(n4110), .Y(n1909) );
  AO22X1_HVT U2073 ( .A1(key_round[86]), .A2(n4532), .A3(n4548), .A4(n1913), 
        .Y(n2211) );
  NAND4X0_HVT U2074 ( .A1(n1914), .A2(n1915), .A3(n1916), .A4(n1917), .Y(n1913) );
  OA222X1_HVT U2075 ( .A1(n1084), .A2(n4239), .A3(n1340), .A4(n4225), .A5(
        n1212), .A6(n4214), .Y(n1917) );
  OA222X1_HVT U2076 ( .A1(n700), .A2(n4201), .A3(n956), .A4(n4188), .A5(n828), 
        .A6(n4175), .Y(n1916) );
  OA222X1_HVT U2077 ( .A1(n316), .A2(n4162), .A3(n572), .A4(n4149), .A5(n444), 
        .A6(n4136), .Y(n1915) );
  OA22X1_HVT U2078 ( .A1(n188), .A2(n4123), .A3(n60), .A4(n4110), .Y(n1914) );
  AO22X1_HVT U2079 ( .A1(key_round[87]), .A2(n4532), .A3(n4548), .A4(n1918), 
        .Y(n2212) );
  NAND4X0_HVT U2080 ( .A1(n1919), .A2(n1920), .A3(n1921), .A4(n1922), .Y(n1918) );
  OA222X1_HVT U2081 ( .A1(n1083), .A2(n4239), .A3(n1339), .A4(n4226), .A5(
        n1211), .A6(n4214), .Y(n1922) );
  OA222X1_HVT U2082 ( .A1(n699), .A2(n4201), .A3(n955), .A4(n4188), .A5(n827), 
        .A6(n4175), .Y(n1921) );
  OA222X1_HVT U2083 ( .A1(n315), .A2(n4162), .A3(n571), .A4(n4149), .A5(n443), 
        .A6(n4136), .Y(n1920) );
  OA22X1_HVT U2084 ( .A1(n187), .A2(n4123), .A3(n59), .A4(n4110), .Y(n1919) );
  AO22X1_HVT U2085 ( .A1(key_round[88]), .A2(n4532), .A3(n4548), .A4(n1923), 
        .Y(n2213) );
  NAND4X0_HVT U2086 ( .A1(n1924), .A2(n1925), .A3(n1926), .A4(n1927), .Y(n1923) );
  OA222X1_HVT U2087 ( .A1(n1082), .A2(n4239), .A3(n1338), .A4(n4226), .A5(
        n1210), .A6(n4214), .Y(n1927) );
  OA222X1_HVT U2088 ( .A1(n698), .A2(n4201), .A3(n954), .A4(n4188), .A5(n826), 
        .A6(n4175), .Y(n1926) );
  OA222X1_HVT U2089 ( .A1(n314), .A2(n4162), .A3(n570), .A4(n4149), .A5(n442), 
        .A6(n4136), .Y(n1925) );
  OA22X1_HVT U2090 ( .A1(n186), .A2(n4123), .A3(n58), .A4(n4110), .Y(n1924) );
  AO22X1_HVT U2091 ( .A1(key_round[89]), .A2(n4532), .A3(n4548), .A4(n1928), 
        .Y(n2214) );
  NAND4X0_HVT U2092 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .Y(n1928) );
  OA222X1_HVT U2093 ( .A1(n1081), .A2(n4239), .A3(n1337), .A4(n4226), .A5(
        n1209), .A6(n4214), .Y(n1932) );
  OA222X1_HVT U2094 ( .A1(n697), .A2(n4201), .A3(n953), .A4(n4188), .A5(n825), 
        .A6(n4175), .Y(n1931) );
  OA222X1_HVT U2095 ( .A1(n313), .A2(n4162), .A3(n569), .A4(n4149), .A5(n441), 
        .A6(n4136), .Y(n1930) );
  OA22X1_HVT U2096 ( .A1(n185), .A2(n4123), .A3(n57), .A4(n4110), .Y(n1929) );
  AO22X1_HVT U2097 ( .A1(key_round[90]), .A2(n4533), .A3(n4548), .A4(n1933), 
        .Y(n2215) );
  NAND4X0_HVT U2098 ( .A1(n1934), .A2(n1935), .A3(n1936), .A4(n1937), .Y(n1933) );
  OA222X1_HVT U2099 ( .A1(n1080), .A2(n4239), .A3(n1336), .A4(n4226), .A5(
        n1208), .A6(n4214), .Y(n1937) );
  OA222X1_HVT U2100 ( .A1(n696), .A2(n4201), .A3(n952), .A4(n4188), .A5(n824), 
        .A6(n4175), .Y(n1936) );
  OA222X1_HVT U2101 ( .A1(n312), .A2(n4162), .A3(n568), .A4(n4149), .A5(n440), 
        .A6(n4136), .Y(n1935) );
  OA22X1_HVT U2102 ( .A1(n184), .A2(n4123), .A3(n56), .A4(n4110), .Y(n1934) );
  AO22X1_HVT U2103 ( .A1(key_round[91]), .A2(n4533), .A3(n4548), .A4(n1938), 
        .Y(n2216) );
  NAND4X0_HVT U2104 ( .A1(n1939), .A2(n1940), .A3(n1941), .A4(n1942), .Y(n1938) );
  OA222X1_HVT U2105 ( .A1(n1079), .A2(n4239), .A3(n1335), .A4(n4226), .A5(
        n1207), .A6(n4214), .Y(n1942) );
  OA222X1_HVT U2106 ( .A1(n695), .A2(n4201), .A3(n951), .A4(n4188), .A5(n823), 
        .A6(n4175), .Y(n1941) );
  OA222X1_HVT U2107 ( .A1(n311), .A2(n4162), .A3(n567), .A4(n4149), .A5(n439), 
        .A6(n4136), .Y(n1940) );
  OA22X1_HVT U2108 ( .A1(n183), .A2(n4123), .A3(n55), .A4(n4110), .Y(n1939) );
  AO22X1_HVT U2109 ( .A1(key_round[92]), .A2(n4533), .A3(n4548), .A4(n1943), 
        .Y(n2217) );
  NAND4X0_HVT U2110 ( .A1(n1944), .A2(n1945), .A3(n1946), .A4(n1947), .Y(n1943) );
  OA222X1_HVT U2111 ( .A1(n1078), .A2(n4239), .A3(n1334), .A4(n4226), .A5(
        n1206), .A6(n4214), .Y(n1947) );
  OA222X1_HVT U2112 ( .A1(n694), .A2(n4201), .A3(n950), .A4(n4188), .A5(n822), 
        .A6(n4175), .Y(n1946) );
  OA222X1_HVT U2113 ( .A1(n310), .A2(n4162), .A3(n566), .A4(n4149), .A5(n438), 
        .A6(n4136), .Y(n1945) );
  OA22X1_HVT U2114 ( .A1(n182), .A2(n4123), .A3(n54), .A4(n4110), .Y(n1944) );
  AO22X1_HVT U2115 ( .A1(key_round[93]), .A2(n4533), .A3(n4548), .A4(n1948), 
        .Y(n2218) );
  NAND4X0_HVT U2116 ( .A1(n1949), .A2(n1950), .A3(n1951), .A4(n1952), .Y(n1948) );
  OA222X1_HVT U2117 ( .A1(n1077), .A2(n4239), .A3(n1333), .A4(n4226), .A5(
        n1205), .A6(n4214), .Y(n1952) );
  OA222X1_HVT U2118 ( .A1(n693), .A2(n4201), .A3(n949), .A4(n4188), .A5(n821), 
        .A6(n4175), .Y(n1951) );
  OA222X1_HVT U2119 ( .A1(n309), .A2(n4162), .A3(n565), .A4(n4149), .A5(n437), 
        .A6(n4136), .Y(n1950) );
  OA22X1_HVT U2120 ( .A1(n181), .A2(n4123), .A3(n53), .A4(n4110), .Y(n1949) );
  AO22X1_HVT U2121 ( .A1(key_round[94]), .A2(n4522), .A3(n4548), .A4(n1953), 
        .Y(n2219) );
  NAND4X0_HVT U2122 ( .A1(n1954), .A2(n1955), .A3(n1956), .A4(n1957), .Y(n1953) );
  OA222X1_HVT U2123 ( .A1(n1076), .A2(n4239), .A3(n1332), .A4(n4226), .A5(
        n1204), .A6(n4214), .Y(n1957) );
  OA222X1_HVT U2124 ( .A1(n692), .A2(n4201), .A3(n948), .A4(n4188), .A5(n820), 
        .A6(n4175), .Y(n1956) );
  OA222X1_HVT U2125 ( .A1(n308), .A2(n4162), .A3(n564), .A4(n4149), .A5(n436), 
        .A6(n4136), .Y(n1955) );
  OA22X1_HVT U2126 ( .A1(n180), .A2(n4123), .A3(n52), .A4(n4110), .Y(n1954) );
  AO22X1_HVT U2127 ( .A1(key_round[95]), .A2(n4525), .A3(n4548), .A4(n1958), 
        .Y(n2220) );
  NAND4X0_HVT U2128 ( .A1(n1959), .A2(n1960), .A3(n1961), .A4(n1962), .Y(n1958) );
  OA222X1_HVT U2129 ( .A1(n1075), .A2(n4239), .A3(n1331), .A4(n4226), .A5(
        n1203), .A6(n4214), .Y(n1962) );
  OA222X1_HVT U2130 ( .A1(n691), .A2(n4201), .A3(n947), .A4(n4188), .A5(n819), 
        .A6(n4175), .Y(n1961) );
  OA222X1_HVT U2131 ( .A1(n307), .A2(n4162), .A3(n563), .A4(n4149), .A5(n435), 
        .A6(n4136), .Y(n1960) );
  OA22X1_HVT U2132 ( .A1(n179), .A2(n4123), .A3(n51), .A4(n4110), .Y(n1959) );
  AO22X1_HVT U2133 ( .A1(key_round[96]), .A2(n4525), .A3(n4548), .A4(n1963), 
        .Y(n2221) );
  NAND4X0_HVT U2134 ( .A1(n1964), .A2(n1965), .A3(n1966), .A4(n1967), .Y(n1963) );
  OA222X1_HVT U2135 ( .A1(n1074), .A2(n4240), .A3(n1330), .A4(n4226), .A5(
        n1202), .A6(n4215), .Y(n1967) );
  OA222X1_HVT U2136 ( .A1(n690), .A2(n4202), .A3(n946), .A4(n4189), .A5(n818), 
        .A6(n4176), .Y(n1966) );
  OA222X1_HVT U2137 ( .A1(n306), .A2(n4163), .A3(n562), .A4(n4150), .A5(n434), 
        .A6(n4137), .Y(n1965) );
  OA22X1_HVT U2138 ( .A1(n178), .A2(n4124), .A3(n50), .A4(n4111), .Y(n1964) );
  AO22X1_HVT U2139 ( .A1(key_round[97]), .A2(n4525), .A3(n4548), .A4(n1968), 
        .Y(n2222) );
  NAND4X0_HVT U2140 ( .A1(n1969), .A2(n1970), .A3(n1971), .A4(n1972), .Y(n1968) );
  OA222X1_HVT U2141 ( .A1(n1073), .A2(n4240), .A3(n1329), .A4(n4226), .A5(
        n1201), .A6(n4215), .Y(n1972) );
  OA222X1_HVT U2142 ( .A1(n689), .A2(n4202), .A3(n945), .A4(n4189), .A5(n817), 
        .A6(n4176), .Y(n1971) );
  OA222X1_HVT U2143 ( .A1(n305), .A2(n4163), .A3(n561), .A4(n4150), .A5(n433), 
        .A6(n4137), .Y(n1970) );
  OA22X1_HVT U2144 ( .A1(n177), .A2(n4124), .A3(n49), .A4(n4111), .Y(n1969) );
  AO22X1_HVT U2145 ( .A1(key_round[98]), .A2(n4525), .A3(n4548), .A4(n1973), 
        .Y(n2223) );
  NAND4X0_HVT U2146 ( .A1(n1974), .A2(n1975), .A3(n1976), .A4(n1977), .Y(n1973) );
  OA222X1_HVT U2147 ( .A1(n1072), .A2(n4240), .A3(n1328), .A4(n4226), .A5(
        n1200), .A6(n4215), .Y(n1977) );
  OA222X1_HVT U2148 ( .A1(n688), .A2(n4202), .A3(n944), .A4(n4189), .A5(n816), 
        .A6(n4176), .Y(n1976) );
  OA222X1_HVT U2149 ( .A1(n304), .A2(n4163), .A3(n560), .A4(n4150), .A5(n432), 
        .A6(n4137), .Y(n1975) );
  OA22X1_HVT U2150 ( .A1(n176), .A2(n4124), .A3(n48), .A4(n4111), .Y(n1974) );
  AO22X1_HVT U2151 ( .A1(key_round[99]), .A2(n4525), .A3(n4548), .A4(n1978), 
        .Y(n2224) );
  NAND4X0_HVT U2152 ( .A1(n1979), .A2(n1980), .A3(n1981), .A4(n1982), .Y(n1978) );
  OA222X1_HVT U2153 ( .A1(n1071), .A2(n4240), .A3(n1327), .A4(n4226), .A5(
        n1199), .A6(n4215), .Y(n1982) );
  OA222X1_HVT U2154 ( .A1(n687), .A2(n4202), .A3(n943), .A4(n4189), .A5(n815), 
        .A6(n4176), .Y(n1981) );
  OA222X1_HVT U2155 ( .A1(n303), .A2(n4163), .A3(n559), .A4(n4150), .A5(n431), 
        .A6(n4137), .Y(n1980) );
  OA22X1_HVT U2156 ( .A1(n175), .A2(n4124), .A3(n47), .A4(n4111), .Y(n1979) );
  AO22X1_HVT U2157 ( .A1(key_round[100]), .A2(n4525), .A3(n4547), .A4(n1983), 
        .Y(n2225) );
  NAND4X0_HVT U2158 ( .A1(n1984), .A2(n1985), .A3(n1986), .A4(n1987), .Y(n1983) );
  OA222X1_HVT U2159 ( .A1(n1070), .A2(n4240), .A3(n1326), .A4(n4227), .A5(
        n1198), .A6(n4215), .Y(n1987) );
  OA222X1_HVT U2160 ( .A1(n686), .A2(n4202), .A3(n942), .A4(n4189), .A5(n814), 
        .A6(n4176), .Y(n1986) );
  OA222X1_HVT U2161 ( .A1(n302), .A2(n4163), .A3(n558), .A4(n4150), .A5(n430), 
        .A6(n4137), .Y(n1985) );
  OA22X1_HVT U2162 ( .A1(n174), .A2(n4124), .A3(n46), .A4(n4111), .Y(n1984) );
  AO22X1_HVT U2163 ( .A1(key_round[101]), .A2(n4524), .A3(n4547), .A4(n1988), 
        .Y(n2226) );
  NAND4X0_HVT U2164 ( .A1(n1989), .A2(n1990), .A3(n1991), .A4(n1992), .Y(n1988) );
  OA222X1_HVT U2165 ( .A1(n1069), .A2(n4240), .A3(n1325), .A4(n4227), .A5(
        n1197), .A6(n4215), .Y(n1992) );
  OA222X1_HVT U2166 ( .A1(n685), .A2(n4202), .A3(n941), .A4(n4189), .A5(n813), 
        .A6(n4176), .Y(n1991) );
  OA222X1_HVT U2167 ( .A1(n301), .A2(n4163), .A3(n557), .A4(n4150), .A5(n429), 
        .A6(n4137), .Y(n1990) );
  OA22X1_HVT U2168 ( .A1(n173), .A2(n4124), .A3(n45), .A4(n4111), .Y(n1989) );
  AO22X1_HVT U2169 ( .A1(key_round[102]), .A2(n4524), .A3(n4547), .A4(n1993), 
        .Y(n2227) );
  NAND4X0_HVT U2170 ( .A1(n1994), .A2(n1995), .A3(n1996), .A4(n1997), .Y(n1993) );
  OA222X1_HVT U2171 ( .A1(n1068), .A2(n4240), .A3(n1324), .A4(n4227), .A5(
        n1196), .A6(n4215), .Y(n1997) );
  OA222X1_HVT U2172 ( .A1(n684), .A2(n4202), .A3(n940), .A4(n4189), .A5(n812), 
        .A6(n4176), .Y(n1996) );
  OA222X1_HVT U2173 ( .A1(n300), .A2(n4163), .A3(n556), .A4(n4150), .A5(n428), 
        .A6(n4137), .Y(n1995) );
  OA22X1_HVT U2174 ( .A1(n172), .A2(n4124), .A3(n44), .A4(n4111), .Y(n1994) );
  AO22X1_HVT U2175 ( .A1(key_round[103]), .A2(n4524), .A3(n4547), .A4(n1998), 
        .Y(n2228) );
  NAND4X0_HVT U2176 ( .A1(n1999), .A2(n2000), .A3(n2001), .A4(n2002), .Y(n1998) );
  OA222X1_HVT U2177 ( .A1(n1067), .A2(n4240), .A3(n1323), .A4(n4227), .A5(
        n1195), .A6(n4215), .Y(n2002) );
  OA222X1_HVT U2178 ( .A1(n683), .A2(n4202), .A3(n939), .A4(n4189), .A5(n811), 
        .A6(n4176), .Y(n2001) );
  OA222X1_HVT U2179 ( .A1(n299), .A2(n4163), .A3(n555), .A4(n4150), .A5(n427), 
        .A6(n4137), .Y(n2000) );
  OA22X1_HVT U2180 ( .A1(n171), .A2(n4124), .A3(n43), .A4(n4111), .Y(n1999) );
  AO22X1_HVT U2181 ( .A1(key_round[104]), .A2(n4524), .A3(n4547), .A4(n2003), 
        .Y(n2229) );
  NAND4X0_HVT U2182 ( .A1(n2004), .A2(n2005), .A3(n2006), .A4(n2007), .Y(n2003) );
  OA222X1_HVT U2183 ( .A1(n1066), .A2(n4240), .A3(n1322), .A4(n4227), .A5(
        n1194), .A6(n4215), .Y(n2007) );
  OA222X1_HVT U2184 ( .A1(n682), .A2(n4202), .A3(n938), .A4(n4189), .A5(n810), 
        .A6(n4176), .Y(n2006) );
  OA222X1_HVT U2185 ( .A1(n298), .A2(n4163), .A3(n554), .A4(n4150), .A5(n426), 
        .A6(n4137), .Y(n2005) );
  OA22X1_HVT U2186 ( .A1(n170), .A2(n4124), .A3(n42), .A4(n4111), .Y(n2004) );
  AO22X1_HVT U2187 ( .A1(key_round[105]), .A2(n4524), .A3(n4547), .A4(n2008), 
        .Y(n2230) );
  NAND4X0_HVT U2188 ( .A1(n2009), .A2(n2010), .A3(n2011), .A4(n2012), .Y(n2008) );
  OA222X1_HVT U2189 ( .A1(n1065), .A2(n4240), .A3(n1321), .A4(n4227), .A5(
        n1193), .A6(n4215), .Y(n2012) );
  OA222X1_HVT U2190 ( .A1(n681), .A2(n4202), .A3(n937), .A4(n4189), .A5(n809), 
        .A6(n4176), .Y(n2011) );
  OA222X1_HVT U2191 ( .A1(n297), .A2(n4163), .A3(n553), .A4(n4150), .A5(n425), 
        .A6(n4137), .Y(n2010) );
  OA22X1_HVT U2192 ( .A1(n169), .A2(n4124), .A3(n41), .A4(n4111), .Y(n2009) );
  AO22X1_HVT U2193 ( .A1(key_round[106]), .A2(n4524), .A3(n4547), .A4(n2013), 
        .Y(n2231) );
  NAND4X0_HVT U2194 ( .A1(n2014), .A2(n2015), .A3(n2016), .A4(n2017), .Y(n2013) );
  OA222X1_HVT U2195 ( .A1(n1064), .A2(n4240), .A3(n1320), .A4(n4227), .A5(
        n1192), .A6(n4215), .Y(n2017) );
  OA222X1_HVT U2196 ( .A1(n680), .A2(n4202), .A3(n936), .A4(n4189), .A5(n808), 
        .A6(n4176), .Y(n2016) );
  OA222X1_HVT U2197 ( .A1(n296), .A2(n4163), .A3(n552), .A4(n4150), .A5(n424), 
        .A6(n4137), .Y(n2015) );
  OA22X1_HVT U2198 ( .A1(n168), .A2(n4124), .A3(n40), .A4(n4111), .Y(n2014) );
  AO22X1_HVT U2199 ( .A1(key_round[107]), .A2(n4524), .A3(n4547), .A4(n2018), 
        .Y(n2232) );
  NAND4X0_HVT U2200 ( .A1(n2019), .A2(n2020), .A3(n2021), .A4(n2022), .Y(n2018) );
  OA222X1_HVT U2201 ( .A1(n1063), .A2(n4240), .A3(n1319), .A4(n4227), .A5(
        n1191), .A6(n4215), .Y(n2022) );
  OA222X1_HVT U2202 ( .A1(n679), .A2(n4202), .A3(n935), .A4(n4189), .A5(n807), 
        .A6(n4176), .Y(n2021) );
  OA222X1_HVT U2203 ( .A1(n295), .A2(n4163), .A3(n551), .A4(n4150), .A5(n423), 
        .A6(n4137), .Y(n2020) );
  OA22X1_HVT U2204 ( .A1(n167), .A2(n4124), .A3(n39), .A4(n4111), .Y(n2019) );
  AO22X1_HVT U2205 ( .A1(key_round[108]), .A2(n4524), .A3(n4547), .A4(n2023), 
        .Y(n2233) );
  NAND4X0_HVT U2206 ( .A1(n2024), .A2(n2025), .A3(n2026), .A4(n2027), .Y(n2023) );
  OA222X1_HVT U2207 ( .A1(n1062), .A2(n4241), .A3(n1318), .A4(n4227), .A5(
        n1190), .A6(n4216), .Y(n2027) );
  OA222X1_HVT U2208 ( .A1(n678), .A2(n4203), .A3(n934), .A4(n4190), .A5(n806), 
        .A6(n4177), .Y(n2026) );
  OA222X1_HVT U2209 ( .A1(n294), .A2(n4164), .A3(n550), .A4(n4151), .A5(n422), 
        .A6(n4138), .Y(n2025) );
  OA22X1_HVT U2210 ( .A1(n166), .A2(n4125), .A3(n38), .A4(n4112), .Y(n2024) );
  AO22X1_HVT U2211 ( .A1(key_round[109]), .A2(n4524), .A3(n4547), .A4(n2028), 
        .Y(n2234) );
  NAND4X0_HVT U2212 ( .A1(n2029), .A2(n2030), .A3(n2031), .A4(n2032), .Y(n2028) );
  OA222X1_HVT U2213 ( .A1(n1061), .A2(n4241), .A3(n1317), .A4(n4227), .A5(
        n1189), .A6(n4216), .Y(n2032) );
  OA222X1_HVT U2214 ( .A1(n677), .A2(n4203), .A3(n933), .A4(n4190), .A5(n805), 
        .A6(n4177), .Y(n2031) );
  OA222X1_HVT U2215 ( .A1(n293), .A2(n4164), .A3(n549), .A4(n4151), .A5(n421), 
        .A6(n4138), .Y(n2030) );
  OA22X1_HVT U2216 ( .A1(n165), .A2(n4125), .A3(n37), .A4(n4112), .Y(n2029) );
  AO22X1_HVT U2217 ( .A1(key_round[110]), .A2(n4524), .A3(n4547), .A4(n2033), 
        .Y(n2235) );
  NAND4X0_HVT U2218 ( .A1(n2034), .A2(n2035), .A3(n2036), .A4(n2037), .Y(n2033) );
  OA222X1_HVT U2219 ( .A1(n1060), .A2(n4241), .A3(n1316), .A4(n4227), .A5(
        n1188), .A6(n4216), .Y(n2037) );
  OA222X1_HVT U2220 ( .A1(n676), .A2(n4203), .A3(n932), .A4(n4190), .A5(n804), 
        .A6(n4177), .Y(n2036) );
  OA222X1_HVT U2221 ( .A1(n292), .A2(n4164), .A3(n548), .A4(n4151), .A5(n420), 
        .A6(n4138), .Y(n2035) );
  OA22X1_HVT U2222 ( .A1(n164), .A2(n4125), .A3(n36), .A4(n4112), .Y(n2034) );
  AO22X1_HVT U2223 ( .A1(key_round[111]), .A2(n4524), .A3(n4547), .A4(n2038), 
        .Y(n2236) );
  NAND4X0_HVT U2224 ( .A1(n2039), .A2(n2040), .A3(n2041), .A4(n2042), .Y(n2038) );
  OA222X1_HVT U2225 ( .A1(n1059), .A2(n4241), .A3(n1315), .A4(n4227), .A5(
        n1187), .A6(n4216), .Y(n2042) );
  OA222X1_HVT U2226 ( .A1(n675), .A2(n4203), .A3(n931), .A4(n4190), .A5(n803), 
        .A6(n4177), .Y(n2041) );
  OA222X1_HVT U2227 ( .A1(n291), .A2(n4164), .A3(n547), .A4(n4151), .A5(n419), 
        .A6(n4138), .Y(n2040) );
  OA22X1_HVT U2228 ( .A1(n163), .A2(n4125), .A3(n35), .A4(n4112), .Y(n2039) );
  AO22X1_HVT U2229 ( .A1(key_round[112]), .A2(n4524), .A3(n4547), .A4(n2043), 
        .Y(n2237) );
  NAND4X0_HVT U2230 ( .A1(n2044), .A2(n2045), .A3(n2046), .A4(n2047), .Y(n2043) );
  OA222X1_HVT U2231 ( .A1(n1058), .A2(n4241), .A3(n1314), .A4(n4227), .A5(
        n1186), .A6(n4216), .Y(n2047) );
  OA222X1_HVT U2232 ( .A1(n674), .A2(n4203), .A3(n930), .A4(n4190), .A5(n802), 
        .A6(n4177), .Y(n2046) );
  OA222X1_HVT U2233 ( .A1(n290), .A2(n4164), .A3(n546), .A4(n4151), .A5(n418), 
        .A6(n4138), .Y(n2045) );
  OA22X1_HVT U2234 ( .A1(n162), .A2(n4125), .A3(n34), .A4(n4112), .Y(n2044) );
  AO22X1_HVT U2235 ( .A1(key_round[113]), .A2(n4523), .A3(n4547), .A4(n2048), 
        .Y(n2238) );
  NAND4X0_HVT U2236 ( .A1(n2049), .A2(n2050), .A3(n2051), .A4(n2052), .Y(n2048) );
  OA222X1_HVT U2237 ( .A1(n1057), .A2(n4241), .A3(n1313), .A4(n4228), .A5(
        n1185), .A6(n4216), .Y(n2052) );
  OA222X1_HVT U2238 ( .A1(n673), .A2(n4203), .A3(n929), .A4(n4190), .A5(n801), 
        .A6(n4177), .Y(n2051) );
  OA222X1_HVT U2239 ( .A1(n289), .A2(n4164), .A3(n545), .A4(n4151), .A5(n417), 
        .A6(n4138), .Y(n2050) );
  OA22X1_HVT U2240 ( .A1(n161), .A2(n4125), .A3(n33), .A4(n4112), .Y(n2049) );
  AO22X1_HVT U2241 ( .A1(key_round[114]), .A2(n4523), .A3(n4547), .A4(n2053), 
        .Y(n2239) );
  NAND4X0_HVT U2242 ( .A1(n2054), .A2(n2055), .A3(n2056), .A4(n2057), .Y(n2053) );
  OA222X1_HVT U2243 ( .A1(n1056), .A2(n4241), .A3(n1312), .A4(n4228), .A5(
        n1184), .A6(n4216), .Y(n2057) );
  OA222X1_HVT U2244 ( .A1(n672), .A2(n4203), .A3(n928), .A4(n4190), .A5(n800), 
        .A6(n4177), .Y(n2056) );
  OA222X1_HVT U2245 ( .A1(n288), .A2(n4164), .A3(n544), .A4(n4151), .A5(n416), 
        .A6(n4138), .Y(n2055) );
  OA22X1_HVT U2246 ( .A1(n160), .A2(n4125), .A3(n32), .A4(n4112), .Y(n2054) );
  AO22X1_HVT U2247 ( .A1(key_round[115]), .A2(n4523), .A3(n4546), .A4(n2058), 
        .Y(n2240) );
  NAND4X0_HVT U2248 ( .A1(n2059), .A2(n2060), .A3(n2061), .A4(n2062), .Y(n2058) );
  OA222X1_HVT U2249 ( .A1(n1055), .A2(n4241), .A3(n1311), .A4(n4228), .A5(
        n1183), .A6(n4216), .Y(n2062) );
  OA222X1_HVT U2250 ( .A1(n671), .A2(n4203), .A3(n927), .A4(n4190), .A5(n799), 
        .A6(n4177), .Y(n2061) );
  OA222X1_HVT U2251 ( .A1(n287), .A2(n4164), .A3(n543), .A4(n4151), .A5(n415), 
        .A6(n4138), .Y(n2060) );
  OA22X1_HVT U2252 ( .A1(n159), .A2(n4125), .A3(n31), .A4(n4112), .Y(n2059) );
  AO22X1_HVT U2253 ( .A1(key_round[116]), .A2(n4523), .A3(n4546), .A4(n2063), 
        .Y(n2241) );
  NAND4X0_HVT U2254 ( .A1(n2064), .A2(n2065), .A3(n2066), .A4(n2067), .Y(n2063) );
  OA222X1_HVT U2255 ( .A1(n1054), .A2(n4241), .A3(n1310), .A4(n4228), .A5(
        n1182), .A6(n4216), .Y(n2067) );
  OA222X1_HVT U2256 ( .A1(n670), .A2(n4203), .A3(n926), .A4(n4190), .A5(n798), 
        .A6(n4177), .Y(n2066) );
  OA222X1_HVT U2257 ( .A1(n286), .A2(n4164), .A3(n542), .A4(n4151), .A5(n414), 
        .A6(n4138), .Y(n2065) );
  OA22X1_HVT U2258 ( .A1(n158), .A2(n4125), .A3(n30), .A4(n4112), .Y(n2064) );
  AO22X1_HVT U2259 ( .A1(key_round[117]), .A2(n4523), .A3(n4546), .A4(n2068), 
        .Y(n2242) );
  NAND4X0_HVT U2260 ( .A1(n2069), .A2(n2070), .A3(n2071), .A4(n2072), .Y(n2068) );
  OA222X1_HVT U2261 ( .A1(n1053), .A2(n4241), .A3(n1309), .A4(n4228), .A5(
        n1181), .A6(n4216), .Y(n2072) );
  OA222X1_HVT U2262 ( .A1(n669), .A2(n4203), .A3(n925), .A4(n4190), .A5(n797), 
        .A6(n4177), .Y(n2071) );
  OA222X1_HVT U2263 ( .A1(n285), .A2(n4164), .A3(n541), .A4(n4151), .A5(n413), 
        .A6(n4138), .Y(n2070) );
  OA22X1_HVT U2264 ( .A1(n157), .A2(n4125), .A3(n29), .A4(n4112), .Y(n2069) );
  AO22X1_HVT U2265 ( .A1(key_round[118]), .A2(n4523), .A3(n4546), .A4(n2073), 
        .Y(n2243) );
  NAND4X0_HVT U2266 ( .A1(n2074), .A2(n2075), .A3(n2076), .A4(n2077), .Y(n2073) );
  OA222X1_HVT U2267 ( .A1(n1052), .A2(n4241), .A3(n1308), .A4(n4228), .A5(
        n1180), .A6(n4216), .Y(n2077) );
  OA222X1_HVT U2268 ( .A1(n668), .A2(n4203), .A3(n924), .A4(n4190), .A5(n796), 
        .A6(n4177), .Y(n2076) );
  OA222X1_HVT U2269 ( .A1(n284), .A2(n4164), .A3(n540), .A4(n4151), .A5(n412), 
        .A6(n4138), .Y(n2075) );
  OA22X1_HVT U2270 ( .A1(n156), .A2(n4125), .A3(n28), .A4(n4112), .Y(n2074) );
  AO22X1_HVT U2271 ( .A1(key_round[119]), .A2(n4523), .A3(n4546), .A4(n2078), 
        .Y(n2244) );
  NAND4X0_HVT U2272 ( .A1(n2079), .A2(n2080), .A3(n2081), .A4(n2082), .Y(n2078) );
  OA222X1_HVT U2273 ( .A1(n1051), .A2(n4241), .A3(n1307), .A4(n4228), .A5(
        n1179), .A6(n4216), .Y(n2082) );
  OA222X1_HVT U2274 ( .A1(n667), .A2(n4203), .A3(n923), .A4(n4190), .A5(n795), 
        .A6(n4177), .Y(n2081) );
  OA222X1_HVT U2275 ( .A1(n283), .A2(n4164), .A3(n539), .A4(n4151), .A5(n411), 
        .A6(n4138), .Y(n2080) );
  OA22X1_HVT U2276 ( .A1(n155), .A2(n4125), .A3(n27), .A4(n4112), .Y(n2079) );
  AO22X1_HVT U2277 ( .A1(key_round[120]), .A2(n4523), .A3(n4546), .A4(n2083), 
        .Y(n2245) );
  NAND4X0_HVT U2278 ( .A1(n2084), .A2(n2085), .A3(n2086), .A4(n2087), .Y(n2083) );
  OA222X1_HVT U2279 ( .A1(n1050), .A2(n4242), .A3(n1306), .A4(n4228), .A5(
        n1178), .A6(n4217), .Y(n2087) );
  OA222X1_HVT U2280 ( .A1(n666), .A2(n4204), .A3(n922), .A4(n4191), .A5(n794), 
        .A6(n4178), .Y(n2086) );
  OA222X1_HVT U2281 ( .A1(n282), .A2(n4165), .A3(n538), .A4(n4152), .A5(n410), 
        .A6(n4139), .Y(n2085) );
  OA22X1_HVT U2282 ( .A1(n154), .A2(n4126), .A3(n26), .A4(n4113), .Y(n2084) );
  AO22X1_HVT U2283 ( .A1(key_round[121]), .A2(n4523), .A3(n4546), .A4(n2088), 
        .Y(n2246) );
  NAND4X0_HVT U2284 ( .A1(n2089), .A2(n2090), .A3(n2091), .A4(n2092), .Y(n2088) );
  OA222X1_HVT U2285 ( .A1(n1049), .A2(n4242), .A3(n1305), .A4(n4228), .A5(
        n1177), .A6(n4217), .Y(n2092) );
  OA222X1_HVT U2286 ( .A1(n665), .A2(n4204), .A3(n921), .A4(n4191), .A5(n793), 
        .A6(n4178), .Y(n2091) );
  OA222X1_HVT U2287 ( .A1(n281), .A2(n4165), .A3(n537), .A4(n4152), .A5(n409), 
        .A6(n4139), .Y(n2090) );
  OA22X1_HVT U2288 ( .A1(n153), .A2(n4126), .A3(n25), .A4(n4113), .Y(n2089) );
  AO22X1_HVT U2289 ( .A1(key_round[122]), .A2(n4523), .A3(n4546), .A4(n2093), 
        .Y(n2247) );
  NAND4X0_HVT U2290 ( .A1(n2094), .A2(n2095), .A3(n2096), .A4(n2097), .Y(n2093) );
  OA222X1_HVT U2291 ( .A1(n1048), .A2(n4242), .A3(n1304), .A4(n4228), .A5(
        n1176), .A6(n4217), .Y(n2097) );
  OA222X1_HVT U2292 ( .A1(n664), .A2(n4204), .A3(n920), .A4(n4191), .A5(n792), 
        .A6(n4178), .Y(n2096) );
  OA222X1_HVT U2293 ( .A1(n280), .A2(n4165), .A3(n536), .A4(n4152), .A5(n408), 
        .A6(n4139), .Y(n2095) );
  OA22X1_HVT U2294 ( .A1(n152), .A2(n4126), .A3(n24), .A4(n4113), .Y(n2094) );
  AO22X1_HVT U2295 ( .A1(key_round[123]), .A2(n4523), .A3(n4546), .A4(n2098), 
        .Y(n2248) );
  NAND4X0_HVT U2296 ( .A1(n2099), .A2(n2100), .A3(n2101), .A4(n2102), .Y(n2098) );
  OA222X1_HVT U2297 ( .A1(n1047), .A2(n4242), .A3(n1303), .A4(n4228), .A5(
        n1175), .A6(n4217), .Y(n2102) );
  OA222X1_HVT U2298 ( .A1(n663), .A2(n4204), .A3(n919), .A4(n4191), .A5(n791), 
        .A6(n4178), .Y(n2101) );
  OA222X1_HVT U2299 ( .A1(n279), .A2(n4165), .A3(n535), .A4(n4152), .A5(n407), 
        .A6(n4139), .Y(n2100) );
  OA22X1_HVT U2300 ( .A1(n151), .A2(n4126), .A3(n23), .A4(n4113), .Y(n2099) );
  AO22X1_HVT U2301 ( .A1(key_round[124]), .A2(n4523), .A3(n4546), .A4(n2103), 
        .Y(n2249) );
  NAND4X0_HVT U2302 ( .A1(n2104), .A2(n2105), .A3(n2106), .A4(n2107), .Y(n2103) );
  OA222X1_HVT U2303 ( .A1(n1046), .A2(n4242), .A3(n1302), .A4(n4228), .A5(
        n1174), .A6(n4217), .Y(n2107) );
  OA222X1_HVT U2304 ( .A1(n662), .A2(n4204), .A3(n918), .A4(n4191), .A5(n790), 
        .A6(n4178), .Y(n2106) );
  OA222X1_HVT U2305 ( .A1(n278), .A2(n4165), .A3(n534), .A4(n4152), .A5(n406), 
        .A6(n4139), .Y(n2105) );
  OA22X1_HVT U2306 ( .A1(n150), .A2(n4126), .A3(n22), .A4(n4113), .Y(n2104) );
  AO22X1_HVT U2307 ( .A1(key_round[125]), .A2(n4522), .A3(n4546), .A4(n2108), 
        .Y(n2250) );
  NAND4X0_HVT U2308 ( .A1(n2109), .A2(n2110), .A3(n2111), .A4(n2112), .Y(n2108) );
  OA222X1_HVT U2309 ( .A1(n1045), .A2(n4242), .A3(n1301), .A4(n4228), .A5(
        n1173), .A6(n4217), .Y(n2112) );
  OA222X1_HVT U2310 ( .A1(n661), .A2(n4204), .A3(n917), .A4(n4191), .A5(n789), 
        .A6(n4178), .Y(n2111) );
  OA222X1_HVT U2311 ( .A1(n277), .A2(n4165), .A3(n533), .A4(n4152), .A5(n405), 
        .A6(n4139), .Y(n2110) );
  OA22X1_HVT U2312 ( .A1(n149), .A2(n4126), .A3(n21), .A4(n4113), .Y(n2109) );
  AO22X1_HVT U2313 ( .A1(key_round[126]), .A2(n4522), .A3(n4546), .A4(n2113), 
        .Y(n2251) );
  NAND4X0_HVT U2314 ( .A1(n2114), .A2(n2115), .A3(n2116), .A4(n2117), .Y(n2113) );
  OA222X1_HVT U2315 ( .A1(n1044), .A2(n4242), .A3(n1300), .A4(n4229), .A5(
        n1172), .A6(n4217), .Y(n2117) );
  OA222X1_HVT U2316 ( .A1(n660), .A2(n4204), .A3(n916), .A4(n4191), .A5(n788), 
        .A6(n4178), .Y(n2116) );
  OA222X1_HVT U2317 ( .A1(n276), .A2(n4165), .A3(n532), .A4(n4152), .A5(n404), 
        .A6(n4139), .Y(n2115) );
  OA22X1_HVT U2318 ( .A1(n148), .A2(n4126), .A3(n20), .A4(n4113), .Y(n2114) );
  AO22X1_HVT U2319 ( .A1(key_round[127]), .A2(n4522), .A3(n4546), .A4(n2118), 
        .Y(n2252) );
  NAND4X0_HVT U2320 ( .A1(n2119), .A2(n2120), .A3(n2121), .A4(n2122), .Y(n2118) );
  OA222X1_HVT U2321 ( .A1(n1043), .A2(n4242), .A3(n1299), .A4(n4229), .A5(
        n1171), .A6(n4217), .Y(n2122) );
  NAND2X0_HVT U2322 ( .A1(rount_no[0]), .A2(rount_no[3]), .Y(n1479) );
  NAND2X0_HVT U2323 ( .A1(rount_no[3]), .A2(rount_no[1]), .Y(n1478) );
  NAND2X0_HVT U2324 ( .A1(n2123), .A2(rount_no[3]), .Y(n1477) );
  OA222X1_HVT U2325 ( .A1(n659), .A2(n4204), .A3(n915), .A4(n4191), .A5(n787), 
        .A6(n4178), .Y(n2121) );
  NAND3X0_HVT U2326 ( .A1(rount_no[1]), .A2(n4557), .A3(rount_no[2]), .Y(n1482) );
  NAND3X0_HVT U2327 ( .A1(rount_no[0]), .A2(rount_no[1]), .A3(rount_no[2]), 
        .Y(n1481) );
  NAND3X0_HVT U2328 ( .A1(rount_no[0]), .A2(n4558), .A3(rount_no[2]), .Y(n1480) );
  OA222X1_HVT U2329 ( .A1(n275), .A2(n4165), .A3(n531), .A4(n4152), .A5(n403), 
        .A6(n4139), .Y(n2120) );
  OR3X1_HVT U2330 ( .A1(n4558), .A2(rount_no[2]), .A3(n4557), .Y(n1485) );
  NAND2X0_HVT U2331 ( .A1(rount_no[2]), .A2(n2123), .Y(n1484) );
  NAND3X0_HVT U2332 ( .A1(rount_no[1]), .A2(n4557), .A3(n2124), .Y(n1483) );
  OA22X1_HVT U2333 ( .A1(n147), .A2(n4126), .A3(n19), .A4(n4113), .Y(n2119) );
  NAND2X0_HVT U2334 ( .A1(n2124), .A2(n2123), .Y(n1487) );
  AND2X1_HVT U2335 ( .A1(n4557), .A2(n4558), .Y(n2123) );
  NAND3X0_HVT U2336 ( .A1(rount_no[0]), .A2(n4558), .A3(n2124), .Y(n1486) );
  NOR2X0_HVT U2337 ( .A1(rount_no[2]), .A2(rount_no[3]), .Y(n2124) );
  AO22X1_HVT U2338 ( .A1(n3998), .A2(n4540), .A3(\keys[10][0] ), .A4(n4522), 
        .Y(n2253) );
  AO22X1_HVT U2339 ( .A1(n4001), .A2(n4540), .A3(\keys[10][1] ), .A4(n4522), 
        .Y(n2254) );
  AO22X1_HVT U2340 ( .A1(keyout[2]), .A2(n4540), .A3(\keys[10][2] ), .A4(n4522), .Y(n2255) );
  AO22X1_HVT U2341 ( .A1(n4005), .A2(n4540), .A3(\keys[10][3] ), .A4(n4522), 
        .Y(n2256) );
  AO22X1_HVT U2342 ( .A1(n4008), .A2(n4540), .A3(\keys[10][4] ), .A4(n4522), 
        .Y(n2257) );
  AO22X1_HVT U2343 ( .A1(n4011), .A2(n4540), .A3(\keys[10][5] ), .A4(n4522), 
        .Y(n2258) );
  AO22X1_HVT U2344 ( .A1(n4014), .A2(n4540), .A3(\keys[10][6] ), .A4(n4522), 
        .Y(n2259) );
  AO22X1_HVT U2345 ( .A1(keyout[7]), .A2(n4540), .A3(\keys[10][7] ), .A4(n4521), .Y(n2260) );
  AO22X1_HVT U2346 ( .A1(n4018), .A2(n4540), .A3(\keys[10][8] ), .A4(n4521), 
        .Y(n2261) );
  AO22X1_HVT U2347 ( .A1(n4021), .A2(n4540), .A3(\keys[10][9] ), .A4(n4521), 
        .Y(n2262) );
  AO22X1_HVT U2348 ( .A1(n4024), .A2(n4539), .A3(\keys[10][10] ), .A4(n4521), 
        .Y(n2263) );
  AO22X1_HVT U2349 ( .A1(n4027), .A2(n4539), .A3(\keys[10][11] ), .A4(n4521), 
        .Y(n2264) );
  AO22X1_HVT U2350 ( .A1(n4030), .A2(n4539), .A3(\keys[10][12] ), .A4(n4521), 
        .Y(n2265) );
  AO22X1_HVT U2351 ( .A1(n4033), .A2(n4543), .A3(\keys[10][13] ), .A4(n4521), 
        .Y(n2266) );
  AO22X1_HVT U2352 ( .A1(n4036), .A2(n4539), .A3(\keys[10][14] ), .A4(n4521), 
        .Y(n2267) );
  AO22X1_HVT U2353 ( .A1(n4039), .A2(n4539), .A3(\keys[10][15] ), .A4(n4521), 
        .Y(n2268) );
  AO22X1_HVT U2354 ( .A1(n4042), .A2(n4539), .A3(\keys[10][16] ), .A4(n4521), 
        .Y(n2269) );
  AO22X1_HVT U2355 ( .A1(n4045), .A2(n4539), .A3(\keys[10][17] ), .A4(n4521), 
        .Y(n2270) );
  AO22X1_HVT U2356 ( .A1(n4048), .A2(n4539), .A3(\keys[10][18] ), .A4(n4521), 
        .Y(n2271) );
  AO22X1_HVT U2357 ( .A1(n4051), .A2(n4539), .A3(\keys[10][19] ), .A4(n4520), 
        .Y(n2272) );
  AO22X1_HVT U2358 ( .A1(n4054), .A2(n4539), .A3(\keys[10][20] ), .A4(n4520), 
        .Y(n2273) );
  AO22X1_HVT U2359 ( .A1(n4057), .A2(n4539), .A3(\keys[10][21] ), .A4(n4520), 
        .Y(n2274) );
  AO22X1_HVT U2360 ( .A1(n4060), .A2(n4539), .A3(\keys[10][22] ), .A4(n4520), 
        .Y(n2275) );
  AO22X1_HVT U2361 ( .A1(n4063), .A2(n4539), .A3(\keys[10][23] ), .A4(n4520), 
        .Y(n2276) );
  AO22X1_HVT U2362 ( .A1(n4066), .A2(n4539), .A3(\keys[10][24] ), .A4(n4520), 
        .Y(n2277) );
  AO22X1_HVT U2363 ( .A1(n4068), .A2(n4538), .A3(\keys[10][25] ), .A4(n4520), 
        .Y(n2278) );
  AO22X1_HVT U2364 ( .A1(n4071), .A2(n4538), .A3(\keys[10][26] ), .A4(n4520), 
        .Y(n2279) );
  AO22X1_HVT U2365 ( .A1(n4074), .A2(n4538), .A3(\keys[10][27] ), .A4(n4520), 
        .Y(n2280) );
  AO22X1_HVT U2366 ( .A1(n4077), .A2(n4538), .A3(\keys[10][28] ), .A4(n4520), 
        .Y(n2281) );
  AO22X1_HVT U2367 ( .A1(n4080), .A2(n4538), .A3(\keys[10][29] ), .A4(n4520), 
        .Y(n2282) );
  AO22X1_HVT U2368 ( .A1(keyout[30]), .A2(n4538), .A3(\keys[10][30] ), .A4(
        n4520), .Y(n2283) );
  AO22X1_HVT U2369 ( .A1(n3852), .A2(n4538), .A3(\keys[10][31] ), .A4(n4519), 
        .Y(n2284) );
  AO22X1_HVT U2370 ( .A1(keyout[32]), .A2(n4538), .A3(\keys[10][32] ), .A4(
        n4519), .Y(n2285) );
  AO22X1_HVT U2371 ( .A1(n3876), .A2(n4538), .A3(\keys[10][33] ), .A4(n4519), 
        .Y(n2286) );
  AO22X1_HVT U2372 ( .A1(n3913), .A2(n4538), .A3(\keys[10][34] ), .A4(n4519), 
        .Y(n2287) );
  AO22X1_HVT U2373 ( .A1(keyout[35]), .A2(n4538), .A3(\keys[10][35] ), .A4(
        n4519), .Y(n2288) );
  AO22X1_HVT U2374 ( .A1(keyout[36]), .A2(n4538), .A3(\keys[10][36] ), .A4(
        n4519), .Y(n2289) );
  AO22X1_HVT U2375 ( .A1(n3911), .A2(n4538), .A3(\keys[10][37] ), .A4(n4519), 
        .Y(n2290) );
  AO22X1_HVT U2376 ( .A1(keyout[38]), .A2(n4538), .A3(\keys[10][38] ), .A4(
        n4519), .Y(n2291) );
  AO22X1_HVT U2377 ( .A1(keyout[39]), .A2(n4538), .A3(\keys[10][39] ), .A4(
        n4519), .Y(n2292) );
  AO22X1_HVT U2378 ( .A1(n3952), .A2(n4537), .A3(\keys[10][40] ), .A4(n4519), 
        .Y(n2293) );
  AO22X1_HVT U2379 ( .A1(n3884), .A2(n4537), .A3(\keys[10][41] ), .A4(n4519), 
        .Y(n2294) );
  AO22X1_HVT U2380 ( .A1(n3973), .A2(n4537), .A3(\keys[10][42] ), .A4(n4519), 
        .Y(n2295) );
  AO22X1_HVT U2381 ( .A1(n3890), .A2(n4537), .A3(\keys[10][43] ), .A4(n4518), 
        .Y(n2296) );
  AO22X1_HVT U2382 ( .A1(n3902), .A2(n4537), .A3(\keys[10][44] ), .A4(n4518), 
        .Y(n2297) );
  AO22X1_HVT U2383 ( .A1(n3935), .A2(n4536), .A3(\keys[10][45] ), .A4(n4518), 
        .Y(n2298) );
  AO22X1_HVT U2384 ( .A1(n3813), .A2(n4535), .A3(\keys[10][46] ), .A4(n4522), 
        .Y(n2299) );
  AO22X1_HVT U2385 ( .A1(n3850), .A2(n4539), .A3(\keys[10][47] ), .A4(n4512), 
        .Y(n2300) );
  NAND4X0_HVT U2386 ( .A1(state[1]), .A2(state[0]), .A3(n1468), .A4(n4559), 
        .Y(n1430) );
  AND2X1_HVT U2387 ( .A1(state[3]), .A2(n16), .Y(n1468) );
  keygen_1 key ( .round_num(round_number), .keyin({prev_key[127:24], n3822, 
        prev_key[22:19], n3933, n9, prev_key[16], n7, prev_key[14:11], n3918, 
        prev_key[9:8], n3900, prev_key[6:3], n3848, prev_key[1:0]}), .keyout(
        keyout) );
  NBUFFX2_HVT U3 ( .A(keyout[85]), .Y(n1) );
  NBUFFX2_HVT U4 ( .A(keyout[85]), .Y(n2) );
  NBUFFX4_HVT U5 ( .A(keyout[78]), .Y(n3947) );
  OAI22X1_HVT U6 ( .A1(n4374), .A2(n3978), .A3(n584), .A4(n4385), .Y(n3095) );
  INVX0_HVT U7 ( .A(n3978), .Y(n3979) );
  INVX2_HVT U8 ( .A(keyout[74]), .Y(n3978) );
  INVX2_HVT U9 ( .A(n6), .Y(n7) );
  INVX1_HVT U10 ( .A(n3936), .Y(n3) );
  INVX1_HVT U11 ( .A(n3815), .Y(n4) );
  OAI22X1_HVT U12 ( .A1(n4352), .A2(n3815), .A3(n439), .A4(n5), .Y(n3240) );
  IBUFFX16_HVT U13 ( .A(n4355), .Y(n5) );
  INVX1_HVT U14 ( .A(n8), .Y(n9) );
  INVX1_HVT U15 ( .A(n3940), .Y(n10) );
  OAI22X1_HVT U16 ( .A1(n4533), .A2(n3948), .A3(n1336), .A4(n4554), .Y(n2343)
         );
  INVX0_HVT U17 ( .A(n4534), .Y(n4533) );
  INVX0_HVT U18 ( .A(n4537), .Y(n4515) );
  INVX0_HVT U19 ( .A(keyout[54]), .Y(n12) );
  INVX0_HVT U62 ( .A(n12), .Y(n13) );
  INVX1_HVT U429 ( .A(n1428), .Y(n14) );
  INVX0_HVT U430 ( .A(keyout[48]), .Y(n15) );
  INVX1_HVT U435 ( .A(n15), .Y(n1427) );
  INVX0_HVT U592 ( .A(keyout[49]), .Y(n1428) );
  INVX0_HVT U667 ( .A(n1428), .Y(n1429) );
  INVX0_HVT U784 ( .A(keyout[50]), .Y(n1431) );
  INVX1_HVT U814 ( .A(n1431), .Y(n1432) );
  INVX0_HVT U815 ( .A(keyout[52]), .Y(n1433) );
  INVX0_HVT U958 ( .A(n1433), .Y(n1434) );
  INVX0_HVT U959 ( .A(keyout[86]), .Y(n1435) );
  INVX1_HVT U1037 ( .A(n1435), .Y(n1436) );
  INVX0_HVT U1041 ( .A(keyout[84]), .Y(n1437) );
  INVX1_HVT U1043 ( .A(n1437), .Y(n1438) );
  NBUFFX2_HVT U1166 ( .A(keyout[28]), .Y(n4076) );
  NBUFFX2_HVT U1167 ( .A(keyout[29]), .Y(n4081) );
  NBUFFX2_HVT U1383 ( .A(keyout[87]), .Y(n1439) );
  NBUFFX2_HVT U1420 ( .A(keyout[87]), .Y(n1440) );
  OAI222X1_HVT U1424 ( .A1(n3798), .A2(n3799), .A3(n4271), .A4(n3800), .A5(
        n3801), .A6(n4256), .Y(n3701) );
  IBUFFX16_HVT U1427 ( .A(n4275), .Y(n3798) );
  IBUFFX16_HVT U1430 ( .A(local_key[87]), .Y(n3799) );
  IBUFFX16_HVT U1431 ( .A(keyout[87]), .Y(n3800) );
  INVX0_HVT U1432 ( .A(keyout[122]), .Y(n3802) );
  INVX1_HVT U1444 ( .A(n3802), .Y(n3803) );
  INVX0_HVT U1446 ( .A(keyout[61]), .Y(n3804) );
  INVX1_HVT U1465 ( .A(n3804), .Y(n3805) );
  OAI222X1_HVT U1470 ( .A1(n4282), .A2(n3806), .A3(n4270), .A4(n3804), .A5(
        n3807), .A6(n4257), .Y(n3727) );
  IBUFFX16_HVT U1522 ( .A(local_key[61]), .Y(n3806) );
  IBUFFX2_HVT U1525 ( .A(n4282), .Y(n4277) );
  INVX1_HVT U1526 ( .A(keyout[123]), .Y(n3808) );
  INVX1_HVT U1529 ( .A(n3808), .Y(n3809) );
  INVX0_HVT U1530 ( .A(keyout[81]), .Y(n3810) );
  INVX1_HVT U1532 ( .A(n3810), .Y(n3811) );
  INVX1_HVT U1533 ( .A(keyout[46]), .Y(n3812) );
  INVX1_HVT U1550 ( .A(n3812), .Y(n3813) );
  OAI22X1_HVT U1552 ( .A1(n4352), .A2(n3948), .A3(n440), .A4(n3814), .Y(n3239)
         );
  IBUFFX16_HVT U1554 ( .A(n4356), .Y(n3814) );
  NBUFFX2_HVT U2388 ( .A(keyout[26]), .Y(n4070) );
  INVX1_HVT U2389 ( .A(keyout[91]), .Y(n3815) );
  INVX1_HVT U2390 ( .A(n3815), .Y(n3816) );
  NBUFFX2_HVT U2391 ( .A(keyout[123]), .Y(n3817) );
  INVX1_HVT U2392 ( .A(n3847), .Y(n3848) );
  INVX1_HVT U2393 ( .A(n3899), .Y(n3900) );
  NBUFFX2_HVT U2394 ( .A(keyout[57]), .Y(n4084) );
  NBUFFX2_HVT U2395 ( .A(keyout[58]), .Y(n4086) );
  INVX1_HVT U2396 ( .A(n1441), .Y(n4282) );
  AND2X1_HVT U2397 ( .A1(n3957), .A2(n3955), .Y(n3818) );
  NBUFFX2_HVT U2398 ( .A(keyout[37]), .Y(n3819) );
  NAND2X0_HVT U2399 ( .A1(n3818), .A2(n3956), .Y(n3713) );
  INVX1_HVT U2400 ( .A(n3821), .Y(n3822) );
  NBUFFX2_HVT U2401 ( .A(keyout[107]), .Y(n3820) );
  NBUFFX2_HVT U2402 ( .A(keyout[125]), .Y(n3823) );
  INVX1_HVT U2403 ( .A(keyout[67]), .Y(n3824) );
  INVX1_HVT U2404 ( .A(n3824), .Y(n3825) );
  INVX1_HVT U2405 ( .A(keyout[89]), .Y(n3826) );
  INVX1_HVT U2406 ( .A(n3826), .Y(n3827) );
  INVX1_HVT U2407 ( .A(keyout[121]), .Y(n3828) );
  INVX1_HVT U2408 ( .A(n3828), .Y(n3829) );
  INVX1_HVT U2409 ( .A(keyout[92]), .Y(n3830) );
  INVX1_HVT U2410 ( .A(n3830), .Y(n3831) );
  NBUFFX2_HVT U2411 ( .A(keyout[62]), .Y(n3832) );
  NBUFFX2_HVT U2412 ( .A(keyout[62]), .Y(n3833) );
  INVX0_HVT U2413 ( .A(n3868), .Y(n3834) );
  INVX1_HVT U2414 ( .A(n3864), .Y(n3835) );
  NAND2X0_HVT U2415 ( .A1(n4323), .A2(n3973), .Y(n3836) );
  NAND2X0_HVT U2416 ( .A1(\keys[1][42] ), .A2(n4311), .Y(n3837) );
  NAND2X0_HVT U2417 ( .A1(n3836), .A2(n3837), .Y(n3447) );
  INVX1_HVT U2418 ( .A(n4306), .Y(n4323) );
  INVX0_HVT U2419 ( .A(keyout[104]), .Y(n3838) );
  INVX0_HVT U2420 ( .A(n3838), .Y(n3839) );
  NAND2X0_HVT U2421 ( .A1(n4272), .A2(local_key[124]), .Y(n3840) );
  NAND2X0_HVT U2422 ( .A1(n4259), .A2(n3844), .Y(n3841) );
  NAND2X0_HVT U2423 ( .A1(prev_key[124]), .A2(n4245), .Y(n3842) );
  NAND3X0_HVT U2424 ( .A1(n3840), .A2(n3841), .A3(n3842), .Y(n3664) );
  INVX1_HVT U2425 ( .A(keyout[124]), .Y(n3843) );
  INVX0_HVT U2426 ( .A(n3843), .Y(n3844) );
  INVX0_HVT U2427 ( .A(n3843), .Y(n3845) );
  INVX0_HVT U2428 ( .A(n3843), .Y(n3846) );
  INVX1_HVT U2429 ( .A(keyout[47]), .Y(n3849) );
  INVX1_HVT U2430 ( .A(n3849), .Y(n3850) );
  INVX1_HVT U2431 ( .A(keyout[31]), .Y(n3851) );
  INVX1_HVT U2432 ( .A(n3851), .Y(n3852) );
  INVX1_HVT U2433 ( .A(keyout[41]), .Y(n3853) );
  INVX1_HVT U2434 ( .A(n3853), .Y(n3854) );
  INVX1_HVT U2435 ( .A(n3917), .Y(n3918) );
  NAND2X0_HVT U2436 ( .A1(n4277), .A2(local_key[63]), .Y(n3855) );
  NAND2X0_HVT U2437 ( .A1(n4264), .A2(n3859), .Y(n3856) );
  NAND2X0_HVT U2438 ( .A1(prev_key[63]), .A2(n4250), .Y(n3857) );
  NAND3X0_HVT U2439 ( .A1(n3855), .A2(n3856), .A3(n3857), .Y(n3725) );
  INVX1_HVT U2440 ( .A(keyout[63]), .Y(n3858) );
  INVX0_HVT U2441 ( .A(n3858), .Y(n3859) );
  INVX0_HVT U2442 ( .A(n3858), .Y(n3860) );
  INVX0_HVT U2443 ( .A(n3858), .Y(n3861) );
  INVX1_HVT U2444 ( .A(keyout[55]), .Y(n3921) );
  INVX1_HVT U2445 ( .A(keyout[43]), .Y(n3889) );
  INVX1_HVT U2446 ( .A(keyout[73]), .Y(n3895) );
  INVX1_HVT U2447 ( .A(keyout[79]), .Y(n3897) );
  INVX0_HVT U2448 ( .A(n3993), .Y(n4374) );
  INVX1_HVT U2449 ( .A(keyout[106]), .Y(n3879) );
  INVX1_HVT U2450 ( .A(n4257), .Y(n4252) );
  INVX1_HVT U2451 ( .A(n4282), .Y(n4279) );
  INVX0_HVT U2452 ( .A(n4401), .Y(n3867) );
  NAND2X0_HVT U2453 ( .A1(n4275), .A2(local_key[83]), .Y(n3923) );
  INVX1_HVT U2454 ( .A(keyout[47]), .Y(n3894) );
  INVX1_HVT U2455 ( .A(keyout[41]), .Y(n3893) );
  INVX1_HVT U2456 ( .A(keyout[72]), .Y(n3950) );
  AND2X1_HVT U2457 ( .A1(n3968), .A2(n3970), .Y(n3862) );
  INVX1_HVT U2458 ( .A(n3826), .Y(n3863) );
  INVX1_HVT U2459 ( .A(keyout[94]), .Y(n3864) );
  INVX1_HVT U2460 ( .A(n3864), .Y(n3865) );
  INVX1_HVT U2461 ( .A(n3921), .Y(n3866) );
  OAI22X1_HVT U2462 ( .A1(n4395), .A2(n3921), .A3(n731), .A4(n3867), .Y(n2948)
         );
  IBUFFX2_HVT U2463 ( .A(n4395), .Y(n4413) );
  INVX1_HVT U2464 ( .A(keyout[95]), .Y(n3868) );
  INVX1_HVT U2465 ( .A(n3868), .Y(n3869) );
  INVX1_HVT U2466 ( .A(keyout[45]), .Y(n3934) );
  NBUFFX2_HVT U2467 ( .A(keyout[65]), .Y(n3870) );
  OAI22X1_HVT U2468 ( .A1(n4374), .A2(n3958), .A3(n583), .A4(n4394), .Y(n3096)
         );
  INVX1_HVT U2469 ( .A(n3934), .Y(n3871) );
  OAI22X1_HVT U2470 ( .A1(n4329), .A2(n3934), .A3(n357), .A4(n4341), .Y(n3322)
         );
  INVX0_HVT U2471 ( .A(n4341), .Y(n4337) );
  INVX1_HVT U2472 ( .A(n3978), .Y(n3872) );
  OAI22X1_HVT U2473 ( .A1(n4441), .A2(n3978), .A3(n968), .A4(n4461), .Y(n2711)
         );
  NBUFFX2_HVT U2474 ( .A(keyout[109]), .Y(n3873) );
  INVX1_HVT U2475 ( .A(n3919), .Y(n3874) );
  INVX1_HVT U2476 ( .A(keyout[33]), .Y(n3875) );
  INVX1_HVT U2477 ( .A(n3875), .Y(n3876) );
  AO22X1_HVT U2478 ( .A1(n4394), .A2(n3888), .A3(n3877), .A4(n4381), .Y(n3065)
         );
  INVX1_HVT U2479 ( .A(keyout[44]), .Y(n3901) );
  INVX0_HVT U2480 ( .A(n3901), .Y(n3888) );
  INVX1_HVT U2481 ( .A(n3889), .Y(n3878) );
  OAI22X1_HVT U2482 ( .A1(n4306), .A2(n3889), .A3(n231), .A4(n4328), .Y(n3448)
         );
  INVX1_HVT U2483 ( .A(n3879), .Y(n3880) );
  INVX1_HVT U2484 ( .A(n3891), .Y(n3881) );
  INVX1_HVT U2485 ( .A(keyout[108]), .Y(n3882) );
  INVX0_HVT U2486 ( .A(keyout[108]), .Y(n3891) );
  INVX1_HVT U2487 ( .A(keyout[37]), .Y(n3909) );
  OAI22X1_HVT U2488 ( .A1(n4429), .A2(n3891), .A3(n806), .A4(n4439), .Y(n2873)
         );
  IBUFFX2_HVT U2489 ( .A(n4419), .Y(n4438) );
  IBUFFX2_HVT U2490 ( .A(n4431), .Y(n4421) );
  NBUFFX2_HVT U2491 ( .A(keyout[65]), .Y(n3883) );
  INVX1_HVT U2492 ( .A(n3893), .Y(n3884) );
  OAI22X1_HVT U2493 ( .A1(n4329), .A2(n3893), .A3(n361), .A4(n4341), .Y(n3318)
         );
  INVX1_HVT U2494 ( .A(n3894), .Y(n3885) );
  OAI22X1_HVT U2495 ( .A1(n4329), .A2(n3894), .A3(n355), .A4(n4350), .Y(n3324)
         );
  IBUFFX2_HVT U2496 ( .A(n4329), .Y(n4345) );
  INVX1_HVT U2497 ( .A(n3895), .Y(n3886) );
  OAI22X1_HVT U2498 ( .A1(n4441), .A2(n3895), .A3(n969), .A4(n4461), .Y(n2710)
         );
  INVX1_HVT U2499 ( .A(n3897), .Y(n3887) );
  OAI22X1_HVT U2500 ( .A1(n4441), .A2(n3897), .A3(n963), .A4(n4461), .Y(n2716)
         );
  IBUFFX2_HVT U2501 ( .A(n4441), .Y(n4458) );
  IBUFFX2_HVT U2502 ( .A(n4373), .Y(n4389) );
  INVX1_HVT U2503 ( .A(n3889), .Y(n3890) );
  INVX1_HVT U2504 ( .A(n3882), .Y(n3892) );
  INVX1_HVT U2505 ( .A(n3895), .Y(n3896) );
  INVX1_HVT U2506 ( .A(n3897), .Y(n3898) );
  INVX1_HVT U2507 ( .A(keyout[42]), .Y(n3971) );
  INVX1_HVT U2508 ( .A(n3901), .Y(n3902) );
  INVX1_HVT U2509 ( .A(keyout[83]), .Y(n3903) );
  INVX1_HVT U2510 ( .A(n3903), .Y(n3904) );
  INVX0_HVT U2511 ( .A(n3976), .Y(n3905) );
  NAND2X1_HVT U2512 ( .A1(n4279), .A2(local_key[37]), .Y(n3906) );
  NAND2X0_HVT U2513 ( .A1(n4266), .A2(n3910), .Y(n3907) );
  NAND2X0_HVT U2514 ( .A1(prev_key[37]), .A2(n4252), .Y(n3908) );
  NAND3X0_HVT U2515 ( .A1(n3906), .A2(n3907), .A3(n3908), .Y(n3751) );
  INVX1_HVT U2516 ( .A(n3909), .Y(n3910) );
  INVX0_HVT U2517 ( .A(n3909), .Y(n3911) );
  INVX1_HVT U2518 ( .A(keyout[34]), .Y(n3912) );
  INVX1_HVT U2519 ( .A(n3912), .Y(n3913) );
  NBUFFX2_HVT U2520 ( .A(keyout[66]), .Y(n3914) );
  NBUFFX2_HVT U2521 ( .A(keyout[115]), .Y(n3915) );
  INVX1_HVT U2522 ( .A(n3926), .Y(n3916) );
  INVX1_HVT U2523 ( .A(keyout[83]), .Y(n3926) );
  INVX1_HVT U2524 ( .A(keyout[53]), .Y(n3919) );
  INVX1_HVT U2525 ( .A(n3919), .Y(n3920) );
  INVX1_HVT U2526 ( .A(n3921), .Y(n3922) );
  NAND2X0_HVT U2527 ( .A1(n4262), .A2(keyout[83]), .Y(n3924) );
  NAND2X0_HVT U2528 ( .A1(prev_key[83]), .A2(n4248), .Y(n3925) );
  NAND3X0_HVT U2529 ( .A1(n3923), .A2(n3924), .A3(n3925), .Y(n3705) );
  INVX1_HVT U2530 ( .A(n3926), .Y(n3927) );
  INVX0_HVT U2531 ( .A(n4256), .Y(n4248) );
  NAND2X0_HVT U2532 ( .A1(n4275), .A2(local_key[80]), .Y(n3928) );
  NAND2X0_HVT U2533 ( .A1(n4262), .A2(keyout[80]), .Y(n3929) );
  NAND2X0_HVT U2534 ( .A1(prev_key[80]), .A2(n4248), .Y(n3930) );
  NAND3X0_HVT U2535 ( .A1(n3928), .A2(n3929), .A3(n3930), .Y(n3708) );
  NBUFFX2_HVT U2536 ( .A(keyout[80]), .Y(n3931) );
  INVX1_HVT U2537 ( .A(n3932), .Y(n3933) );
  INVX1_HVT U2538 ( .A(n3934), .Y(n3935) );
  INVX1_HVT U2539 ( .A(keyout[51]), .Y(n3936) );
  INVX1_HVT U2540 ( .A(n3936), .Y(n3937) );
  INVX1_HVT U2541 ( .A(n3824), .Y(n3938) );
  INVX1_HVT U2542 ( .A(n3950), .Y(n3939) );
  INVX1_HVT U2543 ( .A(keyout[56]), .Y(n3940) );
  INVX1_HVT U2544 ( .A(n3940), .Y(n3941) );
  INVX1_HVT U2545 ( .A(keyout[60]), .Y(n3942) );
  INVX1_HVT U2546 ( .A(n3942), .Y(n3943) );
  NAND2X0_HVT U2547 ( .A1(n3862), .A2(n3969), .Y(n3746) );
  NAND2X0_HVT U2548 ( .A1(n4279), .A2(local_key[42]), .Y(n3968) );
  INVX1_HVT U2549 ( .A(n3971), .Y(n3973) );
  NBUFFX2_HVT U2550 ( .A(keyout[46]), .Y(n3944) );
  NBUFFX2_HVT U2551 ( .A(keyout[46]), .Y(n3945) );
  NBUFFX2_HVT U2552 ( .A(keyout[78]), .Y(n3946) );
  INVX0_HVT U2553 ( .A(n3971), .Y(n3974) );
  INVX1_HVT U2554 ( .A(keyout[90]), .Y(n3948) );
  INVX1_HVT U2555 ( .A(n3948), .Y(n3949) );
  INVX1_HVT U2556 ( .A(n3950), .Y(n3951) );
  NBUFFX2_HVT U2557 ( .A(keyout[40]), .Y(n3952) );
  NBUFFX2_HVT U2558 ( .A(keyout[40]), .Y(n3953) );
  NAND2X0_HVT U2559 ( .A1(n4276), .A2(local_key[75]), .Y(n3955) );
  NAND2X0_HVT U2560 ( .A1(n4263), .A2(keyout[75]), .Y(n3956) );
  NAND2X0_HVT U2561 ( .A1(prev_key[75]), .A2(n4249), .Y(n3957) );
  INVX1_HVT U2562 ( .A(keyout[75]), .Y(n3958) );
  INVX0_HVT U2563 ( .A(n3958), .Y(n3959) );
  INVX0_HVT U2564 ( .A(n3958), .Y(n3960) );
  NAND2X0_HVT U2565 ( .A1(n4276), .A2(local_key[76]), .Y(n3961) );
  NAND2X0_HVT U2566 ( .A1(n4263), .A2(n3965), .Y(n3962) );
  NAND2X0_HVT U2567 ( .A1(prev_key[76]), .A2(n4249), .Y(n3963) );
  NAND3X0_HVT U2568 ( .A1(n3961), .A2(n3962), .A3(n3963), .Y(n3712) );
  INVX1_HVT U2569 ( .A(keyout[76]), .Y(n3964) );
  INVX0_HVT U2570 ( .A(n3964), .Y(n3965) );
  INVX0_HVT U2571 ( .A(n3964), .Y(n3966) );
  INVX0_HVT U2572 ( .A(n3964), .Y(n3967) );
  NAND2X0_HVT U2573 ( .A1(n4266), .A2(n3972), .Y(n3969) );
  NAND2X0_HVT U2574 ( .A1(prev_key[42]), .A2(n4252), .Y(n3970) );
  INVX1_HVT U2575 ( .A(n3971), .Y(n3972) );
  INVX1_HVT U2576 ( .A(keyout[82]), .Y(n3976) );
  INVX1_HVT U2577 ( .A(n3976), .Y(n3977) );
  NAND2X0_HVT U2578 ( .A1(n4276), .A2(local_key[77]), .Y(n3980) );
  NAND2X0_HVT U2579 ( .A1(n4263), .A2(n3984), .Y(n3981) );
  NAND2X0_HVT U2580 ( .A1(prev_key[77]), .A2(n4249), .Y(n3982) );
  NAND3X0_HVT U2581 ( .A1(n3980), .A2(n3981), .A3(n3982), .Y(n3711) );
  INVX1_HVT U2582 ( .A(keyout[77]), .Y(n3983) );
  INVX0_HVT U2583 ( .A(n3983), .Y(n3984) );
  INVX0_HVT U2584 ( .A(n3983), .Y(n3985) );
  INVX0_HVT U2585 ( .A(n3983), .Y(n3986) );
  INVX0_HVT U2586 ( .A(n4507), .Y(n4537) );
  INVX0_HVT U2587 ( .A(n4507), .Y(n4536) );
  INVX0_HVT U2588 ( .A(n4270), .Y(n4269) );
  INVX0_HVT U2589 ( .A(n4091), .Y(n4093) );
  INVX0_HVT U2590 ( .A(n4097), .Y(n4099) );
  INVX0_HVT U2591 ( .A(n4100), .Y(n4102) );
  INVX0_HVT U2592 ( .A(n4094), .Y(n4096) );
  INVX1_HVT U2593 ( .A(n1443), .Y(n4256) );
  INVX0_HVT U2594 ( .A(n1443), .Y(n4257) );
  INVX0_HVT U2595 ( .A(n4140), .Y(n4139) );
  INVX1_HVT U2596 ( .A(n1442), .Y(n4270) );
  INVX0_HVT U2597 ( .A(n3988), .Y(n4330) );
  INVX1_HVT U2598 ( .A(n1485), .Y(n4140) );
  INVX0_HVT U2599 ( .A(n3995), .Y(n4441) );
  INVX0_HVT U2600 ( .A(n3994), .Y(n4463) );
  INVX0_HVT U2601 ( .A(n3996), .Y(n4419) );
  INVX0_HVT U2602 ( .A(n3992), .Y(n4352) );
  INVX0_HVT U2603 ( .A(n4511), .Y(n4510) );
  INVX1_HVT U2604 ( .A(n4319), .Y(n4313) );
  INVX1_HVT U2605 ( .A(n4319), .Y(n4314) );
  INVX1_HVT U2606 ( .A(n4319), .Y(n4315) );
  INVX1_HVT U2607 ( .A(n4319), .Y(n4316) );
  INVX1_HVT U2608 ( .A(n4319), .Y(n4317) );
  INVX1_HVT U2609 ( .A(n4270), .Y(n4264) );
  INVX1_HVT U2610 ( .A(n4270), .Y(n4267) );
  INVX1_HVT U2611 ( .A(n4270), .Y(n4265) );
  INVX1_HVT U2612 ( .A(n4270), .Y(n4266) );
  INVX1_HVT U2613 ( .A(n4271), .Y(n4259) );
  INVX1_HVT U2614 ( .A(n4271), .Y(n4261) );
  INVX1_HVT U2615 ( .A(n4271), .Y(n4262) );
  INVX1_HVT U2616 ( .A(n4271), .Y(n4260) );
  INVX1_HVT U2617 ( .A(n4270), .Y(n4268) );
  INVX1_HVT U2618 ( .A(n4271), .Y(n4263) );
  INVX1_HVT U2619 ( .A(n4296), .Y(n4285) );
  INVX1_HVT U2620 ( .A(n4342), .Y(n4334) );
  INVX1_HVT U2621 ( .A(n4342), .Y(n4333) );
  INVX1_HVT U2622 ( .A(n4342), .Y(n4332) );
  INVX1_HVT U2623 ( .A(n4342), .Y(n4331) );
  INVX1_HVT U2624 ( .A(n4319), .Y(n4318) );
  INVX1_HVT U2625 ( .A(n4296), .Y(n4288) );
  INVX1_HVT U2626 ( .A(n4296), .Y(n4287) );
  INVX1_HVT U2627 ( .A(n4296), .Y(n4286) );
  INVX1_HVT U2628 ( .A(n4295), .Y(n4293) );
  INVX1_HVT U2629 ( .A(n4295), .Y(n4292) );
  INVX1_HVT U2630 ( .A(n4295), .Y(n4291) );
  INVX1_HVT U2631 ( .A(n4295), .Y(n4290) );
  INVX1_HVT U2632 ( .A(n4295), .Y(n4289) );
  INVX1_HVT U2633 ( .A(n4320), .Y(n4310) );
  INVX1_HVT U2634 ( .A(n4320), .Y(n4311) );
  INVX1_HVT U2635 ( .A(n4320), .Y(n4312) );
  INVX1_HVT U2636 ( .A(n4320), .Y(n4308) );
  INVX1_HVT U2637 ( .A(n4320), .Y(n4309) );
  INVX1_HVT U2638 ( .A(n4295), .Y(n4294) );
  INVX1_HVT U2639 ( .A(n4341), .Y(n4338) );
  INVX1_HVT U2640 ( .A(n4341), .Y(n4336) );
  INVX1_HVT U2641 ( .A(n4341), .Y(n4335) );
  INVX1_HVT U2642 ( .A(n4341), .Y(n4339) );
  INVX1_HVT U2643 ( .A(n4341), .Y(n4340) );
  INVX1_HVT U2644 ( .A(n4091), .Y(n4092) );
  INVX1_HVT U2645 ( .A(n4097), .Y(n4098) );
  INVX1_HVT U2646 ( .A(n4100), .Y(n4101) );
  INVX1_HVT U2647 ( .A(n4537), .Y(n4512) );
  INVX1_HVT U2648 ( .A(n4537), .Y(n4513) );
  INVX1_HVT U2649 ( .A(n4537), .Y(n4514) );
  INVX1_HVT U2650 ( .A(n4535), .Y(n4527) );
  INVX1_HVT U2651 ( .A(n4534), .Y(n4528) );
  INVX1_HVT U2652 ( .A(n4535), .Y(n4526) );
  INVX1_HVT U2653 ( .A(n4534), .Y(n4529) );
  INVX1_HVT U2654 ( .A(n4534), .Y(n4530) );
  INVX1_HVT U2655 ( .A(n4534), .Y(n4531) );
  INVX1_HVT U2656 ( .A(n4534), .Y(n4532) );
  INVX1_HVT U2657 ( .A(n4535), .Y(n4525) );
  INVX1_HVT U2658 ( .A(n4535), .Y(n4524) );
  INVX1_HVT U2659 ( .A(n4535), .Y(n4523) );
  INVX1_HVT U2660 ( .A(n4535), .Y(n4522) );
  INVX1_HVT U2661 ( .A(n4536), .Y(n4521) );
  INVX1_HVT U2662 ( .A(n4536), .Y(n4520) );
  INVX1_HVT U2663 ( .A(n4536), .Y(n4519) );
  INVX1_HVT U2664 ( .A(n4536), .Y(n4516) );
  INVX1_HVT U2665 ( .A(n4536), .Y(n4517) );
  INVX1_HVT U2666 ( .A(n4536), .Y(n4518) );
  INVX1_HVT U2667 ( .A(n4497), .Y(n4491) );
  INVX1_HVT U2668 ( .A(n4497), .Y(n4492) );
  INVX1_HVT U2669 ( .A(n4497), .Y(n4493) );
  INVX1_HVT U2670 ( .A(n4497), .Y(n4494) );
  INVX1_HVT U2671 ( .A(n4497), .Y(n4495) );
  INVX1_HVT U2672 ( .A(n4408), .Y(n4402) );
  INVX1_HVT U2673 ( .A(n4408), .Y(n4403) );
  INVX1_HVT U2674 ( .A(n4408), .Y(n4404) );
  INVX1_HVT U2675 ( .A(n4408), .Y(n4405) );
  INVX1_HVT U2676 ( .A(n4408), .Y(n4406) );
  INVX1_HVT U2677 ( .A(n4306), .Y(n4319) );
  INVX1_HVT U2678 ( .A(n4257), .Y(n4254) );
  INVX1_HVT U2679 ( .A(n4257), .Y(n4250) );
  INVX1_HVT U2680 ( .A(n4257), .Y(n4253) );
  INVX1_HVT U2681 ( .A(n4257), .Y(n4251) );
  INVX1_HVT U2682 ( .A(n4114), .Y(n4108) );
  INVX1_HVT U2683 ( .A(n4114), .Y(n4109) );
  INVX1_HVT U2684 ( .A(n4114), .Y(n4110) );
  INVX1_HVT U2685 ( .A(n4114), .Y(n4111) );
  INVX0_HVT U2686 ( .A(n1442), .Y(n4271) );
  INVX1_HVT U2687 ( .A(n4115), .Y(n4103) );
  INVX1_HVT U2688 ( .A(n4115), .Y(n4104) );
  INVX1_HVT U2689 ( .A(n4115), .Y(n4105) );
  INVX1_HVT U2690 ( .A(n4115), .Y(n4106) );
  INVX1_HVT U2691 ( .A(n4114), .Y(n4113) );
  INVX1_HVT U2692 ( .A(n4306), .Y(n4321) );
  INVX1_HVT U2693 ( .A(n4306), .Y(n4322) );
  INVX1_HVT U2694 ( .A(n4329), .Y(n4343) );
  INVX1_HVT U2695 ( .A(n4329), .Y(n4344) );
  INVX1_HVT U2696 ( .A(n4386), .Y(n4375) );
  INVX1_HVT U2697 ( .A(n4364), .Y(n4353) );
  INVX1_HVT U2698 ( .A(n4283), .Y(n4296) );
  INVX1_HVT U2699 ( .A(n4307), .Y(n4325) );
  INVX1_HVT U2700 ( .A(n4307), .Y(n4326) );
  INVX1_HVT U2701 ( .A(n4307), .Y(n4327) );
  INVX1_HVT U2702 ( .A(n4330), .Y(n4347) );
  INVX1_HVT U2703 ( .A(n4330), .Y(n4348) );
  INVX1_HVT U2704 ( .A(n4330), .Y(n4349) );
  INVX1_HVT U2705 ( .A(n4329), .Y(n4342) );
  INVX1_HVT U2706 ( .A(n4364), .Y(n4356) );
  INVX1_HVT U2707 ( .A(n4364), .Y(n4355) );
  INVX1_HVT U2708 ( .A(n4364), .Y(n4354) );
  INVX1_HVT U2709 ( .A(n4386), .Y(n4378) );
  INVX1_HVT U2710 ( .A(n4386), .Y(n4377) );
  INVX1_HVT U2711 ( .A(n4386), .Y(n4376) );
  INVX1_HVT U2712 ( .A(n4475), .Y(n4467) );
  INVX1_HVT U2713 ( .A(n4475), .Y(n4466) );
  INVX1_HVT U2714 ( .A(n4475), .Y(n4465) );
  INVX1_HVT U2715 ( .A(n4431), .Y(n4420) );
  INVX1_HVT U2716 ( .A(n4475), .Y(n4464) );
  INVX1_HVT U2717 ( .A(n4453), .Y(n4442) );
  INVX1_HVT U2718 ( .A(n4256), .Y(n4245) );
  INVX1_HVT U2719 ( .A(n4256), .Y(n4246) );
  INVX1_HVT U2720 ( .A(n4256), .Y(n4247) );
  INVX1_HVT U2721 ( .A(n4497), .Y(n4496) );
  INVX1_HVT U2722 ( .A(n4408), .Y(n4407) );
  INVX1_HVT U2723 ( .A(n4283), .Y(n4295) );
  INVX1_HVT U2724 ( .A(n4453), .Y(n4444) );
  INVX1_HVT U2725 ( .A(n4453), .Y(n4445) );
  INVX1_HVT U2726 ( .A(n4453), .Y(n4443) );
  INVX1_HVT U2727 ( .A(n4431), .Y(n4423) );
  INVX1_HVT U2728 ( .A(n4431), .Y(n4422) );
  INVX1_HVT U2729 ( .A(n4363), .Y(n4360) );
  INVX1_HVT U2730 ( .A(n4363), .Y(n4359) );
  INVX1_HVT U2731 ( .A(n4363), .Y(n4358) );
  INVX1_HVT U2732 ( .A(n4363), .Y(n4357) );
  INVX1_HVT U2733 ( .A(n4363), .Y(n4362) );
  INVX1_HVT U2734 ( .A(n4363), .Y(n4361) );
  INVX1_HVT U2735 ( .A(n4385), .Y(n4382) );
  INVX1_HVT U2736 ( .A(n4385), .Y(n4381) );
  INVX1_HVT U2737 ( .A(n4385), .Y(n4380) );
  INVX1_HVT U2738 ( .A(n4385), .Y(n4379) );
  INVX1_HVT U2739 ( .A(n4385), .Y(n4384) );
  INVX1_HVT U2740 ( .A(n4385), .Y(n4383) );
  INVX1_HVT U2741 ( .A(n4306), .Y(n4324) );
  INVX1_HVT U2742 ( .A(n4329), .Y(n4346) );
  INVX1_HVT U2743 ( .A(n4114), .Y(n4112) );
  INVX1_HVT U2744 ( .A(n4409), .Y(n4397) );
  INVX1_HVT U2745 ( .A(n4409), .Y(n4398) );
  INVX1_HVT U2746 ( .A(n4409), .Y(n4399) );
  INVX1_HVT U2747 ( .A(n4409), .Y(n4400) );
  INVX1_HVT U2748 ( .A(n4409), .Y(n4401) );
  INVX1_HVT U2749 ( .A(n4498), .Y(n4486) );
  INVX1_HVT U2750 ( .A(n4498), .Y(n4487) );
  INVX1_HVT U2751 ( .A(n4498), .Y(n4488) );
  INVX1_HVT U2752 ( .A(n4498), .Y(n4489) );
  INVX1_HVT U2753 ( .A(n4498), .Y(n4490) );
  INVX1_HVT U2754 ( .A(n4306), .Y(n4320) );
  INVX1_HVT U2755 ( .A(n4329), .Y(n4341) );
  INVX1_HVT U2756 ( .A(n4474), .Y(n4471) );
  INVX1_HVT U2757 ( .A(n4474), .Y(n4470) );
  INVX1_HVT U2758 ( .A(n4474), .Y(n4469) );
  INVX1_HVT U2759 ( .A(n4474), .Y(n4468) );
  INVX1_HVT U2760 ( .A(n4474), .Y(n4473) );
  INVX1_HVT U2761 ( .A(n4474), .Y(n4472) );
  INVX1_HVT U2762 ( .A(n4452), .Y(n4451) );
  INVX1_HVT U2763 ( .A(n4452), .Y(n4446) );
  INVX1_HVT U2764 ( .A(n4452), .Y(n4447) );
  INVX1_HVT U2765 ( .A(n4452), .Y(n4448) );
  INVX1_HVT U2766 ( .A(n4452), .Y(n4449) );
  INVX1_HVT U2767 ( .A(n4452), .Y(n4450) );
  INVX1_HVT U2768 ( .A(n4430), .Y(n4427) );
  INVX1_HVT U2769 ( .A(n4430), .Y(n4426) );
  INVX1_HVT U2770 ( .A(n4430), .Y(n4425) );
  INVX1_HVT U2771 ( .A(n4430), .Y(n4424) );
  INVX1_HVT U2772 ( .A(n4430), .Y(n4428) );
  INVX1_HVT U2773 ( .A(n4256), .Y(n4255) );
  INVX1_HVT U2774 ( .A(n4256), .Y(n4249) );
  INVX1_HVT U2775 ( .A(n4115), .Y(n4107) );
  INVX1_HVT U2776 ( .A(n4430), .Y(n4429) );
  INVX1_HVT U2777 ( .A(n4307), .Y(n4328) );
  INVX1_HVT U2778 ( .A(n4330), .Y(n4350) );
  INVX1_HVT U2779 ( .A(n4284), .Y(n4301) );
  INVX1_HVT U2780 ( .A(n4284), .Y(n4302) );
  INVX1_HVT U2781 ( .A(n4284), .Y(n4303) );
  INVX1_HVT U2782 ( .A(n4283), .Y(n4297) );
  INVX1_HVT U2783 ( .A(n4283), .Y(n4298) );
  INVX1_HVT U2784 ( .A(n4283), .Y(n4299) );
  INVX1_HVT U2785 ( .A(n4282), .Y(n4272) );
  INVX1_HVT U2786 ( .A(n4282), .Y(n4273) );
  INVX1_HVT U2787 ( .A(n4282), .Y(n4274) );
  INVX1_HVT U2788 ( .A(n4282), .Y(n4275) );
  INVX1_HVT U2789 ( .A(n4282), .Y(n4278) );
  INVX1_HVT U2790 ( .A(n4282), .Y(n4280) );
  INVX1_HVT U2791 ( .A(n4282), .Y(n4281) );
  INVX1_HVT U2792 ( .A(n4284), .Y(n4305) );
  INVX1_HVT U2793 ( .A(n4283), .Y(n4300) );
  INVX1_HVT U2794 ( .A(n4284), .Y(n4304) );
  INVX1_HVT U2795 ( .A(n4282), .Y(n4276) );
  NBUFFX2_HVT U2796 ( .A(keyout[13]), .Y(n4034) );
  NBUFFX2_HVT U2797 ( .A(keyout[21]), .Y(n4058) );
  NBUFFX2_HVT U2798 ( .A(keyout[13]), .Y(n4033) );
  NBUFFX2_HVT U2799 ( .A(keyout[21]), .Y(n4057) );
  NBUFFX2_HVT U2800 ( .A(keyout[13]), .Y(n4032) );
  NBUFFX2_HVT U2801 ( .A(keyout[21]), .Y(n4056) );
  NBUFFX2_HVT U2802 ( .A(keyout[10]), .Y(n4025) );
  NBUFFX2_HVT U2803 ( .A(keyout[18]), .Y(n4049) );
  NBUFFX2_HVT U2804 ( .A(keyout[10]), .Y(n4024) );
  NBUFFX2_HVT U2805 ( .A(keyout[18]), .Y(n4048) );
  NBUFFX2_HVT U2806 ( .A(keyout[18]), .Y(n4047) );
  NBUFFX2_HVT U2807 ( .A(keyout[10]), .Y(n4023) );
  INVX0_HVT U2808 ( .A(keyout[88]), .Y(n4091) );
  NBUFFX2_HVT U2809 ( .A(keyout[12]), .Y(n4029) );
  NBUFFX2_HVT U2810 ( .A(keyout[20]), .Y(n4053) );
  NBUFFX2_HVT U2811 ( .A(keyout[30]), .Y(n4083) );
  NBUFFX2_HVT U2812 ( .A(keyout[12]), .Y(n4031) );
  NBUFFX2_HVT U2813 ( .A(keyout[20]), .Y(n4055) );
  NBUFFX2_HVT U2814 ( .A(keyout[12]), .Y(n4030) );
  NBUFFX2_HVT U2815 ( .A(keyout[20]), .Y(n4054) );
  NBUFFX2_HVT U2816 ( .A(keyout[30]), .Y(n4082) );
  INVX0_HVT U2817 ( .A(keyout[126]), .Y(n4097) );
  INVX0_HVT U2818 ( .A(keyout[127]), .Y(n4100) );
  NBUFFX2_HVT U2819 ( .A(keyout[11]), .Y(n4028) );
  NBUFFX2_HVT U2820 ( .A(keyout[19]), .Y(n4052) );
  NBUFFX2_HVT U2821 ( .A(keyout[11]), .Y(n4027) );
  NBUFFX2_HVT U2822 ( .A(keyout[19]), .Y(n4051) );
  NBUFFX2_HVT U2823 ( .A(keyout[19]), .Y(n4050) );
  NBUFFX2_HVT U2824 ( .A(keyout[11]), .Y(n4026) );
  INVX1_HVT U2825 ( .A(n4094), .Y(n4095) );
  NBUFFX2_HVT U2826 ( .A(keyout[8]), .Y(n4019) );
  NBUFFX2_HVT U2827 ( .A(keyout[16]), .Y(n4043) );
  NBUFFX2_HVT U2828 ( .A(keyout[8]), .Y(n4018) );
  NBUFFX2_HVT U2829 ( .A(keyout[16]), .Y(n4042) );
  NBUFFX2_HVT U2830 ( .A(keyout[14]), .Y(n4037) );
  NBUFFX2_HVT U2831 ( .A(keyout[22]), .Y(n4061) );
  NBUFFX2_HVT U2832 ( .A(keyout[14]), .Y(n4036) );
  NBUFFX2_HVT U2833 ( .A(keyout[22]), .Y(n4060) );
  NBUFFX2_HVT U2834 ( .A(keyout[15]), .Y(n4040) );
  NBUFFX2_HVT U2835 ( .A(keyout[23]), .Y(n4064) );
  NBUFFX2_HVT U2836 ( .A(keyout[15]), .Y(n4039) );
  NBUFFX2_HVT U2837 ( .A(keyout[23]), .Y(n4063) );
  NBUFFX2_HVT U2838 ( .A(keyout[9]), .Y(n4022) );
  NBUFFX2_HVT U2839 ( .A(keyout[17]), .Y(n4046) );
  NBUFFX2_HVT U2840 ( .A(keyout[9]), .Y(n4021) );
  NBUFFX2_HVT U2841 ( .A(keyout[17]), .Y(n4045) );
  NBUFFX2_HVT U2842 ( .A(keyout[16]), .Y(n4041) );
  NBUFFX2_HVT U2843 ( .A(keyout[8]), .Y(n4017) );
  NBUFFX2_HVT U2844 ( .A(keyout[14]), .Y(n4035) );
  NBUFFX2_HVT U2845 ( .A(keyout[22]), .Y(n4059) );
  NBUFFX2_HVT U2846 ( .A(keyout[15]), .Y(n4038) );
  NBUFFX2_HVT U2847 ( .A(keyout[23]), .Y(n4062) );
  NBUFFX2_HVT U2848 ( .A(keyout[17]), .Y(n4044) );
  NBUFFX2_HVT U2849 ( .A(keyout[9]), .Y(n4020) );
  NBUFFX2_HVT U2850 ( .A(keyout[7]), .Y(n4016) );
  NBUFFX2_HVT U2851 ( .A(keyout[3]), .Y(n4006) );
  NBUFFX2_HVT U2852 ( .A(keyout[3]), .Y(n4005) );
  NBUFFX2_HVT U2853 ( .A(keyout[3]), .Y(n4004) );
  NBUFFX2_HVT U2854 ( .A(keyout[2]), .Y(n4003) );
  NBUFFX2_HVT U2855 ( .A(keyout[6]), .Y(n4015) );
  NBUFFX2_HVT U2856 ( .A(keyout[6]), .Y(n4014) );
  NBUFFX2_HVT U2857 ( .A(keyout[5]), .Y(n4012) );
  NBUFFX2_HVT U2858 ( .A(keyout[5]), .Y(n4011) );
  NBUFFX2_HVT U2859 ( .A(keyout[6]), .Y(n4013) );
  NBUFFX2_HVT U2860 ( .A(keyout[5]), .Y(n4010) );
  NBUFFX2_HVT U2861 ( .A(keyout[1]), .Y(n4000) );
  NBUFFX2_HVT U2862 ( .A(keyout[1]), .Y(n4002) );
  NBUFFX2_HVT U2863 ( .A(keyout[1]), .Y(n4001) );
  NBUFFX2_HVT U2864 ( .A(keyout[4]), .Y(n4009) );
  NBUFFX2_HVT U2865 ( .A(keyout[4]), .Y(n4008) );
  NBUFFX2_HVT U2866 ( .A(keyout[4]), .Y(n4007) );
  NBUFFX2_HVT U2867 ( .A(keyout[0]), .Y(n3999) );
  NBUFFX2_HVT U2868 ( .A(keyout[0]), .Y(n3998) );
  NBUFFX2_HVT U2869 ( .A(keyout[0]), .Y(n3997) );
  INVX1_HVT U2870 ( .A(n4507), .Y(n4535) );
  INVX1_HVT U2871 ( .A(n4507), .Y(n4534) );
  INVX1_HVT U2872 ( .A(n4140), .Y(n4134) );
  INVX1_HVT U2873 ( .A(n4140), .Y(n4135) );
  INVX1_HVT U2874 ( .A(n4140), .Y(n4136) );
  INVX1_HVT U2875 ( .A(n4140), .Y(n4137) );
  INVX1_HVT U2876 ( .A(n4141), .Y(n4129) );
  INVX1_HVT U2877 ( .A(n4141), .Y(n4130) );
  INVX1_HVT U2878 ( .A(n4141), .Y(n4131) );
  INVX1_HVT U2879 ( .A(n4141), .Y(n4132) );
  INVX1_HVT U2880 ( .A(n4484), .Y(n4497) );
  INVX1_HVT U2881 ( .A(n4395), .Y(n4408) );
  INVX1_HVT U2882 ( .A(n3987), .Y(n4306) );
  INVX1_HVT U2883 ( .A(n4128), .Y(n4116) );
  INVX1_HVT U2884 ( .A(n4128), .Y(n4117) );
  INVX1_HVT U2885 ( .A(n4128), .Y(n4118) );
  INVX1_HVT U2886 ( .A(n4128), .Y(n4119) );
  INVX1_HVT U2887 ( .A(n4167), .Y(n4155) );
  INVX1_HVT U2888 ( .A(n4167), .Y(n4156) );
  INVX1_HVT U2889 ( .A(n4167), .Y(n4157) );
  INVX1_HVT U2890 ( .A(n4167), .Y(n4158) );
  INVX1_HVT U2891 ( .A(n4166), .Y(n4160) );
  INVX1_HVT U2892 ( .A(n4166), .Y(n4161) );
  INVX1_HVT U2893 ( .A(n4166), .Y(n4162) );
  INVX1_HVT U2894 ( .A(n4166), .Y(n4163) );
  INVX1_HVT U2895 ( .A(n1487), .Y(n4114) );
  INVX1_HVT U2896 ( .A(n4193), .Y(n4181) );
  INVX1_HVT U2897 ( .A(n4193), .Y(n4182) );
  INVX1_HVT U2898 ( .A(n4193), .Y(n4183) );
  INVX1_HVT U2899 ( .A(n4193), .Y(n4184) );
  INVX1_HVT U2900 ( .A(n4206), .Y(n4194) );
  INVX1_HVT U2901 ( .A(n4206), .Y(n4195) );
  INVX1_HVT U2902 ( .A(n4206), .Y(n4196) );
  INVX1_HVT U2903 ( .A(n4206), .Y(n4197) );
  INVX1_HVT U2904 ( .A(n4180), .Y(n4168) );
  INVX1_HVT U2905 ( .A(n4180), .Y(n4169) );
  INVX1_HVT U2906 ( .A(n4180), .Y(n4170) );
  INVX1_HVT U2907 ( .A(n4180), .Y(n4171) );
  INVX1_HVT U2908 ( .A(n4127), .Y(n4121) );
  INVX1_HVT U2909 ( .A(n4127), .Y(n4122) );
  INVX1_HVT U2910 ( .A(n4127), .Y(n4123) );
  INVX1_HVT U2911 ( .A(n4127), .Y(n4124) );
  INVX1_HVT U2912 ( .A(n4205), .Y(n4199) );
  INVX1_HVT U2913 ( .A(n4205), .Y(n4200) );
  INVX1_HVT U2914 ( .A(n4205), .Y(n4201) );
  INVX1_HVT U2915 ( .A(n4205), .Y(n4202) );
  INVX1_HVT U2916 ( .A(n4179), .Y(n4173) );
  INVX1_HVT U2917 ( .A(n4179), .Y(n4174) );
  INVX1_HVT U2918 ( .A(n4179), .Y(n4175) );
  INVX1_HVT U2919 ( .A(n4179), .Y(n4176) );
  INVX1_HVT U2920 ( .A(n4243), .Y(n4237) );
  INVX1_HVT U2921 ( .A(n4243), .Y(n4238) );
  INVX1_HVT U2922 ( .A(n4243), .Y(n4239) );
  INVX1_HVT U2923 ( .A(n4243), .Y(n4240) );
  INVX1_HVT U2924 ( .A(n4153), .Y(n4147) );
  INVX1_HVT U2925 ( .A(n4153), .Y(n4148) );
  INVX1_HVT U2926 ( .A(n4153), .Y(n4149) );
  INVX1_HVT U2927 ( .A(n4153), .Y(n4150) );
  INVX1_HVT U2928 ( .A(n4153), .Y(n4152) );
  INVX1_HVT U2929 ( .A(n4192), .Y(n4186) );
  INVX1_HVT U2930 ( .A(n4192), .Y(n4187) );
  INVX1_HVT U2931 ( .A(n4192), .Y(n4188) );
  INVX1_HVT U2932 ( .A(n4192), .Y(n4189) );
  INVX0_HVT U2933 ( .A(n1487), .Y(n4115) );
  INVX1_HVT U2934 ( .A(n4243), .Y(n4242) );
  INVX1_HVT U2935 ( .A(n4230), .Y(n4224) );
  INVX1_HVT U2936 ( .A(n4230), .Y(n4225) );
  INVX1_HVT U2937 ( .A(n4230), .Y(n4226) );
  INVX1_HVT U2938 ( .A(n4230), .Y(n4227) );
  INVX1_HVT U2939 ( .A(n4218), .Y(n4217) );
  INVX1_HVT U2940 ( .A(n4218), .Y(n4212) );
  INVX1_HVT U2941 ( .A(n4218), .Y(n4213) );
  INVX1_HVT U2942 ( .A(n4218), .Y(n4214) );
  INVX1_HVT U2943 ( .A(n4218), .Y(n4215) );
  INVX1_HVT U2944 ( .A(n4244), .Y(n4232) );
  INVX1_HVT U2945 ( .A(n4244), .Y(n4233) );
  INVX1_HVT U2946 ( .A(n4244), .Y(n4234) );
  INVX1_HVT U2947 ( .A(n4244), .Y(n4235) );
  INVX1_HVT U2948 ( .A(n4231), .Y(n4220) );
  INVX1_HVT U2949 ( .A(n4231), .Y(n4221) );
  INVX1_HVT U2950 ( .A(n4231), .Y(n4222) );
  INVX1_HVT U2951 ( .A(n4154), .Y(n4142) );
  INVX1_HVT U2952 ( .A(n4154), .Y(n4143) );
  INVX1_HVT U2953 ( .A(n4154), .Y(n4144) );
  INVX1_HVT U2954 ( .A(n4154), .Y(n4145) );
  INVX1_HVT U2955 ( .A(n4351), .Y(n4365) );
  INVX1_HVT U2956 ( .A(n4351), .Y(n4366) );
  INVX1_HVT U2957 ( .A(n4351), .Y(n4367) );
  INVX1_HVT U2958 ( .A(n4373), .Y(n4387) );
  INVX1_HVT U2959 ( .A(n4373), .Y(n4388) );
  INVX1_HVT U2960 ( .A(n4462), .Y(n4476) );
  INVX1_HVT U2961 ( .A(n4462), .Y(n4477) );
  INVX1_HVT U2962 ( .A(n4462), .Y(n4478) );
  INVX1_HVT U2963 ( .A(n4395), .Y(n4410) );
  INVX1_HVT U2964 ( .A(n4395), .Y(n4411) );
  INVX1_HVT U2965 ( .A(n4395), .Y(n4412) );
  INVX1_HVT U2966 ( .A(n4440), .Y(n4454) );
  INVX1_HVT U2967 ( .A(n4440), .Y(n4455) );
  INVX1_HVT U2968 ( .A(n4440), .Y(n4456) );
  INVX1_HVT U2969 ( .A(n4418), .Y(n4432) );
  INVX1_HVT U2970 ( .A(n4418), .Y(n4433) );
  INVX1_HVT U2971 ( .A(n4418), .Y(n4434) );
  INVX1_HVT U2972 ( .A(n4351), .Y(n4364) );
  INVX1_HVT U2973 ( .A(n4373), .Y(n4386) );
  INVX1_HVT U2974 ( .A(n3988), .Y(n4329) );
  INVX1_HVT U2975 ( .A(n4167), .Y(n4159) );
  INVX1_HVT U2976 ( .A(n4166), .Y(n4164) );
  INVX1_HVT U2977 ( .A(n4484), .Y(n4501) );
  INVX1_HVT U2978 ( .A(n4352), .Y(n4369) );
  INVX1_HVT U2979 ( .A(n4352), .Y(n4370) );
  INVX1_HVT U2980 ( .A(n4352), .Y(n4371) );
  INVX1_HVT U2981 ( .A(n4374), .Y(n4391) );
  INVX1_HVT U2982 ( .A(n4374), .Y(n4392) );
  INVX1_HVT U2983 ( .A(n4374), .Y(n4393) );
  INVX1_HVT U2984 ( .A(n4463), .Y(n4480) );
  INVX1_HVT U2985 ( .A(n4463), .Y(n4481) );
  INVX1_HVT U2986 ( .A(n4463), .Y(n4482) );
  INVX1_HVT U2987 ( .A(n4485), .Y(n4503) );
  INVX1_HVT U2988 ( .A(n4485), .Y(n4504) );
  INVX1_HVT U2989 ( .A(n4485), .Y(n4505) );
  INVX1_HVT U2990 ( .A(n4396), .Y(n4414) );
  INVX1_HVT U2991 ( .A(n4396), .Y(n4415) );
  INVX1_HVT U2992 ( .A(n4396), .Y(n4416) );
  INVX1_HVT U2993 ( .A(n4441), .Y(n4459) );
  INVX1_HVT U2994 ( .A(n4441), .Y(n4460) );
  INVX1_HVT U2995 ( .A(n4419), .Y(n4436) );
  INVX1_HVT U2996 ( .A(n4419), .Y(n4437) );
  INVX1_HVT U2997 ( .A(n4484), .Y(n4500) );
  INVX1_HVT U2998 ( .A(n4484), .Y(n4499) );
  INVX1_HVT U2999 ( .A(n4462), .Y(n4475) );
  INVX1_HVT U3000 ( .A(n4440), .Y(n4453) );
  INVX1_HVT U3001 ( .A(n4418), .Y(n4431) );
  INVX1_HVT U3002 ( .A(n3989), .Y(n4283) );
  INVX1_HVT U3003 ( .A(n3987), .Y(n4307) );
  INVX1_HVT U3004 ( .A(n4128), .Y(n4120) );
  INVX1_HVT U3005 ( .A(n4179), .Y(n4177) );
  INVX1_HVT U3006 ( .A(n4127), .Y(n4125) );
  INVX1_HVT U3007 ( .A(n4205), .Y(n4203) );
  INVX1_HVT U3008 ( .A(n4192), .Y(n4190) );
  INVX1_HVT U3009 ( .A(n4166), .Y(n4165) );
  INVX1_HVT U3010 ( .A(n4140), .Y(n4138) );
  INVX1_HVT U3011 ( .A(n4219), .Y(n4207) );
  INVX1_HVT U3012 ( .A(n4219), .Y(n4208) );
  INVX1_HVT U3013 ( .A(n4219), .Y(n4209) );
  INVX1_HVT U3014 ( .A(n4219), .Y(n4210) );
  INVX1_HVT U3015 ( .A(n4507), .Y(n4539) );
  INVX1_HVT U3016 ( .A(n4508), .Y(n4545) );
  INVX1_HVT U3017 ( .A(n4509), .Y(n4551) );
  INVX1_HVT U3018 ( .A(n4351), .Y(n4363) );
  INVX1_HVT U3019 ( .A(n4373), .Y(n4385) );
  INVX1_HVT U3020 ( .A(n4180), .Y(n4172) );
  INVX1_HVT U3021 ( .A(n4206), .Y(n4198) );
  INVX1_HVT U3022 ( .A(n4193), .Y(n4185) );
  INVX1_HVT U3023 ( .A(n4462), .Y(n4479) );
  INVX1_HVT U3024 ( .A(n4484), .Y(n4502) );
  INVX1_HVT U3025 ( .A(n4440), .Y(n4457) );
  INVX1_HVT U3026 ( .A(n4418), .Y(n4435) );
  INVX1_HVT U3027 ( .A(n4373), .Y(n4390) );
  INVX1_HVT U3028 ( .A(n4351), .Y(n4368) );
  INVX1_HVT U3029 ( .A(n4153), .Y(n4151) );
  INVX1_HVT U3030 ( .A(n4127), .Y(n4126) );
  INVX1_HVT U3031 ( .A(n4141), .Y(n4133) );
  INVX1_HVT U3032 ( .A(n4395), .Y(n4409) );
  INVX1_HVT U3033 ( .A(n4484), .Y(n4498) );
  INVX1_HVT U3034 ( .A(n4462), .Y(n4474) );
  INVX1_HVT U3035 ( .A(n4440), .Y(n4452) );
  INVX1_HVT U3036 ( .A(n4418), .Y(n4430) );
  INVX1_HVT U3037 ( .A(n4510), .Y(n4553) );
  INVX1_HVT U3038 ( .A(n4510), .Y(n4552) );
  INVX1_HVT U3039 ( .A(n4230), .Y(n4228) );
  INVX1_HVT U3040 ( .A(n4243), .Y(n4241) );
  INVX1_HVT U3041 ( .A(n4244), .Y(n4236) );
  INVX1_HVT U3042 ( .A(n4154), .Y(n4146) );
  INVX1_HVT U3043 ( .A(n4179), .Y(n4178) );
  INVX1_HVT U3044 ( .A(n4205), .Y(n4204) );
  INVX1_HVT U3045 ( .A(n4192), .Y(n4191) );
  INVX1_HVT U3046 ( .A(n4485), .Y(n4506) );
  INVX1_HVT U3047 ( .A(n4218), .Y(n4216) );
  INVX1_HVT U3048 ( .A(n4231), .Y(n4223) );
  INVX1_HVT U3049 ( .A(n4508), .Y(n4542) );
  INVX1_HVT U3050 ( .A(n4508), .Y(n4540) );
  INVX1_HVT U3051 ( .A(n4508), .Y(n4541) );
  INVX1_HVT U3052 ( .A(n4507), .Y(n4538) );
  INVX1_HVT U3053 ( .A(n4508), .Y(n4544) );
  INVX1_HVT U3054 ( .A(n4508), .Y(n4543) );
  INVX1_HVT U3055 ( .A(n4509), .Y(n4546) );
  INVX1_HVT U3056 ( .A(n4509), .Y(n4550) );
  INVX1_HVT U3057 ( .A(n4509), .Y(n4549) );
  INVX1_HVT U3058 ( .A(n4509), .Y(n4548) );
  INVX1_HVT U3059 ( .A(n4509), .Y(n4547) );
  INVX1_HVT U3060 ( .A(n4219), .Y(n4211) );
  INVX1_HVT U3061 ( .A(n4230), .Y(n4229) );
  INVX1_HVT U3062 ( .A(n4396), .Y(n4417) );
  INVX1_HVT U3063 ( .A(n4510), .Y(n4554) );
  INVX1_HVT U3064 ( .A(n4463), .Y(n4483) );
  INVX1_HVT U3065 ( .A(n4441), .Y(n4461) );
  INVX1_HVT U3066 ( .A(n4419), .Y(n4439) );
  INVX1_HVT U3067 ( .A(n4374), .Y(n4394) );
  INVX1_HVT U3068 ( .A(n4352), .Y(n4372) );
  INVX0_HVT U3069 ( .A(n1443), .Y(n4258) );
  INVX1_HVT U3070 ( .A(n3989), .Y(n4284) );
  NBUFFX2_HVT U3071 ( .A(keyout[29]), .Y(n4080) );
  NBUFFX2_HVT U3072 ( .A(keyout[29]), .Y(n4079) );
  NBUFFX2_HVT U3073 ( .A(keyout[58]), .Y(n4087) );
  NBUFFX2_HVT U3074 ( .A(keyout[26]), .Y(n4072) );
  NBUFFX2_HVT U3075 ( .A(keyout[26]), .Y(n4071) );
  NBUFFX2_HVT U3076 ( .A(keyout[28]), .Y(n4078) );
  NBUFFX2_HVT U3077 ( .A(keyout[28]), .Y(n4077) );
  NBUFFX2_HVT U3078 ( .A(keyout[59]), .Y(n4090) );
  NBUFFX2_HVT U3079 ( .A(keyout[27]), .Y(n4075) );
  NBUFFX2_HVT U3080 ( .A(keyout[27]), .Y(n4074) );
  NBUFFX2_HVT U3081 ( .A(keyout[24]), .Y(n4067) );
  NBUFFX2_HVT U3082 ( .A(keyout[24]), .Y(n4066) );
  NBUFFX2_HVT U3083 ( .A(keyout[59]), .Y(n4089) );
  NBUFFX2_HVT U3084 ( .A(keyout[27]), .Y(n4073) );
  NBUFFX2_HVT U3085 ( .A(keyout[24]), .Y(n4065) );
  NBUFFX2_HVT U3086 ( .A(keyout[59]), .Y(n4088) );
  NBUFFX2_HVT U3087 ( .A(keyout[57]), .Y(n4085) );
  NBUFFX2_HVT U3088 ( .A(keyout[25]), .Y(n4069) );
  NBUFFX2_HVT U3089 ( .A(keyout[25]), .Y(n4068) );
  INVX0_HVT U3090 ( .A(keyout[120]), .Y(n4094) );
  INVX1_HVT U3091 ( .A(n4511), .Y(n4507) );
  INVX1_HVT U3092 ( .A(n3991), .Y(n4395) );
  INVX1_HVT U3093 ( .A(n3990), .Y(n4484) );
  INVX0_HVT U3094 ( .A(n1485), .Y(n4141) );
  AND2X1_HVT U3095 ( .A1(n1469), .A2(n4559), .Y(n3987) );
  INVX1_HVT U3096 ( .A(n1483), .Y(n4167) );
  INVX1_HVT U3097 ( .A(n1486), .Y(n4128) );
  INVX0_HVT U3098 ( .A(n1483), .Y(n4166) );
  INVX1_HVT U3099 ( .A(n1480), .Y(n4206) );
  INVX1_HVT U3100 ( .A(n1482), .Y(n4180) );
  INVX1_HVT U3101 ( .A(n1481), .Y(n4193) );
  INVX0_HVT U3102 ( .A(n1486), .Y(n4127) );
  INVX0_HVT U3103 ( .A(n1480), .Y(n4205) );
  INVX0_HVT U3104 ( .A(n1482), .Y(n4179) );
  INVX0_HVT U3105 ( .A(n1481), .Y(n4192) );
  INVX1_HVT U3106 ( .A(n1477), .Y(n4243) );
  INVX1_HVT U3107 ( .A(n1484), .Y(n4153) );
  INVX1_HVT U3108 ( .A(n1478), .Y(n4230) );
  INVX1_HVT U3109 ( .A(n3994), .Y(n4462) );
  INVX1_HVT U3110 ( .A(n3995), .Y(n4440) );
  INVX1_HVT U3111 ( .A(n3996), .Y(n4418) );
  INVX1_HVT U3112 ( .A(n3993), .Y(n4373) );
  INVX1_HVT U3113 ( .A(n3992), .Y(n4351) );
  INVX1_HVT U3114 ( .A(n1479), .Y(n4218) );
  INVX0_HVT U3115 ( .A(n1478), .Y(n4231) );
  INVX0_HVT U3116 ( .A(n1477), .Y(n4244) );
  INVX0_HVT U3117 ( .A(n1484), .Y(n4154) );
  AND2X1_HVT U3118 ( .A1(n4556), .A2(n4559), .Y(n3988) );
  INVX1_HVT U3119 ( .A(n3990), .Y(n4485) );
  INVX1_HVT U3120 ( .A(n3991), .Y(n4396) );
  AND2X1_HVT U3121 ( .A1(n1454), .A2(n4559), .Y(n3989) );
  INVX1_HVT U3122 ( .A(n4511), .Y(n4508) );
  INVX1_HVT U3123 ( .A(n4511), .Y(n4509) );
  INVX0_HVT U3124 ( .A(n1479), .Y(n4219) );
  INVX1_HVT U3125 ( .A(n1430), .Y(n4511) );
  NOR2X1_HVT U3126 ( .A1(n1447), .A2(rest), .Y(n3990) );
  NOR2X1_HVT U3127 ( .A1(n1450), .A2(rest), .Y(n3991) );
  NOR2X1_HVT U3128 ( .A1(n1449), .A2(rest), .Y(n3992) );
  NOR2X1_HVT U3129 ( .A1(n1457), .A2(rest), .Y(n3993) );
  NOR2X1_HVT U3130 ( .A1(n1456), .A2(rest), .Y(n3994) );
  NOR2X1_HVT U3131 ( .A1(n1466), .A2(rest), .Y(n3995) );
  NOR2X1_HVT U3132 ( .A1(n1458), .A2(rest), .Y(n3996) );
  INVX0_HVT U3133 ( .A(n1452), .Y(n4555) );
  INVX0_HVT U3134 ( .A(n1455), .Y(n4556) );
  INVX0_HVT U3135 ( .A(rount_no[0]), .Y(n4557) );
  INVX0_HVT U3136 ( .A(rount_no[1]), .Y(n4558) );
  INVX0_HVT U3137 ( .A(rest), .Y(n4559) );
endmodule

