
module inv_sbox_0 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n203, n204, n205, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n196, n197,
         n198, n199, n200, n201, n202, n206, n208, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454;

  NAND2X0_HVT U4 ( .A1(n384), .A2(n383), .Y(n4) );
  NAND2X0_HVT U5 ( .A1(n4), .A2(n378), .Y(n5) );
  NAND2X0_HVT U7 ( .A1(n327), .A2(n380), .Y(n8) );
  NAND2X0_HVT U8 ( .A1(n384), .A2(n378), .Y(n9) );
  NAND2X0_HVT U9 ( .A1(n277), .A2(n9), .Y(n10) );
  NAND2X0_HVT U10 ( .A1(n1), .A2(n12), .Y(n11) );
  NAND2X0_HVT U11 ( .A1(n331), .A2(n383), .Y(n13) );
  NAND2X0_HVT U12 ( .A1(n290), .A2(n364), .Y(n14) );
  NAND2X0_HVT U13 ( .A1(n381), .A2(n9), .Y(n15) );
  NAND2X0_HVT U19 ( .A1(n289), .A2(n452), .Y(n22) );
  NAND2X0_HVT U25 ( .A1(in[6]), .A2(n365), .Y(n6) );
  NAND2X0_HVT U32 ( .A1(n367), .A2(n326), .Y(n34) );
  NAND2X0_HVT U35 ( .A1(n9), .A2(n234), .Y(n37) );
  NAND2X0_HVT U38 ( .A1(n364), .A2(n331), .Y(n40) );
  NAND2X0_HVT U42 ( .A1(n7), .A2(n453), .Y(n44) );
  OA21X1_HVT U53 ( .A1(n328), .A2(n52), .A3(n421), .Y(n54) );
  NAND2X0_HVT U55 ( .A1(n381), .A2(n4), .Y(n56) );
  MUX41X1_HVT U56 ( .A1(n329), .A3(n376), .A2(n419), .A4(n56), .S0(n358), .S1(
        n310), .Y(n57) );
  AO21X1_HVT U60 ( .A1(n62), .A2(n361), .A3(n23), .Y(n61) );
  NAND2X0_HVT U66 ( .A1(n387), .A2(n352), .Y(n68) );
  MUX41X1_HVT U67 ( .A1(n410), .A3(n435), .A2(n412), .A4(n68), .S0(n362), .S1(
        n355), .Y(n69) );
  MUX41X1_HVT U68 ( .A1(n410), .A3(n342), .A2(n411), .A4(n1), .S0(n357), .S1(
        n309), .Y(n70) );
  MUX41X1_HVT U71 ( .A1(n305), .A3(n279), .A2(n13), .A4(n406), .S0(n357), .S1(
        n336), .Y(n72) );
  NAND2X0_HVT U72 ( .A1(n375), .A2(n8), .Y(n73) );
  MUX41X1_HVT U74 ( .A1(n11), .A3(n426), .A2(n425), .A4(n416), .S0(n358), .S1(
        n336), .Y(n75) );
  MUX41X1_HVT U78 ( .A1(n78), .A3(n74), .A2(n75), .A4(n72), .S0(n372), .S1(
        n370), .Y(n79) );
  MUX41X1_HVT U79 ( .A1(n422), .A3(n20), .A2(n424), .A4(n19), .S0(n358), .S1(
        n391), .Y(n80) );
  MUX41X1_HVT U80 ( .A1(n437), .A3(n329), .A2(n10), .A4(n303), .S0(n357), .S1(
        n336), .Y(n81) );
  NAND2X0_HVT U81 ( .A1(n260), .A2(n8), .Y(n82) );
  AND2X1_HVT U82 ( .A1(n305), .A2(n379), .Y(n83) );
  MUX41X1_HVT U83 ( .A1(n83), .A3(n423), .A2(n438), .A4(n82), .S0(n357), .S1(
        n336), .Y(n84) );
  MUX41X1_HVT U84 ( .A1(n349), .A3(n294), .A2(n439), .A4(n27), .S0(n358), .S1(
        n336), .Y(n85) );
  MUX41X1_HVT U85 ( .A1(n85), .A3(n81), .A2(n84), .A4(n80), .S0(n372), .S1(
        n369), .Y(n86) );
  MUX41X1_HVT U87 ( .A1(n400), .A3(n349), .A2(n440), .A4(n419), .S0(n356), 
        .S1(n309), .Y(n87) );
  MUX41X1_HVT U88 ( .A1(n412), .A3(n397), .A2(n32), .A4(n48), .S0(n357), .S1(
        n341), .Y(n88) );
  NAND2X0_HVT U89 ( .A1(n326), .A2(n450), .Y(n89) );
  MUX41X1_HVT U90 ( .A1(n279), .A3(n8), .A2(n49), .A4(n89), .S0(n357), .S1(
        n309), .Y(n90) );
  MUX41X1_HVT U95 ( .A1(n94), .A3(n88), .A2(n90), .A4(n87), .S0(n372), .S1(
        n369), .Y(n95) );
  MUX41X1_HVT U96 ( .A1(n435), .A3(n15), .A2(n420), .A4(n441), .S0(n358), .S1(
        n393), .Y(n96) );
  MUX41X1_HVT U98 ( .A1(n97), .A3(n442), .A2(n428), .A4(n30), .S0(n358), .S1(
        n391), .Y(n98) );
  MUX41X1_HVT U99 ( .A1(n34), .A3(n414), .A2(n50), .A4(n375), .S0(n336), .S1(
        n355), .Y(n99) );
  NAND2X0_HVT U100 ( .A1(n326), .A2(n449), .Y(n100) );
  MUX41X1_HVT U101 ( .A1(n443), .A3(n14), .A2(n427), .A4(n100), .S0(n336), 
        .S1(n353), .Y(n101) );
  MUX41X1_HVT U102 ( .A1(n101), .A3(n98), .A2(n99), .A4(n96), .S0(n373), .S1(
        n370), .Y(n102) );
  AND2X1_HVT U104 ( .A1(n8), .A2(n377), .Y(n103) );
  MUX41X1_HVT U105 ( .A1(n16), .A3(n444), .A2(n82), .A4(n103), .S0(n358), .S1(
        n309), .Y(n104) );
  MUX41X1_HVT U108 ( .A1(n416), .A3(n374), .A2(n419), .A4(n382), .S0(n358), 
        .S1(n341), .Y(n107) );
  MUX41X1_HVT U109 ( .A1(n442), .A3(n397), .A2(n439), .A4(n433), .S0(n357), 
        .S1(n341), .Y(n108) );
  MUX41X1_HVT U110 ( .A1(n108), .A3(n106), .A2(n107), .A4(n104), .S0(n373), 
        .S1(n370), .Y(n109) );
  NAND2X0_HVT U114 ( .A1(n277), .A2(n8), .Y(n113) );
  MUX41X1_HVT U115 ( .A1(n113), .A3(n13), .A2(n430), .A4(n379), .S0(n341), 
        .S1(n355), .Y(n114) );
  NAND2X0_HVT U118 ( .A1(n331), .A2(n342), .Y(n117) );
  MUX41X1_HVT U119 ( .A1(n445), .A3(n116), .A2(n39), .A4(n117), .S0(n356), 
        .S1(n341), .Y(n118) );
  MUX41X1_HVT U122 ( .A1(n434), .A3(n346), .A2(n48), .A4(n318), .S0(n356), 
        .S1(n309), .Y(n120) );
  MUX41X1_HVT U124 ( .A1(n348), .A3(n121), .A2(n25), .A4(n332), .S0(n361), 
        .S1(n356), .Y(n122) );
  AOI21X1_HVT U127 ( .A1(n360), .A2(n126), .A3(n404), .Y(n125) );
  NAND2X0_HVT U129 ( .A1(n390), .A2(n1), .Y(n128) );
  MUX41X1_HVT U130 ( .A1(n128), .A3(n127), .A2(n124), .A4(n125), .S0(n362), 
        .S1(n370), .Y(n129) );
  AND2X1_HVT U131 ( .A1(n352), .A2(n331), .Y(n130) );
  MUX41X1_HVT U132 ( .A1(n302), .A3(n130), .A2(n447), .A4(n410), .S0(n336), 
        .S1(n354), .Y(n131) );
  MUX41X1_HVT U133 ( .A1(n448), .A3(n403), .A2(n323), .A4(n402), .S0(n361), 
        .S1(n353), .Y(n132) );
  MUX41X1_HVT U136 ( .A1(n51), .A3(n100), .A2(n134), .A4(n408), .S0(n353), 
        .S1(n310), .Y(n135) );
  MUX41X1_HVT U137 ( .A1(n9), .A3(n31), .A2(n27), .A4(n441), .S0(n362), .S1(
        n353), .Y(n136) );
  MUX41X1_HVT U139 ( .A1(n137), .A3(n133), .A2(n129), .A4(n123), .S0(n373), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n425), .A3(n347), .A2(n418), .A4(n13), .S0(n310), 
        .S1(n355), .Y(n138) );
  NAND2X0_HVT U141 ( .A1(n376), .A2(n326), .Y(n139) );
  MUX41X1_HVT U145 ( .A1(n33), .A3(n444), .A2(n142), .A4(n82), .S0(n360), .S1(
        n309), .Y(n143) );
  OA21X1_HVT U153 ( .A1(n398), .A2(n328), .A3(n407), .Y(n151) );
  MUX41X1_HVT U155 ( .A1(n418), .A3(n13), .A2(n21), .A4(n420), .S0(n359), .S1(
        n310), .Y(n153) );
  MUX41X1_HVT U156 ( .A1(n153), .A3(n149), .A2(n152), .A4(n147), .S0(n373), 
        .S1(n370), .Y(n154) );
  NAND2X0_HVT U159 ( .A1(n157), .A2(n158), .Y(n156) );
  MUX41X1_HVT U162 ( .A1(n304), .A3(n415), .A2(n37), .A4(n160), .S0(n359), 
        .S1(n310), .Y(n161) );
  NAND2X0_HVT U163 ( .A1(n387), .A2(n450), .Y(n162) );
  MUX41X1_HVT U164 ( .A1(n10), .A3(n162), .A2(n39), .A4(n416), .S0(n356), .S1(
        n310), .Y(n163) );
  NAND2X0_HVT U166 ( .A1(n12), .A2(n166), .Y(n165) );
  MUX41X1_HVT U174 ( .A1(n440), .A3(n323), .A2(n448), .A4(n234), .S0(n359), 
        .S1(n393), .Y(n174) );
  NAND2X0_HVT U177 ( .A1(n333), .A2(n342), .Y(n176) );
  MUX41X1_HVT U178 ( .A1(n350), .A3(n176), .A2(n279), .A4(n46), .S0(n359), 
        .S1(n310), .Y(n177) );
  AND2X1_HVT U179 ( .A1(n305), .A2(n377), .Y(n178) );
  MUX41X1_HVT U183 ( .A1(n431), .A3(n329), .A2(n416), .A4(n44), .S0(n361), 
        .S1(n354), .Y(n182) );
  AND2X1_HVT U185 ( .A1(n453), .A2(n331), .Y(n184) );
  OA21X1_HVT U189 ( .A1(n422), .A2(n328), .A3(n62), .Y(n188) );
  NAND2X0_HVT U191 ( .A1(n328), .A2(n409), .Y(n190) );
  AND2X1_HVT U192 ( .A1(n426), .A2(n192), .Y(n191) );
  NAND2X0_HVT U194 ( .A1(n44), .A2(n192), .Y(n194) );
  MUX41X1_HVT U195 ( .A1(n193), .A3(n194), .A2(n191), .A4(n190), .S0(n357), 
        .S1(n369), .Y(n195) );
  NAND2X0_HVT U198 ( .A1(n333), .A2(n234), .Y(n12) );
  NAND2X0_HVT U200 ( .A1(n378), .A2(n326), .Y(n126) );
  AO21X1_HVT U204 ( .A1(n374), .A2(n324), .A3(n328), .Y(n166) );
  AO21X1_HVT U205 ( .A1(n331), .A2(n1), .A3(n328), .Y(n158) );
  NAND2X0_HVT U207 ( .A1(n326), .A2(n279), .Y(n62) );
  MUX21X2_HVT U1 ( .A1(n411), .A2(n420), .S0(n301), .Y(n53) );
  INVX2_HVT U2 ( .A(n330), .Y(n384) );
  INVX0_HVT U3 ( .A(n205), .Y(n436) );
  MUX21X2_HVT U6 ( .A1(n315), .A2(n205), .S0(n317), .Y(n316) );
  INVX1_HVT U14 ( .A(n316), .Y(n187) );
  NAND2X0_HVT U15 ( .A1(n449), .A2(n196), .Y(n197) );
  NAND2X0_HVT U16 ( .A1(n367), .A2(n286), .Y(n198) );
  NAND2X0_HVT U17 ( .A1(n197), .A2(n198), .Y(n28) );
  INVX0_HVT U18 ( .A(n286), .Y(n196) );
  NAND2X0_HVT U20 ( .A1(n175), .A2(n199), .Y(n200) );
  NAND2X0_HVT U21 ( .A1(n168), .A2(n227), .Y(n201) );
  NAND2X0_HVT U22 ( .A1(n200), .A2(n201), .Y(out[6]) );
  INVX1_HVT U23 ( .A(n227), .Y(n199) );
  NBUFFX2_HVT U24 ( .A(n454), .Y(n367) );
  IBUFFX2_HVT U26 ( .A(n333), .Y(n286) );
  MUX21X1_HVT U27 ( .A1(n28), .A2(n25), .S0(n361), .Y(n164) );
  INVX1_HVT U28 ( .A(n272), .Y(n227) );
  MUX21X1_HVT U29 ( .A1(n365), .A2(n367), .S0(n289), .Y(n47) );
  MUX41X1_HVT U30 ( .A1(n188), .A3(n185), .A2(n187), .A4(n186), .S0(n202), 
        .S1(n321), .Y(n189) );
  IBUFFX16_HVT U31 ( .A(n368), .Y(n202) );
  MUX21X2_HVT U33 ( .A1(n102), .A2(n95), .S0(in[7]), .Y(out[2]) );
  MUX21X2_HVT U34 ( .A1(n146), .A2(n145), .S0(n206), .Y(n147) );
  IBUFFX16_HVT U36 ( .A(n355), .Y(n206) );
  IBUFFX2_HVT U37 ( .A(n341), .Y(n246) );
  MUX21X2_HVT U39 ( .A1(n91), .A2(n380), .S0(n386), .Y(n92) );
  NBUFFX4_HVT U40 ( .A(n260), .Y(n383) );
  MUX41X1_HVT U41 ( .A1(n171), .A3(n89), .A2(n24), .A4(n345), .S0(n208), .S1(
        n309), .Y(n172) );
  IBUFFX16_HVT U43 ( .A(n359), .Y(n208) );
  NAND2X0_HVT U44 ( .A1(n416), .A2(n218), .Y(n219) );
  NAND2X0_HVT U45 ( .A1(n65), .A2(n351), .Y(n220) );
  NAND2X0_HVT U46 ( .A1(n219), .A2(n220), .Y(n66) );
  IBUFFX2_HVT U47 ( .A(n351), .Y(n218) );
  NAND2X0_HVT U48 ( .A1(n375), .A2(n221), .Y(n222) );
  NAND2X0_HVT U49 ( .A1(n383), .A2(n385), .Y(n223) );
  NAND2X0_HVT U50 ( .A1(n222), .A2(n223), .Y(n325) );
  IBUFFX2_HVT U51 ( .A(n385), .Y(n221) );
  MUX21X1_HVT U52 ( .A1(n324), .A2(n325), .S0(n321), .Y(n65) );
  INVX0_HVT U54 ( .A(n388), .Y(n385) );
  INVX0_HVT U57 ( .A(n325), .Y(n24) );
  IBUFFX2_HVT U58 ( .A(n394), .Y(n391) );
  IBUFFX2_HVT U59 ( .A(n391), .Y(n297) );
  INVX0_HVT U61 ( .A(n391), .Y(n263) );
  INVX0_HVT U62 ( .A(n391), .Y(n282) );
  MUX41X1_HVT U63 ( .A1(n288), .A3(n436), .A2(n73), .A4(n276), .S0(n354), .S1(
        n341), .Y(n74) );
  NAND2X0_HVT U64 ( .A1(n342), .A2(n224), .Y(n225) );
  NAND2X0_HVT U65 ( .A1(n367), .A2(n271), .Y(n226) );
  NAND2X0_HVT U69 ( .A1(n225), .A2(n226), .Y(n29) );
  INVX0_HVT U70 ( .A(n271), .Y(n224) );
  INVX2_HVT U73 ( .A(n319), .Y(n276) );
  INVX1_HVT U75 ( .A(n240), .Y(n342) );
  IBUFFX2_HVT U76 ( .A(n386), .Y(n271) );
  INVX0_HVT U77 ( .A(n29), .Y(n420) );
  MUX21X2_HVT U86 ( .A1(n278), .A2(n367), .S0(n333), .Y(n171) );
  NAND2X0_HVT U91 ( .A1(n332), .A2(n228), .Y(n229) );
  NAND2X0_HVT U92 ( .A1(n56), .A2(n310), .Y(n230) );
  NAND2X0_HVT U93 ( .A1(n229), .A2(n230), .Y(n60) );
  INVX0_HVT U94 ( .A(n310), .Y(n228) );
  NAND2X0_HVT U97 ( .A1(n61), .A2(n231), .Y(n232) );
  NAND2X0_HVT U103 ( .A1(n60), .A2(n255), .Y(n233) );
  NAND2X0_HVT U106 ( .A1(n232), .A2(n233), .Y(n63) );
  INVX0_HVT U107 ( .A(n255), .Y(n231) );
  MUX21X1_HVT U111 ( .A1(n364), .A2(n382), .S0(n331), .Y(n332) );
  IBUFFX16_HVT U112 ( .A(n394), .Y(n310) );
  IBUFFX2_HVT U113 ( .A(n353), .Y(n255) );
  INVX0_HVT U116 ( .A(n47), .Y(n432) );
  INVX0_HVT U117 ( .A(n28), .Y(n419) );
  INVX0_HVT U120 ( .A(n375), .Y(n234) );
  NAND2X0_HVT U121 ( .A1(n366), .A2(n451), .Y(n237) );
  NAND2X0_HVT U123 ( .A1(n235), .A2(n236), .Y(n238) );
  NAND2X0_HVT U125 ( .A1(n237), .A2(n238), .Y(n18) );
  INVX0_HVT U126 ( .A(n366), .Y(n235) );
  INVX0_HVT U128 ( .A(n451), .Y(n236) );
  INVX0_HVT U134 ( .A(n374), .Y(n453) );
  NBUFFX2_HVT U135 ( .A(n454), .Y(n366) );
  INVX0_HVT U138 ( .A(in[3]), .Y(n451) );
  INVX1_HVT U142 ( .A(n451), .Y(n239) );
  INVX1_HVT U143 ( .A(n239), .Y(n240) );
  NAND2X0_HVT U144 ( .A1(n417), .A2(n241), .Y(n242) );
  NAND2X0_HVT U146 ( .A1(n58), .A2(n351), .Y(n243) );
  NAND2X0_HVT U147 ( .A1(n242), .A2(n243), .Y(n59) );
  INVX0_HVT U148 ( .A(n351), .Y(n241) );
  MUX21X2_HVT U149 ( .A1(n376), .A2(n366), .S0(n244), .Y(n27) );
  IBUFFX16_HVT U150 ( .A(n388), .Y(n244) );
  IBUFFX2_HVT U151 ( .A(n26), .Y(n417) );
  INVX0_HVT U152 ( .A(n41), .Y(n429) );
  MUX41X1_HVT U154 ( .A1(n47), .A3(n178), .A2(n395), .A4(n34), .S0(n245), .S1(
        n246), .Y(n179) );
  IBUFFX16_HVT U157 ( .A(n359), .Y(n245) );
  IBUFFX2_HVT U158 ( .A(n388), .Y(n289) );
  MUX21X1_HVT U160 ( .A1(n374), .A2(n248), .S0(n330), .Y(n247) );
  IBUFFX16_HVT U161 ( .A(n276), .Y(n248) );
  MUX41X1_HVT U165 ( .A1(n148), .A3(n325), .A2(n428), .A4(n438), .S0(n249), 
        .S1(n250), .Y(n149) );
  IBUFFX16_HVT U167 ( .A(n361), .Y(n249) );
  IBUFFX16_HVT U168 ( .A(n353), .Y(n250) );
  IBUFFX2_HVT U169 ( .A(n330), .Y(n320) );
  MUX41X1_HVT U170 ( .A1(n140), .A3(n138), .A2(n143), .A4(n141), .S0(n369), 
        .S1(n251), .Y(n144) );
  IBUFFX16_HVT U171 ( .A(n372), .Y(n251) );
  MUX41X1_HVT U172 ( .A1(n429), .A3(n397), .A2(n294), .A4(n17), .S0(n391), 
        .S1(n356), .Y(n115) );
  NAND2X0_HVT U173 ( .A1(n109), .A2(n252), .Y(n253) );
  NAND2X0_HVT U175 ( .A1(n119), .A2(n311), .Y(n254) );
  NAND2X0_HVT U176 ( .A1(n253), .A2(n254), .Y(out[3]) );
  IBUFFX2_HVT U180 ( .A(n311), .Y(n252) );
  NAND2X2_HVT U181 ( .A1(n376), .A2(n327), .Y(n17) );
  INVX1_HVT U182 ( .A(n385), .Y(n330) );
  INVX0_HVT U184 ( .A(n385), .Y(n331) );
  NAND2X0_HVT U186 ( .A1(n348), .A2(n256), .Y(n257) );
  NAND2X0_HVT U187 ( .A1(n432), .A2(n273), .Y(n258) );
  NAND2X0_HVT U188 ( .A1(n257), .A2(n258), .Y(n193) );
  INVX0_HVT U190 ( .A(n273), .Y(n256) );
  IBUFFX2_HVT U193 ( .A(n361), .Y(n273) );
  MUX21X2_HVT U196 ( .A1(n453), .A2(n365), .S0(n333), .Y(n41) );
  INVX0_HVT U197 ( .A(n2), .Y(n259) );
  INVX1_HVT U199 ( .A(n259), .Y(n260) );
  MUX41X1_HVT U201 ( .A1(n247), .A3(n324), .A2(n400), .A4(n403), .S0(n261), 
        .S1(n275), .Y(n181) );
  IBUFFX16_HVT U202 ( .A(n309), .Y(n261) );
  MUX21X1_HVT U203 ( .A1(n1), .A2(n383), .S0(n327), .Y(n16) );
  IBUFFX2_HVT U206 ( .A(n385), .Y(n326) );
  INVX1_HVT U208 ( .A(n214), .Y(n444) );
  MUX41X1_HVT U209 ( .A1(n418), .A3(n446), .A2(n41), .A4(n139), .S0(n262), 
        .S1(n263), .Y(n140) );
  IBUFFX16_HVT U210 ( .A(n360), .Y(n262) );
  INVX1_HVT U211 ( .A(n247), .Y(n270) );
  INVX1_HVT U212 ( .A(n270), .Y(n438) );
  MUX41X1_HVT U213 ( .A1(n170), .A3(n172), .A2(n173), .A4(n174), .S0(n264), 
        .S1(n265), .Y(n175) );
  IBUFFX16_HVT U214 ( .A(n369), .Y(n264) );
  IBUFFX16_HVT U215 ( .A(n372), .Y(n265) );
  NAND2X0_HVT U216 ( .A1(n54), .A2(n266), .Y(n267) );
  NAND2X0_HVT U217 ( .A1(n53), .A2(n295), .Y(n268) );
  NAND2X0_HVT U218 ( .A1(n267), .A2(n268), .Y(n55) );
  INVX0_HVT U219 ( .A(n295), .Y(n266) );
  IBUFFX2_HVT U220 ( .A(n353), .Y(n295) );
  MUX41X1_HVT U221 ( .A1(n57), .A3(n63), .A2(n55), .A4(n59), .S0(n371), .S1(
        n269), .Y(n64) );
  IBUFFX16_HVT U222 ( .A(n368), .Y(n269) );
  IBUFFX16_HVT U223 ( .A(in[7]), .Y(n272) );
  IBUFFX2_HVT U224 ( .A(n362), .Y(n301) );
  AND2X1_HVT U225 ( .A1(in[3]), .A2(n366), .Y(n274) );
  INVX8_HVT U226 ( .A(n274), .Y(n1) );
  INVX2_HVT U227 ( .A(n274), .Y(n277) );
  INVX0_HVT U228 ( .A(n304), .Y(n46) );
  IBUFFX16_HVT U229 ( .A(n356), .Y(n275) );
  INVX0_HVT U230 ( .A(n364), .Y(n319) );
  IBUFFX2_HVT U231 ( .A(n277), .Y(n278) );
  INVX1_HVT U232 ( .A(n277), .Y(n279) );
  IBUFFX2_HVT U233 ( .A(n277), .Y(n280) );
  NBUFFX2_HVT U234 ( .A(n451), .Y(n363) );
  MUX41X1_HVT U235 ( .A1(n403), .A3(n105), .A2(n379), .A4(n443), .S0(n281), 
        .S1(n282), .Y(n106) );
  IBUFFX16_HVT U236 ( .A(n357), .Y(n281) );
  NAND2X0_HVT U237 ( .A1(n165), .A2(n283), .Y(n284) );
  NAND2X0_HVT U238 ( .A1(n164), .A2(n355), .Y(n285) );
  NAND2X0_HVT U239 ( .A1(n284), .A2(n285), .Y(n167) );
  IBUFFX2_HVT U240 ( .A(n355), .Y(n283) );
  MUX41X1_HVT U241 ( .A1(n180), .A3(n183), .A2(n189), .A4(n195), .S0(n287), 
        .S1(n338), .Y(out[7]) );
  IBUFFX16_HVT U242 ( .A(n373), .Y(n287) );
  INVX0_HVT U243 ( .A(n30), .Y(n421) );
  AO21X2_HVT U244 ( .A1(n362), .A2(n405), .A3(n449), .Y(n146) );
  AO21X1_HVT U245 ( .A1(n387), .A2(n449), .A3(n328), .Y(n192) );
  NBUFFX2_HVT U246 ( .A(n29), .Y(n288) );
  INVX1_HVT U247 ( .A(n388), .Y(n290) );
  NAND2X0_HVT U248 ( .A1(n349), .A2(n291), .Y(n292) );
  NAND2X0_HVT U249 ( .A1(n50), .A2(n362), .Y(n293) );
  NAND2X0_HVT U250 ( .A1(n292), .A2(n293), .Y(n186) );
  IBUFFX2_HVT U251 ( .A(n362), .Y(n291) );
  XOR2X1_HVT U252 ( .A1(n377), .A2(n384), .Y(n50) );
  NBUFFX4_HVT U253 ( .A(n392), .Y(n362) );
  INVX1_HVT U254 ( .A(n31), .Y(n294) );
  MUX41X1_HVT U255 ( .A1(n38), .A3(n382), .A2(n280), .A4(n277), .S0(n296), 
        .S1(n297), .Y(n173) );
  IBUFFX16_HVT U256 ( .A(n359), .Y(n296) );
  INVX1_HVT U257 ( .A(n31), .Y(n422) );
  NAND2X0_HVT U258 ( .A1(n144), .A2(n298), .Y(n299) );
  NAND2X0_HVT U259 ( .A1(n154), .A2(n338), .Y(n300) );
  NAND2X0_HVT U260 ( .A1(n300), .A2(n299), .Y(out[5]) );
  IBUFFX2_HVT U261 ( .A(n338), .Y(n298) );
  NBUFFX2_HVT U262 ( .A(n401), .Y(n302) );
  INVX0_HVT U263 ( .A(n302), .Y(n303) );
  INVX1_HVT U264 ( .A(n216), .Y(n447) );
  MUX21X1_HVT U265 ( .A1(n5), .A2(n418), .S0(n321), .Y(n58) );
  MUX21X1_HVT U266 ( .A1(n377), .A2(n277), .S0(n290), .Y(n304) );
  MUX21X2_HVT U267 ( .A1(n447), .A2(n401), .S0(n361), .Y(n145) );
  INVX1_HVT U268 ( .A(n402), .Y(n305) );
  INVX0_HVT U269 ( .A(n7), .Y(n402) );
  MUX21X2_HVT U270 ( .A1(n376), .A2(n406), .S0(n306), .Y(n93) );
  IBUFFX16_HVT U271 ( .A(n362), .Y(n306) );
  INVX1_HVT U272 ( .A(n315), .Y(n43) );
  MUX21X1_HVT U273 ( .A1(n364), .A2(n452), .S0(n289), .Y(n45) );
  MUX21X1_HVT U274 ( .A1(n452), .A2(n450), .S0(n333), .Y(n116) );
  IBUFFX2_HVT U275 ( .A(n394), .Y(n393) );
  OR2X1_HVT U276 ( .A1(n240), .A2(n454), .Y(n3) );
  IBUFFX2_HVT U277 ( .A(n454), .Y(n352) );
  MUX21X1_HVT U278 ( .A1(n111), .A2(n110), .S0(n360), .Y(n112) );
  MUX41X1_HVT U279 ( .A1(n161), .A3(n167), .A2(n159), .A4(n163), .S0(n307), 
        .S1(n308), .Y(n168) );
  IBUFFX16_HVT U280 ( .A(n373), .Y(n307) );
  IBUFFX16_HVT U281 ( .A(n368), .Y(n308) );
  INVX0_HVT U282 ( .A(n45), .Y(n431) );
  INVX1_HVT U283 ( .A(n388), .Y(n386) );
  MUX21X2_HVT U284 ( .A1(n156), .A2(n155), .S0(n360), .Y(n159) );
  MUX21X2_HVT U285 ( .A1(n318), .A2(n45), .S0(n328), .Y(n155) );
  IBUFFX2_HVT U286 ( .A(n394), .Y(n309) );
  INVX1_HVT U287 ( .A(in[4]), .Y(n394) );
  IBUFFX2_HVT U288 ( .A(n394), .Y(n341) );
  INVX1_HVT U289 ( .A(in[6]), .Y(n454) );
  NBUFFX2_HVT U290 ( .A(n338), .Y(n311) );
  NBUFFX4_HVT U291 ( .A(n392), .Y(n336) );
  INVX2_HVT U292 ( .A(n394), .Y(n392) );
  IBUFFX2_HVT U293 ( .A(n38), .Y(n427) );
  NAND2X0_HVT U294 ( .A1(n181), .A2(n312), .Y(n313) );
  NAND2X0_HVT U295 ( .A1(n182), .A2(n368), .Y(n314) );
  NAND2X0_HVT U296 ( .A1(n313), .A2(n314), .Y(n183) );
  IBUFFX2_HVT U297 ( .A(n368), .Y(n312) );
  INVX0_HVT U298 ( .A(in[7]), .Y(n338) );
  INVX2_HVT U299 ( .A(in[0]), .Y(n388) );
  MUX41X1_HVT U300 ( .A1(n450), .A3(n22), .A2(n431), .A4(n25), .S0(n341), .S1(
        n359), .Y(n141) );
  MUX21X1_HVT U301 ( .A1(n379), .A2(n454), .S0(n388), .Y(n315) );
  IBUFFX16_HVT U302 ( .A(n392), .Y(n317) );
  IBUFFX2_HVT U303 ( .A(n388), .Y(n327) );
  MUX21X1_HVT U304 ( .A1(n379), .A2(n319), .S0(n387), .Y(n318) );
  INVX1_HVT U305 ( .A(n379), .Y(n452) );
  MUX21X1_HVT U306 ( .A1(n404), .A2(n43), .S0(n362), .Y(n110) );
  AO21X1_HVT U307 ( .A1(n430), .A2(n336), .A3(n26), .Y(n111) );
  NAND2X0_HVT U308 ( .A1(n384), .A2(n1), .Y(n7) );
  INVX1_HVT U309 ( .A(in[5]), .Y(n371) );
  INVX1_HVT U310 ( .A(n368), .Y(n369) );
  INVX1_HVT U311 ( .A(n23), .Y(n416) );
  INVX1_HVT U312 ( .A(n392), .Y(n328) );
  INVX0_HVT U313 ( .A(n371), .Y(n373) );
  INVX1_HVT U314 ( .A(n354), .Y(n321) );
  INVX1_HVT U315 ( .A(n368), .Y(n370) );
  INVX1_HVT U316 ( .A(in[1]), .Y(n368) );
  INVX1_HVT U317 ( .A(n388), .Y(n387) );
  INVX0_HVT U318 ( .A(n44), .Y(n403) );
  NBUFFX2_HVT U319 ( .A(n18), .Y(n375) );
  INVX0_HVT U320 ( .A(n400), .Y(n324) );
  MUX21X2_HVT U321 ( .A1(n93), .A2(n92), .S0(n359), .Y(n94) );
  INVX0_HVT U322 ( .A(n56), .Y(n322) );
  INVX0_HVT U323 ( .A(n322), .Y(n323) );
  INVX0_HVT U324 ( .A(n4), .Y(n400) );
  MUX41X1_HVT U325 ( .A1(n66), .A3(n69), .A2(n67), .A4(n70), .S0(n371), .S1(
        n368), .Y(n71) );
  INVX1_HVT U326 ( .A(n371), .Y(n372) );
  MUX41X1_HVT U327 ( .A1(n169), .A3(n348), .A2(n345), .A4(n350), .S0(n337), 
        .S1(n328), .Y(n170) );
  MUX41X1_HVT U328 ( .A1(n112), .A3(n115), .A2(n114), .A4(n118), .S0(n371), 
        .S1(n368), .Y(n119) );
  MUX21X2_HVT U329 ( .A1(n151), .A2(n150), .S0(n360), .Y(n152) );
  MUX21X1_HVT U330 ( .A1(n27), .A2(n349), .S0(n362), .Y(n150) );
  INVX1_HVT U331 ( .A(n27), .Y(n418) );
  INVX1_HVT U332 ( .A(n203), .Y(n329) );
  INVX1_HVT U333 ( .A(n388), .Y(n333) );
  MUX21X2_HVT U334 ( .A1(n184), .A2(n437), .S0(n361), .Y(n185) );
  INVX1_HVT U335 ( .A(n332), .Y(n25) );
  INVX1_HVT U336 ( .A(n207), .Y(n437) );
  OA21X2_HVT U337 ( .A1(n399), .A2(n328), .A3(n23), .Y(n77) );
  MUX21X1_HVT U338 ( .A1(n374), .A2(n364), .S0(n387), .Y(n23) );
  INVX0_HVT U339 ( .A(n358), .Y(n337) );
  MUX21X1_HVT U340 ( .A1(n278), .A2(n452), .S0(n386), .Y(n169) );
  NAND2X0_HVT U341 ( .A1(n79), .A2(in[7]), .Y(n334) );
  NAND2X0_HVT U342 ( .A1(n86), .A2(n311), .Y(n335) );
  NAND2X0_HVT U343 ( .A1(n334), .A2(n335), .Y(out[1]) );
  MUX41X1_HVT U344 ( .A1(n415), .A3(n413), .A2(n40), .A4(n414), .S0(n337), 
        .S1(n391), .Y(n67) );
  NAND2X0_HVT U345 ( .A1(n71), .A2(n311), .Y(n339) );
  NAND2X0_HVT U346 ( .A1(n64), .A2(in[7]), .Y(n340) );
  NAND2X0_HVT U347 ( .A1(n339), .A2(n340), .Y(out[0]) );
  NAND2X0_HVT U348 ( .A1(n179), .A2(n368), .Y(n343) );
  NAND2X0_HVT U349 ( .A1(n177), .A2(n370), .Y(n344) );
  NAND2X0_HVT U350 ( .A1(n344), .A2(n343), .Y(n180) );
  INVX1_HVT U351 ( .A(n382), .Y(n449) );
  NBUFFX2_HVT U352 ( .A(n2), .Y(n382) );
  AND2X1_HVT U353 ( .A1(n7), .A2(n383), .Y(n345) );
  AND2X1_HVT U354 ( .A1(n383), .A2(n17), .Y(n346) );
  MUX21X1_HVT U355 ( .A1(n449), .A2(n453), .S0(n290), .Y(n35) );
  MUX21X1_HVT U356 ( .A1(n367), .A2(n450), .S0(n290), .Y(n148) );
  NAND2X0_HVT U357 ( .A1(n363), .A2(n366), .Y(n2) );
  MUX21X1_HVT U358 ( .A1(n449), .A2(n367), .S0(n327), .Y(n205) );
  MUX21X1_HVT U359 ( .A1(n367), .A2(n453), .S0(n290), .Y(n38) );
  MUX21X1_HVT U360 ( .A1(n449), .A2(n452), .S0(n327), .Y(n52) );
  INVX1_HVT U361 ( .A(n377), .Y(n450) );
  MUX21X1_HVT U362 ( .A1(n278), .A2(n450), .S0(n386), .Y(n30) );
  MUX21X1_HVT U363 ( .A1(n375), .A2(n280), .S0(n333), .Y(n33) );
  MUX21X1_HVT U364 ( .A1(n377), .A2(n380), .S0(n387), .Y(n160) );
  MUX21X1_HVT U365 ( .A1(n382), .A2(n378), .S0(n386), .Y(n142) );
  MUX21X1_HVT U366 ( .A1(n280), .A2(n375), .S0(n320), .Y(n210) );
  MUX21X1_HVT U367 ( .A1(n453), .A2(n367), .S0(n320), .Y(n215) );
  MUX21X1_HVT U368 ( .A1(n377), .A2(n383), .S0(n384), .Y(n216) );
  XNOR2X1_HVT U369 ( .A1(n382), .A2(n384), .Y(n347) );
  MUX21X1_HVT U370 ( .A1(n374), .A2(n450), .S0(n290), .Y(n36) );
  MUX21X1_HVT U371 ( .A1(n364), .A2(n383), .S0(n333), .Y(n207) );
  MUX21X1_HVT U372 ( .A1(n365), .A2(n449), .S0(n290), .Y(n32) );
  MUX21X1_HVT U373 ( .A1(n367), .A2(n260), .S0(n327), .Y(n105) );
  MUX21X1_HVT U374 ( .A1(n381), .A2(n383), .S0(n386), .Y(n20) );
  MUX21X1_HVT U375 ( .A1(n380), .A2(n365), .S0(n327), .Y(n21) );
  XOR2X1_HVT U376 ( .A1(n1), .A2(n384), .Y(n39) );
  MUX21X1_HVT U377 ( .A1(n367), .A2(n375), .S0(n387), .Y(n42) );
  MUX21X1_HVT U378 ( .A1(n35), .A2(n346), .S0(n360), .Y(n127) );
  MUX21X1_HVT U379 ( .A1(n374), .A2(n367), .S0(n392), .Y(n91) );
  MUX21X1_HVT U380 ( .A1(n446), .A2(n347), .S0(n360), .Y(n124) );
  XOR2X1_HVT U381 ( .A1(n379), .A2(n320), .Y(n49) );
  XOR2X1_HVT U382 ( .A1(n376), .A2(n384), .Y(n48) );
  MUX21X1_HVT U383 ( .A1(n276), .A2(n380), .S0(n386), .Y(n213) );
  MUX21X1_HVT U384 ( .A1(n381), .A2(n367), .S0(n387), .Y(n121) );
  NBUFFX2_HVT U385 ( .A(n392), .Y(n361) );
  AND2X1_HVT U386 ( .A1(n386), .A2(n367), .Y(n348) );
  NBUFFX2_HVT U387 ( .A(n451), .Y(n365) );
  NBUFFX2_HVT U388 ( .A(n6), .Y(n377) );
  NBUFFX2_HVT U389 ( .A(n18), .Y(n374) );
  NBUFFX2_HVT U390 ( .A(n18), .Y(n376) );
  AND2X1_HVT U391 ( .A1(n381), .A2(n331), .Y(n349) );
  AND2X1_HVT U392 ( .A1(n452), .A2(n326), .Y(n350) );
  NBUFFX2_HVT U393 ( .A(n6), .Y(n378) );
  NBUFFX2_HVT U394 ( .A(n3), .Y(n379) );
  NBUFFX2_HVT U395 ( .A(n3), .Y(n381) );
  NBUFFX2_HVT U396 ( .A(n3), .Y(n380) );
  MUX21X1_HVT U397 ( .A1(n122), .A2(n120), .S0(n369), .Y(n123) );
  NBUFFX2_HVT U398 ( .A(n240), .Y(n364) );
  MUX21X1_HVT U399 ( .A1(n76), .A2(n77), .S0(n360), .Y(n78) );
  MUX21X1_HVT U400 ( .A1(n318), .A2(n396), .S0(n362), .Y(n76) );
  NBUFFX2_HVT U401 ( .A(n390), .Y(n359) );
  XNOR2X1_HVT U402 ( .A1(n328), .A2(n356), .Y(n351) );
  NBUFFX2_HVT U403 ( .A(n390), .Y(n360) );
  NBUFFX2_HVT U404 ( .A(n389), .Y(n356) );
  NBUFFX2_HVT U405 ( .A(n389), .Y(n355) );
  NBUFFX2_HVT U406 ( .A(n389), .Y(n353) );
  NBUFFX2_HVT U407 ( .A(n389), .Y(n354) );
  NBUFFX2_HVT U408 ( .A(n390), .Y(n357) );
  NBUFFX2_HVT U409 ( .A(n390), .Y(n358) );
  MUX21X1_HVT U410 ( .A1(n280), .A2(n342), .S0(n333), .Y(n217) );
  MUX21X1_HVT U411 ( .A1(n378), .A2(n342), .S0(n289), .Y(n97) );
  MUX21X1_HVT U412 ( .A1(n132), .A2(n131), .S0(n370), .Y(n133) );
  MUX21X1_HVT U413 ( .A1(n136), .A2(n135), .S0(n369), .Y(n137) );
  MUX21X1_HVT U414 ( .A1(n277), .A2(n342), .S0(n320), .Y(n157) );
  MUX21X1_HVT U415 ( .A1(n342), .A2(n378), .S0(n320), .Y(n212) );
  MUX21X1_HVT U416 ( .A1(n342), .A2(n1), .S0(n320), .Y(n211) );
  NBUFFX2_HVT U417 ( .A(in[2]), .Y(n390) );
  NBUFFX2_HVT U418 ( .A(in[2]), .Y(n389) );
  MUX21X1_HVT U419 ( .A1(n276), .A2(n352), .S0(n320), .Y(n214) );
  MUX21X1_HVT U420 ( .A1(n380), .A2(n352), .S0(n289), .Y(n209) );
  MUX21X1_HVT U421 ( .A1(n352), .A2(n381), .S0(n289), .Y(n204) );
  MUX21X1_HVT U422 ( .A1(n352), .A2(n450), .S0(n327), .Y(n203) );
  MUX21X1_HVT U423 ( .A1(n449), .A2(n352), .S0(n289), .Y(n134) );
  XOR2X1_HVT U424 ( .A1(n320), .A2(n352), .Y(n51) );
  MUX21X1_HVT U425 ( .A1(n378), .A2(n352), .S0(n290), .Y(n31) );
  MUX21X1_HVT U426 ( .A1(n352), .A2(n278), .S0(n289), .Y(n26) );
  MUX21X1_HVT U427 ( .A1(n352), .A2(n1), .S0(n387), .Y(n19) );
  INVX0_HVT U428 ( .A(n13), .Y(n395) );
  INVX0_HVT U429 ( .A(n34), .Y(n396) );
  INVX0_HVT U430 ( .A(n40), .Y(n397) );
  INVX0_HVT U431 ( .A(n100), .Y(n398) );
  INVX0_HVT U432 ( .A(n139), .Y(n399) );
  INVX0_HVT U433 ( .A(n5), .Y(n401) );
  INVX0_HVT U434 ( .A(n8), .Y(n404) );
  INVX0_HVT U435 ( .A(n9), .Y(n405) );
  INVX0_HVT U436 ( .A(n37), .Y(n406) );
  INVX0_HVT U437 ( .A(n15), .Y(n407) );
  INVX0_HVT U438 ( .A(n10), .Y(n408) );
  INVX0_HVT U439 ( .A(n14), .Y(n409) );
  INVX0_HVT U440 ( .A(n16), .Y(n410) );
  INVX0_HVT U441 ( .A(n17), .Y(n411) );
  INVX0_HVT U442 ( .A(n19), .Y(n412) );
  INVX0_HVT U443 ( .A(n20), .Y(n413) );
  INVX0_HVT U444 ( .A(n21), .Y(n414) );
  INVX0_HVT U445 ( .A(n22), .Y(n415) );
  INVX0_HVT U446 ( .A(n32), .Y(n423) );
  INVX0_HVT U447 ( .A(n33), .Y(n424) );
  INVX0_HVT U448 ( .A(n35), .Y(n425) );
  INVX0_HVT U449 ( .A(n36), .Y(n426) );
  INVX0_HVT U450 ( .A(n39), .Y(n428) );
  INVX0_HVT U451 ( .A(n42), .Y(n430) );
  INVX0_HVT U452 ( .A(n48), .Y(n433) );
  INVX0_HVT U453 ( .A(n11), .Y(n434) );
  INVX0_HVT U454 ( .A(n204), .Y(n435) );
  INVX0_HVT U455 ( .A(n209), .Y(n439) );
  INVX0_HVT U456 ( .A(n210), .Y(n440) );
  INVX0_HVT U457 ( .A(n211), .Y(n441) );
  INVX0_HVT U458 ( .A(n212), .Y(n442) );
  INVX0_HVT U459 ( .A(n213), .Y(n443) );
  INVX0_HVT U460 ( .A(n157), .Y(n445) );
  INVX0_HVT U461 ( .A(n215), .Y(n446) );
  INVX0_HVT U462 ( .A(n217), .Y(n448) );
endmodule

