
module reg_D_6 ( clk, rst, enable, in, out );
  input [127:0] in;
  output [127:0] out;
  input clk, rst, enable;
  wire   n1, n2, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288;
  tri   clk;
  tri   rst;
  tri   [127:0] in;

  DFFX1_HVT \out_reg[127]  ( .D(n159), .CLK(clk), .Q(out[127]) );
  DFFX1_HVT \out_reg[126]  ( .D(n160), .CLK(clk), .Q(out[126]) );
  DFFX1_HVT \out_reg[125]  ( .D(n161), .CLK(clk), .Q(out[125]) );
  DFFX1_HVT \out_reg[124]  ( .D(n162), .CLK(clk), .Q(out[124]) );
  DFFX1_HVT \out_reg[123]  ( .D(n163), .CLK(clk), .Q(out[123]) );
  DFFX1_HVT \out_reg[122]  ( .D(n164), .CLK(clk), .Q(out[122]) );
  DFFX1_HVT \out_reg[121]  ( .D(n165), .CLK(clk), .Q(out[121]) );
  DFFX1_HVT \out_reg[120]  ( .D(n166), .CLK(clk), .Q(out[120]) );
  DFFX1_HVT \out_reg[119]  ( .D(n167), .CLK(clk), .Q(out[119]) );
  DFFX1_HVT \out_reg[118]  ( .D(n168), .CLK(clk), .Q(out[118]) );
  DFFX1_HVT \out_reg[117]  ( .D(n169), .CLK(clk), .Q(out[117]) );
  DFFX1_HVT \out_reg[116]  ( .D(n170), .CLK(clk), .Q(out[116]) );
  DFFX1_HVT \out_reg[115]  ( .D(n171), .CLK(clk), .Q(out[115]) );
  DFFX1_HVT \out_reg[114]  ( .D(n172), .CLK(clk), .Q(out[114]) );
  DFFX1_HVT \out_reg[113]  ( .D(n173), .CLK(clk), .Q(out[113]) );
  DFFX1_HVT \out_reg[112]  ( .D(n174), .CLK(clk), .Q(out[112]) );
  DFFX1_HVT \out_reg[111]  ( .D(n175), .CLK(clk), .Q(out[111]) );
  DFFX1_HVT \out_reg[110]  ( .D(n176), .CLK(clk), .Q(out[110]) );
  DFFX1_HVT \out_reg[109]  ( .D(n177), .CLK(clk), .Q(out[109]) );
  DFFX1_HVT \out_reg[108]  ( .D(n178), .CLK(clk), .Q(out[108]) );
  DFFX1_HVT \out_reg[107]  ( .D(n179), .CLK(clk), .Q(out[107]) );
  DFFX1_HVT \out_reg[106]  ( .D(n180), .CLK(clk), .Q(out[106]) );
  DFFX1_HVT \out_reg[105]  ( .D(n181), .CLK(clk), .Q(out[105]) );
  DFFX1_HVT \out_reg[104]  ( .D(n182), .CLK(clk), .Q(out[104]) );
  DFFX1_HVT \out_reg[103]  ( .D(n183), .CLK(clk), .Q(out[103]) );
  DFFX1_HVT \out_reg[102]  ( .D(n184), .CLK(clk), .Q(out[102]) );
  DFFX1_HVT \out_reg[101]  ( .D(n185), .CLK(clk), .Q(out[101]) );
  DFFX1_HVT \out_reg[100]  ( .D(n186), .CLK(clk), .Q(out[100]) );
  DFFX1_HVT \out_reg[99]  ( .D(n187), .CLK(clk), .Q(out[99]) );
  DFFX1_HVT \out_reg[98]  ( .D(n188), .CLK(clk), .Q(out[98]) );
  DFFX1_HVT \out_reg[97]  ( .D(n189), .CLK(clk), .Q(out[97]) );
  DFFX1_HVT \out_reg[96]  ( .D(n190), .CLK(clk), .Q(out[96]) );
  DFFX1_HVT \out_reg[95]  ( .D(n191), .CLK(clk), .Q(out[95]) );
  DFFX1_HVT \out_reg[94]  ( .D(n192), .CLK(clk), .Q(out[94]) );
  DFFX1_HVT \out_reg[93]  ( .D(n193), .CLK(clk), .Q(out[93]) );
  DFFX1_HVT \out_reg[92]  ( .D(n194), .CLK(clk), .Q(out[92]) );
  DFFX1_HVT \out_reg[91]  ( .D(n195), .CLK(clk), .Q(out[91]) );
  DFFX1_HVT \out_reg[90]  ( .D(n196), .CLK(clk), .Q(out[90]) );
  DFFX1_HVT \out_reg[89]  ( .D(n197), .CLK(clk), .Q(out[89]) );
  DFFX1_HVT \out_reg[88]  ( .D(n198), .CLK(clk), .Q(out[88]) );
  DFFX1_HVT \out_reg[87]  ( .D(n199), .CLK(clk), .Q(out[87]) );
  DFFX1_HVT \out_reg[86]  ( .D(n200), .CLK(clk), .Q(out[86]) );
  DFFX1_HVT \out_reg[85]  ( .D(n201), .CLK(clk), .Q(out[85]) );
  DFFX1_HVT \out_reg[84]  ( .D(n202), .CLK(clk), .Q(out[84]) );
  DFFX1_HVT \out_reg[83]  ( .D(n203), .CLK(clk), .Q(out[83]) );
  DFFX1_HVT \out_reg[82]  ( .D(n204), .CLK(clk), .Q(out[82]) );
  DFFX1_HVT \out_reg[81]  ( .D(n205), .CLK(clk), .Q(out[81]) );
  DFFX1_HVT \out_reg[80]  ( .D(n206), .CLK(clk), .Q(out[80]) );
  DFFX1_HVT \out_reg[79]  ( .D(n207), .CLK(clk), .Q(out[79]) );
  DFFX1_HVT \out_reg[78]  ( .D(n208), .CLK(clk), .Q(out[78]) );
  DFFX1_HVT \out_reg[77]  ( .D(n209), .CLK(clk), .Q(out[77]) );
  DFFX1_HVT \out_reg[76]  ( .D(n210), .CLK(clk), .Q(out[76]) );
  DFFX1_HVT \out_reg[75]  ( .D(n211), .CLK(clk), .Q(out[75]) );
  DFFX1_HVT \out_reg[74]  ( .D(n212), .CLK(clk), .Q(out[74]) );
  DFFX1_HVT \out_reg[73]  ( .D(n213), .CLK(clk), .Q(out[73]) );
  DFFX1_HVT \out_reg[72]  ( .D(n214), .CLK(clk), .Q(out[72]) );
  DFFX1_HVT \out_reg[71]  ( .D(n215), .CLK(clk), .Q(out[71]) );
  DFFX1_HVT \out_reg[70]  ( .D(n216), .CLK(clk), .Q(out[70]) );
  DFFX1_HVT \out_reg[69]  ( .D(n217), .CLK(clk), .Q(out[69]) );
  DFFX1_HVT \out_reg[68]  ( .D(n218), .CLK(clk), .Q(out[68]) );
  DFFX1_HVT \out_reg[67]  ( .D(n219), .CLK(clk), .Q(out[67]) );
  DFFX1_HVT \out_reg[66]  ( .D(n220), .CLK(clk), .Q(out[66]) );
  DFFX1_HVT \out_reg[65]  ( .D(n221), .CLK(clk), .Q(out[65]) );
  DFFX1_HVT \out_reg[64]  ( .D(n222), .CLK(clk), .Q(out[64]) );
  DFFX1_HVT \out_reg[63]  ( .D(n223), .CLK(clk), .Q(out[63]) );
  DFFX1_HVT \out_reg[62]  ( .D(n224), .CLK(clk), .Q(out[62]) );
  DFFX1_HVT \out_reg[61]  ( .D(n225), .CLK(clk), .Q(out[61]) );
  DFFX1_HVT \out_reg[60]  ( .D(n226), .CLK(clk), .Q(out[60]) );
  DFFX1_HVT \out_reg[59]  ( .D(n227), .CLK(clk), .Q(out[59]) );
  DFFX1_HVT \out_reg[58]  ( .D(n228), .CLK(clk), .Q(out[58]) );
  DFFX1_HVT \out_reg[57]  ( .D(n229), .CLK(clk), .Q(out[57]) );
  DFFX1_HVT \out_reg[56]  ( .D(n230), .CLK(clk), .Q(out[56]) );
  DFFX1_HVT \out_reg[55]  ( .D(n231), .CLK(clk), .Q(out[55]) );
  DFFX1_HVT \out_reg[54]  ( .D(n232), .CLK(clk), .Q(out[54]) );
  DFFX1_HVT \out_reg[53]  ( .D(n233), .CLK(clk), .Q(out[53]) );
  DFFX1_HVT \out_reg[52]  ( .D(n234), .CLK(clk), .Q(out[52]) );
  DFFX1_HVT \out_reg[51]  ( .D(n235), .CLK(clk), .Q(out[51]) );
  DFFX1_HVT \out_reg[50]  ( .D(n236), .CLK(clk), .Q(out[50]) );
  DFFX1_HVT \out_reg[49]  ( .D(n237), .CLK(clk), .Q(out[49]) );
  DFFX1_HVT \out_reg[48]  ( .D(n238), .CLK(clk), .Q(out[48]) );
  DFFX1_HVT \out_reg[47]  ( .D(n239), .CLK(clk), .Q(out[47]) );
  DFFX1_HVT \out_reg[46]  ( .D(n240), .CLK(clk), .Q(out[46]) );
  DFFX1_HVT \out_reg[45]  ( .D(n241), .CLK(clk), .Q(out[45]) );
  DFFX1_HVT \out_reg[44]  ( .D(n242), .CLK(clk), .Q(out[44]) );
  DFFX1_HVT \out_reg[43]  ( .D(n243), .CLK(clk), .Q(out[43]) );
  DFFX1_HVT \out_reg[42]  ( .D(n244), .CLK(clk), .Q(out[42]) );
  DFFX1_HVT \out_reg[41]  ( .D(n245), .CLK(clk), .Q(out[41]) );
  DFFX1_HVT \out_reg[40]  ( .D(n246), .CLK(clk), .Q(out[40]) );
  DFFX1_HVT \out_reg[39]  ( .D(n247), .CLK(clk), .Q(out[39]) );
  DFFX1_HVT \out_reg[38]  ( .D(n248), .CLK(clk), .Q(out[38]) );
  DFFX1_HVT \out_reg[37]  ( .D(n249), .CLK(clk), .Q(out[37]) );
  DFFX1_HVT \out_reg[36]  ( .D(n250), .CLK(clk), .Q(out[36]) );
  DFFX1_HVT \out_reg[35]  ( .D(n251), .CLK(clk), .Q(out[35]) );
  DFFX1_HVT \out_reg[34]  ( .D(n252), .CLK(clk), .Q(out[34]) );
  DFFX1_HVT \out_reg[33]  ( .D(n253), .CLK(clk), .Q(out[33]) );
  DFFX1_HVT \out_reg[32]  ( .D(n254), .CLK(clk), .Q(out[32]) );
  DFFX1_HVT \out_reg[31]  ( .D(n255), .CLK(clk), .Q(out[31]) );
  DFFX1_HVT \out_reg[30]  ( .D(n256), .CLK(clk), .Q(out[30]) );
  DFFX1_HVT \out_reg[29]  ( .D(n257), .CLK(clk), .Q(out[29]) );
  DFFX1_HVT \out_reg[28]  ( .D(n258), .CLK(clk), .Q(out[28]) );
  DFFX1_HVT \out_reg[27]  ( .D(n259), .CLK(clk), .Q(out[27]) );
  DFFX1_HVT \out_reg[26]  ( .D(n260), .CLK(clk), .Q(out[26]) );
  DFFX1_HVT \out_reg[25]  ( .D(n261), .CLK(clk), .Q(out[25]) );
  DFFX1_HVT \out_reg[24]  ( .D(n262), .CLK(clk), .Q(out[24]) );
  DFFX1_HVT \out_reg[23]  ( .D(n263), .CLK(clk), .Q(out[23]) );
  DFFX1_HVT \out_reg[22]  ( .D(n264), .CLK(clk), .Q(out[22]) );
  DFFX1_HVT \out_reg[21]  ( .D(n265), .CLK(clk), .Q(out[21]) );
  DFFX1_HVT \out_reg[20]  ( .D(n266), .CLK(clk), .Q(out[20]) );
  DFFX1_HVT \out_reg[19]  ( .D(n267), .CLK(clk), .Q(out[19]) );
  DFFX1_HVT \out_reg[18]  ( .D(n268), .CLK(clk), .Q(out[18]) );
  DFFX1_HVT \out_reg[17]  ( .D(n269), .CLK(clk), .Q(out[17]) );
  DFFX1_HVT \out_reg[16]  ( .D(n270), .CLK(clk), .Q(out[16]) );
  DFFX1_HVT \out_reg[15]  ( .D(n271), .CLK(clk), .Q(out[15]) );
  DFFX1_HVT \out_reg[14]  ( .D(n272), .CLK(clk), .Q(out[14]) );
  DFFX1_HVT \out_reg[13]  ( .D(n273), .CLK(clk), .Q(out[13]) );
  DFFX1_HVT \out_reg[12]  ( .D(n274), .CLK(clk), .Q(out[12]) );
  DFFX1_HVT \out_reg[11]  ( .D(n275), .CLK(clk), .Q(out[11]) );
  DFFX1_HVT \out_reg[10]  ( .D(n276), .CLK(clk), .Q(out[10]) );
  DFFX1_HVT \out_reg[9]  ( .D(n277), .CLK(clk), .Q(out[9]) );
  DFFX1_HVT \out_reg[8]  ( .D(n278), .CLK(clk), .Q(out[8]) );
  DFFX1_HVT \out_reg[7]  ( .D(n279), .CLK(clk), .Q(out[7]) );
  DFFX1_HVT \out_reg[6]  ( .D(n280), .CLK(clk), .Q(out[6]) );
  DFFX1_HVT \out_reg[5]  ( .D(n281), .CLK(clk), .Q(out[5]) );
  DFFX1_HVT \out_reg[4]  ( .D(n282), .CLK(clk), .Q(out[4]) );
  DFFX1_HVT \out_reg[3]  ( .D(n283), .CLK(clk), .Q(out[3]) );
  DFFX1_HVT \out_reg[2]  ( .D(n284), .CLK(clk), .Q(out[2]) );
  DFFX1_HVT \out_reg[1]  ( .D(n285), .CLK(clk), .Q(out[1]) );
  DFFX1_HVT \out_reg[0]  ( .D(n286), .CLK(clk), .Q(out[0]) );
  AO22X1_HVT U4 ( .A1(out[0]), .A2(n144), .A3(in[0]), .A4(n141), .Y(n286) );
  AO22X1_HVT U5 ( .A1(out[1]), .A2(n144), .A3(in[1]), .A4(n141), .Y(n285) );
  AO22X1_HVT U6 ( .A1(out[2]), .A2(n144), .A3(in[2]), .A4(n141), .Y(n284) );
  AO22X1_HVT U7 ( .A1(out[3]), .A2(n144), .A3(in[3]), .A4(n141), .Y(n283) );
  AO22X1_HVT U8 ( .A1(out[4]), .A2(n144), .A3(in[4]), .A4(n141), .Y(n282) );
  AO22X1_HVT U9 ( .A1(out[5]), .A2(n144), .A3(in[5]), .A4(n141), .Y(n281) );
  AO22X1_HVT U10 ( .A1(out[6]), .A2(n144), .A3(in[6]), .A4(n141), .Y(n280) );
  AO22X1_HVT U11 ( .A1(out[7]), .A2(n144), .A3(in[7]), .A4(n141), .Y(n279) );
  AO22X1_HVT U12 ( .A1(out[8]), .A2(n144), .A3(in[8]), .A4(n140), .Y(n278) );
  AO22X1_HVT U13 ( .A1(out[9]), .A2(n144), .A3(in[9]), .A4(n140), .Y(n277) );
  AO22X1_HVT U14 ( .A1(out[10]), .A2(n144), .A3(in[10]), .A4(n140), .Y(n276)
         );
  AO22X1_HVT U15 ( .A1(out[11]), .A2(n144), .A3(in[11]), .A4(n140), .Y(n275)
         );
  AO22X1_HVT U16 ( .A1(out[12]), .A2(n145), .A3(in[12]), .A4(n140), .Y(n274)
         );
  AO22X1_HVT U17 ( .A1(out[13]), .A2(n145), .A3(in[13]), .A4(n140), .Y(n273)
         );
  AO22X1_HVT U18 ( .A1(out[14]), .A2(n145), .A3(in[14]), .A4(n140), .Y(n272)
         );
  AO22X1_HVT U19 ( .A1(out[15]), .A2(n145), .A3(in[15]), .A4(n140), .Y(n271)
         );
  AO22X1_HVT U20 ( .A1(out[16]), .A2(n145), .A3(in[16]), .A4(n140), .Y(n270)
         );
  AO22X1_HVT U21 ( .A1(out[17]), .A2(n145), .A3(in[17]), .A4(n140), .Y(n269)
         );
  AO22X1_HVT U22 ( .A1(out[18]), .A2(n145), .A3(in[18]), .A4(n140), .Y(n268)
         );
  AO22X1_HVT U23 ( .A1(out[19]), .A2(n145), .A3(in[19]), .A4(n140), .Y(n267)
         );
  AO22X1_HVT U24 ( .A1(out[20]), .A2(n145), .A3(in[20]), .A4(n139), .Y(n266)
         );
  AO22X1_HVT U25 ( .A1(out[21]), .A2(n145), .A3(in[21]), .A4(n139), .Y(n265)
         );
  AO22X1_HVT U26 ( .A1(out[22]), .A2(n145), .A3(in[22]), .A4(n139), .Y(n264)
         );
  AO22X1_HVT U27 ( .A1(out[23]), .A2(n145), .A3(in[23]), .A4(n139), .Y(n263)
         );
  AO22X1_HVT U28 ( .A1(out[24]), .A2(n146), .A3(in[24]), .A4(n139), .Y(n262)
         );
  AO22X1_HVT U29 ( .A1(out[25]), .A2(n146), .A3(in[25]), .A4(n139), .Y(n261)
         );
  AO22X1_HVT U30 ( .A1(out[26]), .A2(n146), .A3(in[26]), .A4(n139), .Y(n260)
         );
  AO22X1_HVT U31 ( .A1(out[27]), .A2(n146), .A3(in[27]), .A4(n139), .Y(n259)
         );
  AO22X1_HVT U32 ( .A1(out[28]), .A2(n146), .A3(in[28]), .A4(n139), .Y(n258)
         );
  AO22X1_HVT U33 ( .A1(out[29]), .A2(n146), .A3(in[29]), .A4(n139), .Y(n257)
         );
  AO22X1_HVT U34 ( .A1(out[30]), .A2(n146), .A3(in[30]), .A4(n139), .Y(n256)
         );
  AO22X1_HVT U35 ( .A1(out[31]), .A2(n146), .A3(in[31]), .A4(n139), .Y(n255)
         );
  AO22X1_HVT U36 ( .A1(out[32]), .A2(n146), .A3(in[32]), .A4(n138), .Y(n254)
         );
  AO22X1_HVT U37 ( .A1(out[33]), .A2(n146), .A3(in[33]), .A4(n138), .Y(n253)
         );
  AO22X1_HVT U38 ( .A1(out[34]), .A2(n146), .A3(in[34]), .A4(n138), .Y(n252)
         );
  AO22X1_HVT U39 ( .A1(out[35]), .A2(n146), .A3(in[35]), .A4(n138), .Y(n251)
         );
  AO22X1_HVT U40 ( .A1(out[36]), .A2(n147), .A3(in[36]), .A4(n138), .Y(n250)
         );
  AO22X1_HVT U41 ( .A1(out[37]), .A2(n147), .A3(in[37]), .A4(n138), .Y(n249)
         );
  AO22X1_HVT U42 ( .A1(out[38]), .A2(n147), .A3(in[38]), .A4(n138), .Y(n248)
         );
  AO22X1_HVT U43 ( .A1(out[39]), .A2(n147), .A3(in[39]), .A4(n138), .Y(n247)
         );
  AO22X1_HVT U44 ( .A1(out[40]), .A2(n147), .A3(in[40]), .A4(n138), .Y(n246)
         );
  AO22X1_HVT U45 ( .A1(out[41]), .A2(n147), .A3(in[41]), .A4(n138), .Y(n245)
         );
  AO22X1_HVT U46 ( .A1(out[42]), .A2(n147), .A3(in[42]), .A4(n138), .Y(n244)
         );
  AO22X1_HVT U47 ( .A1(out[43]), .A2(n147), .A3(in[43]), .A4(n138), .Y(n243)
         );
  AO22X1_HVT U48 ( .A1(out[44]), .A2(n147), .A3(in[44]), .A4(n137), .Y(n242)
         );
  AO22X1_HVT U49 ( .A1(out[45]), .A2(n147), .A3(in[45]), .A4(n137), .Y(n241)
         );
  AO22X1_HVT U50 ( .A1(out[46]), .A2(n147), .A3(in[46]), .A4(n137), .Y(n240)
         );
  AO22X1_HVT U51 ( .A1(out[47]), .A2(n147), .A3(in[47]), .A4(n137), .Y(n239)
         );
  AO22X1_HVT U52 ( .A1(out[48]), .A2(n148), .A3(in[48]), .A4(n137), .Y(n238)
         );
  AO22X1_HVT U53 ( .A1(out[49]), .A2(n148), .A3(in[49]), .A4(n137), .Y(n237)
         );
  AO22X1_HVT U54 ( .A1(out[50]), .A2(n148), .A3(in[50]), .A4(n137), .Y(n236)
         );
  AO22X1_HVT U55 ( .A1(out[51]), .A2(n148), .A3(in[51]), .A4(n137), .Y(n235)
         );
  AO22X1_HVT U56 ( .A1(out[52]), .A2(n148), .A3(in[52]), .A4(n137), .Y(n234)
         );
  AO22X1_HVT U57 ( .A1(out[53]), .A2(n148), .A3(in[53]), .A4(n137), .Y(n233)
         );
  AO22X1_HVT U58 ( .A1(out[54]), .A2(n148), .A3(in[54]), .A4(n137), .Y(n232)
         );
  AO22X1_HVT U59 ( .A1(out[55]), .A2(n148), .A3(in[55]), .A4(n137), .Y(n231)
         );
  AO22X1_HVT U60 ( .A1(out[56]), .A2(n148), .A3(in[56]), .A4(n136), .Y(n230)
         );
  AO22X1_HVT U61 ( .A1(out[57]), .A2(n148), .A3(in[57]), .A4(n136), .Y(n229)
         );
  AO22X1_HVT U62 ( .A1(out[58]), .A2(n148), .A3(in[58]), .A4(n136), .Y(n228)
         );
  AO22X1_HVT U63 ( .A1(out[59]), .A2(n148), .A3(in[59]), .A4(n136), .Y(n227)
         );
  AO22X1_HVT U64 ( .A1(out[60]), .A2(n149), .A3(in[60]), .A4(n136), .Y(n226)
         );
  AO22X1_HVT U65 ( .A1(out[61]), .A2(n149), .A3(in[61]), .A4(n136), .Y(n225)
         );
  AO22X1_HVT U66 ( .A1(out[62]), .A2(n149), .A3(in[62]), .A4(n136), .Y(n224)
         );
  AO22X1_HVT U67 ( .A1(out[63]), .A2(n149), .A3(in[63]), .A4(n136), .Y(n223)
         );
  AO22X1_HVT U68 ( .A1(out[64]), .A2(n149), .A3(in[64]), .A4(n136), .Y(n222)
         );
  AO22X1_HVT U69 ( .A1(out[65]), .A2(n149), .A3(in[65]), .A4(n136), .Y(n221)
         );
  AO22X1_HVT U70 ( .A1(out[66]), .A2(n149), .A3(in[66]), .A4(n136), .Y(n220)
         );
  AO22X1_HVT U71 ( .A1(out[67]), .A2(n149), .A3(in[67]), .A4(n136), .Y(n219)
         );
  AO22X1_HVT U72 ( .A1(out[68]), .A2(n149), .A3(in[68]), .A4(n135), .Y(n218)
         );
  AO22X1_HVT U73 ( .A1(out[69]), .A2(n149), .A3(in[69]), .A4(n135), .Y(n217)
         );
  AO22X1_HVT U74 ( .A1(out[70]), .A2(n149), .A3(in[70]), .A4(n135), .Y(n216)
         );
  AO22X1_HVT U75 ( .A1(out[71]), .A2(n149), .A3(in[71]), .A4(n135), .Y(n215)
         );
  AO22X1_HVT U76 ( .A1(out[72]), .A2(n150), .A3(in[72]), .A4(n135), .Y(n214)
         );
  AO22X1_HVT U77 ( .A1(out[73]), .A2(n150), .A3(in[73]), .A4(n135), .Y(n213)
         );
  AO22X1_HVT U78 ( .A1(out[74]), .A2(n150), .A3(in[74]), .A4(n135), .Y(n212)
         );
  AO22X1_HVT U79 ( .A1(out[75]), .A2(n150), .A3(in[75]), .A4(n135), .Y(n211)
         );
  AO22X1_HVT U80 ( .A1(out[76]), .A2(n150), .A3(in[76]), .A4(n135), .Y(n210)
         );
  AO22X1_HVT U81 ( .A1(out[77]), .A2(n150), .A3(in[77]), .A4(n135), .Y(n209)
         );
  AO22X1_HVT U82 ( .A1(out[78]), .A2(n150), .A3(in[78]), .A4(n135), .Y(n208)
         );
  AO22X1_HVT U83 ( .A1(out[79]), .A2(n150), .A3(in[79]), .A4(n135), .Y(n207)
         );
  AO22X1_HVT U84 ( .A1(out[80]), .A2(n150), .A3(in[80]), .A4(n134), .Y(n206)
         );
  AO22X1_HVT U85 ( .A1(out[81]), .A2(n150), .A3(in[81]), .A4(n134), .Y(n205)
         );
  AO22X1_HVT U86 ( .A1(out[82]), .A2(n150), .A3(in[82]), .A4(n134), .Y(n204)
         );
  AO22X1_HVT U87 ( .A1(out[83]), .A2(n150), .A3(in[83]), .A4(n134), .Y(n203)
         );
  AO22X1_HVT U88 ( .A1(out[84]), .A2(n151), .A3(in[84]), .A4(n134), .Y(n202)
         );
  AO22X1_HVT U89 ( .A1(out[85]), .A2(n151), .A3(in[85]), .A4(n134), .Y(n201)
         );
  AO22X1_HVT U90 ( .A1(out[86]), .A2(n151), .A3(in[86]), .A4(n134), .Y(n200)
         );
  AO22X1_HVT U91 ( .A1(out[87]), .A2(n151), .A3(in[87]), .A4(n134), .Y(n199)
         );
  AO22X1_HVT U92 ( .A1(out[88]), .A2(n151), .A3(in[88]), .A4(n134), .Y(n198)
         );
  AO22X1_HVT U93 ( .A1(out[89]), .A2(n151), .A3(in[89]), .A4(n134), .Y(n197)
         );
  AO22X1_HVT U94 ( .A1(out[90]), .A2(n151), .A3(in[90]), .A4(n134), .Y(n196)
         );
  AO22X1_HVT U95 ( .A1(out[91]), .A2(n151), .A3(in[91]), .A4(n134), .Y(n195)
         );
  AO22X1_HVT U96 ( .A1(out[92]), .A2(n151), .A3(in[92]), .A4(n133), .Y(n194)
         );
  AO22X1_HVT U97 ( .A1(out[93]), .A2(n151), .A3(in[93]), .A4(n133), .Y(n193)
         );
  AO22X1_HVT U98 ( .A1(out[94]), .A2(n151), .A3(in[94]), .A4(n133), .Y(n192)
         );
  AO22X1_HVT U99 ( .A1(out[95]), .A2(n151), .A3(in[95]), .A4(n133), .Y(n191)
         );
  AO22X1_HVT U100 ( .A1(out[96]), .A2(n152), .A3(in[96]), .A4(n133), .Y(n190)
         );
  AO22X1_HVT U101 ( .A1(out[97]), .A2(n152), .A3(in[97]), .A4(n133), .Y(n189)
         );
  AO22X1_HVT U102 ( .A1(out[98]), .A2(n152), .A3(in[98]), .A4(n133), .Y(n188)
         );
  AO22X1_HVT U103 ( .A1(out[99]), .A2(n152), .A3(in[99]), .A4(n133), .Y(n187)
         );
  AO22X1_HVT U104 ( .A1(out[100]), .A2(n152), .A3(in[100]), .A4(n133), .Y(n186) );
  AO22X1_HVT U105 ( .A1(out[101]), .A2(n152), .A3(in[101]), .A4(n133), .Y(n185) );
  AO22X1_HVT U106 ( .A1(out[102]), .A2(n152), .A3(in[102]), .A4(n133), .Y(n184) );
  AO22X1_HVT U107 ( .A1(out[103]), .A2(n152), .A3(in[103]), .A4(n133), .Y(n183) );
  AO22X1_HVT U108 ( .A1(out[104]), .A2(n152), .A3(in[104]), .A4(n2), .Y(n182)
         );
  AO22X1_HVT U109 ( .A1(out[105]), .A2(n152), .A3(in[105]), .A4(n2), .Y(n181)
         );
  AO22X1_HVT U110 ( .A1(out[106]), .A2(n152), .A3(in[106]), .A4(n2), .Y(n180)
         );
  AO22X1_HVT U111 ( .A1(out[107]), .A2(n152), .A3(in[107]), .A4(n2), .Y(n179)
         );
  AO22X1_HVT U112 ( .A1(out[108]), .A2(n153), .A3(in[108]), .A4(n2), .Y(n178)
         );
  AO22X1_HVT U113 ( .A1(out[109]), .A2(n153), .A3(in[109]), .A4(n2), .Y(n177)
         );
  AO22X1_HVT U114 ( .A1(out[110]), .A2(n153), .A3(in[110]), .A4(n2), .Y(n176)
         );
  AO22X1_HVT U115 ( .A1(out[111]), .A2(n153), .A3(in[111]), .A4(n2), .Y(n175)
         );
  AO22X1_HVT U116 ( .A1(out[112]), .A2(n153), .A3(in[112]), .A4(n2), .Y(n174)
         );
  AO22X1_HVT U117 ( .A1(out[113]), .A2(n153), .A3(in[113]), .A4(n2), .Y(n173)
         );
  AO22X1_HVT U118 ( .A1(out[114]), .A2(n153), .A3(in[114]), .A4(n2), .Y(n172)
         );
  AO22X1_HVT U119 ( .A1(out[115]), .A2(n153), .A3(in[115]), .A4(n2), .Y(n171)
         );
  AO22X1_HVT U120 ( .A1(out[116]), .A2(n153), .A3(in[116]), .A4(n1), .Y(n170)
         );
  AO22X1_HVT U121 ( .A1(out[117]), .A2(n153), .A3(in[117]), .A4(n1), .Y(n169)
         );
  AO22X1_HVT U122 ( .A1(out[118]), .A2(n153), .A3(in[118]), .A4(n1), .Y(n168)
         );
  AO22X1_HVT U123 ( .A1(out[119]), .A2(n153), .A3(in[119]), .A4(n1), .Y(n167)
         );
  AO22X1_HVT U124 ( .A1(out[120]), .A2(n154), .A3(in[120]), .A4(n1), .Y(n166)
         );
  AO22X1_HVT U125 ( .A1(out[121]), .A2(n154), .A3(in[121]), .A4(n1), .Y(n165)
         );
  AO22X1_HVT U126 ( .A1(out[122]), .A2(n154), .A3(in[122]), .A4(n1), .Y(n164)
         );
  AO22X1_HVT U127 ( .A1(out[123]), .A2(n154), .A3(in[123]), .A4(n1), .Y(n163)
         );
  AO22X1_HVT U128 ( .A1(out[124]), .A2(n154), .A3(in[124]), .A4(n1), .Y(n162)
         );
  AO22X1_HVT U129 ( .A1(out[125]), .A2(n154), .A3(in[125]), .A4(n1), .Y(n161)
         );
  AO22X1_HVT U130 ( .A1(out[126]), .A2(n154), .A3(in[126]), .A4(n1), .Y(n160)
         );
  AO22X1_HVT U131 ( .A1(out[127]), .A2(n154), .A3(in[127]), .A4(n1), .Y(n159)
         );
  AND2X1_HVT U132 ( .A1(n158), .A2(n287), .Y(n288) );
  NAND2X0_HVT U133 ( .A1(enable), .A2(n158), .Y(n287) );
  INVX1_HVT U2 ( .A(n142), .Y(n139) );
  INVX1_HVT U3 ( .A(n142), .Y(n138) );
  INVX1_HVT U134 ( .A(n142), .Y(n137) );
  INVX1_HVT U135 ( .A(n142), .Y(n136) );
  INVX1_HVT U136 ( .A(n143), .Y(n134) );
  INVX1_HVT U137 ( .A(n143), .Y(n133) );
  INVX1_HVT U138 ( .A(n143), .Y(n2) );
  INVX1_HVT U139 ( .A(n143), .Y(n1) );
  INVX1_HVT U140 ( .A(n142), .Y(n140) );
  INVX1_HVT U141 ( .A(n142), .Y(n141) );
  INVX1_HVT U142 ( .A(n143), .Y(n135) );
  INVX1_HVT U143 ( .A(n157), .Y(n142) );
  INVX0_HVT U144 ( .A(n157), .Y(n143) );
  INVX1_HVT U145 ( .A(n156), .Y(n144) );
  INVX1_HVT U146 ( .A(n156), .Y(n145) );
  INVX1_HVT U147 ( .A(n156), .Y(n146) );
  INVX1_HVT U148 ( .A(n156), .Y(n147) );
  INVX1_HVT U149 ( .A(n155), .Y(n149) );
  INVX1_HVT U150 ( .A(n155), .Y(n150) );
  INVX1_HVT U151 ( .A(n155), .Y(n151) );
  INVX1_HVT U152 ( .A(n155), .Y(n152) );
  INVX1_HVT U153 ( .A(n155), .Y(n154) );
  INVX1_HVT U154 ( .A(n155), .Y(n153) );
  INVX1_HVT U155 ( .A(n156), .Y(n148) );
  INVX1_HVT U156 ( .A(n288), .Y(n155) );
  INVX0_HVT U157 ( .A(n288), .Y(n156) );
  INVX0_HVT U158 ( .A(n287), .Y(n157) );
  INVX0_HVT U159 ( .A(rst), .Y(n158) );
endmodule

