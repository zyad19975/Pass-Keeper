
module sbox_12 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n7, n8, n23, n28, n50, n51, n118, n119, n210, n211, n212, n213, n214,
         n216, n217, n218, n219, n227, n229, n230, n231, n232, n235, n236,
         n238, n241, n242, n245, n246, n249, n252, n253, n254, n261, n264,
         n269, n272, n275, n279, n280, n282, n283, n286, n289, n292, n293,
         n297, n299, n300, n301, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786;

  NAND2X0_HVT U4 ( .A1(n517), .A2(n784), .Y(n783) );
  NAND2X0_HVT U5 ( .A1(n523), .A2(n515), .Y(n781) );
  NAND2X0_HVT U13 ( .A1(n775), .A2(n313), .Y(n776) );
  NAND2X0_HVT U21 ( .A1(n517), .A2(n526), .Y(n767) );
  NAND2X0_HVT U24 ( .A1(n335), .A2(n474), .Y(n765) );
  NAND2X0_HVT U33 ( .A1(n365), .A2(n526), .Y(n757) );
  NAND2X0_HVT U35 ( .A1(n513), .A2(n526), .Y(n755) );
  NAND2X0_HVT U42 ( .A1(n406), .A2(n335), .Y(n748) );
  MUX41X1_HVT U51 ( .A1(n539), .A3(n560), .A2(n333), .A4(n540), .S0(n487), 
        .S1(n529), .Y(n741) );
  NAND2X0_HVT U53 ( .A1(n738), .A2(n747), .Y(n739) );
  NAND2X0_HVT U56 ( .A1(n517), .A2(n734), .Y(n735) );
  MUX41X1_HVT U57 ( .A1(n548), .A3(n769), .A2(n735), .A4(n778), .S0(n487), 
        .S1(n506), .Y(n733) );
  NAND2X0_HVT U58 ( .A1(n522), .A2(n396), .Y(n732) );
  MUX41X1_HVT U59 ( .A1(n498), .A3(n732), .A2(n496), .A4(n551), .S0(n488), 
        .S1(n529), .Y(n731) );
  MUX41X1_HVT U61 ( .A1(n494), .A3(n383), .A2(n544), .A4(n471), .S0(n488), 
        .S1(n506), .Y(n729) );
  NAND2X0_HVT U62 ( .A1(n474), .A2(n520), .Y(n728) );
  MUX41X1_HVT U63 ( .A1(n728), .A3(n542), .A2(n317), .A4(n541), .S0(n488), 
        .S1(n529), .Y(n727) );
  MUX41X1_HVT U68 ( .A1(n388), .A3(n724), .A2(n723), .A4(n725), .S0(n390), 
        .S1(n487), .Y(n722) );
  NAND2X0_HVT U73 ( .A1(n329), .A2(n717), .Y(n718) );
  MUX41X1_HVT U77 ( .A1(n780), .A3(n557), .A2(n714), .A4(n547), .S0(n508), 
        .S1(n376), .Y(n713) );
  AND2X1_HVT U83 ( .A1(n393), .A2(n449), .Y(n706) );
  MUX41X1_HVT U84 ( .A1(n545), .A3(n468), .A2(n772), .A4(n706), .S0(n390), 
        .S1(n532), .Y(n705) );
  NAND2X0_HVT U85 ( .A1(n526), .A2(n572), .Y(n704) );
  MUX41X1_HVT U90 ( .A1(n744), .A3(n748), .A2(n539), .A4(n701), .S0(n501), 
        .S1(n532), .Y(n700) );
  MUX41X1_HVT U97 ( .A1(n570), .A3(n493), .A2(n393), .A4(n773), .S0(n503), 
        .S1(n213), .Y(n692) );
  NAND2X0_HVT U101 ( .A1(n687), .A2(n686), .Y(n688) );
  MUX41X1_HVT U103 ( .A1(n396), .A3(n562), .A2(n448), .A4(n755), .S0(n390), 
        .S1(n532), .Y(n684) );
  MUX41X1_HVT U105 ( .A1(n567), .A3(n742), .A2(n683), .A4(n559), .S0(n390), 
        .S1(n485), .Y(n682) );
  NAND2X0_HVT U110 ( .A1(n519), .A2(n677), .Y(n678) );
  AND2X1_HVT U115 ( .A1(n218), .A2(n473), .Y(n674) );
  MUX41X1_HVT U116 ( .A1(n372), .A3(n674), .A2(n438), .A4(n759), .S0(n501), 
        .S1(n213), .Y(n673) );
  MUX41X1_HVT U136 ( .A1(n491), .A3(n757), .A2(n538), .A4(n754), .S0(n501), 
        .S1(n489), .Y(n652) );
  AND2X1_HVT U140 ( .A1(n331), .A2(n526), .Y(n648) );
  AND2X1_HVT U154 ( .A1(n510), .A2(n424), .Y(n635) );
  NAND2X0_HVT U158 ( .A1(n406), .A2(n572), .Y(n631) );
  MUX41X1_HVT U159 ( .A1(n372), .A3(n473), .A2(n631), .A4(n574), .S0(n501), 
        .S1(n213), .Y(n630) );
  AND2X1_HVT U162 ( .A1(n467), .A2(n238), .Y(n627) );
  MUX41X1_HVT U163 ( .A1(n383), .A3(n627), .A2(n492), .A4(n628), .S0(n241), 
        .S1(n532), .Y(n626) );
  MUX41X1_HVT U165 ( .A1(n767), .A3(n566), .A2(n744), .A4(n625), .S0(n487), 
        .S1(n241), .Y(n624) );
  NAND2X0_HVT U166 ( .A1(n521), .A2(n734), .Y(n623) );
  NAND2X0_HVT U167 ( .A1(n537), .A2(n526), .Y(n622) );
  MUX41X1_HVT U168 ( .A1(n548), .A3(n330), .A2(n622), .A4(n623), .S0(n373), 
        .S1(n311), .Y(n621) );
  NAND2X0_HVT U174 ( .A1(n391), .A2(n468), .Y(n775) );
  NAND2X0_HVT U177 ( .A1(n391), .A2(n513), .Y(n614) );
  MUX41X1_HVT U180 ( .A1(n543), .A3(n780), .A2(n372), .A4(n490), .S0(n508), 
        .S1(n376), .Y(n611) );
  MUX41X1_HVT U182 ( .A1(n554), .A3(n517), .A2(n8), .A4(n563), .S0(n487), .S1(
        n376), .Y(n609) );
  MUX41X1_HVT U189 ( .A1(n603), .A3(n775), .A2(n604), .A4(n559), .S0(n508), 
        .S1(n504), .Y(n602) );
  AO21X1_HVT U197 ( .A1(n495), .A2(n311), .A3(n568), .Y(n595) );
  NAND2X0_HVT U208 ( .A1(n384), .A2(n517), .Y(n677) );
  NAND2X0_HVT U215 ( .A1(n677), .A2(n330), .Y(n585) );
  NAND2X0_HVT U218 ( .A1(n435), .A2(n392), .Y(n638) );
  NAND2X0_HVT U220 ( .A1(n311), .A2(n348), .Y(n709) );
  INVX0_HVT U241 ( .A(n765), .Y(n576) );
  INVX0_HVT U242 ( .A(n748), .Y(n575) );
  INVX0_HVT U245 ( .A(n781), .Y(n574) );
  INVX0_HVT U256 ( .A(n638), .Y(n568) );
  INVX0_HVT U264 ( .A(n755), .Y(n564) );
  INVX0_HVT U265 ( .A(n763), .Y(n563) );
  INVX0_HVT U268 ( .A(n767), .Y(n560) );
  INVX0_HVT U270 ( .A(n585), .Y(n559) );
  INVX0_HVT U284 ( .A(n348), .Y(n549) );
  INVX0_HVT U296 ( .A(n773), .Y(n542) );
  INVX0_HVT U306 ( .A(n622), .Y(n536) );
  MUX21X1_HVT U1 ( .A1(n289), .A2(n486), .S0(n436), .Y(n760) );
  NBUFFX2_HVT U2 ( .A(n316), .Y(n513) );
  NBUFFX2_HVT U3 ( .A(n409), .Y(n521) );
  INVX1_HVT U6 ( .A(n472), .Y(n471) );
  AO21X1_HVT U7 ( .A1(n503), .A2(n330), .A3(n468), .Y(n671) );
  INVX1_HVT U8 ( .A(n356), .Y(n750) );
  MUX21X1_HVT U9 ( .A1(n435), .A2(n537), .S0(n218), .Y(n625) );
  NBUFFX2_HVT U10 ( .A(n445), .Y(n384) );
  NBUFFX2_HVT U11 ( .A(n565), .Y(n512) );
  MUX21X1_HVT U12 ( .A1(n571), .A2(n774), .S0(n376), .Y(n690) );
  AND3X1_HVT U14 ( .A1(n527), .A2(n474), .A3(n326), .Y(n659) );
  MUX21X1_HVT U15 ( .A1(n607), .A2(n608), .S0(n504), .Y(n606) );
  AOI21X1_HVT U16 ( .A1(n423), .A2(n480), .A3(n766), .Y(n607) );
  INVX1_HVT U17 ( .A(n506), .Y(n454) );
  AND2X1_HVT U18 ( .A1(n431), .A2(n432), .Y(n7) );
  AND2X1_HVT U19 ( .A1(n362), .A2(n363), .Y(n8) );
  XNOR2X1_HVT U20 ( .A1(n500), .A2(n436), .Y(n23) );
  AND2X1_HVT U22 ( .A1(n380), .A2(n408), .Y(n28) );
  INVX1_HVT U23 ( .A(n784), .Y(n286) );
  INVX1_HVT U25 ( .A(n480), .Y(n484) );
  INVX1_HVT U26 ( .A(n534), .Y(n485) );
  INVX1_HVT U27 ( .A(n762), .Y(n567) );
  INVX0_HVT U28 ( .A(n407), .Y(n280) );
  INVX1_HVT U29 ( .A(n519), .Y(n537) );
  MUX21X2_HVT U30 ( .A1(n470), .A2(n365), .S0(n392), .Y(n694) );
  NAND2X0_HVT U31 ( .A1(n663), .A2(n505), .Y(n50) );
  NAND2X0_HVT U32 ( .A1(n662), .A2(n531), .Y(n51) );
  NAND2X0_HVT U34 ( .A1(n50), .A2(n51), .Y(n661) );
  AOI21X1_HVT U36 ( .A1(n388), .A2(n489), .A3(n752), .Y(n591) );
  MUX21X1_HVT U37 ( .A1(n521), .A2(n469), .S0(n389), .Y(n388) );
  MUX41X1_HVT U38 ( .A1(n305), .A3(n423), .A2(n776), .A4(n735), .S0(n377), 
        .S1(n458), .Y(n588) );
  NAND2X0_HVT U39 ( .A1(n313), .A2(n118), .Y(n119) );
  NAND2X0_HVT U40 ( .A1(n520), .A2(n436), .Y(n210) );
  NAND2X0_HVT U41 ( .A1(n119), .A2(n210), .Y(n604) );
  INVX0_HVT U43 ( .A(n405), .Y(n118) );
  MUX21X2_HVT U44 ( .A1(n331), .A2(n471), .S0(n391), .Y(n683) );
  INVX1_HVT U45 ( .A(n28), .Y(n467) );
  INVX1_HVT U46 ( .A(n383), .Y(n771) );
  INVX0_HVT U47 ( .A(n475), .Y(n445) );
  INVX1_HVT U48 ( .A(n480), .Y(n534) );
  MUX21X1_HVT U49 ( .A1(n335), .A2(n521), .S0(n384), .Y(n334) );
  MUX21X1_HVT U50 ( .A1(n289), .A2(n323), .S0(n433), .Y(n333) );
  INVX1_HVT U52 ( .A(n757), .Y(n553) );
  INVX1_HVT U54 ( .A(n502), .Y(n318) );
  INVX1_HVT U55 ( .A(n402), .Y(n475) );
  AND3X1_HVT U60 ( .A1(n323), .A2(n734), .A3(n709), .Y(n710) );
  INVX1_HVT U64 ( .A(n332), .Y(n699) );
  XOR2X1_HVT U65 ( .A1(n528), .A2(n489), .Y(n743) );
  INVX1_HVT U66 ( .A(n337), .Y(n672) );
  NBUFFX2_HVT U67 ( .A(n527), .Y(n502) );
  MUX21X1_HVT U69 ( .A1(n435), .A2(n578), .S0(n269), .Y(n434) );
  INVX1_HVT U70 ( .A(n502), .Y(n443) );
  OA21X1_HVT U71 ( .A1(n536), .A2(n484), .A3(n759), .Y(n644) );
  INVX1_HVT U72 ( .A(n282), .Y(n572) );
  MUX21X1_HVT U74 ( .A1(n572), .A2(n471), .S0(n436), .Y(n628) );
  INVX1_HVT U75 ( .A(n321), .Y(n311) );
  INVX1_HVT U76 ( .A(n760), .Y(n566) );
  INVX1_HVT U78 ( .A(n485), .Y(n321) );
  MUX21X1_HVT U79 ( .A1(n424), .A2(n704), .S0(n484), .Y(n608) );
  INVX1_HVT U80 ( .A(n499), .Y(n376) );
  INVX1_HVT U81 ( .A(n573), .Y(n238) );
  NBUFFX2_HVT U82 ( .A(n527), .Y(n390) );
  NAND2X0_HVT U86 ( .A1(n739), .A2(n484), .Y(n446) );
  INVX1_HVT U87 ( .A(n333), .Y(n769) );
  INVX1_HVT U88 ( .A(n503), .Y(n279) );
  OA21X1_HVT U89 ( .A1(n750), .A2(n481), .A3(n638), .Y(n639) );
  INVX1_HVT U91 ( .A(n443), .Y(n214) );
  INVX1_HVT U92 ( .A(n511), .Y(n283) );
  INVX1_HVT U93 ( .A(n504), .Y(n415) );
  INVX1_HVT U94 ( .A(n504), .Y(n377) );
  NBUFFX2_HVT U95 ( .A(n533), .Y(n508) );
  NBUFFX2_HVT U96 ( .A(n530), .Y(n507) );
  INVX0_HVT U98 ( .A(n779), .Y(n328) );
  INVX0_HVT U99 ( .A(n328), .Y(n331) );
  NBUFFX2_HVT U100 ( .A(n533), .Y(n510) );
  NBUFFX2_HVT U102 ( .A(n530), .Y(n506) );
  INVX1_HVT U104 ( .A(n323), .Y(n500) );
  INVX1_HVT U106 ( .A(in[6]), .Y(n385) );
  INVX1_HVT U107 ( .A(n322), .Y(n424) );
  INVX1_HVT U108 ( .A(n346), .Y(n752) );
  INVX0_HVT U109 ( .A(n766), .Y(n545) );
  AND2X1_HVT U111 ( .A1(n440), .A2(n441), .Y(n211) );
  INVX0_HVT U112 ( .A(n438), .Y(n764) );
  INVX1_HVT U113 ( .A(n522), .Y(n312) );
  INVX0_HVT U114 ( .A(n516), .Y(n435) );
  MUX21X1_HVT U117 ( .A1(n329), .A2(n512), .S0(n523), .Y(n719) );
  NBUFFX2_HVT U118 ( .A(n445), .Y(n393) );
  MUX41X1_HVT U119 ( .A1(n654), .A3(n652), .A2(n653), .A4(n650), .S0(n453), 
        .S1(n454), .Y(n649) );
  NBUFFX2_HVT U120 ( .A(n464), .Y(n212) );
  INVX0_HVT U121 ( .A(n777), .Y(n561) );
  INVX1_HVT U122 ( .A(n359), .Y(n241) );
  INVX1_HVT U123 ( .A(n469), .Y(n470) );
  MUX41X1_HVT U124 ( .A1(n599), .A3(n597), .A2(n598), .A4(n594), .S0(n453), 
        .S1(n454), .Y(n593) );
  INVX0_HVT U125 ( .A(n476), .Y(n526) );
  NBUFFX2_HVT U126 ( .A(n485), .Y(n213) );
  MUX41X1_HVT U127 ( .A1(n771), .A3(n614), .A2(n444), .A4(n752), .S0(n214), 
        .S1(n485), .Y(n613) );
  MUX21X2_HVT U128 ( .A1(n522), .A2(n486), .S0(n405), .Y(n762) );
  INVX1_HVT U129 ( .A(n556), .Y(n364) );
  INVX0_HVT U130 ( .A(n525), .Y(n218) );
  INVX0_HVT U131 ( .A(n475), .Y(n406) );
  MUX21X2_HVT U132 ( .A1(n512), .A2(n312), .S0(n445), .Y(n439) );
  MUX41X1_HVT U133 ( .A1(n512), .A3(n616), .A2(n546), .A4(n775), .S0(n487), 
        .S1(n528), .Y(n615) );
  MUX41X1_HVT U134 ( .A1(n388), .A3(n555), .A2(n767), .A4(n498), .S0(n501), 
        .S1(n269), .Y(n662) );
  INVX0_HVT U135 ( .A(n455), .Y(n754) );
  MUX21X1_HVT U137 ( .A1(n518), .A2(n330), .S0(n212), .Y(n701) );
  INVX1_HVT U138 ( .A(n475), .Y(n524) );
  MUX21X1_HVT U139 ( .A1(n515), .A2(n518), .S0(n353), .Y(n777) );
  MUX21X1_HVT U141 ( .A1(n518), .A2(n313), .S0(n523), .Y(n696) );
  MUX41X1_HVT U142 ( .A1(n438), .A3(n569), .A2(n500), .A4(n570), .S0(n481), 
        .S1(n443), .Y(n715) );
  NAND2X0_HVT U143 ( .A1(n461), .A2(n435), .Y(n216) );
  NAND2X0_HVT U144 ( .A1(n218), .A2(n331), .Y(n217) );
  NAND2X0_HVT U145 ( .A1(n216), .A2(n217), .Y(n745) );
  INVX1_HVT U146 ( .A(n509), .Y(n458) );
  INVX0_HVT U147 ( .A(n325), .Y(n326) );
  INVX0_HVT U148 ( .A(n525), .Y(n405) );
  INVX1_HVT U149 ( .A(n402), .Y(n525) );
  INVX1_HVT U150 ( .A(n512), .Y(n486) );
  XNOR2X1_HVT U151 ( .A1(n405), .A2(n289), .Y(n742) );
  MUX41X1_HVT U152 ( .A1(n600), .A3(n755), .A2(n23), .A4(n748), .S0(n458), 
        .S1(n318), .Y(n599) );
  INVX1_HVT U153 ( .A(n768), .Y(n540) );
  MUX21X1_HVT U155 ( .A1(n515), .A2(n329), .S0(n433), .Y(n582) );
  NAND2X0_HVT U156 ( .A1(n280), .A2(n514), .Y(n219) );
  MUX21X1_HVT U157 ( .A1(n466), .A2(n515), .S0(n392), .Y(n772) );
  INVX1_HVT U160 ( .A(n477), .Y(n392) );
  INVX0_HVT U161 ( .A(n334), .Y(n778) );
  MUX21X1_HVT U164 ( .A1(n219), .A2(n465), .S0(n525), .Y(n438) );
  MUX21X1_HVT U169 ( .A1(n516), .A2(n219), .S0(n389), .Y(n774) );
  NAND2X0_HVT U170 ( .A1(n567), .A2(n279), .Y(n227) );
  NAND2X0_HVT U171 ( .A1(n760), .A2(n502), .Y(n229) );
  NAND2X0_HVT U172 ( .A1(n227), .A2(n229), .Y(n660) );
  INVX1_HVT U173 ( .A(in[1]), .Y(n477) );
  INVX0_HVT U175 ( .A(n772), .Y(n544) );
  MUX41X1_HVT U176 ( .A1(n749), .A3(n378), .A2(n7), .A4(n331), .S0(n508), .S1(
        n376), .Y(n598) );
  INVX0_HVT U178 ( .A(n394), .Y(n230) );
  INVX1_HVT U179 ( .A(in[3]), .Y(n394) );
  INVX0_HVT U181 ( .A(n582), .Y(n231) );
  MUX41X1_HVT U183 ( .A1(n602), .A3(n606), .A2(n605), .A4(n609), .S0(n511), 
        .S1(n506), .Y(n601) );
  MUX41X1_HVT U184 ( .A1(n751), .A3(n744), .A2(n493), .A4(n238), .S0(n487), 
        .S1(n318), .Y(n605) );
  MUX21X1_HVT U185 ( .A1(n556), .A2(n335), .S0(n525), .Y(n751) );
  XOR2X1_HVT U186 ( .A1(n518), .A2(n353), .Y(n492) );
  NAND2X0_HVT U187 ( .A1(n666), .A2(n510), .Y(n232) );
  NAND2X0_HVT U188 ( .A1(n667), .A2(n481), .Y(n235) );
  NAND2X0_HVT U190 ( .A1(n232), .A2(n235), .Y(n663) );
  MUX21X2_HVT U191 ( .A1(n585), .A2(n760), .S0(n321), .Y(n579) );
  MUX21X2_HVT U192 ( .A1(n396), .A2(n455), .S0(n359), .Y(n680) );
  INVX0_HVT U193 ( .A(n286), .Y(n396) );
  NAND2X0_HVT U194 ( .A1(n334), .A2(n507), .Y(n236) );
  NAND2X0_HVT U195 ( .A1(n236), .A2(n238), .Y(n724) );
  NBUFFX2_HVT U196 ( .A(n533), .Y(n487) );
  NBUFFX2_HVT U198 ( .A(n533), .Y(n488) );
  NBUFFX2_HVT U199 ( .A(n533), .Y(n489) );
  MUX41X1_HVT U200 ( .A1(n549), .A3(n444), .A2(n762), .A4(n439), .S0(n241), 
        .S1(n321), .Y(n612) );
  NAND2X0_HVT U201 ( .A1(n761), .A2(n401), .Y(n425) );
  INVX0_HVT U202 ( .A(n780), .Y(n562) );
  MUX41X1_HVT U203 ( .A1(n569), .A3(n704), .A2(n495), .A4(n491), .S0(n214), 
        .S1(n532), .Y(n703) );
  AO21X1_HVT U204 ( .A1(n510), .A2(n696), .A3(n568), .Y(n697) );
  INVX1_HVT U205 ( .A(n696), .Y(n557) );
  INVX1_HVT U206 ( .A(n324), .Y(n316) );
  MUX21X1_HVT U207 ( .A1(n562), .A2(n435), .S0(n507), .Y(n723) );
  XOR2X2_HVT U209 ( .A1(n513), .A2(n212), .Y(n763) );
  MUX41X1_HVT U210 ( .A1(n589), .A3(n590), .A2(n587), .A4(n588), .S0(n505), 
        .S1(n453), .Y(n586) );
  INVX0_HVT U211 ( .A(n352), .Y(n465) );
  MUX41X1_HVT U212 ( .A1(n346), .A3(n552), .A2(n764), .A4(n648), .S0(n488), 
        .S1(n443), .Y(n647) );
  INVX0_HVT U213 ( .A(n558), .Y(n242) );
  INVX1_HVT U214 ( .A(n583), .Y(n548) );
  INVX0_HVT U216 ( .A(n477), .Y(n523) );
  NAND2X0_HVT U217 ( .A1(n591), .A2(n279), .Y(n245) );
  NAND2X0_HVT U219 ( .A1(n592), .A2(n504), .Y(n246) );
  NAND2X0_HVT U221 ( .A1(n245), .A2(n246), .Y(n590) );
  MUX41X1_HVT U222 ( .A1(n719), .A3(n718), .A2(n763), .A4(n765), .S0(n487), 
        .S1(n503), .Y(n716) );
  MUX41X1_HVT U223 ( .A1(n777), .A3(n758), .A2(n754), .A4(n356), .S0(n376), 
        .S1(n458), .Y(n589) );
  NAND2X0_HVT U224 ( .A1(n771), .A2(n279), .Y(n249) );
  NAND2X0_HVT U225 ( .A1(n552), .A2(n501), .Y(n252) );
  NAND2X0_HVT U226 ( .A1(n249), .A2(n252), .Y(n657) );
  NBUFFX2_HVT U227 ( .A(n527), .Y(n501) );
  NAND2X0_HVT U228 ( .A1(n571), .A2(n528), .Y(n253) );
  NAND2X0_HVT U229 ( .A1(n439), .A2(n318), .Y(n254) );
  NAND2X0_HVT U230 ( .A1(n253), .A2(n254), .Y(n483) );
  MUX21X1_HVT U231 ( .A1(n482), .A2(n483), .S0(n532), .Y(n587) );
  INVX0_HVT U232 ( .A(n261), .Y(n482) );
  INVX1_HVT U233 ( .A(n464), .Y(n353) );
  MUX21X1_HVT U234 ( .A1(n513), .A2(n286), .S0(n528), .Y(n261) );
  INVX0_HVT U235 ( .A(n485), .Y(n401) );
  NAND2X0_HVT U236 ( .A1(n486), .A2(n406), .Y(n264) );
  NAND2X0_HVT U237 ( .A1(n264), .A2(n299), .Y(n758) );
  INVX0_HVT U238 ( .A(n758), .Y(n552) );
  INVX1_HVT U239 ( .A(n489), .Y(n269) );
  INVX1_HVT U240 ( .A(in[4]), .Y(n325) );
  INVX1_HVT U243 ( .A(n325), .Y(n324) );
  OA21X1_HVT U244 ( .A1(n496), .A2(n401), .A3(n759), .Y(n619) );
  MUX21X1_HVT U246 ( .A1(n282), .A2(n516), .S0(n464), .Y(n759) );
  INVX0_HVT U247 ( .A(n379), .Y(n282) );
  NAND2X0_HVT U248 ( .A1(n620), .A2(n279), .Y(n272) );
  NAND2X0_HVT U249 ( .A1(n619), .A2(n214), .Y(n275) );
  NAND2X0_HVT U250 ( .A1(n272), .A2(n275), .Y(n618) );
  MUX41X1_HVT U251 ( .A1(n494), .A3(n678), .A2(n564), .A4(n519), .S0(n279), 
        .S1(n213), .Y(n636) );
  MUX21X1_HVT U252 ( .A1(n494), .A2(n690), .S0(n743), .Y(n689) );
  INVX1_HVT U253 ( .A(n466), .Y(n472) );
  INVX1_HVT U254 ( .A(n584), .Y(n539) );
  OR2X1_HVT U255 ( .A1(n461), .A2(n328), .Y(n734) );
  INVX0_HVT U257 ( .A(n782), .Y(n556) );
  INVX0_HVT U258 ( .A(n477), .Y(n464) );
  MUX21X1_HVT U259 ( .A1(n512), .A2(n521), .S0(n476), .Y(n455) );
  INVX1_HVT U260 ( .A(n452), .Y(n407) );
  MUX41X1_HVT U261 ( .A1(n661), .A3(n675), .A2(n656), .A4(n669), .S0(in[6]), 
        .S1(n283), .Y(out[3]) );
  INVX1_HVT U262 ( .A(n477), .Y(n476) );
  NBUFFX2_HVT U263 ( .A(n322), .Y(n289) );
  NBUFFX2_HVT U266 ( .A(n322), .Y(n515) );
  INVX0_HVT U267 ( .A(n452), .Y(n322) );
  INVX0_HVT U269 ( .A(n352), .Y(n466) );
  INVX1_HVT U271 ( .A(n534), .Y(n532) );
  NAND2X0_HVT U272 ( .A1(n330), .A2(n508), .Y(n292) );
  NAND2X0_HVT U273 ( .A1(n768), .A2(n481), .Y(n293) );
  NAND2X0_HVT U274 ( .A1(n292), .A2(n293), .Y(n711) );
  INVX0_HVT U275 ( .A(n328), .Y(n330) );
  INVX0_HVT U276 ( .A(n510), .Y(n481) );
  INVX0_HVT U277 ( .A(n476), .Y(n461) );
  NAND2X0_HVT U278 ( .A1(n512), .A2(n406), .Y(n297) );
  NAND2X0_HVT U279 ( .A1(n556), .A2(n433), .Y(n299) );
  NAND2X0_HVT U280 ( .A1(n297), .A2(n299), .Y(n578) );
  NBUFFX2_HVT U281 ( .A(n524), .Y(n436) );
  INVX0_HVT U282 ( .A(n477), .Y(n391) );
  NAND2X0_HVT U283 ( .A1(n575), .A2(n269), .Y(n300) );
  NAND2X0_HVT U285 ( .A1(n444), .A2(n509), .Y(n301) );
  NAND2X0_HVT U286 ( .A1(n300), .A2(n301), .Y(n596) );
  NBUFFX2_HVT U287 ( .A(n533), .Y(n509) );
  INVX1_HVT U288 ( .A(n322), .Y(n335) );
  INVX1_HVT U289 ( .A(n394), .Y(n452) );
  NAND2X0_HVT U290 ( .A1(n639), .A2(n377), .Y(n303) );
  NAND2X0_HVT U291 ( .A1(n640), .A2(n214), .Y(n304) );
  NAND2X0_HVT U292 ( .A1(n303), .A2(n304), .Y(n637) );
  MUX21X1_HVT U293 ( .A1(n547), .A2(n327), .S0(n509), .Y(n640) );
  NAND2X0_HVT U294 ( .A1(n354), .A2(n355), .Y(n305) );
  MUX41X1_HVT U295 ( .A1(n545), .A3(n558), .A2(n470), .A4(n329), .S0(n488), 
        .S1(n501), .Y(n646) );
  INVX0_HVT U297 ( .A(n328), .Y(n329) );
  NAND2X0_HVT U298 ( .A1(n331), .A2(n401), .Y(n306) );
  NAND2X0_HVT U299 ( .A1(n231), .A2(n510), .Y(n307) );
  NAND2X0_HVT U300 ( .A1(n306), .A2(n307), .Y(n620) );
  INVX0_HVT U301 ( .A(n465), .Y(n468) );
  INVX1_HVT U302 ( .A(n336), .Y(n308) );
  INVX1_HVT U303 ( .A(n466), .Y(n336) );
  INVX1_HVT U304 ( .A(n28), .Y(n469) );
  MUX41X1_HVT U305 ( .A1(n613), .A3(n615), .A2(n611), .A4(n612), .S0(n505), 
        .S1(n453), .Y(n610) );
  INVX0_HVT U307 ( .A(n448), .Y(n761) );
  INVX0_HVT U308 ( .A(n336), .Y(n473) );
  INVX0_HVT U309 ( .A(n524), .Y(n389) );
  INVX0_HVT U310 ( .A(n785), .Y(n309) );
  INVX1_HVT U311 ( .A(n309), .Y(n310) );
  INVX0_HVT U312 ( .A(n734), .Y(n570) );
  INVX1_HVT U313 ( .A(n499), .Y(n527) );
  MUX21X1_HVT U314 ( .A1(n517), .A2(n449), .S0(n118), .Y(n448) );
  MUX21X1_HVT U315 ( .A1(n280), .A2(n518), .S0(n389), .Y(n780) );
  NBUFFX2_HVT U316 ( .A(n380), .Y(n313) );
  MUX41X1_HVT U317 ( .A1(n744), .A3(n238), .A2(n570), .A4(n538), .S0(n321), 
        .S1(n359), .Y(n642) );
  NAND2X0_HVT U318 ( .A1(n673), .A2(n505), .Y(n314) );
  NAND2X0_HVT U319 ( .A1(n670), .A2(n454), .Y(n315) );
  NAND2X0_HVT U320 ( .A1(n314), .A2(n315), .Y(n669) );
  NBUFFX2_HVT U321 ( .A(n565), .Y(n514) );
  INVX0_HVT U322 ( .A(n717), .Y(n573) );
  NAND2X0_HVT U323 ( .A1(n218), .A2(n521), .Y(n717) );
  NBUFFX2_HVT U324 ( .A(n380), .Y(n522) );
  INVX1_HVT U325 ( .A(n524), .Y(n433) );
  AND2X1_HVT U326 ( .A1(n775), .A2(n313), .Y(n317) );
  NAND2X0_HVT U327 ( .A1(n553), .A2(n318), .Y(n319) );
  NAND2X0_HVT U328 ( .A1(n668), .A2(n502), .Y(n320) );
  NAND2X0_HVT U329 ( .A1(n319), .A2(n320), .Y(n667) );
  MUX21X1_HVT U330 ( .A1(n519), .A2(n699), .S0(n497), .Y(n698) );
  MUX21X1_HVT U331 ( .A1(n310), .A2(n486), .S0(n353), .Y(n768) );
  XNOR2X1_HVT U332 ( .A1(n484), .A2(n406), .Y(n497) );
  INVX0_HVT U333 ( .A(n513), .Y(n449) );
  NAND2X0_HVT U334 ( .A1(n280), .A2(n514), .Y(n323) );
  INVX1_HVT U335 ( .A(in[2]), .Y(n499) );
  INVX1_HVT U336 ( .A(n581), .Y(n569) );
  NBUFFX2_HVT U337 ( .A(in[1]), .Y(n402) );
  INVX1_HVT U338 ( .A(n516), .Y(n327) );
  XNOR2X2_HVT U339 ( .A1(n308), .A2(n523), .Y(n744) );
  NAND2X0_HVT U340 ( .A1(n421), .A2(n420), .Y(out[6]) );
  MUX21X1_HVT U341 ( .A1(n486), .A2(n289), .S0(n484), .Y(n332) );
  INVX0_HVT U342 ( .A(n395), .Y(n668) );
  INVX0_HVT U343 ( .A(n686), .Y(n546) );
  MUX21X1_HVT U344 ( .A1(n756), .A2(n755), .S0(n415), .Y(n337) );
  INVX0_HVT U345 ( .A(n759), .Y(n571) );
  NAND2X0_HVT U346 ( .A1(n492), .A2(n279), .Y(n338) );
  NAND2X0_HVT U347 ( .A1(n544), .A2(n390), .Y(n339) );
  NAND2X0_HVT U348 ( .A1(n338), .A2(n339), .Y(n658) );
  OR2X1_HVT U349 ( .A1(n286), .A2(n336), .Y(n773) );
  INVX0_HVT U350 ( .A(n774), .Y(n541) );
  NAND2X0_HVT U351 ( .A1(n313), .A2(n433), .Y(n340) );
  NAND2X0_HVT U352 ( .A1(n424), .A2(n391), .Y(n341) );
  NAND2X0_HVT U353 ( .A1(n340), .A2(n341), .Y(n423) );
  NAND2X0_HVT U354 ( .A1(n517), .A2(n461), .Y(n342) );
  NAND2X0_HVT U355 ( .A1(n468), .A2(n392), .Y(n343) );
  NAND2X0_HVT U356 ( .A1(n342), .A2(n343), .Y(n753) );
  NAND2X0_HVT U357 ( .A1(n641), .A2(n385), .Y(n344) );
  NAND2X0_HVT U358 ( .A1(n649), .A2(in[6]), .Y(n345) );
  NAND2X0_HVT U359 ( .A1(n344), .A2(n345), .Y(out[4]) );
  AND2X1_HVT U360 ( .A1(n366), .A2(n367), .Y(n346) );
  INVX0_HVT U361 ( .A(n677), .Y(n558) );
  XNOR2X1_HVT U362 ( .A1(n347), .A2(n484), .Y(n746) );
  AND2X1_HVT U363 ( .A1(n381), .A2(n382), .Y(n347) );
  OA21X1_HVT U364 ( .A1(n550), .A2(n318), .A3(n551), .Y(n679) );
  INVX0_HVT U365 ( .A(n753), .Y(n550) );
  NAND2X0_HVT U366 ( .A1(n468), .A2(n474), .Y(n348) );
  NAND2X0_HVT U367 ( .A1(n513), .A2(n218), .Y(n349) );
  NAND2X0_HVT U368 ( .A1(n348), .A2(n349), .Y(n714) );
  INVX1_HVT U369 ( .A(n437), .Y(n442) );
  NAND2X0_HVT U370 ( .A1(n561), .A2(n531), .Y(n350) );
  NAND2X0_HVT U371 ( .A1(n474), .A2(n507), .Y(n351) );
  NAND2X0_HVT U372 ( .A1(n350), .A2(n351), .Y(n725) );
  INVX0_HVT U373 ( .A(n392), .Y(n474) );
  NAND2X0_HVT U374 ( .A1(n408), .A2(n409), .Y(n352) );
  INVX1_HVT U375 ( .A(n577), .Y(n538) );
  NAND2X0_HVT U376 ( .A1(n470), .A2(n353), .Y(n354) );
  NAND2X0_HVT U377 ( .A1(n424), .A2(n392), .Y(n355) );
  NAND2X0_HVT U378 ( .A1(n355), .A2(n354), .Y(n766) );
  NAND2X0_HVT U379 ( .A1(n721), .A2(n241), .Y(n429) );
  MUX21X1_HVT U380 ( .A1(n230), .A2(n310), .S0(n476), .Y(n356) );
  NAND2X0_HVT U381 ( .A1(n365), .A2(n118), .Y(n357) );
  NAND2X0_HVT U382 ( .A1(n500), .A2(n393), .Y(n358) );
  NAND2X0_HVT U383 ( .A1(n357), .A2(n358), .Y(n616) );
  NAND2X0_HVT U384 ( .A1(n374), .A2(n375), .Y(n594) );
  MUX41X1_HVT U385 ( .A1(n642), .A3(n646), .A2(n643), .A4(n647), .S0(n511), 
        .S1(n505), .Y(n641) );
  NAND2X0_HVT U386 ( .A1(n759), .A2(n359), .Y(n360) );
  NAND2X0_HVT U387 ( .A1(n678), .A2(n502), .Y(n361) );
  NAND2X0_HVT U388 ( .A1(n360), .A2(n361), .Y(n676) );
  INVX0_HVT U389 ( .A(n502), .Y(n359) );
  INVX1_HVT U390 ( .A(n499), .Y(n528) );
  MUX41X1_HVT U391 ( .A1(n722), .A3(n726), .A2(n730), .A4(n736), .S0(n511), 
        .S1(in[6]), .Y(out[0]) );
  NAND2X0_HVT U392 ( .A1(n519), .A2(n433), .Y(n362) );
  NAND2X0_HVT U393 ( .A1(n473), .A2(n436), .Y(n363) );
  NAND2X0_HVT U394 ( .A1(n362), .A2(n363), .Y(n749) );
  MUX41X1_HVT U395 ( .A1(n576), .A3(n745), .A2(n774), .A4(n540), .S0(n401), 
        .S1(n390), .Y(n707) );
  INVX1_HVT U396 ( .A(n364), .Y(n365) );
  NAND2X0_HVT U397 ( .A1(n572), .A2(n526), .Y(n366) );
  NAND2X0_HVT U398 ( .A1(n556), .A2(n406), .Y(n367) );
  NAND2X0_HVT U399 ( .A1(n665), .A2(n664), .Y(n666) );
  NAND2X0_HVT U400 ( .A1(n655), .A2(n241), .Y(n368) );
  NAND2X0_HVT U401 ( .A1(n535), .A2(n377), .Y(n369) );
  NAND2X0_HVT U402 ( .A1(n369), .A2(n368), .Y(n654) );
  NAND2X0_HVT U403 ( .A1(n783), .A2(n373), .Y(n370) );
  NAND2X0_HVT U404 ( .A1(n651), .A2(n377), .Y(n371) );
  NAND2X0_HVT U405 ( .A1(n370), .A2(n371), .Y(n650) );
  INVX1_HVT U406 ( .A(n317), .Y(n372) );
  MUX41X1_HVT U407 ( .A1(n659), .A3(n657), .A2(n660), .A4(n658), .S0(n454), 
        .S1(n488), .Y(n656) );
  NAND2X0_HVT U408 ( .A1(n595), .A2(n373), .Y(n374) );
  NAND2X0_HVT U409 ( .A1(n596), .A2(n415), .Y(n375) );
  INVX0_HVT U410 ( .A(n415), .Y(n373) );
  NAND2X0_HVT U411 ( .A1(n381), .A2(n382), .Y(n378) );
  INVX0_HVT U412 ( .A(n786), .Y(n379) );
  INVX1_HVT U413 ( .A(n379), .Y(n380) );
  NAND2X0_HVT U414 ( .A1(n500), .A2(n461), .Y(n381) );
  NAND2X0_HVT U415 ( .A1(n572), .A2(n523), .Y(n382) );
  OR2X1_HVT U416 ( .A1(n481), .A2(n751), .Y(n478) );
  INVX0_HVT U417 ( .A(n751), .Y(n554) );
  INVX1_HVT U418 ( .A(n534), .Y(n533) );
  MUX41X1_HVT U419 ( .A1(n713), .A3(n716), .A2(n715), .A4(n720), .S0(n511), 
        .S1(n530), .Y(n712) );
  MUX21X1_HVT U420 ( .A1(n512), .A2(n329), .S0(n405), .Y(n383) );
  MUX41X1_HVT U421 ( .A1(n632), .A3(n637), .A2(n630), .A4(n636), .S0(in[0]), 
        .S1(n454), .Y(n629) );
  NAND2X0_HVT U422 ( .A1(n681), .A2(n385), .Y(n386) );
  NAND2X0_HVT U423 ( .A1(n691), .A2(in[6]), .Y(n387) );
  NAND2X0_HVT U424 ( .A1(n386), .A2(n387), .Y(out[2]) );
  MUX41X1_HVT U425 ( .A1(n703), .A3(n707), .A2(n705), .A4(n708), .S0(n511), 
        .S1(n505), .Y(n702) );
  MUX41X1_HVT U426 ( .A1(n689), .A3(n685), .A2(n684), .A4(n682), .S0(n454), 
        .S1(n453), .Y(n681) );
  MUX41X1_HVT U427 ( .A1(n624), .A3(n618), .A2(n626), .A4(n621), .S0(n453), 
        .S1(n505), .Y(n617) );
  NBUFFX2_HVT U428 ( .A(n527), .Y(n503) );
  INVX1_HVT U429 ( .A(n580), .Y(n547) );
  MUX21X1_HVT U430 ( .A1(n424), .A2(n449), .S0(n353), .Y(n395) );
  MUX41X1_HVT U431 ( .A1(n680), .A3(n211), .A2(n679), .A4(n676), .S0(n454), 
        .S1(n488), .Y(n675) );
  NAND2X0_HVT U432 ( .A1(n391), .A2(n310), .Y(n784) );
  NAND2X0_HVT U433 ( .A1(n772), .A2(n458), .Y(n397) );
  NAND2X0_HVT U434 ( .A1(n490), .A2(n508), .Y(n398) );
  NAND2X0_HVT U435 ( .A1(n397), .A2(n398), .Y(n592) );
  NAND2X0_HVT U436 ( .A1(n710), .A2(n214), .Y(n399) );
  NAND2X0_HVT U437 ( .A1(n711), .A2(n279), .Y(n400) );
  NAND2X0_HVT U438 ( .A1(n400), .A2(n399), .Y(n708) );
  MUX41X1_HVT U439 ( .A1(n694), .A3(n231), .A2(n493), .A4(n576), .S0(n318), 
        .S1(n401), .Y(n693) );
  INVX1_HVT U440 ( .A(n410), .Y(n444) );
  INVX0_HVT U441 ( .A(n783), .Y(n543) );
  MUX41X1_HVT U442 ( .A1(n695), .A3(n700), .A2(n692), .A4(n693), .S0(n505), 
        .S1(n453), .Y(n691) );
  NAND2X0_HVT U443 ( .A1(n697), .A2(n279), .Y(n403) );
  NAND2X0_HVT U444 ( .A1(n698), .A2(n214), .Y(n404) );
  NAND2X0_HVT U445 ( .A1(n404), .A2(n403), .Y(n695) );
  INVX1_HVT U446 ( .A(n511), .Y(n453) );
  NAND2X0_HVT U447 ( .A1(n407), .A2(n565), .Y(n408) );
  NAND2X0_HVT U448 ( .A1(n326), .A2(n452), .Y(n409) );
  MUX21X1_HVT U449 ( .A1(n449), .A2(n330), .S0(n392), .Y(n410) );
  NAND2X0_HVT U450 ( .A1(n634), .A2(n373), .Y(n411) );
  NAND2X0_HVT U451 ( .A1(n633), .A2(n377), .Y(n412) );
  NAND2X0_HVT U452 ( .A1(n411), .A2(n412), .Y(n632) );
  MUX21X1_HVT U453 ( .A1(n752), .A2(n557), .S0(n508), .Y(n633) );
  NAND2X0_HVT U454 ( .A1(n741), .A2(n241), .Y(n413) );
  NAND2X0_HVT U455 ( .A1(n737), .A2(n377), .Y(n414) );
  NAND2X0_HVT U456 ( .A1(n413), .A2(n414), .Y(n736) );
  MUX41X1_HVT U457 ( .A1(n231), .A3(n467), .A2(n753), .A4(n282), .S0(n279), 
        .S1(n480), .Y(n597) );
  INVX0_HVT U458 ( .A(n423), .Y(n756) );
  NAND2X0_HVT U459 ( .A1(n727), .A2(n377), .Y(n416) );
  NAND2X0_HVT U460 ( .A1(n729), .A2(n504), .Y(n417) );
  NAND2X0_HVT U461 ( .A1(n416), .A2(n417), .Y(n726) );
  NAND2X0_HVT U462 ( .A1(n645), .A2(n377), .Y(n418) );
  NAND2X0_HVT U463 ( .A1(n644), .A2(n214), .Y(n419) );
  NAND2X0_HVT U464 ( .A1(n418), .A2(n419), .Y(n643) );
  NAND2X0_HVT U465 ( .A1(n601), .A2(n385), .Y(n420) );
  NAND2X0_HVT U466 ( .A1(n610), .A2(in[6]), .Y(n421) );
  INVX0_HVT U467 ( .A(n578), .Y(n555) );
  MUX21X1_HVT U468 ( .A1(n515), .A2(n514), .S0(n502), .Y(n422) );
  NAND2X0_HVT U469 ( .A1(n286), .A2(n510), .Y(n426) );
  NAND2X0_HVT U470 ( .A1(n425), .A2(n426), .Y(n645) );
  NAND2X0_HVT U471 ( .A1(n586), .A2(n385), .Y(n427) );
  NAND2X0_HVT U472 ( .A1(n593), .A2(in[6]), .Y(n428) );
  NAND2X0_HVT U473 ( .A1(n427), .A2(n428), .Y(out[7]) );
  NAND2X0_HVT U474 ( .A1(n746), .A2(n415), .Y(n430) );
  NAND2X0_HVT U475 ( .A1(n429), .A2(n430), .Y(n720) );
  MUX21X1_HVT U476 ( .A1(n572), .A2(n231), .S0(n510), .Y(n721) );
  MUX41X1_HVT U477 ( .A1(n781), .A3(n7), .A2(n378), .A4(n327), .S0(n401), .S1(
        n503), .Y(n653) );
  NAND2X0_HVT U478 ( .A1(n467), .A2(n433), .Y(n431) );
  NAND2X0_HVT U479 ( .A1(n435), .A2(n393), .Y(n432) );
  INVX0_HVT U480 ( .A(n434), .Y(n655) );
  XOR2X1_HVT U481 ( .A1(n476), .A2(n499), .Y(n437) );
  NAND2X0_HVT U482 ( .A1(n422), .A2(n437), .Y(n440) );
  NAND2X0_HVT U483 ( .A1(n537), .A2(n442), .Y(n441) );
  INVX1_HVT U484 ( .A(n324), .Y(n565) );
  NAND2X0_HVT U485 ( .A1(n740), .A2(n508), .Y(n447) );
  NAND2X0_HVT U486 ( .A1(n446), .A2(n447), .Y(n737) );
  MUX21X1_HVT U487 ( .A1(n335), .A2(n755), .S0(n507), .Y(n740) );
  INVX1_HVT U488 ( .A(n579), .Y(n535) );
  MUX21X1_HVT U489 ( .A1(n635), .A2(n520), .S0(n497), .Y(n634) );
  NAND2X0_HVT U490 ( .A1(n731), .A2(n415), .Y(n450) );
  NAND2X0_HVT U491 ( .A1(n733), .A2(n241), .Y(n451) );
  NAND2X0_HVT U492 ( .A1(n450), .A2(n451), .Y(n730) );
  AO21X1_HVT U493 ( .A1(n118), .A2(n327), .A3(n484), .Y(n687) );
  NAND2X0_HVT U494 ( .A1(n463), .A2(n462), .Y(out[5]) );
  NAND2X0_HVT U495 ( .A1(n702), .A2(n385), .Y(n456) );
  NAND2X0_HVT U496 ( .A1(n712), .A2(in[6]), .Y(n457) );
  NAND2X0_HVT U497 ( .A1(n456), .A2(n457), .Y(out[1]) );
  NAND2X0_HVT U498 ( .A1(n671), .A2(n458), .Y(n459) );
  NAND2X0_HVT U499 ( .A1(n672), .A2(n311), .Y(n460) );
  NAND2X0_HVT U500 ( .A1(n459), .A2(n460), .Y(n670) );
  INVX1_HVT U501 ( .A(n770), .Y(n551) );
  NAND2X0_HVT U502 ( .A1(n629), .A2(in[6]), .Y(n462) );
  NAND2X0_HVT U503 ( .A1(n617), .A2(n385), .Y(n463) );
  NAND2X0_HVT U504 ( .A1(n481), .A2(n305), .Y(n479) );
  NAND2X0_HVT U505 ( .A1(n478), .A2(n479), .Y(n651) );
  NBUFFX2_HVT U506 ( .A(in[7]), .Y(n480) );
  INVX1_HVT U507 ( .A(n531), .Y(n530) );
  INVX1_HVT U508 ( .A(in[5]), .Y(n531) );
  AND2X1_HVT U509 ( .A1(n470), .A2(n734), .Y(n490) );
  MUX21X1_HVT U510 ( .A1(n365), .A2(n572), .S0(n507), .Y(n738) );
  NBUFFX2_HVT U511 ( .A(n782), .Y(n517) );
  NBUFFX2_HVT U512 ( .A(n782), .Y(n518) );
  AND2X1_HVT U513 ( .A1(n519), .A2(n717), .Y(n491) );
  MUX21X1_HVT U514 ( .A1(n471), .A2(n513), .S0(n218), .Y(n686) );
  NAND2X0_HVT U515 ( .A1(n316), .A2(n394), .Y(n782) );
  MUX21X1_HVT U516 ( .A1(n289), .A2(n467), .S0(n384), .Y(n580) );
  NBUFFX2_HVT U517 ( .A(n785), .Y(n519) );
  NBUFFX2_HVT U518 ( .A(n310), .Y(n520) );
  MUX21X1_HVT U519 ( .A1(n289), .A2(n282), .S0(n384), .Y(n603) );
  MUX21X1_HVT U520 ( .A1(n327), .A2(n365), .S0(n393), .Y(n770) );
  MUX21X1_HVT U521 ( .A1(n289), .A2(n512), .S0(n391), .Y(n600) );
  AND2X1_HVT U522 ( .A1(n391), .A2(n537), .Y(n493) );
  MUX21X1_HVT U523 ( .A1(n219), .A2(n364), .S0(n384), .Y(n577) );
  MUX21X1_HVT U524 ( .A1(n520), .A2(n513), .S0(n406), .Y(n584) );
  AND2X1_HVT U525 ( .A1(n282), .A2(n242), .Y(n494) );
  XNOR2X1_HVT U526 ( .A1(n313), .A2(n212), .Y(n495) );
  MUX21X1_HVT U527 ( .A1(n331), .A2(n521), .S0(n528), .Y(n665) );
  NBUFFX2_HVT U528 ( .A(n528), .Y(n504) );
  NBUFFX2_HVT U529 ( .A(n529), .Y(n505) );
  MUX21X1_HVT U530 ( .A1(n688), .A2(n535), .S0(n214), .Y(n685) );
  AND2X1_HVT U531 ( .A1(n471), .A2(n474), .Y(n496) );
  NAND2X0_HVT U532 ( .A1(n280), .A2(n316), .Y(n785) );
  XOR2X1_HVT U533 ( .A1(n393), .A2(n506), .Y(n747) );
  MUX21X1_HVT U534 ( .A1(n784), .A2(n525), .S0(n504), .Y(n664) );
  MUX21X1_HVT U535 ( .A1(n335), .A2(n327), .S0(n464), .Y(n581) );
  NBUFFX2_HVT U536 ( .A(n779), .Y(n516) );
  AND2X1_HVT U537 ( .A1(n515), .A2(n474), .Y(n498) );
  NBUFFX2_HVT U538 ( .A(n530), .Y(n529) );
  MUX21X1_HVT U539 ( .A1(n449), .A2(n467), .S0(n523), .Y(n583) );
  NAND2X0_HVT U540 ( .A1(n326), .A2(n230), .Y(n786) );
  NAND2X0_HVT U541 ( .A1(n326), .A2(n394), .Y(n779) );
  NBUFFX2_HVT U542 ( .A(in[0]), .Y(n511) );
endmodule

