
module sbox_16 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n7, n9, n19, n23, n33, n50, n121, n147, n210, n211, n212, n213, n216,
         n217, n218, n219, n226, n227, n229, n230, n231, n232, n235, n236,
         n238, n243, n252, n253, n254, n258, n259, n261, n264, n267, n271,
         n272, n273, n279, n280, n282, n283, n289, n293, n297, n298, n300,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779;

  NAND2X0_HVT U4 ( .A1(n230), .A2(n777), .Y(n776) );
  NAND2X0_HVT U5 ( .A1(n430), .A2(n502), .Y(n774) );
  NAND2X0_HVT U13 ( .A1(n768), .A2(n508), .Y(n769) );
  NAND2X0_HVT U15 ( .A1(n777), .A2(n33), .Y(n766) );
  NAND2X0_HVT U21 ( .A1(n230), .A2(n343), .Y(n761) );
  NAND2X0_HVT U24 ( .A1(n399), .A2(n343), .Y(n759) );
  NAND2X0_HVT U33 ( .A1(n426), .A2(n343), .Y(n751) );
  NAND2X0_HVT U42 ( .A1(n509), .A2(n499), .Y(n742) );
  NAND2X0_HVT U53 ( .A1(n731), .A2(n741), .Y(n732) );
  NAND2X0_HVT U56 ( .A1(n230), .A2(n727), .Y(n728) );
  NAND2X0_HVT U58 ( .A1(n508), .A2(n327), .Y(n725) );
  NAND2X0_HVT U62 ( .A1(n50), .A2(n506), .Y(n721) );
  AO21X1_HVT U66 ( .A1(n563), .A2(n516), .A3(n566), .Y(n717) );
  NAND2X0_HVT U73 ( .A1(n504), .A2(n370), .Y(n711) );
  MUX41X1_HVT U74 ( .A1(n712), .A3(n757), .A2(n711), .A4(n759), .S0(n489), 
        .S1(n457), .Y(n709) );
  MUX41X1_HVT U82 ( .A1(n739), .A3(n531), .A2(n569), .A4(n767), .S0(n490), 
        .S1(n411), .Y(n700) );
  AND2X1_HVT U83 ( .A1(n385), .A2(n402), .Y(n699) );
  MUX41X1_HVT U96 ( .A1(n569), .A3(n475), .A2(n561), .A4(n687), .S0(n489), 
        .S1(n365), .Y(n686) );
  NAND2X0_HVT U101 ( .A1(n680), .A2(n679), .Y(n681) );
  MUX41X1_HVT U103 ( .A1(n327), .A3(n328), .A2(n321), .A4(n749), .S0(n489), 
        .S1(n462), .Y(n677) );
  MUX41X1_HVT U105 ( .A1(n556), .A3(n736), .A2(n676), .A4(n550), .S0(n491), 
        .S1(n462), .Y(n675) );
  MUX41X1_HVT U106 ( .A1(n675), .A3(n678), .A2(n677), .A4(n682), .S0(n498), 
        .S1(n493), .Y(n674) );
  OA21X1_HVT U109 ( .A1(n543), .A2(n371), .A3(n407), .Y(n672) );
  NAND2X0_HVT U110 ( .A1(n507), .A2(n670), .Y(n671) );
  MUX41X1_HVT U114 ( .A1(n667), .A3(n673), .A2(n669), .A4(n672), .S0(n516), 
        .S1(n457), .Y(n666) );
  NAND2X0_HVT U123 ( .A1(n657), .A2(n656), .Y(n658) );
  MUX41X1_HVT U125 ( .A1(n761), .A3(n481), .A2(n535), .A4(n19), .S0(n490), 
        .S1(n495), .Y(n654) );
  MUX41X1_HVT U131 ( .A1(n649), .A3(n651), .A2(n650), .A4(n652), .S0(n516), 
        .S1(n521), .Y(n648) );
  MUX41X1_HVT U135 ( .A1(n9), .A3(n318), .A2(n774), .A4(n756), .S0(n491), .S1(
        n521), .Y(n645) );
  MUX41X1_HVT U147 ( .A1(n528), .A3(n370), .A2(n562), .A4(n738), .S0(n489), 
        .S1(n521), .Y(n635) );
  MUX41X1_HVT U148 ( .A1(n635), .A3(n639), .A2(n636), .A4(n640), .S0(n498), 
        .S1(n493), .Y(n634) );
  AND2X1_HVT U154 ( .A1(n496), .A2(n399), .Y(n628) );
  NAND2X0_HVT U158 ( .A1(n432), .A2(n419), .Y(n624) );
  MUX41X1_HVT U159 ( .A1(n389), .A3(n450), .A2(n624), .A4(n567), .S0(n484), 
        .S1(n411), .Y(n623) );
  AND2X1_HVT U162 ( .A1(n364), .A2(n370), .Y(n620) );
  MUX41X1_HVT U165 ( .A1(n761), .A3(n555), .A2(n738), .A4(n618), .S0(n521), 
        .S1(n484), .Y(n617) );
  NAND2X0_HVT U166 ( .A1(n508), .A2(n406), .Y(n616) );
  NAND2X0_HVT U174 ( .A1(n430), .A2(n448), .Y(n768) );
  MUX41X1_HVT U176 ( .A1(n283), .A3(n609), .A2(n538), .A4(n768), .S0(n521), 
        .S1(n483), .Y(n608) );
  NAND2X0_HVT U177 ( .A1(n510), .A2(n283), .Y(n607) );
  MUX41X1_HVT U178 ( .A1(n764), .A3(n607), .A2(n210), .A4(n746), .S0(n489), 
        .S1(n411), .Y(n606) );
  MUX41X1_HVT U182 ( .A1(n546), .A3(n428), .A2(n530), .A4(n552), .S0(n521), 
        .S1(n483), .Y(n602) );
  MUX41X1_HVT U189 ( .A1(n596), .A3(n768), .A2(n597), .A4(n550), .S0(n497), 
        .S1(n484), .Y(n595) );
  AO21X1_HVT U197 ( .A1(n478), .A2(n497), .A3(n558), .Y(n588) );
  NAND2X0_HVT U208 ( .A1(n417), .A2(n428), .Y(n670) );
  NAND2X0_HVT U212 ( .A1(n433), .A2(n333), .Y(n727) );
  NAND2X0_HVT U214 ( .A1(n448), .A2(n343), .Y(n578) );
  NAND2X0_HVT U215 ( .A1(n670), .A2(n504), .Y(n577) );
  NAND2X0_HVT U218 ( .A1(n318), .A2(n385), .Y(n631) );
  NAND2X0_HVT U220 ( .A1(n497), .A2(n578), .Y(n702) );
  INVX0_HVT U241 ( .A(n759), .Y(n569) );
  INVX0_HVT U245 ( .A(n774), .Y(n567) );
  INVX0_HVT U256 ( .A(n631), .Y(n558) );
  INVX0_HVT U259 ( .A(n753), .Y(n555) );
  INVX0_HVT U264 ( .A(n749), .Y(n553) );
  INVX0_HVT U265 ( .A(n757), .Y(n552) );
  INVX0_HVT U268 ( .A(n761), .Y(n551) );
  INVX0_HVT U270 ( .A(n577), .Y(n550) );
  INVX0_HVT U271 ( .A(n670), .Y(n549) );
  INVX0_HVT U278 ( .A(n751), .Y(n544) );
  INVX0_HVT U284 ( .A(n578), .Y(n541) );
  INVX0_HVT U289 ( .A(n679), .Y(n538) );
  INVX0_HVT U295 ( .A(n776), .Y(n534) );
  INVX0_HVT U296 ( .A(n766), .Y(n533) );
  INVX0_HVT U302 ( .A(n576), .Y(n529) );
  INVX0_HVT U310 ( .A(n571), .Y(n524) );
  NBUFFX2_HVT U1 ( .A(n324), .Y(n499) );
  INVX1_HVT U2 ( .A(n742), .Y(n568) );
  MUX21X1_HVT U3 ( .A1(n507), .A2(n692), .S0(n480), .Y(n691) );
  MUX21X1_HVT U6 ( .A1(n375), .A2(n424), .S0(n385), .Y(n687) );
  OA21X1_HVT U7 ( .A1(n293), .A2(n522), .A3(n752), .Y(n637) );
  NOR2X0_HVT U8 ( .A1(n382), .A2(n432), .Y(n293) );
  MUX21X1_HVT U9 ( .A1(n428), .A2(n446), .S0(n431), .Y(n747) );
  MUX21X1_HVT U10 ( .A1(n386), .A2(n764), .S0(n371), .Y(n649) );
  MUX21X1_HVT U11 ( .A1(n613), .A2(n612), .S0(n491), .Y(n611) );
  OA21X1_HVT U12 ( .A1(n522), .A2(n750), .A3(n537), .Y(n600) );
  INVX1_HVT U14 ( .A(n743), .Y(n530) );
  AND2X1_HVT U16 ( .A1(n375), .A2(n727), .Y(n7) );
  AND2X1_HVT U17 ( .A1(n322), .A2(n323), .Y(n9) );
  AND2X1_HVT U18 ( .A1(n356), .A2(n357), .Y(n19) );
  AND2X1_HVT U19 ( .A1(n313), .A2(n312), .Y(n23) );
  INVX0_HVT U20 ( .A(n775), .Y(n427) );
  INVX0_HVT U22 ( .A(n470), .Y(n640) );
  INVX1_HVT U23 ( .A(n547), .Y(n422) );
  NAND2X0_HVT U25 ( .A1(n387), .A2(n50), .Y(n121) );
  NAND2X0_HVT U26 ( .A1(n33), .A2(n509), .Y(n147) );
  NAND2X0_HVT U27 ( .A1(n121), .A2(n147), .Y(n738) );
  INVX0_HVT U28 ( .A(n387), .Y(n33) );
  INVX0_HVT U29 ( .A(n509), .Y(n50) );
  INVX1_HVT U30 ( .A(n23), .Y(n387) );
  MUX21X1_HVT U31 ( .A1(n654), .A2(n655), .S0(n516), .Y(n653) );
  MUX21X2_HVT U32 ( .A1(n754), .A2(n326), .S0(n497), .Y(n638) );
  MUX41X1_HVT U34 ( .A1(n693), .A3(n688), .A2(n686), .A4(n685), .S0(n437), 
        .S1(n261), .Y(n684) );
  NBUFFX2_HVT U35 ( .A(n325), .Y(n503) );
  INVX1_HVT U36 ( .A(n378), .Y(n510) );
  INVX1_HVT U37 ( .A(n421), .Y(n424) );
  INVX1_HVT U38 ( .A(n310), .Y(n226) );
  INVX2_HVT U39 ( .A(n512), .Y(n482) );
  INVX1_HVT U40 ( .A(n403), .Y(n404) );
  MUX21X2_HVT U41 ( .A1(n499), .A2(n469), .S0(n231), .Y(n668) );
  AND3X1_HVT U43 ( .A1(n506), .A2(n406), .A3(n702), .Y(n703) );
  INVX1_HVT U44 ( .A(n520), .Y(n410) );
  INVX1_HVT U45 ( .A(n410), .Y(n411) );
  INVX1_HVT U46 ( .A(n522), .Y(n457) );
  MUX21X1_HVT U47 ( .A1(n527), .A2(n499), .S0(n430), .Y(n763) );
  NBUFFX2_HVT U48 ( .A(n405), .Y(n496) );
  XOR2X1_HVT U49 ( .A1(n283), .A2(n433), .Y(n757) );
  INVX1_HVT U50 ( .A(n326), .Y(n327) );
  INVX1_HVT U51 ( .A(n755), .Y(n556) );
  MUX21X1_HVT U52 ( .A1(n544), .A2(n660), .S0(n231), .Y(n659) );
  INVX1_HVT U54 ( .A(n371), .Y(n231) );
  NBUFFX2_HVT U55 ( .A(n517), .Y(n516) );
  INVX1_HVT U57 ( .A(n491), .Y(n331) );
  INVX1_HVT U59 ( .A(n405), .Y(n451) );
  INVX1_HVT U60 ( .A(n289), .Y(n480) );
  OA21X1_HVT U61 ( .A1(n744), .A2(n522), .A3(n631), .Y(n632) );
  MUX21X1_HVT U63 ( .A1(n560), .A2(n527), .S0(n460), .Y(n618) );
  INVX1_HVT U64 ( .A(n293), .Y(n615) );
  INVX1_HVT U65 ( .A(n484), .Y(n309) );
  MUX21X1_HVT U67 ( .A1(n352), .A2(n507), .S0(n430), .Y(n597) );
  INVX1_HVT U68 ( .A(n482), .Y(n483) );
  MUX21X1_HVT U69 ( .A1(n343), .A2(n361), .S0(n518), .Y(n718) );
  MUX21X1_HVT U70 ( .A1(n703), .A2(n704), .S0(n331), .Y(n701) );
  AND3X1_HVT U71 ( .A1(n491), .A2(n343), .A3(n402), .Y(n651) );
  NAND2X0_HVT U72 ( .A1(n273), .A2(n279), .Y(n642) );
  NBUFFX2_HVT U75 ( .A(n520), .Y(n462) );
  INVX1_HVT U76 ( .A(n457), .Y(n393) );
  INVX1_HVT U77 ( .A(n523), .Y(n521) );
  INVX0_HVT U78 ( .A(n520), .Y(n522) );
  INVX1_HVT U79 ( .A(n522), .Y(n519) );
  INVX0_HVT U80 ( .A(n379), .Y(n335) );
  INVX0_HVT U81 ( .A(n496), .Y(n394) );
  INVX1_HVT U84 ( .A(n460), .Y(n343) );
  INVX1_HVT U85 ( .A(n494), .Y(n437) );
  INVX1_HVT U86 ( .A(n363), .Y(n340) );
  INVX1_HVT U87 ( .A(n380), .Y(n365) );
  INVX1_HVT U88 ( .A(in[0]), .Y(n261) );
  INVX0_HVT U89 ( .A(n491), .Y(n353) );
  INVX0_HVT U90 ( .A(n378), .Y(n432) );
  NBUFFX2_HVT U91 ( .A(n405), .Y(n497) );
  NBUFFX2_HVT U92 ( .A(in[0]), .Y(n498) );
  NBUFFX2_HVT U93 ( .A(n513), .Y(n492) );
  NBUFFX2_HVT U94 ( .A(n515), .Y(n493) );
  INVX0_HVT U95 ( .A(n504), .Y(n318) );
  INVX0_HVT U97 ( .A(n439), .Y(n433) );
  AND2X1_HVT U98 ( .A1(n359), .A2(n358), .Y(n210) );
  INVX0_HVT U99 ( .A(n744), .Y(n526) );
  MUX41X1_HVT U100 ( .A1(n717), .A3(n535), .A2(n718), .A4(n716), .S0(n309), 
        .S1(n457), .Y(n715) );
  INVX0_HVT U102 ( .A(n361), .Y(n770) );
  INVX0_HVT U104 ( .A(n554), .Y(n369) );
  INVX0_HVT U107 ( .A(n300), .Y(n420) );
  INVX1_HVT U108 ( .A(n523), .Y(n405) );
  MUX41X1_HVT U111 ( .A1(n625), .A3(n623), .A2(n630), .A4(n629), .S0(n418), 
        .S1(n498), .Y(n622) );
  INVX0_HVT U112 ( .A(n542), .Y(n389) );
  MUX21X1_HVT U113 ( .A1(n626), .A2(n627), .S0(n492), .Y(n625) );
  INVX0_HVT U115 ( .A(n324), .Y(n325) );
  INVX1_HVT U116 ( .A(n427), .Y(n428) );
  INVX0_HVT U117 ( .A(n547), .Y(n421) );
  AO21X1_HVT U118 ( .A1(n497), .A2(n689), .A3(n558), .Y(n690) );
  MUX21X2_HVT U119 ( .A1(n388), .A2(n777), .S0(n490), .Y(n673) );
  INVX1_HVT U120 ( .A(n429), .Y(n756) );
  INVX1_HVT U121 ( .A(n752), .Y(n465) );
  INVX1_HVT U122 ( .A(n333), .Y(n560) );
  INVX1_HVT U124 ( .A(n668), .Y(n486) );
  INVX0_HVT U126 ( .A(n574), .Y(n561) );
  NAND2X0_HVT U127 ( .A1(n328), .A2(n437), .Y(n211) );
  NAND2X0_HVT U128 ( .A1(n318), .A2(n516), .Y(n212) );
  NAND2X0_HVT U129 ( .A1(n211), .A2(n212), .Y(n716) );
  INVX0_HVT U130 ( .A(n445), .Y(n446) );
  MUX41X1_HVT U132 ( .A1(n349), .A3(n465), .A2(n402), .A4(n777), .S0(n231), 
        .S1(n410), .Y(n580) );
  INVX1_HVT U133 ( .A(n370), .Y(n566) );
  MUX21X1_HVT U134 ( .A1(n565), .A2(n450), .S0(n460), .Y(n621) );
  MUX41X1_HVT U136 ( .A1(n748), .A3(n751), .A2(n528), .A4(n474), .S0(n451), 
        .S1(n463), .Y(n644) );
  NAND2X0_HVT U137 ( .A1(n671), .A2(n492), .Y(n213) );
  NAND2X0_HVT U138 ( .A1(n752), .A2(n331), .Y(n216) );
  NAND2X0_HVT U139 ( .A1(n213), .A2(n216), .Y(n669) );
  NAND2X0_HVT U140 ( .A1(n404), .A2(n329), .Y(n217) );
  NAND2X0_HVT U141 ( .A1(n348), .A2(n460), .Y(n218) );
  NAND2X0_HVT U142 ( .A1(n217), .A2(n218), .Y(n752) );
  INVX1_HVT U143 ( .A(n378), .Y(n460) );
  INVX0_HVT U144 ( .A(n568), .Y(n219) );
  INVX1_HVT U145 ( .A(n769), .Y(n542) );
  INVX1_HVT U146 ( .A(n280), .Y(n282) );
  NAND2X0_HVT U149 ( .A1(n753), .A2(n231), .Y(n227) );
  NAND2X0_HVT U150 ( .A1(n556), .A2(n463), .Y(n229) );
  NAND2X0_HVT U151 ( .A1(n227), .A2(n229), .Y(n652) );
  MUX41X1_HVT U152 ( .A1(n619), .A3(n614), .A2(n617), .A4(n611), .S0(n261), 
        .S1(n418), .Y(n610) );
  INVX0_HVT U153 ( .A(n427), .Y(n230) );
  INVX0_HVT U155 ( .A(n767), .Y(n532) );
  MUX21X1_HVT U156 ( .A1(n382), .A2(n348), .S0(n432), .Y(n767) );
  MUX21X2_HVT U157 ( .A1(n381), .A2(n23), .S0(n431), .Y(n743) );
  NAND2X0_HVT U160 ( .A1(n312), .A2(n313), .Y(n232) );
  INVX0_HVT U161 ( .A(n779), .Y(n565) );
  INVX0_HVT U163 ( .A(n762), .Y(n531) );
  INVX1_HVT U164 ( .A(n449), .Y(n375) );
  INVX0_HVT U167 ( .A(n378), .Y(n235) );
  NAND2X0_HVT U168 ( .A1(n502), .A2(n340), .Y(n236) );
  NAND2X0_HVT U169 ( .A1(n469), .A2(n461), .Y(n238) );
  NAND2X0_HVT U170 ( .A1(n236), .A2(n238), .Y(n753) );
  INVX0_HVT U171 ( .A(n368), .Y(n469) );
  INVX0_HVT U172 ( .A(n378), .Y(n461) );
  MUX41X1_HVT U173 ( .A1(n715), .A3(n723), .A2(n719), .A4(n729), .S0(in[6]), 
        .S1(n498), .Y(out[0]) );
  NAND2X0_HVT U175 ( .A1(n714), .A2(n490), .Y(n243) );
  NAND2X0_HVT U179 ( .A1(n740), .A2(n353), .Y(n252) );
  NAND2X0_HVT U180 ( .A1(n243), .A2(n252), .Y(n713) );
  XOR2X1_HVT U181 ( .A1(n429), .A2(n519), .Y(n740) );
  INVX0_HVT U183 ( .A(n396), .Y(n527) );
  INVX1_HVT U184 ( .A(n379), .Y(n431) );
  INVX1_HVT U185 ( .A(n330), .Y(n379) );
  INVX0_HVT U186 ( .A(n772), .Y(n253) );
  INVX0_HVT U187 ( .A(n253), .Y(n254) );
  NAND2X0_HVT U188 ( .A1(n568), .A2(n394), .Y(n258) );
  NAND2X0_HVT U190 ( .A1(n210), .A2(n521), .Y(n259) );
  NAND2X0_HVT U191 ( .A1(n258), .A2(n259), .Y(n589) );
  MUX41X1_HVT U192 ( .A1(n653), .A3(n666), .A2(n648), .A4(n661), .S0(n332), 
        .S1(n261), .Y(out[3]) );
  INVX0_HVT U193 ( .A(n763), .Y(n525) );
  MUX41X1_HVT U194 ( .A1(n646), .A3(n645), .A2(n644), .A4(n642), .S0(n418), 
        .S1(n261), .Y(n641) );
  INVX0_HVT U195 ( .A(n388), .Y(n748) );
  INVX1_HVT U196 ( .A(n570), .Y(n528) );
  NAND2X0_HVT U198 ( .A1(n662), .A2(n418), .Y(n264) );
  NAND2X0_HVT U199 ( .A1(n665), .A2(n493), .Y(n267) );
  NAND2X0_HVT U200 ( .A1(n264), .A2(n267), .Y(n661) );
  INVX1_HVT U201 ( .A(n330), .Y(n438) );
  INVX0_HVT U202 ( .A(n438), .Y(n430) );
  INVX0_HVT U203 ( .A(n317), .Y(n613) );
  NBUFFX2_HVT U204 ( .A(n405), .Y(n495) );
  INVX1_HVT U205 ( .A(n750), .Y(n564) );
  MUX21X1_HVT U206 ( .A1(n600), .A2(n601), .S0(n490), .Y(n599) );
  NAND2X0_HVT U207 ( .A1(n760), .A2(n394), .Y(n271) );
  NAND2X0_HVT U209 ( .A1(n546), .A2(n495), .Y(n272) );
  NAND2X0_HVT U210 ( .A1(n271), .A2(n272), .Y(n643) );
  NAND2X0_HVT U211 ( .A1(n776), .A2(n490), .Y(n273) );
  NAND2X0_HVT U213 ( .A1(n643), .A2(n463), .Y(n279) );
  INVX0_HVT U216 ( .A(n503), .Y(n362) );
  MUX21X1_HVT U217 ( .A1(n553), .A2(n564), .S0(n492), .Y(n664) );
  INVX0_HVT U219 ( .A(n396), .Y(n280) );
  INVX0_HVT U221 ( .A(n440), .Y(n283) );
  INVX0_HVT U222 ( .A(n368), .Y(n440) );
  XOR2X2_HVT U223 ( .A1(n282), .A2(n461), .Y(n735) );
  XNOR2X2_HVT U224 ( .A1(n230), .A2(n510), .Y(n477) );
  XNOR2X1_HVT U225 ( .A1(n520), .A2(n511), .Y(n289) );
  INVX1_HVT U226 ( .A(n330), .Y(n439) );
  INVX0_HVT U227 ( .A(n507), .Y(n487) );
  INVX1_HVT U228 ( .A(n758), .Y(n471) );
  INVX1_HVT U229 ( .A(n439), .Y(n417) );
  INVX1_HVT U230 ( .A(n386), .Y(n472) );
  NAND2X0_HVT U231 ( .A1(n690), .A2(n353), .Y(n297) );
  NAND2X0_HVT U232 ( .A1(n691), .A2(n492), .Y(n298) );
  NAND2X0_HVT U233 ( .A1(n297), .A2(n298), .Y(n688) );
  INVX1_HVT U234 ( .A(n438), .Y(n509) );
  INVX0_HVT U235 ( .A(in[3]), .Y(n300) );
  NAND2X0_HVT U236 ( .A1(n633), .A2(n489), .Y(n303) );
  NAND2X0_HVT U237 ( .A1(n632), .A2(n353), .Y(n304) );
  NAND2X0_HVT U238 ( .A1(n303), .A2(n304), .Y(n630) );
  MUX21X1_HVT U239 ( .A1(n424), .A2(n527), .S0(n385), .Y(n609) );
  NAND2X0_HVT U240 ( .A1(n548), .A2(n519), .Y(n376) );
  INVX1_HVT U242 ( .A(n689), .Y(n548) );
  INVX1_HVT U243 ( .A(n464), .Y(n665) );
  NAND2X0_HVT U244 ( .A1(n374), .A2(n497), .Y(n305) );
  AND2X1_HVT U246 ( .A1(n305), .A2(n752), .Y(n612) );
  INVX1_HVT U247 ( .A(n514), .Y(n513) );
  INVX1_HVT U248 ( .A(in[2]), .Y(n514) );
  MUX21X1_HVT U249 ( .A1(n352), .A2(n469), .S0(n363), .Y(n755) );
  INVX1_HVT U250 ( .A(in[5]), .Y(n518) );
  NAND2X0_HVT U251 ( .A1(n345), .A2(n344), .Y(n306) );
  INVX1_HVT U252 ( .A(in[4]), .Y(n368) );
  NAND2X0_HVT U253 ( .A1(n634), .A2(n434), .Y(n467) );
  MUX21X2_HVT U254 ( .A1(n637), .A2(n638), .S0(n331), .Y(n636) );
  MUX21X2_HVT U255 ( .A1(n316), .A2(n395), .S0(n439), .Y(n349) );
  NAND2X0_HVT U257 ( .A1(n565), .A2(n340), .Y(n307) );
  NAND2X0_HVT U258 ( .A1(n424), .A2(n510), .Y(n308) );
  NAND2X0_HVT U260 ( .A1(n307), .A2(n308), .Y(n746) );
  INVX0_HVT U261 ( .A(n746), .Y(n545) );
  MUX41X1_HVT U262 ( .A1(n254), .A3(n540), .A2(n616), .A4(n615), .S0(n309), 
        .S1(n519), .Y(n614) );
  MUX21X1_HVT U263 ( .A1(n503), .A2(n527), .S0(n432), .Y(n744) );
  NAND2X0_HVT U266 ( .A1(n554), .A2(n334), .Y(n312) );
  NAND2X0_HVT U267 ( .A1(n310), .A2(n311), .Y(n313) );
  INVX0_HVT U269 ( .A(n300), .Y(n310) );
  INVX0_HVT U272 ( .A(n554), .Y(n311) );
  INVX0_HVT U273 ( .A(in[4]), .Y(n554) );
  INVX0_HVT U274 ( .A(n232), .Y(n445) );
  NAND2X0_HVT U275 ( .A1(n659), .A2(n393), .Y(n314) );
  NAND2X0_HVT U276 ( .A1(n658), .A2(n365), .Y(n315) );
  NAND2X0_HVT U277 ( .A1(n314), .A2(n315), .Y(n655) );
  INVX0_HVT U279 ( .A(n360), .Y(n316) );
  INVX0_HVT U280 ( .A(in[1]), .Y(n378) );
  MUX41X1_HVT U281 ( .A1(n608), .A3(n606), .A2(n605), .A4(n604), .S0(n418), 
        .S1(n261), .Y(n603) );
  INVX1_HVT U282 ( .A(n482), .Y(n484) );
  INVX0_HVT U283 ( .A(n321), .Y(n754) );
  INVX0_HVT U285 ( .A(n523), .Y(n520) );
  MUX21X1_HVT U286 ( .A1(n697), .A2(n399), .S0(n496), .Y(n601) );
  MUX21X1_HVT U287 ( .A1(n419), .A2(n561), .S0(n496), .Y(n714) );
  MUX21X1_HVT U288 ( .A1(n318), .A2(n574), .S0(n496), .Y(n317) );
  INVX1_HVT U290 ( .A(in[7]), .Y(n523) );
  NAND2X0_HVT U291 ( .A1(n539), .A2(n394), .Y(n319) );
  NAND2X0_HVT U292 ( .A1(n318), .A2(n495), .Y(n320) );
  NAND2X0_HVT U293 ( .A1(n319), .A2(n320), .Y(n633) );
  MUX21X1_HVT U294 ( .A1(n440), .A2(n422), .S0(n433), .Y(n321) );
  INVX0_HVT U297 ( .A(n422), .Y(n425) );
  NAND2X0_HVT U298 ( .A1(n446), .A2(n340), .Y(n322) );
  NAND2X0_HVT U299 ( .A1(n560), .A2(n363), .Y(n323) );
  INVX0_HVT U300 ( .A(n379), .Y(n363) );
  MUX41X1_HVT U301 ( .A1(n738), .A3(n745), .A2(n710), .A4(n475), .S0(n393), 
        .S1(n514), .Y(n598) );
  INVX1_HVT U303 ( .A(n514), .Y(n512) );
  OA21X1_HVT U304 ( .A1(n522), .A2(n773), .A3(n545), .Y(n584) );
  INVX0_HVT U305 ( .A(n773), .Y(n535) );
  INVX1_HVT U306 ( .A(n334), .Y(n324) );
  INVX0_HVT U307 ( .A(n508), .Y(n419) );
  INVX1_HVT U308 ( .A(n777), .Y(n326) );
  INVX0_HVT U309 ( .A(in[3]), .Y(n334) );
  INVX1_HVT U311 ( .A(n575), .Y(n540) );
  MUX21X1_HVT U312 ( .A1(n382), .A2(n404), .S0(n510), .Y(n429) );
  AND2X1_HVT U313 ( .A1(n345), .A2(n344), .Y(n328) );
  INVX0_HVT U314 ( .A(in[1]), .Y(n329) );
  INVX1_HVT U315 ( .A(n329), .Y(n330) );
  INVX1_HVT U316 ( .A(n434), .Y(n332) );
  INVX1_HVT U317 ( .A(in[6]), .Y(n434) );
  MUX41X1_HVT U318 ( .A1(n529), .A3(n551), .A2(n525), .A4(n531), .S0(n365), 
        .S1(n516), .Y(n734) );
  NAND2X0_HVT U319 ( .A1(n325), .A2(n369), .Y(n333) );
  MUX21X1_HVT U320 ( .A1(n565), .A2(n447), .S0(n456), .Y(n773) );
  INVX1_HVT U321 ( .A(n23), .Y(n448) );
  MUX41X1_HVT U322 ( .A1(n581), .A3(n583), .A2(n580), .A4(n582), .S0(n498), 
        .S1(n418), .Y(n579) );
  INVX0_HVT U323 ( .A(n565), .Y(n352) );
  MUX21X1_HVT U324 ( .A1(n421), .A2(n387), .S0(n335), .Y(n336) );
  INVX0_HVT U325 ( .A(n536), .Y(n337) );
  NAND2X0_HVT U326 ( .A1(n765), .A2(n394), .Y(n338) );
  NAND2X0_HVT U327 ( .A1(n7), .A2(n495), .Y(n339) );
  NAND2X0_HVT U328 ( .A1(n338), .A2(n339), .Y(n585) );
  INVX0_HVT U329 ( .A(n765), .Y(n536) );
  OR2X1_HVT U330 ( .A1(n440), .A2(n511), .Y(n749) );
  NAND2X0_HVT U331 ( .A1(n509), .A2(n282), .Y(n777) );
  INVX0_HVT U332 ( .A(n336), .Y(n543) );
  NAND2X0_HVT U333 ( .A1(n499), .A2(n340), .Y(n341) );
  NAND2X0_HVT U334 ( .A1(n425), .A2(n385), .Y(n342) );
  NAND2X0_HVT U335 ( .A1(n341), .A2(n342), .Y(n745) );
  INVX1_HVT U336 ( .A(n379), .Y(n385) );
  NAND2X0_HVT U337 ( .A1(n421), .A2(n343), .Y(n344) );
  NAND2X0_HVT U338 ( .A1(n499), .A2(n432), .Y(n345) );
  NAND2X0_HVT U339 ( .A1(n387), .A2(n50), .Y(n346) );
  NAND2X0_HVT U340 ( .A1(n395), .A2(n385), .Y(n347) );
  NAND2X0_HVT U341 ( .A1(n346), .A2(n347), .Y(n707) );
  INVX1_HVT U342 ( .A(n253), .Y(n348) );
  MUX21X1_HVT U343 ( .A1(n254), .A2(n762), .S0(n380), .Y(n704) );
  AO21X1_HVT U344 ( .A1(n492), .A2(n254), .A3(n364), .Y(n663) );
  MUX21X1_HVT U345 ( .A1(n767), .A2(n465), .S0(n463), .Y(n683) );
  AO21X1_HVT U346 ( .A1(n439), .A2(n560), .A3(n522), .Y(n680) );
  NAND2X0_HVT U347 ( .A1(n628), .A2(n289), .Y(n350) );
  NAND2X0_HVT U348 ( .A1(n507), .A2(n480), .Y(n351) );
  NAND2X0_HVT U349 ( .A1(n350), .A2(n351), .Y(n627) );
  MUX21X1_HVT U350 ( .A1(n469), .A2(n282), .S0(n235), .Y(n762) );
  MUX41X1_HVT U351 ( .A1(n671), .A3(n476), .A2(n506), .A4(n553), .S0(n489), 
        .S1(n462), .Y(n629) );
  INVX1_HVT U352 ( .A(n493), .Y(n418) );
  MUX21X1_HVT U353 ( .A1(n477), .A2(n536), .S0(n231), .Y(n650) );
  MUX21X1_HVT U354 ( .A1(n427), .A2(n362), .S0(n511), .Y(n361) );
  MUX41X1_HVT U355 ( .A1(n701), .A3(n698), .A2(n700), .A4(n696), .S0(n261), 
        .S1(n418), .Y(n695) );
  OR2X1_HVT U356 ( .A1(n335), .A2(n352), .Y(n697) );
  NAND2X0_HVT U357 ( .A1(n524), .A2(n353), .Y(n354) );
  NAND2X0_HVT U358 ( .A1(n647), .A2(n491), .Y(n355) );
  NAND2X0_HVT U359 ( .A1(n354), .A2(n355), .Y(n646) );
  NAND2X0_HVT U360 ( .A1(n425), .A2(n340), .Y(n356) );
  NAND2X0_HVT U361 ( .A1(n500), .A2(n430), .Y(n357) );
  MUX21X1_HVT U362 ( .A1(n19), .A2(n348), .S0(n495), .Y(n647) );
  NAND2X0_HVT U363 ( .A1(n469), .A2(n340), .Y(n358) );
  NAND2X0_HVT U364 ( .A1(n504), .A2(n433), .Y(n359) );
  INVX1_HVT U365 ( .A(n403), .Y(n360) );
  MUX41X1_HVT U366 ( .A1(n620), .A3(n557), .A2(n621), .A4(n477), .S0(n309), 
        .S1(n365), .Y(n619) );
  INVX1_HVT U367 ( .A(n511), .Y(n456) );
  INVX1_HVT U368 ( .A(n438), .Y(n511) );
  INVX1_HVT U369 ( .A(n449), .Y(n447) );
  INVX0_HVT U370 ( .A(n450), .Y(n364) );
  INVX0_HVT U371 ( .A(n496), .Y(n380) );
  INVX0_HVT U372 ( .A(n764), .Y(n557) );
  INVX1_HVT U373 ( .A(n448), .Y(n450) );
  XOR2X1_HVT U374 ( .A1(n417), .A2(n482), .Y(n488) );
  MUX41X1_HVT U375 ( .A1(n763), .A3(n540), .A2(n771), .A4(n728), .S0(n393), 
        .S1(n494), .Y(n726) );
  MUX41X1_HVT U376 ( .A1(n595), .A3(n598), .A2(n599), .A4(n602), .S0(n515), 
        .S1(n498), .Y(n594) );
  NBUFFX2_HVT U377 ( .A(n368), .Y(n500) );
  MUX21X1_HVT U378 ( .A1(n469), .A2(n560), .S0(n363), .Y(n764) );
  NAND2X0_HVT U379 ( .A1(n674), .A2(n434), .Y(n366) );
  NAND2X0_HVT U380 ( .A1(n684), .A2(n332), .Y(n367) );
  NAND2X0_HVT U381 ( .A1(n366), .A2(n367), .Y(out[2]) );
  MUX21X1_HVT U382 ( .A1(n503), .A2(n565), .S0(n417), .Y(n771) );
  INVX0_HVT U383 ( .A(n745), .Y(n546) );
  MUX41X1_HVT U384 ( .A1(n743), .A3(n756), .A2(n9), .A4(n254), .S0(n495), .S1(
        n483), .Y(n591) );
  MUX21X1_HVT U385 ( .A1(n663), .A2(n664), .S0(n495), .Y(n662) );
  MUX41X1_HVT U386 ( .A1(n534), .A3(n306), .A2(n389), .A4(n7), .S0(n519), .S1(
        n512), .Y(n604) );
  NBUFFX2_HVT U387 ( .A(n710), .Y(n370) );
  NAND2X0_HVT U388 ( .A1(n335), .A2(n360), .Y(n710) );
  INVX1_HVT U389 ( .A(n573), .Y(n559) );
  INVX1_HVT U390 ( .A(n513), .Y(n371) );
  INVX0_HVT U391 ( .A(n771), .Y(n563) );
  INVX0_HVT U392 ( .A(n390), .Y(n372) );
  NAND2X0_HVT U393 ( .A1(n499), .A2(n430), .Y(n373) );
  NAND2X0_HVT U394 ( .A1(n447), .A2(n456), .Y(n374) );
  NAND2X0_HVT U395 ( .A1(n373), .A2(n455), .Y(n760) );
  MUX21X1_HVT U396 ( .A1(n502), .A2(n348), .S0(n439), .Y(n574) );
  MUX41X1_HVT U397 ( .A1(n561), .A3(n364), .A2(n747), .A4(n352), .S0(n482), 
        .S1(n462), .Y(n590) );
  NAND2X0_HVT U398 ( .A1(n746), .A2(n394), .Y(n377) );
  NAND2X0_HVT U399 ( .A1(n376), .A2(n377), .Y(n626) );
  INVX1_HVT U400 ( .A(n445), .Y(n449) );
  INVX1_HVT U401 ( .A(n492), .Y(n463) );
  NAND2X0_HVT U402 ( .A1(n420), .A2(n501), .Y(n381) );
  NAND2X0_HVT U403 ( .A1(n420), .A2(n501), .Y(n382) );
  INVX0_HVT U404 ( .A(n760), .Y(n537) );
  NAND2X0_HVT U405 ( .A1(n730), .A2(n353), .Y(n383) );
  NAND2X0_HVT U406 ( .A1(n734), .A2(n491), .Y(n384) );
  NAND2X0_HVT U407 ( .A1(n383), .A2(n384), .Y(n729) );
  MUX21X1_HVT U408 ( .A1(n733), .A2(n732), .S0(n394), .Y(n730) );
  MUX21X1_HVT U409 ( .A1(n500), .A2(n360), .S0(n431), .Y(n388) );
  MUX21X1_HVT U410 ( .A1(n505), .A2(n395), .S0(n235), .Y(n386) );
  MUX41X1_HVT U411 ( .A1(n735), .A3(n742), .A2(n593), .A4(n749), .S0(n394), 
        .S1(n483), .Y(n592) );
  MUX41X1_HVT U412 ( .A1(n306), .A3(n707), .A2(n548), .A4(n539), .S0(n484), 
        .S1(n497), .Y(n706) );
  INVX1_HVT U413 ( .A(n572), .Y(n539) );
  MUX41X1_HVT U414 ( .A1(n475), .A3(n562), .A2(n766), .A4(n432), .S0(n353), 
        .S1(n462), .Y(n685) );
  NAND2X0_HVT U415 ( .A1(n487), .A2(n390), .Y(n391) );
  NAND2X0_HVT U416 ( .A1(n486), .A2(n372), .Y(n392) );
  NAND2X0_HVT U417 ( .A1(n392), .A2(n391), .Y(n485) );
  INVX1_HVT U418 ( .A(n488), .Y(n390) );
  INVX1_HVT U419 ( .A(n440), .Y(n395) );
  NAND2X0_HVT U420 ( .A1(n420), .A2(n368), .Y(n396) );
  NAND2X0_HVT U421 ( .A1(n594), .A2(n434), .Y(n397) );
  NAND2X0_HVT U422 ( .A1(n603), .A2(n332), .Y(n398) );
  NAND2X0_HVT U423 ( .A1(n397), .A2(n398), .Y(out[6]) );
  NBUFFX2_HVT U424 ( .A(n499), .Y(n399) );
  NAND2X0_HVT U425 ( .A1(n724), .A2(n353), .Y(n400) );
  NAND2X0_HVT U426 ( .A1(n726), .A2(n490), .Y(n401) );
  NAND2X0_HVT U427 ( .A1(n401), .A2(n400), .Y(n723) );
  INVX1_HVT U428 ( .A(n500), .Y(n402) );
  MUX21X1_HVT U429 ( .A1(n499), .A2(n283), .S0(n496), .Y(n692) );
  NBUFFX2_HVT U430 ( .A(n368), .Y(n501) );
  INVX0_HVT U431 ( .A(n779), .Y(n403) );
  INVX0_HVT U432 ( .A(n562), .Y(n406) );
  INVX0_HVT U433 ( .A(n727), .Y(n562) );
  MUX21X1_HVT U434 ( .A1(n565), .A2(n502), .S0(n431), .Y(n750) );
  NBUFFX2_HVT U435 ( .A(n300), .Y(n502) );
  MUX41X1_HVT U436 ( .A1(n760), .A3(n564), .A2(n769), .A4(n728), .S0(n331), 
        .S1(n410), .Y(n581) );
  MUX21X1_HVT U437 ( .A1(n504), .A2(n423), .S0(n417), .Y(n407) );
  INVX0_HVT U438 ( .A(n423), .Y(n426) );
  MUX41X1_HVT U439 ( .A1(n587), .A3(n591), .A2(n590), .A4(n592), .S0(n498), 
        .S1(n493), .Y(n586) );
  NAND2X0_HVT U440 ( .A1(n588), .A2(n492), .Y(n408) );
  NAND2X0_HVT U441 ( .A1(n589), .A2(n463), .Y(n409) );
  NAND2X0_HVT U442 ( .A1(n409), .A2(n408), .Y(n587) );
  NAND2X0_HVT U443 ( .A1(n720), .A2(n353), .Y(n412) );
  NAND2X0_HVT U444 ( .A1(n722), .A2(n231), .Y(n413) );
  NAND2X0_HVT U445 ( .A1(n412), .A2(n413), .Y(n719) );
  NAND2X0_HVT U446 ( .A1(n476), .A2(n414), .Y(n415) );
  NAND2X0_HVT U447 ( .A1(n683), .A2(n737), .Y(n416) );
  NAND2X0_HVT U448 ( .A1(n415), .A2(n416), .Y(n682) );
  INVX0_HVT U449 ( .A(n737), .Y(n414) );
  XOR2X1_HVT U450 ( .A1(n371), .A2(n451), .Y(n737) );
  NBUFFX2_HVT U451 ( .A(n404), .Y(n508) );
  MUX41X1_HVT U452 ( .A1(n709), .A3(n706), .A2(n713), .A4(n708), .S0(n261), 
        .S1(n494), .Y(n705) );
  MUX41X1_HVT U453 ( .A1(n526), .A3(n472), .A2(n748), .A4(n770), .S0(n411), 
        .S1(n482), .Y(n582) );
  NBUFFX2_HVT U454 ( .A(n772), .Y(n504) );
  INVX0_HVT U455 ( .A(n547), .Y(n423) );
  INVX1_HVT U456 ( .A(n505), .Y(n547) );
  MUX41X1_HVT U457 ( .A1(n694), .A3(n529), .A2(n219), .A4(n738), .S0(n309), 
        .S1(n451), .Y(n693) );
  MUX41X1_HVT U458 ( .A1(n557), .A3(n476), .A2(n33), .A4(n536), .S0(n393), 
        .S1(n494), .Y(n722) );
  NAND2X0_HVT U459 ( .A1(n695), .A2(n434), .Y(n435) );
  NAND2X0_HVT U460 ( .A1(n705), .A2(n332), .Y(n436) );
  NAND2X0_HVT U461 ( .A1(n435), .A2(n436), .Y(out[1]) );
  MUX41X1_HVT U462 ( .A1(n532), .A3(n542), .A2(n533), .A4(n721), .S0(n410), 
        .S1(n437), .Y(n720) );
  NAND2X0_HVT U463 ( .A1(n441), .A2(n442), .Y(out[5]) );
  MUX21X1_HVT U464 ( .A1(n753), .A2(n577), .S0(n495), .Y(n571) );
  MUX41X1_HVT U465 ( .A1(n407), .A3(n479), .A2(n725), .A4(n481), .S0(n393), 
        .S1(n437), .Y(n724) );
  NAND2X0_HVT U466 ( .A1(n467), .A2(n468), .Y(out[4]) );
  NAND2X0_HVT U467 ( .A1(n586), .A2(n332), .Y(n458) );
  NAND2X0_HVT U468 ( .A1(n610), .A2(n434), .Y(n441) );
  NAND2X0_HVT U469 ( .A1(n622), .A2(n332), .Y(n442) );
  NAND2X0_HVT U470 ( .A1(n399), .A2(n437), .Y(n443) );
  NAND2X0_HVT U471 ( .A1(n749), .A2(n516), .Y(n444) );
  NAND2X0_HVT U472 ( .A1(n443), .A2(n444), .Y(n733) );
  NAND2X0_HVT U473 ( .A1(n584), .A2(n463), .Y(n452) );
  NAND2X0_HVT U474 ( .A1(n585), .A2(n490), .Y(n453) );
  NAND2X0_HVT U475 ( .A1(n452), .A2(n453), .Y(n583) );
  NAND2X0_HVT U476 ( .A1(n502), .A2(n511), .Y(n454) );
  NAND2X0_HVT U477 ( .A1(n375), .A2(n456), .Y(n455) );
  NAND2X0_HVT U478 ( .A1(n374), .A2(n454), .Y(n765) );
  NAND2X0_HVT U479 ( .A1(n579), .A2(n434), .Y(n459) );
  NAND2X0_HVT U480 ( .A1(n459), .A2(n458), .Y(out[7]) );
  MUX41X1_HVT U481 ( .A1(n537), .A3(n364), .A2(n337), .A4(n699), .S0(n489), 
        .S1(n519), .Y(n698) );
  MUX41X1_HVT U482 ( .A1(n559), .A3(n697), .A2(n478), .A4(n474), .S0(n489), 
        .S1(n457), .Y(n696) );
  MUX41X1_HVT U483 ( .A1(n562), .A3(n559), .A2(n487), .A4(n471), .S0(n492), 
        .S1(n411), .Y(n708) );
  MUX41X1_HVT U484 ( .A1(n755), .A3(n349), .A2(n541), .A4(n210), .S0(n484), 
        .S1(n365), .Y(n605) );
  MUX41X1_HVT U485 ( .A1(n465), .A3(n758), .A2(n466), .A4(n542), .S0(n309), 
        .S1(n451), .Y(n464) );
  NAND2X0_HVT U486 ( .A1(n363), .A2(n450), .Y(n466) );
  NAND2X0_HVT U487 ( .A1(n641), .A2(n332), .Y(n468) );
  MUX41X1_HVT U488 ( .A1(n772), .A3(n549), .A2(n33), .A4(n537), .S0(n309), 
        .S1(n451), .Y(n639) );
  MUX41X1_HVT U489 ( .A1(n473), .A3(n472), .A2(n471), .A4(n746), .S0(n489), 
        .S1(n451), .Y(n470) );
  NAND2X0_HVT U490 ( .A1(n254), .A2(n438), .Y(n473) );
  INVX1_HVT U491 ( .A(n518), .Y(n517) );
  NBUFFX2_HVT U492 ( .A(n775), .Y(n505) );
  MUX21X1_HVT U493 ( .A1(n426), .A2(n419), .S0(n516), .Y(n731) );
  AND2X1_HVT U494 ( .A1(n507), .A2(n710), .Y(n474) );
  MUX21X1_HVT U495 ( .A1(n448), .A2(n527), .S0(n510), .Y(n758) );
  MUX21X1_HVT U496 ( .A1(n375), .A2(n395), .S0(n460), .Y(n679) );
  NAND2X0_HVT U497 ( .A1(n368), .A2(n226), .Y(n775) );
  MUX21X1_HVT U498 ( .A1(n230), .A2(n254), .S0(n385), .Y(n694) );
  NBUFFX2_HVT U499 ( .A(n778), .Y(n506) );
  MUX21X1_HVT U500 ( .A1(n502), .A2(n446), .S0(n235), .Y(n572) );
  MUX21X1_HVT U501 ( .A1(n500), .A2(n503), .S0(n509), .Y(n660) );
  MUX21X1_HVT U502 ( .A1(n502), .A2(n500), .S0(n461), .Y(n593) );
  NBUFFX2_HVT U503 ( .A(n778), .Y(n507) );
  MUX21X1_HVT U504 ( .A1(n502), .A2(n360), .S0(n385), .Y(n596) );
  MUX21X1_HVT U505 ( .A1(n507), .A2(n423), .S0(n335), .Y(n570) );
  MUX21X1_HVT U506 ( .A1(n230), .A2(n352), .S0(n430), .Y(n689) );
  XOR2X1_HVT U507 ( .A1(n510), .A2(n560), .Y(n739) );
  MUX21X1_HVT U508 ( .A1(n506), .A2(n283), .S0(n335), .Y(n576) );
  AND2X1_HVT U509 ( .A1(n509), .A2(n487), .Y(n475) );
  AND2X1_HVT U510 ( .A1(n508), .A2(n670), .Y(n476) );
  XNOR2X1_HVT U511 ( .A1(n404), .A2(n432), .Y(n478) );
  MUX21X1_HVT U512 ( .A1(n504), .A2(n283), .S0(n461), .Y(n712) );
  MUX21X1_HVT U513 ( .A1(n254), .A2(n508), .S0(n491), .Y(n657) );
  NBUFFX2_HVT U514 ( .A(n513), .Y(n491) );
  NBUFFX2_HVT U515 ( .A(n513), .Y(n490) );
  NBUFFX2_HVT U516 ( .A(n515), .Y(n494) );
  NBUFFX2_HVT U517 ( .A(n513), .Y(n489) );
  MUX21X1_HVT U518 ( .A1(n681), .A2(n524), .S0(n491), .Y(n678) );
  XOR2X1_HVT U519 ( .A1(n235), .A2(n499), .Y(n736) );
  MUX21X1_HVT U520 ( .A1(n254), .A2(n450), .S0(n335), .Y(n676) );
  NAND2X0_HVT U521 ( .A1(n420), .A2(n501), .Y(n778) );
  AND2X1_HVT U522 ( .A1(n375), .A2(n343), .Y(n479) );
  MUX21X1_HVT U523 ( .A1(n499), .A2(n560), .S0(n509), .Y(n573) );
  XOR2X1_HVT U524 ( .A1(n235), .A2(n515), .Y(n741) );
  MUX21X1_HVT U525 ( .A1(n327), .A2(n439), .S0(n490), .Y(n656) );
  AND2X1_HVT U526 ( .A1(n503), .A2(n50), .Y(n481) );
  NBUFFX2_HVT U527 ( .A(n517), .Y(n515) );
  NAND2X0_HVT U528 ( .A1(n369), .A2(n324), .Y(n779) );
  NAND2X0_HVT U529 ( .A1(n226), .A2(n369), .Y(n772) );
  MUX21X1_HVT U530 ( .A1(n402), .A2(n387), .S0(n460), .Y(n575) );
  INVX0_HVT U531 ( .A(n485), .Y(n667) );
endmodule

