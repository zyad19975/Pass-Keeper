
module inv_sbox_1 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n196, n197, n198, n199, n200, n201, n202, n208, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630;

  NAND2X0_HVT U5 ( .A1(n627), .A2(n345), .Y(n626) );
  NAND2X0_HVT U7 ( .A1(n350), .A2(n347), .Y(n623) );
  NAND2X0_HVT U9 ( .A1(n320), .A2(n622), .Y(n621) );
  NAND2X0_HVT U10 ( .A1(n320), .A2(n619), .Y(n620) );
  NAND2X0_HVT U11 ( .A1(n356), .A2(n348), .Y(n618) );
  NAND2X0_HVT U12 ( .A1(n352), .A2(n334), .Y(n617) );
  NAND2X0_HVT U13 ( .A1(n628), .A2(n622), .Y(n616) );
  NAND2X0_HVT U15 ( .A1(n291), .A2(n352), .Y(n614) );
  NAND2X0_HVT U19 ( .A1(n253), .A2(n420), .Y(n609) );
  NAND2X0_HVT U25 ( .A1(n230), .A2(n333), .Y(n625) );
  NAND2X0_HVT U32 ( .A1(n335), .A2(n356), .Y(n597) );
  NAND2X0_HVT U35 ( .A1(n622), .A2(n300), .Y(n594) );
  NAND2X0_HVT U38 ( .A1(n334), .A2(n356), .Y(n591) );
  NAND2X0_HVT U42 ( .A1(n624), .A2(n421), .Y(n587) );
  OA21X1_HVT U53 ( .A1(n197), .A2(n579), .A3(n390), .Y(n577) );
  NAND2X0_HVT U55 ( .A1(n346), .A2(n627), .Y(n575) );
  AO21X1_HVT U60 ( .A1(n569), .A2(n330), .A3(n608), .Y(n570) );
  MUX41X1_HVT U62 ( .A1(n568), .A3(n574), .A2(n572), .A4(n576), .S0(n341), 
        .S1(n338), .Y(n567) );
  NAND2X0_HVT U66 ( .A1(n277), .A2(n282), .Y(n563) );
  MUX41X1_HVT U67 ( .A1(n378), .A3(n403), .A2(n380), .A4(n563), .S0(n332), 
        .S1(n324), .Y(n562) );
  MUX41X1_HVT U71 ( .A1(n301), .A3(n318), .A2(n618), .A4(n374), .S0(n326), 
        .S1(n358), .Y(n559) );
  NAND2X0_HVT U72 ( .A1(n343), .A2(n623), .Y(n558) );
  MUX41X1_HVT U73 ( .A1(n602), .A3(n558), .A2(n404), .A4(n333), .S0(n331), 
        .S1(n323), .Y(n557) );
  MUX41X1_HVT U78 ( .A1(n553), .A3(n557), .A2(n556), .A4(n559), .S0(n341), 
        .S1(n338), .Y(n552) );
  MUX41X1_HVT U79 ( .A1(n391), .A3(n611), .A2(n393), .A4(n612), .S0(n327), 
        .S1(n360), .Y(n551) );
  MUX41X1_HVT U80 ( .A1(n406), .A3(n402), .A2(n621), .A4(n626), .S0(n326), 
        .S1(n361), .Y(n550) );
  NAND2X0_HVT U81 ( .A1(n219), .A2(n623), .Y(n549) );
  AND2X1_HVT U82 ( .A1(n301), .A2(n628), .Y(n548) );
  MUX41X1_HVT U84 ( .A1(n314), .A3(n391), .A2(n407), .A4(n604), .S0(n327), 
        .S1(n360), .Y(n546) );
  MUX41X1_HVT U88 ( .A1(n380), .A3(n365), .A2(n599), .A4(n583), .S0(n326), 
        .S1(n361), .Y(n543) );
  NAND2X0_HVT U89 ( .A1(n356), .A2(n418), .Y(n542) );
  MUX41X1_HVT U96 ( .A1(n403), .A3(n616), .A2(n389), .A4(n409), .S0(n327), 
        .S1(n361), .Y(n535) );
  MUX41X1_HVT U99 ( .A1(n597), .A3(n382), .A2(n581), .A4(n343), .S0(n270), 
        .S1(n324), .Y(n532) );
  NAND2X0_HVT U100 ( .A1(n356), .A2(n305), .Y(n531) );
  MUX41X1_HVT U101 ( .A1(n411), .A3(n617), .A2(n304), .A4(n531), .S0(n361), 
        .S1(n322), .Y(n530) );
  AND2X1_HVT U104 ( .A1(n623), .A2(n344), .Y(n528) );
  MUX41X1_HVT U105 ( .A1(n615), .A3(n412), .A2(n549), .A4(n528), .S0(n327), 
        .S1(n361), .Y(n527) );
  MUX41X1_HVT U107 ( .A1(n411), .A3(n346), .A2(n526), .A4(n371), .S0(n326), 
        .S1(n358), .Y(n525) );
  MUX41X1_HVT U108 ( .A1(n384), .A3(n342), .A2(n229), .A4(n349), .S0(n327), 
        .S1(n358), .Y(n524) );
  AO21X1_HVT U112 ( .A1(n398), .A2(n331), .A3(n605), .Y(n520) );
  NAND2X0_HVT U114 ( .A1(n316), .A2(n623), .Y(n518) );
  MUX41X1_HVT U115 ( .A1(n518), .A3(n618), .A2(n398), .A4(n346), .S0(n270), 
        .S1(n324), .Y(n517) );
  MUX41X1_HVT U116 ( .A1(n397), .A3(n391), .A2(n365), .A4(n614), .S0(n325), 
        .S1(n360), .Y(n516) );
  NAND2X0_HVT U118 ( .A1(n356), .A2(n307), .Y(n514) );
  MUX41X1_HVT U119 ( .A1(n413), .A3(n515), .A2(n592), .A4(n514), .S0(n325), 
        .S1(n360), .Y(n513) );
  MUX41X1_HVT U120 ( .A1(n513), .A3(n517), .A2(n516), .A4(n519), .S0(in[5]), 
        .S1(n338), .Y(n512) );
  MUX41X1_HVT U122 ( .A1(n401), .A3(n310), .A2(n583), .A4(n405), .S0(n325), 
        .S1(n361), .Y(n511) );
  MUX41X1_HVT U124 ( .A1(n312), .A3(n510), .A2(n606), .A4(n386), .S0(n330), 
        .S1(n325), .Y(n509) );
  AOI21X1_HVT U127 ( .A1(n329), .A2(n505), .A3(n372), .Y(n506) );
  NAND2X0_HVT U129 ( .A1(n328), .A2(n320), .Y(n503) );
  MUX41X1_HVT U130 ( .A1(n503), .A3(n504), .A2(n507), .A4(n506), .S0(n332), 
        .S1(n338), .Y(n502) );
  AND2X1_HVT U131 ( .A1(n282), .A2(n248), .Y(n501) );
  MUX41X1_HVT U132 ( .A1(n369), .A3(n501), .A2(n415), .A4(n378), .S0(n331), 
        .S1(n323), .Y(n500) );
  MUX41X1_HVT U133 ( .A1(n416), .A3(n371), .A2(n299), .A4(n370), .S0(n330), 
        .S1(n322), .Y(n499) );
  MUX41X1_HVT U136 ( .A1(n580), .A3(n531), .A2(n497), .A4(n376), .S0(n324), 
        .S1(n360), .Y(n496) );
  MUX41X1_HVT U140 ( .A1(n394), .A3(n311), .A2(n388), .A4(n618), .S0(n331), 
        .S1(n324), .Y(n493) );
  NAND2X0_HVT U141 ( .A1(n342), .A2(n356), .Y(n492) );
  MUX41X1_HVT U142 ( .A1(n492), .A3(n590), .A2(n414), .A4(n388), .S0(n329), 
        .S1(n358), .Y(n491) );
  MUX41X1_HVT U145 ( .A1(n598), .A3(n412), .A2(n489), .A4(n549), .S0(n329), 
        .S1(n358), .Y(n488) );
  AO21X1_HVT U148 ( .A1(n332), .A2(n373), .A3(n305), .Y(n485) );
  MUX41X1_HVT U151 ( .A1(n308), .A3(n396), .A2(n385), .A4(n483), .S0(n330), 
        .S1(n322), .Y(n482) );
  MUX41X1_HVT U155 ( .A1(n388), .A3(n618), .A2(n610), .A4(n389), .S0(n328), 
        .S1(n360), .Y(n478) );
  NAND2X0_HVT U159 ( .A1(n474), .A2(n473), .Y(n475) );
  MUX41X1_HVT U162 ( .A1(n256), .A3(n383), .A2(n594), .A4(n471), .S0(n328), 
        .S1(n358), .Y(n470) );
  NAND2X0_HVT U163 ( .A1(n268), .A2(n418), .Y(n469) );
  MUX41X1_HVT U164 ( .A1(n621), .A3(n469), .A2(n592), .A4(n384), .S0(n325), 
        .S1(n359), .Y(n468) );
  MUX41X1_HVT U172 ( .A1(n542), .A3(n460), .A2(n309), .A4(n607), .S0(n328), 
        .S1(n361), .Y(n459) );
  MUX41X1_HVT U173 ( .A1(n320), .A3(n318), .A2(n348), .A4(n593), .S0(n328), 
        .S1(n361), .Y(n458) );
  MUX41X1_HVT U175 ( .A1(n457), .A3(n458), .A2(n459), .A4(n461), .S0(n339), 
        .S1(n341), .Y(n456) );
  NAND2X0_HVT U177 ( .A1(n277), .A2(n307), .Y(n455) );
  MUX41X1_HVT U178 ( .A1(n313), .A3(n455), .A2(n317), .A4(n585), .S0(n328), 
        .S1(n360), .Y(n454) );
  AND2X1_HVT U179 ( .A1(n624), .A2(n344), .Y(n453) );
  MUX41X1_HVT U180 ( .A1(n597), .A3(n363), .A2(n453), .A4(n584), .S0(n328), 
        .S1(n359), .Y(n452) );
  MUX41X1_HVT U182 ( .A1(n371), .A3(n627), .A2(n368), .A4(n308), .S0(n325), 
        .S1(n358), .Y(n450) );
  MUX41X1_HVT U183 ( .A1(n399), .A3(n402), .A2(n384), .A4(n587), .S0(n330), 
        .S1(n323), .Y(n449) );
  AND2X1_HVT U185 ( .A1(n421), .A2(n248), .Y(n447) );
  MUX41X1_HVT U190 ( .A1(n444), .A3(n445), .A2(n443), .A4(n446), .S0(n339), 
        .S1(n323), .Y(n442) );
  NAND2X0_HVT U191 ( .A1(n302), .A2(n377), .Y(n441) );
  AND2X1_HVT U192 ( .A1(n395), .A2(n439), .Y(n440) );
  NAND2X0_HVT U194 ( .A1(n587), .A2(n439), .Y(n437) );
  NAND2X0_HVT U198 ( .A1(n354), .A2(n421), .Y(n619) );
  NAND2X0_HVT U200 ( .A1(n345), .A2(n356), .Y(n505) );
  NAND2X0_HVT U207 ( .A1(n356), .A2(n317), .Y(n569) );
  INVX0_HVT U1 ( .A(n335), .Y(n230) );
  INVX1_HVT U2 ( .A(n264), .Y(n196) );
  INVX1_HVT U3 ( .A(n196), .Y(n197) );
  MUX41X1_HVT U4 ( .A1(n441), .A3(n440), .A2(n437), .A4(n438), .S0(n198), .S1(
        n199), .Y(n436) );
  IBUFFX16_HVT U6 ( .A(n326), .Y(n198) );
  IBUFFX16_HVT U8 ( .A(n339), .Y(n199) );
  MUX41X1_HVT U14 ( .A1(n384), .A3(n394), .A2(n395), .A4(n620), .S0(n200), 
        .S1(n245), .Y(n556) );
  IBUFFX16_HVT U16 ( .A(n327), .Y(n200) );
  MUX21X2_HVT U17 ( .A1(n554), .A2(n555), .S0(n201), .Y(n553) );
  IBUFFX16_HVT U18 ( .A(n329), .Y(n201) );
  MUX21X2_HVT U20 ( .A1(n405), .A2(n364), .S0(n332), .Y(n555) );
  NAND2X0_HVT U21 ( .A1(n538), .A2(n202), .Y(n208) );
  NAND2X0_HVT U22 ( .A1(n539), .A2(n238), .Y(n218) );
  NAND2X0_HVT U23 ( .A1(n208), .A2(n218), .Y(n537) );
  INVX0_HVT U24 ( .A(n238), .Y(n202) );
  IBUFFX2_HVT U26 ( .A(n257), .Y(n238) );
  INVX2_HVT U27 ( .A(n347), .Y(n420) );
  NAND2X2_HVT U28 ( .A1(n293), .A2(n294), .Y(n613) );
  XNOR2X2_HVT U29 ( .A1(n197), .A2(n325), .Y(n315) );
  MUX21X1_HVT U30 ( .A1(n384), .A2(n566), .S0(n315), .Y(n565) );
  NBUFFX2_HVT U31 ( .A(n419), .Y(n333) );
  OR2X1_HVT U33 ( .A1(n295), .A2(n292), .Y(n219) );
  MUX21X1_HVT U34 ( .A1(n387), .A2(n573), .S0(n315), .Y(n572) );
  MUX21X2_HVT U36 ( .A1(n454), .A2(n452), .S0(n337), .Y(n451) );
  MUX21X1_HVT U37 ( .A1(n336), .A2(n291), .S0(n267), .Y(n604) );
  MUX21X1_HVT U39 ( .A1(n307), .A2(n417), .S0(n220), .Y(n606) );
  IBUFFX16_HVT U40 ( .A(n277), .Y(n220) );
  INVX0_HVT U41 ( .A(n607), .Y(n385) );
  NAND2X0_HVT U43 ( .A1(n449), .A2(n221), .Y(n222) );
  NAND2X0_HVT U44 ( .A1(n450), .A2(n339), .Y(n223) );
  NAND2X0_HVT U45 ( .A1(n222), .A2(n223), .Y(n448) );
  IBUFFX2_HVT U46 ( .A(n339), .Y(n221) );
  INVX1_HVT U47 ( .A(n337), .Y(n339) );
  MUX21X2_HVT U48 ( .A1(n627), .A2(n385), .S0(n278), .Y(n566) );
  MUX41X2_HVT U49 ( .A1(n313), .A3(n309), .A2(n312), .A4(n462), .S0(n328), 
        .S1(n359), .Y(n461) );
  INVX0_HVT U50 ( .A(n606), .Y(n386) );
  MUX21X1_HVT U51 ( .A1(n476), .A2(n475), .S0(n224), .Y(n472) );
  INVX1_HVT U52 ( .A(n331), .Y(n264) );
  AO21X1_HVT U54 ( .A1(n254), .A2(n305), .A3(n264), .Y(n439) );
  AO21X1_HVT U56 ( .A1(n248), .A2(n316), .A3(n264), .Y(n473) );
  IBUFFX16_HVT U57 ( .A(n329), .Y(n224) );
  NAND2X0_HVT U58 ( .A1(n230), .A2(n225), .Y(n226) );
  NAND2X0_HVT U59 ( .A1(n348), .A2(n254), .Y(n227) );
  NAND2X0_HVT U61 ( .A1(n226), .A2(n227), .Y(n229) );
  IBUFFX2_HVT U63 ( .A(n254), .Y(n225) );
  INVX0_HVT U64 ( .A(n229), .Y(n603) );
  MUX41X1_HVT U65 ( .A1(n392), .A3(n548), .A2(n549), .A4(n308), .S0(n228), 
        .S1(n358), .Y(n547) );
  IBUFFX16_HVT U68 ( .A(n326), .Y(n228) );
  INVX1_HVT U69 ( .A(n348), .Y(n305) );
  NAND2X0_HVT U70 ( .A1(n343), .A2(n231), .Y(n232) );
  NAND2X0_HVT U74 ( .A1(n374), .A2(n269), .Y(n233) );
  NAND2X0_HVT U75 ( .A1(n232), .A2(n233), .Y(n538) );
  INVX0_HVT U76 ( .A(n269), .Y(n231) );
  INVX1_HVT U77 ( .A(n332), .Y(n269) );
  MUX41X1_HVT U83 ( .A1(n470), .A3(n472), .A2(n464), .A4(n468), .S0(n339), 
        .S1(n234), .Y(n463) );
  IBUFFX16_HVT U85 ( .A(n341), .Y(n234) );
  INVX0_HVT U86 ( .A(n332), .Y(n249) );
  INVX0_HVT U87 ( .A(n332), .Y(n302) );
  MUX21X1_HVT U90 ( .A1(n389), .A2(n379), .S0(n332), .Y(n578) );
  NAND2X0_HVT U91 ( .A1(n346), .A2(n235), .Y(n236) );
  NAND2X0_HVT U92 ( .A1(n540), .A2(n244), .Y(n237) );
  NAND2X0_HVT U93 ( .A1(n236), .A2(n237), .Y(n539) );
  INVX0_HVT U94 ( .A(n244), .Y(n235) );
  IBUFFX2_HVT U95 ( .A(n254), .Y(n244) );
  NBUFFX2_HVT U97 ( .A(n628), .Y(n347) );
  IBUFFX2_HVT U98 ( .A(n623), .Y(n372) );
  INVX0_HVT U102 ( .A(n335), .Y(n240) );
  INVX1_HVT U103 ( .A(n429), .Y(n408) );
  MUX41X1_HVT U106 ( .A1(n314), .A3(n368), .A2(n229), .A4(n408), .S0(n239), 
        .S1(n360), .Y(n544) );
  IBUFFX16_HVT U109 ( .A(n325), .Y(n239) );
  OR2X1_HVT U110 ( .A1(n334), .A2(n240), .Y(n630) );
  IBUFFX2_HVT U111 ( .A(n334), .Y(n307) );
  MUX41X1_HVT U113 ( .A1(n550), .A3(n546), .A2(n551), .A4(n547), .S0(n241), 
        .S1(n338), .Y(n545) );
  IBUFFX16_HVT U117 ( .A(n341), .Y(n241) );
  INVX1_HVT U121 ( .A(n592), .Y(n396) );
  IBUFFX2_HVT U123 ( .A(n612), .Y(n380) );
  MUX41X1_HVT U125 ( .A1(n537), .A3(n541), .A2(n543), .A4(n544), .S0(n242), 
        .S1(n243), .Y(n536) );
  IBUFFX16_HVT U126 ( .A(n337), .Y(n242) );
  IBUFFX16_HVT U128 ( .A(n340), .Y(n243) );
  INVX0_HVT U134 ( .A(n358), .Y(n245) );
  MUX21X1_HVT U135 ( .A1(n604), .A2(n314), .S0(n331), .Y(n481) );
  MUX21X2_HVT U137 ( .A1(n536), .A2(n529), .S0(n255), .Y(out[2]) );
  MUX21X2_HVT U138 ( .A1(n601), .A2(n396), .S0(n246), .Y(n272) );
  IBUFFX16_HVT U139 ( .A(n322), .Y(n246) );
  MUX41X1_HVT U143 ( .A1(n533), .A3(n530), .A2(n535), .A4(n532), .S0(n340), 
        .S1(n247), .Y(n529) );
  IBUFFX16_HVT U144 ( .A(n337), .Y(n247) );
  OA21X1_HVT U146 ( .A1(n367), .A2(n302), .A3(n608), .Y(n554) );
  MUX21X2_HVT U147 ( .A1(n271), .A2(n272), .S0(n361), .Y(n533) );
  XOR2X2_HVT U149 ( .A1(n320), .A2(n252), .Y(n592) );
  INVX1_HVT U150 ( .A(n351), .Y(n248) );
  INVX1_HVT U152 ( .A(n355), .Y(n351) );
  MUX21X2_HVT U153 ( .A1(n410), .A2(n534), .S0(n278), .Y(n271) );
  XOR2X2_HVT U154 ( .A1(n344), .A2(n352), .Y(n581) );
  NAND2X0_HVT U156 ( .A1(n372), .A2(n269), .Y(n250) );
  NAND2X0_HVT U157 ( .A1(n588), .A2(n332), .Y(n251) );
  NAND2X0_HVT U158 ( .A1(n250), .A2(n251), .Y(n521) );
  NBUFFX2_HVT U160 ( .A(n351), .Y(n252) );
  NBUFFX2_HVT U161 ( .A(n351), .Y(n253) );
  NBUFFX2_HVT U165 ( .A(n351), .Y(n254) );
  INVX2_HVT U166 ( .A(in[0]), .Y(n355) );
  INVX1_HVT U167 ( .A(n355), .Y(n352) );
  INVX1_HVT U168 ( .A(n248), .Y(n353) );
  NAND2X0_HVT U169 ( .A1(n567), .A2(n273), .Y(n274) );
  INVX0_HVT U170 ( .A(n256), .Y(n585) );
  INVX0_HVT U171 ( .A(n304), .Y(n593) );
  INVX1_HVT U174 ( .A(n608), .Y(n384) );
  OA21X1_HVT U176 ( .A1(n366), .A2(n264), .A3(n375), .Y(n480) );
  INVX1_HVT U181 ( .A(n327), .Y(n278) );
  INVX1_HVT U184 ( .A(in[1]), .Y(n337) );
  INVX1_HVT U186 ( .A(n323), .Y(n257) );
  INVX1_HVT U187 ( .A(in[7]), .Y(n255) );
  INVX1_HVT U188 ( .A(n255), .Y(n273) );
  INVX1_HVT U189 ( .A(in[6]), .Y(n306) );
  INVX1_HVT U193 ( .A(in[5]), .Y(n340) );
  MUX21X1_HVT U195 ( .A1(n282), .A2(n420), .S0(n352), .Y(n588) );
  MUX21X1_HVT U196 ( .A1(n292), .A2(n613), .S0(n276), .Y(n304) );
  INVX1_HVT U197 ( .A(n276), .Y(n356) );
  INVX0_HVT U199 ( .A(n355), .Y(n276) );
  MUX21X1_HVT U201 ( .A1(n344), .A2(n321), .S0(n353), .Y(n256) );
  MUX21X1_HVT U202 ( .A1(n319), .A2(n418), .S0(n277), .Y(n601) );
  IBUFFX2_HVT U203 ( .A(n601), .Y(n390) );
  NAND2X0_HVT U204 ( .A1(n466), .A2(n257), .Y(n258) );
  NAND2X0_HVT U205 ( .A1(n467), .A2(n324), .Y(n259) );
  NAND2X0_HVT U206 ( .A1(n258), .A2(n259), .Y(n464) );
  NAND2X0_HVT U208 ( .A1(n456), .A2(n255), .Y(n260) );
  NAND2X0_HVT U209 ( .A1(n463), .A2(n273), .Y(n261) );
  NAND2X0_HVT U210 ( .A1(n260), .A2(n261), .Y(out[6]) );
  NAND2X0_HVT U211 ( .A1(n619), .A2(n465), .Y(n466) );
  MUX21X1_HVT U212 ( .A1(n603), .A2(n606), .S0(n330), .Y(n467) );
  NAND2X0_HVT U213 ( .A1(n314), .A2(n197), .Y(n262) );
  NAND2X0_HVT U214 ( .A1(n581), .A2(n332), .Y(n263) );
  NAND2X0_HVT U215 ( .A1(n262), .A2(n263), .Y(n445) );
  INVX1_HVT U216 ( .A(n370), .Y(n301) );
  NAND2X0_HVT U217 ( .A1(n404), .A2(n197), .Y(n265) );
  NAND2X0_HVT U218 ( .A1(n588), .A2(n331), .Y(n266) );
  NAND2X0_HVT U219 ( .A1(n265), .A2(n266), .Y(n444) );
  INVX0_HVT U220 ( .A(n433), .Y(n404) );
  MUX21X1_HVT U221 ( .A1(n613), .A2(n334), .S0(n350), .Y(n608) );
  INVX0_HVT U222 ( .A(n276), .Y(n267) );
  INVX1_HVT U223 ( .A(n267), .Y(n268) );
  MUX21X1_HVT U224 ( .A1(n335), .A2(n333), .S0(n267), .Y(n584) );
  OR2X1_HVT U225 ( .A1(n267), .A2(n418), .Y(n622) );
  IBUFFX2_HVT U226 ( .A(n355), .Y(n277) );
  AO21X1_HVT U227 ( .A1(n342), .A2(n627), .A3(n302), .Y(n465) );
  INVX2_HVT U228 ( .A(n362), .Y(n359) );
  IBUFFX4_HVT U229 ( .A(n362), .Y(n358) );
  IBUFFX2_HVT U230 ( .A(n362), .Y(n361) );
  MUX21X2_HVT U231 ( .A1(n512), .A2(n522), .S0(in[7]), .Y(out[3]) );
  MUX21X2_HVT U232 ( .A1(n495), .A2(n496), .S0(n339), .Y(n494) );
  INVX1_HVT U233 ( .A(n249), .Y(n270) );
  IBUFFX2_HVT U234 ( .A(n362), .Y(n360) );
  MUX21X2_HVT U235 ( .A1(n477), .A2(n487), .S0(n273), .Y(out[5]) );
  MUX41X1_HVT U236 ( .A1(n383), .A3(n591), .A2(n381), .A4(n382), .S0(n270), 
        .S1(n278), .Y(n564) );
  NAND2X0_HVT U237 ( .A1(n560), .A2(n255), .Y(n275) );
  NAND2X0_HVT U238 ( .A1(n274), .A2(n275), .Y(out[0]) );
  MUX41X1_HVT U239 ( .A1(n317), .A3(n582), .A2(n623), .A4(n542), .S0(n270), 
        .S1(n326), .Y(n541) );
  IBUFFX2_HVT U240 ( .A(n584), .Y(n400) );
  INVX0_HVT U241 ( .A(n604), .Y(n388) );
  MUX21X2_HVT U242 ( .A1(n545), .A2(n552), .S0(in[7]), .Y(out[1]) );
  MUX41X1_HVT U243 ( .A1(n564), .A3(n561), .A2(n565), .A4(n562), .S0(n340), 
        .S1(n338), .Y(n560) );
  INVX1_HVT U244 ( .A(n340), .Y(n341) );
  NBUFFX2_HVT U245 ( .A(n419), .Y(n334) );
  OA21X1_HVT U246 ( .A1(n391), .A2(n197), .A3(n569), .Y(n443) );
  NBUFFX2_HVT U247 ( .A(n306), .Y(n335) );
  INVX1_HVT U248 ( .A(n615), .Y(n378) );
  MUX21X1_HVT U249 ( .A1(n414), .A2(n311), .S0(n324), .Y(n507) );
  INVX1_HVT U250 ( .A(n283), .Y(n523) );
  INVX0_HVT U251 ( .A(n365), .Y(n284) );
  MUX21X1_HVT U252 ( .A1(n613), .A2(n336), .S0(n331), .Y(n540) );
  INVX1_HVT U253 ( .A(n630), .Y(n319) );
  INVX0_HVT U254 ( .A(n319), .Y(n316) );
  INVX1_HVT U255 ( .A(n316), .Y(n318) );
  INVX1_HVT U256 ( .A(n316), .Y(n317) );
  OR2X1_HVT U257 ( .A1(n334), .A2(n306), .Y(n628) );
  INVX0_HVT U258 ( .A(n333), .Y(n295) );
  INVX0_HVT U259 ( .A(n303), .Y(n462) );
  INVX1_HVT U260 ( .A(in[4]), .Y(n362) );
  IBUFFX2_HVT U261 ( .A(n355), .Y(n354) );
  MUX21X1_HVT U262 ( .A1(n318), .A2(n336), .S0(n353), .Y(n460) );
  NAND2X0_HVT U263 ( .A1(n447), .A2(n302), .Y(n279) );
  NAND2X0_HVT U264 ( .A1(n406), .A2(n330), .Y(n280) );
  NAND2X0_HVT U265 ( .A1(n279), .A2(n280), .Y(n446) );
  INVX1_HVT U266 ( .A(n431), .Y(n406) );
  MUX41X1_HVT U267 ( .A1(n575), .A3(n229), .A2(n281), .A4(n402), .S0(n257), 
        .S1(n249), .Y(n574) );
  MUX41X1_HVT U268 ( .A1(n321), .A3(n379), .A2(n307), .A4(n378), .S0(n278), 
        .S1(n302), .Y(n561) );
  NAND2X0_HVT U269 ( .A1(n293), .A2(n294), .Y(n281) );
  INVX1_HVT U270 ( .A(n306), .Y(n282) );
  INVX1_HVT U271 ( .A(n291), .Y(n421) );
  INVX1_HVT U272 ( .A(n281), .Y(n300) );
  MUX41X1_HVT U273 ( .A1(n583), .A3(n430), .A2(n284), .A4(n427), .S0(n257), 
        .S1(n269), .Y(n283) );
  INVX0_HVT U274 ( .A(n306), .Y(n292) );
  MUX21X1_HVT U275 ( .A1(n321), .A2(n219), .S0(n353), .Y(n615) );
  INVX1_HVT U276 ( .A(n298), .Y(n299) );
  NAND2X0_HVT U277 ( .A1(n276), .A2(n629), .Y(n627) );
  MUX41X1_HVT U278 ( .A1(n527), .A3(n524), .A2(n525), .A4(n523), .S0(n340), 
        .S1(n337), .Y(n522) );
  NAND2X0_HVT U279 ( .A1(n386), .A2(n269), .Y(n285) );
  NAND2X0_HVT U280 ( .A1(n575), .A2(n331), .Y(n286) );
  NAND2X0_HVT U281 ( .A1(n285), .A2(n286), .Y(n571) );
  MUX21X1_HVT U282 ( .A1(n571), .A2(n570), .S0(n328), .Y(n568) );
  NAND2X0_HVT U283 ( .A1(n520), .A2(n257), .Y(n289) );
  NAND2X0_HVT U284 ( .A1(n586), .A2(n249), .Y(n287) );
  NAND2X0_HVT U285 ( .A1(n405), .A2(n331), .Y(n288) );
  NAND2X0_HVT U286 ( .A1(n287), .A2(n288), .Y(n476) );
  MUX21X1_HVT U287 ( .A1(n334), .A2(n420), .S0(n350), .Y(n586) );
  INVX1_HVT U288 ( .A(n432), .Y(n405) );
  NAND2X0_HVT U289 ( .A1(n521), .A2(n329), .Y(n290) );
  NAND2X0_HVT U290 ( .A1(n289), .A2(n290), .Y(n519) );
  NAND2X0_HVT U291 ( .A1(n293), .A2(n294), .Y(n291) );
  MUX41X1_HVT U292 ( .A1(n300), .A3(n416), .A2(n299), .A4(n408), .S0(n278), 
        .S1(n249), .Y(n457) );
  NAND2X0_HVT U293 ( .A1(n306), .A2(n333), .Y(n293) );
  NAND2X0_HVT U294 ( .A1(n292), .A2(in[3]), .Y(n294) );
  MUX41X1_HVT U295 ( .A1(n448), .A3(n436), .A2(n451), .A4(n442), .S0(n255), 
        .S1(n341), .Y(out[7]) );
  OR2X1_HVT U296 ( .A1(n295), .A2(n292), .Y(n629) );
  NAND2X0_HVT U297 ( .A1(n499), .A2(n337), .Y(n296) );
  NAND2X0_HVT U298 ( .A1(n500), .A2(n338), .Y(n297) );
  NAND2X0_HVT U299 ( .A1(n296), .A2(n297), .Y(n498) );
  INVX0_HVT U300 ( .A(n575), .Y(n298) );
  NAND2X0_HVT U301 ( .A1(n252), .A2(n630), .Y(n624) );
  MUX41X1_HVT U302 ( .A1(n409), .A3(n604), .A2(n600), .A4(n622), .S0(n249), 
        .S1(n257), .Y(n495) );
  MUX41X1_HVT U303 ( .A1(n491), .A3(n493), .A2(n488), .A4(n490), .S0(n339), 
        .S1(n340), .Y(n487) );
  INVX1_HVT U304 ( .A(n319), .Y(n321) );
  MUX41X1_HVT U305 ( .A1(n484), .A3(n479), .A2(n482), .A4(n478), .S0(n340), 
        .S1(n337), .Y(n477) );
  INVX1_HVT U306 ( .A(n319), .Y(n320) );
  MUX21X1_HVT U307 ( .A1(n346), .A2(n316), .S0(n267), .Y(n303) );
  INVX1_HVT U308 ( .A(n424), .Y(n414) );
  NBUFFX2_HVT U309 ( .A(n629), .Y(n348) );
  INVX1_HVT U310 ( .A(n348), .Y(n417) );
  INVX0_HVT U311 ( .A(n587), .Y(n371) );
  MUX41X1_HVT U312 ( .A1(n508), .A3(n502), .A2(n498), .A4(n494), .S0(n340), 
        .S1(n255), .Y(out[4]) );
  NBUFFX2_HVT U313 ( .A(n306), .Y(n336) );
  MUX21X1_HVT U314 ( .A1(n417), .A2(n421), .S0(n248), .Y(n607) );
  INVX1_HVT U315 ( .A(n596), .Y(n394) );
  MUX21X2_HVT U316 ( .A1(n509), .A2(n511), .S0(n339), .Y(n508) );
  MUX41X1_HVT U317 ( .A1(n606), .A3(n609), .A2(n399), .A4(n418), .S0(n257), 
        .S1(n269), .Y(n490) );
  INVX0_HVT U318 ( .A(in[3]), .Y(n419) );
  MUX21X1_HVT U319 ( .A1(n281), .A2(n295), .S0(n248), .Y(n308) );
  IBUFFX2_HVT U320 ( .A(n355), .Y(n350) );
  MUX21X2_HVT U321 ( .A1(n415), .A2(n369), .S0(n330), .Y(n486) );
  MUX21X2_HVT U322 ( .A1(n486), .A2(n485), .S0(n324), .Y(n484) );
  MUX21X2_HVT U323 ( .A1(n480), .A2(n481), .S0(n329), .Y(n479) );
  MUX21X2_HVT U324 ( .A1(n578), .A2(n577), .S0(n328), .Y(n576) );
  NBUFFX2_HVT U325 ( .A(n629), .Y(n349) );
  AND2X1_HVT U326 ( .A1(n301), .A2(n219), .Y(n309) );
  AND2X1_HVT U327 ( .A1(n349), .A2(n614), .Y(n310) );
  MUX21X1_HVT U328 ( .A1(n400), .A2(n312), .S0(n330), .Y(n438) );
  MUX21X1_HVT U329 ( .A1(n344), .A2(n346), .S0(n277), .Y(n471) );
  MUX21X1_HVT U330 ( .A1(n421), .A2(n333), .S0(n268), .Y(n590) );
  MUX21X1_HVT U331 ( .A1(n417), .A2(n300), .S0(n353), .Y(n596) );
  MUX21X1_HVT U332 ( .A1(n417), .A2(n335), .S0(n353), .Y(n433) );
  MUX21X1_HVT U333 ( .A1(n306), .A2(n418), .S0(n352), .Y(n483) );
  MUX21X1_HVT U334 ( .A1(n300), .A2(n336), .S0(n354), .Y(n424) );
  MUX21X1_HVT U335 ( .A1(n336), .A2(n349), .S0(n354), .Y(n526) );
  MUX21X1_HVT U336 ( .A1(n317), .A2(n342), .S0(n352), .Y(n429) );
  MUX21X1_HVT U337 ( .A1(n333), .A2(n305), .S0(n254), .Y(n599) );
  MUX21X1_HVT U338 ( .A1(n596), .A2(n310), .S0(n329), .Y(n504) );
  XOR2X1_HVT U339 ( .A1(n613), .A2(n276), .Y(n583) );
  MUX21X1_HVT U340 ( .A1(n306), .A2(n343), .S0(n277), .Y(n589) );
  MUX21X1_HVT U341 ( .A1(n291), .A2(n317), .S0(n354), .Y(n598) );
  MUX21X1_HVT U342 ( .A1(n281), .A2(n418), .S0(n350), .Y(n595) );
  MUX21X1_HVT U343 ( .A1(n420), .A2(n334), .S0(n354), .Y(n432) );
  XNOR2X1_HVT U344 ( .A1(n219), .A2(n350), .Y(n311) );
  INVX1_HVT U345 ( .A(n625), .Y(n418) );
  MUX21X1_HVT U346 ( .A1(n347), .A2(n349), .S0(n268), .Y(n611) );
  MUX21X1_HVT U347 ( .A1(n305), .A2(n420), .S0(n354), .Y(n579) );
  MUX21X1_HVT U348 ( .A1(n344), .A2(n349), .S0(n353), .Y(n423) );
  MUX21X1_HVT U349 ( .A1(n334), .A2(n349), .S0(n277), .Y(n431) );
  MUX21X1_HVT U350 ( .A1(n347), .A2(n333), .S0(n268), .Y(n610) );
  XOR2X1_HVT U351 ( .A1(n347), .A2(n277), .Y(n582) );
  AND2X1_HVT U352 ( .A1(n253), .A2(n336), .Y(n312) );
  MUX21X1_HVT U353 ( .A1(n333), .A2(n346), .S0(n277), .Y(n426) );
  NBUFFX2_HVT U354 ( .A(n359), .Y(n331) );
  NBUFFX2_HVT U355 ( .A(n359), .Y(n330) );
  NBUFFX2_HVT U356 ( .A(n359), .Y(n332) );
  NBUFFX2_HVT U357 ( .A(n613), .Y(n342) );
  NBUFFX2_HVT U358 ( .A(n613), .Y(n343) );
  MUX21X1_HVT U359 ( .A1(n346), .A2(n335), .S0(n352), .Y(n510) );
  AND2X1_HVT U360 ( .A1(n420), .A2(n356), .Y(n313) );
  MUX21X1_HVT U361 ( .A1(n388), .A2(n626), .S0(n329), .Y(n573) );
  MUX21X1_HVT U362 ( .A1(n349), .A2(n345), .S0(n350), .Y(n489) );
  NBUFFX2_HVT U363 ( .A(n625), .Y(n344) );
  NBUFFX2_HVT U364 ( .A(n628), .Y(n346) );
  AND2X1_HVT U365 ( .A1(n628), .A2(n356), .Y(n314) );
  NBUFFX2_HVT U366 ( .A(n625), .Y(n345) );
  NBUFFX2_HVT U367 ( .A(n357), .Y(n328) );
  NBUFFX2_HVT U368 ( .A(n357), .Y(n329) );
  NBUFFX2_HVT U369 ( .A(n357), .Y(n325) );
  NBUFFX2_HVT U370 ( .A(n357), .Y(n327) );
  NBUFFX2_HVT U371 ( .A(n322), .Y(n326) );
  NBUFFX2_HVT U372 ( .A(in[2]), .Y(n323) );
  NBUFFX2_HVT U373 ( .A(n357), .Y(n324) );
  NBUFFX2_HVT U374 ( .A(n357), .Y(n322) );
  INVX1_HVT U375 ( .A(n337), .Y(n338) );
  MUX21X1_HVT U376 ( .A1(n318), .A2(n307), .S0(n350), .Y(n422) );
  MUX21X1_HVT U377 ( .A1(n321), .A2(n307), .S0(n352), .Y(n474) );
  MUX21X1_HVT U378 ( .A1(n345), .A2(n307), .S0(n354), .Y(n534) );
  MUX21X1_HVT U379 ( .A1(n420), .A2(n418), .S0(n253), .Y(n515) );
  MUX21X1_HVT U380 ( .A1(n336), .A2(n307), .S0(n276), .Y(n602) );
  MUX21X1_HVT U381 ( .A1(n307), .A2(n321), .S0(n354), .Y(n428) );
  MUX21X1_HVT U382 ( .A1(n307), .A2(n345), .S0(n354), .Y(n427) );
  NBUFFX2_HVT U383 ( .A(in[2]), .Y(n357) );
  MUX21X1_HVT U384 ( .A1(n417), .A2(n282), .S0(n253), .Y(n497) );
  XOR2X1_HVT U385 ( .A1(n268), .A2(n292), .Y(n580) );
  MUX21X1_HVT U386 ( .A1(n282), .A2(n346), .S0(n353), .Y(n434) );
  MUX21X1_HVT U387 ( .A1(n346), .A2(n282), .S0(n352), .Y(n430) );
  MUX21X1_HVT U388 ( .A1(n333), .A2(n282), .S0(n353), .Y(n425) );
  MUX21X1_HVT U389 ( .A1(n282), .A2(n320), .S0(n353), .Y(n612) );
  MUX21X1_HVT U390 ( .A1(n282), .A2(n317), .S0(n350), .Y(n605) );
  MUX21X1_HVT U391 ( .A1(n345), .A2(n282), .S0(n350), .Y(n600) );
  MUX21X1_HVT U392 ( .A1(n282), .A2(n418), .S0(n352), .Y(n435) );
  INVX0_HVT U393 ( .A(n618), .Y(n363) );
  INVX0_HVT U394 ( .A(n597), .Y(n364) );
  INVX0_HVT U395 ( .A(n591), .Y(n365) );
  INVX0_HVT U396 ( .A(n531), .Y(n366) );
  INVX0_HVT U397 ( .A(n492), .Y(n367) );
  INVX0_HVT U398 ( .A(n627), .Y(n368) );
  INVX0_HVT U399 ( .A(n626), .Y(n369) );
  INVX0_HVT U400 ( .A(n624), .Y(n370) );
  INVX0_HVT U401 ( .A(n622), .Y(n373) );
  INVX0_HVT U402 ( .A(n594), .Y(n374) );
  INVX0_HVT U403 ( .A(n616), .Y(n375) );
  INVX0_HVT U404 ( .A(n621), .Y(n376) );
  INVX0_HVT U405 ( .A(n617), .Y(n377) );
  INVX0_HVT U406 ( .A(n614), .Y(n379) );
  INVX0_HVT U407 ( .A(n611), .Y(n381) );
  INVX0_HVT U408 ( .A(n610), .Y(n382) );
  INVX0_HVT U409 ( .A(n609), .Y(n383) );
  INVX0_HVT U410 ( .A(n605), .Y(n387) );
  INVX0_HVT U411 ( .A(n602), .Y(n389) );
  INVX0_HVT U412 ( .A(n600), .Y(n391) );
  INVX0_HVT U413 ( .A(n599), .Y(n392) );
  INVX0_HVT U414 ( .A(n598), .Y(n393) );
  INVX0_HVT U415 ( .A(n595), .Y(n395) );
  INVX0_HVT U416 ( .A(n590), .Y(n397) );
  INVX0_HVT U417 ( .A(n589), .Y(n398) );
  INVX0_HVT U418 ( .A(n586), .Y(n399) );
  INVX0_HVT U419 ( .A(n620), .Y(n401) );
  INVX0_HVT U420 ( .A(n435), .Y(n402) );
  INVX0_HVT U421 ( .A(n434), .Y(n403) );
  INVX0_HVT U422 ( .A(n430), .Y(n407) );
  INVX0_HVT U423 ( .A(n428), .Y(n409) );
  INVX0_HVT U424 ( .A(n427), .Y(n410) );
  INVX0_HVT U425 ( .A(n426), .Y(n411) );
  INVX0_HVT U426 ( .A(n425), .Y(n412) );
  INVX0_HVT U427 ( .A(n474), .Y(n413) );
  INVX0_HVT U428 ( .A(n423), .Y(n415) );
  INVX0_HVT U429 ( .A(n422), .Y(n416) );
endmodule

