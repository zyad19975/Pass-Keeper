
module keygen ( round_num, keyin, keyout );
  input [0:3] round_num;
  input [0:127] keyin;
  output [0:127] keyout;
  wire   n283, n284, n3, n4, n286, n285, n290, n289, n288, n287, n293, n292,
         n291, n29, n31, n32, n33, n34, n35, n36, n37, n38, n40, n41, n42, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n62, n63, n65, n67, n68, n69, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n108, n109, n110, n111, n112, n113, n115, n117, n118, n1, n2,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n39, n43, n61, n64,
         n66, n70, n71, n84, n107, n114, n116, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n149,
         n151, n153, n154, n155, n157, n160, n162, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n204, n205, n206, n207, n208, n209, n210, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n246, n247, n248, n249,
         n250, n251, n252, n253, n255, n256, n257, n259, n260, n261, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282;
  wire   [0:31] dummy;

  sbox_0 a1 ( .in({keyin[104:106], n194, n196, keyin[109], n220, keyin[111]}), 
        .out(dummy[0:7]) );
  sbox_19 a2 ( .in({n165, keyin[113:119]}), .out(dummy[8:15]) );
  sbox_18 a3 ( .in({n157, n170, keyin[122:123], n200, keyin[125], n255, 
        keyin[127]}), .out(dummy[16:23]) );
  sbox_17 a4 ( .in({n209, n166, keyin[98], n232, keyin[100:103]}), .out(
        dummy[24:31]) );
  XOR2X2_HVT U66 ( .A1(dummy[3]), .A2(keyin[3]), .Y(n38) );
  XNOR2X2_HVT U84 ( .A1(dummy[27]), .A2(keyin[27]), .Y(n95) );
  XNOR2X2_HVT U94 ( .A1(dummy[22]), .A2(keyin[22]), .Y(n100) );
  XNOR2X2_HVT U96 ( .A1(dummy[21]), .A2(keyin[21]), .Y(n101) );
  XNOR2X2_HVT U100 ( .A1(dummy[19]), .A2(keyin[19]), .Y(n103) );
  XNOR2X2_HVT U102 ( .A1(dummy[18]), .A2(keyin[18]), .Y(n104) );
  XNOR2X2_HVT U120 ( .A1(dummy[9]), .A2(keyin[9]), .Y(n80) );
  XOR2X2_HVT U136 ( .A1(dummy[0]), .A2(keyin[0]), .Y(n45) );
  INVX0_HVT U165 ( .A(n87), .Y(n29) );
  INVX0_HVT U167 ( .A(n85), .Y(n31) );
  INVX0_HVT U169 ( .A(n86), .Y(n33) );
  XNOR3X1_HVT U176 ( .A1(keyin[70]), .A2(n1), .A3(n273), .Y(keyout[70]) );
  XNOR3X1_HVT U178 ( .A1(keyin[68]), .A2(n74), .A3(n131), .Y(keyout[68]) );
  XNOR3X1_HVT U179 ( .A1(keyin[32]), .A2(keyin[64]), .A3(n76), .Y(n46) );
  NAND3X0_HVT U180 ( .A1(n86), .A2(n87), .A3(n88), .Y(n82) );
  AO21X1_HVT U182 ( .A1(n92), .A2(round_num[2]), .A3(n33), .Y(n89) );
  XNOR3X1_HVT U196 ( .A1(n59), .A2(n249), .A3(n103), .Y(keyout[115]) );
  AND2X1_HVT U210 ( .A1(n87), .A2(n115), .Y(n72) );
  AND2X1_HVT U213 ( .A1(n86), .A2(n117), .Y(n78) );
  NAND2X0_HVT U215 ( .A1(round_num[2]), .A2(n118), .Y(n86) );
  AO21X1_HVT U217 ( .A1(n92), .A2(n35), .A3(n29), .Y(n79) );
  NAND2X0_HVT U218 ( .A1(round_num[0]), .A2(n113), .Y(n87) );
  NAND2X0_HVT U221 ( .A1(n118), .A2(n35), .Y(n76) );
  INVX1_HVT U1 ( .A(n206), .Y(n157) );
  XOR2X1_HVT U2 ( .A1(dummy[30]), .A2(n190), .Y(n91) );
  XOR2X1_HVT U3 ( .A1(dummy[11]), .A2(n197), .Y(n111) );
  NBUFFX2_HVT U4 ( .A(keyin[108]), .Y(n196) );
  XOR2X1_HVT U5 ( .A1(dummy[26]), .A2(n256), .Y(n114) );
  NBUFFX2_HVT U6 ( .A(keyin[124]), .Y(n200) );
  XNOR2X1_HVT U7 ( .A1(n9), .A2(n269), .Y(keyout[2]) );
  INVX1_HVT U8 ( .A(n89), .Y(n9) );
  XNOR2X1_HVT U9 ( .A1(n276), .A2(n14), .Y(keyout[76]) );
  NBUFFX2_HVT U10 ( .A(keyin[100]), .Y(n149) );
  XOR2X1_HVT U11 ( .A1(dummy[17]), .A2(keyin[17]), .Y(n264) );
  INVX1_HVT U12 ( .A(n77), .Y(n3) );
  INVX1_HVT U13 ( .A(n109), .Y(n225) );
  INVX1_HVT U14 ( .A(n111), .Y(n286) );
  NBUFFX2_HVT U15 ( .A(keyin[107]), .Y(n194) );
  NBUFFX2_HVT U16 ( .A(keyin[110]), .Y(n220) );
  INVX0_HVT U17 ( .A(n255), .Y(n201) );
  XNOR2X1_HVT U18 ( .A1(n293), .A2(n207), .Y(keyout[93]) );
  XNOR2X1_HVT U19 ( .A1(keyout[13]), .A2(n228), .Y(keyout[77]) );
  XOR2X1_HVT U20 ( .A1(n111), .A2(n281), .Y(keyout[75]) );
  XNOR2X1_HVT U21 ( .A1(n94), .A2(keyin[60]), .Y(keyout[60]) );
  XNOR2X1_HVT U22 ( .A1(dummy[28]), .A2(keyin[28]), .Y(n94) );
  XOR2X1_HVT U23 ( .A1(n250), .A2(n63), .Y(keyout[79]) );
  INVX1_HVT U24 ( .A(n78), .Y(n2) );
  XOR3X1_HVT U25 ( .A1(n49), .A2(n204), .A3(n93), .Y(keyout[125]) );
  INVX0_HVT U26 ( .A(keyin[125]), .Y(n204) );
  INVX1_HVT U27 ( .A(n250), .Y(n244) );
  INVX1_HVT U28 ( .A(n271), .Y(n202) );
  INVX1_HVT U29 ( .A(n103), .Y(keyout[19]) );
  INVX1_HVT U30 ( .A(n104), .Y(keyout[18]) );
  INVX1_HVT U31 ( .A(n95), .Y(keyout[27]) );
  INVX1_HVT U32 ( .A(n284), .Y(n146) );
  DELLN1X2_HVT U33 ( .A(keyin[104]), .Y(n247) );
  XNOR3X1_HVT U34 ( .A1(n67), .A2(n194), .A3(n111), .Y(keyout[107]) );
  DELLN1X2_HVT U35 ( .A(n196), .Y(n141) );
  XOR3X1_HVT U36 ( .A1(n60), .A2(n195), .A3(n104), .Y(keyout[114]) );
  NBUFFX2_HVT U37 ( .A(keyin[115]), .Y(n249) );
  DELLN1X2_HVT U38 ( .A(keyin[116]), .Y(n186) );
  DELLN1X2_HVT U39 ( .A(keyin[117]), .Y(n154) );
  INVX1_HVT U40 ( .A(n206), .Y(n11) );
  INVX1_HVT U41 ( .A(n54), .Y(n10) );
  INVX0_HVT U42 ( .A(n200), .Y(n21) );
  XOR2X1_HVT U43 ( .A1(n72), .A2(keyin[38]), .Y(n1) );
  INVX1_HVT U44 ( .A(n98), .Y(n291) );
  XNOR3X1_HVT U45 ( .A1(n65), .A2(keyin[109]), .A3(n109), .Y(keyout[109]) );
  XNOR2X1_HVT U46 ( .A1(n77), .A2(n2), .Y(keyout[5]) );
  NAND2X0_HVT U47 ( .A1(n283), .A2(n251), .Y(n6) );
  NAND2X0_HVT U48 ( .A1(n5), .A2(keyin[32]), .Y(n7) );
  NAND2X0_HVT U49 ( .A1(n6), .A2(n7), .Y(keyout[32]) );
  INVX0_HVT U50 ( .A(n283), .Y(n5) );
  XNOR2X2_HVT U51 ( .A1(n1), .A2(n273), .Y(keyout[38]) );
  XOR2X1_HVT U52 ( .A1(dummy[15]), .A2(keyin[15]), .Y(n250) );
  XNOR2X1_HVT U53 ( .A1(n77), .A2(n8), .Y(keyout[101]) );
  XNOR2X1_HVT U54 ( .A1(n85), .A2(n268), .Y(n8) );
  INVX1_HVT U55 ( .A(n73), .Y(n4) );
  XNOR2X2_HVT U56 ( .A1(n98), .A2(n54), .Y(keyout[88]) );
  XOR3X2_HVT U57 ( .A1(n10), .A2(n11), .A3(n98), .Y(keyout[120]) );
  XNOR2X1_HVT U58 ( .A1(n273), .A2(n72), .Y(keyout[6]) );
  XOR2X1_HVT U59 ( .A1(n143), .A2(n74), .Y(keyout[36]) );
  XOR2X1_HVT U60 ( .A1(n82), .A2(n38), .Y(keyout[3]) );
  NBUFFX2_HVT U61 ( .A(keyin[99]), .Y(n232) );
  XOR2X1_HVT U62 ( .A1(n270), .A2(n64), .Y(keyout[97]) );
  INVX0_HVT U63 ( .A(n102), .Y(n289) );
  XOR2X1_HVT U64 ( .A1(n37), .A2(n38), .Y(keyout[35]) );
  XOR3X2_HVT U65 ( .A1(keyin[68]), .A2(n149), .A3(n282), .Y(keyout[100]) );
  XOR2X1_HVT U67 ( .A1(n273), .A2(n179), .Y(keyout[102]) );
  INVX1_HVT U68 ( .A(n73), .Y(n143) );
  XNOR2X2_HVT U69 ( .A1(n44), .A2(n270), .Y(keyout[65]) );
  INVX1_HVT U70 ( .A(n191), .Y(n171) );
  XOR2X1_HVT U71 ( .A1(n230), .A2(n47), .Y(keyout[95]) );
  XOR2X2_HVT U72 ( .A1(n45), .A2(n46), .Y(keyout[64]) );
  XNOR2X1_HVT U73 ( .A1(n97), .A2(n53), .Y(keyout[89]) );
  XOR2X1_HVT U74 ( .A1(dummy[25]), .A2(n130), .Y(n97) );
  INVX0_HVT U75 ( .A(n97), .Y(n127) );
  INVX1_HVT U76 ( .A(n106), .Y(n287) );
  INVX1_HVT U77 ( .A(round_num[2]), .Y(n35) );
  INVX1_HVT U78 ( .A(keyin[13]), .Y(n172) );
  XOR2X1_HVT U79 ( .A1(dummy[12]), .A2(keyin[12]), .Y(n276) );
  INVX1_HVT U80 ( .A(round_num[0]), .Y(n32) );
  INVX1_HVT U81 ( .A(round_num[1]), .Y(n34) );
  INVX1_HVT U82 ( .A(round_num[3]), .Y(n36) );
  NBUFFX2_HVT U83 ( .A(keyin[126]), .Y(n255) );
  INVX1_HVT U85 ( .A(keyin[23]), .Y(n218) );
  INVX1_HVT U86 ( .A(n75), .Y(n17) );
  INVX1_HVT U87 ( .A(n65), .Y(n228) );
  XOR2X1_HVT U88 ( .A1(dummy[26]), .A2(n256), .Y(n96) );
  INVX1_HVT U89 ( .A(n49), .Y(n207) );
  NBUFFX2_HVT U90 ( .A(keyin[96]), .Y(n209) );
  INVX1_HVT U91 ( .A(keyin[5]), .Y(n184) );
  XNOR2X1_HVT U92 ( .A1(n120), .A2(keyin[39]), .Y(n119) );
  INVX1_HVT U93 ( .A(keyin[16]), .Y(n246) );
  INVX1_HVT U95 ( .A(keyin[24]), .Y(n133) );
  XOR3X1_HVT U97 ( .A1(n241), .A2(n242), .A3(n243), .Y(keyout[111]) );
  INVX1_HVT U98 ( .A(keyin[111]), .Y(n242) );
  INVX1_HVT U99 ( .A(n63), .Y(n241) );
  XNOR2X1_HVT U101 ( .A1(n99), .A2(n55), .Y(keyout[87]) );
  XNOR2X1_HVT U103 ( .A1(n264), .A2(n12), .Y(keyout[81]) );
  INVX1_HVT U104 ( .A(keyin[44]), .Y(n153) );
  XOR2X1_HVT U105 ( .A1(n250), .A2(keyin[47]), .Y(keyout[47]) );
  XNOR2X1_HVT U106 ( .A1(n104), .A2(n60), .Y(keyout[82]) );
  INVX1_HVT U107 ( .A(n96), .Y(keyout[26]) );
  INVX1_HVT U108 ( .A(n109), .Y(keyout[13]) );
  XNOR2X1_HVT U109 ( .A1(n229), .A2(n267), .Y(keyout[40]) );
  INVX1_HVT U110 ( .A(keyin[40]), .Y(n267) );
  XNOR2X1_HVT U111 ( .A1(keyin[41]), .A2(n80), .Y(keyout[41]) );
  XNOR2X1_HVT U112 ( .A1(n108), .A2(keyin[46]), .Y(keyout[46]) );
  INVX1_HVT U113 ( .A(keyin[20]), .Y(n176) );
  XNOR2X1_HVT U114 ( .A1(keyin[53]), .A2(n101), .Y(keyout[53]) );
  INVX1_HVT U115 ( .A(keyin[63]), .Y(n180) );
  XNOR2X1_HVT U116 ( .A1(n81), .A2(n223), .Y(keyout[72]) );
  INVX1_HVT U117 ( .A(n16), .Y(n223) );
  XNOR2X1_HVT U118 ( .A1(n112), .A2(n68), .Y(keyout[74]) );
  XNOR2X1_HVT U119 ( .A1(n100), .A2(n56), .Y(keyout[86]) );
  XNOR2X1_HVT U121 ( .A1(n96), .A2(n52), .Y(keyout[90]) );
  XNOR2X1_HVT U122 ( .A1(n95), .A2(n51), .Y(keyout[91]) );
  XOR2X1_HVT U123 ( .A1(n1), .A2(n208), .Y(n179) );
  XOR3X1_HVT U124 ( .A1(keyin[71]), .A2(n132), .A3(n119), .Y(keyout[103]) );
  INVX1_HVT U125 ( .A(keyin[103]), .Y(n132) );
  INVX1_HVT U126 ( .A(keyin[106]), .Y(n168) );
  INVX1_HVT U127 ( .A(n68), .Y(n167) );
  INVX1_HVT U128 ( .A(keyin[114]), .Y(n195) );
  XOR3X1_HVT U129 ( .A1(n58), .A2(n231), .A3(n102), .Y(keyout[116]) );
  INVX1_HVT U130 ( .A(n186), .Y(n231) );
  INVX1_HVT U131 ( .A(keyin[122]), .Y(n257) );
  AND3X1_HVT U132 ( .A1(n34), .A2(n36), .A3(round_num[0]), .Y(n118) );
  AND3X1_HVT U133 ( .A1(n34), .A2(n35), .A3(round_num[3]), .Y(n113) );
  AND3X1_HVT U134 ( .A1(n32), .A2(n36), .A3(round_num[1]), .Y(n92) );
  INVX1_HVT U135 ( .A(keyin[4]), .Y(n189) );
  NAND4X0_HVT U137 ( .A1(round_num[1]), .A2(round_num[2]), .A3(round_num[3]), 
        .A4(n32), .Y(n75) );
  INVX1_HVT U138 ( .A(keyin[7]), .Y(n252) );
  INVX1_HVT U139 ( .A(n113), .Y(n253) );
  INVX1_HVT U140 ( .A(keyin[26]), .Y(n256) );
  NBUFFX2_HVT U141 ( .A(n42), .Y(n269) );
  NAND4X0_HVT U142 ( .A1(round_num[1]), .A2(round_num[3]), .A3(n32), .A4(n35), 
        .Y(n88) );
  NAND4X0_HVT U143 ( .A1(round_num[2]), .A2(round_num[3]), .A3(n32), .A4(n34), 
        .Y(n117) );
  NAND3X0_HVT U144 ( .A1(n34), .A2(n36), .A3(round_num[2]), .Y(n115) );
  XOR2X1_HVT U145 ( .A1(n79), .A2(keyin[36]), .Y(n74) );
  XNOR2X1_HVT U146 ( .A1(n185), .A2(n221), .Y(n105) );
  INVX1_HVT U147 ( .A(keyin[14]), .Y(n265) );
  INVX0_HVT U148 ( .A(n93), .Y(n293) );
  INVX1_HVT U149 ( .A(keyin[25]), .Y(n130) );
  INVX1_HVT U150 ( .A(keyin[98]), .Y(n274) );
  INVX1_HVT U151 ( .A(n74), .Y(n142) );
  INVX1_HVT U152 ( .A(keyin[11]), .Y(n197) );
  NBUFFX2_HVT U153 ( .A(keyin[112]), .Y(n165) );
  XNOR2X1_HVT U154 ( .A1(n285), .A2(n272), .Y(keyout[73]) );
  INVX1_HVT U155 ( .A(n69), .Y(n272) );
  XNOR2X1_HVT U156 ( .A1(n219), .A2(n264), .Y(keyout[49]) );
  XOR3X1_HVT U157 ( .A1(n55), .A2(keyin[119]), .A3(n290), .Y(keyout[119]) );
  INVX1_HVT U158 ( .A(keyin[45]), .Y(n224) );
  INVX1_HVT U159 ( .A(n105), .Y(keyout[17]) );
  XNOR3X1_HVT U160 ( .A1(n69), .A2(keyin[105]), .A3(n80), .Y(keyout[105]) );
  XOR3X1_HVT U161 ( .A1(keyin[66]), .A2(n41), .A3(n27), .Y(keyout[66]) );
  INVX1_HVT U162 ( .A(n91), .Y(keyout[30]) );
  INVX1_HVT U163 ( .A(keyin[32]), .Y(n251) );
  INVX1_HVT U164 ( .A(keyin[56]), .Y(n136) );
  XOR3X1_HVT U166 ( .A1(n46), .A2(n209), .A3(n24), .Y(keyout[96]) );
  INVX1_HVT U168 ( .A(n274), .Y(n216) );
  XOR3X1_HVT U170 ( .A1(n15), .A2(n220), .A3(n108), .Y(keyout[110]) );
  XOR3X1_HVT U171 ( .A1(n51), .A2(n61), .A3(n95), .Y(keyout[123]) );
  XOR3X1_HVT U172 ( .A1(n50), .A2(n21), .A3(n116), .Y(keyout[124]) );
  XNOR2X1_HVT U173 ( .A1(keyin[49]), .A2(keyin[81]), .Y(n12) );
  INVX0_HVT U174 ( .A(n103), .Y(n288) );
  INVX0_HVT U175 ( .A(n114), .Y(n71) );
  XOR2X1_HVT U177 ( .A1(keyin[69]), .A2(n31), .Y(n13) );
  INVX1_HVT U181 ( .A(keyin[17]), .Y(n221) );
  XNOR2X1_HVT U183 ( .A1(keyin[44]), .A2(keyin[76]), .Y(n14) );
  XNOR2X1_HVT U184 ( .A1(keyin[46]), .A2(keyin[78]), .Y(n15) );
  XNOR2X1_HVT U185 ( .A1(keyin[40]), .A2(keyin[72]), .Y(n16) );
  INVX1_HVT U186 ( .A(keyin[10]), .Y(n210) );
  INVX1_HVT U187 ( .A(n50), .Y(n275) );
  INVX1_HVT U188 ( .A(n59), .Y(n188) );
  INVX1_HVT U189 ( .A(keyin[31]), .Y(n239) );
  IBUFFX2_HVT U190 ( .A(keyin[123]), .Y(n61) );
  XNOR2X2_HVT U191 ( .A1(n276), .A2(n153), .Y(keyout[44]) );
  INVX0_HVT U192 ( .A(n91), .Y(n30) );
  XNOR2X2_HVT U193 ( .A1(dummy[20]), .A2(keyin[20]), .Y(n102) );
  XOR3X2_HVT U194 ( .A1(n56), .A2(n240), .A3(n100), .Y(keyout[118]) );
  INVX0_HVT U195 ( .A(n160), .Y(n155) );
  XOR3X1_HVT U197 ( .A1(n53), .A2(n170), .A3(n160), .Y(keyout[121]) );
  INVX1_HVT U198 ( .A(dummy[1]), .Y(n191) );
  INVX0_HVT U199 ( .A(n42), .Y(n137) );
  XOR2X2_HVT U200 ( .A1(dummy[8]), .A2(n266), .Y(n81) );
  XNOR2X2_HVT U201 ( .A1(n18), .A2(n17), .Y(n164) );
  NAND2X0_HVT U202 ( .A1(n192), .A2(n193), .Y(n18) );
  XNOR3X1_HVT U203 ( .A1(n57), .A2(n154), .A3(n101), .Y(keyout[117]) );
  INVX1_HVT U204 ( .A(n225), .Y(n19) );
  XOR3X1_HVT U205 ( .A1(n16), .A2(n247), .A3(n81), .Y(keyout[104]) );
  XOR3X2_HVT U206 ( .A1(n37), .A2(n20), .A3(n38), .Y(keyout[99]) );
  XOR2X1_HVT U207 ( .A1(keyin[67]), .A2(n232), .Y(n20) );
  XOR2X1_HVT U208 ( .A1(dummy[8]), .A2(keyin[8]), .Y(n229) );
  INVX1_HVT U209 ( .A(n263), .Y(n22) );
  XOR2X1_HVT U211 ( .A1(dummy[10]), .A2(n210), .Y(n112) );
  INVX0_HVT U212 ( .A(n45), .Y(n23) );
  INVX1_HVT U214 ( .A(n23), .Y(n24) );
  INVX0_HVT U216 ( .A(dummy[10]), .Y(n25) );
  XNOR2X1_HVT U219 ( .A1(keyin[12]), .A2(dummy[12]), .Y(n110) );
  INVX0_HVT U220 ( .A(n100), .Y(keyout[22]) );
  INVX0_HVT U222 ( .A(dummy[17]), .Y(n185) );
  INVX1_HVT U223 ( .A(n25), .Y(n26) );
  INVX1_HVT U224 ( .A(n137), .Y(n27) );
  NAND2X0_HVT U225 ( .A1(keyin[62]), .A2(n91), .Y(n39) );
  NAND2X0_HVT U226 ( .A1(n28), .A2(n30), .Y(n43) );
  NAND2X0_HVT U227 ( .A1(n39), .A2(n43), .Y(keyout[62]) );
  INVX0_HVT U228 ( .A(keyin[62]), .Y(n28) );
  INVX1_HVT U229 ( .A(n116), .Y(n292) );
  XNOR2X2_HVT U230 ( .A1(n91), .A2(n48), .Y(keyout[94]) );
  XOR3X1_HVT U231 ( .A1(n48), .A2(n201), .A3(n91), .Y(keyout[126]) );
  XOR2X1_HVT U232 ( .A1(n66), .A2(keyin[97]), .Y(n64) );
  INVX1_HVT U233 ( .A(n44), .Y(n66) );
  INVX0_HVT U234 ( .A(n164), .Y(keyout[1]) );
  NAND2X0_HVT U235 ( .A1(keyin[58]), .A2(n114), .Y(n84) );
  NAND2X0_HVT U236 ( .A1(n70), .A2(n71), .Y(n107) );
  NAND2X0_HVT U237 ( .A1(n84), .A2(n107), .Y(keyout[58]) );
  INVX0_HVT U238 ( .A(keyin[58]), .Y(n70) );
  XNOR2X2_HVT U239 ( .A1(dummy[29]), .A2(keyin[29]), .Y(n93) );
  XNOR2X2_HVT U240 ( .A1(dummy[28]), .A2(keyin[28]), .Y(n116) );
  XOR3X2_HVT U241 ( .A1(n252), .A2(n253), .A3(dummy[7]), .Y(n120) );
  NAND2X0_HVT U242 ( .A1(keyin[54]), .A2(n100), .Y(n123) );
  NAND2X0_HVT U243 ( .A1(n121), .A2(n122), .Y(n124) );
  NAND2X0_HVT U244 ( .A1(n123), .A2(n124), .Y(keyout[54]) );
  INVX0_HVT U245 ( .A(keyin[54]), .Y(n121) );
  INVX0_HVT U246 ( .A(n100), .Y(n122) );
  XOR2X1_HVT U247 ( .A1(dummy[4]), .A2(n189), .Y(n131) );
  INVX0_HVT U248 ( .A(n119), .Y(keyout[39]) );
  XOR2X1_HVT U249 ( .A1(dummy[20]), .A2(n176), .Y(n125) );
  NAND2X0_HVT U250 ( .A1(keyin[57]), .A2(n97), .Y(n128) );
  NAND2X0_HVT U251 ( .A1(n127), .A2(n126), .Y(n129) );
  NAND2X0_HVT U252 ( .A1(n128), .A2(n129), .Y(keyout[57]) );
  INVX0_HVT U253 ( .A(keyin[57]), .Y(n126) );
  INVX0_HVT U254 ( .A(dummy[31]), .Y(n233) );
  XOR3X1_HVT U255 ( .A1(n167), .A2(n168), .A3(n263), .Y(keyout[106]) );
  XOR2X2_HVT U256 ( .A1(n171), .A2(keyin[1]), .Y(n270) );
  XOR2X2_HVT U257 ( .A1(dummy[24]), .A2(n133), .Y(n98) );
  XNOR3X1_HVT U258 ( .A1(n62), .A2(n165), .A3(n106), .Y(keyout[112]) );
  XNOR2X2_HVT U259 ( .A1(dummy[10]), .A2(n210), .Y(n263) );
  INVX1_HVT U260 ( .A(n278), .Y(keyout[11]) );
  XNOR2X2_HVT U261 ( .A1(keyin[59]), .A2(n95), .Y(keyout[59]) );
  XNOR2X2_HVT U262 ( .A1(n83), .A2(keyin[71]), .Y(keyout[71]) );
  NBUFFX2_HVT U263 ( .A(n276), .Y(keyout[12]) );
  XNOR2X2_HVT U264 ( .A1(n136), .A2(n291), .Y(keyout[56]) );
  NAND2X0_HVT U265 ( .A1(n41), .A2(n42), .Y(n139) );
  NAND2X0_HVT U266 ( .A1(n137), .A2(n138), .Y(n140) );
  NAND2X0_HVT U267 ( .A1(n139), .A2(n140), .Y(n40) );
  INVX0_HVT U268 ( .A(n41), .Y(n138) );
  XOR3X2_HVT U269 ( .A1(n216), .A2(n217), .A3(n40), .Y(keyout[98]) );
  NAND2X0_HVT U270 ( .A1(n131), .A2(n74), .Y(n144) );
  NAND2X0_HVT U271 ( .A1(n143), .A2(n142), .Y(n145) );
  NAND2X0_HVT U272 ( .A1(n144), .A2(n145), .Y(n282) );
  XOR3X2_HVT U273 ( .A1(n14), .A2(n141), .A3(n110), .Y(keyout[108]) );
  XNOR2X2_HVT U274 ( .A1(keyin[50]), .A2(n104), .Y(keyout[50]) );
  XNOR2X2_HVT U275 ( .A1(n125), .A2(keyin[52]), .Y(keyout[52]) );
  INVX1_HVT U276 ( .A(keyin[49]), .Y(n219) );
  XNOR2X2_HVT U277 ( .A1(n106), .A2(keyin[48]), .Y(keyout[48]) );
  INVX1_HVT U278 ( .A(n146), .Y(keyout[7]) );
  INVX1_HVT U279 ( .A(n261), .Y(n240) );
  OR2X1_HVT U280 ( .A1(keyin[33]), .A2(n164), .Y(n260) );
  XNOR2X2_HVT U281 ( .A1(n101), .A2(n57), .Y(keyout[85]) );
  IBUFFX2_HVT U282 ( .A(n101), .Y(keyout[21]) );
  NBUFFX2_HVT U283 ( .A(n290), .Y(keyout[23]) );
  INVX1_HVT U284 ( .A(keyin[55]), .Y(n198) );
  XNOR2X1_HVT U285 ( .A1(keyin[51]), .A2(n103), .Y(keyout[51]) );
  INVX0_HVT U286 ( .A(n229), .Y(n151) );
  INVX1_HVT U287 ( .A(n151), .Y(keyout[8]) );
  INVX1_HVT U288 ( .A(n155), .Y(keyout[25]) );
  XOR2X1_HVT U289 ( .A1(dummy[25]), .A2(keyin[25]), .Y(n160) );
  INVX1_HVT U290 ( .A(n212), .Y(keyout[28]) );
  INVX1_HVT U291 ( .A(n292), .Y(n212) );
  XNOR2X1_HVT U292 ( .A1(n26), .A2(n210), .Y(keyout[10]) );
  INVX0_HVT U293 ( .A(n236), .Y(keyout[16]) );
  INVX1_HVT U294 ( .A(n287), .Y(n236) );
  INVX1_HVT U295 ( .A(n293), .Y(n162) );
  INVX1_HVT U296 ( .A(n162), .Y(keyout[29]) );
  XOR3X1_HVT U297 ( .A1(n52), .A2(n257), .A3(n114), .Y(keyout[122]) );
  OR2X1_HVT U298 ( .A1(keyin[1]), .A2(n191), .Y(n192) );
  INVX1_HVT U299 ( .A(keyin[66]), .Y(n217) );
  INVX1_HVT U300 ( .A(keyin[15]), .Y(n205) );
  INVX1_HVT U301 ( .A(keyin[30]), .Y(n190) );
  INVX1_HVT U302 ( .A(n215), .Y(n166) );
  INVX1_HVT U303 ( .A(keyin[97]), .Y(n215) );
  INVX1_HVT U304 ( .A(keyin[121]), .Y(n169) );
  INVX1_HVT U305 ( .A(n169), .Y(n170) );
  INVX1_HVT U306 ( .A(keyin[120]), .Y(n206) );
  XNOR3X1_HVT U307 ( .A1(n47), .A2(keyin[127]), .A3(n90), .Y(keyout[127]) );
  XOR2X2_HVT U308 ( .A1(dummy[13]), .A2(n172), .Y(n109) );
  NAND2X0_HVT U309 ( .A1(n289), .A2(n187), .Y(n174) );
  NAND2X0_HVT U310 ( .A1(n173), .A2(n58), .Y(n175) );
  NAND2X0_HVT U311 ( .A1(n174), .A2(n175), .Y(keyout[84]) );
  INVX0_HVT U312 ( .A(n289), .Y(n173) );
  INVX1_HVT U313 ( .A(n58), .Y(n187) );
  INVX1_HVT U314 ( .A(n99), .Y(n290) );
  NBUFFX2_HVT U315 ( .A(n230), .Y(keyout[31]) );
  NAND2X0_HVT U316 ( .A1(n233), .A2(n239), .Y(n178) );
  XOR3X1_HVT U317 ( .A1(n12), .A2(keyin[113]), .A3(n105), .Y(keyout[113]) );
  XNOR2X2_HVT U318 ( .A1(n180), .A2(n230), .Y(keyout[63]) );
  NAND2X0_HVT U319 ( .A1(n288), .A2(n188), .Y(n182) );
  NAND2X0_HVT U320 ( .A1(n181), .A2(n59), .Y(n183) );
  NAND2X0_HVT U321 ( .A1(n183), .A2(n182), .Y(keyout[83]) );
  INVX0_HVT U322 ( .A(n288), .Y(n181) );
  XOR2X2_HVT U323 ( .A1(dummy[5]), .A2(n184), .Y(n77) );
  XOR2X2_HVT U324 ( .A1(dummy[4]), .A2(n189), .Y(n73) );
  NAND2X0_HVT U325 ( .A1(n191), .A2(keyin[1]), .Y(n193) );
  XNOR2X2_HVT U326 ( .A1(n22), .A2(keyin[42]), .Y(keyout[42]) );
  XNOR2X2_HVT U327 ( .A1(n198), .A2(n290), .Y(keyout[55]) );
  DELLN2X2_HVT U328 ( .A(keyin[102]), .Y(n199) );
  INVX1_HVT U329 ( .A(n202), .Y(keyout[14]) );
  XNOR2X1_HVT U330 ( .A1(n205), .A2(dummy[15]), .Y(n243) );
  XOR3X1_HVT U331 ( .A1(keyin[67]), .A2(n37), .A3(n38), .Y(keyout[67]) );
  XNOR2X1_HVT U332 ( .A1(keyin[70]), .A2(n199), .Y(n208) );
  INVX1_HVT U333 ( .A(n98), .Y(keyout[24]) );
  XNOR2X2_HVT U334 ( .A1(dummy[14]), .A2(keyin[14]), .Y(n108) );
  INVX1_HVT U335 ( .A(n5), .Y(keyout[0]) );
  XOR2X2_HVT U336 ( .A1(dummy[2]), .A2(keyin[2]), .Y(n42) );
  NAND2X0_HVT U337 ( .A1(n292), .A2(n275), .Y(n213) );
  NAND2X0_HVT U338 ( .A1(n212), .A2(n50), .Y(n214) );
  NAND2X0_HVT U339 ( .A1(n214), .A2(n213), .Y(keyout[92]) );
  XOR2X2_HVT U340 ( .A1(dummy[23]), .A2(n218), .Y(n99) );
  XNOR2X2_HVT U341 ( .A1(keyin[61]), .A2(n93), .Y(keyout[61]) );
  XOR2X2_HVT U342 ( .A1(n4), .A2(n79), .Y(keyout[4]) );
  NBUFFX2_HVT U343 ( .A(n285), .Y(keyout[9]) );
  INVX1_HVT U344 ( .A(n80), .Y(n285) );
  XOR2X2_HVT U345 ( .A1(n3), .A2(n85), .Y(keyout[37]) );
  NAND2X0_HVT U346 ( .A1(keyin[45]), .A2(n19), .Y(n226) );
  NAND2X0_HVT U347 ( .A1(n224), .A2(n225), .Y(n227) );
  NAND2X0_HVT U348 ( .A1(n226), .A2(n227), .Y(keyout[45]) );
  INVX1_HVT U349 ( .A(keyin[8]), .Y(n266) );
  AND2X1_HVT U350 ( .A1(n178), .A2(n235), .Y(n230) );
  NAND2X0_HVT U351 ( .A1(n233), .A2(n239), .Y(n234) );
  NAND2X0_HVT U352 ( .A1(dummy[31]), .A2(keyin[31]), .Y(n235) );
  NAND2X0_HVT U353 ( .A1(n234), .A2(n235), .Y(n90) );
  NAND2X0_HVT U354 ( .A1(n287), .A2(n248), .Y(n237) );
  NAND2X0_HVT U355 ( .A1(n236), .A2(n62), .Y(n238) );
  NAND2X0_HVT U356 ( .A1(n237), .A2(n238), .Y(keyout[80]) );
  INVX1_HVT U357 ( .A(n62), .Y(n248) );
  INVX1_HVT U358 ( .A(n244), .Y(keyout[15]) );
  XOR2X2_HVT U359 ( .A1(dummy[16]), .A2(n246), .Y(n106) );
  XOR2X2_HVT U360 ( .A1(n41), .A2(n269), .Y(keyout[34]) );
  XOR3X2_HVT U361 ( .A1(n252), .A2(n253), .A3(dummy[7]), .Y(n284) );
  XOR2X2_HVT U362 ( .A1(dummy[6]), .A2(keyin[6]), .Y(n273) );
  XNOR2X2_HVT U363 ( .A1(dummy[14]), .A2(n265), .Y(n271) );
  NBUFFX2_HVT U364 ( .A(n289), .Y(keyout[20]) );
  XNOR2X2_HVT U365 ( .A1(n284), .A2(keyin[39]), .Y(n83) );
  NAND2X0_HVT U366 ( .A1(keyin[33]), .A2(n164), .Y(n259) );
  NAND2X0_HVT U367 ( .A1(n260), .A2(n259), .Y(keyout[33]) );
  DELLN2X2_HVT U368 ( .A(keyin[118]), .Y(n261) );
  XNOR2X1_HVT U369 ( .A1(keyin[69]), .A2(keyin[101]), .Y(n268) );
  XNOR2X2_HVT U370 ( .A1(n271), .A2(n15), .Y(keyout[78]) );
  XNOR2X2_HVT U371 ( .A1(n3), .A2(n13), .Y(keyout[69]) );
  XNOR2X2_HVT U372 ( .A1(n45), .A2(n76), .Y(n283) );
  INVX1_HVT U373 ( .A(n67), .Y(n281) );
  INVX1_HVT U374 ( .A(keyin[43]), .Y(n277) );
  NAND2X0_HVT U375 ( .A1(keyin[43]), .A2(n278), .Y(n279) );
  NAND2X0_HVT U376 ( .A1(n277), .A2(n286), .Y(n280) );
  NAND2X0_HVT U377 ( .A1(n279), .A2(n280), .Y(keyout[43]) );
  INVX0_HVT U378 ( .A(n286), .Y(n278) );
  XOR2X1_HVT U379 ( .A1(n82), .A2(keyin[35]), .Y(n37) );
  XOR2X1_HVT U380 ( .A1(n89), .A2(keyin[34]), .Y(n41) );
  XNOR2X1_HVT U381 ( .A1(n78), .A2(keyin[37]), .Y(n85) );
  XOR3X1_HVT U382 ( .A1(keyin[65]), .A2(keyin[33]), .A3(n75), .Y(n44) );
  XOR2X1_HVT U383 ( .A1(keyin[41]), .A2(keyin[73]), .Y(n69) );
  XOR2X1_HVT U384 ( .A1(keyin[42]), .A2(keyin[74]), .Y(n68) );
  XOR2X1_HVT U385 ( .A1(keyin[45]), .A2(keyin[77]), .Y(n65) );
  XOR2X1_HVT U386 ( .A1(keyin[47]), .A2(keyin[79]), .Y(n63) );
  XOR2X1_HVT U387 ( .A1(keyin[50]), .A2(keyin[82]), .Y(n60) );
  XOR2X1_HVT U388 ( .A1(keyin[51]), .A2(keyin[83]), .Y(n59) );
  XOR2X1_HVT U389 ( .A1(keyin[52]), .A2(keyin[84]), .Y(n58) );
  XOR2X1_HVT U390 ( .A1(keyin[53]), .A2(keyin[85]), .Y(n57) );
  XOR2X1_HVT U391 ( .A1(keyin[54]), .A2(keyin[86]), .Y(n56) );
  XOR2X1_HVT U392 ( .A1(keyin[55]), .A2(keyin[87]), .Y(n55) );
  XOR2X1_HVT U393 ( .A1(keyin[57]), .A2(keyin[89]), .Y(n53) );
  XOR2X1_HVT U394 ( .A1(keyin[58]), .A2(keyin[90]), .Y(n52) );
  XOR2X1_HVT U395 ( .A1(keyin[59]), .A2(keyin[91]), .Y(n51) );
  XOR2X1_HVT U396 ( .A1(keyin[60]), .A2(keyin[92]), .Y(n50) );
  XOR2X1_HVT U397 ( .A1(keyin[61]), .A2(keyin[93]), .Y(n49) );
  XOR2X1_HVT U398 ( .A1(keyin[62]), .A2(keyin[94]), .Y(n48) );
  XOR2X1_HVT U399 ( .A1(keyin[63]), .A2(keyin[95]), .Y(n47) );
  XOR2X1_HVT U400 ( .A1(keyin[43]), .A2(keyin[75]), .Y(n67) );
  XOR2X1_HVT U401 ( .A1(keyin[48]), .A2(keyin[80]), .Y(n62) );
  XOR2X1_HVT U402 ( .A1(keyin[56]), .A2(keyin[88]), .Y(n54) );
endmodule

