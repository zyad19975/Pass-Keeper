
module sbox_13 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n3, n23, n50, n121, n210, n211, n212, n213, n216, n217, n218, n219,
         n224, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582;

  NAND2X0_HVT U4 ( .A1(n579), .A2(n240), .Y(n580) );
  NAND2X0_HVT U5 ( .A1(n298), .A2(n281), .Y(n578) );
  NAND2X0_HVT U13 ( .A1(n570), .A2(n294), .Y(n571) );
  NAND2X0_HVT U15 ( .A1(n239), .A2(n283), .Y(n568) );
  NAND2X0_HVT U21 ( .A1(n293), .A2(n302), .Y(n562) );
  NAND2X0_HVT U24 ( .A1(n289), .A2(n302), .Y(n560) );
  NAND2X0_HVT U33 ( .A1(n360), .A2(n302), .Y(n551) );
  NAND2X0_HVT U35 ( .A1(n286), .A2(n302), .Y(n549) );
  NAND2X0_HVT U42 ( .A1(n296), .A2(n288), .Y(n542) );
  MUX41X1_HVT U51 ( .A1(n349), .A3(n309), .A2(n326), .A4(n327), .S0(n306), 
        .S1(n303), .Y(n534) );
  NAND2X0_HVT U53 ( .A1(n531), .A2(n541), .Y(n532) );
  NAND2X0_HVT U56 ( .A1(n293), .A2(n527), .Y(n528) );
  MUX41X1_HVT U57 ( .A1(n350), .A3(n564), .A2(n528), .A4(n573), .S0(n306), 
        .S1(n275), .Y(n526) );
  NAND2X0_HVT U58 ( .A1(n294), .A2(n240), .Y(n525) );
  MUX41X1_HVT U59 ( .A1(n271), .A3(n525), .A2(n269), .A4(n325), .S0(n306), 
        .S1(n303), .Y(n524) );
  MUX41X1_HVT U61 ( .A1(n268), .A3(n324), .A2(n323), .A4(n283), .S0(n259), 
        .S1(in[5]), .Y(n522) );
  NAND2X0_HVT U62 ( .A1(n302), .A2(n245), .Y(n521) );
  MUX41X1_HVT U63 ( .A1(n521), .A3(n315), .A2(n255), .A4(n322), .S0(n306), 
        .S1(n303), .Y(n520) );
  AO21X1_HVT U66 ( .A1(n320), .A2(n277), .A3(n344), .Y(n517) );
  MUX41X1_HVT U68 ( .A1(n318), .A3(n517), .A2(n516), .A4(n518), .S0(n272), 
        .S1(n259), .Y(n515) );
  MUX41X1_HVT U69 ( .A1(n515), .A3(n523), .A2(n519), .A4(n529), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n291), .A2(n510), .Y(n511) );
  MUX41X1_HVT U74 ( .A1(n512), .A3(n558), .A2(n511), .A4(n560), .S0(n273), 
        .S1(n259), .Y(n509) );
  MUX41X1_HVT U75 ( .A1(n347), .A3(n352), .A2(n244), .A4(n329), .S0(n272), 
        .S1(n305), .Y(n508) );
  MUX41X1_HVT U82 ( .A1(n539), .A3(n327), .A2(n310), .A4(n569), .S0(n272), 
        .S1(n259), .Y(n500) );
  AND2X1_HVT U83 ( .A1(n299), .A2(n213), .Y(n499) );
  MUX41X1_HVT U84 ( .A1(n328), .A3(n260), .A2(n567), .A4(n499), .S0(n272), 
        .S1(n305), .Y(n498) );
  NAND2X0_HVT U85 ( .A1(n302), .A2(n363), .Y(n497) );
  MUX41X1_HVT U86 ( .A1(n352), .A3(n497), .A2(n266), .A4(n264), .S0(n272), 
        .S1(n304), .Y(n496) );
  MUX41X1_HVT U87 ( .A1(n496), .A3(n500), .A2(n498), .A4(n501), .S0(in[0]), 
        .S1(n275), .Y(n495) );
  MUX41X1_HVT U90 ( .A1(n538), .A3(n542), .A2(n349), .A4(n494), .S0(in[2]), 
        .S1(n305), .Y(n493) );
  AO21X1_HVT U93 ( .A1(n280), .A2(n489), .A3(n348), .Y(n490) );
  MUX41X1_HVT U96 ( .A1(n310), .A3(n267), .A2(n351), .A4(n487), .S0(n272), 
        .S1(n304), .Y(n486) );
  MUX41X1_HVT U97 ( .A1(n347), .A3(n267), .A2(n298), .A4(n568), .S0(n272), 
        .S1(n305), .Y(n485) );
  MUX41X1_HVT U98 ( .A1(n485), .A3(n488), .A2(n486), .A4(n493), .S0(n287), 
        .S1(n275), .Y(n484) );
  NAND2X0_HVT U101 ( .A1(n480), .A2(n479), .Y(n481) );
  MUX41X1_HVT U103 ( .A1(n240), .A3(n319), .A2(n332), .A4(n549), .S0(n272), 
        .S1(n304), .Y(n477) );
  MUX41X1_HVT U105 ( .A1(n331), .A3(n536), .A2(n476), .A4(n346), .S0(n272), 
        .S1(n305), .Y(n475) );
  MUX41X1_HVT U106 ( .A1(n475), .A3(n478), .A2(n477), .A4(n482), .S0(in[0]), 
        .S1(n275), .Y(n474) );
  OA21X1_HVT U109 ( .A1(n338), .A2(n257), .A3(n325), .Y(n472) );
  NAND2X0_HVT U110 ( .A1(n581), .A2(n470), .Y(n471) );
  MUX41X1_HVT U114 ( .A1(n467), .A3(n473), .A2(n469), .A4(n472), .S0(n277), 
        .S1(n304), .Y(n466) );
  NAND2X0_HVT U123 ( .A1(n457), .A2(n456), .Y(n458) );
  MUX41X1_HVT U131 ( .A1(n449), .A3(n451), .A2(n450), .A4(n452), .S0(n277), 
        .S1(n279), .Y(n448) );
  MUX41X1_HVT U132 ( .A1(n448), .A3(n461), .A2(n453), .A4(n466), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  MUX41X1_HVT U135 ( .A1(n356), .A3(n361), .A2(n578), .A4(n557), .S0(n273), 
        .S1(n279), .Y(n445) );
  MUX41X1_HVT U136 ( .A1(n264), .A3(n551), .A2(n357), .A4(n548), .S0(n251), 
        .S1(n279), .Y(n444) );
  AND2X1_HVT U140 ( .A1(n290), .A2(n301), .Y(n440) );
  OA21X1_HVT U144 ( .A1(n313), .A2(n307), .A3(n553), .Y(n436) );
  NAND2X0_HVT U146 ( .A1(n298), .A2(n295), .Y(n510) );
  MUX41X1_HVT U147 ( .A1(n357), .A3(n510), .A2(n347), .A4(n538), .S0(n273), 
        .S1(n280), .Y(n434) );
  MUX41X1_HVT U148 ( .A1(n434), .A3(n438), .A2(n435), .A4(n439), .S0(in[0]), 
        .S1(n275), .Y(n433) );
  OA21X1_HVT U151 ( .A1(n544), .A2(n307), .A3(n430), .Y(n431) );
  MUX41X1_HVT U153 ( .A1(n471), .A3(n268), .A2(n581), .A4(n312), .S0(n274), 
        .S1(n259), .Y(n428) );
  AND2X1_HVT U154 ( .A1(n280), .A2(n289), .Y(n427) );
  NAND2X0_HVT U158 ( .A1(n247), .A2(n363), .Y(n423) );
  MUX41X1_HVT U159 ( .A1(n571), .A3(n283), .A2(n423), .A4(n317), .S0(n238), 
        .S1(n259), .Y(n422) );
  AND2X1_HVT U162 ( .A1(n260), .A2(n510), .Y(n419) );
  NAND2X0_HVT U166 ( .A1(n294), .A2(n527), .Y(n415) );
  NAND2X0_HVT U167 ( .A1(n243), .A2(n302), .Y(n414) );
  MUX41X1_HVT U168 ( .A1(n350), .A3(n290), .A2(n414), .A4(n415), .S0(n238), 
        .S1(n304), .Y(n413) );
  OA21X1_HVT U170 ( .A1(n269), .A2(n307), .A3(n553), .Y(n411) );
  MUX41X1_HVT U172 ( .A1(n410), .A3(n416), .A2(n413), .A4(n418), .S0(in[0]), 
        .S1(n275), .Y(n409) );
  NAND2X0_HVT U174 ( .A1(n297), .A2(n577), .Y(n570) );
  MUX41X1_HVT U176 ( .A1(n284), .A3(n408), .A2(n354), .A4(n570), .S0(n211), 
        .S1(n238), .Y(n407) );
  NAND2X0_HVT U177 ( .A1(n300), .A2(n285), .Y(n406) );
  MUX41X1_HVT U178 ( .A1(n566), .A3(n406), .A2(n358), .A4(n546), .S0(n273), 
        .S1(n259), .Y(n405) );
  MUX41X1_HVT U179 ( .A1(n556), .A3(n359), .A2(n314), .A4(n358), .S0(n238), 
        .S1(n305), .Y(n404) );
  MUX41X1_HVT U180 ( .A1(n316), .A3(n575), .A2(n571), .A4(n263), .S0(n278), 
        .S1(n238), .Y(n403) );
  MUX41X1_HVT U181 ( .A1(n403), .A3(n405), .A2(n404), .A4(n407), .S0(n287), 
        .S1(n276), .Y(n402) );
  MUX41X1_HVT U182 ( .A1(n340), .A3(n579), .A2(n342), .A4(n330), .S0(n211), 
        .S1(n253), .Y(n401) );
  OA21X1_HVT U184 ( .A1(n550), .A2(n307), .A3(n328), .Y(n399) );
  MUX41X1_HVT U186 ( .A1(n267), .A3(n545), .A2(n510), .A4(n538), .S0(n238), 
        .S1(n259), .Y(n397) );
  MUX41X1_HVT U189 ( .A1(n395), .A3(n570), .A2(n396), .A4(n346), .S0(n278), 
        .S1(n238), .Y(n394) );
  MUX41X1_HVT U190 ( .A1(n394), .A3(n397), .A2(n398), .A4(n401), .S0(n276), 
        .S1(n287), .Y(n393) );
  MUX41X1_HVT U195 ( .A1(n260), .A3(n351), .A2(n582), .A4(n547), .S0(n238), 
        .S1(n304), .Y(n389) );
  AO21X1_HVT U197 ( .A1(n266), .A2(n279), .A3(n348), .Y(n387) );
  OA21X1_HVT U201 ( .A1(n576), .A2(n307), .A3(n339), .Y(n383) );
  MUX41X1_HVT U203 ( .A1(n548), .A3(n341), .A2(n572), .A4(n552), .S0(n238), 
        .S1(n305), .Y(n381) );
  MUX41X1_HVT U204 ( .A1(n528), .A3(n571), .A2(n218), .A4(n561), .S0(n253), 
        .S1(n304), .Y(n380) );
  MUX41X1_HVT U205 ( .A1(n213), .A3(n239), .A2(n359), .A4(n335), .S0(n238), 
        .S1(n259), .Y(n379) );
  NAND2X0_HVT U208 ( .A1(n296), .A2(n293), .Y(n470) );
  NAND2X0_HVT U212 ( .A1(n298), .A2(n291), .Y(n527) );
  NAND2X0_HVT U214 ( .A1(n260), .A2(n302), .Y(n377) );
  NAND2X0_HVT U215 ( .A1(n470), .A2(n292), .Y(n376) );
  AO21X1_HVT U216 ( .A1(n301), .A2(n361), .A3(n307), .Y(n480) );
  NAND2X0_HVT U218 ( .A1(n361), .A2(n299), .Y(n430) );
  NAND2X0_HVT U220 ( .A1(n279), .A2(n377), .Y(n502) );
  NAND2X0_HVT U1 ( .A1(n312), .A2(n3), .Y(n23) );
  NAND2X0_HVT U2 ( .A1(n218), .A2(n274), .Y(n50) );
  NAND2X0_HVT U3 ( .A1(n23), .A2(n50), .Y(n464) );
  IBUFFX2_HVT U6 ( .A(n274), .Y(n3) );
  MUX21X1_HVT U7 ( .A1(n288), .A2(n295), .S0(n224), .Y(n218) );
  MUX21X1_HVT U8 ( .A1(n463), .A2(n464), .S0(n279), .Y(n462) );
  INVX2_HVT U9 ( .A(in[7]), .Y(n308) );
  MUX41X1_HVT U10 ( .A1(n429), .A3(n424), .A2(n428), .A4(n422), .S0(n121), 
        .S1(n219), .Y(n421) );
  IBUFFX16_HVT U11 ( .A(n287), .Y(n121) );
  IBUFFX2_HVT U12 ( .A(n307), .Y(n305) );
  IBUFFX2_HVT U14 ( .A(n218), .Y(n550) );
  MUX21X2_HVT U16 ( .A1(n443), .A2(n580), .S0(n251), .Y(n442) );
  IBUFFX2_HVT U17 ( .A(n301), .Y(n297) );
  MUX21X2_HVT U18 ( .A1(n505), .A2(n495), .S0(n210), .Y(out[1]) );
  IBUFFX16_HVT U19 ( .A(in[6]), .Y(n210) );
  INVX1_HVT U20 ( .A(n301), .Y(n298) );
  INVX1_HVT U22 ( .A(n300), .Y(n224) );
  IBUFFX2_HVT U23 ( .A(n301), .Y(n300) );
  INVX2_HVT U25 ( .A(in[1]), .Y(n301) );
  INVX0_HVT U26 ( .A(in[1]), .Y(n302) );
  INVX0_HVT U27 ( .A(n301), .Y(n299) );
  INVX0_HVT U28 ( .A(n301), .Y(n296) );
  INVX0_HVT U29 ( .A(n301), .Y(n247) );
  INVX0_HVT U30 ( .A(n235), .Y(n211) );
  MUX21X1_HVT U31 ( .A1(n561), .A2(n340), .S0(n279), .Y(n443) );
  IBUFFX4_HVT U32 ( .A(n307), .Y(n259) );
  INVX2_HVT U34 ( .A(n308), .Y(n306) );
  INVX1_HVT U36 ( .A(n250), .Y(n579) );
  NBUFFX2_HVT U37 ( .A(n365), .Y(n285) );
  MUX21X1_HVT U38 ( .A1(n289), .A2(n282), .S0(n302), .Y(n561) );
  MUX21X1_HVT U39 ( .A1(n212), .A2(n555), .S0(n235), .Y(n437) );
  MUX21X1_HVT U40 ( .A1(n285), .A2(n281), .S0(n247), .Y(n460) );
  INVX0_HVT U41 ( .A(n212), .Y(n239) );
  MUX21X1_HVT U43 ( .A1(n286), .A2(n360), .S0(n299), .Y(n555) );
  XOR2X1_HVT U44 ( .A1(n307), .A2(n557), .Y(n540) );
  INVX1_HVT U45 ( .A(n231), .Y(n507) );
  INVX0_HVT U46 ( .A(n286), .Y(n232) );
  INVX2_HVT U47 ( .A(n236), .Y(n238) );
  MUX21X1_HVT U48 ( .A1(n363), .A2(n283), .S0(n300), .Y(n420) );
  INVX0_HVT U49 ( .A(n581), .Y(n244) );
  INVX0_HVT U50 ( .A(n261), .Y(n242) );
  AND2X1_HVT U52 ( .A1(n299), .A2(n245), .Y(n212) );
  NBUFFX2_HVT U54 ( .A(n364), .Y(n282) );
  INVX1_HVT U55 ( .A(n278), .Y(n235) );
  INVX1_HVT U60 ( .A(n244), .Y(n246) );
  INVX1_HVT U64 ( .A(in[0]), .Y(n241) );
  INVX0_HVT U65 ( .A(n277), .Y(n219) );
  INVX1_HVT U67 ( .A(in[3]), .Y(n362) );
  MUX21X1_HVT U70 ( .A1(n393), .A2(n402), .S0(in[6]), .Y(out[6]) );
  NBUFFX2_HVT U71 ( .A(in[2]), .Y(n274) );
  INVX1_HVT U72 ( .A(n257), .Y(n251) );
  NBUFFX2_HVT U76 ( .A(in[2]), .Y(n272) );
  DELLN1X2_HVT U77 ( .A(in[2]), .Y(n273) );
  MUX21X1_HVT U78 ( .A1(n334), .A2(n447), .S0(n272), .Y(n446) );
  MUX21X1_HVT U79 ( .A1(n388), .A2(n387), .S0(n274), .Y(n386) );
  MUX21X1_HVT U80 ( .A1(n540), .A2(n514), .S0(n274), .Y(n513) );
  MUX21X1_HVT U81 ( .A1(n504), .A2(n503), .S0(n253), .Y(n501) );
  MUX21X1_HVT U88 ( .A1(n311), .A2(n460), .S0(n273), .Y(n459) );
  INVX1_HVT U89 ( .A(n253), .Y(n236) );
  INVX1_HVT U91 ( .A(n285), .Y(n213) );
  IBUFFX2_HVT U92 ( .A(n575), .Y(n319) );
  NAND2X0_HVT U94 ( .A1(n426), .A2(n251), .Y(n216) );
  NAND2X0_HVT U95 ( .A1(n425), .A2(n252), .Y(n217) );
  NAND2X0_HVT U99 ( .A1(n216), .A2(n217), .Y(n424) );
  MUX21X1_HVT U100 ( .A1(n360), .A2(n363), .S0(n224), .Y(n546) );
  MUX21X1_HVT U102 ( .A1(n353), .A2(n546), .S0(n235), .Y(n425) );
  NBUFFX4_HVT U104 ( .A(n579), .Y(n293) );
  MUX41X1_HVT U107 ( .A1(n444), .A3(n446), .A2(n442), .A4(n445), .S0(n287), 
        .S1(n219), .Y(n441) );
  AND3X1_HVT U108 ( .A1(n246), .A2(n527), .A3(n502), .Y(n503) );
  MUX21X2_HVT U111 ( .A1(n459), .A2(n458), .S0(n280), .Y(n455) );
  INVX1_HVT U112 ( .A(n579), .Y(n360) );
  MUX21X2_HVT U113 ( .A1(n454), .A2(n455), .S0(n277), .Y(n453) );
  INVX0_HVT U115 ( .A(n555), .Y(n332) );
  INVX1_HVT U116 ( .A(n577), .Y(n364) );
  INVX1_HVT U117 ( .A(n371), .Y(n334) );
  INVX0_HVT U118 ( .A(n547), .Y(n338) );
  INVX0_HVT U119 ( .A(n561), .Y(n328) );
  MUX21X2_HVT U120 ( .A1(n465), .A2(n462), .S0(n219), .Y(n461) );
  INVX1_HVT U121 ( .A(n582), .Y(n363) );
  MUX41X1_HVT U122 ( .A1(n345), .A3(n290), .A2(n328), .A4(n283), .S0(in[2]), 
        .S1(n308), .Y(n438) );
  INVX0_HVT U124 ( .A(n546), .Y(n339) );
  MUX21X1_HVT U125 ( .A1(n293), .A2(n577), .S0(n247), .Y(n547) );
  MUX21X2_HVT U126 ( .A1(n436), .A2(n437), .S0(n252), .Y(n435) );
  MUX21X2_HVT U127 ( .A1(n292), .A2(n355), .S0(n235), .Y(n447) );
  MUX21X1_HVT U128 ( .A1(n285), .A2(n360), .S0(n224), .Y(n370) );
  MUX21X1_HVT U129 ( .A1(n232), .A2(n364), .S0(n224), .Y(n231) );
  INVX1_HVT U130 ( .A(n364), .Y(n260) );
  INVX1_HVT U133 ( .A(n576), .Y(n318) );
  INVX1_HVT U134 ( .A(n370), .Y(n355) );
  MUX21X1_HVT U137 ( .A1(n363), .A2(n282), .S0(n224), .Y(n576) );
  NAND2X0_HVT U138 ( .A1(n378), .A2(n261), .Y(n233) );
  NAND2X0_HVT U139 ( .A1(n385), .A2(n242), .Y(n234) );
  NAND2X0_HVT U141 ( .A1(n233), .A2(n234), .Y(out[7]) );
  MUX21X2_HVT U142 ( .A1(n384), .A2(n383), .S0(n252), .Y(n382) );
  AO21X1_HVT U143 ( .A1(n272), .A2(n290), .A3(n260), .Y(n463) );
  MUX41X1_HVT U145 ( .A1(n419), .A3(n324), .A2(n420), .A4(n265), .S0(n236), 
        .S1(n305), .Y(n418) );
  MUX21X1_HVT U149 ( .A1(n282), .A2(n289), .S0(n302), .Y(n237) );
  MUX21X1_HVT U150 ( .A1(n361), .A2(n237), .S0(n235), .Y(n432) );
  NBUFFX4_HVT U152 ( .A(n365), .Y(n284) );
  IBUFFX2_HVT U155 ( .A(n544), .Y(n341) );
  NBUFFX2_HVT U156 ( .A(in[2]), .Y(n253) );
  MUX41X1_HVT U157 ( .A1(n379), .A3(n380), .A2(n381), .A4(n382), .S0(n276), 
        .S1(n287), .Y(n378) );
  IBUFFX2_HVT U160 ( .A(n527), .Y(n347) );
  INVX0_HVT U161 ( .A(n253), .Y(n252) );
  MUX41X1_HVT U163 ( .A1(n513), .A3(n508), .A2(n509), .A4(n506), .S0(n241), 
        .S1(n219), .Y(n505) );
  INVX1_HVT U164 ( .A(n212), .Y(n240) );
  MUX21X2_HVT U165 ( .A1(n432), .A2(n431), .S0(n252), .Y(n429) );
  MUX41X1_HVT U169 ( .A1(n391), .A3(n389), .A2(n390), .A4(n386), .S0(n241), 
        .S1(n219), .Y(n385) );
  MUX41X1_HVT U171 ( .A1(n355), .A3(n318), .A2(n271), .A4(n562), .S0(n252), 
        .S1(n308), .Y(n454) );
  INVX1_HVT U173 ( .A(n581), .Y(n243) );
  INVX1_HVT U175 ( .A(n244), .Y(n245) );
  NAND2X0_HVT U183 ( .A1(n281), .A2(n297), .Y(n248) );
  NAND2X0_HVT U185 ( .A1(n282), .A2(n301), .Y(n249) );
  NAND2X0_HVT U187 ( .A1(n248), .A2(n249), .Y(n567) );
  INVX0_HVT U188 ( .A(n567), .Y(n323) );
  MUX21X1_HVT U191 ( .A1(n567), .A2(n263), .S0(n278), .Y(n384) );
  AND2X1_HVT U192 ( .A1(n284), .A2(n362), .Y(n250) );
  INVX1_HVT U193 ( .A(n367), .Y(n358) );
  MUX41X1_HVT U194 ( .A1(n557), .A3(n543), .A2(n290), .A4(n356), .S0(n235), 
        .S1(n251), .Y(n390) );
  IBUFFX2_HVT U196 ( .A(n543), .Y(n342) );
  MUX41X1_HVT U198 ( .A1(n549), .A3(n542), .A2(n392), .A4(n535), .S0(n252), 
        .S1(n304), .Y(n391) );
  MUX21X2_HVT U199 ( .A1(n409), .A2(n421), .S0(in[6]), .Y(out[5]) );
  INVX0_HVT U200 ( .A(n307), .Y(n304) );
  INVX0_HVT U202 ( .A(n329), .Y(n256) );
  MUX21X1_HVT U206 ( .A1(n335), .A2(n569), .S0(n251), .Y(n483) );
  INVX0_HVT U207 ( .A(in[6]), .Y(n261) );
  INVX1_HVT U209 ( .A(in[2]), .Y(n257) );
  INVX1_HVT U210 ( .A(n553), .Y(n335) );
  INVX0_HVT U211 ( .A(n571), .Y(n255) );
  INVX1_HVT U213 ( .A(n254), .Y(n465) );
  MUX41X1_HVT U217 ( .A1(n335), .A3(n256), .A2(n258), .A4(n255), .S0(n257), 
        .S1(n308), .Y(n254) );
  NAND2X0_HVT U219 ( .A1(n247), .A2(n282), .Y(n258) );
  AND3X2_HVT U221 ( .A1(n272), .A2(n302), .A3(n213), .Y(n451) );
  MUX41X1_HVT U222 ( .A1(n237), .A3(n507), .A2(n353), .A4(n575), .S0(n235), 
        .S1(n257), .Y(n506) );
  INVX2_HVT U223 ( .A(in[7]), .Y(n307) );
  XOR2X2_HVT U224 ( .A1(n284), .A2(n288), .Y(n577) );
  MUX41X1_HVT U225 ( .A1(n336), .A3(n440), .A2(n339), .A4(n559), .S0(n257), 
        .S1(n308), .Y(n439) );
  MUX21X2_HVT U226 ( .A1(n433), .A2(n441), .S0(in[6]), .Y(out[4]) );
  MUX41X1_HVT U227 ( .A1(n417), .A3(n538), .A2(n333), .A4(n562), .S0(n308), 
        .S1(n257), .Y(n416) );
  XOR2X1_HVT U228 ( .A1(n257), .A2(n308), .Y(n537) );
  MUX21X1_HVT U229 ( .A1(n245), .A2(n468), .S0(n262), .Y(n467) );
  XNOR2X1_HVT U230 ( .A1(n302), .A2(n257), .Y(n262) );
  MUX21X2_HVT U231 ( .A1(n268), .A2(n483), .S0(n537), .Y(n482) );
  MUX21X1_HVT U232 ( .A1(n265), .A2(n323), .S0(n274), .Y(n450) );
  NBUFFX2_HVT U233 ( .A(n364), .Y(n283) );
  AND2X1_HVT U234 ( .A1(n283), .A2(n527), .Y(n263) );
  MUX21X1_HVT U235 ( .A1(n360), .A2(n363), .S0(n277), .Y(n531) );
  MUX21X1_HVT U236 ( .A1(n553), .A2(n471), .S0(n274), .Y(n469) );
  MUX21X1_HVT U237 ( .A1(n319), .A2(n361), .S0(n277), .Y(n516) );
  AND2X1_HVT U238 ( .A1(n246), .A2(n510), .Y(n264) );
  MUX21X1_HVT U239 ( .A1(n246), .A2(n283), .S0(n298), .Y(n543) );
  MUX21X1_HVT U240 ( .A1(n283), .A2(n286), .S0(n297), .Y(n479) );
  MUX21X1_HVT U241 ( .A1(n360), .A2(n243), .S0(n300), .Y(n408) );
  MUX21X1_HVT U242 ( .A1(n283), .A2(n360), .S0(n298), .Y(n487) );
  MUX21X1_HVT U243 ( .A1(n260), .A2(n361), .S0(n299), .Y(n369) );
  MUX21X1_HVT U244 ( .A1(n577), .A2(n243), .S0(n297), .Y(n559) );
  XOR2X1_HVT U245 ( .A1(n577), .A2(n296), .Y(n538) );
  MUX21X1_HVT U246 ( .A1(n243), .A2(n363), .S0(n297), .Y(n557) );
  MUX21X1_HVT U247 ( .A1(n281), .A2(n243), .S0(n247), .Y(n544) );
  MUX21X1_HVT U248 ( .A1(n293), .A2(n292), .S0(n247), .Y(n494) );
  XOR2X1_HVT U249 ( .A1(n299), .A2(n361), .Y(n539) );
  MUX21X1_HVT U250 ( .A1(n362), .A2(n295), .S0(n296), .Y(n395) );
  MUX21X1_HVT U251 ( .A1(n295), .A2(n581), .S0(n300), .Y(n396) );
  MUX21X1_HVT U252 ( .A1(n361), .A2(n360), .S0(n298), .Y(n565) );
  INVX1_HVT U253 ( .A(n290), .Y(n361) );
  MUX21X1_HVT U254 ( .A1(n246), .A2(n291), .S0(n298), .Y(n569) );
  MUX21X1_HVT U255 ( .A1(n293), .A2(n295), .S0(n247), .Y(n489) );
  MUX21X1_HVT U256 ( .A1(n281), .A2(n363), .S0(n296), .Y(n573) );
  MUX21X1_HVT U257 ( .A1(n293), .A2(n281), .S0(n300), .Y(n572) );
  MUX21X1_HVT U258 ( .A1(n362), .A2(n286), .S0(n300), .Y(n392) );
  XOR2X1_HVT U259 ( .A1(n246), .A2(n296), .Y(n535) );
  XNOR2X1_HVT U260 ( .A1(n579), .A2(n297), .Y(n265) );
  MUX21X1_HVT U261 ( .A1(n294), .A2(n291), .S0(n298), .Y(n553) );
  MUX21X1_HVT U262 ( .A1(n246), .A2(n285), .S0(n299), .Y(n375) );
  MUX21X1_HVT U263 ( .A1(n245), .A2(n293), .S0(n300), .Y(n368) );
  XNOR2X1_HVT U264 ( .A1(n294), .A2(n299), .Y(n266) );
  AND2X1_HVT U265 ( .A1(n296), .A2(n243), .Y(n267) );
  MUX21X1_HVT U266 ( .A1(n291), .A2(n281), .S0(n247), .Y(n373) );
  AND2X1_HVT U267 ( .A1(n294), .A2(n470), .Y(n268) );
  MUX21X1_HVT U268 ( .A1(n292), .A2(n285), .S0(n296), .Y(n512) );
  MUX21X1_HVT U269 ( .A1(n292), .A2(n295), .S0(n274), .Y(n457) );
  XOR2X1_HVT U270 ( .A1(n284), .A2(n299), .Y(n558) );
  NBUFFX2_HVT U271 ( .A(n306), .Y(n280) );
  NBUFFX2_HVT U272 ( .A(n306), .Y(n278) );
  NBUFFX2_HVT U273 ( .A(n306), .Y(n279) );
  NBUFFX2_HVT U274 ( .A(n362), .Y(n281) );
  NBUFFX2_HVT U275 ( .A(in[5]), .Y(n277) );
  NBUFFX2_HVT U276 ( .A(n303), .Y(n276) );
  NBUFFX2_HVT U277 ( .A(n303), .Y(n275) );
  MUX21X1_HVT U278 ( .A1(n481), .A2(n334), .S0(n251), .Y(n478) );
  MUX21X1_HVT U279 ( .A1(n399), .A2(n400), .S0(n274), .Y(n398) );
  MUX21X1_HVT U280 ( .A1(n497), .A2(n288), .S0(n279), .Y(n400) );
  MUX21X1_HVT U281 ( .A1(n520), .A2(n522), .S0(n274), .Y(n519) );
  XOR2X1_HVT U282 ( .A1(n297), .A2(n289), .Y(n536) );
  MUX21X1_HVT U283 ( .A1(n291), .A2(n364), .S0(n300), .Y(n476) );
  MUX21X1_HVT U284 ( .A1(n563), .A2(n292), .S0(n280), .Y(n504) );
  MUX21X1_HVT U285 ( .A1(n412), .A2(n411), .S0(n253), .Y(n410) );
  MUX21X1_HVT U286 ( .A1(n292), .A2(n351), .S0(n280), .Y(n412) );
  AND2X1_HVT U287 ( .A1(n364), .A2(n302), .Y(n269) );
  MUX21X1_HVT U288 ( .A1(n288), .A2(n360), .S0(n298), .Y(n545) );
  MUX21X1_HVT U289 ( .A1(n363), .A2(n351), .S0(n280), .Y(n514) );
  MUX21X1_HVT U290 ( .A1(n566), .A2(n336), .S0(n273), .Y(n449) );
  MUX21X1_HVT U291 ( .A1(n361), .A2(n243), .S0(n297), .Y(n417) );
  NAND2X0_HVT U292 ( .A1(n289), .A2(n286), .Y(n581) );
  NBUFFX2_HVT U293 ( .A(n365), .Y(n286) );
  MUX21X1_HVT U294 ( .A1(n243), .A2(n288), .S0(n300), .Y(n564) );
  MUX21X1_HVT U295 ( .A1(n337), .A2(n239), .S0(n273), .Y(n473) );
  MUX21X1_HVT U296 ( .A1(n427), .A2(n246), .S0(n270), .Y(n426) );
  MUX21X1_HVT U297 ( .A1(n240), .A2(n301), .S0(n274), .Y(n456) );
  NBUFFX2_HVT U298 ( .A(n574), .Y(n290) );
  MUX21X1_HVT U299 ( .A1(n532), .A2(n533), .S0(n278), .Y(n530) );
  MUX21X1_HVT U300 ( .A1(n289), .A2(n549), .S0(n277), .Y(n533) );
  XOR2X1_HVT U301 ( .A1(n296), .A2(n276), .Y(n541) );
  NBUFFX2_HVT U302 ( .A(n574), .Y(n291) );
  MUX21X1_HVT U303 ( .A1(n288), .A2(n361), .S0(n298), .Y(n372) );
  MUX21X1_HVT U304 ( .A1(n343), .A2(n358), .S0(n306), .Y(n388) );
  MUX21X1_HVT U305 ( .A1(n554), .A2(n376), .S0(n278), .Y(n371) );
  MUX21X1_HVT U306 ( .A1(n293), .A2(n289), .S0(n296), .Y(n575) );
  MUX21X1_HVT U307 ( .A1(n331), .A2(n554), .S0(n273), .Y(n452) );
  MUX21X1_HVT U308 ( .A1(n321), .A2(n302), .S0(n277), .Y(n518) );
  MUX21X1_HVT U309 ( .A1(n245), .A2(n492), .S0(n270), .Y(n491) );
  MUX21X1_HVT U310 ( .A1(n288), .A2(n285), .S0(n280), .Y(n492) );
  NBUFFX2_HVT U311 ( .A(n582), .Y(n295) );
  NBUFFX2_HVT U312 ( .A(n574), .Y(n292) );
  NBUFFX2_HVT U313 ( .A(n582), .Y(n294) );
  XNOR2X1_HVT U314 ( .A1(n307), .A2(n297), .Y(n270) );
  AND2X1_HVT U315 ( .A1(n281), .A2(n302), .Y(n271) );
  NBUFFX2_HVT U316 ( .A(in[5]), .Y(n303) );
  INVX0_HVT U317 ( .A(in[4]), .Y(n365) );
  MUX21X1_HVT U318 ( .A1(n474), .A2(n484), .S0(in[6]), .Y(out[2]) );
  MUX21X1_HVT U319 ( .A1(n490), .A2(n491), .S0(n274), .Y(n488) );
  MUX21X1_HVT U320 ( .A1(n530), .A2(n534), .S0(n251), .Y(n529) );
  MUX21X1_HVT U321 ( .A1(n524), .A2(n526), .S0(n274), .Y(n523) );
  MUX21X1_HVT U322 ( .A1(n360), .A2(n213), .S0(n298), .Y(n552) );
  NAND2X0_HVT U323 ( .A1(in[3]), .A2(in[4]), .Y(n582) );
  MUX21X1_HVT U324 ( .A1(n213), .A2(n260), .S0(n297), .Y(n374) );
  MUX21X1_HVT U325 ( .A1(n213), .A2(n363), .S0(n299), .Y(n548) );
  MUX21X1_HVT U326 ( .A1(n213), .A2(n361), .S0(n247), .Y(n566) );
  NAND2X0_HVT U327 ( .A1(in[4]), .A2(n362), .Y(n574) );
  MUX21X1_HVT U328 ( .A1(n213), .A2(n245), .S0(n296), .Y(n563) );
  MUX21X1_HVT U329 ( .A1(n213), .A2(n291), .S0(n297), .Y(n367) );
  MUX21X1_HVT U330 ( .A1(n295), .A2(n213), .S0(n247), .Y(n556) );
  MUX21X1_HVT U331 ( .A1(n289), .A2(n213), .S0(in[2]), .Y(n468) );
  MUX21X1_HVT U332 ( .A1(n213), .A2(n294), .S0(n247), .Y(n366) );
  MUX21X1_HVT U333 ( .A1(n281), .A2(n213), .S0(n299), .Y(n554) );
  NBUFFX2_HVT U334 ( .A(in[3]), .Y(n288) );
  NBUFFX2_HVT U335 ( .A(in[3]), .Y(n289) );
  NBUFFX2_HVT U336 ( .A(in[0]), .Y(n287) );
  INVX0_HVT U337 ( .A(n562), .Y(n309) );
  INVX0_HVT U338 ( .A(n560), .Y(n310) );
  INVX0_HVT U339 ( .A(n551), .Y(n311) );
  INVX0_HVT U340 ( .A(n549), .Y(n312) );
  INVX0_HVT U341 ( .A(n414), .Y(n313) );
  INVX0_HVT U342 ( .A(n377), .Y(n314) );
  INVX0_HVT U343 ( .A(n568), .Y(n315) );
  INVX0_HVT U344 ( .A(n580), .Y(n316) );
  INVX0_HVT U345 ( .A(n578), .Y(n317) );
  INVX0_HVT U346 ( .A(n573), .Y(n320) );
  INVX0_HVT U347 ( .A(n572), .Y(n321) );
  INVX0_HVT U348 ( .A(n569), .Y(n322) );
  INVX0_HVT U349 ( .A(n566), .Y(n324) );
  INVX0_HVT U350 ( .A(n565), .Y(n325) );
  INVX0_HVT U351 ( .A(n564), .Y(n326) );
  INVX0_HVT U352 ( .A(n563), .Y(n327) );
  INVX0_HVT U353 ( .A(n559), .Y(n329) );
  INVX0_HVT U354 ( .A(n558), .Y(n330) );
  INVX0_HVT U355 ( .A(n556), .Y(n331) );
  INVX0_HVT U356 ( .A(n554), .Y(n333) );
  INVX0_HVT U357 ( .A(n552), .Y(n336) );
  INVX0_HVT U358 ( .A(n548), .Y(n337) );
  INVX0_HVT U359 ( .A(n545), .Y(n340) );
  INVX0_HVT U360 ( .A(n542), .Y(n343) );
  INVX0_HVT U361 ( .A(n510), .Y(n344) );
  INVX0_HVT U362 ( .A(n470), .Y(n345) );
  INVX0_HVT U363 ( .A(n376), .Y(n346) );
  INVX0_HVT U364 ( .A(n430), .Y(n348) );
  INVX0_HVT U365 ( .A(n375), .Y(n349) );
  INVX0_HVT U366 ( .A(n374), .Y(n350) );
  INVX0_HVT U367 ( .A(n373), .Y(n351) );
  INVX0_HVT U368 ( .A(n372), .Y(n352) );
  INVX0_HVT U369 ( .A(n489), .Y(n353) );
  INVX0_HVT U370 ( .A(n479), .Y(n354) );
  INVX0_HVT U371 ( .A(n369), .Y(n356) );
  INVX0_HVT U372 ( .A(n368), .Y(n357) );
  INVX0_HVT U373 ( .A(n366), .Y(n359) );
endmodule

