
module sbox_4 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n5, n19, n23, n33, n50, n118, n119, n210, n211, n212, n213, n216,
         n217, n218, n219, n222, n224, n227, n231, n232, n234, n236, n238,
         n245, n249, n252, n261, n264, n271, n273, n274, n275, n278, n279,
         n280, n282, n283, n285, n289, n291, n293, n296, n297, n300, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768;

  NAND2X0_HVT U4 ( .A1(n411), .A2(n766), .Y(n765) );
  NAND2X0_HVT U5 ( .A1(n231), .A2(n489), .Y(n764) );
  NAND2X0_HVT U15 ( .A1(n766), .A2(n484), .Y(n754) );
  NAND2X0_HVT U21 ( .A1(n357), .A2(n502), .Y(n749) );
  NAND2X0_HVT U24 ( .A1(n395), .A2(n502), .Y(n747) );
  NAND2X0_HVT U33 ( .A1(n410), .A2(n502), .Y(n739) );
  NAND2X0_HVT U42 ( .A1(n401), .A2(n483), .Y(n730) );
  MUX41X1_HVT U51 ( .A1(n516), .A3(n535), .A2(n512), .A4(n436), .S0(n300), 
        .S1(n477), .Y(n722) );
  NAND2X0_HVT U53 ( .A1(n719), .A2(n729), .Y(n720) );
  NAND2X0_HVT U56 ( .A1(n411), .A2(n715), .Y(n716) );
  NAND2X0_HVT U58 ( .A1(n498), .A2(n766), .Y(n713) );
  NAND2X0_HVT U62 ( .A1(n119), .A2(n496), .Y(n709) );
  MUX41X1_HVT U63 ( .A1(n709), .A3(n519), .A2(n449), .A4(n518), .S0(n462), 
        .S1(n477), .Y(n708) );
  NAND2X0_HVT U73 ( .A1(n491), .A2(n698), .Y(n699) );
  AND3X1_HVT U80 ( .A1(n494), .A2(n715), .A3(n690), .Y(n691) );
  AND2X1_HVT U83 ( .A1(n401), .A2(n458), .Y(n687) );
  MUX41X1_HVT U86 ( .A1(n546), .A3(n685), .A2(n469), .A4(n465), .S0(n429), 
        .S1(n508), .Y(n684) );
  MUX41X1_HVT U90 ( .A1(n249), .A3(n730), .A2(n516), .A4(n682), .S0(n347), 
        .S1(n508), .Y(n681) );
  NAND2X0_HVT U101 ( .A1(n668), .A2(n667), .Y(n669) );
  MUX41X1_HVT U103 ( .A1(n766), .A3(n537), .A2(n526), .A4(n737), .S0(n421), 
        .S1(n507), .Y(n665) );
  NAND2X0_HVT U110 ( .A1(n494), .A2(n658), .Y(n659) );
  AND2X1_HVT U115 ( .A1(n453), .A2(n484), .Y(n655) );
  NAND2X0_HVT U123 ( .A1(n646), .A2(n645), .Y(n647) );
  MUX41X1_HVT U125 ( .A1(n749), .A3(n472), .A2(n521), .A4(n530), .S0(n421), 
        .S1(n479), .Y(n643) );
  MUX41X1_HVT U135 ( .A1(n19), .A3(n444), .A2(n764), .A4(n744), .S0(n421), 
        .S1(n422), .Y(n634) );
  AND2X1_HVT U140 ( .A1(n326), .A2(n238), .Y(n629) );
  AND2X1_HVT U154 ( .A1(n461), .A2(n483), .Y(n616) );
  NAND2X0_HVT U158 ( .A1(n231), .A2(n418), .Y(n612) );
  MUX41X1_HVT U159 ( .A1(n757), .A3(n484), .A2(n612), .A4(n554), .S0(n429), 
        .S1(n509), .Y(n611) );
  AND2X1_HVT U162 ( .A1(n381), .A2(n285), .Y(n608) );
  MUX41X1_HVT U165 ( .A1(n749), .A3(n543), .A2(n249), .A4(n606), .S0(n479), 
        .S1(n429), .Y(n605) );
  NAND2X0_HVT U166 ( .A1(n498), .A2(n715), .Y(n604) );
  NAND2X0_HVT U167 ( .A1(n437), .A2(n336), .Y(n603) );
  MUX41X1_HVT U168 ( .A1(n524), .A3(n492), .A2(n603), .A4(n604), .S0(n441), 
        .S1(n509), .Y(n602) );
  NAND2X0_HVT U174 ( .A1(n324), .A2(n311), .Y(n756) );
  NAND2X0_HVT U177 ( .A1(n231), .A2(n487), .Y(n595) );
  MUX41X1_HVT U179 ( .A1(n743), .A3(n541), .A2(n525), .A4(n542), .S0(n441), 
        .S1(n508), .Y(n593) );
  MUX41X1_HVT U182 ( .A1(n529), .A3(n391), .A2(n517), .A4(n538), .S0(n461), 
        .S1(n264), .Y(n590) );
  MUX41X1_HVT U189 ( .A1(n584), .A3(n756), .A2(n585), .A4(n534), .S0(n462), 
        .S1(n441), .Y(n583) );
  AO21X1_HVT U197 ( .A1(n469), .A2(n461), .A3(n545), .Y(n576) );
  NAND2X0_HVT U208 ( .A1(n501), .A2(n357), .Y(n658) );
  NAND2X0_HVT U212 ( .A1(n365), .A2(n493), .Y(n715) );
  NAND2X0_HVT U214 ( .A1(n311), .A2(n502), .Y(n566) );
  NAND2X0_HVT U215 ( .A1(n658), .A2(n325), .Y(n565) );
  NAND2X0_HVT U218 ( .A1(n547), .A2(n231), .Y(n619) );
  NAND2X0_HVT U220 ( .A1(n566), .A2(n463), .Y(n690) );
  INVX0_HVT U241 ( .A(n747), .Y(n556) );
  INVX0_HVT U245 ( .A(n764), .Y(n554) );
  INVX0_HVT U256 ( .A(n619), .Y(n545) );
  INVX0_HVT U262 ( .A(n557), .Y(n541) );
  INVX0_HVT U264 ( .A(n737), .Y(n539) );
  INVX0_HVT U265 ( .A(n745), .Y(n538) );
  INVX0_HVT U268 ( .A(n749), .Y(n535) );
  INVX0_HVT U270 ( .A(n565), .Y(n534) );
  INVX0_HVT U276 ( .A(n733), .Y(n529) );
  INVX0_HVT U277 ( .A(n734), .Y(n528) );
  INVX0_HVT U278 ( .A(n739), .Y(n527) );
  INVX0_HVT U284 ( .A(n566), .Y(n525) );
  INVX0_HVT U294 ( .A(n762), .Y(n521) );
  INVX0_HVT U295 ( .A(n765), .Y(n520) );
  INVX0_HVT U302 ( .A(n564), .Y(n516) );
  INVX0_HVT U306 ( .A(n603), .Y(n514) );
  XOR2X1_HVT U1 ( .A1(n314), .A2(n387), .Y(n446) );
  INVX1_HVT U2 ( .A(n234), .Y(n236) );
  MUX21X1_HVT U3 ( .A1(n410), .A2(n314), .S0(n336), .Y(n675) );
  MUX21X1_HVT U6 ( .A1(n278), .A2(n495), .S0(n335), .Y(n426) );
  INVX1_HVT U7 ( .A(n491), .Y(n444) );
  NBUFFX2_HVT U8 ( .A(n236), .Y(n492) );
  INVX1_HVT U9 ( .A(n303), .Y(n508) );
  MUX21X1_HVT U10 ( .A1(n753), .A2(n464), .S0(n461), .Y(n573) );
  MUX21X1_HVT U11 ( .A1(n490), .A2(n406), .S0(n227), .Y(n758) );
  INVX1_HVT U12 ( .A(n303), .Y(n509) );
  NBUFFX2_HVT U13 ( .A(n503), .Y(n421) );
  INVX1_HVT U14 ( .A(n118), .Y(n577) );
  INVX1_HVT U16 ( .A(n510), .Y(n507) );
  INVX1_HVT U17 ( .A(n507), .Y(n404) );
  INVX0_HVT U18 ( .A(n741), .Y(n543) );
  INVX1_HVT U19 ( .A(n333), .Y(n502) );
  INVX1_HVT U20 ( .A(n378), .Y(n315) );
  INVX1_HVT U22 ( .A(n421), .Y(n455) );
  AND2X1_HVT U23 ( .A1(n216), .A2(n217), .Y(n5) );
  AND2X1_HVT U25 ( .A1(n318), .A2(n319), .Y(n19) );
  AND2X1_HVT U26 ( .A1(n280), .A2(n282), .Y(n23) );
  INVX1_HVT U27 ( .A(in[4]), .Y(n540) );
  INVX1_HVT U28 ( .A(n731), .Y(n517) );
  MUX21X2_HVT U29 ( .A1(n261), .A2(n398), .S0(n500), .Y(n731) );
  INVX1_HVT U30 ( .A(n333), .Y(n349) );
  NAND2X0_HVT U31 ( .A1(n418), .A2(n231), .Y(n33) );
  NAND2X0_HVT U32 ( .A1(n484), .A2(n336), .Y(n50) );
  NAND2X0_HVT U34 ( .A1(n33), .A2(n50), .Y(n762) );
  INVX1_HVT U35 ( .A(n224), .Y(n366) );
  MUX21X1_HVT U36 ( .A1(n730), .A2(n558), .S0(n480), .Y(n118) );
  MUX41X1_HVT U37 ( .A1(n736), .A3(n513), .A2(n758), .A4(n305), .S0(n421), 
        .S1(n509), .Y(n570) );
  MUX41X1_HVT U38 ( .A1(n522), .A3(n533), .A2(n409), .A4(n492), .S0(n479), 
        .S1(n264), .Y(n627) );
  NAND2X0_HVT U39 ( .A1(n278), .A2(n119), .Y(n210) );
  NAND2X0_HVT U40 ( .A1(n483), .A2(n500), .Y(n211) );
  NAND2X0_HVT U41 ( .A1(n210), .A2(n211), .Y(n748) );
  INVX0_HVT U43 ( .A(n500), .Y(n119) );
  MUX21X2_HVT U44 ( .A1(n357), .A2(n763), .S0(n365), .Y(n735) );
  NBUFFX2_HVT U45 ( .A(n236), .Y(n493) );
  MUX21X2_HVT U46 ( .A1(n391), .A2(n483), .S0(n453), .Y(n761) );
  NAND2X0_HVT U47 ( .A1(n444), .A2(n478), .Y(n212) );
  NAND2X0_HVT U48 ( .A1(n537), .A2(n252), .Y(n213) );
  NAND2X0_HVT U49 ( .A1(n212), .A2(n213), .Y(n704) );
  INVX0_HVT U50 ( .A(in[3]), .Y(n555) );
  INVX0_HVT U52 ( .A(n497), .Y(n418) );
  MUX41X1_HVT U54 ( .A1(n656), .A3(n642), .A2(n650), .A4(n637), .S0(n359), 
        .S1(n232), .Y(out[3]) );
  NAND2X0_HVT U55 ( .A1(n483), .A2(n433), .Y(n216) );
  NAND2X0_HVT U57 ( .A1(n458), .A2(n475), .Y(n217) );
  MUX41X1_HVT U59 ( .A1(n694), .A3(n696), .A2(n697), .A4(n701), .S0(n477), 
        .S1(n481), .Y(n693) );
  INVX1_HVT U60 ( .A(n362), .Y(n411) );
  MUX21X1_HVT U61 ( .A1(n485), .A2(n473), .S0(n358), .Y(n436) );
  INVX1_HVT U64 ( .A(n759), .Y(n550) );
  INVX1_HVT U65 ( .A(n505), .Y(n252) );
  MUX21X1_HVT U66 ( .A1(n565), .A2(n741), .S0(n445), .Y(n561) );
  INVX1_HVT U67 ( .A(n455), .Y(n429) );
  INVX0_HVT U68 ( .A(n510), .Y(n506) );
  INVX1_HVT U69 ( .A(n502), .Y(n350) );
  MUX21X1_HVT U70 ( .A1(n497), .A2(n491), .S0(n500), .Y(n740) );
  NBUFFX2_HVT U71 ( .A(n506), .Y(n480) );
  NBUFFX2_HVT U72 ( .A(n400), .Y(n365) );
  INVX1_HVT U74 ( .A(n300), .Y(n303) );
  INVX1_HVT U75 ( .A(n332), .Y(n333) );
  INVX1_HVT U76 ( .A(n475), .Y(n450) );
  MUX21X1_HVT U77 ( .A1(n487), .A2(n531), .S0(n453), .Y(n742) );
  MUX21X1_HVT U78 ( .A1(n551), .A2(n539), .S0(n433), .Y(n653) );
  INVX1_HVT U79 ( .A(n475), .Y(n433) );
  MUX21X1_HVT U81 ( .A1(n527), .A2(n649), .S0(n264), .Y(n648) );
  MUX21X1_HVT U82 ( .A1(n444), .A2(n560), .S0(n382), .Y(n443) );
  OA21X1_HVT U84 ( .A1(n514), .A2(n425), .A3(n377), .Y(n625) );
  OA21X1_HVT U85 ( .A1(n470), .A2(n414), .A3(n377), .Y(n600) );
  MUX21X1_HVT U87 ( .A1(n615), .A2(n614), .S0(n433), .Y(n613) );
  INVX1_HVT U88 ( .A(n751), .Y(n512) );
  INVX1_HVT U89 ( .A(n475), .Y(n344) );
  XOR2X1_HVT U91 ( .A1(n339), .A2(n326), .Y(n727) );
  MUX21X1_HVT U92 ( .A1(n692), .A2(n691), .S0(n476), .Y(n689) );
  XOR2X1_HVT U93 ( .A1(n453), .A2(n395), .Y(n724) );
  AO21X1_HVT U94 ( .A1(n238), .A2(n444), .A3(n382), .Y(n668) );
  INVX1_HVT U95 ( .A(n560), .Y(n530) );
  MUX21X1_HVT U96 ( .A1(n418), .A2(n224), .S0(n500), .Y(n609) );
  MUX21X1_HVT U97 ( .A1(n588), .A2(n589), .S0(n315), .Y(n587) );
  INVX1_HVT U98 ( .A(n297), .Y(n766) );
  INVX1_HVT U99 ( .A(n441), .Y(n454) );
  XOR2X1_HVT U100 ( .A1(n494), .A2(n365), .Y(n723) );
  INVX1_HVT U102 ( .A(n461), .Y(n425) );
  INVX0_HVT U104 ( .A(n365), .Y(n336) );
  INVX1_HVT U105 ( .A(n478), .Y(n245) );
  INVX1_HVT U106 ( .A(in[1]), .Y(n332) );
  INVX1_HVT U107 ( .A(n463), .Y(n430) );
  INVX1_HVT U108 ( .A(n482), .Y(n232) );
  INVX1_HVT U109 ( .A(n227), .Y(n335) );
  INVX0_HVT U111 ( .A(n349), .Y(n453) );
  INVX0_HVT U112 ( .A(n485), .Y(n442) );
  AND2X1_HVT U113 ( .A1(n330), .A2(n331), .Y(n218) );
  INVX1_HVT U114 ( .A(n553), .Y(n285) );
  AND2X1_HVT U116 ( .A1(n388), .A2(n389), .Y(n219) );
  AND2X1_HVT U117 ( .A1(n396), .A2(n397), .Y(n222) );
  INVX0_HVT U118 ( .A(n761), .Y(n537) );
  INVX0_HVT U119 ( .A(n313), .Y(n224) );
  INVX0_HVT U120 ( .A(n313), .Y(n314) );
  INVX0_HVT U121 ( .A(n333), .Y(n227) );
  INVX0_HVT U122 ( .A(n349), .Y(n500) );
  MUX41X1_HVT U124 ( .A1(n583), .A3(n586), .A2(n587), .A4(n590), .S0(n478), 
        .S1(n482), .Y(n582) );
  INVX0_HVT U126 ( .A(n426), .Y(n746) );
  MUX21X1_HVT U127 ( .A1(n669), .A2(n511), .S0(n347), .Y(n666) );
  INVX1_HVT U128 ( .A(n446), .Y(n726) );
  MUX41X1_HVT U129 ( .A1(n753), .A3(n687), .A2(n522), .A4(n381), .S0(n264), 
        .S1(n404), .Y(n686) );
  INVX0_HVT U130 ( .A(n357), .Y(n531) );
  INVX0_HVT U131 ( .A(n373), .Y(n473) );
  NBUFFX2_HVT U132 ( .A(n453), .Y(n231) );
  MUX21X1_HVT U133 ( .A1(n297), .A2(n742), .S0(n414), .Y(n626) );
  OR2X1_HVT U134 ( .A1(n350), .A2(n497), .Y(n685) );
  MUX41X1_HVT U136 ( .A1(n655), .A3(n757), .A2(n740), .A4(n426), .S0(n454), 
        .S1(n462), .Y(n654) );
  INVX1_HVT U137 ( .A(n439), .Y(n428) );
  INVX1_HVT U138 ( .A(n349), .Y(n401) );
  INVX1_HVT U139 ( .A(n732), .Y(n513) );
  INVX1_HVT U141 ( .A(n436), .Y(n750) );
  INVX0_HVT U142 ( .A(n362), .Y(n391) );
  INVX1_HVT U143 ( .A(n748), .Y(n522) );
  INVX0_HVT U144 ( .A(n760), .Y(n234) );
  INVX0_HVT U145 ( .A(n738), .Y(n551) );
  INVX0_HVT U146 ( .A(n510), .Y(n300) );
  INVX0_HVT U147 ( .A(n698), .Y(n553) );
  MUX41X1_HVT U148 ( .A1(n666), .A3(n663), .A2(n670), .A4(n665), .S0(n232), 
        .S1(n504), .Y(n662) );
  MUX41X1_HVT U149 ( .A1(n641), .A3(n639), .A2(n640), .A4(n638), .S0(n245), 
        .S1(n404), .Y(n637) );
  INVX1_HVT U150 ( .A(n324), .Y(n238) );
  INVX1_HVT U151 ( .A(n339), .Y(n324) );
  INVX1_HVT U152 ( .A(n373), .Y(n437) );
  INVX1_HVT U153 ( .A(n667), .Y(n523) );
  MUX41X1_HVT U155 ( .A1(n607), .A3(n602), .A2(n605), .A4(n599), .S0(n232), 
        .S1(n245), .Y(n598) );
  INVX0_HVT U156 ( .A(n490), .Y(n395) );
  INVX0_HVT U157 ( .A(n409), .Y(n381) );
  INVX1_HVT U160 ( .A(n451), .Y(n763) );
  MUX41X1_HVT U161 ( .A1(n751), .A3(n524), .A2(n759), .A4(n716), .S0(n430), 
        .S1(n477), .Y(n714) );
  INVX1_HVT U163 ( .A(n449), .Y(n757) );
  NBUFFX4_HVT U164 ( .A(n427), .Y(n483) );
  MUX41X1_HVT U169 ( .A1(n761), .A3(n464), .A2(n520), .A4(n757), .S0(n315), 
        .S1(n445), .Y(n592) );
  MUX21X1_HVT U170 ( .A1(n490), .A2(n552), .S0(n501), .Y(n759) );
  MUX21X1_HVT U171 ( .A1(n531), .A2(n473), .S0(n501), .Y(n597) );
  INVX0_HVT U172 ( .A(n390), .Y(n736) );
  INVX0_HVT U173 ( .A(n446), .Y(n249) );
  OR2X1_HVT U175 ( .A1(n304), .A2(n540), .Y(n768) );
  NBUFFX2_HVT U176 ( .A(n767), .Y(n261) );
  MUX41X1_HVT U178 ( .A1(n580), .A3(n578), .A2(n579), .A4(n575), .S0(n232), 
        .S1(n252), .Y(n574) );
  INVX0_HVT U180 ( .A(n758), .Y(n536) );
  NAND2X0_HVT U181 ( .A1(n394), .A2(n264), .Y(n271) );
  NAND2X0_HVT U183 ( .A1(n466), .A2(n433), .Y(n273) );
  NAND2X0_HVT U184 ( .A1(n271), .A2(n273), .Y(n639) );
  INVX0_HVT U185 ( .A(n440), .Y(n264) );
  INVX0_HVT U186 ( .A(n400), .Y(n339) );
  XNOR2X1_HVT U187 ( .A1(n462), .A2(n744), .Y(n728) );
  NAND2X0_HVT U188 ( .A1(n439), .A2(n555), .Y(n760) );
  NAND2X0_HVT U190 ( .A1(n601), .A2(n455), .Y(n274) );
  NAND2X0_HVT U191 ( .A1(n600), .A2(n347), .Y(n275) );
  NAND2X0_HVT U192 ( .A1(n274), .A2(n275), .Y(n599) );
  INVX0_HVT U193 ( .A(n740), .Y(n549) );
  MUX21X1_HVT U194 ( .A1(n552), .A2(n489), .S0(n365), .Y(n738) );
  INVX1_HVT U195 ( .A(n497), .Y(n552) );
  MUX41X1_HVT U196 ( .A1(n569), .A3(n568), .A2(n571), .A4(n570), .S0(n252), 
        .S1(n481), .Y(n567) );
  MUX41X1_HVT U198 ( .A1(n595), .A3(n752), .A2(n734), .A4(n542), .S0(n344), 
        .S1(n507), .Y(n594) );
  MUX21X1_HVT U199 ( .A1(n391), .A2(n493), .S0(n452), .Y(n682) );
  MUX21X1_HVT U200 ( .A1(n492), .A2(n409), .S0(n452), .Y(n664) );
  INVX0_HVT U201 ( .A(in[3]), .Y(n304) );
  MUX41X1_HVT U202 ( .A1(n593), .A3(n596), .A2(n592), .A4(n594), .S0(n481), 
        .S1(n245), .Y(n591) );
  INVX0_HVT U203 ( .A(n742), .Y(n526) );
  MUX41X1_HVT U204 ( .A1(n613), .A3(n618), .A2(n611), .A4(n617), .S0(n481), 
        .S1(n245), .Y(n610) );
  INVX0_HVT U205 ( .A(n715), .Y(n548) );
  MUX41X1_HVT U206 ( .A1(n528), .A3(n746), .A2(n222), .A4(n629), .S0(n344), 
        .S1(n463), .Y(n628) );
  NAND2X0_HVT U207 ( .A1(n328), .A2(n329), .Y(n278) );
  INVX1_HVT U209 ( .A(n440), .Y(n503) );
  NAND2X0_HVT U210 ( .A1(n437), .A2(n279), .Y(n280) );
  NAND2X0_HVT U211 ( .A1(n5), .A2(n474), .Y(n282) );
  INVX1_HVT U213 ( .A(n474), .Y(n279) );
  MUX41X1_HVT U216 ( .A1(n581), .A3(n723), .A2(n737), .A4(n730), .S0(n450), 
        .S1(n303), .Y(n580) );
  NAND2X0_HVT U217 ( .A1(n550), .A2(n505), .Y(n283) );
  NAND2X0_HVT U219 ( .A1(n283), .A2(n285), .Y(n705) );
  MUX21X2_HVT U221 ( .A1(n552), .A2(n531), .S0(n358), .Y(n734) );
  NAND2X0_HVT U222 ( .A1(n659), .A2(n347), .Y(n289) );
  NAND2X0_HVT U223 ( .A1(n433), .A2(n740), .Y(n291) );
  NAND2X0_HVT U224 ( .A1(n289), .A2(n291), .Y(n657) );
  NAND2X0_HVT U225 ( .A1(n222), .A2(n264), .Y(n293) );
  NAND2X0_HVT U226 ( .A1(n752), .A2(n433), .Y(n296) );
  NAND2X0_HVT U227 ( .A1(n293), .A2(n296), .Y(n638) );
  INVX0_HVT U228 ( .A(n415), .Y(n752) );
  INVX1_HVT U229 ( .A(n562), .Y(n546) );
  AND2X1_HVT U230 ( .A1(n358), .A2(n495), .Y(n297) );
  MUX41X1_HVT U231 ( .A1(n706), .A3(n705), .A2(n704), .A4(n521), .S0(n312), 
        .S1(n344), .Y(n703) );
  INVX1_HVT U232 ( .A(n509), .Y(n312) );
  INVX1_HVT U233 ( .A(n304), .Y(n405) );
  AO21X1_HVT U234 ( .A1(n463), .A2(n677), .A3(n545), .Y(n678) );
  INVX1_HVT U235 ( .A(n677), .Y(n532) );
  INVX1_HVT U236 ( .A(n414), .Y(n422) );
  MUX41X1_HVT U237 ( .A1(n703), .A3(n711), .A2(n707), .A4(n717), .S0(n334), 
        .S1(n482), .Y(out[0]) );
  MUX41X1_HVT U238 ( .A1(n631), .A3(n633), .A2(n634), .A4(n635), .S0(n505), 
        .S1(n482), .Y(n630) );
  MUX21X1_HVT U239 ( .A1(n492), .A2(n399), .S0(n339), .Y(n415) );
  NAND2X0_HVT U240 ( .A1(n396), .A2(n397), .Y(n305) );
  INVX1_HVT U242 ( .A(n398), .Y(n313) );
  NAND2X0_HVT U243 ( .A1(n467), .A2(n306), .Y(n307) );
  NAND2X0_HVT U244 ( .A1(n671), .A2(n725), .Y(n308) );
  NAND2X0_HVT U246 ( .A1(n307), .A2(n308), .Y(n670) );
  INVX0_HVT U247 ( .A(n725), .Y(n306) );
  NAND2X0_HVT U248 ( .A1(n496), .A2(n119), .Y(n309) );
  NAND2X0_HVT U249 ( .A1(n325), .A2(n350), .Y(n310) );
  NAND2X0_HVT U250 ( .A1(n309), .A2(n310), .Y(n755) );
  MUX21X1_HVT U251 ( .A1(n549), .A2(n755), .S0(n476), .Y(n671) );
  XOR2X1_HVT U252 ( .A1(n476), .A2(n462), .Y(n725) );
  INVX0_HVT U253 ( .A(n755), .Y(n518) );
  INVX0_HVT U254 ( .A(n278), .Y(n311) );
  MUX41X1_HVT U255 ( .A1(n754), .A3(n231), .A2(n468), .A4(n548), .S0(n433), 
        .S1(n312), .Y(n673) );
  MUX41X1_HVT U257 ( .A1(n664), .A3(n534), .A2(n544), .A4(n724), .S0(n476), 
        .S1(n312), .Y(n663) );
  INVX0_HVT U258 ( .A(n743), .Y(n544) );
  INVX1_HVT U259 ( .A(n443), .Y(n636) );
  MUX21X1_HVT U260 ( .A1(n685), .A2(n395), .S0(n479), .Y(n589) );
  INVX0_HVT U261 ( .A(n332), .Y(n400) );
  INVX1_HVT U263 ( .A(n332), .Y(n452) );
  MUX41X1_HVT U266 ( .A1(n219), .A3(n381), .A2(n735), .A4(n499), .S0(n344), 
        .S1(n507), .Y(n578) );
  MUX41X1_HVT U267 ( .A1(n285), .A3(n515), .A2(n726), .A4(n548), .S0(n344), 
        .S1(n461), .Y(n623) );
  XNOR2X1_HVT U269 ( .A1(n411), .A2(n452), .Y(n466) );
  NAND2X0_HVT U271 ( .A1(n765), .A2(n315), .Y(n316) );
  NAND2X0_HVT U272 ( .A1(n632), .A2(n344), .Y(n317) );
  NAND2X0_HVT U273 ( .A1(n316), .A2(n317), .Y(n631) );
  OR2X1_HVT U274 ( .A1(n442), .A2(n350), .Y(n737) );
  NAND2X0_HVT U275 ( .A1(n547), .A2(n324), .Y(n318) );
  NAND2X0_HVT U279 ( .A1(n366), .A2(n238), .Y(n319) );
  INVX1_HVT U280 ( .A(n493), .Y(n547) );
  MUX41X1_HVT U281 ( .A1(n624), .A3(n628), .A2(n623), .A4(n627), .S0(n482), 
        .S1(n252), .Y(n622) );
  INVX1_HVT U282 ( .A(n754), .Y(n519) );
  INVX0_HVT U283 ( .A(n753), .Y(n394) );
  NAND2X0_HVT U285 ( .A1(n582), .A2(n359), .Y(n320) );
  NAND2X0_HVT U286 ( .A1(n591), .A2(n334), .Y(n321) );
  NAND2X0_HVT U287 ( .A1(n321), .A2(n320), .Y(out[6]) );
  NAND2X0_HVT U288 ( .A1(n325), .A2(n462), .Y(n322) );
  NAND2X0_HVT U289 ( .A1(n750), .A2(n382), .Y(n323) );
  NAND2X0_HVT U290 ( .A1(n322), .A2(n323), .Y(n692) );
  MUX41X1_HVT U291 ( .A1(n487), .A3(n597), .A2(n523), .A4(n756), .S0(n422), 
        .S1(n264), .Y(n596) );
  MUX21X1_HVT U292 ( .A1(n224), .A2(n399), .S0(n324), .Y(n667) );
  NBUFFX2_HVT U293 ( .A(n236), .Y(n325) );
  NBUFFX2_HVT U296 ( .A(n760), .Y(n326) );
  NBUFFX2_HVT U297 ( .A(in[5]), .Y(n505) );
  XNOR2X2_HVT U298 ( .A1(n486), .A2(n405), .Y(n398) );
  NBUFFX2_HVT U299 ( .A(n398), .Y(n484) );
  MUX21X1_HVT U300 ( .A1(n489), .A2(n451), .S0(n339), .Y(n753) );
  NAND2X0_HVT U301 ( .A1(n486), .A2(n405), .Y(n328) );
  NAND2X0_HVT U303 ( .A1(n327), .A2(n439), .Y(n329) );
  NAND2X0_HVT U304 ( .A1(n328), .A2(n329), .Y(n451) );
  INVX0_HVT U305 ( .A(n405), .Y(n327) );
  NAND2X0_HVT U307 ( .A1(n489), .A2(n502), .Y(n330) );
  NAND2X0_HVT U308 ( .A1(n311), .A2(n387), .Y(n331) );
  INVX1_HVT U309 ( .A(in[7]), .Y(n510) );
  MUX41X1_HVT U310 ( .A1(n436), .A3(n727), .A2(n755), .A4(n556), .S0(n455), 
        .S1(n422), .Y(n688) );
  INVX1_HVT U311 ( .A(n440), .Y(n441) );
  MUX21X2_HVT U312 ( .A1(n390), .A2(n766), .S0(n421), .Y(n661) );
  AND3X1_HVT U313 ( .A1(n475), .A2(n238), .A3(n458), .Y(n640) );
  INVX0_HVT U314 ( .A(in[2]), .Y(n440) );
  INVX1_HVT U315 ( .A(n359), .Y(n334) );
  INVX1_HVT U316 ( .A(in[6]), .Y(n359) );
  MUX21X1_HVT U317 ( .A1(n547), .A2(n437), .S0(n350), .Y(n606) );
  MUX41X1_HVT U318 ( .A1(n19), .A3(n326), .A2(n731), .A4(n744), .S0(n461), 
        .S1(n378), .Y(n579) );
  MUX41X1_HVT U319 ( .A1(n608), .A3(n415), .A2(n609), .A4(n466), .S0(n455), 
        .S1(n508), .Y(n607) );
  NAND2X0_HVT U320 ( .A1(n647), .A2(n422), .Y(n337) );
  NAND2X0_HVT U321 ( .A1(n648), .A2(n382), .Y(n338) );
  NAND2X0_HVT U322 ( .A1(n337), .A2(n338), .Y(n644) );
  INVX1_HVT U323 ( .A(n555), .Y(n427) );
  MUX41X1_HVT U324 ( .A1(n689), .A3(n686), .A2(n688), .A4(n684), .S0(n232), 
        .S1(n245), .Y(n683) );
  INVX1_HVT U325 ( .A(n540), .Y(n439) );
  MUX41X1_HVT U326 ( .A1(n468), .A3(n556), .A2(n675), .A4(n219), .S0(n378), 
        .S1(n508), .Y(n674) );
  INVX1_HVT U327 ( .A(n763), .Y(n409) );
  NAND2X0_HVT U328 ( .A1(n413), .A2(n412), .Y(n635) );
  NBUFFX2_HVT U329 ( .A(n540), .Y(n485) );
  NBUFFX2_HVT U330 ( .A(n540), .Y(n486) );
  NAND2X0_HVT U331 ( .A1(n399), .A2(n339), .Y(n340) );
  NAND2X0_HVT U332 ( .A1(n497), .A2(n452), .Y(n341) );
  NAND2X0_HVT U333 ( .A1(n340), .A2(n341), .Y(n390) );
  NAND2X0_HVT U334 ( .A1(n491), .A2(n238), .Y(n342) );
  NAND2X0_HVT U335 ( .A1(n391), .A2(n358), .Y(n343) );
  NAND2X0_HVT U336 ( .A1(n342), .A2(n343), .Y(n438) );
  NAND2X0_HVT U337 ( .A1(n501), .A2(n499), .Y(n698) );
  NAND2X0_HVT U338 ( .A1(n544), .A2(n433), .Y(n345) );
  NAND2X0_HVT U339 ( .A1(n741), .A2(n475), .Y(n346) );
  NAND2X0_HVT U340 ( .A1(n345), .A2(n346), .Y(n641) );
  MUX21X1_HVT U341 ( .A1(n489), .A2(n442), .S0(n501), .Y(n741) );
  NAND2X0_HVT U342 ( .A1(n347), .A2(n735), .Y(n348) );
  AND2X1_HVT U343 ( .A1(n348), .A2(n438), .Y(n660) );
  INVX0_HVT U344 ( .A(n454), .Y(n347) );
  XOR2X1_HVT U345 ( .A1(n442), .A2(n502), .Y(n745) );
  MUX21X1_HVT U346 ( .A1(n483), .A2(n410), .S0(n452), .Y(n733) );
  MUX41X1_HVT U347 ( .A1(n713), .A3(n472), .A2(n438), .A4(n470), .S0(n425), 
        .S1(n477), .Y(n712) );
  NAND2X0_HVT U348 ( .A1(n720), .A2(n414), .Y(n351) );
  NAND2X0_HVT U349 ( .A1(n721), .A2(n463), .Y(n352) );
  NAND2X0_HVT U350 ( .A1(n351), .A2(n352), .Y(n718) );
  NAND2X0_HVT U351 ( .A1(n722), .A2(n315), .Y(n353) );
  NAND2X0_HVT U352 ( .A1(n718), .A2(n450), .Y(n354) );
  NAND2X0_HVT U353 ( .A1(n353), .A2(n354), .Y(n717) );
  MUX21X1_HVT U354 ( .A1(n483), .A2(n737), .S0(n505), .Y(n721) );
  NAND2X0_HVT U355 ( .A1(n708), .A2(n344), .Y(n355) );
  NAND2X0_HVT U356 ( .A1(n710), .A2(n315), .Y(n356) );
  NAND2X0_HVT U357 ( .A1(n355), .A2(n356), .Y(n707) );
  INVX0_HVT U358 ( .A(n480), .Y(n382) );
  NAND2X0_HVT U359 ( .A1(n485), .A2(n488), .Y(n357) );
  NBUFFX2_HVT U360 ( .A(n400), .Y(n358) );
  NAND2X0_HVT U361 ( .A1(n567), .A2(n359), .Y(n360) );
  NAND2X0_HVT U362 ( .A1(n574), .A2(n334), .Y(n361) );
  NAND2X0_HVT U363 ( .A1(n360), .A2(n361), .Y(out[7]) );
  AND2X1_HVT U364 ( .A1(n486), .A2(n488), .Y(n362) );
  NAND2X0_HVT U365 ( .A1(n576), .A2(n315), .Y(n363) );
  NAND2X0_HVT U366 ( .A1(n577), .A2(n378), .Y(n364) );
  NAND2X0_HVT U367 ( .A1(n363), .A2(n364), .Y(n575) );
  INVX1_HVT U368 ( .A(n480), .Y(n414) );
  NAND2X0_HVT U369 ( .A1(n610), .A2(in[6]), .Y(n367) );
  NAND2X0_HVT U370 ( .A1(n598), .A2(n359), .Y(n368) );
  NAND2X0_HVT U371 ( .A1(n368), .A2(n367), .Y(out[5]) );
  NAND2X0_HVT U372 ( .A1(n651), .A2(n245), .Y(n369) );
  NAND2X0_HVT U373 ( .A1(n654), .A2(n505), .Y(n370) );
  NAND2X0_HVT U374 ( .A1(n369), .A2(n370), .Y(n650) );
  MUX21X1_HVT U375 ( .A1(n536), .A2(n502), .S0(n505), .Y(n706) );
  MUX41X1_HVT U376 ( .A1(n657), .A3(n660), .A2(n23), .A4(n661), .S0(n505), 
        .S1(n404), .Y(n656) );
  NAND2X0_HVT U377 ( .A1(n620), .A2(n450), .Y(n371) );
  NAND2X0_HVT U378 ( .A1(n621), .A2(n476), .Y(n372) );
  NAND2X0_HVT U379 ( .A1(n371), .A2(n372), .Y(n618) );
  MUX21X1_HVT U380 ( .A1(n218), .A2(n444), .S0(n463), .Y(n621) );
  NAND2X0_HVT U381 ( .A1(n428), .A2(n427), .Y(n373) );
  INVX1_HVT U382 ( .A(n349), .Y(n501) );
  NAND2X0_HVT U383 ( .A1(n616), .A2(n374), .Y(n375) );
  NAND2X0_HVT U384 ( .A1(n496), .A2(n471), .Y(n376) );
  NAND2X0_HVT U385 ( .A1(n375), .A2(n376), .Y(n615) );
  INVX0_HVT U386 ( .A(n471), .Y(n374) );
  INVX1_HVT U387 ( .A(n549), .Y(n377) );
  NAND2X0_HVT U388 ( .A1(n678), .A2(n378), .Y(n379) );
  NAND2X0_HVT U389 ( .A1(n679), .A2(n476), .Y(n380) );
  NAND2X0_HVT U390 ( .A1(n379), .A2(n380), .Y(n676) );
  INVX0_HVT U391 ( .A(n476), .Y(n378) );
  NAND2X0_HVT U392 ( .A1(n622), .A2(n359), .Y(n402) );
  NAND2X0_HVT U393 ( .A1(n492), .A2(n238), .Y(n383) );
  NAND2X0_HVT U394 ( .A1(n399), .A2(n401), .Y(n384) );
  NAND2X0_HVT U395 ( .A1(n383), .A2(n384), .Y(n700) );
  NAND2X0_HVT U396 ( .A1(n728), .A2(n450), .Y(n385) );
  NAND2X0_HVT U397 ( .A1(n702), .A2(n315), .Y(n386) );
  NAND2X0_HVT U398 ( .A1(n385), .A2(n386), .Y(n701) );
  NAND2X0_HVT U399 ( .A1(n489), .A2(n387), .Y(n388) );
  NAND2X0_HVT U400 ( .A1(n325), .A2(n119), .Y(n389) );
  INVX0_HVT U401 ( .A(n339), .Y(n387) );
  MUX21X1_HVT U402 ( .A1(n418), .A2(n219), .S0(n462), .Y(n702) );
  INVX1_HVT U403 ( .A(n487), .Y(n458) );
  MUX21X2_HVT U404 ( .A1(n532), .A2(n734), .S0(n445), .Y(n614) );
  NAND2X0_HVT U405 ( .A1(n496), .A2(n374), .Y(n392) );
  NAND2X0_HVT U406 ( .A1(n680), .A2(n471), .Y(n393) );
  NAND2X0_HVT U407 ( .A1(n393), .A2(n392), .Y(n679) );
  INVX1_HVT U408 ( .A(n480), .Y(n445) );
  NBUFFX2_HVT U409 ( .A(n503), .Y(n475) );
  NAND2X0_HVT U410 ( .A1(n442), .A2(n324), .Y(n396) );
  NAND2X0_HVT U411 ( .A1(n531), .A2(n227), .Y(n397) );
  NBUFFX2_HVT U412 ( .A(n555), .Y(n488) );
  INVX1_HVT U413 ( .A(n558), .Y(n542) );
  OA21X1_HVT U414 ( .A1(n732), .A2(n430), .A3(n619), .Y(n620) );
  NBUFFX2_HVT U415 ( .A(n485), .Y(n399) );
  MUX41X1_HVT U416 ( .A1(n415), .A3(n409), .A2(n467), .A4(n394), .S0(n477), 
        .S1(n425), .Y(n710) );
  NAND2X0_HVT U417 ( .A1(n630), .A2(n334), .Y(n403) );
  NAND2X0_HVT U418 ( .A1(n402), .A2(n403), .Y(out[4]) );
  XOR2X1_HVT U419 ( .A1(n506), .A2(n358), .Y(n471) );
  AO21X1_HVT U420 ( .A1(n476), .A2(n491), .A3(n381), .Y(n652) );
  INVX1_HVT U421 ( .A(n362), .Y(n406) );
  NAND2X0_HVT U422 ( .A1(n714), .A2(n429), .Y(n407) );
  NAND2X0_HVT U423 ( .A1(n712), .A2(n450), .Y(n408) );
  NAND2X0_HVT U424 ( .A1(n407), .A2(n408), .Y(n711) );
  OA21X1_HVT U425 ( .A1(n414), .A2(n762), .A3(n528), .Y(n572) );
  MUX41X1_HVT U426 ( .A1(n757), .A3(n716), .A2(n748), .A4(n551), .S0(n344), 
        .S1(n509), .Y(n569) );
  INVX0_HVT U427 ( .A(n406), .Y(n410) );
  NAND2X0_HVT U428 ( .A1(n636), .A2(n347), .Y(n412) );
  NAND2X0_HVT U429 ( .A1(n511), .A2(n450), .Y(n413) );
  NAND2X0_HVT U430 ( .A1(n625), .A2(n315), .Y(n416) );
  NAND2X0_HVT U431 ( .A1(n626), .A2(n450), .Y(n417) );
  NAND2X0_HVT U432 ( .A1(n416), .A2(n417), .Y(n624) );
  NBUFFX2_HVT U433 ( .A(n768), .Y(n498) );
  INVX1_HVT U434 ( .A(n563), .Y(n524) );
  NAND2X0_HVT U435 ( .A1(n572), .A2(n378), .Y(n419) );
  NAND2X0_HVT U436 ( .A1(n573), .A2(n429), .Y(n420) );
  NAND2X0_HVT U437 ( .A1(n420), .A2(n419), .Y(n571) );
  NAND2X0_HVT U438 ( .A1(n473), .A2(n336), .Y(n423) );
  NAND2X0_HVT U439 ( .A1(n552), .A2(n453), .Y(n424) );
  NAND2X0_HVT U440 ( .A1(n423), .A2(n424), .Y(n744) );
  INVX0_HVT U441 ( .A(n658), .Y(n533) );
  NBUFFX2_HVT U442 ( .A(n540), .Y(n487) );
  INVX1_HVT U443 ( .A(n559), .Y(n515) );
  NAND2X0_HVT U444 ( .A1(n652), .A2(n430), .Y(n431) );
  NAND2X0_HVT U445 ( .A1(n653), .A2(n463), .Y(n432) );
  NAND2X0_HVT U446 ( .A1(n431), .A2(n432), .Y(n651) );
  NAND2X0_HVT U447 ( .A1(n643), .A2(n252), .Y(n434) );
  NAND2X0_HVT U448 ( .A1(n644), .A2(n505), .Y(n435) );
  NAND2X0_HVT U449 ( .A1(n434), .A2(n435), .Y(n642) );
  MUX41X1_HVT U450 ( .A1(n736), .A3(n515), .A2(n739), .A4(n465), .S0(n450), 
        .S1(n382), .Y(n633) );
  MUX41X1_HVT U451 ( .A1(n761), .A3(n532), .A2(n695), .A4(n218), .S0(n479), 
        .S1(n441), .Y(n694) );
  NAND2X0_HVT U452 ( .A1(n447), .A2(n448), .Y(out[1]) );
  INVX1_HVT U453 ( .A(n561), .Y(n511) );
  NAND2X0_HVT U454 ( .A1(n693), .A2(n334), .Y(n447) );
  NAND2X0_HVT U455 ( .A1(n683), .A2(n359), .Y(n448) );
  AND2X1_HVT U456 ( .A1(n756), .A2(n499), .Y(n449) );
  MUX41X1_HVT U457 ( .A1(n546), .A3(n548), .A2(n426), .A4(n437), .S0(n450), 
        .S1(n507), .Y(n696) );
  MUX41X1_HVT U458 ( .A1(n659), .A3(n261), .A2(n467), .A4(n539), .S0(n508), 
        .S1(n421), .Y(n617) );
  MUX41X1_HVT U459 ( .A1(n745), .A3(n700), .A2(n747), .A4(n699), .S0(n450), 
        .S1(n507), .Y(n697) );
  MUX41X1_HVT U460 ( .A1(n549), .A3(n541), .A2(n766), .A4(n458), .S0(n454), 
        .S1(n445), .Y(n568) );
  NAND2X0_HVT U461 ( .A1(n456), .A2(n457), .Y(out[2]) );
  OA21X1_HVT U462 ( .A1(n414), .A2(n738), .A3(n522), .Y(n588) );
  MUX41X1_HVT U463 ( .A1(n726), .A3(n285), .A2(n733), .A4(n468), .S0(n454), 
        .S1(n430), .Y(n586) );
  NAND2X0_HVT U464 ( .A1(n662), .A2(n359), .Y(n456) );
  NAND2X0_HVT U465 ( .A1(n672), .A2(n334), .Y(n457) );
  MUX41X1_HVT U466 ( .A1(n674), .A3(n681), .A2(n673), .A4(n676), .S0(n481), 
        .S1(n245), .Y(n672) );
  NAND2X0_HVT U467 ( .A1(n529), .A2(n463), .Y(n459) );
  NAND2X0_HVT U468 ( .A1(n748), .A2(n425), .Y(n460) );
  NAND2X0_HVT U469 ( .A1(n459), .A2(n460), .Y(n632) );
  NBUFFX2_HVT U470 ( .A(n506), .Y(n461) );
  NBUFFX2_HVT U471 ( .A(n506), .Y(n462) );
  NBUFFX2_HVT U472 ( .A(n506), .Y(n463) );
  AND2X1_HVT U473 ( .A1(n224), .A2(n715), .Y(n464) );
  MUX21X1_HVT U474 ( .A1(n410), .A2(n418), .S0(n505), .Y(n719) );
  AND2X1_HVT U475 ( .A1(n494), .A2(n698), .Y(n465) );
  MUX21X1_HVT U476 ( .A1(n410), .A2(n399), .S0(n401), .Y(n560) );
  NBUFFX2_HVT U477 ( .A(n767), .Y(n494) );
  MUX21X1_HVT U478 ( .A1(n490), .A2(n437), .S0(n401), .Y(n732) );
  MUX21X1_HVT U479 ( .A1(n487), .A2(n490), .S0(n335), .Y(n649) );
  NBUFFX2_HVT U480 ( .A(n767), .Y(n495) );
  MUX21X1_HVT U481 ( .A1(n488), .A2(n485), .S0(n452), .Y(n581) );
  NBUFFX2_HVT U482 ( .A(n373), .Y(n496) );
  MUX21X1_HVT U483 ( .A1(n261), .A2(n411), .S0(n335), .Y(n559) );
  MUX21X1_HVT U484 ( .A1(n391), .A2(n499), .S0(n401), .Y(n677) );
  MUX21X1_HVT U485 ( .A1(n261), .A2(n399), .S0(n365), .Y(n564) );
  AND2X1_HVT U486 ( .A1(n498), .A2(n658), .Y(n467) );
  AND2X1_HVT U487 ( .A1(n452), .A2(n437), .Y(n468) );
  XNOR2X1_HVT U488 ( .A1(n498), .A2(n335), .Y(n469) );
  MUX21X1_HVT U489 ( .A1(n325), .A2(n499), .S0(n503), .Y(n646) );
  NBUFFX2_HVT U490 ( .A(in[2]), .Y(n476) );
  NBUFFX2_HVT U491 ( .A(n327), .Y(n489) );
  NBUFFX2_HVT U492 ( .A(n304), .Y(n490) );
  NBUFFX2_HVT U493 ( .A(n506), .Y(n479) );
  NBUFFX2_HVT U494 ( .A(n504), .Y(n478) );
  NBUFFX2_HVT U495 ( .A(n504), .Y(n477) );
  MUX21X1_HVT U496 ( .A1(n326), .A2(n219), .S0(n479), .Y(n601) );
  NAND2X0_HVT U497 ( .A1(n427), .A2(n428), .Y(n767) );
  AND2X1_HVT U498 ( .A1(n484), .A2(n502), .Y(n470) );
  MUX21X1_HVT U499 ( .A1(n473), .A2(n483), .S0(n335), .Y(n751) );
  MUX21X1_HVT U500 ( .A1(n766), .A2(n238), .S0(n503), .Y(n645) );
  NBUFFX2_HVT U501 ( .A(n768), .Y(n497) );
  NBUFFX2_HVT U502 ( .A(n236), .Y(n491) );
  MUX21X1_HVT U503 ( .A1(n483), .A2(n547), .S0(n387), .Y(n562) );
  XOR2X1_HVT U504 ( .A1(n231), .A2(n478), .Y(n729) );
  NBUFFX2_HVT U505 ( .A(n768), .Y(n499) );
  MUX21X1_HVT U506 ( .A1(n483), .A2(n487), .S0(n480), .Y(n680) );
  AND2X1_HVT U507 ( .A1(n490), .A2(n336), .Y(n472) );
  NBUFFX2_HVT U508 ( .A(in[5]), .Y(n504) );
  MUX21X1_HVT U509 ( .A1(n311), .A2(n487), .S0(n401), .Y(n695) );
  MUX21X1_HVT U510 ( .A1(n458), .A2(n763), .S0(n335), .Y(n563) );
  MUX21X1_HVT U511 ( .A1(n490), .A2(n499), .S0(n500), .Y(n584) );
  MUX21X1_HVT U512 ( .A1(n498), .A2(n261), .S0(n452), .Y(n585) );
  MUX21X1_HVT U513 ( .A1(n498), .A2(n458), .S0(n387), .Y(n743) );
  MUX21X1_HVT U514 ( .A1(n442), .A2(n326), .S0(n358), .Y(n558) );
  MUX21X1_HVT U515 ( .A1(n458), .A2(n499), .S0(n501), .Y(n557) );
  NBUFFX2_HVT U516 ( .A(in[0]), .Y(n481) );
  NBUFFX2_HVT U517 ( .A(in[0]), .Y(n482) );
  XNOR2X1_HVT U518 ( .A1(n501), .A2(n441), .Y(n474) );
endmodule

