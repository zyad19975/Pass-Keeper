
module reg_D_0 ( clk, rst, enable, in, out );
  input [127:0] in;
  output [127:0] out;
  input clk, rst, enable;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n130, n1, n129, n131, n132, n133,
         n134, n135, n136, n137, n138, n139;

  DFFARX1_HVT \out_reg[127]  ( .D(n130), .CLK(clk), .RSTB(n138), .Q(out[127])
         );
  DFFARX1_HVT \out_reg[126]  ( .D(n128), .CLK(clk), .RSTB(n138), .Q(out[126])
         );
  DFFARX1_HVT \out_reg[125]  ( .D(n127), .CLK(clk), .RSTB(n138), .Q(out[125])
         );
  DFFARX1_HVT \out_reg[124]  ( .D(n126), .CLK(clk), .RSTB(n138), .Q(out[124])
         );
  DFFARX1_HVT \out_reg[123]  ( .D(n125), .CLK(clk), .RSTB(n138), .Q(out[123])
         );
  DFFARX1_HVT \out_reg[122]  ( .D(n124), .CLK(clk), .RSTB(n129), .Q(out[122])
         );
  DFFARX1_HVT \out_reg[121]  ( .D(n123), .CLK(clk), .RSTB(n129), .Q(out[121])
         );
  DFFARX1_HVT \out_reg[120]  ( .D(n122), .CLK(clk), .RSTB(n139), .Q(out[120])
         );
  DFFARX1_HVT \out_reg[119]  ( .D(n121), .CLK(clk), .RSTB(n138), .Q(out[119])
         );
  DFFARX1_HVT \out_reg[118]  ( .D(n120), .CLK(clk), .RSTB(n138), .Q(out[118])
         );
  DFFARX1_HVT \out_reg[117]  ( .D(n119), .CLK(clk), .RSTB(n138), .Q(out[117])
         );
  DFFARX1_HVT \out_reg[116]  ( .D(n118), .CLK(clk), .RSTB(n138), .Q(out[116])
         );
  DFFARX1_HVT \out_reg[115]  ( .D(n117), .CLK(clk), .RSTB(n138), .Q(out[115])
         );
  DFFARX1_HVT \out_reg[114]  ( .D(n116), .CLK(clk), .RSTB(n131), .Q(out[114])
         );
  DFFARX1_HVT \out_reg[113]  ( .D(n115), .CLK(clk), .RSTB(n132), .Q(out[113])
         );
  DFFARX1_HVT \out_reg[112]  ( .D(n114), .CLK(clk), .RSTB(n133), .Q(out[112])
         );
  DFFARX1_HVT \out_reg[111]  ( .D(n113), .CLK(clk), .RSTB(n134), .Q(out[111])
         );
  DFFARX1_HVT \out_reg[110]  ( .D(n112), .CLK(clk), .RSTB(n135), .Q(out[110])
         );
  DFFARX1_HVT \out_reg[109]  ( .D(n111), .CLK(clk), .RSTB(n1), .Q(out[109]) );
  DFFARX1_HVT \out_reg[108]  ( .D(n110), .CLK(clk), .RSTB(n1), .Q(out[108]) );
  DFFARX1_HVT \out_reg[107]  ( .D(n109), .CLK(clk), .RSTB(n1), .Q(out[107]) );
  DFFARX1_HVT \out_reg[106]  ( .D(n108), .CLK(clk), .RSTB(n1), .Q(out[106]) );
  DFFARX1_HVT \out_reg[105]  ( .D(n107), .CLK(clk), .RSTB(n1), .Q(out[105]) );
  DFFARX1_HVT \out_reg[104]  ( .D(n106), .CLK(clk), .RSTB(n1), .Q(out[104]) );
  DFFARX1_HVT \out_reg[103]  ( .D(n105), .CLK(clk), .RSTB(n1), .Q(out[103]) );
  DFFARX1_HVT \out_reg[102]  ( .D(n104), .CLK(clk), .RSTB(n1), .Q(out[102]) );
  DFFARX1_HVT \out_reg[101]  ( .D(n103), .CLK(clk), .RSTB(n1), .Q(out[101]) );
  DFFARX1_HVT \out_reg[100]  ( .D(n102), .CLK(clk), .RSTB(n1), .Q(out[100]) );
  DFFARX1_HVT \out_reg[99]  ( .D(n101), .CLK(clk), .RSTB(n138), .Q(out[99]) );
  DFFARX1_HVT \out_reg[98]  ( .D(n100), .CLK(clk), .RSTB(n138), .Q(out[98]) );
  DFFARX1_HVT \out_reg[97]  ( .D(n99), .CLK(clk), .RSTB(n137), .Q(out[97]) );
  DFFARX1_HVT \out_reg[96]  ( .D(n98), .CLK(clk), .RSTB(n137), .Q(out[96]) );
  DFFARX1_HVT \out_reg[95]  ( .D(n97), .CLK(clk), .RSTB(n137), .Q(out[95]) );
  DFFARX1_HVT \out_reg[94]  ( .D(n96), .CLK(clk), .RSTB(n137), .Q(out[94]) );
  DFFARX1_HVT \out_reg[93]  ( .D(n95), .CLK(clk), .RSTB(n137), .Q(out[93]) );
  DFFARX1_HVT \out_reg[92]  ( .D(n94), .CLK(clk), .RSTB(n137), .Q(out[92]) );
  DFFARX1_HVT \out_reg[91]  ( .D(n93), .CLK(clk), .RSTB(n137), .Q(out[91]) );
  DFFARX1_HVT \out_reg[90]  ( .D(n92), .CLK(clk), .RSTB(n137), .Q(out[90]) );
  DFFARX1_HVT \out_reg[89]  ( .D(n91), .CLK(clk), .RSTB(n137), .Q(out[89]) );
  DFFARX1_HVT \out_reg[88]  ( .D(n90), .CLK(clk), .RSTB(n137), .Q(out[88]) );
  DFFARX1_HVT \out_reg[87]  ( .D(n89), .CLK(clk), .RSTB(n137), .Q(out[87]) );
  DFFARX1_HVT \out_reg[86]  ( .D(n88), .CLK(clk), .RSTB(n136), .Q(out[86]) );
  DFFARX1_HVT \out_reg[85]  ( .D(n87), .CLK(clk), .RSTB(n136), .Q(out[85]) );
  DFFARX1_HVT \out_reg[84]  ( .D(n86), .CLK(clk), .RSTB(n136), .Q(out[84]) );
  DFFARX1_HVT \out_reg[83]  ( .D(n85), .CLK(clk), .RSTB(n136), .Q(out[83]) );
  DFFARX1_HVT \out_reg[82]  ( .D(n84), .CLK(clk), .RSTB(n136), .Q(out[82]) );
  DFFARX1_HVT \out_reg[81]  ( .D(n83), .CLK(clk), .RSTB(n136), .Q(out[81]) );
  DFFARX1_HVT \out_reg[80]  ( .D(n82), .CLK(clk), .RSTB(n136), .Q(out[80]) );
  DFFARX1_HVT \out_reg[79]  ( .D(n81), .CLK(clk), .RSTB(n136), .Q(out[79]) );
  DFFARX1_HVT \out_reg[78]  ( .D(n80), .CLK(clk), .RSTB(n136), .Q(out[78]) );
  DFFARX1_HVT \out_reg[77]  ( .D(n79), .CLK(clk), .RSTB(n136), .Q(out[77]) );
  DFFARX1_HVT \out_reg[76]  ( .D(n78), .CLK(clk), .RSTB(n136), .Q(out[76]) );
  DFFARX1_HVT \out_reg[75]  ( .D(n77), .CLK(clk), .RSTB(n135), .Q(out[75]) );
  DFFARX1_HVT \out_reg[74]  ( .D(n76), .CLK(clk), .RSTB(n135), .Q(out[74]) );
  DFFARX1_HVT \out_reg[73]  ( .D(n75), .CLK(clk), .RSTB(n135), .Q(out[73]) );
  DFFARX1_HVT \out_reg[72]  ( .D(n74), .CLK(clk), .RSTB(n135), .Q(out[72]) );
  DFFARX1_HVT \out_reg[71]  ( .D(n73), .CLK(clk), .RSTB(n135), .Q(out[71]) );
  DFFARX1_HVT \out_reg[70]  ( .D(n72), .CLK(clk), .RSTB(n135), .Q(out[70]) );
  DFFARX1_HVT \out_reg[69]  ( .D(n71), .CLK(clk), .RSTB(n135), .Q(out[69]) );
  DFFARX1_HVT \out_reg[68]  ( .D(n70), .CLK(clk), .RSTB(n135), .Q(out[68]) );
  DFFARX1_HVT \out_reg[67]  ( .D(n69), .CLK(clk), .RSTB(n135), .Q(out[67]) );
  DFFARX1_HVT \out_reg[66]  ( .D(n68), .CLK(clk), .RSTB(n135), .Q(out[66]) );
  DFFARX1_HVT \out_reg[65]  ( .D(n67), .CLK(clk), .RSTB(n135), .Q(out[65]) );
  DFFARX1_HVT \out_reg[64]  ( .D(n66), .CLK(clk), .RSTB(n134), .Q(out[64]) );
  DFFARX1_HVT \out_reg[63]  ( .D(n65), .CLK(clk), .RSTB(n134), .Q(out[63]) );
  DFFARX1_HVT \out_reg[62]  ( .D(n64), .CLK(clk), .RSTB(n134), .Q(out[62]) );
  DFFARX1_HVT \out_reg[61]  ( .D(n63), .CLK(clk), .RSTB(n134), .Q(out[61]) );
  DFFARX1_HVT \out_reg[60]  ( .D(n62), .CLK(clk), .RSTB(n134), .Q(out[60]) );
  DFFARX1_HVT \out_reg[59]  ( .D(n61), .CLK(clk), .RSTB(n134), .Q(out[59]) );
  DFFARX1_HVT \out_reg[58]  ( .D(n60), .CLK(clk), .RSTB(n134), .Q(out[58]) );
  DFFARX1_HVT \out_reg[57]  ( .D(n59), .CLK(clk), .RSTB(n134), .Q(out[57]) );
  DFFARX1_HVT \out_reg[56]  ( .D(n58), .CLK(clk), .RSTB(n134), .Q(out[56]) );
  DFFARX1_HVT \out_reg[55]  ( .D(n57), .CLK(clk), .RSTB(n134), .Q(out[55]) );
  DFFARX1_HVT \out_reg[54]  ( .D(n56), .CLK(clk), .RSTB(n134), .Q(out[54]) );
  DFFARX1_HVT \out_reg[53]  ( .D(n55), .CLK(clk), .RSTB(n133), .Q(out[53]) );
  DFFARX1_HVT \out_reg[52]  ( .D(n54), .CLK(clk), .RSTB(n133), .Q(out[52]) );
  DFFARX1_HVT \out_reg[51]  ( .D(n53), .CLK(clk), .RSTB(n133), .Q(out[51]) );
  DFFARX1_HVT \out_reg[50]  ( .D(n52), .CLK(clk), .RSTB(n133), .Q(out[50]) );
  DFFARX1_HVT \out_reg[49]  ( .D(n51), .CLK(clk), .RSTB(n133), .Q(out[49]) );
  DFFARX1_HVT \out_reg[48]  ( .D(n50), .CLK(clk), .RSTB(n133), .Q(out[48]) );
  DFFARX1_HVT \out_reg[47]  ( .D(n49), .CLK(clk), .RSTB(n133), .Q(out[47]) );
  DFFARX1_HVT \out_reg[46]  ( .D(n48), .CLK(clk), .RSTB(n133), .Q(out[46]) );
  DFFARX1_HVT \out_reg[45]  ( .D(n47), .CLK(clk), .RSTB(n133), .Q(out[45]) );
  DFFARX1_HVT \out_reg[44]  ( .D(n46), .CLK(clk), .RSTB(n133), .Q(out[44]) );
  DFFARX1_HVT \out_reg[43]  ( .D(n45), .CLK(clk), .RSTB(n133), .Q(out[43]) );
  DFFARX1_HVT \out_reg[42]  ( .D(n44), .CLK(clk), .RSTB(n132), .Q(out[42]) );
  DFFARX1_HVT \out_reg[41]  ( .D(n43), .CLK(clk), .RSTB(n132), .Q(out[41]) );
  DFFARX1_HVT \out_reg[40]  ( .D(n42), .CLK(clk), .RSTB(n132), .Q(out[40]) );
  DFFARX1_HVT \out_reg[39]  ( .D(n41), .CLK(clk), .RSTB(n132), .Q(out[39]) );
  DFFARX1_HVT \out_reg[38]  ( .D(n40), .CLK(clk), .RSTB(n132), .Q(out[38]) );
  DFFARX1_HVT \out_reg[37]  ( .D(n39), .CLK(clk), .RSTB(n132), .Q(out[37]) );
  DFFARX1_HVT \out_reg[36]  ( .D(n38), .CLK(clk), .RSTB(n132), .Q(out[36]) );
  DFFARX1_HVT \out_reg[35]  ( .D(n37), .CLK(clk), .RSTB(n132), .Q(out[35]) );
  DFFARX1_HVT \out_reg[34]  ( .D(n36), .CLK(clk), .RSTB(n132), .Q(out[34]) );
  DFFARX1_HVT \out_reg[33]  ( .D(n35), .CLK(clk), .RSTB(n132), .Q(out[33]) );
  DFFARX1_HVT \out_reg[32]  ( .D(n34), .CLK(clk), .RSTB(n132), .Q(out[32]) );
  DFFARX1_HVT \out_reg[31]  ( .D(n33), .CLK(clk), .RSTB(n131), .Q(out[31]) );
  DFFARX1_HVT \out_reg[30]  ( .D(n32), .CLK(clk), .RSTB(n131), .Q(out[30]) );
  DFFARX1_HVT \out_reg[29]  ( .D(n31), .CLK(clk), .RSTB(n131), .Q(out[29]) );
  DFFARX1_HVT \out_reg[28]  ( .D(n30), .CLK(clk), .RSTB(n131), .Q(out[28]) );
  DFFARX1_HVT \out_reg[27]  ( .D(n29), .CLK(clk), .RSTB(n131), .Q(out[27]) );
  DFFARX1_HVT \out_reg[26]  ( .D(n28), .CLK(clk), .RSTB(n131), .Q(out[26]) );
  DFFARX1_HVT \out_reg[25]  ( .D(n27), .CLK(clk), .RSTB(n131), .Q(out[25]) );
  DFFARX1_HVT \out_reg[24]  ( .D(n26), .CLK(clk), .RSTB(n131), .Q(out[24]) );
  DFFARX1_HVT \out_reg[23]  ( .D(n25), .CLK(clk), .RSTB(n131), .Q(out[23]) );
  DFFARX1_HVT \out_reg[22]  ( .D(n24), .CLK(clk), .RSTB(n131), .Q(out[22]) );
  DFFARX1_HVT \out_reg[21]  ( .D(n23), .CLK(clk), .RSTB(n131), .Q(out[21]) );
  DFFARX1_HVT \out_reg[20]  ( .D(n22), .CLK(clk), .RSTB(n129), .Q(out[20]) );
  DFFARX1_HVT \out_reg[19]  ( .D(n21), .CLK(clk), .RSTB(n129), .Q(out[19]) );
  DFFARX1_HVT \out_reg[18]  ( .D(n20), .CLK(clk), .RSTB(n129), .Q(out[18]) );
  DFFARX1_HVT \out_reg[17]  ( .D(n19), .CLK(clk), .RSTB(n129), .Q(out[17]) );
  DFFARX1_HVT \out_reg[16]  ( .D(n18), .CLK(clk), .RSTB(n129), .Q(out[16]) );
  DFFARX1_HVT \out_reg[15]  ( .D(n17), .CLK(clk), .RSTB(n129), .Q(out[15]) );
  DFFARX1_HVT \out_reg[14]  ( .D(n16), .CLK(clk), .RSTB(n129), .Q(out[14]) );
  DFFARX1_HVT \out_reg[13]  ( .D(n15), .CLK(clk), .RSTB(n129), .Q(out[13]) );
  DFFARX1_HVT \out_reg[12]  ( .D(n14), .CLK(clk), .RSTB(n129), .Q(out[12]) );
  DFFARX1_HVT \out_reg[11]  ( .D(n13), .CLK(clk), .RSTB(n139), .Q(out[11]) );
  DFFARX1_HVT \out_reg[10]  ( .D(n12), .CLK(clk), .RSTB(n1), .Q(out[10]) );
  DFFARX1_HVT \out_reg[9]  ( .D(n11), .CLK(clk), .RSTB(n138), .Q(out[9]) );
  DFFARX1_HVT \out_reg[8]  ( .D(n10), .CLK(clk), .RSTB(n137), .Q(out[8]) );
  DFFARX1_HVT \out_reg[7]  ( .D(n9), .CLK(clk), .RSTB(n136), .Q(out[7]) );
  DFFARX1_HVT \out_reg[6]  ( .D(n8), .CLK(clk), .RSTB(n135), .Q(out[6]) );
  DFFARX1_HVT \out_reg[5]  ( .D(n7), .CLK(clk), .RSTB(n134), .Q(out[5]) );
  DFFARX1_HVT \out_reg[4]  ( .D(n6), .CLK(clk), .RSTB(n133), .Q(out[4]) );
  DFFARX1_HVT \out_reg[3]  ( .D(n5), .CLK(clk), .RSTB(n132), .Q(out[3]) );
  DFFARX1_HVT \out_reg[2]  ( .D(n4), .CLK(clk), .RSTB(n131), .Q(out[2]) );
  DFFARX1_HVT \out_reg[1]  ( .D(n3), .CLK(clk), .RSTB(n129), .Q(out[1]) );
  DFFARX1_HVT \out_reg[0]  ( .D(n2), .CLK(clk), .RSTB(n1), .Q(out[0]) );
  NBUFFX2_HVT U2 ( .A(n139), .Y(n138) );
  NBUFFX2_HVT U3 ( .A(n139), .Y(n131) );
  NBUFFX2_HVT U4 ( .A(n139), .Y(n132) );
  NBUFFX2_HVT U5 ( .A(n139), .Y(n133) );
  NBUFFX2_HVT U6 ( .A(n139), .Y(n134) );
  NBUFFX2_HVT U7 ( .A(n139), .Y(n135) );
  NBUFFX2_HVT U8 ( .A(n139), .Y(n136) );
  NBUFFX2_HVT U9 ( .A(n139), .Y(n137) );
  NBUFFX2_HVT U10 ( .A(n139), .Y(n1) );
  NBUFFX2_HVT U11 ( .A(n139), .Y(n129) );
  INVX0_HVT U12 ( .A(rst), .Y(n139) );
  MUX21X1_HVT U13 ( .A1(out[97]), .A2(in[97]), .S0(enable), .Y(n99) );
  MUX21X1_HVT U14 ( .A1(out[96]), .A2(in[96]), .S0(enable), .Y(n98) );
  MUX21X1_HVT U15 ( .A1(out[95]), .A2(in[95]), .S0(enable), .Y(n97) );
  MUX21X1_HVT U16 ( .A1(out[94]), .A2(in[94]), .S0(enable), .Y(n96) );
  MUX21X1_HVT U17 ( .A1(out[93]), .A2(in[93]), .S0(enable), .Y(n95) );
  MUX21X1_HVT U18 ( .A1(out[92]), .A2(in[92]), .S0(enable), .Y(n94) );
  MUX21X1_HVT U19 ( .A1(out[91]), .A2(in[91]), .S0(enable), .Y(n93) );
  MUX21X1_HVT U20 ( .A1(out[90]), .A2(in[90]), .S0(enable), .Y(n92) );
  MUX21X1_HVT U21 ( .A1(out[89]), .A2(in[89]), .S0(enable), .Y(n91) );
  MUX21X1_HVT U22 ( .A1(out[88]), .A2(in[88]), .S0(enable), .Y(n90) );
  MUX21X1_HVT U23 ( .A1(out[7]), .A2(in[7]), .S0(enable), .Y(n9) );
  MUX21X1_HVT U24 ( .A1(out[87]), .A2(in[87]), .S0(enable), .Y(n89) );
  MUX21X1_HVT U25 ( .A1(out[86]), .A2(in[86]), .S0(enable), .Y(n88) );
  MUX21X1_HVT U26 ( .A1(out[85]), .A2(in[85]), .S0(enable), .Y(n87) );
  MUX21X1_HVT U27 ( .A1(out[84]), .A2(in[84]), .S0(enable), .Y(n86) );
  MUX21X1_HVT U28 ( .A1(out[83]), .A2(in[83]), .S0(enable), .Y(n85) );
  MUX21X1_HVT U29 ( .A1(out[82]), .A2(in[82]), .S0(enable), .Y(n84) );
  MUX21X1_HVT U30 ( .A1(out[81]), .A2(in[81]), .S0(enable), .Y(n83) );
  MUX21X1_HVT U31 ( .A1(out[80]), .A2(in[80]), .S0(enable), .Y(n82) );
  MUX21X1_HVT U32 ( .A1(out[79]), .A2(in[79]), .S0(enable), .Y(n81) );
  MUX21X1_HVT U33 ( .A1(out[78]), .A2(in[78]), .S0(enable), .Y(n80) );
  MUX21X1_HVT U34 ( .A1(out[6]), .A2(in[6]), .S0(enable), .Y(n8) );
  MUX21X1_HVT U35 ( .A1(out[77]), .A2(in[77]), .S0(enable), .Y(n79) );
  MUX21X1_HVT U36 ( .A1(out[76]), .A2(in[76]), .S0(enable), .Y(n78) );
  MUX21X1_HVT U37 ( .A1(out[75]), .A2(in[75]), .S0(enable), .Y(n77) );
  MUX21X1_HVT U38 ( .A1(out[74]), .A2(in[74]), .S0(enable), .Y(n76) );
  MUX21X1_HVT U39 ( .A1(out[73]), .A2(in[73]), .S0(enable), .Y(n75) );
  MUX21X1_HVT U40 ( .A1(out[72]), .A2(in[72]), .S0(enable), .Y(n74) );
  MUX21X1_HVT U41 ( .A1(out[71]), .A2(in[71]), .S0(enable), .Y(n73) );
  MUX21X1_HVT U42 ( .A1(out[70]), .A2(in[70]), .S0(enable), .Y(n72) );
  MUX21X1_HVT U43 ( .A1(out[69]), .A2(in[69]), .S0(enable), .Y(n71) );
  MUX21X1_HVT U44 ( .A1(out[68]), .A2(in[68]), .S0(enable), .Y(n70) );
  MUX21X1_HVT U45 ( .A1(out[5]), .A2(in[5]), .S0(enable), .Y(n7) );
  MUX21X1_HVT U46 ( .A1(out[67]), .A2(in[67]), .S0(enable), .Y(n69) );
  MUX21X1_HVT U47 ( .A1(out[66]), .A2(in[66]), .S0(enable), .Y(n68) );
  MUX21X1_HVT U48 ( .A1(out[65]), .A2(in[65]), .S0(enable), .Y(n67) );
  MUX21X1_HVT U49 ( .A1(out[64]), .A2(in[64]), .S0(enable), .Y(n66) );
  MUX21X1_HVT U50 ( .A1(out[63]), .A2(in[63]), .S0(enable), .Y(n65) );
  MUX21X1_HVT U51 ( .A1(out[62]), .A2(in[62]), .S0(enable), .Y(n64) );
  MUX21X1_HVT U52 ( .A1(out[61]), .A2(in[61]), .S0(enable), .Y(n63) );
  MUX21X1_HVT U53 ( .A1(out[60]), .A2(in[60]), .S0(enable), .Y(n62) );
  MUX21X1_HVT U54 ( .A1(out[59]), .A2(in[59]), .S0(enable), .Y(n61) );
  MUX21X1_HVT U55 ( .A1(out[58]), .A2(in[58]), .S0(enable), .Y(n60) );
  MUX21X1_HVT U56 ( .A1(out[4]), .A2(in[4]), .S0(enable), .Y(n6) );
  MUX21X1_HVT U57 ( .A1(out[57]), .A2(in[57]), .S0(enable), .Y(n59) );
  MUX21X1_HVT U58 ( .A1(out[56]), .A2(in[56]), .S0(enable), .Y(n58) );
  MUX21X1_HVT U59 ( .A1(out[55]), .A2(in[55]), .S0(enable), .Y(n57) );
  MUX21X1_HVT U60 ( .A1(out[54]), .A2(in[54]), .S0(enable), .Y(n56) );
  MUX21X1_HVT U61 ( .A1(out[53]), .A2(in[53]), .S0(enable), .Y(n55) );
  MUX21X1_HVT U62 ( .A1(out[52]), .A2(in[52]), .S0(enable), .Y(n54) );
  MUX21X1_HVT U63 ( .A1(out[51]), .A2(in[51]), .S0(enable), .Y(n53) );
  MUX21X1_HVT U64 ( .A1(out[50]), .A2(in[50]), .S0(enable), .Y(n52) );
  MUX21X1_HVT U65 ( .A1(out[49]), .A2(in[49]), .S0(enable), .Y(n51) );
  MUX21X1_HVT U66 ( .A1(out[48]), .A2(in[48]), .S0(enable), .Y(n50) );
  MUX21X1_HVT U67 ( .A1(out[3]), .A2(in[3]), .S0(enable), .Y(n5) );
  MUX21X1_HVT U68 ( .A1(out[47]), .A2(in[47]), .S0(enable), .Y(n49) );
  MUX21X1_HVT U69 ( .A1(out[46]), .A2(in[46]), .S0(enable), .Y(n48) );
  MUX21X1_HVT U70 ( .A1(out[45]), .A2(in[45]), .S0(enable), .Y(n47) );
  MUX21X1_HVT U71 ( .A1(out[44]), .A2(in[44]), .S0(enable), .Y(n46) );
  MUX21X1_HVT U72 ( .A1(out[43]), .A2(in[43]), .S0(enable), .Y(n45) );
  MUX21X1_HVT U73 ( .A1(out[42]), .A2(in[42]), .S0(enable), .Y(n44) );
  MUX21X1_HVT U74 ( .A1(out[41]), .A2(in[41]), .S0(enable), .Y(n43) );
  MUX21X1_HVT U75 ( .A1(out[40]), .A2(in[40]), .S0(enable), .Y(n42) );
  MUX21X1_HVT U76 ( .A1(out[39]), .A2(in[39]), .S0(enable), .Y(n41) );
  MUX21X1_HVT U77 ( .A1(out[38]), .A2(in[38]), .S0(enable), .Y(n40) );
  MUX21X1_HVT U78 ( .A1(out[2]), .A2(in[2]), .S0(enable), .Y(n4) );
  MUX21X1_HVT U79 ( .A1(out[37]), .A2(in[37]), .S0(enable), .Y(n39) );
  MUX21X1_HVT U80 ( .A1(out[36]), .A2(in[36]), .S0(enable), .Y(n38) );
  MUX21X1_HVT U81 ( .A1(out[35]), .A2(in[35]), .S0(enable), .Y(n37) );
  MUX21X1_HVT U82 ( .A1(out[34]), .A2(in[34]), .S0(enable), .Y(n36) );
  MUX21X1_HVT U83 ( .A1(out[33]), .A2(in[33]), .S0(enable), .Y(n35) );
  MUX21X1_HVT U84 ( .A1(out[32]), .A2(in[32]), .S0(enable), .Y(n34) );
  MUX21X1_HVT U85 ( .A1(out[31]), .A2(in[31]), .S0(enable), .Y(n33) );
  MUX21X1_HVT U86 ( .A1(out[30]), .A2(in[30]), .S0(enable), .Y(n32) );
  MUX21X1_HVT U87 ( .A1(out[29]), .A2(in[29]), .S0(enable), .Y(n31) );
  MUX21X1_HVT U88 ( .A1(out[28]), .A2(in[28]), .S0(enable), .Y(n30) );
  MUX21X1_HVT U89 ( .A1(out[1]), .A2(in[1]), .S0(enable), .Y(n3) );
  MUX21X1_HVT U90 ( .A1(out[27]), .A2(in[27]), .S0(enable), .Y(n29) );
  MUX21X1_HVT U91 ( .A1(out[26]), .A2(in[26]), .S0(enable), .Y(n28) );
  MUX21X1_HVT U92 ( .A1(out[25]), .A2(in[25]), .S0(enable), .Y(n27) );
  MUX21X1_HVT U93 ( .A1(out[24]), .A2(in[24]), .S0(enable), .Y(n26) );
  MUX21X1_HVT U94 ( .A1(out[23]), .A2(in[23]), .S0(enable), .Y(n25) );
  MUX21X1_HVT U95 ( .A1(out[22]), .A2(in[22]), .S0(enable), .Y(n24) );
  MUX21X1_HVT U96 ( .A1(out[21]), .A2(in[21]), .S0(enable), .Y(n23) );
  MUX21X1_HVT U97 ( .A1(out[20]), .A2(in[20]), .S0(enable), .Y(n22) );
  MUX21X1_HVT U98 ( .A1(out[19]), .A2(in[19]), .S0(enable), .Y(n21) );
  MUX21X1_HVT U99 ( .A1(out[18]), .A2(in[18]), .S0(enable), .Y(n20) );
  MUX21X1_HVT U100 ( .A1(out[0]), .A2(in[0]), .S0(enable), .Y(n2) );
  MUX21X1_HVT U101 ( .A1(out[17]), .A2(in[17]), .S0(enable), .Y(n19) );
  MUX21X1_HVT U102 ( .A1(out[16]), .A2(in[16]), .S0(enable), .Y(n18) );
  MUX21X1_HVT U103 ( .A1(out[15]), .A2(in[15]), .S0(enable), .Y(n17) );
  MUX21X1_HVT U104 ( .A1(out[14]), .A2(in[14]), .S0(enable), .Y(n16) );
  MUX21X1_HVT U105 ( .A1(out[13]), .A2(in[13]), .S0(enable), .Y(n15) );
  MUX21X1_HVT U106 ( .A1(out[12]), .A2(in[12]), .S0(enable), .Y(n14) );
  MUX21X1_HVT U107 ( .A1(out[127]), .A2(in[127]), .S0(enable), .Y(n130) );
  MUX21X1_HVT U108 ( .A1(out[11]), .A2(in[11]), .S0(enable), .Y(n13) );
  MUX21X1_HVT U109 ( .A1(out[126]), .A2(in[126]), .S0(enable), .Y(n128) );
  MUX21X1_HVT U110 ( .A1(out[125]), .A2(in[125]), .S0(enable), .Y(n127) );
  MUX21X1_HVT U111 ( .A1(out[124]), .A2(in[124]), .S0(enable), .Y(n126) );
  MUX21X1_HVT U112 ( .A1(out[123]), .A2(in[123]), .S0(enable), .Y(n125) );
  MUX21X1_HVT U113 ( .A1(out[122]), .A2(in[122]), .S0(enable), .Y(n124) );
  MUX21X1_HVT U114 ( .A1(out[121]), .A2(in[121]), .S0(enable), .Y(n123) );
  MUX21X1_HVT U115 ( .A1(out[120]), .A2(in[120]), .S0(enable), .Y(n122) );
  MUX21X1_HVT U116 ( .A1(out[119]), .A2(in[119]), .S0(enable), .Y(n121) );
  MUX21X1_HVT U117 ( .A1(out[118]), .A2(in[118]), .S0(enable), .Y(n120) );
  MUX21X1_HVT U118 ( .A1(out[10]), .A2(in[10]), .S0(enable), .Y(n12) );
  MUX21X1_HVT U119 ( .A1(out[117]), .A2(in[117]), .S0(enable), .Y(n119) );
  MUX21X1_HVT U120 ( .A1(out[116]), .A2(in[116]), .S0(enable), .Y(n118) );
  MUX21X1_HVT U121 ( .A1(out[115]), .A2(in[115]), .S0(enable), .Y(n117) );
  MUX21X1_HVT U122 ( .A1(out[114]), .A2(in[114]), .S0(enable), .Y(n116) );
  MUX21X1_HVT U123 ( .A1(out[113]), .A2(in[113]), .S0(enable), .Y(n115) );
  MUX21X1_HVT U124 ( .A1(out[112]), .A2(in[112]), .S0(enable), .Y(n114) );
  MUX21X1_HVT U125 ( .A1(out[111]), .A2(in[111]), .S0(enable), .Y(n113) );
  MUX21X1_HVT U126 ( .A1(out[110]), .A2(in[110]), .S0(enable), .Y(n112) );
  MUX21X1_HVT U127 ( .A1(out[109]), .A2(in[109]), .S0(enable), .Y(n111) );
  MUX21X1_HVT U128 ( .A1(out[108]), .A2(in[108]), .S0(enable), .Y(n110) );
  MUX21X1_HVT U129 ( .A1(out[9]), .A2(in[9]), .S0(enable), .Y(n11) );
  MUX21X1_HVT U130 ( .A1(out[107]), .A2(in[107]), .S0(enable), .Y(n109) );
  MUX21X1_HVT U131 ( .A1(out[106]), .A2(in[106]), .S0(enable), .Y(n108) );
  MUX21X1_HVT U132 ( .A1(out[105]), .A2(in[105]), .S0(enable), .Y(n107) );
  MUX21X1_HVT U133 ( .A1(out[104]), .A2(in[104]), .S0(enable), .Y(n106) );
  MUX21X1_HVT U134 ( .A1(out[103]), .A2(in[103]), .S0(enable), .Y(n105) );
  MUX21X1_HVT U135 ( .A1(out[102]), .A2(in[102]), .S0(enable), .Y(n104) );
  MUX21X1_HVT U136 ( .A1(out[101]), .A2(in[101]), .S0(enable), .Y(n103) );
  MUX21X1_HVT U137 ( .A1(out[100]), .A2(in[100]), .S0(enable), .Y(n102) );
  MUX21X1_HVT U138 ( .A1(out[99]), .A2(in[99]), .S0(enable), .Y(n101) );
  MUX21X1_HVT U139 ( .A1(out[98]), .A2(in[98]), .S0(enable), .Y(n100) );
  MUX21X1_HVT U140 ( .A1(out[8]), .A2(in[8]), .S0(enable), .Y(n10) );
endmodule

