
module RAM_memory ( data, addr, we, clk, rst, q );
  input [255:0] data;
  input [3:0] addr;
  output [255:0] q;
  input we, clk, rst;
  wire   N26, N27, N28, N29, \ram[15][255] , \ram[15][254] , \ram[15][253] ,
         \ram[15][252] , \ram[15][251] , \ram[15][250] , \ram[15][249] ,
         \ram[15][248] , \ram[15][247] , \ram[15][246] , \ram[15][245] ,
         \ram[15][244] , \ram[15][243] , \ram[15][242] , \ram[15][241] ,
         \ram[15][240] , \ram[15][239] , \ram[15][238] , \ram[15][237] ,
         \ram[15][236] , \ram[15][235] , \ram[15][234] , \ram[15][233] ,
         \ram[15][232] , \ram[15][231] , \ram[15][230] , \ram[15][229] ,
         \ram[15][228] , \ram[15][227] , \ram[15][226] , \ram[15][225] ,
         \ram[15][224] , \ram[15][223] , \ram[15][222] , \ram[15][221] ,
         \ram[15][220] , \ram[15][219] , \ram[15][218] , \ram[15][217] ,
         \ram[15][216] , \ram[15][215] , \ram[15][214] , \ram[15][213] ,
         \ram[15][212] , \ram[15][211] , \ram[15][210] , \ram[15][209] ,
         \ram[15][208] , \ram[15][207] , \ram[15][206] , \ram[15][205] ,
         \ram[15][204] , \ram[15][203] , \ram[15][202] , \ram[15][201] ,
         \ram[15][200] , \ram[15][199] , \ram[15][198] , \ram[15][197] ,
         \ram[15][196] , \ram[15][195] , \ram[15][194] , \ram[15][193] ,
         \ram[15][192] , \ram[15][191] , \ram[15][190] , \ram[15][189] ,
         \ram[15][188] , \ram[15][187] , \ram[15][186] , \ram[15][185] ,
         \ram[15][184] , \ram[15][183] , \ram[15][182] , \ram[15][181] ,
         \ram[15][180] , \ram[15][179] , \ram[15][178] , \ram[15][177] ,
         \ram[15][176] , \ram[15][175] , \ram[15][174] , \ram[15][173] ,
         \ram[15][172] , \ram[15][171] , \ram[15][170] , \ram[15][169] ,
         \ram[15][168] , \ram[15][167] , \ram[15][166] , \ram[15][165] ,
         \ram[15][164] , \ram[15][163] , \ram[15][162] , \ram[15][161] ,
         \ram[15][160] , \ram[15][159] , \ram[15][158] , \ram[15][157] ,
         \ram[15][156] , \ram[15][155] , \ram[15][154] , \ram[15][153] ,
         \ram[15][152] , \ram[15][151] , \ram[15][150] , \ram[15][149] ,
         \ram[15][148] , \ram[15][147] , \ram[15][146] , \ram[15][145] ,
         \ram[15][144] , \ram[15][143] , \ram[15][142] , \ram[15][141] ,
         \ram[15][140] , \ram[15][139] , \ram[15][138] , \ram[15][137] ,
         \ram[15][136] , \ram[15][135] , \ram[15][134] , \ram[15][133] ,
         \ram[15][132] , \ram[15][131] , \ram[15][130] , \ram[15][129] ,
         \ram[15][128] , \ram[15][127] , \ram[15][126] , \ram[15][125] ,
         \ram[15][124] , \ram[15][123] , \ram[15][122] , \ram[15][121] ,
         \ram[15][120] , \ram[15][119] , \ram[15][118] , \ram[15][117] ,
         \ram[15][116] , \ram[15][115] , \ram[15][114] , \ram[15][113] ,
         \ram[15][112] , \ram[15][111] , \ram[15][110] , \ram[15][109] ,
         \ram[15][108] , \ram[15][107] , \ram[15][106] , \ram[15][105] ,
         \ram[15][104] , \ram[15][103] , \ram[15][102] , \ram[15][101] ,
         \ram[15][100] , \ram[15][99] , \ram[15][98] , \ram[15][97] ,
         \ram[15][96] , \ram[15][95] , \ram[15][94] , \ram[15][93] ,
         \ram[15][92] , \ram[15][91] , \ram[15][90] , \ram[15][89] ,
         \ram[15][88] , \ram[15][87] , \ram[15][86] , \ram[15][85] ,
         \ram[15][84] , \ram[15][83] , \ram[15][82] , \ram[15][81] ,
         \ram[15][80] , \ram[15][79] , \ram[15][78] , \ram[15][77] ,
         \ram[15][76] , \ram[15][75] , \ram[15][74] , \ram[15][73] ,
         \ram[15][72] , \ram[15][71] , \ram[15][70] , \ram[15][69] ,
         \ram[15][68] , \ram[15][67] , \ram[15][66] , \ram[15][65] ,
         \ram[15][64] , \ram[15][63] , \ram[15][62] , \ram[15][61] ,
         \ram[15][60] , \ram[15][59] , \ram[15][58] , \ram[15][57] ,
         \ram[15][56] , \ram[15][55] , \ram[15][54] , \ram[15][53] ,
         \ram[15][52] , \ram[15][51] , \ram[15][50] , \ram[15][49] ,
         \ram[15][48] , \ram[15][47] , \ram[15][46] , \ram[15][45] ,
         \ram[15][44] , \ram[15][43] , \ram[15][42] , \ram[15][41] ,
         \ram[15][40] , \ram[15][39] , \ram[15][38] , \ram[15][37] ,
         \ram[15][36] , \ram[15][35] , \ram[15][34] , \ram[15][33] ,
         \ram[15][32] , \ram[15][31] , \ram[15][30] , \ram[15][29] ,
         \ram[15][28] , \ram[15][27] , \ram[15][26] , \ram[15][25] ,
         \ram[15][24] , \ram[15][23] , \ram[15][22] , \ram[15][21] ,
         \ram[15][20] , \ram[15][19] , \ram[15][18] , \ram[15][17] ,
         \ram[15][16] , \ram[15][15] , \ram[15][14] , \ram[15][13] ,
         \ram[15][12] , \ram[15][11] , \ram[15][10] , \ram[15][9] ,
         \ram[15][8] , \ram[15][7] , \ram[15][6] , \ram[15][5] , \ram[15][4] ,
         \ram[15][3] , \ram[15][2] , \ram[15][1] , \ram[15][0] ,
         \ram[14][255] , \ram[14][254] , \ram[14][253] , \ram[14][252] ,
         \ram[14][251] , \ram[14][250] , \ram[14][249] , \ram[14][248] ,
         \ram[14][247] , \ram[14][246] , \ram[14][245] , \ram[14][244] ,
         \ram[14][243] , \ram[14][242] , \ram[14][241] , \ram[14][240] ,
         \ram[14][239] , \ram[14][238] , \ram[14][237] , \ram[14][236] ,
         \ram[14][235] , \ram[14][234] , \ram[14][233] , \ram[14][232] ,
         \ram[14][231] , \ram[14][230] , \ram[14][229] , \ram[14][228] ,
         \ram[14][227] , \ram[14][226] , \ram[14][225] , \ram[14][224] ,
         \ram[14][223] , \ram[14][222] , \ram[14][221] , \ram[14][220] ,
         \ram[14][219] , \ram[14][218] , \ram[14][217] , \ram[14][216] ,
         \ram[14][215] , \ram[14][214] , \ram[14][213] , \ram[14][212] ,
         \ram[14][211] , \ram[14][210] , \ram[14][209] , \ram[14][208] ,
         \ram[14][207] , \ram[14][206] , \ram[14][205] , \ram[14][204] ,
         \ram[14][203] , \ram[14][202] , \ram[14][201] , \ram[14][200] ,
         \ram[14][199] , \ram[14][198] , \ram[14][197] , \ram[14][196] ,
         \ram[14][195] , \ram[14][194] , \ram[14][193] , \ram[14][192] ,
         \ram[14][191] , \ram[14][190] , \ram[14][189] , \ram[14][188] ,
         \ram[14][187] , \ram[14][186] , \ram[14][185] , \ram[14][184] ,
         \ram[14][183] , \ram[14][182] , \ram[14][181] , \ram[14][180] ,
         \ram[14][179] , \ram[14][178] , \ram[14][177] , \ram[14][176] ,
         \ram[14][175] , \ram[14][174] , \ram[14][173] , \ram[14][172] ,
         \ram[14][171] , \ram[14][170] , \ram[14][169] , \ram[14][168] ,
         \ram[14][167] , \ram[14][166] , \ram[14][165] , \ram[14][164] ,
         \ram[14][163] , \ram[14][162] , \ram[14][161] , \ram[14][160] ,
         \ram[14][159] , \ram[14][158] , \ram[14][157] , \ram[14][156] ,
         \ram[14][155] , \ram[14][154] , \ram[14][153] , \ram[14][152] ,
         \ram[14][151] , \ram[14][150] , \ram[14][149] , \ram[14][148] ,
         \ram[14][147] , \ram[14][146] , \ram[14][145] , \ram[14][144] ,
         \ram[14][143] , \ram[14][142] , \ram[14][141] , \ram[14][140] ,
         \ram[14][139] , \ram[14][138] , \ram[14][137] , \ram[14][136] ,
         \ram[14][135] , \ram[14][134] , \ram[14][133] , \ram[14][132] ,
         \ram[14][131] , \ram[14][130] , \ram[14][129] , \ram[14][128] ,
         \ram[14][127] , \ram[14][126] , \ram[14][125] , \ram[14][124] ,
         \ram[14][123] , \ram[14][122] , \ram[14][121] , \ram[14][120] ,
         \ram[14][119] , \ram[14][118] , \ram[14][117] , \ram[14][116] ,
         \ram[14][115] , \ram[14][114] , \ram[14][113] , \ram[14][112] ,
         \ram[14][111] , \ram[14][110] , \ram[14][109] , \ram[14][108] ,
         \ram[14][107] , \ram[14][106] , \ram[14][105] , \ram[14][104] ,
         \ram[14][103] , \ram[14][102] , \ram[14][101] , \ram[14][100] ,
         \ram[14][99] , \ram[14][98] , \ram[14][97] , \ram[14][96] ,
         \ram[14][95] , \ram[14][94] , \ram[14][93] , \ram[14][92] ,
         \ram[14][91] , \ram[14][90] , \ram[14][89] , \ram[14][88] ,
         \ram[14][87] , \ram[14][86] , \ram[14][85] , \ram[14][84] ,
         \ram[14][83] , \ram[14][82] , \ram[14][81] , \ram[14][80] ,
         \ram[14][79] , \ram[14][78] , \ram[14][77] , \ram[14][76] ,
         \ram[14][75] , \ram[14][74] , \ram[14][73] , \ram[14][72] ,
         \ram[14][71] , \ram[14][70] , \ram[14][69] , \ram[14][68] ,
         \ram[14][67] , \ram[14][66] , \ram[14][65] , \ram[14][64] ,
         \ram[14][63] , \ram[14][62] , \ram[14][61] , \ram[14][60] ,
         \ram[14][59] , \ram[14][58] , \ram[14][57] , \ram[14][56] ,
         \ram[14][55] , \ram[14][54] , \ram[14][53] , \ram[14][52] ,
         \ram[14][51] , \ram[14][50] , \ram[14][49] , \ram[14][48] ,
         \ram[14][47] , \ram[14][46] , \ram[14][45] , \ram[14][44] ,
         \ram[14][43] , \ram[14][42] , \ram[14][41] , \ram[14][40] ,
         \ram[14][39] , \ram[14][38] , \ram[14][37] , \ram[14][36] ,
         \ram[14][35] , \ram[14][34] , \ram[14][33] , \ram[14][32] ,
         \ram[14][31] , \ram[14][30] , \ram[14][29] , \ram[14][28] ,
         \ram[14][27] , \ram[14][26] , \ram[14][25] , \ram[14][24] ,
         \ram[14][23] , \ram[14][22] , \ram[14][21] , \ram[14][20] ,
         \ram[14][19] , \ram[14][18] , \ram[14][17] , \ram[14][16] ,
         \ram[14][15] , \ram[14][14] , \ram[14][13] , \ram[14][12] ,
         \ram[14][11] , \ram[14][10] , \ram[14][9] , \ram[14][8] ,
         \ram[14][7] , \ram[14][6] , \ram[14][5] , \ram[14][4] , \ram[14][3] ,
         \ram[14][2] , \ram[14][1] , \ram[14][0] , \ram[13][255] ,
         \ram[13][254] , \ram[13][253] , \ram[13][252] , \ram[13][251] ,
         \ram[13][250] , \ram[13][249] , \ram[13][248] , \ram[13][247] ,
         \ram[13][246] , \ram[13][245] , \ram[13][244] , \ram[13][243] ,
         \ram[13][242] , \ram[13][241] , \ram[13][240] , \ram[13][239] ,
         \ram[13][238] , \ram[13][237] , \ram[13][236] , \ram[13][235] ,
         \ram[13][234] , \ram[13][233] , \ram[13][232] , \ram[13][231] ,
         \ram[13][230] , \ram[13][229] , \ram[13][228] , \ram[13][227] ,
         \ram[13][226] , \ram[13][225] , \ram[13][224] , \ram[13][223] ,
         \ram[13][222] , \ram[13][221] , \ram[13][220] , \ram[13][219] ,
         \ram[13][218] , \ram[13][217] , \ram[13][216] , \ram[13][215] ,
         \ram[13][214] , \ram[13][213] , \ram[13][212] , \ram[13][211] ,
         \ram[13][210] , \ram[13][209] , \ram[13][208] , \ram[13][207] ,
         \ram[13][206] , \ram[13][205] , \ram[13][204] , \ram[13][203] ,
         \ram[13][202] , \ram[13][201] , \ram[13][200] , \ram[13][199] ,
         \ram[13][198] , \ram[13][197] , \ram[13][196] , \ram[13][195] ,
         \ram[13][194] , \ram[13][193] , \ram[13][192] , \ram[13][191] ,
         \ram[13][190] , \ram[13][189] , \ram[13][188] , \ram[13][187] ,
         \ram[13][186] , \ram[13][185] , \ram[13][184] , \ram[13][183] ,
         \ram[13][182] , \ram[13][181] , \ram[13][180] , \ram[13][179] ,
         \ram[13][178] , \ram[13][177] , \ram[13][176] , \ram[13][175] ,
         \ram[13][174] , \ram[13][173] , \ram[13][172] , \ram[13][171] ,
         \ram[13][170] , \ram[13][169] , \ram[13][168] , \ram[13][167] ,
         \ram[13][166] , \ram[13][165] , \ram[13][164] , \ram[13][163] ,
         \ram[13][162] , \ram[13][161] , \ram[13][160] , \ram[13][159] ,
         \ram[13][158] , \ram[13][157] , \ram[13][156] , \ram[13][155] ,
         \ram[13][154] , \ram[13][153] , \ram[13][152] , \ram[13][151] ,
         \ram[13][150] , \ram[13][149] , \ram[13][148] , \ram[13][147] ,
         \ram[13][146] , \ram[13][145] , \ram[13][144] , \ram[13][143] ,
         \ram[13][142] , \ram[13][141] , \ram[13][140] , \ram[13][139] ,
         \ram[13][138] , \ram[13][137] , \ram[13][136] , \ram[13][135] ,
         \ram[13][134] , \ram[13][133] , \ram[13][132] , \ram[13][131] ,
         \ram[13][130] , \ram[13][129] , \ram[13][128] , \ram[13][127] ,
         \ram[13][126] , \ram[13][125] , \ram[13][124] , \ram[13][123] ,
         \ram[13][122] , \ram[13][121] , \ram[13][120] , \ram[13][119] ,
         \ram[13][118] , \ram[13][117] , \ram[13][116] , \ram[13][115] ,
         \ram[13][114] , \ram[13][113] , \ram[13][112] , \ram[13][111] ,
         \ram[13][110] , \ram[13][109] , \ram[13][108] , \ram[13][107] ,
         \ram[13][106] , \ram[13][105] , \ram[13][104] , \ram[13][103] ,
         \ram[13][102] , \ram[13][101] , \ram[13][100] , \ram[13][99] ,
         \ram[13][98] , \ram[13][97] , \ram[13][96] , \ram[13][95] ,
         \ram[13][94] , \ram[13][93] , \ram[13][92] , \ram[13][91] ,
         \ram[13][90] , \ram[13][89] , \ram[13][88] , \ram[13][87] ,
         \ram[13][86] , \ram[13][85] , \ram[13][84] , \ram[13][83] ,
         \ram[13][82] , \ram[13][81] , \ram[13][80] , \ram[13][79] ,
         \ram[13][78] , \ram[13][77] , \ram[13][76] , \ram[13][75] ,
         \ram[13][74] , \ram[13][73] , \ram[13][72] , \ram[13][71] ,
         \ram[13][70] , \ram[13][69] , \ram[13][68] , \ram[13][67] ,
         \ram[13][66] , \ram[13][65] , \ram[13][64] , \ram[13][63] ,
         \ram[13][62] , \ram[13][61] , \ram[13][60] , \ram[13][59] ,
         \ram[13][58] , \ram[13][57] , \ram[13][56] , \ram[13][55] ,
         \ram[13][54] , \ram[13][53] , \ram[13][52] , \ram[13][51] ,
         \ram[13][50] , \ram[13][49] , \ram[13][48] , \ram[13][47] ,
         \ram[13][46] , \ram[13][45] , \ram[13][44] , \ram[13][43] ,
         \ram[13][42] , \ram[13][41] , \ram[13][40] , \ram[13][39] ,
         \ram[13][38] , \ram[13][37] , \ram[13][36] , \ram[13][35] ,
         \ram[13][34] , \ram[13][33] , \ram[13][32] , \ram[13][31] ,
         \ram[13][30] , \ram[13][29] , \ram[13][28] , \ram[13][27] ,
         \ram[13][26] , \ram[13][25] , \ram[13][24] , \ram[13][23] ,
         \ram[13][22] , \ram[13][21] , \ram[13][20] , \ram[13][19] ,
         \ram[13][18] , \ram[13][17] , \ram[13][16] , \ram[13][15] ,
         \ram[13][14] , \ram[13][13] , \ram[13][12] , \ram[13][11] ,
         \ram[13][10] , \ram[13][9] , \ram[13][8] , \ram[13][7] , \ram[13][6] ,
         \ram[13][5] , \ram[13][4] , \ram[13][3] , \ram[13][2] , \ram[13][1] ,
         \ram[13][0] , \ram[12][255] , \ram[12][254] , \ram[12][253] ,
         \ram[12][252] , \ram[12][251] , \ram[12][250] , \ram[12][249] ,
         \ram[12][248] , \ram[12][247] , \ram[12][246] , \ram[12][245] ,
         \ram[12][244] , \ram[12][243] , \ram[12][242] , \ram[12][241] ,
         \ram[12][240] , \ram[12][239] , \ram[12][238] , \ram[12][237] ,
         \ram[12][236] , \ram[12][235] , \ram[12][234] , \ram[12][233] ,
         \ram[12][232] , \ram[12][231] , \ram[12][230] , \ram[12][229] ,
         \ram[12][228] , \ram[12][227] , \ram[12][226] , \ram[12][225] ,
         \ram[12][224] , \ram[12][223] , \ram[12][222] , \ram[12][221] ,
         \ram[12][220] , \ram[12][219] , \ram[12][218] , \ram[12][217] ,
         \ram[12][216] , \ram[12][215] , \ram[12][214] , \ram[12][213] ,
         \ram[12][212] , \ram[12][211] , \ram[12][210] , \ram[12][209] ,
         \ram[12][208] , \ram[12][207] , \ram[12][206] , \ram[12][205] ,
         \ram[12][204] , \ram[12][203] , \ram[12][202] , \ram[12][201] ,
         \ram[12][200] , \ram[12][199] , \ram[12][198] , \ram[12][197] ,
         \ram[12][196] , \ram[12][195] , \ram[12][194] , \ram[12][193] ,
         \ram[12][192] , \ram[12][191] , \ram[12][190] , \ram[12][189] ,
         \ram[12][188] , \ram[12][187] , \ram[12][186] , \ram[12][185] ,
         \ram[12][184] , \ram[12][183] , \ram[12][182] , \ram[12][181] ,
         \ram[12][180] , \ram[12][179] , \ram[12][178] , \ram[12][177] ,
         \ram[12][176] , \ram[12][175] , \ram[12][174] , \ram[12][173] ,
         \ram[12][172] , \ram[12][171] , \ram[12][170] , \ram[12][169] ,
         \ram[12][168] , \ram[12][167] , \ram[12][166] , \ram[12][165] ,
         \ram[12][164] , \ram[12][163] , \ram[12][162] , \ram[12][161] ,
         \ram[12][160] , \ram[12][159] , \ram[12][158] , \ram[12][157] ,
         \ram[12][156] , \ram[12][155] , \ram[12][154] , \ram[12][153] ,
         \ram[12][152] , \ram[12][151] , \ram[12][150] , \ram[12][149] ,
         \ram[12][148] , \ram[12][147] , \ram[12][146] , \ram[12][145] ,
         \ram[12][144] , \ram[12][143] , \ram[12][142] , \ram[12][141] ,
         \ram[12][140] , \ram[12][139] , \ram[12][138] , \ram[12][137] ,
         \ram[12][136] , \ram[12][135] , \ram[12][134] , \ram[12][133] ,
         \ram[12][132] , \ram[12][131] , \ram[12][130] , \ram[12][129] ,
         \ram[12][128] , \ram[12][127] , \ram[12][126] , \ram[12][125] ,
         \ram[12][124] , \ram[12][123] , \ram[12][122] , \ram[12][121] ,
         \ram[12][120] , \ram[12][119] , \ram[12][118] , \ram[12][117] ,
         \ram[12][116] , \ram[12][115] , \ram[12][114] , \ram[12][113] ,
         \ram[12][112] , \ram[12][111] , \ram[12][110] , \ram[12][109] ,
         \ram[12][108] , \ram[12][107] , \ram[12][106] , \ram[12][105] ,
         \ram[12][104] , \ram[12][103] , \ram[12][102] , \ram[12][101] ,
         \ram[12][100] , \ram[12][99] , \ram[12][98] , \ram[12][97] ,
         \ram[12][96] , \ram[12][95] , \ram[12][94] , \ram[12][93] ,
         \ram[12][92] , \ram[12][91] , \ram[12][90] , \ram[12][89] ,
         \ram[12][88] , \ram[12][87] , \ram[12][86] , \ram[12][85] ,
         \ram[12][84] , \ram[12][83] , \ram[12][82] , \ram[12][81] ,
         \ram[12][80] , \ram[12][79] , \ram[12][78] , \ram[12][77] ,
         \ram[12][76] , \ram[12][75] , \ram[12][74] , \ram[12][73] ,
         \ram[12][72] , \ram[12][71] , \ram[12][70] , \ram[12][69] ,
         \ram[12][68] , \ram[12][67] , \ram[12][66] , \ram[12][65] ,
         \ram[12][64] , \ram[12][63] , \ram[12][62] , \ram[12][61] ,
         \ram[12][60] , \ram[12][59] , \ram[12][58] , \ram[12][57] ,
         \ram[12][56] , \ram[12][55] , \ram[12][54] , \ram[12][53] ,
         \ram[12][52] , \ram[12][51] , \ram[12][50] , \ram[12][49] ,
         \ram[12][48] , \ram[12][47] , \ram[12][46] , \ram[12][45] ,
         \ram[12][44] , \ram[12][43] , \ram[12][42] , \ram[12][41] ,
         \ram[12][40] , \ram[12][39] , \ram[12][38] , \ram[12][37] ,
         \ram[12][36] , \ram[12][35] , \ram[12][34] , \ram[12][33] ,
         \ram[12][32] , \ram[12][31] , \ram[12][30] , \ram[12][29] ,
         \ram[12][28] , \ram[12][27] , \ram[12][26] , \ram[12][25] ,
         \ram[12][24] , \ram[12][23] , \ram[12][22] , \ram[12][21] ,
         \ram[12][20] , \ram[12][19] , \ram[12][18] , \ram[12][17] ,
         \ram[12][16] , \ram[12][15] , \ram[12][14] , \ram[12][13] ,
         \ram[12][12] , \ram[12][11] , \ram[12][10] , \ram[12][9] ,
         \ram[12][8] , \ram[12][7] , \ram[12][6] , \ram[12][5] , \ram[12][4] ,
         \ram[12][3] , \ram[12][2] , \ram[12][1] , \ram[12][0] ,
         \ram[11][255] , \ram[11][254] , \ram[11][253] , \ram[11][252] ,
         \ram[11][251] , \ram[11][250] , \ram[11][249] , \ram[11][248] ,
         \ram[11][247] , \ram[11][246] , \ram[11][245] , \ram[11][244] ,
         \ram[11][243] , \ram[11][242] , \ram[11][241] , \ram[11][240] ,
         \ram[11][239] , \ram[11][238] , \ram[11][237] , \ram[11][236] ,
         \ram[11][235] , \ram[11][234] , \ram[11][233] , \ram[11][232] ,
         \ram[11][231] , \ram[11][230] , \ram[11][229] , \ram[11][228] ,
         \ram[11][227] , \ram[11][226] , \ram[11][225] , \ram[11][224] ,
         \ram[11][223] , \ram[11][222] , \ram[11][221] , \ram[11][220] ,
         \ram[11][219] , \ram[11][218] , \ram[11][217] , \ram[11][216] ,
         \ram[11][215] , \ram[11][214] , \ram[11][213] , \ram[11][212] ,
         \ram[11][211] , \ram[11][210] , \ram[11][209] , \ram[11][208] ,
         \ram[11][207] , \ram[11][206] , \ram[11][205] , \ram[11][204] ,
         \ram[11][203] , \ram[11][202] , \ram[11][201] , \ram[11][200] ,
         \ram[11][199] , \ram[11][198] , \ram[11][197] , \ram[11][196] ,
         \ram[11][195] , \ram[11][194] , \ram[11][193] , \ram[11][192] ,
         \ram[11][191] , \ram[11][190] , \ram[11][189] , \ram[11][188] ,
         \ram[11][187] , \ram[11][186] , \ram[11][185] , \ram[11][184] ,
         \ram[11][183] , \ram[11][182] , \ram[11][181] , \ram[11][180] ,
         \ram[11][179] , \ram[11][178] , \ram[11][177] , \ram[11][176] ,
         \ram[11][175] , \ram[11][174] , \ram[11][173] , \ram[11][172] ,
         \ram[11][171] , \ram[11][170] , \ram[11][169] , \ram[11][168] ,
         \ram[11][167] , \ram[11][166] , \ram[11][165] , \ram[11][164] ,
         \ram[11][163] , \ram[11][162] , \ram[11][161] , \ram[11][160] ,
         \ram[11][159] , \ram[11][158] , \ram[11][157] , \ram[11][156] ,
         \ram[11][155] , \ram[11][154] , \ram[11][153] , \ram[11][152] ,
         \ram[11][151] , \ram[11][150] , \ram[11][149] , \ram[11][148] ,
         \ram[11][147] , \ram[11][146] , \ram[11][145] , \ram[11][144] ,
         \ram[11][143] , \ram[11][142] , \ram[11][141] , \ram[11][140] ,
         \ram[11][139] , \ram[11][138] , \ram[11][137] , \ram[11][136] ,
         \ram[11][135] , \ram[11][134] , \ram[11][133] , \ram[11][132] ,
         \ram[11][131] , \ram[11][130] , \ram[11][129] , \ram[11][128] ,
         \ram[11][127] , \ram[11][126] , \ram[11][125] , \ram[11][124] ,
         \ram[11][123] , \ram[11][122] , \ram[11][121] , \ram[11][120] ,
         \ram[11][119] , \ram[11][118] , \ram[11][117] , \ram[11][116] ,
         \ram[11][115] , \ram[11][114] , \ram[11][113] , \ram[11][112] ,
         \ram[11][111] , \ram[11][110] , \ram[11][109] , \ram[11][108] ,
         \ram[11][107] , \ram[11][106] , \ram[11][105] , \ram[11][104] ,
         \ram[11][103] , \ram[11][102] , \ram[11][101] , \ram[11][100] ,
         \ram[11][99] , \ram[11][98] , \ram[11][97] , \ram[11][96] ,
         \ram[11][95] , \ram[11][94] , \ram[11][93] , \ram[11][92] ,
         \ram[11][91] , \ram[11][90] , \ram[11][89] , \ram[11][88] ,
         \ram[11][87] , \ram[11][86] , \ram[11][85] , \ram[11][84] ,
         \ram[11][83] , \ram[11][82] , \ram[11][81] , \ram[11][80] ,
         \ram[11][79] , \ram[11][78] , \ram[11][77] , \ram[11][76] ,
         \ram[11][75] , \ram[11][74] , \ram[11][73] , \ram[11][72] ,
         \ram[11][71] , \ram[11][70] , \ram[11][69] , \ram[11][68] ,
         \ram[11][67] , \ram[11][66] , \ram[11][65] , \ram[11][64] ,
         \ram[11][63] , \ram[11][62] , \ram[11][61] , \ram[11][60] ,
         \ram[11][59] , \ram[11][58] , \ram[11][57] , \ram[11][56] ,
         \ram[11][55] , \ram[11][54] , \ram[11][53] , \ram[11][52] ,
         \ram[11][51] , \ram[11][50] , \ram[11][49] , \ram[11][48] ,
         \ram[11][47] , \ram[11][46] , \ram[11][45] , \ram[11][44] ,
         \ram[11][43] , \ram[11][42] , \ram[11][41] , \ram[11][40] ,
         \ram[11][39] , \ram[11][38] , \ram[11][37] , \ram[11][36] ,
         \ram[11][35] , \ram[11][34] , \ram[11][33] , \ram[11][32] ,
         \ram[11][31] , \ram[11][30] , \ram[11][29] , \ram[11][28] ,
         \ram[11][27] , \ram[11][26] , \ram[11][25] , \ram[11][24] ,
         \ram[11][23] , \ram[11][22] , \ram[11][21] , \ram[11][20] ,
         \ram[11][19] , \ram[11][18] , \ram[11][17] , \ram[11][16] ,
         \ram[11][15] , \ram[11][14] , \ram[11][13] , \ram[11][12] ,
         \ram[11][11] , \ram[11][10] , \ram[11][9] , \ram[11][8] ,
         \ram[11][7] , \ram[11][6] , \ram[11][5] , \ram[11][4] , \ram[11][3] ,
         \ram[11][2] , \ram[11][1] , \ram[11][0] , \ram[10][255] ,
         \ram[10][254] , \ram[10][253] , \ram[10][252] , \ram[10][251] ,
         \ram[10][250] , \ram[10][249] , \ram[10][248] , \ram[10][247] ,
         \ram[10][246] , \ram[10][245] , \ram[10][244] , \ram[10][243] ,
         \ram[10][242] , \ram[10][241] , \ram[10][240] , \ram[10][239] ,
         \ram[10][238] , \ram[10][237] , \ram[10][236] , \ram[10][235] ,
         \ram[10][234] , \ram[10][233] , \ram[10][232] , \ram[10][231] ,
         \ram[10][230] , \ram[10][229] , \ram[10][228] , \ram[10][227] ,
         \ram[10][226] , \ram[10][225] , \ram[10][224] , \ram[10][223] ,
         \ram[10][222] , \ram[10][221] , \ram[10][220] , \ram[10][219] ,
         \ram[10][218] , \ram[10][217] , \ram[10][216] , \ram[10][215] ,
         \ram[10][214] , \ram[10][213] , \ram[10][212] , \ram[10][211] ,
         \ram[10][210] , \ram[10][209] , \ram[10][208] , \ram[10][207] ,
         \ram[10][206] , \ram[10][205] , \ram[10][204] , \ram[10][203] ,
         \ram[10][202] , \ram[10][201] , \ram[10][200] , \ram[10][199] ,
         \ram[10][198] , \ram[10][197] , \ram[10][196] , \ram[10][195] ,
         \ram[10][194] , \ram[10][193] , \ram[10][192] , \ram[10][191] ,
         \ram[10][190] , \ram[10][189] , \ram[10][188] , \ram[10][187] ,
         \ram[10][186] , \ram[10][185] , \ram[10][184] , \ram[10][183] ,
         \ram[10][182] , \ram[10][181] , \ram[10][180] , \ram[10][179] ,
         \ram[10][178] , \ram[10][177] , \ram[10][176] , \ram[10][175] ,
         \ram[10][174] , \ram[10][173] , \ram[10][172] , \ram[10][171] ,
         \ram[10][170] , \ram[10][169] , \ram[10][168] , \ram[10][167] ,
         \ram[10][166] , \ram[10][165] , \ram[10][164] , \ram[10][163] ,
         \ram[10][162] , \ram[10][161] , \ram[10][160] , \ram[10][159] ,
         \ram[10][158] , \ram[10][157] , \ram[10][156] , \ram[10][155] ,
         \ram[10][154] , \ram[10][153] , \ram[10][152] , \ram[10][151] ,
         \ram[10][150] , \ram[10][149] , \ram[10][148] , \ram[10][147] ,
         \ram[10][146] , \ram[10][145] , \ram[10][144] , \ram[10][143] ,
         \ram[10][142] , \ram[10][141] , \ram[10][140] , \ram[10][139] ,
         \ram[10][138] , \ram[10][137] , \ram[10][136] , \ram[10][135] ,
         \ram[10][134] , \ram[10][133] , \ram[10][132] , \ram[10][131] ,
         \ram[10][130] , \ram[10][129] , \ram[10][128] , \ram[10][127] ,
         \ram[10][126] , \ram[10][125] , \ram[10][124] , \ram[10][123] ,
         \ram[10][122] , \ram[10][121] , \ram[10][120] , \ram[10][119] ,
         \ram[10][118] , \ram[10][117] , \ram[10][116] , \ram[10][115] ,
         \ram[10][114] , \ram[10][113] , \ram[10][112] , \ram[10][111] ,
         \ram[10][110] , \ram[10][109] , \ram[10][108] , \ram[10][107] ,
         \ram[10][106] , \ram[10][105] , \ram[10][104] , \ram[10][103] ,
         \ram[10][102] , \ram[10][101] , \ram[10][100] , \ram[10][99] ,
         \ram[10][98] , \ram[10][97] , \ram[10][96] , \ram[10][95] ,
         \ram[10][94] , \ram[10][93] , \ram[10][92] , \ram[10][91] ,
         \ram[10][90] , \ram[10][89] , \ram[10][88] , \ram[10][87] ,
         \ram[10][86] , \ram[10][85] , \ram[10][84] , \ram[10][83] ,
         \ram[10][82] , \ram[10][81] , \ram[10][80] , \ram[10][79] ,
         \ram[10][78] , \ram[10][77] , \ram[10][76] , \ram[10][75] ,
         \ram[10][74] , \ram[10][73] , \ram[10][72] , \ram[10][71] ,
         \ram[10][70] , \ram[10][69] , \ram[10][68] , \ram[10][67] ,
         \ram[10][66] , \ram[10][65] , \ram[10][64] , \ram[10][63] ,
         \ram[10][62] , \ram[10][61] , \ram[10][60] , \ram[10][59] ,
         \ram[10][58] , \ram[10][57] , \ram[10][56] , \ram[10][55] ,
         \ram[10][54] , \ram[10][53] , \ram[10][52] , \ram[10][51] ,
         \ram[10][50] , \ram[10][49] , \ram[10][48] , \ram[10][47] ,
         \ram[10][46] , \ram[10][45] , \ram[10][44] , \ram[10][43] ,
         \ram[10][42] , \ram[10][41] , \ram[10][40] , \ram[10][39] ,
         \ram[10][38] , \ram[10][37] , \ram[10][36] , \ram[10][35] ,
         \ram[10][34] , \ram[10][33] , \ram[10][32] , \ram[10][31] ,
         \ram[10][30] , \ram[10][29] , \ram[10][28] , \ram[10][27] ,
         \ram[10][26] , \ram[10][25] , \ram[10][24] , \ram[10][23] ,
         \ram[10][22] , \ram[10][21] , \ram[10][20] , \ram[10][19] ,
         \ram[10][18] , \ram[10][17] , \ram[10][16] , \ram[10][15] ,
         \ram[10][14] , \ram[10][13] , \ram[10][12] , \ram[10][11] ,
         \ram[10][10] , \ram[10][9] , \ram[10][8] , \ram[10][7] , \ram[10][6] ,
         \ram[10][5] , \ram[10][4] , \ram[10][3] , \ram[10][2] , \ram[10][1] ,
         \ram[10][0] , \ram[9][255] , \ram[9][254] , \ram[9][253] ,
         \ram[9][252] , \ram[9][251] , \ram[9][250] , \ram[9][249] ,
         \ram[9][248] , \ram[9][247] , \ram[9][246] , \ram[9][245] ,
         \ram[9][244] , \ram[9][243] , \ram[9][242] , \ram[9][241] ,
         \ram[9][240] , \ram[9][239] , \ram[9][238] , \ram[9][237] ,
         \ram[9][236] , \ram[9][235] , \ram[9][234] , \ram[9][233] ,
         \ram[9][232] , \ram[9][231] , \ram[9][230] , \ram[9][229] ,
         \ram[9][228] , \ram[9][227] , \ram[9][226] , \ram[9][225] ,
         \ram[9][224] , \ram[9][223] , \ram[9][222] , \ram[9][221] ,
         \ram[9][220] , \ram[9][219] , \ram[9][218] , \ram[9][217] ,
         \ram[9][216] , \ram[9][215] , \ram[9][214] , \ram[9][213] ,
         \ram[9][212] , \ram[9][211] , \ram[9][210] , \ram[9][209] ,
         \ram[9][208] , \ram[9][207] , \ram[9][206] , \ram[9][205] ,
         \ram[9][204] , \ram[9][203] , \ram[9][202] , \ram[9][201] ,
         \ram[9][200] , \ram[9][199] , \ram[9][198] , \ram[9][197] ,
         \ram[9][196] , \ram[9][195] , \ram[9][194] , \ram[9][193] ,
         \ram[9][192] , \ram[9][191] , \ram[9][190] , \ram[9][189] ,
         \ram[9][188] , \ram[9][187] , \ram[9][186] , \ram[9][185] ,
         \ram[9][184] , \ram[9][183] , \ram[9][182] , \ram[9][181] ,
         \ram[9][180] , \ram[9][179] , \ram[9][178] , \ram[9][177] ,
         \ram[9][176] , \ram[9][175] , \ram[9][174] , \ram[9][173] ,
         \ram[9][172] , \ram[9][171] , \ram[9][170] , \ram[9][169] ,
         \ram[9][168] , \ram[9][167] , \ram[9][166] , \ram[9][165] ,
         \ram[9][164] , \ram[9][163] , \ram[9][162] , \ram[9][161] ,
         \ram[9][160] , \ram[9][159] , \ram[9][158] , \ram[9][157] ,
         \ram[9][156] , \ram[9][155] , \ram[9][154] , \ram[9][153] ,
         \ram[9][152] , \ram[9][151] , \ram[9][150] , \ram[9][149] ,
         \ram[9][148] , \ram[9][147] , \ram[9][146] , \ram[9][145] ,
         \ram[9][144] , \ram[9][143] , \ram[9][142] , \ram[9][141] ,
         \ram[9][140] , \ram[9][139] , \ram[9][138] , \ram[9][137] ,
         \ram[9][136] , \ram[9][135] , \ram[9][134] , \ram[9][133] ,
         \ram[9][132] , \ram[9][131] , \ram[9][130] , \ram[9][129] ,
         \ram[9][128] , \ram[9][127] , \ram[9][126] , \ram[9][125] ,
         \ram[9][124] , \ram[9][123] , \ram[9][122] , \ram[9][121] ,
         \ram[9][120] , \ram[9][119] , \ram[9][118] , \ram[9][117] ,
         \ram[9][116] , \ram[9][115] , \ram[9][114] , \ram[9][113] ,
         \ram[9][112] , \ram[9][111] , \ram[9][110] , \ram[9][109] ,
         \ram[9][108] , \ram[9][107] , \ram[9][106] , \ram[9][105] ,
         \ram[9][104] , \ram[9][103] , \ram[9][102] , \ram[9][101] ,
         \ram[9][100] , \ram[9][99] , \ram[9][98] , \ram[9][97] , \ram[9][96] ,
         \ram[9][95] , \ram[9][94] , \ram[9][93] , \ram[9][92] , \ram[9][91] ,
         \ram[9][90] , \ram[9][89] , \ram[9][88] , \ram[9][87] , \ram[9][86] ,
         \ram[9][85] , \ram[9][84] , \ram[9][83] , \ram[9][82] , \ram[9][81] ,
         \ram[9][80] , \ram[9][79] , \ram[9][78] , \ram[9][77] , \ram[9][76] ,
         \ram[9][75] , \ram[9][74] , \ram[9][73] , \ram[9][72] , \ram[9][71] ,
         \ram[9][70] , \ram[9][69] , \ram[9][68] , \ram[9][67] , \ram[9][66] ,
         \ram[9][65] , \ram[9][64] , \ram[9][63] , \ram[9][62] , \ram[9][61] ,
         \ram[9][60] , \ram[9][59] , \ram[9][58] , \ram[9][57] , \ram[9][56] ,
         \ram[9][55] , \ram[9][54] , \ram[9][53] , \ram[9][52] , \ram[9][51] ,
         \ram[9][50] , \ram[9][49] , \ram[9][48] , \ram[9][47] , \ram[9][46] ,
         \ram[9][45] , \ram[9][44] , \ram[9][43] , \ram[9][42] , \ram[9][41] ,
         \ram[9][40] , \ram[9][39] , \ram[9][38] , \ram[9][37] , \ram[9][36] ,
         \ram[9][35] , \ram[9][34] , \ram[9][33] , \ram[9][32] , \ram[9][31] ,
         \ram[9][30] , \ram[9][29] , \ram[9][28] , \ram[9][27] , \ram[9][26] ,
         \ram[9][25] , \ram[9][24] , \ram[9][23] , \ram[9][22] , \ram[9][21] ,
         \ram[9][20] , \ram[9][19] , \ram[9][18] , \ram[9][17] , \ram[9][16] ,
         \ram[9][15] , \ram[9][14] , \ram[9][13] , \ram[9][12] , \ram[9][11] ,
         \ram[9][10] , \ram[9][9] , \ram[9][8] , \ram[9][7] , \ram[9][6] ,
         \ram[9][5] , \ram[9][4] , \ram[9][3] , \ram[9][2] , \ram[9][1] ,
         \ram[9][0] , \ram[8][255] , \ram[8][254] , \ram[8][253] ,
         \ram[8][252] , \ram[8][251] , \ram[8][250] , \ram[8][249] ,
         \ram[8][248] , \ram[8][247] , \ram[8][246] , \ram[8][245] ,
         \ram[8][244] , \ram[8][243] , \ram[8][242] , \ram[8][241] ,
         \ram[8][240] , \ram[8][239] , \ram[8][238] , \ram[8][237] ,
         \ram[8][236] , \ram[8][235] , \ram[8][234] , \ram[8][233] ,
         \ram[8][232] , \ram[8][231] , \ram[8][230] , \ram[8][229] ,
         \ram[8][228] , \ram[8][227] , \ram[8][226] , \ram[8][225] ,
         \ram[8][224] , \ram[8][223] , \ram[8][222] , \ram[8][221] ,
         \ram[8][220] , \ram[8][219] , \ram[8][218] , \ram[8][217] ,
         \ram[8][216] , \ram[8][215] , \ram[8][214] , \ram[8][213] ,
         \ram[8][212] , \ram[8][211] , \ram[8][210] , \ram[8][209] ,
         \ram[8][208] , \ram[8][207] , \ram[8][206] , \ram[8][205] ,
         \ram[8][204] , \ram[8][203] , \ram[8][202] , \ram[8][201] ,
         \ram[8][200] , \ram[8][199] , \ram[8][198] , \ram[8][197] ,
         \ram[8][196] , \ram[8][195] , \ram[8][194] , \ram[8][193] ,
         \ram[8][192] , \ram[8][191] , \ram[8][190] , \ram[8][189] ,
         \ram[8][188] , \ram[8][187] , \ram[8][186] , \ram[8][185] ,
         \ram[8][184] , \ram[8][183] , \ram[8][182] , \ram[8][181] ,
         \ram[8][180] , \ram[8][179] , \ram[8][178] , \ram[8][177] ,
         \ram[8][176] , \ram[8][175] , \ram[8][174] , \ram[8][173] ,
         \ram[8][172] , \ram[8][171] , \ram[8][170] , \ram[8][169] ,
         \ram[8][168] , \ram[8][167] , \ram[8][166] , \ram[8][165] ,
         \ram[8][164] , \ram[8][163] , \ram[8][162] , \ram[8][161] ,
         \ram[8][160] , \ram[8][159] , \ram[8][158] , \ram[8][157] ,
         \ram[8][156] , \ram[8][155] , \ram[8][154] , \ram[8][153] ,
         \ram[8][152] , \ram[8][151] , \ram[8][150] , \ram[8][149] ,
         \ram[8][148] , \ram[8][147] , \ram[8][146] , \ram[8][145] ,
         \ram[8][144] , \ram[8][143] , \ram[8][142] , \ram[8][141] ,
         \ram[8][140] , \ram[8][139] , \ram[8][138] , \ram[8][137] ,
         \ram[8][136] , \ram[8][135] , \ram[8][134] , \ram[8][133] ,
         \ram[8][132] , \ram[8][131] , \ram[8][130] , \ram[8][129] ,
         \ram[8][128] , \ram[8][127] , \ram[8][126] , \ram[8][125] ,
         \ram[8][124] , \ram[8][123] , \ram[8][122] , \ram[8][121] ,
         \ram[8][120] , \ram[8][119] , \ram[8][118] , \ram[8][117] ,
         \ram[8][116] , \ram[8][115] , \ram[8][114] , \ram[8][113] ,
         \ram[8][112] , \ram[8][111] , \ram[8][110] , \ram[8][109] ,
         \ram[8][108] , \ram[8][107] , \ram[8][106] , \ram[8][105] ,
         \ram[8][104] , \ram[8][103] , \ram[8][102] , \ram[8][101] ,
         \ram[8][100] , \ram[8][99] , \ram[8][98] , \ram[8][97] , \ram[8][96] ,
         \ram[8][95] , \ram[8][94] , \ram[8][93] , \ram[8][92] , \ram[8][91] ,
         \ram[8][90] , \ram[8][89] , \ram[8][88] , \ram[8][87] , \ram[8][86] ,
         \ram[8][85] , \ram[8][84] , \ram[8][83] , \ram[8][82] , \ram[8][81] ,
         \ram[8][80] , \ram[8][79] , \ram[8][78] , \ram[8][77] , \ram[8][76] ,
         \ram[8][75] , \ram[8][74] , \ram[8][73] , \ram[8][72] , \ram[8][71] ,
         \ram[8][70] , \ram[8][69] , \ram[8][68] , \ram[8][67] , \ram[8][66] ,
         \ram[8][65] , \ram[8][64] , \ram[8][63] , \ram[8][62] , \ram[8][61] ,
         \ram[8][60] , \ram[8][59] , \ram[8][58] , \ram[8][57] , \ram[8][56] ,
         \ram[8][55] , \ram[8][54] , \ram[8][53] , \ram[8][52] , \ram[8][51] ,
         \ram[8][50] , \ram[8][49] , \ram[8][48] , \ram[8][47] , \ram[8][46] ,
         \ram[8][45] , \ram[8][44] , \ram[8][43] , \ram[8][42] , \ram[8][41] ,
         \ram[8][40] , \ram[8][39] , \ram[8][38] , \ram[8][37] , \ram[8][36] ,
         \ram[8][35] , \ram[8][34] , \ram[8][33] , \ram[8][32] , \ram[8][31] ,
         \ram[8][30] , \ram[8][29] , \ram[8][28] , \ram[8][27] , \ram[8][26] ,
         \ram[8][25] , \ram[8][24] , \ram[8][23] , \ram[8][22] , \ram[8][21] ,
         \ram[8][20] , \ram[8][19] , \ram[8][18] , \ram[8][17] , \ram[8][16] ,
         \ram[8][15] , \ram[8][14] , \ram[8][13] , \ram[8][12] , \ram[8][11] ,
         \ram[8][10] , \ram[8][9] , \ram[8][8] , \ram[8][7] , \ram[8][6] ,
         \ram[8][5] , \ram[8][4] , \ram[8][3] , \ram[8][2] , \ram[8][1] ,
         \ram[8][0] , \ram[7][255] , \ram[7][254] , \ram[7][253] ,
         \ram[7][252] , \ram[7][251] , \ram[7][250] , \ram[7][249] ,
         \ram[7][248] , \ram[7][247] , \ram[7][246] , \ram[7][245] ,
         \ram[7][244] , \ram[7][243] , \ram[7][242] , \ram[7][241] ,
         \ram[7][240] , \ram[7][239] , \ram[7][238] , \ram[7][237] ,
         \ram[7][236] , \ram[7][235] , \ram[7][234] , \ram[7][233] ,
         \ram[7][232] , \ram[7][231] , \ram[7][230] , \ram[7][229] ,
         \ram[7][228] , \ram[7][227] , \ram[7][226] , \ram[7][225] ,
         \ram[7][224] , \ram[7][223] , \ram[7][222] , \ram[7][221] ,
         \ram[7][220] , \ram[7][219] , \ram[7][218] , \ram[7][217] ,
         \ram[7][216] , \ram[7][215] , \ram[7][214] , \ram[7][213] ,
         \ram[7][212] , \ram[7][211] , \ram[7][210] , \ram[7][209] ,
         \ram[7][208] , \ram[7][207] , \ram[7][206] , \ram[7][205] ,
         \ram[7][204] , \ram[7][203] , \ram[7][202] , \ram[7][201] ,
         \ram[7][200] , \ram[7][199] , \ram[7][198] , \ram[7][197] ,
         \ram[7][196] , \ram[7][195] , \ram[7][194] , \ram[7][193] ,
         \ram[7][192] , \ram[7][191] , \ram[7][190] , \ram[7][189] ,
         \ram[7][188] , \ram[7][187] , \ram[7][186] , \ram[7][185] ,
         \ram[7][184] , \ram[7][183] , \ram[7][182] , \ram[7][181] ,
         \ram[7][180] , \ram[7][179] , \ram[7][178] , \ram[7][177] ,
         \ram[7][176] , \ram[7][175] , \ram[7][174] , \ram[7][173] ,
         \ram[7][172] , \ram[7][171] , \ram[7][170] , \ram[7][169] ,
         \ram[7][168] , \ram[7][167] , \ram[7][166] , \ram[7][165] ,
         \ram[7][164] , \ram[7][163] , \ram[7][162] , \ram[7][161] ,
         \ram[7][160] , \ram[7][159] , \ram[7][158] , \ram[7][157] ,
         \ram[7][156] , \ram[7][155] , \ram[7][154] , \ram[7][153] ,
         \ram[7][152] , \ram[7][151] , \ram[7][150] , \ram[7][149] ,
         \ram[7][148] , \ram[7][147] , \ram[7][146] , \ram[7][145] ,
         \ram[7][144] , \ram[7][143] , \ram[7][142] , \ram[7][141] ,
         \ram[7][140] , \ram[7][139] , \ram[7][138] , \ram[7][137] ,
         \ram[7][136] , \ram[7][135] , \ram[7][134] , \ram[7][133] ,
         \ram[7][132] , \ram[7][131] , \ram[7][130] , \ram[7][129] ,
         \ram[7][128] , \ram[7][127] , \ram[7][126] , \ram[7][125] ,
         \ram[7][124] , \ram[7][123] , \ram[7][122] , \ram[7][121] ,
         \ram[7][120] , \ram[7][119] , \ram[7][118] , \ram[7][117] ,
         \ram[7][116] , \ram[7][115] , \ram[7][114] , \ram[7][113] ,
         \ram[7][112] , \ram[7][111] , \ram[7][110] , \ram[7][109] ,
         \ram[7][108] , \ram[7][107] , \ram[7][106] , \ram[7][105] ,
         \ram[7][104] , \ram[7][103] , \ram[7][102] , \ram[7][101] ,
         \ram[7][100] , \ram[7][99] , \ram[7][98] , \ram[7][97] , \ram[7][96] ,
         \ram[7][95] , \ram[7][94] , \ram[7][93] , \ram[7][92] , \ram[7][91] ,
         \ram[7][90] , \ram[7][89] , \ram[7][88] , \ram[7][87] , \ram[7][86] ,
         \ram[7][85] , \ram[7][84] , \ram[7][83] , \ram[7][82] , \ram[7][81] ,
         \ram[7][80] , \ram[7][79] , \ram[7][78] , \ram[7][77] , \ram[7][76] ,
         \ram[7][75] , \ram[7][74] , \ram[7][73] , \ram[7][72] , \ram[7][71] ,
         \ram[7][70] , \ram[7][69] , \ram[7][68] , \ram[7][67] , \ram[7][66] ,
         \ram[7][65] , \ram[7][64] , \ram[7][63] , \ram[7][62] , \ram[7][61] ,
         \ram[7][60] , \ram[7][59] , \ram[7][58] , \ram[7][57] , \ram[7][56] ,
         \ram[7][55] , \ram[7][54] , \ram[7][53] , \ram[7][52] , \ram[7][51] ,
         \ram[7][50] , \ram[7][49] , \ram[7][48] , \ram[7][47] , \ram[7][46] ,
         \ram[7][45] , \ram[7][44] , \ram[7][43] , \ram[7][42] , \ram[7][41] ,
         \ram[7][40] , \ram[7][39] , \ram[7][38] , \ram[7][37] , \ram[7][36] ,
         \ram[7][35] , \ram[7][34] , \ram[7][33] , \ram[7][32] , \ram[7][31] ,
         \ram[7][30] , \ram[7][29] , \ram[7][28] , \ram[7][27] , \ram[7][26] ,
         \ram[7][25] , \ram[7][24] , \ram[7][23] , \ram[7][22] , \ram[7][21] ,
         \ram[7][20] , \ram[7][19] , \ram[7][18] , \ram[7][17] , \ram[7][16] ,
         \ram[7][15] , \ram[7][14] , \ram[7][13] , \ram[7][12] , \ram[7][11] ,
         \ram[7][10] , \ram[7][9] , \ram[7][8] , \ram[7][7] , \ram[7][6] ,
         \ram[7][5] , \ram[7][4] , \ram[7][3] , \ram[7][2] , \ram[7][1] ,
         \ram[7][0] , \ram[6][255] , \ram[6][254] , \ram[6][253] ,
         \ram[6][252] , \ram[6][251] , \ram[6][250] , \ram[6][249] ,
         \ram[6][248] , \ram[6][247] , \ram[6][246] , \ram[6][245] ,
         \ram[6][244] , \ram[6][243] , \ram[6][242] , \ram[6][241] ,
         \ram[6][240] , \ram[6][239] , \ram[6][238] , \ram[6][237] ,
         \ram[6][236] , \ram[6][235] , \ram[6][234] , \ram[6][233] ,
         \ram[6][232] , \ram[6][231] , \ram[6][230] , \ram[6][229] ,
         \ram[6][228] , \ram[6][227] , \ram[6][226] , \ram[6][225] ,
         \ram[6][224] , \ram[6][223] , \ram[6][222] , \ram[6][221] ,
         \ram[6][220] , \ram[6][219] , \ram[6][218] , \ram[6][217] ,
         \ram[6][216] , \ram[6][215] , \ram[6][214] , \ram[6][213] ,
         \ram[6][212] , \ram[6][211] , \ram[6][210] , \ram[6][209] ,
         \ram[6][208] , \ram[6][207] , \ram[6][206] , \ram[6][205] ,
         \ram[6][204] , \ram[6][203] , \ram[6][202] , \ram[6][201] ,
         \ram[6][200] , \ram[6][199] , \ram[6][198] , \ram[6][197] ,
         \ram[6][196] , \ram[6][195] , \ram[6][194] , \ram[6][193] ,
         \ram[6][192] , \ram[6][191] , \ram[6][190] , \ram[6][189] ,
         \ram[6][188] , \ram[6][187] , \ram[6][186] , \ram[6][185] ,
         \ram[6][184] , \ram[6][183] , \ram[6][182] , \ram[6][181] ,
         \ram[6][180] , \ram[6][179] , \ram[6][178] , \ram[6][177] ,
         \ram[6][176] , \ram[6][175] , \ram[6][174] , \ram[6][173] ,
         \ram[6][172] , \ram[6][171] , \ram[6][170] , \ram[6][169] ,
         \ram[6][168] , \ram[6][167] , \ram[6][166] , \ram[6][165] ,
         \ram[6][164] , \ram[6][163] , \ram[6][162] , \ram[6][161] ,
         \ram[6][160] , \ram[6][159] , \ram[6][158] , \ram[6][157] ,
         \ram[6][156] , \ram[6][155] , \ram[6][154] , \ram[6][153] ,
         \ram[6][152] , \ram[6][151] , \ram[6][150] , \ram[6][149] ,
         \ram[6][148] , \ram[6][147] , \ram[6][146] , \ram[6][145] ,
         \ram[6][144] , \ram[6][143] , \ram[6][142] , \ram[6][141] ,
         \ram[6][140] , \ram[6][139] , \ram[6][138] , \ram[6][137] ,
         \ram[6][136] , \ram[6][135] , \ram[6][134] , \ram[6][133] ,
         \ram[6][132] , \ram[6][131] , \ram[6][130] , \ram[6][129] ,
         \ram[6][128] , \ram[6][127] , \ram[6][126] , \ram[6][125] ,
         \ram[6][124] , \ram[6][123] , \ram[6][122] , \ram[6][121] ,
         \ram[6][120] , \ram[6][119] , \ram[6][118] , \ram[6][117] ,
         \ram[6][116] , \ram[6][115] , \ram[6][114] , \ram[6][113] ,
         \ram[6][112] , \ram[6][111] , \ram[6][110] , \ram[6][109] ,
         \ram[6][108] , \ram[6][107] , \ram[6][106] , \ram[6][105] ,
         \ram[6][104] , \ram[6][103] , \ram[6][102] , \ram[6][101] ,
         \ram[6][100] , \ram[6][99] , \ram[6][98] , \ram[6][97] , \ram[6][96] ,
         \ram[6][95] , \ram[6][94] , \ram[6][93] , \ram[6][92] , \ram[6][91] ,
         \ram[6][90] , \ram[6][89] , \ram[6][88] , \ram[6][87] , \ram[6][86] ,
         \ram[6][85] , \ram[6][84] , \ram[6][83] , \ram[6][82] , \ram[6][81] ,
         \ram[6][80] , \ram[6][79] , \ram[6][78] , \ram[6][77] , \ram[6][76] ,
         \ram[6][75] , \ram[6][74] , \ram[6][73] , \ram[6][72] , \ram[6][71] ,
         \ram[6][70] , \ram[6][69] , \ram[6][68] , \ram[6][67] , \ram[6][66] ,
         \ram[6][65] , \ram[6][64] , \ram[6][63] , \ram[6][62] , \ram[6][61] ,
         \ram[6][60] , \ram[6][59] , \ram[6][58] , \ram[6][57] , \ram[6][56] ,
         \ram[6][55] , \ram[6][54] , \ram[6][53] , \ram[6][52] , \ram[6][51] ,
         \ram[6][50] , \ram[6][49] , \ram[6][48] , \ram[6][47] , \ram[6][46] ,
         \ram[6][45] , \ram[6][44] , \ram[6][43] , \ram[6][42] , \ram[6][41] ,
         \ram[6][40] , \ram[6][39] , \ram[6][38] , \ram[6][37] , \ram[6][36] ,
         \ram[6][35] , \ram[6][34] , \ram[6][33] , \ram[6][32] , \ram[6][31] ,
         \ram[6][30] , \ram[6][29] , \ram[6][28] , \ram[6][27] , \ram[6][26] ,
         \ram[6][25] , \ram[6][24] , \ram[6][23] , \ram[6][22] , \ram[6][21] ,
         \ram[6][20] , \ram[6][19] , \ram[6][18] , \ram[6][17] , \ram[6][16] ,
         \ram[6][15] , \ram[6][14] , \ram[6][13] , \ram[6][12] , \ram[6][11] ,
         \ram[6][10] , \ram[6][9] , \ram[6][8] , \ram[6][7] , \ram[6][6] ,
         \ram[6][5] , \ram[6][4] , \ram[6][3] , \ram[6][2] , \ram[6][1] ,
         \ram[6][0] , \ram[5][255] , \ram[5][254] , \ram[5][253] ,
         \ram[5][252] , \ram[5][251] , \ram[5][250] , \ram[5][249] ,
         \ram[5][248] , \ram[5][247] , \ram[5][246] , \ram[5][245] ,
         \ram[5][244] , \ram[5][243] , \ram[5][242] , \ram[5][241] ,
         \ram[5][240] , \ram[5][239] , \ram[5][238] , \ram[5][237] ,
         \ram[5][236] , \ram[5][235] , \ram[5][234] , \ram[5][233] ,
         \ram[5][232] , \ram[5][231] , \ram[5][230] , \ram[5][229] ,
         \ram[5][228] , \ram[5][227] , \ram[5][226] , \ram[5][225] ,
         \ram[5][224] , \ram[5][223] , \ram[5][222] , \ram[5][221] ,
         \ram[5][220] , \ram[5][219] , \ram[5][218] , \ram[5][217] ,
         \ram[5][216] , \ram[5][215] , \ram[5][214] , \ram[5][213] ,
         \ram[5][212] , \ram[5][211] , \ram[5][210] , \ram[5][209] ,
         \ram[5][208] , \ram[5][207] , \ram[5][206] , \ram[5][205] ,
         \ram[5][204] , \ram[5][203] , \ram[5][202] , \ram[5][201] ,
         \ram[5][200] , \ram[5][199] , \ram[5][198] , \ram[5][197] ,
         \ram[5][196] , \ram[5][195] , \ram[5][194] , \ram[5][193] ,
         \ram[5][192] , \ram[5][191] , \ram[5][190] , \ram[5][189] ,
         \ram[5][188] , \ram[5][187] , \ram[5][186] , \ram[5][185] ,
         \ram[5][184] , \ram[5][183] , \ram[5][182] , \ram[5][181] ,
         \ram[5][180] , \ram[5][179] , \ram[5][178] , \ram[5][177] ,
         \ram[5][176] , \ram[5][175] , \ram[5][174] , \ram[5][173] ,
         \ram[5][172] , \ram[5][171] , \ram[5][170] , \ram[5][169] ,
         \ram[5][168] , \ram[5][167] , \ram[5][166] , \ram[5][165] ,
         \ram[5][164] , \ram[5][163] , \ram[5][162] , \ram[5][161] ,
         \ram[5][160] , \ram[5][159] , \ram[5][158] , \ram[5][157] ,
         \ram[5][156] , \ram[5][155] , \ram[5][154] , \ram[5][153] ,
         \ram[5][152] , \ram[5][151] , \ram[5][150] , \ram[5][149] ,
         \ram[5][148] , \ram[5][147] , \ram[5][146] , \ram[5][145] ,
         \ram[5][144] , \ram[5][143] , \ram[5][142] , \ram[5][141] ,
         \ram[5][140] , \ram[5][139] , \ram[5][138] , \ram[5][137] ,
         \ram[5][136] , \ram[5][135] , \ram[5][134] , \ram[5][133] ,
         \ram[5][132] , \ram[5][131] , \ram[5][130] , \ram[5][129] ,
         \ram[5][128] , \ram[5][127] , \ram[5][126] , \ram[5][125] ,
         \ram[5][124] , \ram[5][123] , \ram[5][122] , \ram[5][121] ,
         \ram[5][120] , \ram[5][119] , \ram[5][118] , \ram[5][117] ,
         \ram[5][116] , \ram[5][115] , \ram[5][114] , \ram[5][113] ,
         \ram[5][112] , \ram[5][111] , \ram[5][110] , \ram[5][109] ,
         \ram[5][108] , \ram[5][107] , \ram[5][106] , \ram[5][105] ,
         \ram[5][104] , \ram[5][103] , \ram[5][102] , \ram[5][101] ,
         \ram[5][100] , \ram[5][99] , \ram[5][98] , \ram[5][97] , \ram[5][96] ,
         \ram[5][95] , \ram[5][94] , \ram[5][93] , \ram[5][92] , \ram[5][91] ,
         \ram[5][90] , \ram[5][89] , \ram[5][88] , \ram[5][87] , \ram[5][86] ,
         \ram[5][85] , \ram[5][84] , \ram[5][83] , \ram[5][82] , \ram[5][81] ,
         \ram[5][80] , \ram[5][79] , \ram[5][78] , \ram[5][77] , \ram[5][76] ,
         \ram[5][75] , \ram[5][74] , \ram[5][73] , \ram[5][72] , \ram[5][71] ,
         \ram[5][70] , \ram[5][69] , \ram[5][68] , \ram[5][67] , \ram[5][66] ,
         \ram[5][65] , \ram[5][64] , \ram[5][63] , \ram[5][62] , \ram[5][61] ,
         \ram[5][60] , \ram[5][59] , \ram[5][58] , \ram[5][57] , \ram[5][56] ,
         \ram[5][55] , \ram[5][54] , \ram[5][53] , \ram[5][52] , \ram[5][51] ,
         \ram[5][50] , \ram[5][49] , \ram[5][48] , \ram[5][47] , \ram[5][46] ,
         \ram[5][45] , \ram[5][44] , \ram[5][43] , \ram[5][42] , \ram[5][41] ,
         \ram[5][40] , \ram[5][39] , \ram[5][38] , \ram[5][37] , \ram[5][36] ,
         \ram[5][35] , \ram[5][34] , \ram[5][33] , \ram[5][32] , \ram[5][31] ,
         \ram[5][30] , \ram[5][29] , \ram[5][28] , \ram[5][27] , \ram[5][26] ,
         \ram[5][25] , \ram[5][24] , \ram[5][23] , \ram[5][22] , \ram[5][21] ,
         \ram[5][20] , \ram[5][19] , \ram[5][18] , \ram[5][17] , \ram[5][16] ,
         \ram[5][15] , \ram[5][14] , \ram[5][13] , \ram[5][12] , \ram[5][11] ,
         \ram[5][10] , \ram[5][9] , \ram[5][8] , \ram[5][7] , \ram[5][6] ,
         \ram[5][5] , \ram[5][4] , \ram[5][3] , \ram[5][2] , \ram[5][1] ,
         \ram[5][0] , \ram[4][255] , \ram[4][254] , \ram[4][253] ,
         \ram[4][252] , \ram[4][251] , \ram[4][250] , \ram[4][249] ,
         \ram[4][248] , \ram[4][247] , \ram[4][246] , \ram[4][245] ,
         \ram[4][244] , \ram[4][243] , \ram[4][242] , \ram[4][241] ,
         \ram[4][240] , \ram[4][239] , \ram[4][238] , \ram[4][237] ,
         \ram[4][236] , \ram[4][235] , \ram[4][234] , \ram[4][233] ,
         \ram[4][232] , \ram[4][231] , \ram[4][230] , \ram[4][229] ,
         \ram[4][228] , \ram[4][227] , \ram[4][226] , \ram[4][225] ,
         \ram[4][224] , \ram[4][223] , \ram[4][222] , \ram[4][221] ,
         \ram[4][220] , \ram[4][219] , \ram[4][218] , \ram[4][217] ,
         \ram[4][216] , \ram[4][215] , \ram[4][214] , \ram[4][213] ,
         \ram[4][212] , \ram[4][211] , \ram[4][210] , \ram[4][209] ,
         \ram[4][208] , \ram[4][207] , \ram[4][206] , \ram[4][205] ,
         \ram[4][204] , \ram[4][203] , \ram[4][202] , \ram[4][201] ,
         \ram[4][200] , \ram[4][199] , \ram[4][198] , \ram[4][197] ,
         \ram[4][196] , \ram[4][195] , \ram[4][194] , \ram[4][193] ,
         \ram[4][192] , \ram[4][191] , \ram[4][190] , \ram[4][189] ,
         \ram[4][188] , \ram[4][187] , \ram[4][186] , \ram[4][185] ,
         \ram[4][184] , \ram[4][183] , \ram[4][182] , \ram[4][181] ,
         \ram[4][180] , \ram[4][179] , \ram[4][178] , \ram[4][177] ,
         \ram[4][176] , \ram[4][175] , \ram[4][174] , \ram[4][173] ,
         \ram[4][172] , \ram[4][171] , \ram[4][170] , \ram[4][169] ,
         \ram[4][168] , \ram[4][167] , \ram[4][166] , \ram[4][165] ,
         \ram[4][164] , \ram[4][163] , \ram[4][162] , \ram[4][161] ,
         \ram[4][160] , \ram[4][159] , \ram[4][158] , \ram[4][157] ,
         \ram[4][156] , \ram[4][155] , \ram[4][154] , \ram[4][153] ,
         \ram[4][152] , \ram[4][151] , \ram[4][150] , \ram[4][149] ,
         \ram[4][148] , \ram[4][147] , \ram[4][146] , \ram[4][145] ,
         \ram[4][144] , \ram[4][143] , \ram[4][142] , \ram[4][141] ,
         \ram[4][140] , \ram[4][139] , \ram[4][138] , \ram[4][137] ,
         \ram[4][136] , \ram[4][135] , \ram[4][134] , \ram[4][133] ,
         \ram[4][132] , \ram[4][131] , \ram[4][130] , \ram[4][129] ,
         \ram[4][128] , \ram[4][127] , \ram[4][126] , \ram[4][125] ,
         \ram[4][124] , \ram[4][123] , \ram[4][122] , \ram[4][121] ,
         \ram[4][120] , \ram[4][119] , \ram[4][118] , \ram[4][117] ,
         \ram[4][116] , \ram[4][115] , \ram[4][114] , \ram[4][113] ,
         \ram[4][112] , \ram[4][111] , \ram[4][110] , \ram[4][109] ,
         \ram[4][108] , \ram[4][107] , \ram[4][106] , \ram[4][105] ,
         \ram[4][104] , \ram[4][103] , \ram[4][102] , \ram[4][101] ,
         \ram[4][100] , \ram[4][99] , \ram[4][98] , \ram[4][97] , \ram[4][96] ,
         \ram[4][95] , \ram[4][94] , \ram[4][93] , \ram[4][92] , \ram[4][91] ,
         \ram[4][90] , \ram[4][89] , \ram[4][88] , \ram[4][87] , \ram[4][86] ,
         \ram[4][85] , \ram[4][84] , \ram[4][83] , \ram[4][82] , \ram[4][81] ,
         \ram[4][80] , \ram[4][79] , \ram[4][78] , \ram[4][77] , \ram[4][76] ,
         \ram[4][75] , \ram[4][74] , \ram[4][73] , \ram[4][72] , \ram[4][71] ,
         \ram[4][70] , \ram[4][69] , \ram[4][68] , \ram[4][67] , \ram[4][66] ,
         \ram[4][65] , \ram[4][64] , \ram[4][63] , \ram[4][62] , \ram[4][61] ,
         \ram[4][60] , \ram[4][59] , \ram[4][58] , \ram[4][57] , \ram[4][56] ,
         \ram[4][55] , \ram[4][54] , \ram[4][53] , \ram[4][52] , \ram[4][51] ,
         \ram[4][50] , \ram[4][49] , \ram[4][48] , \ram[4][47] , \ram[4][46] ,
         \ram[4][45] , \ram[4][44] , \ram[4][43] , \ram[4][42] , \ram[4][41] ,
         \ram[4][40] , \ram[4][39] , \ram[4][38] , \ram[4][37] , \ram[4][36] ,
         \ram[4][35] , \ram[4][34] , \ram[4][33] , \ram[4][32] , \ram[4][31] ,
         \ram[4][30] , \ram[4][29] , \ram[4][28] , \ram[4][27] , \ram[4][26] ,
         \ram[4][25] , \ram[4][24] , \ram[4][23] , \ram[4][22] , \ram[4][21] ,
         \ram[4][20] , \ram[4][19] , \ram[4][18] , \ram[4][17] , \ram[4][16] ,
         \ram[4][15] , \ram[4][14] , \ram[4][13] , \ram[4][12] , \ram[4][11] ,
         \ram[4][10] , \ram[4][9] , \ram[4][8] , \ram[4][7] , \ram[4][6] ,
         \ram[4][5] , \ram[4][4] , \ram[4][3] , \ram[4][2] , \ram[4][1] ,
         \ram[4][0] , \ram[3][255] , \ram[3][254] , \ram[3][253] ,
         \ram[3][252] , \ram[3][251] , \ram[3][250] , \ram[3][249] ,
         \ram[3][248] , \ram[3][247] , \ram[3][246] , \ram[3][245] ,
         \ram[3][244] , \ram[3][243] , \ram[3][242] , \ram[3][241] ,
         \ram[3][240] , \ram[3][239] , \ram[3][238] , \ram[3][237] ,
         \ram[3][236] , \ram[3][235] , \ram[3][234] , \ram[3][233] ,
         \ram[3][232] , \ram[3][231] , \ram[3][230] , \ram[3][229] ,
         \ram[3][228] , \ram[3][227] , \ram[3][226] , \ram[3][225] ,
         \ram[3][224] , \ram[3][223] , \ram[3][222] , \ram[3][221] ,
         \ram[3][220] , \ram[3][219] , \ram[3][218] , \ram[3][217] ,
         \ram[3][216] , \ram[3][215] , \ram[3][214] , \ram[3][213] ,
         \ram[3][212] , \ram[3][211] , \ram[3][210] , \ram[3][209] ,
         \ram[3][208] , \ram[3][207] , \ram[3][206] , \ram[3][205] ,
         \ram[3][204] , \ram[3][203] , \ram[3][202] , \ram[3][201] ,
         \ram[3][200] , \ram[3][199] , \ram[3][198] , \ram[3][197] ,
         \ram[3][196] , \ram[3][195] , \ram[3][194] , \ram[3][193] ,
         \ram[3][192] , \ram[3][191] , \ram[3][190] , \ram[3][189] ,
         \ram[3][188] , \ram[3][187] , \ram[3][186] , \ram[3][185] ,
         \ram[3][184] , \ram[3][183] , \ram[3][182] , \ram[3][181] ,
         \ram[3][180] , \ram[3][179] , \ram[3][178] , \ram[3][177] ,
         \ram[3][176] , \ram[3][175] , \ram[3][174] , \ram[3][173] ,
         \ram[3][172] , \ram[3][171] , \ram[3][170] , \ram[3][169] ,
         \ram[3][168] , \ram[3][167] , \ram[3][166] , \ram[3][165] ,
         \ram[3][164] , \ram[3][163] , \ram[3][162] , \ram[3][161] ,
         \ram[3][160] , \ram[3][159] , \ram[3][158] , \ram[3][157] ,
         \ram[3][156] , \ram[3][155] , \ram[3][154] , \ram[3][153] ,
         \ram[3][152] , \ram[3][151] , \ram[3][150] , \ram[3][149] ,
         \ram[3][148] , \ram[3][147] , \ram[3][146] , \ram[3][145] ,
         \ram[3][144] , \ram[3][143] , \ram[3][142] , \ram[3][141] ,
         \ram[3][140] , \ram[3][139] , \ram[3][138] , \ram[3][137] ,
         \ram[3][136] , \ram[3][135] , \ram[3][134] , \ram[3][133] ,
         \ram[3][132] , \ram[3][131] , \ram[3][130] , \ram[3][129] ,
         \ram[3][128] , \ram[3][127] , \ram[3][126] , \ram[3][125] ,
         \ram[3][124] , \ram[3][123] , \ram[3][122] , \ram[3][121] ,
         \ram[3][120] , \ram[3][119] , \ram[3][118] , \ram[3][117] ,
         \ram[3][116] , \ram[3][115] , \ram[3][114] , \ram[3][113] ,
         \ram[3][112] , \ram[3][111] , \ram[3][110] , \ram[3][109] ,
         \ram[3][108] , \ram[3][107] , \ram[3][106] , \ram[3][105] ,
         \ram[3][104] , \ram[3][103] , \ram[3][102] , \ram[3][101] ,
         \ram[3][100] , \ram[3][99] , \ram[3][98] , \ram[3][97] , \ram[3][96] ,
         \ram[3][95] , \ram[3][94] , \ram[3][93] , \ram[3][92] , \ram[3][91] ,
         \ram[3][90] , \ram[3][89] , \ram[3][88] , \ram[3][87] , \ram[3][86] ,
         \ram[3][85] , \ram[3][84] , \ram[3][83] , \ram[3][82] , \ram[3][81] ,
         \ram[3][80] , \ram[3][79] , \ram[3][78] , \ram[3][77] , \ram[3][76] ,
         \ram[3][75] , \ram[3][74] , \ram[3][73] , \ram[3][72] , \ram[3][71] ,
         \ram[3][70] , \ram[3][69] , \ram[3][68] , \ram[3][67] , \ram[3][66] ,
         \ram[3][65] , \ram[3][64] , \ram[3][63] , \ram[3][62] , \ram[3][61] ,
         \ram[3][60] , \ram[3][59] , \ram[3][58] , \ram[3][57] , \ram[3][56] ,
         \ram[3][55] , \ram[3][54] , \ram[3][53] , \ram[3][52] , \ram[3][51] ,
         \ram[3][50] , \ram[3][49] , \ram[3][48] , \ram[3][47] , \ram[3][46] ,
         \ram[3][45] , \ram[3][44] , \ram[3][43] , \ram[3][42] , \ram[3][41] ,
         \ram[3][40] , \ram[3][39] , \ram[3][38] , \ram[3][37] , \ram[3][36] ,
         \ram[3][35] , \ram[3][34] , \ram[3][33] , \ram[3][32] , \ram[3][31] ,
         \ram[3][30] , \ram[3][29] , \ram[3][28] , \ram[3][27] , \ram[3][26] ,
         \ram[3][25] , \ram[3][24] , \ram[3][23] , \ram[3][22] , \ram[3][21] ,
         \ram[3][20] , \ram[3][19] , \ram[3][18] , \ram[3][17] , \ram[3][16] ,
         \ram[3][15] , \ram[3][14] , \ram[3][13] , \ram[3][12] , \ram[3][11] ,
         \ram[3][10] , \ram[3][9] , \ram[3][8] , \ram[3][7] , \ram[3][6] ,
         \ram[3][5] , \ram[3][4] , \ram[3][3] , \ram[3][2] , \ram[3][1] ,
         \ram[3][0] , \ram[2][255] , \ram[2][254] , \ram[2][253] ,
         \ram[2][252] , \ram[2][251] , \ram[2][250] , \ram[2][249] ,
         \ram[2][248] , \ram[2][247] , \ram[2][246] , \ram[2][245] ,
         \ram[2][244] , \ram[2][243] , \ram[2][242] , \ram[2][241] ,
         \ram[2][240] , \ram[2][239] , \ram[2][238] , \ram[2][237] ,
         \ram[2][236] , \ram[2][235] , \ram[2][234] , \ram[2][233] ,
         \ram[2][232] , \ram[2][231] , \ram[2][230] , \ram[2][229] ,
         \ram[2][228] , \ram[2][227] , \ram[2][226] , \ram[2][225] ,
         \ram[2][224] , \ram[2][223] , \ram[2][222] , \ram[2][221] ,
         \ram[2][220] , \ram[2][219] , \ram[2][218] , \ram[2][217] ,
         \ram[2][216] , \ram[2][215] , \ram[2][214] , \ram[2][213] ,
         \ram[2][212] , \ram[2][211] , \ram[2][210] , \ram[2][209] ,
         \ram[2][208] , \ram[2][207] , \ram[2][206] , \ram[2][205] ,
         \ram[2][204] , \ram[2][203] , \ram[2][202] , \ram[2][201] ,
         \ram[2][200] , \ram[2][199] , \ram[2][198] , \ram[2][197] ,
         \ram[2][196] , \ram[2][195] , \ram[2][194] , \ram[2][193] ,
         \ram[2][192] , \ram[2][191] , \ram[2][190] , \ram[2][189] ,
         \ram[2][188] , \ram[2][187] , \ram[2][186] , \ram[2][185] ,
         \ram[2][184] , \ram[2][183] , \ram[2][182] , \ram[2][181] ,
         \ram[2][180] , \ram[2][179] , \ram[2][178] , \ram[2][177] ,
         \ram[2][176] , \ram[2][175] , \ram[2][174] , \ram[2][173] ,
         \ram[2][172] , \ram[2][171] , \ram[2][170] , \ram[2][169] ,
         \ram[2][168] , \ram[2][167] , \ram[2][166] , \ram[2][165] ,
         \ram[2][164] , \ram[2][163] , \ram[2][162] , \ram[2][161] ,
         \ram[2][160] , \ram[2][159] , \ram[2][158] , \ram[2][157] ,
         \ram[2][156] , \ram[2][155] , \ram[2][154] , \ram[2][153] ,
         \ram[2][152] , \ram[2][151] , \ram[2][150] , \ram[2][149] ,
         \ram[2][148] , \ram[2][147] , \ram[2][146] , \ram[2][145] ,
         \ram[2][144] , \ram[2][143] , \ram[2][142] , \ram[2][141] ,
         \ram[2][140] , \ram[2][139] , \ram[2][138] , \ram[2][137] ,
         \ram[2][136] , \ram[2][135] , \ram[2][134] , \ram[2][133] ,
         \ram[2][132] , \ram[2][131] , \ram[2][130] , \ram[2][129] ,
         \ram[2][128] , \ram[2][127] , \ram[2][126] , \ram[2][125] ,
         \ram[2][124] , \ram[2][123] , \ram[2][122] , \ram[2][121] ,
         \ram[2][120] , \ram[2][119] , \ram[2][118] , \ram[2][117] ,
         \ram[2][116] , \ram[2][115] , \ram[2][114] , \ram[2][113] ,
         \ram[2][112] , \ram[2][111] , \ram[2][110] , \ram[2][109] ,
         \ram[2][108] , \ram[2][107] , \ram[2][106] , \ram[2][105] ,
         \ram[2][104] , \ram[2][103] , \ram[2][102] , \ram[2][101] ,
         \ram[2][100] , \ram[2][99] , \ram[2][98] , \ram[2][97] , \ram[2][96] ,
         \ram[2][95] , \ram[2][94] , \ram[2][93] , \ram[2][92] , \ram[2][91] ,
         \ram[2][90] , \ram[2][89] , \ram[2][88] , \ram[2][87] , \ram[2][86] ,
         \ram[2][85] , \ram[2][84] , \ram[2][83] , \ram[2][82] , \ram[2][81] ,
         \ram[2][80] , \ram[2][79] , \ram[2][78] , \ram[2][77] , \ram[2][76] ,
         \ram[2][75] , \ram[2][74] , \ram[2][73] , \ram[2][72] , \ram[2][71] ,
         \ram[2][70] , \ram[2][69] , \ram[2][68] , \ram[2][67] , \ram[2][66] ,
         \ram[2][65] , \ram[2][64] , \ram[2][63] , \ram[2][62] , \ram[2][61] ,
         \ram[2][60] , \ram[2][59] , \ram[2][58] , \ram[2][57] , \ram[2][56] ,
         \ram[2][55] , \ram[2][54] , \ram[2][53] , \ram[2][52] , \ram[2][51] ,
         \ram[2][50] , \ram[2][49] , \ram[2][48] , \ram[2][47] , \ram[2][46] ,
         \ram[2][45] , \ram[2][44] , \ram[2][43] , \ram[2][42] , \ram[2][41] ,
         \ram[2][40] , \ram[2][39] , \ram[2][38] , \ram[2][37] , \ram[2][36] ,
         \ram[2][35] , \ram[2][34] , \ram[2][33] , \ram[2][32] , \ram[2][31] ,
         \ram[2][30] , \ram[2][29] , \ram[2][28] , \ram[2][27] , \ram[2][26] ,
         \ram[2][25] , \ram[2][24] , \ram[2][23] , \ram[2][22] , \ram[2][21] ,
         \ram[2][20] , \ram[2][19] , \ram[2][18] , \ram[2][17] , \ram[2][16] ,
         \ram[2][15] , \ram[2][14] , \ram[2][13] , \ram[2][12] , \ram[2][11] ,
         \ram[2][10] , \ram[2][9] , \ram[2][8] , \ram[2][7] , \ram[2][6] ,
         \ram[2][5] , \ram[2][4] , \ram[2][3] , \ram[2][2] , \ram[2][1] ,
         \ram[2][0] , \ram[1][255] , \ram[1][254] , \ram[1][253] ,
         \ram[1][252] , \ram[1][251] , \ram[1][250] , \ram[1][249] ,
         \ram[1][248] , \ram[1][247] , \ram[1][246] , \ram[1][245] ,
         \ram[1][244] , \ram[1][243] , \ram[1][242] , \ram[1][241] ,
         \ram[1][240] , \ram[1][239] , \ram[1][238] , \ram[1][237] ,
         \ram[1][236] , \ram[1][235] , \ram[1][234] , \ram[1][233] ,
         \ram[1][232] , \ram[1][231] , \ram[1][230] , \ram[1][229] ,
         \ram[1][228] , \ram[1][227] , \ram[1][226] , \ram[1][225] ,
         \ram[1][224] , \ram[1][223] , \ram[1][222] , \ram[1][221] ,
         \ram[1][220] , \ram[1][219] , \ram[1][218] , \ram[1][217] ,
         \ram[1][216] , \ram[1][215] , \ram[1][214] , \ram[1][213] ,
         \ram[1][212] , \ram[1][211] , \ram[1][210] , \ram[1][209] ,
         \ram[1][208] , \ram[1][207] , \ram[1][206] , \ram[1][205] ,
         \ram[1][204] , \ram[1][203] , \ram[1][202] , \ram[1][201] ,
         \ram[1][200] , \ram[1][199] , \ram[1][198] , \ram[1][197] ,
         \ram[1][196] , \ram[1][195] , \ram[1][194] , \ram[1][193] ,
         \ram[1][192] , \ram[1][191] , \ram[1][190] , \ram[1][189] ,
         \ram[1][188] , \ram[1][187] , \ram[1][186] , \ram[1][185] ,
         \ram[1][184] , \ram[1][183] , \ram[1][182] , \ram[1][181] ,
         \ram[1][180] , \ram[1][179] , \ram[1][178] , \ram[1][177] ,
         \ram[1][176] , \ram[1][175] , \ram[1][174] , \ram[1][173] ,
         \ram[1][172] , \ram[1][171] , \ram[1][170] , \ram[1][169] ,
         \ram[1][168] , \ram[1][167] , \ram[1][166] , \ram[1][165] ,
         \ram[1][164] , \ram[1][163] , \ram[1][162] , \ram[1][161] ,
         \ram[1][160] , \ram[1][159] , \ram[1][158] , \ram[1][157] ,
         \ram[1][156] , \ram[1][155] , \ram[1][154] , \ram[1][153] ,
         \ram[1][152] , \ram[1][151] , \ram[1][150] , \ram[1][149] ,
         \ram[1][148] , \ram[1][147] , \ram[1][146] , \ram[1][145] ,
         \ram[1][144] , \ram[1][143] , \ram[1][142] , \ram[1][141] ,
         \ram[1][140] , \ram[1][139] , \ram[1][138] , \ram[1][137] ,
         \ram[1][136] , \ram[1][135] , \ram[1][134] , \ram[1][133] ,
         \ram[1][132] , \ram[1][131] , \ram[1][130] , \ram[1][129] ,
         \ram[1][128] , \ram[1][127] , \ram[1][126] , \ram[1][125] ,
         \ram[1][124] , \ram[1][123] , \ram[1][122] , \ram[1][121] ,
         \ram[1][120] , \ram[1][119] , \ram[1][118] , \ram[1][117] ,
         \ram[1][116] , \ram[1][115] , \ram[1][114] , \ram[1][113] ,
         \ram[1][112] , \ram[1][111] , \ram[1][110] , \ram[1][109] ,
         \ram[1][108] , \ram[1][107] , \ram[1][106] , \ram[1][105] ,
         \ram[1][104] , \ram[1][103] , \ram[1][102] , \ram[1][101] ,
         \ram[1][100] , \ram[1][99] , \ram[1][98] , \ram[1][97] , \ram[1][96] ,
         \ram[1][95] , \ram[1][94] , \ram[1][93] , \ram[1][92] , \ram[1][91] ,
         \ram[1][90] , \ram[1][89] , \ram[1][88] , \ram[1][87] , \ram[1][86] ,
         \ram[1][85] , \ram[1][84] , \ram[1][83] , \ram[1][82] , \ram[1][81] ,
         \ram[1][80] , \ram[1][79] , \ram[1][78] , \ram[1][77] , \ram[1][76] ,
         \ram[1][75] , \ram[1][74] , \ram[1][73] , \ram[1][72] , \ram[1][71] ,
         \ram[1][70] , \ram[1][69] , \ram[1][68] , \ram[1][67] , \ram[1][66] ,
         \ram[1][65] , \ram[1][64] , \ram[1][63] , \ram[1][62] , \ram[1][61] ,
         \ram[1][60] , \ram[1][59] , \ram[1][58] , \ram[1][57] , \ram[1][56] ,
         \ram[1][55] , \ram[1][54] , \ram[1][53] , \ram[1][52] , \ram[1][51] ,
         \ram[1][50] , \ram[1][49] , \ram[1][48] , \ram[1][47] , \ram[1][46] ,
         \ram[1][45] , \ram[1][44] , \ram[1][43] , \ram[1][42] , \ram[1][41] ,
         \ram[1][40] , \ram[1][39] , \ram[1][38] , \ram[1][37] , \ram[1][36] ,
         \ram[1][35] , \ram[1][34] , \ram[1][33] , \ram[1][32] , \ram[1][31] ,
         \ram[1][30] , \ram[1][29] , \ram[1][28] , \ram[1][27] , \ram[1][26] ,
         \ram[1][25] , \ram[1][24] , \ram[1][23] , \ram[1][22] , \ram[1][21] ,
         \ram[1][20] , \ram[1][19] , \ram[1][18] , \ram[1][17] , \ram[1][16] ,
         \ram[1][15] , \ram[1][14] , \ram[1][13] , \ram[1][12] , \ram[1][11] ,
         \ram[1][10] , \ram[1][9] , \ram[1][8] , \ram[1][7] , \ram[1][6] ,
         \ram[1][5] , \ram[1][4] , \ram[1][3] , \ram[1][2] , \ram[1][1] ,
         \ram[1][0] , \ram[0][255] , \ram[0][254] , \ram[0][253] ,
         \ram[0][252] , \ram[0][251] , \ram[0][250] , \ram[0][249] ,
         \ram[0][248] , \ram[0][247] , \ram[0][246] , \ram[0][245] ,
         \ram[0][244] , \ram[0][243] , \ram[0][242] , \ram[0][241] ,
         \ram[0][240] , \ram[0][239] , \ram[0][238] , \ram[0][237] ,
         \ram[0][236] , \ram[0][235] , \ram[0][234] , \ram[0][233] ,
         \ram[0][232] , \ram[0][231] , \ram[0][230] , \ram[0][229] ,
         \ram[0][228] , \ram[0][227] , \ram[0][226] , \ram[0][225] ,
         \ram[0][224] , \ram[0][223] , \ram[0][222] , \ram[0][221] ,
         \ram[0][220] , \ram[0][219] , \ram[0][218] , \ram[0][217] ,
         \ram[0][216] , \ram[0][215] , \ram[0][214] , \ram[0][213] ,
         \ram[0][212] , \ram[0][211] , \ram[0][210] , \ram[0][209] ,
         \ram[0][208] , \ram[0][207] , \ram[0][206] , \ram[0][205] ,
         \ram[0][204] , \ram[0][203] , \ram[0][202] , \ram[0][201] ,
         \ram[0][200] , \ram[0][199] , \ram[0][198] , \ram[0][197] ,
         \ram[0][196] , \ram[0][195] , \ram[0][194] , \ram[0][193] ,
         \ram[0][192] , \ram[0][191] , \ram[0][190] , \ram[0][189] ,
         \ram[0][188] , \ram[0][187] , \ram[0][186] , \ram[0][185] ,
         \ram[0][184] , \ram[0][183] , \ram[0][182] , \ram[0][181] ,
         \ram[0][180] , \ram[0][179] , \ram[0][178] , \ram[0][177] ,
         \ram[0][176] , \ram[0][175] , \ram[0][174] , \ram[0][173] ,
         \ram[0][172] , \ram[0][171] , \ram[0][170] , \ram[0][169] ,
         \ram[0][168] , \ram[0][167] , \ram[0][166] , \ram[0][165] ,
         \ram[0][164] , \ram[0][163] , \ram[0][162] , \ram[0][161] ,
         \ram[0][160] , \ram[0][159] , \ram[0][158] , \ram[0][157] ,
         \ram[0][156] , \ram[0][155] , \ram[0][154] , \ram[0][153] ,
         \ram[0][152] , \ram[0][151] , \ram[0][150] , \ram[0][149] ,
         \ram[0][148] , \ram[0][147] , \ram[0][146] , \ram[0][145] ,
         \ram[0][144] , \ram[0][143] , \ram[0][142] , \ram[0][141] ,
         \ram[0][140] , \ram[0][139] , \ram[0][138] , \ram[0][137] ,
         \ram[0][136] , \ram[0][135] , \ram[0][134] , \ram[0][133] ,
         \ram[0][132] , \ram[0][131] , \ram[0][130] , \ram[0][129] ,
         \ram[0][128] , \ram[0][127] , \ram[0][126] , \ram[0][125] ,
         \ram[0][124] , \ram[0][123] , \ram[0][122] , \ram[0][121] ,
         \ram[0][120] , \ram[0][119] , \ram[0][118] , \ram[0][117] ,
         \ram[0][116] , \ram[0][115] , \ram[0][114] , \ram[0][113] ,
         \ram[0][112] , \ram[0][111] , \ram[0][110] , \ram[0][109] ,
         \ram[0][108] , \ram[0][107] , \ram[0][106] , \ram[0][105] ,
         \ram[0][104] , \ram[0][103] , \ram[0][102] , \ram[0][101] ,
         \ram[0][100] , \ram[0][99] , \ram[0][98] , \ram[0][97] , \ram[0][96] ,
         \ram[0][95] , \ram[0][94] , \ram[0][93] , \ram[0][92] , \ram[0][91] ,
         \ram[0][90] , \ram[0][89] , \ram[0][88] , \ram[0][87] , \ram[0][86] ,
         \ram[0][85] , \ram[0][84] , \ram[0][83] , \ram[0][82] , \ram[0][81] ,
         \ram[0][80] , \ram[0][79] , \ram[0][78] , \ram[0][77] , \ram[0][76] ,
         \ram[0][75] , \ram[0][74] , \ram[0][73] , \ram[0][72] , \ram[0][71] ,
         \ram[0][70] , \ram[0][69] , \ram[0][68] , \ram[0][67] , \ram[0][66] ,
         \ram[0][65] , \ram[0][64] , \ram[0][63] , \ram[0][62] , \ram[0][61] ,
         \ram[0][60] , \ram[0][59] , \ram[0][58] , \ram[0][57] , \ram[0][56] ,
         \ram[0][55] , \ram[0][54] , \ram[0][53] , \ram[0][52] , \ram[0][51] ,
         \ram[0][50] , \ram[0][49] , \ram[0][48] , \ram[0][47] , \ram[0][46] ,
         \ram[0][45] , \ram[0][44] , \ram[0][43] , \ram[0][42] , \ram[0][41] ,
         \ram[0][40] , \ram[0][39] , \ram[0][38] , \ram[0][37] , \ram[0][36] ,
         \ram[0][35] , \ram[0][34] , \ram[0][33] , \ram[0][32] , \ram[0][31] ,
         \ram[0][30] , \ram[0][29] , \ram[0][28] , \ram[0][27] , \ram[0][26] ,
         \ram[0][25] , \ram[0][24] , \ram[0][23] , \ram[0][22] , \ram[0][21] ,
         \ram[0][20] , \ram[0][19] , \ram[0][18] , \ram[0][17] , \ram[0][16] ,
         \ram[0][15] , \ram[0][14] , \ram[0][13] , \ram[0][12] , \ram[0][11] ,
         \ram[0][10] , \ram[0][9] , \ram[0][8] , \ram[0][7] , \ram[0][6] ,
         \ram[0][5] , \ram[0][4] , \ram[0][3] , \ram[0][2] , \ram[0][1] ,
         \ram[0][0] , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412;
  assign N26 = addr[0];
  assign N27 = addr[1];
  assign N28 = addr[2];
  assign N29 = addr[3];

  DFFX1_HVT \ram_reg[15][255]  ( .D(n4156), .CLK(clk), .Q(\ram[15][255] ) );
  DFFX1_HVT \ram_reg[15][254]  ( .D(n4155), .CLK(clk), .Q(\ram[15][254] ) );
  DFFX1_HVT \ram_reg[15][253]  ( .D(n4154), .CLK(clk), .Q(\ram[15][253] ) );
  DFFX1_HVT \ram_reg[15][252]  ( .D(n4153), .CLK(clk), .Q(\ram[15][252] ) );
  DFFX1_HVT \ram_reg[15][251]  ( .D(n4152), .CLK(clk), .Q(\ram[15][251] ) );
  DFFX1_HVT \ram_reg[15][250]  ( .D(n4151), .CLK(clk), .Q(\ram[15][250] ) );
  DFFX1_HVT \ram_reg[15][249]  ( .D(n4150), .CLK(clk), .Q(\ram[15][249] ) );
  DFFX1_HVT \ram_reg[15][248]  ( .D(n4149), .CLK(clk), .Q(\ram[15][248] ) );
  DFFX1_HVT \ram_reg[15][247]  ( .D(n4148), .CLK(clk), .Q(\ram[15][247] ) );
  DFFX1_HVT \ram_reg[15][246]  ( .D(n4147), .CLK(clk), .Q(\ram[15][246] ) );
  DFFX1_HVT \ram_reg[15][245]  ( .D(n4146), .CLK(clk), .Q(\ram[15][245] ) );
  DFFX1_HVT \ram_reg[15][244]  ( .D(n4145), .CLK(clk), .Q(\ram[15][244] ) );
  DFFX1_HVT \ram_reg[15][243]  ( .D(n4144), .CLK(clk), .Q(\ram[15][243] ) );
  DFFX1_HVT \ram_reg[15][242]  ( .D(n4143), .CLK(clk), .Q(\ram[15][242] ) );
  DFFX1_HVT \ram_reg[15][241]  ( .D(n4142), .CLK(clk), .Q(\ram[15][241] ) );
  DFFX1_HVT \ram_reg[15][240]  ( .D(n4141), .CLK(clk), .Q(\ram[15][240] ) );
  DFFX1_HVT \ram_reg[15][239]  ( .D(n4140), .CLK(clk), .Q(\ram[15][239] ) );
  DFFX1_HVT \ram_reg[15][238]  ( .D(n4139), .CLK(clk), .Q(\ram[15][238] ) );
  DFFX1_HVT \ram_reg[15][237]  ( .D(n4138), .CLK(clk), .Q(\ram[15][237] ) );
  DFFX1_HVT \ram_reg[15][236]  ( .D(n4137), .CLK(clk), .Q(\ram[15][236] ) );
  DFFX1_HVT \ram_reg[15][235]  ( .D(n4136), .CLK(clk), .Q(\ram[15][235] ) );
  DFFX1_HVT \ram_reg[15][234]  ( .D(n4135), .CLK(clk), .Q(\ram[15][234] ) );
  DFFX1_HVT \ram_reg[15][233]  ( .D(n4134), .CLK(clk), .Q(\ram[15][233] ) );
  DFFX1_HVT \ram_reg[15][232]  ( .D(n4133), .CLK(clk), .Q(\ram[15][232] ) );
  DFFX1_HVT \ram_reg[15][231]  ( .D(n4132), .CLK(clk), .Q(\ram[15][231] ) );
  DFFX1_HVT \ram_reg[15][230]  ( .D(n4131), .CLK(clk), .Q(\ram[15][230] ) );
  DFFX1_HVT \ram_reg[15][229]  ( .D(n4130), .CLK(clk), .Q(\ram[15][229] ) );
  DFFX1_HVT \ram_reg[15][228]  ( .D(n4129), .CLK(clk), .Q(\ram[15][228] ) );
  DFFX1_HVT \ram_reg[15][227]  ( .D(n4128), .CLK(clk), .Q(\ram[15][227] ) );
  DFFX1_HVT \ram_reg[15][226]  ( .D(n4127), .CLK(clk), .Q(\ram[15][226] ) );
  DFFX1_HVT \ram_reg[15][225]  ( .D(n4126), .CLK(clk), .Q(\ram[15][225] ) );
  DFFX1_HVT \ram_reg[15][224]  ( .D(n4125), .CLK(clk), .Q(\ram[15][224] ) );
  DFFX1_HVT \ram_reg[15][223]  ( .D(n4124), .CLK(clk), .Q(\ram[15][223] ) );
  DFFX1_HVT \ram_reg[15][222]  ( .D(n4123), .CLK(clk), .Q(\ram[15][222] ) );
  DFFX1_HVT \ram_reg[15][221]  ( .D(n4122), .CLK(clk), .Q(\ram[15][221] ) );
  DFFX1_HVT \ram_reg[15][220]  ( .D(n4121), .CLK(clk), .Q(\ram[15][220] ) );
  DFFX1_HVT \ram_reg[15][219]  ( .D(n4120), .CLK(clk), .Q(\ram[15][219] ) );
  DFFX1_HVT \ram_reg[15][218]  ( .D(n4119), .CLK(clk), .Q(\ram[15][218] ) );
  DFFX1_HVT \ram_reg[15][217]  ( .D(n4118), .CLK(clk), .Q(\ram[15][217] ) );
  DFFX1_HVT \ram_reg[15][216]  ( .D(n4117), .CLK(clk), .Q(\ram[15][216] ) );
  DFFX1_HVT \ram_reg[15][215]  ( .D(n4116), .CLK(clk), .Q(\ram[15][215] ) );
  DFFX1_HVT \ram_reg[15][214]  ( .D(n4115), .CLK(clk), .Q(\ram[15][214] ) );
  DFFX1_HVT \ram_reg[15][213]  ( .D(n4114), .CLK(clk), .Q(\ram[15][213] ) );
  DFFX1_HVT \ram_reg[15][212]  ( .D(n4113), .CLK(clk), .Q(\ram[15][212] ) );
  DFFX1_HVT \ram_reg[15][211]  ( .D(n4112), .CLK(clk), .Q(\ram[15][211] ) );
  DFFX1_HVT \ram_reg[15][210]  ( .D(n4111), .CLK(clk), .Q(\ram[15][210] ) );
  DFFX1_HVT \ram_reg[15][209]  ( .D(n4110), .CLK(clk), .Q(\ram[15][209] ) );
  DFFX1_HVT \ram_reg[15][208]  ( .D(n4109), .CLK(clk), .Q(\ram[15][208] ) );
  DFFX1_HVT \ram_reg[15][207]  ( .D(n4108), .CLK(clk), .Q(\ram[15][207] ) );
  DFFX1_HVT \ram_reg[15][206]  ( .D(n4107), .CLK(clk), .Q(\ram[15][206] ) );
  DFFX1_HVT \ram_reg[15][205]  ( .D(n4106), .CLK(clk), .Q(\ram[15][205] ) );
  DFFX1_HVT \ram_reg[15][204]  ( .D(n4105), .CLK(clk), .Q(\ram[15][204] ) );
  DFFX1_HVT \ram_reg[15][203]  ( .D(n4104), .CLK(clk), .Q(\ram[15][203] ) );
  DFFX1_HVT \ram_reg[15][202]  ( .D(n4103), .CLK(clk), .Q(\ram[15][202] ) );
  DFFX1_HVT \ram_reg[15][201]  ( .D(n4102), .CLK(clk), .Q(\ram[15][201] ) );
  DFFX1_HVT \ram_reg[15][200]  ( .D(n4101), .CLK(clk), .Q(\ram[15][200] ) );
  DFFX1_HVT \ram_reg[15][199]  ( .D(n4100), .CLK(clk), .Q(\ram[15][199] ) );
  DFFX1_HVT \ram_reg[15][198]  ( .D(n4099), .CLK(clk), .Q(\ram[15][198] ) );
  DFFX1_HVT \ram_reg[15][197]  ( .D(n4098), .CLK(clk), .Q(\ram[15][197] ) );
  DFFX1_HVT \ram_reg[15][196]  ( .D(n4097), .CLK(clk), .Q(\ram[15][196] ) );
  DFFX1_HVT \ram_reg[15][195]  ( .D(n4096), .CLK(clk), .Q(\ram[15][195] ) );
  DFFX1_HVT \ram_reg[15][194]  ( .D(n4095), .CLK(clk), .Q(\ram[15][194] ) );
  DFFX1_HVT \ram_reg[15][193]  ( .D(n4094), .CLK(clk), .Q(\ram[15][193] ) );
  DFFX1_HVT \ram_reg[15][192]  ( .D(n4093), .CLK(clk), .Q(\ram[15][192] ) );
  DFFX1_HVT \ram_reg[15][191]  ( .D(n4092), .CLK(clk), .Q(\ram[15][191] ) );
  DFFX1_HVT \ram_reg[15][190]  ( .D(n4091), .CLK(clk), .Q(\ram[15][190] ) );
  DFFX1_HVT \ram_reg[15][189]  ( .D(n4090), .CLK(clk), .Q(\ram[15][189] ) );
  DFFX1_HVT \ram_reg[15][188]  ( .D(n4089), .CLK(clk), .Q(\ram[15][188] ) );
  DFFX1_HVT \ram_reg[15][187]  ( .D(n4088), .CLK(clk), .Q(\ram[15][187] ) );
  DFFX1_HVT \ram_reg[15][186]  ( .D(n4087), .CLK(clk), .Q(\ram[15][186] ) );
  DFFX1_HVT \ram_reg[15][185]  ( .D(n4086), .CLK(clk), .Q(\ram[15][185] ) );
  DFFX1_HVT \ram_reg[15][184]  ( .D(n4085), .CLK(clk), .Q(\ram[15][184] ) );
  DFFX1_HVT \ram_reg[15][183]  ( .D(n4084), .CLK(clk), .Q(\ram[15][183] ) );
  DFFX1_HVT \ram_reg[15][182]  ( .D(n4083), .CLK(clk), .Q(\ram[15][182] ) );
  DFFX1_HVT \ram_reg[15][181]  ( .D(n4082), .CLK(clk), .Q(\ram[15][181] ) );
  DFFX1_HVT \ram_reg[15][180]  ( .D(n4081), .CLK(clk), .Q(\ram[15][180] ) );
  DFFX1_HVT \ram_reg[15][179]  ( .D(n4080), .CLK(clk), .Q(\ram[15][179] ) );
  DFFX1_HVT \ram_reg[15][178]  ( .D(n4079), .CLK(clk), .Q(\ram[15][178] ) );
  DFFX1_HVT \ram_reg[15][177]  ( .D(n4078), .CLK(clk), .Q(\ram[15][177] ) );
  DFFX1_HVT \ram_reg[15][176]  ( .D(n4077), .CLK(clk), .Q(\ram[15][176] ) );
  DFFX1_HVT \ram_reg[15][175]  ( .D(n4076), .CLK(clk), .Q(\ram[15][175] ) );
  DFFX1_HVT \ram_reg[15][174]  ( .D(n4075), .CLK(clk), .Q(\ram[15][174] ) );
  DFFX1_HVT \ram_reg[15][173]  ( .D(n4074), .CLK(clk), .Q(\ram[15][173] ) );
  DFFX1_HVT \ram_reg[15][172]  ( .D(n4073), .CLK(clk), .Q(\ram[15][172] ) );
  DFFX1_HVT \ram_reg[15][171]  ( .D(n4072), .CLK(clk), .Q(\ram[15][171] ) );
  DFFX1_HVT \ram_reg[15][170]  ( .D(n4071), .CLK(clk), .Q(\ram[15][170] ) );
  DFFX1_HVT \ram_reg[15][169]  ( .D(n4070), .CLK(clk), .Q(\ram[15][169] ) );
  DFFX1_HVT \ram_reg[15][168]  ( .D(n4069), .CLK(clk), .Q(\ram[15][168] ) );
  DFFX1_HVT \ram_reg[15][167]  ( .D(n4068), .CLK(clk), .Q(\ram[15][167] ) );
  DFFX1_HVT \ram_reg[15][166]  ( .D(n4067), .CLK(clk), .Q(\ram[15][166] ) );
  DFFX1_HVT \ram_reg[15][165]  ( .D(n4066), .CLK(clk), .Q(\ram[15][165] ) );
  DFFX1_HVT \ram_reg[15][164]  ( .D(n4065), .CLK(clk), .Q(\ram[15][164] ) );
  DFFX1_HVT \ram_reg[15][163]  ( .D(n4064), .CLK(clk), .Q(\ram[15][163] ) );
  DFFX1_HVT \ram_reg[15][162]  ( .D(n4063), .CLK(clk), .Q(\ram[15][162] ) );
  DFFX1_HVT \ram_reg[15][161]  ( .D(n4062), .CLK(clk), .Q(\ram[15][161] ) );
  DFFX1_HVT \ram_reg[15][160]  ( .D(n4061), .CLK(clk), .Q(\ram[15][160] ) );
  DFFX1_HVT \ram_reg[15][159]  ( .D(n4060), .CLK(clk), .Q(\ram[15][159] ) );
  DFFX1_HVT \ram_reg[15][158]  ( .D(n4059), .CLK(clk), .Q(\ram[15][158] ) );
  DFFX1_HVT \ram_reg[15][157]  ( .D(n4058), .CLK(clk), .Q(\ram[15][157] ) );
  DFFX1_HVT \ram_reg[15][156]  ( .D(n4057), .CLK(clk), .Q(\ram[15][156] ) );
  DFFX1_HVT \ram_reg[15][155]  ( .D(n4056), .CLK(clk), .Q(\ram[15][155] ) );
  DFFX1_HVT \ram_reg[15][154]  ( .D(n4055), .CLK(clk), .Q(\ram[15][154] ) );
  DFFX1_HVT \ram_reg[15][153]  ( .D(n4054), .CLK(clk), .Q(\ram[15][153] ) );
  DFFX1_HVT \ram_reg[15][152]  ( .D(n4053), .CLK(clk), .Q(\ram[15][152] ) );
  DFFX1_HVT \ram_reg[15][151]  ( .D(n4052), .CLK(clk), .Q(\ram[15][151] ) );
  DFFX1_HVT \ram_reg[15][150]  ( .D(n4051), .CLK(clk), .Q(\ram[15][150] ) );
  DFFX1_HVT \ram_reg[15][149]  ( .D(n4050), .CLK(clk), .Q(\ram[15][149] ) );
  DFFX1_HVT \ram_reg[15][148]  ( .D(n4049), .CLK(clk), .Q(\ram[15][148] ) );
  DFFX1_HVT \ram_reg[15][147]  ( .D(n4048), .CLK(clk), .Q(\ram[15][147] ) );
  DFFX1_HVT \ram_reg[15][146]  ( .D(n4047), .CLK(clk), .Q(\ram[15][146] ) );
  DFFX1_HVT \ram_reg[15][145]  ( .D(n4046), .CLK(clk), .Q(\ram[15][145] ) );
  DFFX1_HVT \ram_reg[15][144]  ( .D(n4045), .CLK(clk), .Q(\ram[15][144] ) );
  DFFX1_HVT \ram_reg[15][143]  ( .D(n4044), .CLK(clk), .Q(\ram[15][143] ) );
  DFFX1_HVT \ram_reg[15][142]  ( .D(n4043), .CLK(clk), .Q(\ram[15][142] ) );
  DFFX1_HVT \ram_reg[15][141]  ( .D(n4042), .CLK(clk), .Q(\ram[15][141] ) );
  DFFX1_HVT \ram_reg[15][140]  ( .D(n4041), .CLK(clk), .Q(\ram[15][140] ) );
  DFFX1_HVT \ram_reg[15][139]  ( .D(n4040), .CLK(clk), .Q(\ram[15][139] ) );
  DFFX1_HVT \ram_reg[15][138]  ( .D(n4039), .CLK(clk), .Q(\ram[15][138] ) );
  DFFX1_HVT \ram_reg[15][137]  ( .D(n4038), .CLK(clk), .Q(\ram[15][137] ) );
  DFFX1_HVT \ram_reg[15][136]  ( .D(n4037), .CLK(clk), .Q(\ram[15][136] ) );
  DFFX1_HVT \ram_reg[15][135]  ( .D(n4036), .CLK(clk), .Q(\ram[15][135] ) );
  DFFX1_HVT \ram_reg[15][134]  ( .D(n4035), .CLK(clk), .Q(\ram[15][134] ) );
  DFFX1_HVT \ram_reg[15][133]  ( .D(n4034), .CLK(clk), .Q(\ram[15][133] ) );
  DFFX1_HVT \ram_reg[15][132]  ( .D(n4033), .CLK(clk), .Q(\ram[15][132] ) );
  DFFX1_HVT \ram_reg[15][131]  ( .D(n4032), .CLK(clk), .Q(\ram[15][131] ) );
  DFFX1_HVT \ram_reg[15][130]  ( .D(n4031), .CLK(clk), .Q(\ram[15][130] ) );
  DFFX1_HVT \ram_reg[15][129]  ( .D(n4030), .CLK(clk), .Q(\ram[15][129] ) );
  DFFX1_HVT \ram_reg[15][128]  ( .D(n4029), .CLK(clk), .Q(\ram[15][128] ) );
  DFFX1_HVT \ram_reg[15][127]  ( .D(n4028), .CLK(clk), .Q(\ram[15][127] ) );
  DFFX1_HVT \ram_reg[15][126]  ( .D(n4027), .CLK(clk), .Q(\ram[15][126] ) );
  DFFX1_HVT \ram_reg[15][125]  ( .D(n4026), .CLK(clk), .Q(\ram[15][125] ) );
  DFFX1_HVT \ram_reg[15][124]  ( .D(n4025), .CLK(clk), .Q(\ram[15][124] ) );
  DFFX1_HVT \ram_reg[15][123]  ( .D(n4024), .CLK(clk), .Q(\ram[15][123] ) );
  DFFX1_HVT \ram_reg[15][122]  ( .D(n4023), .CLK(clk), .Q(\ram[15][122] ) );
  DFFX1_HVT \ram_reg[15][121]  ( .D(n4022), .CLK(clk), .Q(\ram[15][121] ) );
  DFFX1_HVT \ram_reg[15][120]  ( .D(n4021), .CLK(clk), .Q(\ram[15][120] ) );
  DFFX1_HVT \ram_reg[15][119]  ( .D(n4020), .CLK(clk), .Q(\ram[15][119] ) );
  DFFX1_HVT \ram_reg[15][118]  ( .D(n4019), .CLK(clk), .Q(\ram[15][118] ) );
  DFFX1_HVT \ram_reg[15][117]  ( .D(n4018), .CLK(clk), .Q(\ram[15][117] ) );
  DFFX1_HVT \ram_reg[15][116]  ( .D(n4017), .CLK(clk), .Q(\ram[15][116] ) );
  DFFX1_HVT \ram_reg[15][115]  ( .D(n4016), .CLK(clk), .Q(\ram[15][115] ) );
  DFFX1_HVT \ram_reg[15][114]  ( .D(n4015), .CLK(clk), .Q(\ram[15][114] ) );
  DFFX1_HVT \ram_reg[15][113]  ( .D(n4014), .CLK(clk), .Q(\ram[15][113] ) );
  DFFX1_HVT \ram_reg[15][112]  ( .D(n4013), .CLK(clk), .Q(\ram[15][112] ) );
  DFFX1_HVT \ram_reg[15][111]  ( .D(n4012), .CLK(clk), .Q(\ram[15][111] ) );
  DFFX1_HVT \ram_reg[15][110]  ( .D(n4011), .CLK(clk), .Q(\ram[15][110] ) );
  DFFX1_HVT \ram_reg[15][109]  ( .D(n4010), .CLK(clk), .Q(\ram[15][109] ) );
  DFFX1_HVT \ram_reg[15][108]  ( .D(n4009), .CLK(clk), .Q(\ram[15][108] ) );
  DFFX1_HVT \ram_reg[15][107]  ( .D(n4008), .CLK(clk), .Q(\ram[15][107] ) );
  DFFX1_HVT \ram_reg[15][106]  ( .D(n4007), .CLK(clk), .Q(\ram[15][106] ) );
  DFFX1_HVT \ram_reg[15][105]  ( .D(n4006), .CLK(clk), .Q(\ram[15][105] ) );
  DFFX1_HVT \ram_reg[15][104]  ( .D(n4005), .CLK(clk), .Q(\ram[15][104] ) );
  DFFX1_HVT \ram_reg[15][103]  ( .D(n4004), .CLK(clk), .Q(\ram[15][103] ) );
  DFFX1_HVT \ram_reg[15][102]  ( .D(n4003), .CLK(clk), .Q(\ram[15][102] ) );
  DFFX1_HVT \ram_reg[15][101]  ( .D(n4002), .CLK(clk), .Q(\ram[15][101] ) );
  DFFX1_HVT \ram_reg[15][100]  ( .D(n4001), .CLK(clk), .Q(\ram[15][100] ) );
  DFFX1_HVT \ram_reg[15][99]  ( .D(n4000), .CLK(clk), .Q(\ram[15][99] ) );
  DFFX1_HVT \ram_reg[15][98]  ( .D(n3999), .CLK(clk), .Q(\ram[15][98] ) );
  DFFX1_HVT \ram_reg[15][97]  ( .D(n3998), .CLK(clk), .Q(\ram[15][97] ) );
  DFFX1_HVT \ram_reg[15][96]  ( .D(n3997), .CLK(clk), .Q(\ram[15][96] ) );
  DFFX1_HVT \ram_reg[15][95]  ( .D(n3996), .CLK(clk), .Q(\ram[15][95] ) );
  DFFX1_HVT \ram_reg[15][94]  ( .D(n3995), .CLK(clk), .Q(\ram[15][94] ) );
  DFFX1_HVT \ram_reg[15][93]  ( .D(n3994), .CLK(clk), .Q(\ram[15][93] ) );
  DFFX1_HVT \ram_reg[15][92]  ( .D(n3993), .CLK(clk), .Q(\ram[15][92] ) );
  DFFX1_HVT \ram_reg[15][91]  ( .D(n3992), .CLK(clk), .Q(\ram[15][91] ) );
  DFFX1_HVT \ram_reg[15][90]  ( .D(n3991), .CLK(clk), .Q(\ram[15][90] ) );
  DFFX1_HVT \ram_reg[15][89]  ( .D(n3990), .CLK(clk), .Q(\ram[15][89] ) );
  DFFX1_HVT \ram_reg[15][88]  ( .D(n3989), .CLK(clk), .Q(\ram[15][88] ) );
  DFFX1_HVT \ram_reg[15][87]  ( .D(n3988), .CLK(clk), .Q(\ram[15][87] ) );
  DFFX1_HVT \ram_reg[15][86]  ( .D(n3987), .CLK(clk), .Q(\ram[15][86] ) );
  DFFX1_HVT \ram_reg[15][85]  ( .D(n3986), .CLK(clk), .Q(\ram[15][85] ) );
  DFFX1_HVT \ram_reg[15][84]  ( .D(n3985), .CLK(clk), .Q(\ram[15][84] ) );
  DFFX1_HVT \ram_reg[15][83]  ( .D(n3984), .CLK(clk), .Q(\ram[15][83] ) );
  DFFX1_HVT \ram_reg[15][82]  ( .D(n3983), .CLK(clk), .Q(\ram[15][82] ) );
  DFFX1_HVT \ram_reg[15][81]  ( .D(n3982), .CLK(clk), .Q(\ram[15][81] ) );
  DFFX1_HVT \ram_reg[15][80]  ( .D(n3981), .CLK(clk), .Q(\ram[15][80] ) );
  DFFX1_HVT \ram_reg[15][79]  ( .D(n3980), .CLK(clk), .Q(\ram[15][79] ) );
  DFFX1_HVT \ram_reg[15][78]  ( .D(n3979), .CLK(clk), .Q(\ram[15][78] ) );
  DFFX1_HVT \ram_reg[15][77]  ( .D(n3978), .CLK(clk), .Q(\ram[15][77] ) );
  DFFX1_HVT \ram_reg[15][76]  ( .D(n3977), .CLK(clk), .Q(\ram[15][76] ) );
  DFFX1_HVT \ram_reg[15][75]  ( .D(n3976), .CLK(clk), .Q(\ram[15][75] ) );
  DFFX1_HVT \ram_reg[15][74]  ( .D(n3975), .CLK(clk), .Q(\ram[15][74] ) );
  DFFX1_HVT \ram_reg[15][73]  ( .D(n3974), .CLK(clk), .Q(\ram[15][73] ) );
  DFFX1_HVT \ram_reg[15][72]  ( .D(n3973), .CLK(clk), .Q(\ram[15][72] ) );
  DFFX1_HVT \ram_reg[15][71]  ( .D(n3972), .CLK(clk), .Q(\ram[15][71] ) );
  DFFX1_HVT \ram_reg[15][70]  ( .D(n3971), .CLK(clk), .Q(\ram[15][70] ) );
  DFFX1_HVT \ram_reg[15][69]  ( .D(n3970), .CLK(clk), .Q(\ram[15][69] ) );
  DFFX1_HVT \ram_reg[15][68]  ( .D(n3969), .CLK(clk), .Q(\ram[15][68] ) );
  DFFX1_HVT \ram_reg[15][67]  ( .D(n3968), .CLK(clk), .Q(\ram[15][67] ) );
  DFFX1_HVT \ram_reg[15][66]  ( .D(n3967), .CLK(clk), .Q(\ram[15][66] ) );
  DFFX1_HVT \ram_reg[15][65]  ( .D(n3966), .CLK(clk), .Q(\ram[15][65] ) );
  DFFX1_HVT \ram_reg[15][64]  ( .D(n3965), .CLK(clk), .Q(\ram[15][64] ) );
  DFFX1_HVT \ram_reg[15][63]  ( .D(n3964), .CLK(clk), .Q(\ram[15][63] ) );
  DFFX1_HVT \ram_reg[15][62]  ( .D(n3963), .CLK(clk), .Q(\ram[15][62] ) );
  DFFX1_HVT \ram_reg[15][61]  ( .D(n3962), .CLK(clk), .Q(\ram[15][61] ) );
  DFFX1_HVT \ram_reg[15][60]  ( .D(n3961), .CLK(clk), .Q(\ram[15][60] ) );
  DFFX1_HVT \ram_reg[15][59]  ( .D(n3960), .CLK(clk), .Q(\ram[15][59] ) );
  DFFX1_HVT \ram_reg[15][58]  ( .D(n3959), .CLK(clk), .Q(\ram[15][58] ) );
  DFFX1_HVT \ram_reg[15][57]  ( .D(n3958), .CLK(clk), .Q(\ram[15][57] ) );
  DFFX1_HVT \ram_reg[15][56]  ( .D(n3957), .CLK(clk), .Q(\ram[15][56] ) );
  DFFX1_HVT \ram_reg[15][55]  ( .D(n3956), .CLK(clk), .Q(\ram[15][55] ) );
  DFFX1_HVT \ram_reg[15][54]  ( .D(n3955), .CLK(clk), .Q(\ram[15][54] ) );
  DFFX1_HVT \ram_reg[15][53]  ( .D(n3954), .CLK(clk), .Q(\ram[15][53] ) );
  DFFX1_HVT \ram_reg[15][52]  ( .D(n3953), .CLK(clk), .Q(\ram[15][52] ) );
  DFFX1_HVT \ram_reg[15][51]  ( .D(n3952), .CLK(clk), .Q(\ram[15][51] ) );
  DFFX1_HVT \ram_reg[15][50]  ( .D(n3951), .CLK(clk), .Q(\ram[15][50] ) );
  DFFX1_HVT \ram_reg[15][49]  ( .D(n3950), .CLK(clk), .Q(\ram[15][49] ) );
  DFFX1_HVT \ram_reg[15][48]  ( .D(n3949), .CLK(clk), .Q(\ram[15][48] ) );
  DFFX1_HVT \ram_reg[15][47]  ( .D(n3948), .CLK(clk), .Q(\ram[15][47] ) );
  DFFX1_HVT \ram_reg[15][46]  ( .D(n3947), .CLK(clk), .Q(\ram[15][46] ) );
  DFFX1_HVT \ram_reg[15][45]  ( .D(n3946), .CLK(clk), .Q(\ram[15][45] ) );
  DFFX1_HVT \ram_reg[15][44]  ( .D(n3945), .CLK(clk), .Q(\ram[15][44] ) );
  DFFX1_HVT \ram_reg[15][43]  ( .D(n3944), .CLK(clk), .Q(\ram[15][43] ) );
  DFFX1_HVT \ram_reg[15][42]  ( .D(n3943), .CLK(clk), .Q(\ram[15][42] ) );
  DFFX1_HVT \ram_reg[15][41]  ( .D(n3942), .CLK(clk), .Q(\ram[15][41] ) );
  DFFX1_HVT \ram_reg[15][40]  ( .D(n3941), .CLK(clk), .Q(\ram[15][40] ) );
  DFFX1_HVT \ram_reg[15][39]  ( .D(n3940), .CLK(clk), .Q(\ram[15][39] ) );
  DFFX1_HVT \ram_reg[15][38]  ( .D(n3939), .CLK(clk), .Q(\ram[15][38] ) );
  DFFX1_HVT \ram_reg[15][37]  ( .D(n3938), .CLK(clk), .Q(\ram[15][37] ) );
  DFFX1_HVT \ram_reg[15][36]  ( .D(n3937), .CLK(clk), .Q(\ram[15][36] ) );
  DFFX1_HVT \ram_reg[15][35]  ( .D(n3936), .CLK(clk), .Q(\ram[15][35] ) );
  DFFX1_HVT \ram_reg[15][34]  ( .D(n3935), .CLK(clk), .Q(\ram[15][34] ) );
  DFFX1_HVT \ram_reg[15][33]  ( .D(n3934), .CLK(clk), .Q(\ram[15][33] ) );
  DFFX1_HVT \ram_reg[15][32]  ( .D(n3933), .CLK(clk), .Q(\ram[15][32] ) );
  DFFX1_HVT \ram_reg[15][31]  ( .D(n3932), .CLK(clk), .Q(\ram[15][31] ) );
  DFFX1_HVT \ram_reg[15][30]  ( .D(n3931), .CLK(clk), .Q(\ram[15][30] ) );
  DFFX1_HVT \ram_reg[15][29]  ( .D(n3930), .CLK(clk), .Q(\ram[15][29] ) );
  DFFX1_HVT \ram_reg[15][28]  ( .D(n3929), .CLK(clk), .Q(\ram[15][28] ) );
  DFFX1_HVT \ram_reg[15][27]  ( .D(n3928), .CLK(clk), .Q(\ram[15][27] ) );
  DFFX1_HVT \ram_reg[15][26]  ( .D(n3927), .CLK(clk), .Q(\ram[15][26] ) );
  DFFX1_HVT \ram_reg[15][25]  ( .D(n3926), .CLK(clk), .Q(\ram[15][25] ) );
  DFFX1_HVT \ram_reg[15][24]  ( .D(n3925), .CLK(clk), .Q(\ram[15][24] ) );
  DFFX1_HVT \ram_reg[15][23]  ( .D(n3924), .CLK(clk), .Q(\ram[15][23] ) );
  DFFX1_HVT \ram_reg[15][22]  ( .D(n3923), .CLK(clk), .Q(\ram[15][22] ) );
  DFFX1_HVT \ram_reg[15][21]  ( .D(n3922), .CLK(clk), .Q(\ram[15][21] ) );
  DFFX1_HVT \ram_reg[15][20]  ( .D(n3921), .CLK(clk), .Q(\ram[15][20] ) );
  DFFX1_HVT \ram_reg[15][19]  ( .D(n3920), .CLK(clk), .Q(\ram[15][19] ) );
  DFFX1_HVT \ram_reg[15][18]  ( .D(n3919), .CLK(clk), .Q(\ram[15][18] ) );
  DFFX1_HVT \ram_reg[15][17]  ( .D(n3918), .CLK(clk), .Q(\ram[15][17] ) );
  DFFX1_HVT \ram_reg[15][16]  ( .D(n3917), .CLK(clk), .Q(\ram[15][16] ) );
  DFFX1_HVT \ram_reg[15][15]  ( .D(n3916), .CLK(clk), .Q(\ram[15][15] ) );
  DFFX1_HVT \ram_reg[15][14]  ( .D(n3915), .CLK(clk), .Q(\ram[15][14] ) );
  DFFX1_HVT \ram_reg[15][13]  ( .D(n3914), .CLK(clk), .Q(\ram[15][13] ) );
  DFFX1_HVT \ram_reg[15][12]  ( .D(n3913), .CLK(clk), .Q(\ram[15][12] ) );
  DFFX1_HVT \ram_reg[15][11]  ( .D(n3912), .CLK(clk), .Q(\ram[15][11] ) );
  DFFX1_HVT \ram_reg[15][10]  ( .D(n3911), .CLK(clk), .Q(\ram[15][10] ) );
  DFFX1_HVT \ram_reg[15][9]  ( .D(n3910), .CLK(clk), .Q(\ram[15][9] ) );
  DFFX1_HVT \ram_reg[15][8]  ( .D(n3909), .CLK(clk), .Q(\ram[15][8] ) );
  DFFX1_HVT \ram_reg[15][7]  ( .D(n3908), .CLK(clk), .Q(\ram[15][7] ) );
  DFFX1_HVT \ram_reg[15][6]  ( .D(n3907), .CLK(clk), .Q(\ram[15][6] ) );
  DFFX1_HVT \ram_reg[15][5]  ( .D(n3906), .CLK(clk), .Q(\ram[15][5] ) );
  DFFX1_HVT \ram_reg[15][4]  ( .D(n3905), .CLK(clk), .Q(\ram[15][4] ) );
  DFFX1_HVT \ram_reg[15][3]  ( .D(n3904), .CLK(clk), .Q(\ram[15][3] ) );
  DFFX1_HVT \ram_reg[15][2]  ( .D(n3903), .CLK(clk), .Q(\ram[15][2] ) );
  DFFX1_HVT \ram_reg[15][1]  ( .D(n3902), .CLK(clk), .Q(\ram[15][1] ) );
  DFFX1_HVT \ram_reg[15][0]  ( .D(n3901), .CLK(clk), .Q(\ram[15][0] ) );
  DFFX1_HVT \ram_reg[14][255]  ( .D(n3900), .CLK(clk), .Q(\ram[14][255] ) );
  DFFX1_HVT \ram_reg[14][254]  ( .D(n3899), .CLK(clk), .Q(\ram[14][254] ) );
  DFFX1_HVT \ram_reg[14][253]  ( .D(n3898), .CLK(clk), .Q(\ram[14][253] ) );
  DFFX1_HVT \ram_reg[14][252]  ( .D(n3897), .CLK(clk), .Q(\ram[14][252] ) );
  DFFX1_HVT \ram_reg[14][251]  ( .D(n3896), .CLK(clk), .Q(\ram[14][251] ) );
  DFFX1_HVT \ram_reg[14][250]  ( .D(n3895), .CLK(clk), .Q(\ram[14][250] ) );
  DFFX1_HVT \ram_reg[14][249]  ( .D(n3894), .CLK(clk), .Q(\ram[14][249] ) );
  DFFX1_HVT \ram_reg[14][248]  ( .D(n3893), .CLK(clk), .Q(\ram[14][248] ) );
  DFFX1_HVT \ram_reg[14][247]  ( .D(n3892), .CLK(clk), .Q(\ram[14][247] ) );
  DFFX1_HVT \ram_reg[14][246]  ( .D(n3891), .CLK(clk), .Q(\ram[14][246] ) );
  DFFX1_HVT \ram_reg[14][245]  ( .D(n3890), .CLK(clk), .Q(\ram[14][245] ) );
  DFFX1_HVT \ram_reg[14][244]  ( .D(n3889), .CLK(clk), .Q(\ram[14][244] ) );
  DFFX1_HVT \ram_reg[14][243]  ( .D(n3888), .CLK(clk), .Q(\ram[14][243] ) );
  DFFX1_HVT \ram_reg[14][242]  ( .D(n3887), .CLK(clk), .Q(\ram[14][242] ) );
  DFFX1_HVT \ram_reg[14][241]  ( .D(n3886), .CLK(clk), .Q(\ram[14][241] ) );
  DFFX1_HVT \ram_reg[14][240]  ( .D(n3885), .CLK(clk), .Q(\ram[14][240] ) );
  DFFX1_HVT \ram_reg[14][239]  ( .D(n3884), .CLK(clk), .Q(\ram[14][239] ) );
  DFFX1_HVT \ram_reg[14][238]  ( .D(n3883), .CLK(clk), .Q(\ram[14][238] ) );
  DFFX1_HVT \ram_reg[14][237]  ( .D(n3882), .CLK(clk), .Q(\ram[14][237] ) );
  DFFX1_HVT \ram_reg[14][236]  ( .D(n3881), .CLK(clk), .Q(\ram[14][236] ) );
  DFFX1_HVT \ram_reg[14][235]  ( .D(n3880), .CLK(clk), .Q(\ram[14][235] ) );
  DFFX1_HVT \ram_reg[14][234]  ( .D(n3879), .CLK(clk), .Q(\ram[14][234] ) );
  DFFX1_HVT \ram_reg[14][233]  ( .D(n3878), .CLK(clk), .Q(\ram[14][233] ) );
  DFFX1_HVT \ram_reg[14][232]  ( .D(n3877), .CLK(clk), .Q(\ram[14][232] ) );
  DFFX1_HVT \ram_reg[14][231]  ( .D(n3876), .CLK(clk), .Q(\ram[14][231] ) );
  DFFX1_HVT \ram_reg[14][230]  ( .D(n3875), .CLK(clk), .Q(\ram[14][230] ) );
  DFFX1_HVT \ram_reg[14][229]  ( .D(n3874), .CLK(clk), .Q(\ram[14][229] ) );
  DFFX1_HVT \ram_reg[14][228]  ( .D(n3873), .CLK(clk), .Q(\ram[14][228] ) );
  DFFX1_HVT \ram_reg[14][227]  ( .D(n3872), .CLK(clk), .Q(\ram[14][227] ) );
  DFFX1_HVT \ram_reg[14][226]  ( .D(n3871), .CLK(clk), .Q(\ram[14][226] ) );
  DFFX1_HVT \ram_reg[14][225]  ( .D(n3870), .CLK(clk), .Q(\ram[14][225] ) );
  DFFX1_HVT \ram_reg[14][224]  ( .D(n3869), .CLK(clk), .Q(\ram[14][224] ) );
  DFFX1_HVT \ram_reg[14][223]  ( .D(n3868), .CLK(clk), .Q(\ram[14][223] ) );
  DFFX1_HVT \ram_reg[14][222]  ( .D(n3867), .CLK(clk), .Q(\ram[14][222] ) );
  DFFX1_HVT \ram_reg[14][221]  ( .D(n3866), .CLK(clk), .Q(\ram[14][221] ) );
  DFFX1_HVT \ram_reg[14][220]  ( .D(n3865), .CLK(clk), .Q(\ram[14][220] ) );
  DFFX1_HVT \ram_reg[14][219]  ( .D(n3864), .CLK(clk), .Q(\ram[14][219] ) );
  DFFX1_HVT \ram_reg[14][218]  ( .D(n3863), .CLK(clk), .Q(\ram[14][218] ) );
  DFFX1_HVT \ram_reg[14][217]  ( .D(n3862), .CLK(clk), .Q(\ram[14][217] ) );
  DFFX1_HVT \ram_reg[14][216]  ( .D(n3861), .CLK(clk), .Q(\ram[14][216] ) );
  DFFX1_HVT \ram_reg[14][215]  ( .D(n3860), .CLK(clk), .Q(\ram[14][215] ) );
  DFFX1_HVT \ram_reg[14][214]  ( .D(n3859), .CLK(clk), .Q(\ram[14][214] ) );
  DFFX1_HVT \ram_reg[14][213]  ( .D(n3858), .CLK(clk), .Q(\ram[14][213] ) );
  DFFX1_HVT \ram_reg[14][212]  ( .D(n3857), .CLK(clk), .Q(\ram[14][212] ) );
  DFFX1_HVT \ram_reg[14][211]  ( .D(n3856), .CLK(clk), .Q(\ram[14][211] ) );
  DFFX1_HVT \ram_reg[14][210]  ( .D(n3855), .CLK(clk), .Q(\ram[14][210] ) );
  DFFX1_HVT \ram_reg[14][209]  ( .D(n3854), .CLK(clk), .Q(\ram[14][209] ) );
  DFFX1_HVT \ram_reg[14][208]  ( .D(n3853), .CLK(clk), .Q(\ram[14][208] ) );
  DFFX1_HVT \ram_reg[14][207]  ( .D(n3852), .CLK(clk), .Q(\ram[14][207] ) );
  DFFX1_HVT \ram_reg[14][206]  ( .D(n3851), .CLK(clk), .Q(\ram[14][206] ) );
  DFFX1_HVT \ram_reg[14][205]  ( .D(n3850), .CLK(clk), .Q(\ram[14][205] ) );
  DFFX1_HVT \ram_reg[14][204]  ( .D(n3849), .CLK(clk), .Q(\ram[14][204] ) );
  DFFX1_HVT \ram_reg[14][203]  ( .D(n3848), .CLK(clk), .Q(\ram[14][203] ) );
  DFFX1_HVT \ram_reg[14][202]  ( .D(n3847), .CLK(clk), .Q(\ram[14][202] ) );
  DFFX1_HVT \ram_reg[14][201]  ( .D(n3846), .CLK(clk), .Q(\ram[14][201] ) );
  DFFX1_HVT \ram_reg[14][200]  ( .D(n3845), .CLK(clk), .Q(\ram[14][200] ) );
  DFFX1_HVT \ram_reg[14][199]  ( .D(n3844), .CLK(clk), .Q(\ram[14][199] ) );
  DFFX1_HVT \ram_reg[14][198]  ( .D(n3843), .CLK(clk), .Q(\ram[14][198] ) );
  DFFX1_HVT \ram_reg[14][197]  ( .D(n3842), .CLK(clk), .Q(\ram[14][197] ) );
  DFFX1_HVT \ram_reg[14][196]  ( .D(n3841), .CLK(clk), .Q(\ram[14][196] ) );
  DFFX1_HVT \ram_reg[14][195]  ( .D(n3840), .CLK(clk), .Q(\ram[14][195] ) );
  DFFX1_HVT \ram_reg[14][194]  ( .D(n3839), .CLK(clk), .Q(\ram[14][194] ) );
  DFFX1_HVT \ram_reg[14][193]  ( .D(n3838), .CLK(clk), .Q(\ram[14][193] ) );
  DFFX1_HVT \ram_reg[14][192]  ( .D(n3837), .CLK(clk), .Q(\ram[14][192] ) );
  DFFX1_HVT \ram_reg[14][191]  ( .D(n3836), .CLK(clk), .Q(\ram[14][191] ) );
  DFFX1_HVT \ram_reg[14][190]  ( .D(n3835), .CLK(clk), .Q(\ram[14][190] ) );
  DFFX1_HVT \ram_reg[14][189]  ( .D(n3834), .CLK(clk), .Q(\ram[14][189] ) );
  DFFX1_HVT \ram_reg[14][188]  ( .D(n3833), .CLK(clk), .Q(\ram[14][188] ) );
  DFFX1_HVT \ram_reg[14][187]  ( .D(n3832), .CLK(clk), .Q(\ram[14][187] ) );
  DFFX1_HVT \ram_reg[14][186]  ( .D(n3831), .CLK(clk), .Q(\ram[14][186] ) );
  DFFX1_HVT \ram_reg[14][185]  ( .D(n3830), .CLK(clk), .Q(\ram[14][185] ) );
  DFFX1_HVT \ram_reg[14][184]  ( .D(n3829), .CLK(clk), .Q(\ram[14][184] ) );
  DFFX1_HVT \ram_reg[14][183]  ( .D(n3828), .CLK(clk), .Q(\ram[14][183] ) );
  DFFX1_HVT \ram_reg[14][182]  ( .D(n3827), .CLK(clk), .Q(\ram[14][182] ) );
  DFFX1_HVT \ram_reg[14][181]  ( .D(n3826), .CLK(clk), .Q(\ram[14][181] ) );
  DFFX1_HVT \ram_reg[14][180]  ( .D(n3825), .CLK(clk), .Q(\ram[14][180] ) );
  DFFX1_HVT \ram_reg[14][179]  ( .D(n3824), .CLK(clk), .Q(\ram[14][179] ) );
  DFFX1_HVT \ram_reg[14][178]  ( .D(n3823), .CLK(clk), .Q(\ram[14][178] ) );
  DFFX1_HVT \ram_reg[14][177]  ( .D(n3822), .CLK(clk), .Q(\ram[14][177] ) );
  DFFX1_HVT \ram_reg[14][176]  ( .D(n3821), .CLK(clk), .Q(\ram[14][176] ) );
  DFFX1_HVT \ram_reg[14][175]  ( .D(n3820), .CLK(clk), .Q(\ram[14][175] ) );
  DFFX1_HVT \ram_reg[14][174]  ( .D(n3819), .CLK(clk), .Q(\ram[14][174] ) );
  DFFX1_HVT \ram_reg[14][173]  ( .D(n3818), .CLK(clk), .Q(\ram[14][173] ) );
  DFFX1_HVT \ram_reg[14][172]  ( .D(n3817), .CLK(clk), .Q(\ram[14][172] ) );
  DFFX1_HVT \ram_reg[14][171]  ( .D(n3816), .CLK(clk), .Q(\ram[14][171] ) );
  DFFX1_HVT \ram_reg[14][170]  ( .D(n3815), .CLK(clk), .Q(\ram[14][170] ) );
  DFFX1_HVT \ram_reg[14][169]  ( .D(n3814), .CLK(clk), .Q(\ram[14][169] ) );
  DFFX1_HVT \ram_reg[14][168]  ( .D(n3813), .CLK(clk), .Q(\ram[14][168] ) );
  DFFX1_HVT \ram_reg[14][167]  ( .D(n3812), .CLK(clk), .Q(\ram[14][167] ) );
  DFFX1_HVT \ram_reg[14][166]  ( .D(n3811), .CLK(clk), .Q(\ram[14][166] ) );
  DFFX1_HVT \ram_reg[14][165]  ( .D(n3810), .CLK(clk), .Q(\ram[14][165] ) );
  DFFX1_HVT \ram_reg[14][164]  ( .D(n3809), .CLK(clk), .Q(\ram[14][164] ) );
  DFFX1_HVT \ram_reg[14][163]  ( .D(n3808), .CLK(clk), .Q(\ram[14][163] ) );
  DFFX1_HVT \ram_reg[14][162]  ( .D(n3807), .CLK(clk), .Q(\ram[14][162] ) );
  DFFX1_HVT \ram_reg[14][161]  ( .D(n3806), .CLK(clk), .Q(\ram[14][161] ) );
  DFFX1_HVT \ram_reg[14][160]  ( .D(n3805), .CLK(clk), .Q(\ram[14][160] ) );
  DFFX1_HVT \ram_reg[14][159]  ( .D(n3804), .CLK(clk), .Q(\ram[14][159] ) );
  DFFX1_HVT \ram_reg[14][158]  ( .D(n3803), .CLK(clk), .Q(\ram[14][158] ) );
  DFFX1_HVT \ram_reg[14][157]  ( .D(n3802), .CLK(clk), .Q(\ram[14][157] ) );
  DFFX1_HVT \ram_reg[14][156]  ( .D(n3801), .CLK(clk), .Q(\ram[14][156] ) );
  DFFX1_HVT \ram_reg[14][155]  ( .D(n3800), .CLK(clk), .Q(\ram[14][155] ) );
  DFFX1_HVT \ram_reg[14][154]  ( .D(n3799), .CLK(clk), .Q(\ram[14][154] ) );
  DFFX1_HVT \ram_reg[14][153]  ( .D(n3798), .CLK(clk), .Q(\ram[14][153] ) );
  DFFX1_HVT \ram_reg[14][152]  ( .D(n3797), .CLK(clk), .Q(\ram[14][152] ) );
  DFFX1_HVT \ram_reg[14][151]  ( .D(n3796), .CLK(clk), .Q(\ram[14][151] ) );
  DFFX1_HVT \ram_reg[14][150]  ( .D(n3795), .CLK(clk), .Q(\ram[14][150] ) );
  DFFX1_HVT \ram_reg[14][149]  ( .D(n3794), .CLK(clk), .Q(\ram[14][149] ) );
  DFFX1_HVT \ram_reg[14][148]  ( .D(n3793), .CLK(clk), .Q(\ram[14][148] ) );
  DFFX1_HVT \ram_reg[14][147]  ( .D(n3792), .CLK(clk), .Q(\ram[14][147] ) );
  DFFX1_HVT \ram_reg[14][146]  ( .D(n3791), .CLK(clk), .Q(\ram[14][146] ) );
  DFFX1_HVT \ram_reg[14][145]  ( .D(n3790), .CLK(clk), .Q(\ram[14][145] ) );
  DFFX1_HVT \ram_reg[14][144]  ( .D(n3789), .CLK(clk), .Q(\ram[14][144] ) );
  DFFX1_HVT \ram_reg[14][143]  ( .D(n3788), .CLK(clk), .Q(\ram[14][143] ) );
  DFFX1_HVT \ram_reg[14][142]  ( .D(n3787), .CLK(clk), .Q(\ram[14][142] ) );
  DFFX1_HVT \ram_reg[14][141]  ( .D(n3786), .CLK(clk), .Q(\ram[14][141] ) );
  DFFX1_HVT \ram_reg[14][140]  ( .D(n3785), .CLK(clk), .Q(\ram[14][140] ) );
  DFFX1_HVT \ram_reg[14][139]  ( .D(n3784), .CLK(clk), .Q(\ram[14][139] ) );
  DFFX1_HVT \ram_reg[14][138]  ( .D(n3783), .CLK(clk), .Q(\ram[14][138] ) );
  DFFX1_HVT \ram_reg[14][137]  ( .D(n3782), .CLK(clk), .Q(\ram[14][137] ) );
  DFFX1_HVT \ram_reg[14][136]  ( .D(n3781), .CLK(clk), .Q(\ram[14][136] ) );
  DFFX1_HVT \ram_reg[14][135]  ( .D(n3780), .CLK(clk), .Q(\ram[14][135] ) );
  DFFX1_HVT \ram_reg[14][134]  ( .D(n3779), .CLK(clk), .Q(\ram[14][134] ) );
  DFFX1_HVT \ram_reg[14][133]  ( .D(n3778), .CLK(clk), .Q(\ram[14][133] ) );
  DFFX1_HVT \ram_reg[14][132]  ( .D(n3777), .CLK(clk), .Q(\ram[14][132] ) );
  DFFX1_HVT \ram_reg[14][131]  ( .D(n3776), .CLK(clk), .Q(\ram[14][131] ) );
  DFFX1_HVT \ram_reg[14][130]  ( .D(n3775), .CLK(clk), .Q(\ram[14][130] ) );
  DFFX1_HVT \ram_reg[14][129]  ( .D(n3774), .CLK(clk), .Q(\ram[14][129] ) );
  DFFX1_HVT \ram_reg[14][128]  ( .D(n3773), .CLK(clk), .Q(\ram[14][128] ) );
  DFFX1_HVT \ram_reg[14][127]  ( .D(n3772), .CLK(clk), .Q(\ram[14][127] ) );
  DFFX1_HVT \ram_reg[14][126]  ( .D(n3771), .CLK(clk), .Q(\ram[14][126] ) );
  DFFX1_HVT \ram_reg[14][125]  ( .D(n3770), .CLK(clk), .Q(\ram[14][125] ) );
  DFFX1_HVT \ram_reg[14][124]  ( .D(n3769), .CLK(clk), .Q(\ram[14][124] ) );
  DFFX1_HVT \ram_reg[14][123]  ( .D(n3768), .CLK(clk), .Q(\ram[14][123] ) );
  DFFX1_HVT \ram_reg[14][122]  ( .D(n3767), .CLK(clk), .Q(\ram[14][122] ) );
  DFFX1_HVT \ram_reg[14][121]  ( .D(n3766), .CLK(clk), .Q(\ram[14][121] ) );
  DFFX1_HVT \ram_reg[14][120]  ( .D(n3765), .CLK(clk), .Q(\ram[14][120] ) );
  DFFX1_HVT \ram_reg[14][119]  ( .D(n3764), .CLK(clk), .Q(\ram[14][119] ) );
  DFFX1_HVT \ram_reg[14][118]  ( .D(n3763), .CLK(clk), .Q(\ram[14][118] ) );
  DFFX1_HVT \ram_reg[14][117]  ( .D(n3762), .CLK(clk), .Q(\ram[14][117] ) );
  DFFX1_HVT \ram_reg[14][116]  ( .D(n3761), .CLK(clk), .Q(\ram[14][116] ) );
  DFFX1_HVT \ram_reg[14][115]  ( .D(n3760), .CLK(clk), .Q(\ram[14][115] ) );
  DFFX1_HVT \ram_reg[14][114]  ( .D(n3759), .CLK(clk), .Q(\ram[14][114] ) );
  DFFX1_HVT \ram_reg[14][113]  ( .D(n3758), .CLK(clk), .Q(\ram[14][113] ) );
  DFFX1_HVT \ram_reg[14][112]  ( .D(n3757), .CLK(clk), .Q(\ram[14][112] ) );
  DFFX1_HVT \ram_reg[14][111]  ( .D(n3756), .CLK(clk), .Q(\ram[14][111] ) );
  DFFX1_HVT \ram_reg[14][110]  ( .D(n3755), .CLK(clk), .Q(\ram[14][110] ) );
  DFFX1_HVT \ram_reg[14][109]  ( .D(n3754), .CLK(clk), .Q(\ram[14][109] ) );
  DFFX1_HVT \ram_reg[14][108]  ( .D(n3753), .CLK(clk), .Q(\ram[14][108] ) );
  DFFX1_HVT \ram_reg[14][107]  ( .D(n3752), .CLK(clk), .Q(\ram[14][107] ) );
  DFFX1_HVT \ram_reg[14][106]  ( .D(n3751), .CLK(clk), .Q(\ram[14][106] ) );
  DFFX1_HVT \ram_reg[14][105]  ( .D(n3750), .CLK(clk), .Q(\ram[14][105] ) );
  DFFX1_HVT \ram_reg[14][104]  ( .D(n3749), .CLK(clk), .Q(\ram[14][104] ) );
  DFFX1_HVT \ram_reg[14][103]  ( .D(n3748), .CLK(clk), .Q(\ram[14][103] ) );
  DFFX1_HVT \ram_reg[14][102]  ( .D(n3747), .CLK(clk), .Q(\ram[14][102] ) );
  DFFX1_HVT \ram_reg[14][101]  ( .D(n3746), .CLK(clk), .Q(\ram[14][101] ) );
  DFFX1_HVT \ram_reg[14][100]  ( .D(n3745), .CLK(clk), .Q(\ram[14][100] ) );
  DFFX1_HVT \ram_reg[14][99]  ( .D(n3744), .CLK(clk), .Q(\ram[14][99] ) );
  DFFX1_HVT \ram_reg[14][98]  ( .D(n3743), .CLK(clk), .Q(\ram[14][98] ) );
  DFFX1_HVT \ram_reg[14][97]  ( .D(n3742), .CLK(clk), .Q(\ram[14][97] ) );
  DFFX1_HVT \ram_reg[14][96]  ( .D(n3741), .CLK(clk), .Q(\ram[14][96] ) );
  DFFX1_HVT \ram_reg[14][95]  ( .D(n3740), .CLK(clk), .Q(\ram[14][95] ) );
  DFFX1_HVT \ram_reg[14][94]  ( .D(n3739), .CLK(clk), .Q(\ram[14][94] ) );
  DFFX1_HVT \ram_reg[14][93]  ( .D(n3738), .CLK(clk), .Q(\ram[14][93] ) );
  DFFX1_HVT \ram_reg[14][92]  ( .D(n3737), .CLK(clk), .Q(\ram[14][92] ) );
  DFFX1_HVT \ram_reg[14][91]  ( .D(n3736), .CLK(clk), .Q(\ram[14][91] ) );
  DFFX1_HVT \ram_reg[14][90]  ( .D(n3735), .CLK(clk), .Q(\ram[14][90] ) );
  DFFX1_HVT \ram_reg[14][89]  ( .D(n3734), .CLK(clk), .Q(\ram[14][89] ) );
  DFFX1_HVT \ram_reg[14][88]  ( .D(n3733), .CLK(clk), .Q(\ram[14][88] ) );
  DFFX1_HVT \ram_reg[14][87]  ( .D(n3732), .CLK(clk), .Q(\ram[14][87] ) );
  DFFX1_HVT \ram_reg[14][86]  ( .D(n3731), .CLK(clk), .Q(\ram[14][86] ) );
  DFFX1_HVT \ram_reg[14][85]  ( .D(n3730), .CLK(clk), .Q(\ram[14][85] ) );
  DFFX1_HVT \ram_reg[14][84]  ( .D(n3729), .CLK(clk), .Q(\ram[14][84] ) );
  DFFX1_HVT \ram_reg[14][83]  ( .D(n3728), .CLK(clk), .Q(\ram[14][83] ) );
  DFFX1_HVT \ram_reg[14][82]  ( .D(n3727), .CLK(clk), .Q(\ram[14][82] ) );
  DFFX1_HVT \ram_reg[14][81]  ( .D(n3726), .CLK(clk), .Q(\ram[14][81] ) );
  DFFX1_HVT \ram_reg[14][80]  ( .D(n3725), .CLK(clk), .Q(\ram[14][80] ) );
  DFFX1_HVT \ram_reg[14][79]  ( .D(n3724), .CLK(clk), .Q(\ram[14][79] ) );
  DFFX1_HVT \ram_reg[14][78]  ( .D(n3723), .CLK(clk), .Q(\ram[14][78] ) );
  DFFX1_HVT \ram_reg[14][77]  ( .D(n3722), .CLK(clk), .Q(\ram[14][77] ) );
  DFFX1_HVT \ram_reg[14][76]  ( .D(n3721), .CLK(clk), .Q(\ram[14][76] ) );
  DFFX1_HVT \ram_reg[14][75]  ( .D(n3720), .CLK(clk), .Q(\ram[14][75] ) );
  DFFX1_HVT \ram_reg[14][74]  ( .D(n3719), .CLK(clk), .Q(\ram[14][74] ) );
  DFFX1_HVT \ram_reg[14][73]  ( .D(n3718), .CLK(clk), .Q(\ram[14][73] ) );
  DFFX1_HVT \ram_reg[14][72]  ( .D(n3717), .CLK(clk), .Q(\ram[14][72] ) );
  DFFX1_HVT \ram_reg[14][71]  ( .D(n3716), .CLK(clk), .Q(\ram[14][71] ) );
  DFFX1_HVT \ram_reg[14][70]  ( .D(n3715), .CLK(clk), .Q(\ram[14][70] ) );
  DFFX1_HVT \ram_reg[14][69]  ( .D(n3714), .CLK(clk), .Q(\ram[14][69] ) );
  DFFX1_HVT \ram_reg[14][68]  ( .D(n3713), .CLK(clk), .Q(\ram[14][68] ) );
  DFFX1_HVT \ram_reg[14][67]  ( .D(n3712), .CLK(clk), .Q(\ram[14][67] ) );
  DFFX1_HVT \ram_reg[14][66]  ( .D(n3711), .CLK(clk), .Q(\ram[14][66] ) );
  DFFX1_HVT \ram_reg[14][65]  ( .D(n3710), .CLK(clk), .Q(\ram[14][65] ) );
  DFFX1_HVT \ram_reg[14][64]  ( .D(n3709), .CLK(clk), .Q(\ram[14][64] ) );
  DFFX1_HVT \ram_reg[14][63]  ( .D(n3708), .CLK(clk), .Q(\ram[14][63] ) );
  DFFX1_HVT \ram_reg[14][62]  ( .D(n3707), .CLK(clk), .Q(\ram[14][62] ) );
  DFFX1_HVT \ram_reg[14][61]  ( .D(n3706), .CLK(clk), .Q(\ram[14][61] ) );
  DFFX1_HVT \ram_reg[14][60]  ( .D(n3705), .CLK(clk), .Q(\ram[14][60] ) );
  DFFX1_HVT \ram_reg[14][59]  ( .D(n3704), .CLK(clk), .Q(\ram[14][59] ) );
  DFFX1_HVT \ram_reg[14][58]  ( .D(n3703), .CLK(clk), .Q(\ram[14][58] ) );
  DFFX1_HVT \ram_reg[14][57]  ( .D(n3702), .CLK(clk), .Q(\ram[14][57] ) );
  DFFX1_HVT \ram_reg[14][56]  ( .D(n3701), .CLK(clk), .Q(\ram[14][56] ) );
  DFFX1_HVT \ram_reg[14][55]  ( .D(n3700), .CLK(clk), .Q(\ram[14][55] ) );
  DFFX1_HVT \ram_reg[14][54]  ( .D(n3699), .CLK(clk), .Q(\ram[14][54] ) );
  DFFX1_HVT \ram_reg[14][53]  ( .D(n3698), .CLK(clk), .Q(\ram[14][53] ) );
  DFFX1_HVT \ram_reg[14][52]  ( .D(n3697), .CLK(clk), .Q(\ram[14][52] ) );
  DFFX1_HVT \ram_reg[14][51]  ( .D(n3696), .CLK(clk), .Q(\ram[14][51] ) );
  DFFX1_HVT \ram_reg[14][50]  ( .D(n3695), .CLK(clk), .Q(\ram[14][50] ) );
  DFFX1_HVT \ram_reg[14][49]  ( .D(n3694), .CLK(clk), .Q(\ram[14][49] ) );
  DFFX1_HVT \ram_reg[14][48]  ( .D(n3693), .CLK(clk), .Q(\ram[14][48] ) );
  DFFX1_HVT \ram_reg[14][47]  ( .D(n3692), .CLK(clk), .Q(\ram[14][47] ) );
  DFFX1_HVT \ram_reg[14][46]  ( .D(n3691), .CLK(clk), .Q(\ram[14][46] ) );
  DFFX1_HVT \ram_reg[14][45]  ( .D(n3690), .CLK(clk), .Q(\ram[14][45] ) );
  DFFX1_HVT \ram_reg[14][44]  ( .D(n3689), .CLK(clk), .Q(\ram[14][44] ) );
  DFFX1_HVT \ram_reg[14][43]  ( .D(n3688), .CLK(clk), .Q(\ram[14][43] ) );
  DFFX1_HVT \ram_reg[14][42]  ( .D(n3687), .CLK(clk), .Q(\ram[14][42] ) );
  DFFX1_HVT \ram_reg[14][41]  ( .D(n3686), .CLK(clk), .Q(\ram[14][41] ) );
  DFFX1_HVT \ram_reg[14][40]  ( .D(n3685), .CLK(clk), .Q(\ram[14][40] ) );
  DFFX1_HVT \ram_reg[14][39]  ( .D(n3684), .CLK(clk), .Q(\ram[14][39] ) );
  DFFX1_HVT \ram_reg[14][38]  ( .D(n3683), .CLK(clk), .Q(\ram[14][38] ) );
  DFFX1_HVT \ram_reg[14][37]  ( .D(n3682), .CLK(clk), .Q(\ram[14][37] ) );
  DFFX1_HVT \ram_reg[14][36]  ( .D(n3681), .CLK(clk), .Q(\ram[14][36] ) );
  DFFX1_HVT \ram_reg[14][35]  ( .D(n3680), .CLK(clk), .Q(\ram[14][35] ) );
  DFFX1_HVT \ram_reg[14][34]  ( .D(n3679), .CLK(clk), .Q(\ram[14][34] ) );
  DFFX1_HVT \ram_reg[14][33]  ( .D(n3678), .CLK(clk), .Q(\ram[14][33] ) );
  DFFX1_HVT \ram_reg[14][32]  ( .D(n3677), .CLK(clk), .Q(\ram[14][32] ) );
  DFFX1_HVT \ram_reg[14][31]  ( .D(n3676), .CLK(clk), .Q(\ram[14][31] ) );
  DFFX1_HVT \ram_reg[14][30]  ( .D(n3675), .CLK(clk), .Q(\ram[14][30] ) );
  DFFX1_HVT \ram_reg[14][29]  ( .D(n3674), .CLK(clk), .Q(\ram[14][29] ) );
  DFFX1_HVT \ram_reg[14][28]  ( .D(n3673), .CLK(clk), .Q(\ram[14][28] ) );
  DFFX1_HVT \ram_reg[14][27]  ( .D(n3672), .CLK(clk), .Q(\ram[14][27] ) );
  DFFX1_HVT \ram_reg[14][26]  ( .D(n3671), .CLK(clk), .Q(\ram[14][26] ) );
  DFFX1_HVT \ram_reg[14][25]  ( .D(n3670), .CLK(clk), .Q(\ram[14][25] ) );
  DFFX1_HVT \ram_reg[14][24]  ( .D(n3669), .CLK(clk), .Q(\ram[14][24] ) );
  DFFX1_HVT \ram_reg[14][23]  ( .D(n3668), .CLK(clk), .Q(\ram[14][23] ) );
  DFFX1_HVT \ram_reg[14][22]  ( .D(n3667), .CLK(clk), .Q(\ram[14][22] ) );
  DFFX1_HVT \ram_reg[14][21]  ( .D(n3666), .CLK(clk), .Q(\ram[14][21] ) );
  DFFX1_HVT \ram_reg[14][20]  ( .D(n3665), .CLK(clk), .Q(\ram[14][20] ) );
  DFFX1_HVT \ram_reg[14][19]  ( .D(n3664), .CLK(clk), .Q(\ram[14][19] ) );
  DFFX1_HVT \ram_reg[14][18]  ( .D(n3663), .CLK(clk), .Q(\ram[14][18] ) );
  DFFX1_HVT \ram_reg[14][17]  ( .D(n3662), .CLK(clk), .Q(\ram[14][17] ) );
  DFFX1_HVT \ram_reg[14][16]  ( .D(n3661), .CLK(clk), .Q(\ram[14][16] ) );
  DFFX1_HVT \ram_reg[14][15]  ( .D(n3660), .CLK(clk), .Q(\ram[14][15] ) );
  DFFX1_HVT \ram_reg[14][14]  ( .D(n3659), .CLK(clk), .Q(\ram[14][14] ) );
  DFFX1_HVT \ram_reg[14][13]  ( .D(n3658), .CLK(clk), .Q(\ram[14][13] ) );
  DFFX1_HVT \ram_reg[14][12]  ( .D(n3657), .CLK(clk), .Q(\ram[14][12] ) );
  DFFX1_HVT \ram_reg[14][11]  ( .D(n3656), .CLK(clk), .Q(\ram[14][11] ) );
  DFFX1_HVT \ram_reg[14][10]  ( .D(n3655), .CLK(clk), .Q(\ram[14][10] ) );
  DFFX1_HVT \ram_reg[14][9]  ( .D(n3654), .CLK(clk), .Q(\ram[14][9] ) );
  DFFX1_HVT \ram_reg[14][8]  ( .D(n3653), .CLK(clk), .Q(\ram[14][8] ) );
  DFFX1_HVT \ram_reg[14][7]  ( .D(n3652), .CLK(clk), .Q(\ram[14][7] ) );
  DFFX1_HVT \ram_reg[14][6]  ( .D(n3651), .CLK(clk), .Q(\ram[14][6] ) );
  DFFX1_HVT \ram_reg[14][5]  ( .D(n3650), .CLK(clk), .Q(\ram[14][5] ) );
  DFFX1_HVT \ram_reg[14][4]  ( .D(n3649), .CLK(clk), .Q(\ram[14][4] ) );
  DFFX1_HVT \ram_reg[14][3]  ( .D(n3648), .CLK(clk), .Q(\ram[14][3] ) );
  DFFX1_HVT \ram_reg[14][2]  ( .D(n3647), .CLK(clk), .Q(\ram[14][2] ) );
  DFFX1_HVT \ram_reg[14][1]  ( .D(n3646), .CLK(clk), .Q(\ram[14][1] ) );
  DFFX1_HVT \ram_reg[14][0]  ( .D(n3645), .CLK(clk), .Q(\ram[14][0] ) );
  DFFX1_HVT \ram_reg[13][255]  ( .D(n3644), .CLK(clk), .Q(\ram[13][255] ) );
  DFFX1_HVT \ram_reg[13][254]  ( .D(n3643), .CLK(clk), .Q(\ram[13][254] ) );
  DFFX1_HVT \ram_reg[13][253]  ( .D(n3642), .CLK(clk), .Q(\ram[13][253] ) );
  DFFX1_HVT \ram_reg[13][252]  ( .D(n3641), .CLK(clk), .Q(\ram[13][252] ) );
  DFFX1_HVT \ram_reg[13][251]  ( .D(n3640), .CLK(clk), .Q(\ram[13][251] ) );
  DFFX1_HVT \ram_reg[13][250]  ( .D(n3639), .CLK(clk), .Q(\ram[13][250] ) );
  DFFX1_HVT \ram_reg[13][249]  ( .D(n3638), .CLK(clk), .Q(\ram[13][249] ) );
  DFFX1_HVT \ram_reg[13][248]  ( .D(n3637), .CLK(clk), .Q(\ram[13][248] ) );
  DFFX1_HVT \ram_reg[13][247]  ( .D(n3636), .CLK(clk), .Q(\ram[13][247] ) );
  DFFX1_HVT \ram_reg[13][246]  ( .D(n3635), .CLK(clk), .Q(\ram[13][246] ) );
  DFFX1_HVT \ram_reg[13][245]  ( .D(n3634), .CLK(clk), .Q(\ram[13][245] ) );
  DFFX1_HVT \ram_reg[13][244]  ( .D(n3633), .CLK(clk), .Q(\ram[13][244] ) );
  DFFX1_HVT \ram_reg[13][243]  ( .D(n3632), .CLK(clk), .Q(\ram[13][243] ) );
  DFFX1_HVT \ram_reg[13][242]  ( .D(n3631), .CLK(clk), .Q(\ram[13][242] ) );
  DFFX1_HVT \ram_reg[13][241]  ( .D(n3630), .CLK(clk), .Q(\ram[13][241] ) );
  DFFX1_HVT \ram_reg[13][240]  ( .D(n3629), .CLK(clk), .Q(\ram[13][240] ) );
  DFFX1_HVT \ram_reg[13][239]  ( .D(n3628), .CLK(clk), .Q(\ram[13][239] ) );
  DFFX1_HVT \ram_reg[13][238]  ( .D(n3627), .CLK(clk), .Q(\ram[13][238] ) );
  DFFX1_HVT \ram_reg[13][237]  ( .D(n3626), .CLK(clk), .Q(\ram[13][237] ) );
  DFFX1_HVT \ram_reg[13][236]  ( .D(n3625), .CLK(clk), .Q(\ram[13][236] ) );
  DFFX1_HVT \ram_reg[13][235]  ( .D(n3624), .CLK(clk), .Q(\ram[13][235] ) );
  DFFX1_HVT \ram_reg[13][234]  ( .D(n3623), .CLK(clk), .Q(\ram[13][234] ) );
  DFFX1_HVT \ram_reg[13][233]  ( .D(n3622), .CLK(clk), .Q(\ram[13][233] ) );
  DFFX1_HVT \ram_reg[13][232]  ( .D(n3621), .CLK(clk), .Q(\ram[13][232] ) );
  DFFX1_HVT \ram_reg[13][231]  ( .D(n3620), .CLK(clk), .Q(\ram[13][231] ) );
  DFFX1_HVT \ram_reg[13][230]  ( .D(n3619), .CLK(clk), .Q(\ram[13][230] ) );
  DFFX1_HVT \ram_reg[13][229]  ( .D(n3618), .CLK(clk), .Q(\ram[13][229] ) );
  DFFX1_HVT \ram_reg[13][228]  ( .D(n3617), .CLK(clk), .Q(\ram[13][228] ) );
  DFFX1_HVT \ram_reg[13][227]  ( .D(n3616), .CLK(clk), .Q(\ram[13][227] ) );
  DFFX1_HVT \ram_reg[13][226]  ( .D(n3615), .CLK(clk), .Q(\ram[13][226] ) );
  DFFX1_HVT \ram_reg[13][225]  ( .D(n3614), .CLK(clk), .Q(\ram[13][225] ) );
  DFFX1_HVT \ram_reg[13][224]  ( .D(n3613), .CLK(clk), .Q(\ram[13][224] ) );
  DFFX1_HVT \ram_reg[13][223]  ( .D(n3612), .CLK(clk), .Q(\ram[13][223] ) );
  DFFX1_HVT \ram_reg[13][222]  ( .D(n3611), .CLK(clk), .Q(\ram[13][222] ) );
  DFFX1_HVT \ram_reg[13][221]  ( .D(n3610), .CLK(clk), .Q(\ram[13][221] ) );
  DFFX1_HVT \ram_reg[13][220]  ( .D(n3609), .CLK(clk), .Q(\ram[13][220] ) );
  DFFX1_HVT \ram_reg[13][219]  ( .D(n3608), .CLK(clk), .Q(\ram[13][219] ) );
  DFFX1_HVT \ram_reg[13][218]  ( .D(n3607), .CLK(clk), .Q(\ram[13][218] ) );
  DFFX1_HVT \ram_reg[13][217]  ( .D(n3606), .CLK(clk), .Q(\ram[13][217] ) );
  DFFX1_HVT \ram_reg[13][216]  ( .D(n3605), .CLK(clk), .Q(\ram[13][216] ) );
  DFFX1_HVT \ram_reg[13][215]  ( .D(n3604), .CLK(clk), .Q(\ram[13][215] ) );
  DFFX1_HVT \ram_reg[13][214]  ( .D(n3603), .CLK(clk), .Q(\ram[13][214] ) );
  DFFX1_HVT \ram_reg[13][213]  ( .D(n3602), .CLK(clk), .Q(\ram[13][213] ) );
  DFFX1_HVT \ram_reg[13][212]  ( .D(n3601), .CLK(clk), .Q(\ram[13][212] ) );
  DFFX1_HVT \ram_reg[13][211]  ( .D(n3600), .CLK(clk), .Q(\ram[13][211] ) );
  DFFX1_HVT \ram_reg[13][210]  ( .D(n3599), .CLK(clk), .Q(\ram[13][210] ) );
  DFFX1_HVT \ram_reg[13][209]  ( .D(n3598), .CLK(clk), .Q(\ram[13][209] ) );
  DFFX1_HVT \ram_reg[13][208]  ( .D(n3597), .CLK(clk), .Q(\ram[13][208] ) );
  DFFX1_HVT \ram_reg[13][207]  ( .D(n3596), .CLK(clk), .Q(\ram[13][207] ) );
  DFFX1_HVT \ram_reg[13][206]  ( .D(n3595), .CLK(clk), .Q(\ram[13][206] ) );
  DFFX1_HVT \ram_reg[13][205]  ( .D(n3594), .CLK(clk), .Q(\ram[13][205] ) );
  DFFX1_HVT \ram_reg[13][204]  ( .D(n3593), .CLK(clk), .Q(\ram[13][204] ) );
  DFFX1_HVT \ram_reg[13][203]  ( .D(n3592), .CLK(clk), .Q(\ram[13][203] ) );
  DFFX1_HVT \ram_reg[13][202]  ( .D(n3591), .CLK(clk), .Q(\ram[13][202] ) );
  DFFX1_HVT \ram_reg[13][201]  ( .D(n3590), .CLK(clk), .Q(\ram[13][201] ) );
  DFFX1_HVT \ram_reg[13][200]  ( .D(n3589), .CLK(clk), .Q(\ram[13][200] ) );
  DFFX1_HVT \ram_reg[13][199]  ( .D(n3588), .CLK(clk), .Q(\ram[13][199] ) );
  DFFX1_HVT \ram_reg[13][198]  ( .D(n3587), .CLK(clk), .Q(\ram[13][198] ) );
  DFFX1_HVT \ram_reg[13][197]  ( .D(n3586), .CLK(clk), .Q(\ram[13][197] ) );
  DFFX1_HVT \ram_reg[13][196]  ( .D(n3585), .CLK(clk), .Q(\ram[13][196] ) );
  DFFX1_HVT \ram_reg[13][195]  ( .D(n3584), .CLK(clk), .Q(\ram[13][195] ) );
  DFFX1_HVT \ram_reg[13][194]  ( .D(n3583), .CLK(clk), .Q(\ram[13][194] ) );
  DFFX1_HVT \ram_reg[13][193]  ( .D(n3582), .CLK(clk), .Q(\ram[13][193] ) );
  DFFX1_HVT \ram_reg[13][192]  ( .D(n3581), .CLK(clk), .Q(\ram[13][192] ) );
  DFFX1_HVT \ram_reg[13][191]  ( .D(n3580), .CLK(clk), .Q(\ram[13][191] ) );
  DFFX1_HVT \ram_reg[13][190]  ( .D(n3579), .CLK(clk), .Q(\ram[13][190] ) );
  DFFX1_HVT \ram_reg[13][189]  ( .D(n3578), .CLK(clk), .Q(\ram[13][189] ) );
  DFFX1_HVT \ram_reg[13][188]  ( .D(n3577), .CLK(clk), .Q(\ram[13][188] ) );
  DFFX1_HVT \ram_reg[13][187]  ( .D(n3576), .CLK(clk), .Q(\ram[13][187] ) );
  DFFX1_HVT \ram_reg[13][186]  ( .D(n3575), .CLK(clk), .Q(\ram[13][186] ) );
  DFFX1_HVT \ram_reg[13][185]  ( .D(n3574), .CLK(clk), .Q(\ram[13][185] ) );
  DFFX1_HVT \ram_reg[13][184]  ( .D(n3573), .CLK(clk), .Q(\ram[13][184] ) );
  DFFX1_HVT \ram_reg[13][183]  ( .D(n3572), .CLK(clk), .Q(\ram[13][183] ) );
  DFFX1_HVT \ram_reg[13][182]  ( .D(n3571), .CLK(clk), .Q(\ram[13][182] ) );
  DFFX1_HVT \ram_reg[13][181]  ( .D(n3570), .CLK(clk), .Q(\ram[13][181] ) );
  DFFX1_HVT \ram_reg[13][180]  ( .D(n3569), .CLK(clk), .Q(\ram[13][180] ) );
  DFFX1_HVT \ram_reg[13][179]  ( .D(n3568), .CLK(clk), .Q(\ram[13][179] ) );
  DFFX1_HVT \ram_reg[13][178]  ( .D(n3567), .CLK(clk), .Q(\ram[13][178] ) );
  DFFX1_HVT \ram_reg[13][177]  ( .D(n3566), .CLK(clk), .Q(\ram[13][177] ) );
  DFFX1_HVT \ram_reg[13][176]  ( .D(n3565), .CLK(clk), .Q(\ram[13][176] ) );
  DFFX1_HVT \ram_reg[13][175]  ( .D(n3564), .CLK(clk), .Q(\ram[13][175] ) );
  DFFX1_HVT \ram_reg[13][174]  ( .D(n3563), .CLK(clk), .Q(\ram[13][174] ) );
  DFFX1_HVT \ram_reg[13][173]  ( .D(n3562), .CLK(clk), .Q(\ram[13][173] ) );
  DFFX1_HVT \ram_reg[13][172]  ( .D(n3561), .CLK(clk), .Q(\ram[13][172] ) );
  DFFX1_HVT \ram_reg[13][171]  ( .D(n3560), .CLK(clk), .Q(\ram[13][171] ) );
  DFFX1_HVT \ram_reg[13][170]  ( .D(n3559), .CLK(clk), .Q(\ram[13][170] ) );
  DFFX1_HVT \ram_reg[13][169]  ( .D(n3558), .CLK(clk), .Q(\ram[13][169] ) );
  DFFX1_HVT \ram_reg[13][168]  ( .D(n3557), .CLK(clk), .Q(\ram[13][168] ) );
  DFFX1_HVT \ram_reg[13][167]  ( .D(n3556), .CLK(clk), .Q(\ram[13][167] ) );
  DFFX1_HVT \ram_reg[13][166]  ( .D(n3555), .CLK(clk), .Q(\ram[13][166] ) );
  DFFX1_HVT \ram_reg[13][165]  ( .D(n3554), .CLK(clk), .Q(\ram[13][165] ) );
  DFFX1_HVT \ram_reg[13][164]  ( .D(n3553), .CLK(clk), .Q(\ram[13][164] ) );
  DFFX1_HVT \ram_reg[13][163]  ( .D(n3552), .CLK(clk), .Q(\ram[13][163] ) );
  DFFX1_HVT \ram_reg[13][162]  ( .D(n3551), .CLK(clk), .Q(\ram[13][162] ) );
  DFFX1_HVT \ram_reg[13][161]  ( .D(n3550), .CLK(clk), .Q(\ram[13][161] ) );
  DFFX1_HVT \ram_reg[13][160]  ( .D(n3549), .CLK(clk), .Q(\ram[13][160] ) );
  DFFX1_HVT \ram_reg[13][159]  ( .D(n3548), .CLK(clk), .Q(\ram[13][159] ) );
  DFFX1_HVT \ram_reg[13][158]  ( .D(n3547), .CLK(clk), .Q(\ram[13][158] ) );
  DFFX1_HVT \ram_reg[13][157]  ( .D(n3546), .CLK(clk), .Q(\ram[13][157] ) );
  DFFX1_HVT \ram_reg[13][156]  ( .D(n3545), .CLK(clk), .Q(\ram[13][156] ) );
  DFFX1_HVT \ram_reg[13][155]  ( .D(n3544), .CLK(clk), .Q(\ram[13][155] ) );
  DFFX1_HVT \ram_reg[13][154]  ( .D(n3543), .CLK(clk), .Q(\ram[13][154] ) );
  DFFX1_HVT \ram_reg[13][153]  ( .D(n3542), .CLK(clk), .Q(\ram[13][153] ) );
  DFFX1_HVT \ram_reg[13][152]  ( .D(n3541), .CLK(clk), .Q(\ram[13][152] ) );
  DFFX1_HVT \ram_reg[13][151]  ( .D(n3540), .CLK(clk), .Q(\ram[13][151] ) );
  DFFX1_HVT \ram_reg[13][150]  ( .D(n3539), .CLK(clk), .Q(\ram[13][150] ) );
  DFFX1_HVT \ram_reg[13][149]  ( .D(n3538), .CLK(clk), .Q(\ram[13][149] ) );
  DFFX1_HVT \ram_reg[13][148]  ( .D(n3537), .CLK(clk), .Q(\ram[13][148] ) );
  DFFX1_HVT \ram_reg[13][147]  ( .D(n3536), .CLK(clk), .Q(\ram[13][147] ) );
  DFFX1_HVT \ram_reg[13][146]  ( .D(n3535), .CLK(clk), .Q(\ram[13][146] ) );
  DFFX1_HVT \ram_reg[13][145]  ( .D(n3534), .CLK(clk), .Q(\ram[13][145] ) );
  DFFX1_HVT \ram_reg[13][144]  ( .D(n3533), .CLK(clk), .Q(\ram[13][144] ) );
  DFFX1_HVT \ram_reg[13][143]  ( .D(n3532), .CLK(clk), .Q(\ram[13][143] ) );
  DFFX1_HVT \ram_reg[13][142]  ( .D(n3531), .CLK(clk), .Q(\ram[13][142] ) );
  DFFX1_HVT \ram_reg[13][141]  ( .D(n3530), .CLK(clk), .Q(\ram[13][141] ) );
  DFFX1_HVT \ram_reg[13][140]  ( .D(n3529), .CLK(clk), .Q(\ram[13][140] ) );
  DFFX1_HVT \ram_reg[13][139]  ( .D(n3528), .CLK(clk), .Q(\ram[13][139] ) );
  DFFX1_HVT \ram_reg[13][138]  ( .D(n3527), .CLK(clk), .Q(\ram[13][138] ) );
  DFFX1_HVT \ram_reg[13][137]  ( .D(n3526), .CLK(clk), .Q(\ram[13][137] ) );
  DFFX1_HVT \ram_reg[13][136]  ( .D(n3525), .CLK(clk), .Q(\ram[13][136] ) );
  DFFX1_HVT \ram_reg[13][135]  ( .D(n3524), .CLK(clk), .Q(\ram[13][135] ) );
  DFFX1_HVT \ram_reg[13][134]  ( .D(n3523), .CLK(clk), .Q(\ram[13][134] ) );
  DFFX1_HVT \ram_reg[13][133]  ( .D(n3522), .CLK(clk), .Q(\ram[13][133] ) );
  DFFX1_HVT \ram_reg[13][132]  ( .D(n3521), .CLK(clk), .Q(\ram[13][132] ) );
  DFFX1_HVT \ram_reg[13][131]  ( .D(n3520), .CLK(clk), .Q(\ram[13][131] ) );
  DFFX1_HVT \ram_reg[13][130]  ( .D(n3519), .CLK(clk), .Q(\ram[13][130] ) );
  DFFX1_HVT \ram_reg[13][129]  ( .D(n3518), .CLK(clk), .Q(\ram[13][129] ) );
  DFFX1_HVT \ram_reg[13][128]  ( .D(n3517), .CLK(clk), .Q(\ram[13][128] ) );
  DFFX1_HVT \ram_reg[13][127]  ( .D(n3516), .CLK(clk), .Q(\ram[13][127] ) );
  DFFX1_HVT \ram_reg[13][126]  ( .D(n3515), .CLK(clk), .Q(\ram[13][126] ) );
  DFFX1_HVT \ram_reg[13][125]  ( .D(n3514), .CLK(clk), .Q(\ram[13][125] ) );
  DFFX1_HVT \ram_reg[13][124]  ( .D(n3513), .CLK(clk), .Q(\ram[13][124] ) );
  DFFX1_HVT \ram_reg[13][123]  ( .D(n3512), .CLK(clk), .Q(\ram[13][123] ) );
  DFFX1_HVT \ram_reg[13][122]  ( .D(n3511), .CLK(clk), .Q(\ram[13][122] ) );
  DFFX1_HVT \ram_reg[13][121]  ( .D(n3510), .CLK(clk), .Q(\ram[13][121] ) );
  DFFX1_HVT \ram_reg[13][120]  ( .D(n3509), .CLK(clk), .Q(\ram[13][120] ) );
  DFFX1_HVT \ram_reg[13][119]  ( .D(n3508), .CLK(clk), .Q(\ram[13][119] ) );
  DFFX1_HVT \ram_reg[13][118]  ( .D(n3507), .CLK(clk), .Q(\ram[13][118] ) );
  DFFX1_HVT \ram_reg[13][117]  ( .D(n3506), .CLK(clk), .Q(\ram[13][117] ) );
  DFFX1_HVT \ram_reg[13][116]  ( .D(n3505), .CLK(clk), .Q(\ram[13][116] ) );
  DFFX1_HVT \ram_reg[13][115]  ( .D(n3504), .CLK(clk), .Q(\ram[13][115] ) );
  DFFX1_HVT \ram_reg[13][114]  ( .D(n3503), .CLK(clk), .Q(\ram[13][114] ) );
  DFFX1_HVT \ram_reg[13][113]  ( .D(n3502), .CLK(clk), .Q(\ram[13][113] ) );
  DFFX1_HVT \ram_reg[13][112]  ( .D(n3501), .CLK(clk), .Q(\ram[13][112] ) );
  DFFX1_HVT \ram_reg[13][111]  ( .D(n3500), .CLK(clk), .Q(\ram[13][111] ) );
  DFFX1_HVT \ram_reg[13][110]  ( .D(n3499), .CLK(clk), .Q(\ram[13][110] ) );
  DFFX1_HVT \ram_reg[13][109]  ( .D(n3498), .CLK(clk), .Q(\ram[13][109] ) );
  DFFX1_HVT \ram_reg[13][108]  ( .D(n3497), .CLK(clk), .Q(\ram[13][108] ) );
  DFFX1_HVT \ram_reg[13][107]  ( .D(n3496), .CLK(clk), .Q(\ram[13][107] ) );
  DFFX1_HVT \ram_reg[13][106]  ( .D(n3495), .CLK(clk), .Q(\ram[13][106] ) );
  DFFX1_HVT \ram_reg[13][105]  ( .D(n3494), .CLK(clk), .Q(\ram[13][105] ) );
  DFFX1_HVT \ram_reg[13][104]  ( .D(n3493), .CLK(clk), .Q(\ram[13][104] ) );
  DFFX1_HVT \ram_reg[13][103]  ( .D(n3492), .CLK(clk), .Q(\ram[13][103] ) );
  DFFX1_HVT \ram_reg[13][102]  ( .D(n3491), .CLK(clk), .Q(\ram[13][102] ) );
  DFFX1_HVT \ram_reg[13][101]  ( .D(n3490), .CLK(clk), .Q(\ram[13][101] ) );
  DFFX1_HVT \ram_reg[13][100]  ( .D(n3489), .CLK(clk), .Q(\ram[13][100] ) );
  DFFX1_HVT \ram_reg[13][99]  ( .D(n3488), .CLK(clk), .Q(\ram[13][99] ) );
  DFFX1_HVT \ram_reg[13][98]  ( .D(n3487), .CLK(clk), .Q(\ram[13][98] ) );
  DFFX1_HVT \ram_reg[13][97]  ( .D(n3486), .CLK(clk), .Q(\ram[13][97] ) );
  DFFX1_HVT \ram_reg[13][96]  ( .D(n3485), .CLK(clk), .Q(\ram[13][96] ) );
  DFFX1_HVT \ram_reg[13][95]  ( .D(n3484), .CLK(clk), .Q(\ram[13][95] ) );
  DFFX1_HVT \ram_reg[13][94]  ( .D(n3483), .CLK(clk), .Q(\ram[13][94] ) );
  DFFX1_HVT \ram_reg[13][93]  ( .D(n3482), .CLK(clk), .Q(\ram[13][93] ) );
  DFFX1_HVT \ram_reg[13][92]  ( .D(n3481), .CLK(clk), .Q(\ram[13][92] ) );
  DFFX1_HVT \ram_reg[13][91]  ( .D(n3480), .CLK(clk), .Q(\ram[13][91] ) );
  DFFX1_HVT \ram_reg[13][90]  ( .D(n3479), .CLK(clk), .Q(\ram[13][90] ) );
  DFFX1_HVT \ram_reg[13][89]  ( .D(n3478), .CLK(clk), .Q(\ram[13][89] ) );
  DFFX1_HVT \ram_reg[13][88]  ( .D(n3477), .CLK(clk), .Q(\ram[13][88] ) );
  DFFX1_HVT \ram_reg[13][87]  ( .D(n3476), .CLK(clk), .Q(\ram[13][87] ) );
  DFFX1_HVT \ram_reg[13][86]  ( .D(n3475), .CLK(clk), .Q(\ram[13][86] ) );
  DFFX1_HVT \ram_reg[13][85]  ( .D(n3474), .CLK(clk), .Q(\ram[13][85] ) );
  DFFX1_HVT \ram_reg[13][84]  ( .D(n3473), .CLK(clk), .Q(\ram[13][84] ) );
  DFFX1_HVT \ram_reg[13][83]  ( .D(n3472), .CLK(clk), .Q(\ram[13][83] ) );
  DFFX1_HVT \ram_reg[13][82]  ( .D(n3471), .CLK(clk), .Q(\ram[13][82] ) );
  DFFX1_HVT \ram_reg[13][81]  ( .D(n3470), .CLK(clk), .Q(\ram[13][81] ) );
  DFFX1_HVT \ram_reg[13][80]  ( .D(n3469), .CLK(clk), .Q(\ram[13][80] ) );
  DFFX1_HVT \ram_reg[13][79]  ( .D(n3468), .CLK(clk), .Q(\ram[13][79] ) );
  DFFX1_HVT \ram_reg[13][78]  ( .D(n3467), .CLK(clk), .Q(\ram[13][78] ) );
  DFFX1_HVT \ram_reg[13][77]  ( .D(n3466), .CLK(clk), .Q(\ram[13][77] ) );
  DFFX1_HVT \ram_reg[13][76]  ( .D(n3465), .CLK(clk), .Q(\ram[13][76] ) );
  DFFX1_HVT \ram_reg[13][75]  ( .D(n3464), .CLK(clk), .Q(\ram[13][75] ) );
  DFFX1_HVT \ram_reg[13][74]  ( .D(n3463), .CLK(clk), .Q(\ram[13][74] ) );
  DFFX1_HVT \ram_reg[13][73]  ( .D(n3462), .CLK(clk), .Q(\ram[13][73] ) );
  DFFX1_HVT \ram_reg[13][72]  ( .D(n3461), .CLK(clk), .Q(\ram[13][72] ) );
  DFFX1_HVT \ram_reg[13][71]  ( .D(n3460), .CLK(clk), .Q(\ram[13][71] ) );
  DFFX1_HVT \ram_reg[13][70]  ( .D(n3459), .CLK(clk), .Q(\ram[13][70] ) );
  DFFX1_HVT \ram_reg[13][69]  ( .D(n3458), .CLK(clk), .Q(\ram[13][69] ) );
  DFFX1_HVT \ram_reg[13][68]  ( .D(n3457), .CLK(clk), .Q(\ram[13][68] ) );
  DFFX1_HVT \ram_reg[13][67]  ( .D(n3456), .CLK(clk), .Q(\ram[13][67] ) );
  DFFX1_HVT \ram_reg[13][66]  ( .D(n3455), .CLK(clk), .Q(\ram[13][66] ) );
  DFFX1_HVT \ram_reg[13][65]  ( .D(n3454), .CLK(clk), .Q(\ram[13][65] ) );
  DFFX1_HVT \ram_reg[13][64]  ( .D(n3453), .CLK(clk), .Q(\ram[13][64] ) );
  DFFX1_HVT \ram_reg[13][63]  ( .D(n3452), .CLK(clk), .Q(\ram[13][63] ) );
  DFFX1_HVT \ram_reg[13][62]  ( .D(n3451), .CLK(clk), .Q(\ram[13][62] ) );
  DFFX1_HVT \ram_reg[13][61]  ( .D(n3450), .CLK(clk), .Q(\ram[13][61] ) );
  DFFX1_HVT \ram_reg[13][60]  ( .D(n3449), .CLK(clk), .Q(\ram[13][60] ) );
  DFFX1_HVT \ram_reg[13][59]  ( .D(n3448), .CLK(clk), .Q(\ram[13][59] ) );
  DFFX1_HVT \ram_reg[13][58]  ( .D(n3447), .CLK(clk), .Q(\ram[13][58] ) );
  DFFX1_HVT \ram_reg[13][57]  ( .D(n3446), .CLK(clk), .Q(\ram[13][57] ) );
  DFFX1_HVT \ram_reg[13][56]  ( .D(n3445), .CLK(clk), .Q(\ram[13][56] ) );
  DFFX1_HVT \ram_reg[13][55]  ( .D(n3444), .CLK(clk), .Q(\ram[13][55] ) );
  DFFX1_HVT \ram_reg[13][54]  ( .D(n3443), .CLK(clk), .Q(\ram[13][54] ) );
  DFFX1_HVT \ram_reg[13][53]  ( .D(n3442), .CLK(clk), .Q(\ram[13][53] ) );
  DFFX1_HVT \ram_reg[13][52]  ( .D(n3441), .CLK(clk), .Q(\ram[13][52] ) );
  DFFX1_HVT \ram_reg[13][51]  ( .D(n3440), .CLK(clk), .Q(\ram[13][51] ) );
  DFFX1_HVT \ram_reg[13][50]  ( .D(n3439), .CLK(clk), .Q(\ram[13][50] ) );
  DFFX1_HVT \ram_reg[13][49]  ( .D(n3438), .CLK(clk), .Q(\ram[13][49] ) );
  DFFX1_HVT \ram_reg[13][48]  ( .D(n3437), .CLK(clk), .Q(\ram[13][48] ) );
  DFFX1_HVT \ram_reg[13][47]  ( .D(n3436), .CLK(clk), .Q(\ram[13][47] ) );
  DFFX1_HVT \ram_reg[13][46]  ( .D(n3435), .CLK(clk), .Q(\ram[13][46] ) );
  DFFX1_HVT \ram_reg[13][45]  ( .D(n3434), .CLK(clk), .Q(\ram[13][45] ) );
  DFFX1_HVT \ram_reg[13][44]  ( .D(n3433), .CLK(clk), .Q(\ram[13][44] ) );
  DFFX1_HVT \ram_reg[13][43]  ( .D(n3432), .CLK(clk), .Q(\ram[13][43] ) );
  DFFX1_HVT \ram_reg[13][42]  ( .D(n3431), .CLK(clk), .Q(\ram[13][42] ) );
  DFFX1_HVT \ram_reg[13][41]  ( .D(n3430), .CLK(clk), .Q(\ram[13][41] ) );
  DFFX1_HVT \ram_reg[13][40]  ( .D(n3429), .CLK(clk), .Q(\ram[13][40] ) );
  DFFX1_HVT \ram_reg[13][39]  ( .D(n3428), .CLK(clk), .Q(\ram[13][39] ) );
  DFFX1_HVT \ram_reg[13][38]  ( .D(n3427), .CLK(clk), .Q(\ram[13][38] ) );
  DFFX1_HVT \ram_reg[13][37]  ( .D(n3426), .CLK(clk), .Q(\ram[13][37] ) );
  DFFX1_HVT \ram_reg[13][36]  ( .D(n3425), .CLK(clk), .Q(\ram[13][36] ) );
  DFFX1_HVT \ram_reg[13][35]  ( .D(n3424), .CLK(clk), .Q(\ram[13][35] ) );
  DFFX1_HVT \ram_reg[13][34]  ( .D(n3423), .CLK(clk), .Q(\ram[13][34] ) );
  DFFX1_HVT \ram_reg[13][33]  ( .D(n3422), .CLK(clk), .Q(\ram[13][33] ) );
  DFFX1_HVT \ram_reg[13][32]  ( .D(n3421), .CLK(clk), .Q(\ram[13][32] ) );
  DFFX1_HVT \ram_reg[13][31]  ( .D(n3420), .CLK(clk), .Q(\ram[13][31] ) );
  DFFX1_HVT \ram_reg[13][30]  ( .D(n3419), .CLK(clk), .Q(\ram[13][30] ) );
  DFFX1_HVT \ram_reg[13][29]  ( .D(n3418), .CLK(clk), .Q(\ram[13][29] ) );
  DFFX1_HVT \ram_reg[13][28]  ( .D(n3417), .CLK(clk), .Q(\ram[13][28] ) );
  DFFX1_HVT \ram_reg[13][27]  ( .D(n3416), .CLK(clk), .Q(\ram[13][27] ) );
  DFFX1_HVT \ram_reg[13][26]  ( .D(n3415), .CLK(clk), .Q(\ram[13][26] ) );
  DFFX1_HVT \ram_reg[13][25]  ( .D(n3414), .CLK(clk), .Q(\ram[13][25] ) );
  DFFX1_HVT \ram_reg[13][24]  ( .D(n3413), .CLK(clk), .Q(\ram[13][24] ) );
  DFFX1_HVT \ram_reg[13][23]  ( .D(n3412), .CLK(clk), .Q(\ram[13][23] ) );
  DFFX1_HVT \ram_reg[13][22]  ( .D(n3411), .CLK(clk), .Q(\ram[13][22] ) );
  DFFX1_HVT \ram_reg[13][21]  ( .D(n3410), .CLK(clk), .Q(\ram[13][21] ) );
  DFFX1_HVT \ram_reg[13][20]  ( .D(n3409), .CLK(clk), .Q(\ram[13][20] ) );
  DFFX1_HVT \ram_reg[13][19]  ( .D(n3408), .CLK(clk), .Q(\ram[13][19] ) );
  DFFX1_HVT \ram_reg[13][18]  ( .D(n3407), .CLK(clk), .Q(\ram[13][18] ) );
  DFFX1_HVT \ram_reg[13][17]  ( .D(n3406), .CLK(clk), .Q(\ram[13][17] ) );
  DFFX1_HVT \ram_reg[13][16]  ( .D(n3405), .CLK(clk), .Q(\ram[13][16] ) );
  DFFX1_HVT \ram_reg[13][15]  ( .D(n3404), .CLK(clk), .Q(\ram[13][15] ) );
  DFFX1_HVT \ram_reg[13][14]  ( .D(n3403), .CLK(clk), .Q(\ram[13][14] ) );
  DFFX1_HVT \ram_reg[13][13]  ( .D(n3402), .CLK(clk), .Q(\ram[13][13] ) );
  DFFX1_HVT \ram_reg[13][12]  ( .D(n3401), .CLK(clk), .Q(\ram[13][12] ) );
  DFFX1_HVT \ram_reg[13][11]  ( .D(n3400), .CLK(clk), .Q(\ram[13][11] ) );
  DFFX1_HVT \ram_reg[13][10]  ( .D(n3399), .CLK(clk), .Q(\ram[13][10] ) );
  DFFX1_HVT \ram_reg[13][9]  ( .D(n3398), .CLK(clk), .Q(\ram[13][9] ) );
  DFFX1_HVT \ram_reg[13][8]  ( .D(n3397), .CLK(clk), .Q(\ram[13][8] ) );
  DFFX1_HVT \ram_reg[13][7]  ( .D(n3396), .CLK(clk), .Q(\ram[13][7] ) );
  DFFX1_HVT \ram_reg[13][6]  ( .D(n3395), .CLK(clk), .Q(\ram[13][6] ) );
  DFFX1_HVT \ram_reg[13][5]  ( .D(n3394), .CLK(clk), .Q(\ram[13][5] ) );
  DFFX1_HVT \ram_reg[13][4]  ( .D(n3393), .CLK(clk), .Q(\ram[13][4] ) );
  DFFX1_HVT \ram_reg[13][3]  ( .D(n3392), .CLK(clk), .Q(\ram[13][3] ) );
  DFFX1_HVT \ram_reg[13][2]  ( .D(n3391), .CLK(clk), .Q(\ram[13][2] ) );
  DFFX1_HVT \ram_reg[13][1]  ( .D(n3390), .CLK(clk), .Q(\ram[13][1] ) );
  DFFX1_HVT \ram_reg[13][0]  ( .D(n3389), .CLK(clk), .Q(\ram[13][0] ) );
  DFFX1_HVT \ram_reg[12][255]  ( .D(n3388), .CLK(clk), .Q(\ram[12][255] ) );
  DFFX1_HVT \ram_reg[12][254]  ( .D(n3387), .CLK(clk), .Q(\ram[12][254] ) );
  DFFX1_HVT \ram_reg[12][253]  ( .D(n3386), .CLK(clk), .Q(\ram[12][253] ) );
  DFFX1_HVT \ram_reg[12][252]  ( .D(n3385), .CLK(clk), .Q(\ram[12][252] ) );
  DFFX1_HVT \ram_reg[12][251]  ( .D(n3384), .CLK(clk), .Q(\ram[12][251] ) );
  DFFX1_HVT \ram_reg[12][250]  ( .D(n3383), .CLK(clk), .Q(\ram[12][250] ) );
  DFFX1_HVT \ram_reg[12][249]  ( .D(n3382), .CLK(clk), .Q(\ram[12][249] ) );
  DFFX1_HVT \ram_reg[12][248]  ( .D(n3381), .CLK(clk), .Q(\ram[12][248] ) );
  DFFX1_HVT \ram_reg[12][247]  ( .D(n3380), .CLK(clk), .Q(\ram[12][247] ) );
  DFFX1_HVT \ram_reg[12][246]  ( .D(n3379), .CLK(clk), .Q(\ram[12][246] ) );
  DFFX1_HVT \ram_reg[12][245]  ( .D(n3378), .CLK(clk), .Q(\ram[12][245] ) );
  DFFX1_HVT \ram_reg[12][244]  ( .D(n3377), .CLK(clk), .Q(\ram[12][244] ) );
  DFFX1_HVT \ram_reg[12][243]  ( .D(n3376), .CLK(clk), .Q(\ram[12][243] ) );
  DFFX1_HVT \ram_reg[12][242]  ( .D(n3375), .CLK(clk), .Q(\ram[12][242] ) );
  DFFX1_HVT \ram_reg[12][241]  ( .D(n3374), .CLK(clk), .Q(\ram[12][241] ) );
  DFFX1_HVT \ram_reg[12][240]  ( .D(n3373), .CLK(clk), .Q(\ram[12][240] ) );
  DFFX1_HVT \ram_reg[12][239]  ( .D(n3372), .CLK(clk), .Q(\ram[12][239] ) );
  DFFX1_HVT \ram_reg[12][238]  ( .D(n3371), .CLK(clk), .Q(\ram[12][238] ) );
  DFFX1_HVT \ram_reg[12][237]  ( .D(n3370), .CLK(clk), .Q(\ram[12][237] ) );
  DFFX1_HVT \ram_reg[12][236]  ( .D(n3369), .CLK(clk), .Q(\ram[12][236] ) );
  DFFX1_HVT \ram_reg[12][235]  ( .D(n3368), .CLK(clk), .Q(\ram[12][235] ) );
  DFFX1_HVT \ram_reg[12][234]  ( .D(n3367), .CLK(clk), .Q(\ram[12][234] ) );
  DFFX1_HVT \ram_reg[12][233]  ( .D(n3366), .CLK(clk), .Q(\ram[12][233] ) );
  DFFX1_HVT \ram_reg[12][232]  ( .D(n3365), .CLK(clk), .Q(\ram[12][232] ) );
  DFFX1_HVT \ram_reg[12][231]  ( .D(n3364), .CLK(clk), .Q(\ram[12][231] ) );
  DFFX1_HVT \ram_reg[12][230]  ( .D(n3363), .CLK(clk), .Q(\ram[12][230] ) );
  DFFX1_HVT \ram_reg[12][229]  ( .D(n3362), .CLK(clk), .Q(\ram[12][229] ) );
  DFFX1_HVT \ram_reg[12][228]  ( .D(n3361), .CLK(clk), .Q(\ram[12][228] ) );
  DFFX1_HVT \ram_reg[12][227]  ( .D(n3360), .CLK(clk), .Q(\ram[12][227] ) );
  DFFX1_HVT \ram_reg[12][226]  ( .D(n3359), .CLK(clk), .Q(\ram[12][226] ) );
  DFFX1_HVT \ram_reg[12][225]  ( .D(n3358), .CLK(clk), .Q(\ram[12][225] ) );
  DFFX1_HVT \ram_reg[12][224]  ( .D(n3357), .CLK(clk), .Q(\ram[12][224] ) );
  DFFX1_HVT \ram_reg[12][223]  ( .D(n3356), .CLK(clk), .Q(\ram[12][223] ) );
  DFFX1_HVT \ram_reg[12][222]  ( .D(n3355), .CLK(clk), .Q(\ram[12][222] ) );
  DFFX1_HVT \ram_reg[12][221]  ( .D(n3354), .CLK(clk), .Q(\ram[12][221] ) );
  DFFX1_HVT \ram_reg[12][220]  ( .D(n3353), .CLK(clk), .Q(\ram[12][220] ) );
  DFFX1_HVT \ram_reg[12][219]  ( .D(n3352), .CLK(clk), .Q(\ram[12][219] ) );
  DFFX1_HVT \ram_reg[12][218]  ( .D(n3351), .CLK(clk), .Q(\ram[12][218] ) );
  DFFX1_HVT \ram_reg[12][217]  ( .D(n3350), .CLK(clk), .Q(\ram[12][217] ) );
  DFFX1_HVT \ram_reg[12][216]  ( .D(n3349), .CLK(clk), .Q(\ram[12][216] ) );
  DFFX1_HVT \ram_reg[12][215]  ( .D(n3348), .CLK(clk), .Q(\ram[12][215] ) );
  DFFX1_HVT \ram_reg[12][214]  ( .D(n3347), .CLK(clk), .Q(\ram[12][214] ) );
  DFFX1_HVT \ram_reg[12][213]  ( .D(n3346), .CLK(clk), .Q(\ram[12][213] ) );
  DFFX1_HVT \ram_reg[12][212]  ( .D(n3345), .CLK(clk), .Q(\ram[12][212] ) );
  DFFX1_HVT \ram_reg[12][211]  ( .D(n3344), .CLK(clk), .Q(\ram[12][211] ) );
  DFFX1_HVT \ram_reg[12][210]  ( .D(n3343), .CLK(clk), .Q(\ram[12][210] ) );
  DFFX1_HVT \ram_reg[12][209]  ( .D(n3342), .CLK(clk), .Q(\ram[12][209] ) );
  DFFX1_HVT \ram_reg[12][208]  ( .D(n3341), .CLK(clk), .Q(\ram[12][208] ) );
  DFFX1_HVT \ram_reg[12][207]  ( .D(n3340), .CLK(clk), .Q(\ram[12][207] ) );
  DFFX1_HVT \ram_reg[12][206]  ( .D(n3339), .CLK(clk), .Q(\ram[12][206] ) );
  DFFX1_HVT \ram_reg[12][205]  ( .D(n3338), .CLK(clk), .Q(\ram[12][205] ) );
  DFFX1_HVT \ram_reg[12][204]  ( .D(n3337), .CLK(clk), .Q(\ram[12][204] ) );
  DFFX1_HVT \ram_reg[12][203]  ( .D(n3336), .CLK(clk), .Q(\ram[12][203] ) );
  DFFX1_HVT \ram_reg[12][202]  ( .D(n3335), .CLK(clk), .Q(\ram[12][202] ) );
  DFFX1_HVT \ram_reg[12][201]  ( .D(n3334), .CLK(clk), .Q(\ram[12][201] ) );
  DFFX1_HVT \ram_reg[12][200]  ( .D(n3333), .CLK(clk), .Q(\ram[12][200] ) );
  DFFX1_HVT \ram_reg[12][199]  ( .D(n3332), .CLK(clk), .Q(\ram[12][199] ) );
  DFFX1_HVT \ram_reg[12][198]  ( .D(n3331), .CLK(clk), .Q(\ram[12][198] ) );
  DFFX1_HVT \ram_reg[12][197]  ( .D(n3330), .CLK(clk), .Q(\ram[12][197] ) );
  DFFX1_HVT \ram_reg[12][196]  ( .D(n3329), .CLK(clk), .Q(\ram[12][196] ) );
  DFFX1_HVT \ram_reg[12][195]  ( .D(n3328), .CLK(clk), .Q(\ram[12][195] ) );
  DFFX1_HVT \ram_reg[12][194]  ( .D(n3327), .CLK(clk), .Q(\ram[12][194] ) );
  DFFX1_HVT \ram_reg[12][193]  ( .D(n3326), .CLK(clk), .Q(\ram[12][193] ) );
  DFFX1_HVT \ram_reg[12][192]  ( .D(n3325), .CLK(clk), .Q(\ram[12][192] ) );
  DFFX1_HVT \ram_reg[12][191]  ( .D(n3324), .CLK(clk), .Q(\ram[12][191] ) );
  DFFX1_HVT \ram_reg[12][190]  ( .D(n3323), .CLK(clk), .Q(\ram[12][190] ) );
  DFFX1_HVT \ram_reg[12][189]  ( .D(n3322), .CLK(clk), .Q(\ram[12][189] ) );
  DFFX1_HVT \ram_reg[12][188]  ( .D(n3321), .CLK(clk), .Q(\ram[12][188] ) );
  DFFX1_HVT \ram_reg[12][187]  ( .D(n3320), .CLK(clk), .Q(\ram[12][187] ) );
  DFFX1_HVT \ram_reg[12][186]  ( .D(n3319), .CLK(clk), .Q(\ram[12][186] ) );
  DFFX1_HVT \ram_reg[12][185]  ( .D(n3318), .CLK(clk), .Q(\ram[12][185] ) );
  DFFX1_HVT \ram_reg[12][184]  ( .D(n3317), .CLK(clk), .Q(\ram[12][184] ) );
  DFFX1_HVT \ram_reg[12][183]  ( .D(n3316), .CLK(clk), .Q(\ram[12][183] ) );
  DFFX1_HVT \ram_reg[12][182]  ( .D(n3315), .CLK(clk), .Q(\ram[12][182] ) );
  DFFX1_HVT \ram_reg[12][181]  ( .D(n3314), .CLK(clk), .Q(\ram[12][181] ) );
  DFFX1_HVT \ram_reg[12][180]  ( .D(n3313), .CLK(clk), .Q(\ram[12][180] ) );
  DFFX1_HVT \ram_reg[12][179]  ( .D(n3312), .CLK(clk), .Q(\ram[12][179] ) );
  DFFX1_HVT \ram_reg[12][178]  ( .D(n3311), .CLK(clk), .Q(\ram[12][178] ) );
  DFFX1_HVT \ram_reg[12][177]  ( .D(n3310), .CLK(clk), .Q(\ram[12][177] ) );
  DFFX1_HVT \ram_reg[12][176]  ( .D(n3309), .CLK(clk), .Q(\ram[12][176] ) );
  DFFX1_HVT \ram_reg[12][175]  ( .D(n3308), .CLK(clk), .Q(\ram[12][175] ) );
  DFFX1_HVT \ram_reg[12][174]  ( .D(n3307), .CLK(clk), .Q(\ram[12][174] ) );
  DFFX1_HVT \ram_reg[12][173]  ( .D(n3306), .CLK(clk), .Q(\ram[12][173] ) );
  DFFX1_HVT \ram_reg[12][172]  ( .D(n3305), .CLK(clk), .Q(\ram[12][172] ) );
  DFFX1_HVT \ram_reg[12][171]  ( .D(n3304), .CLK(clk), .Q(\ram[12][171] ) );
  DFFX1_HVT \ram_reg[12][170]  ( .D(n3303), .CLK(clk), .Q(\ram[12][170] ) );
  DFFX1_HVT \ram_reg[12][169]  ( .D(n3302), .CLK(clk), .Q(\ram[12][169] ) );
  DFFX1_HVT \ram_reg[12][168]  ( .D(n3301), .CLK(clk), .Q(\ram[12][168] ) );
  DFFX1_HVT \ram_reg[12][167]  ( .D(n3300), .CLK(clk), .Q(\ram[12][167] ) );
  DFFX1_HVT \ram_reg[12][166]  ( .D(n3299), .CLK(clk), .Q(\ram[12][166] ) );
  DFFX1_HVT \ram_reg[12][165]  ( .D(n3298), .CLK(clk), .Q(\ram[12][165] ) );
  DFFX1_HVT \ram_reg[12][164]  ( .D(n3297), .CLK(clk), .Q(\ram[12][164] ) );
  DFFX1_HVT \ram_reg[12][163]  ( .D(n3296), .CLK(clk), .Q(\ram[12][163] ) );
  DFFX1_HVT \ram_reg[12][162]  ( .D(n3295), .CLK(clk), .Q(\ram[12][162] ) );
  DFFX1_HVT \ram_reg[12][161]  ( .D(n3294), .CLK(clk), .Q(\ram[12][161] ) );
  DFFX1_HVT \ram_reg[12][160]  ( .D(n3293), .CLK(clk), .Q(\ram[12][160] ) );
  DFFX1_HVT \ram_reg[12][159]  ( .D(n3292), .CLK(clk), .Q(\ram[12][159] ) );
  DFFX1_HVT \ram_reg[12][158]  ( .D(n3291), .CLK(clk), .Q(\ram[12][158] ) );
  DFFX1_HVT \ram_reg[12][157]  ( .D(n3290), .CLK(clk), .Q(\ram[12][157] ) );
  DFFX1_HVT \ram_reg[12][156]  ( .D(n3289), .CLK(clk), .Q(\ram[12][156] ) );
  DFFX1_HVT \ram_reg[12][155]  ( .D(n3288), .CLK(clk), .Q(\ram[12][155] ) );
  DFFX1_HVT \ram_reg[12][154]  ( .D(n3287), .CLK(clk), .Q(\ram[12][154] ) );
  DFFX1_HVT \ram_reg[12][153]  ( .D(n3286), .CLK(clk), .Q(\ram[12][153] ) );
  DFFX1_HVT \ram_reg[12][152]  ( .D(n3285), .CLK(clk), .Q(\ram[12][152] ) );
  DFFX1_HVT \ram_reg[12][151]  ( .D(n3284), .CLK(clk), .Q(\ram[12][151] ) );
  DFFX1_HVT \ram_reg[12][150]  ( .D(n3283), .CLK(clk), .Q(\ram[12][150] ) );
  DFFX1_HVT \ram_reg[12][149]  ( .D(n3282), .CLK(clk), .Q(\ram[12][149] ) );
  DFFX1_HVT \ram_reg[12][148]  ( .D(n3281), .CLK(clk), .Q(\ram[12][148] ) );
  DFFX1_HVT \ram_reg[12][147]  ( .D(n3280), .CLK(clk), .Q(\ram[12][147] ) );
  DFFX1_HVT \ram_reg[12][146]  ( .D(n3279), .CLK(clk), .Q(\ram[12][146] ) );
  DFFX1_HVT \ram_reg[12][145]  ( .D(n3278), .CLK(clk), .Q(\ram[12][145] ) );
  DFFX1_HVT \ram_reg[12][144]  ( .D(n3277), .CLK(clk), .Q(\ram[12][144] ) );
  DFFX1_HVT \ram_reg[12][143]  ( .D(n3276), .CLK(clk), .Q(\ram[12][143] ) );
  DFFX1_HVT \ram_reg[12][142]  ( .D(n3275), .CLK(clk), .Q(\ram[12][142] ) );
  DFFX1_HVT \ram_reg[12][141]  ( .D(n3274), .CLK(clk), .Q(\ram[12][141] ) );
  DFFX1_HVT \ram_reg[12][140]  ( .D(n3273), .CLK(clk), .Q(\ram[12][140] ) );
  DFFX1_HVT \ram_reg[12][139]  ( .D(n3272), .CLK(clk), .Q(\ram[12][139] ) );
  DFFX1_HVT \ram_reg[12][138]  ( .D(n3271), .CLK(clk), .Q(\ram[12][138] ) );
  DFFX1_HVT \ram_reg[12][137]  ( .D(n3270), .CLK(clk), .Q(\ram[12][137] ) );
  DFFX1_HVT \ram_reg[12][136]  ( .D(n3269), .CLK(clk), .Q(\ram[12][136] ) );
  DFFX1_HVT \ram_reg[12][135]  ( .D(n3268), .CLK(clk), .Q(\ram[12][135] ) );
  DFFX1_HVT \ram_reg[12][134]  ( .D(n3267), .CLK(clk), .Q(\ram[12][134] ) );
  DFFX1_HVT \ram_reg[12][133]  ( .D(n3266), .CLK(clk), .Q(\ram[12][133] ) );
  DFFX1_HVT \ram_reg[12][132]  ( .D(n3265), .CLK(clk), .Q(\ram[12][132] ) );
  DFFX1_HVT \ram_reg[12][131]  ( .D(n3264), .CLK(clk), .Q(\ram[12][131] ) );
  DFFX1_HVT \ram_reg[12][130]  ( .D(n3263), .CLK(clk), .Q(\ram[12][130] ) );
  DFFX1_HVT \ram_reg[12][129]  ( .D(n3262), .CLK(clk), .Q(\ram[12][129] ) );
  DFFX1_HVT \ram_reg[12][128]  ( .D(n3261), .CLK(clk), .Q(\ram[12][128] ) );
  DFFX1_HVT \ram_reg[12][127]  ( .D(n3260), .CLK(clk), .Q(\ram[12][127] ) );
  DFFX1_HVT \ram_reg[12][126]  ( .D(n3259), .CLK(clk), .Q(\ram[12][126] ) );
  DFFX1_HVT \ram_reg[12][125]  ( .D(n3258), .CLK(clk), .Q(\ram[12][125] ) );
  DFFX1_HVT \ram_reg[12][124]  ( .D(n3257), .CLK(clk), .Q(\ram[12][124] ) );
  DFFX1_HVT \ram_reg[12][123]  ( .D(n3256), .CLK(clk), .Q(\ram[12][123] ) );
  DFFX1_HVT \ram_reg[12][122]  ( .D(n3255), .CLK(clk), .Q(\ram[12][122] ) );
  DFFX1_HVT \ram_reg[12][121]  ( .D(n3254), .CLK(clk), .Q(\ram[12][121] ) );
  DFFX1_HVT \ram_reg[12][120]  ( .D(n3253), .CLK(clk), .Q(\ram[12][120] ) );
  DFFX1_HVT \ram_reg[12][119]  ( .D(n3252), .CLK(clk), .Q(\ram[12][119] ) );
  DFFX1_HVT \ram_reg[12][118]  ( .D(n3251), .CLK(clk), .Q(\ram[12][118] ) );
  DFFX1_HVT \ram_reg[12][117]  ( .D(n3250), .CLK(clk), .Q(\ram[12][117] ) );
  DFFX1_HVT \ram_reg[12][116]  ( .D(n3249), .CLK(clk), .Q(\ram[12][116] ) );
  DFFX1_HVT \ram_reg[12][115]  ( .D(n3248), .CLK(clk), .Q(\ram[12][115] ) );
  DFFX1_HVT \ram_reg[12][114]  ( .D(n3247), .CLK(clk), .Q(\ram[12][114] ) );
  DFFX1_HVT \ram_reg[12][113]  ( .D(n3246), .CLK(clk), .Q(\ram[12][113] ) );
  DFFX1_HVT \ram_reg[12][112]  ( .D(n3245), .CLK(clk), .Q(\ram[12][112] ) );
  DFFX1_HVT \ram_reg[12][111]  ( .D(n3244), .CLK(clk), .Q(\ram[12][111] ) );
  DFFX1_HVT \ram_reg[12][110]  ( .D(n3243), .CLK(clk), .Q(\ram[12][110] ) );
  DFFX1_HVT \ram_reg[12][109]  ( .D(n3242), .CLK(clk), .Q(\ram[12][109] ) );
  DFFX1_HVT \ram_reg[12][108]  ( .D(n3241), .CLK(clk), .Q(\ram[12][108] ) );
  DFFX1_HVT \ram_reg[12][107]  ( .D(n3240), .CLK(clk), .Q(\ram[12][107] ) );
  DFFX1_HVT \ram_reg[12][106]  ( .D(n3239), .CLK(clk), .Q(\ram[12][106] ) );
  DFFX1_HVT \ram_reg[12][105]  ( .D(n3238), .CLK(clk), .Q(\ram[12][105] ) );
  DFFX1_HVT \ram_reg[12][104]  ( .D(n3237), .CLK(clk), .Q(\ram[12][104] ) );
  DFFX1_HVT \ram_reg[12][103]  ( .D(n3236), .CLK(clk), .Q(\ram[12][103] ) );
  DFFX1_HVT \ram_reg[12][102]  ( .D(n3235), .CLK(clk), .Q(\ram[12][102] ) );
  DFFX1_HVT \ram_reg[12][101]  ( .D(n3234), .CLK(clk), .Q(\ram[12][101] ) );
  DFFX1_HVT \ram_reg[12][100]  ( .D(n3233), .CLK(clk), .Q(\ram[12][100] ) );
  DFFX1_HVT \ram_reg[12][99]  ( .D(n3232), .CLK(clk), .Q(\ram[12][99] ) );
  DFFX1_HVT \ram_reg[12][98]  ( .D(n3231), .CLK(clk), .Q(\ram[12][98] ) );
  DFFX1_HVT \ram_reg[12][97]  ( .D(n3230), .CLK(clk), .Q(\ram[12][97] ) );
  DFFX1_HVT \ram_reg[12][96]  ( .D(n3229), .CLK(clk), .Q(\ram[12][96] ) );
  DFFX1_HVT \ram_reg[12][95]  ( .D(n3228), .CLK(clk), .Q(\ram[12][95] ) );
  DFFX1_HVT \ram_reg[12][94]  ( .D(n3227), .CLK(clk), .Q(\ram[12][94] ) );
  DFFX1_HVT \ram_reg[12][93]  ( .D(n3226), .CLK(clk), .Q(\ram[12][93] ) );
  DFFX1_HVT \ram_reg[12][92]  ( .D(n3225), .CLK(clk), .Q(\ram[12][92] ) );
  DFFX1_HVT \ram_reg[12][91]  ( .D(n3224), .CLK(clk), .Q(\ram[12][91] ) );
  DFFX1_HVT \ram_reg[12][90]  ( .D(n3223), .CLK(clk), .Q(\ram[12][90] ) );
  DFFX1_HVT \ram_reg[12][89]  ( .D(n3222), .CLK(clk), .Q(\ram[12][89] ) );
  DFFX1_HVT \ram_reg[12][88]  ( .D(n3221), .CLK(clk), .Q(\ram[12][88] ) );
  DFFX1_HVT \ram_reg[12][87]  ( .D(n3220), .CLK(clk), .Q(\ram[12][87] ) );
  DFFX1_HVT \ram_reg[12][86]  ( .D(n3219), .CLK(clk), .Q(\ram[12][86] ) );
  DFFX1_HVT \ram_reg[12][85]  ( .D(n3218), .CLK(clk), .Q(\ram[12][85] ) );
  DFFX1_HVT \ram_reg[12][84]  ( .D(n3217), .CLK(clk), .Q(\ram[12][84] ) );
  DFFX1_HVT \ram_reg[12][83]  ( .D(n3216), .CLK(clk), .Q(\ram[12][83] ) );
  DFFX1_HVT \ram_reg[12][82]  ( .D(n3215), .CLK(clk), .Q(\ram[12][82] ) );
  DFFX1_HVT \ram_reg[12][81]  ( .D(n3214), .CLK(clk), .Q(\ram[12][81] ) );
  DFFX1_HVT \ram_reg[12][80]  ( .D(n3213), .CLK(clk), .Q(\ram[12][80] ) );
  DFFX1_HVT \ram_reg[12][79]  ( .D(n3212), .CLK(clk), .Q(\ram[12][79] ) );
  DFFX1_HVT \ram_reg[12][78]  ( .D(n3211), .CLK(clk), .Q(\ram[12][78] ) );
  DFFX1_HVT \ram_reg[12][77]  ( .D(n3210), .CLK(clk), .Q(\ram[12][77] ) );
  DFFX1_HVT \ram_reg[12][76]  ( .D(n3209), .CLK(clk), .Q(\ram[12][76] ) );
  DFFX1_HVT \ram_reg[12][75]  ( .D(n3208), .CLK(clk), .Q(\ram[12][75] ) );
  DFFX1_HVT \ram_reg[12][74]  ( .D(n3207), .CLK(clk), .Q(\ram[12][74] ) );
  DFFX1_HVT \ram_reg[12][73]  ( .D(n3206), .CLK(clk), .Q(\ram[12][73] ) );
  DFFX1_HVT \ram_reg[12][72]  ( .D(n3205), .CLK(clk), .Q(\ram[12][72] ) );
  DFFX1_HVT \ram_reg[12][71]  ( .D(n3204), .CLK(clk), .Q(\ram[12][71] ) );
  DFFX1_HVT \ram_reg[12][70]  ( .D(n3203), .CLK(clk), .Q(\ram[12][70] ) );
  DFFX1_HVT \ram_reg[12][69]  ( .D(n3202), .CLK(clk), .Q(\ram[12][69] ) );
  DFFX1_HVT \ram_reg[12][68]  ( .D(n3201), .CLK(clk), .Q(\ram[12][68] ) );
  DFFX1_HVT \ram_reg[12][67]  ( .D(n3200), .CLK(clk), .Q(\ram[12][67] ) );
  DFFX1_HVT \ram_reg[12][66]  ( .D(n3199), .CLK(clk), .Q(\ram[12][66] ) );
  DFFX1_HVT \ram_reg[12][65]  ( .D(n3198), .CLK(clk), .Q(\ram[12][65] ) );
  DFFX1_HVT \ram_reg[12][64]  ( .D(n3197), .CLK(clk), .Q(\ram[12][64] ) );
  DFFX1_HVT \ram_reg[12][63]  ( .D(n3196), .CLK(clk), .Q(\ram[12][63] ) );
  DFFX1_HVT \ram_reg[12][62]  ( .D(n3195), .CLK(clk), .Q(\ram[12][62] ) );
  DFFX1_HVT \ram_reg[12][61]  ( .D(n3194), .CLK(clk), .Q(\ram[12][61] ) );
  DFFX1_HVT \ram_reg[12][60]  ( .D(n3193), .CLK(clk), .Q(\ram[12][60] ) );
  DFFX1_HVT \ram_reg[12][59]  ( .D(n3192), .CLK(clk), .Q(\ram[12][59] ) );
  DFFX1_HVT \ram_reg[12][58]  ( .D(n3191), .CLK(clk), .Q(\ram[12][58] ) );
  DFFX1_HVT \ram_reg[12][57]  ( .D(n3190), .CLK(clk), .Q(\ram[12][57] ) );
  DFFX1_HVT \ram_reg[12][56]  ( .D(n3189), .CLK(clk), .Q(\ram[12][56] ) );
  DFFX1_HVT \ram_reg[12][55]  ( .D(n3188), .CLK(clk), .Q(\ram[12][55] ) );
  DFFX1_HVT \ram_reg[12][54]  ( .D(n3187), .CLK(clk), .Q(\ram[12][54] ) );
  DFFX1_HVT \ram_reg[12][53]  ( .D(n3186), .CLK(clk), .Q(\ram[12][53] ) );
  DFFX1_HVT \ram_reg[12][52]  ( .D(n3185), .CLK(clk), .Q(\ram[12][52] ) );
  DFFX1_HVT \ram_reg[12][51]  ( .D(n3184), .CLK(clk), .Q(\ram[12][51] ) );
  DFFX1_HVT \ram_reg[12][50]  ( .D(n3183), .CLK(clk), .Q(\ram[12][50] ) );
  DFFX1_HVT \ram_reg[12][49]  ( .D(n3182), .CLK(clk), .Q(\ram[12][49] ) );
  DFFX1_HVT \ram_reg[12][48]  ( .D(n3181), .CLK(clk), .Q(\ram[12][48] ) );
  DFFX1_HVT \ram_reg[12][47]  ( .D(n3180), .CLK(clk), .Q(\ram[12][47] ) );
  DFFX1_HVT \ram_reg[12][46]  ( .D(n3179), .CLK(clk), .Q(\ram[12][46] ) );
  DFFX1_HVT \ram_reg[12][45]  ( .D(n3178), .CLK(clk), .Q(\ram[12][45] ) );
  DFFX1_HVT \ram_reg[12][44]  ( .D(n3177), .CLK(clk), .Q(\ram[12][44] ) );
  DFFX1_HVT \ram_reg[12][43]  ( .D(n3176), .CLK(clk), .Q(\ram[12][43] ) );
  DFFX1_HVT \ram_reg[12][42]  ( .D(n3175), .CLK(clk), .Q(\ram[12][42] ) );
  DFFX1_HVT \ram_reg[12][41]  ( .D(n3174), .CLK(clk), .Q(\ram[12][41] ) );
  DFFX1_HVT \ram_reg[12][40]  ( .D(n3173), .CLK(clk), .Q(\ram[12][40] ) );
  DFFX1_HVT \ram_reg[12][39]  ( .D(n3172), .CLK(clk), .Q(\ram[12][39] ) );
  DFFX1_HVT \ram_reg[12][38]  ( .D(n3171), .CLK(clk), .Q(\ram[12][38] ) );
  DFFX1_HVT \ram_reg[12][37]  ( .D(n3170), .CLK(clk), .Q(\ram[12][37] ) );
  DFFX1_HVT \ram_reg[12][36]  ( .D(n3169), .CLK(clk), .Q(\ram[12][36] ) );
  DFFX1_HVT \ram_reg[12][35]  ( .D(n3168), .CLK(clk), .Q(\ram[12][35] ) );
  DFFX1_HVT \ram_reg[12][34]  ( .D(n3167), .CLK(clk), .Q(\ram[12][34] ) );
  DFFX1_HVT \ram_reg[12][33]  ( .D(n3166), .CLK(clk), .Q(\ram[12][33] ) );
  DFFX1_HVT \ram_reg[12][32]  ( .D(n3165), .CLK(clk), .Q(\ram[12][32] ) );
  DFFX1_HVT \ram_reg[12][31]  ( .D(n3164), .CLK(clk), .Q(\ram[12][31] ) );
  DFFX1_HVT \ram_reg[12][30]  ( .D(n3163), .CLK(clk), .Q(\ram[12][30] ) );
  DFFX1_HVT \ram_reg[12][29]  ( .D(n3162), .CLK(clk), .Q(\ram[12][29] ) );
  DFFX1_HVT \ram_reg[12][28]  ( .D(n3161), .CLK(clk), .Q(\ram[12][28] ) );
  DFFX1_HVT \ram_reg[12][27]  ( .D(n3160), .CLK(clk), .Q(\ram[12][27] ) );
  DFFX1_HVT \ram_reg[12][26]  ( .D(n3159), .CLK(clk), .Q(\ram[12][26] ) );
  DFFX1_HVT \ram_reg[12][25]  ( .D(n3158), .CLK(clk), .Q(\ram[12][25] ) );
  DFFX1_HVT \ram_reg[12][24]  ( .D(n3157), .CLK(clk), .Q(\ram[12][24] ) );
  DFFX1_HVT \ram_reg[12][23]  ( .D(n3156), .CLK(clk), .Q(\ram[12][23] ) );
  DFFX1_HVT \ram_reg[12][22]  ( .D(n3155), .CLK(clk), .Q(\ram[12][22] ) );
  DFFX1_HVT \ram_reg[12][21]  ( .D(n3154), .CLK(clk), .Q(\ram[12][21] ) );
  DFFX1_HVT \ram_reg[12][20]  ( .D(n3153), .CLK(clk), .Q(\ram[12][20] ) );
  DFFX1_HVT \ram_reg[12][19]  ( .D(n3152), .CLK(clk), .Q(\ram[12][19] ) );
  DFFX1_HVT \ram_reg[12][18]  ( .D(n3151), .CLK(clk), .Q(\ram[12][18] ) );
  DFFX1_HVT \ram_reg[12][17]  ( .D(n3150), .CLK(clk), .Q(\ram[12][17] ) );
  DFFX1_HVT \ram_reg[12][16]  ( .D(n3149), .CLK(clk), .Q(\ram[12][16] ) );
  DFFX1_HVT \ram_reg[12][15]  ( .D(n3148), .CLK(clk), .Q(\ram[12][15] ) );
  DFFX1_HVT \ram_reg[12][14]  ( .D(n3147), .CLK(clk), .Q(\ram[12][14] ) );
  DFFX1_HVT \ram_reg[12][13]  ( .D(n3146), .CLK(clk), .Q(\ram[12][13] ) );
  DFFX1_HVT \ram_reg[12][12]  ( .D(n3145), .CLK(clk), .Q(\ram[12][12] ) );
  DFFX1_HVT \ram_reg[12][11]  ( .D(n3144), .CLK(clk), .Q(\ram[12][11] ) );
  DFFX1_HVT \ram_reg[12][10]  ( .D(n3143), .CLK(clk), .Q(\ram[12][10] ) );
  DFFX1_HVT \ram_reg[12][9]  ( .D(n3142), .CLK(clk), .Q(\ram[12][9] ) );
  DFFX1_HVT \ram_reg[12][8]  ( .D(n3141), .CLK(clk), .Q(\ram[12][8] ) );
  DFFX1_HVT \ram_reg[12][7]  ( .D(n3140), .CLK(clk), .Q(\ram[12][7] ) );
  DFFX1_HVT \ram_reg[12][6]  ( .D(n3139), .CLK(clk), .Q(\ram[12][6] ) );
  DFFX1_HVT \ram_reg[12][5]  ( .D(n3138), .CLK(clk), .Q(\ram[12][5] ) );
  DFFX1_HVT \ram_reg[12][4]  ( .D(n3137), .CLK(clk), .Q(\ram[12][4] ) );
  DFFX1_HVT \ram_reg[12][3]  ( .D(n3136), .CLK(clk), .Q(\ram[12][3] ) );
  DFFX1_HVT \ram_reg[12][2]  ( .D(n3135), .CLK(clk), .Q(\ram[12][2] ) );
  DFFX1_HVT \ram_reg[12][1]  ( .D(n3134), .CLK(clk), .Q(\ram[12][1] ) );
  DFFX1_HVT \ram_reg[12][0]  ( .D(n3133), .CLK(clk), .Q(\ram[12][0] ) );
  DFFX1_HVT \ram_reg[11][255]  ( .D(n3132), .CLK(clk), .Q(\ram[11][255] ) );
  DFFX1_HVT \ram_reg[11][254]  ( .D(n3131), .CLK(clk), .Q(\ram[11][254] ) );
  DFFX1_HVT \ram_reg[11][253]  ( .D(n3130), .CLK(clk), .Q(\ram[11][253] ) );
  DFFX1_HVT \ram_reg[11][252]  ( .D(n3129), .CLK(clk), .Q(\ram[11][252] ) );
  DFFX1_HVT \ram_reg[11][251]  ( .D(n3128), .CLK(clk), .Q(\ram[11][251] ) );
  DFFX1_HVT \ram_reg[11][250]  ( .D(n3127), .CLK(clk), .Q(\ram[11][250] ) );
  DFFX1_HVT \ram_reg[11][249]  ( .D(n3126), .CLK(clk), .Q(\ram[11][249] ) );
  DFFX1_HVT \ram_reg[11][248]  ( .D(n3125), .CLK(clk), .Q(\ram[11][248] ) );
  DFFX1_HVT \ram_reg[11][247]  ( .D(n3124), .CLK(clk), .Q(\ram[11][247] ) );
  DFFX1_HVT \ram_reg[11][246]  ( .D(n3123), .CLK(clk), .Q(\ram[11][246] ) );
  DFFX1_HVT \ram_reg[11][245]  ( .D(n3122), .CLK(clk), .Q(\ram[11][245] ) );
  DFFX1_HVT \ram_reg[11][244]  ( .D(n3121), .CLK(clk), .Q(\ram[11][244] ) );
  DFFX1_HVT \ram_reg[11][243]  ( .D(n3120), .CLK(clk), .Q(\ram[11][243] ) );
  DFFX1_HVT \ram_reg[11][242]  ( .D(n3119), .CLK(clk), .Q(\ram[11][242] ) );
  DFFX1_HVT \ram_reg[11][241]  ( .D(n3118), .CLK(clk), .Q(\ram[11][241] ) );
  DFFX1_HVT \ram_reg[11][240]  ( .D(n3117), .CLK(clk), .Q(\ram[11][240] ) );
  DFFX1_HVT \ram_reg[11][239]  ( .D(n3116), .CLK(clk), .Q(\ram[11][239] ) );
  DFFX1_HVT \ram_reg[11][238]  ( .D(n3115), .CLK(clk), .Q(\ram[11][238] ) );
  DFFX1_HVT \ram_reg[11][237]  ( .D(n3114), .CLK(clk), .Q(\ram[11][237] ) );
  DFFX1_HVT \ram_reg[11][236]  ( .D(n3113), .CLK(clk), .Q(\ram[11][236] ) );
  DFFX1_HVT \ram_reg[11][235]  ( .D(n3112), .CLK(clk), .Q(\ram[11][235] ) );
  DFFX1_HVT \ram_reg[11][234]  ( .D(n3111), .CLK(clk), .Q(\ram[11][234] ) );
  DFFX1_HVT \ram_reg[11][233]  ( .D(n3110), .CLK(clk), .Q(\ram[11][233] ) );
  DFFX1_HVT \ram_reg[11][232]  ( .D(n3109), .CLK(clk), .Q(\ram[11][232] ) );
  DFFX1_HVT \ram_reg[11][231]  ( .D(n3108), .CLK(clk), .Q(\ram[11][231] ) );
  DFFX1_HVT \ram_reg[11][230]  ( .D(n3107), .CLK(clk), .Q(\ram[11][230] ) );
  DFFX1_HVT \ram_reg[11][229]  ( .D(n3106), .CLK(clk), .Q(\ram[11][229] ) );
  DFFX1_HVT \ram_reg[11][228]  ( .D(n3105), .CLK(clk), .Q(\ram[11][228] ) );
  DFFX1_HVT \ram_reg[11][227]  ( .D(n3104), .CLK(clk), .Q(\ram[11][227] ) );
  DFFX1_HVT \ram_reg[11][226]  ( .D(n3103), .CLK(clk), .Q(\ram[11][226] ) );
  DFFX1_HVT \ram_reg[11][225]  ( .D(n3102), .CLK(clk), .Q(\ram[11][225] ) );
  DFFX1_HVT \ram_reg[11][224]  ( .D(n3101), .CLK(clk), .Q(\ram[11][224] ) );
  DFFX1_HVT \ram_reg[11][223]  ( .D(n3100), .CLK(clk), .Q(\ram[11][223] ) );
  DFFX1_HVT \ram_reg[11][222]  ( .D(n3099), .CLK(clk), .Q(\ram[11][222] ) );
  DFFX1_HVT \ram_reg[11][221]  ( .D(n3098), .CLK(clk), .Q(\ram[11][221] ) );
  DFFX1_HVT \ram_reg[11][220]  ( .D(n3097), .CLK(clk), .Q(\ram[11][220] ) );
  DFFX1_HVT \ram_reg[11][219]  ( .D(n3096), .CLK(clk), .Q(\ram[11][219] ) );
  DFFX1_HVT \ram_reg[11][218]  ( .D(n3095), .CLK(clk), .Q(\ram[11][218] ) );
  DFFX1_HVT \ram_reg[11][217]  ( .D(n3094), .CLK(clk), .Q(\ram[11][217] ) );
  DFFX1_HVT \ram_reg[11][216]  ( .D(n3093), .CLK(clk), .Q(\ram[11][216] ) );
  DFFX1_HVT \ram_reg[11][215]  ( .D(n3092), .CLK(clk), .Q(\ram[11][215] ) );
  DFFX1_HVT \ram_reg[11][214]  ( .D(n3091), .CLK(clk), .Q(\ram[11][214] ) );
  DFFX1_HVT \ram_reg[11][213]  ( .D(n3090), .CLK(clk), .Q(\ram[11][213] ) );
  DFFX1_HVT \ram_reg[11][212]  ( .D(n3089), .CLK(clk), .Q(\ram[11][212] ) );
  DFFX1_HVT \ram_reg[11][211]  ( .D(n3088), .CLK(clk), .Q(\ram[11][211] ) );
  DFFX1_HVT \ram_reg[11][210]  ( .D(n3087), .CLK(clk), .Q(\ram[11][210] ) );
  DFFX1_HVT \ram_reg[11][209]  ( .D(n3086), .CLK(clk), .Q(\ram[11][209] ) );
  DFFX1_HVT \ram_reg[11][208]  ( .D(n3085), .CLK(clk), .Q(\ram[11][208] ) );
  DFFX1_HVT \ram_reg[11][207]  ( .D(n3084), .CLK(clk), .Q(\ram[11][207] ) );
  DFFX1_HVT \ram_reg[11][206]  ( .D(n3083), .CLK(clk), .Q(\ram[11][206] ) );
  DFFX1_HVT \ram_reg[11][205]  ( .D(n3082), .CLK(clk), .Q(\ram[11][205] ) );
  DFFX1_HVT \ram_reg[11][204]  ( .D(n3081), .CLK(clk), .Q(\ram[11][204] ) );
  DFFX1_HVT \ram_reg[11][203]  ( .D(n3080), .CLK(clk), .Q(\ram[11][203] ) );
  DFFX1_HVT \ram_reg[11][202]  ( .D(n3079), .CLK(clk), .Q(\ram[11][202] ) );
  DFFX1_HVT \ram_reg[11][201]  ( .D(n3078), .CLK(clk), .Q(\ram[11][201] ) );
  DFFX1_HVT \ram_reg[11][200]  ( .D(n3077), .CLK(clk), .Q(\ram[11][200] ) );
  DFFX1_HVT \ram_reg[11][199]  ( .D(n3076), .CLK(clk), .Q(\ram[11][199] ) );
  DFFX1_HVT \ram_reg[11][198]  ( .D(n3075), .CLK(clk), .Q(\ram[11][198] ) );
  DFFX1_HVT \ram_reg[11][197]  ( .D(n3074), .CLK(clk), .Q(\ram[11][197] ) );
  DFFX1_HVT \ram_reg[11][196]  ( .D(n3073), .CLK(clk), .Q(\ram[11][196] ) );
  DFFX1_HVT \ram_reg[11][195]  ( .D(n3072), .CLK(clk), .Q(\ram[11][195] ) );
  DFFX1_HVT \ram_reg[11][194]  ( .D(n3071), .CLK(clk), .Q(\ram[11][194] ) );
  DFFX1_HVT \ram_reg[11][193]  ( .D(n3070), .CLK(clk), .Q(\ram[11][193] ) );
  DFFX1_HVT \ram_reg[11][192]  ( .D(n3069), .CLK(clk), .Q(\ram[11][192] ) );
  DFFX1_HVT \ram_reg[11][191]  ( .D(n3068), .CLK(clk), .Q(\ram[11][191] ) );
  DFFX1_HVT \ram_reg[11][190]  ( .D(n3067), .CLK(clk), .Q(\ram[11][190] ) );
  DFFX1_HVT \ram_reg[11][189]  ( .D(n3066), .CLK(clk), .Q(\ram[11][189] ) );
  DFFX1_HVT \ram_reg[11][188]  ( .D(n3065), .CLK(clk), .Q(\ram[11][188] ) );
  DFFX1_HVT \ram_reg[11][187]  ( .D(n3064), .CLK(clk), .Q(\ram[11][187] ) );
  DFFX1_HVT \ram_reg[11][186]  ( .D(n3063), .CLK(clk), .Q(\ram[11][186] ) );
  DFFX1_HVT \ram_reg[11][185]  ( .D(n3062), .CLK(clk), .Q(\ram[11][185] ) );
  DFFX1_HVT \ram_reg[11][184]  ( .D(n3061), .CLK(clk), .Q(\ram[11][184] ) );
  DFFX1_HVT \ram_reg[11][183]  ( .D(n3060), .CLK(clk), .Q(\ram[11][183] ) );
  DFFX1_HVT \ram_reg[11][182]  ( .D(n3059), .CLK(clk), .Q(\ram[11][182] ) );
  DFFX1_HVT \ram_reg[11][181]  ( .D(n3058), .CLK(clk), .Q(\ram[11][181] ) );
  DFFX1_HVT \ram_reg[11][180]  ( .D(n3057), .CLK(clk), .Q(\ram[11][180] ) );
  DFFX1_HVT \ram_reg[11][179]  ( .D(n3056), .CLK(clk), .Q(\ram[11][179] ) );
  DFFX1_HVT \ram_reg[11][178]  ( .D(n3055), .CLK(clk), .Q(\ram[11][178] ) );
  DFFX1_HVT \ram_reg[11][177]  ( .D(n3054), .CLK(clk), .Q(\ram[11][177] ) );
  DFFX1_HVT \ram_reg[11][176]  ( .D(n3053), .CLK(clk), .Q(\ram[11][176] ) );
  DFFX1_HVT \ram_reg[11][175]  ( .D(n3052), .CLK(clk), .Q(\ram[11][175] ) );
  DFFX1_HVT \ram_reg[11][174]  ( .D(n3051), .CLK(clk), .Q(\ram[11][174] ) );
  DFFX1_HVT \ram_reg[11][173]  ( .D(n3050), .CLK(clk), .Q(\ram[11][173] ) );
  DFFX1_HVT \ram_reg[11][172]  ( .D(n3049), .CLK(clk), .Q(\ram[11][172] ) );
  DFFX1_HVT \ram_reg[11][171]  ( .D(n3048), .CLK(clk), .Q(\ram[11][171] ) );
  DFFX1_HVT \ram_reg[11][170]  ( .D(n3047), .CLK(clk), .Q(\ram[11][170] ) );
  DFFX1_HVT \ram_reg[11][169]  ( .D(n3046), .CLK(clk), .Q(\ram[11][169] ) );
  DFFX1_HVT \ram_reg[11][168]  ( .D(n3045), .CLK(clk), .Q(\ram[11][168] ) );
  DFFX1_HVT \ram_reg[11][167]  ( .D(n3044), .CLK(clk), .Q(\ram[11][167] ) );
  DFFX1_HVT \ram_reg[11][166]  ( .D(n3043), .CLK(clk), .Q(\ram[11][166] ) );
  DFFX1_HVT \ram_reg[11][165]  ( .D(n3042), .CLK(clk), .Q(\ram[11][165] ) );
  DFFX1_HVT \ram_reg[11][164]  ( .D(n3041), .CLK(clk), .Q(\ram[11][164] ) );
  DFFX1_HVT \ram_reg[11][163]  ( .D(n3040), .CLK(clk), .Q(\ram[11][163] ) );
  DFFX1_HVT \ram_reg[11][162]  ( .D(n3039), .CLK(clk), .Q(\ram[11][162] ) );
  DFFX1_HVT \ram_reg[11][161]  ( .D(n3038), .CLK(clk), .Q(\ram[11][161] ) );
  DFFX1_HVT \ram_reg[11][160]  ( .D(n3037), .CLK(clk), .Q(\ram[11][160] ) );
  DFFX1_HVT \ram_reg[11][159]  ( .D(n3036), .CLK(clk), .Q(\ram[11][159] ) );
  DFFX1_HVT \ram_reg[11][158]  ( .D(n3035), .CLK(clk), .Q(\ram[11][158] ) );
  DFFX1_HVT \ram_reg[11][157]  ( .D(n3034), .CLK(clk), .Q(\ram[11][157] ) );
  DFFX1_HVT \ram_reg[11][156]  ( .D(n3033), .CLK(clk), .Q(\ram[11][156] ) );
  DFFX1_HVT \ram_reg[11][155]  ( .D(n3032), .CLK(clk), .Q(\ram[11][155] ) );
  DFFX1_HVT \ram_reg[11][154]  ( .D(n3031), .CLK(clk), .Q(\ram[11][154] ) );
  DFFX1_HVT \ram_reg[11][153]  ( .D(n3030), .CLK(clk), .Q(\ram[11][153] ) );
  DFFX1_HVT \ram_reg[11][152]  ( .D(n3029), .CLK(clk), .Q(\ram[11][152] ) );
  DFFX1_HVT \ram_reg[11][151]  ( .D(n3028), .CLK(clk), .Q(\ram[11][151] ) );
  DFFX1_HVT \ram_reg[11][150]  ( .D(n3027), .CLK(clk), .Q(\ram[11][150] ) );
  DFFX1_HVT \ram_reg[11][149]  ( .D(n3026), .CLK(clk), .Q(\ram[11][149] ) );
  DFFX1_HVT \ram_reg[11][148]  ( .D(n3025), .CLK(clk), .Q(\ram[11][148] ) );
  DFFX1_HVT \ram_reg[11][147]  ( .D(n3024), .CLK(clk), .Q(\ram[11][147] ) );
  DFFX1_HVT \ram_reg[11][146]  ( .D(n3023), .CLK(clk), .Q(\ram[11][146] ) );
  DFFX1_HVT \ram_reg[11][145]  ( .D(n3022), .CLK(clk), .Q(\ram[11][145] ) );
  DFFX1_HVT \ram_reg[11][144]  ( .D(n3021), .CLK(clk), .Q(\ram[11][144] ) );
  DFFX1_HVT \ram_reg[11][143]  ( .D(n3020), .CLK(clk), .Q(\ram[11][143] ) );
  DFFX1_HVT \ram_reg[11][142]  ( .D(n3019), .CLK(clk), .Q(\ram[11][142] ) );
  DFFX1_HVT \ram_reg[11][141]  ( .D(n3018), .CLK(clk), .Q(\ram[11][141] ) );
  DFFX1_HVT \ram_reg[11][140]  ( .D(n3017), .CLK(clk), .Q(\ram[11][140] ) );
  DFFX1_HVT \ram_reg[11][139]  ( .D(n3016), .CLK(clk), .Q(\ram[11][139] ) );
  DFFX1_HVT \ram_reg[11][138]  ( .D(n3015), .CLK(clk), .Q(\ram[11][138] ) );
  DFFX1_HVT \ram_reg[11][137]  ( .D(n3014), .CLK(clk), .Q(\ram[11][137] ) );
  DFFX1_HVT \ram_reg[11][136]  ( .D(n3013), .CLK(clk), .Q(\ram[11][136] ) );
  DFFX1_HVT \ram_reg[11][135]  ( .D(n3012), .CLK(clk), .Q(\ram[11][135] ) );
  DFFX1_HVT \ram_reg[11][134]  ( .D(n3011), .CLK(clk), .Q(\ram[11][134] ) );
  DFFX1_HVT \ram_reg[11][133]  ( .D(n3010), .CLK(clk), .Q(\ram[11][133] ) );
  DFFX1_HVT \ram_reg[11][132]  ( .D(n3009), .CLK(clk), .Q(\ram[11][132] ) );
  DFFX1_HVT \ram_reg[11][131]  ( .D(n3008), .CLK(clk), .Q(\ram[11][131] ) );
  DFFX1_HVT \ram_reg[11][130]  ( .D(n3007), .CLK(clk), .Q(\ram[11][130] ) );
  DFFX1_HVT \ram_reg[11][129]  ( .D(n3006), .CLK(clk), .Q(\ram[11][129] ) );
  DFFX1_HVT \ram_reg[11][128]  ( .D(n3005), .CLK(clk), .Q(\ram[11][128] ) );
  DFFX1_HVT \ram_reg[11][127]  ( .D(n3004), .CLK(clk), .Q(\ram[11][127] ) );
  DFFX1_HVT \ram_reg[11][126]  ( .D(n3003), .CLK(clk), .Q(\ram[11][126] ) );
  DFFX1_HVT \ram_reg[11][125]  ( .D(n3002), .CLK(clk), .Q(\ram[11][125] ) );
  DFFX1_HVT \ram_reg[11][124]  ( .D(n3001), .CLK(clk), .Q(\ram[11][124] ) );
  DFFX1_HVT \ram_reg[11][123]  ( .D(n3000), .CLK(clk), .Q(\ram[11][123] ) );
  DFFX1_HVT \ram_reg[11][122]  ( .D(n2999), .CLK(clk), .Q(\ram[11][122] ) );
  DFFX1_HVT \ram_reg[11][121]  ( .D(n2998), .CLK(clk), .Q(\ram[11][121] ) );
  DFFX1_HVT \ram_reg[11][120]  ( .D(n2997), .CLK(clk), .Q(\ram[11][120] ) );
  DFFX1_HVT \ram_reg[11][119]  ( .D(n2996), .CLK(clk), .Q(\ram[11][119] ) );
  DFFX1_HVT \ram_reg[11][118]  ( .D(n2995), .CLK(clk), .Q(\ram[11][118] ) );
  DFFX1_HVT \ram_reg[11][117]  ( .D(n2994), .CLK(clk), .Q(\ram[11][117] ) );
  DFFX1_HVT \ram_reg[11][116]  ( .D(n2993), .CLK(clk), .Q(\ram[11][116] ) );
  DFFX1_HVT \ram_reg[11][115]  ( .D(n2992), .CLK(clk), .Q(\ram[11][115] ) );
  DFFX1_HVT \ram_reg[11][114]  ( .D(n2991), .CLK(clk), .Q(\ram[11][114] ) );
  DFFX1_HVT \ram_reg[11][113]  ( .D(n2990), .CLK(clk), .Q(\ram[11][113] ) );
  DFFX1_HVT \ram_reg[11][112]  ( .D(n2989), .CLK(clk), .Q(\ram[11][112] ) );
  DFFX1_HVT \ram_reg[11][111]  ( .D(n2988), .CLK(clk), .Q(\ram[11][111] ) );
  DFFX1_HVT \ram_reg[11][110]  ( .D(n2987), .CLK(clk), .Q(\ram[11][110] ) );
  DFFX1_HVT \ram_reg[11][109]  ( .D(n2986), .CLK(clk), .Q(\ram[11][109] ) );
  DFFX1_HVT \ram_reg[11][108]  ( .D(n2985), .CLK(clk), .Q(\ram[11][108] ) );
  DFFX1_HVT \ram_reg[11][107]  ( .D(n2984), .CLK(clk), .Q(\ram[11][107] ) );
  DFFX1_HVT \ram_reg[11][106]  ( .D(n2983), .CLK(clk), .Q(\ram[11][106] ) );
  DFFX1_HVT \ram_reg[11][105]  ( .D(n2982), .CLK(clk), .Q(\ram[11][105] ) );
  DFFX1_HVT \ram_reg[11][104]  ( .D(n2981), .CLK(clk), .Q(\ram[11][104] ) );
  DFFX1_HVT \ram_reg[11][103]  ( .D(n2980), .CLK(clk), .Q(\ram[11][103] ) );
  DFFX1_HVT \ram_reg[11][102]  ( .D(n2979), .CLK(clk), .Q(\ram[11][102] ) );
  DFFX1_HVT \ram_reg[11][101]  ( .D(n2978), .CLK(clk), .Q(\ram[11][101] ) );
  DFFX1_HVT \ram_reg[11][100]  ( .D(n2977), .CLK(clk), .Q(\ram[11][100] ) );
  DFFX1_HVT \ram_reg[11][99]  ( .D(n2976), .CLK(clk), .Q(\ram[11][99] ) );
  DFFX1_HVT \ram_reg[11][98]  ( .D(n2975), .CLK(clk), .Q(\ram[11][98] ) );
  DFFX1_HVT \ram_reg[11][97]  ( .D(n2974), .CLK(clk), .Q(\ram[11][97] ) );
  DFFX1_HVT \ram_reg[11][96]  ( .D(n2973), .CLK(clk), .Q(\ram[11][96] ) );
  DFFX1_HVT \ram_reg[11][95]  ( .D(n2972), .CLK(clk), .Q(\ram[11][95] ) );
  DFFX1_HVT \ram_reg[11][94]  ( .D(n2971), .CLK(clk), .Q(\ram[11][94] ) );
  DFFX1_HVT \ram_reg[11][93]  ( .D(n2970), .CLK(clk), .Q(\ram[11][93] ) );
  DFFX1_HVT \ram_reg[11][92]  ( .D(n2969), .CLK(clk), .Q(\ram[11][92] ) );
  DFFX1_HVT \ram_reg[11][91]  ( .D(n2968), .CLK(clk), .Q(\ram[11][91] ) );
  DFFX1_HVT \ram_reg[11][90]  ( .D(n2967), .CLK(clk), .Q(\ram[11][90] ) );
  DFFX1_HVT \ram_reg[11][89]  ( .D(n2966), .CLK(clk), .Q(\ram[11][89] ) );
  DFFX1_HVT \ram_reg[11][88]  ( .D(n2965), .CLK(clk), .Q(\ram[11][88] ) );
  DFFX1_HVT \ram_reg[11][87]  ( .D(n2964), .CLK(clk), .Q(\ram[11][87] ) );
  DFFX1_HVT \ram_reg[11][86]  ( .D(n2963), .CLK(clk), .Q(\ram[11][86] ) );
  DFFX1_HVT \ram_reg[11][85]  ( .D(n2962), .CLK(clk), .Q(\ram[11][85] ) );
  DFFX1_HVT \ram_reg[11][84]  ( .D(n2961), .CLK(clk), .Q(\ram[11][84] ) );
  DFFX1_HVT \ram_reg[11][83]  ( .D(n2960), .CLK(clk), .Q(\ram[11][83] ) );
  DFFX1_HVT \ram_reg[11][82]  ( .D(n2959), .CLK(clk), .Q(\ram[11][82] ) );
  DFFX1_HVT \ram_reg[11][81]  ( .D(n2958), .CLK(clk), .Q(\ram[11][81] ) );
  DFFX1_HVT \ram_reg[11][80]  ( .D(n2957), .CLK(clk), .Q(\ram[11][80] ) );
  DFFX1_HVT \ram_reg[11][79]  ( .D(n2956), .CLK(clk), .Q(\ram[11][79] ) );
  DFFX1_HVT \ram_reg[11][78]  ( .D(n2955), .CLK(clk), .Q(\ram[11][78] ) );
  DFFX1_HVT \ram_reg[11][77]  ( .D(n2954), .CLK(clk), .Q(\ram[11][77] ) );
  DFFX1_HVT \ram_reg[11][76]  ( .D(n2953), .CLK(clk), .Q(\ram[11][76] ) );
  DFFX1_HVT \ram_reg[11][75]  ( .D(n2952), .CLK(clk), .Q(\ram[11][75] ) );
  DFFX1_HVT \ram_reg[11][74]  ( .D(n2951), .CLK(clk), .Q(\ram[11][74] ) );
  DFFX1_HVT \ram_reg[11][73]  ( .D(n2950), .CLK(clk), .Q(\ram[11][73] ) );
  DFFX1_HVT \ram_reg[11][72]  ( .D(n2949), .CLK(clk), .Q(\ram[11][72] ) );
  DFFX1_HVT \ram_reg[11][71]  ( .D(n2948), .CLK(clk), .Q(\ram[11][71] ) );
  DFFX1_HVT \ram_reg[11][70]  ( .D(n2947), .CLK(clk), .Q(\ram[11][70] ) );
  DFFX1_HVT \ram_reg[11][69]  ( .D(n2946), .CLK(clk), .Q(\ram[11][69] ) );
  DFFX1_HVT \ram_reg[11][68]  ( .D(n2945), .CLK(clk), .Q(\ram[11][68] ) );
  DFFX1_HVT \ram_reg[11][67]  ( .D(n2944), .CLK(clk), .Q(\ram[11][67] ) );
  DFFX1_HVT \ram_reg[11][66]  ( .D(n2943), .CLK(clk), .Q(\ram[11][66] ) );
  DFFX1_HVT \ram_reg[11][65]  ( .D(n2942), .CLK(clk), .Q(\ram[11][65] ) );
  DFFX1_HVT \ram_reg[11][64]  ( .D(n2941), .CLK(clk), .Q(\ram[11][64] ) );
  DFFX1_HVT \ram_reg[11][63]  ( .D(n2940), .CLK(clk), .Q(\ram[11][63] ) );
  DFFX1_HVT \ram_reg[11][62]  ( .D(n2939), .CLK(clk), .Q(\ram[11][62] ) );
  DFFX1_HVT \ram_reg[11][61]  ( .D(n2938), .CLK(clk), .Q(\ram[11][61] ) );
  DFFX1_HVT \ram_reg[11][60]  ( .D(n2937), .CLK(clk), .Q(\ram[11][60] ) );
  DFFX1_HVT \ram_reg[11][59]  ( .D(n2936), .CLK(clk), .Q(\ram[11][59] ) );
  DFFX1_HVT \ram_reg[11][58]  ( .D(n2935), .CLK(clk), .Q(\ram[11][58] ) );
  DFFX1_HVT \ram_reg[11][57]  ( .D(n2934), .CLK(clk), .Q(\ram[11][57] ) );
  DFFX1_HVT \ram_reg[11][56]  ( .D(n2933), .CLK(clk), .Q(\ram[11][56] ) );
  DFFX1_HVT \ram_reg[11][55]  ( .D(n2932), .CLK(clk), .Q(\ram[11][55] ) );
  DFFX1_HVT \ram_reg[11][54]  ( .D(n2931), .CLK(clk), .Q(\ram[11][54] ) );
  DFFX1_HVT \ram_reg[11][53]  ( .D(n2930), .CLK(clk), .Q(\ram[11][53] ) );
  DFFX1_HVT \ram_reg[11][52]  ( .D(n2929), .CLK(clk), .Q(\ram[11][52] ) );
  DFFX1_HVT \ram_reg[11][51]  ( .D(n2928), .CLK(clk), .Q(\ram[11][51] ) );
  DFFX1_HVT \ram_reg[11][50]  ( .D(n2927), .CLK(clk), .Q(\ram[11][50] ) );
  DFFX1_HVT \ram_reg[11][49]  ( .D(n2926), .CLK(clk), .Q(\ram[11][49] ) );
  DFFX1_HVT \ram_reg[11][48]  ( .D(n2925), .CLK(clk), .Q(\ram[11][48] ) );
  DFFX1_HVT \ram_reg[11][47]  ( .D(n2924), .CLK(clk), .Q(\ram[11][47] ) );
  DFFX1_HVT \ram_reg[11][46]  ( .D(n2923), .CLK(clk), .Q(\ram[11][46] ) );
  DFFX1_HVT \ram_reg[11][45]  ( .D(n2922), .CLK(clk), .Q(\ram[11][45] ) );
  DFFX1_HVT \ram_reg[11][44]  ( .D(n2921), .CLK(clk), .Q(\ram[11][44] ) );
  DFFX1_HVT \ram_reg[11][43]  ( .D(n2920), .CLK(clk), .Q(\ram[11][43] ) );
  DFFX1_HVT \ram_reg[11][42]  ( .D(n2919), .CLK(clk), .Q(\ram[11][42] ) );
  DFFX1_HVT \ram_reg[11][41]  ( .D(n2918), .CLK(clk), .Q(\ram[11][41] ) );
  DFFX1_HVT \ram_reg[11][40]  ( .D(n2917), .CLK(clk), .Q(\ram[11][40] ) );
  DFFX1_HVT \ram_reg[11][39]  ( .D(n2916), .CLK(clk), .Q(\ram[11][39] ) );
  DFFX1_HVT \ram_reg[11][38]  ( .D(n2915), .CLK(clk), .Q(\ram[11][38] ) );
  DFFX1_HVT \ram_reg[11][37]  ( .D(n2914), .CLK(clk), .Q(\ram[11][37] ) );
  DFFX1_HVT \ram_reg[11][36]  ( .D(n2913), .CLK(clk), .Q(\ram[11][36] ) );
  DFFX1_HVT \ram_reg[11][35]  ( .D(n2912), .CLK(clk), .Q(\ram[11][35] ) );
  DFFX1_HVT \ram_reg[11][34]  ( .D(n2911), .CLK(clk), .Q(\ram[11][34] ) );
  DFFX1_HVT \ram_reg[11][33]  ( .D(n2910), .CLK(clk), .Q(\ram[11][33] ) );
  DFFX1_HVT \ram_reg[11][32]  ( .D(n2909), .CLK(clk), .Q(\ram[11][32] ) );
  DFFX1_HVT \ram_reg[11][31]  ( .D(n2908), .CLK(clk), .Q(\ram[11][31] ) );
  DFFX1_HVT \ram_reg[11][30]  ( .D(n2907), .CLK(clk), .Q(\ram[11][30] ) );
  DFFX1_HVT \ram_reg[11][29]  ( .D(n2906), .CLK(clk), .Q(\ram[11][29] ) );
  DFFX1_HVT \ram_reg[11][28]  ( .D(n2905), .CLK(clk), .Q(\ram[11][28] ) );
  DFFX1_HVT \ram_reg[11][27]  ( .D(n2904), .CLK(clk), .Q(\ram[11][27] ) );
  DFFX1_HVT \ram_reg[11][26]  ( .D(n2903), .CLK(clk), .Q(\ram[11][26] ) );
  DFFX1_HVT \ram_reg[11][25]  ( .D(n2902), .CLK(clk), .Q(\ram[11][25] ) );
  DFFX1_HVT \ram_reg[11][24]  ( .D(n2901), .CLK(clk), .Q(\ram[11][24] ) );
  DFFX1_HVT \ram_reg[11][23]  ( .D(n2900), .CLK(clk), .Q(\ram[11][23] ) );
  DFFX1_HVT \ram_reg[11][22]  ( .D(n2899), .CLK(clk), .Q(\ram[11][22] ) );
  DFFX1_HVT \ram_reg[11][21]  ( .D(n2898), .CLK(clk), .Q(\ram[11][21] ) );
  DFFX1_HVT \ram_reg[11][20]  ( .D(n2897), .CLK(clk), .Q(\ram[11][20] ) );
  DFFX1_HVT \ram_reg[11][19]  ( .D(n2896), .CLK(clk), .Q(\ram[11][19] ) );
  DFFX1_HVT \ram_reg[11][18]  ( .D(n2895), .CLK(clk), .Q(\ram[11][18] ) );
  DFFX1_HVT \ram_reg[11][17]  ( .D(n2894), .CLK(clk), .Q(\ram[11][17] ) );
  DFFX1_HVT \ram_reg[11][16]  ( .D(n2893), .CLK(clk), .Q(\ram[11][16] ) );
  DFFX1_HVT \ram_reg[11][15]  ( .D(n2892), .CLK(clk), .Q(\ram[11][15] ) );
  DFFX1_HVT \ram_reg[11][14]  ( .D(n2891), .CLK(clk), .Q(\ram[11][14] ) );
  DFFX1_HVT \ram_reg[11][13]  ( .D(n2890), .CLK(clk), .Q(\ram[11][13] ) );
  DFFX1_HVT \ram_reg[11][12]  ( .D(n2889), .CLK(clk), .Q(\ram[11][12] ) );
  DFFX1_HVT \ram_reg[11][11]  ( .D(n2888), .CLK(clk), .Q(\ram[11][11] ) );
  DFFX1_HVT \ram_reg[11][10]  ( .D(n2887), .CLK(clk), .Q(\ram[11][10] ) );
  DFFX1_HVT \ram_reg[11][9]  ( .D(n2886), .CLK(clk), .Q(\ram[11][9] ) );
  DFFX1_HVT \ram_reg[11][8]  ( .D(n2885), .CLK(clk), .Q(\ram[11][8] ) );
  DFFX1_HVT \ram_reg[11][7]  ( .D(n2884), .CLK(clk), .Q(\ram[11][7] ) );
  DFFX1_HVT \ram_reg[11][6]  ( .D(n2883), .CLK(clk), .Q(\ram[11][6] ) );
  DFFX1_HVT \ram_reg[11][5]  ( .D(n2882), .CLK(clk), .Q(\ram[11][5] ) );
  DFFX1_HVT \ram_reg[11][4]  ( .D(n2881), .CLK(clk), .Q(\ram[11][4] ) );
  DFFX1_HVT \ram_reg[11][3]  ( .D(n2880), .CLK(clk), .Q(\ram[11][3] ) );
  DFFX1_HVT \ram_reg[11][2]  ( .D(n2879), .CLK(clk), .Q(\ram[11][2] ) );
  DFFX1_HVT \ram_reg[11][1]  ( .D(n2878), .CLK(clk), .Q(\ram[11][1] ) );
  DFFX1_HVT \ram_reg[11][0]  ( .D(n2877), .CLK(clk), .Q(\ram[11][0] ) );
  DFFX1_HVT \ram_reg[10][255]  ( .D(n2876), .CLK(clk), .Q(\ram[10][255] ) );
  DFFX1_HVT \ram_reg[10][254]  ( .D(n2875), .CLK(clk), .Q(\ram[10][254] ) );
  DFFX1_HVT \ram_reg[10][253]  ( .D(n2874), .CLK(clk), .Q(\ram[10][253] ) );
  DFFX1_HVT \ram_reg[10][252]  ( .D(n2873), .CLK(clk), .Q(\ram[10][252] ) );
  DFFX1_HVT \ram_reg[10][251]  ( .D(n2872), .CLK(clk), .Q(\ram[10][251] ) );
  DFFX1_HVT \ram_reg[10][250]  ( .D(n2871), .CLK(clk), .Q(\ram[10][250] ) );
  DFFX1_HVT \ram_reg[10][249]  ( .D(n2870), .CLK(clk), .Q(\ram[10][249] ) );
  DFFX1_HVT \ram_reg[10][248]  ( .D(n2869), .CLK(clk), .Q(\ram[10][248] ) );
  DFFX1_HVT \ram_reg[10][247]  ( .D(n2868), .CLK(clk), .Q(\ram[10][247] ) );
  DFFX1_HVT \ram_reg[10][246]  ( .D(n2867), .CLK(clk), .Q(\ram[10][246] ) );
  DFFX1_HVT \ram_reg[10][245]  ( .D(n2866), .CLK(clk), .Q(\ram[10][245] ) );
  DFFX1_HVT \ram_reg[10][244]  ( .D(n2865), .CLK(clk), .Q(\ram[10][244] ) );
  DFFX1_HVT \ram_reg[10][243]  ( .D(n2864), .CLK(clk), .Q(\ram[10][243] ) );
  DFFX1_HVT \ram_reg[10][242]  ( .D(n2863), .CLK(clk), .Q(\ram[10][242] ) );
  DFFX1_HVT \ram_reg[10][241]  ( .D(n2862), .CLK(clk), .Q(\ram[10][241] ) );
  DFFX1_HVT \ram_reg[10][240]  ( .D(n2861), .CLK(clk), .Q(\ram[10][240] ) );
  DFFX1_HVT \ram_reg[10][239]  ( .D(n2860), .CLK(clk), .Q(\ram[10][239] ) );
  DFFX1_HVT \ram_reg[10][238]  ( .D(n2859), .CLK(clk), .Q(\ram[10][238] ) );
  DFFX1_HVT \ram_reg[10][237]  ( .D(n2858), .CLK(clk), .Q(\ram[10][237] ) );
  DFFX1_HVT \ram_reg[10][236]  ( .D(n2857), .CLK(clk), .Q(\ram[10][236] ) );
  DFFX1_HVT \ram_reg[10][235]  ( .D(n2856), .CLK(clk), .Q(\ram[10][235] ) );
  DFFX1_HVT \ram_reg[10][234]  ( .D(n2855), .CLK(clk), .Q(\ram[10][234] ) );
  DFFX1_HVT \ram_reg[10][233]  ( .D(n2854), .CLK(clk), .Q(\ram[10][233] ) );
  DFFX1_HVT \ram_reg[10][232]  ( .D(n2853), .CLK(clk), .Q(\ram[10][232] ) );
  DFFX1_HVT \ram_reg[10][231]  ( .D(n2852), .CLK(clk), .Q(\ram[10][231] ) );
  DFFX1_HVT \ram_reg[10][230]  ( .D(n2851), .CLK(clk), .Q(\ram[10][230] ) );
  DFFX1_HVT \ram_reg[10][229]  ( .D(n2850), .CLK(clk), .Q(\ram[10][229] ) );
  DFFX1_HVT \ram_reg[10][228]  ( .D(n2849), .CLK(clk), .Q(\ram[10][228] ) );
  DFFX1_HVT \ram_reg[10][227]  ( .D(n2848), .CLK(clk), .Q(\ram[10][227] ) );
  DFFX1_HVT \ram_reg[10][226]  ( .D(n2847), .CLK(clk), .Q(\ram[10][226] ) );
  DFFX1_HVT \ram_reg[10][225]  ( .D(n2846), .CLK(clk), .Q(\ram[10][225] ) );
  DFFX1_HVT \ram_reg[10][224]  ( .D(n2845), .CLK(clk), .Q(\ram[10][224] ) );
  DFFX1_HVT \ram_reg[10][223]  ( .D(n2844), .CLK(clk), .Q(\ram[10][223] ) );
  DFFX1_HVT \ram_reg[10][222]  ( .D(n2843), .CLK(clk), .Q(\ram[10][222] ) );
  DFFX1_HVT \ram_reg[10][221]  ( .D(n2842), .CLK(clk), .Q(\ram[10][221] ) );
  DFFX1_HVT \ram_reg[10][220]  ( .D(n2841), .CLK(clk), .Q(\ram[10][220] ) );
  DFFX1_HVT \ram_reg[10][219]  ( .D(n2840), .CLK(clk), .Q(\ram[10][219] ) );
  DFFX1_HVT \ram_reg[10][218]  ( .D(n2839), .CLK(clk), .Q(\ram[10][218] ) );
  DFFX1_HVT \ram_reg[10][217]  ( .D(n2838), .CLK(clk), .Q(\ram[10][217] ) );
  DFFX1_HVT \ram_reg[10][216]  ( .D(n2837), .CLK(clk), .Q(\ram[10][216] ) );
  DFFX1_HVT \ram_reg[10][215]  ( .D(n2836), .CLK(clk), .Q(\ram[10][215] ) );
  DFFX1_HVT \ram_reg[10][214]  ( .D(n2835), .CLK(clk), .Q(\ram[10][214] ) );
  DFFX1_HVT \ram_reg[10][213]  ( .D(n2834), .CLK(clk), .Q(\ram[10][213] ) );
  DFFX1_HVT \ram_reg[10][212]  ( .D(n2833), .CLK(clk), .Q(\ram[10][212] ) );
  DFFX1_HVT \ram_reg[10][211]  ( .D(n2832), .CLK(clk), .Q(\ram[10][211] ) );
  DFFX1_HVT \ram_reg[10][210]  ( .D(n2831), .CLK(clk), .Q(\ram[10][210] ) );
  DFFX1_HVT \ram_reg[10][209]  ( .D(n2830), .CLK(clk), .Q(\ram[10][209] ) );
  DFFX1_HVT \ram_reg[10][208]  ( .D(n2829), .CLK(clk), .Q(\ram[10][208] ) );
  DFFX1_HVT \ram_reg[10][207]  ( .D(n2828), .CLK(clk), .Q(\ram[10][207] ) );
  DFFX1_HVT \ram_reg[10][206]  ( .D(n2827), .CLK(clk), .Q(\ram[10][206] ) );
  DFFX1_HVT \ram_reg[10][205]  ( .D(n2826), .CLK(clk), .Q(\ram[10][205] ) );
  DFFX1_HVT \ram_reg[10][204]  ( .D(n2825), .CLK(clk), .Q(\ram[10][204] ) );
  DFFX1_HVT \ram_reg[10][203]  ( .D(n2824), .CLK(clk), .Q(\ram[10][203] ) );
  DFFX1_HVT \ram_reg[10][202]  ( .D(n2823), .CLK(clk), .Q(\ram[10][202] ) );
  DFFX1_HVT \ram_reg[10][201]  ( .D(n2822), .CLK(clk), .Q(\ram[10][201] ) );
  DFFX1_HVT \ram_reg[10][200]  ( .D(n2821), .CLK(clk), .Q(\ram[10][200] ) );
  DFFX1_HVT \ram_reg[10][199]  ( .D(n2820), .CLK(clk), .Q(\ram[10][199] ) );
  DFFX1_HVT \ram_reg[10][198]  ( .D(n2819), .CLK(clk), .Q(\ram[10][198] ) );
  DFFX1_HVT \ram_reg[10][197]  ( .D(n2818), .CLK(clk), .Q(\ram[10][197] ) );
  DFFX1_HVT \ram_reg[10][196]  ( .D(n2817), .CLK(clk), .Q(\ram[10][196] ) );
  DFFX1_HVT \ram_reg[10][195]  ( .D(n2816), .CLK(clk), .Q(\ram[10][195] ) );
  DFFX1_HVT \ram_reg[10][194]  ( .D(n2815), .CLK(clk), .Q(\ram[10][194] ) );
  DFFX1_HVT \ram_reg[10][193]  ( .D(n2814), .CLK(clk), .Q(\ram[10][193] ) );
  DFFX1_HVT \ram_reg[10][192]  ( .D(n2813), .CLK(clk), .Q(\ram[10][192] ) );
  DFFX1_HVT \ram_reg[10][191]  ( .D(n2812), .CLK(clk), .Q(\ram[10][191] ) );
  DFFX1_HVT \ram_reg[10][190]  ( .D(n2811), .CLK(clk), .Q(\ram[10][190] ) );
  DFFX1_HVT \ram_reg[10][189]  ( .D(n2810), .CLK(clk), .Q(\ram[10][189] ) );
  DFFX1_HVT \ram_reg[10][188]  ( .D(n2809), .CLK(clk), .Q(\ram[10][188] ) );
  DFFX1_HVT \ram_reg[10][187]  ( .D(n2808), .CLK(clk), .Q(\ram[10][187] ) );
  DFFX1_HVT \ram_reg[10][186]  ( .D(n2807), .CLK(clk), .Q(\ram[10][186] ) );
  DFFX1_HVT \ram_reg[10][185]  ( .D(n2806), .CLK(clk), .Q(\ram[10][185] ) );
  DFFX1_HVT \ram_reg[10][184]  ( .D(n2805), .CLK(clk), .Q(\ram[10][184] ) );
  DFFX1_HVT \ram_reg[10][183]  ( .D(n2804), .CLK(clk), .Q(\ram[10][183] ) );
  DFFX1_HVT \ram_reg[10][182]  ( .D(n2803), .CLK(clk), .Q(\ram[10][182] ) );
  DFFX1_HVT \ram_reg[10][181]  ( .D(n2802), .CLK(clk), .Q(\ram[10][181] ) );
  DFFX1_HVT \ram_reg[10][180]  ( .D(n2801), .CLK(clk), .Q(\ram[10][180] ) );
  DFFX1_HVT \ram_reg[10][179]  ( .D(n2800), .CLK(clk), .Q(\ram[10][179] ) );
  DFFX1_HVT \ram_reg[10][178]  ( .D(n2799), .CLK(clk), .Q(\ram[10][178] ) );
  DFFX1_HVT \ram_reg[10][177]  ( .D(n2798), .CLK(clk), .Q(\ram[10][177] ) );
  DFFX1_HVT \ram_reg[10][176]  ( .D(n2797), .CLK(clk), .Q(\ram[10][176] ) );
  DFFX1_HVT \ram_reg[10][175]  ( .D(n2796), .CLK(clk), .Q(\ram[10][175] ) );
  DFFX1_HVT \ram_reg[10][174]  ( .D(n2795), .CLK(clk), .Q(\ram[10][174] ) );
  DFFX1_HVT \ram_reg[10][173]  ( .D(n2794), .CLK(clk), .Q(\ram[10][173] ) );
  DFFX1_HVT \ram_reg[10][172]  ( .D(n2793), .CLK(clk), .Q(\ram[10][172] ) );
  DFFX1_HVT \ram_reg[10][171]  ( .D(n2792), .CLK(clk), .Q(\ram[10][171] ) );
  DFFX1_HVT \ram_reg[10][170]  ( .D(n2791), .CLK(clk), .Q(\ram[10][170] ) );
  DFFX1_HVT \ram_reg[10][169]  ( .D(n2790), .CLK(clk), .Q(\ram[10][169] ) );
  DFFX1_HVT \ram_reg[10][168]  ( .D(n2789), .CLK(clk), .Q(\ram[10][168] ) );
  DFFX1_HVT \ram_reg[10][167]  ( .D(n2788), .CLK(clk), .Q(\ram[10][167] ) );
  DFFX1_HVT \ram_reg[10][166]  ( .D(n2787), .CLK(clk), .Q(\ram[10][166] ) );
  DFFX1_HVT \ram_reg[10][165]  ( .D(n2786), .CLK(clk), .Q(\ram[10][165] ) );
  DFFX1_HVT \ram_reg[10][164]  ( .D(n2785), .CLK(clk), .Q(\ram[10][164] ) );
  DFFX1_HVT \ram_reg[10][163]  ( .D(n2784), .CLK(clk), .Q(\ram[10][163] ) );
  DFFX1_HVT \ram_reg[10][162]  ( .D(n2783), .CLK(clk), .Q(\ram[10][162] ) );
  DFFX1_HVT \ram_reg[10][161]  ( .D(n2782), .CLK(clk), .Q(\ram[10][161] ) );
  DFFX1_HVT \ram_reg[10][160]  ( .D(n2781), .CLK(clk), .Q(\ram[10][160] ) );
  DFFX1_HVT \ram_reg[10][159]  ( .D(n2780), .CLK(clk), .Q(\ram[10][159] ) );
  DFFX1_HVT \ram_reg[10][158]  ( .D(n2779), .CLK(clk), .Q(\ram[10][158] ) );
  DFFX1_HVT \ram_reg[10][157]  ( .D(n2778), .CLK(clk), .Q(\ram[10][157] ) );
  DFFX1_HVT \ram_reg[10][156]  ( .D(n2777), .CLK(clk), .Q(\ram[10][156] ) );
  DFFX1_HVT \ram_reg[10][155]  ( .D(n2776), .CLK(clk), .Q(\ram[10][155] ) );
  DFFX1_HVT \ram_reg[10][154]  ( .D(n2775), .CLK(clk), .Q(\ram[10][154] ) );
  DFFX1_HVT \ram_reg[10][153]  ( .D(n2774), .CLK(clk), .Q(\ram[10][153] ) );
  DFFX1_HVT \ram_reg[10][152]  ( .D(n2773), .CLK(clk), .Q(\ram[10][152] ) );
  DFFX1_HVT \ram_reg[10][151]  ( .D(n2772), .CLK(clk), .Q(\ram[10][151] ) );
  DFFX1_HVT \ram_reg[10][150]  ( .D(n2771), .CLK(clk), .Q(\ram[10][150] ) );
  DFFX1_HVT \ram_reg[10][149]  ( .D(n2770), .CLK(clk), .Q(\ram[10][149] ) );
  DFFX1_HVT \ram_reg[10][148]  ( .D(n2769), .CLK(clk), .Q(\ram[10][148] ) );
  DFFX1_HVT \ram_reg[10][147]  ( .D(n2768), .CLK(clk), .Q(\ram[10][147] ) );
  DFFX1_HVT \ram_reg[10][146]  ( .D(n2767), .CLK(clk), .Q(\ram[10][146] ) );
  DFFX1_HVT \ram_reg[10][145]  ( .D(n2766), .CLK(clk), .Q(\ram[10][145] ) );
  DFFX1_HVT \ram_reg[10][144]  ( .D(n2765), .CLK(clk), .Q(\ram[10][144] ) );
  DFFX1_HVT \ram_reg[10][143]  ( .D(n2764), .CLK(clk), .Q(\ram[10][143] ) );
  DFFX1_HVT \ram_reg[10][142]  ( .D(n2763), .CLK(clk), .Q(\ram[10][142] ) );
  DFFX1_HVT \ram_reg[10][141]  ( .D(n2762), .CLK(clk), .Q(\ram[10][141] ) );
  DFFX1_HVT \ram_reg[10][140]  ( .D(n2761), .CLK(clk), .Q(\ram[10][140] ) );
  DFFX1_HVT \ram_reg[10][139]  ( .D(n2760), .CLK(clk), .Q(\ram[10][139] ) );
  DFFX1_HVT \ram_reg[10][138]  ( .D(n2759), .CLK(clk), .Q(\ram[10][138] ) );
  DFFX1_HVT \ram_reg[10][137]  ( .D(n2758), .CLK(clk), .Q(\ram[10][137] ) );
  DFFX1_HVT \ram_reg[10][136]  ( .D(n2757), .CLK(clk), .Q(\ram[10][136] ) );
  DFFX1_HVT \ram_reg[10][135]  ( .D(n2756), .CLK(clk), .Q(\ram[10][135] ) );
  DFFX1_HVT \ram_reg[10][134]  ( .D(n2755), .CLK(clk), .Q(\ram[10][134] ) );
  DFFX1_HVT \ram_reg[10][133]  ( .D(n2754), .CLK(clk), .Q(\ram[10][133] ) );
  DFFX1_HVT \ram_reg[10][132]  ( .D(n2753), .CLK(clk), .Q(\ram[10][132] ) );
  DFFX1_HVT \ram_reg[10][131]  ( .D(n2752), .CLK(clk), .Q(\ram[10][131] ) );
  DFFX1_HVT \ram_reg[10][130]  ( .D(n2751), .CLK(clk), .Q(\ram[10][130] ) );
  DFFX1_HVT \ram_reg[10][129]  ( .D(n2750), .CLK(clk), .Q(\ram[10][129] ) );
  DFFX1_HVT \ram_reg[10][128]  ( .D(n2749), .CLK(clk), .Q(\ram[10][128] ) );
  DFFX1_HVT \ram_reg[10][127]  ( .D(n2748), .CLK(clk), .Q(\ram[10][127] ) );
  DFFX1_HVT \ram_reg[10][126]  ( .D(n2747), .CLK(clk), .Q(\ram[10][126] ) );
  DFFX1_HVT \ram_reg[10][125]  ( .D(n2746), .CLK(clk), .Q(\ram[10][125] ) );
  DFFX1_HVT \ram_reg[10][124]  ( .D(n2745), .CLK(clk), .Q(\ram[10][124] ) );
  DFFX1_HVT \ram_reg[10][123]  ( .D(n2744), .CLK(clk), .Q(\ram[10][123] ) );
  DFFX1_HVT \ram_reg[10][122]  ( .D(n2743), .CLK(clk), .Q(\ram[10][122] ) );
  DFFX1_HVT \ram_reg[10][121]  ( .D(n2742), .CLK(clk), .Q(\ram[10][121] ) );
  DFFX1_HVT \ram_reg[10][120]  ( .D(n2741), .CLK(clk), .Q(\ram[10][120] ) );
  DFFX1_HVT \ram_reg[10][119]  ( .D(n2740), .CLK(clk), .Q(\ram[10][119] ) );
  DFFX1_HVT \ram_reg[10][118]  ( .D(n2739), .CLK(clk), .Q(\ram[10][118] ) );
  DFFX1_HVT \ram_reg[10][117]  ( .D(n2738), .CLK(clk), .Q(\ram[10][117] ) );
  DFFX1_HVT \ram_reg[10][116]  ( .D(n2737), .CLK(clk), .Q(\ram[10][116] ) );
  DFFX1_HVT \ram_reg[10][115]  ( .D(n2736), .CLK(clk), .Q(\ram[10][115] ) );
  DFFX1_HVT \ram_reg[10][114]  ( .D(n2735), .CLK(clk), .Q(\ram[10][114] ) );
  DFFX1_HVT \ram_reg[10][113]  ( .D(n2734), .CLK(clk), .Q(\ram[10][113] ) );
  DFFX1_HVT \ram_reg[10][112]  ( .D(n2733), .CLK(clk), .Q(\ram[10][112] ) );
  DFFX1_HVT \ram_reg[10][111]  ( .D(n2732), .CLK(clk), .Q(\ram[10][111] ) );
  DFFX1_HVT \ram_reg[10][110]  ( .D(n2731), .CLK(clk), .Q(\ram[10][110] ) );
  DFFX1_HVT \ram_reg[10][109]  ( .D(n2730), .CLK(clk), .Q(\ram[10][109] ) );
  DFFX1_HVT \ram_reg[10][108]  ( .D(n2729), .CLK(clk), .Q(\ram[10][108] ) );
  DFFX1_HVT \ram_reg[10][107]  ( .D(n2728), .CLK(clk), .Q(\ram[10][107] ) );
  DFFX1_HVT \ram_reg[10][106]  ( .D(n2727), .CLK(clk), .Q(\ram[10][106] ) );
  DFFX1_HVT \ram_reg[10][105]  ( .D(n2726), .CLK(clk), .Q(\ram[10][105] ) );
  DFFX1_HVT \ram_reg[10][104]  ( .D(n2725), .CLK(clk), .Q(\ram[10][104] ) );
  DFFX1_HVT \ram_reg[10][103]  ( .D(n2724), .CLK(clk), .Q(\ram[10][103] ) );
  DFFX1_HVT \ram_reg[10][102]  ( .D(n2723), .CLK(clk), .Q(\ram[10][102] ) );
  DFFX1_HVT \ram_reg[10][101]  ( .D(n2722), .CLK(clk), .Q(\ram[10][101] ) );
  DFFX1_HVT \ram_reg[10][100]  ( .D(n2721), .CLK(clk), .Q(\ram[10][100] ) );
  DFFX1_HVT \ram_reg[10][99]  ( .D(n2720), .CLK(clk), .Q(\ram[10][99] ) );
  DFFX1_HVT \ram_reg[10][98]  ( .D(n2719), .CLK(clk), .Q(\ram[10][98] ) );
  DFFX1_HVT \ram_reg[10][97]  ( .D(n2718), .CLK(clk), .Q(\ram[10][97] ) );
  DFFX1_HVT \ram_reg[10][96]  ( .D(n2717), .CLK(clk), .Q(\ram[10][96] ) );
  DFFX1_HVT \ram_reg[10][95]  ( .D(n2716), .CLK(clk), .Q(\ram[10][95] ) );
  DFFX1_HVT \ram_reg[10][94]  ( .D(n2715), .CLK(clk), .Q(\ram[10][94] ) );
  DFFX1_HVT \ram_reg[10][93]  ( .D(n2714), .CLK(clk), .Q(\ram[10][93] ) );
  DFFX1_HVT \ram_reg[10][92]  ( .D(n2713), .CLK(clk), .Q(\ram[10][92] ) );
  DFFX1_HVT \ram_reg[10][91]  ( .D(n2712), .CLK(clk), .Q(\ram[10][91] ) );
  DFFX1_HVT \ram_reg[10][90]  ( .D(n2711), .CLK(clk), .Q(\ram[10][90] ) );
  DFFX1_HVT \ram_reg[10][89]  ( .D(n2710), .CLK(clk), .Q(\ram[10][89] ) );
  DFFX1_HVT \ram_reg[10][88]  ( .D(n2709), .CLK(clk), .Q(\ram[10][88] ) );
  DFFX1_HVT \ram_reg[10][87]  ( .D(n2708), .CLK(clk), .Q(\ram[10][87] ) );
  DFFX1_HVT \ram_reg[10][86]  ( .D(n2707), .CLK(clk), .Q(\ram[10][86] ) );
  DFFX1_HVT \ram_reg[10][85]  ( .D(n2706), .CLK(clk), .Q(\ram[10][85] ) );
  DFFX1_HVT \ram_reg[10][84]  ( .D(n2705), .CLK(clk), .Q(\ram[10][84] ) );
  DFFX1_HVT \ram_reg[10][83]  ( .D(n2704), .CLK(clk), .Q(\ram[10][83] ) );
  DFFX1_HVT \ram_reg[10][82]  ( .D(n2703), .CLK(clk), .Q(\ram[10][82] ) );
  DFFX1_HVT \ram_reg[10][81]  ( .D(n2702), .CLK(clk), .Q(\ram[10][81] ) );
  DFFX1_HVT \ram_reg[10][80]  ( .D(n2701), .CLK(clk), .Q(\ram[10][80] ) );
  DFFX1_HVT \ram_reg[10][79]  ( .D(n2700), .CLK(clk), .Q(\ram[10][79] ) );
  DFFX1_HVT \ram_reg[10][78]  ( .D(n2699), .CLK(clk), .Q(\ram[10][78] ) );
  DFFX1_HVT \ram_reg[10][77]  ( .D(n2698), .CLK(clk), .Q(\ram[10][77] ) );
  DFFX1_HVT \ram_reg[10][76]  ( .D(n2697), .CLK(clk), .Q(\ram[10][76] ) );
  DFFX1_HVT \ram_reg[10][75]  ( .D(n2696), .CLK(clk), .Q(\ram[10][75] ) );
  DFFX1_HVT \ram_reg[10][74]  ( .D(n2695), .CLK(clk), .Q(\ram[10][74] ) );
  DFFX1_HVT \ram_reg[10][73]  ( .D(n2694), .CLK(clk), .Q(\ram[10][73] ) );
  DFFX1_HVT \ram_reg[10][72]  ( .D(n2693), .CLK(clk), .Q(\ram[10][72] ) );
  DFFX1_HVT \ram_reg[10][71]  ( .D(n2692), .CLK(clk), .Q(\ram[10][71] ) );
  DFFX1_HVT \ram_reg[10][70]  ( .D(n2691), .CLK(clk), .Q(\ram[10][70] ) );
  DFFX1_HVT \ram_reg[10][69]  ( .D(n2690), .CLK(clk), .Q(\ram[10][69] ) );
  DFFX1_HVT \ram_reg[10][68]  ( .D(n2689), .CLK(clk), .Q(\ram[10][68] ) );
  DFFX1_HVT \ram_reg[10][67]  ( .D(n2688), .CLK(clk), .Q(\ram[10][67] ) );
  DFFX1_HVT \ram_reg[10][66]  ( .D(n2687), .CLK(clk), .Q(\ram[10][66] ) );
  DFFX1_HVT \ram_reg[10][65]  ( .D(n2686), .CLK(clk), .Q(\ram[10][65] ) );
  DFFX1_HVT \ram_reg[10][64]  ( .D(n2685), .CLK(clk), .Q(\ram[10][64] ) );
  DFFX1_HVT \ram_reg[10][63]  ( .D(n2684), .CLK(clk), .Q(\ram[10][63] ) );
  DFFX1_HVT \ram_reg[10][62]  ( .D(n2683), .CLK(clk), .Q(\ram[10][62] ) );
  DFFX1_HVT \ram_reg[10][61]  ( .D(n2682), .CLK(clk), .Q(\ram[10][61] ) );
  DFFX1_HVT \ram_reg[10][60]  ( .D(n2681), .CLK(clk), .Q(\ram[10][60] ) );
  DFFX1_HVT \ram_reg[10][59]  ( .D(n2680), .CLK(clk), .Q(\ram[10][59] ) );
  DFFX1_HVT \ram_reg[10][58]  ( .D(n2679), .CLK(clk), .Q(\ram[10][58] ) );
  DFFX1_HVT \ram_reg[10][57]  ( .D(n2678), .CLK(clk), .Q(\ram[10][57] ) );
  DFFX1_HVT \ram_reg[10][56]  ( .D(n2677), .CLK(clk), .Q(\ram[10][56] ) );
  DFFX1_HVT \ram_reg[10][55]  ( .D(n2676), .CLK(clk), .Q(\ram[10][55] ) );
  DFFX1_HVT \ram_reg[10][54]  ( .D(n2675), .CLK(clk), .Q(\ram[10][54] ) );
  DFFX1_HVT \ram_reg[10][53]  ( .D(n2674), .CLK(clk), .Q(\ram[10][53] ) );
  DFFX1_HVT \ram_reg[10][52]  ( .D(n2673), .CLK(clk), .Q(\ram[10][52] ) );
  DFFX1_HVT \ram_reg[10][51]  ( .D(n2672), .CLK(clk), .Q(\ram[10][51] ) );
  DFFX1_HVT \ram_reg[10][50]  ( .D(n2671), .CLK(clk), .Q(\ram[10][50] ) );
  DFFX1_HVT \ram_reg[10][49]  ( .D(n2670), .CLK(clk), .Q(\ram[10][49] ) );
  DFFX1_HVT \ram_reg[10][48]  ( .D(n2669), .CLK(clk), .Q(\ram[10][48] ) );
  DFFX1_HVT \ram_reg[10][47]  ( .D(n2668), .CLK(clk), .Q(\ram[10][47] ) );
  DFFX1_HVT \ram_reg[10][46]  ( .D(n2667), .CLK(clk), .Q(\ram[10][46] ) );
  DFFX1_HVT \ram_reg[10][45]  ( .D(n2666), .CLK(clk), .Q(\ram[10][45] ) );
  DFFX1_HVT \ram_reg[10][44]  ( .D(n2665), .CLK(clk), .Q(\ram[10][44] ) );
  DFFX1_HVT \ram_reg[10][43]  ( .D(n2664), .CLK(clk), .Q(\ram[10][43] ) );
  DFFX1_HVT \ram_reg[10][42]  ( .D(n2663), .CLK(clk), .Q(\ram[10][42] ) );
  DFFX1_HVT \ram_reg[10][41]  ( .D(n2662), .CLK(clk), .Q(\ram[10][41] ) );
  DFFX1_HVT \ram_reg[10][40]  ( .D(n2661), .CLK(clk), .Q(\ram[10][40] ) );
  DFFX1_HVT \ram_reg[10][39]  ( .D(n2660), .CLK(clk), .Q(\ram[10][39] ) );
  DFFX1_HVT \ram_reg[10][38]  ( .D(n2659), .CLK(clk), .Q(\ram[10][38] ) );
  DFFX1_HVT \ram_reg[10][37]  ( .D(n2658), .CLK(clk), .Q(\ram[10][37] ) );
  DFFX1_HVT \ram_reg[10][36]  ( .D(n2657), .CLK(clk), .Q(\ram[10][36] ) );
  DFFX1_HVT \ram_reg[10][35]  ( .D(n2656), .CLK(clk), .Q(\ram[10][35] ) );
  DFFX1_HVT \ram_reg[10][34]  ( .D(n2655), .CLK(clk), .Q(\ram[10][34] ) );
  DFFX1_HVT \ram_reg[10][33]  ( .D(n2654), .CLK(clk), .Q(\ram[10][33] ) );
  DFFX1_HVT \ram_reg[10][32]  ( .D(n2653), .CLK(clk), .Q(\ram[10][32] ) );
  DFFX1_HVT \ram_reg[10][31]  ( .D(n2652), .CLK(clk), .Q(\ram[10][31] ) );
  DFFX1_HVT \ram_reg[10][30]  ( .D(n2651), .CLK(clk), .Q(\ram[10][30] ) );
  DFFX1_HVT \ram_reg[10][29]  ( .D(n2650), .CLK(clk), .Q(\ram[10][29] ) );
  DFFX1_HVT \ram_reg[10][28]  ( .D(n2649), .CLK(clk), .Q(\ram[10][28] ) );
  DFFX1_HVT \ram_reg[10][27]  ( .D(n2648), .CLK(clk), .Q(\ram[10][27] ) );
  DFFX1_HVT \ram_reg[10][26]  ( .D(n2647), .CLK(clk), .Q(\ram[10][26] ) );
  DFFX1_HVT \ram_reg[10][25]  ( .D(n2646), .CLK(clk), .Q(\ram[10][25] ) );
  DFFX1_HVT \ram_reg[10][24]  ( .D(n2645), .CLK(clk), .Q(\ram[10][24] ) );
  DFFX1_HVT \ram_reg[10][23]  ( .D(n2644), .CLK(clk), .Q(\ram[10][23] ) );
  DFFX1_HVT \ram_reg[10][22]  ( .D(n2643), .CLK(clk), .Q(\ram[10][22] ) );
  DFFX1_HVT \ram_reg[10][21]  ( .D(n2642), .CLK(clk), .Q(\ram[10][21] ) );
  DFFX1_HVT \ram_reg[10][20]  ( .D(n2641), .CLK(clk), .Q(\ram[10][20] ) );
  DFFX1_HVT \ram_reg[10][19]  ( .D(n2640), .CLK(clk), .Q(\ram[10][19] ) );
  DFFX1_HVT \ram_reg[10][18]  ( .D(n2639), .CLK(clk), .Q(\ram[10][18] ) );
  DFFX1_HVT \ram_reg[10][17]  ( .D(n2638), .CLK(clk), .Q(\ram[10][17] ) );
  DFFX1_HVT \ram_reg[10][16]  ( .D(n2637), .CLK(clk), .Q(\ram[10][16] ) );
  DFFX1_HVT \ram_reg[10][15]  ( .D(n2636), .CLK(clk), .Q(\ram[10][15] ) );
  DFFX1_HVT \ram_reg[10][14]  ( .D(n2635), .CLK(clk), .Q(\ram[10][14] ) );
  DFFX1_HVT \ram_reg[10][13]  ( .D(n2634), .CLK(clk), .Q(\ram[10][13] ) );
  DFFX1_HVT \ram_reg[10][12]  ( .D(n2633), .CLK(clk), .Q(\ram[10][12] ) );
  DFFX1_HVT \ram_reg[10][11]  ( .D(n2632), .CLK(clk), .Q(\ram[10][11] ) );
  DFFX1_HVT \ram_reg[10][10]  ( .D(n2631), .CLK(clk), .Q(\ram[10][10] ) );
  DFFX1_HVT \ram_reg[10][9]  ( .D(n2630), .CLK(clk), .Q(\ram[10][9] ) );
  DFFX1_HVT \ram_reg[10][8]  ( .D(n2629), .CLK(clk), .Q(\ram[10][8] ) );
  DFFX1_HVT \ram_reg[10][7]  ( .D(n2628), .CLK(clk), .Q(\ram[10][7] ) );
  DFFX1_HVT \ram_reg[10][6]  ( .D(n2627), .CLK(clk), .Q(\ram[10][6] ) );
  DFFX1_HVT \ram_reg[10][5]  ( .D(n2626), .CLK(clk), .Q(\ram[10][5] ) );
  DFFX1_HVT \ram_reg[10][4]  ( .D(n2625), .CLK(clk), .Q(\ram[10][4] ) );
  DFFX1_HVT \ram_reg[10][3]  ( .D(n2624), .CLK(clk), .Q(\ram[10][3] ) );
  DFFX1_HVT \ram_reg[10][2]  ( .D(n2623), .CLK(clk), .Q(\ram[10][2] ) );
  DFFX1_HVT \ram_reg[10][1]  ( .D(n2622), .CLK(clk), .Q(\ram[10][1] ) );
  DFFX1_HVT \ram_reg[10][0]  ( .D(n2621), .CLK(clk), .Q(\ram[10][0] ) );
  DFFX1_HVT \ram_reg[9][255]  ( .D(n2620), .CLK(clk), .Q(\ram[9][255] ) );
  DFFX1_HVT \ram_reg[9][254]  ( .D(n2619), .CLK(clk), .Q(\ram[9][254] ) );
  DFFX1_HVT \ram_reg[9][253]  ( .D(n2618), .CLK(clk), .Q(\ram[9][253] ) );
  DFFX1_HVT \ram_reg[9][252]  ( .D(n2617), .CLK(clk), .Q(\ram[9][252] ) );
  DFFX1_HVT \ram_reg[9][251]  ( .D(n2616), .CLK(clk), .Q(\ram[9][251] ) );
  DFFX1_HVT \ram_reg[9][250]  ( .D(n2615), .CLK(clk), .Q(\ram[9][250] ) );
  DFFX1_HVT \ram_reg[9][249]  ( .D(n2614), .CLK(clk), .Q(\ram[9][249] ) );
  DFFX1_HVT \ram_reg[9][248]  ( .D(n2613), .CLK(clk), .Q(\ram[9][248] ) );
  DFFX1_HVT \ram_reg[9][247]  ( .D(n2612), .CLK(clk), .Q(\ram[9][247] ) );
  DFFX1_HVT \ram_reg[9][246]  ( .D(n2611), .CLK(clk), .Q(\ram[9][246] ) );
  DFFX1_HVT \ram_reg[9][245]  ( .D(n2610), .CLK(clk), .Q(\ram[9][245] ) );
  DFFX1_HVT \ram_reg[9][244]  ( .D(n2609), .CLK(clk), .Q(\ram[9][244] ) );
  DFFX1_HVT \ram_reg[9][243]  ( .D(n2608), .CLK(clk), .Q(\ram[9][243] ) );
  DFFX1_HVT \ram_reg[9][242]  ( .D(n2607), .CLK(clk), .Q(\ram[9][242] ) );
  DFFX1_HVT \ram_reg[9][241]  ( .D(n2606), .CLK(clk), .Q(\ram[9][241] ) );
  DFFX1_HVT \ram_reg[9][240]  ( .D(n2605), .CLK(clk), .Q(\ram[9][240] ) );
  DFFX1_HVT \ram_reg[9][239]  ( .D(n2604), .CLK(clk), .Q(\ram[9][239] ) );
  DFFX1_HVT \ram_reg[9][238]  ( .D(n2603), .CLK(clk), .Q(\ram[9][238] ) );
  DFFX1_HVT \ram_reg[9][237]  ( .D(n2602), .CLK(clk), .Q(\ram[9][237] ) );
  DFFX1_HVT \ram_reg[9][236]  ( .D(n2601), .CLK(clk), .Q(\ram[9][236] ) );
  DFFX1_HVT \ram_reg[9][235]  ( .D(n2600), .CLK(clk), .Q(\ram[9][235] ) );
  DFFX1_HVT \ram_reg[9][234]  ( .D(n2599), .CLK(clk), .Q(\ram[9][234] ) );
  DFFX1_HVT \ram_reg[9][233]  ( .D(n2598), .CLK(clk), .Q(\ram[9][233] ) );
  DFFX1_HVT \ram_reg[9][232]  ( .D(n2597), .CLK(clk), .Q(\ram[9][232] ) );
  DFFX1_HVT \ram_reg[9][231]  ( .D(n2596), .CLK(clk), .Q(\ram[9][231] ) );
  DFFX1_HVT \ram_reg[9][230]  ( .D(n2595), .CLK(clk), .Q(\ram[9][230] ) );
  DFFX1_HVT \ram_reg[9][229]  ( .D(n2594), .CLK(clk), .Q(\ram[9][229] ) );
  DFFX1_HVT \ram_reg[9][228]  ( .D(n2593), .CLK(clk), .Q(\ram[9][228] ) );
  DFFX1_HVT \ram_reg[9][227]  ( .D(n2592), .CLK(clk), .Q(\ram[9][227] ) );
  DFFX1_HVT \ram_reg[9][226]  ( .D(n2591), .CLK(clk), .Q(\ram[9][226] ) );
  DFFX1_HVT \ram_reg[9][225]  ( .D(n2590), .CLK(clk), .Q(\ram[9][225] ) );
  DFFX1_HVT \ram_reg[9][224]  ( .D(n2589), .CLK(clk), .Q(\ram[9][224] ) );
  DFFX1_HVT \ram_reg[9][223]  ( .D(n2588), .CLK(clk), .Q(\ram[9][223] ) );
  DFFX1_HVT \ram_reg[9][222]  ( .D(n2587), .CLK(clk), .Q(\ram[9][222] ) );
  DFFX1_HVT \ram_reg[9][221]  ( .D(n2586), .CLK(clk), .Q(\ram[9][221] ) );
  DFFX1_HVT \ram_reg[9][220]  ( .D(n2585), .CLK(clk), .Q(\ram[9][220] ) );
  DFFX1_HVT \ram_reg[9][219]  ( .D(n2584), .CLK(clk), .Q(\ram[9][219] ) );
  DFFX1_HVT \ram_reg[9][218]  ( .D(n2583), .CLK(clk), .Q(\ram[9][218] ) );
  DFFX1_HVT \ram_reg[9][217]  ( .D(n2582), .CLK(clk), .Q(\ram[9][217] ) );
  DFFX1_HVT \ram_reg[9][216]  ( .D(n2581), .CLK(clk), .Q(\ram[9][216] ) );
  DFFX1_HVT \ram_reg[9][215]  ( .D(n2580), .CLK(clk), .Q(\ram[9][215] ) );
  DFFX1_HVT \ram_reg[9][214]  ( .D(n2579), .CLK(clk), .Q(\ram[9][214] ) );
  DFFX1_HVT \ram_reg[9][213]  ( .D(n2578), .CLK(clk), .Q(\ram[9][213] ) );
  DFFX1_HVT \ram_reg[9][212]  ( .D(n2577), .CLK(clk), .Q(\ram[9][212] ) );
  DFFX1_HVT \ram_reg[9][211]  ( .D(n2576), .CLK(clk), .Q(\ram[9][211] ) );
  DFFX1_HVT \ram_reg[9][210]  ( .D(n2575), .CLK(clk), .Q(\ram[9][210] ) );
  DFFX1_HVT \ram_reg[9][209]  ( .D(n2574), .CLK(clk), .Q(\ram[9][209] ) );
  DFFX1_HVT \ram_reg[9][208]  ( .D(n2573), .CLK(clk), .Q(\ram[9][208] ) );
  DFFX1_HVT \ram_reg[9][207]  ( .D(n2572), .CLK(clk), .Q(\ram[9][207] ) );
  DFFX1_HVT \ram_reg[9][206]  ( .D(n2571), .CLK(clk), .Q(\ram[9][206] ) );
  DFFX1_HVT \ram_reg[9][205]  ( .D(n2570), .CLK(clk), .Q(\ram[9][205] ) );
  DFFX1_HVT \ram_reg[9][204]  ( .D(n2569), .CLK(clk), .Q(\ram[9][204] ) );
  DFFX1_HVT \ram_reg[9][203]  ( .D(n2568), .CLK(clk), .Q(\ram[9][203] ) );
  DFFX1_HVT \ram_reg[9][202]  ( .D(n2567), .CLK(clk), .Q(\ram[9][202] ) );
  DFFX1_HVT \ram_reg[9][201]  ( .D(n2566), .CLK(clk), .Q(\ram[9][201] ) );
  DFFX1_HVT \ram_reg[9][200]  ( .D(n2565), .CLK(clk), .Q(\ram[9][200] ) );
  DFFX1_HVT \ram_reg[9][199]  ( .D(n2564), .CLK(clk), .Q(\ram[9][199] ) );
  DFFX1_HVT \ram_reg[9][198]  ( .D(n2563), .CLK(clk), .Q(\ram[9][198] ) );
  DFFX1_HVT \ram_reg[9][197]  ( .D(n2562), .CLK(clk), .Q(\ram[9][197] ) );
  DFFX1_HVT \ram_reg[9][196]  ( .D(n2561), .CLK(clk), .Q(\ram[9][196] ) );
  DFFX1_HVT \ram_reg[9][195]  ( .D(n2560), .CLK(clk), .Q(\ram[9][195] ) );
  DFFX1_HVT \ram_reg[9][194]  ( .D(n2559), .CLK(clk), .Q(\ram[9][194] ) );
  DFFX1_HVT \ram_reg[9][193]  ( .D(n2558), .CLK(clk), .Q(\ram[9][193] ) );
  DFFX1_HVT \ram_reg[9][192]  ( .D(n2557), .CLK(clk), .Q(\ram[9][192] ) );
  DFFX1_HVT \ram_reg[9][191]  ( .D(n2556), .CLK(clk), .Q(\ram[9][191] ) );
  DFFX1_HVT \ram_reg[9][190]  ( .D(n2555), .CLK(clk), .Q(\ram[9][190] ) );
  DFFX1_HVT \ram_reg[9][189]  ( .D(n2554), .CLK(clk), .Q(\ram[9][189] ) );
  DFFX1_HVT \ram_reg[9][188]  ( .D(n2553), .CLK(clk), .Q(\ram[9][188] ) );
  DFFX1_HVT \ram_reg[9][187]  ( .D(n2552), .CLK(clk), .Q(\ram[9][187] ) );
  DFFX1_HVT \ram_reg[9][186]  ( .D(n2551), .CLK(clk), .Q(\ram[9][186] ) );
  DFFX1_HVT \ram_reg[9][185]  ( .D(n2550), .CLK(clk), .Q(\ram[9][185] ) );
  DFFX1_HVT \ram_reg[9][184]  ( .D(n2549), .CLK(clk), .Q(\ram[9][184] ) );
  DFFX1_HVT \ram_reg[9][183]  ( .D(n2548), .CLK(clk), .Q(\ram[9][183] ) );
  DFFX1_HVT \ram_reg[9][182]  ( .D(n2547), .CLK(clk), .Q(\ram[9][182] ) );
  DFFX1_HVT \ram_reg[9][181]  ( .D(n2546), .CLK(clk), .Q(\ram[9][181] ) );
  DFFX1_HVT \ram_reg[9][180]  ( .D(n2545), .CLK(clk), .Q(\ram[9][180] ) );
  DFFX1_HVT \ram_reg[9][179]  ( .D(n2544), .CLK(clk), .Q(\ram[9][179] ) );
  DFFX1_HVT \ram_reg[9][178]  ( .D(n2543), .CLK(clk), .Q(\ram[9][178] ) );
  DFFX1_HVT \ram_reg[9][177]  ( .D(n2542), .CLK(clk), .Q(\ram[9][177] ) );
  DFFX1_HVT \ram_reg[9][176]  ( .D(n2541), .CLK(clk), .Q(\ram[9][176] ) );
  DFFX1_HVT \ram_reg[9][175]  ( .D(n2540), .CLK(clk), .Q(\ram[9][175] ) );
  DFFX1_HVT \ram_reg[9][174]  ( .D(n2539), .CLK(clk), .Q(\ram[9][174] ) );
  DFFX1_HVT \ram_reg[9][173]  ( .D(n2538), .CLK(clk), .Q(\ram[9][173] ) );
  DFFX1_HVT \ram_reg[9][172]  ( .D(n2537), .CLK(clk), .Q(\ram[9][172] ) );
  DFFX1_HVT \ram_reg[9][171]  ( .D(n2536), .CLK(clk), .Q(\ram[9][171] ) );
  DFFX1_HVT \ram_reg[9][170]  ( .D(n2535), .CLK(clk), .Q(\ram[9][170] ) );
  DFFX1_HVT \ram_reg[9][169]  ( .D(n2534), .CLK(clk), .Q(\ram[9][169] ) );
  DFFX1_HVT \ram_reg[9][168]  ( .D(n2533), .CLK(clk), .Q(\ram[9][168] ) );
  DFFX1_HVT \ram_reg[9][167]  ( .D(n2532), .CLK(clk), .Q(\ram[9][167] ) );
  DFFX1_HVT \ram_reg[9][166]  ( .D(n2531), .CLK(clk), .Q(\ram[9][166] ) );
  DFFX1_HVT \ram_reg[9][165]  ( .D(n2530), .CLK(clk), .Q(\ram[9][165] ) );
  DFFX1_HVT \ram_reg[9][164]  ( .D(n2529), .CLK(clk), .Q(\ram[9][164] ) );
  DFFX1_HVT \ram_reg[9][163]  ( .D(n2528), .CLK(clk), .Q(\ram[9][163] ) );
  DFFX1_HVT \ram_reg[9][162]  ( .D(n2527), .CLK(clk), .Q(\ram[9][162] ) );
  DFFX1_HVT \ram_reg[9][161]  ( .D(n2526), .CLK(clk), .Q(\ram[9][161] ) );
  DFFX1_HVT \ram_reg[9][160]  ( .D(n2525), .CLK(clk), .Q(\ram[9][160] ) );
  DFFX1_HVT \ram_reg[9][159]  ( .D(n2524), .CLK(clk), .Q(\ram[9][159] ) );
  DFFX1_HVT \ram_reg[9][158]  ( .D(n2523), .CLK(clk), .Q(\ram[9][158] ) );
  DFFX1_HVT \ram_reg[9][157]  ( .D(n2522), .CLK(clk), .Q(\ram[9][157] ) );
  DFFX1_HVT \ram_reg[9][156]  ( .D(n2521), .CLK(clk), .Q(\ram[9][156] ) );
  DFFX1_HVT \ram_reg[9][155]  ( .D(n2520), .CLK(clk), .Q(\ram[9][155] ) );
  DFFX1_HVT \ram_reg[9][154]  ( .D(n2519), .CLK(clk), .Q(\ram[9][154] ) );
  DFFX1_HVT \ram_reg[9][153]  ( .D(n2518), .CLK(clk), .Q(\ram[9][153] ) );
  DFFX1_HVT \ram_reg[9][152]  ( .D(n2517), .CLK(clk), .Q(\ram[9][152] ) );
  DFFX1_HVT \ram_reg[9][151]  ( .D(n2516), .CLK(clk), .Q(\ram[9][151] ) );
  DFFX1_HVT \ram_reg[9][150]  ( .D(n2515), .CLK(clk), .Q(\ram[9][150] ) );
  DFFX1_HVT \ram_reg[9][149]  ( .D(n2514), .CLK(clk), .Q(\ram[9][149] ) );
  DFFX1_HVT \ram_reg[9][148]  ( .D(n2513), .CLK(clk), .Q(\ram[9][148] ) );
  DFFX1_HVT \ram_reg[9][147]  ( .D(n2512), .CLK(clk), .Q(\ram[9][147] ) );
  DFFX1_HVT \ram_reg[9][146]  ( .D(n2511), .CLK(clk), .Q(\ram[9][146] ) );
  DFFX1_HVT \ram_reg[9][145]  ( .D(n2510), .CLK(clk), .Q(\ram[9][145] ) );
  DFFX1_HVT \ram_reg[9][144]  ( .D(n2509), .CLK(clk), .Q(\ram[9][144] ) );
  DFFX1_HVT \ram_reg[9][143]  ( .D(n2508), .CLK(clk), .Q(\ram[9][143] ) );
  DFFX1_HVT \ram_reg[9][142]  ( .D(n2507), .CLK(clk), .Q(\ram[9][142] ) );
  DFFX1_HVT \ram_reg[9][141]  ( .D(n2506), .CLK(clk), .Q(\ram[9][141] ) );
  DFFX1_HVT \ram_reg[9][140]  ( .D(n2505), .CLK(clk), .Q(\ram[9][140] ) );
  DFFX1_HVT \ram_reg[9][139]  ( .D(n2504), .CLK(clk), .Q(\ram[9][139] ) );
  DFFX1_HVT \ram_reg[9][138]  ( .D(n2503), .CLK(clk), .Q(\ram[9][138] ) );
  DFFX1_HVT \ram_reg[9][137]  ( .D(n2502), .CLK(clk), .Q(\ram[9][137] ) );
  DFFX1_HVT \ram_reg[9][136]  ( .D(n2501), .CLK(clk), .Q(\ram[9][136] ) );
  DFFX1_HVT \ram_reg[9][135]  ( .D(n2500), .CLK(clk), .Q(\ram[9][135] ) );
  DFFX1_HVT \ram_reg[9][134]  ( .D(n2499), .CLK(clk), .Q(\ram[9][134] ) );
  DFFX1_HVT \ram_reg[9][133]  ( .D(n2498), .CLK(clk), .Q(\ram[9][133] ) );
  DFFX1_HVT \ram_reg[9][132]  ( .D(n2497), .CLK(clk), .Q(\ram[9][132] ) );
  DFFX1_HVT \ram_reg[9][131]  ( .D(n2496), .CLK(clk), .Q(\ram[9][131] ) );
  DFFX1_HVT \ram_reg[9][130]  ( .D(n2495), .CLK(clk), .Q(\ram[9][130] ) );
  DFFX1_HVT \ram_reg[9][129]  ( .D(n2494), .CLK(clk), .Q(\ram[9][129] ) );
  DFFX1_HVT \ram_reg[9][128]  ( .D(n2493), .CLK(clk), .Q(\ram[9][128] ) );
  DFFX1_HVT \ram_reg[9][127]  ( .D(n2492), .CLK(clk), .Q(\ram[9][127] ) );
  DFFX1_HVT \ram_reg[9][126]  ( .D(n2491), .CLK(clk), .Q(\ram[9][126] ) );
  DFFX1_HVT \ram_reg[9][125]  ( .D(n2490), .CLK(clk), .Q(\ram[9][125] ) );
  DFFX1_HVT \ram_reg[9][124]  ( .D(n2489), .CLK(clk), .Q(\ram[9][124] ) );
  DFFX1_HVT \ram_reg[9][123]  ( .D(n2488), .CLK(clk), .Q(\ram[9][123] ) );
  DFFX1_HVT \ram_reg[9][122]  ( .D(n2487), .CLK(clk), .Q(\ram[9][122] ) );
  DFFX1_HVT \ram_reg[9][121]  ( .D(n2486), .CLK(clk), .Q(\ram[9][121] ) );
  DFFX1_HVT \ram_reg[9][120]  ( .D(n2485), .CLK(clk), .Q(\ram[9][120] ) );
  DFFX1_HVT \ram_reg[9][119]  ( .D(n2484), .CLK(clk), .Q(\ram[9][119] ) );
  DFFX1_HVT \ram_reg[9][118]  ( .D(n2483), .CLK(clk), .Q(\ram[9][118] ) );
  DFFX1_HVT \ram_reg[9][117]  ( .D(n2482), .CLK(clk), .Q(\ram[9][117] ) );
  DFFX1_HVT \ram_reg[9][116]  ( .D(n2481), .CLK(clk), .Q(\ram[9][116] ) );
  DFFX1_HVT \ram_reg[9][115]  ( .D(n2480), .CLK(clk), .Q(\ram[9][115] ) );
  DFFX1_HVT \ram_reg[9][114]  ( .D(n2479), .CLK(clk), .Q(\ram[9][114] ) );
  DFFX1_HVT \ram_reg[9][113]  ( .D(n2478), .CLK(clk), .Q(\ram[9][113] ) );
  DFFX1_HVT \ram_reg[9][112]  ( .D(n2477), .CLK(clk), .Q(\ram[9][112] ) );
  DFFX1_HVT \ram_reg[9][111]  ( .D(n2476), .CLK(clk), .Q(\ram[9][111] ) );
  DFFX1_HVT \ram_reg[9][110]  ( .D(n2475), .CLK(clk), .Q(\ram[9][110] ) );
  DFFX1_HVT \ram_reg[9][109]  ( .D(n2474), .CLK(clk), .Q(\ram[9][109] ) );
  DFFX1_HVT \ram_reg[9][108]  ( .D(n2473), .CLK(clk), .Q(\ram[9][108] ) );
  DFFX1_HVT \ram_reg[9][107]  ( .D(n2472), .CLK(clk), .Q(\ram[9][107] ) );
  DFFX1_HVT \ram_reg[9][106]  ( .D(n2471), .CLK(clk), .Q(\ram[9][106] ) );
  DFFX1_HVT \ram_reg[9][105]  ( .D(n2470), .CLK(clk), .Q(\ram[9][105] ) );
  DFFX1_HVT \ram_reg[9][104]  ( .D(n2469), .CLK(clk), .Q(\ram[9][104] ) );
  DFFX1_HVT \ram_reg[9][103]  ( .D(n2468), .CLK(clk), .Q(\ram[9][103] ) );
  DFFX1_HVT \ram_reg[9][102]  ( .D(n2467), .CLK(clk), .Q(\ram[9][102] ) );
  DFFX1_HVT \ram_reg[9][101]  ( .D(n2466), .CLK(clk), .Q(\ram[9][101] ) );
  DFFX1_HVT \ram_reg[9][100]  ( .D(n2465), .CLK(clk), .Q(\ram[9][100] ) );
  DFFX1_HVT \ram_reg[9][99]  ( .D(n2464), .CLK(clk), .Q(\ram[9][99] ) );
  DFFX1_HVT \ram_reg[9][98]  ( .D(n2463), .CLK(clk), .Q(\ram[9][98] ) );
  DFFX1_HVT \ram_reg[9][97]  ( .D(n2462), .CLK(clk), .Q(\ram[9][97] ) );
  DFFX1_HVT \ram_reg[9][96]  ( .D(n2461), .CLK(clk), .Q(\ram[9][96] ) );
  DFFX1_HVT \ram_reg[9][95]  ( .D(n2460), .CLK(clk), .Q(\ram[9][95] ) );
  DFFX1_HVT \ram_reg[9][94]  ( .D(n2459), .CLK(clk), .Q(\ram[9][94] ) );
  DFFX1_HVT \ram_reg[9][93]  ( .D(n2458), .CLK(clk), .Q(\ram[9][93] ) );
  DFFX1_HVT \ram_reg[9][92]  ( .D(n2457), .CLK(clk), .Q(\ram[9][92] ) );
  DFFX1_HVT \ram_reg[9][91]  ( .D(n2456), .CLK(clk), .Q(\ram[9][91] ) );
  DFFX1_HVT \ram_reg[9][90]  ( .D(n2455), .CLK(clk), .Q(\ram[9][90] ) );
  DFFX1_HVT \ram_reg[9][89]  ( .D(n2454), .CLK(clk), .Q(\ram[9][89] ) );
  DFFX1_HVT \ram_reg[9][88]  ( .D(n2453), .CLK(clk), .Q(\ram[9][88] ) );
  DFFX1_HVT \ram_reg[9][87]  ( .D(n2452), .CLK(clk), .Q(\ram[9][87] ) );
  DFFX1_HVT \ram_reg[9][86]  ( .D(n2451), .CLK(clk), .Q(\ram[9][86] ) );
  DFFX1_HVT \ram_reg[9][85]  ( .D(n2450), .CLK(clk), .Q(\ram[9][85] ) );
  DFFX1_HVT \ram_reg[9][84]  ( .D(n2449), .CLK(clk), .Q(\ram[9][84] ) );
  DFFX1_HVT \ram_reg[9][83]  ( .D(n2448), .CLK(clk), .Q(\ram[9][83] ) );
  DFFX1_HVT \ram_reg[9][82]  ( .D(n2447), .CLK(clk), .Q(\ram[9][82] ) );
  DFFX1_HVT \ram_reg[9][81]  ( .D(n2446), .CLK(clk), .Q(\ram[9][81] ) );
  DFFX1_HVT \ram_reg[9][80]  ( .D(n2445), .CLK(clk), .Q(\ram[9][80] ) );
  DFFX1_HVT \ram_reg[9][79]  ( .D(n2444), .CLK(clk), .Q(\ram[9][79] ) );
  DFFX1_HVT \ram_reg[9][78]  ( .D(n2443), .CLK(clk), .Q(\ram[9][78] ) );
  DFFX1_HVT \ram_reg[9][77]  ( .D(n2442), .CLK(clk), .Q(\ram[9][77] ) );
  DFFX1_HVT \ram_reg[9][76]  ( .D(n2441), .CLK(clk), .Q(\ram[9][76] ) );
  DFFX1_HVT \ram_reg[9][75]  ( .D(n2440), .CLK(clk), .Q(\ram[9][75] ) );
  DFFX1_HVT \ram_reg[9][74]  ( .D(n2439), .CLK(clk), .Q(\ram[9][74] ) );
  DFFX1_HVT \ram_reg[9][73]  ( .D(n2438), .CLK(clk), .Q(\ram[9][73] ) );
  DFFX1_HVT \ram_reg[9][72]  ( .D(n2437), .CLK(clk), .Q(\ram[9][72] ) );
  DFFX1_HVT \ram_reg[9][71]  ( .D(n2436), .CLK(clk), .Q(\ram[9][71] ) );
  DFFX1_HVT \ram_reg[9][70]  ( .D(n2435), .CLK(clk), .Q(\ram[9][70] ) );
  DFFX1_HVT \ram_reg[9][69]  ( .D(n2434), .CLK(clk), .Q(\ram[9][69] ) );
  DFFX1_HVT \ram_reg[9][68]  ( .D(n2433), .CLK(clk), .Q(\ram[9][68] ) );
  DFFX1_HVT \ram_reg[9][67]  ( .D(n2432), .CLK(clk), .Q(\ram[9][67] ) );
  DFFX1_HVT \ram_reg[9][66]  ( .D(n2431), .CLK(clk), .Q(\ram[9][66] ) );
  DFFX1_HVT \ram_reg[9][65]  ( .D(n2430), .CLK(clk), .Q(\ram[9][65] ) );
  DFFX1_HVT \ram_reg[9][64]  ( .D(n2429), .CLK(clk), .Q(\ram[9][64] ) );
  DFFX1_HVT \ram_reg[9][63]  ( .D(n2428), .CLK(clk), .Q(\ram[9][63] ) );
  DFFX1_HVT \ram_reg[9][62]  ( .D(n2427), .CLK(clk), .Q(\ram[9][62] ) );
  DFFX1_HVT \ram_reg[9][61]  ( .D(n2426), .CLK(clk), .Q(\ram[9][61] ) );
  DFFX1_HVT \ram_reg[9][60]  ( .D(n2425), .CLK(clk), .Q(\ram[9][60] ) );
  DFFX1_HVT \ram_reg[9][59]  ( .D(n2424), .CLK(clk), .Q(\ram[9][59] ) );
  DFFX1_HVT \ram_reg[9][58]  ( .D(n2423), .CLK(clk), .Q(\ram[9][58] ) );
  DFFX1_HVT \ram_reg[9][57]  ( .D(n2422), .CLK(clk), .Q(\ram[9][57] ) );
  DFFX1_HVT \ram_reg[9][56]  ( .D(n2421), .CLK(clk), .Q(\ram[9][56] ) );
  DFFX1_HVT \ram_reg[9][55]  ( .D(n2420), .CLK(clk), .Q(\ram[9][55] ) );
  DFFX1_HVT \ram_reg[9][54]  ( .D(n2419), .CLK(clk), .Q(\ram[9][54] ) );
  DFFX1_HVT \ram_reg[9][53]  ( .D(n2418), .CLK(clk), .Q(\ram[9][53] ) );
  DFFX1_HVT \ram_reg[9][52]  ( .D(n2417), .CLK(clk), .Q(\ram[9][52] ) );
  DFFX1_HVT \ram_reg[9][51]  ( .D(n2416), .CLK(clk), .Q(\ram[9][51] ) );
  DFFX1_HVT \ram_reg[9][50]  ( .D(n2415), .CLK(clk), .Q(\ram[9][50] ) );
  DFFX1_HVT \ram_reg[9][49]  ( .D(n2414), .CLK(clk), .Q(\ram[9][49] ) );
  DFFX1_HVT \ram_reg[9][48]  ( .D(n2413), .CLK(clk), .Q(\ram[9][48] ) );
  DFFX1_HVT \ram_reg[9][47]  ( .D(n2412), .CLK(clk), .Q(\ram[9][47] ) );
  DFFX1_HVT \ram_reg[9][46]  ( .D(n2411), .CLK(clk), .Q(\ram[9][46] ) );
  DFFX1_HVT \ram_reg[9][45]  ( .D(n2410), .CLK(clk), .Q(\ram[9][45] ) );
  DFFX1_HVT \ram_reg[9][44]  ( .D(n2409), .CLK(clk), .Q(\ram[9][44] ) );
  DFFX1_HVT \ram_reg[9][43]  ( .D(n2408), .CLK(clk), .Q(\ram[9][43] ) );
  DFFX1_HVT \ram_reg[9][42]  ( .D(n2407), .CLK(clk), .Q(\ram[9][42] ) );
  DFFX1_HVT \ram_reg[9][41]  ( .D(n2406), .CLK(clk), .Q(\ram[9][41] ) );
  DFFX1_HVT \ram_reg[9][40]  ( .D(n2405), .CLK(clk), .Q(\ram[9][40] ) );
  DFFX1_HVT \ram_reg[9][39]  ( .D(n2404), .CLK(clk), .Q(\ram[9][39] ) );
  DFFX1_HVT \ram_reg[9][38]  ( .D(n2403), .CLK(clk), .Q(\ram[9][38] ) );
  DFFX1_HVT \ram_reg[9][37]  ( .D(n2402), .CLK(clk), .Q(\ram[9][37] ) );
  DFFX1_HVT \ram_reg[9][36]  ( .D(n2401), .CLK(clk), .Q(\ram[9][36] ) );
  DFFX1_HVT \ram_reg[9][35]  ( .D(n2400), .CLK(clk), .Q(\ram[9][35] ) );
  DFFX1_HVT \ram_reg[9][34]  ( .D(n2399), .CLK(clk), .Q(\ram[9][34] ) );
  DFFX1_HVT \ram_reg[9][33]  ( .D(n2398), .CLK(clk), .Q(\ram[9][33] ) );
  DFFX1_HVT \ram_reg[9][32]  ( .D(n2397), .CLK(clk), .Q(\ram[9][32] ) );
  DFFX1_HVT \ram_reg[9][31]  ( .D(n2396), .CLK(clk), .Q(\ram[9][31] ) );
  DFFX1_HVT \ram_reg[9][30]  ( .D(n2395), .CLK(clk), .Q(\ram[9][30] ) );
  DFFX1_HVT \ram_reg[9][29]  ( .D(n2394), .CLK(clk), .Q(\ram[9][29] ) );
  DFFX1_HVT \ram_reg[9][28]  ( .D(n2393), .CLK(clk), .Q(\ram[9][28] ) );
  DFFX1_HVT \ram_reg[9][27]  ( .D(n2392), .CLK(clk), .Q(\ram[9][27] ) );
  DFFX1_HVT \ram_reg[9][26]  ( .D(n2391), .CLK(clk), .Q(\ram[9][26] ) );
  DFFX1_HVT \ram_reg[9][25]  ( .D(n2390), .CLK(clk), .Q(\ram[9][25] ) );
  DFFX1_HVT \ram_reg[9][24]  ( .D(n2389), .CLK(clk), .Q(\ram[9][24] ) );
  DFFX1_HVT \ram_reg[9][23]  ( .D(n2388), .CLK(clk), .Q(\ram[9][23] ) );
  DFFX1_HVT \ram_reg[9][22]  ( .D(n2387), .CLK(clk), .Q(\ram[9][22] ) );
  DFFX1_HVT \ram_reg[9][21]  ( .D(n2386), .CLK(clk), .Q(\ram[9][21] ) );
  DFFX1_HVT \ram_reg[9][20]  ( .D(n2385), .CLK(clk), .Q(\ram[9][20] ) );
  DFFX1_HVT \ram_reg[9][19]  ( .D(n2384), .CLK(clk), .Q(\ram[9][19] ) );
  DFFX1_HVT \ram_reg[9][18]  ( .D(n2383), .CLK(clk), .Q(\ram[9][18] ) );
  DFFX1_HVT \ram_reg[9][17]  ( .D(n2382), .CLK(clk), .Q(\ram[9][17] ) );
  DFFX1_HVT \ram_reg[9][16]  ( .D(n2381), .CLK(clk), .Q(\ram[9][16] ) );
  DFFX1_HVT \ram_reg[9][15]  ( .D(n2380), .CLK(clk), .Q(\ram[9][15] ) );
  DFFX1_HVT \ram_reg[9][14]  ( .D(n2379), .CLK(clk), .Q(\ram[9][14] ) );
  DFFX1_HVT \ram_reg[9][13]  ( .D(n2378), .CLK(clk), .Q(\ram[9][13] ) );
  DFFX1_HVT \ram_reg[9][12]  ( .D(n2377), .CLK(clk), .Q(\ram[9][12] ) );
  DFFX1_HVT \ram_reg[9][11]  ( .D(n2376), .CLK(clk), .Q(\ram[9][11] ) );
  DFFX1_HVT \ram_reg[9][10]  ( .D(n2375), .CLK(clk), .Q(\ram[9][10] ) );
  DFFX1_HVT \ram_reg[9][9]  ( .D(n2374), .CLK(clk), .Q(\ram[9][9] ) );
  DFFX1_HVT \ram_reg[9][8]  ( .D(n2373), .CLK(clk), .Q(\ram[9][8] ) );
  DFFX1_HVT \ram_reg[9][7]  ( .D(n2372), .CLK(clk), .Q(\ram[9][7] ) );
  DFFX1_HVT \ram_reg[9][6]  ( .D(n2371), .CLK(clk), .Q(\ram[9][6] ) );
  DFFX1_HVT \ram_reg[9][5]  ( .D(n2370), .CLK(clk), .Q(\ram[9][5] ) );
  DFFX1_HVT \ram_reg[9][4]  ( .D(n2369), .CLK(clk), .Q(\ram[9][4] ) );
  DFFX1_HVT \ram_reg[9][3]  ( .D(n2368), .CLK(clk), .Q(\ram[9][3] ) );
  DFFX1_HVT \ram_reg[9][2]  ( .D(n2367), .CLK(clk), .Q(\ram[9][2] ) );
  DFFX1_HVT \ram_reg[9][1]  ( .D(n2366), .CLK(clk), .Q(\ram[9][1] ) );
  DFFX1_HVT \ram_reg[9][0]  ( .D(n2365), .CLK(clk), .Q(\ram[9][0] ) );
  DFFX1_HVT \ram_reg[8][255]  ( .D(n2364), .CLK(clk), .Q(\ram[8][255] ) );
  DFFX1_HVT \ram_reg[8][254]  ( .D(n2363), .CLK(clk), .Q(\ram[8][254] ) );
  DFFX1_HVT \ram_reg[8][253]  ( .D(n2362), .CLK(clk), .Q(\ram[8][253] ) );
  DFFX1_HVT \ram_reg[8][252]  ( .D(n2361), .CLK(clk), .Q(\ram[8][252] ) );
  DFFX1_HVT \ram_reg[8][251]  ( .D(n2360), .CLK(clk), .Q(\ram[8][251] ) );
  DFFX1_HVT \ram_reg[8][250]  ( .D(n2359), .CLK(clk), .Q(\ram[8][250] ) );
  DFFX1_HVT \ram_reg[8][249]  ( .D(n2358), .CLK(clk), .Q(\ram[8][249] ) );
  DFFX1_HVT \ram_reg[8][248]  ( .D(n2357), .CLK(clk), .Q(\ram[8][248] ) );
  DFFX1_HVT \ram_reg[8][247]  ( .D(n2356), .CLK(clk), .Q(\ram[8][247] ) );
  DFFX1_HVT \ram_reg[8][246]  ( .D(n2355), .CLK(clk), .Q(\ram[8][246] ) );
  DFFX1_HVT \ram_reg[8][245]  ( .D(n2354), .CLK(clk), .Q(\ram[8][245] ) );
  DFFX1_HVT \ram_reg[8][244]  ( .D(n2353), .CLK(clk), .Q(\ram[8][244] ) );
  DFFX1_HVT \ram_reg[8][243]  ( .D(n2352), .CLK(clk), .Q(\ram[8][243] ) );
  DFFX1_HVT \ram_reg[8][242]  ( .D(n2351), .CLK(clk), .Q(\ram[8][242] ) );
  DFFX1_HVT \ram_reg[8][241]  ( .D(n2350), .CLK(clk), .Q(\ram[8][241] ) );
  DFFX1_HVT \ram_reg[8][240]  ( .D(n2349), .CLK(clk), .Q(\ram[8][240] ) );
  DFFX1_HVT \ram_reg[8][239]  ( .D(n2348), .CLK(clk), .Q(\ram[8][239] ) );
  DFFX1_HVT \ram_reg[8][238]  ( .D(n2347), .CLK(clk), .Q(\ram[8][238] ) );
  DFFX1_HVT \ram_reg[8][237]  ( .D(n2346), .CLK(clk), .Q(\ram[8][237] ) );
  DFFX1_HVT \ram_reg[8][236]  ( .D(n2345), .CLK(clk), .Q(\ram[8][236] ) );
  DFFX1_HVT \ram_reg[8][235]  ( .D(n2344), .CLK(clk), .Q(\ram[8][235] ) );
  DFFX1_HVT \ram_reg[8][234]  ( .D(n2343), .CLK(clk), .Q(\ram[8][234] ) );
  DFFX1_HVT \ram_reg[8][233]  ( .D(n2342), .CLK(clk), .Q(\ram[8][233] ) );
  DFFX1_HVT \ram_reg[8][232]  ( .D(n2341), .CLK(clk), .Q(\ram[8][232] ) );
  DFFX1_HVT \ram_reg[8][231]  ( .D(n2340), .CLK(clk), .Q(\ram[8][231] ) );
  DFFX1_HVT \ram_reg[8][230]  ( .D(n2339), .CLK(clk), .Q(\ram[8][230] ) );
  DFFX1_HVT \ram_reg[8][229]  ( .D(n2338), .CLK(clk), .Q(\ram[8][229] ) );
  DFFX1_HVT \ram_reg[8][228]  ( .D(n2337), .CLK(clk), .Q(\ram[8][228] ) );
  DFFX1_HVT \ram_reg[8][227]  ( .D(n2336), .CLK(clk), .Q(\ram[8][227] ) );
  DFFX1_HVT \ram_reg[8][226]  ( .D(n2335), .CLK(clk), .Q(\ram[8][226] ) );
  DFFX1_HVT \ram_reg[8][225]  ( .D(n2334), .CLK(clk), .Q(\ram[8][225] ) );
  DFFX1_HVT \ram_reg[8][224]  ( .D(n2333), .CLK(clk), .Q(\ram[8][224] ) );
  DFFX1_HVT \ram_reg[8][223]  ( .D(n2332), .CLK(clk), .Q(\ram[8][223] ) );
  DFFX1_HVT \ram_reg[8][222]  ( .D(n2331), .CLK(clk), .Q(\ram[8][222] ) );
  DFFX1_HVT \ram_reg[8][221]  ( .D(n2330), .CLK(clk), .Q(\ram[8][221] ) );
  DFFX1_HVT \ram_reg[8][220]  ( .D(n2329), .CLK(clk), .Q(\ram[8][220] ) );
  DFFX1_HVT \ram_reg[8][219]  ( .D(n2328), .CLK(clk), .Q(\ram[8][219] ) );
  DFFX1_HVT \ram_reg[8][218]  ( .D(n2327), .CLK(clk), .Q(\ram[8][218] ) );
  DFFX1_HVT \ram_reg[8][217]  ( .D(n2326), .CLK(clk), .Q(\ram[8][217] ) );
  DFFX1_HVT \ram_reg[8][216]  ( .D(n2325), .CLK(clk), .Q(\ram[8][216] ) );
  DFFX1_HVT \ram_reg[8][215]  ( .D(n2324), .CLK(clk), .Q(\ram[8][215] ) );
  DFFX1_HVT \ram_reg[8][214]  ( .D(n2323), .CLK(clk), .Q(\ram[8][214] ) );
  DFFX1_HVT \ram_reg[8][213]  ( .D(n2322), .CLK(clk), .Q(\ram[8][213] ) );
  DFFX1_HVT \ram_reg[8][212]  ( .D(n2321), .CLK(clk), .Q(\ram[8][212] ) );
  DFFX1_HVT \ram_reg[8][211]  ( .D(n2320), .CLK(clk), .Q(\ram[8][211] ) );
  DFFX1_HVT \ram_reg[8][210]  ( .D(n2319), .CLK(clk), .Q(\ram[8][210] ) );
  DFFX1_HVT \ram_reg[8][209]  ( .D(n2318), .CLK(clk), .Q(\ram[8][209] ) );
  DFFX1_HVT \ram_reg[8][208]  ( .D(n2317), .CLK(clk), .Q(\ram[8][208] ) );
  DFFX1_HVT \ram_reg[8][207]  ( .D(n2316), .CLK(clk), .Q(\ram[8][207] ) );
  DFFX1_HVT \ram_reg[8][206]  ( .D(n2315), .CLK(clk), .Q(\ram[8][206] ) );
  DFFX1_HVT \ram_reg[8][205]  ( .D(n2314), .CLK(clk), .Q(\ram[8][205] ) );
  DFFX1_HVT \ram_reg[8][204]  ( .D(n2313), .CLK(clk), .Q(\ram[8][204] ) );
  DFFX1_HVT \ram_reg[8][203]  ( .D(n2312), .CLK(clk), .Q(\ram[8][203] ) );
  DFFX1_HVT \ram_reg[8][202]  ( .D(n2311), .CLK(clk), .Q(\ram[8][202] ) );
  DFFX1_HVT \ram_reg[8][201]  ( .D(n2310), .CLK(clk), .Q(\ram[8][201] ) );
  DFFX1_HVT \ram_reg[8][200]  ( .D(n2309), .CLK(clk), .Q(\ram[8][200] ) );
  DFFX1_HVT \ram_reg[8][199]  ( .D(n2308), .CLK(clk), .Q(\ram[8][199] ) );
  DFFX1_HVT \ram_reg[8][198]  ( .D(n2307), .CLK(clk), .Q(\ram[8][198] ) );
  DFFX1_HVT \ram_reg[8][197]  ( .D(n2306), .CLK(clk), .Q(\ram[8][197] ) );
  DFFX1_HVT \ram_reg[8][196]  ( .D(n2305), .CLK(clk), .Q(\ram[8][196] ) );
  DFFX1_HVT \ram_reg[8][195]  ( .D(n2304), .CLK(clk), .Q(\ram[8][195] ) );
  DFFX1_HVT \ram_reg[8][194]  ( .D(n2303), .CLK(clk), .Q(\ram[8][194] ) );
  DFFX1_HVT \ram_reg[8][193]  ( .D(n2302), .CLK(clk), .Q(\ram[8][193] ) );
  DFFX1_HVT \ram_reg[8][192]  ( .D(n2301), .CLK(clk), .Q(\ram[8][192] ) );
  DFFX1_HVT \ram_reg[8][191]  ( .D(n2300), .CLK(clk), .Q(\ram[8][191] ) );
  DFFX1_HVT \ram_reg[8][190]  ( .D(n2299), .CLK(clk), .Q(\ram[8][190] ) );
  DFFX1_HVT \ram_reg[8][189]  ( .D(n2298), .CLK(clk), .Q(\ram[8][189] ) );
  DFFX1_HVT \ram_reg[8][188]  ( .D(n2297), .CLK(clk), .Q(\ram[8][188] ) );
  DFFX1_HVT \ram_reg[8][187]  ( .D(n2296), .CLK(clk), .Q(\ram[8][187] ) );
  DFFX1_HVT \ram_reg[8][186]  ( .D(n2295), .CLK(clk), .Q(\ram[8][186] ) );
  DFFX1_HVT \ram_reg[8][185]  ( .D(n2294), .CLK(clk), .Q(\ram[8][185] ) );
  DFFX1_HVT \ram_reg[8][184]  ( .D(n2293), .CLK(clk), .Q(\ram[8][184] ) );
  DFFX1_HVT \ram_reg[8][183]  ( .D(n2292), .CLK(clk), .Q(\ram[8][183] ) );
  DFFX1_HVT \ram_reg[8][182]  ( .D(n2291), .CLK(clk), .Q(\ram[8][182] ) );
  DFFX1_HVT \ram_reg[8][181]  ( .D(n2290), .CLK(clk), .Q(\ram[8][181] ) );
  DFFX1_HVT \ram_reg[8][180]  ( .D(n2289), .CLK(clk), .Q(\ram[8][180] ) );
  DFFX1_HVT \ram_reg[8][179]  ( .D(n2288), .CLK(clk), .Q(\ram[8][179] ) );
  DFFX1_HVT \ram_reg[8][178]  ( .D(n2287), .CLK(clk), .Q(\ram[8][178] ) );
  DFFX1_HVT \ram_reg[8][177]  ( .D(n2286), .CLK(clk), .Q(\ram[8][177] ) );
  DFFX1_HVT \ram_reg[8][176]  ( .D(n2285), .CLK(clk), .Q(\ram[8][176] ) );
  DFFX1_HVT \ram_reg[8][175]  ( .D(n2284), .CLK(clk), .Q(\ram[8][175] ) );
  DFFX1_HVT \ram_reg[8][174]  ( .D(n2283), .CLK(clk), .Q(\ram[8][174] ) );
  DFFX1_HVT \ram_reg[8][173]  ( .D(n2282), .CLK(clk), .Q(\ram[8][173] ) );
  DFFX1_HVT \ram_reg[8][172]  ( .D(n2281), .CLK(clk), .Q(\ram[8][172] ) );
  DFFX1_HVT \ram_reg[8][171]  ( .D(n2280), .CLK(clk), .Q(\ram[8][171] ) );
  DFFX1_HVT \ram_reg[8][170]  ( .D(n2279), .CLK(clk), .Q(\ram[8][170] ) );
  DFFX1_HVT \ram_reg[8][169]  ( .D(n2278), .CLK(clk), .Q(\ram[8][169] ) );
  DFFX1_HVT \ram_reg[8][168]  ( .D(n2277), .CLK(clk), .Q(\ram[8][168] ) );
  DFFX1_HVT \ram_reg[8][167]  ( .D(n2276), .CLK(clk), .Q(\ram[8][167] ) );
  DFFX1_HVT \ram_reg[8][166]  ( .D(n2275), .CLK(clk), .Q(\ram[8][166] ) );
  DFFX1_HVT \ram_reg[8][165]  ( .D(n2274), .CLK(clk), .Q(\ram[8][165] ) );
  DFFX1_HVT \ram_reg[8][164]  ( .D(n2273), .CLK(clk), .Q(\ram[8][164] ) );
  DFFX1_HVT \ram_reg[8][163]  ( .D(n2272), .CLK(clk), .Q(\ram[8][163] ) );
  DFFX1_HVT \ram_reg[8][162]  ( .D(n2271), .CLK(clk), .Q(\ram[8][162] ) );
  DFFX1_HVT \ram_reg[8][161]  ( .D(n2270), .CLK(clk), .Q(\ram[8][161] ) );
  DFFX1_HVT \ram_reg[8][160]  ( .D(n2269), .CLK(clk), .Q(\ram[8][160] ) );
  DFFX1_HVT \ram_reg[8][159]  ( .D(n2268), .CLK(clk), .Q(\ram[8][159] ) );
  DFFX1_HVT \ram_reg[8][158]  ( .D(n2267), .CLK(clk), .Q(\ram[8][158] ) );
  DFFX1_HVT \ram_reg[8][157]  ( .D(n2266), .CLK(clk), .Q(\ram[8][157] ) );
  DFFX1_HVT \ram_reg[8][156]  ( .D(n2265), .CLK(clk), .Q(\ram[8][156] ) );
  DFFX1_HVT \ram_reg[8][155]  ( .D(n2264), .CLK(clk), .Q(\ram[8][155] ) );
  DFFX1_HVT \ram_reg[8][154]  ( .D(n2263), .CLK(clk), .Q(\ram[8][154] ) );
  DFFX1_HVT \ram_reg[8][153]  ( .D(n2262), .CLK(clk), .Q(\ram[8][153] ) );
  DFFX1_HVT \ram_reg[8][152]  ( .D(n2261), .CLK(clk), .Q(\ram[8][152] ) );
  DFFX1_HVT \ram_reg[8][151]  ( .D(n2260), .CLK(clk), .Q(\ram[8][151] ) );
  DFFX1_HVT \ram_reg[8][150]  ( .D(n2259), .CLK(clk), .Q(\ram[8][150] ) );
  DFFX1_HVT \ram_reg[8][149]  ( .D(n2258), .CLK(clk), .Q(\ram[8][149] ) );
  DFFX1_HVT \ram_reg[8][148]  ( .D(n2257), .CLK(clk), .Q(\ram[8][148] ) );
  DFFX1_HVT \ram_reg[8][147]  ( .D(n2256), .CLK(clk), .Q(\ram[8][147] ) );
  DFFX1_HVT \ram_reg[8][146]  ( .D(n2255), .CLK(clk), .Q(\ram[8][146] ) );
  DFFX1_HVT \ram_reg[8][145]  ( .D(n2254), .CLK(clk), .Q(\ram[8][145] ) );
  DFFX1_HVT \ram_reg[8][144]  ( .D(n2253), .CLK(clk), .Q(\ram[8][144] ) );
  DFFX1_HVT \ram_reg[8][143]  ( .D(n2252), .CLK(clk), .Q(\ram[8][143] ) );
  DFFX1_HVT \ram_reg[8][142]  ( .D(n2251), .CLK(clk), .Q(\ram[8][142] ) );
  DFFX1_HVT \ram_reg[8][141]  ( .D(n2250), .CLK(clk), .Q(\ram[8][141] ) );
  DFFX1_HVT \ram_reg[8][140]  ( .D(n2249), .CLK(clk), .Q(\ram[8][140] ) );
  DFFX1_HVT \ram_reg[8][139]  ( .D(n2248), .CLK(clk), .Q(\ram[8][139] ) );
  DFFX1_HVT \ram_reg[8][138]  ( .D(n2247), .CLK(clk), .Q(\ram[8][138] ) );
  DFFX1_HVT \ram_reg[8][137]  ( .D(n2246), .CLK(clk), .Q(\ram[8][137] ) );
  DFFX1_HVT \ram_reg[8][136]  ( .D(n2245), .CLK(clk), .Q(\ram[8][136] ) );
  DFFX1_HVT \ram_reg[8][135]  ( .D(n2244), .CLK(clk), .Q(\ram[8][135] ) );
  DFFX1_HVT \ram_reg[8][134]  ( .D(n2243), .CLK(clk), .Q(\ram[8][134] ) );
  DFFX1_HVT \ram_reg[8][133]  ( .D(n2242), .CLK(clk), .Q(\ram[8][133] ) );
  DFFX1_HVT \ram_reg[8][132]  ( .D(n2241), .CLK(clk), .Q(\ram[8][132] ) );
  DFFX1_HVT \ram_reg[8][131]  ( .D(n2240), .CLK(clk), .Q(\ram[8][131] ) );
  DFFX1_HVT \ram_reg[8][130]  ( .D(n2239), .CLK(clk), .Q(\ram[8][130] ) );
  DFFX1_HVT \ram_reg[8][129]  ( .D(n2238), .CLK(clk), .Q(\ram[8][129] ) );
  DFFX1_HVT \ram_reg[8][128]  ( .D(n2237), .CLK(clk), .Q(\ram[8][128] ) );
  DFFX1_HVT \ram_reg[8][127]  ( .D(n2236), .CLK(clk), .Q(\ram[8][127] ) );
  DFFX1_HVT \ram_reg[8][126]  ( .D(n2235), .CLK(clk), .Q(\ram[8][126] ) );
  DFFX1_HVT \ram_reg[8][125]  ( .D(n2234), .CLK(clk), .Q(\ram[8][125] ) );
  DFFX1_HVT \ram_reg[8][124]  ( .D(n2233), .CLK(clk), .Q(\ram[8][124] ) );
  DFFX1_HVT \ram_reg[8][123]  ( .D(n2232), .CLK(clk), .Q(\ram[8][123] ) );
  DFFX1_HVT \ram_reg[8][122]  ( .D(n2231), .CLK(clk), .Q(\ram[8][122] ) );
  DFFX1_HVT \ram_reg[8][121]  ( .D(n2230), .CLK(clk), .Q(\ram[8][121] ) );
  DFFX1_HVT \ram_reg[8][120]  ( .D(n2229), .CLK(clk), .Q(\ram[8][120] ) );
  DFFX1_HVT \ram_reg[8][119]  ( .D(n2228), .CLK(clk), .Q(\ram[8][119] ) );
  DFFX1_HVT \ram_reg[8][118]  ( .D(n2227), .CLK(clk), .Q(\ram[8][118] ) );
  DFFX1_HVT \ram_reg[8][117]  ( .D(n2226), .CLK(clk), .Q(\ram[8][117] ) );
  DFFX1_HVT \ram_reg[8][116]  ( .D(n2225), .CLK(clk), .Q(\ram[8][116] ) );
  DFFX1_HVT \ram_reg[8][115]  ( .D(n2224), .CLK(clk), .Q(\ram[8][115] ) );
  DFFX1_HVT \ram_reg[8][114]  ( .D(n2223), .CLK(clk), .Q(\ram[8][114] ) );
  DFFX1_HVT \ram_reg[8][113]  ( .D(n2222), .CLK(clk), .Q(\ram[8][113] ) );
  DFFX1_HVT \ram_reg[8][112]  ( .D(n2221), .CLK(clk), .Q(\ram[8][112] ) );
  DFFX1_HVT \ram_reg[8][111]  ( .D(n2220), .CLK(clk), .Q(\ram[8][111] ) );
  DFFX1_HVT \ram_reg[8][110]  ( .D(n2219), .CLK(clk), .Q(\ram[8][110] ) );
  DFFX1_HVT \ram_reg[8][109]  ( .D(n2218), .CLK(clk), .Q(\ram[8][109] ) );
  DFFX1_HVT \ram_reg[8][108]  ( .D(n2217), .CLK(clk), .Q(\ram[8][108] ) );
  DFFX1_HVT \ram_reg[8][107]  ( .D(n2216), .CLK(clk), .Q(\ram[8][107] ) );
  DFFX1_HVT \ram_reg[8][106]  ( .D(n2215), .CLK(clk), .Q(\ram[8][106] ) );
  DFFX1_HVT \ram_reg[8][105]  ( .D(n2214), .CLK(clk), .Q(\ram[8][105] ) );
  DFFX1_HVT \ram_reg[8][104]  ( .D(n2213), .CLK(clk), .Q(\ram[8][104] ) );
  DFFX1_HVT \ram_reg[8][103]  ( .D(n2212), .CLK(clk), .Q(\ram[8][103] ) );
  DFFX1_HVT \ram_reg[8][102]  ( .D(n2211), .CLK(clk), .Q(\ram[8][102] ) );
  DFFX1_HVT \ram_reg[8][101]  ( .D(n2210), .CLK(clk), .Q(\ram[8][101] ) );
  DFFX1_HVT \ram_reg[8][100]  ( .D(n2209), .CLK(clk), .Q(\ram[8][100] ) );
  DFFX1_HVT \ram_reg[8][99]  ( .D(n2208), .CLK(clk), .Q(\ram[8][99] ) );
  DFFX1_HVT \ram_reg[8][98]  ( .D(n2207), .CLK(clk), .Q(\ram[8][98] ) );
  DFFX1_HVT \ram_reg[8][97]  ( .D(n2206), .CLK(clk), .Q(\ram[8][97] ) );
  DFFX1_HVT \ram_reg[8][96]  ( .D(n2205), .CLK(clk), .Q(\ram[8][96] ) );
  DFFX1_HVT \ram_reg[8][95]  ( .D(n2204), .CLK(clk), .Q(\ram[8][95] ) );
  DFFX1_HVT \ram_reg[8][94]  ( .D(n2203), .CLK(clk), .Q(\ram[8][94] ) );
  DFFX1_HVT \ram_reg[8][93]  ( .D(n2202), .CLK(clk), .Q(\ram[8][93] ) );
  DFFX1_HVT \ram_reg[8][92]  ( .D(n2201), .CLK(clk), .Q(\ram[8][92] ) );
  DFFX1_HVT \ram_reg[8][91]  ( .D(n2200), .CLK(clk), .Q(\ram[8][91] ) );
  DFFX1_HVT \ram_reg[8][90]  ( .D(n2199), .CLK(clk), .Q(\ram[8][90] ) );
  DFFX1_HVT \ram_reg[8][89]  ( .D(n2198), .CLK(clk), .Q(\ram[8][89] ) );
  DFFX1_HVT \ram_reg[8][88]  ( .D(n2197), .CLK(clk), .Q(\ram[8][88] ) );
  DFFX1_HVT \ram_reg[8][87]  ( .D(n2196), .CLK(clk), .Q(\ram[8][87] ) );
  DFFX1_HVT \ram_reg[8][86]  ( .D(n2195), .CLK(clk), .Q(\ram[8][86] ) );
  DFFX1_HVT \ram_reg[8][85]  ( .D(n2194), .CLK(clk), .Q(\ram[8][85] ) );
  DFFX1_HVT \ram_reg[8][84]  ( .D(n2193), .CLK(clk), .Q(\ram[8][84] ) );
  DFFX1_HVT \ram_reg[8][83]  ( .D(n2192), .CLK(clk), .Q(\ram[8][83] ) );
  DFFX1_HVT \ram_reg[8][82]  ( .D(n2191), .CLK(clk), .Q(\ram[8][82] ) );
  DFFX1_HVT \ram_reg[8][81]  ( .D(n2190), .CLK(clk), .Q(\ram[8][81] ) );
  DFFX1_HVT \ram_reg[8][80]  ( .D(n2189), .CLK(clk), .Q(\ram[8][80] ) );
  DFFX1_HVT \ram_reg[8][79]  ( .D(n2188), .CLK(clk), .Q(\ram[8][79] ) );
  DFFX1_HVT \ram_reg[8][78]  ( .D(n2187), .CLK(clk), .Q(\ram[8][78] ) );
  DFFX1_HVT \ram_reg[8][77]  ( .D(n2186), .CLK(clk), .Q(\ram[8][77] ) );
  DFFX1_HVT \ram_reg[8][76]  ( .D(n2185), .CLK(clk), .Q(\ram[8][76] ) );
  DFFX1_HVT \ram_reg[8][75]  ( .D(n2184), .CLK(clk), .Q(\ram[8][75] ) );
  DFFX1_HVT \ram_reg[8][74]  ( .D(n2183), .CLK(clk), .Q(\ram[8][74] ) );
  DFFX1_HVT \ram_reg[8][73]  ( .D(n2182), .CLK(clk), .Q(\ram[8][73] ) );
  DFFX1_HVT \ram_reg[8][72]  ( .D(n2181), .CLK(clk), .Q(\ram[8][72] ) );
  DFFX1_HVT \ram_reg[8][71]  ( .D(n2180), .CLK(clk), .Q(\ram[8][71] ) );
  DFFX1_HVT \ram_reg[8][70]  ( .D(n2179), .CLK(clk), .Q(\ram[8][70] ) );
  DFFX1_HVT \ram_reg[8][69]  ( .D(n2178), .CLK(clk), .Q(\ram[8][69] ) );
  DFFX1_HVT \ram_reg[8][68]  ( .D(n2177), .CLK(clk), .Q(\ram[8][68] ) );
  DFFX1_HVT \ram_reg[8][67]  ( .D(n2176), .CLK(clk), .Q(\ram[8][67] ) );
  DFFX1_HVT \ram_reg[8][66]  ( .D(n2175), .CLK(clk), .Q(\ram[8][66] ) );
  DFFX1_HVT \ram_reg[8][65]  ( .D(n2174), .CLK(clk), .Q(\ram[8][65] ) );
  DFFX1_HVT \ram_reg[8][64]  ( .D(n2173), .CLK(clk), .Q(\ram[8][64] ) );
  DFFX1_HVT \ram_reg[8][63]  ( .D(n2172), .CLK(clk), .Q(\ram[8][63] ) );
  DFFX1_HVT \ram_reg[8][62]  ( .D(n2171), .CLK(clk), .Q(\ram[8][62] ) );
  DFFX1_HVT \ram_reg[8][61]  ( .D(n2170), .CLK(clk), .Q(\ram[8][61] ) );
  DFFX1_HVT \ram_reg[8][60]  ( .D(n2169), .CLK(clk), .Q(\ram[8][60] ) );
  DFFX1_HVT \ram_reg[8][59]  ( .D(n2168), .CLK(clk), .Q(\ram[8][59] ) );
  DFFX1_HVT \ram_reg[8][58]  ( .D(n2167), .CLK(clk), .Q(\ram[8][58] ) );
  DFFX1_HVT \ram_reg[8][57]  ( .D(n2166), .CLK(clk), .Q(\ram[8][57] ) );
  DFFX1_HVT \ram_reg[8][56]  ( .D(n2165), .CLK(clk), .Q(\ram[8][56] ) );
  DFFX1_HVT \ram_reg[8][55]  ( .D(n2164), .CLK(clk), .Q(\ram[8][55] ) );
  DFFX1_HVT \ram_reg[8][54]  ( .D(n2163), .CLK(clk), .Q(\ram[8][54] ) );
  DFFX1_HVT \ram_reg[8][53]  ( .D(n2162), .CLK(clk), .Q(\ram[8][53] ) );
  DFFX1_HVT \ram_reg[8][52]  ( .D(n2161), .CLK(clk), .Q(\ram[8][52] ) );
  DFFX1_HVT \ram_reg[8][51]  ( .D(n2160), .CLK(clk), .Q(\ram[8][51] ) );
  DFFX1_HVT \ram_reg[8][50]  ( .D(n2159), .CLK(clk), .Q(\ram[8][50] ) );
  DFFX1_HVT \ram_reg[8][49]  ( .D(n2158), .CLK(clk), .Q(\ram[8][49] ) );
  DFFX1_HVT \ram_reg[8][48]  ( .D(n2157), .CLK(clk), .Q(\ram[8][48] ) );
  DFFX1_HVT \ram_reg[8][47]  ( .D(n2156), .CLK(clk), .Q(\ram[8][47] ) );
  DFFX1_HVT \ram_reg[8][46]  ( .D(n2155), .CLK(clk), .Q(\ram[8][46] ) );
  DFFX1_HVT \ram_reg[8][45]  ( .D(n2154), .CLK(clk), .Q(\ram[8][45] ) );
  DFFX1_HVT \ram_reg[8][44]  ( .D(n2153), .CLK(clk), .Q(\ram[8][44] ) );
  DFFX1_HVT \ram_reg[8][43]  ( .D(n2152), .CLK(clk), .Q(\ram[8][43] ) );
  DFFX1_HVT \ram_reg[8][42]  ( .D(n2151), .CLK(clk), .Q(\ram[8][42] ) );
  DFFX1_HVT \ram_reg[8][41]  ( .D(n2150), .CLK(clk), .Q(\ram[8][41] ) );
  DFFX1_HVT \ram_reg[8][40]  ( .D(n2149), .CLK(clk), .Q(\ram[8][40] ) );
  DFFX1_HVT \ram_reg[8][39]  ( .D(n2148), .CLK(clk), .Q(\ram[8][39] ) );
  DFFX1_HVT \ram_reg[8][38]  ( .D(n2147), .CLK(clk), .Q(\ram[8][38] ) );
  DFFX1_HVT \ram_reg[8][37]  ( .D(n2146), .CLK(clk), .Q(\ram[8][37] ) );
  DFFX1_HVT \ram_reg[8][36]  ( .D(n2145), .CLK(clk), .Q(\ram[8][36] ) );
  DFFX1_HVT \ram_reg[8][35]  ( .D(n2144), .CLK(clk), .Q(\ram[8][35] ) );
  DFFX1_HVT \ram_reg[8][34]  ( .D(n2143), .CLK(clk), .Q(\ram[8][34] ) );
  DFFX1_HVT \ram_reg[8][33]  ( .D(n2142), .CLK(clk), .Q(\ram[8][33] ) );
  DFFX1_HVT \ram_reg[8][32]  ( .D(n2141), .CLK(clk), .Q(\ram[8][32] ) );
  DFFX1_HVT \ram_reg[8][31]  ( .D(n2140), .CLK(clk), .Q(\ram[8][31] ) );
  DFFX1_HVT \ram_reg[8][30]  ( .D(n2139), .CLK(clk), .Q(\ram[8][30] ) );
  DFFX1_HVT \ram_reg[8][29]  ( .D(n2138), .CLK(clk), .Q(\ram[8][29] ) );
  DFFX1_HVT \ram_reg[8][28]  ( .D(n2137), .CLK(clk), .Q(\ram[8][28] ) );
  DFFX1_HVT \ram_reg[8][27]  ( .D(n2136), .CLK(clk), .Q(\ram[8][27] ) );
  DFFX1_HVT \ram_reg[8][26]  ( .D(n2135), .CLK(clk), .Q(\ram[8][26] ) );
  DFFX1_HVT \ram_reg[8][25]  ( .D(n2134), .CLK(clk), .Q(\ram[8][25] ) );
  DFFX1_HVT \ram_reg[8][24]  ( .D(n2133), .CLK(clk), .Q(\ram[8][24] ) );
  DFFX1_HVT \ram_reg[8][23]  ( .D(n2132), .CLK(clk), .Q(\ram[8][23] ) );
  DFFX1_HVT \ram_reg[8][22]  ( .D(n2131), .CLK(clk), .Q(\ram[8][22] ) );
  DFFX1_HVT \ram_reg[8][21]  ( .D(n2130), .CLK(clk), .Q(\ram[8][21] ) );
  DFFX1_HVT \ram_reg[8][20]  ( .D(n2129), .CLK(clk), .Q(\ram[8][20] ) );
  DFFX1_HVT \ram_reg[8][19]  ( .D(n2128), .CLK(clk), .Q(\ram[8][19] ) );
  DFFX1_HVT \ram_reg[8][18]  ( .D(n2127), .CLK(clk), .Q(\ram[8][18] ) );
  DFFX1_HVT \ram_reg[8][17]  ( .D(n2126), .CLK(clk), .Q(\ram[8][17] ) );
  DFFX1_HVT \ram_reg[8][16]  ( .D(n2125), .CLK(clk), .Q(\ram[8][16] ) );
  DFFX1_HVT \ram_reg[8][15]  ( .D(n2124), .CLK(clk), .Q(\ram[8][15] ) );
  DFFX1_HVT \ram_reg[8][14]  ( .D(n2123), .CLK(clk), .Q(\ram[8][14] ) );
  DFFX1_HVT \ram_reg[8][13]  ( .D(n2122), .CLK(clk), .Q(\ram[8][13] ) );
  DFFX1_HVT \ram_reg[8][12]  ( .D(n2121), .CLK(clk), .Q(\ram[8][12] ) );
  DFFX1_HVT \ram_reg[8][11]  ( .D(n2120), .CLK(clk), .Q(\ram[8][11] ) );
  DFFX1_HVT \ram_reg[8][10]  ( .D(n2119), .CLK(clk), .Q(\ram[8][10] ) );
  DFFX1_HVT \ram_reg[8][9]  ( .D(n2118), .CLK(clk), .Q(\ram[8][9] ) );
  DFFX1_HVT \ram_reg[8][8]  ( .D(n2117), .CLK(clk), .Q(\ram[8][8] ) );
  DFFX1_HVT \ram_reg[8][7]  ( .D(n2116), .CLK(clk), .Q(\ram[8][7] ) );
  DFFX1_HVT \ram_reg[8][6]  ( .D(n2115), .CLK(clk), .Q(\ram[8][6] ) );
  DFFX1_HVT \ram_reg[8][5]  ( .D(n2114), .CLK(clk), .Q(\ram[8][5] ) );
  DFFX1_HVT \ram_reg[8][4]  ( .D(n2113), .CLK(clk), .Q(\ram[8][4] ) );
  DFFX1_HVT \ram_reg[8][3]  ( .D(n2112), .CLK(clk), .Q(\ram[8][3] ) );
  DFFX1_HVT \ram_reg[8][2]  ( .D(n2111), .CLK(clk), .Q(\ram[8][2] ) );
  DFFX1_HVT \ram_reg[8][1]  ( .D(n2110), .CLK(clk), .Q(\ram[8][1] ) );
  DFFX1_HVT \ram_reg[8][0]  ( .D(n2109), .CLK(clk), .Q(\ram[8][0] ) );
  DFFX1_HVT \ram_reg[7][255]  ( .D(n2108), .CLK(clk), .Q(\ram[7][255] ) );
  DFFX1_HVT \ram_reg[7][254]  ( .D(n2107), .CLK(clk), .Q(\ram[7][254] ) );
  DFFX1_HVT \ram_reg[7][253]  ( .D(n2106), .CLK(clk), .Q(\ram[7][253] ) );
  DFFX1_HVT \ram_reg[7][252]  ( .D(n2105), .CLK(clk), .Q(\ram[7][252] ) );
  DFFX1_HVT \ram_reg[7][251]  ( .D(n2104), .CLK(clk), .Q(\ram[7][251] ) );
  DFFX1_HVT \ram_reg[7][250]  ( .D(n2103), .CLK(clk), .Q(\ram[7][250] ) );
  DFFX1_HVT \ram_reg[7][249]  ( .D(n2102), .CLK(clk), .Q(\ram[7][249] ) );
  DFFX1_HVT \ram_reg[7][248]  ( .D(n2101), .CLK(clk), .Q(\ram[7][248] ) );
  DFFX1_HVT \ram_reg[7][247]  ( .D(n2100), .CLK(clk), .Q(\ram[7][247] ) );
  DFFX1_HVT \ram_reg[7][246]  ( .D(n2099), .CLK(clk), .Q(\ram[7][246] ) );
  DFFX1_HVT \ram_reg[7][245]  ( .D(n2098), .CLK(clk), .Q(\ram[7][245] ) );
  DFFX1_HVT \ram_reg[7][244]  ( .D(n2097), .CLK(clk), .Q(\ram[7][244] ) );
  DFFX1_HVT \ram_reg[7][243]  ( .D(n2096), .CLK(clk), .Q(\ram[7][243] ) );
  DFFX1_HVT \ram_reg[7][242]  ( .D(n2095), .CLK(clk), .Q(\ram[7][242] ) );
  DFFX1_HVT \ram_reg[7][241]  ( .D(n2094), .CLK(clk), .Q(\ram[7][241] ) );
  DFFX1_HVT \ram_reg[7][240]  ( .D(n2093), .CLK(clk), .Q(\ram[7][240] ) );
  DFFX1_HVT \ram_reg[7][239]  ( .D(n2092), .CLK(clk), .Q(\ram[7][239] ) );
  DFFX1_HVT \ram_reg[7][238]  ( .D(n2091), .CLK(clk), .Q(\ram[7][238] ) );
  DFFX1_HVT \ram_reg[7][237]  ( .D(n2090), .CLK(clk), .Q(\ram[7][237] ) );
  DFFX1_HVT \ram_reg[7][236]  ( .D(n2089), .CLK(clk), .Q(\ram[7][236] ) );
  DFFX1_HVT \ram_reg[7][235]  ( .D(n2088), .CLK(clk), .Q(\ram[7][235] ) );
  DFFX1_HVT \ram_reg[7][234]  ( .D(n2087), .CLK(clk), .Q(\ram[7][234] ) );
  DFFX1_HVT \ram_reg[7][233]  ( .D(n2086), .CLK(clk), .Q(\ram[7][233] ) );
  DFFX1_HVT \ram_reg[7][232]  ( .D(n2085), .CLK(clk), .Q(\ram[7][232] ) );
  DFFX1_HVT \ram_reg[7][231]  ( .D(n2084), .CLK(clk), .Q(\ram[7][231] ) );
  DFFX1_HVT \ram_reg[7][230]  ( .D(n2083), .CLK(clk), .Q(\ram[7][230] ) );
  DFFX1_HVT \ram_reg[7][229]  ( .D(n2082), .CLK(clk), .Q(\ram[7][229] ) );
  DFFX1_HVT \ram_reg[7][228]  ( .D(n2081), .CLK(clk), .Q(\ram[7][228] ) );
  DFFX1_HVT \ram_reg[7][227]  ( .D(n2080), .CLK(clk), .Q(\ram[7][227] ) );
  DFFX1_HVT \ram_reg[7][226]  ( .D(n2079), .CLK(clk), .Q(\ram[7][226] ) );
  DFFX1_HVT \ram_reg[7][225]  ( .D(n2078), .CLK(clk), .Q(\ram[7][225] ) );
  DFFX1_HVT \ram_reg[7][224]  ( .D(n2077), .CLK(clk), .Q(\ram[7][224] ) );
  DFFX1_HVT \ram_reg[7][223]  ( .D(n2076), .CLK(clk), .Q(\ram[7][223] ) );
  DFFX1_HVT \ram_reg[7][222]  ( .D(n2075), .CLK(clk), .Q(\ram[7][222] ) );
  DFFX1_HVT \ram_reg[7][221]  ( .D(n2074), .CLK(clk), .Q(\ram[7][221] ) );
  DFFX1_HVT \ram_reg[7][220]  ( .D(n2073), .CLK(clk), .Q(\ram[7][220] ) );
  DFFX1_HVT \ram_reg[7][219]  ( .D(n2072), .CLK(clk), .Q(\ram[7][219] ) );
  DFFX1_HVT \ram_reg[7][218]  ( .D(n2071), .CLK(clk), .Q(\ram[7][218] ) );
  DFFX1_HVT \ram_reg[7][217]  ( .D(n2070), .CLK(clk), .Q(\ram[7][217] ) );
  DFFX1_HVT \ram_reg[7][216]  ( .D(n2069), .CLK(clk), .Q(\ram[7][216] ) );
  DFFX1_HVT \ram_reg[7][215]  ( .D(n2068), .CLK(clk), .Q(\ram[7][215] ) );
  DFFX1_HVT \ram_reg[7][214]  ( .D(n2067), .CLK(clk), .Q(\ram[7][214] ) );
  DFFX1_HVT \ram_reg[7][213]  ( .D(n2066), .CLK(clk), .Q(\ram[7][213] ) );
  DFFX1_HVT \ram_reg[7][212]  ( .D(n2065), .CLK(clk), .Q(\ram[7][212] ) );
  DFFX1_HVT \ram_reg[7][211]  ( .D(n2064), .CLK(clk), .Q(\ram[7][211] ) );
  DFFX1_HVT \ram_reg[7][210]  ( .D(n2063), .CLK(clk), .Q(\ram[7][210] ) );
  DFFX1_HVT \ram_reg[7][209]  ( .D(n2062), .CLK(clk), .Q(\ram[7][209] ) );
  DFFX1_HVT \ram_reg[7][208]  ( .D(n2061), .CLK(clk), .Q(\ram[7][208] ) );
  DFFX1_HVT \ram_reg[7][207]  ( .D(n2060), .CLK(clk), .Q(\ram[7][207] ) );
  DFFX1_HVT \ram_reg[7][206]  ( .D(n2059), .CLK(clk), .Q(\ram[7][206] ) );
  DFFX1_HVT \ram_reg[7][205]  ( .D(n2058), .CLK(clk), .Q(\ram[7][205] ) );
  DFFX1_HVT \ram_reg[7][204]  ( .D(n2057), .CLK(clk), .Q(\ram[7][204] ) );
  DFFX1_HVT \ram_reg[7][203]  ( .D(n2056), .CLK(clk), .Q(\ram[7][203] ) );
  DFFX1_HVT \ram_reg[7][202]  ( .D(n2055), .CLK(clk), .Q(\ram[7][202] ) );
  DFFX1_HVT \ram_reg[7][201]  ( .D(n2054), .CLK(clk), .Q(\ram[7][201] ) );
  DFFX1_HVT \ram_reg[7][200]  ( .D(n2053), .CLK(clk), .Q(\ram[7][200] ) );
  DFFX1_HVT \ram_reg[7][199]  ( .D(n2052), .CLK(clk), .Q(\ram[7][199] ) );
  DFFX1_HVT \ram_reg[7][198]  ( .D(n2051), .CLK(clk), .Q(\ram[7][198] ) );
  DFFX1_HVT \ram_reg[7][197]  ( .D(n2050), .CLK(clk), .Q(\ram[7][197] ) );
  DFFX1_HVT \ram_reg[7][196]  ( .D(n2049), .CLK(clk), .Q(\ram[7][196] ) );
  DFFX1_HVT \ram_reg[7][195]  ( .D(n2048), .CLK(clk), .Q(\ram[7][195] ) );
  DFFX1_HVT \ram_reg[7][194]  ( .D(n2047), .CLK(clk), .Q(\ram[7][194] ) );
  DFFX1_HVT \ram_reg[7][193]  ( .D(n2046), .CLK(clk), .Q(\ram[7][193] ) );
  DFFX1_HVT \ram_reg[7][192]  ( .D(n2045), .CLK(clk), .Q(\ram[7][192] ) );
  DFFX1_HVT \ram_reg[7][191]  ( .D(n2044), .CLK(clk), .Q(\ram[7][191] ) );
  DFFX1_HVT \ram_reg[7][190]  ( .D(n2043), .CLK(clk), .Q(\ram[7][190] ) );
  DFFX1_HVT \ram_reg[7][189]  ( .D(n2042), .CLK(clk), .Q(\ram[7][189] ) );
  DFFX1_HVT \ram_reg[7][188]  ( .D(n2041), .CLK(clk), .Q(\ram[7][188] ) );
  DFFX1_HVT \ram_reg[7][187]  ( .D(n2040), .CLK(clk), .Q(\ram[7][187] ) );
  DFFX1_HVT \ram_reg[7][186]  ( .D(n2039), .CLK(clk), .Q(\ram[7][186] ) );
  DFFX1_HVT \ram_reg[7][185]  ( .D(n2038), .CLK(clk), .Q(\ram[7][185] ) );
  DFFX1_HVT \ram_reg[7][184]  ( .D(n2037), .CLK(clk), .Q(\ram[7][184] ) );
  DFFX1_HVT \ram_reg[7][183]  ( .D(n2036), .CLK(clk), .Q(\ram[7][183] ) );
  DFFX1_HVT \ram_reg[7][182]  ( .D(n2035), .CLK(clk), .Q(\ram[7][182] ) );
  DFFX1_HVT \ram_reg[7][181]  ( .D(n2034), .CLK(clk), .Q(\ram[7][181] ) );
  DFFX1_HVT \ram_reg[7][180]  ( .D(n2033), .CLK(clk), .Q(\ram[7][180] ) );
  DFFX1_HVT \ram_reg[7][179]  ( .D(n2032), .CLK(clk), .Q(\ram[7][179] ) );
  DFFX1_HVT \ram_reg[7][178]  ( .D(n2031), .CLK(clk), .Q(\ram[7][178] ) );
  DFFX1_HVT \ram_reg[7][177]  ( .D(n2030), .CLK(clk), .Q(\ram[7][177] ) );
  DFFX1_HVT \ram_reg[7][176]  ( .D(n2029), .CLK(clk), .Q(\ram[7][176] ) );
  DFFX1_HVT \ram_reg[7][175]  ( .D(n2028), .CLK(clk), .Q(\ram[7][175] ) );
  DFFX1_HVT \ram_reg[7][174]  ( .D(n2027), .CLK(clk), .Q(\ram[7][174] ) );
  DFFX1_HVT \ram_reg[7][173]  ( .D(n2026), .CLK(clk), .Q(\ram[7][173] ) );
  DFFX1_HVT \ram_reg[7][172]  ( .D(n2025), .CLK(clk), .Q(\ram[7][172] ) );
  DFFX1_HVT \ram_reg[7][171]  ( .D(n2024), .CLK(clk), .Q(\ram[7][171] ) );
  DFFX1_HVT \ram_reg[7][170]  ( .D(n2023), .CLK(clk), .Q(\ram[7][170] ) );
  DFFX1_HVT \ram_reg[7][169]  ( .D(n2022), .CLK(clk), .Q(\ram[7][169] ) );
  DFFX1_HVT \ram_reg[7][168]  ( .D(n2021), .CLK(clk), .Q(\ram[7][168] ) );
  DFFX1_HVT \ram_reg[7][167]  ( .D(n2020), .CLK(clk), .Q(\ram[7][167] ) );
  DFFX1_HVT \ram_reg[7][166]  ( .D(n2019), .CLK(clk), .Q(\ram[7][166] ) );
  DFFX1_HVT \ram_reg[7][165]  ( .D(n2018), .CLK(clk), .Q(\ram[7][165] ) );
  DFFX1_HVT \ram_reg[7][164]  ( .D(n2017), .CLK(clk), .Q(\ram[7][164] ) );
  DFFX1_HVT \ram_reg[7][163]  ( .D(n2016), .CLK(clk), .Q(\ram[7][163] ) );
  DFFX1_HVT \ram_reg[7][162]  ( .D(n2015), .CLK(clk), .Q(\ram[7][162] ) );
  DFFX1_HVT \ram_reg[7][161]  ( .D(n2014), .CLK(clk), .Q(\ram[7][161] ) );
  DFFX1_HVT \ram_reg[7][160]  ( .D(n2013), .CLK(clk), .Q(\ram[7][160] ) );
  DFFX1_HVT \ram_reg[7][159]  ( .D(n2012), .CLK(clk), .Q(\ram[7][159] ) );
  DFFX1_HVT \ram_reg[7][158]  ( .D(n2011), .CLK(clk), .Q(\ram[7][158] ) );
  DFFX1_HVT \ram_reg[7][157]  ( .D(n2010), .CLK(clk), .Q(\ram[7][157] ) );
  DFFX1_HVT \ram_reg[7][156]  ( .D(n2009), .CLK(clk), .Q(\ram[7][156] ) );
  DFFX1_HVT \ram_reg[7][155]  ( .D(n2008), .CLK(clk), .Q(\ram[7][155] ) );
  DFFX1_HVT \ram_reg[7][154]  ( .D(n2007), .CLK(clk), .Q(\ram[7][154] ) );
  DFFX1_HVT \ram_reg[7][153]  ( .D(n2006), .CLK(clk), .Q(\ram[7][153] ) );
  DFFX1_HVT \ram_reg[7][152]  ( .D(n2005), .CLK(clk), .Q(\ram[7][152] ) );
  DFFX1_HVT \ram_reg[7][151]  ( .D(n2004), .CLK(clk), .Q(\ram[7][151] ) );
  DFFX1_HVT \ram_reg[7][150]  ( .D(n2003), .CLK(clk), .Q(\ram[7][150] ) );
  DFFX1_HVT \ram_reg[7][149]  ( .D(n2002), .CLK(clk), .Q(\ram[7][149] ) );
  DFFX1_HVT \ram_reg[7][148]  ( .D(n2001), .CLK(clk), .Q(\ram[7][148] ) );
  DFFX1_HVT \ram_reg[7][147]  ( .D(n2000), .CLK(clk), .Q(\ram[7][147] ) );
  DFFX1_HVT \ram_reg[7][146]  ( .D(n1999), .CLK(clk), .Q(\ram[7][146] ) );
  DFFX1_HVT \ram_reg[7][145]  ( .D(n1998), .CLK(clk), .Q(\ram[7][145] ) );
  DFFX1_HVT \ram_reg[7][144]  ( .D(n1997), .CLK(clk), .Q(\ram[7][144] ) );
  DFFX1_HVT \ram_reg[7][143]  ( .D(n1996), .CLK(clk), .Q(\ram[7][143] ) );
  DFFX1_HVT \ram_reg[7][142]  ( .D(n1995), .CLK(clk), .Q(\ram[7][142] ) );
  DFFX1_HVT \ram_reg[7][141]  ( .D(n1994), .CLK(clk), .Q(\ram[7][141] ) );
  DFFX1_HVT \ram_reg[7][140]  ( .D(n1993), .CLK(clk), .Q(\ram[7][140] ) );
  DFFX1_HVT \ram_reg[7][139]  ( .D(n1992), .CLK(clk), .Q(\ram[7][139] ) );
  DFFX1_HVT \ram_reg[7][138]  ( .D(n1991), .CLK(clk), .Q(\ram[7][138] ) );
  DFFX1_HVT \ram_reg[7][137]  ( .D(n1990), .CLK(clk), .Q(\ram[7][137] ) );
  DFFX1_HVT \ram_reg[7][136]  ( .D(n1989), .CLK(clk), .Q(\ram[7][136] ) );
  DFFX1_HVT \ram_reg[7][135]  ( .D(n1988), .CLK(clk), .Q(\ram[7][135] ) );
  DFFX1_HVT \ram_reg[7][134]  ( .D(n1987), .CLK(clk), .Q(\ram[7][134] ) );
  DFFX1_HVT \ram_reg[7][133]  ( .D(n1986), .CLK(clk), .Q(\ram[7][133] ) );
  DFFX1_HVT \ram_reg[7][132]  ( .D(n1985), .CLK(clk), .Q(\ram[7][132] ) );
  DFFX1_HVT \ram_reg[7][131]  ( .D(n1984), .CLK(clk), .Q(\ram[7][131] ) );
  DFFX1_HVT \ram_reg[7][130]  ( .D(n1983), .CLK(clk), .Q(\ram[7][130] ) );
  DFFX1_HVT \ram_reg[7][129]  ( .D(n1982), .CLK(clk), .Q(\ram[7][129] ) );
  DFFX1_HVT \ram_reg[7][128]  ( .D(n1981), .CLK(clk), .Q(\ram[7][128] ) );
  DFFX1_HVT \ram_reg[7][127]  ( .D(n1980), .CLK(clk), .Q(\ram[7][127] ) );
  DFFX1_HVT \ram_reg[7][126]  ( .D(n1979), .CLK(clk), .Q(\ram[7][126] ) );
  DFFX1_HVT \ram_reg[7][125]  ( .D(n1978), .CLK(clk), .Q(\ram[7][125] ) );
  DFFX1_HVT \ram_reg[7][124]  ( .D(n1977), .CLK(clk), .Q(\ram[7][124] ) );
  DFFX1_HVT \ram_reg[7][123]  ( .D(n1976), .CLK(clk), .Q(\ram[7][123] ) );
  DFFX1_HVT \ram_reg[7][122]  ( .D(n1975), .CLK(clk), .Q(\ram[7][122] ) );
  DFFX1_HVT \ram_reg[7][121]  ( .D(n1974), .CLK(clk), .Q(\ram[7][121] ) );
  DFFX1_HVT \ram_reg[7][120]  ( .D(n1973), .CLK(clk), .Q(\ram[7][120] ) );
  DFFX1_HVT \ram_reg[7][119]  ( .D(n1972), .CLK(clk), .Q(\ram[7][119] ) );
  DFFX1_HVT \ram_reg[7][118]  ( .D(n1971), .CLK(clk), .Q(\ram[7][118] ) );
  DFFX1_HVT \ram_reg[7][117]  ( .D(n1970), .CLK(clk), .Q(\ram[7][117] ) );
  DFFX1_HVT \ram_reg[7][116]  ( .D(n1969), .CLK(clk), .Q(\ram[7][116] ) );
  DFFX1_HVT \ram_reg[7][115]  ( .D(n1968), .CLK(clk), .Q(\ram[7][115] ) );
  DFFX1_HVT \ram_reg[7][114]  ( .D(n1967), .CLK(clk), .Q(\ram[7][114] ) );
  DFFX1_HVT \ram_reg[7][113]  ( .D(n1966), .CLK(clk), .Q(\ram[7][113] ) );
  DFFX1_HVT \ram_reg[7][112]  ( .D(n1965), .CLK(clk), .Q(\ram[7][112] ) );
  DFFX1_HVT \ram_reg[7][111]  ( .D(n1964), .CLK(clk), .Q(\ram[7][111] ) );
  DFFX1_HVT \ram_reg[7][110]  ( .D(n1963), .CLK(clk), .Q(\ram[7][110] ) );
  DFFX1_HVT \ram_reg[7][109]  ( .D(n1962), .CLK(clk), .Q(\ram[7][109] ) );
  DFFX1_HVT \ram_reg[7][108]  ( .D(n1961), .CLK(clk), .Q(\ram[7][108] ) );
  DFFX1_HVT \ram_reg[7][107]  ( .D(n1960), .CLK(clk), .Q(\ram[7][107] ) );
  DFFX1_HVT \ram_reg[7][106]  ( .D(n1959), .CLK(clk), .Q(\ram[7][106] ) );
  DFFX1_HVT \ram_reg[7][105]  ( .D(n1958), .CLK(clk), .Q(\ram[7][105] ) );
  DFFX1_HVT \ram_reg[7][104]  ( .D(n1957), .CLK(clk), .Q(\ram[7][104] ) );
  DFFX1_HVT \ram_reg[7][103]  ( .D(n1956), .CLK(clk), .Q(\ram[7][103] ) );
  DFFX1_HVT \ram_reg[7][102]  ( .D(n1955), .CLK(clk), .Q(\ram[7][102] ) );
  DFFX1_HVT \ram_reg[7][101]  ( .D(n1954), .CLK(clk), .Q(\ram[7][101] ) );
  DFFX1_HVT \ram_reg[7][100]  ( .D(n1953), .CLK(clk), .Q(\ram[7][100] ) );
  DFFX1_HVT \ram_reg[7][99]  ( .D(n1952), .CLK(clk), .Q(\ram[7][99] ) );
  DFFX1_HVT \ram_reg[7][98]  ( .D(n1951), .CLK(clk), .Q(\ram[7][98] ) );
  DFFX1_HVT \ram_reg[7][97]  ( .D(n1950), .CLK(clk), .Q(\ram[7][97] ) );
  DFFX1_HVT \ram_reg[7][96]  ( .D(n1949), .CLK(clk), .Q(\ram[7][96] ) );
  DFFX1_HVT \ram_reg[7][95]  ( .D(n1948), .CLK(clk), .Q(\ram[7][95] ) );
  DFFX1_HVT \ram_reg[7][94]  ( .D(n1947), .CLK(clk), .Q(\ram[7][94] ) );
  DFFX1_HVT \ram_reg[7][93]  ( .D(n1946), .CLK(clk), .Q(\ram[7][93] ) );
  DFFX1_HVT \ram_reg[7][92]  ( .D(n1945), .CLK(clk), .Q(\ram[7][92] ) );
  DFFX1_HVT \ram_reg[7][91]  ( .D(n1944), .CLK(clk), .Q(\ram[7][91] ) );
  DFFX1_HVT \ram_reg[7][90]  ( .D(n1943), .CLK(clk), .Q(\ram[7][90] ) );
  DFFX1_HVT \ram_reg[7][89]  ( .D(n1942), .CLK(clk), .Q(\ram[7][89] ) );
  DFFX1_HVT \ram_reg[7][88]  ( .D(n1941), .CLK(clk), .Q(\ram[7][88] ) );
  DFFX1_HVT \ram_reg[7][87]  ( .D(n1940), .CLK(clk), .Q(\ram[7][87] ) );
  DFFX1_HVT \ram_reg[7][86]  ( .D(n1939), .CLK(clk), .Q(\ram[7][86] ) );
  DFFX1_HVT \ram_reg[7][85]  ( .D(n1938), .CLK(clk), .Q(\ram[7][85] ) );
  DFFX1_HVT \ram_reg[7][84]  ( .D(n1937), .CLK(clk), .Q(\ram[7][84] ) );
  DFFX1_HVT \ram_reg[7][83]  ( .D(n1936), .CLK(clk), .Q(\ram[7][83] ) );
  DFFX1_HVT \ram_reg[7][82]  ( .D(n1935), .CLK(clk), .Q(\ram[7][82] ) );
  DFFX1_HVT \ram_reg[7][81]  ( .D(n1934), .CLK(clk), .Q(\ram[7][81] ) );
  DFFX1_HVT \ram_reg[7][80]  ( .D(n1933), .CLK(clk), .Q(\ram[7][80] ) );
  DFFX1_HVT \ram_reg[7][79]  ( .D(n1932), .CLK(clk), .Q(\ram[7][79] ) );
  DFFX1_HVT \ram_reg[7][78]  ( .D(n1931), .CLK(clk), .Q(\ram[7][78] ) );
  DFFX1_HVT \ram_reg[7][77]  ( .D(n1930), .CLK(clk), .Q(\ram[7][77] ) );
  DFFX1_HVT \ram_reg[7][76]  ( .D(n1929), .CLK(clk), .Q(\ram[7][76] ) );
  DFFX1_HVT \ram_reg[7][75]  ( .D(n1928), .CLK(clk), .Q(\ram[7][75] ) );
  DFFX1_HVT \ram_reg[7][74]  ( .D(n1927), .CLK(clk), .Q(\ram[7][74] ) );
  DFFX1_HVT \ram_reg[7][73]  ( .D(n1926), .CLK(clk), .Q(\ram[7][73] ) );
  DFFX1_HVT \ram_reg[7][72]  ( .D(n1925), .CLK(clk), .Q(\ram[7][72] ) );
  DFFX1_HVT \ram_reg[7][71]  ( .D(n1924), .CLK(clk), .Q(\ram[7][71] ) );
  DFFX1_HVT \ram_reg[7][70]  ( .D(n1923), .CLK(clk), .Q(\ram[7][70] ) );
  DFFX1_HVT \ram_reg[7][69]  ( .D(n1922), .CLK(clk), .Q(\ram[7][69] ) );
  DFFX1_HVT \ram_reg[7][68]  ( .D(n1921), .CLK(clk), .Q(\ram[7][68] ) );
  DFFX1_HVT \ram_reg[7][67]  ( .D(n1920), .CLK(clk), .Q(\ram[7][67] ) );
  DFFX1_HVT \ram_reg[7][66]  ( .D(n1919), .CLK(clk), .Q(\ram[7][66] ) );
  DFFX1_HVT \ram_reg[7][65]  ( .D(n1918), .CLK(clk), .Q(\ram[7][65] ) );
  DFFX1_HVT \ram_reg[7][64]  ( .D(n1917), .CLK(clk), .Q(\ram[7][64] ) );
  DFFX1_HVT \ram_reg[7][63]  ( .D(n1916), .CLK(clk), .Q(\ram[7][63] ) );
  DFFX1_HVT \ram_reg[7][62]  ( .D(n1915), .CLK(clk), .Q(\ram[7][62] ) );
  DFFX1_HVT \ram_reg[7][61]  ( .D(n1914), .CLK(clk), .Q(\ram[7][61] ) );
  DFFX1_HVT \ram_reg[7][60]  ( .D(n1913), .CLK(clk), .Q(\ram[7][60] ) );
  DFFX1_HVT \ram_reg[7][59]  ( .D(n1912), .CLK(clk), .Q(\ram[7][59] ) );
  DFFX1_HVT \ram_reg[7][58]  ( .D(n1911), .CLK(clk), .Q(\ram[7][58] ) );
  DFFX1_HVT \ram_reg[7][57]  ( .D(n1910), .CLK(clk), .Q(\ram[7][57] ) );
  DFFX1_HVT \ram_reg[7][56]  ( .D(n1909), .CLK(clk), .Q(\ram[7][56] ) );
  DFFX1_HVT \ram_reg[7][55]  ( .D(n1908), .CLK(clk), .Q(\ram[7][55] ) );
  DFFX1_HVT \ram_reg[7][54]  ( .D(n1907), .CLK(clk), .Q(\ram[7][54] ) );
  DFFX1_HVT \ram_reg[7][53]  ( .D(n1906), .CLK(clk), .Q(\ram[7][53] ) );
  DFFX1_HVT \ram_reg[7][52]  ( .D(n1905), .CLK(clk), .Q(\ram[7][52] ) );
  DFFX1_HVT \ram_reg[7][51]  ( .D(n1904), .CLK(clk), .Q(\ram[7][51] ) );
  DFFX1_HVT \ram_reg[7][50]  ( .D(n1903), .CLK(clk), .Q(\ram[7][50] ) );
  DFFX1_HVT \ram_reg[7][49]  ( .D(n1902), .CLK(clk), .Q(\ram[7][49] ) );
  DFFX1_HVT \ram_reg[7][48]  ( .D(n1901), .CLK(clk), .Q(\ram[7][48] ) );
  DFFX1_HVT \ram_reg[7][47]  ( .D(n1900), .CLK(clk), .Q(\ram[7][47] ) );
  DFFX1_HVT \ram_reg[7][46]  ( .D(n1899), .CLK(clk), .Q(\ram[7][46] ) );
  DFFX1_HVT \ram_reg[7][45]  ( .D(n1898), .CLK(clk), .Q(\ram[7][45] ) );
  DFFX1_HVT \ram_reg[7][44]  ( .D(n1897), .CLK(clk), .Q(\ram[7][44] ) );
  DFFX1_HVT \ram_reg[7][43]  ( .D(n1896), .CLK(clk), .Q(\ram[7][43] ) );
  DFFX1_HVT \ram_reg[7][42]  ( .D(n1895), .CLK(clk), .Q(\ram[7][42] ) );
  DFFX1_HVT \ram_reg[7][41]  ( .D(n1894), .CLK(clk), .Q(\ram[7][41] ) );
  DFFX1_HVT \ram_reg[7][40]  ( .D(n1893), .CLK(clk), .Q(\ram[7][40] ) );
  DFFX1_HVT \ram_reg[7][39]  ( .D(n1892), .CLK(clk), .Q(\ram[7][39] ) );
  DFFX1_HVT \ram_reg[7][38]  ( .D(n1891), .CLK(clk), .Q(\ram[7][38] ) );
  DFFX1_HVT \ram_reg[7][37]  ( .D(n1890), .CLK(clk), .Q(\ram[7][37] ) );
  DFFX1_HVT \ram_reg[7][36]  ( .D(n1889), .CLK(clk), .Q(\ram[7][36] ) );
  DFFX1_HVT \ram_reg[7][35]  ( .D(n1888), .CLK(clk), .Q(\ram[7][35] ) );
  DFFX1_HVT \ram_reg[7][34]  ( .D(n1887), .CLK(clk), .Q(\ram[7][34] ) );
  DFFX1_HVT \ram_reg[7][33]  ( .D(n1886), .CLK(clk), .Q(\ram[7][33] ) );
  DFFX1_HVT \ram_reg[7][32]  ( .D(n1885), .CLK(clk), .Q(\ram[7][32] ) );
  DFFX1_HVT \ram_reg[7][31]  ( .D(n1884), .CLK(clk), .Q(\ram[7][31] ) );
  DFFX1_HVT \ram_reg[7][30]  ( .D(n1883), .CLK(clk), .Q(\ram[7][30] ) );
  DFFX1_HVT \ram_reg[7][29]  ( .D(n1882), .CLK(clk), .Q(\ram[7][29] ) );
  DFFX1_HVT \ram_reg[7][28]  ( .D(n1881), .CLK(clk), .Q(\ram[7][28] ) );
  DFFX1_HVT \ram_reg[7][27]  ( .D(n1880), .CLK(clk), .Q(\ram[7][27] ) );
  DFFX1_HVT \ram_reg[7][26]  ( .D(n1879), .CLK(clk), .Q(\ram[7][26] ) );
  DFFX1_HVT \ram_reg[7][25]  ( .D(n1878), .CLK(clk), .Q(\ram[7][25] ) );
  DFFX1_HVT \ram_reg[7][24]  ( .D(n1877), .CLK(clk), .Q(\ram[7][24] ) );
  DFFX1_HVT \ram_reg[7][23]  ( .D(n1876), .CLK(clk), .Q(\ram[7][23] ) );
  DFFX1_HVT \ram_reg[7][22]  ( .D(n1875), .CLK(clk), .Q(\ram[7][22] ) );
  DFFX1_HVT \ram_reg[7][21]  ( .D(n1874), .CLK(clk), .Q(\ram[7][21] ) );
  DFFX1_HVT \ram_reg[7][20]  ( .D(n1873), .CLK(clk), .Q(\ram[7][20] ) );
  DFFX1_HVT \ram_reg[7][19]  ( .D(n1872), .CLK(clk), .Q(\ram[7][19] ) );
  DFFX1_HVT \ram_reg[7][18]  ( .D(n1871), .CLK(clk), .Q(\ram[7][18] ) );
  DFFX1_HVT \ram_reg[7][17]  ( .D(n1870), .CLK(clk), .Q(\ram[7][17] ) );
  DFFX1_HVT \ram_reg[7][16]  ( .D(n1869), .CLK(clk), .Q(\ram[7][16] ) );
  DFFX1_HVT \ram_reg[7][15]  ( .D(n1868), .CLK(clk), .Q(\ram[7][15] ) );
  DFFX1_HVT \ram_reg[7][14]  ( .D(n1867), .CLK(clk), .Q(\ram[7][14] ) );
  DFFX1_HVT \ram_reg[7][13]  ( .D(n1866), .CLK(clk), .Q(\ram[7][13] ) );
  DFFX1_HVT \ram_reg[7][12]  ( .D(n1865), .CLK(clk), .Q(\ram[7][12] ) );
  DFFX1_HVT \ram_reg[7][11]  ( .D(n1864), .CLK(clk), .Q(\ram[7][11] ) );
  DFFX1_HVT \ram_reg[7][10]  ( .D(n1863), .CLK(clk), .Q(\ram[7][10] ) );
  DFFX1_HVT \ram_reg[7][9]  ( .D(n1862), .CLK(clk), .Q(\ram[7][9] ) );
  DFFX1_HVT \ram_reg[7][8]  ( .D(n1861), .CLK(clk), .Q(\ram[7][8] ) );
  DFFX1_HVT \ram_reg[7][7]  ( .D(n1860), .CLK(clk), .Q(\ram[7][7] ) );
  DFFX1_HVT \ram_reg[7][6]  ( .D(n1859), .CLK(clk), .Q(\ram[7][6] ) );
  DFFX1_HVT \ram_reg[7][5]  ( .D(n1858), .CLK(clk), .Q(\ram[7][5] ) );
  DFFX1_HVT \ram_reg[7][4]  ( .D(n1857), .CLK(clk), .Q(\ram[7][4] ) );
  DFFX1_HVT \ram_reg[7][3]  ( .D(n1856), .CLK(clk), .Q(\ram[7][3] ) );
  DFFX1_HVT \ram_reg[7][2]  ( .D(n1855), .CLK(clk), .Q(\ram[7][2] ) );
  DFFX1_HVT \ram_reg[7][1]  ( .D(n1854), .CLK(clk), .Q(\ram[7][1] ) );
  DFFX1_HVT \ram_reg[7][0]  ( .D(n1853), .CLK(clk), .Q(\ram[7][0] ) );
  DFFX1_HVT \ram_reg[6][255]  ( .D(n1852), .CLK(clk), .Q(\ram[6][255] ) );
  DFFX1_HVT \ram_reg[6][254]  ( .D(n1851), .CLK(clk), .Q(\ram[6][254] ) );
  DFFX1_HVT \ram_reg[6][253]  ( .D(n1850), .CLK(clk), .Q(\ram[6][253] ) );
  DFFX1_HVT \ram_reg[6][252]  ( .D(n1849), .CLK(clk), .Q(\ram[6][252] ) );
  DFFX1_HVT \ram_reg[6][251]  ( .D(n1848), .CLK(clk), .Q(\ram[6][251] ) );
  DFFX1_HVT \ram_reg[6][250]  ( .D(n1847), .CLK(clk), .Q(\ram[6][250] ) );
  DFFX1_HVT \ram_reg[6][249]  ( .D(n1846), .CLK(clk), .Q(\ram[6][249] ) );
  DFFX1_HVT \ram_reg[6][248]  ( .D(n1845), .CLK(clk), .Q(\ram[6][248] ) );
  DFFX1_HVT \ram_reg[6][247]  ( .D(n1844), .CLK(clk), .Q(\ram[6][247] ) );
  DFFX1_HVT \ram_reg[6][246]  ( .D(n1843), .CLK(clk), .Q(\ram[6][246] ) );
  DFFX1_HVT \ram_reg[6][245]  ( .D(n1842), .CLK(clk), .Q(\ram[6][245] ) );
  DFFX1_HVT \ram_reg[6][244]  ( .D(n1841), .CLK(clk), .Q(\ram[6][244] ) );
  DFFX1_HVT \ram_reg[6][243]  ( .D(n1840), .CLK(clk), .Q(\ram[6][243] ) );
  DFFX1_HVT \ram_reg[6][242]  ( .D(n1839), .CLK(clk), .Q(\ram[6][242] ) );
  DFFX1_HVT \ram_reg[6][241]  ( .D(n1838), .CLK(clk), .Q(\ram[6][241] ) );
  DFFX1_HVT \ram_reg[6][240]  ( .D(n1837), .CLK(clk), .Q(\ram[6][240] ) );
  DFFX1_HVT \ram_reg[6][239]  ( .D(n1836), .CLK(clk), .Q(\ram[6][239] ) );
  DFFX1_HVT \ram_reg[6][238]  ( .D(n1835), .CLK(clk), .Q(\ram[6][238] ) );
  DFFX1_HVT \ram_reg[6][237]  ( .D(n1834), .CLK(clk), .Q(\ram[6][237] ) );
  DFFX1_HVT \ram_reg[6][236]  ( .D(n1833), .CLK(clk), .Q(\ram[6][236] ) );
  DFFX1_HVT \ram_reg[6][235]  ( .D(n1832), .CLK(clk), .Q(\ram[6][235] ) );
  DFFX1_HVT \ram_reg[6][234]  ( .D(n1831), .CLK(clk), .Q(\ram[6][234] ) );
  DFFX1_HVT \ram_reg[6][233]  ( .D(n1830), .CLK(clk), .Q(\ram[6][233] ) );
  DFFX1_HVT \ram_reg[6][232]  ( .D(n1829), .CLK(clk), .Q(\ram[6][232] ) );
  DFFX1_HVT \ram_reg[6][231]  ( .D(n1828), .CLK(clk), .Q(\ram[6][231] ) );
  DFFX1_HVT \ram_reg[6][230]  ( .D(n1827), .CLK(clk), .Q(\ram[6][230] ) );
  DFFX1_HVT \ram_reg[6][229]  ( .D(n1826), .CLK(clk), .Q(\ram[6][229] ) );
  DFFX1_HVT \ram_reg[6][228]  ( .D(n1825), .CLK(clk), .Q(\ram[6][228] ) );
  DFFX1_HVT \ram_reg[6][227]  ( .D(n1824), .CLK(clk), .Q(\ram[6][227] ) );
  DFFX1_HVT \ram_reg[6][226]  ( .D(n1823), .CLK(clk), .Q(\ram[6][226] ) );
  DFFX1_HVT \ram_reg[6][225]  ( .D(n1822), .CLK(clk), .Q(\ram[6][225] ) );
  DFFX1_HVT \ram_reg[6][224]  ( .D(n1821), .CLK(clk), .Q(\ram[6][224] ) );
  DFFX1_HVT \ram_reg[6][223]  ( .D(n1820), .CLK(clk), .Q(\ram[6][223] ) );
  DFFX1_HVT \ram_reg[6][222]  ( .D(n1819), .CLK(clk), .Q(\ram[6][222] ) );
  DFFX1_HVT \ram_reg[6][221]  ( .D(n1818), .CLK(clk), .Q(\ram[6][221] ) );
  DFFX1_HVT \ram_reg[6][220]  ( .D(n1817), .CLK(clk), .Q(\ram[6][220] ) );
  DFFX1_HVT \ram_reg[6][219]  ( .D(n1816), .CLK(clk), .Q(\ram[6][219] ) );
  DFFX1_HVT \ram_reg[6][218]  ( .D(n1815), .CLK(clk), .Q(\ram[6][218] ) );
  DFFX1_HVT \ram_reg[6][217]  ( .D(n1814), .CLK(clk), .Q(\ram[6][217] ) );
  DFFX1_HVT \ram_reg[6][216]  ( .D(n1813), .CLK(clk), .Q(\ram[6][216] ) );
  DFFX1_HVT \ram_reg[6][215]  ( .D(n1812), .CLK(clk), .Q(\ram[6][215] ) );
  DFFX1_HVT \ram_reg[6][214]  ( .D(n1811), .CLK(clk), .Q(\ram[6][214] ) );
  DFFX1_HVT \ram_reg[6][213]  ( .D(n1810), .CLK(clk), .Q(\ram[6][213] ) );
  DFFX1_HVT \ram_reg[6][212]  ( .D(n1809), .CLK(clk), .Q(\ram[6][212] ) );
  DFFX1_HVT \ram_reg[6][211]  ( .D(n1808), .CLK(clk), .Q(\ram[6][211] ) );
  DFFX1_HVT \ram_reg[6][210]  ( .D(n1807), .CLK(clk), .Q(\ram[6][210] ) );
  DFFX1_HVT \ram_reg[6][209]  ( .D(n1806), .CLK(clk), .Q(\ram[6][209] ) );
  DFFX1_HVT \ram_reg[6][208]  ( .D(n1805), .CLK(clk), .Q(\ram[6][208] ) );
  DFFX1_HVT \ram_reg[6][207]  ( .D(n1804), .CLK(clk), .Q(\ram[6][207] ) );
  DFFX1_HVT \ram_reg[6][206]  ( .D(n1803), .CLK(clk), .Q(\ram[6][206] ) );
  DFFX1_HVT \ram_reg[6][205]  ( .D(n1802), .CLK(clk), .Q(\ram[6][205] ) );
  DFFX1_HVT \ram_reg[6][204]  ( .D(n1801), .CLK(clk), .Q(\ram[6][204] ) );
  DFFX1_HVT \ram_reg[6][203]  ( .D(n1800), .CLK(clk), .Q(\ram[6][203] ) );
  DFFX1_HVT \ram_reg[6][202]  ( .D(n1799), .CLK(clk), .Q(\ram[6][202] ) );
  DFFX1_HVT \ram_reg[6][201]  ( .D(n1798), .CLK(clk), .Q(\ram[6][201] ) );
  DFFX1_HVT \ram_reg[6][200]  ( .D(n1797), .CLK(clk), .Q(\ram[6][200] ) );
  DFFX1_HVT \ram_reg[6][199]  ( .D(n1796), .CLK(clk), .Q(\ram[6][199] ) );
  DFFX1_HVT \ram_reg[6][198]  ( .D(n1795), .CLK(clk), .Q(\ram[6][198] ) );
  DFFX1_HVT \ram_reg[6][197]  ( .D(n1794), .CLK(clk), .Q(\ram[6][197] ) );
  DFFX1_HVT \ram_reg[6][196]  ( .D(n1793), .CLK(clk), .Q(\ram[6][196] ) );
  DFFX1_HVT \ram_reg[6][195]  ( .D(n1792), .CLK(clk), .Q(\ram[6][195] ) );
  DFFX1_HVT \ram_reg[6][194]  ( .D(n1791), .CLK(clk), .Q(\ram[6][194] ) );
  DFFX1_HVT \ram_reg[6][193]  ( .D(n1790), .CLK(clk), .Q(\ram[6][193] ) );
  DFFX1_HVT \ram_reg[6][192]  ( .D(n1789), .CLK(clk), .Q(\ram[6][192] ) );
  DFFX1_HVT \ram_reg[6][191]  ( .D(n1788), .CLK(clk), .Q(\ram[6][191] ) );
  DFFX1_HVT \ram_reg[6][190]  ( .D(n1787), .CLK(clk), .Q(\ram[6][190] ) );
  DFFX1_HVT \ram_reg[6][189]  ( .D(n1786), .CLK(clk), .Q(\ram[6][189] ) );
  DFFX1_HVT \ram_reg[6][188]  ( .D(n1785), .CLK(clk), .Q(\ram[6][188] ) );
  DFFX1_HVT \ram_reg[6][187]  ( .D(n1784), .CLK(clk), .Q(\ram[6][187] ) );
  DFFX1_HVT \ram_reg[6][186]  ( .D(n1783), .CLK(clk), .Q(\ram[6][186] ) );
  DFFX1_HVT \ram_reg[6][185]  ( .D(n1782), .CLK(clk), .Q(\ram[6][185] ) );
  DFFX1_HVT \ram_reg[6][184]  ( .D(n1781), .CLK(clk), .Q(\ram[6][184] ) );
  DFFX1_HVT \ram_reg[6][183]  ( .D(n1780), .CLK(clk), .Q(\ram[6][183] ) );
  DFFX1_HVT \ram_reg[6][182]  ( .D(n1779), .CLK(clk), .Q(\ram[6][182] ) );
  DFFX1_HVT \ram_reg[6][181]  ( .D(n1778), .CLK(clk), .Q(\ram[6][181] ) );
  DFFX1_HVT \ram_reg[6][180]  ( .D(n1777), .CLK(clk), .Q(\ram[6][180] ) );
  DFFX1_HVT \ram_reg[6][179]  ( .D(n1776), .CLK(clk), .Q(\ram[6][179] ) );
  DFFX1_HVT \ram_reg[6][178]  ( .D(n1775), .CLK(clk), .Q(\ram[6][178] ) );
  DFFX1_HVT \ram_reg[6][177]  ( .D(n1774), .CLK(clk), .Q(\ram[6][177] ) );
  DFFX1_HVT \ram_reg[6][176]  ( .D(n1773), .CLK(clk), .Q(\ram[6][176] ) );
  DFFX1_HVT \ram_reg[6][175]  ( .D(n1772), .CLK(clk), .Q(\ram[6][175] ) );
  DFFX1_HVT \ram_reg[6][174]  ( .D(n1771), .CLK(clk), .Q(\ram[6][174] ) );
  DFFX1_HVT \ram_reg[6][173]  ( .D(n1770), .CLK(clk), .Q(\ram[6][173] ) );
  DFFX1_HVT \ram_reg[6][172]  ( .D(n1769), .CLK(clk), .Q(\ram[6][172] ) );
  DFFX1_HVT \ram_reg[6][171]  ( .D(n1768), .CLK(clk), .Q(\ram[6][171] ) );
  DFFX1_HVT \ram_reg[6][170]  ( .D(n1767), .CLK(clk), .Q(\ram[6][170] ) );
  DFFX1_HVT \ram_reg[6][169]  ( .D(n1766), .CLK(clk), .Q(\ram[6][169] ) );
  DFFX1_HVT \ram_reg[6][168]  ( .D(n1765), .CLK(clk), .Q(\ram[6][168] ) );
  DFFX1_HVT \ram_reg[6][167]  ( .D(n1764), .CLK(clk), .Q(\ram[6][167] ) );
  DFFX1_HVT \ram_reg[6][166]  ( .D(n1763), .CLK(clk), .Q(\ram[6][166] ) );
  DFFX1_HVT \ram_reg[6][165]  ( .D(n1762), .CLK(clk), .Q(\ram[6][165] ) );
  DFFX1_HVT \ram_reg[6][164]  ( .D(n1761), .CLK(clk), .Q(\ram[6][164] ) );
  DFFX1_HVT \ram_reg[6][163]  ( .D(n1760), .CLK(clk), .Q(\ram[6][163] ) );
  DFFX1_HVT \ram_reg[6][162]  ( .D(n1759), .CLK(clk), .Q(\ram[6][162] ) );
  DFFX1_HVT \ram_reg[6][161]  ( .D(n1758), .CLK(clk), .Q(\ram[6][161] ) );
  DFFX1_HVT \ram_reg[6][160]  ( .D(n1757), .CLK(clk), .Q(\ram[6][160] ) );
  DFFX1_HVT \ram_reg[6][159]  ( .D(n1756), .CLK(clk), .Q(\ram[6][159] ) );
  DFFX1_HVT \ram_reg[6][158]  ( .D(n1755), .CLK(clk), .Q(\ram[6][158] ) );
  DFFX1_HVT \ram_reg[6][157]  ( .D(n1754), .CLK(clk), .Q(\ram[6][157] ) );
  DFFX1_HVT \ram_reg[6][156]  ( .D(n1753), .CLK(clk), .Q(\ram[6][156] ) );
  DFFX1_HVT \ram_reg[6][155]  ( .D(n1752), .CLK(clk), .Q(\ram[6][155] ) );
  DFFX1_HVT \ram_reg[6][154]  ( .D(n1751), .CLK(clk), .Q(\ram[6][154] ) );
  DFFX1_HVT \ram_reg[6][153]  ( .D(n1750), .CLK(clk), .Q(\ram[6][153] ) );
  DFFX1_HVT \ram_reg[6][152]  ( .D(n1749), .CLK(clk), .Q(\ram[6][152] ) );
  DFFX1_HVT \ram_reg[6][151]  ( .D(n1748), .CLK(clk), .Q(\ram[6][151] ) );
  DFFX1_HVT \ram_reg[6][150]  ( .D(n1747), .CLK(clk), .Q(\ram[6][150] ) );
  DFFX1_HVT \ram_reg[6][149]  ( .D(n1746), .CLK(clk), .Q(\ram[6][149] ) );
  DFFX1_HVT \ram_reg[6][148]  ( .D(n1745), .CLK(clk), .Q(\ram[6][148] ) );
  DFFX1_HVT \ram_reg[6][147]  ( .D(n1744), .CLK(clk), .Q(\ram[6][147] ) );
  DFFX1_HVT \ram_reg[6][146]  ( .D(n1743), .CLK(clk), .Q(\ram[6][146] ) );
  DFFX1_HVT \ram_reg[6][145]  ( .D(n1742), .CLK(clk), .Q(\ram[6][145] ) );
  DFFX1_HVT \ram_reg[6][144]  ( .D(n1741), .CLK(clk), .Q(\ram[6][144] ) );
  DFFX1_HVT \ram_reg[6][143]  ( .D(n1740), .CLK(clk), .Q(\ram[6][143] ) );
  DFFX1_HVT \ram_reg[6][142]  ( .D(n1739), .CLK(clk), .Q(\ram[6][142] ) );
  DFFX1_HVT \ram_reg[6][141]  ( .D(n1738), .CLK(clk), .Q(\ram[6][141] ) );
  DFFX1_HVT \ram_reg[6][140]  ( .D(n1737), .CLK(clk), .Q(\ram[6][140] ) );
  DFFX1_HVT \ram_reg[6][139]  ( .D(n1736), .CLK(clk), .Q(\ram[6][139] ) );
  DFFX1_HVT \ram_reg[6][138]  ( .D(n1735), .CLK(clk), .Q(\ram[6][138] ) );
  DFFX1_HVT \ram_reg[6][137]  ( .D(n1734), .CLK(clk), .Q(\ram[6][137] ) );
  DFFX1_HVT \ram_reg[6][136]  ( .D(n1733), .CLK(clk), .Q(\ram[6][136] ) );
  DFFX1_HVT \ram_reg[6][135]  ( .D(n1732), .CLK(clk), .Q(\ram[6][135] ) );
  DFFX1_HVT \ram_reg[6][134]  ( .D(n1731), .CLK(clk), .Q(\ram[6][134] ) );
  DFFX1_HVT \ram_reg[6][133]  ( .D(n1730), .CLK(clk), .Q(\ram[6][133] ) );
  DFFX1_HVT \ram_reg[6][132]  ( .D(n1729), .CLK(clk), .Q(\ram[6][132] ) );
  DFFX1_HVT \ram_reg[6][131]  ( .D(n1728), .CLK(clk), .Q(\ram[6][131] ) );
  DFFX1_HVT \ram_reg[6][130]  ( .D(n1727), .CLK(clk), .Q(\ram[6][130] ) );
  DFFX1_HVT \ram_reg[6][129]  ( .D(n1726), .CLK(clk), .Q(\ram[6][129] ) );
  DFFX1_HVT \ram_reg[6][128]  ( .D(n1725), .CLK(clk), .Q(\ram[6][128] ) );
  DFFX1_HVT \ram_reg[6][127]  ( .D(n1724), .CLK(clk), .Q(\ram[6][127] ) );
  DFFX1_HVT \ram_reg[6][126]  ( .D(n1723), .CLK(clk), .Q(\ram[6][126] ) );
  DFFX1_HVT \ram_reg[6][125]  ( .D(n1722), .CLK(clk), .Q(\ram[6][125] ) );
  DFFX1_HVT \ram_reg[6][124]  ( .D(n1721), .CLK(clk), .Q(\ram[6][124] ) );
  DFFX1_HVT \ram_reg[6][123]  ( .D(n1720), .CLK(clk), .Q(\ram[6][123] ) );
  DFFX1_HVT \ram_reg[6][122]  ( .D(n1719), .CLK(clk), .Q(\ram[6][122] ) );
  DFFX1_HVT \ram_reg[6][121]  ( .D(n1718), .CLK(clk), .Q(\ram[6][121] ) );
  DFFX1_HVT \ram_reg[6][120]  ( .D(n1717), .CLK(clk), .Q(\ram[6][120] ) );
  DFFX1_HVT \ram_reg[6][119]  ( .D(n1716), .CLK(clk), .Q(\ram[6][119] ) );
  DFFX1_HVT \ram_reg[6][118]  ( .D(n1715), .CLK(clk), .Q(\ram[6][118] ) );
  DFFX1_HVT \ram_reg[6][117]  ( .D(n1714), .CLK(clk), .Q(\ram[6][117] ) );
  DFFX1_HVT \ram_reg[6][116]  ( .D(n1713), .CLK(clk), .Q(\ram[6][116] ) );
  DFFX1_HVT \ram_reg[6][115]  ( .D(n1712), .CLK(clk), .Q(\ram[6][115] ) );
  DFFX1_HVT \ram_reg[6][114]  ( .D(n1711), .CLK(clk), .Q(\ram[6][114] ) );
  DFFX1_HVT \ram_reg[6][113]  ( .D(n1710), .CLK(clk), .Q(\ram[6][113] ) );
  DFFX1_HVT \ram_reg[6][112]  ( .D(n1709), .CLK(clk), .Q(\ram[6][112] ) );
  DFFX1_HVT \ram_reg[6][111]  ( .D(n1708), .CLK(clk), .Q(\ram[6][111] ) );
  DFFX1_HVT \ram_reg[6][110]  ( .D(n1707), .CLK(clk), .Q(\ram[6][110] ) );
  DFFX1_HVT \ram_reg[6][109]  ( .D(n1706), .CLK(clk), .Q(\ram[6][109] ) );
  DFFX1_HVT \ram_reg[6][108]  ( .D(n1705), .CLK(clk), .Q(\ram[6][108] ) );
  DFFX1_HVT \ram_reg[6][107]  ( .D(n1704), .CLK(clk), .Q(\ram[6][107] ) );
  DFFX1_HVT \ram_reg[6][106]  ( .D(n1703), .CLK(clk), .Q(\ram[6][106] ) );
  DFFX1_HVT \ram_reg[6][105]  ( .D(n1702), .CLK(clk), .Q(\ram[6][105] ) );
  DFFX1_HVT \ram_reg[6][104]  ( .D(n1701), .CLK(clk), .Q(\ram[6][104] ) );
  DFFX1_HVT \ram_reg[6][103]  ( .D(n1700), .CLK(clk), .Q(\ram[6][103] ) );
  DFFX1_HVT \ram_reg[6][102]  ( .D(n1699), .CLK(clk), .Q(\ram[6][102] ) );
  DFFX1_HVT \ram_reg[6][101]  ( .D(n1698), .CLK(clk), .Q(\ram[6][101] ) );
  DFFX1_HVT \ram_reg[6][100]  ( .D(n1697), .CLK(clk), .Q(\ram[6][100] ) );
  DFFX1_HVT \ram_reg[6][99]  ( .D(n1696), .CLK(clk), .Q(\ram[6][99] ) );
  DFFX1_HVT \ram_reg[6][98]  ( .D(n1695), .CLK(clk), .Q(\ram[6][98] ) );
  DFFX1_HVT \ram_reg[6][97]  ( .D(n1694), .CLK(clk), .Q(\ram[6][97] ) );
  DFFX1_HVT \ram_reg[6][96]  ( .D(n1693), .CLK(clk), .Q(\ram[6][96] ) );
  DFFX1_HVT \ram_reg[6][95]  ( .D(n1692), .CLK(clk), .Q(\ram[6][95] ) );
  DFFX1_HVT \ram_reg[6][94]  ( .D(n1691), .CLK(clk), .Q(\ram[6][94] ) );
  DFFX1_HVT \ram_reg[6][93]  ( .D(n1690), .CLK(clk), .Q(\ram[6][93] ) );
  DFFX1_HVT \ram_reg[6][92]  ( .D(n1689), .CLK(clk), .Q(\ram[6][92] ) );
  DFFX1_HVT \ram_reg[6][91]  ( .D(n1688), .CLK(clk), .Q(\ram[6][91] ) );
  DFFX1_HVT \ram_reg[6][90]  ( .D(n1687), .CLK(clk), .Q(\ram[6][90] ) );
  DFFX1_HVT \ram_reg[6][89]  ( .D(n1686), .CLK(clk), .Q(\ram[6][89] ) );
  DFFX1_HVT \ram_reg[6][88]  ( .D(n1685), .CLK(clk), .Q(\ram[6][88] ) );
  DFFX1_HVT \ram_reg[6][87]  ( .D(n1684), .CLK(clk), .Q(\ram[6][87] ) );
  DFFX1_HVT \ram_reg[6][86]  ( .D(n1683), .CLK(clk), .Q(\ram[6][86] ) );
  DFFX1_HVT \ram_reg[6][85]  ( .D(n1682), .CLK(clk), .Q(\ram[6][85] ) );
  DFFX1_HVT \ram_reg[6][84]  ( .D(n1681), .CLK(clk), .Q(\ram[6][84] ) );
  DFFX1_HVT \ram_reg[6][83]  ( .D(n1680), .CLK(clk), .Q(\ram[6][83] ) );
  DFFX1_HVT \ram_reg[6][82]  ( .D(n1679), .CLK(clk), .Q(\ram[6][82] ) );
  DFFX1_HVT \ram_reg[6][81]  ( .D(n1678), .CLK(clk), .Q(\ram[6][81] ) );
  DFFX1_HVT \ram_reg[6][80]  ( .D(n1677), .CLK(clk), .Q(\ram[6][80] ) );
  DFFX1_HVT \ram_reg[6][79]  ( .D(n1676), .CLK(clk), .Q(\ram[6][79] ) );
  DFFX1_HVT \ram_reg[6][78]  ( .D(n1675), .CLK(clk), .Q(\ram[6][78] ) );
  DFFX1_HVT \ram_reg[6][77]  ( .D(n1674), .CLK(clk), .Q(\ram[6][77] ) );
  DFFX1_HVT \ram_reg[6][76]  ( .D(n1673), .CLK(clk), .Q(\ram[6][76] ) );
  DFFX1_HVT \ram_reg[6][75]  ( .D(n1672), .CLK(clk), .Q(\ram[6][75] ) );
  DFFX1_HVT \ram_reg[6][74]  ( .D(n1671), .CLK(clk), .Q(\ram[6][74] ) );
  DFFX1_HVT \ram_reg[6][73]  ( .D(n1670), .CLK(clk), .Q(\ram[6][73] ) );
  DFFX1_HVT \ram_reg[6][72]  ( .D(n1669), .CLK(clk), .Q(\ram[6][72] ) );
  DFFX1_HVT \ram_reg[6][71]  ( .D(n1668), .CLK(clk), .Q(\ram[6][71] ) );
  DFFX1_HVT \ram_reg[6][70]  ( .D(n1667), .CLK(clk), .Q(\ram[6][70] ) );
  DFFX1_HVT \ram_reg[6][69]  ( .D(n1666), .CLK(clk), .Q(\ram[6][69] ) );
  DFFX1_HVT \ram_reg[6][68]  ( .D(n1665), .CLK(clk), .Q(\ram[6][68] ) );
  DFFX1_HVT \ram_reg[6][67]  ( .D(n1664), .CLK(clk), .Q(\ram[6][67] ) );
  DFFX1_HVT \ram_reg[6][66]  ( .D(n1663), .CLK(clk), .Q(\ram[6][66] ) );
  DFFX1_HVT \ram_reg[6][65]  ( .D(n1662), .CLK(clk), .Q(\ram[6][65] ) );
  DFFX1_HVT \ram_reg[6][64]  ( .D(n1661), .CLK(clk), .Q(\ram[6][64] ) );
  DFFX1_HVT \ram_reg[6][63]  ( .D(n1660), .CLK(clk), .Q(\ram[6][63] ) );
  DFFX1_HVT \ram_reg[6][62]  ( .D(n1659), .CLK(clk), .Q(\ram[6][62] ) );
  DFFX1_HVT \ram_reg[6][61]  ( .D(n1658), .CLK(clk), .Q(\ram[6][61] ) );
  DFFX1_HVT \ram_reg[6][60]  ( .D(n1657), .CLK(clk), .Q(\ram[6][60] ) );
  DFFX1_HVT \ram_reg[6][59]  ( .D(n1656), .CLK(clk), .Q(\ram[6][59] ) );
  DFFX1_HVT \ram_reg[6][58]  ( .D(n1655), .CLK(clk), .Q(\ram[6][58] ) );
  DFFX1_HVT \ram_reg[6][57]  ( .D(n1654), .CLK(clk), .Q(\ram[6][57] ) );
  DFFX1_HVT \ram_reg[6][56]  ( .D(n1653), .CLK(clk), .Q(\ram[6][56] ) );
  DFFX1_HVT \ram_reg[6][55]  ( .D(n1652), .CLK(clk), .Q(\ram[6][55] ) );
  DFFX1_HVT \ram_reg[6][54]  ( .D(n1651), .CLK(clk), .Q(\ram[6][54] ) );
  DFFX1_HVT \ram_reg[6][53]  ( .D(n1650), .CLK(clk), .Q(\ram[6][53] ) );
  DFFX1_HVT \ram_reg[6][52]  ( .D(n1649), .CLK(clk), .Q(\ram[6][52] ) );
  DFFX1_HVT \ram_reg[6][51]  ( .D(n1648), .CLK(clk), .Q(\ram[6][51] ) );
  DFFX1_HVT \ram_reg[6][50]  ( .D(n1647), .CLK(clk), .Q(\ram[6][50] ) );
  DFFX1_HVT \ram_reg[6][49]  ( .D(n1646), .CLK(clk), .Q(\ram[6][49] ) );
  DFFX1_HVT \ram_reg[6][48]  ( .D(n1645), .CLK(clk), .Q(\ram[6][48] ) );
  DFFX1_HVT \ram_reg[6][47]  ( .D(n1644), .CLK(clk), .Q(\ram[6][47] ) );
  DFFX1_HVT \ram_reg[6][46]  ( .D(n1643), .CLK(clk), .Q(\ram[6][46] ) );
  DFFX1_HVT \ram_reg[6][45]  ( .D(n1642), .CLK(clk), .Q(\ram[6][45] ) );
  DFFX1_HVT \ram_reg[6][44]  ( .D(n1641), .CLK(clk), .Q(\ram[6][44] ) );
  DFFX1_HVT \ram_reg[6][43]  ( .D(n1640), .CLK(clk), .Q(\ram[6][43] ) );
  DFFX1_HVT \ram_reg[6][42]  ( .D(n1639), .CLK(clk), .Q(\ram[6][42] ) );
  DFFX1_HVT \ram_reg[6][41]  ( .D(n1638), .CLK(clk), .Q(\ram[6][41] ) );
  DFFX1_HVT \ram_reg[6][40]  ( .D(n1637), .CLK(clk), .Q(\ram[6][40] ) );
  DFFX1_HVT \ram_reg[6][39]  ( .D(n1636), .CLK(clk), .Q(\ram[6][39] ) );
  DFFX1_HVT \ram_reg[6][38]  ( .D(n1635), .CLK(clk), .Q(\ram[6][38] ) );
  DFFX1_HVT \ram_reg[6][37]  ( .D(n1634), .CLK(clk), .Q(\ram[6][37] ) );
  DFFX1_HVT \ram_reg[6][36]  ( .D(n1633), .CLK(clk), .Q(\ram[6][36] ) );
  DFFX1_HVT \ram_reg[6][35]  ( .D(n1632), .CLK(clk), .Q(\ram[6][35] ) );
  DFFX1_HVT \ram_reg[6][34]  ( .D(n1631), .CLK(clk), .Q(\ram[6][34] ) );
  DFFX1_HVT \ram_reg[6][33]  ( .D(n1630), .CLK(clk), .Q(\ram[6][33] ) );
  DFFX1_HVT \ram_reg[6][32]  ( .D(n1629), .CLK(clk), .Q(\ram[6][32] ) );
  DFFX1_HVT \ram_reg[6][31]  ( .D(n1628), .CLK(clk), .Q(\ram[6][31] ) );
  DFFX1_HVT \ram_reg[6][30]  ( .D(n1627), .CLK(clk), .Q(\ram[6][30] ) );
  DFFX1_HVT \ram_reg[6][29]  ( .D(n1626), .CLK(clk), .Q(\ram[6][29] ) );
  DFFX1_HVT \ram_reg[6][28]  ( .D(n1625), .CLK(clk), .Q(\ram[6][28] ) );
  DFFX1_HVT \ram_reg[6][27]  ( .D(n1624), .CLK(clk), .Q(\ram[6][27] ) );
  DFFX1_HVT \ram_reg[6][26]  ( .D(n1623), .CLK(clk), .Q(\ram[6][26] ) );
  DFFX1_HVT \ram_reg[6][25]  ( .D(n1622), .CLK(clk), .Q(\ram[6][25] ) );
  DFFX1_HVT \ram_reg[6][24]  ( .D(n1621), .CLK(clk), .Q(\ram[6][24] ) );
  DFFX1_HVT \ram_reg[6][23]  ( .D(n1620), .CLK(clk), .Q(\ram[6][23] ) );
  DFFX1_HVT \ram_reg[6][22]  ( .D(n1619), .CLK(clk), .Q(\ram[6][22] ) );
  DFFX1_HVT \ram_reg[6][21]  ( .D(n1618), .CLK(clk), .Q(\ram[6][21] ) );
  DFFX1_HVT \ram_reg[6][20]  ( .D(n1617), .CLK(clk), .Q(\ram[6][20] ) );
  DFFX1_HVT \ram_reg[6][19]  ( .D(n1616), .CLK(clk), .Q(\ram[6][19] ) );
  DFFX1_HVT \ram_reg[6][18]  ( .D(n1615), .CLK(clk), .Q(\ram[6][18] ) );
  DFFX1_HVT \ram_reg[6][17]  ( .D(n1614), .CLK(clk), .Q(\ram[6][17] ) );
  DFFX1_HVT \ram_reg[6][16]  ( .D(n1613), .CLK(clk), .Q(\ram[6][16] ) );
  DFFX1_HVT \ram_reg[6][15]  ( .D(n1612), .CLK(clk), .Q(\ram[6][15] ) );
  DFFX1_HVT \ram_reg[6][14]  ( .D(n1611), .CLK(clk), .Q(\ram[6][14] ) );
  DFFX1_HVT \ram_reg[6][13]  ( .D(n1610), .CLK(clk), .Q(\ram[6][13] ) );
  DFFX1_HVT \ram_reg[6][12]  ( .D(n1609), .CLK(clk), .Q(\ram[6][12] ) );
  DFFX1_HVT \ram_reg[6][11]  ( .D(n1608), .CLK(clk), .Q(\ram[6][11] ) );
  DFFX1_HVT \ram_reg[6][10]  ( .D(n1607), .CLK(clk), .Q(\ram[6][10] ) );
  DFFX1_HVT \ram_reg[6][9]  ( .D(n1606), .CLK(clk), .Q(\ram[6][9] ) );
  DFFX1_HVT \ram_reg[6][8]  ( .D(n1605), .CLK(clk), .Q(\ram[6][8] ) );
  DFFX1_HVT \ram_reg[6][7]  ( .D(n1604), .CLK(clk), .Q(\ram[6][7] ) );
  DFFX1_HVT \ram_reg[6][6]  ( .D(n1603), .CLK(clk), .Q(\ram[6][6] ) );
  DFFX1_HVT \ram_reg[6][5]  ( .D(n1602), .CLK(clk), .Q(\ram[6][5] ) );
  DFFX1_HVT \ram_reg[6][4]  ( .D(n1601), .CLK(clk), .Q(\ram[6][4] ) );
  DFFX1_HVT \ram_reg[6][3]  ( .D(n1600), .CLK(clk), .Q(\ram[6][3] ) );
  DFFX1_HVT \ram_reg[6][2]  ( .D(n1599), .CLK(clk), .Q(\ram[6][2] ) );
  DFFX1_HVT \ram_reg[6][1]  ( .D(n1598), .CLK(clk), .Q(\ram[6][1] ) );
  DFFX1_HVT \ram_reg[6][0]  ( .D(n1597), .CLK(clk), .Q(\ram[6][0] ) );
  DFFX1_HVT \ram_reg[5][255]  ( .D(n1596), .CLK(clk), .Q(\ram[5][255] ) );
  DFFX1_HVT \ram_reg[5][254]  ( .D(n1595), .CLK(clk), .Q(\ram[5][254] ) );
  DFFX1_HVT \ram_reg[5][253]  ( .D(n1594), .CLK(clk), .Q(\ram[5][253] ) );
  DFFX1_HVT \ram_reg[5][252]  ( .D(n1593), .CLK(clk), .Q(\ram[5][252] ) );
  DFFX1_HVT \ram_reg[5][251]  ( .D(n1592), .CLK(clk), .Q(\ram[5][251] ) );
  DFFX1_HVT \ram_reg[5][250]  ( .D(n1591), .CLK(clk), .Q(\ram[5][250] ) );
  DFFX1_HVT \ram_reg[5][249]  ( .D(n1590), .CLK(clk), .Q(\ram[5][249] ) );
  DFFX1_HVT \ram_reg[5][248]  ( .D(n1589), .CLK(clk), .Q(\ram[5][248] ) );
  DFFX1_HVT \ram_reg[5][247]  ( .D(n1588), .CLK(clk), .Q(\ram[5][247] ) );
  DFFX1_HVT \ram_reg[5][246]  ( .D(n1587), .CLK(clk), .Q(\ram[5][246] ) );
  DFFX1_HVT \ram_reg[5][245]  ( .D(n1586), .CLK(clk), .Q(\ram[5][245] ) );
  DFFX1_HVT \ram_reg[5][244]  ( .D(n1585), .CLK(clk), .Q(\ram[5][244] ) );
  DFFX1_HVT \ram_reg[5][243]  ( .D(n1584), .CLK(clk), .Q(\ram[5][243] ) );
  DFFX1_HVT \ram_reg[5][242]  ( .D(n1583), .CLK(clk), .Q(\ram[5][242] ) );
  DFFX1_HVT \ram_reg[5][241]  ( .D(n1582), .CLK(clk), .Q(\ram[5][241] ) );
  DFFX1_HVT \ram_reg[5][240]  ( .D(n1581), .CLK(clk), .Q(\ram[5][240] ) );
  DFFX1_HVT \ram_reg[5][239]  ( .D(n1580), .CLK(clk), .Q(\ram[5][239] ) );
  DFFX1_HVT \ram_reg[5][238]  ( .D(n1579), .CLK(clk), .Q(\ram[5][238] ) );
  DFFX1_HVT \ram_reg[5][237]  ( .D(n1578), .CLK(clk), .Q(\ram[5][237] ) );
  DFFX1_HVT \ram_reg[5][236]  ( .D(n1577), .CLK(clk), .Q(\ram[5][236] ) );
  DFFX1_HVT \ram_reg[5][235]  ( .D(n1576), .CLK(clk), .Q(\ram[5][235] ) );
  DFFX1_HVT \ram_reg[5][234]  ( .D(n1575), .CLK(clk), .Q(\ram[5][234] ) );
  DFFX1_HVT \ram_reg[5][233]  ( .D(n1574), .CLK(clk), .Q(\ram[5][233] ) );
  DFFX1_HVT \ram_reg[5][232]  ( .D(n1573), .CLK(clk), .Q(\ram[5][232] ) );
  DFFX1_HVT \ram_reg[5][231]  ( .D(n1572), .CLK(clk), .Q(\ram[5][231] ) );
  DFFX1_HVT \ram_reg[5][230]  ( .D(n1571), .CLK(clk), .Q(\ram[5][230] ) );
  DFFX1_HVT \ram_reg[5][229]  ( .D(n1570), .CLK(clk), .Q(\ram[5][229] ) );
  DFFX1_HVT \ram_reg[5][228]  ( .D(n1569), .CLK(clk), .Q(\ram[5][228] ) );
  DFFX1_HVT \ram_reg[5][227]  ( .D(n1568), .CLK(clk), .Q(\ram[5][227] ) );
  DFFX1_HVT \ram_reg[5][226]  ( .D(n1567), .CLK(clk), .Q(\ram[5][226] ) );
  DFFX1_HVT \ram_reg[5][225]  ( .D(n1566), .CLK(clk), .Q(\ram[5][225] ) );
  DFFX1_HVT \ram_reg[5][224]  ( .D(n1565), .CLK(clk), .Q(\ram[5][224] ) );
  DFFX1_HVT \ram_reg[5][223]  ( .D(n1564), .CLK(clk), .Q(\ram[5][223] ) );
  DFFX1_HVT \ram_reg[5][222]  ( .D(n1563), .CLK(clk), .Q(\ram[5][222] ) );
  DFFX1_HVT \ram_reg[5][221]  ( .D(n1562), .CLK(clk), .Q(\ram[5][221] ) );
  DFFX1_HVT \ram_reg[5][220]  ( .D(n1561), .CLK(clk), .Q(\ram[5][220] ) );
  DFFX1_HVT \ram_reg[5][219]  ( .D(n1560), .CLK(clk), .Q(\ram[5][219] ) );
  DFFX1_HVT \ram_reg[5][218]  ( .D(n1559), .CLK(clk), .Q(\ram[5][218] ) );
  DFFX1_HVT \ram_reg[5][217]  ( .D(n1558), .CLK(clk), .Q(\ram[5][217] ) );
  DFFX1_HVT \ram_reg[5][216]  ( .D(n1557), .CLK(clk), .Q(\ram[5][216] ) );
  DFFX1_HVT \ram_reg[5][215]  ( .D(n1556), .CLK(clk), .Q(\ram[5][215] ) );
  DFFX1_HVT \ram_reg[5][214]  ( .D(n1555), .CLK(clk), .Q(\ram[5][214] ) );
  DFFX1_HVT \ram_reg[5][213]  ( .D(n1554), .CLK(clk), .Q(\ram[5][213] ) );
  DFFX1_HVT \ram_reg[5][212]  ( .D(n1553), .CLK(clk), .Q(\ram[5][212] ) );
  DFFX1_HVT \ram_reg[5][211]  ( .D(n1552), .CLK(clk), .Q(\ram[5][211] ) );
  DFFX1_HVT \ram_reg[5][210]  ( .D(n1551), .CLK(clk), .Q(\ram[5][210] ) );
  DFFX1_HVT \ram_reg[5][209]  ( .D(n1550), .CLK(clk), .Q(\ram[5][209] ) );
  DFFX1_HVT \ram_reg[5][208]  ( .D(n1549), .CLK(clk), .Q(\ram[5][208] ) );
  DFFX1_HVT \ram_reg[5][207]  ( .D(n1548), .CLK(clk), .Q(\ram[5][207] ) );
  DFFX1_HVT \ram_reg[5][206]  ( .D(n1547), .CLK(clk), .Q(\ram[5][206] ) );
  DFFX1_HVT \ram_reg[5][205]  ( .D(n1546), .CLK(clk), .Q(\ram[5][205] ) );
  DFFX1_HVT \ram_reg[5][204]  ( .D(n1545), .CLK(clk), .Q(\ram[5][204] ) );
  DFFX1_HVT \ram_reg[5][203]  ( .D(n1544), .CLK(clk), .Q(\ram[5][203] ) );
  DFFX1_HVT \ram_reg[5][202]  ( .D(n1543), .CLK(clk), .Q(\ram[5][202] ) );
  DFFX1_HVT \ram_reg[5][201]  ( .D(n1542), .CLK(clk), .Q(\ram[5][201] ) );
  DFFX1_HVT \ram_reg[5][200]  ( .D(n1541), .CLK(clk), .Q(\ram[5][200] ) );
  DFFX1_HVT \ram_reg[5][199]  ( .D(n1540), .CLK(clk), .Q(\ram[5][199] ) );
  DFFX1_HVT \ram_reg[5][198]  ( .D(n1539), .CLK(clk), .Q(\ram[5][198] ) );
  DFFX1_HVT \ram_reg[5][197]  ( .D(n1538), .CLK(clk), .Q(\ram[5][197] ) );
  DFFX1_HVT \ram_reg[5][196]  ( .D(n1537), .CLK(clk), .Q(\ram[5][196] ) );
  DFFX1_HVT \ram_reg[5][195]  ( .D(n1536), .CLK(clk), .Q(\ram[5][195] ) );
  DFFX1_HVT \ram_reg[5][194]  ( .D(n1535), .CLK(clk), .Q(\ram[5][194] ) );
  DFFX1_HVT \ram_reg[5][193]  ( .D(n1534), .CLK(clk), .Q(\ram[5][193] ) );
  DFFX1_HVT \ram_reg[5][192]  ( .D(n1533), .CLK(clk), .Q(\ram[5][192] ) );
  DFFX1_HVT \ram_reg[5][191]  ( .D(n1532), .CLK(clk), .Q(\ram[5][191] ) );
  DFFX1_HVT \ram_reg[5][190]  ( .D(n1531), .CLK(clk), .Q(\ram[5][190] ) );
  DFFX1_HVT \ram_reg[5][189]  ( .D(n1530), .CLK(clk), .Q(\ram[5][189] ) );
  DFFX1_HVT \ram_reg[5][188]  ( .D(n1529), .CLK(clk), .Q(\ram[5][188] ) );
  DFFX1_HVT \ram_reg[5][187]  ( .D(n1528), .CLK(clk), .Q(\ram[5][187] ) );
  DFFX1_HVT \ram_reg[5][186]  ( .D(n1527), .CLK(clk), .Q(\ram[5][186] ) );
  DFFX1_HVT \ram_reg[5][185]  ( .D(n1526), .CLK(clk), .Q(\ram[5][185] ) );
  DFFX1_HVT \ram_reg[5][184]  ( .D(n1525), .CLK(clk), .Q(\ram[5][184] ) );
  DFFX1_HVT \ram_reg[5][183]  ( .D(n1524), .CLK(clk), .Q(\ram[5][183] ) );
  DFFX1_HVT \ram_reg[5][182]  ( .D(n1523), .CLK(clk), .Q(\ram[5][182] ) );
  DFFX1_HVT \ram_reg[5][181]  ( .D(n1522), .CLK(clk), .Q(\ram[5][181] ) );
  DFFX1_HVT \ram_reg[5][180]  ( .D(n1521), .CLK(clk), .Q(\ram[5][180] ) );
  DFFX1_HVT \ram_reg[5][179]  ( .D(n1520), .CLK(clk), .Q(\ram[5][179] ) );
  DFFX1_HVT \ram_reg[5][178]  ( .D(n1519), .CLK(clk), .Q(\ram[5][178] ) );
  DFFX1_HVT \ram_reg[5][177]  ( .D(n1518), .CLK(clk), .Q(\ram[5][177] ) );
  DFFX1_HVT \ram_reg[5][176]  ( .D(n1517), .CLK(clk), .Q(\ram[5][176] ) );
  DFFX1_HVT \ram_reg[5][175]  ( .D(n1516), .CLK(clk), .Q(\ram[5][175] ) );
  DFFX1_HVT \ram_reg[5][174]  ( .D(n1515), .CLK(clk), .Q(\ram[5][174] ) );
  DFFX1_HVT \ram_reg[5][173]  ( .D(n1514), .CLK(clk), .Q(\ram[5][173] ) );
  DFFX1_HVT \ram_reg[5][172]  ( .D(n1513), .CLK(clk), .Q(\ram[5][172] ) );
  DFFX1_HVT \ram_reg[5][171]  ( .D(n1512), .CLK(clk), .Q(\ram[5][171] ) );
  DFFX1_HVT \ram_reg[5][170]  ( .D(n1511), .CLK(clk), .Q(\ram[5][170] ) );
  DFFX1_HVT \ram_reg[5][169]  ( .D(n1510), .CLK(clk), .Q(\ram[5][169] ) );
  DFFX1_HVT \ram_reg[5][168]  ( .D(n1509), .CLK(clk), .Q(\ram[5][168] ) );
  DFFX1_HVT \ram_reg[5][167]  ( .D(n1508), .CLK(clk), .Q(\ram[5][167] ) );
  DFFX1_HVT \ram_reg[5][166]  ( .D(n1507), .CLK(clk), .Q(\ram[5][166] ) );
  DFFX1_HVT \ram_reg[5][165]  ( .D(n1506), .CLK(clk), .Q(\ram[5][165] ) );
  DFFX1_HVT \ram_reg[5][164]  ( .D(n1505), .CLK(clk), .Q(\ram[5][164] ) );
  DFFX1_HVT \ram_reg[5][163]  ( .D(n1504), .CLK(clk), .Q(\ram[5][163] ) );
  DFFX1_HVT \ram_reg[5][162]  ( .D(n1503), .CLK(clk), .Q(\ram[5][162] ) );
  DFFX1_HVT \ram_reg[5][161]  ( .D(n1502), .CLK(clk), .Q(\ram[5][161] ) );
  DFFX1_HVT \ram_reg[5][160]  ( .D(n1501), .CLK(clk), .Q(\ram[5][160] ) );
  DFFX1_HVT \ram_reg[5][159]  ( .D(n1500), .CLK(clk), .Q(\ram[5][159] ) );
  DFFX1_HVT \ram_reg[5][158]  ( .D(n1499), .CLK(clk), .Q(\ram[5][158] ) );
  DFFX1_HVT \ram_reg[5][157]  ( .D(n1498), .CLK(clk), .Q(\ram[5][157] ) );
  DFFX1_HVT \ram_reg[5][156]  ( .D(n1497), .CLK(clk), .Q(\ram[5][156] ) );
  DFFX1_HVT \ram_reg[5][155]  ( .D(n1496), .CLK(clk), .Q(\ram[5][155] ) );
  DFFX1_HVT \ram_reg[5][154]  ( .D(n1495), .CLK(clk), .Q(\ram[5][154] ) );
  DFFX1_HVT \ram_reg[5][153]  ( .D(n1494), .CLK(clk), .Q(\ram[5][153] ) );
  DFFX1_HVT \ram_reg[5][152]  ( .D(n1493), .CLK(clk), .Q(\ram[5][152] ) );
  DFFX1_HVT \ram_reg[5][151]  ( .D(n1492), .CLK(clk), .Q(\ram[5][151] ) );
  DFFX1_HVT \ram_reg[5][150]  ( .D(n1491), .CLK(clk), .Q(\ram[5][150] ) );
  DFFX1_HVT \ram_reg[5][149]  ( .D(n1490), .CLK(clk), .Q(\ram[5][149] ) );
  DFFX1_HVT \ram_reg[5][148]  ( .D(n1489), .CLK(clk), .Q(\ram[5][148] ) );
  DFFX1_HVT \ram_reg[5][147]  ( .D(n1488), .CLK(clk), .Q(\ram[5][147] ) );
  DFFX1_HVT \ram_reg[5][146]  ( .D(n1487), .CLK(clk), .Q(\ram[5][146] ) );
  DFFX1_HVT \ram_reg[5][145]  ( .D(n1486), .CLK(clk), .Q(\ram[5][145] ) );
  DFFX1_HVT \ram_reg[5][144]  ( .D(n1485), .CLK(clk), .Q(\ram[5][144] ) );
  DFFX1_HVT \ram_reg[5][143]  ( .D(n1484), .CLK(clk), .Q(\ram[5][143] ) );
  DFFX1_HVT \ram_reg[5][142]  ( .D(n1483), .CLK(clk), .Q(\ram[5][142] ) );
  DFFX1_HVT \ram_reg[5][141]  ( .D(n1482), .CLK(clk), .Q(\ram[5][141] ) );
  DFFX1_HVT \ram_reg[5][140]  ( .D(n1481), .CLK(clk), .Q(\ram[5][140] ) );
  DFFX1_HVT \ram_reg[5][139]  ( .D(n1480), .CLK(clk), .Q(\ram[5][139] ) );
  DFFX1_HVT \ram_reg[5][138]  ( .D(n1479), .CLK(clk), .Q(\ram[5][138] ) );
  DFFX1_HVT \ram_reg[5][137]  ( .D(n1478), .CLK(clk), .Q(\ram[5][137] ) );
  DFFX1_HVT \ram_reg[5][136]  ( .D(n1477), .CLK(clk), .Q(\ram[5][136] ) );
  DFFX1_HVT \ram_reg[5][135]  ( .D(n1476), .CLK(clk), .Q(\ram[5][135] ) );
  DFFX1_HVT \ram_reg[5][134]  ( .D(n1475), .CLK(clk), .Q(\ram[5][134] ) );
  DFFX1_HVT \ram_reg[5][133]  ( .D(n1474), .CLK(clk), .Q(\ram[5][133] ) );
  DFFX1_HVT \ram_reg[5][132]  ( .D(n1473), .CLK(clk), .Q(\ram[5][132] ) );
  DFFX1_HVT \ram_reg[5][131]  ( .D(n1472), .CLK(clk), .Q(\ram[5][131] ) );
  DFFX1_HVT \ram_reg[5][130]  ( .D(n1471), .CLK(clk), .Q(\ram[5][130] ) );
  DFFX1_HVT \ram_reg[5][129]  ( .D(n1470), .CLK(clk), .Q(\ram[5][129] ) );
  DFFX1_HVT \ram_reg[5][128]  ( .D(n1469), .CLK(clk), .Q(\ram[5][128] ) );
  DFFX1_HVT \ram_reg[5][127]  ( .D(n1468), .CLK(clk), .Q(\ram[5][127] ) );
  DFFX1_HVT \ram_reg[5][126]  ( .D(n1467), .CLK(clk), .Q(\ram[5][126] ) );
  DFFX1_HVT \ram_reg[5][125]  ( .D(n1466), .CLK(clk), .Q(\ram[5][125] ) );
  DFFX1_HVT \ram_reg[5][124]  ( .D(n1465), .CLK(clk), .Q(\ram[5][124] ) );
  DFFX1_HVT \ram_reg[5][123]  ( .D(n1464), .CLK(clk), .Q(\ram[5][123] ) );
  DFFX1_HVT \ram_reg[5][122]  ( .D(n1463), .CLK(clk), .Q(\ram[5][122] ) );
  DFFX1_HVT \ram_reg[5][121]  ( .D(n1462), .CLK(clk), .Q(\ram[5][121] ) );
  DFFX1_HVT \ram_reg[5][120]  ( .D(n1461), .CLK(clk), .Q(\ram[5][120] ) );
  DFFX1_HVT \ram_reg[5][119]  ( .D(n1460), .CLK(clk), .Q(\ram[5][119] ) );
  DFFX1_HVT \ram_reg[5][118]  ( .D(n1459), .CLK(clk), .Q(\ram[5][118] ) );
  DFFX1_HVT \ram_reg[5][117]  ( .D(n1458), .CLK(clk), .Q(\ram[5][117] ) );
  DFFX1_HVT \ram_reg[5][116]  ( .D(n1457), .CLK(clk), .Q(\ram[5][116] ) );
  DFFX1_HVT \ram_reg[5][115]  ( .D(n1456), .CLK(clk), .Q(\ram[5][115] ) );
  DFFX1_HVT \ram_reg[5][114]  ( .D(n1455), .CLK(clk), .Q(\ram[5][114] ) );
  DFFX1_HVT \ram_reg[5][113]  ( .D(n1454), .CLK(clk), .Q(\ram[5][113] ) );
  DFFX1_HVT \ram_reg[5][112]  ( .D(n1453), .CLK(clk), .Q(\ram[5][112] ) );
  DFFX1_HVT \ram_reg[5][111]  ( .D(n1452), .CLK(clk), .Q(\ram[5][111] ) );
  DFFX1_HVT \ram_reg[5][110]  ( .D(n1451), .CLK(clk), .Q(\ram[5][110] ) );
  DFFX1_HVT \ram_reg[5][109]  ( .D(n1450), .CLK(clk), .Q(\ram[5][109] ) );
  DFFX1_HVT \ram_reg[5][108]  ( .D(n1449), .CLK(clk), .Q(\ram[5][108] ) );
  DFFX1_HVT \ram_reg[5][107]  ( .D(n1448), .CLK(clk), .Q(\ram[5][107] ) );
  DFFX1_HVT \ram_reg[5][106]  ( .D(n1447), .CLK(clk), .Q(\ram[5][106] ) );
  DFFX1_HVT \ram_reg[5][105]  ( .D(n1446), .CLK(clk), .Q(\ram[5][105] ) );
  DFFX1_HVT \ram_reg[5][104]  ( .D(n1445), .CLK(clk), .Q(\ram[5][104] ) );
  DFFX1_HVT \ram_reg[5][103]  ( .D(n1444), .CLK(clk), .Q(\ram[5][103] ) );
  DFFX1_HVT \ram_reg[5][102]  ( .D(n1443), .CLK(clk), .Q(\ram[5][102] ) );
  DFFX1_HVT \ram_reg[5][101]  ( .D(n1442), .CLK(clk), .Q(\ram[5][101] ) );
  DFFX1_HVT \ram_reg[5][100]  ( .D(n1441), .CLK(clk), .Q(\ram[5][100] ) );
  DFFX1_HVT \ram_reg[5][99]  ( .D(n1440), .CLK(clk), .Q(\ram[5][99] ) );
  DFFX1_HVT \ram_reg[5][98]  ( .D(n1439), .CLK(clk), .Q(\ram[5][98] ) );
  DFFX1_HVT \ram_reg[5][97]  ( .D(n1438), .CLK(clk), .Q(\ram[5][97] ) );
  DFFX1_HVT \ram_reg[5][96]  ( .D(n1437), .CLK(clk), .Q(\ram[5][96] ) );
  DFFX1_HVT \ram_reg[5][95]  ( .D(n1436), .CLK(clk), .Q(\ram[5][95] ) );
  DFFX1_HVT \ram_reg[5][94]  ( .D(n1435), .CLK(clk), .Q(\ram[5][94] ) );
  DFFX1_HVT \ram_reg[5][93]  ( .D(n1434), .CLK(clk), .Q(\ram[5][93] ) );
  DFFX1_HVT \ram_reg[5][92]  ( .D(n1433), .CLK(clk), .Q(\ram[5][92] ) );
  DFFX1_HVT \ram_reg[5][91]  ( .D(n1432), .CLK(clk), .Q(\ram[5][91] ) );
  DFFX1_HVT \ram_reg[5][90]  ( .D(n1431), .CLK(clk), .Q(\ram[5][90] ) );
  DFFX1_HVT \ram_reg[5][89]  ( .D(n1430), .CLK(clk), .Q(\ram[5][89] ) );
  DFFX1_HVT \ram_reg[5][88]  ( .D(n1429), .CLK(clk), .Q(\ram[5][88] ) );
  DFFX1_HVT \ram_reg[5][87]  ( .D(n1428), .CLK(clk), .Q(\ram[5][87] ) );
  DFFX1_HVT \ram_reg[5][86]  ( .D(n1427), .CLK(clk), .Q(\ram[5][86] ) );
  DFFX1_HVT \ram_reg[5][85]  ( .D(n1426), .CLK(clk), .Q(\ram[5][85] ) );
  DFFX1_HVT \ram_reg[5][84]  ( .D(n1425), .CLK(clk), .Q(\ram[5][84] ) );
  DFFX1_HVT \ram_reg[5][83]  ( .D(n1424), .CLK(clk), .Q(\ram[5][83] ) );
  DFFX1_HVT \ram_reg[5][82]  ( .D(n1423), .CLK(clk), .Q(\ram[5][82] ) );
  DFFX1_HVT \ram_reg[5][81]  ( .D(n1422), .CLK(clk), .Q(\ram[5][81] ) );
  DFFX1_HVT \ram_reg[5][80]  ( .D(n1421), .CLK(clk), .Q(\ram[5][80] ) );
  DFFX1_HVT \ram_reg[5][79]  ( .D(n1420), .CLK(clk), .Q(\ram[5][79] ) );
  DFFX1_HVT \ram_reg[5][78]  ( .D(n1419), .CLK(clk), .Q(\ram[5][78] ) );
  DFFX1_HVT \ram_reg[5][77]  ( .D(n1418), .CLK(clk), .Q(\ram[5][77] ) );
  DFFX1_HVT \ram_reg[5][76]  ( .D(n1417), .CLK(clk), .Q(\ram[5][76] ) );
  DFFX1_HVT \ram_reg[5][75]  ( .D(n1416), .CLK(clk), .Q(\ram[5][75] ) );
  DFFX1_HVT \ram_reg[5][74]  ( .D(n1415), .CLK(clk), .Q(\ram[5][74] ) );
  DFFX1_HVT \ram_reg[5][73]  ( .D(n1414), .CLK(clk), .Q(\ram[5][73] ) );
  DFFX1_HVT \ram_reg[5][72]  ( .D(n1413), .CLK(clk), .Q(\ram[5][72] ) );
  DFFX1_HVT \ram_reg[5][71]  ( .D(n1412), .CLK(clk), .Q(\ram[5][71] ) );
  DFFX1_HVT \ram_reg[5][70]  ( .D(n1411), .CLK(clk), .Q(\ram[5][70] ) );
  DFFX1_HVT \ram_reg[5][69]  ( .D(n1410), .CLK(clk), .Q(\ram[5][69] ) );
  DFFX1_HVT \ram_reg[5][68]  ( .D(n1409), .CLK(clk), .Q(\ram[5][68] ) );
  DFFX1_HVT \ram_reg[5][67]  ( .D(n1408), .CLK(clk), .Q(\ram[5][67] ) );
  DFFX1_HVT \ram_reg[5][66]  ( .D(n1407), .CLK(clk), .Q(\ram[5][66] ) );
  DFFX1_HVT \ram_reg[5][65]  ( .D(n1406), .CLK(clk), .Q(\ram[5][65] ) );
  DFFX1_HVT \ram_reg[5][64]  ( .D(n1405), .CLK(clk), .Q(\ram[5][64] ) );
  DFFX1_HVT \ram_reg[5][63]  ( .D(n1404), .CLK(clk), .Q(\ram[5][63] ) );
  DFFX1_HVT \ram_reg[5][62]  ( .D(n1403), .CLK(clk), .Q(\ram[5][62] ) );
  DFFX1_HVT \ram_reg[5][61]  ( .D(n1402), .CLK(clk), .Q(\ram[5][61] ) );
  DFFX1_HVT \ram_reg[5][60]  ( .D(n1401), .CLK(clk), .Q(\ram[5][60] ) );
  DFFX1_HVT \ram_reg[5][59]  ( .D(n1400), .CLK(clk), .Q(\ram[5][59] ) );
  DFFX1_HVT \ram_reg[5][58]  ( .D(n1399), .CLK(clk), .Q(\ram[5][58] ) );
  DFFX1_HVT \ram_reg[5][57]  ( .D(n1398), .CLK(clk), .Q(\ram[5][57] ) );
  DFFX1_HVT \ram_reg[5][56]  ( .D(n1397), .CLK(clk), .Q(\ram[5][56] ) );
  DFFX1_HVT \ram_reg[5][55]  ( .D(n1396), .CLK(clk), .Q(\ram[5][55] ) );
  DFFX1_HVT \ram_reg[5][54]  ( .D(n1395), .CLK(clk), .Q(\ram[5][54] ) );
  DFFX1_HVT \ram_reg[5][53]  ( .D(n1394), .CLK(clk), .Q(\ram[5][53] ) );
  DFFX1_HVT \ram_reg[5][52]  ( .D(n1393), .CLK(clk), .Q(\ram[5][52] ) );
  DFFX1_HVT \ram_reg[5][51]  ( .D(n1392), .CLK(clk), .Q(\ram[5][51] ) );
  DFFX1_HVT \ram_reg[5][50]  ( .D(n1391), .CLK(clk), .Q(\ram[5][50] ) );
  DFFX1_HVT \ram_reg[5][49]  ( .D(n1390), .CLK(clk), .Q(\ram[5][49] ) );
  DFFX1_HVT \ram_reg[5][48]  ( .D(n1389), .CLK(clk), .Q(\ram[5][48] ) );
  DFFX1_HVT \ram_reg[5][47]  ( .D(n1388), .CLK(clk), .Q(\ram[5][47] ) );
  DFFX1_HVT \ram_reg[5][46]  ( .D(n1387), .CLK(clk), .Q(\ram[5][46] ) );
  DFFX1_HVT \ram_reg[5][45]  ( .D(n1386), .CLK(clk), .Q(\ram[5][45] ) );
  DFFX1_HVT \ram_reg[5][44]  ( .D(n1385), .CLK(clk), .Q(\ram[5][44] ) );
  DFFX1_HVT \ram_reg[5][43]  ( .D(n1384), .CLK(clk), .Q(\ram[5][43] ) );
  DFFX1_HVT \ram_reg[5][42]  ( .D(n1383), .CLK(clk), .Q(\ram[5][42] ) );
  DFFX1_HVT \ram_reg[5][41]  ( .D(n1382), .CLK(clk), .Q(\ram[5][41] ) );
  DFFX1_HVT \ram_reg[5][40]  ( .D(n1381), .CLK(clk), .Q(\ram[5][40] ) );
  DFFX1_HVT \ram_reg[5][39]  ( .D(n1380), .CLK(clk), .Q(\ram[5][39] ) );
  DFFX1_HVT \ram_reg[5][38]  ( .D(n1379), .CLK(clk), .Q(\ram[5][38] ) );
  DFFX1_HVT \ram_reg[5][37]  ( .D(n1378), .CLK(clk), .Q(\ram[5][37] ) );
  DFFX1_HVT \ram_reg[5][36]  ( .D(n1377), .CLK(clk), .Q(\ram[5][36] ) );
  DFFX1_HVT \ram_reg[5][35]  ( .D(n1376), .CLK(clk), .Q(\ram[5][35] ) );
  DFFX1_HVT \ram_reg[5][34]  ( .D(n1375), .CLK(clk), .Q(\ram[5][34] ) );
  DFFX1_HVT \ram_reg[5][33]  ( .D(n1374), .CLK(clk), .Q(\ram[5][33] ) );
  DFFX1_HVT \ram_reg[5][32]  ( .D(n1373), .CLK(clk), .Q(\ram[5][32] ) );
  DFFX1_HVT \ram_reg[5][31]  ( .D(n1372), .CLK(clk), .Q(\ram[5][31] ) );
  DFFX1_HVT \ram_reg[5][30]  ( .D(n1371), .CLK(clk), .Q(\ram[5][30] ) );
  DFFX1_HVT \ram_reg[5][29]  ( .D(n1370), .CLK(clk), .Q(\ram[5][29] ) );
  DFFX1_HVT \ram_reg[5][28]  ( .D(n1369), .CLK(clk), .Q(\ram[5][28] ) );
  DFFX1_HVT \ram_reg[5][27]  ( .D(n1368), .CLK(clk), .Q(\ram[5][27] ) );
  DFFX1_HVT \ram_reg[5][26]  ( .D(n1367), .CLK(clk), .Q(\ram[5][26] ) );
  DFFX1_HVT \ram_reg[5][25]  ( .D(n1366), .CLK(clk), .Q(\ram[5][25] ) );
  DFFX1_HVT \ram_reg[5][24]  ( .D(n1365), .CLK(clk), .Q(\ram[5][24] ) );
  DFFX1_HVT \ram_reg[5][23]  ( .D(n1364), .CLK(clk), .Q(\ram[5][23] ) );
  DFFX1_HVT \ram_reg[5][22]  ( .D(n1363), .CLK(clk), .Q(\ram[5][22] ) );
  DFFX1_HVT \ram_reg[5][21]  ( .D(n1362), .CLK(clk), .Q(\ram[5][21] ) );
  DFFX1_HVT \ram_reg[5][20]  ( .D(n1361), .CLK(clk), .Q(\ram[5][20] ) );
  DFFX1_HVT \ram_reg[5][19]  ( .D(n1360), .CLK(clk), .Q(\ram[5][19] ) );
  DFFX1_HVT \ram_reg[5][18]  ( .D(n1359), .CLK(clk), .Q(\ram[5][18] ) );
  DFFX1_HVT \ram_reg[5][17]  ( .D(n1358), .CLK(clk), .Q(\ram[5][17] ) );
  DFFX1_HVT \ram_reg[5][16]  ( .D(n1357), .CLK(clk), .Q(\ram[5][16] ) );
  DFFX1_HVT \ram_reg[5][15]  ( .D(n1356), .CLK(clk), .Q(\ram[5][15] ) );
  DFFX1_HVT \ram_reg[5][14]  ( .D(n1355), .CLK(clk), .Q(\ram[5][14] ) );
  DFFX1_HVT \ram_reg[5][13]  ( .D(n1354), .CLK(clk), .Q(\ram[5][13] ) );
  DFFX1_HVT \ram_reg[5][12]  ( .D(n1353), .CLK(clk), .Q(\ram[5][12] ) );
  DFFX1_HVT \ram_reg[5][11]  ( .D(n1352), .CLK(clk), .Q(\ram[5][11] ) );
  DFFX1_HVT \ram_reg[5][10]  ( .D(n1351), .CLK(clk), .Q(\ram[5][10] ) );
  DFFX1_HVT \ram_reg[5][9]  ( .D(n1350), .CLK(clk), .Q(\ram[5][9] ) );
  DFFX1_HVT \ram_reg[5][8]  ( .D(n1349), .CLK(clk), .Q(\ram[5][8] ) );
  DFFX1_HVT \ram_reg[5][7]  ( .D(n1348), .CLK(clk), .Q(\ram[5][7] ) );
  DFFX1_HVT \ram_reg[5][6]  ( .D(n1347), .CLK(clk), .Q(\ram[5][6] ) );
  DFFX1_HVT \ram_reg[5][5]  ( .D(n1346), .CLK(clk), .Q(\ram[5][5] ) );
  DFFX1_HVT \ram_reg[5][4]  ( .D(n1345), .CLK(clk), .Q(\ram[5][4] ) );
  DFFX1_HVT \ram_reg[5][3]  ( .D(n1344), .CLK(clk), .Q(\ram[5][3] ) );
  DFFX1_HVT \ram_reg[5][2]  ( .D(n1343), .CLK(clk), .Q(\ram[5][2] ) );
  DFFX1_HVT \ram_reg[5][1]  ( .D(n1342), .CLK(clk), .Q(\ram[5][1] ) );
  DFFX1_HVT \ram_reg[5][0]  ( .D(n1341), .CLK(clk), .Q(\ram[5][0] ) );
  DFFX1_HVT \ram_reg[4][255]  ( .D(n1340), .CLK(clk), .Q(\ram[4][255] ) );
  DFFX1_HVT \ram_reg[4][254]  ( .D(n1339), .CLK(clk), .Q(\ram[4][254] ) );
  DFFX1_HVT \ram_reg[4][253]  ( .D(n1338), .CLK(clk), .Q(\ram[4][253] ) );
  DFFX1_HVT \ram_reg[4][252]  ( .D(n1337), .CLK(clk), .Q(\ram[4][252] ) );
  DFFX1_HVT \ram_reg[4][251]  ( .D(n1336), .CLK(clk), .Q(\ram[4][251] ) );
  DFFX1_HVT \ram_reg[4][250]  ( .D(n1335), .CLK(clk), .Q(\ram[4][250] ) );
  DFFX1_HVT \ram_reg[4][249]  ( .D(n1334), .CLK(clk), .Q(\ram[4][249] ) );
  DFFX1_HVT \ram_reg[4][248]  ( .D(n1333), .CLK(clk), .Q(\ram[4][248] ) );
  DFFX1_HVT \ram_reg[4][247]  ( .D(n1332), .CLK(clk), .Q(\ram[4][247] ) );
  DFFX1_HVT \ram_reg[4][246]  ( .D(n1331), .CLK(clk), .Q(\ram[4][246] ) );
  DFFX1_HVT \ram_reg[4][245]  ( .D(n1330), .CLK(clk), .Q(\ram[4][245] ) );
  DFFX1_HVT \ram_reg[4][244]  ( .D(n1329), .CLK(clk), .Q(\ram[4][244] ) );
  DFFX1_HVT \ram_reg[4][243]  ( .D(n1328), .CLK(clk), .Q(\ram[4][243] ) );
  DFFX1_HVT \ram_reg[4][242]  ( .D(n1327), .CLK(clk), .Q(\ram[4][242] ) );
  DFFX1_HVT \ram_reg[4][241]  ( .D(n1326), .CLK(clk), .Q(\ram[4][241] ) );
  DFFX1_HVT \ram_reg[4][240]  ( .D(n1325), .CLK(clk), .Q(\ram[4][240] ) );
  DFFX1_HVT \ram_reg[4][239]  ( .D(n1324), .CLK(clk), .Q(\ram[4][239] ) );
  DFFX1_HVT \ram_reg[4][238]  ( .D(n1323), .CLK(clk), .Q(\ram[4][238] ) );
  DFFX1_HVT \ram_reg[4][237]  ( .D(n1322), .CLK(clk), .Q(\ram[4][237] ) );
  DFFX1_HVT \ram_reg[4][236]  ( .D(n1321), .CLK(clk), .Q(\ram[4][236] ) );
  DFFX1_HVT \ram_reg[4][235]  ( .D(n1320), .CLK(clk), .Q(\ram[4][235] ) );
  DFFX1_HVT \ram_reg[4][234]  ( .D(n1319), .CLK(clk), .Q(\ram[4][234] ) );
  DFFX1_HVT \ram_reg[4][233]  ( .D(n1318), .CLK(clk), .Q(\ram[4][233] ) );
  DFFX1_HVT \ram_reg[4][232]  ( .D(n1317), .CLK(clk), .Q(\ram[4][232] ) );
  DFFX1_HVT \ram_reg[4][231]  ( .D(n1316), .CLK(clk), .Q(\ram[4][231] ) );
  DFFX1_HVT \ram_reg[4][230]  ( .D(n1315), .CLK(clk), .Q(\ram[4][230] ) );
  DFFX1_HVT \ram_reg[4][229]  ( .D(n1314), .CLK(clk), .Q(\ram[4][229] ) );
  DFFX1_HVT \ram_reg[4][228]  ( .D(n1313), .CLK(clk), .Q(\ram[4][228] ) );
  DFFX1_HVT \ram_reg[4][227]  ( .D(n1312), .CLK(clk), .Q(\ram[4][227] ) );
  DFFX1_HVT \ram_reg[4][226]  ( .D(n1311), .CLK(clk), .Q(\ram[4][226] ) );
  DFFX1_HVT \ram_reg[4][225]  ( .D(n1310), .CLK(clk), .Q(\ram[4][225] ) );
  DFFX1_HVT \ram_reg[4][224]  ( .D(n1309), .CLK(clk), .Q(\ram[4][224] ) );
  DFFX1_HVT \ram_reg[4][223]  ( .D(n1308), .CLK(clk), .Q(\ram[4][223] ) );
  DFFX1_HVT \ram_reg[4][222]  ( .D(n1307), .CLK(clk), .Q(\ram[4][222] ) );
  DFFX1_HVT \ram_reg[4][221]  ( .D(n1306), .CLK(clk), .Q(\ram[4][221] ) );
  DFFX1_HVT \ram_reg[4][220]  ( .D(n1305), .CLK(clk), .Q(\ram[4][220] ) );
  DFFX1_HVT \ram_reg[4][219]  ( .D(n1304), .CLK(clk), .Q(\ram[4][219] ) );
  DFFX1_HVT \ram_reg[4][218]  ( .D(n1303), .CLK(clk), .Q(\ram[4][218] ) );
  DFFX1_HVT \ram_reg[4][217]  ( .D(n1302), .CLK(clk), .Q(\ram[4][217] ) );
  DFFX1_HVT \ram_reg[4][216]  ( .D(n1301), .CLK(clk), .Q(\ram[4][216] ) );
  DFFX1_HVT \ram_reg[4][215]  ( .D(n1300), .CLK(clk), .Q(\ram[4][215] ) );
  DFFX1_HVT \ram_reg[4][214]  ( .D(n1299), .CLK(clk), .Q(\ram[4][214] ) );
  DFFX1_HVT \ram_reg[4][213]  ( .D(n1298), .CLK(clk), .Q(\ram[4][213] ) );
  DFFX1_HVT \ram_reg[4][212]  ( .D(n1297), .CLK(clk), .Q(\ram[4][212] ) );
  DFFX1_HVT \ram_reg[4][211]  ( .D(n1296), .CLK(clk), .Q(\ram[4][211] ) );
  DFFX1_HVT \ram_reg[4][210]  ( .D(n1295), .CLK(clk), .Q(\ram[4][210] ) );
  DFFX1_HVT \ram_reg[4][209]  ( .D(n1294), .CLK(clk), .Q(\ram[4][209] ) );
  DFFX1_HVT \ram_reg[4][208]  ( .D(n1293), .CLK(clk), .Q(\ram[4][208] ) );
  DFFX1_HVT \ram_reg[4][207]  ( .D(n1292), .CLK(clk), .Q(\ram[4][207] ) );
  DFFX1_HVT \ram_reg[4][206]  ( .D(n1291), .CLK(clk), .Q(\ram[4][206] ) );
  DFFX1_HVT \ram_reg[4][205]  ( .D(n1290), .CLK(clk), .Q(\ram[4][205] ) );
  DFFX1_HVT \ram_reg[4][204]  ( .D(n1289), .CLK(clk), .Q(\ram[4][204] ) );
  DFFX1_HVT \ram_reg[4][203]  ( .D(n1288), .CLK(clk), .Q(\ram[4][203] ) );
  DFFX1_HVT \ram_reg[4][202]  ( .D(n1287), .CLK(clk), .Q(\ram[4][202] ) );
  DFFX1_HVT \ram_reg[4][201]  ( .D(n1286), .CLK(clk), .Q(\ram[4][201] ) );
  DFFX1_HVT \ram_reg[4][200]  ( .D(n1285), .CLK(clk), .Q(\ram[4][200] ) );
  DFFX1_HVT \ram_reg[4][199]  ( .D(n1284), .CLK(clk), .Q(\ram[4][199] ) );
  DFFX1_HVT \ram_reg[4][198]  ( .D(n1283), .CLK(clk), .Q(\ram[4][198] ) );
  DFFX1_HVT \ram_reg[4][197]  ( .D(n1282), .CLK(clk), .Q(\ram[4][197] ) );
  DFFX1_HVT \ram_reg[4][196]  ( .D(n1281), .CLK(clk), .Q(\ram[4][196] ) );
  DFFX1_HVT \ram_reg[4][195]  ( .D(n1280), .CLK(clk), .Q(\ram[4][195] ) );
  DFFX1_HVT \ram_reg[4][194]  ( .D(n1279), .CLK(clk), .Q(\ram[4][194] ) );
  DFFX1_HVT \ram_reg[4][193]  ( .D(n1278), .CLK(clk), .Q(\ram[4][193] ) );
  DFFX1_HVT \ram_reg[4][192]  ( .D(n1277), .CLK(clk), .Q(\ram[4][192] ) );
  DFFX1_HVT \ram_reg[4][191]  ( .D(n1276), .CLK(clk), .Q(\ram[4][191] ) );
  DFFX1_HVT \ram_reg[4][190]  ( .D(n1275), .CLK(clk), .Q(\ram[4][190] ) );
  DFFX1_HVT \ram_reg[4][189]  ( .D(n1274), .CLK(clk), .Q(\ram[4][189] ) );
  DFFX1_HVT \ram_reg[4][188]  ( .D(n1273), .CLK(clk), .Q(\ram[4][188] ) );
  DFFX1_HVT \ram_reg[4][187]  ( .D(n1272), .CLK(clk), .Q(\ram[4][187] ) );
  DFFX1_HVT \ram_reg[4][186]  ( .D(n1271), .CLK(clk), .Q(\ram[4][186] ) );
  DFFX1_HVT \ram_reg[4][185]  ( .D(n1270), .CLK(clk), .Q(\ram[4][185] ) );
  DFFX1_HVT \ram_reg[4][184]  ( .D(n1269), .CLK(clk), .Q(\ram[4][184] ) );
  DFFX1_HVT \ram_reg[4][183]  ( .D(n1268), .CLK(clk), .Q(\ram[4][183] ) );
  DFFX1_HVT \ram_reg[4][182]  ( .D(n1267), .CLK(clk), .Q(\ram[4][182] ) );
  DFFX1_HVT \ram_reg[4][181]  ( .D(n1266), .CLK(clk), .Q(\ram[4][181] ) );
  DFFX1_HVT \ram_reg[4][180]  ( .D(n1265), .CLK(clk), .Q(\ram[4][180] ) );
  DFFX1_HVT \ram_reg[4][179]  ( .D(n1264), .CLK(clk), .Q(\ram[4][179] ) );
  DFFX1_HVT \ram_reg[4][178]  ( .D(n1263), .CLK(clk), .Q(\ram[4][178] ) );
  DFFX1_HVT \ram_reg[4][177]  ( .D(n1262), .CLK(clk), .Q(\ram[4][177] ) );
  DFFX1_HVT \ram_reg[4][176]  ( .D(n1261), .CLK(clk), .Q(\ram[4][176] ) );
  DFFX1_HVT \ram_reg[4][175]  ( .D(n1260), .CLK(clk), .Q(\ram[4][175] ) );
  DFFX1_HVT \ram_reg[4][174]  ( .D(n1259), .CLK(clk), .Q(\ram[4][174] ) );
  DFFX1_HVT \ram_reg[4][173]  ( .D(n1258), .CLK(clk), .Q(\ram[4][173] ) );
  DFFX1_HVT \ram_reg[4][172]  ( .D(n1257), .CLK(clk), .Q(\ram[4][172] ) );
  DFFX1_HVT \ram_reg[4][171]  ( .D(n1256), .CLK(clk), .Q(\ram[4][171] ) );
  DFFX1_HVT \ram_reg[4][170]  ( .D(n1255), .CLK(clk), .Q(\ram[4][170] ) );
  DFFX1_HVT \ram_reg[4][169]  ( .D(n1254), .CLK(clk), .Q(\ram[4][169] ) );
  DFFX1_HVT \ram_reg[4][168]  ( .D(n1253), .CLK(clk), .Q(\ram[4][168] ) );
  DFFX1_HVT \ram_reg[4][167]  ( .D(n1252), .CLK(clk), .Q(\ram[4][167] ) );
  DFFX1_HVT \ram_reg[4][166]  ( .D(n1251), .CLK(clk), .Q(\ram[4][166] ) );
  DFFX1_HVT \ram_reg[4][165]  ( .D(n1250), .CLK(clk), .Q(\ram[4][165] ) );
  DFFX1_HVT \ram_reg[4][164]  ( .D(n1249), .CLK(clk), .Q(\ram[4][164] ) );
  DFFX1_HVT \ram_reg[4][163]  ( .D(n1248), .CLK(clk), .Q(\ram[4][163] ) );
  DFFX1_HVT \ram_reg[4][162]  ( .D(n1247), .CLK(clk), .Q(\ram[4][162] ) );
  DFFX1_HVT \ram_reg[4][161]  ( .D(n1246), .CLK(clk), .Q(\ram[4][161] ) );
  DFFX1_HVT \ram_reg[4][160]  ( .D(n1245), .CLK(clk), .Q(\ram[4][160] ) );
  DFFX1_HVT \ram_reg[4][159]  ( .D(n1244), .CLK(clk), .Q(\ram[4][159] ) );
  DFFX1_HVT \ram_reg[4][158]  ( .D(n1243), .CLK(clk), .Q(\ram[4][158] ) );
  DFFX1_HVT \ram_reg[4][157]  ( .D(n1242), .CLK(clk), .Q(\ram[4][157] ) );
  DFFX1_HVT \ram_reg[4][156]  ( .D(n1241), .CLK(clk), .Q(\ram[4][156] ) );
  DFFX1_HVT \ram_reg[4][155]  ( .D(n1240), .CLK(clk), .Q(\ram[4][155] ) );
  DFFX1_HVT \ram_reg[4][154]  ( .D(n1239), .CLK(clk), .Q(\ram[4][154] ) );
  DFFX1_HVT \ram_reg[4][153]  ( .D(n1238), .CLK(clk), .Q(\ram[4][153] ) );
  DFFX1_HVT \ram_reg[4][152]  ( .D(n1237), .CLK(clk), .Q(\ram[4][152] ) );
  DFFX1_HVT \ram_reg[4][151]  ( .D(n1236), .CLK(clk), .Q(\ram[4][151] ) );
  DFFX1_HVT \ram_reg[4][150]  ( .D(n1235), .CLK(clk), .Q(\ram[4][150] ) );
  DFFX1_HVT \ram_reg[4][149]  ( .D(n1234), .CLK(clk), .Q(\ram[4][149] ) );
  DFFX1_HVT \ram_reg[4][148]  ( .D(n1233), .CLK(clk), .Q(\ram[4][148] ) );
  DFFX1_HVT \ram_reg[4][147]  ( .D(n1232), .CLK(clk), .Q(\ram[4][147] ) );
  DFFX1_HVT \ram_reg[4][146]  ( .D(n1231), .CLK(clk), .Q(\ram[4][146] ) );
  DFFX1_HVT \ram_reg[4][145]  ( .D(n1230), .CLK(clk), .Q(\ram[4][145] ) );
  DFFX1_HVT \ram_reg[4][144]  ( .D(n1229), .CLK(clk), .Q(\ram[4][144] ) );
  DFFX1_HVT \ram_reg[4][143]  ( .D(n1228), .CLK(clk), .Q(\ram[4][143] ) );
  DFFX1_HVT \ram_reg[4][142]  ( .D(n1227), .CLK(clk), .Q(\ram[4][142] ) );
  DFFX1_HVT \ram_reg[4][141]  ( .D(n1226), .CLK(clk), .Q(\ram[4][141] ) );
  DFFX1_HVT \ram_reg[4][140]  ( .D(n1225), .CLK(clk), .Q(\ram[4][140] ) );
  DFFX1_HVT \ram_reg[4][139]  ( .D(n1224), .CLK(clk), .Q(\ram[4][139] ) );
  DFFX1_HVT \ram_reg[4][138]  ( .D(n1223), .CLK(clk), .Q(\ram[4][138] ) );
  DFFX1_HVT \ram_reg[4][137]  ( .D(n1222), .CLK(clk), .Q(\ram[4][137] ) );
  DFFX1_HVT \ram_reg[4][136]  ( .D(n1221), .CLK(clk), .Q(\ram[4][136] ) );
  DFFX1_HVT \ram_reg[4][135]  ( .D(n1220), .CLK(clk), .Q(\ram[4][135] ) );
  DFFX1_HVT \ram_reg[4][134]  ( .D(n1219), .CLK(clk), .Q(\ram[4][134] ) );
  DFFX1_HVT \ram_reg[4][133]  ( .D(n1218), .CLK(clk), .Q(\ram[4][133] ) );
  DFFX1_HVT \ram_reg[4][132]  ( .D(n1217), .CLK(clk), .Q(\ram[4][132] ) );
  DFFX1_HVT \ram_reg[4][131]  ( .D(n1216), .CLK(clk), .Q(\ram[4][131] ) );
  DFFX1_HVT \ram_reg[4][130]  ( .D(n1215), .CLK(clk), .Q(\ram[4][130] ) );
  DFFX1_HVT \ram_reg[4][129]  ( .D(n1214), .CLK(clk), .Q(\ram[4][129] ) );
  DFFX1_HVT \ram_reg[4][128]  ( .D(n1213), .CLK(clk), .Q(\ram[4][128] ) );
  DFFX1_HVT \ram_reg[4][127]  ( .D(n1212), .CLK(clk), .Q(\ram[4][127] ) );
  DFFX1_HVT \ram_reg[4][126]  ( .D(n1211), .CLK(clk), .Q(\ram[4][126] ) );
  DFFX1_HVT \ram_reg[4][125]  ( .D(n1210), .CLK(clk), .Q(\ram[4][125] ) );
  DFFX1_HVT \ram_reg[4][124]  ( .D(n1209), .CLK(clk), .Q(\ram[4][124] ) );
  DFFX1_HVT \ram_reg[4][123]  ( .D(n1208), .CLK(clk), .Q(\ram[4][123] ) );
  DFFX1_HVT \ram_reg[4][122]  ( .D(n1207), .CLK(clk), .Q(\ram[4][122] ) );
  DFFX1_HVT \ram_reg[4][121]  ( .D(n1206), .CLK(clk), .Q(\ram[4][121] ) );
  DFFX1_HVT \ram_reg[4][120]  ( .D(n1205), .CLK(clk), .Q(\ram[4][120] ) );
  DFFX1_HVT \ram_reg[4][119]  ( .D(n1204), .CLK(clk), .Q(\ram[4][119] ) );
  DFFX1_HVT \ram_reg[4][118]  ( .D(n1203), .CLK(clk), .Q(\ram[4][118] ) );
  DFFX1_HVT \ram_reg[4][117]  ( .D(n1202), .CLK(clk), .Q(\ram[4][117] ) );
  DFFX1_HVT \ram_reg[4][116]  ( .D(n1201), .CLK(clk), .Q(\ram[4][116] ) );
  DFFX1_HVT \ram_reg[4][115]  ( .D(n1200), .CLK(clk), .Q(\ram[4][115] ) );
  DFFX1_HVT \ram_reg[4][114]  ( .D(n1199), .CLK(clk), .Q(\ram[4][114] ) );
  DFFX1_HVT \ram_reg[4][113]  ( .D(n1198), .CLK(clk), .Q(\ram[4][113] ) );
  DFFX1_HVT \ram_reg[4][112]  ( .D(n1197), .CLK(clk), .Q(\ram[4][112] ) );
  DFFX1_HVT \ram_reg[4][111]  ( .D(n1196), .CLK(clk), .Q(\ram[4][111] ) );
  DFFX1_HVT \ram_reg[4][110]  ( .D(n1195), .CLK(clk), .Q(\ram[4][110] ) );
  DFFX1_HVT \ram_reg[4][109]  ( .D(n1194), .CLK(clk), .Q(\ram[4][109] ) );
  DFFX1_HVT \ram_reg[4][108]  ( .D(n1193), .CLK(clk), .Q(\ram[4][108] ) );
  DFFX1_HVT \ram_reg[4][107]  ( .D(n1192), .CLK(clk), .Q(\ram[4][107] ) );
  DFFX1_HVT \ram_reg[4][106]  ( .D(n1191), .CLK(clk), .Q(\ram[4][106] ) );
  DFFX1_HVT \ram_reg[4][105]  ( .D(n1190), .CLK(clk), .Q(\ram[4][105] ) );
  DFFX1_HVT \ram_reg[4][104]  ( .D(n1189), .CLK(clk), .Q(\ram[4][104] ) );
  DFFX1_HVT \ram_reg[4][103]  ( .D(n1188), .CLK(clk), .Q(\ram[4][103] ) );
  DFFX1_HVT \ram_reg[4][102]  ( .D(n1187), .CLK(clk), .Q(\ram[4][102] ) );
  DFFX1_HVT \ram_reg[4][101]  ( .D(n1186), .CLK(clk), .Q(\ram[4][101] ) );
  DFFX1_HVT \ram_reg[4][100]  ( .D(n1185), .CLK(clk), .Q(\ram[4][100] ) );
  DFFX1_HVT \ram_reg[4][99]  ( .D(n1184), .CLK(clk), .Q(\ram[4][99] ) );
  DFFX1_HVT \ram_reg[4][98]  ( .D(n1183), .CLK(clk), .Q(\ram[4][98] ) );
  DFFX1_HVT \ram_reg[4][97]  ( .D(n1182), .CLK(clk), .Q(\ram[4][97] ) );
  DFFX1_HVT \ram_reg[4][96]  ( .D(n1181), .CLK(clk), .Q(\ram[4][96] ) );
  DFFX1_HVT \ram_reg[4][95]  ( .D(n1180), .CLK(clk), .Q(\ram[4][95] ) );
  DFFX1_HVT \ram_reg[4][94]  ( .D(n1179), .CLK(clk), .Q(\ram[4][94] ) );
  DFFX1_HVT \ram_reg[4][93]  ( .D(n1178), .CLK(clk), .Q(\ram[4][93] ) );
  DFFX1_HVT \ram_reg[4][92]  ( .D(n1177), .CLK(clk), .Q(\ram[4][92] ) );
  DFFX1_HVT \ram_reg[4][91]  ( .D(n1176), .CLK(clk), .Q(\ram[4][91] ) );
  DFFX1_HVT \ram_reg[4][90]  ( .D(n1175), .CLK(clk), .Q(\ram[4][90] ) );
  DFFX1_HVT \ram_reg[4][89]  ( .D(n1174), .CLK(clk), .Q(\ram[4][89] ) );
  DFFX1_HVT \ram_reg[4][88]  ( .D(n1173), .CLK(clk), .Q(\ram[4][88] ) );
  DFFX1_HVT \ram_reg[4][87]  ( .D(n1172), .CLK(clk), .Q(\ram[4][87] ) );
  DFFX1_HVT \ram_reg[4][86]  ( .D(n1171), .CLK(clk), .Q(\ram[4][86] ) );
  DFFX1_HVT \ram_reg[4][85]  ( .D(n1170), .CLK(clk), .Q(\ram[4][85] ) );
  DFFX1_HVT \ram_reg[4][84]  ( .D(n1169), .CLK(clk), .Q(\ram[4][84] ) );
  DFFX1_HVT \ram_reg[4][83]  ( .D(n1168), .CLK(clk), .Q(\ram[4][83] ) );
  DFFX1_HVT \ram_reg[4][82]  ( .D(n1167), .CLK(clk), .Q(\ram[4][82] ) );
  DFFX1_HVT \ram_reg[4][81]  ( .D(n1166), .CLK(clk), .Q(\ram[4][81] ) );
  DFFX1_HVT \ram_reg[4][80]  ( .D(n1165), .CLK(clk), .Q(\ram[4][80] ) );
  DFFX1_HVT \ram_reg[4][79]  ( .D(n1164), .CLK(clk), .Q(\ram[4][79] ) );
  DFFX1_HVT \ram_reg[4][78]  ( .D(n1163), .CLK(clk), .Q(\ram[4][78] ) );
  DFFX1_HVT \ram_reg[4][77]  ( .D(n1162), .CLK(clk), .Q(\ram[4][77] ) );
  DFFX1_HVT \ram_reg[4][76]  ( .D(n1161), .CLK(clk), .Q(\ram[4][76] ) );
  DFFX1_HVT \ram_reg[4][75]  ( .D(n1160), .CLK(clk), .Q(\ram[4][75] ) );
  DFFX1_HVT \ram_reg[4][74]  ( .D(n1159), .CLK(clk), .Q(\ram[4][74] ) );
  DFFX1_HVT \ram_reg[4][73]  ( .D(n1158), .CLK(clk), .Q(\ram[4][73] ) );
  DFFX1_HVT \ram_reg[4][72]  ( .D(n1157), .CLK(clk), .Q(\ram[4][72] ) );
  DFFX1_HVT \ram_reg[4][71]  ( .D(n1156), .CLK(clk), .Q(\ram[4][71] ) );
  DFFX1_HVT \ram_reg[4][70]  ( .D(n1155), .CLK(clk), .Q(\ram[4][70] ) );
  DFFX1_HVT \ram_reg[4][69]  ( .D(n1154), .CLK(clk), .Q(\ram[4][69] ) );
  DFFX1_HVT \ram_reg[4][68]  ( .D(n1153), .CLK(clk), .Q(\ram[4][68] ) );
  DFFX1_HVT \ram_reg[4][67]  ( .D(n1152), .CLK(clk), .Q(\ram[4][67] ) );
  DFFX1_HVT \ram_reg[4][66]  ( .D(n1151), .CLK(clk), .Q(\ram[4][66] ) );
  DFFX1_HVT \ram_reg[4][65]  ( .D(n1150), .CLK(clk), .Q(\ram[4][65] ) );
  DFFX1_HVT \ram_reg[4][64]  ( .D(n1149), .CLK(clk), .Q(\ram[4][64] ) );
  DFFX1_HVT \ram_reg[4][63]  ( .D(n1148), .CLK(clk), .Q(\ram[4][63] ) );
  DFFX1_HVT \ram_reg[4][62]  ( .D(n1147), .CLK(clk), .Q(\ram[4][62] ) );
  DFFX1_HVT \ram_reg[4][61]  ( .D(n1146), .CLK(clk), .Q(\ram[4][61] ) );
  DFFX1_HVT \ram_reg[4][60]  ( .D(n1145), .CLK(clk), .Q(\ram[4][60] ) );
  DFFX1_HVT \ram_reg[4][59]  ( .D(n1144), .CLK(clk), .Q(\ram[4][59] ) );
  DFFX1_HVT \ram_reg[4][58]  ( .D(n1143), .CLK(clk), .Q(\ram[4][58] ) );
  DFFX1_HVT \ram_reg[4][57]  ( .D(n1142), .CLK(clk), .Q(\ram[4][57] ) );
  DFFX1_HVT \ram_reg[4][56]  ( .D(n1141), .CLK(clk), .Q(\ram[4][56] ) );
  DFFX1_HVT \ram_reg[4][55]  ( .D(n1140), .CLK(clk), .Q(\ram[4][55] ) );
  DFFX1_HVT \ram_reg[4][54]  ( .D(n1139), .CLK(clk), .Q(\ram[4][54] ) );
  DFFX1_HVT \ram_reg[4][53]  ( .D(n1138), .CLK(clk), .Q(\ram[4][53] ) );
  DFFX1_HVT \ram_reg[4][52]  ( .D(n1137), .CLK(clk), .Q(\ram[4][52] ) );
  DFFX1_HVT \ram_reg[4][51]  ( .D(n1136), .CLK(clk), .Q(\ram[4][51] ) );
  DFFX1_HVT \ram_reg[4][50]  ( .D(n1135), .CLK(clk), .Q(\ram[4][50] ) );
  DFFX1_HVT \ram_reg[4][49]  ( .D(n1134), .CLK(clk), .Q(\ram[4][49] ) );
  DFFX1_HVT \ram_reg[4][48]  ( .D(n1133), .CLK(clk), .Q(\ram[4][48] ) );
  DFFX1_HVT \ram_reg[4][47]  ( .D(n1132), .CLK(clk), .Q(\ram[4][47] ) );
  DFFX1_HVT \ram_reg[4][46]  ( .D(n1131), .CLK(clk), .Q(\ram[4][46] ) );
  DFFX1_HVT \ram_reg[4][45]  ( .D(n1130), .CLK(clk), .Q(\ram[4][45] ) );
  DFFX1_HVT \ram_reg[4][44]  ( .D(n1129), .CLK(clk), .Q(\ram[4][44] ) );
  DFFX1_HVT \ram_reg[4][43]  ( .D(n1128), .CLK(clk), .Q(\ram[4][43] ) );
  DFFX1_HVT \ram_reg[4][42]  ( .D(n1127), .CLK(clk), .Q(\ram[4][42] ) );
  DFFX1_HVT \ram_reg[4][41]  ( .D(n1126), .CLK(clk), .Q(\ram[4][41] ) );
  DFFX1_HVT \ram_reg[4][40]  ( .D(n1125), .CLK(clk), .Q(\ram[4][40] ) );
  DFFX1_HVT \ram_reg[4][39]  ( .D(n1124), .CLK(clk), .Q(\ram[4][39] ) );
  DFFX1_HVT \ram_reg[4][38]  ( .D(n1123), .CLK(clk), .Q(\ram[4][38] ) );
  DFFX1_HVT \ram_reg[4][37]  ( .D(n1122), .CLK(clk), .Q(\ram[4][37] ) );
  DFFX1_HVT \ram_reg[4][36]  ( .D(n1121), .CLK(clk), .Q(\ram[4][36] ) );
  DFFX1_HVT \ram_reg[4][35]  ( .D(n1120), .CLK(clk), .Q(\ram[4][35] ) );
  DFFX1_HVT \ram_reg[4][34]  ( .D(n1119), .CLK(clk), .Q(\ram[4][34] ) );
  DFFX1_HVT \ram_reg[4][33]  ( .D(n1118), .CLK(clk), .Q(\ram[4][33] ) );
  DFFX1_HVT \ram_reg[4][32]  ( .D(n1117), .CLK(clk), .Q(\ram[4][32] ) );
  DFFX1_HVT \ram_reg[4][31]  ( .D(n1116), .CLK(clk), .Q(\ram[4][31] ) );
  DFFX1_HVT \ram_reg[4][30]  ( .D(n1115), .CLK(clk), .Q(\ram[4][30] ) );
  DFFX1_HVT \ram_reg[4][29]  ( .D(n1114), .CLK(clk), .Q(\ram[4][29] ) );
  DFFX1_HVT \ram_reg[4][28]  ( .D(n1113), .CLK(clk), .Q(\ram[4][28] ) );
  DFFX1_HVT \ram_reg[4][27]  ( .D(n1112), .CLK(clk), .Q(\ram[4][27] ) );
  DFFX1_HVT \ram_reg[4][26]  ( .D(n1111), .CLK(clk), .Q(\ram[4][26] ) );
  DFFX1_HVT \ram_reg[4][25]  ( .D(n1110), .CLK(clk), .Q(\ram[4][25] ) );
  DFFX1_HVT \ram_reg[4][24]  ( .D(n1109), .CLK(clk), .Q(\ram[4][24] ) );
  DFFX1_HVT \ram_reg[4][23]  ( .D(n1108), .CLK(clk), .Q(\ram[4][23] ) );
  DFFX1_HVT \ram_reg[4][22]  ( .D(n1107), .CLK(clk), .Q(\ram[4][22] ) );
  DFFX1_HVT \ram_reg[4][21]  ( .D(n1106), .CLK(clk), .Q(\ram[4][21] ) );
  DFFX1_HVT \ram_reg[4][20]  ( .D(n1105), .CLK(clk), .Q(\ram[4][20] ) );
  DFFX1_HVT \ram_reg[4][19]  ( .D(n1104), .CLK(clk), .Q(\ram[4][19] ) );
  DFFX1_HVT \ram_reg[4][18]  ( .D(n1103), .CLK(clk), .Q(\ram[4][18] ) );
  DFFX1_HVT \ram_reg[4][17]  ( .D(n1102), .CLK(clk), .Q(\ram[4][17] ) );
  DFFX1_HVT \ram_reg[4][16]  ( .D(n1101), .CLK(clk), .Q(\ram[4][16] ) );
  DFFX1_HVT \ram_reg[4][15]  ( .D(n1100), .CLK(clk), .Q(\ram[4][15] ) );
  DFFX1_HVT \ram_reg[4][14]  ( .D(n1099), .CLK(clk), .Q(\ram[4][14] ) );
  DFFX1_HVT \ram_reg[4][13]  ( .D(n1098), .CLK(clk), .Q(\ram[4][13] ) );
  DFFX1_HVT \ram_reg[4][12]  ( .D(n1097), .CLK(clk), .Q(\ram[4][12] ) );
  DFFX1_HVT \ram_reg[4][11]  ( .D(n1096), .CLK(clk), .Q(\ram[4][11] ) );
  DFFX1_HVT \ram_reg[4][10]  ( .D(n1095), .CLK(clk), .Q(\ram[4][10] ) );
  DFFX1_HVT \ram_reg[4][9]  ( .D(n1094), .CLK(clk), .Q(\ram[4][9] ) );
  DFFX1_HVT \ram_reg[4][8]  ( .D(n1093), .CLK(clk), .Q(\ram[4][8] ) );
  DFFX1_HVT \ram_reg[4][7]  ( .D(n1092), .CLK(clk), .Q(\ram[4][7] ) );
  DFFX1_HVT \ram_reg[4][6]  ( .D(n1091), .CLK(clk), .Q(\ram[4][6] ) );
  DFFX1_HVT \ram_reg[4][5]  ( .D(n1090), .CLK(clk), .Q(\ram[4][5] ) );
  DFFX1_HVT \ram_reg[4][4]  ( .D(n1089), .CLK(clk), .Q(\ram[4][4] ) );
  DFFX1_HVT \ram_reg[4][3]  ( .D(n1088), .CLK(clk), .Q(\ram[4][3] ) );
  DFFX1_HVT \ram_reg[4][2]  ( .D(n1087), .CLK(clk), .Q(\ram[4][2] ) );
  DFFX1_HVT \ram_reg[4][1]  ( .D(n1086), .CLK(clk), .Q(\ram[4][1] ) );
  DFFX1_HVT \ram_reg[4][0]  ( .D(n1085), .CLK(clk), .Q(\ram[4][0] ) );
  DFFX1_HVT \ram_reg[3][255]  ( .D(n1084), .CLK(clk), .Q(\ram[3][255] ) );
  DFFX1_HVT \ram_reg[3][254]  ( .D(n1083), .CLK(clk), .Q(\ram[3][254] ) );
  DFFX1_HVT \ram_reg[3][253]  ( .D(n1082), .CLK(clk), .Q(\ram[3][253] ) );
  DFFX1_HVT \ram_reg[3][252]  ( .D(n1081), .CLK(clk), .Q(\ram[3][252] ) );
  DFFX1_HVT \ram_reg[3][251]  ( .D(n1080), .CLK(clk), .Q(\ram[3][251] ) );
  DFFX1_HVT \ram_reg[3][250]  ( .D(n1079), .CLK(clk), .Q(\ram[3][250] ) );
  DFFX1_HVT \ram_reg[3][249]  ( .D(n1078), .CLK(clk), .Q(\ram[3][249] ) );
  DFFX1_HVT \ram_reg[3][248]  ( .D(n1077), .CLK(clk), .Q(\ram[3][248] ) );
  DFFX1_HVT \ram_reg[3][247]  ( .D(n1076), .CLK(clk), .Q(\ram[3][247] ) );
  DFFX1_HVT \ram_reg[3][246]  ( .D(n1075), .CLK(clk), .Q(\ram[3][246] ) );
  DFFX1_HVT \ram_reg[3][245]  ( .D(n1074), .CLK(clk), .Q(\ram[3][245] ) );
  DFFX1_HVT \ram_reg[3][244]  ( .D(n1073), .CLK(clk), .Q(\ram[3][244] ) );
  DFFX1_HVT \ram_reg[3][243]  ( .D(n1072), .CLK(clk), .Q(\ram[3][243] ) );
  DFFX1_HVT \ram_reg[3][242]  ( .D(n1071), .CLK(clk), .Q(\ram[3][242] ) );
  DFFX1_HVT \ram_reg[3][241]  ( .D(n1070), .CLK(clk), .Q(\ram[3][241] ) );
  DFFX1_HVT \ram_reg[3][240]  ( .D(n1069), .CLK(clk), .Q(\ram[3][240] ) );
  DFFX1_HVT \ram_reg[3][239]  ( .D(n1068), .CLK(clk), .Q(\ram[3][239] ) );
  DFFX1_HVT \ram_reg[3][238]  ( .D(n1067), .CLK(clk), .Q(\ram[3][238] ) );
  DFFX1_HVT \ram_reg[3][237]  ( .D(n1066), .CLK(clk), .Q(\ram[3][237] ) );
  DFFX1_HVT \ram_reg[3][236]  ( .D(n1065), .CLK(clk), .Q(\ram[3][236] ) );
  DFFX1_HVT \ram_reg[3][235]  ( .D(n1064), .CLK(clk), .Q(\ram[3][235] ) );
  DFFX1_HVT \ram_reg[3][234]  ( .D(n1063), .CLK(clk), .Q(\ram[3][234] ) );
  DFFX1_HVT \ram_reg[3][233]  ( .D(n1062), .CLK(clk), .Q(\ram[3][233] ) );
  DFFX1_HVT \ram_reg[3][232]  ( .D(n1061), .CLK(clk), .Q(\ram[3][232] ) );
  DFFX1_HVT \ram_reg[3][231]  ( .D(n1060), .CLK(clk), .Q(\ram[3][231] ) );
  DFFX1_HVT \ram_reg[3][230]  ( .D(n1059), .CLK(clk), .Q(\ram[3][230] ) );
  DFFX1_HVT \ram_reg[3][229]  ( .D(n1058), .CLK(clk), .Q(\ram[3][229] ) );
  DFFX1_HVT \ram_reg[3][228]  ( .D(n1057), .CLK(clk), .Q(\ram[3][228] ) );
  DFFX1_HVT \ram_reg[3][227]  ( .D(n1056), .CLK(clk), .Q(\ram[3][227] ) );
  DFFX1_HVT \ram_reg[3][226]  ( .D(n1055), .CLK(clk), .Q(\ram[3][226] ) );
  DFFX1_HVT \ram_reg[3][225]  ( .D(n1054), .CLK(clk), .Q(\ram[3][225] ) );
  DFFX1_HVT \ram_reg[3][224]  ( .D(n1053), .CLK(clk), .Q(\ram[3][224] ) );
  DFFX1_HVT \ram_reg[3][223]  ( .D(n1052), .CLK(clk), .Q(\ram[3][223] ) );
  DFFX1_HVT \ram_reg[3][222]  ( .D(n1051), .CLK(clk), .Q(\ram[3][222] ) );
  DFFX1_HVT \ram_reg[3][221]  ( .D(n1050), .CLK(clk), .Q(\ram[3][221] ) );
  DFFX1_HVT \ram_reg[3][220]  ( .D(n1049), .CLK(clk), .Q(\ram[3][220] ) );
  DFFX1_HVT \ram_reg[3][219]  ( .D(n1048), .CLK(clk), .Q(\ram[3][219] ) );
  DFFX1_HVT \ram_reg[3][218]  ( .D(n1047), .CLK(clk), .Q(\ram[3][218] ) );
  DFFX1_HVT \ram_reg[3][217]  ( .D(n1046), .CLK(clk), .Q(\ram[3][217] ) );
  DFFX1_HVT \ram_reg[3][216]  ( .D(n1045), .CLK(clk), .Q(\ram[3][216] ) );
  DFFX1_HVT \ram_reg[3][215]  ( .D(n1044), .CLK(clk), .Q(\ram[3][215] ) );
  DFFX1_HVT \ram_reg[3][214]  ( .D(n1043), .CLK(clk), .Q(\ram[3][214] ) );
  DFFX1_HVT \ram_reg[3][213]  ( .D(n1042), .CLK(clk), .Q(\ram[3][213] ) );
  DFFX1_HVT \ram_reg[3][212]  ( .D(n1041), .CLK(clk), .Q(\ram[3][212] ) );
  DFFX1_HVT \ram_reg[3][211]  ( .D(n1040), .CLK(clk), .Q(\ram[3][211] ) );
  DFFX1_HVT \ram_reg[3][210]  ( .D(n1039), .CLK(clk), .Q(\ram[3][210] ) );
  DFFX1_HVT \ram_reg[3][209]  ( .D(n1038), .CLK(clk), .Q(\ram[3][209] ) );
  DFFX1_HVT \ram_reg[3][208]  ( .D(n1037), .CLK(clk), .Q(\ram[3][208] ) );
  DFFX1_HVT \ram_reg[3][207]  ( .D(n1036), .CLK(clk), .Q(\ram[3][207] ) );
  DFFX1_HVT \ram_reg[3][206]  ( .D(n1035), .CLK(clk), .Q(\ram[3][206] ) );
  DFFX1_HVT \ram_reg[3][205]  ( .D(n1034), .CLK(clk), .Q(\ram[3][205] ) );
  DFFX1_HVT \ram_reg[3][204]  ( .D(n1033), .CLK(clk), .Q(\ram[3][204] ) );
  DFFX1_HVT \ram_reg[3][203]  ( .D(n1032), .CLK(clk), .Q(\ram[3][203] ) );
  DFFX1_HVT \ram_reg[3][202]  ( .D(n1031), .CLK(clk), .Q(\ram[3][202] ) );
  DFFX1_HVT \ram_reg[3][201]  ( .D(n1030), .CLK(clk), .Q(\ram[3][201] ) );
  DFFX1_HVT \ram_reg[3][200]  ( .D(n1029), .CLK(clk), .Q(\ram[3][200] ) );
  DFFX1_HVT \ram_reg[3][199]  ( .D(n1028), .CLK(clk), .Q(\ram[3][199] ) );
  DFFX1_HVT \ram_reg[3][198]  ( .D(n1027), .CLK(clk), .Q(\ram[3][198] ) );
  DFFX1_HVT \ram_reg[3][197]  ( .D(n1026), .CLK(clk), .Q(\ram[3][197] ) );
  DFFX1_HVT \ram_reg[3][196]  ( .D(n1025), .CLK(clk), .Q(\ram[3][196] ) );
  DFFX1_HVT \ram_reg[3][195]  ( .D(n1024), .CLK(clk), .Q(\ram[3][195] ) );
  DFFX1_HVT \ram_reg[3][194]  ( .D(n1023), .CLK(clk), .Q(\ram[3][194] ) );
  DFFX1_HVT \ram_reg[3][193]  ( .D(n1022), .CLK(clk), .Q(\ram[3][193] ) );
  DFFX1_HVT \ram_reg[3][192]  ( .D(n1021), .CLK(clk), .Q(\ram[3][192] ) );
  DFFX1_HVT \ram_reg[3][191]  ( .D(n1020), .CLK(clk), .Q(\ram[3][191] ) );
  DFFX1_HVT \ram_reg[3][190]  ( .D(n1019), .CLK(clk), .Q(\ram[3][190] ) );
  DFFX1_HVT \ram_reg[3][189]  ( .D(n1018), .CLK(clk), .Q(\ram[3][189] ) );
  DFFX1_HVT \ram_reg[3][188]  ( .D(n1017), .CLK(clk), .Q(\ram[3][188] ) );
  DFFX1_HVT \ram_reg[3][187]  ( .D(n1016), .CLK(clk), .Q(\ram[3][187] ) );
  DFFX1_HVT \ram_reg[3][186]  ( .D(n1015), .CLK(clk), .Q(\ram[3][186] ) );
  DFFX1_HVT \ram_reg[3][185]  ( .D(n1014), .CLK(clk), .Q(\ram[3][185] ) );
  DFFX1_HVT \ram_reg[3][184]  ( .D(n1013), .CLK(clk), .Q(\ram[3][184] ) );
  DFFX1_HVT \ram_reg[3][183]  ( .D(n1012), .CLK(clk), .Q(\ram[3][183] ) );
  DFFX1_HVT \ram_reg[3][182]  ( .D(n1011), .CLK(clk), .Q(\ram[3][182] ) );
  DFFX1_HVT \ram_reg[3][181]  ( .D(n1010), .CLK(clk), .Q(\ram[3][181] ) );
  DFFX1_HVT \ram_reg[3][180]  ( .D(n1009), .CLK(clk), .Q(\ram[3][180] ) );
  DFFX1_HVT \ram_reg[3][179]  ( .D(n1008), .CLK(clk), .Q(\ram[3][179] ) );
  DFFX1_HVT \ram_reg[3][178]  ( .D(n1007), .CLK(clk), .Q(\ram[3][178] ) );
  DFFX1_HVT \ram_reg[3][177]  ( .D(n1006), .CLK(clk), .Q(\ram[3][177] ) );
  DFFX1_HVT \ram_reg[3][176]  ( .D(n1005), .CLK(clk), .Q(\ram[3][176] ) );
  DFFX1_HVT \ram_reg[3][175]  ( .D(n1004), .CLK(clk), .Q(\ram[3][175] ) );
  DFFX1_HVT \ram_reg[3][174]  ( .D(n1003), .CLK(clk), .Q(\ram[3][174] ) );
  DFFX1_HVT \ram_reg[3][173]  ( .D(n1002), .CLK(clk), .Q(\ram[3][173] ) );
  DFFX1_HVT \ram_reg[3][172]  ( .D(n1001), .CLK(clk), .Q(\ram[3][172] ) );
  DFFX1_HVT \ram_reg[3][171]  ( .D(n1000), .CLK(clk), .Q(\ram[3][171] ) );
  DFFX1_HVT \ram_reg[3][170]  ( .D(n999), .CLK(clk), .Q(\ram[3][170] ) );
  DFFX1_HVT \ram_reg[3][169]  ( .D(n998), .CLK(clk), .Q(\ram[3][169] ) );
  DFFX1_HVT \ram_reg[3][168]  ( .D(n997), .CLK(clk), .Q(\ram[3][168] ) );
  DFFX1_HVT \ram_reg[3][167]  ( .D(n996), .CLK(clk), .Q(\ram[3][167] ) );
  DFFX1_HVT \ram_reg[3][166]  ( .D(n995), .CLK(clk), .Q(\ram[3][166] ) );
  DFFX1_HVT \ram_reg[3][165]  ( .D(n994), .CLK(clk), .Q(\ram[3][165] ) );
  DFFX1_HVT \ram_reg[3][164]  ( .D(n993), .CLK(clk), .Q(\ram[3][164] ) );
  DFFX1_HVT \ram_reg[3][163]  ( .D(n992), .CLK(clk), .Q(\ram[3][163] ) );
  DFFX1_HVT \ram_reg[3][162]  ( .D(n991), .CLK(clk), .Q(\ram[3][162] ) );
  DFFX1_HVT \ram_reg[3][161]  ( .D(n990), .CLK(clk), .Q(\ram[3][161] ) );
  DFFX1_HVT \ram_reg[3][160]  ( .D(n989), .CLK(clk), .Q(\ram[3][160] ) );
  DFFX1_HVT \ram_reg[3][159]  ( .D(n988), .CLK(clk), .Q(\ram[3][159] ) );
  DFFX1_HVT \ram_reg[3][158]  ( .D(n987), .CLK(clk), .Q(\ram[3][158] ) );
  DFFX1_HVT \ram_reg[3][157]  ( .D(n986), .CLK(clk), .Q(\ram[3][157] ) );
  DFFX1_HVT \ram_reg[3][156]  ( .D(n985), .CLK(clk), .Q(\ram[3][156] ) );
  DFFX1_HVT \ram_reg[3][155]  ( .D(n984), .CLK(clk), .Q(\ram[3][155] ) );
  DFFX1_HVT \ram_reg[3][154]  ( .D(n983), .CLK(clk), .Q(\ram[3][154] ) );
  DFFX1_HVT \ram_reg[3][153]  ( .D(n982), .CLK(clk), .Q(\ram[3][153] ) );
  DFFX1_HVT \ram_reg[3][152]  ( .D(n981), .CLK(clk), .Q(\ram[3][152] ) );
  DFFX1_HVT \ram_reg[3][151]  ( .D(n980), .CLK(clk), .Q(\ram[3][151] ) );
  DFFX1_HVT \ram_reg[3][150]  ( .D(n979), .CLK(clk), .Q(\ram[3][150] ) );
  DFFX1_HVT \ram_reg[3][149]  ( .D(n978), .CLK(clk), .Q(\ram[3][149] ) );
  DFFX1_HVT \ram_reg[3][148]  ( .D(n977), .CLK(clk), .Q(\ram[3][148] ) );
  DFFX1_HVT \ram_reg[3][147]  ( .D(n976), .CLK(clk), .Q(\ram[3][147] ) );
  DFFX1_HVT \ram_reg[3][146]  ( .D(n975), .CLK(clk), .Q(\ram[3][146] ) );
  DFFX1_HVT \ram_reg[3][145]  ( .D(n974), .CLK(clk), .Q(\ram[3][145] ) );
  DFFX1_HVT \ram_reg[3][144]  ( .D(n973), .CLK(clk), .Q(\ram[3][144] ) );
  DFFX1_HVT \ram_reg[3][143]  ( .D(n972), .CLK(clk), .Q(\ram[3][143] ) );
  DFFX1_HVT \ram_reg[3][142]  ( .D(n971), .CLK(clk), .Q(\ram[3][142] ) );
  DFFX1_HVT \ram_reg[3][141]  ( .D(n970), .CLK(clk), .Q(\ram[3][141] ) );
  DFFX1_HVT \ram_reg[3][140]  ( .D(n969), .CLK(clk), .Q(\ram[3][140] ) );
  DFFX1_HVT \ram_reg[3][139]  ( .D(n968), .CLK(clk), .Q(\ram[3][139] ) );
  DFFX1_HVT \ram_reg[3][138]  ( .D(n967), .CLK(clk), .Q(\ram[3][138] ) );
  DFFX1_HVT \ram_reg[3][137]  ( .D(n966), .CLK(clk), .Q(\ram[3][137] ) );
  DFFX1_HVT \ram_reg[3][136]  ( .D(n965), .CLK(clk), .Q(\ram[3][136] ) );
  DFFX1_HVT \ram_reg[3][135]  ( .D(n964), .CLK(clk), .Q(\ram[3][135] ) );
  DFFX1_HVT \ram_reg[3][134]  ( .D(n963), .CLK(clk), .Q(\ram[3][134] ) );
  DFFX1_HVT \ram_reg[3][133]  ( .D(n962), .CLK(clk), .Q(\ram[3][133] ) );
  DFFX1_HVT \ram_reg[3][132]  ( .D(n961), .CLK(clk), .Q(\ram[3][132] ) );
  DFFX1_HVT \ram_reg[3][131]  ( .D(n960), .CLK(clk), .Q(\ram[3][131] ) );
  DFFX1_HVT \ram_reg[3][130]  ( .D(n959), .CLK(clk), .Q(\ram[3][130] ) );
  DFFX1_HVT \ram_reg[3][129]  ( .D(n958), .CLK(clk), .Q(\ram[3][129] ) );
  DFFX1_HVT \ram_reg[3][128]  ( .D(n957), .CLK(clk), .Q(\ram[3][128] ) );
  DFFX1_HVT \ram_reg[3][127]  ( .D(n956), .CLK(clk), .Q(\ram[3][127] ) );
  DFFX1_HVT \ram_reg[3][126]  ( .D(n955), .CLK(clk), .Q(\ram[3][126] ) );
  DFFX1_HVT \ram_reg[3][125]  ( .D(n954), .CLK(clk), .Q(\ram[3][125] ) );
  DFFX1_HVT \ram_reg[3][124]  ( .D(n953), .CLK(clk), .Q(\ram[3][124] ) );
  DFFX1_HVT \ram_reg[3][123]  ( .D(n952), .CLK(clk), .Q(\ram[3][123] ) );
  DFFX1_HVT \ram_reg[3][122]  ( .D(n951), .CLK(clk), .Q(\ram[3][122] ) );
  DFFX1_HVT \ram_reg[3][121]  ( .D(n950), .CLK(clk), .Q(\ram[3][121] ) );
  DFFX1_HVT \ram_reg[3][120]  ( .D(n949), .CLK(clk), .Q(\ram[3][120] ) );
  DFFX1_HVT \ram_reg[3][119]  ( .D(n948), .CLK(clk), .Q(\ram[3][119] ) );
  DFFX1_HVT \ram_reg[3][118]  ( .D(n947), .CLK(clk), .Q(\ram[3][118] ) );
  DFFX1_HVT \ram_reg[3][117]  ( .D(n946), .CLK(clk), .Q(\ram[3][117] ) );
  DFFX1_HVT \ram_reg[3][116]  ( .D(n945), .CLK(clk), .Q(\ram[3][116] ) );
  DFFX1_HVT \ram_reg[3][115]  ( .D(n944), .CLK(clk), .Q(\ram[3][115] ) );
  DFFX1_HVT \ram_reg[3][114]  ( .D(n943), .CLK(clk), .Q(\ram[3][114] ) );
  DFFX1_HVT \ram_reg[3][113]  ( .D(n942), .CLK(clk), .Q(\ram[3][113] ) );
  DFFX1_HVT \ram_reg[3][112]  ( .D(n941), .CLK(clk), .Q(\ram[3][112] ) );
  DFFX1_HVT \ram_reg[3][111]  ( .D(n940), .CLK(clk), .Q(\ram[3][111] ) );
  DFFX1_HVT \ram_reg[3][110]  ( .D(n939), .CLK(clk), .Q(\ram[3][110] ) );
  DFFX1_HVT \ram_reg[3][109]  ( .D(n938), .CLK(clk), .Q(\ram[3][109] ) );
  DFFX1_HVT \ram_reg[3][108]  ( .D(n937), .CLK(clk), .Q(\ram[3][108] ) );
  DFFX1_HVT \ram_reg[3][107]  ( .D(n936), .CLK(clk), .Q(\ram[3][107] ) );
  DFFX1_HVT \ram_reg[3][106]  ( .D(n935), .CLK(clk), .Q(\ram[3][106] ) );
  DFFX1_HVT \ram_reg[3][105]  ( .D(n934), .CLK(clk), .Q(\ram[3][105] ) );
  DFFX1_HVT \ram_reg[3][104]  ( .D(n933), .CLK(clk), .Q(\ram[3][104] ) );
  DFFX1_HVT \ram_reg[3][103]  ( .D(n932), .CLK(clk), .Q(\ram[3][103] ) );
  DFFX1_HVT \ram_reg[3][102]  ( .D(n931), .CLK(clk), .Q(\ram[3][102] ) );
  DFFX1_HVT \ram_reg[3][101]  ( .D(n930), .CLK(clk), .Q(\ram[3][101] ) );
  DFFX1_HVT \ram_reg[3][100]  ( .D(n929), .CLK(clk), .Q(\ram[3][100] ) );
  DFFX1_HVT \ram_reg[3][99]  ( .D(n928), .CLK(clk), .Q(\ram[3][99] ) );
  DFFX1_HVT \ram_reg[3][98]  ( .D(n927), .CLK(clk), .Q(\ram[3][98] ) );
  DFFX1_HVT \ram_reg[3][97]  ( .D(n926), .CLK(clk), .Q(\ram[3][97] ) );
  DFFX1_HVT \ram_reg[3][96]  ( .D(n925), .CLK(clk), .Q(\ram[3][96] ) );
  DFFX1_HVT \ram_reg[3][95]  ( .D(n924), .CLK(clk), .Q(\ram[3][95] ) );
  DFFX1_HVT \ram_reg[3][94]  ( .D(n923), .CLK(clk), .Q(\ram[3][94] ) );
  DFFX1_HVT \ram_reg[3][93]  ( .D(n922), .CLK(clk), .Q(\ram[3][93] ) );
  DFFX1_HVT \ram_reg[3][92]  ( .D(n921), .CLK(clk), .Q(\ram[3][92] ) );
  DFFX1_HVT \ram_reg[3][91]  ( .D(n920), .CLK(clk), .Q(\ram[3][91] ) );
  DFFX1_HVT \ram_reg[3][90]  ( .D(n919), .CLK(clk), .Q(\ram[3][90] ) );
  DFFX1_HVT \ram_reg[3][89]  ( .D(n918), .CLK(clk), .Q(\ram[3][89] ) );
  DFFX1_HVT \ram_reg[3][88]  ( .D(n917), .CLK(clk), .Q(\ram[3][88] ) );
  DFFX1_HVT \ram_reg[3][87]  ( .D(n916), .CLK(clk), .Q(\ram[3][87] ) );
  DFFX1_HVT \ram_reg[3][86]  ( .D(n915), .CLK(clk), .Q(\ram[3][86] ) );
  DFFX1_HVT \ram_reg[3][85]  ( .D(n914), .CLK(clk), .Q(\ram[3][85] ) );
  DFFX1_HVT \ram_reg[3][84]  ( .D(n913), .CLK(clk), .Q(\ram[3][84] ) );
  DFFX1_HVT \ram_reg[3][83]  ( .D(n912), .CLK(clk), .Q(\ram[3][83] ) );
  DFFX1_HVT \ram_reg[3][82]  ( .D(n911), .CLK(clk), .Q(\ram[3][82] ) );
  DFFX1_HVT \ram_reg[3][81]  ( .D(n910), .CLK(clk), .Q(\ram[3][81] ) );
  DFFX1_HVT \ram_reg[3][80]  ( .D(n909), .CLK(clk), .Q(\ram[3][80] ) );
  DFFX1_HVT \ram_reg[3][79]  ( .D(n908), .CLK(clk), .Q(\ram[3][79] ) );
  DFFX1_HVT \ram_reg[3][78]  ( .D(n907), .CLK(clk), .Q(\ram[3][78] ) );
  DFFX1_HVT \ram_reg[3][77]  ( .D(n906), .CLK(clk), .Q(\ram[3][77] ) );
  DFFX1_HVT \ram_reg[3][76]  ( .D(n905), .CLK(clk), .Q(\ram[3][76] ) );
  DFFX1_HVT \ram_reg[3][75]  ( .D(n904), .CLK(clk), .Q(\ram[3][75] ) );
  DFFX1_HVT \ram_reg[3][74]  ( .D(n903), .CLK(clk), .Q(\ram[3][74] ) );
  DFFX1_HVT \ram_reg[3][73]  ( .D(n902), .CLK(clk), .Q(\ram[3][73] ) );
  DFFX1_HVT \ram_reg[3][72]  ( .D(n901), .CLK(clk), .Q(\ram[3][72] ) );
  DFFX1_HVT \ram_reg[3][71]  ( .D(n900), .CLK(clk), .Q(\ram[3][71] ) );
  DFFX1_HVT \ram_reg[3][70]  ( .D(n899), .CLK(clk), .Q(\ram[3][70] ) );
  DFFX1_HVT \ram_reg[3][69]  ( .D(n898), .CLK(clk), .Q(\ram[3][69] ) );
  DFFX1_HVT \ram_reg[3][68]  ( .D(n897), .CLK(clk), .Q(\ram[3][68] ) );
  DFFX1_HVT \ram_reg[3][67]  ( .D(n896), .CLK(clk), .Q(\ram[3][67] ) );
  DFFX1_HVT \ram_reg[3][66]  ( .D(n895), .CLK(clk), .Q(\ram[3][66] ) );
  DFFX1_HVT \ram_reg[3][65]  ( .D(n894), .CLK(clk), .Q(\ram[3][65] ) );
  DFFX1_HVT \ram_reg[3][64]  ( .D(n893), .CLK(clk), .Q(\ram[3][64] ) );
  DFFX1_HVT \ram_reg[3][63]  ( .D(n892), .CLK(clk), .Q(\ram[3][63] ) );
  DFFX1_HVT \ram_reg[3][62]  ( .D(n891), .CLK(clk), .Q(\ram[3][62] ) );
  DFFX1_HVT \ram_reg[3][61]  ( .D(n890), .CLK(clk), .Q(\ram[3][61] ) );
  DFFX1_HVT \ram_reg[3][60]  ( .D(n889), .CLK(clk), .Q(\ram[3][60] ) );
  DFFX1_HVT \ram_reg[3][59]  ( .D(n888), .CLK(clk), .Q(\ram[3][59] ) );
  DFFX1_HVT \ram_reg[3][58]  ( .D(n887), .CLK(clk), .Q(\ram[3][58] ) );
  DFFX1_HVT \ram_reg[3][57]  ( .D(n886), .CLK(clk), .Q(\ram[3][57] ) );
  DFFX1_HVT \ram_reg[3][56]  ( .D(n885), .CLK(clk), .Q(\ram[3][56] ) );
  DFFX1_HVT \ram_reg[3][55]  ( .D(n884), .CLK(clk), .Q(\ram[3][55] ) );
  DFFX1_HVT \ram_reg[3][54]  ( .D(n883), .CLK(clk), .Q(\ram[3][54] ) );
  DFFX1_HVT \ram_reg[3][53]  ( .D(n882), .CLK(clk), .Q(\ram[3][53] ) );
  DFFX1_HVT \ram_reg[3][52]  ( .D(n881), .CLK(clk), .Q(\ram[3][52] ) );
  DFFX1_HVT \ram_reg[3][51]  ( .D(n880), .CLK(clk), .Q(\ram[3][51] ) );
  DFFX1_HVT \ram_reg[3][50]  ( .D(n879), .CLK(clk), .Q(\ram[3][50] ) );
  DFFX1_HVT \ram_reg[3][49]  ( .D(n878), .CLK(clk), .Q(\ram[3][49] ) );
  DFFX1_HVT \ram_reg[3][48]  ( .D(n877), .CLK(clk), .Q(\ram[3][48] ) );
  DFFX1_HVT \ram_reg[3][47]  ( .D(n876), .CLK(clk), .Q(\ram[3][47] ) );
  DFFX1_HVT \ram_reg[3][46]  ( .D(n875), .CLK(clk), .Q(\ram[3][46] ) );
  DFFX1_HVT \ram_reg[3][45]  ( .D(n874), .CLK(clk), .Q(\ram[3][45] ) );
  DFFX1_HVT \ram_reg[3][44]  ( .D(n873), .CLK(clk), .Q(\ram[3][44] ) );
  DFFX1_HVT \ram_reg[3][43]  ( .D(n872), .CLK(clk), .Q(\ram[3][43] ) );
  DFFX1_HVT \ram_reg[3][42]  ( .D(n871), .CLK(clk), .Q(\ram[3][42] ) );
  DFFX1_HVT \ram_reg[3][41]  ( .D(n870), .CLK(clk), .Q(\ram[3][41] ) );
  DFFX1_HVT \ram_reg[3][40]  ( .D(n869), .CLK(clk), .Q(\ram[3][40] ) );
  DFFX1_HVT \ram_reg[3][39]  ( .D(n868), .CLK(clk), .Q(\ram[3][39] ) );
  DFFX1_HVT \ram_reg[3][38]  ( .D(n867), .CLK(clk), .Q(\ram[3][38] ) );
  DFFX1_HVT \ram_reg[3][37]  ( .D(n866), .CLK(clk), .Q(\ram[3][37] ) );
  DFFX1_HVT \ram_reg[3][36]  ( .D(n865), .CLK(clk), .Q(\ram[3][36] ) );
  DFFX1_HVT \ram_reg[3][35]  ( .D(n864), .CLK(clk), .Q(\ram[3][35] ) );
  DFFX1_HVT \ram_reg[3][34]  ( .D(n863), .CLK(clk), .Q(\ram[3][34] ) );
  DFFX1_HVT \ram_reg[3][33]  ( .D(n862), .CLK(clk), .Q(\ram[3][33] ) );
  DFFX1_HVT \ram_reg[3][32]  ( .D(n861), .CLK(clk), .Q(\ram[3][32] ) );
  DFFX1_HVT \ram_reg[3][31]  ( .D(n860), .CLK(clk), .Q(\ram[3][31] ) );
  DFFX1_HVT \ram_reg[3][30]  ( .D(n859), .CLK(clk), .Q(\ram[3][30] ) );
  DFFX1_HVT \ram_reg[3][29]  ( .D(n858), .CLK(clk), .Q(\ram[3][29] ) );
  DFFX1_HVT \ram_reg[3][28]  ( .D(n857), .CLK(clk), .Q(\ram[3][28] ) );
  DFFX1_HVT \ram_reg[3][27]  ( .D(n856), .CLK(clk), .Q(\ram[3][27] ) );
  DFFX1_HVT \ram_reg[3][26]  ( .D(n855), .CLK(clk), .Q(\ram[3][26] ) );
  DFFX1_HVT \ram_reg[3][25]  ( .D(n854), .CLK(clk), .Q(\ram[3][25] ) );
  DFFX1_HVT \ram_reg[3][24]  ( .D(n853), .CLK(clk), .Q(\ram[3][24] ) );
  DFFX1_HVT \ram_reg[3][23]  ( .D(n852), .CLK(clk), .Q(\ram[3][23] ) );
  DFFX1_HVT \ram_reg[3][22]  ( .D(n851), .CLK(clk), .Q(\ram[3][22] ) );
  DFFX1_HVT \ram_reg[3][21]  ( .D(n850), .CLK(clk), .Q(\ram[3][21] ) );
  DFFX1_HVT \ram_reg[3][20]  ( .D(n849), .CLK(clk), .Q(\ram[3][20] ) );
  DFFX1_HVT \ram_reg[3][19]  ( .D(n848), .CLK(clk), .Q(\ram[3][19] ) );
  DFFX1_HVT \ram_reg[3][18]  ( .D(n847), .CLK(clk), .Q(\ram[3][18] ) );
  DFFX1_HVT \ram_reg[3][17]  ( .D(n846), .CLK(clk), .Q(\ram[3][17] ) );
  DFFX1_HVT \ram_reg[3][16]  ( .D(n845), .CLK(clk), .Q(\ram[3][16] ) );
  DFFX1_HVT \ram_reg[3][15]  ( .D(n844), .CLK(clk), .Q(\ram[3][15] ) );
  DFFX1_HVT \ram_reg[3][14]  ( .D(n843), .CLK(clk), .Q(\ram[3][14] ) );
  DFFX1_HVT \ram_reg[3][13]  ( .D(n842), .CLK(clk), .Q(\ram[3][13] ) );
  DFFX1_HVT \ram_reg[3][12]  ( .D(n841), .CLK(clk), .Q(\ram[3][12] ) );
  DFFX1_HVT \ram_reg[3][11]  ( .D(n840), .CLK(clk), .Q(\ram[3][11] ) );
  DFFX1_HVT \ram_reg[3][10]  ( .D(n839), .CLK(clk), .Q(\ram[3][10] ) );
  DFFX1_HVT \ram_reg[3][9]  ( .D(n838), .CLK(clk), .Q(\ram[3][9] ) );
  DFFX1_HVT \ram_reg[3][8]  ( .D(n837), .CLK(clk), .Q(\ram[3][8] ) );
  DFFX1_HVT \ram_reg[3][7]  ( .D(n836), .CLK(clk), .Q(\ram[3][7] ) );
  DFFX1_HVT \ram_reg[3][6]  ( .D(n835), .CLK(clk), .Q(\ram[3][6] ) );
  DFFX1_HVT \ram_reg[3][5]  ( .D(n834), .CLK(clk), .Q(\ram[3][5] ) );
  DFFX1_HVT \ram_reg[3][4]  ( .D(n833), .CLK(clk), .Q(\ram[3][4] ) );
  DFFX1_HVT \ram_reg[3][3]  ( .D(n832), .CLK(clk), .Q(\ram[3][3] ) );
  DFFX1_HVT \ram_reg[3][2]  ( .D(n831), .CLK(clk), .Q(\ram[3][2] ) );
  DFFX1_HVT \ram_reg[3][1]  ( .D(n830), .CLK(clk), .Q(\ram[3][1] ) );
  DFFX1_HVT \ram_reg[3][0]  ( .D(n829), .CLK(clk), .Q(\ram[3][0] ) );
  DFFX1_HVT \ram_reg[2][255]  ( .D(n828), .CLK(clk), .Q(\ram[2][255] ) );
  DFFX1_HVT \ram_reg[2][254]  ( .D(n827), .CLK(clk), .Q(\ram[2][254] ) );
  DFFX1_HVT \ram_reg[2][253]  ( .D(n826), .CLK(clk), .Q(\ram[2][253] ) );
  DFFX1_HVT \ram_reg[2][252]  ( .D(n825), .CLK(clk), .Q(\ram[2][252] ) );
  DFFX1_HVT \ram_reg[2][251]  ( .D(n824), .CLK(clk), .Q(\ram[2][251] ) );
  DFFX1_HVT \ram_reg[2][250]  ( .D(n823), .CLK(clk), .Q(\ram[2][250] ) );
  DFFX1_HVT \ram_reg[2][249]  ( .D(n822), .CLK(clk), .Q(\ram[2][249] ) );
  DFFX1_HVT \ram_reg[2][248]  ( .D(n821), .CLK(clk), .Q(\ram[2][248] ) );
  DFFX1_HVT \ram_reg[2][247]  ( .D(n820), .CLK(clk), .Q(\ram[2][247] ) );
  DFFX1_HVT \ram_reg[2][246]  ( .D(n819), .CLK(clk), .Q(\ram[2][246] ) );
  DFFX1_HVT \ram_reg[2][245]  ( .D(n818), .CLK(clk), .Q(\ram[2][245] ) );
  DFFX1_HVT \ram_reg[2][244]  ( .D(n817), .CLK(clk), .Q(\ram[2][244] ) );
  DFFX1_HVT \ram_reg[2][243]  ( .D(n816), .CLK(clk), .Q(\ram[2][243] ) );
  DFFX1_HVT \ram_reg[2][242]  ( .D(n815), .CLK(clk), .Q(\ram[2][242] ) );
  DFFX1_HVT \ram_reg[2][241]  ( .D(n814), .CLK(clk), .Q(\ram[2][241] ) );
  DFFX1_HVT \ram_reg[2][240]  ( .D(n813), .CLK(clk), .Q(\ram[2][240] ) );
  DFFX1_HVT \ram_reg[2][239]  ( .D(n812), .CLK(clk), .Q(\ram[2][239] ) );
  DFFX1_HVT \ram_reg[2][238]  ( .D(n811), .CLK(clk), .Q(\ram[2][238] ) );
  DFFX1_HVT \ram_reg[2][237]  ( .D(n810), .CLK(clk), .Q(\ram[2][237] ) );
  DFFX1_HVT \ram_reg[2][236]  ( .D(n809), .CLK(clk), .Q(\ram[2][236] ) );
  DFFX1_HVT \ram_reg[2][235]  ( .D(n808), .CLK(clk), .Q(\ram[2][235] ) );
  DFFX1_HVT \ram_reg[2][234]  ( .D(n807), .CLK(clk), .Q(\ram[2][234] ) );
  DFFX1_HVT \ram_reg[2][233]  ( .D(n806), .CLK(clk), .Q(\ram[2][233] ) );
  DFFX1_HVT \ram_reg[2][232]  ( .D(n805), .CLK(clk), .Q(\ram[2][232] ) );
  DFFX1_HVT \ram_reg[2][231]  ( .D(n804), .CLK(clk), .Q(\ram[2][231] ) );
  DFFX1_HVT \ram_reg[2][230]  ( .D(n803), .CLK(clk), .Q(\ram[2][230] ) );
  DFFX1_HVT \ram_reg[2][229]  ( .D(n802), .CLK(clk), .Q(\ram[2][229] ) );
  DFFX1_HVT \ram_reg[2][228]  ( .D(n801), .CLK(clk), .Q(\ram[2][228] ) );
  DFFX1_HVT \ram_reg[2][227]  ( .D(n800), .CLK(clk), .Q(\ram[2][227] ) );
  DFFX1_HVT \ram_reg[2][226]  ( .D(n799), .CLK(clk), .Q(\ram[2][226] ) );
  DFFX1_HVT \ram_reg[2][225]  ( .D(n798), .CLK(clk), .Q(\ram[2][225] ) );
  DFFX1_HVT \ram_reg[2][224]  ( .D(n797), .CLK(clk), .Q(\ram[2][224] ) );
  DFFX1_HVT \ram_reg[2][223]  ( .D(n796), .CLK(clk), .Q(\ram[2][223] ) );
  DFFX1_HVT \ram_reg[2][222]  ( .D(n795), .CLK(clk), .Q(\ram[2][222] ) );
  DFFX1_HVT \ram_reg[2][221]  ( .D(n794), .CLK(clk), .Q(\ram[2][221] ) );
  DFFX1_HVT \ram_reg[2][220]  ( .D(n793), .CLK(clk), .Q(\ram[2][220] ) );
  DFFX1_HVT \ram_reg[2][219]  ( .D(n792), .CLK(clk), .Q(\ram[2][219] ) );
  DFFX1_HVT \ram_reg[2][218]  ( .D(n791), .CLK(clk), .Q(\ram[2][218] ) );
  DFFX1_HVT \ram_reg[2][217]  ( .D(n790), .CLK(clk), .Q(\ram[2][217] ) );
  DFFX1_HVT \ram_reg[2][216]  ( .D(n789), .CLK(clk), .Q(\ram[2][216] ) );
  DFFX1_HVT \ram_reg[2][215]  ( .D(n788), .CLK(clk), .Q(\ram[2][215] ) );
  DFFX1_HVT \ram_reg[2][214]  ( .D(n787), .CLK(clk), .Q(\ram[2][214] ) );
  DFFX1_HVT \ram_reg[2][213]  ( .D(n786), .CLK(clk), .Q(\ram[2][213] ) );
  DFFX1_HVT \ram_reg[2][212]  ( .D(n785), .CLK(clk), .Q(\ram[2][212] ) );
  DFFX1_HVT \ram_reg[2][211]  ( .D(n784), .CLK(clk), .Q(\ram[2][211] ) );
  DFFX1_HVT \ram_reg[2][210]  ( .D(n783), .CLK(clk), .Q(\ram[2][210] ) );
  DFFX1_HVT \ram_reg[2][209]  ( .D(n782), .CLK(clk), .Q(\ram[2][209] ) );
  DFFX1_HVT \ram_reg[2][208]  ( .D(n781), .CLK(clk), .Q(\ram[2][208] ) );
  DFFX1_HVT \ram_reg[2][207]  ( .D(n780), .CLK(clk), .Q(\ram[2][207] ) );
  DFFX1_HVT \ram_reg[2][206]  ( .D(n779), .CLK(clk), .Q(\ram[2][206] ) );
  DFFX1_HVT \ram_reg[2][205]  ( .D(n778), .CLK(clk), .Q(\ram[2][205] ) );
  DFFX1_HVT \ram_reg[2][204]  ( .D(n777), .CLK(clk), .Q(\ram[2][204] ) );
  DFFX1_HVT \ram_reg[2][203]  ( .D(n776), .CLK(clk), .Q(\ram[2][203] ) );
  DFFX1_HVT \ram_reg[2][202]  ( .D(n775), .CLK(clk), .Q(\ram[2][202] ) );
  DFFX1_HVT \ram_reg[2][201]  ( .D(n774), .CLK(clk), .Q(\ram[2][201] ) );
  DFFX1_HVT \ram_reg[2][200]  ( .D(n773), .CLK(clk), .Q(\ram[2][200] ) );
  DFFX1_HVT \ram_reg[2][199]  ( .D(n772), .CLK(clk), .Q(\ram[2][199] ) );
  DFFX1_HVT \ram_reg[2][198]  ( .D(n771), .CLK(clk), .Q(\ram[2][198] ) );
  DFFX1_HVT \ram_reg[2][197]  ( .D(n770), .CLK(clk), .Q(\ram[2][197] ) );
  DFFX1_HVT \ram_reg[2][196]  ( .D(n769), .CLK(clk), .Q(\ram[2][196] ) );
  DFFX1_HVT \ram_reg[2][195]  ( .D(n768), .CLK(clk), .Q(\ram[2][195] ) );
  DFFX1_HVT \ram_reg[2][194]  ( .D(n767), .CLK(clk), .Q(\ram[2][194] ) );
  DFFX1_HVT \ram_reg[2][193]  ( .D(n766), .CLK(clk), .Q(\ram[2][193] ) );
  DFFX1_HVT \ram_reg[2][192]  ( .D(n765), .CLK(clk), .Q(\ram[2][192] ) );
  DFFX1_HVT \ram_reg[2][191]  ( .D(n764), .CLK(clk), .Q(\ram[2][191] ) );
  DFFX1_HVT \ram_reg[2][190]  ( .D(n763), .CLK(clk), .Q(\ram[2][190] ) );
  DFFX1_HVT \ram_reg[2][189]  ( .D(n762), .CLK(clk), .Q(\ram[2][189] ) );
  DFFX1_HVT \ram_reg[2][188]  ( .D(n761), .CLK(clk), .Q(\ram[2][188] ) );
  DFFX1_HVT \ram_reg[2][187]  ( .D(n760), .CLK(clk), .Q(\ram[2][187] ) );
  DFFX1_HVT \ram_reg[2][186]  ( .D(n759), .CLK(clk), .Q(\ram[2][186] ) );
  DFFX1_HVT \ram_reg[2][185]  ( .D(n758), .CLK(clk), .Q(\ram[2][185] ) );
  DFFX1_HVT \ram_reg[2][184]  ( .D(n757), .CLK(clk), .Q(\ram[2][184] ) );
  DFFX1_HVT \ram_reg[2][183]  ( .D(n756), .CLK(clk), .Q(\ram[2][183] ) );
  DFFX1_HVT \ram_reg[2][182]  ( .D(n755), .CLK(clk), .Q(\ram[2][182] ) );
  DFFX1_HVT \ram_reg[2][181]  ( .D(n754), .CLK(clk), .Q(\ram[2][181] ) );
  DFFX1_HVT \ram_reg[2][180]  ( .D(n753), .CLK(clk), .Q(\ram[2][180] ) );
  DFFX1_HVT \ram_reg[2][179]  ( .D(n752), .CLK(clk), .Q(\ram[2][179] ) );
  DFFX1_HVT \ram_reg[2][178]  ( .D(n751), .CLK(clk), .Q(\ram[2][178] ) );
  DFFX1_HVT \ram_reg[2][177]  ( .D(n750), .CLK(clk), .Q(\ram[2][177] ) );
  DFFX1_HVT \ram_reg[2][176]  ( .D(n749), .CLK(clk), .Q(\ram[2][176] ) );
  DFFX1_HVT \ram_reg[2][175]  ( .D(n748), .CLK(clk), .Q(\ram[2][175] ) );
  DFFX1_HVT \ram_reg[2][174]  ( .D(n747), .CLK(clk), .Q(\ram[2][174] ) );
  DFFX1_HVT \ram_reg[2][173]  ( .D(n746), .CLK(clk), .Q(\ram[2][173] ) );
  DFFX1_HVT \ram_reg[2][172]  ( .D(n745), .CLK(clk), .Q(\ram[2][172] ) );
  DFFX1_HVT \ram_reg[2][171]  ( .D(n744), .CLK(clk), .Q(\ram[2][171] ) );
  DFFX1_HVT \ram_reg[2][170]  ( .D(n743), .CLK(clk), .Q(\ram[2][170] ) );
  DFFX1_HVT \ram_reg[2][169]  ( .D(n742), .CLK(clk), .Q(\ram[2][169] ) );
  DFFX1_HVT \ram_reg[2][168]  ( .D(n741), .CLK(clk), .Q(\ram[2][168] ) );
  DFFX1_HVT \ram_reg[2][167]  ( .D(n740), .CLK(clk), .Q(\ram[2][167] ) );
  DFFX1_HVT \ram_reg[2][166]  ( .D(n739), .CLK(clk), .Q(\ram[2][166] ) );
  DFFX1_HVT \ram_reg[2][165]  ( .D(n738), .CLK(clk), .Q(\ram[2][165] ) );
  DFFX1_HVT \ram_reg[2][164]  ( .D(n737), .CLK(clk), .Q(\ram[2][164] ) );
  DFFX1_HVT \ram_reg[2][163]  ( .D(n736), .CLK(clk), .Q(\ram[2][163] ) );
  DFFX1_HVT \ram_reg[2][162]  ( .D(n735), .CLK(clk), .Q(\ram[2][162] ) );
  DFFX1_HVT \ram_reg[2][161]  ( .D(n734), .CLK(clk), .Q(\ram[2][161] ) );
  DFFX1_HVT \ram_reg[2][160]  ( .D(n733), .CLK(clk), .Q(\ram[2][160] ) );
  DFFX1_HVT \ram_reg[2][159]  ( .D(n732), .CLK(clk), .Q(\ram[2][159] ) );
  DFFX1_HVT \ram_reg[2][158]  ( .D(n731), .CLK(clk), .Q(\ram[2][158] ) );
  DFFX1_HVT \ram_reg[2][157]  ( .D(n730), .CLK(clk), .Q(\ram[2][157] ) );
  DFFX1_HVT \ram_reg[2][156]  ( .D(n729), .CLK(clk), .Q(\ram[2][156] ) );
  DFFX1_HVT \ram_reg[2][155]  ( .D(n728), .CLK(clk), .Q(\ram[2][155] ) );
  DFFX1_HVT \ram_reg[2][154]  ( .D(n727), .CLK(clk), .Q(\ram[2][154] ) );
  DFFX1_HVT \ram_reg[2][153]  ( .D(n726), .CLK(clk), .Q(\ram[2][153] ) );
  DFFX1_HVT \ram_reg[2][152]  ( .D(n725), .CLK(clk), .Q(\ram[2][152] ) );
  DFFX1_HVT \ram_reg[2][151]  ( .D(n724), .CLK(clk), .Q(\ram[2][151] ) );
  DFFX1_HVT \ram_reg[2][150]  ( .D(n723), .CLK(clk), .Q(\ram[2][150] ) );
  DFFX1_HVT \ram_reg[2][149]  ( .D(n722), .CLK(clk), .Q(\ram[2][149] ) );
  DFFX1_HVT \ram_reg[2][148]  ( .D(n721), .CLK(clk), .Q(\ram[2][148] ) );
  DFFX1_HVT \ram_reg[2][147]  ( .D(n720), .CLK(clk), .Q(\ram[2][147] ) );
  DFFX1_HVT \ram_reg[2][146]  ( .D(n719), .CLK(clk), .Q(\ram[2][146] ) );
  DFFX1_HVT \ram_reg[2][145]  ( .D(n718), .CLK(clk), .Q(\ram[2][145] ) );
  DFFX1_HVT \ram_reg[2][144]  ( .D(n717), .CLK(clk), .Q(\ram[2][144] ) );
  DFFX1_HVT \ram_reg[2][143]  ( .D(n716), .CLK(clk), .Q(\ram[2][143] ) );
  DFFX1_HVT \ram_reg[2][142]  ( .D(n715), .CLK(clk), .Q(\ram[2][142] ) );
  DFFX1_HVT \ram_reg[2][141]  ( .D(n714), .CLK(clk), .Q(\ram[2][141] ) );
  DFFX1_HVT \ram_reg[2][140]  ( .D(n713), .CLK(clk), .Q(\ram[2][140] ) );
  DFFX1_HVT \ram_reg[2][139]  ( .D(n712), .CLK(clk), .Q(\ram[2][139] ) );
  DFFX1_HVT \ram_reg[2][138]  ( .D(n711), .CLK(clk), .Q(\ram[2][138] ) );
  DFFX1_HVT \ram_reg[2][137]  ( .D(n710), .CLK(clk), .Q(\ram[2][137] ) );
  DFFX1_HVT \ram_reg[2][136]  ( .D(n709), .CLK(clk), .Q(\ram[2][136] ) );
  DFFX1_HVT \ram_reg[2][135]  ( .D(n708), .CLK(clk), .Q(\ram[2][135] ) );
  DFFX1_HVT \ram_reg[2][134]  ( .D(n707), .CLK(clk), .Q(\ram[2][134] ) );
  DFFX1_HVT \ram_reg[2][133]  ( .D(n706), .CLK(clk), .Q(\ram[2][133] ) );
  DFFX1_HVT \ram_reg[2][132]  ( .D(n705), .CLK(clk), .Q(\ram[2][132] ) );
  DFFX1_HVT \ram_reg[2][131]  ( .D(n704), .CLK(clk), .Q(\ram[2][131] ) );
  DFFX1_HVT \ram_reg[2][130]  ( .D(n703), .CLK(clk), .Q(\ram[2][130] ) );
  DFFX1_HVT \ram_reg[2][129]  ( .D(n702), .CLK(clk), .Q(\ram[2][129] ) );
  DFFX1_HVT \ram_reg[2][128]  ( .D(n701), .CLK(clk), .Q(\ram[2][128] ) );
  DFFX1_HVT \ram_reg[2][127]  ( .D(n700), .CLK(clk), .Q(\ram[2][127] ) );
  DFFX1_HVT \ram_reg[2][126]  ( .D(n699), .CLK(clk), .Q(\ram[2][126] ) );
  DFFX1_HVT \ram_reg[2][125]  ( .D(n698), .CLK(clk), .Q(\ram[2][125] ) );
  DFFX1_HVT \ram_reg[2][124]  ( .D(n697), .CLK(clk), .Q(\ram[2][124] ) );
  DFFX1_HVT \ram_reg[2][123]  ( .D(n696), .CLK(clk), .Q(\ram[2][123] ) );
  DFFX1_HVT \ram_reg[2][122]  ( .D(n695), .CLK(clk), .Q(\ram[2][122] ) );
  DFFX1_HVT \ram_reg[2][121]  ( .D(n694), .CLK(clk), .Q(\ram[2][121] ) );
  DFFX1_HVT \ram_reg[2][120]  ( .D(n693), .CLK(clk), .Q(\ram[2][120] ) );
  DFFX1_HVT \ram_reg[2][119]  ( .D(n692), .CLK(clk), .Q(\ram[2][119] ) );
  DFFX1_HVT \ram_reg[2][118]  ( .D(n691), .CLK(clk), .Q(\ram[2][118] ) );
  DFFX1_HVT \ram_reg[2][117]  ( .D(n690), .CLK(clk), .Q(\ram[2][117] ) );
  DFFX1_HVT \ram_reg[2][116]  ( .D(n689), .CLK(clk), .Q(\ram[2][116] ) );
  DFFX1_HVT \ram_reg[2][115]  ( .D(n688), .CLK(clk), .Q(\ram[2][115] ) );
  DFFX1_HVT \ram_reg[2][114]  ( .D(n687), .CLK(clk), .Q(\ram[2][114] ) );
  DFFX1_HVT \ram_reg[2][113]  ( .D(n686), .CLK(clk), .Q(\ram[2][113] ) );
  DFFX1_HVT \ram_reg[2][112]  ( .D(n685), .CLK(clk), .Q(\ram[2][112] ) );
  DFFX1_HVT \ram_reg[2][111]  ( .D(n684), .CLK(clk), .Q(\ram[2][111] ) );
  DFFX1_HVT \ram_reg[2][110]  ( .D(n683), .CLK(clk), .Q(\ram[2][110] ) );
  DFFX1_HVT \ram_reg[2][109]  ( .D(n682), .CLK(clk), .Q(\ram[2][109] ) );
  DFFX1_HVT \ram_reg[2][108]  ( .D(n681), .CLK(clk), .Q(\ram[2][108] ) );
  DFFX1_HVT \ram_reg[2][107]  ( .D(n680), .CLK(clk), .Q(\ram[2][107] ) );
  DFFX1_HVT \ram_reg[2][106]  ( .D(n679), .CLK(clk), .Q(\ram[2][106] ) );
  DFFX1_HVT \ram_reg[2][105]  ( .D(n678), .CLK(clk), .Q(\ram[2][105] ) );
  DFFX1_HVT \ram_reg[2][104]  ( .D(n677), .CLK(clk), .Q(\ram[2][104] ) );
  DFFX1_HVT \ram_reg[2][103]  ( .D(n676), .CLK(clk), .Q(\ram[2][103] ) );
  DFFX1_HVT \ram_reg[2][102]  ( .D(n675), .CLK(clk), .Q(\ram[2][102] ) );
  DFFX1_HVT \ram_reg[2][101]  ( .D(n674), .CLK(clk), .Q(\ram[2][101] ) );
  DFFX1_HVT \ram_reg[2][100]  ( .D(n673), .CLK(clk), .Q(\ram[2][100] ) );
  DFFX1_HVT \ram_reg[2][99]  ( .D(n672), .CLK(clk), .Q(\ram[2][99] ) );
  DFFX1_HVT \ram_reg[2][98]  ( .D(n671), .CLK(clk), .Q(\ram[2][98] ) );
  DFFX1_HVT \ram_reg[2][97]  ( .D(n670), .CLK(clk), .Q(\ram[2][97] ) );
  DFFX1_HVT \ram_reg[2][96]  ( .D(n669), .CLK(clk), .Q(\ram[2][96] ) );
  DFFX1_HVT \ram_reg[2][95]  ( .D(n668), .CLK(clk), .Q(\ram[2][95] ) );
  DFFX1_HVT \ram_reg[2][94]  ( .D(n667), .CLK(clk), .Q(\ram[2][94] ) );
  DFFX1_HVT \ram_reg[2][93]  ( .D(n666), .CLK(clk), .Q(\ram[2][93] ) );
  DFFX1_HVT \ram_reg[2][92]  ( .D(n665), .CLK(clk), .Q(\ram[2][92] ) );
  DFFX1_HVT \ram_reg[2][91]  ( .D(n664), .CLK(clk), .Q(\ram[2][91] ) );
  DFFX1_HVT \ram_reg[2][90]  ( .D(n663), .CLK(clk), .Q(\ram[2][90] ) );
  DFFX1_HVT \ram_reg[2][89]  ( .D(n662), .CLK(clk), .Q(\ram[2][89] ) );
  DFFX1_HVT \ram_reg[2][88]  ( .D(n661), .CLK(clk), .Q(\ram[2][88] ) );
  DFFX1_HVT \ram_reg[2][87]  ( .D(n660), .CLK(clk), .Q(\ram[2][87] ) );
  DFFX1_HVT \ram_reg[2][86]  ( .D(n659), .CLK(clk), .Q(\ram[2][86] ) );
  DFFX1_HVT \ram_reg[2][85]  ( .D(n658), .CLK(clk), .Q(\ram[2][85] ) );
  DFFX1_HVT \ram_reg[2][84]  ( .D(n657), .CLK(clk), .Q(\ram[2][84] ) );
  DFFX1_HVT \ram_reg[2][83]  ( .D(n656), .CLK(clk), .Q(\ram[2][83] ) );
  DFFX1_HVT \ram_reg[2][82]  ( .D(n655), .CLK(clk), .Q(\ram[2][82] ) );
  DFFX1_HVT \ram_reg[2][81]  ( .D(n654), .CLK(clk), .Q(\ram[2][81] ) );
  DFFX1_HVT \ram_reg[2][80]  ( .D(n653), .CLK(clk), .Q(\ram[2][80] ) );
  DFFX1_HVT \ram_reg[2][79]  ( .D(n652), .CLK(clk), .Q(\ram[2][79] ) );
  DFFX1_HVT \ram_reg[2][78]  ( .D(n651), .CLK(clk), .Q(\ram[2][78] ) );
  DFFX1_HVT \ram_reg[2][77]  ( .D(n650), .CLK(clk), .Q(\ram[2][77] ) );
  DFFX1_HVT \ram_reg[2][76]  ( .D(n649), .CLK(clk), .Q(\ram[2][76] ) );
  DFFX1_HVT \ram_reg[2][75]  ( .D(n648), .CLK(clk), .Q(\ram[2][75] ) );
  DFFX1_HVT \ram_reg[2][74]  ( .D(n647), .CLK(clk), .Q(\ram[2][74] ) );
  DFFX1_HVT \ram_reg[2][73]  ( .D(n646), .CLK(clk), .Q(\ram[2][73] ) );
  DFFX1_HVT \ram_reg[2][72]  ( .D(n645), .CLK(clk), .Q(\ram[2][72] ) );
  DFFX1_HVT \ram_reg[2][71]  ( .D(n644), .CLK(clk), .Q(\ram[2][71] ) );
  DFFX1_HVT \ram_reg[2][70]  ( .D(n643), .CLK(clk), .Q(\ram[2][70] ) );
  DFFX1_HVT \ram_reg[2][69]  ( .D(n642), .CLK(clk), .Q(\ram[2][69] ) );
  DFFX1_HVT \ram_reg[2][68]  ( .D(n641), .CLK(clk), .Q(\ram[2][68] ) );
  DFFX1_HVT \ram_reg[2][67]  ( .D(n640), .CLK(clk), .Q(\ram[2][67] ) );
  DFFX1_HVT \ram_reg[2][66]  ( .D(n639), .CLK(clk), .Q(\ram[2][66] ) );
  DFFX1_HVT \ram_reg[2][65]  ( .D(n638), .CLK(clk), .Q(\ram[2][65] ) );
  DFFX1_HVT \ram_reg[2][64]  ( .D(n637), .CLK(clk), .Q(\ram[2][64] ) );
  DFFX1_HVT \ram_reg[2][63]  ( .D(n636), .CLK(clk), .Q(\ram[2][63] ) );
  DFFX1_HVT \ram_reg[2][62]  ( .D(n635), .CLK(clk), .Q(\ram[2][62] ) );
  DFFX1_HVT \ram_reg[2][61]  ( .D(n634), .CLK(clk), .Q(\ram[2][61] ) );
  DFFX1_HVT \ram_reg[2][60]  ( .D(n633), .CLK(clk), .Q(\ram[2][60] ) );
  DFFX1_HVT \ram_reg[2][59]  ( .D(n632), .CLK(clk), .Q(\ram[2][59] ) );
  DFFX1_HVT \ram_reg[2][58]  ( .D(n631), .CLK(clk), .Q(\ram[2][58] ) );
  DFFX1_HVT \ram_reg[2][57]  ( .D(n630), .CLK(clk), .Q(\ram[2][57] ) );
  DFFX1_HVT \ram_reg[2][56]  ( .D(n629), .CLK(clk), .Q(\ram[2][56] ) );
  DFFX1_HVT \ram_reg[2][55]  ( .D(n628), .CLK(clk), .Q(\ram[2][55] ) );
  DFFX1_HVT \ram_reg[2][54]  ( .D(n627), .CLK(clk), .Q(\ram[2][54] ) );
  DFFX1_HVT \ram_reg[2][53]  ( .D(n626), .CLK(clk), .Q(\ram[2][53] ) );
  DFFX1_HVT \ram_reg[2][52]  ( .D(n625), .CLK(clk), .Q(\ram[2][52] ) );
  DFFX1_HVT \ram_reg[2][51]  ( .D(n624), .CLK(clk), .Q(\ram[2][51] ) );
  DFFX1_HVT \ram_reg[2][50]  ( .D(n623), .CLK(clk), .Q(\ram[2][50] ) );
  DFFX1_HVT \ram_reg[2][49]  ( .D(n622), .CLK(clk), .Q(\ram[2][49] ) );
  DFFX1_HVT \ram_reg[2][48]  ( .D(n621), .CLK(clk), .Q(\ram[2][48] ) );
  DFFX1_HVT \ram_reg[2][47]  ( .D(n620), .CLK(clk), .Q(\ram[2][47] ) );
  DFFX1_HVT \ram_reg[2][46]  ( .D(n619), .CLK(clk), .Q(\ram[2][46] ) );
  DFFX1_HVT \ram_reg[2][45]  ( .D(n618), .CLK(clk), .Q(\ram[2][45] ) );
  DFFX1_HVT \ram_reg[2][44]  ( .D(n617), .CLK(clk), .Q(\ram[2][44] ) );
  DFFX1_HVT \ram_reg[2][43]  ( .D(n616), .CLK(clk), .Q(\ram[2][43] ) );
  DFFX1_HVT \ram_reg[2][42]  ( .D(n615), .CLK(clk), .Q(\ram[2][42] ) );
  DFFX1_HVT \ram_reg[2][41]  ( .D(n614), .CLK(clk), .Q(\ram[2][41] ) );
  DFFX1_HVT \ram_reg[2][40]  ( .D(n613), .CLK(clk), .Q(\ram[2][40] ) );
  DFFX1_HVT \ram_reg[2][39]  ( .D(n612), .CLK(clk), .Q(\ram[2][39] ) );
  DFFX1_HVT \ram_reg[2][38]  ( .D(n611), .CLK(clk), .Q(\ram[2][38] ) );
  DFFX1_HVT \ram_reg[2][37]  ( .D(n610), .CLK(clk), .Q(\ram[2][37] ) );
  DFFX1_HVT \ram_reg[2][36]  ( .D(n609), .CLK(clk), .Q(\ram[2][36] ) );
  DFFX1_HVT \ram_reg[2][35]  ( .D(n608), .CLK(clk), .Q(\ram[2][35] ) );
  DFFX1_HVT \ram_reg[2][34]  ( .D(n607), .CLK(clk), .Q(\ram[2][34] ) );
  DFFX1_HVT \ram_reg[2][33]  ( .D(n606), .CLK(clk), .Q(\ram[2][33] ) );
  DFFX1_HVT \ram_reg[2][32]  ( .D(n605), .CLK(clk), .Q(\ram[2][32] ) );
  DFFX1_HVT \ram_reg[2][31]  ( .D(n604), .CLK(clk), .Q(\ram[2][31] ) );
  DFFX1_HVT \ram_reg[2][30]  ( .D(n603), .CLK(clk), .Q(\ram[2][30] ) );
  DFFX1_HVT \ram_reg[2][29]  ( .D(n602), .CLK(clk), .Q(\ram[2][29] ) );
  DFFX1_HVT \ram_reg[2][28]  ( .D(n601), .CLK(clk), .Q(\ram[2][28] ) );
  DFFX1_HVT \ram_reg[2][27]  ( .D(n600), .CLK(clk), .Q(\ram[2][27] ) );
  DFFX1_HVT \ram_reg[2][26]  ( .D(n599), .CLK(clk), .Q(\ram[2][26] ) );
  DFFX1_HVT \ram_reg[2][25]  ( .D(n598), .CLK(clk), .Q(\ram[2][25] ) );
  DFFX1_HVT \ram_reg[2][24]  ( .D(n597), .CLK(clk), .Q(\ram[2][24] ) );
  DFFX1_HVT \ram_reg[2][23]  ( .D(n596), .CLK(clk), .Q(\ram[2][23] ) );
  DFFX1_HVT \ram_reg[2][22]  ( .D(n595), .CLK(clk), .Q(\ram[2][22] ) );
  DFFX1_HVT \ram_reg[2][21]  ( .D(n594), .CLK(clk), .Q(\ram[2][21] ) );
  DFFX1_HVT \ram_reg[2][20]  ( .D(n593), .CLK(clk), .Q(\ram[2][20] ) );
  DFFX1_HVT \ram_reg[2][19]  ( .D(n592), .CLK(clk), .Q(\ram[2][19] ) );
  DFFX1_HVT \ram_reg[2][18]  ( .D(n591), .CLK(clk), .Q(\ram[2][18] ) );
  DFFX1_HVT \ram_reg[2][17]  ( .D(n590), .CLK(clk), .Q(\ram[2][17] ) );
  DFFX1_HVT \ram_reg[2][16]  ( .D(n589), .CLK(clk), .Q(\ram[2][16] ) );
  DFFX1_HVT \ram_reg[2][15]  ( .D(n588), .CLK(clk), .Q(\ram[2][15] ) );
  DFFX1_HVT \ram_reg[2][14]  ( .D(n587), .CLK(clk), .Q(\ram[2][14] ) );
  DFFX1_HVT \ram_reg[2][13]  ( .D(n586), .CLK(clk), .Q(\ram[2][13] ) );
  DFFX1_HVT \ram_reg[2][12]  ( .D(n585), .CLK(clk), .Q(\ram[2][12] ) );
  DFFX1_HVT \ram_reg[2][11]  ( .D(n584), .CLK(clk), .Q(\ram[2][11] ) );
  DFFX1_HVT \ram_reg[2][10]  ( .D(n583), .CLK(clk), .Q(\ram[2][10] ) );
  DFFX1_HVT \ram_reg[2][9]  ( .D(n582), .CLK(clk), .Q(\ram[2][9] ) );
  DFFX1_HVT \ram_reg[2][8]  ( .D(n581), .CLK(clk), .Q(\ram[2][8] ) );
  DFFX1_HVT \ram_reg[2][7]  ( .D(n580), .CLK(clk), .Q(\ram[2][7] ) );
  DFFX1_HVT \ram_reg[2][6]  ( .D(n579), .CLK(clk), .Q(\ram[2][6] ) );
  DFFX1_HVT \ram_reg[2][5]  ( .D(n578), .CLK(clk), .Q(\ram[2][5] ) );
  DFFX1_HVT \ram_reg[2][4]  ( .D(n577), .CLK(clk), .Q(\ram[2][4] ) );
  DFFX1_HVT \ram_reg[2][3]  ( .D(n576), .CLK(clk), .Q(\ram[2][3] ) );
  DFFX1_HVT \ram_reg[2][2]  ( .D(n575), .CLK(clk), .Q(\ram[2][2] ) );
  DFFX1_HVT \ram_reg[2][1]  ( .D(n574), .CLK(clk), .Q(\ram[2][1] ) );
  DFFX1_HVT \ram_reg[2][0]  ( .D(n573), .CLK(clk), .Q(\ram[2][0] ) );
  DFFX1_HVT \ram_reg[1][255]  ( .D(n572), .CLK(clk), .Q(\ram[1][255] ) );
  DFFX1_HVT \ram_reg[1][254]  ( .D(n571), .CLK(clk), .Q(\ram[1][254] ) );
  DFFX1_HVT \ram_reg[1][253]  ( .D(n570), .CLK(clk), .Q(\ram[1][253] ) );
  DFFX1_HVT \ram_reg[1][252]  ( .D(n569), .CLK(clk), .Q(\ram[1][252] ) );
  DFFX1_HVT \ram_reg[1][251]  ( .D(n568), .CLK(clk), .Q(\ram[1][251] ) );
  DFFX1_HVT \ram_reg[1][250]  ( .D(n567), .CLK(clk), .Q(\ram[1][250] ) );
  DFFX1_HVT \ram_reg[1][249]  ( .D(n566), .CLK(clk), .Q(\ram[1][249] ) );
  DFFX1_HVT \ram_reg[1][248]  ( .D(n565), .CLK(clk), .Q(\ram[1][248] ) );
  DFFX1_HVT \ram_reg[1][247]  ( .D(n564), .CLK(clk), .Q(\ram[1][247] ) );
  DFFX1_HVT \ram_reg[1][246]  ( .D(n563), .CLK(clk), .Q(\ram[1][246] ) );
  DFFX1_HVT \ram_reg[1][245]  ( .D(n562), .CLK(clk), .Q(\ram[1][245] ) );
  DFFX1_HVT \ram_reg[1][244]  ( .D(n561), .CLK(clk), .Q(\ram[1][244] ) );
  DFFX1_HVT \ram_reg[1][243]  ( .D(n560), .CLK(clk), .Q(\ram[1][243] ) );
  DFFX1_HVT \ram_reg[1][242]  ( .D(n559), .CLK(clk), .Q(\ram[1][242] ) );
  DFFX1_HVT \ram_reg[1][241]  ( .D(n558), .CLK(clk), .Q(\ram[1][241] ) );
  DFFX1_HVT \ram_reg[1][240]  ( .D(n557), .CLK(clk), .Q(\ram[1][240] ) );
  DFFX1_HVT \ram_reg[1][239]  ( .D(n556), .CLK(clk), .Q(\ram[1][239] ) );
  DFFX1_HVT \ram_reg[1][238]  ( .D(n555), .CLK(clk), .Q(\ram[1][238] ) );
  DFFX1_HVT \ram_reg[1][237]  ( .D(n554), .CLK(clk), .Q(\ram[1][237] ) );
  DFFX1_HVT \ram_reg[1][236]  ( .D(n553), .CLK(clk), .Q(\ram[1][236] ) );
  DFFX1_HVT \ram_reg[1][235]  ( .D(n552), .CLK(clk), .Q(\ram[1][235] ) );
  DFFX1_HVT \ram_reg[1][234]  ( .D(n551), .CLK(clk), .Q(\ram[1][234] ) );
  DFFX1_HVT \ram_reg[1][233]  ( .D(n550), .CLK(clk), .Q(\ram[1][233] ) );
  DFFX1_HVT \ram_reg[1][232]  ( .D(n549), .CLK(clk), .Q(\ram[1][232] ) );
  DFFX1_HVT \ram_reg[1][231]  ( .D(n548), .CLK(clk), .Q(\ram[1][231] ) );
  DFFX1_HVT \ram_reg[1][230]  ( .D(n547), .CLK(clk), .Q(\ram[1][230] ) );
  DFFX1_HVT \ram_reg[1][229]  ( .D(n546), .CLK(clk), .Q(\ram[1][229] ) );
  DFFX1_HVT \ram_reg[1][228]  ( .D(n545), .CLK(clk), .Q(\ram[1][228] ) );
  DFFX1_HVT \ram_reg[1][227]  ( .D(n544), .CLK(clk), .Q(\ram[1][227] ) );
  DFFX1_HVT \ram_reg[1][226]  ( .D(n543), .CLK(clk), .Q(\ram[1][226] ) );
  DFFX1_HVT \ram_reg[1][225]  ( .D(n542), .CLK(clk), .Q(\ram[1][225] ) );
  DFFX1_HVT \ram_reg[1][224]  ( .D(n541), .CLK(clk), .Q(\ram[1][224] ) );
  DFFX1_HVT \ram_reg[1][223]  ( .D(n540), .CLK(clk), .Q(\ram[1][223] ) );
  DFFX1_HVT \ram_reg[1][222]  ( .D(n539), .CLK(clk), .Q(\ram[1][222] ) );
  DFFX1_HVT \ram_reg[1][221]  ( .D(n538), .CLK(clk), .Q(\ram[1][221] ) );
  DFFX1_HVT \ram_reg[1][220]  ( .D(n537), .CLK(clk), .Q(\ram[1][220] ) );
  DFFX1_HVT \ram_reg[1][219]  ( .D(n536), .CLK(clk), .Q(\ram[1][219] ) );
  DFFX1_HVT \ram_reg[1][218]  ( .D(n535), .CLK(clk), .Q(\ram[1][218] ) );
  DFFX1_HVT \ram_reg[1][217]  ( .D(n534), .CLK(clk), .Q(\ram[1][217] ) );
  DFFX1_HVT \ram_reg[1][216]  ( .D(n533), .CLK(clk), .Q(\ram[1][216] ) );
  DFFX1_HVT \ram_reg[1][215]  ( .D(n532), .CLK(clk), .Q(\ram[1][215] ) );
  DFFX1_HVT \ram_reg[1][214]  ( .D(n531), .CLK(clk), .Q(\ram[1][214] ) );
  DFFX1_HVT \ram_reg[1][213]  ( .D(n530), .CLK(clk), .Q(\ram[1][213] ) );
  DFFX1_HVT \ram_reg[1][212]  ( .D(n529), .CLK(clk), .Q(\ram[1][212] ) );
  DFFX1_HVT \ram_reg[1][211]  ( .D(n528), .CLK(clk), .Q(\ram[1][211] ) );
  DFFX1_HVT \ram_reg[1][210]  ( .D(n527), .CLK(clk), .Q(\ram[1][210] ) );
  DFFX1_HVT \ram_reg[1][209]  ( .D(n526), .CLK(clk), .Q(\ram[1][209] ) );
  DFFX1_HVT \ram_reg[1][208]  ( .D(n525), .CLK(clk), .Q(\ram[1][208] ) );
  DFFX1_HVT \ram_reg[1][207]  ( .D(n524), .CLK(clk), .Q(\ram[1][207] ) );
  DFFX1_HVT \ram_reg[1][206]  ( .D(n523), .CLK(clk), .Q(\ram[1][206] ) );
  DFFX1_HVT \ram_reg[1][205]  ( .D(n522), .CLK(clk), .Q(\ram[1][205] ) );
  DFFX1_HVT \ram_reg[1][204]  ( .D(n521), .CLK(clk), .Q(\ram[1][204] ) );
  DFFX1_HVT \ram_reg[1][203]  ( .D(n520), .CLK(clk), .Q(\ram[1][203] ) );
  DFFX1_HVT \ram_reg[1][202]  ( .D(n519), .CLK(clk), .Q(\ram[1][202] ) );
  DFFX1_HVT \ram_reg[1][201]  ( .D(n518), .CLK(clk), .Q(\ram[1][201] ) );
  DFFX1_HVT \ram_reg[1][200]  ( .D(n517), .CLK(clk), .Q(\ram[1][200] ) );
  DFFX1_HVT \ram_reg[1][199]  ( .D(n516), .CLK(clk), .Q(\ram[1][199] ) );
  DFFX1_HVT \ram_reg[1][198]  ( .D(n515), .CLK(clk), .Q(\ram[1][198] ) );
  DFFX1_HVT \ram_reg[1][197]  ( .D(n514), .CLK(clk), .Q(\ram[1][197] ) );
  DFFX1_HVT \ram_reg[1][196]  ( .D(n513), .CLK(clk), .Q(\ram[1][196] ) );
  DFFX1_HVT \ram_reg[1][195]  ( .D(n512), .CLK(clk), .Q(\ram[1][195] ) );
  DFFX1_HVT \ram_reg[1][194]  ( .D(n511), .CLK(clk), .Q(\ram[1][194] ) );
  DFFX1_HVT \ram_reg[1][193]  ( .D(n510), .CLK(clk), .Q(\ram[1][193] ) );
  DFFX1_HVT \ram_reg[1][192]  ( .D(n509), .CLK(clk), .Q(\ram[1][192] ) );
  DFFX1_HVT \ram_reg[1][191]  ( .D(n508), .CLK(clk), .Q(\ram[1][191] ) );
  DFFX1_HVT \ram_reg[1][190]  ( .D(n507), .CLK(clk), .Q(\ram[1][190] ) );
  DFFX1_HVT \ram_reg[1][189]  ( .D(n506), .CLK(clk), .Q(\ram[1][189] ) );
  DFFX1_HVT \ram_reg[1][188]  ( .D(n505), .CLK(clk), .Q(\ram[1][188] ) );
  DFFX1_HVT \ram_reg[1][187]  ( .D(n504), .CLK(clk), .Q(\ram[1][187] ) );
  DFFX1_HVT \ram_reg[1][186]  ( .D(n503), .CLK(clk), .Q(\ram[1][186] ) );
  DFFX1_HVT \ram_reg[1][185]  ( .D(n502), .CLK(clk), .Q(\ram[1][185] ) );
  DFFX1_HVT \ram_reg[1][184]  ( .D(n501), .CLK(clk), .Q(\ram[1][184] ) );
  DFFX1_HVT \ram_reg[1][183]  ( .D(n500), .CLK(clk), .Q(\ram[1][183] ) );
  DFFX1_HVT \ram_reg[1][182]  ( .D(n499), .CLK(clk), .Q(\ram[1][182] ) );
  DFFX1_HVT \ram_reg[1][181]  ( .D(n498), .CLK(clk), .Q(\ram[1][181] ) );
  DFFX1_HVT \ram_reg[1][180]  ( .D(n497), .CLK(clk), .Q(\ram[1][180] ) );
  DFFX1_HVT \ram_reg[1][179]  ( .D(n496), .CLK(clk), .Q(\ram[1][179] ) );
  DFFX1_HVT \ram_reg[1][178]  ( .D(n495), .CLK(clk), .Q(\ram[1][178] ) );
  DFFX1_HVT \ram_reg[1][177]  ( .D(n494), .CLK(clk), .Q(\ram[1][177] ) );
  DFFX1_HVT \ram_reg[1][176]  ( .D(n493), .CLK(clk), .Q(\ram[1][176] ) );
  DFFX1_HVT \ram_reg[1][175]  ( .D(n492), .CLK(clk), .Q(\ram[1][175] ) );
  DFFX1_HVT \ram_reg[1][174]  ( .D(n491), .CLK(clk), .Q(\ram[1][174] ) );
  DFFX1_HVT \ram_reg[1][173]  ( .D(n490), .CLK(clk), .Q(\ram[1][173] ) );
  DFFX1_HVT \ram_reg[1][172]  ( .D(n489), .CLK(clk), .Q(\ram[1][172] ) );
  DFFX1_HVT \ram_reg[1][171]  ( .D(n488), .CLK(clk), .Q(\ram[1][171] ) );
  DFFX1_HVT \ram_reg[1][170]  ( .D(n487), .CLK(clk), .Q(\ram[1][170] ) );
  DFFX1_HVT \ram_reg[1][169]  ( .D(n486), .CLK(clk), .Q(\ram[1][169] ) );
  DFFX1_HVT \ram_reg[1][168]  ( .D(n485), .CLK(clk), .Q(\ram[1][168] ) );
  DFFX1_HVT \ram_reg[1][167]  ( .D(n484), .CLK(clk), .Q(\ram[1][167] ) );
  DFFX1_HVT \ram_reg[1][166]  ( .D(n483), .CLK(clk), .Q(\ram[1][166] ) );
  DFFX1_HVT \ram_reg[1][165]  ( .D(n482), .CLK(clk), .Q(\ram[1][165] ) );
  DFFX1_HVT \ram_reg[1][164]  ( .D(n481), .CLK(clk), .Q(\ram[1][164] ) );
  DFFX1_HVT \ram_reg[1][163]  ( .D(n480), .CLK(clk), .Q(\ram[1][163] ) );
  DFFX1_HVT \ram_reg[1][162]  ( .D(n479), .CLK(clk), .Q(\ram[1][162] ) );
  DFFX1_HVT \ram_reg[1][161]  ( .D(n478), .CLK(clk), .Q(\ram[1][161] ) );
  DFFX1_HVT \ram_reg[1][160]  ( .D(n477), .CLK(clk), .Q(\ram[1][160] ) );
  DFFX1_HVT \ram_reg[1][159]  ( .D(n476), .CLK(clk), .Q(\ram[1][159] ) );
  DFFX1_HVT \ram_reg[1][158]  ( .D(n475), .CLK(clk), .Q(\ram[1][158] ) );
  DFFX1_HVT \ram_reg[1][157]  ( .D(n474), .CLK(clk), .Q(\ram[1][157] ) );
  DFFX1_HVT \ram_reg[1][156]  ( .D(n473), .CLK(clk), .Q(\ram[1][156] ) );
  DFFX1_HVT \ram_reg[1][155]  ( .D(n472), .CLK(clk), .Q(\ram[1][155] ) );
  DFFX1_HVT \ram_reg[1][154]  ( .D(n471), .CLK(clk), .Q(\ram[1][154] ) );
  DFFX1_HVT \ram_reg[1][153]  ( .D(n470), .CLK(clk), .Q(\ram[1][153] ) );
  DFFX1_HVT \ram_reg[1][152]  ( .D(n469), .CLK(clk), .Q(\ram[1][152] ) );
  DFFX1_HVT \ram_reg[1][151]  ( .D(n468), .CLK(clk), .Q(\ram[1][151] ) );
  DFFX1_HVT \ram_reg[1][150]  ( .D(n467), .CLK(clk), .Q(\ram[1][150] ) );
  DFFX1_HVT \ram_reg[1][149]  ( .D(n466), .CLK(clk), .Q(\ram[1][149] ) );
  DFFX1_HVT \ram_reg[1][148]  ( .D(n465), .CLK(clk), .Q(\ram[1][148] ) );
  DFFX1_HVT \ram_reg[1][147]  ( .D(n464), .CLK(clk), .Q(\ram[1][147] ) );
  DFFX1_HVT \ram_reg[1][146]  ( .D(n463), .CLK(clk), .Q(\ram[1][146] ) );
  DFFX1_HVT \ram_reg[1][145]  ( .D(n462), .CLK(clk), .Q(\ram[1][145] ) );
  DFFX1_HVT \ram_reg[1][144]  ( .D(n461), .CLK(clk), .Q(\ram[1][144] ) );
  DFFX1_HVT \ram_reg[1][143]  ( .D(n460), .CLK(clk), .Q(\ram[1][143] ) );
  DFFX1_HVT \ram_reg[1][142]  ( .D(n459), .CLK(clk), .Q(\ram[1][142] ) );
  DFFX1_HVT \ram_reg[1][141]  ( .D(n458), .CLK(clk), .Q(\ram[1][141] ) );
  DFFX1_HVT \ram_reg[1][140]  ( .D(n457), .CLK(clk), .Q(\ram[1][140] ) );
  DFFX1_HVT \ram_reg[1][139]  ( .D(n456), .CLK(clk), .Q(\ram[1][139] ) );
  DFFX1_HVT \ram_reg[1][138]  ( .D(n455), .CLK(clk), .Q(\ram[1][138] ) );
  DFFX1_HVT \ram_reg[1][137]  ( .D(n454), .CLK(clk), .Q(\ram[1][137] ) );
  DFFX1_HVT \ram_reg[1][136]  ( .D(n453), .CLK(clk), .Q(\ram[1][136] ) );
  DFFX1_HVT \ram_reg[1][135]  ( .D(n452), .CLK(clk), .Q(\ram[1][135] ) );
  DFFX1_HVT \ram_reg[1][134]  ( .D(n451), .CLK(clk), .Q(\ram[1][134] ) );
  DFFX1_HVT \ram_reg[1][133]  ( .D(n450), .CLK(clk), .Q(\ram[1][133] ) );
  DFFX1_HVT \ram_reg[1][132]  ( .D(n449), .CLK(clk), .Q(\ram[1][132] ) );
  DFFX1_HVT \ram_reg[1][131]  ( .D(n448), .CLK(clk), .Q(\ram[1][131] ) );
  DFFX1_HVT \ram_reg[1][130]  ( .D(n447), .CLK(clk), .Q(\ram[1][130] ) );
  DFFX1_HVT \ram_reg[1][129]  ( .D(n446), .CLK(clk), .Q(\ram[1][129] ) );
  DFFX1_HVT \ram_reg[1][128]  ( .D(n445), .CLK(clk), .Q(\ram[1][128] ) );
  DFFX1_HVT \ram_reg[1][127]  ( .D(n444), .CLK(clk), .Q(\ram[1][127] ) );
  DFFX1_HVT \ram_reg[1][126]  ( .D(n443), .CLK(clk), .Q(\ram[1][126] ) );
  DFFX1_HVT \ram_reg[1][125]  ( .D(n442), .CLK(clk), .Q(\ram[1][125] ) );
  DFFX1_HVT \ram_reg[1][124]  ( .D(n441), .CLK(clk), .Q(\ram[1][124] ) );
  DFFX1_HVT \ram_reg[1][123]  ( .D(n440), .CLK(clk), .Q(\ram[1][123] ) );
  DFFX1_HVT \ram_reg[1][122]  ( .D(n439), .CLK(clk), .Q(\ram[1][122] ) );
  DFFX1_HVT \ram_reg[1][121]  ( .D(n438), .CLK(clk), .Q(\ram[1][121] ) );
  DFFX1_HVT \ram_reg[1][120]  ( .D(n437), .CLK(clk), .Q(\ram[1][120] ) );
  DFFX1_HVT \ram_reg[1][119]  ( .D(n436), .CLK(clk), .Q(\ram[1][119] ) );
  DFFX1_HVT \ram_reg[1][118]  ( .D(n435), .CLK(clk), .Q(\ram[1][118] ) );
  DFFX1_HVT \ram_reg[1][117]  ( .D(n434), .CLK(clk), .Q(\ram[1][117] ) );
  DFFX1_HVT \ram_reg[1][116]  ( .D(n433), .CLK(clk), .Q(\ram[1][116] ) );
  DFFX1_HVT \ram_reg[1][115]  ( .D(n432), .CLK(clk), .Q(\ram[1][115] ) );
  DFFX1_HVT \ram_reg[1][114]  ( .D(n431), .CLK(clk), .Q(\ram[1][114] ) );
  DFFX1_HVT \ram_reg[1][113]  ( .D(n430), .CLK(clk), .Q(\ram[1][113] ) );
  DFFX1_HVT \ram_reg[1][112]  ( .D(n429), .CLK(clk), .Q(\ram[1][112] ) );
  DFFX1_HVT \ram_reg[1][111]  ( .D(n428), .CLK(clk), .Q(\ram[1][111] ) );
  DFFX1_HVT \ram_reg[1][110]  ( .D(n427), .CLK(clk), .Q(\ram[1][110] ) );
  DFFX1_HVT \ram_reg[1][109]  ( .D(n426), .CLK(clk), .Q(\ram[1][109] ) );
  DFFX1_HVT \ram_reg[1][108]  ( .D(n425), .CLK(clk), .Q(\ram[1][108] ) );
  DFFX1_HVT \ram_reg[1][107]  ( .D(n424), .CLK(clk), .Q(\ram[1][107] ) );
  DFFX1_HVT \ram_reg[1][106]  ( .D(n423), .CLK(clk), .Q(\ram[1][106] ) );
  DFFX1_HVT \ram_reg[1][105]  ( .D(n422), .CLK(clk), .Q(\ram[1][105] ) );
  DFFX1_HVT \ram_reg[1][104]  ( .D(n421), .CLK(clk), .Q(\ram[1][104] ) );
  DFFX1_HVT \ram_reg[1][103]  ( .D(n420), .CLK(clk), .Q(\ram[1][103] ) );
  DFFX1_HVT \ram_reg[1][102]  ( .D(n419), .CLK(clk), .Q(\ram[1][102] ) );
  DFFX1_HVT \ram_reg[1][101]  ( .D(n418), .CLK(clk), .Q(\ram[1][101] ) );
  DFFX1_HVT \ram_reg[1][100]  ( .D(n417), .CLK(clk), .Q(\ram[1][100] ) );
  DFFX1_HVT \ram_reg[1][99]  ( .D(n416), .CLK(clk), .Q(\ram[1][99] ) );
  DFFX1_HVT \ram_reg[1][98]  ( .D(n415), .CLK(clk), .Q(\ram[1][98] ) );
  DFFX1_HVT \ram_reg[1][97]  ( .D(n414), .CLK(clk), .Q(\ram[1][97] ) );
  DFFX1_HVT \ram_reg[1][96]  ( .D(n413), .CLK(clk), .Q(\ram[1][96] ) );
  DFFX1_HVT \ram_reg[1][95]  ( .D(n412), .CLK(clk), .Q(\ram[1][95] ) );
  DFFX1_HVT \ram_reg[1][94]  ( .D(n411), .CLK(clk), .Q(\ram[1][94] ) );
  DFFX1_HVT \ram_reg[1][93]  ( .D(n410), .CLK(clk), .Q(\ram[1][93] ) );
  DFFX1_HVT \ram_reg[1][92]  ( .D(n409), .CLK(clk), .Q(\ram[1][92] ) );
  DFFX1_HVT \ram_reg[1][91]  ( .D(n408), .CLK(clk), .Q(\ram[1][91] ) );
  DFFX1_HVT \ram_reg[1][90]  ( .D(n407), .CLK(clk), .Q(\ram[1][90] ) );
  DFFX1_HVT \ram_reg[1][89]  ( .D(n406), .CLK(clk), .Q(\ram[1][89] ) );
  DFFX1_HVT \ram_reg[1][88]  ( .D(n405), .CLK(clk), .Q(\ram[1][88] ) );
  DFFX1_HVT \ram_reg[1][87]  ( .D(n404), .CLK(clk), .Q(\ram[1][87] ) );
  DFFX1_HVT \ram_reg[1][86]  ( .D(n403), .CLK(clk), .Q(\ram[1][86] ) );
  DFFX1_HVT \ram_reg[1][85]  ( .D(n402), .CLK(clk), .Q(\ram[1][85] ) );
  DFFX1_HVT \ram_reg[1][84]  ( .D(n401), .CLK(clk), .Q(\ram[1][84] ) );
  DFFX1_HVT \ram_reg[1][83]  ( .D(n400), .CLK(clk), .Q(\ram[1][83] ) );
  DFFX1_HVT \ram_reg[1][82]  ( .D(n399), .CLK(clk), .Q(\ram[1][82] ) );
  DFFX1_HVT \ram_reg[1][81]  ( .D(n398), .CLK(clk), .Q(\ram[1][81] ) );
  DFFX1_HVT \ram_reg[1][80]  ( .D(n397), .CLK(clk), .Q(\ram[1][80] ) );
  DFFX1_HVT \ram_reg[1][79]  ( .D(n396), .CLK(clk), .Q(\ram[1][79] ) );
  DFFX1_HVT \ram_reg[1][78]  ( .D(n395), .CLK(clk), .Q(\ram[1][78] ) );
  DFFX1_HVT \ram_reg[1][77]  ( .D(n394), .CLK(clk), .Q(\ram[1][77] ) );
  DFFX1_HVT \ram_reg[1][76]  ( .D(n393), .CLK(clk), .Q(\ram[1][76] ) );
  DFFX1_HVT \ram_reg[1][75]  ( .D(n392), .CLK(clk), .Q(\ram[1][75] ) );
  DFFX1_HVT \ram_reg[1][74]  ( .D(n391), .CLK(clk), .Q(\ram[1][74] ) );
  DFFX1_HVT \ram_reg[1][73]  ( .D(n390), .CLK(clk), .Q(\ram[1][73] ) );
  DFFX1_HVT \ram_reg[1][72]  ( .D(n389), .CLK(clk), .Q(\ram[1][72] ) );
  DFFX1_HVT \ram_reg[1][71]  ( .D(n388), .CLK(clk), .Q(\ram[1][71] ) );
  DFFX1_HVT \ram_reg[1][70]  ( .D(n387), .CLK(clk), .Q(\ram[1][70] ) );
  DFFX1_HVT \ram_reg[1][69]  ( .D(n386), .CLK(clk), .Q(\ram[1][69] ) );
  DFFX1_HVT \ram_reg[1][68]  ( .D(n385), .CLK(clk), .Q(\ram[1][68] ) );
  DFFX1_HVT \ram_reg[1][67]  ( .D(n384), .CLK(clk), .Q(\ram[1][67] ) );
  DFFX1_HVT \ram_reg[1][66]  ( .D(n383), .CLK(clk), .Q(\ram[1][66] ) );
  DFFX1_HVT \ram_reg[1][65]  ( .D(n382), .CLK(clk), .Q(\ram[1][65] ) );
  DFFX1_HVT \ram_reg[1][64]  ( .D(n381), .CLK(clk), .Q(\ram[1][64] ) );
  DFFX1_HVT \ram_reg[1][63]  ( .D(n380), .CLK(clk), .Q(\ram[1][63] ) );
  DFFX1_HVT \ram_reg[1][62]  ( .D(n379), .CLK(clk), .Q(\ram[1][62] ) );
  DFFX1_HVT \ram_reg[1][61]  ( .D(n378), .CLK(clk), .Q(\ram[1][61] ) );
  DFFX1_HVT \ram_reg[1][60]  ( .D(n377), .CLK(clk), .Q(\ram[1][60] ) );
  DFFX1_HVT \ram_reg[1][59]  ( .D(n376), .CLK(clk), .Q(\ram[1][59] ) );
  DFFX1_HVT \ram_reg[1][58]  ( .D(n375), .CLK(clk), .Q(\ram[1][58] ) );
  DFFX1_HVT \ram_reg[1][57]  ( .D(n374), .CLK(clk), .Q(\ram[1][57] ) );
  DFFX1_HVT \ram_reg[1][56]  ( .D(n373), .CLK(clk), .Q(\ram[1][56] ) );
  DFFX1_HVT \ram_reg[1][55]  ( .D(n372), .CLK(clk), .Q(\ram[1][55] ) );
  DFFX1_HVT \ram_reg[1][54]  ( .D(n371), .CLK(clk), .Q(\ram[1][54] ) );
  DFFX1_HVT \ram_reg[1][53]  ( .D(n370), .CLK(clk), .Q(\ram[1][53] ) );
  DFFX1_HVT \ram_reg[1][52]  ( .D(n369), .CLK(clk), .Q(\ram[1][52] ) );
  DFFX1_HVT \ram_reg[1][51]  ( .D(n368), .CLK(clk), .Q(\ram[1][51] ) );
  DFFX1_HVT \ram_reg[1][50]  ( .D(n367), .CLK(clk), .Q(\ram[1][50] ) );
  DFFX1_HVT \ram_reg[1][49]  ( .D(n366), .CLK(clk), .Q(\ram[1][49] ) );
  DFFX1_HVT \ram_reg[1][48]  ( .D(n365), .CLK(clk), .Q(\ram[1][48] ) );
  DFFX1_HVT \ram_reg[1][47]  ( .D(n364), .CLK(clk), .Q(\ram[1][47] ) );
  DFFX1_HVT \ram_reg[1][46]  ( .D(n363), .CLK(clk), .Q(\ram[1][46] ) );
  DFFX1_HVT \ram_reg[1][45]  ( .D(n362), .CLK(clk), .Q(\ram[1][45] ) );
  DFFX1_HVT \ram_reg[1][44]  ( .D(n361), .CLK(clk), .Q(\ram[1][44] ) );
  DFFX1_HVT \ram_reg[1][43]  ( .D(n360), .CLK(clk), .Q(\ram[1][43] ) );
  DFFX1_HVT \ram_reg[1][42]  ( .D(n359), .CLK(clk), .Q(\ram[1][42] ) );
  DFFX1_HVT \ram_reg[1][41]  ( .D(n358), .CLK(clk), .Q(\ram[1][41] ) );
  DFFX1_HVT \ram_reg[1][40]  ( .D(n357), .CLK(clk), .Q(\ram[1][40] ) );
  DFFX1_HVT \ram_reg[1][39]  ( .D(n356), .CLK(clk), .Q(\ram[1][39] ) );
  DFFX1_HVT \ram_reg[1][38]  ( .D(n355), .CLK(clk), .Q(\ram[1][38] ) );
  DFFX1_HVT \ram_reg[1][37]  ( .D(n354), .CLK(clk), .Q(\ram[1][37] ) );
  DFFX1_HVT \ram_reg[1][36]  ( .D(n353), .CLK(clk), .Q(\ram[1][36] ) );
  DFFX1_HVT \ram_reg[1][35]  ( .D(n352), .CLK(clk), .Q(\ram[1][35] ) );
  DFFX1_HVT \ram_reg[1][34]  ( .D(n351), .CLK(clk), .Q(\ram[1][34] ) );
  DFFX1_HVT \ram_reg[1][33]  ( .D(n350), .CLK(clk), .Q(\ram[1][33] ) );
  DFFX1_HVT \ram_reg[1][32]  ( .D(n349), .CLK(clk), .Q(\ram[1][32] ) );
  DFFX1_HVT \ram_reg[1][31]  ( .D(n348), .CLK(clk), .Q(\ram[1][31] ) );
  DFFX1_HVT \ram_reg[1][30]  ( .D(n347), .CLK(clk), .Q(\ram[1][30] ) );
  DFFX1_HVT \ram_reg[1][29]  ( .D(n346), .CLK(clk), .Q(\ram[1][29] ) );
  DFFX1_HVT \ram_reg[1][28]  ( .D(n345), .CLK(clk), .Q(\ram[1][28] ) );
  DFFX1_HVT \ram_reg[1][27]  ( .D(n344), .CLK(clk), .Q(\ram[1][27] ) );
  DFFX1_HVT \ram_reg[1][26]  ( .D(n343), .CLK(clk), .Q(\ram[1][26] ) );
  DFFX1_HVT \ram_reg[1][25]  ( .D(n342), .CLK(clk), .Q(\ram[1][25] ) );
  DFFX1_HVT \ram_reg[1][24]  ( .D(n341), .CLK(clk), .Q(\ram[1][24] ) );
  DFFX1_HVT \ram_reg[1][23]  ( .D(n340), .CLK(clk), .Q(\ram[1][23] ) );
  DFFX1_HVT \ram_reg[1][22]  ( .D(n339), .CLK(clk), .Q(\ram[1][22] ) );
  DFFX1_HVT \ram_reg[1][21]  ( .D(n338), .CLK(clk), .Q(\ram[1][21] ) );
  DFFX1_HVT \ram_reg[1][20]  ( .D(n337), .CLK(clk), .Q(\ram[1][20] ) );
  DFFX1_HVT \ram_reg[1][19]  ( .D(n336), .CLK(clk), .Q(\ram[1][19] ) );
  DFFX1_HVT \ram_reg[1][18]  ( .D(n335), .CLK(clk), .Q(\ram[1][18] ) );
  DFFX1_HVT \ram_reg[1][17]  ( .D(n334), .CLK(clk), .Q(\ram[1][17] ) );
  DFFX1_HVT \ram_reg[1][16]  ( .D(n333), .CLK(clk), .Q(\ram[1][16] ) );
  DFFX1_HVT \ram_reg[1][15]  ( .D(n332), .CLK(clk), .Q(\ram[1][15] ) );
  DFFX1_HVT \ram_reg[1][14]  ( .D(n331), .CLK(clk), .Q(\ram[1][14] ) );
  DFFX1_HVT \ram_reg[1][13]  ( .D(n330), .CLK(clk), .Q(\ram[1][13] ) );
  DFFX1_HVT \ram_reg[1][12]  ( .D(n329), .CLK(clk), .Q(\ram[1][12] ) );
  DFFX1_HVT \ram_reg[1][11]  ( .D(n328), .CLK(clk), .Q(\ram[1][11] ) );
  DFFX1_HVT \ram_reg[1][10]  ( .D(n327), .CLK(clk), .Q(\ram[1][10] ) );
  DFFX1_HVT \ram_reg[1][9]  ( .D(n326), .CLK(clk), .Q(\ram[1][9] ) );
  DFFX1_HVT \ram_reg[1][8]  ( .D(n325), .CLK(clk), .Q(\ram[1][8] ) );
  DFFX1_HVT \ram_reg[1][7]  ( .D(n324), .CLK(clk), .Q(\ram[1][7] ) );
  DFFX1_HVT \ram_reg[1][6]  ( .D(n323), .CLK(clk), .Q(\ram[1][6] ) );
  DFFX1_HVT \ram_reg[1][5]  ( .D(n322), .CLK(clk), .Q(\ram[1][5] ) );
  DFFX1_HVT \ram_reg[1][4]  ( .D(n321), .CLK(clk), .Q(\ram[1][4] ) );
  DFFX1_HVT \ram_reg[1][3]  ( .D(n320), .CLK(clk), .Q(\ram[1][3] ) );
  DFFX1_HVT \ram_reg[1][2]  ( .D(n319), .CLK(clk), .Q(\ram[1][2] ) );
  DFFX1_HVT \ram_reg[1][1]  ( .D(n318), .CLK(clk), .Q(\ram[1][1] ) );
  DFFX1_HVT \ram_reg[1][0]  ( .D(n317), .CLK(clk), .Q(\ram[1][0] ) );
  DFFX1_HVT \ram_reg[0][255]  ( .D(n316), .CLK(clk), .Q(\ram[0][255] ) );
  DFFX1_HVT \ram_reg[0][254]  ( .D(n315), .CLK(clk), .Q(\ram[0][254] ) );
  DFFX1_HVT \ram_reg[0][253]  ( .D(n314), .CLK(clk), .Q(\ram[0][253] ) );
  DFFX1_HVT \ram_reg[0][252]  ( .D(n313), .CLK(clk), .Q(\ram[0][252] ) );
  DFFX1_HVT \ram_reg[0][251]  ( .D(n312), .CLK(clk), .Q(\ram[0][251] ) );
  DFFX1_HVT \ram_reg[0][250]  ( .D(n311), .CLK(clk), .Q(\ram[0][250] ) );
  DFFX1_HVT \ram_reg[0][249]  ( .D(n310), .CLK(clk), .Q(\ram[0][249] ) );
  DFFX1_HVT \ram_reg[0][248]  ( .D(n309), .CLK(clk), .Q(\ram[0][248] ) );
  DFFX1_HVT \ram_reg[0][247]  ( .D(n308), .CLK(clk), .Q(\ram[0][247] ) );
  DFFX1_HVT \ram_reg[0][246]  ( .D(n307), .CLK(clk), .Q(\ram[0][246] ) );
  DFFX1_HVT \ram_reg[0][245]  ( .D(n306), .CLK(clk), .Q(\ram[0][245] ) );
  DFFX1_HVT \ram_reg[0][244]  ( .D(n305), .CLK(clk), .Q(\ram[0][244] ) );
  DFFX1_HVT \ram_reg[0][243]  ( .D(n304), .CLK(clk), .Q(\ram[0][243] ) );
  DFFX1_HVT \ram_reg[0][242]  ( .D(n303), .CLK(clk), .Q(\ram[0][242] ) );
  DFFX1_HVT \ram_reg[0][241]  ( .D(n302), .CLK(clk), .Q(\ram[0][241] ) );
  DFFX1_HVT \ram_reg[0][240]  ( .D(n301), .CLK(clk), .Q(\ram[0][240] ) );
  DFFX1_HVT \ram_reg[0][239]  ( .D(n300), .CLK(clk), .Q(\ram[0][239] ) );
  DFFX1_HVT \ram_reg[0][238]  ( .D(n299), .CLK(clk), .Q(\ram[0][238] ) );
  DFFX1_HVT \ram_reg[0][237]  ( .D(n298), .CLK(clk), .Q(\ram[0][237] ) );
  DFFX1_HVT \ram_reg[0][236]  ( .D(n297), .CLK(clk), .Q(\ram[0][236] ) );
  DFFX1_HVT \ram_reg[0][235]  ( .D(n296), .CLK(clk), .Q(\ram[0][235] ) );
  DFFX1_HVT \ram_reg[0][234]  ( .D(n295), .CLK(clk), .Q(\ram[0][234] ) );
  DFFX1_HVT \ram_reg[0][233]  ( .D(n294), .CLK(clk), .Q(\ram[0][233] ) );
  DFFX1_HVT \ram_reg[0][232]  ( .D(n293), .CLK(clk), .Q(\ram[0][232] ) );
  DFFX1_HVT \ram_reg[0][231]  ( .D(n292), .CLK(clk), .Q(\ram[0][231] ) );
  DFFX1_HVT \ram_reg[0][230]  ( .D(n291), .CLK(clk), .Q(\ram[0][230] ) );
  DFFX1_HVT \ram_reg[0][229]  ( .D(n290), .CLK(clk), .Q(\ram[0][229] ) );
  DFFX1_HVT \ram_reg[0][228]  ( .D(n289), .CLK(clk), .Q(\ram[0][228] ) );
  DFFX1_HVT \ram_reg[0][227]  ( .D(n288), .CLK(clk), .Q(\ram[0][227] ) );
  DFFX1_HVT \ram_reg[0][226]  ( .D(n287), .CLK(clk), .Q(\ram[0][226] ) );
  DFFX1_HVT \ram_reg[0][225]  ( .D(n286), .CLK(clk), .Q(\ram[0][225] ) );
  DFFX1_HVT \ram_reg[0][224]  ( .D(n285), .CLK(clk), .Q(\ram[0][224] ) );
  DFFX1_HVT \ram_reg[0][223]  ( .D(n284), .CLK(clk), .Q(\ram[0][223] ) );
  DFFX1_HVT \ram_reg[0][222]  ( .D(n283), .CLK(clk), .Q(\ram[0][222] ) );
  DFFX1_HVT \ram_reg[0][221]  ( .D(n282), .CLK(clk), .Q(\ram[0][221] ) );
  DFFX1_HVT \ram_reg[0][220]  ( .D(n281), .CLK(clk), .Q(\ram[0][220] ) );
  DFFX1_HVT \ram_reg[0][219]  ( .D(n280), .CLK(clk), .Q(\ram[0][219] ) );
  DFFX1_HVT \ram_reg[0][218]  ( .D(n279), .CLK(clk), .Q(\ram[0][218] ) );
  DFFX1_HVT \ram_reg[0][217]  ( .D(n278), .CLK(clk), .Q(\ram[0][217] ) );
  DFFX1_HVT \ram_reg[0][216]  ( .D(n277), .CLK(clk), .Q(\ram[0][216] ) );
  DFFX1_HVT \ram_reg[0][215]  ( .D(n276), .CLK(clk), .Q(\ram[0][215] ) );
  DFFX1_HVT \ram_reg[0][214]  ( .D(n275), .CLK(clk), .Q(\ram[0][214] ) );
  DFFX1_HVT \ram_reg[0][213]  ( .D(n274), .CLK(clk), .Q(\ram[0][213] ) );
  DFFX1_HVT \ram_reg[0][212]  ( .D(n273), .CLK(clk), .Q(\ram[0][212] ) );
  DFFX1_HVT \ram_reg[0][211]  ( .D(n272), .CLK(clk), .Q(\ram[0][211] ) );
  DFFX1_HVT \ram_reg[0][210]  ( .D(n271), .CLK(clk), .Q(\ram[0][210] ) );
  DFFX1_HVT \ram_reg[0][209]  ( .D(n270), .CLK(clk), .Q(\ram[0][209] ) );
  DFFX1_HVT \ram_reg[0][208]  ( .D(n269), .CLK(clk), .Q(\ram[0][208] ) );
  DFFX1_HVT \ram_reg[0][207]  ( .D(n268), .CLK(clk), .Q(\ram[0][207] ) );
  DFFX1_HVT \ram_reg[0][206]  ( .D(n267), .CLK(clk), .Q(\ram[0][206] ) );
  DFFX1_HVT \ram_reg[0][205]  ( .D(n266), .CLK(clk), .Q(\ram[0][205] ) );
  DFFX1_HVT \ram_reg[0][204]  ( .D(n265), .CLK(clk), .Q(\ram[0][204] ) );
  DFFX1_HVT \ram_reg[0][203]  ( .D(n264), .CLK(clk), .Q(\ram[0][203] ) );
  DFFX1_HVT \ram_reg[0][202]  ( .D(n263), .CLK(clk), .Q(\ram[0][202] ) );
  DFFX1_HVT \ram_reg[0][201]  ( .D(n262), .CLK(clk), .Q(\ram[0][201] ) );
  DFFX1_HVT \ram_reg[0][200]  ( .D(n261), .CLK(clk), .Q(\ram[0][200] ) );
  DFFX1_HVT \ram_reg[0][199]  ( .D(n260), .CLK(clk), .Q(\ram[0][199] ) );
  DFFX1_HVT \ram_reg[0][198]  ( .D(n259), .CLK(clk), .Q(\ram[0][198] ) );
  DFFX1_HVT \ram_reg[0][197]  ( .D(n258), .CLK(clk), .Q(\ram[0][197] ) );
  DFFX1_HVT \ram_reg[0][196]  ( .D(n257), .CLK(clk), .Q(\ram[0][196] ) );
  DFFX1_HVT \ram_reg[0][195]  ( .D(n256), .CLK(clk), .Q(\ram[0][195] ) );
  DFFX1_HVT \ram_reg[0][194]  ( .D(n255), .CLK(clk), .Q(\ram[0][194] ) );
  DFFX1_HVT \ram_reg[0][193]  ( .D(n254), .CLK(clk), .Q(\ram[0][193] ) );
  DFFX1_HVT \ram_reg[0][192]  ( .D(n253), .CLK(clk), .Q(\ram[0][192] ) );
  DFFX1_HVT \ram_reg[0][191]  ( .D(n252), .CLK(clk), .Q(\ram[0][191] ) );
  DFFX1_HVT \ram_reg[0][190]  ( .D(n251), .CLK(clk), .Q(\ram[0][190] ) );
  DFFX1_HVT \ram_reg[0][189]  ( .D(n250), .CLK(clk), .Q(\ram[0][189] ) );
  DFFX1_HVT \ram_reg[0][188]  ( .D(n249), .CLK(clk), .Q(\ram[0][188] ) );
  DFFX1_HVT \ram_reg[0][187]  ( .D(n248), .CLK(clk), .Q(\ram[0][187] ) );
  DFFX1_HVT \ram_reg[0][186]  ( .D(n247), .CLK(clk), .Q(\ram[0][186] ) );
  DFFX1_HVT \ram_reg[0][185]  ( .D(n246), .CLK(clk), .Q(\ram[0][185] ) );
  DFFX1_HVT \ram_reg[0][184]  ( .D(n245), .CLK(clk), .Q(\ram[0][184] ) );
  DFFX1_HVT \ram_reg[0][183]  ( .D(n244), .CLK(clk), .Q(\ram[0][183] ) );
  DFFX1_HVT \ram_reg[0][182]  ( .D(n243), .CLK(clk), .Q(\ram[0][182] ) );
  DFFX1_HVT \ram_reg[0][181]  ( .D(n242), .CLK(clk), .Q(\ram[0][181] ) );
  DFFX1_HVT \ram_reg[0][180]  ( .D(n241), .CLK(clk), .Q(\ram[0][180] ) );
  DFFX1_HVT \ram_reg[0][179]  ( .D(n240), .CLK(clk), .Q(\ram[0][179] ) );
  DFFX1_HVT \ram_reg[0][178]  ( .D(n239), .CLK(clk), .Q(\ram[0][178] ) );
  DFFX1_HVT \ram_reg[0][177]  ( .D(n238), .CLK(clk), .Q(\ram[0][177] ) );
  DFFX1_HVT \ram_reg[0][176]  ( .D(n237), .CLK(clk), .Q(\ram[0][176] ) );
  DFFX1_HVT \ram_reg[0][175]  ( .D(n236), .CLK(clk), .Q(\ram[0][175] ) );
  DFFX1_HVT \ram_reg[0][174]  ( .D(n235), .CLK(clk), .Q(\ram[0][174] ) );
  DFFX1_HVT \ram_reg[0][173]  ( .D(n234), .CLK(clk), .Q(\ram[0][173] ) );
  DFFX1_HVT \ram_reg[0][172]  ( .D(n233), .CLK(clk), .Q(\ram[0][172] ) );
  DFFX1_HVT \ram_reg[0][171]  ( .D(n232), .CLK(clk), .Q(\ram[0][171] ) );
  DFFX1_HVT \ram_reg[0][170]  ( .D(n231), .CLK(clk), .Q(\ram[0][170] ) );
  DFFX1_HVT \ram_reg[0][169]  ( .D(n230), .CLK(clk), .Q(\ram[0][169] ) );
  DFFX1_HVT \ram_reg[0][168]  ( .D(n229), .CLK(clk), .Q(\ram[0][168] ) );
  DFFX1_HVT \ram_reg[0][167]  ( .D(n228), .CLK(clk), .Q(\ram[0][167] ) );
  DFFX1_HVT \ram_reg[0][166]  ( .D(n227), .CLK(clk), .Q(\ram[0][166] ) );
  DFFX1_HVT \ram_reg[0][165]  ( .D(n226), .CLK(clk), .Q(\ram[0][165] ) );
  DFFX1_HVT \ram_reg[0][164]  ( .D(n225), .CLK(clk), .Q(\ram[0][164] ) );
  DFFX1_HVT \ram_reg[0][163]  ( .D(n224), .CLK(clk), .Q(\ram[0][163] ) );
  DFFX1_HVT \ram_reg[0][162]  ( .D(n223), .CLK(clk), .Q(\ram[0][162] ) );
  DFFX1_HVT \ram_reg[0][161]  ( .D(n222), .CLK(clk), .Q(\ram[0][161] ) );
  DFFX1_HVT \ram_reg[0][160]  ( .D(n221), .CLK(clk), .Q(\ram[0][160] ) );
  DFFX1_HVT \ram_reg[0][159]  ( .D(n220), .CLK(clk), .Q(\ram[0][159] ) );
  DFFX1_HVT \ram_reg[0][158]  ( .D(n219), .CLK(clk), .Q(\ram[0][158] ) );
  DFFX1_HVT \ram_reg[0][157]  ( .D(n218), .CLK(clk), .Q(\ram[0][157] ) );
  DFFX1_HVT \ram_reg[0][156]  ( .D(n217), .CLK(clk), .Q(\ram[0][156] ) );
  DFFX1_HVT \ram_reg[0][155]  ( .D(n216), .CLK(clk), .Q(\ram[0][155] ) );
  DFFX1_HVT \ram_reg[0][154]  ( .D(n215), .CLK(clk), .Q(\ram[0][154] ) );
  DFFX1_HVT \ram_reg[0][153]  ( .D(n214), .CLK(clk), .Q(\ram[0][153] ) );
  DFFX1_HVT \ram_reg[0][152]  ( .D(n213), .CLK(clk), .Q(\ram[0][152] ) );
  DFFX1_HVT \ram_reg[0][151]  ( .D(n212), .CLK(clk), .Q(\ram[0][151] ) );
  DFFX1_HVT \ram_reg[0][150]  ( .D(n211), .CLK(clk), .Q(\ram[0][150] ) );
  DFFX1_HVT \ram_reg[0][149]  ( .D(n210), .CLK(clk), .Q(\ram[0][149] ) );
  DFFX1_HVT \ram_reg[0][148]  ( .D(n209), .CLK(clk), .Q(\ram[0][148] ) );
  DFFX1_HVT \ram_reg[0][147]  ( .D(n208), .CLK(clk), .Q(\ram[0][147] ) );
  DFFX1_HVT \ram_reg[0][146]  ( .D(n207), .CLK(clk), .Q(\ram[0][146] ) );
  DFFX1_HVT \ram_reg[0][145]  ( .D(n206), .CLK(clk), .Q(\ram[0][145] ) );
  DFFX1_HVT \ram_reg[0][144]  ( .D(n205), .CLK(clk), .Q(\ram[0][144] ) );
  DFFX1_HVT \ram_reg[0][143]  ( .D(n204), .CLK(clk), .Q(\ram[0][143] ) );
  DFFX1_HVT \ram_reg[0][142]  ( .D(n203), .CLK(clk), .Q(\ram[0][142] ) );
  DFFX1_HVT \ram_reg[0][141]  ( .D(n202), .CLK(clk), .Q(\ram[0][141] ) );
  DFFX1_HVT \ram_reg[0][140]  ( .D(n201), .CLK(clk), .Q(\ram[0][140] ) );
  DFFX1_HVT \ram_reg[0][139]  ( .D(n200), .CLK(clk), .Q(\ram[0][139] ) );
  DFFX1_HVT \ram_reg[0][138]  ( .D(n199), .CLK(clk), .Q(\ram[0][138] ) );
  DFFX1_HVT \ram_reg[0][137]  ( .D(n198), .CLK(clk), .Q(\ram[0][137] ) );
  DFFX1_HVT \ram_reg[0][136]  ( .D(n197), .CLK(clk), .Q(\ram[0][136] ) );
  DFFX1_HVT \ram_reg[0][135]  ( .D(n196), .CLK(clk), .Q(\ram[0][135] ) );
  DFFX1_HVT \ram_reg[0][134]  ( .D(n195), .CLK(clk), .Q(\ram[0][134] ) );
  DFFX1_HVT \ram_reg[0][133]  ( .D(n194), .CLK(clk), .Q(\ram[0][133] ) );
  DFFX1_HVT \ram_reg[0][132]  ( .D(n193), .CLK(clk), .Q(\ram[0][132] ) );
  DFFX1_HVT \ram_reg[0][131]  ( .D(n192), .CLK(clk), .Q(\ram[0][131] ) );
  DFFX1_HVT \ram_reg[0][130]  ( .D(n191), .CLK(clk), .Q(\ram[0][130] ) );
  DFFX1_HVT \ram_reg[0][129]  ( .D(n190), .CLK(clk), .Q(\ram[0][129] ) );
  DFFX1_HVT \ram_reg[0][128]  ( .D(n189), .CLK(clk), .Q(\ram[0][128] ) );
  DFFX1_HVT \ram_reg[0][127]  ( .D(n188), .CLK(clk), .Q(\ram[0][127] ) );
  DFFX1_HVT \ram_reg[0][126]  ( .D(n187), .CLK(clk), .Q(\ram[0][126] ) );
  DFFX1_HVT \ram_reg[0][125]  ( .D(n186), .CLK(clk), .Q(\ram[0][125] ) );
  DFFX1_HVT \ram_reg[0][124]  ( .D(n185), .CLK(clk), .Q(\ram[0][124] ) );
  DFFX1_HVT \ram_reg[0][123]  ( .D(n184), .CLK(clk), .Q(\ram[0][123] ) );
  DFFX1_HVT \ram_reg[0][122]  ( .D(n183), .CLK(clk), .Q(\ram[0][122] ) );
  DFFX1_HVT \ram_reg[0][121]  ( .D(n182), .CLK(clk), .Q(\ram[0][121] ) );
  DFFX1_HVT \ram_reg[0][120]  ( .D(n181), .CLK(clk), .Q(\ram[0][120] ) );
  DFFX1_HVT \ram_reg[0][119]  ( .D(n180), .CLK(clk), .Q(\ram[0][119] ) );
  DFFX1_HVT \ram_reg[0][118]  ( .D(n179), .CLK(clk), .Q(\ram[0][118] ) );
  DFFX1_HVT \ram_reg[0][117]  ( .D(n178), .CLK(clk), .Q(\ram[0][117] ) );
  DFFX1_HVT \ram_reg[0][116]  ( .D(n177), .CLK(clk), .Q(\ram[0][116] ) );
  DFFX1_HVT \ram_reg[0][115]  ( .D(n176), .CLK(clk), .Q(\ram[0][115] ) );
  DFFX1_HVT \ram_reg[0][114]  ( .D(n175), .CLK(clk), .Q(\ram[0][114] ) );
  DFFX1_HVT \ram_reg[0][113]  ( .D(n174), .CLK(clk), .Q(\ram[0][113] ) );
  DFFX1_HVT \ram_reg[0][112]  ( .D(n173), .CLK(clk), .Q(\ram[0][112] ) );
  DFFX1_HVT \ram_reg[0][111]  ( .D(n172), .CLK(clk), .Q(\ram[0][111] ) );
  DFFX1_HVT \ram_reg[0][110]  ( .D(n171), .CLK(clk), .Q(\ram[0][110] ) );
  DFFX1_HVT \ram_reg[0][109]  ( .D(n170), .CLK(clk), .Q(\ram[0][109] ) );
  DFFX1_HVT \ram_reg[0][108]  ( .D(n169), .CLK(clk), .Q(\ram[0][108] ) );
  DFFX1_HVT \ram_reg[0][107]  ( .D(n168), .CLK(clk), .Q(\ram[0][107] ) );
  DFFX1_HVT \ram_reg[0][106]  ( .D(n167), .CLK(clk), .Q(\ram[0][106] ) );
  DFFX1_HVT \ram_reg[0][105]  ( .D(n166), .CLK(clk), .Q(\ram[0][105] ) );
  DFFX1_HVT \ram_reg[0][104]  ( .D(n165), .CLK(clk), .Q(\ram[0][104] ) );
  DFFX1_HVT \ram_reg[0][103]  ( .D(n164), .CLK(clk), .Q(\ram[0][103] ) );
  DFFX1_HVT \ram_reg[0][102]  ( .D(n163), .CLK(clk), .Q(\ram[0][102] ) );
  DFFX1_HVT \ram_reg[0][101]  ( .D(n162), .CLK(clk), .Q(\ram[0][101] ) );
  DFFX1_HVT \ram_reg[0][100]  ( .D(n161), .CLK(clk), .Q(\ram[0][100] ) );
  DFFX1_HVT \ram_reg[0][99]  ( .D(n160), .CLK(clk), .Q(\ram[0][99] ) );
  DFFX1_HVT \ram_reg[0][98]  ( .D(n159), .CLK(clk), .Q(\ram[0][98] ) );
  DFFX1_HVT \ram_reg[0][97]  ( .D(n158), .CLK(clk), .Q(\ram[0][97] ) );
  DFFX1_HVT \ram_reg[0][96]  ( .D(n157), .CLK(clk), .Q(\ram[0][96] ) );
  DFFX1_HVT \ram_reg[0][95]  ( .D(n156), .CLK(clk), .Q(\ram[0][95] ) );
  DFFX1_HVT \ram_reg[0][94]  ( .D(n155), .CLK(clk), .Q(\ram[0][94] ) );
  DFFX1_HVT \ram_reg[0][93]  ( .D(n154), .CLK(clk), .Q(\ram[0][93] ) );
  DFFX1_HVT \ram_reg[0][92]  ( .D(n153), .CLK(clk), .Q(\ram[0][92] ) );
  DFFX1_HVT \ram_reg[0][91]  ( .D(n152), .CLK(clk), .Q(\ram[0][91] ) );
  DFFX1_HVT \ram_reg[0][90]  ( .D(n151), .CLK(clk), .Q(\ram[0][90] ) );
  DFFX1_HVT \ram_reg[0][89]  ( .D(n150), .CLK(clk), .Q(\ram[0][89] ) );
  DFFX1_HVT \ram_reg[0][88]  ( .D(n149), .CLK(clk), .Q(\ram[0][88] ) );
  DFFX1_HVT \ram_reg[0][87]  ( .D(n148), .CLK(clk), .Q(\ram[0][87] ) );
  DFFX1_HVT \ram_reg[0][86]  ( .D(n147), .CLK(clk), .Q(\ram[0][86] ) );
  DFFX1_HVT \ram_reg[0][85]  ( .D(n146), .CLK(clk), .Q(\ram[0][85] ) );
  DFFX1_HVT \ram_reg[0][84]  ( .D(n145), .CLK(clk), .Q(\ram[0][84] ) );
  DFFX1_HVT \ram_reg[0][83]  ( .D(n144), .CLK(clk), .Q(\ram[0][83] ) );
  DFFX1_HVT \ram_reg[0][82]  ( .D(n143), .CLK(clk), .Q(\ram[0][82] ) );
  DFFX1_HVT \ram_reg[0][81]  ( .D(n142), .CLK(clk), .Q(\ram[0][81] ) );
  DFFX1_HVT \ram_reg[0][80]  ( .D(n141), .CLK(clk), .Q(\ram[0][80] ) );
  DFFX1_HVT \ram_reg[0][79]  ( .D(n140), .CLK(clk), .Q(\ram[0][79] ) );
  DFFX1_HVT \ram_reg[0][78]  ( .D(n139), .CLK(clk), .Q(\ram[0][78] ) );
  DFFX1_HVT \ram_reg[0][77]  ( .D(n138), .CLK(clk), .Q(\ram[0][77] ) );
  DFFX1_HVT \ram_reg[0][76]  ( .D(n137), .CLK(clk), .Q(\ram[0][76] ) );
  DFFX1_HVT \ram_reg[0][75]  ( .D(n136), .CLK(clk), .Q(\ram[0][75] ) );
  DFFX1_HVT \ram_reg[0][74]  ( .D(n135), .CLK(clk), .Q(\ram[0][74] ) );
  DFFX1_HVT \ram_reg[0][73]  ( .D(n134), .CLK(clk), .Q(\ram[0][73] ) );
  DFFX1_HVT \ram_reg[0][72]  ( .D(n133), .CLK(clk), .Q(\ram[0][72] ) );
  DFFX1_HVT \ram_reg[0][71]  ( .D(n132), .CLK(clk), .Q(\ram[0][71] ) );
  DFFX1_HVT \ram_reg[0][70]  ( .D(n131), .CLK(clk), .Q(\ram[0][70] ) );
  DFFX1_HVT \ram_reg[0][69]  ( .D(n130), .CLK(clk), .Q(\ram[0][69] ) );
  DFFX1_HVT \ram_reg[0][68]  ( .D(n129), .CLK(clk), .Q(\ram[0][68] ) );
  DFFX1_HVT \ram_reg[0][67]  ( .D(n128), .CLK(clk), .Q(\ram[0][67] ) );
  DFFX1_HVT \ram_reg[0][66]  ( .D(n127), .CLK(clk), .Q(\ram[0][66] ) );
  DFFX1_HVT \ram_reg[0][65]  ( .D(n126), .CLK(clk), .Q(\ram[0][65] ) );
  DFFX1_HVT \ram_reg[0][64]  ( .D(n125), .CLK(clk), .Q(\ram[0][64] ) );
  DFFX1_HVT \ram_reg[0][63]  ( .D(n124), .CLK(clk), .Q(\ram[0][63] ) );
  DFFX1_HVT \ram_reg[0][62]  ( .D(n123), .CLK(clk), .Q(\ram[0][62] ) );
  DFFX1_HVT \ram_reg[0][61]  ( .D(n122), .CLK(clk), .Q(\ram[0][61] ) );
  DFFX1_HVT \ram_reg[0][60]  ( .D(n121), .CLK(clk), .Q(\ram[0][60] ) );
  DFFX1_HVT \ram_reg[0][59]  ( .D(n120), .CLK(clk), .Q(\ram[0][59] ) );
  DFFX1_HVT \ram_reg[0][58]  ( .D(n119), .CLK(clk), .Q(\ram[0][58] ) );
  DFFX1_HVT \ram_reg[0][57]  ( .D(n118), .CLK(clk), .Q(\ram[0][57] ) );
  DFFX1_HVT \ram_reg[0][56]  ( .D(n117), .CLK(clk), .Q(\ram[0][56] ) );
  DFFX1_HVT \ram_reg[0][55]  ( .D(n116), .CLK(clk), .Q(\ram[0][55] ) );
  DFFX1_HVT \ram_reg[0][54]  ( .D(n115), .CLK(clk), .Q(\ram[0][54] ) );
  DFFX1_HVT \ram_reg[0][53]  ( .D(n114), .CLK(clk), .Q(\ram[0][53] ) );
  DFFX1_HVT \ram_reg[0][52]  ( .D(n113), .CLK(clk), .Q(\ram[0][52] ) );
  DFFX1_HVT \ram_reg[0][51]  ( .D(n112), .CLK(clk), .Q(\ram[0][51] ) );
  DFFX1_HVT \ram_reg[0][50]  ( .D(n111), .CLK(clk), .Q(\ram[0][50] ) );
  DFFX1_HVT \ram_reg[0][49]  ( .D(n110), .CLK(clk), .Q(\ram[0][49] ) );
  DFFX1_HVT \ram_reg[0][48]  ( .D(n109), .CLK(clk), .Q(\ram[0][48] ) );
  DFFX1_HVT \ram_reg[0][47]  ( .D(n108), .CLK(clk), .Q(\ram[0][47] ) );
  DFFX1_HVT \ram_reg[0][46]  ( .D(n107), .CLK(clk), .Q(\ram[0][46] ) );
  DFFX1_HVT \ram_reg[0][45]  ( .D(n106), .CLK(clk), .Q(\ram[0][45] ) );
  DFFX1_HVT \ram_reg[0][44]  ( .D(n105), .CLK(clk), .Q(\ram[0][44] ) );
  DFFX1_HVT \ram_reg[0][43]  ( .D(n104), .CLK(clk), .Q(\ram[0][43] ) );
  DFFX1_HVT \ram_reg[0][42]  ( .D(n103), .CLK(clk), .Q(\ram[0][42] ) );
  DFFX1_HVT \ram_reg[0][41]  ( .D(n102), .CLK(clk), .Q(\ram[0][41] ) );
  DFFX1_HVT \ram_reg[0][40]  ( .D(n101), .CLK(clk), .Q(\ram[0][40] ) );
  DFFX1_HVT \ram_reg[0][39]  ( .D(n100), .CLK(clk), .Q(\ram[0][39] ) );
  DFFX1_HVT \ram_reg[0][38]  ( .D(n99), .CLK(clk), .Q(\ram[0][38] ) );
  DFFX1_HVT \ram_reg[0][37]  ( .D(n98), .CLK(clk), .Q(\ram[0][37] ) );
  DFFX1_HVT \ram_reg[0][36]  ( .D(n97), .CLK(clk), .Q(\ram[0][36] ) );
  DFFX1_HVT \ram_reg[0][35]  ( .D(n96), .CLK(clk), .Q(\ram[0][35] ) );
  DFFX1_HVT \ram_reg[0][34]  ( .D(n95), .CLK(clk), .Q(\ram[0][34] ) );
  DFFX1_HVT \ram_reg[0][33]  ( .D(n94), .CLK(clk), .Q(\ram[0][33] ) );
  DFFX1_HVT \ram_reg[0][32]  ( .D(n93), .CLK(clk), .Q(\ram[0][32] ) );
  DFFX1_HVT \ram_reg[0][31]  ( .D(n92), .CLK(clk), .Q(\ram[0][31] ) );
  DFFX1_HVT \ram_reg[0][30]  ( .D(n91), .CLK(clk), .Q(\ram[0][30] ) );
  DFFX1_HVT \ram_reg[0][29]  ( .D(n90), .CLK(clk), .Q(\ram[0][29] ) );
  DFFX1_HVT \ram_reg[0][28]  ( .D(n89), .CLK(clk), .Q(\ram[0][28] ) );
  DFFX1_HVT \ram_reg[0][27]  ( .D(n88), .CLK(clk), .Q(\ram[0][27] ) );
  DFFX1_HVT \ram_reg[0][26]  ( .D(n87), .CLK(clk), .Q(\ram[0][26] ) );
  DFFX1_HVT \ram_reg[0][25]  ( .D(n86), .CLK(clk), .Q(\ram[0][25] ) );
  DFFX1_HVT \ram_reg[0][24]  ( .D(n85), .CLK(clk), .Q(\ram[0][24] ) );
  DFFX1_HVT \ram_reg[0][23]  ( .D(n84), .CLK(clk), .Q(\ram[0][23] ) );
  DFFX1_HVT \ram_reg[0][22]  ( .D(n83), .CLK(clk), .Q(\ram[0][22] ) );
  DFFX1_HVT \ram_reg[0][21]  ( .D(n82), .CLK(clk), .Q(\ram[0][21] ) );
  DFFX1_HVT \ram_reg[0][20]  ( .D(n81), .CLK(clk), .Q(\ram[0][20] ) );
  DFFX1_HVT \ram_reg[0][19]  ( .D(n80), .CLK(clk), .Q(\ram[0][19] ) );
  DFFX1_HVT \ram_reg[0][18]  ( .D(n79), .CLK(clk), .Q(\ram[0][18] ) );
  DFFX1_HVT \ram_reg[0][17]  ( .D(n78), .CLK(clk), .Q(\ram[0][17] ) );
  DFFX1_HVT \ram_reg[0][16]  ( .D(n77), .CLK(clk), .Q(\ram[0][16] ) );
  DFFX1_HVT \ram_reg[0][15]  ( .D(n76), .CLK(clk), .Q(\ram[0][15] ) );
  DFFX1_HVT \ram_reg[0][14]  ( .D(n75), .CLK(clk), .Q(\ram[0][14] ) );
  DFFX1_HVT \ram_reg[0][13]  ( .D(n74), .CLK(clk), .Q(\ram[0][13] ) );
  DFFX1_HVT \ram_reg[0][12]  ( .D(n73), .CLK(clk), .Q(\ram[0][12] ) );
  DFFX1_HVT \ram_reg[0][11]  ( .D(n72), .CLK(clk), .Q(\ram[0][11] ) );
  DFFX1_HVT \ram_reg[0][10]  ( .D(n71), .CLK(clk), .Q(\ram[0][10] ) );
  DFFX1_HVT \ram_reg[0][9]  ( .D(n70), .CLK(clk), .Q(\ram[0][9] ) );
  DFFX1_HVT \ram_reg[0][8]  ( .D(n69), .CLK(clk), .Q(\ram[0][8] ) );
  DFFX1_HVT \ram_reg[0][7]  ( .D(n68), .CLK(clk), .Q(\ram[0][7] ) );
  DFFX1_HVT \ram_reg[0][6]  ( .D(n67), .CLK(clk), .Q(\ram[0][6] ) );
  DFFX1_HVT \ram_reg[0][5]  ( .D(n66), .CLK(clk), .Q(\ram[0][5] ) );
  DFFX1_HVT \ram_reg[0][4]  ( .D(n65), .CLK(clk), .Q(\ram[0][4] ) );
  DFFX1_HVT \ram_reg[0][3]  ( .D(n64), .CLK(clk), .Q(\ram[0][3] ) );
  DFFX1_HVT \ram_reg[0][2]  ( .D(n63), .CLK(clk), .Q(\ram[0][2] ) );
  DFFX1_HVT \ram_reg[0][1]  ( .D(n62), .CLK(clk), .Q(\ram[0][1] ) );
  DFFX1_HVT \ram_reg[0][0]  ( .D(n61), .CLK(clk), .Q(\ram[0][0] ) );
  INVX1_HVT U3 ( .A(n4277), .Y(n4276) );
  INVX1_HVT U4 ( .A(n4285), .Y(n4191) );
  INVX1_HVT U5 ( .A(n4286), .Y(n4192) );
  INVX1_HVT U6 ( .A(n4332), .Y(n4310) );
  INVX1_HVT U7 ( .A(n4333), .Y(n4311) );
  INVX1_HVT U8 ( .A(n4331), .Y(n4312) );
  INVX1_HVT U9 ( .A(n4332), .Y(n4313) );
  INVX1_HVT U10 ( .A(n4332), .Y(n4321) );
  INVX1_HVT U11 ( .A(n4332), .Y(n4322) );
  INVX1_HVT U12 ( .A(n4332), .Y(n4323) );
  INVX1_HVT U13 ( .A(n4332), .Y(n4324) );
  INVX1_HVT U14 ( .A(n4332), .Y(n4325) );
  INVX1_HVT U15 ( .A(n4333), .Y(n4314) );
  INVX1_HVT U16 ( .A(n4333), .Y(n4315) );
  INVX1_HVT U17 ( .A(n4333), .Y(n4316) );
  INVX1_HVT U18 ( .A(n4333), .Y(n4317) );
  INVX1_HVT U19 ( .A(n4333), .Y(n4318) );
  INVX1_HVT U20 ( .A(n4333), .Y(n4319) );
  INVX1_HVT U21 ( .A(n4332), .Y(n4320) );
  INVX1_HVT U22 ( .A(n4331), .Y(n4326) );
  INVX1_HVT U23 ( .A(n4331), .Y(n4327) );
  INVX1_HVT U24 ( .A(n4331), .Y(n4328) );
  INVX1_HVT U25 ( .A(n4331), .Y(n4329) );
  INVX1_HVT U26 ( .A(n4331), .Y(n4330) );
  INVX1_HVT U27 ( .A(n4183), .Y(n1) );
  INVX1_HVT U28 ( .A(n4183), .Y(n2) );
  INVX1_HVT U29 ( .A(n4183), .Y(n4) );
  INVX1_HVT U30 ( .A(n4183), .Y(n5) );
  INVX1_HVT U31 ( .A(n4184), .Y(n12) );
  INVX1_HVT U32 ( .A(n4184), .Y(n13) );
  INVX1_HVT U33 ( .A(n4184), .Y(n14) );
  INVX1_HVT U34 ( .A(n4186), .Y(n15) );
  INVX1_HVT U35 ( .A(n4184), .Y(n16) );
  INVX1_HVT U36 ( .A(n4184), .Y(n17) );
  INVX1_HVT U37 ( .A(n4184), .Y(n18) );
  INVX1_HVT U38 ( .A(n4185), .Y(n19) );
  INVX1_HVT U39 ( .A(n4185), .Y(n20) );
  INVX1_HVT U40 ( .A(n4185), .Y(n21) );
  INVX1_HVT U41 ( .A(n4184), .Y(n3) );
  INVX1_HVT U42 ( .A(n4184), .Y(n6) );
  INVX1_HVT U43 ( .A(n4184), .Y(n7) );
  INVX1_HVT U44 ( .A(n4184), .Y(n8) );
  INVX1_HVT U45 ( .A(n4184), .Y(n9) );
  INVX1_HVT U46 ( .A(n4184), .Y(n10) );
  INVX1_HVT U47 ( .A(n4184), .Y(n11) );
  INVX1_HVT U48 ( .A(n4186), .Y(n34) );
  INVX1_HVT U49 ( .A(n4186), .Y(n35) );
  INVX1_HVT U50 ( .A(n4186), .Y(n36) );
  INVX1_HVT U51 ( .A(n4186), .Y(n37) );
  INVX1_HVT U52 ( .A(n4186), .Y(n38) );
  INVX1_HVT U53 ( .A(n4186), .Y(n39) );
  INVX1_HVT U54 ( .A(n4186), .Y(n40) );
  INVX1_HVT U55 ( .A(n4186), .Y(n41) );
  INVX1_HVT U56 ( .A(n4186), .Y(n42) );
  INVX1_HVT U57 ( .A(n4185), .Y(n22) );
  INVX1_HVT U58 ( .A(n4185), .Y(n23) );
  INVX1_HVT U59 ( .A(n4185), .Y(n24) );
  INVX1_HVT U60 ( .A(n4185), .Y(n25) );
  INVX1_HVT U61 ( .A(n4185), .Y(n26) );
  INVX1_HVT U62 ( .A(n4185), .Y(n27) );
  INVX1_HVT U63 ( .A(n4185), .Y(n28) );
  INVX1_HVT U64 ( .A(n4185), .Y(n29) );
  INVX1_HVT U65 ( .A(n4185), .Y(n30) );
  INVX1_HVT U66 ( .A(n4185), .Y(n31) );
  INVX1_HVT U67 ( .A(n4186), .Y(n33) );
  INVX1_HVT U68 ( .A(n4186), .Y(n32) );
  INVX1_HVT U69 ( .A(n4187), .Y(n55) );
  INVX1_HVT U70 ( .A(n4187), .Y(n56) );
  INVX1_HVT U71 ( .A(n4188), .Y(n57) );
  INVX1_HVT U72 ( .A(n4188), .Y(n58) );
  INVX1_HVT U73 ( .A(n4188), .Y(n59) );
  INVX1_HVT U74 ( .A(n4188), .Y(n60) );
  INVX1_HVT U75 ( .A(n4188), .Y(n4157) );
  INVX1_HVT U76 ( .A(n4188), .Y(n4158) );
  INVX1_HVT U77 ( .A(n4188), .Y(n4159) );
  INVX1_HVT U78 ( .A(n4188), .Y(n4160) );
  INVX1_HVT U79 ( .A(n4186), .Y(n43) );
  INVX1_HVT U80 ( .A(n4187), .Y(n44) );
  INVX1_HVT U81 ( .A(n4187), .Y(n45) );
  INVX1_HVT U82 ( .A(n4187), .Y(n46) );
  INVX1_HVT U83 ( .A(n4187), .Y(n47) );
  INVX1_HVT U84 ( .A(n4187), .Y(n48) );
  INVX1_HVT U85 ( .A(n4187), .Y(n49) );
  INVX1_HVT U86 ( .A(n4187), .Y(n50) );
  INVX1_HVT U87 ( .A(n4187), .Y(n51) );
  INVX1_HVT U88 ( .A(n4187), .Y(n52) );
  INVX1_HVT U89 ( .A(n4187), .Y(n53) );
  INVX1_HVT U90 ( .A(n4187), .Y(n54) );
  INVX1_HVT U91 ( .A(n4189), .Y(n4172) );
  INVX1_HVT U92 ( .A(n4189), .Y(n4173) );
  INVX1_HVT U93 ( .A(n4189), .Y(n4174) );
  INVX1_HVT U94 ( .A(n4189), .Y(n4175) );
  INVX1_HVT U95 ( .A(n4189), .Y(n4176) );
  INVX1_HVT U96 ( .A(n4189), .Y(n4177) );
  INVX1_HVT U97 ( .A(n4189), .Y(n4178) );
  INVX1_HVT U98 ( .A(n4188), .Y(n4161) );
  INVX1_HVT U99 ( .A(n4188), .Y(n4162) );
  INVX1_HVT U100 ( .A(n4188), .Y(n4163) );
  INVX1_HVT U101 ( .A(n4188), .Y(n4164) );
  INVX1_HVT U102 ( .A(n4188), .Y(n4165) );
  INVX1_HVT U103 ( .A(n4189), .Y(n4166) );
  INVX1_HVT U104 ( .A(n4189), .Y(n4167) );
  INVX1_HVT U105 ( .A(n4189), .Y(n4168) );
  INVX1_HVT U106 ( .A(n4189), .Y(n4169) );
  INVX1_HVT U107 ( .A(n4189), .Y(n4170) );
  INVX1_HVT U108 ( .A(n4189), .Y(n4171) );
  INVX1_HVT U109 ( .A(n4190), .Y(n4179) );
  INVX1_HVT U110 ( .A(n4190), .Y(n4180) );
  INVX1_HVT U111 ( .A(n4190), .Y(n4181) );
  INVX1_HVT U112 ( .A(n4309), .Y(n4298) );
  INVX1_HVT U113 ( .A(n4309), .Y(n4299) );
  INVX1_HVT U114 ( .A(n4309), .Y(n4300) );
  INVX1_HVT U115 ( .A(n4309), .Y(n4301) );
  INVX1_HVT U116 ( .A(n4309), .Y(n4302) );
  INVX1_HVT U117 ( .A(n4309), .Y(n4303) );
  INVX1_HVT U118 ( .A(n4309), .Y(n4304) );
  INVX1_HVT U119 ( .A(n4309), .Y(n4305) );
  INVX1_HVT U120 ( .A(n4309), .Y(n4306) );
  INVX1_HVT U121 ( .A(n4309), .Y(n4307) );
  INVX1_HVT U122 ( .A(n4308), .Y(n4287) );
  INVX1_HVT U123 ( .A(n4308), .Y(n4288) );
  INVX1_HVT U124 ( .A(n4308), .Y(n4289) );
  INVX1_HVT U125 ( .A(n4308), .Y(n4290) );
  INVX1_HVT U126 ( .A(n4308), .Y(n4291) );
  INVX1_HVT U127 ( .A(n4308), .Y(n4292) );
  INVX1_HVT U128 ( .A(n4308), .Y(n4293) );
  INVX1_HVT U129 ( .A(n4308), .Y(n4294) );
  INVX1_HVT U130 ( .A(n4308), .Y(n4295) );
  INVX1_HVT U131 ( .A(n4308), .Y(n4296) );
  INVX1_HVT U132 ( .A(n4308), .Y(n4297) );
  INVX1_HVT U133 ( .A(n4277), .Y(n4271) );
  INVX1_HVT U134 ( .A(n4277), .Y(n4272) );
  INVX1_HVT U135 ( .A(n4277), .Y(n4273) );
  INVX1_HVT U136 ( .A(n4277), .Y(n4274) );
  INVX1_HVT U137 ( .A(n4277), .Y(n4275) );
  INVX1_HVT U138 ( .A(n4280), .Y(n4247) );
  INVX1_HVT U139 ( .A(n4280), .Y(n4248) );
  INVX1_HVT U140 ( .A(n4280), .Y(n4249) );
  INVX1_HVT U141 ( .A(n4280), .Y(n4250) );
  INVX1_HVT U142 ( .A(n4280), .Y(n4251) );
  INVX1_HVT U143 ( .A(n4280), .Y(n4252) );
  INVX1_HVT U144 ( .A(n4279), .Y(n4253) );
  INVX1_HVT U145 ( .A(n4279), .Y(n4254) );
  INVX1_HVT U146 ( .A(n4280), .Y(n4266) );
  INVX1_HVT U147 ( .A(n4279), .Y(n4267) );
  INVX1_HVT U148 ( .A(n4278), .Y(n4268) );
  INVX1_HVT U149 ( .A(n4277), .Y(n4269) );
  INVX1_HVT U150 ( .A(n4285), .Y(n4270) );
  INVX1_HVT U151 ( .A(n4279), .Y(n4255) );
  INVX1_HVT U152 ( .A(n4279), .Y(n4256) );
  INVX1_HVT U153 ( .A(n4279), .Y(n4257) );
  INVX1_HVT U154 ( .A(n4279), .Y(n4258) );
  INVX1_HVT U155 ( .A(n4278), .Y(n4259) );
  INVX1_HVT U156 ( .A(n4278), .Y(n4260) );
  INVX1_HVT U157 ( .A(n4278), .Y(n4261) );
  INVX1_HVT U158 ( .A(n4278), .Y(n4262) );
  INVX1_HVT U159 ( .A(n4278), .Y(n4263) );
  INVX1_HVT U160 ( .A(n4278), .Y(n4264) );
  INVX1_HVT U161 ( .A(n4286), .Y(n4265) );
  INVX1_HVT U162 ( .A(n4183), .Y(n4182) );
  INVX1_HVT U163 ( .A(n4285), .Y(n4202) );
  INVX1_HVT U164 ( .A(n4286), .Y(n4203) );
  INVX1_HVT U165 ( .A(n4283), .Y(n4204) );
  INVX1_HVT U166 ( .A(n4285), .Y(n4205) );
  INVX1_HVT U167 ( .A(n4285), .Y(n4206) );
  INVX1_HVT U168 ( .A(n4285), .Y(n4207) );
  INVX1_HVT U169 ( .A(n4285), .Y(n4208) );
  INVX1_HVT U170 ( .A(n4285), .Y(n4209) );
  INVX1_HVT U171 ( .A(n4285), .Y(n4210) );
  INVX1_HVT U172 ( .A(n4284), .Y(n4211) );
  INVX1_HVT U173 ( .A(n4286), .Y(n4193) );
  INVX1_HVT U174 ( .A(n4286), .Y(n4194) );
  INVX1_HVT U175 ( .A(n4286), .Y(n4195) );
  INVX1_HVT U176 ( .A(n4286), .Y(n4196) );
  INVX1_HVT U177 ( .A(n4286), .Y(n4197) );
  INVX1_HVT U178 ( .A(n4286), .Y(n4198) );
  INVX1_HVT U179 ( .A(n4284), .Y(n4199) );
  INVX1_HVT U180 ( .A(n4282), .Y(n4200) );
  INVX1_HVT U181 ( .A(n4281), .Y(n4201) );
  INVX1_HVT U182 ( .A(n4277), .Y(n4224) );
  INVX1_HVT U183 ( .A(n4283), .Y(n4225) );
  INVX1_HVT U184 ( .A(n4284), .Y(n4226) );
  INVX1_HVT U185 ( .A(n4283), .Y(n4227) );
  INVX1_HVT U186 ( .A(n4282), .Y(n4228) );
  INVX1_HVT U187 ( .A(n4283), .Y(n4229) );
  INVX1_HVT U188 ( .A(n4283), .Y(n4230) );
  INVX1_HVT U189 ( .A(n4283), .Y(n4231) );
  INVX1_HVT U190 ( .A(n4283), .Y(n4232) );
  INVX1_HVT U191 ( .A(n4284), .Y(n4212) );
  INVX1_HVT U192 ( .A(n4284), .Y(n4213) );
  INVX1_HVT U193 ( .A(n4284), .Y(n4214) );
  INVX1_HVT U194 ( .A(n4284), .Y(n4215) );
  INVX1_HVT U195 ( .A(n4284), .Y(n4216) );
  INVX1_HVT U196 ( .A(n4284), .Y(n4217) );
  INVX1_HVT U197 ( .A(n4282), .Y(n4218) );
  INVX1_HVT U198 ( .A(n4281), .Y(n4219) );
  INVX1_HVT U199 ( .A(n4280), .Y(n4220) );
  INVX1_HVT U200 ( .A(n4279), .Y(n4221) );
  INVX1_HVT U201 ( .A(n4281), .Y(n4223) );
  INVX1_HVT U202 ( .A(n4278), .Y(n4222) );
  INVX1_HVT U203 ( .A(n4281), .Y(n4245) );
  INVX1_HVT U204 ( .A(n4281), .Y(n4246) );
  INVX1_HVT U205 ( .A(n4283), .Y(n4233) );
  INVX1_HVT U206 ( .A(n4283), .Y(n4234) );
  INVX1_HVT U207 ( .A(n4282), .Y(n4235) );
  INVX1_HVT U208 ( .A(n4282), .Y(n4236) );
  INVX1_HVT U209 ( .A(n4282), .Y(n4237) );
  INVX1_HVT U210 ( .A(n4282), .Y(n4238) );
  INVX1_HVT U211 ( .A(n4282), .Y(n4239) );
  INVX1_HVT U212 ( .A(n4282), .Y(n4240) );
  INVX1_HVT U213 ( .A(n4281), .Y(n4241) );
  INVX1_HVT U214 ( .A(n4281), .Y(n4242) );
  INVX1_HVT U215 ( .A(n4281), .Y(n4243) );
  INVX1_HVT U216 ( .A(n4281), .Y(n4244) );
  INVX1_HVT U217 ( .A(N28), .Y(n4309) );
  INVX1_HVT U218 ( .A(N28), .Y(n4308) );
  INVX1_HVT U219 ( .A(N29), .Y(n4332) );
  INVX1_HVT U220 ( .A(N29), .Y(n4333) );
  INVX1_HVT U221 ( .A(N29), .Y(n4331) );
  INVX1_HVT U222 ( .A(N26), .Y(n4184) );
  INVX1_HVT U223 ( .A(N26), .Y(n4185) );
  INVX1_HVT U224 ( .A(N26), .Y(n4186) );
  INVX1_HVT U225 ( .A(N26), .Y(n4187) );
  INVX1_HVT U226 ( .A(N26), .Y(n4188) );
  INVX1_HVT U227 ( .A(N26), .Y(n4189) );
  INVX1_HVT U228 ( .A(N26), .Y(n4183) );
  INVX1_HVT U229 ( .A(N26), .Y(n4190) );
  INVX1_HVT U230 ( .A(N27), .Y(n4277) );
  INVX1_HVT U231 ( .A(N27), .Y(n4280) );
  INVX1_HVT U232 ( .A(N27), .Y(n4279) );
  INVX1_HVT U233 ( .A(N27), .Y(n4278) );
  INVX1_HVT U234 ( .A(N27), .Y(n4285) );
  INVX1_HVT U235 ( .A(N27), .Y(n4286) );
  INVX1_HVT U236 ( .A(N27), .Y(n4283) );
  INVX1_HVT U237 ( .A(N27), .Y(n4284) );
  INVX1_HVT U238 ( .A(N27), .Y(n4282) );
  INVX1_HVT U239 ( .A(N27), .Y(n4281) );
  MUX41X1_HVT U240 ( .A1(\ram[12][0] ), .A3(\ram[14][0] ), .A2(\ram[13][0] ), 
        .A4(\ram[15][0] ), .S0(n4191), .S1(n1), .Y(n4334) );
  MUX41X1_HVT U241 ( .A1(\ram[8][0] ), .A3(\ram[10][0] ), .A2(\ram[9][0] ), 
        .A4(\ram[11][0] ), .S0(n4255), .S1(n4161), .Y(n4335) );
  MUX41X1_HVT U242 ( .A1(\ram[4][0] ), .A3(\ram[6][0] ), .A2(\ram[5][0] ), 
        .A4(\ram[7][0] ), .S0(n4249), .S1(n59), .Y(n4336) );
  MUX41X1_HVT U243 ( .A1(\ram[0][0] ), .A3(\ram[2][0] ), .A2(\ram[1][0] ), 
        .A4(\ram[3][0] ), .S0(n4244), .S1(n54), .Y(n4337) );
  MUX41X1_HVT U244 ( .A1(n4337), .A3(n4335), .A2(n4336), .A4(n4334), .S0(n4310), .S1(n4287), .Y(q[0]) );
  MUX41X1_HVT U245 ( .A1(\ram[12][1] ), .A3(\ram[14][1] ), .A2(\ram[13][1] ), 
        .A4(\ram[15][1] ), .S0(n4244), .S1(n54), .Y(n4338) );
  MUX41X1_HVT U246 ( .A1(\ram[8][1] ), .A3(\ram[10][1] ), .A2(\ram[9][1] ), 
        .A4(\ram[11][1] ), .S0(n4244), .S1(n54), .Y(n4339) );
  MUX41X1_HVT U247 ( .A1(\ram[4][1] ), .A3(\ram[6][1] ), .A2(\ram[5][1] ), 
        .A4(\ram[7][1] ), .S0(n4244), .S1(n54), .Y(n4340) );
  MUX41X1_HVT U248 ( .A1(\ram[0][1] ), .A3(\ram[2][1] ), .A2(\ram[1][1] ), 
        .A4(\ram[3][1] ), .S0(n4244), .S1(n54), .Y(n4341) );
  MUX41X1_HVT U249 ( .A1(n4341), .A3(n4339), .A2(n4340), .A4(n4338), .S0(n4310), .S1(n4287), .Y(q[1]) );
  MUX41X1_HVT U250 ( .A1(\ram[12][2] ), .A3(\ram[14][2] ), .A2(\ram[13][2] ), 
        .A4(\ram[15][2] ), .S0(n4244), .S1(n54), .Y(n4342) );
  MUX41X1_HVT U251 ( .A1(\ram[8][2] ), .A3(\ram[10][2] ), .A2(\ram[9][2] ), 
        .A4(\ram[11][2] ), .S0(n4244), .S1(n54), .Y(n4343) );
  MUX41X1_HVT U252 ( .A1(\ram[4][2] ), .A3(\ram[6][2] ), .A2(\ram[5][2] ), 
        .A4(\ram[7][2] ), .S0(n4245), .S1(n55), .Y(n4344) );
  MUX41X1_HVT U253 ( .A1(\ram[0][2] ), .A3(\ram[2][2] ), .A2(\ram[1][2] ), 
        .A4(\ram[3][2] ), .S0(n4245), .S1(n55), .Y(n4345) );
  MUX41X1_HVT U254 ( .A1(n4345), .A3(n4343), .A2(n4344), .A4(n4342), .S0(n4310), .S1(n4287), .Y(q[2]) );
  MUX41X1_HVT U255 ( .A1(\ram[12][3] ), .A3(\ram[14][3] ), .A2(\ram[13][3] ), 
        .A4(\ram[15][3] ), .S0(n4245), .S1(n55), .Y(n4346) );
  MUX41X1_HVT U256 ( .A1(\ram[8][3] ), .A3(\ram[10][3] ), .A2(\ram[9][3] ), 
        .A4(\ram[11][3] ), .S0(n4245), .S1(n55), .Y(n4347) );
  MUX41X1_HVT U257 ( .A1(\ram[4][3] ), .A3(\ram[6][3] ), .A2(\ram[5][3] ), 
        .A4(\ram[7][3] ), .S0(n4245), .S1(n55), .Y(n4348) );
  MUX41X1_HVT U258 ( .A1(\ram[0][3] ), .A3(\ram[2][3] ), .A2(\ram[1][3] ), 
        .A4(\ram[3][3] ), .S0(n4245), .S1(n55), .Y(n4349) );
  MUX41X1_HVT U259 ( .A1(n4349), .A3(n4347), .A2(n4348), .A4(n4346), .S0(n4310), .S1(n4287), .Y(q[3]) );
  MUX41X1_HVT U260 ( .A1(\ram[12][4] ), .A3(\ram[14][4] ), .A2(\ram[13][4] ), 
        .A4(\ram[15][4] ), .S0(n4245), .S1(n55), .Y(n4350) );
  MUX41X1_HVT U261 ( .A1(\ram[8][4] ), .A3(\ram[10][4] ), .A2(\ram[9][4] ), 
        .A4(\ram[11][4] ), .S0(n4245), .S1(n55), .Y(n4351) );
  MUX41X1_HVT U262 ( .A1(\ram[4][4] ), .A3(\ram[6][4] ), .A2(\ram[5][4] ), 
        .A4(\ram[7][4] ), .S0(n4245), .S1(n55), .Y(n4352) );
  MUX41X1_HVT U263 ( .A1(\ram[0][4] ), .A3(\ram[2][4] ), .A2(\ram[1][4] ), 
        .A4(\ram[3][4] ), .S0(n4245), .S1(n55), .Y(n4353) );
  MUX41X1_HVT U264 ( .A1(n4353), .A3(n4351), .A2(n4352), .A4(n4350), .S0(n4310), .S1(n4287), .Y(q[4]) );
  MUX41X1_HVT U265 ( .A1(\ram[12][5] ), .A3(\ram[14][5] ), .A2(\ram[13][5] ), 
        .A4(\ram[15][5] ), .S0(n4245), .S1(n55), .Y(n4354) );
  MUX41X1_HVT U266 ( .A1(\ram[8][5] ), .A3(\ram[10][5] ), .A2(\ram[9][5] ), 
        .A4(\ram[11][5] ), .S0(n4245), .S1(n55), .Y(n4355) );
  MUX41X1_HVT U267 ( .A1(\ram[4][5] ), .A3(\ram[6][5] ), .A2(\ram[5][5] ), 
        .A4(\ram[7][5] ), .S0(n4246), .S1(n56), .Y(n4356) );
  MUX41X1_HVT U268 ( .A1(\ram[0][5] ), .A3(\ram[2][5] ), .A2(\ram[1][5] ), 
        .A4(\ram[3][5] ), .S0(n4246), .S1(n56), .Y(n4357) );
  MUX41X1_HVT U269 ( .A1(n4357), .A3(n4355), .A2(n4356), .A4(n4354), .S0(n4310), .S1(n4287), .Y(q[5]) );
  MUX41X1_HVT U270 ( .A1(\ram[12][6] ), .A3(\ram[14][6] ), .A2(\ram[13][6] ), 
        .A4(\ram[15][6] ), .S0(n4246), .S1(n56), .Y(n4358) );
  MUX41X1_HVT U271 ( .A1(\ram[8][6] ), .A3(\ram[10][6] ), .A2(\ram[9][6] ), 
        .A4(\ram[11][6] ), .S0(n4246), .S1(n56), .Y(n4359) );
  MUX41X1_HVT U272 ( .A1(\ram[4][6] ), .A3(\ram[6][6] ), .A2(\ram[5][6] ), 
        .A4(\ram[7][6] ), .S0(n4246), .S1(n56), .Y(n4360) );
  MUX41X1_HVT U273 ( .A1(\ram[0][6] ), .A3(\ram[2][6] ), .A2(\ram[1][6] ), 
        .A4(\ram[3][6] ), .S0(n4246), .S1(n56), .Y(n4361) );
  MUX41X1_HVT U274 ( .A1(n4361), .A3(n4359), .A2(n4360), .A4(n4358), .S0(n4310), .S1(n4287), .Y(q[6]) );
  MUX41X1_HVT U275 ( .A1(\ram[12][7] ), .A3(\ram[14][7] ), .A2(\ram[13][7] ), 
        .A4(\ram[15][7] ), .S0(n4246), .S1(n56), .Y(n4362) );
  MUX41X1_HVT U276 ( .A1(\ram[8][7] ), .A3(\ram[10][7] ), .A2(\ram[9][7] ), 
        .A4(\ram[11][7] ), .S0(n4246), .S1(n56), .Y(n4363) );
  MUX41X1_HVT U277 ( .A1(\ram[4][7] ), .A3(\ram[6][7] ), .A2(\ram[5][7] ), 
        .A4(\ram[7][7] ), .S0(n4246), .S1(n56), .Y(n4364) );
  MUX41X1_HVT U278 ( .A1(\ram[0][7] ), .A3(\ram[2][7] ), .A2(\ram[1][7] ), 
        .A4(\ram[3][7] ), .S0(n4246), .S1(n56), .Y(n4365) );
  MUX41X1_HVT U279 ( .A1(n4365), .A3(n4363), .A2(n4364), .A4(n4362), .S0(n4310), .S1(n4287), .Y(q[7]) );
  MUX41X1_HVT U280 ( .A1(\ram[12][8] ), .A3(\ram[14][8] ), .A2(\ram[13][8] ), 
        .A4(\ram[15][8] ), .S0(n4246), .S1(n56), .Y(n4366) );
  MUX41X1_HVT U281 ( .A1(\ram[8][8] ), .A3(\ram[10][8] ), .A2(\ram[9][8] ), 
        .A4(\ram[11][8] ), .S0(n4246), .S1(n56), .Y(n4367) );
  MUX41X1_HVT U282 ( .A1(\ram[4][8] ), .A3(\ram[6][8] ), .A2(\ram[5][8] ), 
        .A4(\ram[7][8] ), .S0(n4247), .S1(n57), .Y(n4368) );
  MUX41X1_HVT U283 ( .A1(\ram[0][8] ), .A3(\ram[2][8] ), .A2(\ram[1][8] ), 
        .A4(\ram[3][8] ), .S0(n4247), .S1(n57), .Y(n4369) );
  MUX41X1_HVT U284 ( .A1(n4369), .A3(n4367), .A2(n4368), .A4(n4366), .S0(n4310), .S1(n4287), .Y(q[8]) );
  MUX41X1_HVT U285 ( .A1(\ram[12][9] ), .A3(\ram[14][9] ), .A2(\ram[13][9] ), 
        .A4(\ram[15][9] ), .S0(n4247), .S1(n57), .Y(n4370) );
  MUX41X1_HVT U286 ( .A1(\ram[8][9] ), .A3(\ram[10][9] ), .A2(\ram[9][9] ), 
        .A4(\ram[11][9] ), .S0(n4247), .S1(n57), .Y(n4371) );
  MUX41X1_HVT U287 ( .A1(\ram[4][9] ), .A3(\ram[6][9] ), .A2(\ram[5][9] ), 
        .A4(\ram[7][9] ), .S0(n4247), .S1(n57), .Y(n4372) );
  MUX41X1_HVT U288 ( .A1(\ram[0][9] ), .A3(\ram[2][9] ), .A2(\ram[1][9] ), 
        .A4(\ram[3][9] ), .S0(n4247), .S1(n57), .Y(n4373) );
  MUX41X1_HVT U289 ( .A1(n4373), .A3(n4371), .A2(n4372), .A4(n4370), .S0(n4310), .S1(n4287), .Y(q[9]) );
  MUX41X1_HVT U290 ( .A1(\ram[12][10] ), .A3(\ram[14][10] ), .A2(\ram[13][10] ), .A4(\ram[15][10] ), .S0(n4247), .S1(n57), .Y(n4374) );
  MUX41X1_HVT U291 ( .A1(\ram[8][10] ), .A3(\ram[10][10] ), .A2(\ram[9][10] ), 
        .A4(\ram[11][10] ), .S0(n4247), .S1(n57), .Y(n4375) );
  MUX41X1_HVT U292 ( .A1(\ram[4][10] ), .A3(\ram[6][10] ), .A2(\ram[5][10] ), 
        .A4(\ram[7][10] ), .S0(n4247), .S1(n57), .Y(n4376) );
  MUX41X1_HVT U293 ( .A1(\ram[0][10] ), .A3(\ram[2][10] ), .A2(\ram[1][10] ), 
        .A4(\ram[3][10] ), .S0(n4247), .S1(n57), .Y(n4377) );
  MUX41X1_HVT U294 ( .A1(n4377), .A3(n4375), .A2(n4376), .A4(n4374), .S0(n4310), .S1(n4287), .Y(q[10]) );
  MUX41X1_HVT U295 ( .A1(\ram[12][11] ), .A3(\ram[14][11] ), .A2(\ram[13][11] ), .A4(\ram[15][11] ), .S0(n4247), .S1(n57), .Y(n4378) );
  MUX41X1_HVT U296 ( .A1(\ram[8][11] ), .A3(\ram[10][11] ), .A2(\ram[9][11] ), 
        .A4(\ram[11][11] ), .S0(n4247), .S1(n57), .Y(n4379) );
  MUX41X1_HVT U297 ( .A1(\ram[4][11] ), .A3(\ram[6][11] ), .A2(\ram[5][11] ), 
        .A4(\ram[7][11] ), .S0(n4248), .S1(n58), .Y(n4380) );
  MUX41X1_HVT U298 ( .A1(\ram[0][11] ), .A3(\ram[2][11] ), .A2(\ram[1][11] ), 
        .A4(\ram[3][11] ), .S0(n4248), .S1(n58), .Y(n4381) );
  MUX41X1_HVT U299 ( .A1(n4381), .A3(n4379), .A2(n4380), .A4(n4378), .S0(n4310), .S1(n4287), .Y(q[11]) );
  MUX41X1_HVT U300 ( .A1(\ram[12][12] ), .A3(\ram[14][12] ), .A2(\ram[13][12] ), .A4(\ram[15][12] ), .S0(n4248), .S1(n58), .Y(n4382) );
  MUX41X1_HVT U301 ( .A1(\ram[8][12] ), .A3(\ram[10][12] ), .A2(\ram[9][12] ), 
        .A4(\ram[11][12] ), .S0(n4248), .S1(n58), .Y(n4383) );
  MUX41X1_HVT U302 ( .A1(\ram[4][12] ), .A3(\ram[6][12] ), .A2(\ram[5][12] ), 
        .A4(\ram[7][12] ), .S0(n4248), .S1(n58), .Y(n4384) );
  MUX41X1_HVT U303 ( .A1(\ram[0][12] ), .A3(\ram[2][12] ), .A2(\ram[1][12] ), 
        .A4(\ram[3][12] ), .S0(n4248), .S1(n58), .Y(n4385) );
  MUX41X1_HVT U304 ( .A1(n4385), .A3(n4383), .A2(n4384), .A4(n4382), .S0(n4311), .S1(n4288), .Y(q[12]) );
  MUX41X1_HVT U305 ( .A1(\ram[12][13] ), .A3(\ram[14][13] ), .A2(\ram[13][13] ), .A4(\ram[15][13] ), .S0(n4248), .S1(n58), .Y(n4386) );
  MUX41X1_HVT U306 ( .A1(\ram[8][13] ), .A3(\ram[10][13] ), .A2(\ram[9][13] ), 
        .A4(\ram[11][13] ), .S0(n4248), .S1(n58), .Y(n4387) );
  MUX41X1_HVT U307 ( .A1(\ram[4][13] ), .A3(\ram[6][13] ), .A2(\ram[5][13] ), 
        .A4(\ram[7][13] ), .S0(n4248), .S1(n58), .Y(n4388) );
  MUX41X1_HVT U308 ( .A1(\ram[0][13] ), .A3(\ram[2][13] ), .A2(\ram[1][13] ), 
        .A4(\ram[3][13] ), .S0(n4248), .S1(n58), .Y(n4389) );
  MUX41X1_HVT U309 ( .A1(n4389), .A3(n4387), .A2(n4388), .A4(n4386), .S0(n4311), .S1(n4288), .Y(q[13]) );
  MUX41X1_HVT U310 ( .A1(\ram[12][14] ), .A3(\ram[14][14] ), .A2(\ram[13][14] ), .A4(\ram[15][14] ), .S0(n4248), .S1(n58), .Y(n4390) );
  MUX41X1_HVT U311 ( .A1(\ram[8][14] ), .A3(\ram[10][14] ), .A2(\ram[9][14] ), 
        .A4(\ram[11][14] ), .S0(n4248), .S1(n58), .Y(n4391) );
  MUX41X1_HVT U312 ( .A1(\ram[4][14] ), .A3(\ram[6][14] ), .A2(\ram[5][14] ), 
        .A4(\ram[7][14] ), .S0(n4249), .S1(n59), .Y(n4392) );
  MUX41X1_HVT U313 ( .A1(\ram[0][14] ), .A3(\ram[2][14] ), .A2(\ram[1][14] ), 
        .A4(\ram[3][14] ), .S0(n4249), .S1(n59), .Y(n4393) );
  MUX41X1_HVT U314 ( .A1(n4393), .A3(n4391), .A2(n4392), .A4(n4390), .S0(n4311), .S1(n4288), .Y(q[14]) );
  MUX41X1_HVT U315 ( .A1(\ram[12][15] ), .A3(\ram[14][15] ), .A2(\ram[13][15] ), .A4(\ram[15][15] ), .S0(n4249), .S1(n59), .Y(n4394) );
  MUX41X1_HVT U316 ( .A1(\ram[8][15] ), .A3(\ram[10][15] ), .A2(\ram[9][15] ), 
        .A4(\ram[11][15] ), .S0(n4249), .S1(n59), .Y(n4395) );
  MUX41X1_HVT U317 ( .A1(\ram[4][15] ), .A3(\ram[6][15] ), .A2(\ram[5][15] ), 
        .A4(\ram[7][15] ), .S0(n4249), .S1(n59), .Y(n4396) );
  MUX41X1_HVT U318 ( .A1(\ram[0][15] ), .A3(\ram[2][15] ), .A2(\ram[1][15] ), 
        .A4(\ram[3][15] ), .S0(n4249), .S1(n59), .Y(n4397) );
  MUX41X1_HVT U319 ( .A1(n4397), .A3(n4395), .A2(n4396), .A4(n4394), .S0(n4311), .S1(n4288), .Y(q[15]) );
  MUX41X1_HVT U320 ( .A1(\ram[12][16] ), .A3(\ram[14][16] ), .A2(\ram[13][16] ), .A4(\ram[15][16] ), .S0(n4249), .S1(n59), .Y(n4398) );
  MUX41X1_HVT U321 ( .A1(\ram[8][16] ), .A3(\ram[10][16] ), .A2(\ram[9][16] ), 
        .A4(\ram[11][16] ), .S0(n4249), .S1(n59), .Y(n4399) );
  MUX41X1_HVT U322 ( .A1(\ram[4][16] ), .A3(\ram[6][16] ), .A2(\ram[5][16] ), 
        .A4(\ram[7][16] ), .S0(n4249), .S1(n59), .Y(n4400) );
  MUX41X1_HVT U323 ( .A1(\ram[0][16] ), .A3(\ram[2][16] ), .A2(\ram[1][16] ), 
        .A4(\ram[3][16] ), .S0(n4249), .S1(n59), .Y(n4401) );
  MUX41X1_HVT U324 ( .A1(n4401), .A3(n4399), .A2(n4400), .A4(n4398), .S0(n4311), .S1(n4288), .Y(q[16]) );
  MUX41X1_HVT U325 ( .A1(\ram[12][17] ), .A3(\ram[14][17] ), .A2(\ram[13][17] ), .A4(\ram[15][17] ), .S0(n4249), .S1(n59), .Y(n4402) );
  MUX41X1_HVT U326 ( .A1(\ram[8][17] ), .A3(\ram[10][17] ), .A2(\ram[9][17] ), 
        .A4(\ram[11][17] ), .S0(n4250), .S1(n60), .Y(n4403) );
  MUX41X1_HVT U327 ( .A1(\ram[4][17] ), .A3(\ram[6][17] ), .A2(\ram[5][17] ), 
        .A4(\ram[7][17] ), .S0(n4250), .S1(n60), .Y(n4404) );
  MUX41X1_HVT U328 ( .A1(\ram[0][17] ), .A3(\ram[2][17] ), .A2(\ram[1][17] ), 
        .A4(\ram[3][17] ), .S0(n4250), .S1(n60), .Y(n4405) );
  MUX41X1_HVT U329 ( .A1(n4405), .A3(n4403), .A2(n4404), .A4(n4402), .S0(n4311), .S1(n4288), .Y(q[17]) );
  MUX41X1_HVT U330 ( .A1(\ram[12][18] ), .A3(\ram[14][18] ), .A2(\ram[13][18] ), .A4(\ram[15][18] ), .S0(n4250), .S1(n60), .Y(n4406) );
  MUX41X1_HVT U331 ( .A1(\ram[8][18] ), .A3(\ram[10][18] ), .A2(\ram[9][18] ), 
        .A4(\ram[11][18] ), .S0(n4250), .S1(n60), .Y(n4407) );
  MUX41X1_HVT U332 ( .A1(\ram[4][18] ), .A3(\ram[6][18] ), .A2(\ram[5][18] ), 
        .A4(\ram[7][18] ), .S0(n4250), .S1(n60), .Y(n4408) );
  MUX41X1_HVT U333 ( .A1(\ram[0][18] ), .A3(\ram[2][18] ), .A2(\ram[1][18] ), 
        .A4(\ram[3][18] ), .S0(n4250), .S1(n60), .Y(n4409) );
  MUX41X1_HVT U334 ( .A1(n4409), .A3(n4407), .A2(n4408), .A4(n4406), .S0(n4311), .S1(n4288), .Y(q[18]) );
  MUX41X1_HVT U335 ( .A1(\ram[12][19] ), .A3(\ram[14][19] ), .A2(\ram[13][19] ), .A4(\ram[15][19] ), .S0(n4250), .S1(n60), .Y(n4410) );
  MUX41X1_HVT U336 ( .A1(\ram[8][19] ), .A3(\ram[10][19] ), .A2(\ram[9][19] ), 
        .A4(\ram[11][19] ), .S0(n4250), .S1(n60), .Y(n4411) );
  MUX41X1_HVT U337 ( .A1(\ram[4][19] ), .A3(\ram[6][19] ), .A2(\ram[5][19] ), 
        .A4(\ram[7][19] ), .S0(n4250), .S1(n60), .Y(n4412) );
  MUX41X1_HVT U338 ( .A1(\ram[0][19] ), .A3(\ram[2][19] ), .A2(\ram[1][19] ), 
        .A4(\ram[3][19] ), .S0(n4250), .S1(n60), .Y(n4413) );
  MUX41X1_HVT U339 ( .A1(n4413), .A3(n4411), .A2(n4412), .A4(n4410), .S0(n4311), .S1(n4288), .Y(q[19]) );
  MUX41X1_HVT U340 ( .A1(\ram[12][20] ), .A3(\ram[14][20] ), .A2(\ram[13][20] ), .A4(\ram[15][20] ), .S0(n4250), .S1(n60), .Y(n4414) );
  MUX41X1_HVT U341 ( .A1(\ram[8][20] ), .A3(\ram[10][20] ), .A2(\ram[9][20] ), 
        .A4(\ram[11][20] ), .S0(n4251), .S1(n4157), .Y(n4415) );
  MUX41X1_HVT U342 ( .A1(\ram[4][20] ), .A3(\ram[6][20] ), .A2(\ram[5][20] ), 
        .A4(\ram[7][20] ), .S0(n4251), .S1(n4157), .Y(n4416) );
  MUX41X1_HVT U343 ( .A1(\ram[0][20] ), .A3(\ram[2][20] ), .A2(\ram[1][20] ), 
        .A4(\ram[3][20] ), .S0(n4251), .S1(n4157), .Y(n4417) );
  MUX41X1_HVT U344 ( .A1(n4417), .A3(n4415), .A2(n4416), .A4(n4414), .S0(n4311), .S1(n4288), .Y(q[20]) );
  MUX41X1_HVT U345 ( .A1(\ram[12][21] ), .A3(\ram[14][21] ), .A2(\ram[13][21] ), .A4(\ram[15][21] ), .S0(n4251), .S1(n4157), .Y(n4418) );
  MUX41X1_HVT U346 ( .A1(\ram[8][21] ), .A3(\ram[10][21] ), .A2(\ram[9][21] ), 
        .A4(\ram[11][21] ), .S0(n4251), .S1(n4157), .Y(n4419) );
  MUX41X1_HVT U347 ( .A1(\ram[4][21] ), .A3(\ram[6][21] ), .A2(\ram[5][21] ), 
        .A4(\ram[7][21] ), .S0(n4251), .S1(n4157), .Y(n4420) );
  MUX41X1_HVT U348 ( .A1(\ram[0][21] ), .A3(\ram[2][21] ), .A2(\ram[1][21] ), 
        .A4(\ram[3][21] ), .S0(n4251), .S1(n4157), .Y(n4421) );
  MUX41X1_HVT U349 ( .A1(n4421), .A3(n4419), .A2(n4420), .A4(n4418), .S0(n4311), .S1(n4288), .Y(q[21]) );
  MUX41X1_HVT U350 ( .A1(\ram[12][22] ), .A3(\ram[14][22] ), .A2(\ram[13][22] ), .A4(\ram[15][22] ), .S0(n4251), .S1(n4157), .Y(n4422) );
  MUX41X1_HVT U351 ( .A1(\ram[8][22] ), .A3(\ram[10][22] ), .A2(\ram[9][22] ), 
        .A4(\ram[11][22] ), .S0(n4251), .S1(n4157), .Y(n4423) );
  MUX41X1_HVT U352 ( .A1(\ram[4][22] ), .A3(\ram[6][22] ), .A2(\ram[5][22] ), 
        .A4(\ram[7][22] ), .S0(n4251), .S1(n4157), .Y(n4424) );
  MUX41X1_HVT U353 ( .A1(\ram[0][22] ), .A3(\ram[2][22] ), .A2(\ram[1][22] ), 
        .A4(\ram[3][22] ), .S0(n4251), .S1(n4157), .Y(n4425) );
  MUX41X1_HVT U354 ( .A1(n4425), .A3(n4423), .A2(n4424), .A4(n4422), .S0(n4311), .S1(n4288), .Y(q[22]) );
  MUX41X1_HVT U355 ( .A1(\ram[12][23] ), .A3(\ram[14][23] ), .A2(\ram[13][23] ), .A4(\ram[15][23] ), .S0(n4251), .S1(n4157), .Y(n4426) );
  MUX41X1_HVT U356 ( .A1(\ram[8][23] ), .A3(\ram[10][23] ), .A2(\ram[9][23] ), 
        .A4(\ram[11][23] ), .S0(n4252), .S1(n4158), .Y(n4427) );
  MUX41X1_HVT U357 ( .A1(\ram[4][23] ), .A3(\ram[6][23] ), .A2(\ram[5][23] ), 
        .A4(\ram[7][23] ), .S0(n4252), .S1(n4158), .Y(n4428) );
  MUX41X1_HVT U358 ( .A1(\ram[0][23] ), .A3(\ram[2][23] ), .A2(\ram[1][23] ), 
        .A4(\ram[3][23] ), .S0(n4252), .S1(n4158), .Y(n4429) );
  MUX41X1_HVT U359 ( .A1(n4429), .A3(n4427), .A2(n4428), .A4(n4426), .S0(n4311), .S1(n4288), .Y(q[23]) );
  MUX41X1_HVT U360 ( .A1(\ram[12][24] ), .A3(\ram[14][24] ), .A2(\ram[13][24] ), .A4(\ram[15][24] ), .S0(n4252), .S1(n4158), .Y(n4430) );
  MUX41X1_HVT U361 ( .A1(\ram[8][24] ), .A3(\ram[10][24] ), .A2(\ram[9][24] ), 
        .A4(\ram[11][24] ), .S0(n4252), .S1(n4158), .Y(n4431) );
  MUX41X1_HVT U362 ( .A1(\ram[4][24] ), .A3(\ram[6][24] ), .A2(\ram[5][24] ), 
        .A4(\ram[7][24] ), .S0(n4252), .S1(n4158), .Y(n4432) );
  MUX41X1_HVT U363 ( .A1(\ram[0][24] ), .A3(\ram[2][24] ), .A2(\ram[1][24] ), 
        .A4(\ram[3][24] ), .S0(n4252), .S1(n4158), .Y(n4433) );
  MUX41X1_HVT U364 ( .A1(n4433), .A3(n4431), .A2(n4432), .A4(n4430), .S0(n4312), .S1(n4289), .Y(q[24]) );
  MUX41X1_HVT U365 ( .A1(\ram[12][25] ), .A3(\ram[14][25] ), .A2(\ram[13][25] ), .A4(\ram[15][25] ), .S0(n4252), .S1(n4158), .Y(n4434) );
  MUX41X1_HVT U366 ( .A1(\ram[8][25] ), .A3(\ram[10][25] ), .A2(\ram[9][25] ), 
        .A4(\ram[11][25] ), .S0(n4252), .S1(n4158), .Y(n4435) );
  MUX41X1_HVT U367 ( .A1(\ram[4][25] ), .A3(\ram[6][25] ), .A2(\ram[5][25] ), 
        .A4(\ram[7][25] ), .S0(n4252), .S1(n4158), .Y(n4436) );
  MUX41X1_HVT U368 ( .A1(\ram[0][25] ), .A3(\ram[2][25] ), .A2(\ram[1][25] ), 
        .A4(\ram[3][25] ), .S0(n4252), .S1(n4158), .Y(n4437) );
  MUX41X1_HVT U369 ( .A1(n4437), .A3(n4435), .A2(n4436), .A4(n4434), .S0(n4312), .S1(n4289), .Y(q[25]) );
  MUX41X1_HVT U370 ( .A1(\ram[12][26] ), .A3(\ram[14][26] ), .A2(\ram[13][26] ), .A4(\ram[15][26] ), .S0(n4252), .S1(n4158), .Y(n4438) );
  MUX41X1_HVT U371 ( .A1(\ram[8][26] ), .A3(\ram[10][26] ), .A2(\ram[9][26] ), 
        .A4(\ram[11][26] ), .S0(n4253), .S1(n4159), .Y(n4439) );
  MUX41X1_HVT U372 ( .A1(\ram[4][26] ), .A3(\ram[6][26] ), .A2(\ram[5][26] ), 
        .A4(\ram[7][26] ), .S0(n4253), .S1(n4159), .Y(n4440) );
  MUX41X1_HVT U373 ( .A1(\ram[0][26] ), .A3(\ram[2][26] ), .A2(\ram[1][26] ), 
        .A4(\ram[3][26] ), .S0(n4253), .S1(n4159), .Y(n4441) );
  MUX41X1_HVT U374 ( .A1(n4441), .A3(n4439), .A2(n4440), .A4(n4438), .S0(n4312), .S1(n4289), .Y(q[26]) );
  MUX41X1_HVT U375 ( .A1(\ram[12][27] ), .A3(\ram[14][27] ), .A2(\ram[13][27] ), .A4(\ram[15][27] ), .S0(n4253), .S1(n4159), .Y(n4442) );
  MUX41X1_HVT U376 ( .A1(\ram[8][27] ), .A3(\ram[10][27] ), .A2(\ram[9][27] ), 
        .A4(\ram[11][27] ), .S0(n4253), .S1(n4159), .Y(n4443) );
  MUX41X1_HVT U377 ( .A1(\ram[4][27] ), .A3(\ram[6][27] ), .A2(\ram[5][27] ), 
        .A4(\ram[7][27] ), .S0(n4253), .S1(n4159), .Y(n4444) );
  MUX41X1_HVT U378 ( .A1(\ram[0][27] ), .A3(\ram[2][27] ), .A2(\ram[1][27] ), 
        .A4(\ram[3][27] ), .S0(n4253), .S1(n4159), .Y(n4445) );
  MUX41X1_HVT U379 ( .A1(n4445), .A3(n4443), .A2(n4444), .A4(n4442), .S0(n4312), .S1(n4289), .Y(q[27]) );
  MUX41X1_HVT U380 ( .A1(\ram[12][28] ), .A3(\ram[14][28] ), .A2(\ram[13][28] ), .A4(\ram[15][28] ), .S0(n4253), .S1(n4159), .Y(n4446) );
  MUX41X1_HVT U381 ( .A1(\ram[8][28] ), .A3(\ram[10][28] ), .A2(\ram[9][28] ), 
        .A4(\ram[11][28] ), .S0(n4253), .S1(n4159), .Y(n4447) );
  MUX41X1_HVT U382 ( .A1(\ram[4][28] ), .A3(\ram[6][28] ), .A2(\ram[5][28] ), 
        .A4(\ram[7][28] ), .S0(n4253), .S1(n4159), .Y(n4448) );
  MUX41X1_HVT U383 ( .A1(\ram[0][28] ), .A3(\ram[2][28] ), .A2(\ram[1][28] ), 
        .A4(\ram[3][28] ), .S0(n4253), .S1(n4159), .Y(n4449) );
  MUX41X1_HVT U384 ( .A1(n4449), .A3(n4447), .A2(n4448), .A4(n4446), .S0(n4312), .S1(n4289), .Y(q[28]) );
  MUX41X1_HVT U385 ( .A1(\ram[12][29] ), .A3(\ram[14][29] ), .A2(\ram[13][29] ), .A4(\ram[15][29] ), .S0(n4253), .S1(n4159), .Y(n4450) );
  MUX41X1_HVT U386 ( .A1(\ram[8][29] ), .A3(\ram[10][29] ), .A2(\ram[9][29] ), 
        .A4(\ram[11][29] ), .S0(n4254), .S1(n4160), .Y(n4451) );
  MUX41X1_HVT U387 ( .A1(\ram[4][29] ), .A3(\ram[6][29] ), .A2(\ram[5][29] ), 
        .A4(\ram[7][29] ), .S0(n4254), .S1(n4160), .Y(n4452) );
  MUX41X1_HVT U388 ( .A1(\ram[0][29] ), .A3(\ram[2][29] ), .A2(\ram[1][29] ), 
        .A4(\ram[3][29] ), .S0(n4254), .S1(n4160), .Y(n4453) );
  MUX41X1_HVT U389 ( .A1(n4453), .A3(n4451), .A2(n4452), .A4(n4450), .S0(n4312), .S1(n4289), .Y(q[29]) );
  MUX41X1_HVT U390 ( .A1(\ram[12][30] ), .A3(\ram[14][30] ), .A2(\ram[13][30] ), .A4(\ram[15][30] ), .S0(n4254), .S1(n4160), .Y(n4454) );
  MUX41X1_HVT U391 ( .A1(\ram[8][30] ), .A3(\ram[10][30] ), .A2(\ram[9][30] ), 
        .A4(\ram[11][30] ), .S0(n4254), .S1(n4160), .Y(n4455) );
  MUX41X1_HVT U392 ( .A1(\ram[4][30] ), .A3(\ram[6][30] ), .A2(\ram[5][30] ), 
        .A4(\ram[7][30] ), .S0(n4254), .S1(n4160), .Y(n4456) );
  MUX41X1_HVT U393 ( .A1(\ram[0][30] ), .A3(\ram[2][30] ), .A2(\ram[1][30] ), 
        .A4(\ram[3][30] ), .S0(n4254), .S1(n4160), .Y(n4457) );
  MUX41X1_HVT U394 ( .A1(n4457), .A3(n4455), .A2(n4456), .A4(n4454), .S0(n4312), .S1(n4289), .Y(q[30]) );
  MUX41X1_HVT U395 ( .A1(\ram[12][31] ), .A3(\ram[14][31] ), .A2(\ram[13][31] ), .A4(\ram[15][31] ), .S0(n4254), .S1(n4160), .Y(n4458) );
  MUX41X1_HVT U396 ( .A1(\ram[8][31] ), .A3(\ram[10][31] ), .A2(\ram[9][31] ), 
        .A4(\ram[11][31] ), .S0(n4254), .S1(n4160), .Y(n4459) );
  MUX41X1_HVT U397 ( .A1(\ram[4][31] ), .A3(\ram[6][31] ), .A2(\ram[5][31] ), 
        .A4(\ram[7][31] ), .S0(n4254), .S1(n4160), .Y(n4460) );
  MUX41X1_HVT U398 ( .A1(\ram[0][31] ), .A3(\ram[2][31] ), .A2(\ram[1][31] ), 
        .A4(\ram[3][31] ), .S0(n4254), .S1(n4160), .Y(n4461) );
  MUX41X1_HVT U399 ( .A1(n4461), .A3(n4459), .A2(n4460), .A4(n4458), .S0(n4312), .S1(n4289), .Y(q[31]) );
  MUX41X1_HVT U400 ( .A1(\ram[12][32] ), .A3(\ram[14][32] ), .A2(\ram[13][32] ), .A4(\ram[15][32] ), .S0(n4254), .S1(n4160), .Y(n4462) );
  MUX41X1_HVT U401 ( .A1(\ram[8][32] ), .A3(\ram[10][32] ), .A2(\ram[9][32] ), 
        .A4(\ram[11][32] ), .S0(n4239), .S1(n49), .Y(n4463) );
  MUX41X1_HVT U402 ( .A1(\ram[4][32] ), .A3(\ram[6][32] ), .A2(\ram[5][32] ), 
        .A4(\ram[7][32] ), .S0(n4233), .S1(n43), .Y(n4464) );
  MUX41X1_HVT U403 ( .A1(\ram[0][32] ), .A3(\ram[2][32] ), .A2(\ram[1][32] ), 
        .A4(\ram[3][32] ), .S0(n4233), .S1(n43), .Y(n4465) );
  MUX41X1_HVT U404 ( .A1(n4465), .A3(n4463), .A2(n4464), .A4(n4462), .S0(n4312), .S1(n4289), .Y(q[32]) );
  MUX41X1_HVT U405 ( .A1(\ram[12][33] ), .A3(\ram[14][33] ), .A2(\ram[13][33] ), .A4(\ram[15][33] ), .S0(n4233), .S1(n43), .Y(n4466) );
  MUX41X1_HVT U406 ( .A1(\ram[8][33] ), .A3(\ram[10][33] ), .A2(\ram[9][33] ), 
        .A4(\ram[11][33] ), .S0(n4234), .S1(n44), .Y(n4467) );
  MUX41X1_HVT U407 ( .A1(\ram[4][33] ), .A3(\ram[6][33] ), .A2(\ram[5][33] ), 
        .A4(\ram[7][33] ), .S0(n4234), .S1(n44), .Y(n4468) );
  MUX41X1_HVT U408 ( .A1(\ram[0][33] ), .A3(\ram[2][33] ), .A2(\ram[1][33] ), 
        .A4(\ram[3][33] ), .S0(n4234), .S1(n44), .Y(n4469) );
  MUX41X1_HVT U409 ( .A1(n4469), .A3(n4467), .A2(n4468), .A4(n4466), .S0(n4312), .S1(n4289), .Y(q[33]) );
  MUX41X1_HVT U410 ( .A1(\ram[12][34] ), .A3(\ram[14][34] ), .A2(\ram[13][34] ), .A4(\ram[15][34] ), .S0(n4234), .S1(n44), .Y(n4470) );
  MUX41X1_HVT U411 ( .A1(\ram[8][34] ), .A3(\ram[10][34] ), .A2(\ram[9][34] ), 
        .A4(\ram[11][34] ), .S0(n4234), .S1(n44), .Y(n4471) );
  MUX41X1_HVT U412 ( .A1(\ram[4][34] ), .A3(\ram[6][34] ), .A2(\ram[5][34] ), 
        .A4(\ram[7][34] ), .S0(n4234), .S1(n44), .Y(n4472) );
  MUX41X1_HVT U413 ( .A1(\ram[0][34] ), .A3(\ram[2][34] ), .A2(\ram[1][34] ), 
        .A4(\ram[3][34] ), .S0(n4234), .S1(n44), .Y(n4473) );
  MUX41X1_HVT U414 ( .A1(n4473), .A3(n4471), .A2(n4472), .A4(n4470), .S0(n4312), .S1(n4289), .Y(q[34]) );
  MUX41X1_HVT U415 ( .A1(\ram[12][35] ), .A3(\ram[14][35] ), .A2(\ram[13][35] ), .A4(\ram[15][35] ), .S0(n4234), .S1(n44), .Y(n4474) );
  MUX41X1_HVT U416 ( .A1(\ram[8][35] ), .A3(\ram[10][35] ), .A2(\ram[9][35] ), 
        .A4(\ram[11][35] ), .S0(n4234), .S1(n44), .Y(n4475) );
  MUX41X1_HVT U417 ( .A1(\ram[4][35] ), .A3(\ram[6][35] ), .A2(\ram[5][35] ), 
        .A4(\ram[7][35] ), .S0(n4234), .S1(n44), .Y(n4476) );
  MUX41X1_HVT U418 ( .A1(\ram[0][35] ), .A3(\ram[2][35] ), .A2(\ram[1][35] ), 
        .A4(\ram[3][35] ), .S0(n4234), .S1(n44), .Y(n4477) );
  MUX41X1_HVT U419 ( .A1(n4477), .A3(n4475), .A2(n4476), .A4(n4474), .S0(n4312), .S1(n4289), .Y(q[35]) );
  MUX41X1_HVT U420 ( .A1(\ram[12][36] ), .A3(\ram[14][36] ), .A2(\ram[13][36] ), .A4(\ram[15][36] ), .S0(n4234), .S1(n44), .Y(n4478) );
  MUX41X1_HVT U421 ( .A1(\ram[8][36] ), .A3(\ram[10][36] ), .A2(\ram[9][36] ), 
        .A4(\ram[11][36] ), .S0(n4235), .S1(n45), .Y(n4479) );
  MUX41X1_HVT U422 ( .A1(\ram[4][36] ), .A3(\ram[6][36] ), .A2(\ram[5][36] ), 
        .A4(\ram[7][36] ), .S0(n4235), .S1(n45), .Y(n4480) );
  MUX41X1_HVT U423 ( .A1(\ram[0][36] ), .A3(\ram[2][36] ), .A2(\ram[1][36] ), 
        .A4(\ram[3][36] ), .S0(n4235), .S1(n45), .Y(n4481) );
  MUX41X1_HVT U424 ( .A1(n4481), .A3(n4479), .A2(n4480), .A4(n4478), .S0(n4313), .S1(n4290), .Y(q[36]) );
  MUX41X1_HVT U425 ( .A1(\ram[12][37] ), .A3(\ram[14][37] ), .A2(\ram[13][37] ), .A4(\ram[15][37] ), .S0(n4235), .S1(n45), .Y(n4482) );
  MUX41X1_HVT U426 ( .A1(\ram[8][37] ), .A3(\ram[10][37] ), .A2(\ram[9][37] ), 
        .A4(\ram[11][37] ), .S0(n4235), .S1(n45), .Y(n4483) );
  MUX41X1_HVT U427 ( .A1(\ram[4][37] ), .A3(\ram[6][37] ), .A2(\ram[5][37] ), 
        .A4(\ram[7][37] ), .S0(n4235), .S1(n45), .Y(n4484) );
  MUX41X1_HVT U428 ( .A1(\ram[0][37] ), .A3(\ram[2][37] ), .A2(\ram[1][37] ), 
        .A4(\ram[3][37] ), .S0(n4235), .S1(n45), .Y(n4485) );
  MUX41X1_HVT U429 ( .A1(n4485), .A3(n4483), .A2(n4484), .A4(n4482), .S0(n4313), .S1(n4290), .Y(q[37]) );
  MUX41X1_HVT U430 ( .A1(\ram[12][38] ), .A3(\ram[14][38] ), .A2(\ram[13][38] ), .A4(\ram[15][38] ), .S0(n4235), .S1(n45), .Y(n4486) );
  MUX41X1_HVT U431 ( .A1(\ram[8][38] ), .A3(\ram[10][38] ), .A2(\ram[9][38] ), 
        .A4(\ram[11][38] ), .S0(n4235), .S1(n45), .Y(n4487) );
  MUX41X1_HVT U432 ( .A1(\ram[4][38] ), .A3(\ram[6][38] ), .A2(\ram[5][38] ), 
        .A4(\ram[7][38] ), .S0(n4235), .S1(n45), .Y(n4488) );
  MUX41X1_HVT U433 ( .A1(\ram[0][38] ), .A3(\ram[2][38] ), .A2(\ram[1][38] ), 
        .A4(\ram[3][38] ), .S0(n4235), .S1(n45), .Y(n4489) );
  MUX41X1_HVT U434 ( .A1(n4489), .A3(n4487), .A2(n4488), .A4(n4486), .S0(n4313), .S1(n4290), .Y(q[38]) );
  MUX41X1_HVT U435 ( .A1(\ram[12][39] ), .A3(\ram[14][39] ), .A2(\ram[13][39] ), .A4(\ram[15][39] ), .S0(n4235), .S1(n45), .Y(n4490) );
  MUX41X1_HVT U436 ( .A1(\ram[8][39] ), .A3(\ram[10][39] ), .A2(\ram[9][39] ), 
        .A4(\ram[11][39] ), .S0(n4236), .S1(n46), .Y(n4491) );
  MUX41X1_HVT U437 ( .A1(\ram[4][39] ), .A3(\ram[6][39] ), .A2(\ram[5][39] ), 
        .A4(\ram[7][39] ), .S0(n4236), .S1(n46), .Y(n4492) );
  MUX41X1_HVT U438 ( .A1(\ram[0][39] ), .A3(\ram[2][39] ), .A2(\ram[1][39] ), 
        .A4(\ram[3][39] ), .S0(n4236), .S1(n46), .Y(n4493) );
  MUX41X1_HVT U439 ( .A1(n4493), .A3(n4491), .A2(n4492), .A4(n4490), .S0(n4313), .S1(n4290), .Y(q[39]) );
  MUX41X1_HVT U440 ( .A1(\ram[12][40] ), .A3(\ram[14][40] ), .A2(\ram[13][40] ), .A4(\ram[15][40] ), .S0(n4236), .S1(n46), .Y(n4494) );
  MUX41X1_HVT U441 ( .A1(\ram[8][40] ), .A3(\ram[10][40] ), .A2(\ram[9][40] ), 
        .A4(\ram[11][40] ), .S0(n4236), .S1(n46), .Y(n4495) );
  MUX41X1_HVT U442 ( .A1(\ram[4][40] ), .A3(\ram[6][40] ), .A2(\ram[5][40] ), 
        .A4(\ram[7][40] ), .S0(n4236), .S1(n46), .Y(n4496) );
  MUX41X1_HVT U443 ( .A1(\ram[0][40] ), .A3(\ram[2][40] ), .A2(\ram[1][40] ), 
        .A4(\ram[3][40] ), .S0(n4236), .S1(n46), .Y(n4497) );
  MUX41X1_HVT U444 ( .A1(n4497), .A3(n4495), .A2(n4496), .A4(n4494), .S0(n4313), .S1(n4290), .Y(q[40]) );
  MUX41X1_HVT U445 ( .A1(\ram[12][41] ), .A3(\ram[14][41] ), .A2(\ram[13][41] ), .A4(\ram[15][41] ), .S0(n4236), .S1(n46), .Y(n4498) );
  MUX41X1_HVT U446 ( .A1(\ram[8][41] ), .A3(\ram[10][41] ), .A2(\ram[9][41] ), 
        .A4(\ram[11][41] ), .S0(n4236), .S1(n46), .Y(n4499) );
  MUX41X1_HVT U447 ( .A1(\ram[4][41] ), .A3(\ram[6][41] ), .A2(\ram[5][41] ), 
        .A4(\ram[7][41] ), .S0(n4236), .S1(n46), .Y(n4500) );
  MUX41X1_HVT U448 ( .A1(\ram[0][41] ), .A3(\ram[2][41] ), .A2(\ram[1][41] ), 
        .A4(\ram[3][41] ), .S0(n4236), .S1(n46), .Y(n4501) );
  MUX41X1_HVT U449 ( .A1(n4501), .A3(n4499), .A2(n4500), .A4(n4498), .S0(n4313), .S1(n4290), .Y(q[41]) );
  MUX41X1_HVT U450 ( .A1(\ram[12][42] ), .A3(\ram[14][42] ), .A2(\ram[13][42] ), .A4(\ram[15][42] ), .S0(n4236), .S1(n46), .Y(n4502) );
  MUX41X1_HVT U451 ( .A1(\ram[8][42] ), .A3(\ram[10][42] ), .A2(\ram[9][42] ), 
        .A4(\ram[11][42] ), .S0(n4237), .S1(n47), .Y(n4503) );
  MUX41X1_HVT U452 ( .A1(\ram[4][42] ), .A3(\ram[6][42] ), .A2(\ram[5][42] ), 
        .A4(\ram[7][42] ), .S0(n4237), .S1(n47), .Y(n4504) );
  MUX41X1_HVT U453 ( .A1(\ram[0][42] ), .A3(\ram[2][42] ), .A2(\ram[1][42] ), 
        .A4(\ram[3][42] ), .S0(n4237), .S1(n47), .Y(n4505) );
  MUX41X1_HVT U454 ( .A1(n4505), .A3(n4503), .A2(n4504), .A4(n4502), .S0(n4313), .S1(n4290), .Y(q[42]) );
  MUX41X1_HVT U455 ( .A1(\ram[12][43] ), .A3(\ram[14][43] ), .A2(\ram[13][43] ), .A4(\ram[15][43] ), .S0(n4237), .S1(n47), .Y(n4506) );
  MUX41X1_HVT U456 ( .A1(\ram[8][43] ), .A3(\ram[10][43] ), .A2(\ram[9][43] ), 
        .A4(\ram[11][43] ), .S0(n4237), .S1(n47), .Y(n4507) );
  MUX41X1_HVT U457 ( .A1(\ram[4][43] ), .A3(\ram[6][43] ), .A2(\ram[5][43] ), 
        .A4(\ram[7][43] ), .S0(n4237), .S1(n47), .Y(n4508) );
  MUX41X1_HVT U458 ( .A1(\ram[0][43] ), .A3(\ram[2][43] ), .A2(\ram[1][43] ), 
        .A4(\ram[3][43] ), .S0(n4237), .S1(n47), .Y(n4509) );
  MUX41X1_HVT U459 ( .A1(n4509), .A3(n4507), .A2(n4508), .A4(n4506), .S0(n4313), .S1(n4290), .Y(q[43]) );
  MUX41X1_HVT U460 ( .A1(\ram[12][44] ), .A3(\ram[14][44] ), .A2(\ram[13][44] ), .A4(\ram[15][44] ), .S0(n4237), .S1(n47), .Y(n4510) );
  MUX41X1_HVT U461 ( .A1(\ram[8][44] ), .A3(\ram[10][44] ), .A2(\ram[9][44] ), 
        .A4(\ram[11][44] ), .S0(n4237), .S1(n47), .Y(n4511) );
  MUX41X1_HVT U462 ( .A1(\ram[4][44] ), .A3(\ram[6][44] ), .A2(\ram[5][44] ), 
        .A4(\ram[7][44] ), .S0(n4237), .S1(n47), .Y(n4512) );
  MUX41X1_HVT U463 ( .A1(\ram[0][44] ), .A3(\ram[2][44] ), .A2(\ram[1][44] ), 
        .A4(\ram[3][44] ), .S0(n4237), .S1(n47), .Y(n4513) );
  MUX41X1_HVT U464 ( .A1(n4513), .A3(n4511), .A2(n4512), .A4(n4510), .S0(n4313), .S1(n4290), .Y(q[44]) );
  MUX41X1_HVT U465 ( .A1(\ram[12][45] ), .A3(\ram[14][45] ), .A2(\ram[13][45] ), .A4(\ram[15][45] ), .S0(n4237), .S1(n47), .Y(n4514) );
  MUX41X1_HVT U466 ( .A1(\ram[8][45] ), .A3(\ram[10][45] ), .A2(\ram[9][45] ), 
        .A4(\ram[11][45] ), .S0(n4238), .S1(n48), .Y(n4515) );
  MUX41X1_HVT U467 ( .A1(\ram[4][45] ), .A3(\ram[6][45] ), .A2(\ram[5][45] ), 
        .A4(\ram[7][45] ), .S0(n4238), .S1(n48), .Y(n4516) );
  MUX41X1_HVT U468 ( .A1(\ram[0][45] ), .A3(\ram[2][45] ), .A2(\ram[1][45] ), 
        .A4(\ram[3][45] ), .S0(n4238), .S1(n48), .Y(n4517) );
  MUX41X1_HVT U469 ( .A1(n4517), .A3(n4515), .A2(n4516), .A4(n4514), .S0(n4313), .S1(n4290), .Y(q[45]) );
  MUX41X1_HVT U470 ( .A1(\ram[12][46] ), .A3(\ram[14][46] ), .A2(\ram[13][46] ), .A4(\ram[15][46] ), .S0(n4238), .S1(n48), .Y(n4518) );
  MUX41X1_HVT U471 ( .A1(\ram[8][46] ), .A3(\ram[10][46] ), .A2(\ram[9][46] ), 
        .A4(\ram[11][46] ), .S0(n4238), .S1(n48), .Y(n4519) );
  MUX41X1_HVT U472 ( .A1(\ram[4][46] ), .A3(\ram[6][46] ), .A2(\ram[5][46] ), 
        .A4(\ram[7][46] ), .S0(n4238), .S1(n48), .Y(n4520) );
  MUX41X1_HVT U473 ( .A1(\ram[0][46] ), .A3(\ram[2][46] ), .A2(\ram[1][46] ), 
        .A4(\ram[3][46] ), .S0(n4238), .S1(n48), .Y(n4521) );
  MUX41X1_HVT U474 ( .A1(n4521), .A3(n4519), .A2(n4520), .A4(n4518), .S0(n4313), .S1(n4290), .Y(q[46]) );
  MUX41X1_HVT U475 ( .A1(\ram[12][47] ), .A3(\ram[14][47] ), .A2(\ram[13][47] ), .A4(\ram[15][47] ), .S0(n4238), .S1(n48), .Y(n4522) );
  MUX41X1_HVT U476 ( .A1(\ram[8][47] ), .A3(\ram[10][47] ), .A2(\ram[9][47] ), 
        .A4(\ram[11][47] ), .S0(n4238), .S1(n48), .Y(n4523) );
  MUX41X1_HVT U477 ( .A1(\ram[4][47] ), .A3(\ram[6][47] ), .A2(\ram[5][47] ), 
        .A4(\ram[7][47] ), .S0(n4238), .S1(n48), .Y(n4524) );
  MUX41X1_HVT U478 ( .A1(\ram[0][47] ), .A3(\ram[2][47] ), .A2(\ram[1][47] ), 
        .A4(\ram[3][47] ), .S0(n4238), .S1(n48), .Y(n4525) );
  MUX41X1_HVT U479 ( .A1(n4525), .A3(n4523), .A2(n4524), .A4(n4522), .S0(n4313), .S1(n4290), .Y(q[47]) );
  MUX41X1_HVT U480 ( .A1(\ram[12][48] ), .A3(\ram[14][48] ), .A2(\ram[13][48] ), .A4(\ram[15][48] ), .S0(n4238), .S1(n48), .Y(n4526) );
  MUX41X1_HVT U481 ( .A1(\ram[8][48] ), .A3(\ram[10][48] ), .A2(\ram[9][48] ), 
        .A4(\ram[11][48] ), .S0(n4239), .S1(n49), .Y(n4527) );
  MUX41X1_HVT U482 ( .A1(\ram[4][48] ), .A3(\ram[6][48] ), .A2(\ram[5][48] ), 
        .A4(\ram[7][48] ), .S0(n4239), .S1(n49), .Y(n4528) );
  MUX41X1_HVT U483 ( .A1(\ram[0][48] ), .A3(\ram[2][48] ), .A2(\ram[1][48] ), 
        .A4(\ram[3][48] ), .S0(n4239), .S1(n49), .Y(n4529) );
  MUX41X1_HVT U484 ( .A1(n4529), .A3(n4527), .A2(n4528), .A4(n4526), .S0(n4314), .S1(n4291), .Y(q[48]) );
  MUX41X1_HVT U485 ( .A1(\ram[12][49] ), .A3(\ram[14][49] ), .A2(\ram[13][49] ), .A4(\ram[15][49] ), .S0(n4239), .S1(n49), .Y(n4530) );
  MUX41X1_HVT U486 ( .A1(\ram[8][49] ), .A3(\ram[10][49] ), .A2(\ram[9][49] ), 
        .A4(\ram[11][49] ), .S0(n4239), .S1(n49), .Y(n4531) );
  MUX41X1_HVT U487 ( .A1(\ram[4][49] ), .A3(\ram[6][49] ), .A2(\ram[5][49] ), 
        .A4(\ram[7][49] ), .S0(n4239), .S1(n49), .Y(n4532) );
  MUX41X1_HVT U488 ( .A1(\ram[0][49] ), .A3(\ram[2][49] ), .A2(\ram[1][49] ), 
        .A4(\ram[3][49] ), .S0(n4239), .S1(n49), .Y(n4533) );
  MUX41X1_HVT U489 ( .A1(n4533), .A3(n4531), .A2(n4532), .A4(n4530), .S0(n4314), .S1(n4291), .Y(q[49]) );
  MUX41X1_HVT U490 ( .A1(\ram[12][50] ), .A3(\ram[14][50] ), .A2(\ram[13][50] ), .A4(\ram[15][50] ), .S0(n4239), .S1(n49), .Y(n4534) );
  MUX41X1_HVT U491 ( .A1(\ram[8][50] ), .A3(\ram[10][50] ), .A2(\ram[9][50] ), 
        .A4(\ram[11][50] ), .S0(n4239), .S1(n49), .Y(n4535) );
  MUX41X1_HVT U492 ( .A1(\ram[4][50] ), .A3(\ram[6][50] ), .A2(\ram[5][50] ), 
        .A4(\ram[7][50] ), .S0(n4239), .S1(n49), .Y(n4536) );
  MUX41X1_HVT U493 ( .A1(\ram[0][50] ), .A3(\ram[2][50] ), .A2(\ram[1][50] ), 
        .A4(\ram[3][50] ), .S0(n4239), .S1(n49), .Y(n4537) );
  MUX41X1_HVT U494 ( .A1(n4537), .A3(n4535), .A2(n4536), .A4(n4534), .S0(n4314), .S1(n4291), .Y(q[50]) );
  MUX41X1_HVT U495 ( .A1(\ram[12][51] ), .A3(\ram[14][51] ), .A2(\ram[13][51] ), .A4(\ram[15][51] ), .S0(n4240), .S1(n50), .Y(n4538) );
  MUX41X1_HVT U496 ( .A1(\ram[8][51] ), .A3(\ram[10][51] ), .A2(\ram[9][51] ), 
        .A4(\ram[11][51] ), .S0(n4240), .S1(n50), .Y(n4539) );
  MUX41X1_HVT U497 ( .A1(\ram[4][51] ), .A3(\ram[6][51] ), .A2(\ram[5][51] ), 
        .A4(\ram[7][51] ), .S0(n4240), .S1(n50), .Y(n4540) );
  MUX41X1_HVT U498 ( .A1(\ram[0][51] ), .A3(\ram[2][51] ), .A2(\ram[1][51] ), 
        .A4(\ram[3][51] ), .S0(n4240), .S1(n50), .Y(n4541) );
  MUX41X1_HVT U499 ( .A1(n4541), .A3(n4539), .A2(n4540), .A4(n4538), .S0(n4314), .S1(n4291), .Y(q[51]) );
  MUX41X1_HVT U500 ( .A1(\ram[12][52] ), .A3(\ram[14][52] ), .A2(\ram[13][52] ), .A4(\ram[15][52] ), .S0(n4240), .S1(n50), .Y(n4542) );
  MUX41X1_HVT U501 ( .A1(\ram[8][52] ), .A3(\ram[10][52] ), .A2(\ram[9][52] ), 
        .A4(\ram[11][52] ), .S0(n4240), .S1(n50), .Y(n4543) );
  MUX41X1_HVT U502 ( .A1(\ram[4][52] ), .A3(\ram[6][52] ), .A2(\ram[5][52] ), 
        .A4(\ram[7][52] ), .S0(n4240), .S1(n50), .Y(n4544) );
  MUX41X1_HVT U503 ( .A1(\ram[0][52] ), .A3(\ram[2][52] ), .A2(\ram[1][52] ), 
        .A4(\ram[3][52] ), .S0(n4240), .S1(n50), .Y(n4545) );
  MUX41X1_HVT U504 ( .A1(n4545), .A3(n4543), .A2(n4544), .A4(n4542), .S0(n4314), .S1(n4291), .Y(q[52]) );
  MUX41X1_HVT U505 ( .A1(\ram[12][53] ), .A3(\ram[14][53] ), .A2(\ram[13][53] ), .A4(\ram[15][53] ), .S0(n4240), .S1(n50), .Y(n4546) );
  MUX41X1_HVT U506 ( .A1(\ram[8][53] ), .A3(\ram[10][53] ), .A2(\ram[9][53] ), 
        .A4(\ram[11][53] ), .S0(n4240), .S1(n50), .Y(n4547) );
  MUX41X1_HVT U507 ( .A1(\ram[4][53] ), .A3(\ram[6][53] ), .A2(\ram[5][53] ), 
        .A4(\ram[7][53] ), .S0(n4240), .S1(n50), .Y(n4548) );
  MUX41X1_HVT U508 ( .A1(\ram[0][53] ), .A3(\ram[2][53] ), .A2(\ram[1][53] ), 
        .A4(\ram[3][53] ), .S0(n4240), .S1(n50), .Y(n4549) );
  MUX41X1_HVT U509 ( .A1(n4549), .A3(n4547), .A2(n4548), .A4(n4546), .S0(n4314), .S1(n4291), .Y(q[53]) );
  MUX41X1_HVT U510 ( .A1(\ram[12][54] ), .A3(\ram[14][54] ), .A2(\ram[13][54] ), .A4(\ram[15][54] ), .S0(n4241), .S1(n51), .Y(n4550) );
  MUX41X1_HVT U511 ( .A1(\ram[8][54] ), .A3(\ram[10][54] ), .A2(\ram[9][54] ), 
        .A4(\ram[11][54] ), .S0(n4241), .S1(n51), .Y(n4551) );
  MUX41X1_HVT U512 ( .A1(\ram[4][54] ), .A3(\ram[6][54] ), .A2(\ram[5][54] ), 
        .A4(\ram[7][54] ), .S0(n4241), .S1(n51), .Y(n4552) );
  MUX41X1_HVT U513 ( .A1(\ram[0][54] ), .A3(\ram[2][54] ), .A2(\ram[1][54] ), 
        .A4(\ram[3][54] ), .S0(n4241), .S1(n51), .Y(n4553) );
  MUX41X1_HVT U514 ( .A1(n4553), .A3(n4551), .A2(n4552), .A4(n4550), .S0(n4314), .S1(n4291), .Y(q[54]) );
  MUX41X1_HVT U515 ( .A1(\ram[12][55] ), .A3(\ram[14][55] ), .A2(\ram[13][55] ), .A4(\ram[15][55] ), .S0(n4241), .S1(n51), .Y(n4554) );
  MUX41X1_HVT U516 ( .A1(\ram[8][55] ), .A3(\ram[10][55] ), .A2(\ram[9][55] ), 
        .A4(\ram[11][55] ), .S0(n4241), .S1(n51), .Y(n4555) );
  MUX41X1_HVT U517 ( .A1(\ram[4][55] ), .A3(\ram[6][55] ), .A2(\ram[5][55] ), 
        .A4(\ram[7][55] ), .S0(n4241), .S1(n51), .Y(n4556) );
  MUX41X1_HVT U518 ( .A1(\ram[0][55] ), .A3(\ram[2][55] ), .A2(\ram[1][55] ), 
        .A4(\ram[3][55] ), .S0(n4241), .S1(n51), .Y(n4557) );
  MUX41X1_HVT U519 ( .A1(n4557), .A3(n4555), .A2(n4556), .A4(n4554), .S0(n4314), .S1(n4291), .Y(q[55]) );
  MUX41X1_HVT U520 ( .A1(\ram[12][56] ), .A3(\ram[14][56] ), .A2(\ram[13][56] ), .A4(\ram[15][56] ), .S0(n4241), .S1(n51), .Y(n4558) );
  MUX41X1_HVT U521 ( .A1(\ram[8][56] ), .A3(\ram[10][56] ), .A2(\ram[9][56] ), 
        .A4(\ram[11][56] ), .S0(n4241), .S1(n51), .Y(n4559) );
  MUX41X1_HVT U522 ( .A1(\ram[4][56] ), .A3(\ram[6][56] ), .A2(\ram[5][56] ), 
        .A4(\ram[7][56] ), .S0(n4241), .S1(n51), .Y(n4560) );
  MUX41X1_HVT U523 ( .A1(\ram[0][56] ), .A3(\ram[2][56] ), .A2(\ram[1][56] ), 
        .A4(\ram[3][56] ), .S0(n4241), .S1(n51), .Y(n4561) );
  MUX41X1_HVT U524 ( .A1(n4561), .A3(n4559), .A2(n4560), .A4(n4558), .S0(n4314), .S1(n4291), .Y(q[56]) );
  MUX41X1_HVT U525 ( .A1(\ram[12][57] ), .A3(\ram[14][57] ), .A2(\ram[13][57] ), .A4(\ram[15][57] ), .S0(n4242), .S1(n52), .Y(n4562) );
  MUX41X1_HVT U526 ( .A1(\ram[8][57] ), .A3(\ram[10][57] ), .A2(\ram[9][57] ), 
        .A4(\ram[11][57] ), .S0(n4242), .S1(n52), .Y(n4563) );
  MUX41X1_HVT U527 ( .A1(\ram[4][57] ), .A3(\ram[6][57] ), .A2(\ram[5][57] ), 
        .A4(\ram[7][57] ), .S0(n4242), .S1(n52), .Y(n4564) );
  MUX41X1_HVT U528 ( .A1(\ram[0][57] ), .A3(\ram[2][57] ), .A2(\ram[1][57] ), 
        .A4(\ram[3][57] ), .S0(n4242), .S1(n52), .Y(n4565) );
  MUX41X1_HVT U529 ( .A1(n4565), .A3(n4563), .A2(n4564), .A4(n4562), .S0(n4314), .S1(n4291), .Y(q[57]) );
  MUX41X1_HVT U530 ( .A1(\ram[12][58] ), .A3(\ram[14][58] ), .A2(\ram[13][58] ), .A4(\ram[15][58] ), .S0(n4242), .S1(n52), .Y(n4566) );
  MUX41X1_HVT U531 ( .A1(\ram[8][58] ), .A3(\ram[10][58] ), .A2(\ram[9][58] ), 
        .A4(\ram[11][58] ), .S0(n4242), .S1(n52), .Y(n4567) );
  MUX41X1_HVT U532 ( .A1(\ram[4][58] ), .A3(\ram[6][58] ), .A2(\ram[5][58] ), 
        .A4(\ram[7][58] ), .S0(n4242), .S1(n52), .Y(n4568) );
  MUX41X1_HVT U533 ( .A1(\ram[0][58] ), .A3(\ram[2][58] ), .A2(\ram[1][58] ), 
        .A4(\ram[3][58] ), .S0(n4242), .S1(n52), .Y(n4569) );
  MUX41X1_HVT U534 ( .A1(n4569), .A3(n4567), .A2(n4568), .A4(n4566), .S0(n4314), .S1(n4291), .Y(q[58]) );
  MUX41X1_HVT U535 ( .A1(\ram[12][59] ), .A3(\ram[14][59] ), .A2(\ram[13][59] ), .A4(\ram[15][59] ), .S0(n4242), .S1(n52), .Y(n4570) );
  MUX41X1_HVT U536 ( .A1(\ram[8][59] ), .A3(\ram[10][59] ), .A2(\ram[9][59] ), 
        .A4(\ram[11][59] ), .S0(n4242), .S1(n52), .Y(n4571) );
  MUX41X1_HVT U537 ( .A1(\ram[4][59] ), .A3(\ram[6][59] ), .A2(\ram[5][59] ), 
        .A4(\ram[7][59] ), .S0(n4242), .S1(n52), .Y(n4572) );
  MUX41X1_HVT U538 ( .A1(\ram[0][59] ), .A3(\ram[2][59] ), .A2(\ram[1][59] ), 
        .A4(\ram[3][59] ), .S0(n4242), .S1(n52), .Y(n4573) );
  MUX41X1_HVT U539 ( .A1(n4573), .A3(n4571), .A2(n4572), .A4(n4570), .S0(n4314), .S1(n4291), .Y(q[59]) );
  MUX41X1_HVT U540 ( .A1(\ram[12][60] ), .A3(\ram[14][60] ), .A2(\ram[13][60] ), .A4(\ram[15][60] ), .S0(n4243), .S1(n53), .Y(n4574) );
  MUX41X1_HVT U541 ( .A1(\ram[8][60] ), .A3(\ram[10][60] ), .A2(\ram[9][60] ), 
        .A4(\ram[11][60] ), .S0(n4243), .S1(n53), .Y(n4575) );
  MUX41X1_HVT U542 ( .A1(\ram[4][60] ), .A3(\ram[6][60] ), .A2(\ram[5][60] ), 
        .A4(\ram[7][60] ), .S0(n4243), .S1(n53), .Y(n4576) );
  MUX41X1_HVT U543 ( .A1(\ram[0][60] ), .A3(\ram[2][60] ), .A2(\ram[1][60] ), 
        .A4(\ram[3][60] ), .S0(n4243), .S1(n53), .Y(n4577) );
  MUX41X1_HVT U544 ( .A1(n4577), .A3(n4575), .A2(n4576), .A4(n4574), .S0(n4315), .S1(n4292), .Y(q[60]) );
  MUX41X1_HVT U545 ( .A1(\ram[12][61] ), .A3(\ram[14][61] ), .A2(\ram[13][61] ), .A4(\ram[15][61] ), .S0(n4243), .S1(n53), .Y(n4578) );
  MUX41X1_HVT U546 ( .A1(\ram[8][61] ), .A3(\ram[10][61] ), .A2(\ram[9][61] ), 
        .A4(\ram[11][61] ), .S0(n4243), .S1(n53), .Y(n4579) );
  MUX41X1_HVT U547 ( .A1(\ram[4][61] ), .A3(\ram[6][61] ), .A2(\ram[5][61] ), 
        .A4(\ram[7][61] ), .S0(n4243), .S1(n53), .Y(n4580) );
  MUX41X1_HVT U548 ( .A1(\ram[0][61] ), .A3(\ram[2][61] ), .A2(\ram[1][61] ), 
        .A4(\ram[3][61] ), .S0(n4243), .S1(n53), .Y(n4581) );
  MUX41X1_HVT U549 ( .A1(n4581), .A3(n4579), .A2(n4580), .A4(n4578), .S0(n4315), .S1(n4292), .Y(q[61]) );
  MUX41X1_HVT U550 ( .A1(\ram[12][62] ), .A3(\ram[14][62] ), .A2(\ram[13][62] ), .A4(\ram[15][62] ), .S0(n4243), .S1(n53), .Y(n4582) );
  MUX41X1_HVT U551 ( .A1(\ram[8][62] ), .A3(\ram[10][62] ), .A2(\ram[9][62] ), 
        .A4(\ram[11][62] ), .S0(n4243), .S1(n53), .Y(n4583) );
  MUX41X1_HVT U552 ( .A1(\ram[4][62] ), .A3(\ram[6][62] ), .A2(\ram[5][62] ), 
        .A4(\ram[7][62] ), .S0(n4243), .S1(n53), .Y(n4584) );
  MUX41X1_HVT U553 ( .A1(\ram[0][62] ), .A3(\ram[2][62] ), .A2(\ram[1][62] ), 
        .A4(\ram[3][62] ), .S0(n4243), .S1(n53), .Y(n4585) );
  MUX41X1_HVT U554 ( .A1(n4585), .A3(n4583), .A2(n4584), .A4(n4582), .S0(n4315), .S1(n4292), .Y(q[62]) );
  MUX41X1_HVT U555 ( .A1(\ram[12][63] ), .A3(\ram[14][63] ), .A2(\ram[13][63] ), .A4(\ram[15][63] ), .S0(n4244), .S1(n54), .Y(n4586) );
  MUX41X1_HVT U556 ( .A1(\ram[8][63] ), .A3(\ram[10][63] ), .A2(\ram[9][63] ), 
        .A4(\ram[11][63] ), .S0(n4244), .S1(n54), .Y(n4587) );
  MUX41X1_HVT U557 ( .A1(\ram[4][63] ), .A3(\ram[6][63] ), .A2(\ram[5][63] ), 
        .A4(\ram[7][63] ), .S0(n4244), .S1(n54), .Y(n4588) );
  MUX41X1_HVT U558 ( .A1(\ram[0][63] ), .A3(\ram[2][63] ), .A2(\ram[1][63] ), 
        .A4(\ram[3][63] ), .S0(n4244), .S1(n54), .Y(n4589) );
  MUX41X1_HVT U559 ( .A1(n4589), .A3(n4587), .A2(n4588), .A4(n4586), .S0(n4315), .S1(n4292), .Y(q[63]) );
  MUX41X1_HVT U560 ( .A1(\ram[12][64] ), .A3(\ram[14][64] ), .A2(\ram[13][64] ), .A4(\ram[15][64] ), .S0(n4244), .S1(n54), .Y(n4590) );
  MUX41X1_HVT U561 ( .A1(\ram[8][64] ), .A3(\ram[10][64] ), .A2(\ram[9][64] ), 
        .A4(\ram[11][64] ), .S0(n4271), .S1(n4177), .Y(n4591) );
  MUX41X1_HVT U562 ( .A1(\ram[4][64] ), .A3(\ram[6][64] ), .A2(\ram[5][64] ), 
        .A4(\ram[7][64] ), .S0(n4265), .S1(n4171), .Y(n4592) );
  MUX41X1_HVT U563 ( .A1(\ram[0][64] ), .A3(\ram[2][64] ), .A2(\ram[1][64] ), 
        .A4(\ram[3][64] ), .S0(n4265), .S1(n4171), .Y(n4593) );
  MUX41X1_HVT U564 ( .A1(n4593), .A3(n4591), .A2(n4592), .A4(n4590), .S0(n4315), .S1(n4292), .Y(q[64]) );
  MUX41X1_HVT U565 ( .A1(\ram[12][65] ), .A3(\ram[14][65] ), .A2(\ram[13][65] ), .A4(\ram[15][65] ), .S0(n4265), .S1(n4171), .Y(n4594) );
  MUX41X1_HVT U566 ( .A1(\ram[8][65] ), .A3(\ram[10][65] ), .A2(\ram[9][65] ), 
        .A4(\ram[11][65] ), .S0(n4266), .S1(n4172), .Y(n4595) );
  MUX41X1_HVT U567 ( .A1(\ram[4][65] ), .A3(\ram[6][65] ), .A2(\ram[5][65] ), 
        .A4(\ram[7][65] ), .S0(n4266), .S1(n4172), .Y(n4596) );
  MUX41X1_HVT U568 ( .A1(\ram[0][65] ), .A3(\ram[2][65] ), .A2(\ram[1][65] ), 
        .A4(\ram[3][65] ), .S0(n4266), .S1(n4172), .Y(n4597) );
  MUX41X1_HVT U569 ( .A1(n4597), .A3(n4595), .A2(n4596), .A4(n4594), .S0(n4315), .S1(n4292), .Y(q[65]) );
  MUX41X1_HVT U570 ( .A1(\ram[12][66] ), .A3(\ram[14][66] ), .A2(\ram[13][66] ), .A4(\ram[15][66] ), .S0(n4266), .S1(n4172), .Y(n4598) );
  MUX41X1_HVT U571 ( .A1(\ram[8][66] ), .A3(\ram[10][66] ), .A2(\ram[9][66] ), 
        .A4(\ram[11][66] ), .S0(n4266), .S1(n4172), .Y(n4599) );
  MUX41X1_HVT U572 ( .A1(\ram[4][66] ), .A3(\ram[6][66] ), .A2(\ram[5][66] ), 
        .A4(\ram[7][66] ), .S0(n4266), .S1(n4172), .Y(n4600) );
  MUX41X1_HVT U573 ( .A1(\ram[0][66] ), .A3(\ram[2][66] ), .A2(\ram[1][66] ), 
        .A4(\ram[3][66] ), .S0(n4266), .S1(n4172), .Y(n4601) );
  MUX41X1_HVT U574 ( .A1(n4601), .A3(n4599), .A2(n4600), .A4(n4598), .S0(n4315), .S1(n4292), .Y(q[66]) );
  MUX41X1_HVT U575 ( .A1(\ram[12][67] ), .A3(\ram[14][67] ), .A2(\ram[13][67] ), .A4(\ram[15][67] ), .S0(n4266), .S1(n4172), .Y(n4602) );
  MUX41X1_HVT U576 ( .A1(\ram[8][67] ), .A3(\ram[10][67] ), .A2(\ram[9][67] ), 
        .A4(\ram[11][67] ), .S0(n4266), .S1(n4172), .Y(n4603) );
  MUX41X1_HVT U577 ( .A1(\ram[4][67] ), .A3(\ram[6][67] ), .A2(\ram[5][67] ), 
        .A4(\ram[7][67] ), .S0(n4266), .S1(n4172), .Y(n4604) );
  MUX41X1_HVT U578 ( .A1(\ram[0][67] ), .A3(\ram[2][67] ), .A2(\ram[1][67] ), 
        .A4(\ram[3][67] ), .S0(n4266), .S1(n4172), .Y(n4605) );
  MUX41X1_HVT U579 ( .A1(n4605), .A3(n4603), .A2(n4604), .A4(n4602), .S0(n4315), .S1(n4292), .Y(q[67]) );
  MUX41X1_HVT U580 ( .A1(\ram[12][68] ), .A3(\ram[14][68] ), .A2(\ram[13][68] ), .A4(\ram[15][68] ), .S0(n4266), .S1(n4172), .Y(n4606) );
  MUX41X1_HVT U581 ( .A1(\ram[8][68] ), .A3(\ram[10][68] ), .A2(\ram[9][68] ), 
        .A4(\ram[11][68] ), .S0(n4267), .S1(n4173), .Y(n4607) );
  MUX41X1_HVT U582 ( .A1(\ram[4][68] ), .A3(\ram[6][68] ), .A2(\ram[5][68] ), 
        .A4(\ram[7][68] ), .S0(n4267), .S1(n4173), .Y(n4608) );
  MUX41X1_HVT U583 ( .A1(\ram[0][68] ), .A3(\ram[2][68] ), .A2(\ram[1][68] ), 
        .A4(\ram[3][68] ), .S0(n4267), .S1(n4173), .Y(n4609) );
  MUX41X1_HVT U584 ( .A1(n4609), .A3(n4607), .A2(n4608), .A4(n4606), .S0(n4315), .S1(n4292), .Y(q[68]) );
  MUX41X1_HVT U585 ( .A1(\ram[12][69] ), .A3(\ram[14][69] ), .A2(\ram[13][69] ), .A4(\ram[15][69] ), .S0(n4267), .S1(n4173), .Y(n4610) );
  MUX41X1_HVT U586 ( .A1(\ram[8][69] ), .A3(\ram[10][69] ), .A2(\ram[9][69] ), 
        .A4(\ram[11][69] ), .S0(n4267), .S1(n4173), .Y(n4611) );
  MUX41X1_HVT U587 ( .A1(\ram[4][69] ), .A3(\ram[6][69] ), .A2(\ram[5][69] ), 
        .A4(\ram[7][69] ), .S0(n4267), .S1(n4173), .Y(n4612) );
  MUX41X1_HVT U588 ( .A1(\ram[0][69] ), .A3(\ram[2][69] ), .A2(\ram[1][69] ), 
        .A4(\ram[3][69] ), .S0(n4267), .S1(n4173), .Y(n4613) );
  MUX41X1_HVT U589 ( .A1(n4613), .A3(n4611), .A2(n4612), .A4(n4610), .S0(n4315), .S1(n4292), .Y(q[69]) );
  MUX41X1_HVT U590 ( .A1(\ram[12][70] ), .A3(\ram[14][70] ), .A2(\ram[13][70] ), .A4(\ram[15][70] ), .S0(n4267), .S1(n4173), .Y(n4614) );
  MUX41X1_HVT U591 ( .A1(\ram[8][70] ), .A3(\ram[10][70] ), .A2(\ram[9][70] ), 
        .A4(\ram[11][70] ), .S0(n4267), .S1(n4173), .Y(n4615) );
  MUX41X1_HVT U592 ( .A1(\ram[4][70] ), .A3(\ram[6][70] ), .A2(\ram[5][70] ), 
        .A4(\ram[7][70] ), .S0(n4267), .S1(n4173), .Y(n4616) );
  MUX41X1_HVT U593 ( .A1(\ram[0][70] ), .A3(\ram[2][70] ), .A2(\ram[1][70] ), 
        .A4(\ram[3][70] ), .S0(n4267), .S1(n4173), .Y(n4617) );
  MUX41X1_HVT U594 ( .A1(n4617), .A3(n4615), .A2(n4616), .A4(n4614), .S0(n4315), .S1(n4292), .Y(q[70]) );
  MUX41X1_HVT U595 ( .A1(\ram[12][71] ), .A3(\ram[14][71] ), .A2(\ram[13][71] ), .A4(\ram[15][71] ), .S0(n4267), .S1(n4173), .Y(n4618) );
  MUX41X1_HVT U596 ( .A1(\ram[8][71] ), .A3(\ram[10][71] ), .A2(\ram[9][71] ), 
        .A4(\ram[11][71] ), .S0(n4268), .S1(n4174), .Y(n4619) );
  MUX41X1_HVT U597 ( .A1(\ram[4][71] ), .A3(\ram[6][71] ), .A2(\ram[5][71] ), 
        .A4(\ram[7][71] ), .S0(n4268), .S1(n4174), .Y(n4620) );
  MUX41X1_HVT U598 ( .A1(\ram[0][71] ), .A3(\ram[2][71] ), .A2(\ram[1][71] ), 
        .A4(\ram[3][71] ), .S0(n4268), .S1(n4174), .Y(n4621) );
  MUX41X1_HVT U599 ( .A1(n4621), .A3(n4619), .A2(n4620), .A4(n4618), .S0(n4315), .S1(n4292), .Y(q[71]) );
  MUX41X1_HVT U600 ( .A1(\ram[12][72] ), .A3(\ram[14][72] ), .A2(\ram[13][72] ), .A4(\ram[15][72] ), .S0(n4268), .S1(n4174), .Y(n4622) );
  MUX41X1_HVT U601 ( .A1(\ram[8][72] ), .A3(\ram[10][72] ), .A2(\ram[9][72] ), 
        .A4(\ram[11][72] ), .S0(n4268), .S1(n4174), .Y(n4623) );
  MUX41X1_HVT U602 ( .A1(\ram[4][72] ), .A3(\ram[6][72] ), .A2(\ram[5][72] ), 
        .A4(\ram[7][72] ), .S0(n4268), .S1(n4174), .Y(n4624) );
  MUX41X1_HVT U603 ( .A1(\ram[0][72] ), .A3(\ram[2][72] ), .A2(\ram[1][72] ), 
        .A4(\ram[3][72] ), .S0(n4268), .S1(n4174), .Y(n4625) );
  MUX41X1_HVT U604 ( .A1(n4625), .A3(n4623), .A2(n4624), .A4(n4622), .S0(n4316), .S1(n4293), .Y(q[72]) );
  MUX41X1_HVT U605 ( .A1(\ram[12][73] ), .A3(\ram[14][73] ), .A2(\ram[13][73] ), .A4(\ram[15][73] ), .S0(n4268), .S1(n4174), .Y(n4626) );
  MUX41X1_HVT U606 ( .A1(\ram[8][73] ), .A3(\ram[10][73] ), .A2(\ram[9][73] ), 
        .A4(\ram[11][73] ), .S0(n4268), .S1(n4174), .Y(n4627) );
  MUX41X1_HVT U607 ( .A1(\ram[4][73] ), .A3(\ram[6][73] ), .A2(\ram[5][73] ), 
        .A4(\ram[7][73] ), .S0(n4268), .S1(n4174), .Y(n4628) );
  MUX41X1_HVT U608 ( .A1(\ram[0][73] ), .A3(\ram[2][73] ), .A2(\ram[1][73] ), 
        .A4(\ram[3][73] ), .S0(n4268), .S1(n4174), .Y(n4629) );
  MUX41X1_HVT U609 ( .A1(n4629), .A3(n4627), .A2(n4628), .A4(n4626), .S0(n4316), .S1(n4293), .Y(q[73]) );
  MUX41X1_HVT U610 ( .A1(\ram[12][74] ), .A3(\ram[14][74] ), .A2(\ram[13][74] ), .A4(\ram[15][74] ), .S0(n4268), .S1(n4174), .Y(n4630) );
  MUX41X1_HVT U611 ( .A1(\ram[8][74] ), .A3(\ram[10][74] ), .A2(\ram[9][74] ), 
        .A4(\ram[11][74] ), .S0(n4269), .S1(n4175), .Y(n4631) );
  MUX41X1_HVT U612 ( .A1(\ram[4][74] ), .A3(\ram[6][74] ), .A2(\ram[5][74] ), 
        .A4(\ram[7][74] ), .S0(n4269), .S1(n4175), .Y(n4632) );
  MUX41X1_HVT U613 ( .A1(\ram[0][74] ), .A3(\ram[2][74] ), .A2(\ram[1][74] ), 
        .A4(\ram[3][74] ), .S0(n4269), .S1(n4175), .Y(n4633) );
  MUX41X1_HVT U614 ( .A1(n4633), .A3(n4631), .A2(n4632), .A4(n4630), .S0(n4316), .S1(n4293), .Y(q[74]) );
  MUX41X1_HVT U615 ( .A1(\ram[12][75] ), .A3(\ram[14][75] ), .A2(\ram[13][75] ), .A4(\ram[15][75] ), .S0(n4269), .S1(n4175), .Y(n4634) );
  MUX41X1_HVT U616 ( .A1(\ram[8][75] ), .A3(\ram[10][75] ), .A2(\ram[9][75] ), 
        .A4(\ram[11][75] ), .S0(n4269), .S1(n4175), .Y(n4635) );
  MUX41X1_HVT U617 ( .A1(\ram[4][75] ), .A3(\ram[6][75] ), .A2(\ram[5][75] ), 
        .A4(\ram[7][75] ), .S0(n4269), .S1(n4175), .Y(n4636) );
  MUX41X1_HVT U618 ( .A1(\ram[0][75] ), .A3(\ram[2][75] ), .A2(\ram[1][75] ), 
        .A4(\ram[3][75] ), .S0(n4269), .S1(n4175), .Y(n4637) );
  MUX41X1_HVT U619 ( .A1(n4637), .A3(n4635), .A2(n4636), .A4(n4634), .S0(n4316), .S1(n4293), .Y(q[75]) );
  MUX41X1_HVT U620 ( .A1(\ram[12][76] ), .A3(\ram[14][76] ), .A2(\ram[13][76] ), .A4(\ram[15][76] ), .S0(n4269), .S1(n4175), .Y(n4638) );
  MUX41X1_HVT U621 ( .A1(\ram[8][76] ), .A3(\ram[10][76] ), .A2(\ram[9][76] ), 
        .A4(\ram[11][76] ), .S0(n4269), .S1(n4175), .Y(n4639) );
  MUX41X1_HVT U622 ( .A1(\ram[4][76] ), .A3(\ram[6][76] ), .A2(\ram[5][76] ), 
        .A4(\ram[7][76] ), .S0(n4269), .S1(n4175), .Y(n4640) );
  MUX41X1_HVT U623 ( .A1(\ram[0][76] ), .A3(\ram[2][76] ), .A2(\ram[1][76] ), 
        .A4(\ram[3][76] ), .S0(n4269), .S1(n4175), .Y(n4641) );
  MUX41X1_HVT U624 ( .A1(n4641), .A3(n4639), .A2(n4640), .A4(n4638), .S0(n4316), .S1(n4293), .Y(q[76]) );
  MUX41X1_HVT U625 ( .A1(\ram[12][77] ), .A3(\ram[14][77] ), .A2(\ram[13][77] ), .A4(\ram[15][77] ), .S0(n4269), .S1(n4175), .Y(n4642) );
  MUX41X1_HVT U626 ( .A1(\ram[8][77] ), .A3(\ram[10][77] ), .A2(\ram[9][77] ), 
        .A4(\ram[11][77] ), .S0(n4270), .S1(n4176), .Y(n4643) );
  MUX41X1_HVT U627 ( .A1(\ram[4][77] ), .A3(\ram[6][77] ), .A2(\ram[5][77] ), 
        .A4(\ram[7][77] ), .S0(n4270), .S1(n4176), .Y(n4644) );
  MUX41X1_HVT U628 ( .A1(\ram[0][77] ), .A3(\ram[2][77] ), .A2(\ram[1][77] ), 
        .A4(\ram[3][77] ), .S0(n4270), .S1(n4176), .Y(n4645) );
  MUX41X1_HVT U629 ( .A1(n4645), .A3(n4643), .A2(n4644), .A4(n4642), .S0(n4316), .S1(n4293), .Y(q[77]) );
  MUX41X1_HVT U630 ( .A1(\ram[12][78] ), .A3(\ram[14][78] ), .A2(\ram[13][78] ), .A4(\ram[15][78] ), .S0(n4270), .S1(n4176), .Y(n4646) );
  MUX41X1_HVT U631 ( .A1(\ram[8][78] ), .A3(\ram[10][78] ), .A2(\ram[9][78] ), 
        .A4(\ram[11][78] ), .S0(n4270), .S1(n4176), .Y(n4647) );
  MUX41X1_HVT U632 ( .A1(\ram[4][78] ), .A3(\ram[6][78] ), .A2(\ram[5][78] ), 
        .A4(\ram[7][78] ), .S0(n4270), .S1(n4176), .Y(n4648) );
  MUX41X1_HVT U633 ( .A1(\ram[0][78] ), .A3(\ram[2][78] ), .A2(\ram[1][78] ), 
        .A4(\ram[3][78] ), .S0(n4270), .S1(n4176), .Y(n4649) );
  MUX41X1_HVT U634 ( .A1(n4649), .A3(n4647), .A2(n4648), .A4(n4646), .S0(n4316), .S1(n4293), .Y(q[78]) );
  MUX41X1_HVT U635 ( .A1(\ram[12][79] ), .A3(\ram[14][79] ), .A2(\ram[13][79] ), .A4(\ram[15][79] ), .S0(n4270), .S1(n4176), .Y(n4650) );
  MUX41X1_HVT U636 ( .A1(\ram[8][79] ), .A3(\ram[10][79] ), .A2(\ram[9][79] ), 
        .A4(\ram[11][79] ), .S0(n4270), .S1(n4176), .Y(n4651) );
  MUX41X1_HVT U637 ( .A1(\ram[4][79] ), .A3(\ram[6][79] ), .A2(\ram[5][79] ), 
        .A4(\ram[7][79] ), .S0(n4270), .S1(n4176), .Y(n4652) );
  MUX41X1_HVT U638 ( .A1(\ram[0][79] ), .A3(\ram[2][79] ), .A2(\ram[1][79] ), 
        .A4(\ram[3][79] ), .S0(n4270), .S1(n4176), .Y(n4653) );
  MUX41X1_HVT U639 ( .A1(n4653), .A3(n4651), .A2(n4652), .A4(n4650), .S0(n4316), .S1(n4293), .Y(q[79]) );
  MUX41X1_HVT U640 ( .A1(\ram[12][80] ), .A3(\ram[14][80] ), .A2(\ram[13][80] ), .A4(\ram[15][80] ), .S0(n4270), .S1(n4176), .Y(n4654) );
  MUX41X1_HVT U641 ( .A1(\ram[8][80] ), .A3(\ram[10][80] ), .A2(\ram[9][80] ), 
        .A4(\ram[11][80] ), .S0(n4271), .S1(n4177), .Y(n4655) );
  MUX41X1_HVT U642 ( .A1(\ram[4][80] ), .A3(\ram[6][80] ), .A2(\ram[5][80] ), 
        .A4(\ram[7][80] ), .S0(n4271), .S1(n4177), .Y(n4656) );
  MUX41X1_HVT U643 ( .A1(\ram[0][80] ), .A3(\ram[2][80] ), .A2(\ram[1][80] ), 
        .A4(\ram[3][80] ), .S0(n4271), .S1(n4177), .Y(n4657) );
  MUX41X1_HVT U644 ( .A1(n4657), .A3(n4655), .A2(n4656), .A4(n4654), .S0(n4316), .S1(n4293), .Y(q[80]) );
  MUX41X1_HVT U645 ( .A1(\ram[12][81] ), .A3(\ram[14][81] ), .A2(\ram[13][81] ), .A4(\ram[15][81] ), .S0(n4271), .S1(n4177), .Y(n4658) );
  MUX41X1_HVT U646 ( .A1(\ram[8][81] ), .A3(\ram[10][81] ), .A2(\ram[9][81] ), 
        .A4(\ram[11][81] ), .S0(n4271), .S1(n4177), .Y(n4659) );
  MUX41X1_HVT U647 ( .A1(\ram[4][81] ), .A3(\ram[6][81] ), .A2(\ram[5][81] ), 
        .A4(\ram[7][81] ), .S0(n4271), .S1(n4177), .Y(n4660) );
  MUX41X1_HVT U648 ( .A1(\ram[0][81] ), .A3(\ram[2][81] ), .A2(\ram[1][81] ), 
        .A4(\ram[3][81] ), .S0(n4271), .S1(n4177), .Y(n4661) );
  MUX41X1_HVT U649 ( .A1(n4661), .A3(n4659), .A2(n4660), .A4(n4658), .S0(n4316), .S1(n4293), .Y(q[81]) );
  MUX41X1_HVT U650 ( .A1(\ram[12][82] ), .A3(\ram[14][82] ), .A2(\ram[13][82] ), .A4(\ram[15][82] ), .S0(n4271), .S1(n4177), .Y(n4662) );
  MUX41X1_HVT U651 ( .A1(\ram[8][82] ), .A3(\ram[10][82] ), .A2(\ram[9][82] ), 
        .A4(\ram[11][82] ), .S0(n4271), .S1(n4177), .Y(n4663) );
  MUX41X1_HVT U652 ( .A1(\ram[4][82] ), .A3(\ram[6][82] ), .A2(\ram[5][82] ), 
        .A4(\ram[7][82] ), .S0(n4271), .S1(n4177), .Y(n4664) );
  MUX41X1_HVT U653 ( .A1(\ram[0][82] ), .A3(\ram[2][82] ), .A2(\ram[1][82] ), 
        .A4(\ram[3][82] ), .S0(n4271), .S1(n4177), .Y(n4665) );
  MUX41X1_HVT U654 ( .A1(n4665), .A3(n4663), .A2(n4664), .A4(n4662), .S0(n4316), .S1(n4293), .Y(q[82]) );
  MUX41X1_HVT U655 ( .A1(\ram[12][83] ), .A3(\ram[14][83] ), .A2(\ram[13][83] ), .A4(\ram[15][83] ), .S0(n4272), .S1(n4178), .Y(n4666) );
  MUX41X1_HVT U656 ( .A1(\ram[8][83] ), .A3(\ram[10][83] ), .A2(\ram[9][83] ), 
        .A4(\ram[11][83] ), .S0(n4272), .S1(n4178), .Y(n4667) );
  MUX41X1_HVT U657 ( .A1(\ram[4][83] ), .A3(\ram[6][83] ), .A2(\ram[5][83] ), 
        .A4(\ram[7][83] ), .S0(n4272), .S1(n4178), .Y(n4668) );
  MUX41X1_HVT U658 ( .A1(\ram[0][83] ), .A3(\ram[2][83] ), .A2(\ram[1][83] ), 
        .A4(\ram[3][83] ), .S0(n4272), .S1(n4178), .Y(n4669) );
  MUX41X1_HVT U659 ( .A1(n4669), .A3(n4667), .A2(n4668), .A4(n4666), .S0(n4316), .S1(n4293), .Y(q[83]) );
  MUX41X1_HVT U660 ( .A1(\ram[12][84] ), .A3(\ram[14][84] ), .A2(\ram[13][84] ), .A4(\ram[15][84] ), .S0(n4272), .S1(n4178), .Y(n4670) );
  MUX41X1_HVT U661 ( .A1(\ram[8][84] ), .A3(\ram[10][84] ), .A2(\ram[9][84] ), 
        .A4(\ram[11][84] ), .S0(n4272), .S1(n4178), .Y(n4671) );
  MUX41X1_HVT U662 ( .A1(\ram[4][84] ), .A3(\ram[6][84] ), .A2(\ram[5][84] ), 
        .A4(\ram[7][84] ), .S0(n4272), .S1(n4178), .Y(n4672) );
  MUX41X1_HVT U663 ( .A1(\ram[0][84] ), .A3(\ram[2][84] ), .A2(\ram[1][84] ), 
        .A4(\ram[3][84] ), .S0(n4272), .S1(n4178), .Y(n4673) );
  MUX41X1_HVT U664 ( .A1(n4673), .A3(n4671), .A2(n4672), .A4(n4670), .S0(n4317), .S1(n4294), .Y(q[84]) );
  MUX41X1_HVT U665 ( .A1(\ram[12][85] ), .A3(\ram[14][85] ), .A2(\ram[13][85] ), .A4(\ram[15][85] ), .S0(n4272), .S1(n4178), .Y(n4674) );
  MUX41X1_HVT U666 ( .A1(\ram[8][85] ), .A3(\ram[10][85] ), .A2(\ram[9][85] ), 
        .A4(\ram[11][85] ), .S0(n4272), .S1(n4178), .Y(n4675) );
  MUX41X1_HVT U667 ( .A1(\ram[4][85] ), .A3(\ram[6][85] ), .A2(\ram[5][85] ), 
        .A4(\ram[7][85] ), .S0(n4272), .S1(n4178), .Y(n4676) );
  MUX41X1_HVT U668 ( .A1(\ram[0][85] ), .A3(\ram[2][85] ), .A2(\ram[1][85] ), 
        .A4(\ram[3][85] ), .S0(n4272), .S1(n4178), .Y(n4677) );
  MUX41X1_HVT U669 ( .A1(n4677), .A3(n4675), .A2(n4676), .A4(n4674), .S0(n4317), .S1(n4294), .Y(q[85]) );
  MUX41X1_HVT U670 ( .A1(\ram[12][86] ), .A3(\ram[14][86] ), .A2(\ram[13][86] ), .A4(\ram[15][86] ), .S0(n4273), .S1(n4179), .Y(n4678) );
  MUX41X1_HVT U671 ( .A1(\ram[8][86] ), .A3(\ram[10][86] ), .A2(\ram[9][86] ), 
        .A4(\ram[11][86] ), .S0(n4273), .S1(n4179), .Y(n4679) );
  MUX41X1_HVT U672 ( .A1(\ram[4][86] ), .A3(\ram[6][86] ), .A2(\ram[5][86] ), 
        .A4(\ram[7][86] ), .S0(n4273), .S1(n4179), .Y(n4680) );
  MUX41X1_HVT U673 ( .A1(\ram[0][86] ), .A3(\ram[2][86] ), .A2(\ram[1][86] ), 
        .A4(\ram[3][86] ), .S0(n4273), .S1(n4179), .Y(n4681) );
  MUX41X1_HVT U674 ( .A1(n4681), .A3(n4679), .A2(n4680), .A4(n4678), .S0(n4317), .S1(n4294), .Y(q[86]) );
  MUX41X1_HVT U675 ( .A1(\ram[12][87] ), .A3(\ram[14][87] ), .A2(\ram[13][87] ), .A4(\ram[15][87] ), .S0(n4273), .S1(n4179), .Y(n4682) );
  MUX41X1_HVT U676 ( .A1(\ram[8][87] ), .A3(\ram[10][87] ), .A2(\ram[9][87] ), 
        .A4(\ram[11][87] ), .S0(n4273), .S1(n4179), .Y(n4683) );
  MUX41X1_HVT U677 ( .A1(\ram[4][87] ), .A3(\ram[6][87] ), .A2(\ram[5][87] ), 
        .A4(\ram[7][87] ), .S0(n4273), .S1(n4179), .Y(n4684) );
  MUX41X1_HVT U678 ( .A1(\ram[0][87] ), .A3(\ram[2][87] ), .A2(\ram[1][87] ), 
        .A4(\ram[3][87] ), .S0(n4273), .S1(n4179), .Y(n4685) );
  MUX41X1_HVT U679 ( .A1(n4685), .A3(n4683), .A2(n4684), .A4(n4682), .S0(n4317), .S1(n4294), .Y(q[87]) );
  MUX41X1_HVT U680 ( .A1(\ram[12][88] ), .A3(\ram[14][88] ), .A2(\ram[13][88] ), .A4(\ram[15][88] ), .S0(n4273), .S1(n4179), .Y(n4686) );
  MUX41X1_HVT U681 ( .A1(\ram[8][88] ), .A3(\ram[10][88] ), .A2(\ram[9][88] ), 
        .A4(\ram[11][88] ), .S0(n4273), .S1(n4179), .Y(n4687) );
  MUX41X1_HVT U682 ( .A1(\ram[4][88] ), .A3(\ram[6][88] ), .A2(\ram[5][88] ), 
        .A4(\ram[7][88] ), .S0(n4273), .S1(n4179), .Y(n4688) );
  MUX41X1_HVT U683 ( .A1(\ram[0][88] ), .A3(\ram[2][88] ), .A2(\ram[1][88] ), 
        .A4(\ram[3][88] ), .S0(n4273), .S1(n4179), .Y(n4689) );
  MUX41X1_HVT U684 ( .A1(n4689), .A3(n4687), .A2(n4688), .A4(n4686), .S0(n4317), .S1(n4294), .Y(q[88]) );
  MUX41X1_HVT U685 ( .A1(\ram[12][89] ), .A3(\ram[14][89] ), .A2(\ram[13][89] ), .A4(\ram[15][89] ), .S0(n4274), .S1(n4180), .Y(n4690) );
  MUX41X1_HVT U686 ( .A1(\ram[8][89] ), .A3(\ram[10][89] ), .A2(\ram[9][89] ), 
        .A4(\ram[11][89] ), .S0(n4274), .S1(n4180), .Y(n4691) );
  MUX41X1_HVT U687 ( .A1(\ram[4][89] ), .A3(\ram[6][89] ), .A2(\ram[5][89] ), 
        .A4(\ram[7][89] ), .S0(n4274), .S1(n4180), .Y(n4692) );
  MUX41X1_HVT U688 ( .A1(\ram[0][89] ), .A3(\ram[2][89] ), .A2(\ram[1][89] ), 
        .A4(\ram[3][89] ), .S0(n4274), .S1(n4180), .Y(n4693) );
  MUX41X1_HVT U689 ( .A1(n4693), .A3(n4691), .A2(n4692), .A4(n4690), .S0(n4317), .S1(n4294), .Y(q[89]) );
  MUX41X1_HVT U690 ( .A1(\ram[12][90] ), .A3(\ram[14][90] ), .A2(\ram[13][90] ), .A4(\ram[15][90] ), .S0(n4274), .S1(n4180), .Y(n4694) );
  MUX41X1_HVT U691 ( .A1(\ram[8][90] ), .A3(\ram[10][90] ), .A2(\ram[9][90] ), 
        .A4(\ram[11][90] ), .S0(n4274), .S1(n4180), .Y(n4695) );
  MUX41X1_HVT U692 ( .A1(\ram[4][90] ), .A3(\ram[6][90] ), .A2(\ram[5][90] ), 
        .A4(\ram[7][90] ), .S0(n4274), .S1(n4180), .Y(n4696) );
  MUX41X1_HVT U693 ( .A1(\ram[0][90] ), .A3(\ram[2][90] ), .A2(\ram[1][90] ), 
        .A4(\ram[3][90] ), .S0(n4274), .S1(n4180), .Y(n4697) );
  MUX41X1_HVT U694 ( .A1(n4697), .A3(n4695), .A2(n4696), .A4(n4694), .S0(n4317), .S1(n4294), .Y(q[90]) );
  MUX41X1_HVT U695 ( .A1(\ram[12][91] ), .A3(\ram[14][91] ), .A2(\ram[13][91] ), .A4(\ram[15][91] ), .S0(n4274), .S1(n4180), .Y(n4698) );
  MUX41X1_HVT U696 ( .A1(\ram[8][91] ), .A3(\ram[10][91] ), .A2(\ram[9][91] ), 
        .A4(\ram[11][91] ), .S0(n4274), .S1(n4180), .Y(n4699) );
  MUX41X1_HVT U697 ( .A1(\ram[4][91] ), .A3(\ram[6][91] ), .A2(\ram[5][91] ), 
        .A4(\ram[7][91] ), .S0(n4274), .S1(n4180), .Y(n4700) );
  MUX41X1_HVT U698 ( .A1(\ram[0][91] ), .A3(\ram[2][91] ), .A2(\ram[1][91] ), 
        .A4(\ram[3][91] ), .S0(n4274), .S1(n4180), .Y(n4701) );
  MUX41X1_HVT U699 ( .A1(n4701), .A3(n4699), .A2(n4700), .A4(n4698), .S0(n4317), .S1(n4294), .Y(q[91]) );
  MUX41X1_HVT U700 ( .A1(\ram[12][92] ), .A3(\ram[14][92] ), .A2(\ram[13][92] ), .A4(\ram[15][92] ), .S0(n4275), .S1(n4181), .Y(n4702) );
  MUX41X1_HVT U701 ( .A1(\ram[8][92] ), .A3(\ram[10][92] ), .A2(\ram[9][92] ), 
        .A4(\ram[11][92] ), .S0(n4275), .S1(n4181), .Y(n4703) );
  MUX41X1_HVT U702 ( .A1(\ram[4][92] ), .A3(\ram[6][92] ), .A2(\ram[5][92] ), 
        .A4(\ram[7][92] ), .S0(n4275), .S1(n4181), .Y(n4704) );
  MUX41X1_HVT U703 ( .A1(\ram[0][92] ), .A3(\ram[2][92] ), .A2(\ram[1][92] ), 
        .A4(\ram[3][92] ), .S0(n4275), .S1(n4181), .Y(n4705) );
  MUX41X1_HVT U704 ( .A1(n4705), .A3(n4703), .A2(n4704), .A4(n4702), .S0(n4317), .S1(n4294), .Y(q[92]) );
  MUX41X1_HVT U705 ( .A1(\ram[12][93] ), .A3(\ram[14][93] ), .A2(\ram[13][93] ), .A4(\ram[15][93] ), .S0(n4275), .S1(n4181), .Y(n4706) );
  MUX41X1_HVT U706 ( .A1(\ram[8][93] ), .A3(\ram[10][93] ), .A2(\ram[9][93] ), 
        .A4(\ram[11][93] ), .S0(n4275), .S1(n4181), .Y(n4707) );
  MUX41X1_HVT U707 ( .A1(\ram[4][93] ), .A3(\ram[6][93] ), .A2(\ram[5][93] ), 
        .A4(\ram[7][93] ), .S0(n4275), .S1(n4181), .Y(n4708) );
  MUX41X1_HVT U708 ( .A1(\ram[0][93] ), .A3(\ram[2][93] ), .A2(\ram[1][93] ), 
        .A4(\ram[3][93] ), .S0(n4275), .S1(n4181), .Y(n4709) );
  MUX41X1_HVT U709 ( .A1(n4709), .A3(n4707), .A2(n4708), .A4(n4706), .S0(n4317), .S1(n4294), .Y(q[93]) );
  MUX41X1_HVT U710 ( .A1(\ram[12][94] ), .A3(\ram[14][94] ), .A2(\ram[13][94] ), .A4(\ram[15][94] ), .S0(n4275), .S1(n4181), .Y(n4710) );
  MUX41X1_HVT U711 ( .A1(\ram[8][94] ), .A3(\ram[10][94] ), .A2(\ram[9][94] ), 
        .A4(\ram[11][94] ), .S0(n4275), .S1(n4181), .Y(n4711) );
  MUX41X1_HVT U712 ( .A1(\ram[4][94] ), .A3(\ram[6][94] ), .A2(\ram[5][94] ), 
        .A4(\ram[7][94] ), .S0(n4275), .S1(n4181), .Y(n4712) );
  MUX41X1_HVT U713 ( .A1(\ram[0][94] ), .A3(\ram[2][94] ), .A2(\ram[1][94] ), 
        .A4(\ram[3][94] ), .S0(n4275), .S1(n4181), .Y(n4713) );
  MUX41X1_HVT U714 ( .A1(n4713), .A3(n4711), .A2(n4712), .A4(n4710), .S0(n4317), .S1(n4294), .Y(q[94]) );
  MUX41X1_HVT U715 ( .A1(\ram[12][95] ), .A3(\ram[14][95] ), .A2(\ram[13][95] ), .A4(\ram[15][95] ), .S0(n4276), .S1(n4182), .Y(n4714) );
  MUX41X1_HVT U716 ( .A1(\ram[8][95] ), .A3(\ram[10][95] ), .A2(\ram[9][95] ), 
        .A4(\ram[11][95] ), .S0(n4276), .S1(n4182), .Y(n4715) );
  MUX41X1_HVT U717 ( .A1(\ram[4][95] ), .A3(\ram[6][95] ), .A2(\ram[5][95] ), 
        .A4(\ram[7][95] ), .S0(n4276), .S1(n4182), .Y(n4716) );
  MUX41X1_HVT U718 ( .A1(\ram[0][95] ), .A3(\ram[2][95] ), .A2(\ram[1][95] ), 
        .A4(\ram[3][95] ), .S0(n4276), .S1(n4182), .Y(n4717) );
  MUX41X1_HVT U719 ( .A1(n4717), .A3(n4715), .A2(n4716), .A4(n4714), .S0(n4317), .S1(n4294), .Y(q[95]) );
  MUX41X1_HVT U720 ( .A1(\ram[12][96] ), .A3(\ram[14][96] ), .A2(\ram[13][96] ), .A4(\ram[15][96] ), .S0(n4260), .S1(n4166), .Y(n4718) );
  MUX41X1_HVT U721 ( .A1(\ram[8][96] ), .A3(\ram[10][96] ), .A2(\ram[9][96] ), 
        .A4(\ram[11][96] ), .S0(n4255), .S1(n4161), .Y(n4719) );
  MUX41X1_HVT U722 ( .A1(\ram[4][96] ), .A3(\ram[6][96] ), .A2(\ram[5][96] ), 
        .A4(\ram[7][96] ), .S0(n4255), .S1(n4161), .Y(n4720) );
  MUX41X1_HVT U723 ( .A1(\ram[0][96] ), .A3(\ram[2][96] ), .A2(\ram[1][96] ), 
        .A4(\ram[3][96] ), .S0(n4255), .S1(n4161), .Y(n4721) );
  MUX41X1_HVT U724 ( .A1(n4721), .A3(n4719), .A2(n4720), .A4(n4718), .S0(n4318), .S1(n4295), .Y(q[96]) );
  MUX41X1_HVT U725 ( .A1(\ram[12][97] ), .A3(\ram[14][97] ), .A2(\ram[13][97] ), .A4(\ram[15][97] ), .S0(n4255), .S1(n4161), .Y(n4722) );
  MUX41X1_HVT U726 ( .A1(\ram[8][97] ), .A3(\ram[10][97] ), .A2(\ram[9][97] ), 
        .A4(\ram[11][97] ), .S0(n4255), .S1(n4161), .Y(n4723) );
  MUX41X1_HVT U727 ( .A1(\ram[4][97] ), .A3(\ram[6][97] ), .A2(\ram[5][97] ), 
        .A4(\ram[7][97] ), .S0(n4255), .S1(n4161), .Y(n4724) );
  MUX41X1_HVT U728 ( .A1(\ram[0][97] ), .A3(\ram[2][97] ), .A2(\ram[1][97] ), 
        .A4(\ram[3][97] ), .S0(n4255), .S1(n4161), .Y(n4725) );
  MUX41X1_HVT U729 ( .A1(n4725), .A3(n4723), .A2(n4724), .A4(n4722), .S0(n4318), .S1(n4295), .Y(q[97]) );
  MUX41X1_HVT U730 ( .A1(\ram[12][98] ), .A3(\ram[14][98] ), .A2(\ram[13][98] ), .A4(\ram[15][98] ), .S0(n4255), .S1(n4161), .Y(n4726) );
  MUX41X1_HVT U731 ( .A1(\ram[8][98] ), .A3(\ram[10][98] ), .A2(\ram[9][98] ), 
        .A4(\ram[11][98] ), .S0(n4255), .S1(n4161), .Y(n4727) );
  MUX41X1_HVT U732 ( .A1(\ram[4][98] ), .A3(\ram[6][98] ), .A2(\ram[5][98] ), 
        .A4(\ram[7][98] ), .S0(n4255), .S1(n4161), .Y(n4728) );
  MUX41X1_HVT U733 ( .A1(\ram[0][98] ), .A3(\ram[2][98] ), .A2(\ram[1][98] ), 
        .A4(\ram[3][98] ), .S0(n4255), .S1(n4161), .Y(n4729) );
  MUX41X1_HVT U734 ( .A1(n4729), .A3(n4727), .A2(n4728), .A4(n4726), .S0(n4318), .S1(n4295), .Y(q[98]) );
  MUX41X1_HVT U735 ( .A1(\ram[12][99] ), .A3(\ram[14][99] ), .A2(\ram[13][99] ), .A4(\ram[15][99] ), .S0(n4256), .S1(n4162), .Y(n4730) );
  MUX41X1_HVT U736 ( .A1(\ram[8][99] ), .A3(\ram[10][99] ), .A2(\ram[9][99] ), 
        .A4(\ram[11][99] ), .S0(n4256), .S1(n4162), .Y(n4731) );
  MUX41X1_HVT U737 ( .A1(\ram[4][99] ), .A3(\ram[6][99] ), .A2(\ram[5][99] ), 
        .A4(\ram[7][99] ), .S0(n4256), .S1(n4162), .Y(n4732) );
  MUX41X1_HVT U738 ( .A1(\ram[0][99] ), .A3(\ram[2][99] ), .A2(\ram[1][99] ), 
        .A4(\ram[3][99] ), .S0(n4256), .S1(n4162), .Y(n4733) );
  MUX41X1_HVT U739 ( .A1(n4733), .A3(n4731), .A2(n4732), .A4(n4730), .S0(n4318), .S1(n4295), .Y(q[99]) );
  MUX41X1_HVT U740 ( .A1(\ram[12][100] ), .A3(\ram[14][100] ), .A2(
        \ram[13][100] ), .A4(\ram[15][100] ), .S0(n4256), .S1(n4162), .Y(n4734) );
  MUX41X1_HVT U741 ( .A1(\ram[8][100] ), .A3(\ram[10][100] ), .A2(
        \ram[9][100] ), .A4(\ram[11][100] ), .S0(n4256), .S1(n4162), .Y(n4735)
         );
  MUX41X1_HVT U742 ( .A1(\ram[4][100] ), .A3(\ram[6][100] ), .A2(\ram[5][100] ), .A4(\ram[7][100] ), .S0(n4256), .S1(n4162), .Y(n4736) );
  MUX41X1_HVT U743 ( .A1(\ram[0][100] ), .A3(\ram[2][100] ), .A2(\ram[1][100] ), .A4(\ram[3][100] ), .S0(n4256), .S1(n4162), .Y(n4737) );
  MUX41X1_HVT U744 ( .A1(n4737), .A3(n4735), .A2(n4736), .A4(n4734), .S0(n4318), .S1(n4295), .Y(q[100]) );
  MUX41X1_HVT U745 ( .A1(\ram[12][101] ), .A3(\ram[14][101] ), .A2(
        \ram[13][101] ), .A4(\ram[15][101] ), .S0(n4256), .S1(n4162), .Y(n4738) );
  MUX41X1_HVT U746 ( .A1(\ram[8][101] ), .A3(\ram[10][101] ), .A2(
        \ram[9][101] ), .A4(\ram[11][101] ), .S0(n4256), .S1(n4162), .Y(n4739)
         );
  MUX41X1_HVT U747 ( .A1(\ram[4][101] ), .A3(\ram[6][101] ), .A2(\ram[5][101] ), .A4(\ram[7][101] ), .S0(n4256), .S1(n4162), .Y(n4740) );
  MUX41X1_HVT U748 ( .A1(\ram[0][101] ), .A3(\ram[2][101] ), .A2(\ram[1][101] ), .A4(\ram[3][101] ), .S0(n4256), .S1(n4162), .Y(n4741) );
  MUX41X1_HVT U749 ( .A1(n4741), .A3(n4739), .A2(n4740), .A4(n4738), .S0(n4318), .S1(n4295), .Y(q[101]) );
  MUX41X1_HVT U750 ( .A1(\ram[12][102] ), .A3(\ram[14][102] ), .A2(
        \ram[13][102] ), .A4(\ram[15][102] ), .S0(n4257), .S1(n4163), .Y(n4742) );
  MUX41X1_HVT U751 ( .A1(\ram[8][102] ), .A3(\ram[10][102] ), .A2(
        \ram[9][102] ), .A4(\ram[11][102] ), .S0(n4257), .S1(n4163), .Y(n4743)
         );
  MUX41X1_HVT U752 ( .A1(\ram[4][102] ), .A3(\ram[6][102] ), .A2(\ram[5][102] ), .A4(\ram[7][102] ), .S0(n4257), .S1(n4163), .Y(n4744) );
  MUX41X1_HVT U753 ( .A1(\ram[0][102] ), .A3(\ram[2][102] ), .A2(\ram[1][102] ), .A4(\ram[3][102] ), .S0(n4257), .S1(n4163), .Y(n4745) );
  MUX41X1_HVT U754 ( .A1(n4745), .A3(n4743), .A2(n4744), .A4(n4742), .S0(n4318), .S1(n4295), .Y(q[102]) );
  MUX41X1_HVT U755 ( .A1(\ram[12][103] ), .A3(\ram[14][103] ), .A2(
        \ram[13][103] ), .A4(\ram[15][103] ), .S0(n4257), .S1(n4163), .Y(n4746) );
  MUX41X1_HVT U756 ( .A1(\ram[8][103] ), .A3(\ram[10][103] ), .A2(
        \ram[9][103] ), .A4(\ram[11][103] ), .S0(n4257), .S1(n4163), .Y(n4747)
         );
  MUX41X1_HVT U757 ( .A1(\ram[4][103] ), .A3(\ram[6][103] ), .A2(\ram[5][103] ), .A4(\ram[7][103] ), .S0(n4257), .S1(n4163), .Y(n4748) );
  MUX41X1_HVT U758 ( .A1(\ram[0][103] ), .A3(\ram[2][103] ), .A2(\ram[1][103] ), .A4(\ram[3][103] ), .S0(n4257), .S1(n4163), .Y(n4749) );
  MUX41X1_HVT U759 ( .A1(n4749), .A3(n4747), .A2(n4748), .A4(n4746), .S0(n4318), .S1(n4295), .Y(q[103]) );
  MUX41X1_HVT U760 ( .A1(\ram[12][104] ), .A3(\ram[14][104] ), .A2(
        \ram[13][104] ), .A4(\ram[15][104] ), .S0(n4257), .S1(n4163), .Y(n4750) );
  MUX41X1_HVT U761 ( .A1(\ram[8][104] ), .A3(\ram[10][104] ), .A2(
        \ram[9][104] ), .A4(\ram[11][104] ), .S0(n4257), .S1(n4163), .Y(n4751)
         );
  MUX41X1_HVT U762 ( .A1(\ram[4][104] ), .A3(\ram[6][104] ), .A2(\ram[5][104] ), .A4(\ram[7][104] ), .S0(n4257), .S1(n4163), .Y(n4752) );
  MUX41X1_HVT U763 ( .A1(\ram[0][104] ), .A3(\ram[2][104] ), .A2(\ram[1][104] ), .A4(\ram[3][104] ), .S0(n4257), .S1(n4163), .Y(n4753) );
  MUX41X1_HVT U764 ( .A1(n4753), .A3(n4751), .A2(n4752), .A4(n4750), .S0(n4318), .S1(n4295), .Y(q[104]) );
  MUX41X1_HVT U765 ( .A1(\ram[12][105] ), .A3(\ram[14][105] ), .A2(
        \ram[13][105] ), .A4(\ram[15][105] ), .S0(n4258), .S1(n4164), .Y(n4754) );
  MUX41X1_HVT U766 ( .A1(\ram[8][105] ), .A3(\ram[10][105] ), .A2(
        \ram[9][105] ), .A4(\ram[11][105] ), .S0(n4258), .S1(n4164), .Y(n4755)
         );
  MUX41X1_HVT U767 ( .A1(\ram[4][105] ), .A3(\ram[6][105] ), .A2(\ram[5][105] ), .A4(\ram[7][105] ), .S0(n4258), .S1(n4164), .Y(n4756) );
  MUX41X1_HVT U768 ( .A1(\ram[0][105] ), .A3(\ram[2][105] ), .A2(\ram[1][105] ), .A4(\ram[3][105] ), .S0(n4258), .S1(n4164), .Y(n4757) );
  MUX41X1_HVT U769 ( .A1(n4757), .A3(n4755), .A2(n4756), .A4(n4754), .S0(n4318), .S1(n4295), .Y(q[105]) );
  MUX41X1_HVT U770 ( .A1(\ram[12][106] ), .A3(\ram[14][106] ), .A2(
        \ram[13][106] ), .A4(\ram[15][106] ), .S0(n4258), .S1(n4164), .Y(n4758) );
  MUX41X1_HVT U771 ( .A1(\ram[8][106] ), .A3(\ram[10][106] ), .A2(
        \ram[9][106] ), .A4(\ram[11][106] ), .S0(n4258), .S1(n4164), .Y(n4759)
         );
  MUX41X1_HVT U772 ( .A1(\ram[4][106] ), .A3(\ram[6][106] ), .A2(\ram[5][106] ), .A4(\ram[7][106] ), .S0(n4258), .S1(n4164), .Y(n4760) );
  MUX41X1_HVT U773 ( .A1(\ram[0][106] ), .A3(\ram[2][106] ), .A2(\ram[1][106] ), .A4(\ram[3][106] ), .S0(n4258), .S1(n4164), .Y(n4761) );
  MUX41X1_HVT U774 ( .A1(n4761), .A3(n4759), .A2(n4760), .A4(n4758), .S0(n4318), .S1(n4295), .Y(q[106]) );
  MUX41X1_HVT U775 ( .A1(\ram[12][107] ), .A3(\ram[14][107] ), .A2(
        \ram[13][107] ), .A4(\ram[15][107] ), .S0(n4258), .S1(n4164), .Y(n4762) );
  MUX41X1_HVT U776 ( .A1(\ram[8][107] ), .A3(\ram[10][107] ), .A2(
        \ram[9][107] ), .A4(\ram[11][107] ), .S0(n4258), .S1(n4164), .Y(n4763)
         );
  MUX41X1_HVT U777 ( .A1(\ram[4][107] ), .A3(\ram[6][107] ), .A2(\ram[5][107] ), .A4(\ram[7][107] ), .S0(n4258), .S1(n4164), .Y(n4764) );
  MUX41X1_HVT U778 ( .A1(\ram[0][107] ), .A3(\ram[2][107] ), .A2(\ram[1][107] ), .A4(\ram[3][107] ), .S0(n4258), .S1(n4164), .Y(n4765) );
  MUX41X1_HVT U779 ( .A1(n4765), .A3(n4763), .A2(n4764), .A4(n4762), .S0(n4318), .S1(n4295), .Y(q[107]) );
  MUX41X1_HVT U780 ( .A1(\ram[12][108] ), .A3(\ram[14][108] ), .A2(
        \ram[13][108] ), .A4(\ram[15][108] ), .S0(n4259), .S1(n4165), .Y(n4766) );
  MUX41X1_HVT U781 ( .A1(\ram[8][108] ), .A3(\ram[10][108] ), .A2(
        \ram[9][108] ), .A4(\ram[11][108] ), .S0(n4259), .S1(n4165), .Y(n4767)
         );
  MUX41X1_HVT U782 ( .A1(\ram[4][108] ), .A3(\ram[6][108] ), .A2(\ram[5][108] ), .A4(\ram[7][108] ), .S0(n4259), .S1(n4165), .Y(n4768) );
  MUX41X1_HVT U783 ( .A1(\ram[0][108] ), .A3(\ram[2][108] ), .A2(\ram[1][108] ), .A4(\ram[3][108] ), .S0(n4259), .S1(n4165), .Y(n4769) );
  MUX41X1_HVT U784 ( .A1(n4769), .A3(n4767), .A2(n4768), .A4(n4766), .S0(n4319), .S1(n4296), .Y(q[108]) );
  MUX41X1_HVT U785 ( .A1(\ram[12][109] ), .A3(\ram[14][109] ), .A2(
        \ram[13][109] ), .A4(\ram[15][109] ), .S0(n4259), .S1(n4165), .Y(n4770) );
  MUX41X1_HVT U786 ( .A1(\ram[8][109] ), .A3(\ram[10][109] ), .A2(
        \ram[9][109] ), .A4(\ram[11][109] ), .S0(n4259), .S1(n4165), .Y(n4771)
         );
  MUX41X1_HVT U787 ( .A1(\ram[4][109] ), .A3(\ram[6][109] ), .A2(\ram[5][109] ), .A4(\ram[7][109] ), .S0(n4259), .S1(n4165), .Y(n4772) );
  MUX41X1_HVT U788 ( .A1(\ram[0][109] ), .A3(\ram[2][109] ), .A2(\ram[1][109] ), .A4(\ram[3][109] ), .S0(n4259), .S1(n4165), .Y(n4773) );
  MUX41X1_HVT U789 ( .A1(n4773), .A3(n4771), .A2(n4772), .A4(n4770), .S0(n4319), .S1(n4296), .Y(q[109]) );
  MUX41X1_HVT U790 ( .A1(\ram[12][110] ), .A3(\ram[14][110] ), .A2(
        \ram[13][110] ), .A4(\ram[15][110] ), .S0(n4259), .S1(n4165), .Y(n4774) );
  MUX41X1_HVT U791 ( .A1(\ram[8][110] ), .A3(\ram[10][110] ), .A2(
        \ram[9][110] ), .A4(\ram[11][110] ), .S0(n4259), .S1(n4165), .Y(n4775)
         );
  MUX41X1_HVT U792 ( .A1(\ram[4][110] ), .A3(\ram[6][110] ), .A2(\ram[5][110] ), .A4(\ram[7][110] ), .S0(n4259), .S1(n4165), .Y(n4776) );
  MUX41X1_HVT U793 ( .A1(\ram[0][110] ), .A3(\ram[2][110] ), .A2(\ram[1][110] ), .A4(\ram[3][110] ), .S0(n4259), .S1(n4165), .Y(n4777) );
  MUX41X1_HVT U794 ( .A1(n4777), .A3(n4775), .A2(n4776), .A4(n4774), .S0(n4319), .S1(n4296), .Y(q[110]) );
  MUX41X1_HVT U795 ( .A1(\ram[12][111] ), .A3(\ram[14][111] ), .A2(
        \ram[13][111] ), .A4(\ram[15][111] ), .S0(n4260), .S1(n4166), .Y(n4778) );
  MUX41X1_HVT U796 ( .A1(\ram[8][111] ), .A3(\ram[10][111] ), .A2(
        \ram[9][111] ), .A4(\ram[11][111] ), .S0(n4260), .S1(n4166), .Y(n4779)
         );
  MUX41X1_HVT U797 ( .A1(\ram[4][111] ), .A3(\ram[6][111] ), .A2(\ram[5][111] ), .A4(\ram[7][111] ), .S0(n4260), .S1(n4166), .Y(n4780) );
  MUX41X1_HVT U798 ( .A1(\ram[0][111] ), .A3(\ram[2][111] ), .A2(\ram[1][111] ), .A4(\ram[3][111] ), .S0(n4260), .S1(n4166), .Y(n4781) );
  MUX41X1_HVT U799 ( .A1(n4781), .A3(n4779), .A2(n4780), .A4(n4778), .S0(n4319), .S1(n4296), .Y(q[111]) );
  MUX41X1_HVT U800 ( .A1(\ram[12][112] ), .A3(\ram[14][112] ), .A2(
        \ram[13][112] ), .A4(\ram[15][112] ), .S0(n4260), .S1(n4166), .Y(n4782) );
  MUX41X1_HVT U801 ( .A1(\ram[8][112] ), .A3(\ram[10][112] ), .A2(
        \ram[9][112] ), .A4(\ram[11][112] ), .S0(n4260), .S1(n4166), .Y(n4783)
         );
  MUX41X1_HVT U802 ( .A1(\ram[4][112] ), .A3(\ram[6][112] ), .A2(\ram[5][112] ), .A4(\ram[7][112] ), .S0(n4260), .S1(n4166), .Y(n4784) );
  MUX41X1_HVT U803 ( .A1(\ram[0][112] ), .A3(\ram[2][112] ), .A2(\ram[1][112] ), .A4(\ram[3][112] ), .S0(n4260), .S1(n4166), .Y(n4785) );
  MUX41X1_HVT U804 ( .A1(n4785), .A3(n4783), .A2(n4784), .A4(n4782), .S0(n4319), .S1(n4296), .Y(q[112]) );
  MUX41X1_HVT U805 ( .A1(\ram[12][113] ), .A3(\ram[14][113] ), .A2(
        \ram[13][113] ), .A4(\ram[15][113] ), .S0(n4260), .S1(n4166), .Y(n4786) );
  MUX41X1_HVT U806 ( .A1(\ram[8][113] ), .A3(\ram[10][113] ), .A2(
        \ram[9][113] ), .A4(\ram[11][113] ), .S0(n4260), .S1(n4166), .Y(n4787)
         );
  MUX41X1_HVT U807 ( .A1(\ram[4][113] ), .A3(\ram[6][113] ), .A2(\ram[5][113] ), .A4(\ram[7][113] ), .S0(n4260), .S1(n4166), .Y(n4788) );
  MUX41X1_HVT U808 ( .A1(\ram[0][113] ), .A3(\ram[2][113] ), .A2(\ram[1][113] ), .A4(\ram[3][113] ), .S0(n4261), .S1(n4167), .Y(n4789) );
  MUX41X1_HVT U809 ( .A1(n4789), .A3(n4787), .A2(n4788), .A4(n4786), .S0(n4319), .S1(n4296), .Y(q[113]) );
  MUX41X1_HVT U810 ( .A1(\ram[12][114] ), .A3(\ram[14][114] ), .A2(
        \ram[13][114] ), .A4(\ram[15][114] ), .S0(n4261), .S1(n4167), .Y(n4790) );
  MUX41X1_HVT U811 ( .A1(\ram[8][114] ), .A3(\ram[10][114] ), .A2(
        \ram[9][114] ), .A4(\ram[11][114] ), .S0(n4261), .S1(n4167), .Y(n4791)
         );
  MUX41X1_HVT U812 ( .A1(\ram[4][114] ), .A3(\ram[6][114] ), .A2(\ram[5][114] ), .A4(\ram[7][114] ), .S0(n4261), .S1(n4167), .Y(n4792) );
  MUX41X1_HVT U813 ( .A1(\ram[0][114] ), .A3(\ram[2][114] ), .A2(\ram[1][114] ), .A4(\ram[3][114] ), .S0(n4261), .S1(n4167), .Y(n4793) );
  MUX41X1_HVT U814 ( .A1(n4793), .A3(n4791), .A2(n4792), .A4(n4790), .S0(n4319), .S1(n4296), .Y(q[114]) );
  MUX41X1_HVT U815 ( .A1(\ram[12][115] ), .A3(\ram[14][115] ), .A2(
        \ram[13][115] ), .A4(\ram[15][115] ), .S0(n4261), .S1(n4167), .Y(n4794) );
  MUX41X1_HVT U816 ( .A1(\ram[8][115] ), .A3(\ram[10][115] ), .A2(
        \ram[9][115] ), .A4(\ram[11][115] ), .S0(n4261), .S1(n4167), .Y(n4795)
         );
  MUX41X1_HVT U817 ( .A1(\ram[4][115] ), .A3(\ram[6][115] ), .A2(\ram[5][115] ), .A4(\ram[7][115] ), .S0(n4261), .S1(n4167), .Y(n4796) );
  MUX41X1_HVT U818 ( .A1(\ram[0][115] ), .A3(\ram[2][115] ), .A2(\ram[1][115] ), .A4(\ram[3][115] ), .S0(n4261), .S1(n4167), .Y(n4797) );
  MUX41X1_HVT U819 ( .A1(n4797), .A3(n4795), .A2(n4796), .A4(n4794), .S0(n4319), .S1(n4296), .Y(q[115]) );
  MUX41X1_HVT U820 ( .A1(\ram[12][116] ), .A3(\ram[14][116] ), .A2(
        \ram[13][116] ), .A4(\ram[15][116] ), .S0(n4261), .S1(n4167), .Y(n4798) );
  MUX41X1_HVT U821 ( .A1(\ram[8][116] ), .A3(\ram[10][116] ), .A2(
        \ram[9][116] ), .A4(\ram[11][116] ), .S0(n4261), .S1(n4167), .Y(n4799)
         );
  MUX41X1_HVT U822 ( .A1(\ram[4][116] ), .A3(\ram[6][116] ), .A2(\ram[5][116] ), .A4(\ram[7][116] ), .S0(n4261), .S1(n4167), .Y(n4800) );
  MUX41X1_HVT U823 ( .A1(\ram[0][116] ), .A3(\ram[2][116] ), .A2(\ram[1][116] ), .A4(\ram[3][116] ), .S0(n4262), .S1(n4168), .Y(n4801) );
  MUX41X1_HVT U824 ( .A1(n4801), .A3(n4799), .A2(n4800), .A4(n4798), .S0(n4319), .S1(n4296), .Y(q[116]) );
  MUX41X1_HVT U825 ( .A1(\ram[12][117] ), .A3(\ram[14][117] ), .A2(
        \ram[13][117] ), .A4(\ram[15][117] ), .S0(n4262), .S1(n4168), .Y(n4802) );
  MUX41X1_HVT U826 ( .A1(\ram[8][117] ), .A3(\ram[10][117] ), .A2(
        \ram[9][117] ), .A4(\ram[11][117] ), .S0(n4262), .S1(n4168), .Y(n4803)
         );
  MUX41X1_HVT U827 ( .A1(\ram[4][117] ), .A3(\ram[6][117] ), .A2(\ram[5][117] ), .A4(\ram[7][117] ), .S0(n4262), .S1(n4168), .Y(n4804) );
  MUX41X1_HVT U828 ( .A1(\ram[0][117] ), .A3(\ram[2][117] ), .A2(\ram[1][117] ), .A4(\ram[3][117] ), .S0(n4262), .S1(n4168), .Y(n4805) );
  MUX41X1_HVT U829 ( .A1(n4805), .A3(n4803), .A2(n4804), .A4(n4802), .S0(n4319), .S1(n4296), .Y(q[117]) );
  MUX41X1_HVT U830 ( .A1(\ram[12][118] ), .A3(\ram[14][118] ), .A2(
        \ram[13][118] ), .A4(\ram[15][118] ), .S0(n4262), .S1(n4168), .Y(n4806) );
  MUX41X1_HVT U831 ( .A1(\ram[8][118] ), .A3(\ram[10][118] ), .A2(
        \ram[9][118] ), .A4(\ram[11][118] ), .S0(n4262), .S1(n4168), .Y(n4807)
         );
  MUX41X1_HVT U832 ( .A1(\ram[4][118] ), .A3(\ram[6][118] ), .A2(\ram[5][118] ), .A4(\ram[7][118] ), .S0(n4262), .S1(n4168), .Y(n4808) );
  MUX41X1_HVT U833 ( .A1(\ram[0][118] ), .A3(\ram[2][118] ), .A2(\ram[1][118] ), .A4(\ram[3][118] ), .S0(n4262), .S1(n4168), .Y(n4809) );
  MUX41X1_HVT U834 ( .A1(n4809), .A3(n4807), .A2(n4808), .A4(n4806), .S0(n4319), .S1(n4296), .Y(q[118]) );
  MUX41X1_HVT U835 ( .A1(\ram[12][119] ), .A3(\ram[14][119] ), .A2(
        \ram[13][119] ), .A4(\ram[15][119] ), .S0(n4262), .S1(n4168), .Y(n4810) );
  MUX41X1_HVT U836 ( .A1(\ram[8][119] ), .A3(\ram[10][119] ), .A2(
        \ram[9][119] ), .A4(\ram[11][119] ), .S0(n4262), .S1(n4168), .Y(n4811)
         );
  MUX41X1_HVT U837 ( .A1(\ram[4][119] ), .A3(\ram[6][119] ), .A2(\ram[5][119] ), .A4(\ram[7][119] ), .S0(n4262), .S1(n4168), .Y(n4812) );
  MUX41X1_HVT U838 ( .A1(\ram[0][119] ), .A3(\ram[2][119] ), .A2(\ram[1][119] ), .A4(\ram[3][119] ), .S0(n4263), .S1(n4169), .Y(n4813) );
  MUX41X1_HVT U839 ( .A1(n4813), .A3(n4811), .A2(n4812), .A4(n4810), .S0(n4319), .S1(n4296), .Y(q[119]) );
  MUX41X1_HVT U840 ( .A1(\ram[12][120] ), .A3(\ram[14][120] ), .A2(
        \ram[13][120] ), .A4(\ram[15][120] ), .S0(n4263), .S1(n4169), .Y(n4814) );
  MUX41X1_HVT U841 ( .A1(\ram[8][120] ), .A3(\ram[10][120] ), .A2(
        \ram[9][120] ), .A4(\ram[11][120] ), .S0(n4263), .S1(n4169), .Y(n4815)
         );
  MUX41X1_HVT U842 ( .A1(\ram[4][120] ), .A3(\ram[6][120] ), .A2(\ram[5][120] ), .A4(\ram[7][120] ), .S0(n4263), .S1(n4169), .Y(n4816) );
  MUX41X1_HVT U843 ( .A1(\ram[0][120] ), .A3(\ram[2][120] ), .A2(\ram[1][120] ), .A4(\ram[3][120] ), .S0(n4263), .S1(n4169), .Y(n4817) );
  MUX41X1_HVT U844 ( .A1(n4817), .A3(n4815), .A2(n4816), .A4(n4814), .S0(n4320), .S1(n4297), .Y(q[120]) );
  MUX41X1_HVT U845 ( .A1(\ram[12][121] ), .A3(\ram[14][121] ), .A2(
        \ram[13][121] ), .A4(\ram[15][121] ), .S0(n4263), .S1(n4169), .Y(n4818) );
  MUX41X1_HVT U846 ( .A1(\ram[8][121] ), .A3(\ram[10][121] ), .A2(
        \ram[9][121] ), .A4(\ram[11][121] ), .S0(n4263), .S1(n4169), .Y(n4819)
         );
  MUX41X1_HVT U847 ( .A1(\ram[4][121] ), .A3(\ram[6][121] ), .A2(\ram[5][121] ), .A4(\ram[7][121] ), .S0(n4263), .S1(n4169), .Y(n4820) );
  MUX41X1_HVT U848 ( .A1(\ram[0][121] ), .A3(\ram[2][121] ), .A2(\ram[1][121] ), .A4(\ram[3][121] ), .S0(n4263), .S1(n4169), .Y(n4821) );
  MUX41X1_HVT U849 ( .A1(n4821), .A3(n4819), .A2(n4820), .A4(n4818), .S0(n4320), .S1(n4297), .Y(q[121]) );
  MUX41X1_HVT U850 ( .A1(\ram[12][122] ), .A3(\ram[14][122] ), .A2(
        \ram[13][122] ), .A4(\ram[15][122] ), .S0(n4263), .S1(n4169), .Y(n4822) );
  MUX41X1_HVT U851 ( .A1(\ram[8][122] ), .A3(\ram[10][122] ), .A2(
        \ram[9][122] ), .A4(\ram[11][122] ), .S0(n4263), .S1(n4169), .Y(n4823)
         );
  MUX41X1_HVT U852 ( .A1(\ram[4][122] ), .A3(\ram[6][122] ), .A2(\ram[5][122] ), .A4(\ram[7][122] ), .S0(n4263), .S1(n4169), .Y(n4824) );
  MUX41X1_HVT U853 ( .A1(\ram[0][122] ), .A3(\ram[2][122] ), .A2(\ram[1][122] ), .A4(\ram[3][122] ), .S0(n4264), .S1(n4170), .Y(n4825) );
  MUX41X1_HVT U854 ( .A1(n4825), .A3(n4823), .A2(n4824), .A4(n4822), .S0(n4320), .S1(n4297), .Y(q[122]) );
  MUX41X1_HVT U855 ( .A1(\ram[12][123] ), .A3(\ram[14][123] ), .A2(
        \ram[13][123] ), .A4(\ram[15][123] ), .S0(n4264), .S1(n4170), .Y(n4826) );
  MUX41X1_HVT U856 ( .A1(\ram[8][123] ), .A3(\ram[10][123] ), .A2(
        \ram[9][123] ), .A4(\ram[11][123] ), .S0(n4264), .S1(n4170), .Y(n4827)
         );
  MUX41X1_HVT U857 ( .A1(\ram[4][123] ), .A3(\ram[6][123] ), .A2(\ram[5][123] ), .A4(\ram[7][123] ), .S0(n4264), .S1(n4170), .Y(n4828) );
  MUX41X1_HVT U858 ( .A1(\ram[0][123] ), .A3(\ram[2][123] ), .A2(\ram[1][123] ), .A4(\ram[3][123] ), .S0(n4264), .S1(n4170), .Y(n4829) );
  MUX41X1_HVT U859 ( .A1(n4829), .A3(n4827), .A2(n4828), .A4(n4826), .S0(n4320), .S1(n4297), .Y(q[123]) );
  MUX41X1_HVT U860 ( .A1(\ram[12][124] ), .A3(\ram[14][124] ), .A2(
        \ram[13][124] ), .A4(\ram[15][124] ), .S0(n4264), .S1(n4170), .Y(n4830) );
  MUX41X1_HVT U861 ( .A1(\ram[8][124] ), .A3(\ram[10][124] ), .A2(
        \ram[9][124] ), .A4(\ram[11][124] ), .S0(n4264), .S1(n4170), .Y(n4831)
         );
  MUX41X1_HVT U862 ( .A1(\ram[4][124] ), .A3(\ram[6][124] ), .A2(\ram[5][124] ), .A4(\ram[7][124] ), .S0(n4264), .S1(n4170), .Y(n4832) );
  MUX41X1_HVT U863 ( .A1(\ram[0][124] ), .A3(\ram[2][124] ), .A2(\ram[1][124] ), .A4(\ram[3][124] ), .S0(n4264), .S1(n4170), .Y(n4833) );
  MUX41X1_HVT U864 ( .A1(n4833), .A3(n4831), .A2(n4832), .A4(n4830), .S0(n4320), .S1(n4297), .Y(q[124]) );
  MUX41X1_HVT U865 ( .A1(\ram[12][125] ), .A3(\ram[14][125] ), .A2(
        \ram[13][125] ), .A4(\ram[15][125] ), .S0(n4264), .S1(n4170), .Y(n4834) );
  MUX41X1_HVT U866 ( .A1(\ram[8][125] ), .A3(\ram[10][125] ), .A2(
        \ram[9][125] ), .A4(\ram[11][125] ), .S0(n4264), .S1(n4170), .Y(n4835)
         );
  MUX41X1_HVT U867 ( .A1(\ram[4][125] ), .A3(\ram[6][125] ), .A2(\ram[5][125] ), .A4(\ram[7][125] ), .S0(n4264), .S1(n4170), .Y(n4836) );
  MUX41X1_HVT U868 ( .A1(\ram[0][125] ), .A3(\ram[2][125] ), .A2(\ram[1][125] ), .A4(\ram[3][125] ), .S0(n4265), .S1(n4171), .Y(n4837) );
  MUX41X1_HVT U869 ( .A1(n4837), .A3(n4835), .A2(n4836), .A4(n4834), .S0(n4320), .S1(n4297), .Y(q[125]) );
  MUX41X1_HVT U870 ( .A1(\ram[12][126] ), .A3(\ram[14][126] ), .A2(
        \ram[13][126] ), .A4(\ram[15][126] ), .S0(n4265), .S1(n4171), .Y(n4838) );
  MUX41X1_HVT U871 ( .A1(\ram[8][126] ), .A3(\ram[10][126] ), .A2(
        \ram[9][126] ), .A4(\ram[11][126] ), .S0(n4265), .S1(n4171), .Y(n4839)
         );
  MUX41X1_HVT U872 ( .A1(\ram[4][126] ), .A3(\ram[6][126] ), .A2(\ram[5][126] ), .A4(\ram[7][126] ), .S0(n4265), .S1(n4171), .Y(n4840) );
  MUX41X1_HVT U873 ( .A1(\ram[0][126] ), .A3(\ram[2][126] ), .A2(\ram[1][126] ), .A4(\ram[3][126] ), .S0(n4265), .S1(n4171), .Y(n4841) );
  MUX41X1_HVT U874 ( .A1(n4841), .A3(n4839), .A2(n4840), .A4(n4838), .S0(n4320), .S1(n4297), .Y(q[126]) );
  MUX41X1_HVT U875 ( .A1(\ram[12][127] ), .A3(\ram[14][127] ), .A2(
        \ram[13][127] ), .A4(\ram[15][127] ), .S0(n4265), .S1(n4171), .Y(n4842) );
  MUX41X1_HVT U876 ( .A1(\ram[8][127] ), .A3(\ram[10][127] ), .A2(
        \ram[9][127] ), .A4(\ram[11][127] ), .S0(n4265), .S1(n4171), .Y(n4843)
         );
  MUX41X1_HVT U877 ( .A1(\ram[4][127] ), .A3(\ram[6][127] ), .A2(\ram[5][127] ), .A4(\ram[7][127] ), .S0(n4265), .S1(n4171), .Y(n4844) );
  MUX41X1_HVT U878 ( .A1(\ram[0][127] ), .A3(\ram[2][127] ), .A2(\ram[1][127] ), .A4(\ram[3][127] ), .S0(n4265), .S1(n4171), .Y(n4845) );
  MUX41X1_HVT U879 ( .A1(n4845), .A3(n4843), .A2(n4844), .A4(n4842), .S0(n4320), .S1(n4297), .Y(q[127]) );
  MUX41X1_HVT U880 ( .A1(\ram[12][128] ), .A3(\ram[14][128] ), .A2(
        \ram[13][128] ), .A4(\ram[15][128] ), .S0(n4212), .S1(n22), .Y(n4846)
         );
  MUX41X1_HVT U881 ( .A1(\ram[8][128] ), .A3(\ram[10][128] ), .A2(
        \ram[9][128] ), .A4(\ram[11][128] ), .S0(n4207), .S1(n17), .Y(n4847)
         );
  MUX41X1_HVT U882 ( .A1(\ram[4][128] ), .A3(\ram[6][128] ), .A2(\ram[5][128] ), .A4(\ram[7][128] ), .S0(n4201), .S1(n11), .Y(n4848) );
  MUX41X1_HVT U883 ( .A1(\ram[0][128] ), .A3(\ram[2][128] ), .A2(\ram[1][128] ), .A4(\ram[3][128] ), .S0(n4201), .S1(n11), .Y(n4849) );
  MUX41X1_HVT U884 ( .A1(n4849), .A3(n4847), .A2(n4848), .A4(n4846), .S0(n4320), .S1(n4297), .Y(q[128]) );
  MUX41X1_HVT U885 ( .A1(\ram[12][129] ), .A3(\ram[14][129] ), .A2(
        \ram[13][129] ), .A4(\ram[15][129] ), .S0(n4201), .S1(n11), .Y(n4850)
         );
  MUX41X1_HVT U886 ( .A1(\ram[8][129] ), .A3(\ram[10][129] ), .A2(
        \ram[9][129] ), .A4(\ram[11][129] ), .S0(n4202), .S1(n12), .Y(n4851)
         );
  MUX41X1_HVT U887 ( .A1(\ram[4][129] ), .A3(\ram[6][129] ), .A2(\ram[5][129] ), .A4(\ram[7][129] ), .S0(n4202), .S1(n12), .Y(n4852) );
  MUX41X1_HVT U888 ( .A1(\ram[0][129] ), .A3(\ram[2][129] ), .A2(\ram[1][129] ), .A4(\ram[3][129] ), .S0(n4202), .S1(n12), .Y(n4853) );
  MUX41X1_HVT U889 ( .A1(n4853), .A3(n4851), .A2(n4852), .A4(n4850), .S0(n4320), .S1(n4297), .Y(q[129]) );
  MUX41X1_HVT U890 ( .A1(\ram[12][130] ), .A3(\ram[14][130] ), .A2(
        \ram[13][130] ), .A4(\ram[15][130] ), .S0(n4202), .S1(n12), .Y(n4854)
         );
  MUX41X1_HVT U891 ( .A1(\ram[8][130] ), .A3(\ram[10][130] ), .A2(
        \ram[9][130] ), .A4(\ram[11][130] ), .S0(n4202), .S1(n12), .Y(n4855)
         );
  MUX41X1_HVT U892 ( .A1(\ram[4][130] ), .A3(\ram[6][130] ), .A2(\ram[5][130] ), .A4(\ram[7][130] ), .S0(n4202), .S1(n12), .Y(n4856) );
  MUX41X1_HVT U893 ( .A1(\ram[0][130] ), .A3(\ram[2][130] ), .A2(\ram[1][130] ), .A4(\ram[3][130] ), .S0(n4202), .S1(n12), .Y(n4857) );
  MUX41X1_HVT U894 ( .A1(n4857), .A3(n4855), .A2(n4856), .A4(n4854), .S0(n4320), .S1(n4297), .Y(q[130]) );
  MUX41X1_HVT U895 ( .A1(\ram[12][131] ), .A3(\ram[14][131] ), .A2(
        \ram[13][131] ), .A4(\ram[15][131] ), .S0(n4202), .S1(n12), .Y(n4858)
         );
  MUX41X1_HVT U896 ( .A1(\ram[8][131] ), .A3(\ram[10][131] ), .A2(
        \ram[9][131] ), .A4(\ram[11][131] ), .S0(n4202), .S1(n12), .Y(n4859)
         );
  MUX41X1_HVT U897 ( .A1(\ram[4][131] ), .A3(\ram[6][131] ), .A2(\ram[5][131] ), .A4(\ram[7][131] ), .S0(n4202), .S1(n12), .Y(n4860) );
  MUX41X1_HVT U898 ( .A1(\ram[0][131] ), .A3(\ram[2][131] ), .A2(\ram[1][131] ), .A4(\ram[3][131] ), .S0(n4202), .S1(n12), .Y(n4861) );
  MUX41X1_HVT U899 ( .A1(n4861), .A3(n4859), .A2(n4860), .A4(n4858), .S0(n4320), .S1(n4297), .Y(q[131]) );
  MUX41X1_HVT U900 ( .A1(\ram[12][132] ), .A3(\ram[14][132] ), .A2(
        \ram[13][132] ), .A4(\ram[15][132] ), .S0(n4202), .S1(n12), .Y(n4862)
         );
  MUX41X1_HVT U901 ( .A1(\ram[8][132] ), .A3(\ram[10][132] ), .A2(
        \ram[9][132] ), .A4(\ram[11][132] ), .S0(n4203), .S1(n13), .Y(n4863)
         );
  MUX41X1_HVT U902 ( .A1(\ram[4][132] ), .A3(\ram[6][132] ), .A2(\ram[5][132] ), .A4(\ram[7][132] ), .S0(n4203), .S1(n13), .Y(n4864) );
  MUX41X1_HVT U903 ( .A1(\ram[0][132] ), .A3(\ram[2][132] ), .A2(\ram[1][132] ), .A4(\ram[3][132] ), .S0(n4203), .S1(n13), .Y(n4865) );
  MUX41X1_HVT U904 ( .A1(n4865), .A3(n4863), .A2(n4864), .A4(n4862), .S0(n4321), .S1(n4298), .Y(q[132]) );
  MUX41X1_HVT U905 ( .A1(\ram[12][133] ), .A3(\ram[14][133] ), .A2(
        \ram[13][133] ), .A4(\ram[15][133] ), .S0(n4203), .S1(n13), .Y(n4866)
         );
  MUX41X1_HVT U906 ( .A1(\ram[8][133] ), .A3(\ram[10][133] ), .A2(
        \ram[9][133] ), .A4(\ram[11][133] ), .S0(n4203), .S1(n13), .Y(n4867)
         );
  MUX41X1_HVT U907 ( .A1(\ram[4][133] ), .A3(\ram[6][133] ), .A2(\ram[5][133] ), .A4(\ram[7][133] ), .S0(n4203), .S1(n13), .Y(n4868) );
  MUX41X1_HVT U908 ( .A1(\ram[0][133] ), .A3(\ram[2][133] ), .A2(\ram[1][133] ), .A4(\ram[3][133] ), .S0(n4203), .S1(n13), .Y(n4869) );
  MUX41X1_HVT U909 ( .A1(n4869), .A3(n4867), .A2(n4868), .A4(n4866), .S0(n4321), .S1(n4298), .Y(q[133]) );
  MUX41X1_HVT U910 ( .A1(\ram[12][134] ), .A3(\ram[14][134] ), .A2(
        \ram[13][134] ), .A4(\ram[15][134] ), .S0(n4203), .S1(n13), .Y(n4870)
         );
  MUX41X1_HVT U911 ( .A1(\ram[8][134] ), .A3(\ram[10][134] ), .A2(
        \ram[9][134] ), .A4(\ram[11][134] ), .S0(n4203), .S1(n13), .Y(n4871)
         );
  MUX41X1_HVT U912 ( .A1(\ram[4][134] ), .A3(\ram[6][134] ), .A2(\ram[5][134] ), .A4(\ram[7][134] ), .S0(n4203), .S1(n13), .Y(n4872) );
  MUX41X1_HVT U913 ( .A1(\ram[0][134] ), .A3(\ram[2][134] ), .A2(\ram[1][134] ), .A4(\ram[3][134] ), .S0(n4203), .S1(n13), .Y(n4873) );
  MUX41X1_HVT U914 ( .A1(n4873), .A3(n4871), .A2(n4872), .A4(n4870), .S0(n4321), .S1(n4298), .Y(q[134]) );
  MUX41X1_HVT U915 ( .A1(\ram[12][135] ), .A3(\ram[14][135] ), .A2(
        \ram[13][135] ), .A4(\ram[15][135] ), .S0(n4203), .S1(n13), .Y(n4874)
         );
  MUX41X1_HVT U916 ( .A1(\ram[8][135] ), .A3(\ram[10][135] ), .A2(
        \ram[9][135] ), .A4(\ram[11][135] ), .S0(n4204), .S1(n14), .Y(n4875)
         );
  MUX41X1_HVT U917 ( .A1(\ram[4][135] ), .A3(\ram[6][135] ), .A2(\ram[5][135] ), .A4(\ram[7][135] ), .S0(n4204), .S1(n14), .Y(n4876) );
  MUX41X1_HVT U918 ( .A1(\ram[0][135] ), .A3(\ram[2][135] ), .A2(\ram[1][135] ), .A4(\ram[3][135] ), .S0(n4204), .S1(n14), .Y(n4877) );
  MUX41X1_HVT U919 ( .A1(n4877), .A3(n4875), .A2(n4876), .A4(n4874), .S0(n4321), .S1(n4298), .Y(q[135]) );
  MUX41X1_HVT U920 ( .A1(\ram[12][136] ), .A3(\ram[14][136] ), .A2(
        \ram[13][136] ), .A4(\ram[15][136] ), .S0(n4204), .S1(n14), .Y(n4878)
         );
  MUX41X1_HVT U921 ( .A1(\ram[8][136] ), .A3(\ram[10][136] ), .A2(
        \ram[9][136] ), .A4(\ram[11][136] ), .S0(n4204), .S1(n14), .Y(n4879)
         );
  MUX41X1_HVT U922 ( .A1(\ram[4][136] ), .A3(\ram[6][136] ), .A2(\ram[5][136] ), .A4(\ram[7][136] ), .S0(n4204), .S1(n14), .Y(n4880) );
  MUX41X1_HVT U923 ( .A1(\ram[0][136] ), .A3(\ram[2][136] ), .A2(\ram[1][136] ), .A4(\ram[3][136] ), .S0(n4204), .S1(n14), .Y(n4881) );
  MUX41X1_HVT U924 ( .A1(n4881), .A3(n4879), .A2(n4880), .A4(n4878), .S0(n4321), .S1(n4298), .Y(q[136]) );
  MUX41X1_HVT U925 ( .A1(\ram[12][137] ), .A3(\ram[14][137] ), .A2(
        \ram[13][137] ), .A4(\ram[15][137] ), .S0(n4204), .S1(n14), .Y(n4882)
         );
  MUX41X1_HVT U926 ( .A1(\ram[8][137] ), .A3(\ram[10][137] ), .A2(
        \ram[9][137] ), .A4(\ram[11][137] ), .S0(n4204), .S1(n14), .Y(n4883)
         );
  MUX41X1_HVT U927 ( .A1(\ram[4][137] ), .A3(\ram[6][137] ), .A2(\ram[5][137] ), .A4(\ram[7][137] ), .S0(n4204), .S1(n14), .Y(n4884) );
  MUX41X1_HVT U928 ( .A1(\ram[0][137] ), .A3(\ram[2][137] ), .A2(\ram[1][137] ), .A4(\ram[3][137] ), .S0(n4204), .S1(n14), .Y(n4885) );
  MUX41X1_HVT U929 ( .A1(n4885), .A3(n4883), .A2(n4884), .A4(n4882), .S0(n4321), .S1(n4298), .Y(q[137]) );
  MUX41X1_HVT U930 ( .A1(\ram[12][138] ), .A3(\ram[14][138] ), .A2(
        \ram[13][138] ), .A4(\ram[15][138] ), .S0(n4204), .S1(n14), .Y(n4886)
         );
  MUX41X1_HVT U931 ( .A1(\ram[8][138] ), .A3(\ram[10][138] ), .A2(
        \ram[9][138] ), .A4(\ram[11][138] ), .S0(n4205), .S1(n15), .Y(n4887)
         );
  MUX41X1_HVT U932 ( .A1(\ram[4][138] ), .A3(\ram[6][138] ), .A2(\ram[5][138] ), .A4(\ram[7][138] ), .S0(n4205), .S1(n15), .Y(n4888) );
  MUX41X1_HVT U933 ( .A1(\ram[0][138] ), .A3(\ram[2][138] ), .A2(\ram[1][138] ), .A4(\ram[3][138] ), .S0(n4205), .S1(n15), .Y(n4889) );
  MUX41X1_HVT U934 ( .A1(n4889), .A3(n4887), .A2(n4888), .A4(n4886), .S0(n4321), .S1(n4298), .Y(q[138]) );
  MUX41X1_HVT U935 ( .A1(\ram[12][139] ), .A3(\ram[14][139] ), .A2(
        \ram[13][139] ), .A4(\ram[15][139] ), .S0(n4205), .S1(n15), .Y(n4890)
         );
  MUX41X1_HVT U936 ( .A1(\ram[8][139] ), .A3(\ram[10][139] ), .A2(
        \ram[9][139] ), .A4(\ram[11][139] ), .S0(n4205), .S1(n15), .Y(n4891)
         );
  MUX41X1_HVT U937 ( .A1(\ram[4][139] ), .A3(\ram[6][139] ), .A2(\ram[5][139] ), .A4(\ram[7][139] ), .S0(n4205), .S1(n15), .Y(n4892) );
  MUX41X1_HVT U938 ( .A1(\ram[0][139] ), .A3(\ram[2][139] ), .A2(\ram[1][139] ), .A4(\ram[3][139] ), .S0(n4205), .S1(n15), .Y(n4893) );
  MUX41X1_HVT U939 ( .A1(n4893), .A3(n4891), .A2(n4892), .A4(n4890), .S0(n4321), .S1(n4298), .Y(q[139]) );
  MUX41X1_HVT U940 ( .A1(\ram[12][140] ), .A3(\ram[14][140] ), .A2(
        \ram[13][140] ), .A4(\ram[15][140] ), .S0(n4205), .S1(n15), .Y(n4894)
         );
  MUX41X1_HVT U941 ( .A1(\ram[8][140] ), .A3(\ram[10][140] ), .A2(
        \ram[9][140] ), .A4(\ram[11][140] ), .S0(n4205), .S1(n15), .Y(n4895)
         );
  MUX41X1_HVT U942 ( .A1(\ram[4][140] ), .A3(\ram[6][140] ), .A2(\ram[5][140] ), .A4(\ram[7][140] ), .S0(n4205), .S1(n15), .Y(n4896) );
  MUX41X1_HVT U943 ( .A1(\ram[0][140] ), .A3(\ram[2][140] ), .A2(\ram[1][140] ), .A4(\ram[3][140] ), .S0(n4205), .S1(n15), .Y(n4897) );
  MUX41X1_HVT U944 ( .A1(n4897), .A3(n4895), .A2(n4896), .A4(n4894), .S0(n4321), .S1(n4298), .Y(q[140]) );
  MUX41X1_HVT U945 ( .A1(\ram[12][141] ), .A3(\ram[14][141] ), .A2(
        \ram[13][141] ), .A4(\ram[15][141] ), .S0(n4205), .S1(n15), .Y(n4898)
         );
  MUX41X1_HVT U946 ( .A1(\ram[8][141] ), .A3(\ram[10][141] ), .A2(
        \ram[9][141] ), .A4(\ram[11][141] ), .S0(n4206), .S1(n16), .Y(n4899)
         );
  MUX41X1_HVT U947 ( .A1(\ram[4][141] ), .A3(\ram[6][141] ), .A2(\ram[5][141] ), .A4(\ram[7][141] ), .S0(n4206), .S1(n16), .Y(n4900) );
  MUX41X1_HVT U948 ( .A1(\ram[0][141] ), .A3(\ram[2][141] ), .A2(\ram[1][141] ), .A4(\ram[3][141] ), .S0(n4206), .S1(n16), .Y(n4901) );
  MUX41X1_HVT U949 ( .A1(n4901), .A3(n4899), .A2(n4900), .A4(n4898), .S0(n4321), .S1(n4298), .Y(q[141]) );
  MUX41X1_HVT U950 ( .A1(\ram[12][142] ), .A3(\ram[14][142] ), .A2(
        \ram[13][142] ), .A4(\ram[15][142] ), .S0(n4206), .S1(n16), .Y(n4902)
         );
  MUX41X1_HVT U951 ( .A1(\ram[8][142] ), .A3(\ram[10][142] ), .A2(
        \ram[9][142] ), .A4(\ram[11][142] ), .S0(n4206), .S1(n16), .Y(n4903)
         );
  MUX41X1_HVT U952 ( .A1(\ram[4][142] ), .A3(\ram[6][142] ), .A2(\ram[5][142] ), .A4(\ram[7][142] ), .S0(n4206), .S1(n16), .Y(n4904) );
  MUX41X1_HVT U953 ( .A1(\ram[0][142] ), .A3(\ram[2][142] ), .A2(\ram[1][142] ), .A4(\ram[3][142] ), .S0(n4206), .S1(n16), .Y(n4905) );
  MUX41X1_HVT U954 ( .A1(n4905), .A3(n4903), .A2(n4904), .A4(n4902), .S0(n4321), .S1(n4298), .Y(q[142]) );
  MUX41X1_HVT U955 ( .A1(\ram[12][143] ), .A3(\ram[14][143] ), .A2(
        \ram[13][143] ), .A4(\ram[15][143] ), .S0(n4206), .S1(n16), .Y(n4906)
         );
  MUX41X1_HVT U956 ( .A1(\ram[8][143] ), .A3(\ram[10][143] ), .A2(
        \ram[9][143] ), .A4(\ram[11][143] ), .S0(n4206), .S1(n16), .Y(n4907)
         );
  MUX41X1_HVT U957 ( .A1(\ram[4][143] ), .A3(\ram[6][143] ), .A2(\ram[5][143] ), .A4(\ram[7][143] ), .S0(n4206), .S1(n16), .Y(n4908) );
  MUX41X1_HVT U958 ( .A1(\ram[0][143] ), .A3(\ram[2][143] ), .A2(\ram[1][143] ), .A4(\ram[3][143] ), .S0(n4206), .S1(n16), .Y(n4909) );
  MUX41X1_HVT U959 ( .A1(n4909), .A3(n4907), .A2(n4908), .A4(n4906), .S0(n4321), .S1(n4298), .Y(q[143]) );
  MUX41X1_HVT U960 ( .A1(\ram[12][144] ), .A3(\ram[14][144] ), .A2(
        \ram[13][144] ), .A4(\ram[15][144] ), .S0(n4206), .S1(n16), .Y(n4910)
         );
  MUX41X1_HVT U961 ( .A1(\ram[8][144] ), .A3(\ram[10][144] ), .A2(
        \ram[9][144] ), .A4(\ram[11][144] ), .S0(n4207), .S1(n17), .Y(n4911)
         );
  MUX41X1_HVT U962 ( .A1(\ram[4][144] ), .A3(\ram[6][144] ), .A2(\ram[5][144] ), .A4(\ram[7][144] ), .S0(n4207), .S1(n17), .Y(n4912) );
  MUX41X1_HVT U963 ( .A1(\ram[0][144] ), .A3(\ram[2][144] ), .A2(\ram[1][144] ), .A4(\ram[3][144] ), .S0(n4207), .S1(n17), .Y(n4913) );
  MUX41X1_HVT U964 ( .A1(n4913), .A3(n4911), .A2(n4912), .A4(n4910), .S0(n4322), .S1(n4299), .Y(q[144]) );
  MUX41X1_HVT U965 ( .A1(\ram[12][145] ), .A3(\ram[14][145] ), .A2(
        \ram[13][145] ), .A4(\ram[15][145] ), .S0(n4207), .S1(n17), .Y(n4914)
         );
  MUX41X1_HVT U966 ( .A1(\ram[8][145] ), .A3(\ram[10][145] ), .A2(
        \ram[9][145] ), .A4(\ram[11][145] ), .S0(n4207), .S1(n17), .Y(n4915)
         );
  MUX41X1_HVT U967 ( .A1(\ram[4][145] ), .A3(\ram[6][145] ), .A2(\ram[5][145] ), .A4(\ram[7][145] ), .S0(n4207), .S1(n17), .Y(n4916) );
  MUX41X1_HVT U968 ( .A1(\ram[0][145] ), .A3(\ram[2][145] ), .A2(\ram[1][145] ), .A4(\ram[3][145] ), .S0(n4207), .S1(n17), .Y(n4917) );
  MUX41X1_HVT U969 ( .A1(n4917), .A3(n4915), .A2(n4916), .A4(n4914), .S0(n4322), .S1(n4299), .Y(q[145]) );
  MUX41X1_HVT U970 ( .A1(\ram[12][146] ), .A3(\ram[14][146] ), .A2(
        \ram[13][146] ), .A4(\ram[15][146] ), .S0(n4207), .S1(n17), .Y(n4918)
         );
  MUX41X1_HVT U971 ( .A1(\ram[8][146] ), .A3(\ram[10][146] ), .A2(
        \ram[9][146] ), .A4(\ram[11][146] ), .S0(n4207), .S1(n17), .Y(n4919)
         );
  MUX41X1_HVT U972 ( .A1(\ram[4][146] ), .A3(\ram[6][146] ), .A2(\ram[5][146] ), .A4(\ram[7][146] ), .S0(n4207), .S1(n17), .Y(n4920) );
  MUX41X1_HVT U973 ( .A1(\ram[0][146] ), .A3(\ram[2][146] ), .A2(\ram[1][146] ), .A4(\ram[3][146] ), .S0(n4207), .S1(n17), .Y(n4921) );
  MUX41X1_HVT U974 ( .A1(n4921), .A3(n4919), .A2(n4920), .A4(n4918), .S0(n4322), .S1(n4299), .Y(q[146]) );
  MUX41X1_HVT U975 ( .A1(\ram[12][147] ), .A3(\ram[14][147] ), .A2(
        \ram[13][147] ), .A4(\ram[15][147] ), .S0(n4208), .S1(n18), .Y(n4922)
         );
  MUX41X1_HVT U976 ( .A1(\ram[8][147] ), .A3(\ram[10][147] ), .A2(
        \ram[9][147] ), .A4(\ram[11][147] ), .S0(n4208), .S1(n18), .Y(n4923)
         );
  MUX41X1_HVT U977 ( .A1(\ram[4][147] ), .A3(\ram[6][147] ), .A2(\ram[5][147] ), .A4(\ram[7][147] ), .S0(n4208), .S1(n18), .Y(n4924) );
  MUX41X1_HVT U978 ( .A1(\ram[0][147] ), .A3(\ram[2][147] ), .A2(\ram[1][147] ), .A4(\ram[3][147] ), .S0(n4208), .S1(n18), .Y(n4925) );
  MUX41X1_HVT U979 ( .A1(n4925), .A3(n4923), .A2(n4924), .A4(n4922), .S0(n4322), .S1(n4299), .Y(q[147]) );
  MUX41X1_HVT U980 ( .A1(\ram[12][148] ), .A3(\ram[14][148] ), .A2(
        \ram[13][148] ), .A4(\ram[15][148] ), .S0(n4208), .S1(n18), .Y(n4926)
         );
  MUX41X1_HVT U981 ( .A1(\ram[8][148] ), .A3(\ram[10][148] ), .A2(
        \ram[9][148] ), .A4(\ram[11][148] ), .S0(n4208), .S1(n18), .Y(n4927)
         );
  MUX41X1_HVT U982 ( .A1(\ram[4][148] ), .A3(\ram[6][148] ), .A2(\ram[5][148] ), .A4(\ram[7][148] ), .S0(n4208), .S1(n18), .Y(n4928) );
  MUX41X1_HVT U983 ( .A1(\ram[0][148] ), .A3(\ram[2][148] ), .A2(\ram[1][148] ), .A4(\ram[3][148] ), .S0(n4208), .S1(n18), .Y(n4929) );
  MUX41X1_HVT U984 ( .A1(n4929), .A3(n4927), .A2(n4928), .A4(n4926), .S0(n4322), .S1(n4299), .Y(q[148]) );
  MUX41X1_HVT U985 ( .A1(\ram[12][149] ), .A3(\ram[14][149] ), .A2(
        \ram[13][149] ), .A4(\ram[15][149] ), .S0(n4208), .S1(n18), .Y(n4930)
         );
  MUX41X1_HVT U986 ( .A1(\ram[8][149] ), .A3(\ram[10][149] ), .A2(
        \ram[9][149] ), .A4(\ram[11][149] ), .S0(n4208), .S1(n18), .Y(n4931)
         );
  MUX41X1_HVT U987 ( .A1(\ram[4][149] ), .A3(\ram[6][149] ), .A2(\ram[5][149] ), .A4(\ram[7][149] ), .S0(n4208), .S1(n18), .Y(n4932) );
  MUX41X1_HVT U988 ( .A1(\ram[0][149] ), .A3(\ram[2][149] ), .A2(\ram[1][149] ), .A4(\ram[3][149] ), .S0(n4208), .S1(n18), .Y(n4933) );
  MUX41X1_HVT U989 ( .A1(n4933), .A3(n4931), .A2(n4932), .A4(n4930), .S0(n4322), .S1(n4299), .Y(q[149]) );
  MUX41X1_HVT U990 ( .A1(\ram[12][150] ), .A3(\ram[14][150] ), .A2(
        \ram[13][150] ), .A4(\ram[15][150] ), .S0(n4209), .S1(n19), .Y(n4934)
         );
  MUX41X1_HVT U991 ( .A1(\ram[8][150] ), .A3(\ram[10][150] ), .A2(
        \ram[9][150] ), .A4(\ram[11][150] ), .S0(n4209), .S1(n19), .Y(n4935)
         );
  MUX41X1_HVT U992 ( .A1(\ram[4][150] ), .A3(\ram[6][150] ), .A2(\ram[5][150] ), .A4(\ram[7][150] ), .S0(n4209), .S1(n19), .Y(n4936) );
  MUX41X1_HVT U993 ( .A1(\ram[0][150] ), .A3(\ram[2][150] ), .A2(\ram[1][150] ), .A4(\ram[3][150] ), .S0(n4209), .S1(n19), .Y(n4937) );
  MUX41X1_HVT U994 ( .A1(n4937), .A3(n4935), .A2(n4936), .A4(n4934), .S0(n4322), .S1(n4299), .Y(q[150]) );
  MUX41X1_HVT U995 ( .A1(\ram[12][151] ), .A3(\ram[14][151] ), .A2(
        \ram[13][151] ), .A4(\ram[15][151] ), .S0(n4209), .S1(n19), .Y(n4938)
         );
  MUX41X1_HVT U996 ( .A1(\ram[8][151] ), .A3(\ram[10][151] ), .A2(
        \ram[9][151] ), .A4(\ram[11][151] ), .S0(n4209), .S1(n19), .Y(n4939)
         );
  MUX41X1_HVT U997 ( .A1(\ram[4][151] ), .A3(\ram[6][151] ), .A2(\ram[5][151] ), .A4(\ram[7][151] ), .S0(n4209), .S1(n19), .Y(n4940) );
  MUX41X1_HVT U998 ( .A1(\ram[0][151] ), .A3(\ram[2][151] ), .A2(\ram[1][151] ), .A4(\ram[3][151] ), .S0(n4209), .S1(n19), .Y(n4941) );
  MUX41X1_HVT U999 ( .A1(n4941), .A3(n4939), .A2(n4940), .A4(n4938), .S0(n4322), .S1(n4299), .Y(q[151]) );
  MUX41X1_HVT U1000 ( .A1(\ram[12][152] ), .A3(\ram[14][152] ), .A2(
        \ram[13][152] ), .A4(\ram[15][152] ), .S0(n4209), .S1(n19), .Y(n4942)
         );
  MUX41X1_HVT U1001 ( .A1(\ram[8][152] ), .A3(\ram[10][152] ), .A2(
        \ram[9][152] ), .A4(\ram[11][152] ), .S0(n4209), .S1(n19), .Y(n4943)
         );
  MUX41X1_HVT U1002 ( .A1(\ram[4][152] ), .A3(\ram[6][152] ), .A2(
        \ram[5][152] ), .A4(\ram[7][152] ), .S0(n4209), .S1(n19), .Y(n4944) );
  MUX41X1_HVT U1003 ( .A1(\ram[0][152] ), .A3(\ram[2][152] ), .A2(
        \ram[1][152] ), .A4(\ram[3][152] ), .S0(n4209), .S1(n19), .Y(n4945) );
  MUX41X1_HVT U1004 ( .A1(n4945), .A3(n4943), .A2(n4944), .A4(n4942), .S0(
        n4322), .S1(n4299), .Y(q[152]) );
  MUX41X1_HVT U1005 ( .A1(\ram[12][153] ), .A3(\ram[14][153] ), .A2(
        \ram[13][153] ), .A4(\ram[15][153] ), .S0(n4210), .S1(n20), .Y(n4946)
         );
  MUX41X1_HVT U1006 ( .A1(\ram[8][153] ), .A3(\ram[10][153] ), .A2(
        \ram[9][153] ), .A4(\ram[11][153] ), .S0(n4210), .S1(n20), .Y(n4947)
         );
  MUX41X1_HVT U1007 ( .A1(\ram[4][153] ), .A3(\ram[6][153] ), .A2(
        \ram[5][153] ), .A4(\ram[7][153] ), .S0(n4210), .S1(n20), .Y(n4948) );
  MUX41X1_HVT U1008 ( .A1(\ram[0][153] ), .A3(\ram[2][153] ), .A2(
        \ram[1][153] ), .A4(\ram[3][153] ), .S0(n4210), .S1(n20), .Y(n4949) );
  MUX41X1_HVT U1009 ( .A1(n4949), .A3(n4947), .A2(n4948), .A4(n4946), .S0(
        n4322), .S1(n4299), .Y(q[153]) );
  MUX41X1_HVT U1010 ( .A1(\ram[12][154] ), .A3(\ram[14][154] ), .A2(
        \ram[13][154] ), .A4(\ram[15][154] ), .S0(n4210), .S1(n20), .Y(n4950)
         );
  MUX41X1_HVT U1011 ( .A1(\ram[8][154] ), .A3(\ram[10][154] ), .A2(
        \ram[9][154] ), .A4(\ram[11][154] ), .S0(n4210), .S1(n20), .Y(n4951)
         );
  MUX41X1_HVT U1012 ( .A1(\ram[4][154] ), .A3(\ram[6][154] ), .A2(
        \ram[5][154] ), .A4(\ram[7][154] ), .S0(n4210), .S1(n20), .Y(n4952) );
  MUX41X1_HVT U1013 ( .A1(\ram[0][154] ), .A3(\ram[2][154] ), .A2(
        \ram[1][154] ), .A4(\ram[3][154] ), .S0(n4210), .S1(n20), .Y(n4953) );
  MUX41X1_HVT U1014 ( .A1(n4953), .A3(n4951), .A2(n4952), .A4(n4950), .S0(
        n4322), .S1(n4299), .Y(q[154]) );
  MUX41X1_HVT U1015 ( .A1(\ram[12][155] ), .A3(\ram[14][155] ), .A2(
        \ram[13][155] ), .A4(\ram[15][155] ), .S0(n4210), .S1(n20), .Y(n4954)
         );
  MUX41X1_HVT U1016 ( .A1(\ram[8][155] ), .A3(\ram[10][155] ), .A2(
        \ram[9][155] ), .A4(\ram[11][155] ), .S0(n4210), .S1(n20), .Y(n4955)
         );
  MUX41X1_HVT U1017 ( .A1(\ram[4][155] ), .A3(\ram[6][155] ), .A2(
        \ram[5][155] ), .A4(\ram[7][155] ), .S0(n4210), .S1(n20), .Y(n4956) );
  MUX41X1_HVT U1018 ( .A1(\ram[0][155] ), .A3(\ram[2][155] ), .A2(
        \ram[1][155] ), .A4(\ram[3][155] ), .S0(n4210), .S1(n20), .Y(n4957) );
  MUX41X1_HVT U1019 ( .A1(n4957), .A3(n4955), .A2(n4956), .A4(n4954), .S0(
        n4322), .S1(n4299), .Y(q[155]) );
  MUX41X1_HVT U1020 ( .A1(\ram[12][156] ), .A3(\ram[14][156] ), .A2(
        \ram[13][156] ), .A4(\ram[15][156] ), .S0(n4211), .S1(n21), .Y(n4958)
         );
  MUX41X1_HVT U1021 ( .A1(\ram[8][156] ), .A3(\ram[10][156] ), .A2(
        \ram[9][156] ), .A4(\ram[11][156] ), .S0(n4211), .S1(n21), .Y(n4959)
         );
  MUX41X1_HVT U1022 ( .A1(\ram[4][156] ), .A3(\ram[6][156] ), .A2(
        \ram[5][156] ), .A4(\ram[7][156] ), .S0(n4211), .S1(n21), .Y(n4960) );
  MUX41X1_HVT U1023 ( .A1(\ram[0][156] ), .A3(\ram[2][156] ), .A2(
        \ram[1][156] ), .A4(\ram[3][156] ), .S0(n4211), .S1(n21), .Y(n4961) );
  MUX41X1_HVT U1024 ( .A1(n4961), .A3(n4959), .A2(n4960), .A4(n4958), .S0(
        n4323), .S1(n4300), .Y(q[156]) );
  MUX41X1_HVT U1025 ( .A1(\ram[12][157] ), .A3(\ram[14][157] ), .A2(
        \ram[13][157] ), .A4(\ram[15][157] ), .S0(n4211), .S1(n21), .Y(n4962)
         );
  MUX41X1_HVT U1026 ( .A1(\ram[8][157] ), .A3(\ram[10][157] ), .A2(
        \ram[9][157] ), .A4(\ram[11][157] ), .S0(n4211), .S1(n21), .Y(n4963)
         );
  MUX41X1_HVT U1027 ( .A1(\ram[4][157] ), .A3(\ram[6][157] ), .A2(
        \ram[5][157] ), .A4(\ram[7][157] ), .S0(n4211), .S1(n21), .Y(n4964) );
  MUX41X1_HVT U1028 ( .A1(\ram[0][157] ), .A3(\ram[2][157] ), .A2(
        \ram[1][157] ), .A4(\ram[3][157] ), .S0(n4211), .S1(n21), .Y(n4965) );
  MUX41X1_HVT U1029 ( .A1(n4965), .A3(n4963), .A2(n4964), .A4(n4962), .S0(
        n4323), .S1(n4300), .Y(q[157]) );
  MUX41X1_HVT U1030 ( .A1(\ram[12][158] ), .A3(\ram[14][158] ), .A2(
        \ram[13][158] ), .A4(\ram[15][158] ), .S0(n4211), .S1(n21), .Y(n4966)
         );
  MUX41X1_HVT U1031 ( .A1(\ram[8][158] ), .A3(\ram[10][158] ), .A2(
        \ram[9][158] ), .A4(\ram[11][158] ), .S0(n4211), .S1(n21), .Y(n4967)
         );
  MUX41X1_HVT U1032 ( .A1(\ram[4][158] ), .A3(\ram[6][158] ), .A2(
        \ram[5][158] ), .A4(\ram[7][158] ), .S0(n4211), .S1(n21), .Y(n4968) );
  MUX41X1_HVT U1033 ( .A1(\ram[0][158] ), .A3(\ram[2][158] ), .A2(
        \ram[1][158] ), .A4(\ram[3][158] ), .S0(n4211), .S1(n21), .Y(n4969) );
  MUX41X1_HVT U1034 ( .A1(n4969), .A3(n4967), .A2(n4968), .A4(n4966), .S0(
        n4323), .S1(n4300), .Y(q[158]) );
  MUX41X1_HVT U1035 ( .A1(\ram[12][159] ), .A3(\ram[14][159] ), .A2(
        \ram[13][159] ), .A4(\ram[15][159] ), .S0(n4212), .S1(n22), .Y(n4970)
         );
  MUX41X1_HVT U1036 ( .A1(\ram[8][159] ), .A3(\ram[10][159] ), .A2(
        \ram[9][159] ), .A4(\ram[11][159] ), .S0(n4212), .S1(n22), .Y(n4971)
         );
  MUX41X1_HVT U1037 ( .A1(\ram[4][159] ), .A3(\ram[6][159] ), .A2(
        \ram[5][159] ), .A4(\ram[7][159] ), .S0(n4212), .S1(n22), .Y(n4972) );
  MUX41X1_HVT U1038 ( .A1(\ram[0][159] ), .A3(\ram[2][159] ), .A2(
        \ram[1][159] ), .A4(\ram[3][159] ), .S0(n4212), .S1(n22), .Y(n4973) );
  MUX41X1_HVT U1039 ( .A1(n4973), .A3(n4971), .A2(n4972), .A4(n4970), .S0(
        n4323), .S1(n4300), .Y(q[159]) );
  MUX41X1_HVT U1040 ( .A1(\ram[12][160] ), .A3(\ram[14][160] ), .A2(
        \ram[13][160] ), .A4(\ram[15][160] ), .S0(n4196), .S1(n6), .Y(n4974)
         );
  MUX41X1_HVT U1041 ( .A1(\ram[8][160] ), .A3(\ram[10][160] ), .A2(
        \ram[9][160] ), .A4(\ram[11][160] ), .S0(n4191), .S1(n1), .Y(n4975) );
  MUX41X1_HVT U1042 ( .A1(\ram[4][160] ), .A3(\ram[6][160] ), .A2(
        \ram[5][160] ), .A4(\ram[7][160] ), .S0(n4191), .S1(n1), .Y(n4976) );
  MUX41X1_HVT U1043 ( .A1(\ram[0][160] ), .A3(\ram[2][160] ), .A2(
        \ram[1][160] ), .A4(\ram[3][160] ), .S0(n4191), .S1(n1), .Y(n4977) );
  MUX41X1_HVT U1044 ( .A1(n4977), .A3(n4975), .A2(n4976), .A4(n4974), .S0(
        n4323), .S1(n4300), .Y(q[160]) );
  MUX41X1_HVT U1045 ( .A1(\ram[12][161] ), .A3(\ram[14][161] ), .A2(
        \ram[13][161] ), .A4(\ram[15][161] ), .S0(n4191), .S1(n1), .Y(n4978)
         );
  MUX41X1_HVT U1046 ( .A1(\ram[8][161] ), .A3(\ram[10][161] ), .A2(
        \ram[9][161] ), .A4(\ram[11][161] ), .S0(n4191), .S1(n1), .Y(n4979) );
  MUX41X1_HVT U1047 ( .A1(\ram[4][161] ), .A3(\ram[6][161] ), .A2(
        \ram[5][161] ), .A4(\ram[7][161] ), .S0(n4191), .S1(n1), .Y(n4980) );
  MUX41X1_HVT U1048 ( .A1(\ram[0][161] ), .A3(\ram[2][161] ), .A2(
        \ram[1][161] ), .A4(\ram[3][161] ), .S0(n4191), .S1(n1), .Y(n4981) );
  MUX41X1_HVT U1049 ( .A1(n4981), .A3(n4979), .A2(n4980), .A4(n4978), .S0(
        n4323), .S1(n4300), .Y(q[161]) );
  MUX41X1_HVT U1050 ( .A1(\ram[12][162] ), .A3(\ram[14][162] ), .A2(
        \ram[13][162] ), .A4(\ram[15][162] ), .S0(n4191), .S1(n1), .Y(n4982)
         );
  MUX41X1_HVT U1051 ( .A1(\ram[8][162] ), .A3(\ram[10][162] ), .A2(
        \ram[9][162] ), .A4(\ram[11][162] ), .S0(n4191), .S1(n1), .Y(n4983) );
  MUX41X1_HVT U1052 ( .A1(\ram[4][162] ), .A3(\ram[6][162] ), .A2(
        \ram[5][162] ), .A4(\ram[7][162] ), .S0(n4191), .S1(n1), .Y(n4984) );
  MUX41X1_HVT U1053 ( .A1(\ram[0][162] ), .A3(\ram[2][162] ), .A2(
        \ram[1][162] ), .A4(\ram[3][162] ), .S0(n4191), .S1(n1), .Y(n4985) );
  MUX41X1_HVT U1054 ( .A1(n4985), .A3(n4983), .A2(n4984), .A4(n4982), .S0(
        n4323), .S1(n4300), .Y(q[162]) );
  MUX41X1_HVT U1055 ( .A1(\ram[12][163] ), .A3(\ram[14][163] ), .A2(
        \ram[13][163] ), .A4(\ram[15][163] ), .S0(n4192), .S1(n2), .Y(n4986)
         );
  MUX41X1_HVT U1056 ( .A1(\ram[8][163] ), .A3(\ram[10][163] ), .A2(
        \ram[9][163] ), .A4(\ram[11][163] ), .S0(n4192), .S1(n2), .Y(n4987) );
  MUX41X1_HVT U1057 ( .A1(\ram[4][163] ), .A3(\ram[6][163] ), .A2(
        \ram[5][163] ), .A4(\ram[7][163] ), .S0(n4192), .S1(n2), .Y(n4988) );
  MUX41X1_HVT U1058 ( .A1(\ram[0][163] ), .A3(\ram[2][163] ), .A2(
        \ram[1][163] ), .A4(\ram[3][163] ), .S0(n4192), .S1(n2), .Y(n4989) );
  MUX41X1_HVT U1059 ( .A1(n4989), .A3(n4987), .A2(n4988), .A4(n4986), .S0(
        n4323), .S1(n4300), .Y(q[163]) );
  MUX41X1_HVT U1060 ( .A1(\ram[12][164] ), .A3(\ram[14][164] ), .A2(
        \ram[13][164] ), .A4(\ram[15][164] ), .S0(n4192), .S1(n2), .Y(n4990)
         );
  MUX41X1_HVT U1061 ( .A1(\ram[8][164] ), .A3(\ram[10][164] ), .A2(
        \ram[9][164] ), .A4(\ram[11][164] ), .S0(n4192), .S1(n2), .Y(n4991) );
  MUX41X1_HVT U1062 ( .A1(\ram[4][164] ), .A3(\ram[6][164] ), .A2(
        \ram[5][164] ), .A4(\ram[7][164] ), .S0(n4192), .S1(n2), .Y(n4992) );
  MUX41X1_HVT U1063 ( .A1(\ram[0][164] ), .A3(\ram[2][164] ), .A2(
        \ram[1][164] ), .A4(\ram[3][164] ), .S0(n4192), .S1(n2), .Y(n4993) );
  MUX41X1_HVT U1064 ( .A1(n4993), .A3(n4991), .A2(n4992), .A4(n4990), .S0(
        n4323), .S1(n4300), .Y(q[164]) );
  MUX41X1_HVT U1065 ( .A1(\ram[12][165] ), .A3(\ram[14][165] ), .A2(
        \ram[13][165] ), .A4(\ram[15][165] ), .S0(n4192), .S1(n2), .Y(n4994)
         );
  MUX41X1_HVT U1066 ( .A1(\ram[8][165] ), .A3(\ram[10][165] ), .A2(
        \ram[9][165] ), .A4(\ram[11][165] ), .S0(n4192), .S1(n2), .Y(n4995) );
  MUX41X1_HVT U1067 ( .A1(\ram[4][165] ), .A3(\ram[6][165] ), .A2(
        \ram[5][165] ), .A4(\ram[7][165] ), .S0(n4192), .S1(n2), .Y(n4996) );
  MUX41X1_HVT U1068 ( .A1(\ram[0][165] ), .A3(\ram[2][165] ), .A2(
        \ram[1][165] ), .A4(\ram[3][165] ), .S0(n4192), .S1(n2), .Y(n4997) );
  MUX41X1_HVT U1069 ( .A1(n4997), .A3(n4995), .A2(n4996), .A4(n4994), .S0(
        n4323), .S1(n4300), .Y(q[165]) );
  MUX41X1_HVT U1070 ( .A1(\ram[12][166] ), .A3(\ram[14][166] ), .A2(
        \ram[13][166] ), .A4(\ram[15][166] ), .S0(n4193), .S1(n3), .Y(n4998)
         );
  MUX41X1_HVT U1071 ( .A1(\ram[8][166] ), .A3(\ram[10][166] ), .A2(
        \ram[9][166] ), .A4(\ram[11][166] ), .S0(n4193), .S1(n3), .Y(n4999) );
  MUX41X1_HVT U1072 ( .A1(\ram[4][166] ), .A3(\ram[6][166] ), .A2(
        \ram[5][166] ), .A4(\ram[7][166] ), .S0(n4193), .S1(n3), .Y(n5000) );
  MUX41X1_HVT U1073 ( .A1(\ram[0][166] ), .A3(\ram[2][166] ), .A2(
        \ram[1][166] ), .A4(\ram[3][166] ), .S0(n4193), .S1(n3), .Y(n5001) );
  MUX41X1_HVT U1074 ( .A1(n5001), .A3(n4999), .A2(n5000), .A4(n4998), .S0(
        n4323), .S1(n4300), .Y(q[166]) );
  MUX41X1_HVT U1075 ( .A1(\ram[12][167] ), .A3(\ram[14][167] ), .A2(
        \ram[13][167] ), .A4(\ram[15][167] ), .S0(n4193), .S1(n3), .Y(n5002)
         );
  MUX41X1_HVT U1076 ( .A1(\ram[8][167] ), .A3(\ram[10][167] ), .A2(
        \ram[9][167] ), .A4(\ram[11][167] ), .S0(n4193), .S1(n3), .Y(n5003) );
  MUX41X1_HVT U1077 ( .A1(\ram[4][167] ), .A3(\ram[6][167] ), .A2(
        \ram[5][167] ), .A4(\ram[7][167] ), .S0(n4193), .S1(n3), .Y(n5004) );
  MUX41X1_HVT U1078 ( .A1(\ram[0][167] ), .A3(\ram[2][167] ), .A2(
        \ram[1][167] ), .A4(\ram[3][167] ), .S0(n4193), .S1(n3), .Y(n5005) );
  MUX41X1_HVT U1079 ( .A1(n5005), .A3(n5003), .A2(n5004), .A4(n5002), .S0(
        n4323), .S1(n4300), .Y(q[167]) );
  MUX41X1_HVT U1080 ( .A1(\ram[12][168] ), .A3(\ram[14][168] ), .A2(
        \ram[13][168] ), .A4(\ram[15][168] ), .S0(n4193), .S1(n3), .Y(n5006)
         );
  MUX41X1_HVT U1081 ( .A1(\ram[8][168] ), .A3(\ram[10][168] ), .A2(
        \ram[9][168] ), .A4(\ram[11][168] ), .S0(n4193), .S1(n3), .Y(n5007) );
  MUX41X1_HVT U1082 ( .A1(\ram[4][168] ), .A3(\ram[6][168] ), .A2(
        \ram[5][168] ), .A4(\ram[7][168] ), .S0(n4193), .S1(n3), .Y(n5008) );
  MUX41X1_HVT U1083 ( .A1(\ram[0][168] ), .A3(\ram[2][168] ), .A2(
        \ram[1][168] ), .A4(\ram[3][168] ), .S0(n4193), .S1(n3), .Y(n5009) );
  MUX41X1_HVT U1084 ( .A1(n5009), .A3(n5007), .A2(n5008), .A4(n5006), .S0(
        n4324), .S1(n4301), .Y(q[168]) );
  MUX41X1_HVT U1085 ( .A1(\ram[12][169] ), .A3(\ram[14][169] ), .A2(
        \ram[13][169] ), .A4(\ram[15][169] ), .S0(n4194), .S1(n4), .Y(n5010)
         );
  MUX41X1_HVT U1086 ( .A1(\ram[8][169] ), .A3(\ram[10][169] ), .A2(
        \ram[9][169] ), .A4(\ram[11][169] ), .S0(n4194), .S1(n4), .Y(n5011) );
  MUX41X1_HVT U1087 ( .A1(\ram[4][169] ), .A3(\ram[6][169] ), .A2(
        \ram[5][169] ), .A4(\ram[7][169] ), .S0(n4194), .S1(n4), .Y(n5012) );
  MUX41X1_HVT U1088 ( .A1(\ram[0][169] ), .A3(\ram[2][169] ), .A2(
        \ram[1][169] ), .A4(\ram[3][169] ), .S0(n4194), .S1(n4), .Y(n5013) );
  MUX41X1_HVT U1089 ( .A1(n5013), .A3(n5011), .A2(n5012), .A4(n5010), .S0(
        n4324), .S1(n4301), .Y(q[169]) );
  MUX41X1_HVT U1090 ( .A1(\ram[12][170] ), .A3(\ram[14][170] ), .A2(
        \ram[13][170] ), .A4(\ram[15][170] ), .S0(n4194), .S1(n4), .Y(n5014)
         );
  MUX41X1_HVT U1091 ( .A1(\ram[8][170] ), .A3(\ram[10][170] ), .A2(
        \ram[9][170] ), .A4(\ram[11][170] ), .S0(n4194), .S1(n4), .Y(n5015) );
  MUX41X1_HVT U1092 ( .A1(\ram[4][170] ), .A3(\ram[6][170] ), .A2(
        \ram[5][170] ), .A4(\ram[7][170] ), .S0(n4194), .S1(n4), .Y(n5016) );
  MUX41X1_HVT U1093 ( .A1(\ram[0][170] ), .A3(\ram[2][170] ), .A2(
        \ram[1][170] ), .A4(\ram[3][170] ), .S0(n4194), .S1(n4), .Y(n5017) );
  MUX41X1_HVT U1094 ( .A1(n5017), .A3(n5015), .A2(n5016), .A4(n5014), .S0(
        n4324), .S1(n4301), .Y(q[170]) );
  MUX41X1_HVT U1095 ( .A1(\ram[12][171] ), .A3(\ram[14][171] ), .A2(
        \ram[13][171] ), .A4(\ram[15][171] ), .S0(n4194), .S1(n4), .Y(n5018)
         );
  MUX41X1_HVT U1096 ( .A1(\ram[8][171] ), .A3(\ram[10][171] ), .A2(
        \ram[9][171] ), .A4(\ram[11][171] ), .S0(n4194), .S1(n4), .Y(n5019) );
  MUX41X1_HVT U1097 ( .A1(\ram[4][171] ), .A3(\ram[6][171] ), .A2(
        \ram[5][171] ), .A4(\ram[7][171] ), .S0(n4194), .S1(n4), .Y(n5020) );
  MUX41X1_HVT U1098 ( .A1(\ram[0][171] ), .A3(\ram[2][171] ), .A2(
        \ram[1][171] ), .A4(\ram[3][171] ), .S0(n4194), .S1(n4), .Y(n5021) );
  MUX41X1_HVT U1099 ( .A1(n5021), .A3(n5019), .A2(n5020), .A4(n5018), .S0(
        n4324), .S1(n4301), .Y(q[171]) );
  MUX41X1_HVT U1100 ( .A1(\ram[12][172] ), .A3(\ram[14][172] ), .A2(
        \ram[13][172] ), .A4(\ram[15][172] ), .S0(n4195), .S1(n5), .Y(n5022)
         );
  MUX41X1_HVT U1101 ( .A1(\ram[8][172] ), .A3(\ram[10][172] ), .A2(
        \ram[9][172] ), .A4(\ram[11][172] ), .S0(n4195), .S1(n5), .Y(n5023) );
  MUX41X1_HVT U1102 ( .A1(\ram[4][172] ), .A3(\ram[6][172] ), .A2(
        \ram[5][172] ), .A4(\ram[7][172] ), .S0(n4195), .S1(n5), .Y(n5024) );
  MUX41X1_HVT U1103 ( .A1(\ram[0][172] ), .A3(\ram[2][172] ), .A2(
        \ram[1][172] ), .A4(\ram[3][172] ), .S0(n4195), .S1(n5), .Y(n5025) );
  MUX41X1_HVT U1104 ( .A1(n5025), .A3(n5023), .A2(n5024), .A4(n5022), .S0(
        n4324), .S1(n4301), .Y(q[172]) );
  MUX41X1_HVT U1105 ( .A1(\ram[12][173] ), .A3(\ram[14][173] ), .A2(
        \ram[13][173] ), .A4(\ram[15][173] ), .S0(n4195), .S1(n5), .Y(n5026)
         );
  MUX41X1_HVT U1106 ( .A1(\ram[8][173] ), .A3(\ram[10][173] ), .A2(
        \ram[9][173] ), .A4(\ram[11][173] ), .S0(n4195), .S1(n5), .Y(n5027) );
  MUX41X1_HVT U1107 ( .A1(\ram[4][173] ), .A3(\ram[6][173] ), .A2(
        \ram[5][173] ), .A4(\ram[7][173] ), .S0(n4195), .S1(n5), .Y(n5028) );
  MUX41X1_HVT U1108 ( .A1(\ram[0][173] ), .A3(\ram[2][173] ), .A2(
        \ram[1][173] ), .A4(\ram[3][173] ), .S0(n4195), .S1(n5), .Y(n5029) );
  MUX41X1_HVT U1109 ( .A1(n5029), .A3(n5027), .A2(n5028), .A4(n5026), .S0(
        n4324), .S1(n4301), .Y(q[173]) );
  MUX41X1_HVT U1110 ( .A1(\ram[12][174] ), .A3(\ram[14][174] ), .A2(
        \ram[13][174] ), .A4(\ram[15][174] ), .S0(n4195), .S1(n5), .Y(n5030)
         );
  MUX41X1_HVT U1111 ( .A1(\ram[8][174] ), .A3(\ram[10][174] ), .A2(
        \ram[9][174] ), .A4(\ram[11][174] ), .S0(n4195), .S1(n5), .Y(n5031) );
  MUX41X1_HVT U1112 ( .A1(\ram[4][174] ), .A3(\ram[6][174] ), .A2(
        \ram[5][174] ), .A4(\ram[7][174] ), .S0(n4195), .S1(n5), .Y(n5032) );
  MUX41X1_HVT U1113 ( .A1(\ram[0][174] ), .A3(\ram[2][174] ), .A2(
        \ram[1][174] ), .A4(\ram[3][174] ), .S0(n4195), .S1(n5), .Y(n5033) );
  MUX41X1_HVT U1114 ( .A1(n5033), .A3(n5031), .A2(n5032), .A4(n5030), .S0(
        n4324), .S1(n4301), .Y(q[174]) );
  MUX41X1_HVT U1115 ( .A1(\ram[12][175] ), .A3(\ram[14][175] ), .A2(
        \ram[13][175] ), .A4(\ram[15][175] ), .S0(n4196), .S1(n6), .Y(n5034)
         );
  MUX41X1_HVT U1116 ( .A1(\ram[8][175] ), .A3(\ram[10][175] ), .A2(
        \ram[9][175] ), .A4(\ram[11][175] ), .S0(n4196), .S1(n6), .Y(n5035) );
  MUX41X1_HVT U1117 ( .A1(\ram[4][175] ), .A3(\ram[6][175] ), .A2(
        \ram[5][175] ), .A4(\ram[7][175] ), .S0(n4196), .S1(n6), .Y(n5036) );
  MUX41X1_HVT U1118 ( .A1(\ram[0][175] ), .A3(\ram[2][175] ), .A2(
        \ram[1][175] ), .A4(\ram[3][175] ), .S0(n4196), .S1(n6), .Y(n5037) );
  MUX41X1_HVT U1119 ( .A1(n5037), .A3(n5035), .A2(n5036), .A4(n5034), .S0(
        n4324), .S1(n4301), .Y(q[175]) );
  MUX41X1_HVT U1120 ( .A1(\ram[12][176] ), .A3(\ram[14][176] ), .A2(
        \ram[13][176] ), .A4(\ram[15][176] ), .S0(n4196), .S1(n6), .Y(n5038)
         );
  MUX41X1_HVT U1121 ( .A1(\ram[8][176] ), .A3(\ram[10][176] ), .A2(
        \ram[9][176] ), .A4(\ram[11][176] ), .S0(n4196), .S1(n6), .Y(n5039) );
  MUX41X1_HVT U1122 ( .A1(\ram[4][176] ), .A3(\ram[6][176] ), .A2(
        \ram[5][176] ), .A4(\ram[7][176] ), .S0(n4196), .S1(n6), .Y(n5040) );
  MUX41X1_HVT U1123 ( .A1(\ram[0][176] ), .A3(\ram[2][176] ), .A2(
        \ram[1][176] ), .A4(\ram[3][176] ), .S0(n4196), .S1(n6), .Y(n5041) );
  MUX41X1_HVT U1124 ( .A1(n5041), .A3(n5039), .A2(n5040), .A4(n5038), .S0(
        n4324), .S1(n4301), .Y(q[176]) );
  MUX41X1_HVT U1125 ( .A1(\ram[12][177] ), .A3(\ram[14][177] ), .A2(
        \ram[13][177] ), .A4(\ram[15][177] ), .S0(n4196), .S1(n6), .Y(n5042)
         );
  MUX41X1_HVT U1126 ( .A1(\ram[8][177] ), .A3(\ram[10][177] ), .A2(
        \ram[9][177] ), .A4(\ram[11][177] ), .S0(n4196), .S1(n6), .Y(n5043) );
  MUX41X1_HVT U1127 ( .A1(\ram[4][177] ), .A3(\ram[6][177] ), .A2(
        \ram[5][177] ), .A4(\ram[7][177] ), .S0(n4196), .S1(n6), .Y(n5044) );
  MUX41X1_HVT U1128 ( .A1(\ram[0][177] ), .A3(\ram[2][177] ), .A2(
        \ram[1][177] ), .A4(\ram[3][177] ), .S0(n4197), .S1(n7), .Y(n5045) );
  MUX41X1_HVT U1129 ( .A1(n5045), .A3(n5043), .A2(n5044), .A4(n5042), .S0(
        n4324), .S1(n4301), .Y(q[177]) );
  MUX41X1_HVT U1130 ( .A1(\ram[12][178] ), .A3(\ram[14][178] ), .A2(
        \ram[13][178] ), .A4(\ram[15][178] ), .S0(n4197), .S1(n7), .Y(n5046)
         );
  MUX41X1_HVT U1131 ( .A1(\ram[8][178] ), .A3(\ram[10][178] ), .A2(
        \ram[9][178] ), .A4(\ram[11][178] ), .S0(n4197), .S1(n7), .Y(n5047) );
  MUX41X1_HVT U1132 ( .A1(\ram[4][178] ), .A3(\ram[6][178] ), .A2(
        \ram[5][178] ), .A4(\ram[7][178] ), .S0(n4197), .S1(n7), .Y(n5048) );
  MUX41X1_HVT U1133 ( .A1(\ram[0][178] ), .A3(\ram[2][178] ), .A2(
        \ram[1][178] ), .A4(\ram[3][178] ), .S0(n4197), .S1(n7), .Y(n5049) );
  MUX41X1_HVT U1134 ( .A1(n5049), .A3(n5047), .A2(n5048), .A4(n5046), .S0(
        n4324), .S1(n4301), .Y(q[178]) );
  MUX41X1_HVT U1135 ( .A1(\ram[12][179] ), .A3(\ram[14][179] ), .A2(
        \ram[13][179] ), .A4(\ram[15][179] ), .S0(n4197), .S1(n7), .Y(n5050)
         );
  MUX41X1_HVT U1136 ( .A1(\ram[8][179] ), .A3(\ram[10][179] ), .A2(
        \ram[9][179] ), .A4(\ram[11][179] ), .S0(n4197), .S1(n7), .Y(n5051) );
  MUX41X1_HVT U1137 ( .A1(\ram[4][179] ), .A3(\ram[6][179] ), .A2(
        \ram[5][179] ), .A4(\ram[7][179] ), .S0(n4197), .S1(n7), .Y(n5052) );
  MUX41X1_HVT U1138 ( .A1(\ram[0][179] ), .A3(\ram[2][179] ), .A2(
        \ram[1][179] ), .A4(\ram[3][179] ), .S0(n4197), .S1(n7), .Y(n5053) );
  MUX41X1_HVT U1139 ( .A1(n5053), .A3(n5051), .A2(n5052), .A4(n5050), .S0(
        n4324), .S1(n4301), .Y(q[179]) );
  MUX41X1_HVT U1140 ( .A1(\ram[12][180] ), .A3(\ram[14][180] ), .A2(
        \ram[13][180] ), .A4(\ram[15][180] ), .S0(n4197), .S1(n7), .Y(n5054)
         );
  MUX41X1_HVT U1141 ( .A1(\ram[8][180] ), .A3(\ram[10][180] ), .A2(
        \ram[9][180] ), .A4(\ram[11][180] ), .S0(n4197), .S1(n7), .Y(n5055) );
  MUX41X1_HVT U1142 ( .A1(\ram[4][180] ), .A3(\ram[6][180] ), .A2(
        \ram[5][180] ), .A4(\ram[7][180] ), .S0(n4197), .S1(n7), .Y(n5056) );
  MUX41X1_HVT U1143 ( .A1(\ram[0][180] ), .A3(\ram[2][180] ), .A2(
        \ram[1][180] ), .A4(\ram[3][180] ), .S0(n4198), .S1(n8), .Y(n5057) );
  MUX41X1_HVT U1144 ( .A1(n5057), .A3(n5055), .A2(n5056), .A4(n5054), .S0(
        n4325), .S1(n4302), .Y(q[180]) );
  MUX41X1_HVT U1145 ( .A1(\ram[12][181] ), .A3(\ram[14][181] ), .A2(
        \ram[13][181] ), .A4(\ram[15][181] ), .S0(n4198), .S1(n8), .Y(n5058)
         );
  MUX41X1_HVT U1146 ( .A1(\ram[8][181] ), .A3(\ram[10][181] ), .A2(
        \ram[9][181] ), .A4(\ram[11][181] ), .S0(n4198), .S1(n8), .Y(n5059) );
  MUX41X1_HVT U1147 ( .A1(\ram[4][181] ), .A3(\ram[6][181] ), .A2(
        \ram[5][181] ), .A4(\ram[7][181] ), .S0(n4198), .S1(n8), .Y(n5060) );
  MUX41X1_HVT U1148 ( .A1(\ram[0][181] ), .A3(\ram[2][181] ), .A2(
        \ram[1][181] ), .A4(\ram[3][181] ), .S0(n4198), .S1(n8), .Y(n5061) );
  MUX41X1_HVT U1149 ( .A1(n5061), .A3(n5059), .A2(n5060), .A4(n5058), .S0(
        n4325), .S1(n4302), .Y(q[181]) );
  MUX41X1_HVT U1150 ( .A1(\ram[12][182] ), .A3(\ram[14][182] ), .A2(
        \ram[13][182] ), .A4(\ram[15][182] ), .S0(n4198), .S1(n8), .Y(n5062)
         );
  MUX41X1_HVT U1151 ( .A1(\ram[8][182] ), .A3(\ram[10][182] ), .A2(
        \ram[9][182] ), .A4(\ram[11][182] ), .S0(n4198), .S1(n8), .Y(n5063) );
  MUX41X1_HVT U1152 ( .A1(\ram[4][182] ), .A3(\ram[6][182] ), .A2(
        \ram[5][182] ), .A4(\ram[7][182] ), .S0(n4198), .S1(n8), .Y(n5064) );
  MUX41X1_HVT U1153 ( .A1(\ram[0][182] ), .A3(\ram[2][182] ), .A2(
        \ram[1][182] ), .A4(\ram[3][182] ), .S0(n4198), .S1(n8), .Y(n5065) );
  MUX41X1_HVT U1154 ( .A1(n5065), .A3(n5063), .A2(n5064), .A4(n5062), .S0(
        n4325), .S1(n4302), .Y(q[182]) );
  MUX41X1_HVT U1155 ( .A1(\ram[12][183] ), .A3(\ram[14][183] ), .A2(
        \ram[13][183] ), .A4(\ram[15][183] ), .S0(n4198), .S1(n8), .Y(n5066)
         );
  MUX41X1_HVT U1156 ( .A1(\ram[8][183] ), .A3(\ram[10][183] ), .A2(
        \ram[9][183] ), .A4(\ram[11][183] ), .S0(n4198), .S1(n8), .Y(n5067) );
  MUX41X1_HVT U1157 ( .A1(\ram[4][183] ), .A3(\ram[6][183] ), .A2(
        \ram[5][183] ), .A4(\ram[7][183] ), .S0(n4198), .S1(n8), .Y(n5068) );
  MUX41X1_HVT U1158 ( .A1(\ram[0][183] ), .A3(\ram[2][183] ), .A2(
        \ram[1][183] ), .A4(\ram[3][183] ), .S0(n4199), .S1(n9), .Y(n5069) );
  MUX41X1_HVT U1159 ( .A1(n5069), .A3(n5067), .A2(n5068), .A4(n5066), .S0(
        n4325), .S1(n4302), .Y(q[183]) );
  MUX41X1_HVT U1160 ( .A1(\ram[12][184] ), .A3(\ram[14][184] ), .A2(
        \ram[13][184] ), .A4(\ram[15][184] ), .S0(n4199), .S1(n9), .Y(n5070)
         );
  MUX41X1_HVT U1161 ( .A1(\ram[8][184] ), .A3(\ram[10][184] ), .A2(
        \ram[9][184] ), .A4(\ram[11][184] ), .S0(n4199), .S1(n9), .Y(n5071) );
  MUX41X1_HVT U1162 ( .A1(\ram[4][184] ), .A3(\ram[6][184] ), .A2(
        \ram[5][184] ), .A4(\ram[7][184] ), .S0(n4199), .S1(n9), .Y(n5072) );
  MUX41X1_HVT U1163 ( .A1(\ram[0][184] ), .A3(\ram[2][184] ), .A2(
        \ram[1][184] ), .A4(\ram[3][184] ), .S0(n4199), .S1(n9), .Y(n5073) );
  MUX41X1_HVT U1164 ( .A1(n5073), .A3(n5071), .A2(n5072), .A4(n5070), .S0(
        n4325), .S1(n4302), .Y(q[184]) );
  MUX41X1_HVT U1165 ( .A1(\ram[12][185] ), .A3(\ram[14][185] ), .A2(
        \ram[13][185] ), .A4(\ram[15][185] ), .S0(n4199), .S1(n9), .Y(n5074)
         );
  MUX41X1_HVT U1166 ( .A1(\ram[8][185] ), .A3(\ram[10][185] ), .A2(
        \ram[9][185] ), .A4(\ram[11][185] ), .S0(n4199), .S1(n9), .Y(n5075) );
  MUX41X1_HVT U1167 ( .A1(\ram[4][185] ), .A3(\ram[6][185] ), .A2(
        \ram[5][185] ), .A4(\ram[7][185] ), .S0(n4199), .S1(n9), .Y(n5076) );
  MUX41X1_HVT U1168 ( .A1(\ram[0][185] ), .A3(\ram[2][185] ), .A2(
        \ram[1][185] ), .A4(\ram[3][185] ), .S0(n4199), .S1(n9), .Y(n5077) );
  MUX41X1_HVT U1169 ( .A1(n5077), .A3(n5075), .A2(n5076), .A4(n5074), .S0(
        n4325), .S1(n4302), .Y(q[185]) );
  MUX41X1_HVT U1170 ( .A1(\ram[12][186] ), .A3(\ram[14][186] ), .A2(
        \ram[13][186] ), .A4(\ram[15][186] ), .S0(n4199), .S1(n9), .Y(n5078)
         );
  MUX41X1_HVT U1171 ( .A1(\ram[8][186] ), .A3(\ram[10][186] ), .A2(
        \ram[9][186] ), .A4(\ram[11][186] ), .S0(n4199), .S1(n9), .Y(n5079) );
  MUX41X1_HVT U1172 ( .A1(\ram[4][186] ), .A3(\ram[6][186] ), .A2(
        \ram[5][186] ), .A4(\ram[7][186] ), .S0(n4199), .S1(n9), .Y(n5080) );
  MUX41X1_HVT U1173 ( .A1(\ram[0][186] ), .A3(\ram[2][186] ), .A2(
        \ram[1][186] ), .A4(\ram[3][186] ), .S0(n4200), .S1(n10), .Y(n5081) );
  MUX41X1_HVT U1174 ( .A1(n5081), .A3(n5079), .A2(n5080), .A4(n5078), .S0(
        n4325), .S1(n4302), .Y(q[186]) );
  MUX41X1_HVT U1175 ( .A1(\ram[12][187] ), .A3(\ram[14][187] ), .A2(
        \ram[13][187] ), .A4(\ram[15][187] ), .S0(n4200), .S1(n10), .Y(n5082)
         );
  MUX41X1_HVT U1176 ( .A1(\ram[8][187] ), .A3(\ram[10][187] ), .A2(
        \ram[9][187] ), .A4(\ram[11][187] ), .S0(n4200), .S1(n10), .Y(n5083)
         );
  MUX41X1_HVT U1177 ( .A1(\ram[4][187] ), .A3(\ram[6][187] ), .A2(
        \ram[5][187] ), .A4(\ram[7][187] ), .S0(n4200), .S1(n10), .Y(n5084) );
  MUX41X1_HVT U1178 ( .A1(\ram[0][187] ), .A3(\ram[2][187] ), .A2(
        \ram[1][187] ), .A4(\ram[3][187] ), .S0(n4200), .S1(n10), .Y(n5085) );
  MUX41X1_HVT U1179 ( .A1(n5085), .A3(n5083), .A2(n5084), .A4(n5082), .S0(
        n4325), .S1(n4302), .Y(q[187]) );
  MUX41X1_HVT U1180 ( .A1(\ram[12][188] ), .A3(\ram[14][188] ), .A2(
        \ram[13][188] ), .A4(\ram[15][188] ), .S0(n4200), .S1(n10), .Y(n5086)
         );
  MUX41X1_HVT U1181 ( .A1(\ram[8][188] ), .A3(\ram[10][188] ), .A2(
        \ram[9][188] ), .A4(\ram[11][188] ), .S0(n4200), .S1(n10), .Y(n5087)
         );
  MUX41X1_HVT U1182 ( .A1(\ram[4][188] ), .A3(\ram[6][188] ), .A2(
        \ram[5][188] ), .A4(\ram[7][188] ), .S0(n4200), .S1(n10), .Y(n5088) );
  MUX41X1_HVT U1183 ( .A1(\ram[0][188] ), .A3(\ram[2][188] ), .A2(
        \ram[1][188] ), .A4(\ram[3][188] ), .S0(n4200), .S1(n10), .Y(n5089) );
  MUX41X1_HVT U1184 ( .A1(n5089), .A3(n5087), .A2(n5088), .A4(n5086), .S0(
        n4325), .S1(n4302), .Y(q[188]) );
  MUX41X1_HVT U1185 ( .A1(\ram[12][189] ), .A3(\ram[14][189] ), .A2(
        \ram[13][189] ), .A4(\ram[15][189] ), .S0(n4200), .S1(n10), .Y(n5090)
         );
  MUX41X1_HVT U1186 ( .A1(\ram[8][189] ), .A3(\ram[10][189] ), .A2(
        \ram[9][189] ), .A4(\ram[11][189] ), .S0(n4200), .S1(n10), .Y(n5091)
         );
  MUX41X1_HVT U1187 ( .A1(\ram[4][189] ), .A3(\ram[6][189] ), .A2(
        \ram[5][189] ), .A4(\ram[7][189] ), .S0(n4200), .S1(n10), .Y(n5092) );
  MUX41X1_HVT U1188 ( .A1(\ram[0][189] ), .A3(\ram[2][189] ), .A2(
        \ram[1][189] ), .A4(\ram[3][189] ), .S0(n4201), .S1(n11), .Y(n5093) );
  MUX41X1_HVT U1189 ( .A1(n5093), .A3(n5091), .A2(n5092), .A4(n5090), .S0(
        n4325), .S1(n4302), .Y(q[189]) );
  MUX41X1_HVT U1190 ( .A1(\ram[12][190] ), .A3(\ram[14][190] ), .A2(
        \ram[13][190] ), .A4(\ram[15][190] ), .S0(n4201), .S1(n11), .Y(n5094)
         );
  MUX41X1_HVT U1191 ( .A1(\ram[8][190] ), .A3(\ram[10][190] ), .A2(
        \ram[9][190] ), .A4(\ram[11][190] ), .S0(n4201), .S1(n11), .Y(n5095)
         );
  MUX41X1_HVT U1192 ( .A1(\ram[4][190] ), .A3(\ram[6][190] ), .A2(
        \ram[5][190] ), .A4(\ram[7][190] ), .S0(n4201), .S1(n11), .Y(n5096) );
  MUX41X1_HVT U1193 ( .A1(\ram[0][190] ), .A3(\ram[2][190] ), .A2(
        \ram[1][190] ), .A4(\ram[3][190] ), .S0(n4201), .S1(n11), .Y(n5097) );
  MUX41X1_HVT U1194 ( .A1(n5097), .A3(n5095), .A2(n5096), .A4(n5094), .S0(
        n4325), .S1(n4302), .Y(q[190]) );
  MUX41X1_HVT U1195 ( .A1(\ram[12][191] ), .A3(\ram[14][191] ), .A2(
        \ram[13][191] ), .A4(\ram[15][191] ), .S0(n4201), .S1(n11), .Y(n5098)
         );
  MUX41X1_HVT U1196 ( .A1(\ram[8][191] ), .A3(\ram[10][191] ), .A2(
        \ram[9][191] ), .A4(\ram[11][191] ), .S0(n4201), .S1(n11), .Y(n5099)
         );
  MUX41X1_HVT U1197 ( .A1(\ram[4][191] ), .A3(\ram[6][191] ), .A2(
        \ram[5][191] ), .A4(\ram[7][191] ), .S0(n4201), .S1(n11), .Y(n5100) );
  MUX41X1_HVT U1198 ( .A1(\ram[0][191] ), .A3(\ram[2][191] ), .A2(
        \ram[1][191] ), .A4(\ram[3][191] ), .S0(n4201), .S1(n11), .Y(n5101) );
  MUX41X1_HVT U1199 ( .A1(n5101), .A3(n5099), .A2(n5100), .A4(n5098), .S0(
        n4325), .S1(n4302), .Y(q[191]) );
  MUX41X1_HVT U1200 ( .A1(\ram[12][192] ), .A3(\ram[14][192] ), .A2(
        \ram[13][192] ), .A4(\ram[15][192] ), .S0(n4228), .S1(n38), .Y(n5102)
         );
  MUX41X1_HVT U1201 ( .A1(\ram[8][192] ), .A3(\ram[10][192] ), .A2(
        \ram[9][192] ), .A4(\ram[11][192] ), .S0(n4223), .S1(n33), .Y(n5103)
         );
  MUX41X1_HVT U1202 ( .A1(\ram[4][192] ), .A3(\ram[6][192] ), .A2(
        \ram[5][192] ), .A4(\ram[7][192] ), .S0(n4223), .S1(n33), .Y(n5104) );
  MUX41X1_HVT U1203 ( .A1(\ram[0][192] ), .A3(\ram[2][192] ), .A2(
        \ram[1][192] ), .A4(\ram[3][192] ), .S0(n4223), .S1(n33), .Y(n5105) );
  MUX41X1_HVT U1204 ( .A1(n5105), .A3(n5103), .A2(n5104), .A4(n5102), .S0(
        n4326), .S1(n4303), .Y(q[192]) );
  MUX41X1_HVT U1205 ( .A1(\ram[12][193] ), .A3(\ram[14][193] ), .A2(
        \ram[13][193] ), .A4(\ram[15][193] ), .S0(n4233), .S1(n33), .Y(n5106)
         );
  MUX41X1_HVT U1206 ( .A1(\ram[8][193] ), .A3(\ram[10][193] ), .A2(
        \ram[9][193] ), .A4(\ram[11][193] ), .S0(n4223), .S1(n43), .Y(n5107)
         );
  MUX41X1_HVT U1207 ( .A1(\ram[4][193] ), .A3(\ram[6][193] ), .A2(
        \ram[5][193] ), .A4(\ram[7][193] ), .S0(n4223), .S1(n33), .Y(n5108) );
  MUX41X1_HVT U1208 ( .A1(\ram[0][193] ), .A3(\ram[2][193] ), .A2(
        \ram[1][193] ), .A4(\ram[3][193] ), .S0(n4223), .S1(n33), .Y(n5109) );
  MUX41X1_HVT U1209 ( .A1(n5109), .A3(n5107), .A2(n5108), .A4(n5106), .S0(
        n4326), .S1(n4303), .Y(q[193]) );
  MUX41X1_HVT U1210 ( .A1(\ram[12][194] ), .A3(\ram[14][194] ), .A2(
        \ram[13][194] ), .A4(\ram[15][194] ), .S0(n4223), .S1(n33), .Y(n5110)
         );
  MUX41X1_HVT U1211 ( .A1(\ram[8][194] ), .A3(\ram[10][194] ), .A2(
        \ram[9][194] ), .A4(\ram[11][194] ), .S0(n4223), .S1(n33), .Y(n5111)
         );
  MUX41X1_HVT U1212 ( .A1(\ram[4][194] ), .A3(\ram[6][194] ), .A2(
        \ram[5][194] ), .A4(\ram[7][194] ), .S0(n4223), .S1(n33), .Y(n5112) );
  MUX41X1_HVT U1213 ( .A1(\ram[0][194] ), .A3(\ram[2][194] ), .A2(
        \ram[1][194] ), .A4(\ram[3][194] ), .S0(n4223), .S1(n33), .Y(n5113) );
  MUX41X1_HVT U1214 ( .A1(n5113), .A3(n5111), .A2(n5112), .A4(n5110), .S0(
        n4326), .S1(n4303), .Y(q[194]) );
  MUX41X1_HVT U1215 ( .A1(\ram[12][195] ), .A3(\ram[14][195] ), .A2(
        \ram[13][195] ), .A4(\ram[15][195] ), .S0(n4223), .S1(n33), .Y(n5114)
         );
  MUX41X1_HVT U1216 ( .A1(\ram[8][195] ), .A3(\ram[10][195] ), .A2(
        \ram[9][195] ), .A4(\ram[11][195] ), .S0(n4224), .S1(n34), .Y(n5115)
         );
  MUX41X1_HVT U1217 ( .A1(\ram[4][195] ), .A3(\ram[6][195] ), .A2(
        \ram[5][195] ), .A4(\ram[7][195] ), .S0(n4224), .S1(n34), .Y(n5116) );
  MUX41X1_HVT U1218 ( .A1(\ram[0][195] ), .A3(\ram[2][195] ), .A2(
        \ram[1][195] ), .A4(\ram[3][195] ), .S0(n4224), .S1(n34), .Y(n5117) );
  MUX41X1_HVT U1219 ( .A1(n5117), .A3(n5115), .A2(n5116), .A4(n5114), .S0(
        n4326), .S1(n4303), .Y(q[195]) );
  MUX41X1_HVT U1220 ( .A1(\ram[12][196] ), .A3(\ram[14][196] ), .A2(
        \ram[13][196] ), .A4(\ram[15][196] ), .S0(n4224), .S1(n34), .Y(n5118)
         );
  MUX41X1_HVT U1221 ( .A1(\ram[8][196] ), .A3(\ram[10][196] ), .A2(
        \ram[9][196] ), .A4(\ram[11][196] ), .S0(n4224), .S1(n34), .Y(n5119)
         );
  MUX41X1_HVT U1222 ( .A1(\ram[4][196] ), .A3(\ram[6][196] ), .A2(
        \ram[5][196] ), .A4(\ram[7][196] ), .S0(n4224), .S1(n34), .Y(n5120) );
  MUX41X1_HVT U1223 ( .A1(\ram[0][196] ), .A3(\ram[2][196] ), .A2(
        \ram[1][196] ), .A4(\ram[3][196] ), .S0(n4224), .S1(n34), .Y(n5121) );
  MUX41X1_HVT U1224 ( .A1(n5121), .A3(n5119), .A2(n5120), .A4(n5118), .S0(
        n4326), .S1(n4303), .Y(q[196]) );
  MUX41X1_HVT U1225 ( .A1(\ram[12][197] ), .A3(\ram[14][197] ), .A2(
        \ram[13][197] ), .A4(\ram[15][197] ), .S0(n4224), .S1(n34), .Y(n5122)
         );
  MUX41X1_HVT U1226 ( .A1(\ram[8][197] ), .A3(\ram[10][197] ), .A2(
        \ram[9][197] ), .A4(\ram[11][197] ), .S0(n4224), .S1(n34), .Y(n5123)
         );
  MUX41X1_HVT U1227 ( .A1(\ram[4][197] ), .A3(\ram[6][197] ), .A2(
        \ram[5][197] ), .A4(\ram[7][197] ), .S0(n4224), .S1(n34), .Y(n5124) );
  MUX41X1_HVT U1228 ( .A1(\ram[0][197] ), .A3(\ram[2][197] ), .A2(
        \ram[1][197] ), .A4(\ram[3][197] ), .S0(n4224), .S1(n34), .Y(n5125) );
  MUX41X1_HVT U1229 ( .A1(n5125), .A3(n5123), .A2(n5124), .A4(n5122), .S0(
        n4326), .S1(n4303), .Y(q[197]) );
  MUX41X1_HVT U1230 ( .A1(\ram[12][198] ), .A3(\ram[14][198] ), .A2(
        \ram[13][198] ), .A4(\ram[15][198] ), .S0(n4224), .S1(n34), .Y(n5126)
         );
  MUX41X1_HVT U1231 ( .A1(\ram[8][198] ), .A3(\ram[10][198] ), .A2(
        \ram[9][198] ), .A4(\ram[11][198] ), .S0(n4225), .S1(n35), .Y(n5127)
         );
  MUX41X1_HVT U1232 ( .A1(\ram[4][198] ), .A3(\ram[6][198] ), .A2(
        \ram[5][198] ), .A4(\ram[7][198] ), .S0(n4225), .S1(n35), .Y(n5128) );
  MUX41X1_HVT U1233 ( .A1(\ram[0][198] ), .A3(\ram[2][198] ), .A2(
        \ram[1][198] ), .A4(\ram[3][198] ), .S0(n4225), .S1(n35), .Y(n5129) );
  MUX41X1_HVT U1234 ( .A1(n5129), .A3(n5127), .A2(n5128), .A4(n5126), .S0(
        n4326), .S1(n4303), .Y(q[198]) );
  MUX41X1_HVT U1235 ( .A1(\ram[12][199] ), .A3(\ram[14][199] ), .A2(
        \ram[13][199] ), .A4(\ram[15][199] ), .S0(n4225), .S1(n35), .Y(n5130)
         );
  MUX41X1_HVT U1236 ( .A1(\ram[8][199] ), .A3(\ram[10][199] ), .A2(
        \ram[9][199] ), .A4(\ram[11][199] ), .S0(n4225), .S1(n35), .Y(n5131)
         );
  MUX41X1_HVT U1237 ( .A1(\ram[4][199] ), .A3(\ram[6][199] ), .A2(
        \ram[5][199] ), .A4(\ram[7][199] ), .S0(n4225), .S1(n35), .Y(n5132) );
  MUX41X1_HVT U1238 ( .A1(\ram[0][199] ), .A3(\ram[2][199] ), .A2(
        \ram[1][199] ), .A4(\ram[3][199] ), .S0(n4225), .S1(n35), .Y(n5133) );
  MUX41X1_HVT U1239 ( .A1(n5133), .A3(n5131), .A2(n5132), .A4(n5130), .S0(
        n4326), .S1(n4303), .Y(q[199]) );
  MUX41X1_HVT U1240 ( .A1(\ram[12][200] ), .A3(\ram[14][200] ), .A2(
        \ram[13][200] ), .A4(\ram[15][200] ), .S0(n4225), .S1(n35), .Y(n5134)
         );
  MUX41X1_HVT U1241 ( .A1(\ram[8][200] ), .A3(\ram[10][200] ), .A2(
        \ram[9][200] ), .A4(\ram[11][200] ), .S0(n4225), .S1(n35), .Y(n5135)
         );
  MUX41X1_HVT U1242 ( .A1(\ram[4][200] ), .A3(\ram[6][200] ), .A2(
        \ram[5][200] ), .A4(\ram[7][200] ), .S0(n4225), .S1(n35), .Y(n5136) );
  MUX41X1_HVT U1243 ( .A1(\ram[0][200] ), .A3(\ram[2][200] ), .A2(
        \ram[1][200] ), .A4(\ram[3][200] ), .S0(n4225), .S1(n35), .Y(n5137) );
  MUX41X1_HVT U1244 ( .A1(n5137), .A3(n5135), .A2(n5136), .A4(n5134), .S0(
        n4326), .S1(n4303), .Y(q[200]) );
  MUX41X1_HVT U1245 ( .A1(\ram[12][201] ), .A3(\ram[14][201] ), .A2(
        \ram[13][201] ), .A4(\ram[15][201] ), .S0(n4225), .S1(n35), .Y(n5138)
         );
  MUX41X1_HVT U1246 ( .A1(\ram[8][201] ), .A3(\ram[10][201] ), .A2(
        \ram[9][201] ), .A4(\ram[11][201] ), .S0(n4226), .S1(n36), .Y(n5139)
         );
  MUX41X1_HVT U1247 ( .A1(\ram[4][201] ), .A3(\ram[6][201] ), .A2(
        \ram[5][201] ), .A4(\ram[7][201] ), .S0(n4226), .S1(n36), .Y(n5140) );
  MUX41X1_HVT U1248 ( .A1(\ram[0][201] ), .A3(\ram[2][201] ), .A2(
        \ram[1][201] ), .A4(\ram[3][201] ), .S0(n4226), .S1(n36), .Y(n5141) );
  MUX41X1_HVT U1249 ( .A1(n5141), .A3(n5139), .A2(n5140), .A4(n5138), .S0(
        n4326), .S1(n4303), .Y(q[201]) );
  MUX41X1_HVT U1250 ( .A1(\ram[12][202] ), .A3(\ram[14][202] ), .A2(
        \ram[13][202] ), .A4(\ram[15][202] ), .S0(n4226), .S1(n36), .Y(n5142)
         );
  MUX41X1_HVT U1251 ( .A1(\ram[8][202] ), .A3(\ram[10][202] ), .A2(
        \ram[9][202] ), .A4(\ram[11][202] ), .S0(n4226), .S1(n36), .Y(n5143)
         );
  MUX41X1_HVT U1252 ( .A1(\ram[4][202] ), .A3(\ram[6][202] ), .A2(
        \ram[5][202] ), .A4(\ram[7][202] ), .S0(n4226), .S1(n36), .Y(n5144) );
  MUX41X1_HVT U1253 ( .A1(\ram[0][202] ), .A3(\ram[2][202] ), .A2(
        \ram[1][202] ), .A4(\ram[3][202] ), .S0(n4226), .S1(n36), .Y(n5145) );
  MUX41X1_HVT U1254 ( .A1(n5145), .A3(n5143), .A2(n5144), .A4(n5142), .S0(
        n4326), .S1(n4303), .Y(q[202]) );
  MUX41X1_HVT U1255 ( .A1(\ram[12][203] ), .A3(\ram[14][203] ), .A2(
        \ram[13][203] ), .A4(\ram[15][203] ), .S0(n4226), .S1(n36), .Y(n5146)
         );
  MUX41X1_HVT U1256 ( .A1(\ram[8][203] ), .A3(\ram[10][203] ), .A2(
        \ram[9][203] ), .A4(\ram[11][203] ), .S0(n4226), .S1(n36), .Y(n5147)
         );
  MUX41X1_HVT U1257 ( .A1(\ram[4][203] ), .A3(\ram[6][203] ), .A2(
        \ram[5][203] ), .A4(\ram[7][203] ), .S0(n4226), .S1(n36), .Y(n5148) );
  MUX41X1_HVT U1258 ( .A1(\ram[0][203] ), .A3(\ram[2][203] ), .A2(
        \ram[1][203] ), .A4(\ram[3][203] ), .S0(n4226), .S1(n36), .Y(n5149) );
  MUX41X1_HVT U1259 ( .A1(n5149), .A3(n5147), .A2(n5148), .A4(n5146), .S0(
        n4326), .S1(n4303), .Y(q[203]) );
  MUX41X1_HVT U1260 ( .A1(\ram[12][204] ), .A3(\ram[14][204] ), .A2(
        \ram[13][204] ), .A4(\ram[15][204] ), .S0(n4226), .S1(n36), .Y(n5150)
         );
  MUX41X1_HVT U1261 ( .A1(\ram[8][204] ), .A3(\ram[10][204] ), .A2(
        \ram[9][204] ), .A4(\ram[11][204] ), .S0(n4227), .S1(n37), .Y(n5151)
         );
  MUX41X1_HVT U1262 ( .A1(\ram[4][204] ), .A3(\ram[6][204] ), .A2(
        \ram[5][204] ), .A4(\ram[7][204] ), .S0(n4227), .S1(n37), .Y(n5152) );
  MUX41X1_HVT U1263 ( .A1(\ram[0][204] ), .A3(\ram[2][204] ), .A2(
        \ram[1][204] ), .A4(\ram[3][204] ), .S0(n4227), .S1(n37), .Y(n5153) );
  MUX41X1_HVT U1264 ( .A1(n5153), .A3(n5151), .A2(n5152), .A4(n5150), .S0(
        n4327), .S1(n4304), .Y(q[204]) );
  MUX41X1_HVT U1265 ( .A1(\ram[12][205] ), .A3(\ram[14][205] ), .A2(
        \ram[13][205] ), .A4(\ram[15][205] ), .S0(n4227), .S1(n37), .Y(n5154)
         );
  MUX41X1_HVT U1266 ( .A1(\ram[8][205] ), .A3(\ram[10][205] ), .A2(
        \ram[9][205] ), .A4(\ram[11][205] ), .S0(n4227), .S1(n37), .Y(n5155)
         );
  MUX41X1_HVT U1267 ( .A1(\ram[4][205] ), .A3(\ram[6][205] ), .A2(
        \ram[5][205] ), .A4(\ram[7][205] ), .S0(n4227), .S1(n37), .Y(n5156) );
  MUX41X1_HVT U1268 ( .A1(\ram[0][205] ), .A3(\ram[2][205] ), .A2(
        \ram[1][205] ), .A4(\ram[3][205] ), .S0(n4227), .S1(n37), .Y(n5157) );
  MUX41X1_HVT U1269 ( .A1(n5157), .A3(n5155), .A2(n5156), .A4(n5154), .S0(
        n4327), .S1(n4304), .Y(q[205]) );
  MUX41X1_HVT U1270 ( .A1(\ram[12][206] ), .A3(\ram[14][206] ), .A2(
        \ram[13][206] ), .A4(\ram[15][206] ), .S0(n4227), .S1(n37), .Y(n5158)
         );
  MUX41X1_HVT U1271 ( .A1(\ram[8][206] ), .A3(\ram[10][206] ), .A2(
        \ram[9][206] ), .A4(\ram[11][206] ), .S0(n4227), .S1(n37), .Y(n5159)
         );
  MUX41X1_HVT U1272 ( .A1(\ram[4][206] ), .A3(\ram[6][206] ), .A2(
        \ram[5][206] ), .A4(\ram[7][206] ), .S0(n4227), .S1(n37), .Y(n5160) );
  MUX41X1_HVT U1273 ( .A1(\ram[0][206] ), .A3(\ram[2][206] ), .A2(
        \ram[1][206] ), .A4(\ram[3][206] ), .S0(n4227), .S1(n37), .Y(n5161) );
  MUX41X1_HVT U1274 ( .A1(n5161), .A3(n5159), .A2(n5160), .A4(n5158), .S0(
        n4327), .S1(n4304), .Y(q[206]) );
  MUX41X1_HVT U1275 ( .A1(\ram[12][207] ), .A3(\ram[14][207] ), .A2(
        \ram[13][207] ), .A4(\ram[15][207] ), .S0(n4227), .S1(n37), .Y(n5162)
         );
  MUX41X1_HVT U1276 ( .A1(\ram[8][207] ), .A3(\ram[10][207] ), .A2(
        \ram[9][207] ), .A4(\ram[11][207] ), .S0(n4228), .S1(n38), .Y(n5163)
         );
  MUX41X1_HVT U1277 ( .A1(\ram[4][207] ), .A3(\ram[6][207] ), .A2(
        \ram[5][207] ), .A4(\ram[7][207] ), .S0(n4228), .S1(n38), .Y(n5164) );
  MUX41X1_HVT U1278 ( .A1(\ram[0][207] ), .A3(\ram[2][207] ), .A2(
        \ram[1][207] ), .A4(\ram[3][207] ), .S0(n4228), .S1(n38), .Y(n5165) );
  MUX41X1_HVT U1279 ( .A1(n5165), .A3(n5163), .A2(n5164), .A4(n5162), .S0(
        n4327), .S1(n4304), .Y(q[207]) );
  MUX41X1_HVT U1280 ( .A1(\ram[12][208] ), .A3(\ram[14][208] ), .A2(
        \ram[13][208] ), .A4(\ram[15][208] ), .S0(n4228), .S1(n38), .Y(n5166)
         );
  MUX41X1_HVT U1281 ( .A1(\ram[8][208] ), .A3(\ram[10][208] ), .A2(
        \ram[9][208] ), .A4(\ram[11][208] ), .S0(n4228), .S1(n38), .Y(n5167)
         );
  MUX41X1_HVT U1282 ( .A1(\ram[4][208] ), .A3(\ram[6][208] ), .A2(
        \ram[5][208] ), .A4(\ram[7][208] ), .S0(n4228), .S1(n38), .Y(n5168) );
  MUX41X1_HVT U1283 ( .A1(\ram[0][208] ), .A3(\ram[2][208] ), .A2(
        \ram[1][208] ), .A4(\ram[3][208] ), .S0(n4228), .S1(n38), .Y(n5169) );
  MUX41X1_HVT U1284 ( .A1(n5169), .A3(n5167), .A2(n5168), .A4(n5166), .S0(
        n4327), .S1(n4304), .Y(q[208]) );
  MUX41X1_HVT U1285 ( .A1(\ram[12][209] ), .A3(\ram[14][209] ), .A2(
        \ram[13][209] ), .A4(\ram[15][209] ), .S0(n4228), .S1(n38), .Y(n5170)
         );
  MUX41X1_HVT U1286 ( .A1(\ram[8][209] ), .A3(\ram[10][209] ), .A2(
        \ram[9][209] ), .A4(\ram[11][209] ), .S0(n4228), .S1(n38), .Y(n5171)
         );
  MUX41X1_HVT U1287 ( .A1(\ram[4][209] ), .A3(\ram[6][209] ), .A2(
        \ram[5][209] ), .A4(\ram[7][209] ), .S0(n4228), .S1(n38), .Y(n5172) );
  MUX41X1_HVT U1288 ( .A1(\ram[0][209] ), .A3(\ram[2][209] ), .A2(
        \ram[1][209] ), .A4(\ram[3][209] ), .S0(n4228), .S1(n38), .Y(n5173) );
  MUX41X1_HVT U1289 ( .A1(n5173), .A3(n5171), .A2(n5172), .A4(n5170), .S0(
        n4327), .S1(n4304), .Y(q[209]) );
  MUX41X1_HVT U1290 ( .A1(\ram[12][210] ), .A3(\ram[14][210] ), .A2(
        \ram[13][210] ), .A4(\ram[15][210] ), .S0(n4229), .S1(n39), .Y(n5174)
         );
  MUX41X1_HVT U1291 ( .A1(\ram[8][210] ), .A3(\ram[10][210] ), .A2(
        \ram[9][210] ), .A4(\ram[11][210] ), .S0(n4229), .S1(n39), .Y(n5175)
         );
  MUX41X1_HVT U1292 ( .A1(\ram[4][210] ), .A3(\ram[6][210] ), .A2(
        \ram[5][210] ), .A4(\ram[7][210] ), .S0(n4229), .S1(n39), .Y(n5176) );
  MUX41X1_HVT U1293 ( .A1(\ram[0][210] ), .A3(\ram[2][210] ), .A2(
        \ram[1][210] ), .A4(\ram[3][210] ), .S0(n4229), .S1(n39), .Y(n5177) );
  MUX41X1_HVT U1294 ( .A1(n5177), .A3(n5175), .A2(n5176), .A4(n5174), .S0(
        n4327), .S1(n4304), .Y(q[210]) );
  MUX41X1_HVT U1295 ( .A1(\ram[12][211] ), .A3(\ram[14][211] ), .A2(
        \ram[13][211] ), .A4(\ram[15][211] ), .S0(n4229), .S1(n39), .Y(n5178)
         );
  MUX41X1_HVT U1296 ( .A1(\ram[8][211] ), .A3(\ram[10][211] ), .A2(
        \ram[9][211] ), .A4(\ram[11][211] ), .S0(n4229), .S1(n39), .Y(n5179)
         );
  MUX41X1_HVT U1297 ( .A1(\ram[4][211] ), .A3(\ram[6][211] ), .A2(
        \ram[5][211] ), .A4(\ram[7][211] ), .S0(n4229), .S1(n39), .Y(n5180) );
  MUX41X1_HVT U1298 ( .A1(\ram[0][211] ), .A3(\ram[2][211] ), .A2(
        \ram[1][211] ), .A4(\ram[3][211] ), .S0(n4229), .S1(n39), .Y(n5181) );
  MUX41X1_HVT U1299 ( .A1(n5181), .A3(n5179), .A2(n5180), .A4(n5178), .S0(
        n4327), .S1(n4304), .Y(q[211]) );
  MUX41X1_HVT U1300 ( .A1(\ram[12][212] ), .A3(\ram[14][212] ), .A2(
        \ram[13][212] ), .A4(\ram[15][212] ), .S0(n4229), .S1(n39), .Y(n5182)
         );
  MUX41X1_HVT U1301 ( .A1(\ram[8][212] ), .A3(\ram[10][212] ), .A2(
        \ram[9][212] ), .A4(\ram[11][212] ), .S0(n4229), .S1(n39), .Y(n5183)
         );
  MUX41X1_HVT U1302 ( .A1(\ram[4][212] ), .A3(\ram[6][212] ), .A2(
        \ram[5][212] ), .A4(\ram[7][212] ), .S0(n4229), .S1(n39), .Y(n5184) );
  MUX41X1_HVT U1303 ( .A1(\ram[0][212] ), .A3(\ram[2][212] ), .A2(
        \ram[1][212] ), .A4(\ram[3][212] ), .S0(n4229), .S1(n39), .Y(n5185) );
  MUX41X1_HVT U1304 ( .A1(n5185), .A3(n5183), .A2(n5184), .A4(n5182), .S0(
        n4327), .S1(n4304), .Y(q[212]) );
  MUX41X1_HVT U1305 ( .A1(\ram[12][213] ), .A3(\ram[14][213] ), .A2(
        \ram[13][213] ), .A4(\ram[15][213] ), .S0(n4230), .S1(n40), .Y(n5186)
         );
  MUX41X1_HVT U1306 ( .A1(\ram[8][213] ), .A3(\ram[10][213] ), .A2(
        \ram[9][213] ), .A4(\ram[11][213] ), .S0(n4230), .S1(n40), .Y(n5187)
         );
  MUX41X1_HVT U1307 ( .A1(\ram[4][213] ), .A3(\ram[6][213] ), .A2(
        \ram[5][213] ), .A4(\ram[7][213] ), .S0(n4230), .S1(n40), .Y(n5188) );
  MUX41X1_HVT U1308 ( .A1(\ram[0][213] ), .A3(\ram[2][213] ), .A2(
        \ram[1][213] ), .A4(\ram[3][213] ), .S0(n4230), .S1(n40), .Y(n5189) );
  MUX41X1_HVT U1309 ( .A1(n5189), .A3(n5187), .A2(n5188), .A4(n5186), .S0(
        n4327), .S1(n4304), .Y(q[213]) );
  MUX41X1_HVT U1310 ( .A1(\ram[12][214] ), .A3(\ram[14][214] ), .A2(
        \ram[13][214] ), .A4(\ram[15][214] ), .S0(n4230), .S1(n40), .Y(n5190)
         );
  MUX41X1_HVT U1311 ( .A1(\ram[8][214] ), .A3(\ram[10][214] ), .A2(
        \ram[9][214] ), .A4(\ram[11][214] ), .S0(n4230), .S1(n40), .Y(n5191)
         );
  MUX41X1_HVT U1312 ( .A1(\ram[4][214] ), .A3(\ram[6][214] ), .A2(
        \ram[5][214] ), .A4(\ram[7][214] ), .S0(n4230), .S1(n40), .Y(n5192) );
  MUX41X1_HVT U1313 ( .A1(\ram[0][214] ), .A3(\ram[2][214] ), .A2(
        \ram[1][214] ), .A4(\ram[3][214] ), .S0(n4230), .S1(n40), .Y(n5193) );
  MUX41X1_HVT U1314 ( .A1(n5193), .A3(n5191), .A2(n5192), .A4(n5190), .S0(
        n4327), .S1(n4304), .Y(q[214]) );
  MUX41X1_HVT U1315 ( .A1(\ram[12][215] ), .A3(\ram[14][215] ), .A2(
        \ram[13][215] ), .A4(\ram[15][215] ), .S0(n4230), .S1(n40), .Y(n5194)
         );
  MUX41X1_HVT U1316 ( .A1(\ram[8][215] ), .A3(\ram[10][215] ), .A2(
        \ram[9][215] ), .A4(\ram[11][215] ), .S0(n4230), .S1(n40), .Y(n5195)
         );
  MUX41X1_HVT U1317 ( .A1(\ram[4][215] ), .A3(\ram[6][215] ), .A2(
        \ram[5][215] ), .A4(\ram[7][215] ), .S0(n4230), .S1(n40), .Y(n5196) );
  MUX41X1_HVT U1318 ( .A1(\ram[0][215] ), .A3(\ram[2][215] ), .A2(
        \ram[1][215] ), .A4(\ram[3][215] ), .S0(n4230), .S1(n40), .Y(n5197) );
  MUX41X1_HVT U1319 ( .A1(n5197), .A3(n5195), .A2(n5196), .A4(n5194), .S0(
        n4327), .S1(n4304), .Y(q[215]) );
  MUX41X1_HVT U1320 ( .A1(\ram[12][216] ), .A3(\ram[14][216] ), .A2(
        \ram[13][216] ), .A4(\ram[15][216] ), .S0(n4231), .S1(n41), .Y(n5198)
         );
  MUX41X1_HVT U1321 ( .A1(\ram[8][216] ), .A3(\ram[10][216] ), .A2(
        \ram[9][216] ), .A4(\ram[11][216] ), .S0(n4231), .S1(n41), .Y(n5199)
         );
  MUX41X1_HVT U1322 ( .A1(\ram[4][216] ), .A3(\ram[6][216] ), .A2(
        \ram[5][216] ), .A4(\ram[7][216] ), .S0(n4231), .S1(n41), .Y(n5200) );
  MUX41X1_HVT U1323 ( .A1(\ram[0][216] ), .A3(\ram[2][216] ), .A2(
        \ram[1][216] ), .A4(\ram[3][216] ), .S0(n4231), .S1(n41), .Y(n5201) );
  MUX41X1_HVT U1324 ( .A1(n5201), .A3(n5199), .A2(n5200), .A4(n5198), .S0(
        n4328), .S1(n4305), .Y(q[216]) );
  MUX41X1_HVT U1325 ( .A1(\ram[12][217] ), .A3(\ram[14][217] ), .A2(
        \ram[13][217] ), .A4(\ram[15][217] ), .S0(n4231), .S1(n41), .Y(n5202)
         );
  MUX41X1_HVT U1326 ( .A1(\ram[8][217] ), .A3(\ram[10][217] ), .A2(
        \ram[9][217] ), .A4(\ram[11][217] ), .S0(n4231), .S1(n41), .Y(n5203)
         );
  MUX41X1_HVT U1327 ( .A1(\ram[4][217] ), .A3(\ram[6][217] ), .A2(
        \ram[5][217] ), .A4(\ram[7][217] ), .S0(n4231), .S1(n41), .Y(n5204) );
  MUX41X1_HVT U1328 ( .A1(\ram[0][217] ), .A3(\ram[2][217] ), .A2(
        \ram[1][217] ), .A4(\ram[3][217] ), .S0(n4231), .S1(n41), .Y(n5205) );
  MUX41X1_HVT U1329 ( .A1(n5205), .A3(n5203), .A2(n5204), .A4(n5202), .S0(
        n4328), .S1(n4305), .Y(q[217]) );
  MUX41X1_HVT U1330 ( .A1(\ram[12][218] ), .A3(\ram[14][218] ), .A2(
        \ram[13][218] ), .A4(\ram[15][218] ), .S0(n4231), .S1(n41), .Y(n5206)
         );
  MUX41X1_HVT U1331 ( .A1(\ram[8][218] ), .A3(\ram[10][218] ), .A2(
        \ram[9][218] ), .A4(\ram[11][218] ), .S0(n4231), .S1(n41), .Y(n5207)
         );
  MUX41X1_HVT U1332 ( .A1(\ram[4][218] ), .A3(\ram[6][218] ), .A2(
        \ram[5][218] ), .A4(\ram[7][218] ), .S0(n4231), .S1(n41), .Y(n5208) );
  MUX41X1_HVT U1333 ( .A1(\ram[0][218] ), .A3(\ram[2][218] ), .A2(
        \ram[1][218] ), .A4(\ram[3][218] ), .S0(n4231), .S1(n41), .Y(n5209) );
  MUX41X1_HVT U1334 ( .A1(n5209), .A3(n5207), .A2(n5208), .A4(n5206), .S0(
        n4328), .S1(n4305), .Y(q[218]) );
  MUX41X1_HVT U1335 ( .A1(\ram[12][219] ), .A3(\ram[14][219] ), .A2(
        \ram[13][219] ), .A4(\ram[15][219] ), .S0(n4232), .S1(n42), .Y(n5210)
         );
  MUX41X1_HVT U1336 ( .A1(\ram[8][219] ), .A3(\ram[10][219] ), .A2(
        \ram[9][219] ), .A4(\ram[11][219] ), .S0(n4232), .S1(n42), .Y(n5211)
         );
  MUX41X1_HVT U1337 ( .A1(\ram[4][219] ), .A3(\ram[6][219] ), .A2(
        \ram[5][219] ), .A4(\ram[7][219] ), .S0(n4232), .S1(n42), .Y(n5212) );
  MUX41X1_HVT U1338 ( .A1(\ram[0][219] ), .A3(\ram[2][219] ), .A2(
        \ram[1][219] ), .A4(\ram[3][219] ), .S0(n4232), .S1(n42), .Y(n5213) );
  MUX41X1_HVT U1339 ( .A1(n5213), .A3(n5211), .A2(n5212), .A4(n5210), .S0(
        n4328), .S1(n4305), .Y(q[219]) );
  MUX41X1_HVT U1340 ( .A1(\ram[12][220] ), .A3(\ram[14][220] ), .A2(
        \ram[13][220] ), .A4(\ram[15][220] ), .S0(n4232), .S1(n42), .Y(n5214)
         );
  MUX41X1_HVT U1341 ( .A1(\ram[8][220] ), .A3(\ram[10][220] ), .A2(
        \ram[9][220] ), .A4(\ram[11][220] ), .S0(n4232), .S1(n42), .Y(n5215)
         );
  MUX41X1_HVT U1342 ( .A1(\ram[4][220] ), .A3(\ram[6][220] ), .A2(
        \ram[5][220] ), .A4(\ram[7][220] ), .S0(n4232), .S1(n42), .Y(n5216) );
  MUX41X1_HVT U1343 ( .A1(\ram[0][220] ), .A3(\ram[2][220] ), .A2(
        \ram[1][220] ), .A4(\ram[3][220] ), .S0(n4232), .S1(n42), .Y(n5217) );
  MUX41X1_HVT U1344 ( .A1(n5217), .A3(n5215), .A2(n5216), .A4(n5214), .S0(
        n4328), .S1(n4305), .Y(q[220]) );
  MUX41X1_HVT U1345 ( .A1(\ram[12][221] ), .A3(\ram[14][221] ), .A2(
        \ram[13][221] ), .A4(\ram[15][221] ), .S0(n4232), .S1(n42), .Y(n5218)
         );
  MUX41X1_HVT U1346 ( .A1(\ram[8][221] ), .A3(\ram[10][221] ), .A2(
        \ram[9][221] ), .A4(\ram[11][221] ), .S0(n4232), .S1(n42), .Y(n5219)
         );
  MUX41X1_HVT U1347 ( .A1(\ram[4][221] ), .A3(\ram[6][221] ), .A2(
        \ram[5][221] ), .A4(\ram[7][221] ), .S0(n4232), .S1(n42), .Y(n5220) );
  MUX41X1_HVT U1348 ( .A1(\ram[0][221] ), .A3(\ram[2][221] ), .A2(
        \ram[1][221] ), .A4(\ram[3][221] ), .S0(n4232), .S1(n42), .Y(n5221) );
  MUX41X1_HVT U1349 ( .A1(n5221), .A3(n5219), .A2(n5220), .A4(n5218), .S0(
        n4328), .S1(n4305), .Y(q[221]) );
  MUX41X1_HVT U1350 ( .A1(\ram[12][222] ), .A3(\ram[14][222] ), .A2(
        \ram[13][222] ), .A4(\ram[15][222] ), .S0(n4233), .S1(n43), .Y(n5222)
         );
  MUX41X1_HVT U1351 ( .A1(\ram[8][222] ), .A3(\ram[10][222] ), .A2(
        \ram[9][222] ), .A4(\ram[11][222] ), .S0(n4233), .S1(n43), .Y(n5223)
         );
  MUX41X1_HVT U1352 ( .A1(\ram[4][222] ), .A3(\ram[6][222] ), .A2(
        \ram[5][222] ), .A4(\ram[7][222] ), .S0(n4233), .S1(n43), .Y(n5224) );
  MUX41X1_HVT U1353 ( .A1(\ram[0][222] ), .A3(\ram[2][222] ), .A2(
        \ram[1][222] ), .A4(\ram[3][222] ), .S0(n4233), .S1(n43), .Y(n5225) );
  MUX41X1_HVT U1354 ( .A1(n5225), .A3(n5223), .A2(n5224), .A4(n5222), .S0(
        n4328), .S1(n4305), .Y(q[222]) );
  MUX41X1_HVT U1355 ( .A1(\ram[12][223] ), .A3(\ram[14][223] ), .A2(
        \ram[13][223] ), .A4(\ram[15][223] ), .S0(n4233), .S1(n43), .Y(n5226)
         );
  MUX41X1_HVT U1356 ( .A1(\ram[8][223] ), .A3(\ram[10][223] ), .A2(
        \ram[9][223] ), .A4(\ram[11][223] ), .S0(n4233), .S1(n43), .Y(n5227)
         );
  MUX41X1_HVT U1357 ( .A1(\ram[4][223] ), .A3(\ram[6][223] ), .A2(
        \ram[5][223] ), .A4(\ram[7][223] ), .S0(n4233), .S1(n43), .Y(n5228) );
  MUX41X1_HVT U1358 ( .A1(\ram[0][223] ), .A3(\ram[2][223] ), .A2(
        \ram[1][223] ), .A4(\ram[3][223] ), .S0(n4233), .S1(n43), .Y(n5229) );
  MUX41X1_HVT U1359 ( .A1(n5229), .A3(n5227), .A2(n5228), .A4(n5226), .S0(
        n4328), .S1(n4305), .Y(q[223]) );
  MUX41X1_HVT U1360 ( .A1(\ram[12][224] ), .A3(\ram[14][224] ), .A2(
        \ram[13][224] ), .A4(\ram[15][224] ), .S0(n4217), .S1(n27), .Y(n5230)
         );
  MUX41X1_HVT U1361 ( .A1(\ram[8][224] ), .A3(\ram[10][224] ), .A2(
        \ram[9][224] ), .A4(\ram[11][224] ), .S0(n4212), .S1(n22), .Y(n5231)
         );
  MUX41X1_HVT U1362 ( .A1(\ram[4][224] ), .A3(\ram[6][224] ), .A2(
        \ram[5][224] ), .A4(\ram[7][224] ), .S0(n4212), .S1(n22), .Y(n5232) );
  MUX41X1_HVT U1363 ( .A1(\ram[0][224] ), .A3(\ram[2][224] ), .A2(
        \ram[1][224] ), .A4(\ram[3][224] ), .S0(n4212), .S1(n22), .Y(n5233) );
  MUX41X1_HVT U1364 ( .A1(n5233), .A3(n5231), .A2(n5232), .A4(n5230), .S0(
        n4328), .S1(n4305), .Y(q[224]) );
  MUX41X1_HVT U1365 ( .A1(\ram[12][225] ), .A3(\ram[14][225] ), .A2(
        \ram[13][225] ), .A4(\ram[15][225] ), .S0(n4212), .S1(n22), .Y(n5234)
         );
  MUX41X1_HVT U1366 ( .A1(\ram[8][225] ), .A3(\ram[10][225] ), .A2(
        \ram[9][225] ), .A4(\ram[11][225] ), .S0(n4212), .S1(n22), .Y(n5235)
         );
  MUX41X1_HVT U1367 ( .A1(\ram[4][225] ), .A3(\ram[6][225] ), .A2(
        \ram[5][225] ), .A4(\ram[7][225] ), .S0(n4212), .S1(n22), .Y(n5236) );
  MUX41X1_HVT U1368 ( .A1(\ram[0][225] ), .A3(\ram[2][225] ), .A2(
        \ram[1][225] ), .A4(\ram[3][225] ), .S0(n4212), .S1(n22), .Y(n5237) );
  MUX41X1_HVT U1369 ( .A1(n5237), .A3(n5235), .A2(n5236), .A4(n5234), .S0(
        n4328), .S1(n4305), .Y(q[225]) );
  MUX41X1_HVT U1370 ( .A1(\ram[12][226] ), .A3(\ram[14][226] ), .A2(
        \ram[13][226] ), .A4(\ram[15][226] ), .S0(n4213), .S1(n23), .Y(n5238)
         );
  MUX41X1_HVT U1371 ( .A1(\ram[8][226] ), .A3(\ram[10][226] ), .A2(
        \ram[9][226] ), .A4(\ram[11][226] ), .S0(n4213), .S1(n23), .Y(n5239)
         );
  MUX41X1_HVT U1372 ( .A1(\ram[4][226] ), .A3(\ram[6][226] ), .A2(
        \ram[5][226] ), .A4(\ram[7][226] ), .S0(n4213), .S1(n23), .Y(n5240) );
  MUX41X1_HVT U1373 ( .A1(\ram[0][226] ), .A3(\ram[2][226] ), .A2(
        \ram[1][226] ), .A4(\ram[3][226] ), .S0(n4213), .S1(n23), .Y(n5241) );
  MUX41X1_HVT U1374 ( .A1(n5241), .A3(n5239), .A2(n5240), .A4(n5238), .S0(
        n4328), .S1(n4305), .Y(q[226]) );
  MUX41X1_HVT U1375 ( .A1(\ram[12][227] ), .A3(\ram[14][227] ), .A2(
        \ram[13][227] ), .A4(\ram[15][227] ), .S0(n4213), .S1(n23), .Y(n5242)
         );
  MUX41X1_HVT U1376 ( .A1(\ram[8][227] ), .A3(\ram[10][227] ), .A2(
        \ram[9][227] ), .A4(\ram[11][227] ), .S0(n4213), .S1(n23), .Y(n5243)
         );
  MUX41X1_HVT U1377 ( .A1(\ram[4][227] ), .A3(\ram[6][227] ), .A2(
        \ram[5][227] ), .A4(\ram[7][227] ), .S0(n4213), .S1(n23), .Y(n5244) );
  MUX41X1_HVT U1378 ( .A1(\ram[0][227] ), .A3(\ram[2][227] ), .A2(
        \ram[1][227] ), .A4(\ram[3][227] ), .S0(n4213), .S1(n23), .Y(n5245) );
  MUX41X1_HVT U1379 ( .A1(n5245), .A3(n5243), .A2(n5244), .A4(n5242), .S0(
        n4328), .S1(n4305), .Y(q[227]) );
  MUX41X1_HVT U1380 ( .A1(\ram[12][228] ), .A3(\ram[14][228] ), .A2(
        \ram[13][228] ), .A4(\ram[15][228] ), .S0(n4213), .S1(n23), .Y(n5246)
         );
  MUX41X1_HVT U1381 ( .A1(\ram[8][228] ), .A3(\ram[10][228] ), .A2(
        \ram[9][228] ), .A4(\ram[11][228] ), .S0(n4213), .S1(n23), .Y(n5247)
         );
  MUX41X1_HVT U1382 ( .A1(\ram[4][228] ), .A3(\ram[6][228] ), .A2(
        \ram[5][228] ), .A4(\ram[7][228] ), .S0(n4213), .S1(n23), .Y(n5248) );
  MUX41X1_HVT U1383 ( .A1(\ram[0][228] ), .A3(\ram[2][228] ), .A2(
        \ram[1][228] ), .A4(\ram[3][228] ), .S0(n4213), .S1(n23), .Y(n5249) );
  MUX41X1_HVT U1384 ( .A1(n5249), .A3(n5247), .A2(n5248), .A4(n5246), .S0(
        n4329), .S1(n4306), .Y(q[228]) );
  MUX41X1_HVT U1385 ( .A1(\ram[12][229] ), .A3(\ram[14][229] ), .A2(
        \ram[13][229] ), .A4(\ram[15][229] ), .S0(n4214), .S1(n24), .Y(n5250)
         );
  MUX41X1_HVT U1386 ( .A1(\ram[8][229] ), .A3(\ram[10][229] ), .A2(
        \ram[9][229] ), .A4(\ram[11][229] ), .S0(n4214), .S1(n24), .Y(n5251)
         );
  MUX41X1_HVT U1387 ( .A1(\ram[4][229] ), .A3(\ram[6][229] ), .A2(
        \ram[5][229] ), .A4(\ram[7][229] ), .S0(n4214), .S1(n24), .Y(n5252) );
  MUX41X1_HVT U1388 ( .A1(\ram[0][229] ), .A3(\ram[2][229] ), .A2(
        \ram[1][229] ), .A4(\ram[3][229] ), .S0(n4214), .S1(n24), .Y(n5253) );
  MUX41X1_HVT U1389 ( .A1(n5253), .A3(n5251), .A2(n5252), .A4(n5250), .S0(
        n4329), .S1(n4306), .Y(q[229]) );
  MUX41X1_HVT U1390 ( .A1(\ram[12][230] ), .A3(\ram[14][230] ), .A2(
        \ram[13][230] ), .A4(\ram[15][230] ), .S0(n4214), .S1(n24), .Y(n5254)
         );
  MUX41X1_HVT U1391 ( .A1(\ram[8][230] ), .A3(\ram[10][230] ), .A2(
        \ram[9][230] ), .A4(\ram[11][230] ), .S0(n4214), .S1(n24), .Y(n5255)
         );
  MUX41X1_HVT U1392 ( .A1(\ram[4][230] ), .A3(\ram[6][230] ), .A2(
        \ram[5][230] ), .A4(\ram[7][230] ), .S0(n4214), .S1(n24), .Y(n5256) );
  MUX41X1_HVT U1393 ( .A1(\ram[0][230] ), .A3(\ram[2][230] ), .A2(
        \ram[1][230] ), .A4(\ram[3][230] ), .S0(n4214), .S1(n24), .Y(n5257) );
  MUX41X1_HVT U1394 ( .A1(n5257), .A3(n5255), .A2(n5256), .A4(n5254), .S0(
        n4329), .S1(n4306), .Y(q[230]) );
  MUX41X1_HVT U1395 ( .A1(\ram[12][231] ), .A3(\ram[14][231] ), .A2(
        \ram[13][231] ), .A4(\ram[15][231] ), .S0(n4214), .S1(n24), .Y(n5258)
         );
  MUX41X1_HVT U1396 ( .A1(\ram[8][231] ), .A3(\ram[10][231] ), .A2(
        \ram[9][231] ), .A4(\ram[11][231] ), .S0(n4214), .S1(n24), .Y(n5259)
         );
  MUX41X1_HVT U1397 ( .A1(\ram[4][231] ), .A3(\ram[6][231] ), .A2(
        \ram[5][231] ), .A4(\ram[7][231] ), .S0(n4214), .S1(n24), .Y(n5260) );
  MUX41X1_HVT U1398 ( .A1(\ram[0][231] ), .A3(\ram[2][231] ), .A2(
        \ram[1][231] ), .A4(\ram[3][231] ), .S0(n4214), .S1(n24), .Y(n5261) );
  MUX41X1_HVT U1399 ( .A1(n5261), .A3(n5259), .A2(n5260), .A4(n5258), .S0(
        n4329), .S1(n4306), .Y(q[231]) );
  MUX41X1_HVT U1400 ( .A1(\ram[12][232] ), .A3(\ram[14][232] ), .A2(
        \ram[13][232] ), .A4(\ram[15][232] ), .S0(n4215), .S1(n25), .Y(n5262)
         );
  MUX41X1_HVT U1401 ( .A1(\ram[8][232] ), .A3(\ram[10][232] ), .A2(
        \ram[9][232] ), .A4(\ram[11][232] ), .S0(n4215), .S1(n25), .Y(n5263)
         );
  MUX41X1_HVT U1402 ( .A1(\ram[4][232] ), .A3(\ram[6][232] ), .A2(
        \ram[5][232] ), .A4(\ram[7][232] ), .S0(n4215), .S1(n25), .Y(n5264) );
  MUX41X1_HVT U1403 ( .A1(\ram[0][232] ), .A3(\ram[2][232] ), .A2(
        \ram[1][232] ), .A4(\ram[3][232] ), .S0(n4215), .S1(n25), .Y(n5265) );
  MUX41X1_HVT U1404 ( .A1(n5265), .A3(n5263), .A2(n5264), .A4(n5262), .S0(
        n4329), .S1(n4306), .Y(q[232]) );
  MUX41X1_HVT U1405 ( .A1(\ram[12][233] ), .A3(\ram[14][233] ), .A2(
        \ram[13][233] ), .A4(\ram[15][233] ), .S0(n4215), .S1(n25), .Y(n5266)
         );
  MUX41X1_HVT U1406 ( .A1(\ram[8][233] ), .A3(\ram[10][233] ), .A2(
        \ram[9][233] ), .A4(\ram[11][233] ), .S0(n4215), .S1(n25), .Y(n5267)
         );
  MUX41X1_HVT U1407 ( .A1(\ram[4][233] ), .A3(\ram[6][233] ), .A2(
        \ram[5][233] ), .A4(\ram[7][233] ), .S0(n4215), .S1(n25), .Y(n5268) );
  MUX41X1_HVT U1408 ( .A1(\ram[0][233] ), .A3(\ram[2][233] ), .A2(
        \ram[1][233] ), .A4(\ram[3][233] ), .S0(n4215), .S1(n25), .Y(n5269) );
  MUX41X1_HVT U1409 ( .A1(n5269), .A3(n5267), .A2(n5268), .A4(n5266), .S0(
        n4329), .S1(n4306), .Y(q[233]) );
  MUX41X1_HVT U1410 ( .A1(\ram[12][234] ), .A3(\ram[14][234] ), .A2(
        \ram[13][234] ), .A4(\ram[15][234] ), .S0(n4215), .S1(n25), .Y(n5270)
         );
  MUX41X1_HVT U1411 ( .A1(\ram[8][234] ), .A3(\ram[10][234] ), .A2(
        \ram[9][234] ), .A4(\ram[11][234] ), .S0(n4215), .S1(n25), .Y(n5271)
         );
  MUX41X1_HVT U1412 ( .A1(\ram[4][234] ), .A3(\ram[6][234] ), .A2(
        \ram[5][234] ), .A4(\ram[7][234] ), .S0(n4215), .S1(n25), .Y(n5272) );
  MUX41X1_HVT U1413 ( .A1(\ram[0][234] ), .A3(\ram[2][234] ), .A2(
        \ram[1][234] ), .A4(\ram[3][234] ), .S0(n4215), .S1(n25), .Y(n5273) );
  MUX41X1_HVT U1414 ( .A1(n5273), .A3(n5271), .A2(n5272), .A4(n5270), .S0(
        n4329), .S1(n4306), .Y(q[234]) );
  MUX41X1_HVT U1415 ( .A1(\ram[12][235] ), .A3(\ram[14][235] ), .A2(
        \ram[13][235] ), .A4(\ram[15][235] ), .S0(n4216), .S1(n26), .Y(n5274)
         );
  MUX41X1_HVT U1416 ( .A1(\ram[8][235] ), .A3(\ram[10][235] ), .A2(
        \ram[9][235] ), .A4(\ram[11][235] ), .S0(n4216), .S1(n26), .Y(n5275)
         );
  MUX41X1_HVT U1417 ( .A1(\ram[4][235] ), .A3(\ram[6][235] ), .A2(
        \ram[5][235] ), .A4(\ram[7][235] ), .S0(n4216), .S1(n26), .Y(n5276) );
  MUX41X1_HVT U1418 ( .A1(\ram[0][235] ), .A3(\ram[2][235] ), .A2(
        \ram[1][235] ), .A4(\ram[3][235] ), .S0(n4216), .S1(n26), .Y(n5277) );
  MUX41X1_HVT U1419 ( .A1(n5277), .A3(n5275), .A2(n5276), .A4(n5274), .S0(
        n4329), .S1(n4306), .Y(q[235]) );
  MUX41X1_HVT U1420 ( .A1(\ram[12][236] ), .A3(\ram[14][236] ), .A2(
        \ram[13][236] ), .A4(\ram[15][236] ), .S0(n4216), .S1(n26), .Y(n5278)
         );
  MUX41X1_HVT U1421 ( .A1(\ram[8][236] ), .A3(\ram[10][236] ), .A2(
        \ram[9][236] ), .A4(\ram[11][236] ), .S0(n4216), .S1(n26), .Y(n5279)
         );
  MUX41X1_HVT U1422 ( .A1(\ram[4][236] ), .A3(\ram[6][236] ), .A2(
        \ram[5][236] ), .A4(\ram[7][236] ), .S0(n4216), .S1(n26), .Y(n5280) );
  MUX41X1_HVT U1423 ( .A1(\ram[0][236] ), .A3(\ram[2][236] ), .A2(
        \ram[1][236] ), .A4(\ram[3][236] ), .S0(n4216), .S1(n26), .Y(n5281) );
  MUX41X1_HVT U1424 ( .A1(n5281), .A3(n5279), .A2(n5280), .A4(n5278), .S0(
        n4329), .S1(n4306), .Y(q[236]) );
  MUX41X1_HVT U1425 ( .A1(\ram[12][237] ), .A3(\ram[14][237] ), .A2(
        \ram[13][237] ), .A4(\ram[15][237] ), .S0(n4216), .S1(n26), .Y(n5282)
         );
  MUX41X1_HVT U1426 ( .A1(\ram[8][237] ), .A3(\ram[10][237] ), .A2(
        \ram[9][237] ), .A4(\ram[11][237] ), .S0(n4216), .S1(n26), .Y(n5283)
         );
  MUX41X1_HVT U1427 ( .A1(\ram[4][237] ), .A3(\ram[6][237] ), .A2(
        \ram[5][237] ), .A4(\ram[7][237] ), .S0(n4216), .S1(n26), .Y(n5284) );
  MUX41X1_HVT U1428 ( .A1(\ram[0][237] ), .A3(\ram[2][237] ), .A2(
        \ram[1][237] ), .A4(\ram[3][237] ), .S0(n4216), .S1(n26), .Y(n5285) );
  MUX41X1_HVT U1429 ( .A1(n5285), .A3(n5283), .A2(n5284), .A4(n5282), .S0(
        n4329), .S1(n4306), .Y(q[237]) );
  MUX41X1_HVT U1430 ( .A1(\ram[12][238] ), .A3(\ram[14][238] ), .A2(
        \ram[13][238] ), .A4(\ram[15][238] ), .S0(n4217), .S1(n27), .Y(n5286)
         );
  MUX41X1_HVT U1431 ( .A1(\ram[8][238] ), .A3(\ram[10][238] ), .A2(
        \ram[9][238] ), .A4(\ram[11][238] ), .S0(n4217), .S1(n27), .Y(n5287)
         );
  MUX41X1_HVT U1432 ( .A1(\ram[4][238] ), .A3(\ram[6][238] ), .A2(
        \ram[5][238] ), .A4(\ram[7][238] ), .S0(n4217), .S1(n27), .Y(n5288) );
  MUX41X1_HVT U1433 ( .A1(\ram[0][238] ), .A3(\ram[2][238] ), .A2(
        \ram[1][238] ), .A4(\ram[3][238] ), .S0(n4217), .S1(n27), .Y(n5289) );
  MUX41X1_HVT U1434 ( .A1(n5289), .A3(n5287), .A2(n5288), .A4(n5286), .S0(
        n4329), .S1(n4306), .Y(q[238]) );
  MUX41X1_HVT U1435 ( .A1(\ram[12][239] ), .A3(\ram[14][239] ), .A2(
        \ram[13][239] ), .A4(\ram[15][239] ), .S0(n4217), .S1(n27), .Y(n5290)
         );
  MUX41X1_HVT U1436 ( .A1(\ram[8][239] ), .A3(\ram[10][239] ), .A2(
        \ram[9][239] ), .A4(\ram[11][239] ), .S0(n4217), .S1(n27), .Y(n5291)
         );
  MUX41X1_HVT U1437 ( .A1(\ram[4][239] ), .A3(\ram[6][239] ), .A2(
        \ram[5][239] ), .A4(\ram[7][239] ), .S0(n4217), .S1(n27), .Y(n5292) );
  MUX41X1_HVT U1438 ( .A1(\ram[0][239] ), .A3(\ram[2][239] ), .A2(
        \ram[1][239] ), .A4(\ram[3][239] ), .S0(n4217), .S1(n27), .Y(n5293) );
  MUX41X1_HVT U1439 ( .A1(n5293), .A3(n5291), .A2(n5292), .A4(n5290), .S0(
        n4329), .S1(n4306), .Y(q[239]) );
  MUX41X1_HVT U1440 ( .A1(\ram[12][240] ), .A3(\ram[14][240] ), .A2(
        \ram[13][240] ), .A4(\ram[15][240] ), .S0(n4217), .S1(n27), .Y(n5294)
         );
  MUX41X1_HVT U1441 ( .A1(\ram[8][240] ), .A3(\ram[10][240] ), .A2(
        \ram[9][240] ), .A4(\ram[11][240] ), .S0(n4217), .S1(n27), .Y(n5295)
         );
  MUX41X1_HVT U1442 ( .A1(\ram[4][240] ), .A3(\ram[6][240] ), .A2(
        \ram[5][240] ), .A4(\ram[7][240] ), .S0(n4217), .S1(n27), .Y(n5296) );
  MUX41X1_HVT U1443 ( .A1(\ram[0][240] ), .A3(\ram[2][240] ), .A2(
        \ram[1][240] ), .A4(\ram[3][240] ), .S0(n4218), .S1(n28), .Y(n5297) );
  MUX41X1_HVT U1444 ( .A1(n5297), .A3(n5295), .A2(n5296), .A4(n5294), .S0(
        n4330), .S1(n4307), .Y(q[240]) );
  MUX41X1_HVT U1445 ( .A1(\ram[12][241] ), .A3(\ram[14][241] ), .A2(
        \ram[13][241] ), .A4(\ram[15][241] ), .S0(n4218), .S1(n28), .Y(n5298)
         );
  MUX41X1_HVT U1446 ( .A1(\ram[8][241] ), .A3(\ram[10][241] ), .A2(
        \ram[9][241] ), .A4(\ram[11][241] ), .S0(n4218), .S1(n28), .Y(n5299)
         );
  MUX41X1_HVT U1447 ( .A1(\ram[4][241] ), .A3(\ram[6][241] ), .A2(
        \ram[5][241] ), .A4(\ram[7][241] ), .S0(n4218), .S1(n28), .Y(n5300) );
  MUX41X1_HVT U1448 ( .A1(\ram[0][241] ), .A3(\ram[2][241] ), .A2(
        \ram[1][241] ), .A4(\ram[3][241] ), .S0(n4218), .S1(n28), .Y(n5301) );
  MUX41X1_HVT U1449 ( .A1(n5301), .A3(n5299), .A2(n5300), .A4(n5298), .S0(
        n4330), .S1(n4307), .Y(q[241]) );
  MUX41X1_HVT U1450 ( .A1(\ram[12][242] ), .A3(\ram[14][242] ), .A2(
        \ram[13][242] ), .A4(\ram[15][242] ), .S0(n4218), .S1(n28), .Y(n5302)
         );
  MUX41X1_HVT U1451 ( .A1(\ram[8][242] ), .A3(\ram[10][242] ), .A2(
        \ram[9][242] ), .A4(\ram[11][242] ), .S0(n4218), .S1(n28), .Y(n5303)
         );
  MUX41X1_HVT U1452 ( .A1(\ram[4][242] ), .A3(\ram[6][242] ), .A2(
        \ram[5][242] ), .A4(\ram[7][242] ), .S0(n4218), .S1(n28), .Y(n5304) );
  MUX41X1_HVT U1453 ( .A1(\ram[0][242] ), .A3(\ram[2][242] ), .A2(
        \ram[1][242] ), .A4(\ram[3][242] ), .S0(n4218), .S1(n28), .Y(n5305) );
  MUX41X1_HVT U1454 ( .A1(n5305), .A3(n5303), .A2(n5304), .A4(n5302), .S0(
        n4330), .S1(n4307), .Y(q[242]) );
  MUX41X1_HVT U1455 ( .A1(\ram[12][243] ), .A3(\ram[14][243] ), .A2(
        \ram[13][243] ), .A4(\ram[15][243] ), .S0(n4218), .S1(n28), .Y(n5306)
         );
  MUX41X1_HVT U1456 ( .A1(\ram[8][243] ), .A3(\ram[10][243] ), .A2(
        \ram[9][243] ), .A4(\ram[11][243] ), .S0(n4218), .S1(n28), .Y(n5307)
         );
  MUX41X1_HVT U1457 ( .A1(\ram[4][243] ), .A3(\ram[6][243] ), .A2(
        \ram[5][243] ), .A4(\ram[7][243] ), .S0(n4218), .S1(n28), .Y(n5308) );
  MUX41X1_HVT U1458 ( .A1(\ram[0][243] ), .A3(\ram[2][243] ), .A2(
        \ram[1][243] ), .A4(\ram[3][243] ), .S0(n4219), .S1(n29), .Y(n5309) );
  MUX41X1_HVT U1459 ( .A1(n5309), .A3(n5307), .A2(n5308), .A4(n5306), .S0(
        n4330), .S1(n4307), .Y(q[243]) );
  MUX41X1_HVT U1460 ( .A1(\ram[12][244] ), .A3(\ram[14][244] ), .A2(
        \ram[13][244] ), .A4(\ram[15][244] ), .S0(n4219), .S1(n29), .Y(n5310)
         );
  MUX41X1_HVT U1461 ( .A1(\ram[8][244] ), .A3(\ram[10][244] ), .A2(
        \ram[9][244] ), .A4(\ram[11][244] ), .S0(n4219), .S1(n29), .Y(n5311)
         );
  MUX41X1_HVT U1462 ( .A1(\ram[4][244] ), .A3(\ram[6][244] ), .A2(
        \ram[5][244] ), .A4(\ram[7][244] ), .S0(n4219), .S1(n29), .Y(n5312) );
  MUX41X1_HVT U1463 ( .A1(\ram[0][244] ), .A3(\ram[2][244] ), .A2(
        \ram[1][244] ), .A4(\ram[3][244] ), .S0(n4219), .S1(n29), .Y(n5313) );
  MUX41X1_HVT U1464 ( .A1(n5313), .A3(n5311), .A2(n5312), .A4(n5310), .S0(
        n4330), .S1(n4307), .Y(q[244]) );
  MUX41X1_HVT U1465 ( .A1(\ram[12][245] ), .A3(\ram[14][245] ), .A2(
        \ram[13][245] ), .A4(\ram[15][245] ), .S0(n4219), .S1(n29), .Y(n5314)
         );
  MUX41X1_HVT U1466 ( .A1(\ram[8][245] ), .A3(\ram[10][245] ), .A2(
        \ram[9][245] ), .A4(\ram[11][245] ), .S0(n4219), .S1(n29), .Y(n5315)
         );
  MUX41X1_HVT U1467 ( .A1(\ram[4][245] ), .A3(\ram[6][245] ), .A2(
        \ram[5][245] ), .A4(\ram[7][245] ), .S0(n4219), .S1(n29), .Y(n5316) );
  MUX41X1_HVT U1468 ( .A1(\ram[0][245] ), .A3(\ram[2][245] ), .A2(
        \ram[1][245] ), .A4(\ram[3][245] ), .S0(n4219), .S1(n29), .Y(n5317) );
  MUX41X1_HVT U1469 ( .A1(n5317), .A3(n5315), .A2(n5316), .A4(n5314), .S0(
        n4330), .S1(n4307), .Y(q[245]) );
  MUX41X1_HVT U1470 ( .A1(\ram[12][246] ), .A3(\ram[14][246] ), .A2(
        \ram[13][246] ), .A4(\ram[15][246] ), .S0(n4219), .S1(n29), .Y(n5318)
         );
  MUX41X1_HVT U1471 ( .A1(\ram[8][246] ), .A3(\ram[10][246] ), .A2(
        \ram[9][246] ), .A4(\ram[11][246] ), .S0(n4219), .S1(n29), .Y(n5319)
         );
  MUX41X1_HVT U1472 ( .A1(\ram[4][246] ), .A3(\ram[6][246] ), .A2(
        \ram[5][246] ), .A4(\ram[7][246] ), .S0(n4219), .S1(n29), .Y(n5320) );
  MUX41X1_HVT U1473 ( .A1(\ram[0][246] ), .A3(\ram[2][246] ), .A2(
        \ram[1][246] ), .A4(\ram[3][246] ), .S0(n4220), .S1(n30), .Y(n5321) );
  MUX41X1_HVT U1474 ( .A1(n5321), .A3(n5319), .A2(n5320), .A4(n5318), .S0(
        n4330), .S1(n4307), .Y(q[246]) );
  MUX41X1_HVT U1475 ( .A1(\ram[12][247] ), .A3(\ram[14][247] ), .A2(
        \ram[13][247] ), .A4(\ram[15][247] ), .S0(n4220), .S1(n30), .Y(n5322)
         );
  MUX41X1_HVT U1476 ( .A1(\ram[8][247] ), .A3(\ram[10][247] ), .A2(
        \ram[9][247] ), .A4(\ram[11][247] ), .S0(n4220), .S1(n30), .Y(n5323)
         );
  MUX41X1_HVT U1477 ( .A1(\ram[4][247] ), .A3(\ram[6][247] ), .A2(
        \ram[5][247] ), .A4(\ram[7][247] ), .S0(n4220), .S1(n30), .Y(n5324) );
  MUX41X1_HVT U1478 ( .A1(\ram[0][247] ), .A3(\ram[2][247] ), .A2(
        \ram[1][247] ), .A4(\ram[3][247] ), .S0(n4220), .S1(n30), .Y(n5325) );
  MUX41X1_HVT U1479 ( .A1(n5325), .A3(n5323), .A2(n5324), .A4(n5322), .S0(
        n4330), .S1(n4307), .Y(q[247]) );
  MUX41X1_HVT U1480 ( .A1(\ram[12][248] ), .A3(\ram[14][248] ), .A2(
        \ram[13][248] ), .A4(\ram[15][248] ), .S0(n4220), .S1(n30), .Y(n5326)
         );
  MUX41X1_HVT U1481 ( .A1(\ram[8][248] ), .A3(\ram[10][248] ), .A2(
        \ram[9][248] ), .A4(\ram[11][248] ), .S0(n4220), .S1(n30), .Y(n5327)
         );
  MUX41X1_HVT U1482 ( .A1(\ram[4][248] ), .A3(\ram[6][248] ), .A2(
        \ram[5][248] ), .A4(\ram[7][248] ), .S0(n4220), .S1(n30), .Y(n5328) );
  MUX41X1_HVT U1483 ( .A1(\ram[0][248] ), .A3(\ram[2][248] ), .A2(
        \ram[1][248] ), .A4(\ram[3][248] ), .S0(n4220), .S1(n30), .Y(n5329) );
  MUX41X1_HVT U1484 ( .A1(n5329), .A3(n5327), .A2(n5328), .A4(n5326), .S0(
        n4330), .S1(n4307), .Y(q[248]) );
  MUX41X1_HVT U1485 ( .A1(\ram[12][249] ), .A3(\ram[14][249] ), .A2(
        \ram[13][249] ), .A4(\ram[15][249] ), .S0(n4220), .S1(n30), .Y(n5330)
         );
  MUX41X1_HVT U1486 ( .A1(\ram[8][249] ), .A3(\ram[10][249] ), .A2(
        \ram[9][249] ), .A4(\ram[11][249] ), .S0(n4220), .S1(n30), .Y(n5331)
         );
  MUX41X1_HVT U1487 ( .A1(\ram[4][249] ), .A3(\ram[6][249] ), .A2(
        \ram[5][249] ), .A4(\ram[7][249] ), .S0(n4220), .S1(n30), .Y(n5332) );
  MUX41X1_HVT U1488 ( .A1(\ram[0][249] ), .A3(\ram[2][249] ), .A2(
        \ram[1][249] ), .A4(\ram[3][249] ), .S0(n4221), .S1(n31), .Y(n5333) );
  MUX41X1_HVT U1489 ( .A1(n5333), .A3(n5331), .A2(n5332), .A4(n5330), .S0(
        n4330), .S1(n4307), .Y(q[249]) );
  MUX41X1_HVT U1490 ( .A1(\ram[12][250] ), .A3(\ram[14][250] ), .A2(
        \ram[13][250] ), .A4(\ram[15][250] ), .S0(n4221), .S1(n31), .Y(n5334)
         );
  MUX41X1_HVT U1491 ( .A1(\ram[8][250] ), .A3(\ram[10][250] ), .A2(
        \ram[9][250] ), .A4(\ram[11][250] ), .S0(n4221), .S1(n31), .Y(n5335)
         );
  MUX41X1_HVT U1492 ( .A1(\ram[4][250] ), .A3(\ram[6][250] ), .A2(
        \ram[5][250] ), .A4(\ram[7][250] ), .S0(n4221), .S1(n31), .Y(n5336) );
  MUX41X1_HVT U1493 ( .A1(\ram[0][250] ), .A3(\ram[2][250] ), .A2(
        \ram[1][250] ), .A4(\ram[3][250] ), .S0(n4221), .S1(n31), .Y(n5337) );
  MUX41X1_HVT U1494 ( .A1(n5337), .A3(n5335), .A2(n5336), .A4(n5334), .S0(
        n4330), .S1(n4307), .Y(q[250]) );
  MUX41X1_HVT U1495 ( .A1(\ram[12][251] ), .A3(\ram[14][251] ), .A2(
        \ram[13][251] ), .A4(\ram[15][251] ), .S0(n4221), .S1(n31), .Y(n5338)
         );
  MUX41X1_HVT U1496 ( .A1(\ram[8][251] ), .A3(\ram[10][251] ), .A2(
        \ram[9][251] ), .A4(\ram[11][251] ), .S0(n4221), .S1(n31), .Y(n5339)
         );
  MUX41X1_HVT U1497 ( .A1(\ram[4][251] ), .A3(\ram[6][251] ), .A2(
        \ram[5][251] ), .A4(\ram[7][251] ), .S0(n4221), .S1(n31), .Y(n5340) );
  MUX41X1_HVT U1498 ( .A1(\ram[0][251] ), .A3(\ram[2][251] ), .A2(
        \ram[1][251] ), .A4(\ram[3][251] ), .S0(n4221), .S1(n31), .Y(n5341) );
  MUX41X1_HVT U1499 ( .A1(n5341), .A3(n5339), .A2(n5340), .A4(n5338), .S0(
        n4330), .S1(n4307), .Y(q[251]) );
  MUX41X1_HVT U1500 ( .A1(\ram[12][252] ), .A3(\ram[14][252] ), .A2(
        \ram[13][252] ), .A4(\ram[15][252] ), .S0(n4221), .S1(n31), .Y(n5342)
         );
  MUX41X1_HVT U1501 ( .A1(\ram[8][252] ), .A3(\ram[10][252] ), .A2(
        \ram[9][252] ), .A4(\ram[11][252] ), .S0(n4221), .S1(n31), .Y(n5343)
         );
  MUX41X1_HVT U1502 ( .A1(\ram[4][252] ), .A3(\ram[6][252] ), .A2(
        \ram[5][252] ), .A4(\ram[7][252] ), .S0(n4221), .S1(n31), .Y(n5344) );
  MUX41X1_HVT U1503 ( .A1(\ram[0][252] ), .A3(\ram[2][252] ), .A2(
        \ram[1][252] ), .A4(\ram[3][252] ), .S0(n4222), .S1(n32), .Y(n5345) );
  MUX41X1_HVT U1504 ( .A1(n5345), .A3(n5343), .A2(n5344), .A4(n5342), .S0(N29), 
        .S1(N28), .Y(q[252]) );
  MUX41X1_HVT U1505 ( .A1(\ram[12][253] ), .A3(\ram[14][253] ), .A2(
        \ram[13][253] ), .A4(\ram[15][253] ), .S0(n4222), .S1(n32), .Y(n5346)
         );
  MUX41X1_HVT U1506 ( .A1(\ram[8][253] ), .A3(\ram[10][253] ), .A2(
        \ram[9][253] ), .A4(\ram[11][253] ), .S0(n4222), .S1(n32), .Y(n5347)
         );
  MUX41X1_HVT U1507 ( .A1(\ram[4][253] ), .A3(\ram[6][253] ), .A2(
        \ram[5][253] ), .A4(\ram[7][253] ), .S0(n4222), .S1(n32), .Y(n5348) );
  MUX41X1_HVT U1508 ( .A1(\ram[0][253] ), .A3(\ram[2][253] ), .A2(
        \ram[1][253] ), .A4(\ram[3][253] ), .S0(n4222), .S1(n32), .Y(n5349) );
  MUX41X1_HVT U1509 ( .A1(n5349), .A3(n5347), .A2(n5348), .A4(n5346), .S0(N29), 
        .S1(N28), .Y(q[253]) );
  MUX41X1_HVT U1510 ( .A1(\ram[12][254] ), .A3(\ram[14][254] ), .A2(
        \ram[13][254] ), .A4(\ram[15][254] ), .S0(n4222), .S1(n32), .Y(n5350)
         );
  MUX41X1_HVT U1511 ( .A1(\ram[8][254] ), .A3(\ram[10][254] ), .A2(
        \ram[9][254] ), .A4(\ram[11][254] ), .S0(n4222), .S1(n32), .Y(n5351)
         );
  MUX41X1_HVT U1512 ( .A1(\ram[4][254] ), .A3(\ram[6][254] ), .A2(
        \ram[5][254] ), .A4(\ram[7][254] ), .S0(n4222), .S1(n32), .Y(n5352) );
  MUX41X1_HVT U1513 ( .A1(\ram[0][254] ), .A3(\ram[2][254] ), .A2(
        \ram[1][254] ), .A4(\ram[3][254] ), .S0(n4222), .S1(n32), .Y(n5353) );
  MUX41X1_HVT U1514 ( .A1(n5353), .A3(n5351), .A2(n5352), .A4(n5350), .S0(N29), 
        .S1(N28), .Y(q[254]) );
  MUX41X1_HVT U1515 ( .A1(\ram[12][255] ), .A3(\ram[14][255] ), .A2(
        \ram[13][255] ), .A4(\ram[15][255] ), .S0(n4222), .S1(n32), .Y(n5354)
         );
  MUX41X1_HVT U1516 ( .A1(\ram[8][255] ), .A3(\ram[10][255] ), .A2(
        \ram[9][255] ), .A4(\ram[11][255] ), .S0(n4222), .S1(n32), .Y(n5355)
         );
  MUX41X1_HVT U1517 ( .A1(\ram[4][255] ), .A3(\ram[6][255] ), .A2(
        \ram[5][255] ), .A4(\ram[7][255] ), .S0(n4222), .S1(n32), .Y(n5356) );
  MUX41X1_HVT U1518 ( .A1(\ram[0][255] ), .A3(\ram[2][255] ), .A2(
        \ram[1][255] ), .A4(\ram[3][255] ), .S0(n4223), .S1(n33), .Y(n5357) );
  MUX41X1_HVT U1519 ( .A1(n5357), .A3(n5355), .A2(n5356), .A4(n5354), .S0(N29), 
        .S1(N28), .Y(q[255]) );
  AO22X1_HVT U1520 ( .A1(\ram[3][170] ), .A2(n5358), .A3(data[170]), .A4(n5359), .Y(n999) );
  AO22X1_HVT U1521 ( .A1(\ram[3][169] ), .A2(n5358), .A3(data[169]), .A4(n5359), .Y(n998) );
  AO22X1_HVT U1522 ( .A1(\ram[3][168] ), .A2(n5358), .A3(data[168]), .A4(n5359), .Y(n997) );
  AO22X1_HVT U1523 ( .A1(\ram[3][167] ), .A2(n5358), .A3(data[167]), .A4(n5359), .Y(n996) );
  AO22X1_HVT U1524 ( .A1(\ram[3][166] ), .A2(n5358), .A3(data[166]), .A4(n5359), .Y(n995) );
  AO22X1_HVT U1525 ( .A1(\ram[3][165] ), .A2(n5358), .A3(data[165]), .A4(n5359), .Y(n994) );
  AO22X1_HVT U1526 ( .A1(\ram[3][164] ), .A2(n5358), .A3(data[164]), .A4(n5359), .Y(n993) );
  AO22X1_HVT U1527 ( .A1(\ram[3][163] ), .A2(n5358), .A3(data[163]), .A4(n5359), .Y(n992) );
  AO22X1_HVT U1528 ( .A1(\ram[3][162] ), .A2(n5358), .A3(data[162]), .A4(n5359), .Y(n991) );
  AO22X1_HVT U1529 ( .A1(\ram[3][161] ), .A2(n5358), .A3(data[161]), .A4(n5359), .Y(n990) );
  AO22X1_HVT U1530 ( .A1(\ram[0][38] ), .A2(n5360), .A3(data[38]), .A4(n5361), 
        .Y(n99) );
  AO22X1_HVT U1531 ( .A1(\ram[3][160] ), .A2(n5358), .A3(data[160]), .A4(n5359), .Y(n989) );
  AO22X1_HVT U1532 ( .A1(\ram[3][159] ), .A2(n5358), .A3(data[159]), .A4(n5359), .Y(n988) );
  AO22X1_HVT U1533 ( .A1(\ram[3][158] ), .A2(n5358), .A3(data[158]), .A4(n5359), .Y(n987) );
  AO22X1_HVT U1534 ( .A1(\ram[3][157] ), .A2(n5358), .A3(data[157]), .A4(n5359), .Y(n986) );
  AO22X1_HVT U1535 ( .A1(\ram[3][156] ), .A2(n5358), .A3(data[156]), .A4(n5359), .Y(n985) );
  AO22X1_HVT U1536 ( .A1(\ram[3][155] ), .A2(n5358), .A3(data[155]), .A4(n5359), .Y(n984) );
  AO22X1_HVT U1537 ( .A1(\ram[3][154] ), .A2(n5358), .A3(data[154]), .A4(n5359), .Y(n983) );
  AO22X1_HVT U1538 ( .A1(\ram[3][153] ), .A2(n5358), .A3(data[153]), .A4(n5359), .Y(n982) );
  AO22X1_HVT U1539 ( .A1(\ram[3][152] ), .A2(n5358), .A3(data[152]), .A4(n5359), .Y(n981) );
  AO22X1_HVT U1540 ( .A1(\ram[3][151] ), .A2(n5358), .A3(data[151]), .A4(n5359), .Y(n980) );
  AO22X1_HVT U1541 ( .A1(\ram[0][37] ), .A2(n5360), .A3(data[37]), .A4(n5361), 
        .Y(n98) );
  AO22X1_HVT U1542 ( .A1(\ram[3][150] ), .A2(n5358), .A3(data[150]), .A4(n5359), .Y(n979) );
  AO22X1_HVT U1543 ( .A1(\ram[3][149] ), .A2(n5358), .A3(data[149]), .A4(n5359), .Y(n978) );
  AO22X1_HVT U1544 ( .A1(\ram[3][148] ), .A2(n5358), .A3(data[148]), .A4(n5359), .Y(n977) );
  AO22X1_HVT U1545 ( .A1(\ram[3][147] ), .A2(n5358), .A3(data[147]), .A4(n5359), .Y(n976) );
  AO22X1_HVT U1546 ( .A1(\ram[3][146] ), .A2(n5358), .A3(data[146]), .A4(n5359), .Y(n975) );
  AO22X1_HVT U1547 ( .A1(\ram[3][145] ), .A2(n5358), .A3(data[145]), .A4(n5359), .Y(n974) );
  AO22X1_HVT U1548 ( .A1(\ram[3][144] ), .A2(n5358), .A3(data[144]), .A4(n5359), .Y(n973) );
  AO22X1_HVT U1549 ( .A1(\ram[3][143] ), .A2(n5358), .A3(data[143]), .A4(n5359), .Y(n972) );
  AO22X1_HVT U1550 ( .A1(\ram[3][142] ), .A2(n5358), .A3(data[142]), .A4(n5359), .Y(n971) );
  AO22X1_HVT U1551 ( .A1(\ram[3][141] ), .A2(n5358), .A3(data[141]), .A4(n5359), .Y(n970) );
  AO22X1_HVT U1552 ( .A1(\ram[0][36] ), .A2(n5360), .A3(data[36]), .A4(n5361), 
        .Y(n97) );
  AO22X1_HVT U1553 ( .A1(\ram[3][140] ), .A2(n5358), .A3(data[140]), .A4(n5359), .Y(n969) );
  AO22X1_HVT U1554 ( .A1(\ram[3][139] ), .A2(n5358), .A3(data[139]), .A4(n5359), .Y(n968) );
  AO22X1_HVT U1555 ( .A1(\ram[3][138] ), .A2(n5358), .A3(data[138]), .A4(n5359), .Y(n967) );
  AO22X1_HVT U1556 ( .A1(\ram[3][137] ), .A2(n5358), .A3(data[137]), .A4(n5359), .Y(n966) );
  AO22X1_HVT U1557 ( .A1(\ram[3][136] ), .A2(n5358), .A3(data[136]), .A4(n5359), .Y(n965) );
  AO22X1_HVT U1558 ( .A1(\ram[3][135] ), .A2(n5358), .A3(data[135]), .A4(n5359), .Y(n964) );
  AO22X1_HVT U1559 ( .A1(\ram[3][134] ), .A2(n5358), .A3(data[134]), .A4(n5359), .Y(n963) );
  AO22X1_HVT U1560 ( .A1(\ram[3][133] ), .A2(n5358), .A3(data[133]), .A4(n5359), .Y(n962) );
  AO22X1_HVT U1561 ( .A1(\ram[3][132] ), .A2(n5358), .A3(data[132]), .A4(n5359), .Y(n961) );
  AO22X1_HVT U1562 ( .A1(\ram[3][131] ), .A2(n5358), .A3(data[131]), .A4(n5359), .Y(n960) );
  AO22X1_HVT U1563 ( .A1(\ram[0][35] ), .A2(n5360), .A3(data[35]), .A4(n5361), 
        .Y(n96) );
  AO22X1_HVT U1564 ( .A1(\ram[3][130] ), .A2(n5358), .A3(data[130]), .A4(n5359), .Y(n959) );
  AO22X1_HVT U1565 ( .A1(\ram[3][129] ), .A2(n5358), .A3(data[129]), .A4(n5359), .Y(n958) );
  AO22X1_HVT U1566 ( .A1(\ram[3][128] ), .A2(n5358), .A3(data[128]), .A4(n5359), .Y(n957) );
  AO22X1_HVT U1567 ( .A1(\ram[3][127] ), .A2(n5358), .A3(data[127]), .A4(n5359), .Y(n956) );
  AO22X1_HVT U1568 ( .A1(\ram[3][126] ), .A2(n5358), .A3(data[126]), .A4(n5359), .Y(n955) );
  AO22X1_HVT U1569 ( .A1(\ram[3][125] ), .A2(n5358), .A3(data[125]), .A4(n5359), .Y(n954) );
  AO22X1_HVT U1570 ( .A1(\ram[3][124] ), .A2(n5358), .A3(data[124]), .A4(n5359), .Y(n953) );
  AO22X1_HVT U1571 ( .A1(\ram[3][123] ), .A2(n5358), .A3(data[123]), .A4(n5359), .Y(n952) );
  AO22X1_HVT U1572 ( .A1(\ram[3][122] ), .A2(n5358), .A3(data[122]), .A4(n5359), .Y(n951) );
  AO22X1_HVT U1573 ( .A1(\ram[3][121] ), .A2(n5358), .A3(data[121]), .A4(n5359), .Y(n950) );
  AO22X1_HVT U1574 ( .A1(\ram[0][34] ), .A2(n5360), .A3(data[34]), .A4(n5361), 
        .Y(n95) );
  AO22X1_HVT U1575 ( .A1(\ram[3][120] ), .A2(n5358), .A3(data[120]), .A4(n5359), .Y(n949) );
  AO22X1_HVT U1576 ( .A1(\ram[3][119] ), .A2(n5358), .A3(data[119]), .A4(n5359), .Y(n948) );
  AO22X1_HVT U1577 ( .A1(\ram[3][118] ), .A2(n5358), .A3(data[118]), .A4(n5359), .Y(n947) );
  AO22X1_HVT U1578 ( .A1(\ram[3][117] ), .A2(n5358), .A3(data[117]), .A4(n5359), .Y(n946) );
  AO22X1_HVT U1579 ( .A1(\ram[3][116] ), .A2(n5358), .A3(data[116]), .A4(n5359), .Y(n945) );
  AO22X1_HVT U1580 ( .A1(\ram[3][115] ), .A2(n5358), .A3(data[115]), .A4(n5359), .Y(n944) );
  AO22X1_HVT U1581 ( .A1(\ram[3][114] ), .A2(n5358), .A3(data[114]), .A4(n5359), .Y(n943) );
  AO22X1_HVT U1582 ( .A1(\ram[3][113] ), .A2(n5358), .A3(data[113]), .A4(n5359), .Y(n942) );
  AO22X1_HVT U1583 ( .A1(\ram[3][112] ), .A2(n5358), .A3(data[112]), .A4(n5359), .Y(n941) );
  AO22X1_HVT U1584 ( .A1(\ram[3][111] ), .A2(n5358), .A3(data[111]), .A4(n5359), .Y(n940) );
  AO22X1_HVT U1585 ( .A1(\ram[0][33] ), .A2(n5360), .A3(data[33]), .A4(n5361), 
        .Y(n94) );
  AO22X1_HVT U1586 ( .A1(\ram[3][110] ), .A2(n5358), .A3(data[110]), .A4(n5359), .Y(n939) );
  AO22X1_HVT U1587 ( .A1(\ram[3][109] ), .A2(n5358), .A3(data[109]), .A4(n5359), .Y(n938) );
  AO22X1_HVT U1588 ( .A1(\ram[3][108] ), .A2(n5358), .A3(data[108]), .A4(n5359), .Y(n937) );
  AO22X1_HVT U1589 ( .A1(\ram[3][107] ), .A2(n5358), .A3(data[107]), .A4(n5359), .Y(n936) );
  AO22X1_HVT U1590 ( .A1(\ram[3][106] ), .A2(n5358), .A3(data[106]), .A4(n5359), .Y(n935) );
  AO22X1_HVT U1591 ( .A1(\ram[3][105] ), .A2(n5358), .A3(data[105]), .A4(n5359), .Y(n934) );
  AO22X1_HVT U1592 ( .A1(\ram[3][104] ), .A2(n5358), .A3(data[104]), .A4(n5359), .Y(n933) );
  AO22X1_HVT U1593 ( .A1(\ram[3][103] ), .A2(n5358), .A3(data[103]), .A4(n5359), .Y(n932) );
  AO22X1_HVT U1594 ( .A1(\ram[3][102] ), .A2(n5358), .A3(data[102]), .A4(n5359), .Y(n931) );
  AO22X1_HVT U1595 ( .A1(\ram[3][101] ), .A2(n5358), .A3(data[101]), .A4(n5359), .Y(n930) );
  AO22X1_HVT U1596 ( .A1(\ram[0][32] ), .A2(n5360), .A3(data[32]), .A4(n5361), 
        .Y(n93) );
  AO22X1_HVT U1597 ( .A1(\ram[3][100] ), .A2(n5358), .A3(data[100]), .A4(n5359), .Y(n929) );
  AO22X1_HVT U1598 ( .A1(\ram[3][99] ), .A2(n5358), .A3(data[99]), .A4(n5359), 
        .Y(n928) );
  AO22X1_HVT U1599 ( .A1(\ram[3][98] ), .A2(n5358), .A3(data[98]), .A4(n5359), 
        .Y(n927) );
  AO22X1_HVT U1600 ( .A1(\ram[3][97] ), .A2(n5358), .A3(data[97]), .A4(n5359), 
        .Y(n926) );
  AO22X1_HVT U1601 ( .A1(\ram[3][96] ), .A2(n5358), .A3(data[96]), .A4(n5359), 
        .Y(n925) );
  AO22X1_HVT U1602 ( .A1(\ram[3][95] ), .A2(n5358), .A3(data[95]), .A4(n5359), 
        .Y(n924) );
  AO22X1_HVT U1603 ( .A1(\ram[3][94] ), .A2(n5358), .A3(data[94]), .A4(n5359), 
        .Y(n923) );
  AO22X1_HVT U1604 ( .A1(\ram[3][93] ), .A2(n5358), .A3(data[93]), .A4(n5359), 
        .Y(n922) );
  AO22X1_HVT U1605 ( .A1(\ram[3][92] ), .A2(n5358), .A3(data[92]), .A4(n5359), 
        .Y(n921) );
  AO22X1_HVT U1606 ( .A1(\ram[3][91] ), .A2(n5358), .A3(data[91]), .A4(n5359), 
        .Y(n920) );
  AO22X1_HVT U1607 ( .A1(\ram[0][31] ), .A2(n5360), .A3(data[31]), .A4(n5361), 
        .Y(n92) );
  AO22X1_HVT U1608 ( .A1(\ram[3][90] ), .A2(n5358), .A3(data[90]), .A4(n5359), 
        .Y(n919) );
  AO22X1_HVT U1609 ( .A1(\ram[3][89] ), .A2(n5358), .A3(data[89]), .A4(n5359), 
        .Y(n918) );
  AO22X1_HVT U1610 ( .A1(\ram[3][88] ), .A2(n5358), .A3(data[88]), .A4(n5359), 
        .Y(n917) );
  AO22X1_HVT U1611 ( .A1(\ram[3][87] ), .A2(n5358), .A3(data[87]), .A4(n5359), 
        .Y(n916) );
  AO22X1_HVT U1612 ( .A1(\ram[3][86] ), .A2(n5358), .A3(data[86]), .A4(n5359), 
        .Y(n915) );
  AO22X1_HVT U1613 ( .A1(\ram[3][85] ), .A2(n5358), .A3(data[85]), .A4(n5359), 
        .Y(n914) );
  AO22X1_HVT U1614 ( .A1(\ram[3][84] ), .A2(n5358), .A3(data[84]), .A4(n5359), 
        .Y(n913) );
  AO22X1_HVT U1615 ( .A1(\ram[3][83] ), .A2(n5358), .A3(data[83]), .A4(n5359), 
        .Y(n912) );
  AO22X1_HVT U1616 ( .A1(\ram[3][82] ), .A2(n5358), .A3(data[82]), .A4(n5359), 
        .Y(n911) );
  AO22X1_HVT U1617 ( .A1(\ram[3][81] ), .A2(n5358), .A3(data[81]), .A4(n5359), 
        .Y(n910) );
  AO22X1_HVT U1618 ( .A1(\ram[0][30] ), .A2(n5360), .A3(data[30]), .A4(n5361), 
        .Y(n91) );
  AO22X1_HVT U1619 ( .A1(\ram[3][80] ), .A2(n5358), .A3(data[80]), .A4(n5359), 
        .Y(n909) );
  AO22X1_HVT U1620 ( .A1(\ram[3][79] ), .A2(n5358), .A3(data[79]), .A4(n5359), 
        .Y(n908) );
  AO22X1_HVT U1621 ( .A1(\ram[3][78] ), .A2(n5358), .A3(data[78]), .A4(n5359), 
        .Y(n907) );
  AO22X1_HVT U1622 ( .A1(\ram[3][77] ), .A2(n5358), .A3(data[77]), .A4(n5359), 
        .Y(n906) );
  AO22X1_HVT U1623 ( .A1(\ram[3][76] ), .A2(n5358), .A3(data[76]), .A4(n5359), 
        .Y(n905) );
  AO22X1_HVT U1624 ( .A1(\ram[3][75] ), .A2(n5358), .A3(data[75]), .A4(n5359), 
        .Y(n904) );
  AO22X1_HVT U1625 ( .A1(\ram[3][74] ), .A2(n5358), .A3(data[74]), .A4(n5359), 
        .Y(n903) );
  AO22X1_HVT U1626 ( .A1(\ram[3][73] ), .A2(n5358), .A3(data[73]), .A4(n5359), 
        .Y(n902) );
  AO22X1_HVT U1627 ( .A1(\ram[3][72] ), .A2(n5358), .A3(data[72]), .A4(n5359), 
        .Y(n901) );
  AO22X1_HVT U1628 ( .A1(\ram[3][71] ), .A2(n5358), .A3(data[71]), .A4(n5359), 
        .Y(n900) );
  AO22X1_HVT U1629 ( .A1(\ram[0][29] ), .A2(n5360), .A3(data[29]), .A4(n5361), 
        .Y(n90) );
  AO22X1_HVT U1630 ( .A1(\ram[3][70] ), .A2(n5358), .A3(data[70]), .A4(n5359), 
        .Y(n899) );
  AO22X1_HVT U1631 ( .A1(\ram[3][69] ), .A2(n5358), .A3(data[69]), .A4(n5359), 
        .Y(n898) );
  AO22X1_HVT U1632 ( .A1(\ram[3][68] ), .A2(n5358), .A3(data[68]), .A4(n5359), 
        .Y(n897) );
  AO22X1_HVT U1633 ( .A1(\ram[3][67] ), .A2(n5358), .A3(data[67]), .A4(n5359), 
        .Y(n896) );
  AO22X1_HVT U1634 ( .A1(\ram[3][66] ), .A2(n5358), .A3(data[66]), .A4(n5359), 
        .Y(n895) );
  AO22X1_HVT U1635 ( .A1(\ram[3][65] ), .A2(n5358), .A3(data[65]), .A4(n5359), 
        .Y(n894) );
  AO22X1_HVT U1636 ( .A1(\ram[3][64] ), .A2(n5358), .A3(data[64]), .A4(n5359), 
        .Y(n893) );
  AO22X1_HVT U1637 ( .A1(\ram[3][63] ), .A2(n5358), .A3(data[63]), .A4(n5359), 
        .Y(n892) );
  AO22X1_HVT U1638 ( .A1(\ram[3][62] ), .A2(n5358), .A3(data[62]), .A4(n5359), 
        .Y(n891) );
  AO22X1_HVT U1639 ( .A1(\ram[3][61] ), .A2(n5358), .A3(data[61]), .A4(n5359), 
        .Y(n890) );
  AO22X1_HVT U1640 ( .A1(\ram[0][28] ), .A2(n5360), .A3(data[28]), .A4(n5361), 
        .Y(n89) );
  AO22X1_HVT U1641 ( .A1(\ram[3][60] ), .A2(n5358), .A3(data[60]), .A4(n5359), 
        .Y(n889) );
  AO22X1_HVT U1642 ( .A1(\ram[3][59] ), .A2(n5358), .A3(data[59]), .A4(n5359), 
        .Y(n888) );
  AO22X1_HVT U1643 ( .A1(\ram[3][58] ), .A2(n5358), .A3(data[58]), .A4(n5359), 
        .Y(n887) );
  AO22X1_HVT U1644 ( .A1(\ram[3][57] ), .A2(n5358), .A3(data[57]), .A4(n5359), 
        .Y(n886) );
  AO22X1_HVT U1645 ( .A1(\ram[3][56] ), .A2(n5358), .A3(data[56]), .A4(n5359), 
        .Y(n885) );
  AO22X1_HVT U1646 ( .A1(\ram[3][55] ), .A2(n5358), .A3(data[55]), .A4(n5359), 
        .Y(n884) );
  AO22X1_HVT U1647 ( .A1(\ram[3][54] ), .A2(n5358), .A3(data[54]), .A4(n5359), 
        .Y(n883) );
  AO22X1_HVT U1648 ( .A1(\ram[3][53] ), .A2(n5358), .A3(data[53]), .A4(n5359), 
        .Y(n882) );
  AO22X1_HVT U1649 ( .A1(\ram[3][52] ), .A2(n5358), .A3(data[52]), .A4(n5359), 
        .Y(n881) );
  AO22X1_HVT U1650 ( .A1(\ram[3][51] ), .A2(n5358), .A3(data[51]), .A4(n5359), 
        .Y(n880) );
  AO22X1_HVT U1651 ( .A1(\ram[0][27] ), .A2(n5360), .A3(data[27]), .A4(n5361), 
        .Y(n88) );
  AO22X1_HVT U1652 ( .A1(\ram[3][50] ), .A2(n5358), .A3(data[50]), .A4(n5359), 
        .Y(n879) );
  AO22X1_HVT U1653 ( .A1(\ram[3][49] ), .A2(n5358), .A3(data[49]), .A4(n5359), 
        .Y(n878) );
  AO22X1_HVT U1654 ( .A1(\ram[3][48] ), .A2(n5358), .A3(data[48]), .A4(n5359), 
        .Y(n877) );
  AO22X1_HVT U1655 ( .A1(\ram[3][47] ), .A2(n5358), .A3(data[47]), .A4(n5359), 
        .Y(n876) );
  AO22X1_HVT U1656 ( .A1(\ram[3][46] ), .A2(n5358), .A3(data[46]), .A4(n5359), 
        .Y(n875) );
  AO22X1_HVT U1657 ( .A1(\ram[3][45] ), .A2(n5358), .A3(data[45]), .A4(n5359), 
        .Y(n874) );
  AO22X1_HVT U1658 ( .A1(\ram[3][44] ), .A2(n5358), .A3(data[44]), .A4(n5359), 
        .Y(n873) );
  AO22X1_HVT U1659 ( .A1(\ram[3][43] ), .A2(n5358), .A3(data[43]), .A4(n5359), 
        .Y(n872) );
  AO22X1_HVT U1660 ( .A1(\ram[3][42] ), .A2(n5358), .A3(data[42]), .A4(n5359), 
        .Y(n871) );
  AO22X1_HVT U1661 ( .A1(\ram[3][41] ), .A2(n5358), .A3(data[41]), .A4(n5359), 
        .Y(n870) );
  AO22X1_HVT U1662 ( .A1(\ram[0][26] ), .A2(n5360), .A3(data[26]), .A4(n5361), 
        .Y(n87) );
  AO22X1_HVT U1663 ( .A1(\ram[3][40] ), .A2(n5358), .A3(data[40]), .A4(n5359), 
        .Y(n869) );
  AO22X1_HVT U1664 ( .A1(\ram[3][39] ), .A2(n5358), .A3(data[39]), .A4(n5359), 
        .Y(n868) );
  AO22X1_HVT U1665 ( .A1(\ram[3][38] ), .A2(n5358), .A3(data[38]), .A4(n5359), 
        .Y(n867) );
  AO22X1_HVT U1666 ( .A1(\ram[3][37] ), .A2(n5358), .A3(data[37]), .A4(n5359), 
        .Y(n866) );
  AO22X1_HVT U1667 ( .A1(\ram[3][36] ), .A2(n5358), .A3(data[36]), .A4(n5359), 
        .Y(n865) );
  AO22X1_HVT U1668 ( .A1(\ram[3][35] ), .A2(n5358), .A3(data[35]), .A4(n5359), 
        .Y(n864) );
  AO22X1_HVT U1669 ( .A1(\ram[3][34] ), .A2(n5358), .A3(data[34]), .A4(n5359), 
        .Y(n863) );
  AO22X1_HVT U1670 ( .A1(\ram[3][33] ), .A2(n5358), .A3(data[33]), .A4(n5359), 
        .Y(n862) );
  AO22X1_HVT U1671 ( .A1(\ram[3][32] ), .A2(n5358), .A3(data[32]), .A4(n5359), 
        .Y(n861) );
  AO22X1_HVT U1672 ( .A1(\ram[3][31] ), .A2(n5358), .A3(data[31]), .A4(n5359), 
        .Y(n860) );
  AO22X1_HVT U1673 ( .A1(\ram[0][25] ), .A2(n5360), .A3(data[25]), .A4(n5361), 
        .Y(n86) );
  AO22X1_HVT U1674 ( .A1(\ram[3][30] ), .A2(n5358), .A3(data[30]), .A4(n5359), 
        .Y(n859) );
  AO22X1_HVT U1675 ( .A1(\ram[3][29] ), .A2(n5358), .A3(data[29]), .A4(n5359), 
        .Y(n858) );
  AO22X1_HVT U1676 ( .A1(\ram[3][28] ), .A2(n5358), .A3(data[28]), .A4(n5359), 
        .Y(n857) );
  AO22X1_HVT U1677 ( .A1(\ram[3][27] ), .A2(n5358), .A3(data[27]), .A4(n5359), 
        .Y(n856) );
  AO22X1_HVT U1678 ( .A1(\ram[3][26] ), .A2(n5358), .A3(data[26]), .A4(n5359), 
        .Y(n855) );
  AO22X1_HVT U1679 ( .A1(\ram[3][25] ), .A2(n5358), .A3(data[25]), .A4(n5359), 
        .Y(n854) );
  AO22X1_HVT U1680 ( .A1(\ram[3][24] ), .A2(n5358), .A3(data[24]), .A4(n5359), 
        .Y(n853) );
  AO22X1_HVT U1681 ( .A1(\ram[3][23] ), .A2(n5358), .A3(data[23]), .A4(n5359), 
        .Y(n852) );
  AO22X1_HVT U1682 ( .A1(\ram[3][22] ), .A2(n5358), .A3(data[22]), .A4(n5359), 
        .Y(n851) );
  AO22X1_HVT U1683 ( .A1(\ram[3][21] ), .A2(n5358), .A3(data[21]), .A4(n5359), 
        .Y(n850) );
  AO22X1_HVT U1684 ( .A1(\ram[0][24] ), .A2(n5360), .A3(data[24]), .A4(n5361), 
        .Y(n85) );
  AO22X1_HVT U1685 ( .A1(\ram[3][20] ), .A2(n5358), .A3(data[20]), .A4(n5359), 
        .Y(n849) );
  AO22X1_HVT U1686 ( .A1(\ram[3][19] ), .A2(n5358), .A3(data[19]), .A4(n5359), 
        .Y(n848) );
  AO22X1_HVT U1687 ( .A1(\ram[3][18] ), .A2(n5358), .A3(data[18]), .A4(n5359), 
        .Y(n847) );
  AO22X1_HVT U1688 ( .A1(\ram[3][17] ), .A2(n5358), .A3(data[17]), .A4(n5359), 
        .Y(n846) );
  AO22X1_HVT U1689 ( .A1(\ram[3][16] ), .A2(n5358), .A3(data[16]), .A4(n5359), 
        .Y(n845) );
  AO22X1_HVT U1690 ( .A1(\ram[3][15] ), .A2(n5358), .A3(data[15]), .A4(n5359), 
        .Y(n844) );
  AO22X1_HVT U1691 ( .A1(\ram[3][14] ), .A2(n5358), .A3(data[14]), .A4(n5359), 
        .Y(n843) );
  AO22X1_HVT U1692 ( .A1(\ram[3][13] ), .A2(n5358), .A3(data[13]), .A4(n5359), 
        .Y(n842) );
  AO22X1_HVT U1693 ( .A1(\ram[3][12] ), .A2(n5358), .A3(data[12]), .A4(n5359), 
        .Y(n841) );
  AO22X1_HVT U1694 ( .A1(\ram[3][11] ), .A2(n5358), .A3(data[11]), .A4(n5359), 
        .Y(n840) );
  AO22X1_HVT U1695 ( .A1(\ram[0][23] ), .A2(n5360), .A3(data[23]), .A4(n5361), 
        .Y(n84) );
  AO22X1_HVT U1696 ( .A1(\ram[3][10] ), .A2(n5358), .A3(data[10]), .A4(n5359), 
        .Y(n839) );
  AO22X1_HVT U1697 ( .A1(\ram[3][9] ), .A2(n5358), .A3(data[9]), .A4(n5359), 
        .Y(n838) );
  AO22X1_HVT U1698 ( .A1(\ram[3][8] ), .A2(n5358), .A3(data[8]), .A4(n5359), 
        .Y(n837) );
  AO22X1_HVT U1699 ( .A1(\ram[3][7] ), .A2(n5358), .A3(data[7]), .A4(n5359), 
        .Y(n836) );
  AO22X1_HVT U1700 ( .A1(\ram[3][6] ), .A2(n5358), .A3(data[6]), .A4(n5359), 
        .Y(n835) );
  AO22X1_HVT U1701 ( .A1(\ram[3][5] ), .A2(n5358), .A3(data[5]), .A4(n5359), 
        .Y(n834) );
  AO22X1_HVT U1702 ( .A1(\ram[3][4] ), .A2(n5358), .A3(data[4]), .A4(n5359), 
        .Y(n833) );
  AO22X1_HVT U1703 ( .A1(\ram[3][3] ), .A2(n5358), .A3(data[3]), .A4(n5359), 
        .Y(n832) );
  AO22X1_HVT U1704 ( .A1(\ram[3][2] ), .A2(n5358), .A3(data[2]), .A4(n5359), 
        .Y(n831) );
  AO22X1_HVT U1705 ( .A1(\ram[3][1] ), .A2(n5358), .A3(data[1]), .A4(n5359), 
        .Y(n830) );
  AO22X1_HVT U1706 ( .A1(\ram[0][22] ), .A2(n5360), .A3(data[22]), .A4(n5361), 
        .Y(n83) );
  AO22X1_HVT U1707 ( .A1(\ram[3][0] ), .A2(n5358), .A3(data[0]), .A4(n5359), 
        .Y(n829) );
  AO22X1_HVT U1708 ( .A1(\ram[2][255] ), .A2(n5362), .A3(data[255]), .A4(n5363), .Y(n828) );
  AO22X1_HVT U1709 ( .A1(\ram[2][254] ), .A2(n5362), .A3(data[254]), .A4(n5363), .Y(n827) );
  AO22X1_HVT U1710 ( .A1(\ram[2][253] ), .A2(n5362), .A3(data[253]), .A4(n5363), .Y(n826) );
  AO22X1_HVT U1711 ( .A1(\ram[2][252] ), .A2(n5362), .A3(data[252]), .A4(n5363), .Y(n825) );
  AO22X1_HVT U1712 ( .A1(\ram[2][251] ), .A2(n5362), .A3(data[251]), .A4(n5363), .Y(n824) );
  AO22X1_HVT U1713 ( .A1(\ram[2][250] ), .A2(n5362), .A3(data[250]), .A4(n5363), .Y(n823) );
  AO22X1_HVT U1714 ( .A1(\ram[2][249] ), .A2(n5362), .A3(data[249]), .A4(n5363), .Y(n822) );
  AO22X1_HVT U1715 ( .A1(\ram[2][248] ), .A2(n5362), .A3(data[248]), .A4(n5363), .Y(n821) );
  AO22X1_HVT U1716 ( .A1(\ram[2][247] ), .A2(n5362), .A3(data[247]), .A4(n5363), .Y(n820) );
  AO22X1_HVT U1717 ( .A1(\ram[0][21] ), .A2(n5360), .A3(data[21]), .A4(n5361), 
        .Y(n82) );
  AO22X1_HVT U1718 ( .A1(\ram[2][246] ), .A2(n5362), .A3(data[246]), .A4(n5363), .Y(n819) );
  AO22X1_HVT U1719 ( .A1(\ram[2][245] ), .A2(n5362), .A3(data[245]), .A4(n5363), .Y(n818) );
  AO22X1_HVT U1720 ( .A1(\ram[2][244] ), .A2(n5362), .A3(data[244]), .A4(n5363), .Y(n817) );
  AO22X1_HVT U1721 ( .A1(\ram[2][243] ), .A2(n5362), .A3(data[243]), .A4(n5363), .Y(n816) );
  AO22X1_HVT U1722 ( .A1(\ram[2][242] ), .A2(n5362), .A3(data[242]), .A4(n5363), .Y(n815) );
  AO22X1_HVT U1723 ( .A1(\ram[2][241] ), .A2(n5362), .A3(data[241]), .A4(n5363), .Y(n814) );
  AO22X1_HVT U1724 ( .A1(\ram[2][240] ), .A2(n5362), .A3(data[240]), .A4(n5363), .Y(n813) );
  AO22X1_HVT U1725 ( .A1(\ram[2][239] ), .A2(n5362), .A3(data[239]), .A4(n5363), .Y(n812) );
  AO22X1_HVT U1726 ( .A1(\ram[2][238] ), .A2(n5362), .A3(data[238]), .A4(n5363), .Y(n811) );
  AO22X1_HVT U1727 ( .A1(\ram[2][237] ), .A2(n5362), .A3(data[237]), .A4(n5363), .Y(n810) );
  AO22X1_HVT U1728 ( .A1(\ram[0][20] ), .A2(n5360), .A3(data[20]), .A4(n5361), 
        .Y(n81) );
  AO22X1_HVT U1729 ( .A1(\ram[2][236] ), .A2(n5362), .A3(data[236]), .A4(n5363), .Y(n809) );
  AO22X1_HVT U1730 ( .A1(\ram[2][235] ), .A2(n5362), .A3(data[235]), .A4(n5363), .Y(n808) );
  AO22X1_HVT U1731 ( .A1(\ram[2][234] ), .A2(n5362), .A3(data[234]), .A4(n5363), .Y(n807) );
  AO22X1_HVT U1732 ( .A1(\ram[2][233] ), .A2(n5362), .A3(data[233]), .A4(n5363), .Y(n806) );
  AO22X1_HVT U1733 ( .A1(\ram[2][232] ), .A2(n5362), .A3(data[232]), .A4(n5363), .Y(n805) );
  AO22X1_HVT U1734 ( .A1(\ram[2][231] ), .A2(n5362), .A3(data[231]), .A4(n5363), .Y(n804) );
  AO22X1_HVT U1735 ( .A1(\ram[2][230] ), .A2(n5362), .A3(data[230]), .A4(n5363), .Y(n803) );
  AO22X1_HVT U1736 ( .A1(\ram[2][229] ), .A2(n5362), .A3(data[229]), .A4(n5363), .Y(n802) );
  AO22X1_HVT U1737 ( .A1(\ram[2][228] ), .A2(n5362), .A3(data[228]), .A4(n5363), .Y(n801) );
  AO22X1_HVT U1738 ( .A1(\ram[2][227] ), .A2(n5362), .A3(data[227]), .A4(n5363), .Y(n800) );
  AO22X1_HVT U1739 ( .A1(\ram[0][19] ), .A2(n5360), .A3(data[19]), .A4(n5361), 
        .Y(n80) );
  AO22X1_HVT U1740 ( .A1(\ram[2][226] ), .A2(n5362), .A3(data[226]), .A4(n5363), .Y(n799) );
  AO22X1_HVT U1741 ( .A1(\ram[2][225] ), .A2(n5362), .A3(data[225]), .A4(n5363), .Y(n798) );
  AO22X1_HVT U1742 ( .A1(\ram[2][224] ), .A2(n5362), .A3(data[224]), .A4(n5363), .Y(n797) );
  AO22X1_HVT U1743 ( .A1(\ram[2][223] ), .A2(n5362), .A3(data[223]), .A4(n5363), .Y(n796) );
  AO22X1_HVT U1744 ( .A1(\ram[2][222] ), .A2(n5362), .A3(data[222]), .A4(n5363), .Y(n795) );
  AO22X1_HVT U1745 ( .A1(\ram[2][221] ), .A2(n5362), .A3(data[221]), .A4(n5363), .Y(n794) );
  AO22X1_HVT U1746 ( .A1(\ram[2][220] ), .A2(n5362), .A3(data[220]), .A4(n5363), .Y(n793) );
  AO22X1_HVT U1747 ( .A1(\ram[2][219] ), .A2(n5362), .A3(data[219]), .A4(n5363), .Y(n792) );
  AO22X1_HVT U1748 ( .A1(\ram[2][218] ), .A2(n5362), .A3(data[218]), .A4(n5363), .Y(n791) );
  AO22X1_HVT U1749 ( .A1(\ram[2][217] ), .A2(n5362), .A3(data[217]), .A4(n5363), .Y(n790) );
  AO22X1_HVT U1750 ( .A1(\ram[0][18] ), .A2(n5360), .A3(data[18]), .A4(n5361), 
        .Y(n79) );
  AO22X1_HVT U1751 ( .A1(\ram[2][216] ), .A2(n5362), .A3(data[216]), .A4(n5363), .Y(n789) );
  AO22X1_HVT U1752 ( .A1(\ram[2][215] ), .A2(n5362), .A3(data[215]), .A4(n5363), .Y(n788) );
  AO22X1_HVT U1753 ( .A1(\ram[2][214] ), .A2(n5362), .A3(data[214]), .A4(n5363), .Y(n787) );
  AO22X1_HVT U1754 ( .A1(\ram[2][213] ), .A2(n5362), .A3(data[213]), .A4(n5363), .Y(n786) );
  AO22X1_HVT U1755 ( .A1(\ram[2][212] ), .A2(n5362), .A3(data[212]), .A4(n5363), .Y(n785) );
  AO22X1_HVT U1756 ( .A1(\ram[2][211] ), .A2(n5362), .A3(data[211]), .A4(n5363), .Y(n784) );
  AO22X1_HVT U1757 ( .A1(\ram[2][210] ), .A2(n5362), .A3(data[210]), .A4(n5363), .Y(n783) );
  AO22X1_HVT U1758 ( .A1(\ram[2][209] ), .A2(n5362), .A3(data[209]), .A4(n5363), .Y(n782) );
  AO22X1_HVT U1759 ( .A1(\ram[2][208] ), .A2(n5362), .A3(data[208]), .A4(n5363), .Y(n781) );
  AO22X1_HVT U1760 ( .A1(\ram[2][207] ), .A2(n5362), .A3(data[207]), .A4(n5363), .Y(n780) );
  AO22X1_HVT U1761 ( .A1(\ram[0][17] ), .A2(n5360), .A3(data[17]), .A4(n5361), 
        .Y(n78) );
  AO22X1_HVT U1762 ( .A1(\ram[2][206] ), .A2(n5362), .A3(data[206]), .A4(n5363), .Y(n779) );
  AO22X1_HVT U1763 ( .A1(\ram[2][205] ), .A2(n5362), .A3(data[205]), .A4(n5363), .Y(n778) );
  AO22X1_HVT U1764 ( .A1(\ram[2][204] ), .A2(n5362), .A3(data[204]), .A4(n5363), .Y(n777) );
  AO22X1_HVT U1765 ( .A1(\ram[2][203] ), .A2(n5362), .A3(data[203]), .A4(n5363), .Y(n776) );
  AO22X1_HVT U1766 ( .A1(\ram[2][202] ), .A2(n5362), .A3(data[202]), .A4(n5363), .Y(n775) );
  AO22X1_HVT U1767 ( .A1(\ram[2][201] ), .A2(n5362), .A3(data[201]), .A4(n5363), .Y(n774) );
  AO22X1_HVT U1768 ( .A1(\ram[2][200] ), .A2(n5362), .A3(data[200]), .A4(n5363), .Y(n773) );
  AO22X1_HVT U1769 ( .A1(\ram[2][199] ), .A2(n5362), .A3(data[199]), .A4(n5363), .Y(n772) );
  AO22X1_HVT U1770 ( .A1(\ram[2][198] ), .A2(n5362), .A3(data[198]), .A4(n5363), .Y(n771) );
  AO22X1_HVT U1771 ( .A1(\ram[2][197] ), .A2(n5362), .A3(data[197]), .A4(n5363), .Y(n770) );
  AO22X1_HVT U1772 ( .A1(\ram[0][16] ), .A2(n5360), .A3(data[16]), .A4(n5361), 
        .Y(n77) );
  AO22X1_HVT U1773 ( .A1(\ram[2][196] ), .A2(n5362), .A3(data[196]), .A4(n5363), .Y(n769) );
  AO22X1_HVT U1774 ( .A1(\ram[2][195] ), .A2(n5362), .A3(data[195]), .A4(n5363), .Y(n768) );
  AO22X1_HVT U1775 ( .A1(\ram[2][194] ), .A2(n5362), .A3(data[194]), .A4(n5363), .Y(n767) );
  AO22X1_HVT U1776 ( .A1(\ram[2][193] ), .A2(n5362), .A3(data[193]), .A4(n5363), .Y(n766) );
  AO22X1_HVT U1777 ( .A1(\ram[2][192] ), .A2(n5362), .A3(data[192]), .A4(n5363), .Y(n765) );
  AO22X1_HVT U1778 ( .A1(\ram[2][191] ), .A2(n5362), .A3(data[191]), .A4(n5363), .Y(n764) );
  AO22X1_HVT U1779 ( .A1(\ram[2][190] ), .A2(n5362), .A3(data[190]), .A4(n5363), .Y(n763) );
  AO22X1_HVT U1780 ( .A1(\ram[2][189] ), .A2(n5362), .A3(data[189]), .A4(n5363), .Y(n762) );
  AO22X1_HVT U1781 ( .A1(\ram[2][188] ), .A2(n5362), .A3(data[188]), .A4(n5363), .Y(n761) );
  AO22X1_HVT U1782 ( .A1(\ram[2][187] ), .A2(n5362), .A3(data[187]), .A4(n5363), .Y(n760) );
  AO22X1_HVT U1783 ( .A1(\ram[0][15] ), .A2(n5360), .A3(data[15]), .A4(n5361), 
        .Y(n76) );
  AO22X1_HVT U1784 ( .A1(\ram[2][186] ), .A2(n5362), .A3(data[186]), .A4(n5363), .Y(n759) );
  AO22X1_HVT U1785 ( .A1(\ram[2][185] ), .A2(n5362), .A3(data[185]), .A4(n5363), .Y(n758) );
  AO22X1_HVT U1786 ( .A1(\ram[2][184] ), .A2(n5362), .A3(data[184]), .A4(n5363), .Y(n757) );
  AO22X1_HVT U1787 ( .A1(\ram[2][183] ), .A2(n5362), .A3(data[183]), .A4(n5363), .Y(n756) );
  AO22X1_HVT U1788 ( .A1(\ram[2][182] ), .A2(n5362), .A3(data[182]), .A4(n5363), .Y(n755) );
  AO22X1_HVT U1789 ( .A1(\ram[2][181] ), .A2(n5362), .A3(data[181]), .A4(n5363), .Y(n754) );
  AO22X1_HVT U1790 ( .A1(\ram[2][180] ), .A2(n5362), .A3(data[180]), .A4(n5363), .Y(n753) );
  AO22X1_HVT U1791 ( .A1(\ram[2][179] ), .A2(n5362), .A3(data[179]), .A4(n5363), .Y(n752) );
  AO22X1_HVT U1792 ( .A1(\ram[2][178] ), .A2(n5362), .A3(data[178]), .A4(n5363), .Y(n751) );
  AO22X1_HVT U1793 ( .A1(\ram[2][177] ), .A2(n5362), .A3(data[177]), .A4(n5363), .Y(n750) );
  AO22X1_HVT U1794 ( .A1(\ram[0][14] ), .A2(n5360), .A3(data[14]), .A4(n5361), 
        .Y(n75) );
  AO22X1_HVT U1795 ( .A1(\ram[2][176] ), .A2(n5362), .A3(data[176]), .A4(n5363), .Y(n749) );
  AO22X1_HVT U1796 ( .A1(\ram[2][175] ), .A2(n5362), .A3(data[175]), .A4(n5363), .Y(n748) );
  AO22X1_HVT U1797 ( .A1(\ram[2][174] ), .A2(n5362), .A3(data[174]), .A4(n5363), .Y(n747) );
  AO22X1_HVT U1798 ( .A1(\ram[2][173] ), .A2(n5362), .A3(data[173]), .A4(n5363), .Y(n746) );
  AO22X1_HVT U1799 ( .A1(\ram[2][172] ), .A2(n5362), .A3(data[172]), .A4(n5363), .Y(n745) );
  AO22X1_HVT U1800 ( .A1(\ram[2][171] ), .A2(n5362), .A3(data[171]), .A4(n5363), .Y(n744) );
  AO22X1_HVT U1801 ( .A1(\ram[2][170] ), .A2(n5362), .A3(n5363), .A4(data[170]), .Y(n743) );
  AO22X1_HVT U1802 ( .A1(\ram[2][169] ), .A2(n5362), .A3(n5363), .A4(data[169]), .Y(n742) );
  AO22X1_HVT U1803 ( .A1(\ram[2][168] ), .A2(n5362), .A3(n5363), .A4(data[168]), .Y(n741) );
  AO22X1_HVT U1804 ( .A1(\ram[2][167] ), .A2(n5362), .A3(n5363), .A4(data[167]), .Y(n740) );
  AO22X1_HVT U1805 ( .A1(\ram[0][13] ), .A2(n5360), .A3(data[13]), .A4(n5361), 
        .Y(n74) );
  AO22X1_HVT U1806 ( .A1(\ram[2][166] ), .A2(n5362), .A3(n5363), .A4(data[166]), .Y(n739) );
  AO22X1_HVT U1807 ( .A1(\ram[2][165] ), .A2(n5362), .A3(n5363), .A4(data[165]), .Y(n738) );
  AO22X1_HVT U1808 ( .A1(\ram[2][164] ), .A2(n5362), .A3(n5363), .A4(data[164]), .Y(n737) );
  AO22X1_HVT U1809 ( .A1(\ram[2][163] ), .A2(n5362), .A3(n5363), .A4(data[163]), .Y(n736) );
  AO22X1_HVT U1810 ( .A1(\ram[2][162] ), .A2(n5362), .A3(n5363), .A4(data[162]), .Y(n735) );
  AO22X1_HVT U1811 ( .A1(\ram[2][161] ), .A2(n5362), .A3(n5363), .A4(data[161]), .Y(n734) );
  AO22X1_HVT U1812 ( .A1(\ram[2][160] ), .A2(n5362), .A3(n5363), .A4(data[160]), .Y(n733) );
  AO22X1_HVT U1813 ( .A1(\ram[2][159] ), .A2(n5362), .A3(n5363), .A4(data[159]), .Y(n732) );
  AO22X1_HVT U1814 ( .A1(\ram[2][158] ), .A2(n5362), .A3(n5363), .A4(data[158]), .Y(n731) );
  AO22X1_HVT U1815 ( .A1(\ram[2][157] ), .A2(n5362), .A3(n5363), .A4(data[157]), .Y(n730) );
  AO22X1_HVT U1816 ( .A1(\ram[0][12] ), .A2(n5360), .A3(data[12]), .A4(n5361), 
        .Y(n73) );
  AO22X1_HVT U1817 ( .A1(\ram[2][156] ), .A2(n5362), .A3(n5363), .A4(data[156]), .Y(n729) );
  AO22X1_HVT U1818 ( .A1(\ram[2][155] ), .A2(n5362), .A3(n5363), .A4(data[155]), .Y(n728) );
  AO22X1_HVT U1819 ( .A1(\ram[2][154] ), .A2(n5362), .A3(n5363), .A4(data[154]), .Y(n727) );
  AO22X1_HVT U1820 ( .A1(\ram[2][153] ), .A2(n5362), .A3(n5363), .A4(data[153]), .Y(n726) );
  AO22X1_HVT U1821 ( .A1(\ram[2][152] ), .A2(n5362), .A3(n5363), .A4(data[152]), .Y(n725) );
  AO22X1_HVT U1822 ( .A1(\ram[2][151] ), .A2(n5362), .A3(n5363), .A4(data[151]), .Y(n724) );
  AO22X1_HVT U1823 ( .A1(\ram[2][150] ), .A2(n5362), .A3(n5363), .A4(data[150]), .Y(n723) );
  AO22X1_HVT U1824 ( .A1(\ram[2][149] ), .A2(n5362), .A3(n5363), .A4(data[149]), .Y(n722) );
  AO22X1_HVT U1825 ( .A1(\ram[2][148] ), .A2(n5362), .A3(n5363), .A4(data[148]), .Y(n721) );
  AO22X1_HVT U1826 ( .A1(\ram[2][147] ), .A2(n5362), .A3(n5363), .A4(data[147]), .Y(n720) );
  AO22X1_HVT U1827 ( .A1(\ram[0][11] ), .A2(n5360), .A3(data[11]), .A4(n5361), 
        .Y(n72) );
  AO22X1_HVT U1828 ( .A1(\ram[2][146] ), .A2(n5362), .A3(n5363), .A4(data[146]), .Y(n719) );
  AO22X1_HVT U1829 ( .A1(\ram[2][145] ), .A2(n5362), .A3(n5363), .A4(data[145]), .Y(n718) );
  AO22X1_HVT U1830 ( .A1(\ram[2][144] ), .A2(n5362), .A3(n5363), .A4(data[144]), .Y(n717) );
  AO22X1_HVT U1831 ( .A1(\ram[2][143] ), .A2(n5362), .A3(n5363), .A4(data[143]), .Y(n716) );
  AO22X1_HVT U1832 ( .A1(\ram[2][142] ), .A2(n5362), .A3(n5363), .A4(data[142]), .Y(n715) );
  AO22X1_HVT U1833 ( .A1(\ram[2][141] ), .A2(n5362), .A3(n5363), .A4(data[141]), .Y(n714) );
  AO22X1_HVT U1834 ( .A1(\ram[2][140] ), .A2(n5362), .A3(n5363), .A4(data[140]), .Y(n713) );
  AO22X1_HVT U1835 ( .A1(\ram[2][139] ), .A2(n5362), .A3(n5363), .A4(data[139]), .Y(n712) );
  AO22X1_HVT U1836 ( .A1(\ram[2][138] ), .A2(n5362), .A3(n5363), .A4(data[138]), .Y(n711) );
  AO22X1_HVT U1837 ( .A1(\ram[2][137] ), .A2(n5362), .A3(n5363), .A4(data[137]), .Y(n710) );
  AO22X1_HVT U1838 ( .A1(\ram[0][10] ), .A2(n5360), .A3(data[10]), .A4(n5361), 
        .Y(n71) );
  AO22X1_HVT U1839 ( .A1(\ram[2][136] ), .A2(n5362), .A3(n5363), .A4(data[136]), .Y(n709) );
  AO22X1_HVT U1840 ( .A1(\ram[2][135] ), .A2(n5362), .A3(n5363), .A4(data[135]), .Y(n708) );
  AO22X1_HVT U1841 ( .A1(\ram[2][134] ), .A2(n5362), .A3(n5363), .A4(data[134]), .Y(n707) );
  AO22X1_HVT U1842 ( .A1(\ram[2][133] ), .A2(n5362), .A3(n5363), .A4(data[133]), .Y(n706) );
  AO22X1_HVT U1843 ( .A1(\ram[2][132] ), .A2(n5362), .A3(n5363), .A4(data[132]), .Y(n705) );
  AO22X1_HVT U1844 ( .A1(\ram[2][131] ), .A2(n5362), .A3(n5363), .A4(data[131]), .Y(n704) );
  AO22X1_HVT U1845 ( .A1(\ram[2][130] ), .A2(n5362), .A3(n5363), .A4(data[130]), .Y(n703) );
  AO22X1_HVT U1846 ( .A1(\ram[2][129] ), .A2(n5362), .A3(n5363), .A4(data[129]), .Y(n702) );
  AO22X1_HVT U1847 ( .A1(\ram[2][128] ), .A2(n5362), .A3(n5363), .A4(data[128]), .Y(n701) );
  AO22X1_HVT U1848 ( .A1(\ram[2][127] ), .A2(n5362), .A3(n5363), .A4(data[127]), .Y(n700) );
  AO22X1_HVT U1849 ( .A1(\ram[0][9] ), .A2(n5360), .A3(data[9]), .A4(n5361), 
        .Y(n70) );
  AO22X1_HVT U1850 ( .A1(\ram[2][126] ), .A2(n5362), .A3(n5363), .A4(data[126]), .Y(n699) );
  AO22X1_HVT U1851 ( .A1(\ram[2][125] ), .A2(n5362), .A3(n5363), .A4(data[125]), .Y(n698) );
  AO22X1_HVT U1852 ( .A1(\ram[2][124] ), .A2(n5362), .A3(n5363), .A4(data[124]), .Y(n697) );
  AO22X1_HVT U1853 ( .A1(\ram[2][123] ), .A2(n5362), .A3(n5363), .A4(data[123]), .Y(n696) );
  AO22X1_HVT U1854 ( .A1(\ram[2][122] ), .A2(n5362), .A3(n5363), .A4(data[122]), .Y(n695) );
  AO22X1_HVT U1855 ( .A1(\ram[2][121] ), .A2(n5362), .A3(n5363), .A4(data[121]), .Y(n694) );
  AO22X1_HVT U1856 ( .A1(\ram[2][120] ), .A2(n5362), .A3(n5363), .A4(data[120]), .Y(n693) );
  AO22X1_HVT U1857 ( .A1(\ram[2][119] ), .A2(n5362), .A3(n5363), .A4(data[119]), .Y(n692) );
  AO22X1_HVT U1858 ( .A1(\ram[2][118] ), .A2(n5362), .A3(n5363), .A4(data[118]), .Y(n691) );
  AO22X1_HVT U1859 ( .A1(\ram[2][117] ), .A2(n5362), .A3(n5363), .A4(data[117]), .Y(n690) );
  AO22X1_HVT U1860 ( .A1(\ram[0][8] ), .A2(n5360), .A3(data[8]), .A4(n5361), 
        .Y(n69) );
  AO22X1_HVT U1861 ( .A1(\ram[2][116] ), .A2(n5362), .A3(n5363), .A4(data[116]), .Y(n689) );
  AO22X1_HVT U1862 ( .A1(\ram[2][115] ), .A2(n5362), .A3(n5363), .A4(data[115]), .Y(n688) );
  AO22X1_HVT U1863 ( .A1(\ram[2][114] ), .A2(n5362), .A3(n5363), .A4(data[114]), .Y(n687) );
  AO22X1_HVT U1864 ( .A1(\ram[2][113] ), .A2(n5362), .A3(n5363), .A4(data[113]), .Y(n686) );
  AO22X1_HVT U1865 ( .A1(\ram[2][112] ), .A2(n5362), .A3(n5363), .A4(data[112]), .Y(n685) );
  AO22X1_HVT U1866 ( .A1(\ram[2][111] ), .A2(n5362), .A3(n5363), .A4(data[111]), .Y(n684) );
  AO22X1_HVT U1867 ( .A1(\ram[2][110] ), .A2(n5362), .A3(n5363), .A4(data[110]), .Y(n683) );
  AO22X1_HVT U1868 ( .A1(\ram[2][109] ), .A2(n5362), .A3(n5363), .A4(data[109]), .Y(n682) );
  AO22X1_HVT U1869 ( .A1(\ram[2][108] ), .A2(n5362), .A3(n5363), .A4(data[108]), .Y(n681) );
  AO22X1_HVT U1870 ( .A1(\ram[2][107] ), .A2(n5362), .A3(n5363), .A4(data[107]), .Y(n680) );
  AO22X1_HVT U1871 ( .A1(\ram[0][7] ), .A2(n5360), .A3(data[7]), .A4(n5361), 
        .Y(n68) );
  AO22X1_HVT U1872 ( .A1(\ram[2][106] ), .A2(n5362), .A3(n5363), .A4(data[106]), .Y(n679) );
  AO22X1_HVT U1873 ( .A1(\ram[2][105] ), .A2(n5362), .A3(n5363), .A4(data[105]), .Y(n678) );
  AO22X1_HVT U1874 ( .A1(\ram[2][104] ), .A2(n5362), .A3(n5363), .A4(data[104]), .Y(n677) );
  AO22X1_HVT U1875 ( .A1(\ram[2][103] ), .A2(n5362), .A3(n5363), .A4(data[103]), .Y(n676) );
  AO22X1_HVT U1876 ( .A1(\ram[2][102] ), .A2(n5362), .A3(n5363), .A4(data[102]), .Y(n675) );
  AO22X1_HVT U1877 ( .A1(\ram[2][101] ), .A2(n5362), .A3(n5363), .A4(data[101]), .Y(n674) );
  AO22X1_HVT U1878 ( .A1(\ram[2][100] ), .A2(n5362), .A3(n5363), .A4(data[100]), .Y(n673) );
  AO22X1_HVT U1879 ( .A1(\ram[2][99] ), .A2(n5362), .A3(n5363), .A4(data[99]), 
        .Y(n672) );
  AO22X1_HVT U1880 ( .A1(\ram[2][98] ), .A2(n5362), .A3(n5363), .A4(data[98]), 
        .Y(n671) );
  AO22X1_HVT U1881 ( .A1(\ram[2][97] ), .A2(n5362), .A3(n5363), .A4(data[97]), 
        .Y(n670) );
  AO22X1_HVT U1882 ( .A1(\ram[0][6] ), .A2(n5360), .A3(data[6]), .A4(n5361), 
        .Y(n67) );
  AO22X1_HVT U1883 ( .A1(\ram[2][96] ), .A2(n5362), .A3(n5363), .A4(data[96]), 
        .Y(n669) );
  AO22X1_HVT U1884 ( .A1(\ram[2][95] ), .A2(n5362), .A3(n5363), .A4(data[95]), 
        .Y(n668) );
  AO22X1_HVT U1885 ( .A1(\ram[2][94] ), .A2(n5362), .A3(n5363), .A4(data[94]), 
        .Y(n667) );
  AO22X1_HVT U1886 ( .A1(\ram[2][93] ), .A2(n5362), .A3(n5363), .A4(data[93]), 
        .Y(n666) );
  AO22X1_HVT U1887 ( .A1(\ram[2][92] ), .A2(n5362), .A3(n5363), .A4(data[92]), 
        .Y(n665) );
  AO22X1_HVT U1888 ( .A1(\ram[2][91] ), .A2(n5362), .A3(n5363), .A4(data[91]), 
        .Y(n664) );
  AO22X1_HVT U1889 ( .A1(\ram[2][90] ), .A2(n5362), .A3(n5363), .A4(data[90]), 
        .Y(n663) );
  AO22X1_HVT U1890 ( .A1(\ram[2][89] ), .A2(n5362), .A3(n5363), .A4(data[89]), 
        .Y(n662) );
  AO22X1_HVT U1891 ( .A1(\ram[2][88] ), .A2(n5362), .A3(n5363), .A4(data[88]), 
        .Y(n661) );
  AO22X1_HVT U1892 ( .A1(\ram[2][87] ), .A2(n5362), .A3(n5363), .A4(data[87]), 
        .Y(n660) );
  AO22X1_HVT U1893 ( .A1(\ram[0][5] ), .A2(n5360), .A3(data[5]), .A4(n5361), 
        .Y(n66) );
  AO22X1_HVT U1894 ( .A1(\ram[2][86] ), .A2(n5362), .A3(n5363), .A4(data[86]), 
        .Y(n659) );
  AO22X1_HVT U1895 ( .A1(\ram[2][85] ), .A2(n5362), .A3(n5363), .A4(data[85]), 
        .Y(n658) );
  AO22X1_HVT U1896 ( .A1(\ram[2][84] ), .A2(n5362), .A3(n5363), .A4(data[84]), 
        .Y(n657) );
  AO22X1_HVT U1897 ( .A1(\ram[2][83] ), .A2(n5362), .A3(n5363), .A4(data[83]), 
        .Y(n656) );
  AO22X1_HVT U1898 ( .A1(\ram[2][82] ), .A2(n5362), .A3(n5363), .A4(data[82]), 
        .Y(n655) );
  AO22X1_HVT U1899 ( .A1(\ram[2][81] ), .A2(n5362), .A3(n5363), .A4(data[81]), 
        .Y(n654) );
  AO22X1_HVT U1900 ( .A1(\ram[2][80] ), .A2(n5362), .A3(n5363), .A4(data[80]), 
        .Y(n653) );
  AO22X1_HVT U1901 ( .A1(\ram[2][79] ), .A2(n5362), .A3(n5363), .A4(data[79]), 
        .Y(n652) );
  AO22X1_HVT U1902 ( .A1(\ram[2][78] ), .A2(n5362), .A3(n5363), .A4(data[78]), 
        .Y(n651) );
  AO22X1_HVT U1903 ( .A1(\ram[2][77] ), .A2(n5362), .A3(n5363), .A4(data[77]), 
        .Y(n650) );
  AO22X1_HVT U1904 ( .A1(\ram[0][4] ), .A2(n5360), .A3(data[4]), .A4(n5361), 
        .Y(n65) );
  AO22X1_HVT U1905 ( .A1(\ram[2][76] ), .A2(n5362), .A3(n5363), .A4(data[76]), 
        .Y(n649) );
  AO22X1_HVT U1906 ( .A1(\ram[2][75] ), .A2(n5362), .A3(n5363), .A4(data[75]), 
        .Y(n648) );
  AO22X1_HVT U1907 ( .A1(\ram[2][74] ), .A2(n5362), .A3(n5363), .A4(data[74]), 
        .Y(n647) );
  AO22X1_HVT U1908 ( .A1(\ram[2][73] ), .A2(n5362), .A3(n5363), .A4(data[73]), 
        .Y(n646) );
  AO22X1_HVT U1909 ( .A1(\ram[2][72] ), .A2(n5362), .A3(n5363), .A4(data[72]), 
        .Y(n645) );
  AO22X1_HVT U1910 ( .A1(\ram[2][71] ), .A2(n5362), .A3(n5363), .A4(data[71]), 
        .Y(n644) );
  AO22X1_HVT U1911 ( .A1(\ram[2][70] ), .A2(n5362), .A3(n5363), .A4(data[70]), 
        .Y(n643) );
  AO22X1_HVT U1912 ( .A1(\ram[2][69] ), .A2(n5362), .A3(n5363), .A4(data[69]), 
        .Y(n642) );
  AO22X1_HVT U1913 ( .A1(\ram[2][68] ), .A2(n5362), .A3(n5363), .A4(data[68]), 
        .Y(n641) );
  AO22X1_HVT U1914 ( .A1(\ram[2][67] ), .A2(n5362), .A3(n5363), .A4(data[67]), 
        .Y(n640) );
  AO22X1_HVT U1915 ( .A1(\ram[0][3] ), .A2(n5360), .A3(data[3]), .A4(n5361), 
        .Y(n64) );
  AO22X1_HVT U1916 ( .A1(\ram[2][66] ), .A2(n5362), .A3(n5363), .A4(data[66]), 
        .Y(n639) );
  AO22X1_HVT U1917 ( .A1(\ram[2][65] ), .A2(n5362), .A3(n5363), .A4(data[65]), 
        .Y(n638) );
  AO22X1_HVT U1918 ( .A1(\ram[2][64] ), .A2(n5362), .A3(n5363), .A4(data[64]), 
        .Y(n637) );
  AO22X1_HVT U1919 ( .A1(\ram[2][63] ), .A2(n5362), .A3(n5363), .A4(data[63]), 
        .Y(n636) );
  AO22X1_HVT U1920 ( .A1(\ram[2][62] ), .A2(n5362), .A3(n5363), .A4(data[62]), 
        .Y(n635) );
  AO22X1_HVT U1921 ( .A1(\ram[2][61] ), .A2(n5362), .A3(n5363), .A4(data[61]), 
        .Y(n634) );
  AO22X1_HVT U1922 ( .A1(\ram[2][60] ), .A2(n5362), .A3(n5363), .A4(data[60]), 
        .Y(n633) );
  AO22X1_HVT U1923 ( .A1(\ram[2][59] ), .A2(n5362), .A3(n5363), .A4(data[59]), 
        .Y(n632) );
  AO22X1_HVT U1924 ( .A1(\ram[2][58] ), .A2(n5362), .A3(n5363), .A4(data[58]), 
        .Y(n631) );
  AO22X1_HVT U1925 ( .A1(\ram[2][57] ), .A2(n5362), .A3(n5363), .A4(data[57]), 
        .Y(n630) );
  AO22X1_HVT U1926 ( .A1(\ram[0][2] ), .A2(n5360), .A3(data[2]), .A4(n5361), 
        .Y(n63) );
  AO22X1_HVT U1927 ( .A1(\ram[2][56] ), .A2(n5362), .A3(n5363), .A4(data[56]), 
        .Y(n629) );
  AO22X1_HVT U1928 ( .A1(\ram[2][55] ), .A2(n5362), .A3(n5363), .A4(data[55]), 
        .Y(n628) );
  AO22X1_HVT U1929 ( .A1(\ram[2][54] ), .A2(n5362), .A3(n5363), .A4(data[54]), 
        .Y(n627) );
  AO22X1_HVT U1930 ( .A1(\ram[2][53] ), .A2(n5362), .A3(n5363), .A4(data[53]), 
        .Y(n626) );
  AO22X1_HVT U1931 ( .A1(\ram[2][52] ), .A2(n5362), .A3(n5363), .A4(data[52]), 
        .Y(n625) );
  AO22X1_HVT U1932 ( .A1(\ram[2][51] ), .A2(n5362), .A3(n5363), .A4(data[51]), 
        .Y(n624) );
  AO22X1_HVT U1933 ( .A1(\ram[2][50] ), .A2(n5362), .A3(n5363), .A4(data[50]), 
        .Y(n623) );
  AO22X1_HVT U1934 ( .A1(\ram[2][49] ), .A2(n5362), .A3(n5363), .A4(data[49]), 
        .Y(n622) );
  AO22X1_HVT U1935 ( .A1(\ram[2][48] ), .A2(n5362), .A3(n5363), .A4(data[48]), 
        .Y(n621) );
  AO22X1_HVT U1936 ( .A1(\ram[2][47] ), .A2(n5362), .A3(n5363), .A4(data[47]), 
        .Y(n620) );
  AO22X1_HVT U1937 ( .A1(\ram[0][1] ), .A2(n5360), .A3(data[1]), .A4(n5361), 
        .Y(n62) );
  AO22X1_HVT U1938 ( .A1(\ram[2][46] ), .A2(n5362), .A3(n5363), .A4(data[46]), 
        .Y(n619) );
  AO22X1_HVT U1939 ( .A1(\ram[2][45] ), .A2(n5362), .A3(n5363), .A4(data[45]), 
        .Y(n618) );
  AO22X1_HVT U1940 ( .A1(\ram[2][44] ), .A2(n5362), .A3(n5363), .A4(data[44]), 
        .Y(n617) );
  AO22X1_HVT U1941 ( .A1(\ram[2][43] ), .A2(n5362), .A3(n5363), .A4(data[43]), 
        .Y(n616) );
  AO22X1_HVT U1942 ( .A1(\ram[2][42] ), .A2(n5362), .A3(n5363), .A4(data[42]), 
        .Y(n615) );
  AO22X1_HVT U1943 ( .A1(\ram[2][41] ), .A2(n5362), .A3(n5363), .A4(data[41]), 
        .Y(n614) );
  AO22X1_HVT U1944 ( .A1(\ram[2][40] ), .A2(n5362), .A3(n5363), .A4(data[40]), 
        .Y(n613) );
  AO22X1_HVT U1945 ( .A1(\ram[2][39] ), .A2(n5362), .A3(n5363), .A4(data[39]), 
        .Y(n612) );
  AO22X1_HVT U1946 ( .A1(\ram[2][38] ), .A2(n5362), .A3(n5363), .A4(data[38]), 
        .Y(n611) );
  AO22X1_HVT U1947 ( .A1(\ram[2][37] ), .A2(n5362), .A3(n5363), .A4(data[37]), 
        .Y(n610) );
  AO22X1_HVT U1948 ( .A1(\ram[0][0] ), .A2(n5360), .A3(data[0]), .A4(n5361), 
        .Y(n61) );
  AO22X1_HVT U1949 ( .A1(\ram[2][36] ), .A2(n5362), .A3(n5363), .A4(data[36]), 
        .Y(n609) );
  AO22X1_HVT U1950 ( .A1(\ram[2][35] ), .A2(n5362), .A3(n5363), .A4(data[35]), 
        .Y(n608) );
  AO22X1_HVT U1951 ( .A1(\ram[2][34] ), .A2(n5362), .A3(n5363), .A4(data[34]), 
        .Y(n607) );
  AO22X1_HVT U1952 ( .A1(\ram[2][33] ), .A2(n5362), .A3(n5363), .A4(data[33]), 
        .Y(n606) );
  AO22X1_HVT U1953 ( .A1(\ram[2][32] ), .A2(n5362), .A3(n5363), .A4(data[32]), 
        .Y(n605) );
  AO22X1_HVT U1954 ( .A1(\ram[2][31] ), .A2(n5362), .A3(n5363), .A4(data[31]), 
        .Y(n604) );
  AO22X1_HVT U1955 ( .A1(\ram[2][30] ), .A2(n5362), .A3(n5363), .A4(data[30]), 
        .Y(n603) );
  AO22X1_HVT U1956 ( .A1(\ram[2][29] ), .A2(n5362), .A3(n5363), .A4(data[29]), 
        .Y(n602) );
  AO22X1_HVT U1957 ( .A1(\ram[2][28] ), .A2(n5362), .A3(n5363), .A4(data[28]), 
        .Y(n601) );
  AO22X1_HVT U1958 ( .A1(\ram[2][27] ), .A2(n5362), .A3(n5363), .A4(data[27]), 
        .Y(n600) );
  AO22X1_HVT U1959 ( .A1(\ram[2][26] ), .A2(n5362), .A3(n5363), .A4(data[26]), 
        .Y(n599) );
  AO22X1_HVT U1960 ( .A1(\ram[2][25] ), .A2(n5362), .A3(n5363), .A4(data[25]), 
        .Y(n598) );
  AO22X1_HVT U1961 ( .A1(\ram[2][24] ), .A2(n5362), .A3(n5363), .A4(data[24]), 
        .Y(n597) );
  AO22X1_HVT U1962 ( .A1(\ram[2][23] ), .A2(n5362), .A3(n5363), .A4(data[23]), 
        .Y(n596) );
  AO22X1_HVT U1963 ( .A1(\ram[2][22] ), .A2(n5362), .A3(n5363), .A4(data[22]), 
        .Y(n595) );
  AO22X1_HVT U1964 ( .A1(\ram[2][21] ), .A2(n5362), .A3(n5363), .A4(data[21]), 
        .Y(n594) );
  AO22X1_HVT U1965 ( .A1(\ram[2][20] ), .A2(n5362), .A3(n5363), .A4(data[20]), 
        .Y(n593) );
  AO22X1_HVT U1966 ( .A1(\ram[2][19] ), .A2(n5362), .A3(n5363), .A4(data[19]), 
        .Y(n592) );
  AO22X1_HVT U1967 ( .A1(\ram[2][18] ), .A2(n5362), .A3(n5363), .A4(data[18]), 
        .Y(n591) );
  AO22X1_HVT U1968 ( .A1(\ram[2][17] ), .A2(n5362), .A3(n5363), .A4(data[17]), 
        .Y(n590) );
  AO22X1_HVT U1969 ( .A1(\ram[2][16] ), .A2(n5362), .A3(n5363), .A4(data[16]), 
        .Y(n589) );
  AO22X1_HVT U1970 ( .A1(\ram[2][15] ), .A2(n5362), .A3(n5363), .A4(data[15]), 
        .Y(n588) );
  AO22X1_HVT U1971 ( .A1(\ram[2][14] ), .A2(n5362), .A3(n5363), .A4(data[14]), 
        .Y(n587) );
  AO22X1_HVT U1972 ( .A1(\ram[2][13] ), .A2(n5362), .A3(n5363), .A4(data[13]), 
        .Y(n586) );
  AO22X1_HVT U1973 ( .A1(\ram[2][12] ), .A2(n5362), .A3(n5363), .A4(data[12]), 
        .Y(n585) );
  AO22X1_HVT U1974 ( .A1(\ram[2][11] ), .A2(n5362), .A3(n5363), .A4(data[11]), 
        .Y(n584) );
  AO22X1_HVT U1975 ( .A1(\ram[2][10] ), .A2(n5362), .A3(n5363), .A4(data[10]), 
        .Y(n583) );
  AO22X1_HVT U1976 ( .A1(\ram[2][9] ), .A2(n5362), .A3(n5363), .A4(data[9]), 
        .Y(n582) );
  AO22X1_HVT U1977 ( .A1(\ram[2][8] ), .A2(n5362), .A3(n5363), .A4(data[8]), 
        .Y(n581) );
  AO22X1_HVT U1978 ( .A1(\ram[2][7] ), .A2(n5362), .A3(n5363), .A4(data[7]), 
        .Y(n580) );
  AO22X1_HVT U1979 ( .A1(\ram[2][6] ), .A2(n5362), .A3(n5363), .A4(data[6]), 
        .Y(n579) );
  AO22X1_HVT U1980 ( .A1(\ram[2][5] ), .A2(n5362), .A3(n5363), .A4(data[5]), 
        .Y(n578) );
  AO22X1_HVT U1981 ( .A1(\ram[2][4] ), .A2(n5362), .A3(n5363), .A4(data[4]), 
        .Y(n577) );
  AO22X1_HVT U1982 ( .A1(\ram[2][3] ), .A2(n5362), .A3(n5363), .A4(data[3]), 
        .Y(n576) );
  AO22X1_HVT U1983 ( .A1(\ram[2][2] ), .A2(n5362), .A3(n5363), .A4(data[2]), 
        .Y(n575) );
  AO22X1_HVT U1984 ( .A1(\ram[2][1] ), .A2(n5362), .A3(n5363), .A4(data[1]), 
        .Y(n574) );
  AO22X1_HVT U1985 ( .A1(\ram[2][0] ), .A2(n5362), .A3(n5363), .A4(data[0]), 
        .Y(n573) );
  INVX0_HVT U1986 ( .A(n5364), .Y(n5363) );
  AND2X1_HVT U1987 ( .A1(n5364), .A2(n5365), .Y(n5362) );
  NAND3X0_HVT U1988 ( .A1(n5366), .A2(n4183), .A3(n5367), .Y(n5364) );
  AO22X1_HVT U1989 ( .A1(\ram[1][255] ), .A2(n5368), .A3(n5369), .A4(data[255]), .Y(n572) );
  AO22X1_HVT U1990 ( .A1(\ram[1][254] ), .A2(n5368), .A3(n5369), .A4(data[254]), .Y(n571) );
  AO22X1_HVT U1991 ( .A1(\ram[1][253] ), .A2(n5368), .A3(n5369), .A4(data[253]), .Y(n570) );
  AO22X1_HVT U1992 ( .A1(\ram[1][252] ), .A2(n5368), .A3(n5369), .A4(data[252]), .Y(n569) );
  AO22X1_HVT U1993 ( .A1(\ram[1][251] ), .A2(n5368), .A3(n5369), .A4(data[251]), .Y(n568) );
  AO22X1_HVT U1994 ( .A1(\ram[1][250] ), .A2(n5368), .A3(n5369), .A4(data[250]), .Y(n567) );
  AO22X1_HVT U1995 ( .A1(\ram[1][249] ), .A2(n5368), .A3(n5369), .A4(data[249]), .Y(n566) );
  AO22X1_HVT U1996 ( .A1(\ram[1][248] ), .A2(n5368), .A3(n5369), .A4(data[248]), .Y(n565) );
  AO22X1_HVT U1997 ( .A1(\ram[1][247] ), .A2(n5368), .A3(n5369), .A4(data[247]), .Y(n564) );
  AO22X1_HVT U1998 ( .A1(\ram[1][246] ), .A2(n5368), .A3(n5369), .A4(data[246]), .Y(n563) );
  AO22X1_HVT U1999 ( .A1(\ram[1][245] ), .A2(n5368), .A3(n5369), .A4(data[245]), .Y(n562) );
  AO22X1_HVT U2000 ( .A1(\ram[1][244] ), .A2(n5368), .A3(n5369), .A4(data[244]), .Y(n561) );
  AO22X1_HVT U2001 ( .A1(\ram[1][243] ), .A2(n5368), .A3(n5369), .A4(data[243]), .Y(n560) );
  AO22X1_HVT U2002 ( .A1(\ram[1][242] ), .A2(n5368), .A3(n5369), .A4(data[242]), .Y(n559) );
  AO22X1_HVT U2003 ( .A1(\ram[1][241] ), .A2(n5368), .A3(n5369), .A4(data[241]), .Y(n558) );
  AO22X1_HVT U2004 ( .A1(\ram[1][240] ), .A2(n5368), .A3(n5369), .A4(data[240]), .Y(n557) );
  AO22X1_HVT U2005 ( .A1(\ram[1][239] ), .A2(n5368), .A3(n5369), .A4(data[239]), .Y(n556) );
  AO22X1_HVT U2006 ( .A1(\ram[1][238] ), .A2(n5368), .A3(n5369), .A4(data[238]), .Y(n555) );
  AO22X1_HVT U2007 ( .A1(\ram[1][237] ), .A2(n5368), .A3(n5369), .A4(data[237]), .Y(n554) );
  AO22X1_HVT U2008 ( .A1(\ram[1][236] ), .A2(n5368), .A3(n5369), .A4(data[236]), .Y(n553) );
  AO22X1_HVT U2009 ( .A1(\ram[1][235] ), .A2(n5368), .A3(n5369), .A4(data[235]), .Y(n552) );
  AO22X1_HVT U2010 ( .A1(\ram[1][234] ), .A2(n5368), .A3(n5369), .A4(data[234]), .Y(n551) );
  AO22X1_HVT U2011 ( .A1(\ram[1][233] ), .A2(n5368), .A3(n5369), .A4(data[233]), .Y(n550) );
  AO22X1_HVT U2012 ( .A1(\ram[1][232] ), .A2(n5368), .A3(n5369), .A4(data[232]), .Y(n549) );
  AO22X1_HVT U2013 ( .A1(\ram[1][231] ), .A2(n5368), .A3(n5369), .A4(data[231]), .Y(n548) );
  AO22X1_HVT U2014 ( .A1(\ram[1][230] ), .A2(n5368), .A3(n5369), .A4(data[230]), .Y(n547) );
  AO22X1_HVT U2015 ( .A1(\ram[1][229] ), .A2(n5368), .A3(n5369), .A4(data[229]), .Y(n546) );
  AO22X1_HVT U2016 ( .A1(\ram[1][228] ), .A2(n5368), .A3(n5369), .A4(data[228]), .Y(n545) );
  AO22X1_HVT U2017 ( .A1(\ram[1][227] ), .A2(n5368), .A3(n5369), .A4(data[227]), .Y(n544) );
  AO22X1_HVT U2018 ( .A1(\ram[1][226] ), .A2(n5368), .A3(n5369), .A4(data[226]), .Y(n543) );
  AO22X1_HVT U2019 ( .A1(\ram[1][225] ), .A2(n5368), .A3(n5369), .A4(data[225]), .Y(n542) );
  AO22X1_HVT U2020 ( .A1(\ram[1][224] ), .A2(n5368), .A3(n5369), .A4(data[224]), .Y(n541) );
  AO22X1_HVT U2021 ( .A1(\ram[1][223] ), .A2(n5368), .A3(n5369), .A4(data[223]), .Y(n540) );
  AO22X1_HVT U2022 ( .A1(\ram[1][222] ), .A2(n5368), .A3(n5369), .A4(data[222]), .Y(n539) );
  AO22X1_HVT U2023 ( .A1(\ram[1][221] ), .A2(n5368), .A3(n5369), .A4(data[221]), .Y(n538) );
  AO22X1_HVT U2024 ( .A1(\ram[1][220] ), .A2(n5368), .A3(n5369), .A4(data[220]), .Y(n537) );
  AO22X1_HVT U2025 ( .A1(\ram[1][219] ), .A2(n5368), .A3(n5369), .A4(data[219]), .Y(n536) );
  AO22X1_HVT U2026 ( .A1(\ram[1][218] ), .A2(n5368), .A3(n5369), .A4(data[218]), .Y(n535) );
  AO22X1_HVT U2027 ( .A1(\ram[1][217] ), .A2(n5368), .A3(n5369), .A4(data[217]), .Y(n534) );
  AO22X1_HVT U2028 ( .A1(\ram[1][216] ), .A2(n5368), .A3(n5369), .A4(data[216]), .Y(n533) );
  AO22X1_HVT U2029 ( .A1(\ram[1][215] ), .A2(n5368), .A3(n5369), .A4(data[215]), .Y(n532) );
  AO22X1_HVT U2030 ( .A1(\ram[1][214] ), .A2(n5368), .A3(n5369), .A4(data[214]), .Y(n531) );
  AO22X1_HVT U2031 ( .A1(\ram[1][213] ), .A2(n5368), .A3(n5369), .A4(data[213]), .Y(n530) );
  AO22X1_HVT U2032 ( .A1(\ram[1][212] ), .A2(n5368), .A3(n5369), .A4(data[212]), .Y(n529) );
  AO22X1_HVT U2033 ( .A1(\ram[1][211] ), .A2(n5368), .A3(n5369), .A4(data[211]), .Y(n528) );
  AO22X1_HVT U2034 ( .A1(\ram[1][210] ), .A2(n5368), .A3(n5369), .A4(data[210]), .Y(n527) );
  AO22X1_HVT U2035 ( .A1(\ram[1][209] ), .A2(n5368), .A3(n5369), .A4(data[209]), .Y(n526) );
  AO22X1_HVT U2036 ( .A1(\ram[1][208] ), .A2(n5368), .A3(n5369), .A4(data[208]), .Y(n525) );
  AO22X1_HVT U2037 ( .A1(\ram[1][207] ), .A2(n5368), .A3(n5369), .A4(data[207]), .Y(n524) );
  AO22X1_HVT U2038 ( .A1(\ram[1][206] ), .A2(n5368), .A3(n5369), .A4(data[206]), .Y(n523) );
  AO22X1_HVT U2039 ( .A1(\ram[1][205] ), .A2(n5368), .A3(n5369), .A4(data[205]), .Y(n522) );
  AO22X1_HVT U2040 ( .A1(\ram[1][204] ), .A2(n5368), .A3(n5369), .A4(data[204]), .Y(n521) );
  AO22X1_HVT U2041 ( .A1(\ram[1][203] ), .A2(n5368), .A3(n5369), .A4(data[203]), .Y(n520) );
  AO22X1_HVT U2042 ( .A1(\ram[1][202] ), .A2(n5368), .A3(n5369), .A4(data[202]), .Y(n519) );
  AO22X1_HVT U2043 ( .A1(\ram[1][201] ), .A2(n5368), .A3(n5369), .A4(data[201]), .Y(n518) );
  AO22X1_HVT U2044 ( .A1(\ram[1][200] ), .A2(n5368), .A3(n5369), .A4(data[200]), .Y(n517) );
  AO22X1_HVT U2045 ( .A1(\ram[1][199] ), .A2(n5368), .A3(n5369), .A4(data[199]), .Y(n516) );
  AO22X1_HVT U2046 ( .A1(\ram[1][198] ), .A2(n5368), .A3(n5369), .A4(data[198]), .Y(n515) );
  AO22X1_HVT U2047 ( .A1(\ram[1][197] ), .A2(n5368), .A3(n5369), .A4(data[197]), .Y(n514) );
  AO22X1_HVT U2048 ( .A1(\ram[1][196] ), .A2(n5368), .A3(n5369), .A4(data[196]), .Y(n513) );
  AO22X1_HVT U2049 ( .A1(\ram[1][195] ), .A2(n5368), .A3(n5369), .A4(data[195]), .Y(n512) );
  AO22X1_HVT U2050 ( .A1(\ram[1][194] ), .A2(n5368), .A3(n5369), .A4(data[194]), .Y(n511) );
  AO22X1_HVT U2051 ( .A1(\ram[1][193] ), .A2(n5368), .A3(n5369), .A4(data[193]), .Y(n510) );
  AO22X1_HVT U2052 ( .A1(\ram[1][192] ), .A2(n5368), .A3(n5369), .A4(data[192]), .Y(n509) );
  AO22X1_HVT U2053 ( .A1(\ram[1][191] ), .A2(n5368), .A3(n5369), .A4(data[191]), .Y(n508) );
  AO22X1_HVT U2054 ( .A1(\ram[1][190] ), .A2(n5368), .A3(n5369), .A4(data[190]), .Y(n507) );
  AO22X1_HVT U2055 ( .A1(\ram[1][189] ), .A2(n5368), .A3(n5369), .A4(data[189]), .Y(n506) );
  AO22X1_HVT U2056 ( .A1(\ram[1][188] ), .A2(n5368), .A3(n5369), .A4(data[188]), .Y(n505) );
  AO22X1_HVT U2057 ( .A1(\ram[1][187] ), .A2(n5368), .A3(n5369), .A4(data[187]), .Y(n504) );
  AO22X1_HVT U2058 ( .A1(\ram[1][186] ), .A2(n5368), .A3(n5369), .A4(data[186]), .Y(n503) );
  AO22X1_HVT U2059 ( .A1(\ram[1][185] ), .A2(n5368), .A3(n5369), .A4(data[185]), .Y(n502) );
  AO22X1_HVT U2060 ( .A1(\ram[1][184] ), .A2(n5368), .A3(n5369), .A4(data[184]), .Y(n501) );
  AO22X1_HVT U2061 ( .A1(\ram[1][183] ), .A2(n5368), .A3(n5369), .A4(data[183]), .Y(n500) );
  AO22X1_HVT U2062 ( .A1(\ram[1][182] ), .A2(n5368), .A3(n5369), .A4(data[182]), .Y(n499) );
  AO22X1_HVT U2063 ( .A1(\ram[1][181] ), .A2(n5368), .A3(n5369), .A4(data[181]), .Y(n498) );
  AO22X1_HVT U2064 ( .A1(\ram[1][180] ), .A2(n5368), .A3(n5369), .A4(data[180]), .Y(n497) );
  AO22X1_HVT U2065 ( .A1(\ram[1][179] ), .A2(n5368), .A3(n5369), .A4(data[179]), .Y(n496) );
  AO22X1_HVT U2066 ( .A1(\ram[1][178] ), .A2(n5368), .A3(n5369), .A4(data[178]), .Y(n495) );
  AO22X1_HVT U2067 ( .A1(\ram[1][177] ), .A2(n5368), .A3(n5369), .A4(data[177]), .Y(n494) );
  AO22X1_HVT U2068 ( .A1(\ram[1][176] ), .A2(n5368), .A3(n5369), .A4(data[176]), .Y(n493) );
  AO22X1_HVT U2069 ( .A1(\ram[1][175] ), .A2(n5368), .A3(n5369), .A4(data[175]), .Y(n492) );
  AO22X1_HVT U2070 ( .A1(\ram[1][174] ), .A2(n5368), .A3(n5369), .A4(data[174]), .Y(n491) );
  AO22X1_HVT U2071 ( .A1(\ram[1][173] ), .A2(n5368), .A3(n5369), .A4(data[173]), .Y(n490) );
  AO22X1_HVT U2072 ( .A1(\ram[1][172] ), .A2(n5368), .A3(n5369), .A4(data[172]), .Y(n489) );
  AO22X1_HVT U2073 ( .A1(\ram[1][171] ), .A2(n5368), .A3(n5369), .A4(data[171]), .Y(n488) );
  AO22X1_HVT U2074 ( .A1(\ram[1][170] ), .A2(n5368), .A3(n5369), .A4(data[170]), .Y(n487) );
  AO22X1_HVT U2075 ( .A1(\ram[1][169] ), .A2(n5368), .A3(n5369), .A4(data[169]), .Y(n486) );
  AO22X1_HVT U2076 ( .A1(\ram[1][168] ), .A2(n5368), .A3(n5369), .A4(data[168]), .Y(n485) );
  AO22X1_HVT U2077 ( .A1(\ram[1][167] ), .A2(n5368), .A3(n5369), .A4(data[167]), .Y(n484) );
  AO22X1_HVT U2078 ( .A1(\ram[1][166] ), .A2(n5368), .A3(n5369), .A4(data[166]), .Y(n483) );
  AO22X1_HVT U2079 ( .A1(\ram[1][165] ), .A2(n5368), .A3(n5369), .A4(data[165]), .Y(n482) );
  AO22X1_HVT U2080 ( .A1(\ram[1][164] ), .A2(n5368), .A3(n5369), .A4(data[164]), .Y(n481) );
  AO22X1_HVT U2081 ( .A1(\ram[1][163] ), .A2(n5368), .A3(n5369), .A4(data[163]), .Y(n480) );
  AO22X1_HVT U2082 ( .A1(\ram[1][162] ), .A2(n5368), .A3(n5369), .A4(data[162]), .Y(n479) );
  AO22X1_HVT U2083 ( .A1(\ram[1][161] ), .A2(n5368), .A3(n5369), .A4(data[161]), .Y(n478) );
  AO22X1_HVT U2084 ( .A1(\ram[1][160] ), .A2(n5368), .A3(n5369), .A4(data[160]), .Y(n477) );
  AO22X1_HVT U2085 ( .A1(\ram[1][159] ), .A2(n5368), .A3(n5369), .A4(data[159]), .Y(n476) );
  AO22X1_HVT U2086 ( .A1(\ram[1][158] ), .A2(n5368), .A3(n5369), .A4(data[158]), .Y(n475) );
  AO22X1_HVT U2087 ( .A1(\ram[1][157] ), .A2(n5368), .A3(n5369), .A4(data[157]), .Y(n474) );
  AO22X1_HVT U2088 ( .A1(\ram[1][156] ), .A2(n5368), .A3(n5369), .A4(data[156]), .Y(n473) );
  AO22X1_HVT U2089 ( .A1(\ram[1][155] ), .A2(n5368), .A3(n5369), .A4(data[155]), .Y(n472) );
  AO22X1_HVT U2090 ( .A1(\ram[1][154] ), .A2(n5368), .A3(n5369), .A4(data[154]), .Y(n471) );
  AO22X1_HVT U2091 ( .A1(\ram[1][153] ), .A2(n5368), .A3(n5369), .A4(data[153]), .Y(n470) );
  AO22X1_HVT U2092 ( .A1(\ram[1][152] ), .A2(n5368), .A3(n5369), .A4(data[152]), .Y(n469) );
  AO22X1_HVT U2093 ( .A1(\ram[1][151] ), .A2(n5368), .A3(n5369), .A4(data[151]), .Y(n468) );
  AO22X1_HVT U2094 ( .A1(\ram[1][150] ), .A2(n5368), .A3(n5369), .A4(data[150]), .Y(n467) );
  AO22X1_HVT U2095 ( .A1(\ram[1][149] ), .A2(n5368), .A3(n5369), .A4(data[149]), .Y(n466) );
  AO22X1_HVT U2096 ( .A1(\ram[1][148] ), .A2(n5368), .A3(n5369), .A4(data[148]), .Y(n465) );
  AO22X1_HVT U2097 ( .A1(\ram[1][147] ), .A2(n5368), .A3(n5369), .A4(data[147]), .Y(n464) );
  AO22X1_HVT U2098 ( .A1(\ram[1][146] ), .A2(n5368), .A3(n5369), .A4(data[146]), .Y(n463) );
  AO22X1_HVT U2099 ( .A1(\ram[1][145] ), .A2(n5368), .A3(n5369), .A4(data[145]), .Y(n462) );
  AO22X1_HVT U2100 ( .A1(\ram[1][144] ), .A2(n5368), .A3(n5369), .A4(data[144]), .Y(n461) );
  AO22X1_HVT U2101 ( .A1(\ram[1][143] ), .A2(n5368), .A3(n5369), .A4(data[143]), .Y(n460) );
  AO22X1_HVT U2102 ( .A1(\ram[1][142] ), .A2(n5368), .A3(n5369), .A4(data[142]), .Y(n459) );
  AO22X1_HVT U2103 ( .A1(\ram[1][141] ), .A2(n5368), .A3(n5369), .A4(data[141]), .Y(n458) );
  AO22X1_HVT U2104 ( .A1(\ram[1][140] ), .A2(n5368), .A3(n5369), .A4(data[140]), .Y(n457) );
  AO22X1_HVT U2105 ( .A1(\ram[1][139] ), .A2(n5368), .A3(n5369), .A4(data[139]), .Y(n456) );
  AO22X1_HVT U2106 ( .A1(\ram[1][138] ), .A2(n5368), .A3(n5369), .A4(data[138]), .Y(n455) );
  AO22X1_HVT U2107 ( .A1(\ram[1][137] ), .A2(n5368), .A3(n5369), .A4(data[137]), .Y(n454) );
  AO22X1_HVT U2108 ( .A1(\ram[1][136] ), .A2(n5368), .A3(n5369), .A4(data[136]), .Y(n453) );
  AO22X1_HVT U2109 ( .A1(\ram[1][135] ), .A2(n5368), .A3(n5369), .A4(data[135]), .Y(n452) );
  AO22X1_HVT U2110 ( .A1(\ram[1][134] ), .A2(n5368), .A3(n5369), .A4(data[134]), .Y(n451) );
  AO22X1_HVT U2111 ( .A1(\ram[1][133] ), .A2(n5368), .A3(n5369), .A4(data[133]), .Y(n450) );
  AO22X1_HVT U2112 ( .A1(\ram[1][132] ), .A2(n5368), .A3(n5369), .A4(data[132]), .Y(n449) );
  AO22X1_HVT U2113 ( .A1(\ram[1][131] ), .A2(n5368), .A3(n5369), .A4(data[131]), .Y(n448) );
  AO22X1_HVT U2114 ( .A1(\ram[1][130] ), .A2(n5368), .A3(n5369), .A4(data[130]), .Y(n447) );
  AO22X1_HVT U2115 ( .A1(\ram[1][129] ), .A2(n5368), .A3(n5369), .A4(data[129]), .Y(n446) );
  AO22X1_HVT U2116 ( .A1(\ram[1][128] ), .A2(n5368), .A3(n5369), .A4(data[128]), .Y(n445) );
  AO22X1_HVT U2117 ( .A1(\ram[1][127] ), .A2(n5368), .A3(n5369), .A4(data[127]), .Y(n444) );
  AO22X1_HVT U2118 ( .A1(\ram[1][126] ), .A2(n5368), .A3(n5369), .A4(data[126]), .Y(n443) );
  AO22X1_HVT U2119 ( .A1(\ram[1][125] ), .A2(n5368), .A3(n5369), .A4(data[125]), .Y(n442) );
  AO22X1_HVT U2120 ( .A1(\ram[1][124] ), .A2(n5368), .A3(n5369), .A4(data[124]), .Y(n441) );
  AO22X1_HVT U2121 ( .A1(\ram[1][123] ), .A2(n5368), .A3(n5369), .A4(data[123]), .Y(n440) );
  AO22X1_HVT U2122 ( .A1(\ram[1][122] ), .A2(n5368), .A3(n5369), .A4(data[122]), .Y(n439) );
  AO22X1_HVT U2123 ( .A1(\ram[1][121] ), .A2(n5368), .A3(n5369), .A4(data[121]), .Y(n438) );
  AO22X1_HVT U2124 ( .A1(\ram[1][120] ), .A2(n5368), .A3(n5369), .A4(data[120]), .Y(n437) );
  AO22X1_HVT U2125 ( .A1(\ram[1][119] ), .A2(n5368), .A3(n5369), .A4(data[119]), .Y(n436) );
  AO22X1_HVT U2126 ( .A1(\ram[1][118] ), .A2(n5368), .A3(n5369), .A4(data[118]), .Y(n435) );
  AO22X1_HVT U2127 ( .A1(\ram[1][117] ), .A2(n5368), .A3(n5369), .A4(data[117]), .Y(n434) );
  AO22X1_HVT U2128 ( .A1(\ram[1][116] ), .A2(n5368), .A3(n5369), .A4(data[116]), .Y(n433) );
  AO22X1_HVT U2129 ( .A1(\ram[1][115] ), .A2(n5368), .A3(n5369), .A4(data[115]), .Y(n432) );
  AO22X1_HVT U2130 ( .A1(\ram[1][114] ), .A2(n5368), .A3(n5369), .A4(data[114]), .Y(n431) );
  AO22X1_HVT U2131 ( .A1(\ram[1][113] ), .A2(n5368), .A3(n5369), .A4(data[113]), .Y(n430) );
  AO22X1_HVT U2132 ( .A1(\ram[1][112] ), .A2(n5368), .A3(n5369), .A4(data[112]), .Y(n429) );
  AO22X1_HVT U2133 ( .A1(\ram[1][111] ), .A2(n5368), .A3(n5369), .A4(data[111]), .Y(n428) );
  AO22X1_HVT U2134 ( .A1(\ram[1][110] ), .A2(n5368), .A3(n5369), .A4(data[110]), .Y(n427) );
  AO22X1_HVT U2135 ( .A1(\ram[1][109] ), .A2(n5368), .A3(n5369), .A4(data[109]), .Y(n426) );
  AO22X1_HVT U2136 ( .A1(\ram[1][108] ), .A2(n5368), .A3(n5369), .A4(data[108]), .Y(n425) );
  AO22X1_HVT U2137 ( .A1(\ram[1][107] ), .A2(n5368), .A3(n5369), .A4(data[107]), .Y(n424) );
  AO22X1_HVT U2138 ( .A1(\ram[1][106] ), .A2(n5368), .A3(n5369), .A4(data[106]), .Y(n423) );
  AO22X1_HVT U2139 ( .A1(\ram[1][105] ), .A2(n5368), .A3(n5369), .A4(data[105]), .Y(n422) );
  AO22X1_HVT U2140 ( .A1(\ram[1][104] ), .A2(n5368), .A3(n5369), .A4(data[104]), .Y(n421) );
  AO22X1_HVT U2141 ( .A1(\ram[1][103] ), .A2(n5368), .A3(n5369), .A4(data[103]), .Y(n420) );
  AO22X1_HVT U2142 ( .A1(\ram[1][102] ), .A2(n5368), .A3(n5369), .A4(data[102]), .Y(n419) );
  AO22X1_HVT U2143 ( .A1(\ram[1][101] ), .A2(n5368), .A3(n5369), .A4(data[101]), .Y(n418) );
  AO22X1_HVT U2144 ( .A1(\ram[1][100] ), .A2(n5368), .A3(n5369), .A4(data[100]), .Y(n417) );
  AO22X1_HVT U2145 ( .A1(\ram[1][99] ), .A2(n5368), .A3(n5369), .A4(data[99]), 
        .Y(n416) );
  AO22X1_HVT U2146 ( .A1(\ram[15][255] ), .A2(n5370), .A3(n5371), .A4(
        data[255]), .Y(n4156) );
  AO22X1_HVT U2147 ( .A1(\ram[15][254] ), .A2(n5370), .A3(n5371), .A4(
        data[254]), .Y(n4155) );
  AO22X1_HVT U2148 ( .A1(\ram[15][253] ), .A2(n5370), .A3(n5371), .A4(
        data[253]), .Y(n4154) );
  AO22X1_HVT U2149 ( .A1(\ram[15][252] ), .A2(n5370), .A3(n5371), .A4(
        data[252]), .Y(n4153) );
  AO22X1_HVT U2150 ( .A1(\ram[15][251] ), .A2(n5370), .A3(n5371), .A4(
        data[251]), .Y(n4152) );
  AO22X1_HVT U2151 ( .A1(\ram[15][250] ), .A2(n5370), .A3(n5371), .A4(
        data[250]), .Y(n4151) );
  AO22X1_HVT U2152 ( .A1(\ram[15][249] ), .A2(n5370), .A3(n5371), .A4(
        data[249]), .Y(n4150) );
  AO22X1_HVT U2153 ( .A1(\ram[1][98] ), .A2(n5368), .A3(n5369), .A4(data[98]), 
        .Y(n415) );
  AO22X1_HVT U2154 ( .A1(\ram[15][248] ), .A2(n5370), .A3(n5371), .A4(
        data[248]), .Y(n4149) );
  AO22X1_HVT U2155 ( .A1(\ram[15][247] ), .A2(n5370), .A3(n5371), .A4(
        data[247]), .Y(n4148) );
  AO22X1_HVT U2156 ( .A1(\ram[15][246] ), .A2(n5370), .A3(n5371), .A4(
        data[246]), .Y(n4147) );
  AO22X1_HVT U2157 ( .A1(\ram[15][245] ), .A2(n5370), .A3(n5371), .A4(
        data[245]), .Y(n4146) );
  AO22X1_HVT U2158 ( .A1(\ram[15][244] ), .A2(n5370), .A3(n5371), .A4(
        data[244]), .Y(n4145) );
  AO22X1_HVT U2159 ( .A1(\ram[15][243] ), .A2(n5370), .A3(n5371), .A4(
        data[243]), .Y(n4144) );
  AO22X1_HVT U2160 ( .A1(\ram[15][242] ), .A2(n5370), .A3(n5371), .A4(
        data[242]), .Y(n4143) );
  AO22X1_HVT U2161 ( .A1(\ram[15][241] ), .A2(n5370), .A3(n5371), .A4(
        data[241]), .Y(n4142) );
  AO22X1_HVT U2162 ( .A1(\ram[15][240] ), .A2(n5370), .A3(n5371), .A4(
        data[240]), .Y(n4141) );
  AO22X1_HVT U2163 ( .A1(\ram[15][239] ), .A2(n5370), .A3(n5371), .A4(
        data[239]), .Y(n4140) );
  AO22X1_HVT U2164 ( .A1(\ram[1][97] ), .A2(n5368), .A3(n5369), .A4(data[97]), 
        .Y(n414) );
  AO22X1_HVT U2165 ( .A1(\ram[15][238] ), .A2(n5370), .A3(n5371), .A4(
        data[238]), .Y(n4139) );
  AO22X1_HVT U2166 ( .A1(\ram[15][237] ), .A2(n5370), .A3(n5371), .A4(
        data[237]), .Y(n4138) );
  AO22X1_HVT U2167 ( .A1(\ram[15][236] ), .A2(n5370), .A3(n5371), .A4(
        data[236]), .Y(n4137) );
  AO22X1_HVT U2168 ( .A1(\ram[15][235] ), .A2(n5370), .A3(n5371), .A4(
        data[235]), .Y(n4136) );
  AO22X1_HVT U2169 ( .A1(\ram[15][234] ), .A2(n5370), .A3(n5371), .A4(
        data[234]), .Y(n4135) );
  AO22X1_HVT U2170 ( .A1(\ram[15][233] ), .A2(n5370), .A3(n5371), .A4(
        data[233]), .Y(n4134) );
  AO22X1_HVT U2171 ( .A1(\ram[15][232] ), .A2(n5370), .A3(n5371), .A4(
        data[232]), .Y(n4133) );
  AO22X1_HVT U2172 ( .A1(\ram[15][231] ), .A2(n5370), .A3(n5371), .A4(
        data[231]), .Y(n4132) );
  AO22X1_HVT U2173 ( .A1(\ram[15][230] ), .A2(n5370), .A3(n5371), .A4(
        data[230]), .Y(n4131) );
  AO22X1_HVT U2174 ( .A1(\ram[15][229] ), .A2(n5370), .A3(n5371), .A4(
        data[229]), .Y(n4130) );
  AO22X1_HVT U2175 ( .A1(\ram[1][96] ), .A2(n5368), .A3(n5369), .A4(data[96]), 
        .Y(n413) );
  AO22X1_HVT U2176 ( .A1(\ram[15][228] ), .A2(n5370), .A3(n5371), .A4(
        data[228]), .Y(n4129) );
  AO22X1_HVT U2177 ( .A1(\ram[15][227] ), .A2(n5370), .A3(n5371), .A4(
        data[227]), .Y(n4128) );
  AO22X1_HVT U2178 ( .A1(\ram[15][226] ), .A2(n5370), .A3(n5371), .A4(
        data[226]), .Y(n4127) );
  AO22X1_HVT U2179 ( .A1(\ram[15][225] ), .A2(n5370), .A3(n5371), .A4(
        data[225]), .Y(n4126) );
  AO22X1_HVT U2180 ( .A1(\ram[15][224] ), .A2(n5370), .A3(n5371), .A4(
        data[224]), .Y(n4125) );
  AO22X1_HVT U2181 ( .A1(\ram[15][223] ), .A2(n5370), .A3(n5371), .A4(
        data[223]), .Y(n4124) );
  AO22X1_HVT U2182 ( .A1(\ram[15][222] ), .A2(n5370), .A3(n5371), .A4(
        data[222]), .Y(n4123) );
  AO22X1_HVT U2183 ( .A1(\ram[15][221] ), .A2(n5370), .A3(n5371), .A4(
        data[221]), .Y(n4122) );
  AO22X1_HVT U2184 ( .A1(\ram[15][220] ), .A2(n5370), .A3(n5371), .A4(
        data[220]), .Y(n4121) );
  AO22X1_HVT U2185 ( .A1(\ram[15][219] ), .A2(n5370), .A3(n5371), .A4(
        data[219]), .Y(n4120) );
  AO22X1_HVT U2186 ( .A1(\ram[1][95] ), .A2(n5368), .A3(n5369), .A4(data[95]), 
        .Y(n412) );
  AO22X1_HVT U2187 ( .A1(\ram[15][218] ), .A2(n5370), .A3(n5371), .A4(
        data[218]), .Y(n4119) );
  AO22X1_HVT U2188 ( .A1(\ram[15][217] ), .A2(n5370), .A3(n5371), .A4(
        data[217]), .Y(n4118) );
  AO22X1_HVT U2189 ( .A1(\ram[15][216] ), .A2(n5370), .A3(n5371), .A4(
        data[216]), .Y(n4117) );
  AO22X1_HVT U2190 ( .A1(\ram[15][215] ), .A2(n5370), .A3(n5371), .A4(
        data[215]), .Y(n4116) );
  AO22X1_HVT U2191 ( .A1(\ram[15][214] ), .A2(n5370), .A3(n5371), .A4(
        data[214]), .Y(n4115) );
  AO22X1_HVT U2192 ( .A1(\ram[15][213] ), .A2(n5370), .A3(n5371), .A4(
        data[213]), .Y(n4114) );
  AO22X1_HVT U2193 ( .A1(\ram[15][212] ), .A2(n5370), .A3(n5371), .A4(
        data[212]), .Y(n4113) );
  AO22X1_HVT U2194 ( .A1(\ram[15][211] ), .A2(n5370), .A3(n5371), .A4(
        data[211]), .Y(n4112) );
  AO22X1_HVT U2195 ( .A1(\ram[15][210] ), .A2(n5370), .A3(n5371), .A4(
        data[210]), .Y(n4111) );
  AO22X1_HVT U2196 ( .A1(\ram[15][209] ), .A2(n5370), .A3(n5371), .A4(
        data[209]), .Y(n4110) );
  AO22X1_HVT U2197 ( .A1(\ram[1][94] ), .A2(n5368), .A3(n5369), .A4(data[94]), 
        .Y(n411) );
  AO22X1_HVT U2198 ( .A1(\ram[15][208] ), .A2(n5370), .A3(n5371), .A4(
        data[208]), .Y(n4109) );
  AO22X1_HVT U2199 ( .A1(\ram[15][207] ), .A2(n5370), .A3(n5371), .A4(
        data[207]), .Y(n4108) );
  AO22X1_HVT U2200 ( .A1(\ram[15][206] ), .A2(n5370), .A3(n5371), .A4(
        data[206]), .Y(n4107) );
  AO22X1_HVT U2201 ( .A1(\ram[15][205] ), .A2(n5370), .A3(n5371), .A4(
        data[205]), .Y(n4106) );
  AO22X1_HVT U2202 ( .A1(\ram[15][204] ), .A2(n5370), .A3(n5371), .A4(
        data[204]), .Y(n4105) );
  AO22X1_HVT U2203 ( .A1(\ram[15][203] ), .A2(n5370), .A3(n5371), .A4(
        data[203]), .Y(n4104) );
  AO22X1_HVT U2204 ( .A1(\ram[15][202] ), .A2(n5370), .A3(n5371), .A4(
        data[202]), .Y(n4103) );
  AO22X1_HVT U2205 ( .A1(\ram[15][201] ), .A2(n5370), .A3(n5371), .A4(
        data[201]), .Y(n4102) );
  AO22X1_HVT U2206 ( .A1(\ram[15][200] ), .A2(n5370), .A3(n5371), .A4(
        data[200]), .Y(n4101) );
  AO22X1_HVT U2207 ( .A1(\ram[15][199] ), .A2(n5370), .A3(n5371), .A4(
        data[199]), .Y(n4100) );
  AO22X1_HVT U2208 ( .A1(\ram[1][93] ), .A2(n5368), .A3(n5369), .A4(data[93]), 
        .Y(n410) );
  AO22X1_HVT U2209 ( .A1(\ram[15][198] ), .A2(n5370), .A3(n5371), .A4(
        data[198]), .Y(n4099) );
  AO22X1_HVT U2210 ( .A1(\ram[15][197] ), .A2(n5370), .A3(n5371), .A4(
        data[197]), .Y(n4098) );
  AO22X1_HVT U2211 ( .A1(\ram[15][196] ), .A2(n5370), .A3(n5371), .A4(
        data[196]), .Y(n4097) );
  AO22X1_HVT U2212 ( .A1(\ram[15][195] ), .A2(n5370), .A3(n5371), .A4(
        data[195]), .Y(n4096) );
  AO22X1_HVT U2213 ( .A1(\ram[15][194] ), .A2(n5370), .A3(n5371), .A4(
        data[194]), .Y(n4095) );
  AO22X1_HVT U2214 ( .A1(\ram[15][193] ), .A2(n5370), .A3(n5371), .A4(
        data[193]), .Y(n4094) );
  AO22X1_HVT U2215 ( .A1(\ram[15][192] ), .A2(n5370), .A3(n5371), .A4(
        data[192]), .Y(n4093) );
  AO22X1_HVT U2216 ( .A1(\ram[15][191] ), .A2(n5370), .A3(n5371), .A4(
        data[191]), .Y(n4092) );
  AO22X1_HVT U2217 ( .A1(\ram[15][190] ), .A2(n5370), .A3(n5371), .A4(
        data[190]), .Y(n4091) );
  AO22X1_HVT U2218 ( .A1(\ram[15][189] ), .A2(n5370), .A3(n5371), .A4(
        data[189]), .Y(n4090) );
  AO22X1_HVT U2219 ( .A1(\ram[1][92] ), .A2(n5368), .A3(n5369), .A4(data[92]), 
        .Y(n409) );
  AO22X1_HVT U2220 ( .A1(\ram[15][188] ), .A2(n5370), .A3(n5371), .A4(
        data[188]), .Y(n4089) );
  AO22X1_HVT U2221 ( .A1(\ram[15][187] ), .A2(n5370), .A3(n5371), .A4(
        data[187]), .Y(n4088) );
  AO22X1_HVT U2222 ( .A1(\ram[15][186] ), .A2(n5370), .A3(n5371), .A4(
        data[186]), .Y(n4087) );
  AO22X1_HVT U2223 ( .A1(\ram[15][185] ), .A2(n5370), .A3(n5371), .A4(
        data[185]), .Y(n4086) );
  AO22X1_HVT U2224 ( .A1(\ram[15][184] ), .A2(n5370), .A3(n5371), .A4(
        data[184]), .Y(n4085) );
  AO22X1_HVT U2225 ( .A1(\ram[15][183] ), .A2(n5370), .A3(n5371), .A4(
        data[183]), .Y(n4084) );
  AO22X1_HVT U2226 ( .A1(\ram[15][182] ), .A2(n5370), .A3(n5371), .A4(
        data[182]), .Y(n4083) );
  AO22X1_HVT U2227 ( .A1(\ram[15][181] ), .A2(n5370), .A3(n5371), .A4(
        data[181]), .Y(n4082) );
  AO22X1_HVT U2228 ( .A1(\ram[15][180] ), .A2(n5370), .A3(n5371), .A4(
        data[180]), .Y(n4081) );
  AO22X1_HVT U2229 ( .A1(\ram[15][179] ), .A2(n5370), .A3(n5371), .A4(
        data[179]), .Y(n4080) );
  AO22X1_HVT U2230 ( .A1(\ram[1][91] ), .A2(n5368), .A3(n5369), .A4(data[91]), 
        .Y(n408) );
  AO22X1_HVT U2231 ( .A1(\ram[15][178] ), .A2(n5370), .A3(n5371), .A4(
        data[178]), .Y(n4079) );
  AO22X1_HVT U2232 ( .A1(\ram[15][177] ), .A2(n5370), .A3(n5371), .A4(
        data[177]), .Y(n4078) );
  AO22X1_HVT U2233 ( .A1(\ram[15][176] ), .A2(n5370), .A3(n5371), .A4(
        data[176]), .Y(n4077) );
  AO22X1_HVT U2234 ( .A1(\ram[15][175] ), .A2(n5370), .A3(n5371), .A4(
        data[175]), .Y(n4076) );
  AO22X1_HVT U2235 ( .A1(\ram[15][174] ), .A2(n5370), .A3(n5371), .A4(
        data[174]), .Y(n4075) );
  AO22X1_HVT U2236 ( .A1(\ram[15][173] ), .A2(n5370), .A3(n5371), .A4(
        data[173]), .Y(n4074) );
  AO22X1_HVT U2237 ( .A1(\ram[15][172] ), .A2(n5370), .A3(n5371), .A4(
        data[172]), .Y(n4073) );
  AO22X1_HVT U2238 ( .A1(\ram[15][171] ), .A2(n5370), .A3(n5371), .A4(
        data[171]), .Y(n4072) );
  AO22X1_HVT U2239 ( .A1(\ram[15][170] ), .A2(n5370), .A3(n5371), .A4(
        data[170]), .Y(n4071) );
  AO22X1_HVT U2240 ( .A1(\ram[15][169] ), .A2(n5370), .A3(n5371), .A4(
        data[169]), .Y(n4070) );
  AO22X1_HVT U2241 ( .A1(\ram[1][90] ), .A2(n5368), .A3(n5369), .A4(data[90]), 
        .Y(n407) );
  AO22X1_HVT U2242 ( .A1(\ram[15][168] ), .A2(n5370), .A3(n5371), .A4(
        data[168]), .Y(n4069) );
  AO22X1_HVT U2243 ( .A1(\ram[15][167] ), .A2(n5370), .A3(n5371), .A4(
        data[167]), .Y(n4068) );
  AO22X1_HVT U2244 ( .A1(\ram[15][166] ), .A2(n5370), .A3(n5371), .A4(
        data[166]), .Y(n4067) );
  AO22X1_HVT U2245 ( .A1(\ram[15][165] ), .A2(n5370), .A3(n5371), .A4(
        data[165]), .Y(n4066) );
  AO22X1_HVT U2246 ( .A1(\ram[15][164] ), .A2(n5370), .A3(n5371), .A4(
        data[164]), .Y(n4065) );
  AO22X1_HVT U2247 ( .A1(\ram[15][163] ), .A2(n5370), .A3(n5371), .A4(
        data[163]), .Y(n4064) );
  AO22X1_HVT U2248 ( .A1(\ram[15][162] ), .A2(n5370), .A3(n5371), .A4(
        data[162]), .Y(n4063) );
  AO22X1_HVT U2249 ( .A1(\ram[15][161] ), .A2(n5370), .A3(n5371), .A4(
        data[161]), .Y(n4062) );
  AO22X1_HVT U2250 ( .A1(\ram[15][160] ), .A2(n5370), .A3(n5371), .A4(
        data[160]), .Y(n4061) );
  AO22X1_HVT U2251 ( .A1(\ram[15][159] ), .A2(n5370), .A3(n5371), .A4(
        data[159]), .Y(n4060) );
  AO22X1_HVT U2252 ( .A1(\ram[1][89] ), .A2(n5368), .A3(n5369), .A4(data[89]), 
        .Y(n406) );
  AO22X1_HVT U2253 ( .A1(\ram[15][158] ), .A2(n5370), .A3(n5371), .A4(
        data[158]), .Y(n4059) );
  AO22X1_HVT U2254 ( .A1(\ram[15][157] ), .A2(n5370), .A3(n5371), .A4(
        data[157]), .Y(n4058) );
  AO22X1_HVT U2255 ( .A1(\ram[15][156] ), .A2(n5370), .A3(n5371), .A4(
        data[156]), .Y(n4057) );
  AO22X1_HVT U2256 ( .A1(\ram[15][155] ), .A2(n5370), .A3(n5371), .A4(
        data[155]), .Y(n4056) );
  AO22X1_HVT U2257 ( .A1(\ram[15][154] ), .A2(n5370), .A3(n5371), .A4(
        data[154]), .Y(n4055) );
  AO22X1_HVT U2258 ( .A1(\ram[15][153] ), .A2(n5370), .A3(n5371), .A4(
        data[153]), .Y(n4054) );
  AO22X1_HVT U2259 ( .A1(\ram[15][152] ), .A2(n5370), .A3(n5371), .A4(
        data[152]), .Y(n4053) );
  AO22X1_HVT U2260 ( .A1(\ram[15][151] ), .A2(n5370), .A3(n5371), .A4(
        data[151]), .Y(n4052) );
  AO22X1_HVT U2261 ( .A1(\ram[15][150] ), .A2(n5370), .A3(n5371), .A4(
        data[150]), .Y(n4051) );
  AO22X1_HVT U2262 ( .A1(\ram[15][149] ), .A2(n5370), .A3(n5371), .A4(
        data[149]), .Y(n4050) );
  AO22X1_HVT U2263 ( .A1(\ram[1][88] ), .A2(n5368), .A3(n5369), .A4(data[88]), 
        .Y(n405) );
  AO22X1_HVT U2264 ( .A1(\ram[15][148] ), .A2(n5370), .A3(n5371), .A4(
        data[148]), .Y(n4049) );
  AO22X1_HVT U2265 ( .A1(\ram[15][147] ), .A2(n5370), .A3(n5371), .A4(
        data[147]), .Y(n4048) );
  AO22X1_HVT U2266 ( .A1(\ram[15][146] ), .A2(n5370), .A3(n5371), .A4(
        data[146]), .Y(n4047) );
  AO22X1_HVT U2267 ( .A1(\ram[15][145] ), .A2(n5370), .A3(n5371), .A4(
        data[145]), .Y(n4046) );
  AO22X1_HVT U2268 ( .A1(\ram[15][144] ), .A2(n5370), .A3(n5371), .A4(
        data[144]), .Y(n4045) );
  AO22X1_HVT U2269 ( .A1(\ram[15][143] ), .A2(n5370), .A3(n5371), .A4(
        data[143]), .Y(n4044) );
  AO22X1_HVT U2270 ( .A1(\ram[15][142] ), .A2(n5370), .A3(n5371), .A4(
        data[142]), .Y(n4043) );
  AO22X1_HVT U2271 ( .A1(\ram[15][141] ), .A2(n5370), .A3(n5371), .A4(
        data[141]), .Y(n4042) );
  AO22X1_HVT U2272 ( .A1(\ram[15][140] ), .A2(n5370), .A3(n5371), .A4(
        data[140]), .Y(n4041) );
  AO22X1_HVT U2273 ( .A1(\ram[15][139] ), .A2(n5370), .A3(n5371), .A4(
        data[139]), .Y(n4040) );
  AO22X1_HVT U2274 ( .A1(\ram[1][87] ), .A2(n5368), .A3(n5369), .A4(data[87]), 
        .Y(n404) );
  AO22X1_HVT U2275 ( .A1(\ram[15][138] ), .A2(n5370), .A3(n5371), .A4(
        data[138]), .Y(n4039) );
  AO22X1_HVT U2276 ( .A1(\ram[15][137] ), .A2(n5370), .A3(n5371), .A4(
        data[137]), .Y(n4038) );
  AO22X1_HVT U2277 ( .A1(\ram[15][136] ), .A2(n5370), .A3(n5371), .A4(
        data[136]), .Y(n4037) );
  AO22X1_HVT U2278 ( .A1(\ram[15][135] ), .A2(n5370), .A3(n5371), .A4(
        data[135]), .Y(n4036) );
  AO22X1_HVT U2279 ( .A1(\ram[15][134] ), .A2(n5370), .A3(n5371), .A4(
        data[134]), .Y(n4035) );
  AO22X1_HVT U2280 ( .A1(\ram[15][133] ), .A2(n5370), .A3(n5371), .A4(
        data[133]), .Y(n4034) );
  AO22X1_HVT U2281 ( .A1(\ram[15][132] ), .A2(n5370), .A3(n5371), .A4(
        data[132]), .Y(n4033) );
  AO22X1_HVT U2282 ( .A1(\ram[15][131] ), .A2(n5370), .A3(n5371), .A4(
        data[131]), .Y(n4032) );
  AO22X1_HVT U2283 ( .A1(\ram[15][130] ), .A2(n5370), .A3(n5371), .A4(
        data[130]), .Y(n4031) );
  AO22X1_HVT U2284 ( .A1(\ram[15][129] ), .A2(n5370), .A3(n5371), .A4(
        data[129]), .Y(n4030) );
  AO22X1_HVT U2285 ( .A1(\ram[1][86] ), .A2(n5368), .A3(n5369), .A4(data[86]), 
        .Y(n403) );
  AO22X1_HVT U2286 ( .A1(\ram[15][128] ), .A2(n5370), .A3(n5371), .A4(
        data[128]), .Y(n4029) );
  AO22X1_HVT U2287 ( .A1(\ram[15][127] ), .A2(n5370), .A3(n5371), .A4(
        data[127]), .Y(n4028) );
  AO22X1_HVT U2288 ( .A1(\ram[15][126] ), .A2(n5370), .A3(n5371), .A4(
        data[126]), .Y(n4027) );
  AO22X1_HVT U2289 ( .A1(\ram[15][125] ), .A2(n5370), .A3(n5371), .A4(
        data[125]), .Y(n4026) );
  AO22X1_HVT U2290 ( .A1(\ram[15][124] ), .A2(n5370), .A3(n5371), .A4(
        data[124]), .Y(n4025) );
  AO22X1_HVT U2291 ( .A1(\ram[15][123] ), .A2(n5370), .A3(n5371), .A4(
        data[123]), .Y(n4024) );
  AO22X1_HVT U2292 ( .A1(\ram[15][122] ), .A2(n5370), .A3(n5371), .A4(
        data[122]), .Y(n4023) );
  AO22X1_HVT U2293 ( .A1(\ram[15][121] ), .A2(n5370), .A3(n5371), .A4(
        data[121]), .Y(n4022) );
  AO22X1_HVT U2294 ( .A1(\ram[15][120] ), .A2(n5370), .A3(n5371), .A4(
        data[120]), .Y(n4021) );
  AO22X1_HVT U2295 ( .A1(\ram[15][119] ), .A2(n5370), .A3(n5371), .A4(
        data[119]), .Y(n4020) );
  AO22X1_HVT U2296 ( .A1(\ram[1][85] ), .A2(n5368), .A3(n5369), .A4(data[85]), 
        .Y(n402) );
  AO22X1_HVT U2297 ( .A1(\ram[15][118] ), .A2(n5370), .A3(n5371), .A4(
        data[118]), .Y(n4019) );
  AO22X1_HVT U2298 ( .A1(\ram[15][117] ), .A2(n5370), .A3(n5371), .A4(
        data[117]), .Y(n4018) );
  AO22X1_HVT U2299 ( .A1(\ram[15][116] ), .A2(n5370), .A3(n5371), .A4(
        data[116]), .Y(n4017) );
  AO22X1_HVT U2300 ( .A1(\ram[15][115] ), .A2(n5370), .A3(n5371), .A4(
        data[115]), .Y(n4016) );
  AO22X1_HVT U2301 ( .A1(\ram[15][114] ), .A2(n5370), .A3(n5371), .A4(
        data[114]), .Y(n4015) );
  AO22X1_HVT U2302 ( .A1(\ram[15][113] ), .A2(n5370), .A3(n5371), .A4(
        data[113]), .Y(n4014) );
  AO22X1_HVT U2303 ( .A1(\ram[15][112] ), .A2(n5370), .A3(n5371), .A4(
        data[112]), .Y(n4013) );
  AO22X1_HVT U2304 ( .A1(\ram[15][111] ), .A2(n5370), .A3(n5371), .A4(
        data[111]), .Y(n4012) );
  AO22X1_HVT U2305 ( .A1(\ram[15][110] ), .A2(n5370), .A3(n5371), .A4(
        data[110]), .Y(n4011) );
  AO22X1_HVT U2306 ( .A1(\ram[15][109] ), .A2(n5370), .A3(n5371), .A4(
        data[109]), .Y(n4010) );
  AO22X1_HVT U2307 ( .A1(\ram[1][84] ), .A2(n5368), .A3(n5369), .A4(data[84]), 
        .Y(n401) );
  AO22X1_HVT U2308 ( .A1(\ram[15][108] ), .A2(n5370), .A3(n5371), .A4(
        data[108]), .Y(n4009) );
  AO22X1_HVT U2309 ( .A1(\ram[15][107] ), .A2(n5370), .A3(n5371), .A4(
        data[107]), .Y(n4008) );
  AO22X1_HVT U2310 ( .A1(\ram[15][106] ), .A2(n5370), .A3(n5371), .A4(
        data[106]), .Y(n4007) );
  AO22X1_HVT U2311 ( .A1(\ram[15][105] ), .A2(n5370), .A3(n5371), .A4(
        data[105]), .Y(n4006) );
  AO22X1_HVT U2312 ( .A1(\ram[15][104] ), .A2(n5370), .A3(n5371), .A4(
        data[104]), .Y(n4005) );
  AO22X1_HVT U2313 ( .A1(\ram[15][103] ), .A2(n5370), .A3(n5371), .A4(
        data[103]), .Y(n4004) );
  AO22X1_HVT U2314 ( .A1(\ram[15][102] ), .A2(n5370), .A3(n5371), .A4(
        data[102]), .Y(n4003) );
  AO22X1_HVT U2315 ( .A1(\ram[15][101] ), .A2(n5370), .A3(n5371), .A4(
        data[101]), .Y(n4002) );
  AO22X1_HVT U2316 ( .A1(\ram[15][100] ), .A2(n5370), .A3(n5371), .A4(
        data[100]), .Y(n4001) );
  AO22X1_HVT U2317 ( .A1(\ram[15][99] ), .A2(n5370), .A3(n5371), .A4(data[99]), 
        .Y(n4000) );
  AO22X1_HVT U2318 ( .A1(\ram[1][83] ), .A2(n5368), .A3(n5369), .A4(data[83]), 
        .Y(n400) );
  AO22X1_HVT U2319 ( .A1(\ram[15][98] ), .A2(n5370), .A3(n5371), .A4(data[98]), 
        .Y(n3999) );
  AO22X1_HVT U2320 ( .A1(\ram[15][97] ), .A2(n5370), .A3(n5371), .A4(data[97]), 
        .Y(n3998) );
  AO22X1_HVT U2321 ( .A1(\ram[15][96] ), .A2(n5370), .A3(n5371), .A4(data[96]), 
        .Y(n3997) );
  AO22X1_HVT U2322 ( .A1(\ram[15][95] ), .A2(n5370), .A3(n5371), .A4(data[95]), 
        .Y(n3996) );
  AO22X1_HVT U2323 ( .A1(\ram[15][94] ), .A2(n5370), .A3(n5371), .A4(data[94]), 
        .Y(n3995) );
  AO22X1_HVT U2324 ( .A1(\ram[15][93] ), .A2(n5370), .A3(n5371), .A4(data[93]), 
        .Y(n3994) );
  AO22X1_HVT U2325 ( .A1(\ram[15][92] ), .A2(n5370), .A3(n5371), .A4(data[92]), 
        .Y(n3993) );
  AO22X1_HVT U2326 ( .A1(\ram[15][91] ), .A2(n5370), .A3(n5371), .A4(data[91]), 
        .Y(n3992) );
  AO22X1_HVT U2327 ( .A1(\ram[15][90] ), .A2(n5370), .A3(n5371), .A4(data[90]), 
        .Y(n3991) );
  AO22X1_HVT U2328 ( .A1(\ram[15][89] ), .A2(n5370), .A3(n5371), .A4(data[89]), 
        .Y(n3990) );
  AO22X1_HVT U2329 ( .A1(\ram[1][82] ), .A2(n5368), .A3(n5369), .A4(data[82]), 
        .Y(n399) );
  AO22X1_HVT U2330 ( .A1(\ram[15][88] ), .A2(n5370), .A3(n5371), .A4(data[88]), 
        .Y(n3989) );
  AO22X1_HVT U2331 ( .A1(\ram[15][87] ), .A2(n5370), .A3(n5371), .A4(data[87]), 
        .Y(n3988) );
  AO22X1_HVT U2332 ( .A1(\ram[15][86] ), .A2(n5370), .A3(n5371), .A4(data[86]), 
        .Y(n3987) );
  AO22X1_HVT U2333 ( .A1(\ram[15][85] ), .A2(n5370), .A3(n5371), .A4(data[85]), 
        .Y(n3986) );
  AO22X1_HVT U2334 ( .A1(\ram[15][84] ), .A2(n5370), .A3(n5371), .A4(data[84]), 
        .Y(n3985) );
  AO22X1_HVT U2335 ( .A1(\ram[15][83] ), .A2(n5370), .A3(n5371), .A4(data[83]), 
        .Y(n3984) );
  AO22X1_HVT U2336 ( .A1(\ram[15][82] ), .A2(n5370), .A3(n5371), .A4(data[82]), 
        .Y(n3983) );
  AO22X1_HVT U2337 ( .A1(\ram[15][81] ), .A2(n5370), .A3(n5371), .A4(data[81]), 
        .Y(n3982) );
  AO22X1_HVT U2338 ( .A1(\ram[15][80] ), .A2(n5370), .A3(n5371), .A4(data[80]), 
        .Y(n3981) );
  AO22X1_HVT U2339 ( .A1(\ram[15][79] ), .A2(n5370), .A3(n5371), .A4(data[79]), 
        .Y(n3980) );
  AO22X1_HVT U2340 ( .A1(\ram[1][81] ), .A2(n5368), .A3(n5369), .A4(data[81]), 
        .Y(n398) );
  AO22X1_HVT U2341 ( .A1(\ram[15][78] ), .A2(n5370), .A3(n5371), .A4(data[78]), 
        .Y(n3979) );
  AO22X1_HVT U2342 ( .A1(\ram[15][77] ), .A2(n5370), .A3(n5371), .A4(data[77]), 
        .Y(n3978) );
  AO22X1_HVT U2343 ( .A1(\ram[15][76] ), .A2(n5370), .A3(n5371), .A4(data[76]), 
        .Y(n3977) );
  AO22X1_HVT U2344 ( .A1(\ram[15][75] ), .A2(n5370), .A3(n5371), .A4(data[75]), 
        .Y(n3976) );
  AO22X1_HVT U2345 ( .A1(\ram[15][74] ), .A2(n5370), .A3(n5371), .A4(data[74]), 
        .Y(n3975) );
  AO22X1_HVT U2346 ( .A1(\ram[15][73] ), .A2(n5370), .A3(n5371), .A4(data[73]), 
        .Y(n3974) );
  AO22X1_HVT U2347 ( .A1(\ram[15][72] ), .A2(n5370), .A3(n5371), .A4(data[72]), 
        .Y(n3973) );
  AO22X1_HVT U2348 ( .A1(\ram[15][71] ), .A2(n5370), .A3(n5371), .A4(data[71]), 
        .Y(n3972) );
  AO22X1_HVT U2349 ( .A1(\ram[15][70] ), .A2(n5370), .A3(n5371), .A4(data[70]), 
        .Y(n3971) );
  AO22X1_HVT U2350 ( .A1(\ram[15][69] ), .A2(n5370), .A3(n5371), .A4(data[69]), 
        .Y(n3970) );
  AO22X1_HVT U2351 ( .A1(\ram[1][80] ), .A2(n5368), .A3(n5369), .A4(data[80]), 
        .Y(n397) );
  AO22X1_HVT U2352 ( .A1(\ram[15][68] ), .A2(n5370), .A3(n5371), .A4(data[68]), 
        .Y(n3969) );
  AO22X1_HVT U2353 ( .A1(\ram[15][67] ), .A2(n5370), .A3(n5371), .A4(data[67]), 
        .Y(n3968) );
  AO22X1_HVT U2354 ( .A1(\ram[15][66] ), .A2(n5370), .A3(n5371), .A4(data[66]), 
        .Y(n3967) );
  AO22X1_HVT U2355 ( .A1(\ram[15][65] ), .A2(n5370), .A3(n5371), .A4(data[65]), 
        .Y(n3966) );
  AO22X1_HVT U2356 ( .A1(\ram[15][64] ), .A2(n5370), .A3(n5371), .A4(data[64]), 
        .Y(n3965) );
  AO22X1_HVT U2357 ( .A1(\ram[15][63] ), .A2(n5370), .A3(n5371), .A4(data[63]), 
        .Y(n3964) );
  AO22X1_HVT U2358 ( .A1(\ram[15][62] ), .A2(n5370), .A3(n5371), .A4(data[62]), 
        .Y(n3963) );
  AO22X1_HVT U2359 ( .A1(\ram[15][61] ), .A2(n5370), .A3(n5371), .A4(data[61]), 
        .Y(n3962) );
  AO22X1_HVT U2360 ( .A1(\ram[15][60] ), .A2(n5370), .A3(n5371), .A4(data[60]), 
        .Y(n3961) );
  AO22X1_HVT U2361 ( .A1(\ram[15][59] ), .A2(n5370), .A3(n5371), .A4(data[59]), 
        .Y(n3960) );
  AO22X1_HVT U2362 ( .A1(\ram[1][79] ), .A2(n5368), .A3(n5369), .A4(data[79]), 
        .Y(n396) );
  AO22X1_HVT U2363 ( .A1(\ram[15][58] ), .A2(n5370), .A3(n5371), .A4(data[58]), 
        .Y(n3959) );
  AO22X1_HVT U2364 ( .A1(\ram[15][57] ), .A2(n5370), .A3(n5371), .A4(data[57]), 
        .Y(n3958) );
  AO22X1_HVT U2365 ( .A1(\ram[15][56] ), .A2(n5370), .A3(n5371), .A4(data[56]), 
        .Y(n3957) );
  AO22X1_HVT U2366 ( .A1(\ram[15][55] ), .A2(n5370), .A3(n5371), .A4(data[55]), 
        .Y(n3956) );
  AO22X1_HVT U2367 ( .A1(\ram[15][54] ), .A2(n5370), .A3(n5371), .A4(data[54]), 
        .Y(n3955) );
  AO22X1_HVT U2368 ( .A1(\ram[15][53] ), .A2(n5370), .A3(n5371), .A4(data[53]), 
        .Y(n3954) );
  AO22X1_HVT U2369 ( .A1(\ram[15][52] ), .A2(n5370), .A3(n5371), .A4(data[52]), 
        .Y(n3953) );
  AO22X1_HVT U2370 ( .A1(\ram[15][51] ), .A2(n5370), .A3(n5371), .A4(data[51]), 
        .Y(n3952) );
  AO22X1_HVT U2371 ( .A1(\ram[15][50] ), .A2(n5370), .A3(n5371), .A4(data[50]), 
        .Y(n3951) );
  AO22X1_HVT U2372 ( .A1(\ram[15][49] ), .A2(n5370), .A3(n5371), .A4(data[49]), 
        .Y(n3950) );
  AO22X1_HVT U2373 ( .A1(\ram[1][78] ), .A2(n5368), .A3(n5369), .A4(data[78]), 
        .Y(n395) );
  AO22X1_HVT U2374 ( .A1(\ram[15][48] ), .A2(n5370), .A3(n5371), .A4(data[48]), 
        .Y(n3949) );
  AO22X1_HVT U2375 ( .A1(\ram[15][47] ), .A2(n5370), .A3(n5371), .A4(data[47]), 
        .Y(n3948) );
  AO22X1_HVT U2376 ( .A1(\ram[15][46] ), .A2(n5370), .A3(n5371), .A4(data[46]), 
        .Y(n3947) );
  AO22X1_HVT U2377 ( .A1(\ram[15][45] ), .A2(n5370), .A3(n5371), .A4(data[45]), 
        .Y(n3946) );
  AO22X1_HVT U2378 ( .A1(\ram[15][44] ), .A2(n5370), .A3(n5371), .A4(data[44]), 
        .Y(n3945) );
  AO22X1_HVT U2379 ( .A1(\ram[15][43] ), .A2(n5370), .A3(n5371), .A4(data[43]), 
        .Y(n3944) );
  AO22X1_HVT U2380 ( .A1(\ram[15][42] ), .A2(n5370), .A3(n5371), .A4(data[42]), 
        .Y(n3943) );
  AO22X1_HVT U2381 ( .A1(\ram[15][41] ), .A2(n5370), .A3(n5371), .A4(data[41]), 
        .Y(n3942) );
  AO22X1_HVT U2382 ( .A1(\ram[15][40] ), .A2(n5370), .A3(n5371), .A4(data[40]), 
        .Y(n3941) );
  AO22X1_HVT U2383 ( .A1(\ram[15][39] ), .A2(n5370), .A3(n5371), .A4(data[39]), 
        .Y(n3940) );
  AO22X1_HVT U2384 ( .A1(\ram[1][77] ), .A2(n5368), .A3(n5369), .A4(data[77]), 
        .Y(n394) );
  AO22X1_HVT U2385 ( .A1(\ram[15][38] ), .A2(n5370), .A3(n5371), .A4(data[38]), 
        .Y(n3939) );
  AO22X1_HVT U2386 ( .A1(\ram[15][37] ), .A2(n5370), .A3(n5371), .A4(data[37]), 
        .Y(n3938) );
  AO22X1_HVT U2387 ( .A1(\ram[15][36] ), .A2(n5370), .A3(n5371), .A4(data[36]), 
        .Y(n3937) );
  AO22X1_HVT U2388 ( .A1(\ram[15][35] ), .A2(n5370), .A3(n5371), .A4(data[35]), 
        .Y(n3936) );
  AO22X1_HVT U2389 ( .A1(\ram[15][34] ), .A2(n5370), .A3(n5371), .A4(data[34]), 
        .Y(n3935) );
  AO22X1_HVT U2390 ( .A1(\ram[15][33] ), .A2(n5370), .A3(n5371), .A4(data[33]), 
        .Y(n3934) );
  AO22X1_HVT U2391 ( .A1(\ram[15][32] ), .A2(n5370), .A3(n5371), .A4(data[32]), 
        .Y(n3933) );
  AO22X1_HVT U2392 ( .A1(\ram[15][31] ), .A2(n5370), .A3(n5371), .A4(data[31]), 
        .Y(n3932) );
  AO22X1_HVT U2393 ( .A1(\ram[15][30] ), .A2(n5370), .A3(n5371), .A4(data[30]), 
        .Y(n3931) );
  AO22X1_HVT U2394 ( .A1(\ram[15][29] ), .A2(n5370), .A3(n5371), .A4(data[29]), 
        .Y(n3930) );
  AO22X1_HVT U2395 ( .A1(\ram[1][76] ), .A2(n5368), .A3(n5369), .A4(data[76]), 
        .Y(n393) );
  AO22X1_HVT U2396 ( .A1(\ram[15][28] ), .A2(n5370), .A3(n5371), .A4(data[28]), 
        .Y(n3929) );
  AO22X1_HVT U2397 ( .A1(\ram[15][27] ), .A2(n5370), .A3(n5371), .A4(data[27]), 
        .Y(n3928) );
  AO22X1_HVT U2398 ( .A1(\ram[15][26] ), .A2(n5370), .A3(n5371), .A4(data[26]), 
        .Y(n3927) );
  AO22X1_HVT U2399 ( .A1(\ram[15][25] ), .A2(n5370), .A3(n5371), .A4(data[25]), 
        .Y(n3926) );
  AO22X1_HVT U2400 ( .A1(\ram[15][24] ), .A2(n5370), .A3(n5371), .A4(data[24]), 
        .Y(n3925) );
  AO22X1_HVT U2401 ( .A1(\ram[15][23] ), .A2(n5370), .A3(n5371), .A4(data[23]), 
        .Y(n3924) );
  AO22X1_HVT U2402 ( .A1(\ram[15][22] ), .A2(n5370), .A3(n5371), .A4(data[22]), 
        .Y(n3923) );
  AO22X1_HVT U2403 ( .A1(\ram[15][21] ), .A2(n5370), .A3(n5371), .A4(data[21]), 
        .Y(n3922) );
  AO22X1_HVT U2404 ( .A1(\ram[15][20] ), .A2(n5370), .A3(n5371), .A4(data[20]), 
        .Y(n3921) );
  AO22X1_HVT U2405 ( .A1(\ram[15][19] ), .A2(n5370), .A3(n5371), .A4(data[19]), 
        .Y(n3920) );
  AO22X1_HVT U2406 ( .A1(\ram[1][75] ), .A2(n5368), .A3(n5369), .A4(data[75]), 
        .Y(n392) );
  AO22X1_HVT U2407 ( .A1(\ram[15][18] ), .A2(n5370), .A3(n5371), .A4(data[18]), 
        .Y(n3919) );
  AO22X1_HVT U2408 ( .A1(\ram[15][17] ), .A2(n5370), .A3(n5371), .A4(data[17]), 
        .Y(n3918) );
  AO22X1_HVT U2409 ( .A1(\ram[15][16] ), .A2(n5370), .A3(n5371), .A4(data[16]), 
        .Y(n3917) );
  AO22X1_HVT U2410 ( .A1(\ram[15][15] ), .A2(n5370), .A3(n5371), .A4(data[15]), 
        .Y(n3916) );
  AO22X1_HVT U2411 ( .A1(\ram[15][14] ), .A2(n5370), .A3(n5371), .A4(data[14]), 
        .Y(n3915) );
  AO22X1_HVT U2412 ( .A1(\ram[15][13] ), .A2(n5370), .A3(n5371), .A4(data[13]), 
        .Y(n3914) );
  AO22X1_HVT U2413 ( .A1(\ram[15][12] ), .A2(n5370), .A3(n5371), .A4(data[12]), 
        .Y(n3913) );
  AO22X1_HVT U2414 ( .A1(\ram[15][11] ), .A2(n5370), .A3(n5371), .A4(data[11]), 
        .Y(n3912) );
  AO22X1_HVT U2415 ( .A1(\ram[15][10] ), .A2(n5370), .A3(n5371), .A4(data[10]), 
        .Y(n3911) );
  AO22X1_HVT U2416 ( .A1(\ram[15][9] ), .A2(n5370), .A3(n5371), .A4(data[9]), 
        .Y(n3910) );
  AO22X1_HVT U2417 ( .A1(\ram[1][74] ), .A2(n5368), .A3(n5369), .A4(data[74]), 
        .Y(n391) );
  AO22X1_HVT U2418 ( .A1(\ram[15][8] ), .A2(n5370), .A3(n5371), .A4(data[8]), 
        .Y(n3909) );
  AO22X1_HVT U2419 ( .A1(\ram[15][7] ), .A2(n5370), .A3(n5371), .A4(data[7]), 
        .Y(n3908) );
  AO22X1_HVT U2420 ( .A1(\ram[15][6] ), .A2(n5370), .A3(n5371), .A4(data[6]), 
        .Y(n3907) );
  AO22X1_HVT U2421 ( .A1(\ram[15][5] ), .A2(n5370), .A3(n5371), .A4(data[5]), 
        .Y(n3906) );
  AO22X1_HVT U2422 ( .A1(\ram[15][4] ), .A2(n5370), .A3(n5371), .A4(data[4]), 
        .Y(n3905) );
  AO22X1_HVT U2423 ( .A1(\ram[15][3] ), .A2(n5370), .A3(n5371), .A4(data[3]), 
        .Y(n3904) );
  AO22X1_HVT U2424 ( .A1(\ram[15][2] ), .A2(n5370), .A3(n5371), .A4(data[2]), 
        .Y(n3903) );
  AO22X1_HVT U2425 ( .A1(\ram[15][1] ), .A2(n5370), .A3(n5371), .A4(data[1]), 
        .Y(n3902) );
  AO22X1_HVT U2426 ( .A1(\ram[15][0] ), .A2(n5370), .A3(n5371), .A4(data[0]), 
        .Y(n3901) );
  INVX0_HVT U2427 ( .A(n5372), .Y(n5371) );
  AND2X1_HVT U2428 ( .A1(n5372), .A2(n5365), .Y(n5370) );
  NAND3X0_HVT U2429 ( .A1(n4182), .A2(n4276), .A3(n5373), .Y(n5372) );
  AO22X1_HVT U2430 ( .A1(\ram[14][255] ), .A2(n5374), .A3(n5375), .A4(
        data[255]), .Y(n3900) );
  AO22X1_HVT U2431 ( .A1(\ram[1][73] ), .A2(n5368), .A3(n5369), .A4(data[73]), 
        .Y(n390) );
  AO22X1_HVT U2432 ( .A1(\ram[14][254] ), .A2(n5374), .A3(n5375), .A4(
        data[254]), .Y(n3899) );
  AO22X1_HVT U2433 ( .A1(\ram[14][253] ), .A2(n5374), .A3(n5375), .A4(
        data[253]), .Y(n3898) );
  AO22X1_HVT U2434 ( .A1(\ram[14][252] ), .A2(n5374), .A3(n5375), .A4(
        data[252]), .Y(n3897) );
  AO22X1_HVT U2435 ( .A1(\ram[14][251] ), .A2(n5374), .A3(n5375), .A4(
        data[251]), .Y(n3896) );
  AO22X1_HVT U2436 ( .A1(\ram[14][250] ), .A2(n5374), .A3(n5375), .A4(
        data[250]), .Y(n3895) );
  AO22X1_HVT U2437 ( .A1(\ram[14][249] ), .A2(n5374), .A3(n5375), .A4(
        data[249]), .Y(n3894) );
  AO22X1_HVT U2438 ( .A1(\ram[14][248] ), .A2(n5374), .A3(n5375), .A4(
        data[248]), .Y(n3893) );
  AO22X1_HVT U2439 ( .A1(\ram[14][247] ), .A2(n5374), .A3(n5375), .A4(
        data[247]), .Y(n3892) );
  AO22X1_HVT U2440 ( .A1(\ram[14][246] ), .A2(n5374), .A3(n5375), .A4(
        data[246]), .Y(n3891) );
  AO22X1_HVT U2441 ( .A1(\ram[14][245] ), .A2(n5374), .A3(n5375), .A4(
        data[245]), .Y(n3890) );
  AO22X1_HVT U2442 ( .A1(\ram[1][72] ), .A2(n5368), .A3(n5369), .A4(data[72]), 
        .Y(n389) );
  AO22X1_HVT U2443 ( .A1(\ram[14][244] ), .A2(n5374), .A3(n5375), .A4(
        data[244]), .Y(n3889) );
  AO22X1_HVT U2444 ( .A1(\ram[14][243] ), .A2(n5374), .A3(n5375), .A4(
        data[243]), .Y(n3888) );
  AO22X1_HVT U2445 ( .A1(\ram[14][242] ), .A2(n5374), .A3(n5375), .A4(
        data[242]), .Y(n3887) );
  AO22X1_HVT U2446 ( .A1(\ram[14][241] ), .A2(n5374), .A3(n5375), .A4(
        data[241]), .Y(n3886) );
  AO22X1_HVT U2447 ( .A1(\ram[14][240] ), .A2(n5374), .A3(n5375), .A4(
        data[240]), .Y(n3885) );
  AO22X1_HVT U2448 ( .A1(\ram[14][239] ), .A2(n5374), .A3(n5375), .A4(
        data[239]), .Y(n3884) );
  AO22X1_HVT U2449 ( .A1(\ram[14][238] ), .A2(n5374), .A3(n5375), .A4(
        data[238]), .Y(n3883) );
  AO22X1_HVT U2450 ( .A1(\ram[14][237] ), .A2(n5374), .A3(n5375), .A4(
        data[237]), .Y(n3882) );
  AO22X1_HVT U2451 ( .A1(\ram[14][236] ), .A2(n5374), .A3(n5375), .A4(
        data[236]), .Y(n3881) );
  AO22X1_HVT U2452 ( .A1(\ram[14][235] ), .A2(n5374), .A3(n5375), .A4(
        data[235]), .Y(n3880) );
  AO22X1_HVT U2453 ( .A1(\ram[1][71] ), .A2(n5368), .A3(n5369), .A4(data[71]), 
        .Y(n388) );
  AO22X1_HVT U2454 ( .A1(\ram[14][234] ), .A2(n5374), .A3(n5375), .A4(
        data[234]), .Y(n3879) );
  AO22X1_HVT U2455 ( .A1(\ram[14][233] ), .A2(n5374), .A3(n5375), .A4(
        data[233]), .Y(n3878) );
  AO22X1_HVT U2456 ( .A1(\ram[14][232] ), .A2(n5374), .A3(n5375), .A4(
        data[232]), .Y(n3877) );
  AO22X1_HVT U2457 ( .A1(\ram[14][231] ), .A2(n5374), .A3(n5375), .A4(
        data[231]), .Y(n3876) );
  AO22X1_HVT U2458 ( .A1(\ram[14][230] ), .A2(n5374), .A3(n5375), .A4(
        data[230]), .Y(n3875) );
  AO22X1_HVT U2459 ( .A1(\ram[14][229] ), .A2(n5374), .A3(n5375), .A4(
        data[229]), .Y(n3874) );
  AO22X1_HVT U2460 ( .A1(\ram[14][228] ), .A2(n5374), .A3(n5375), .A4(
        data[228]), .Y(n3873) );
  AO22X1_HVT U2461 ( .A1(\ram[14][227] ), .A2(n5374), .A3(n5375), .A4(
        data[227]), .Y(n3872) );
  AO22X1_HVT U2462 ( .A1(\ram[14][226] ), .A2(n5374), .A3(n5375), .A4(
        data[226]), .Y(n3871) );
  AO22X1_HVT U2463 ( .A1(\ram[14][225] ), .A2(n5374), .A3(n5375), .A4(
        data[225]), .Y(n3870) );
  AO22X1_HVT U2464 ( .A1(\ram[1][70] ), .A2(n5368), .A3(n5369), .A4(data[70]), 
        .Y(n387) );
  AO22X1_HVT U2465 ( .A1(\ram[14][224] ), .A2(n5374), .A3(n5375), .A4(
        data[224]), .Y(n3869) );
  AO22X1_HVT U2466 ( .A1(\ram[14][223] ), .A2(n5374), .A3(n5375), .A4(
        data[223]), .Y(n3868) );
  AO22X1_HVT U2467 ( .A1(\ram[14][222] ), .A2(n5374), .A3(n5375), .A4(
        data[222]), .Y(n3867) );
  AO22X1_HVT U2468 ( .A1(\ram[14][221] ), .A2(n5374), .A3(n5375), .A4(
        data[221]), .Y(n3866) );
  AO22X1_HVT U2469 ( .A1(\ram[14][220] ), .A2(n5374), .A3(n5375), .A4(
        data[220]), .Y(n3865) );
  AO22X1_HVT U2470 ( .A1(\ram[14][219] ), .A2(n5374), .A3(n5375), .A4(
        data[219]), .Y(n3864) );
  AO22X1_HVT U2471 ( .A1(\ram[14][218] ), .A2(n5374), .A3(n5375), .A4(
        data[218]), .Y(n3863) );
  AO22X1_HVT U2472 ( .A1(\ram[14][217] ), .A2(n5374), .A3(n5375), .A4(
        data[217]), .Y(n3862) );
  AO22X1_HVT U2473 ( .A1(\ram[14][216] ), .A2(n5374), .A3(n5375), .A4(
        data[216]), .Y(n3861) );
  AO22X1_HVT U2474 ( .A1(\ram[14][215] ), .A2(n5374), .A3(n5375), .A4(
        data[215]), .Y(n3860) );
  AO22X1_HVT U2475 ( .A1(\ram[1][69] ), .A2(n5368), .A3(n5369), .A4(data[69]), 
        .Y(n386) );
  AO22X1_HVT U2476 ( .A1(\ram[14][214] ), .A2(n5374), .A3(n5375), .A4(
        data[214]), .Y(n3859) );
  AO22X1_HVT U2477 ( .A1(\ram[14][213] ), .A2(n5374), .A3(n5375), .A4(
        data[213]), .Y(n3858) );
  AO22X1_HVT U2478 ( .A1(\ram[14][212] ), .A2(n5374), .A3(n5375), .A4(
        data[212]), .Y(n3857) );
  AO22X1_HVT U2479 ( .A1(\ram[14][211] ), .A2(n5374), .A3(n5375), .A4(
        data[211]), .Y(n3856) );
  AO22X1_HVT U2480 ( .A1(\ram[14][210] ), .A2(n5374), .A3(n5375), .A4(
        data[210]), .Y(n3855) );
  AO22X1_HVT U2481 ( .A1(\ram[14][209] ), .A2(n5374), .A3(n5375), .A4(
        data[209]), .Y(n3854) );
  AO22X1_HVT U2482 ( .A1(\ram[14][208] ), .A2(n5374), .A3(n5375), .A4(
        data[208]), .Y(n3853) );
  AO22X1_HVT U2483 ( .A1(\ram[14][207] ), .A2(n5374), .A3(n5375), .A4(
        data[207]), .Y(n3852) );
  AO22X1_HVT U2484 ( .A1(\ram[14][206] ), .A2(n5374), .A3(n5375), .A4(
        data[206]), .Y(n3851) );
  AO22X1_HVT U2485 ( .A1(\ram[14][205] ), .A2(n5374), .A3(n5375), .A4(
        data[205]), .Y(n3850) );
  AO22X1_HVT U2486 ( .A1(\ram[1][68] ), .A2(n5368), .A3(n5369), .A4(data[68]), 
        .Y(n385) );
  AO22X1_HVT U2487 ( .A1(\ram[14][204] ), .A2(n5374), .A3(n5375), .A4(
        data[204]), .Y(n3849) );
  AO22X1_HVT U2488 ( .A1(\ram[14][203] ), .A2(n5374), .A3(n5375), .A4(
        data[203]), .Y(n3848) );
  AO22X1_HVT U2489 ( .A1(\ram[14][202] ), .A2(n5374), .A3(n5375), .A4(
        data[202]), .Y(n3847) );
  AO22X1_HVT U2490 ( .A1(\ram[14][201] ), .A2(n5374), .A3(n5375), .A4(
        data[201]), .Y(n3846) );
  AO22X1_HVT U2491 ( .A1(\ram[14][200] ), .A2(n5374), .A3(n5375), .A4(
        data[200]), .Y(n3845) );
  AO22X1_HVT U2492 ( .A1(\ram[14][199] ), .A2(n5374), .A3(n5375), .A4(
        data[199]), .Y(n3844) );
  AO22X1_HVT U2493 ( .A1(\ram[14][198] ), .A2(n5374), .A3(n5375), .A4(
        data[198]), .Y(n3843) );
  AO22X1_HVT U2494 ( .A1(\ram[14][197] ), .A2(n5374), .A3(n5375), .A4(
        data[197]), .Y(n3842) );
  AO22X1_HVT U2495 ( .A1(\ram[14][196] ), .A2(n5374), .A3(n5375), .A4(
        data[196]), .Y(n3841) );
  AO22X1_HVT U2496 ( .A1(\ram[14][195] ), .A2(n5374), .A3(n5375), .A4(
        data[195]), .Y(n3840) );
  AO22X1_HVT U2497 ( .A1(\ram[1][67] ), .A2(n5368), .A3(n5369), .A4(data[67]), 
        .Y(n384) );
  AO22X1_HVT U2498 ( .A1(\ram[14][194] ), .A2(n5374), .A3(n5375), .A4(
        data[194]), .Y(n3839) );
  AO22X1_HVT U2499 ( .A1(\ram[14][193] ), .A2(n5374), .A3(n5375), .A4(
        data[193]), .Y(n3838) );
  AO22X1_HVT U2500 ( .A1(\ram[14][192] ), .A2(n5374), .A3(n5375), .A4(
        data[192]), .Y(n3837) );
  AO22X1_HVT U2501 ( .A1(\ram[14][191] ), .A2(n5374), .A3(n5375), .A4(
        data[191]), .Y(n3836) );
  AO22X1_HVT U2502 ( .A1(\ram[14][190] ), .A2(n5374), .A3(n5375), .A4(
        data[190]), .Y(n3835) );
  AO22X1_HVT U2503 ( .A1(\ram[14][189] ), .A2(n5374), .A3(n5375), .A4(
        data[189]), .Y(n3834) );
  AO22X1_HVT U2504 ( .A1(\ram[14][188] ), .A2(n5374), .A3(n5375), .A4(
        data[188]), .Y(n3833) );
  AO22X1_HVT U2505 ( .A1(\ram[14][187] ), .A2(n5374), .A3(n5375), .A4(
        data[187]), .Y(n3832) );
  AO22X1_HVT U2506 ( .A1(\ram[14][186] ), .A2(n5374), .A3(n5375), .A4(
        data[186]), .Y(n3831) );
  AO22X1_HVT U2507 ( .A1(\ram[14][185] ), .A2(n5374), .A3(n5375), .A4(
        data[185]), .Y(n3830) );
  AO22X1_HVT U2508 ( .A1(\ram[1][66] ), .A2(n5368), .A3(n5369), .A4(data[66]), 
        .Y(n383) );
  AO22X1_HVT U2509 ( .A1(\ram[14][184] ), .A2(n5374), .A3(n5375), .A4(
        data[184]), .Y(n3829) );
  AO22X1_HVT U2510 ( .A1(\ram[14][183] ), .A2(n5374), .A3(n5375), .A4(
        data[183]), .Y(n3828) );
  AO22X1_HVT U2511 ( .A1(\ram[14][182] ), .A2(n5374), .A3(n5375), .A4(
        data[182]), .Y(n3827) );
  AO22X1_HVT U2512 ( .A1(\ram[14][181] ), .A2(n5374), .A3(n5375), .A4(
        data[181]), .Y(n3826) );
  AO22X1_HVT U2513 ( .A1(\ram[14][180] ), .A2(n5374), .A3(n5375), .A4(
        data[180]), .Y(n3825) );
  AO22X1_HVT U2514 ( .A1(\ram[14][179] ), .A2(n5374), .A3(n5375), .A4(
        data[179]), .Y(n3824) );
  AO22X1_HVT U2515 ( .A1(\ram[14][178] ), .A2(n5374), .A3(n5375), .A4(
        data[178]), .Y(n3823) );
  AO22X1_HVT U2516 ( .A1(\ram[14][177] ), .A2(n5374), .A3(n5375), .A4(
        data[177]), .Y(n3822) );
  AO22X1_HVT U2517 ( .A1(\ram[14][176] ), .A2(n5374), .A3(n5375), .A4(
        data[176]), .Y(n3821) );
  AO22X1_HVT U2518 ( .A1(\ram[14][175] ), .A2(n5374), .A3(n5375), .A4(
        data[175]), .Y(n3820) );
  AO22X1_HVT U2519 ( .A1(\ram[1][65] ), .A2(n5368), .A3(n5369), .A4(data[65]), 
        .Y(n382) );
  AO22X1_HVT U2520 ( .A1(\ram[14][174] ), .A2(n5374), .A3(n5375), .A4(
        data[174]), .Y(n3819) );
  AO22X1_HVT U2521 ( .A1(\ram[14][173] ), .A2(n5374), .A3(n5375), .A4(
        data[173]), .Y(n3818) );
  AO22X1_HVT U2522 ( .A1(\ram[14][172] ), .A2(n5374), .A3(n5375), .A4(
        data[172]), .Y(n3817) );
  AO22X1_HVT U2523 ( .A1(\ram[14][171] ), .A2(n5374), .A3(n5375), .A4(
        data[171]), .Y(n3816) );
  AO22X1_HVT U2524 ( .A1(\ram[14][170] ), .A2(n5374), .A3(n5375), .A4(
        data[170]), .Y(n3815) );
  AO22X1_HVT U2525 ( .A1(\ram[14][169] ), .A2(n5374), .A3(n5375), .A4(
        data[169]), .Y(n3814) );
  AO22X1_HVT U2526 ( .A1(\ram[14][168] ), .A2(n5374), .A3(n5375), .A4(
        data[168]), .Y(n3813) );
  AO22X1_HVT U2527 ( .A1(\ram[14][167] ), .A2(n5374), .A3(n5375), .A4(
        data[167]), .Y(n3812) );
  AO22X1_HVT U2528 ( .A1(\ram[14][166] ), .A2(n5374), .A3(n5375), .A4(
        data[166]), .Y(n3811) );
  AO22X1_HVT U2529 ( .A1(\ram[14][165] ), .A2(n5374), .A3(n5375), .A4(
        data[165]), .Y(n3810) );
  AO22X1_HVT U2530 ( .A1(\ram[1][64] ), .A2(n5368), .A3(n5369), .A4(data[64]), 
        .Y(n381) );
  AO22X1_HVT U2531 ( .A1(\ram[14][164] ), .A2(n5374), .A3(n5375), .A4(
        data[164]), .Y(n3809) );
  AO22X1_HVT U2532 ( .A1(\ram[14][163] ), .A2(n5374), .A3(n5375), .A4(
        data[163]), .Y(n3808) );
  AO22X1_HVT U2533 ( .A1(\ram[14][162] ), .A2(n5374), .A3(n5375), .A4(
        data[162]), .Y(n3807) );
  AO22X1_HVT U2534 ( .A1(\ram[14][161] ), .A2(n5374), .A3(n5375), .A4(
        data[161]), .Y(n3806) );
  AO22X1_HVT U2535 ( .A1(\ram[14][160] ), .A2(n5374), .A3(n5375), .A4(
        data[160]), .Y(n3805) );
  AO22X1_HVT U2536 ( .A1(\ram[14][159] ), .A2(n5374), .A3(n5375), .A4(
        data[159]), .Y(n3804) );
  AO22X1_HVT U2537 ( .A1(\ram[14][158] ), .A2(n5374), .A3(n5375), .A4(
        data[158]), .Y(n3803) );
  AO22X1_HVT U2538 ( .A1(\ram[14][157] ), .A2(n5374), .A3(n5375), .A4(
        data[157]), .Y(n3802) );
  AO22X1_HVT U2539 ( .A1(\ram[14][156] ), .A2(n5374), .A3(n5375), .A4(
        data[156]), .Y(n3801) );
  AO22X1_HVT U2540 ( .A1(\ram[14][155] ), .A2(n5374), .A3(n5375), .A4(
        data[155]), .Y(n3800) );
  AO22X1_HVT U2541 ( .A1(\ram[1][63] ), .A2(n5368), .A3(n5369), .A4(data[63]), 
        .Y(n380) );
  AO22X1_HVT U2542 ( .A1(\ram[14][154] ), .A2(n5374), .A3(n5375), .A4(
        data[154]), .Y(n3799) );
  AO22X1_HVT U2543 ( .A1(\ram[14][153] ), .A2(n5374), .A3(n5375), .A4(
        data[153]), .Y(n3798) );
  AO22X1_HVT U2544 ( .A1(\ram[14][152] ), .A2(n5374), .A3(n5375), .A4(
        data[152]), .Y(n3797) );
  AO22X1_HVT U2545 ( .A1(\ram[14][151] ), .A2(n5374), .A3(n5375), .A4(
        data[151]), .Y(n3796) );
  AO22X1_HVT U2546 ( .A1(\ram[14][150] ), .A2(n5374), .A3(n5375), .A4(
        data[150]), .Y(n3795) );
  AO22X1_HVT U2547 ( .A1(\ram[14][149] ), .A2(n5374), .A3(n5375), .A4(
        data[149]), .Y(n3794) );
  AO22X1_HVT U2548 ( .A1(\ram[14][148] ), .A2(n5374), .A3(n5375), .A4(
        data[148]), .Y(n3793) );
  AO22X1_HVT U2549 ( .A1(\ram[14][147] ), .A2(n5374), .A3(n5375), .A4(
        data[147]), .Y(n3792) );
  AO22X1_HVT U2550 ( .A1(\ram[14][146] ), .A2(n5374), .A3(n5375), .A4(
        data[146]), .Y(n3791) );
  AO22X1_HVT U2551 ( .A1(\ram[14][145] ), .A2(n5374), .A3(n5375), .A4(
        data[145]), .Y(n3790) );
  AO22X1_HVT U2552 ( .A1(\ram[1][62] ), .A2(n5368), .A3(n5369), .A4(data[62]), 
        .Y(n379) );
  AO22X1_HVT U2553 ( .A1(\ram[14][144] ), .A2(n5374), .A3(n5375), .A4(
        data[144]), .Y(n3789) );
  AO22X1_HVT U2554 ( .A1(\ram[14][143] ), .A2(n5374), .A3(n5375), .A4(
        data[143]), .Y(n3788) );
  AO22X1_HVT U2555 ( .A1(\ram[14][142] ), .A2(n5374), .A3(n5375), .A4(
        data[142]), .Y(n3787) );
  AO22X1_HVT U2556 ( .A1(\ram[14][141] ), .A2(n5374), .A3(n5375), .A4(
        data[141]), .Y(n3786) );
  AO22X1_HVT U2557 ( .A1(\ram[14][140] ), .A2(n5374), .A3(n5375), .A4(
        data[140]), .Y(n3785) );
  AO22X1_HVT U2558 ( .A1(\ram[14][139] ), .A2(n5374), .A3(n5375), .A4(
        data[139]), .Y(n3784) );
  AO22X1_HVT U2559 ( .A1(\ram[14][138] ), .A2(n5374), .A3(n5375), .A4(
        data[138]), .Y(n3783) );
  AO22X1_HVT U2560 ( .A1(\ram[14][137] ), .A2(n5374), .A3(n5375), .A4(
        data[137]), .Y(n3782) );
  AO22X1_HVT U2561 ( .A1(\ram[14][136] ), .A2(n5374), .A3(n5375), .A4(
        data[136]), .Y(n3781) );
  AO22X1_HVT U2562 ( .A1(\ram[14][135] ), .A2(n5374), .A3(n5375), .A4(
        data[135]), .Y(n3780) );
  AO22X1_HVT U2563 ( .A1(\ram[1][61] ), .A2(n5368), .A3(n5369), .A4(data[61]), 
        .Y(n378) );
  AO22X1_HVT U2564 ( .A1(\ram[14][134] ), .A2(n5374), .A3(n5375), .A4(
        data[134]), .Y(n3779) );
  AO22X1_HVT U2565 ( .A1(\ram[14][133] ), .A2(n5374), .A3(n5375), .A4(
        data[133]), .Y(n3778) );
  AO22X1_HVT U2566 ( .A1(\ram[14][132] ), .A2(n5374), .A3(n5375), .A4(
        data[132]), .Y(n3777) );
  AO22X1_HVT U2567 ( .A1(\ram[14][131] ), .A2(n5374), .A3(n5375), .A4(
        data[131]), .Y(n3776) );
  AO22X1_HVT U2568 ( .A1(\ram[14][130] ), .A2(n5374), .A3(n5375), .A4(
        data[130]), .Y(n3775) );
  AO22X1_HVT U2569 ( .A1(\ram[14][129] ), .A2(n5374), .A3(n5375), .A4(
        data[129]), .Y(n3774) );
  AO22X1_HVT U2570 ( .A1(\ram[14][128] ), .A2(n5374), .A3(n5375), .A4(
        data[128]), .Y(n3773) );
  AO22X1_HVT U2571 ( .A1(\ram[14][127] ), .A2(n5374), .A3(n5375), .A4(
        data[127]), .Y(n3772) );
  AO22X1_HVT U2572 ( .A1(\ram[14][126] ), .A2(n5374), .A3(n5375), .A4(
        data[126]), .Y(n3771) );
  AO22X1_HVT U2573 ( .A1(\ram[14][125] ), .A2(n5374), .A3(n5375), .A4(
        data[125]), .Y(n3770) );
  AO22X1_HVT U2574 ( .A1(\ram[1][60] ), .A2(n5368), .A3(n5369), .A4(data[60]), 
        .Y(n377) );
  AO22X1_HVT U2575 ( .A1(\ram[14][124] ), .A2(n5374), .A3(n5375), .A4(
        data[124]), .Y(n3769) );
  AO22X1_HVT U2576 ( .A1(\ram[14][123] ), .A2(n5374), .A3(n5375), .A4(
        data[123]), .Y(n3768) );
  AO22X1_HVT U2577 ( .A1(\ram[14][122] ), .A2(n5374), .A3(n5375), .A4(
        data[122]), .Y(n3767) );
  AO22X1_HVT U2578 ( .A1(\ram[14][121] ), .A2(n5374), .A3(n5375), .A4(
        data[121]), .Y(n3766) );
  AO22X1_HVT U2579 ( .A1(\ram[14][120] ), .A2(n5374), .A3(n5375), .A4(
        data[120]), .Y(n3765) );
  AO22X1_HVT U2580 ( .A1(\ram[14][119] ), .A2(n5374), .A3(n5375), .A4(
        data[119]), .Y(n3764) );
  AO22X1_HVT U2581 ( .A1(\ram[14][118] ), .A2(n5374), .A3(n5375), .A4(
        data[118]), .Y(n3763) );
  AO22X1_HVT U2582 ( .A1(\ram[14][117] ), .A2(n5374), .A3(n5375), .A4(
        data[117]), .Y(n3762) );
  AO22X1_HVT U2583 ( .A1(\ram[14][116] ), .A2(n5374), .A3(n5375), .A4(
        data[116]), .Y(n3761) );
  AO22X1_HVT U2584 ( .A1(\ram[14][115] ), .A2(n5374), .A3(n5375), .A4(
        data[115]), .Y(n3760) );
  AO22X1_HVT U2585 ( .A1(\ram[1][59] ), .A2(n5368), .A3(n5369), .A4(data[59]), 
        .Y(n376) );
  AO22X1_HVT U2586 ( .A1(\ram[14][114] ), .A2(n5374), .A3(n5375), .A4(
        data[114]), .Y(n3759) );
  AO22X1_HVT U2587 ( .A1(\ram[14][113] ), .A2(n5374), .A3(n5375), .A4(
        data[113]), .Y(n3758) );
  AO22X1_HVT U2588 ( .A1(\ram[14][112] ), .A2(n5374), .A3(n5375), .A4(
        data[112]), .Y(n3757) );
  AO22X1_HVT U2589 ( .A1(\ram[14][111] ), .A2(n5374), .A3(n5375), .A4(
        data[111]), .Y(n3756) );
  AO22X1_HVT U2590 ( .A1(\ram[14][110] ), .A2(n5374), .A3(n5375), .A4(
        data[110]), .Y(n3755) );
  AO22X1_HVT U2591 ( .A1(\ram[14][109] ), .A2(n5374), .A3(n5375), .A4(
        data[109]), .Y(n3754) );
  AO22X1_HVT U2592 ( .A1(\ram[14][108] ), .A2(n5374), .A3(n5375), .A4(
        data[108]), .Y(n3753) );
  AO22X1_HVT U2593 ( .A1(\ram[14][107] ), .A2(n5374), .A3(n5375), .A4(
        data[107]), .Y(n3752) );
  AO22X1_HVT U2594 ( .A1(\ram[14][106] ), .A2(n5374), .A3(n5375), .A4(
        data[106]), .Y(n3751) );
  AO22X1_HVT U2595 ( .A1(\ram[14][105] ), .A2(n5374), .A3(n5375), .A4(
        data[105]), .Y(n3750) );
  AO22X1_HVT U2596 ( .A1(\ram[1][58] ), .A2(n5368), .A3(n5369), .A4(data[58]), 
        .Y(n375) );
  AO22X1_HVT U2597 ( .A1(\ram[14][104] ), .A2(n5374), .A3(n5375), .A4(
        data[104]), .Y(n3749) );
  AO22X1_HVT U2598 ( .A1(\ram[14][103] ), .A2(n5374), .A3(n5375), .A4(
        data[103]), .Y(n3748) );
  AO22X1_HVT U2599 ( .A1(\ram[14][102] ), .A2(n5374), .A3(n5375), .A4(
        data[102]), .Y(n3747) );
  AO22X1_HVT U2600 ( .A1(\ram[14][101] ), .A2(n5374), .A3(n5375), .A4(
        data[101]), .Y(n3746) );
  AO22X1_HVT U2601 ( .A1(\ram[14][100] ), .A2(n5374), .A3(n5375), .A4(
        data[100]), .Y(n3745) );
  AO22X1_HVT U2602 ( .A1(\ram[14][99] ), .A2(n5374), .A3(n5375), .A4(data[99]), 
        .Y(n3744) );
  AO22X1_HVT U2603 ( .A1(\ram[14][98] ), .A2(n5374), .A3(n5375), .A4(data[98]), 
        .Y(n3743) );
  AO22X1_HVT U2604 ( .A1(\ram[14][97] ), .A2(n5374), .A3(n5375), .A4(data[97]), 
        .Y(n3742) );
  AO22X1_HVT U2605 ( .A1(\ram[14][96] ), .A2(n5374), .A3(n5375), .A4(data[96]), 
        .Y(n3741) );
  AO22X1_HVT U2606 ( .A1(\ram[14][95] ), .A2(n5374), .A3(n5375), .A4(data[95]), 
        .Y(n3740) );
  AO22X1_HVT U2607 ( .A1(\ram[1][57] ), .A2(n5368), .A3(n5369), .A4(data[57]), 
        .Y(n374) );
  AO22X1_HVT U2608 ( .A1(\ram[14][94] ), .A2(n5374), .A3(n5375), .A4(data[94]), 
        .Y(n3739) );
  AO22X1_HVT U2609 ( .A1(\ram[14][93] ), .A2(n5374), .A3(n5375), .A4(data[93]), 
        .Y(n3738) );
  AO22X1_HVT U2610 ( .A1(\ram[14][92] ), .A2(n5374), .A3(n5375), .A4(data[92]), 
        .Y(n3737) );
  AO22X1_HVT U2611 ( .A1(\ram[14][91] ), .A2(n5374), .A3(n5375), .A4(data[91]), 
        .Y(n3736) );
  AO22X1_HVT U2612 ( .A1(\ram[14][90] ), .A2(n5374), .A3(n5375), .A4(data[90]), 
        .Y(n3735) );
  AO22X1_HVT U2613 ( .A1(\ram[14][89] ), .A2(n5374), .A3(n5375), .A4(data[89]), 
        .Y(n3734) );
  AO22X1_HVT U2614 ( .A1(\ram[14][88] ), .A2(n5374), .A3(n5375), .A4(data[88]), 
        .Y(n3733) );
  AO22X1_HVT U2615 ( .A1(\ram[14][87] ), .A2(n5374), .A3(n5375), .A4(data[87]), 
        .Y(n3732) );
  AO22X1_HVT U2616 ( .A1(\ram[14][86] ), .A2(n5374), .A3(n5375), .A4(data[86]), 
        .Y(n3731) );
  AO22X1_HVT U2617 ( .A1(\ram[14][85] ), .A2(n5374), .A3(n5375), .A4(data[85]), 
        .Y(n3730) );
  AO22X1_HVT U2618 ( .A1(\ram[1][56] ), .A2(n5368), .A3(n5369), .A4(data[56]), 
        .Y(n373) );
  AO22X1_HVT U2619 ( .A1(\ram[14][84] ), .A2(n5374), .A3(n5375), .A4(data[84]), 
        .Y(n3729) );
  AO22X1_HVT U2620 ( .A1(\ram[14][83] ), .A2(n5374), .A3(n5375), .A4(data[83]), 
        .Y(n3728) );
  AO22X1_HVT U2621 ( .A1(\ram[14][82] ), .A2(n5374), .A3(n5375), .A4(data[82]), 
        .Y(n3727) );
  AO22X1_HVT U2622 ( .A1(\ram[14][81] ), .A2(n5374), .A3(n5375), .A4(data[81]), 
        .Y(n3726) );
  AO22X1_HVT U2623 ( .A1(\ram[14][80] ), .A2(n5374), .A3(n5375), .A4(data[80]), 
        .Y(n3725) );
  AO22X1_HVT U2624 ( .A1(\ram[14][79] ), .A2(n5374), .A3(n5375), .A4(data[79]), 
        .Y(n3724) );
  AO22X1_HVT U2625 ( .A1(\ram[14][78] ), .A2(n5374), .A3(n5375), .A4(data[78]), 
        .Y(n3723) );
  AO22X1_HVT U2626 ( .A1(\ram[14][77] ), .A2(n5374), .A3(n5375), .A4(data[77]), 
        .Y(n3722) );
  AO22X1_HVT U2627 ( .A1(\ram[14][76] ), .A2(n5374), .A3(n5375), .A4(data[76]), 
        .Y(n3721) );
  AO22X1_HVT U2628 ( .A1(\ram[14][75] ), .A2(n5374), .A3(n5375), .A4(data[75]), 
        .Y(n3720) );
  AO22X1_HVT U2629 ( .A1(\ram[1][55] ), .A2(n5368), .A3(n5369), .A4(data[55]), 
        .Y(n372) );
  AO22X1_HVT U2630 ( .A1(\ram[14][74] ), .A2(n5374), .A3(n5375), .A4(data[74]), 
        .Y(n3719) );
  AO22X1_HVT U2631 ( .A1(\ram[14][73] ), .A2(n5374), .A3(n5375), .A4(data[73]), 
        .Y(n3718) );
  AO22X1_HVT U2632 ( .A1(\ram[14][72] ), .A2(n5374), .A3(n5375), .A4(data[72]), 
        .Y(n3717) );
  AO22X1_HVT U2633 ( .A1(\ram[14][71] ), .A2(n5374), .A3(n5375), .A4(data[71]), 
        .Y(n3716) );
  AO22X1_HVT U2634 ( .A1(\ram[14][70] ), .A2(n5374), .A3(n5375), .A4(data[70]), 
        .Y(n3715) );
  AO22X1_HVT U2635 ( .A1(\ram[14][69] ), .A2(n5374), .A3(n5375), .A4(data[69]), 
        .Y(n3714) );
  AO22X1_HVT U2636 ( .A1(\ram[14][68] ), .A2(n5374), .A3(n5375), .A4(data[68]), 
        .Y(n3713) );
  AO22X1_HVT U2637 ( .A1(\ram[14][67] ), .A2(n5374), .A3(n5375), .A4(data[67]), 
        .Y(n3712) );
  AO22X1_HVT U2638 ( .A1(\ram[14][66] ), .A2(n5374), .A3(n5375), .A4(data[66]), 
        .Y(n3711) );
  AO22X1_HVT U2639 ( .A1(\ram[14][65] ), .A2(n5374), .A3(n5375), .A4(data[65]), 
        .Y(n3710) );
  AO22X1_HVT U2640 ( .A1(\ram[1][54] ), .A2(n5368), .A3(n5369), .A4(data[54]), 
        .Y(n371) );
  AO22X1_HVT U2641 ( .A1(\ram[14][64] ), .A2(n5374), .A3(n5375), .A4(data[64]), 
        .Y(n3709) );
  AO22X1_HVT U2642 ( .A1(\ram[14][63] ), .A2(n5374), .A3(n5375), .A4(data[63]), 
        .Y(n3708) );
  AO22X1_HVT U2643 ( .A1(\ram[14][62] ), .A2(n5374), .A3(n5375), .A4(data[62]), 
        .Y(n3707) );
  AO22X1_HVT U2644 ( .A1(\ram[14][61] ), .A2(n5374), .A3(n5375), .A4(data[61]), 
        .Y(n3706) );
  AO22X1_HVT U2645 ( .A1(\ram[14][60] ), .A2(n5374), .A3(n5375), .A4(data[60]), 
        .Y(n3705) );
  AO22X1_HVT U2646 ( .A1(\ram[14][59] ), .A2(n5374), .A3(n5375), .A4(data[59]), 
        .Y(n3704) );
  AO22X1_HVT U2647 ( .A1(\ram[14][58] ), .A2(n5374), .A3(n5375), .A4(data[58]), 
        .Y(n3703) );
  AO22X1_HVT U2648 ( .A1(\ram[14][57] ), .A2(n5374), .A3(n5375), .A4(data[57]), 
        .Y(n3702) );
  AO22X1_HVT U2649 ( .A1(\ram[14][56] ), .A2(n5374), .A3(n5375), .A4(data[56]), 
        .Y(n3701) );
  AO22X1_HVT U2650 ( .A1(\ram[14][55] ), .A2(n5374), .A3(n5375), .A4(data[55]), 
        .Y(n3700) );
  AO22X1_HVT U2651 ( .A1(\ram[1][53] ), .A2(n5368), .A3(n5369), .A4(data[53]), 
        .Y(n370) );
  AO22X1_HVT U2652 ( .A1(\ram[14][54] ), .A2(n5374), .A3(n5375), .A4(data[54]), 
        .Y(n3699) );
  AO22X1_HVT U2653 ( .A1(\ram[14][53] ), .A2(n5374), .A3(n5375), .A4(data[53]), 
        .Y(n3698) );
  AO22X1_HVT U2654 ( .A1(\ram[14][52] ), .A2(n5374), .A3(n5375), .A4(data[52]), 
        .Y(n3697) );
  AO22X1_HVT U2655 ( .A1(\ram[14][51] ), .A2(n5374), .A3(n5375), .A4(data[51]), 
        .Y(n3696) );
  AO22X1_HVT U2656 ( .A1(\ram[14][50] ), .A2(n5374), .A3(n5375), .A4(data[50]), 
        .Y(n3695) );
  AO22X1_HVT U2657 ( .A1(\ram[14][49] ), .A2(n5374), .A3(n5375), .A4(data[49]), 
        .Y(n3694) );
  AO22X1_HVT U2658 ( .A1(\ram[14][48] ), .A2(n5374), .A3(n5375), .A4(data[48]), 
        .Y(n3693) );
  AO22X1_HVT U2659 ( .A1(\ram[14][47] ), .A2(n5374), .A3(n5375), .A4(data[47]), 
        .Y(n3692) );
  AO22X1_HVT U2660 ( .A1(\ram[14][46] ), .A2(n5374), .A3(n5375), .A4(data[46]), 
        .Y(n3691) );
  AO22X1_HVT U2661 ( .A1(\ram[14][45] ), .A2(n5374), .A3(n5375), .A4(data[45]), 
        .Y(n3690) );
  AO22X1_HVT U2662 ( .A1(\ram[1][52] ), .A2(n5368), .A3(n5369), .A4(data[52]), 
        .Y(n369) );
  AO22X1_HVT U2663 ( .A1(\ram[14][44] ), .A2(n5374), .A3(n5375), .A4(data[44]), 
        .Y(n3689) );
  AO22X1_HVT U2664 ( .A1(\ram[14][43] ), .A2(n5374), .A3(n5375), .A4(data[43]), 
        .Y(n3688) );
  AO22X1_HVT U2665 ( .A1(\ram[14][42] ), .A2(n5374), .A3(n5375), .A4(data[42]), 
        .Y(n3687) );
  AO22X1_HVT U2666 ( .A1(\ram[14][41] ), .A2(n5374), .A3(n5375), .A4(data[41]), 
        .Y(n3686) );
  AO22X1_HVT U2667 ( .A1(\ram[14][40] ), .A2(n5374), .A3(n5375), .A4(data[40]), 
        .Y(n3685) );
  AO22X1_HVT U2668 ( .A1(\ram[14][39] ), .A2(n5374), .A3(n5375), .A4(data[39]), 
        .Y(n3684) );
  AO22X1_HVT U2669 ( .A1(\ram[14][38] ), .A2(n5374), .A3(n5375), .A4(data[38]), 
        .Y(n3683) );
  AO22X1_HVT U2670 ( .A1(\ram[14][37] ), .A2(n5374), .A3(n5375), .A4(data[37]), 
        .Y(n3682) );
  AO22X1_HVT U2671 ( .A1(\ram[14][36] ), .A2(n5374), .A3(n5375), .A4(data[36]), 
        .Y(n3681) );
  AO22X1_HVT U2672 ( .A1(\ram[14][35] ), .A2(n5374), .A3(n5375), .A4(data[35]), 
        .Y(n3680) );
  AO22X1_HVT U2673 ( .A1(\ram[1][51] ), .A2(n5368), .A3(n5369), .A4(data[51]), 
        .Y(n368) );
  AO22X1_HVT U2674 ( .A1(\ram[14][34] ), .A2(n5374), .A3(n5375), .A4(data[34]), 
        .Y(n3679) );
  AO22X1_HVT U2675 ( .A1(\ram[14][33] ), .A2(n5374), .A3(n5375), .A4(data[33]), 
        .Y(n3678) );
  AO22X1_HVT U2676 ( .A1(\ram[14][32] ), .A2(n5374), .A3(n5375), .A4(data[32]), 
        .Y(n3677) );
  AO22X1_HVT U2677 ( .A1(\ram[14][31] ), .A2(n5374), .A3(n5375), .A4(data[31]), 
        .Y(n3676) );
  AO22X1_HVT U2678 ( .A1(\ram[14][30] ), .A2(n5374), .A3(n5375), .A4(data[30]), 
        .Y(n3675) );
  AO22X1_HVT U2679 ( .A1(\ram[14][29] ), .A2(n5374), .A3(n5375), .A4(data[29]), 
        .Y(n3674) );
  AO22X1_HVT U2680 ( .A1(\ram[14][28] ), .A2(n5374), .A3(n5375), .A4(data[28]), 
        .Y(n3673) );
  AO22X1_HVT U2681 ( .A1(\ram[14][27] ), .A2(n5374), .A3(n5375), .A4(data[27]), 
        .Y(n3672) );
  AO22X1_HVT U2682 ( .A1(\ram[14][26] ), .A2(n5374), .A3(n5375), .A4(data[26]), 
        .Y(n3671) );
  AO22X1_HVT U2683 ( .A1(\ram[14][25] ), .A2(n5374), .A3(n5375), .A4(data[25]), 
        .Y(n3670) );
  AO22X1_HVT U2684 ( .A1(\ram[1][50] ), .A2(n5368), .A3(n5369), .A4(data[50]), 
        .Y(n367) );
  AO22X1_HVT U2685 ( .A1(\ram[14][24] ), .A2(n5374), .A3(n5375), .A4(data[24]), 
        .Y(n3669) );
  AO22X1_HVT U2686 ( .A1(\ram[14][23] ), .A2(n5374), .A3(n5375), .A4(data[23]), 
        .Y(n3668) );
  AO22X1_HVT U2687 ( .A1(\ram[14][22] ), .A2(n5374), .A3(n5375), .A4(data[22]), 
        .Y(n3667) );
  AO22X1_HVT U2688 ( .A1(\ram[14][21] ), .A2(n5374), .A3(n5375), .A4(data[21]), 
        .Y(n3666) );
  AO22X1_HVT U2689 ( .A1(\ram[14][20] ), .A2(n5374), .A3(n5375), .A4(data[20]), 
        .Y(n3665) );
  AO22X1_HVT U2690 ( .A1(\ram[14][19] ), .A2(n5374), .A3(n5375), .A4(data[19]), 
        .Y(n3664) );
  AO22X1_HVT U2691 ( .A1(\ram[14][18] ), .A2(n5374), .A3(n5375), .A4(data[18]), 
        .Y(n3663) );
  AO22X1_HVT U2692 ( .A1(\ram[14][17] ), .A2(n5374), .A3(n5375), .A4(data[17]), 
        .Y(n3662) );
  AO22X1_HVT U2693 ( .A1(\ram[14][16] ), .A2(n5374), .A3(n5375), .A4(data[16]), 
        .Y(n3661) );
  AO22X1_HVT U2694 ( .A1(\ram[14][15] ), .A2(n5374), .A3(n5375), .A4(data[15]), 
        .Y(n3660) );
  AO22X1_HVT U2695 ( .A1(\ram[1][49] ), .A2(n5368), .A3(n5369), .A4(data[49]), 
        .Y(n366) );
  AO22X1_HVT U2696 ( .A1(\ram[14][14] ), .A2(n5374), .A3(n5375), .A4(data[14]), 
        .Y(n3659) );
  AO22X1_HVT U2697 ( .A1(\ram[14][13] ), .A2(n5374), .A3(n5375), .A4(data[13]), 
        .Y(n3658) );
  AO22X1_HVT U2698 ( .A1(\ram[14][12] ), .A2(n5374), .A3(n5375), .A4(data[12]), 
        .Y(n3657) );
  AO22X1_HVT U2699 ( .A1(\ram[14][11] ), .A2(n5374), .A3(n5375), .A4(data[11]), 
        .Y(n3656) );
  AO22X1_HVT U2700 ( .A1(\ram[14][10] ), .A2(n5374), .A3(n5375), .A4(data[10]), 
        .Y(n3655) );
  AO22X1_HVT U2701 ( .A1(\ram[14][9] ), .A2(n5374), .A3(n5375), .A4(data[9]), 
        .Y(n3654) );
  AO22X1_HVT U2702 ( .A1(\ram[14][8] ), .A2(n5374), .A3(n5375), .A4(data[8]), 
        .Y(n3653) );
  AO22X1_HVT U2703 ( .A1(\ram[14][7] ), .A2(n5374), .A3(n5375), .A4(data[7]), 
        .Y(n3652) );
  AO22X1_HVT U2704 ( .A1(\ram[14][6] ), .A2(n5374), .A3(n5375), .A4(data[6]), 
        .Y(n3651) );
  AO22X1_HVT U2705 ( .A1(\ram[14][5] ), .A2(n5374), .A3(n5375), .A4(data[5]), 
        .Y(n3650) );
  AO22X1_HVT U2706 ( .A1(\ram[1][48] ), .A2(n5368), .A3(n5369), .A4(data[48]), 
        .Y(n365) );
  AO22X1_HVT U2707 ( .A1(\ram[14][4] ), .A2(n5374), .A3(n5375), .A4(data[4]), 
        .Y(n3649) );
  AO22X1_HVT U2708 ( .A1(\ram[14][3] ), .A2(n5374), .A3(n5375), .A4(data[3]), 
        .Y(n3648) );
  AO22X1_HVT U2709 ( .A1(\ram[14][2] ), .A2(n5374), .A3(n5375), .A4(data[2]), 
        .Y(n3647) );
  AO22X1_HVT U2710 ( .A1(\ram[14][1] ), .A2(n5374), .A3(n5375), .A4(data[1]), 
        .Y(n3646) );
  AO22X1_HVT U2711 ( .A1(\ram[14][0] ), .A2(n5374), .A3(n5375), .A4(data[0]), 
        .Y(n3645) );
  INVX0_HVT U2712 ( .A(n5376), .Y(n5375) );
  AND2X1_HVT U2713 ( .A1(n5376), .A2(n5365), .Y(n5374) );
  NAND3X0_HVT U2714 ( .A1(n4276), .A2(n4183), .A3(n5373), .Y(n5376) );
  AO22X1_HVT U2715 ( .A1(\ram[13][255] ), .A2(n5377), .A3(n5378), .A4(
        data[255]), .Y(n3644) );
  AO22X1_HVT U2716 ( .A1(\ram[13][254] ), .A2(n5377), .A3(n5378), .A4(
        data[254]), .Y(n3643) );
  AO22X1_HVT U2717 ( .A1(\ram[13][253] ), .A2(n5377), .A3(n5378), .A4(
        data[253]), .Y(n3642) );
  AO22X1_HVT U2718 ( .A1(\ram[13][252] ), .A2(n5377), .A3(n5378), .A4(
        data[252]), .Y(n3641) );
  AO22X1_HVT U2719 ( .A1(\ram[13][251] ), .A2(n5377), .A3(n5378), .A4(
        data[251]), .Y(n3640) );
  AO22X1_HVT U2720 ( .A1(\ram[1][47] ), .A2(n5368), .A3(n5369), .A4(data[47]), 
        .Y(n364) );
  AO22X1_HVT U2721 ( .A1(\ram[13][250] ), .A2(n5377), .A3(n5378), .A4(
        data[250]), .Y(n3639) );
  AO22X1_HVT U2722 ( .A1(\ram[13][249] ), .A2(n5377), .A3(n5378), .A4(
        data[249]), .Y(n3638) );
  AO22X1_HVT U2723 ( .A1(\ram[13][248] ), .A2(n5377), .A3(n5378), .A4(
        data[248]), .Y(n3637) );
  AO22X1_HVT U2724 ( .A1(\ram[13][247] ), .A2(n5377), .A3(n5378), .A4(
        data[247]), .Y(n3636) );
  AO22X1_HVT U2725 ( .A1(\ram[13][246] ), .A2(n5377), .A3(n5378), .A4(
        data[246]), .Y(n3635) );
  AO22X1_HVT U2726 ( .A1(\ram[13][245] ), .A2(n5377), .A3(n5378), .A4(
        data[245]), .Y(n3634) );
  AO22X1_HVT U2727 ( .A1(\ram[13][244] ), .A2(n5377), .A3(n5378), .A4(
        data[244]), .Y(n3633) );
  AO22X1_HVT U2728 ( .A1(\ram[13][243] ), .A2(n5377), .A3(n5378), .A4(
        data[243]), .Y(n3632) );
  AO22X1_HVT U2729 ( .A1(\ram[13][242] ), .A2(n5377), .A3(n5378), .A4(
        data[242]), .Y(n3631) );
  AO22X1_HVT U2730 ( .A1(\ram[13][241] ), .A2(n5377), .A3(n5378), .A4(
        data[241]), .Y(n3630) );
  AO22X1_HVT U2731 ( .A1(\ram[1][46] ), .A2(n5368), .A3(n5369), .A4(data[46]), 
        .Y(n363) );
  AO22X1_HVT U2732 ( .A1(\ram[13][240] ), .A2(n5377), .A3(n5378), .A4(
        data[240]), .Y(n3629) );
  AO22X1_HVT U2733 ( .A1(\ram[13][239] ), .A2(n5377), .A3(n5378), .A4(
        data[239]), .Y(n3628) );
  AO22X1_HVT U2734 ( .A1(\ram[13][238] ), .A2(n5377), .A3(n5378), .A4(
        data[238]), .Y(n3627) );
  AO22X1_HVT U2735 ( .A1(\ram[13][237] ), .A2(n5377), .A3(n5378), .A4(
        data[237]), .Y(n3626) );
  AO22X1_HVT U2736 ( .A1(\ram[13][236] ), .A2(n5377), .A3(n5378), .A4(
        data[236]), .Y(n3625) );
  AO22X1_HVT U2737 ( .A1(\ram[13][235] ), .A2(n5377), .A3(n5378), .A4(
        data[235]), .Y(n3624) );
  AO22X1_HVT U2738 ( .A1(\ram[13][234] ), .A2(n5377), .A3(n5378), .A4(
        data[234]), .Y(n3623) );
  AO22X1_HVT U2739 ( .A1(\ram[13][233] ), .A2(n5377), .A3(n5378), .A4(
        data[233]), .Y(n3622) );
  AO22X1_HVT U2740 ( .A1(\ram[13][232] ), .A2(n5377), .A3(n5378), .A4(
        data[232]), .Y(n3621) );
  AO22X1_HVT U2741 ( .A1(\ram[13][231] ), .A2(n5377), .A3(n5378), .A4(
        data[231]), .Y(n3620) );
  AO22X1_HVT U2742 ( .A1(\ram[1][45] ), .A2(n5368), .A3(n5369), .A4(data[45]), 
        .Y(n362) );
  AO22X1_HVT U2743 ( .A1(\ram[13][230] ), .A2(n5377), .A3(n5378), .A4(
        data[230]), .Y(n3619) );
  AO22X1_HVT U2744 ( .A1(\ram[13][229] ), .A2(n5377), .A3(n5378), .A4(
        data[229]), .Y(n3618) );
  AO22X1_HVT U2745 ( .A1(\ram[13][228] ), .A2(n5377), .A3(n5378), .A4(
        data[228]), .Y(n3617) );
  AO22X1_HVT U2746 ( .A1(\ram[13][227] ), .A2(n5377), .A3(n5378), .A4(
        data[227]), .Y(n3616) );
  AO22X1_HVT U2747 ( .A1(\ram[13][226] ), .A2(n5377), .A3(n5378), .A4(
        data[226]), .Y(n3615) );
  AO22X1_HVT U2748 ( .A1(\ram[13][225] ), .A2(n5377), .A3(n5378), .A4(
        data[225]), .Y(n3614) );
  AO22X1_HVT U2749 ( .A1(\ram[13][224] ), .A2(n5377), .A3(n5378), .A4(
        data[224]), .Y(n3613) );
  AO22X1_HVT U2750 ( .A1(\ram[13][223] ), .A2(n5377), .A3(n5378), .A4(
        data[223]), .Y(n3612) );
  AO22X1_HVT U2751 ( .A1(\ram[13][222] ), .A2(n5377), .A3(n5378), .A4(
        data[222]), .Y(n3611) );
  AO22X1_HVT U2752 ( .A1(\ram[13][221] ), .A2(n5377), .A3(n5378), .A4(
        data[221]), .Y(n3610) );
  AO22X1_HVT U2753 ( .A1(\ram[1][44] ), .A2(n5368), .A3(n5369), .A4(data[44]), 
        .Y(n361) );
  AO22X1_HVT U2754 ( .A1(\ram[13][220] ), .A2(n5377), .A3(n5378), .A4(
        data[220]), .Y(n3609) );
  AO22X1_HVT U2755 ( .A1(\ram[13][219] ), .A2(n5377), .A3(n5378), .A4(
        data[219]), .Y(n3608) );
  AO22X1_HVT U2756 ( .A1(\ram[13][218] ), .A2(n5377), .A3(n5378), .A4(
        data[218]), .Y(n3607) );
  AO22X1_HVT U2757 ( .A1(\ram[13][217] ), .A2(n5377), .A3(n5378), .A4(
        data[217]), .Y(n3606) );
  AO22X1_HVT U2758 ( .A1(\ram[13][216] ), .A2(n5377), .A3(n5378), .A4(
        data[216]), .Y(n3605) );
  AO22X1_HVT U2759 ( .A1(\ram[13][215] ), .A2(n5377), .A3(n5378), .A4(
        data[215]), .Y(n3604) );
  AO22X1_HVT U2760 ( .A1(\ram[13][214] ), .A2(n5377), .A3(n5378), .A4(
        data[214]), .Y(n3603) );
  AO22X1_HVT U2761 ( .A1(\ram[13][213] ), .A2(n5377), .A3(n5378), .A4(
        data[213]), .Y(n3602) );
  AO22X1_HVT U2762 ( .A1(\ram[13][212] ), .A2(n5377), .A3(n5378), .A4(
        data[212]), .Y(n3601) );
  AO22X1_HVT U2763 ( .A1(\ram[13][211] ), .A2(n5377), .A3(n5378), .A4(
        data[211]), .Y(n3600) );
  AO22X1_HVT U2764 ( .A1(\ram[1][43] ), .A2(n5368), .A3(n5369), .A4(data[43]), 
        .Y(n360) );
  AO22X1_HVT U2765 ( .A1(\ram[13][210] ), .A2(n5377), .A3(n5378), .A4(
        data[210]), .Y(n3599) );
  AO22X1_HVT U2766 ( .A1(\ram[13][209] ), .A2(n5377), .A3(n5378), .A4(
        data[209]), .Y(n3598) );
  AO22X1_HVT U2767 ( .A1(\ram[13][208] ), .A2(n5377), .A3(n5378), .A4(
        data[208]), .Y(n3597) );
  AO22X1_HVT U2768 ( .A1(\ram[13][207] ), .A2(n5377), .A3(n5378), .A4(
        data[207]), .Y(n3596) );
  AO22X1_HVT U2769 ( .A1(\ram[13][206] ), .A2(n5377), .A3(n5378), .A4(
        data[206]), .Y(n3595) );
  AO22X1_HVT U2770 ( .A1(\ram[13][205] ), .A2(n5377), .A3(n5378), .A4(
        data[205]), .Y(n3594) );
  AO22X1_HVT U2771 ( .A1(\ram[13][204] ), .A2(n5377), .A3(n5378), .A4(
        data[204]), .Y(n3593) );
  AO22X1_HVT U2772 ( .A1(\ram[13][203] ), .A2(n5377), .A3(n5378), .A4(
        data[203]), .Y(n3592) );
  AO22X1_HVT U2773 ( .A1(\ram[13][202] ), .A2(n5377), .A3(n5378), .A4(
        data[202]), .Y(n3591) );
  AO22X1_HVT U2774 ( .A1(\ram[13][201] ), .A2(n5377), .A3(n5378), .A4(
        data[201]), .Y(n3590) );
  AO22X1_HVT U2775 ( .A1(\ram[1][42] ), .A2(n5368), .A3(n5369), .A4(data[42]), 
        .Y(n359) );
  AO22X1_HVT U2776 ( .A1(\ram[13][200] ), .A2(n5377), .A3(n5378), .A4(
        data[200]), .Y(n3589) );
  AO22X1_HVT U2777 ( .A1(\ram[13][199] ), .A2(n5377), .A3(n5378), .A4(
        data[199]), .Y(n3588) );
  AO22X1_HVT U2778 ( .A1(\ram[13][198] ), .A2(n5377), .A3(n5378), .A4(
        data[198]), .Y(n3587) );
  AO22X1_HVT U2779 ( .A1(\ram[13][197] ), .A2(n5377), .A3(n5378), .A4(
        data[197]), .Y(n3586) );
  AO22X1_HVT U2780 ( .A1(\ram[13][196] ), .A2(n5377), .A3(n5378), .A4(
        data[196]), .Y(n3585) );
  AO22X1_HVT U2781 ( .A1(\ram[13][195] ), .A2(n5377), .A3(n5378), .A4(
        data[195]), .Y(n3584) );
  AO22X1_HVT U2782 ( .A1(\ram[13][194] ), .A2(n5377), .A3(n5378), .A4(
        data[194]), .Y(n3583) );
  AO22X1_HVT U2783 ( .A1(\ram[13][193] ), .A2(n5377), .A3(n5378), .A4(
        data[193]), .Y(n3582) );
  AO22X1_HVT U2784 ( .A1(\ram[13][192] ), .A2(n5377), .A3(n5378), .A4(
        data[192]), .Y(n3581) );
  AO22X1_HVT U2785 ( .A1(\ram[13][191] ), .A2(n5377), .A3(n5378), .A4(
        data[191]), .Y(n3580) );
  AO22X1_HVT U2786 ( .A1(\ram[1][41] ), .A2(n5368), .A3(n5369), .A4(data[41]), 
        .Y(n358) );
  AO22X1_HVT U2787 ( .A1(\ram[13][190] ), .A2(n5377), .A3(n5378), .A4(
        data[190]), .Y(n3579) );
  AO22X1_HVT U2788 ( .A1(\ram[13][189] ), .A2(n5377), .A3(n5378), .A4(
        data[189]), .Y(n3578) );
  AO22X1_HVT U2789 ( .A1(\ram[13][188] ), .A2(n5377), .A3(n5378), .A4(
        data[188]), .Y(n3577) );
  AO22X1_HVT U2790 ( .A1(\ram[13][187] ), .A2(n5377), .A3(n5378), .A4(
        data[187]), .Y(n3576) );
  AO22X1_HVT U2791 ( .A1(\ram[13][186] ), .A2(n5377), .A3(n5378), .A4(
        data[186]), .Y(n3575) );
  AO22X1_HVT U2792 ( .A1(\ram[13][185] ), .A2(n5377), .A3(n5378), .A4(
        data[185]), .Y(n3574) );
  AO22X1_HVT U2793 ( .A1(\ram[13][184] ), .A2(n5377), .A3(n5378), .A4(
        data[184]), .Y(n3573) );
  AO22X1_HVT U2794 ( .A1(\ram[13][183] ), .A2(n5377), .A3(n5378), .A4(
        data[183]), .Y(n3572) );
  AO22X1_HVT U2795 ( .A1(\ram[13][182] ), .A2(n5377), .A3(n5378), .A4(
        data[182]), .Y(n3571) );
  AO22X1_HVT U2796 ( .A1(\ram[13][181] ), .A2(n5377), .A3(n5378), .A4(
        data[181]), .Y(n3570) );
  AO22X1_HVT U2797 ( .A1(\ram[1][40] ), .A2(n5368), .A3(n5369), .A4(data[40]), 
        .Y(n357) );
  AO22X1_HVT U2798 ( .A1(\ram[13][180] ), .A2(n5377), .A3(n5378), .A4(
        data[180]), .Y(n3569) );
  AO22X1_HVT U2799 ( .A1(\ram[13][179] ), .A2(n5377), .A3(n5378), .A4(
        data[179]), .Y(n3568) );
  AO22X1_HVT U2800 ( .A1(\ram[13][178] ), .A2(n5377), .A3(n5378), .A4(
        data[178]), .Y(n3567) );
  AO22X1_HVT U2801 ( .A1(\ram[13][177] ), .A2(n5377), .A3(n5378), .A4(
        data[177]), .Y(n3566) );
  AO22X1_HVT U2802 ( .A1(\ram[13][176] ), .A2(n5377), .A3(n5378), .A4(
        data[176]), .Y(n3565) );
  AO22X1_HVT U2803 ( .A1(\ram[13][175] ), .A2(n5377), .A3(n5378), .A4(
        data[175]), .Y(n3564) );
  AO22X1_HVT U2804 ( .A1(\ram[13][174] ), .A2(n5377), .A3(n5378), .A4(
        data[174]), .Y(n3563) );
  AO22X1_HVT U2805 ( .A1(\ram[13][173] ), .A2(n5377), .A3(n5378), .A4(
        data[173]), .Y(n3562) );
  AO22X1_HVT U2806 ( .A1(\ram[13][172] ), .A2(n5377), .A3(n5378), .A4(
        data[172]), .Y(n3561) );
  AO22X1_HVT U2807 ( .A1(\ram[13][171] ), .A2(n5377), .A3(n5378), .A4(
        data[171]), .Y(n3560) );
  AO22X1_HVT U2808 ( .A1(\ram[1][39] ), .A2(n5368), .A3(n5369), .A4(data[39]), 
        .Y(n356) );
  AO22X1_HVT U2809 ( .A1(\ram[13][170] ), .A2(n5377), .A3(n5378), .A4(
        data[170]), .Y(n3559) );
  AO22X1_HVT U2810 ( .A1(\ram[13][169] ), .A2(n5377), .A3(n5378), .A4(
        data[169]), .Y(n3558) );
  AO22X1_HVT U2811 ( .A1(\ram[13][168] ), .A2(n5377), .A3(n5378), .A4(
        data[168]), .Y(n3557) );
  AO22X1_HVT U2812 ( .A1(\ram[13][167] ), .A2(n5377), .A3(n5378), .A4(
        data[167]), .Y(n3556) );
  AO22X1_HVT U2813 ( .A1(\ram[13][166] ), .A2(n5377), .A3(n5378), .A4(
        data[166]), .Y(n3555) );
  AO22X1_HVT U2814 ( .A1(\ram[13][165] ), .A2(n5377), .A3(n5378), .A4(
        data[165]), .Y(n3554) );
  AO22X1_HVT U2815 ( .A1(\ram[13][164] ), .A2(n5377), .A3(n5378), .A4(
        data[164]), .Y(n3553) );
  AO22X1_HVT U2816 ( .A1(\ram[13][163] ), .A2(n5377), .A3(n5378), .A4(
        data[163]), .Y(n3552) );
  AO22X1_HVT U2817 ( .A1(\ram[13][162] ), .A2(n5377), .A3(n5378), .A4(
        data[162]), .Y(n3551) );
  AO22X1_HVT U2818 ( .A1(\ram[13][161] ), .A2(n5377), .A3(n5378), .A4(
        data[161]), .Y(n3550) );
  AO22X1_HVT U2819 ( .A1(\ram[1][38] ), .A2(n5368), .A3(n5369), .A4(data[38]), 
        .Y(n355) );
  AO22X1_HVT U2820 ( .A1(\ram[13][160] ), .A2(n5377), .A3(n5378), .A4(
        data[160]), .Y(n3549) );
  AO22X1_HVT U2821 ( .A1(\ram[13][159] ), .A2(n5377), .A3(n5378), .A4(
        data[159]), .Y(n3548) );
  AO22X1_HVT U2822 ( .A1(\ram[13][158] ), .A2(n5377), .A3(n5378), .A4(
        data[158]), .Y(n3547) );
  AO22X1_HVT U2823 ( .A1(\ram[13][157] ), .A2(n5377), .A3(n5378), .A4(
        data[157]), .Y(n3546) );
  AO22X1_HVT U2824 ( .A1(\ram[13][156] ), .A2(n5377), .A3(n5378), .A4(
        data[156]), .Y(n3545) );
  AO22X1_HVT U2825 ( .A1(\ram[13][155] ), .A2(n5377), .A3(n5378), .A4(
        data[155]), .Y(n3544) );
  AO22X1_HVT U2826 ( .A1(\ram[13][154] ), .A2(n5377), .A3(n5378), .A4(
        data[154]), .Y(n3543) );
  AO22X1_HVT U2827 ( .A1(\ram[13][153] ), .A2(n5377), .A3(n5378), .A4(
        data[153]), .Y(n3542) );
  AO22X1_HVT U2828 ( .A1(\ram[13][152] ), .A2(n5377), .A3(n5378), .A4(
        data[152]), .Y(n3541) );
  AO22X1_HVT U2829 ( .A1(\ram[13][151] ), .A2(n5377), .A3(n5378), .A4(
        data[151]), .Y(n3540) );
  AO22X1_HVT U2830 ( .A1(\ram[1][37] ), .A2(n5368), .A3(n5369), .A4(data[37]), 
        .Y(n354) );
  AO22X1_HVT U2831 ( .A1(\ram[13][150] ), .A2(n5377), .A3(n5378), .A4(
        data[150]), .Y(n3539) );
  AO22X1_HVT U2832 ( .A1(\ram[13][149] ), .A2(n5377), .A3(n5378), .A4(
        data[149]), .Y(n3538) );
  AO22X1_HVT U2833 ( .A1(\ram[13][148] ), .A2(n5377), .A3(n5378), .A4(
        data[148]), .Y(n3537) );
  AO22X1_HVT U2834 ( .A1(\ram[13][147] ), .A2(n5377), .A3(n5378), .A4(
        data[147]), .Y(n3536) );
  AO22X1_HVT U2835 ( .A1(\ram[13][146] ), .A2(n5377), .A3(n5378), .A4(
        data[146]), .Y(n3535) );
  AO22X1_HVT U2836 ( .A1(\ram[13][145] ), .A2(n5377), .A3(n5378), .A4(
        data[145]), .Y(n3534) );
  AO22X1_HVT U2837 ( .A1(\ram[13][144] ), .A2(n5377), .A3(n5378), .A4(
        data[144]), .Y(n3533) );
  AO22X1_HVT U2838 ( .A1(\ram[13][143] ), .A2(n5377), .A3(n5378), .A4(
        data[143]), .Y(n3532) );
  AO22X1_HVT U2839 ( .A1(\ram[13][142] ), .A2(n5377), .A3(n5378), .A4(
        data[142]), .Y(n3531) );
  AO22X1_HVT U2840 ( .A1(\ram[13][141] ), .A2(n5377), .A3(n5378), .A4(
        data[141]), .Y(n3530) );
  AO22X1_HVT U2841 ( .A1(\ram[1][36] ), .A2(n5368), .A3(n5369), .A4(data[36]), 
        .Y(n353) );
  AO22X1_HVT U2842 ( .A1(\ram[13][140] ), .A2(n5377), .A3(n5378), .A4(
        data[140]), .Y(n3529) );
  AO22X1_HVT U2843 ( .A1(\ram[13][139] ), .A2(n5377), .A3(n5378), .A4(
        data[139]), .Y(n3528) );
  AO22X1_HVT U2844 ( .A1(\ram[13][138] ), .A2(n5377), .A3(n5378), .A4(
        data[138]), .Y(n3527) );
  AO22X1_HVT U2845 ( .A1(\ram[13][137] ), .A2(n5377), .A3(n5378), .A4(
        data[137]), .Y(n3526) );
  AO22X1_HVT U2846 ( .A1(\ram[13][136] ), .A2(n5377), .A3(n5378), .A4(
        data[136]), .Y(n3525) );
  AO22X1_HVT U2847 ( .A1(\ram[13][135] ), .A2(n5377), .A3(n5378), .A4(
        data[135]), .Y(n3524) );
  AO22X1_HVT U2848 ( .A1(\ram[13][134] ), .A2(n5377), .A3(n5378), .A4(
        data[134]), .Y(n3523) );
  AO22X1_HVT U2849 ( .A1(\ram[13][133] ), .A2(n5377), .A3(n5378), .A4(
        data[133]), .Y(n3522) );
  AO22X1_HVT U2850 ( .A1(\ram[13][132] ), .A2(n5377), .A3(n5378), .A4(
        data[132]), .Y(n3521) );
  AO22X1_HVT U2851 ( .A1(\ram[13][131] ), .A2(n5377), .A3(n5378), .A4(
        data[131]), .Y(n3520) );
  AO22X1_HVT U2852 ( .A1(\ram[1][35] ), .A2(n5368), .A3(n5369), .A4(data[35]), 
        .Y(n352) );
  AO22X1_HVT U2853 ( .A1(\ram[13][130] ), .A2(n5377), .A3(n5378), .A4(
        data[130]), .Y(n3519) );
  AO22X1_HVT U2854 ( .A1(\ram[13][129] ), .A2(n5377), .A3(n5378), .A4(
        data[129]), .Y(n3518) );
  AO22X1_HVT U2855 ( .A1(\ram[13][128] ), .A2(n5377), .A3(n5378), .A4(
        data[128]), .Y(n3517) );
  AO22X1_HVT U2856 ( .A1(\ram[13][127] ), .A2(n5377), .A3(n5378), .A4(
        data[127]), .Y(n3516) );
  AO22X1_HVT U2857 ( .A1(\ram[13][126] ), .A2(n5377), .A3(n5378), .A4(
        data[126]), .Y(n3515) );
  AO22X1_HVT U2858 ( .A1(\ram[13][125] ), .A2(n5377), .A3(n5378), .A4(
        data[125]), .Y(n3514) );
  AO22X1_HVT U2859 ( .A1(\ram[13][124] ), .A2(n5377), .A3(n5378), .A4(
        data[124]), .Y(n3513) );
  AO22X1_HVT U2860 ( .A1(\ram[13][123] ), .A2(n5377), .A3(n5378), .A4(
        data[123]), .Y(n3512) );
  AO22X1_HVT U2861 ( .A1(\ram[13][122] ), .A2(n5377), .A3(n5378), .A4(
        data[122]), .Y(n3511) );
  AO22X1_HVT U2862 ( .A1(\ram[13][121] ), .A2(n5377), .A3(n5378), .A4(
        data[121]), .Y(n3510) );
  AO22X1_HVT U2863 ( .A1(\ram[1][34] ), .A2(n5368), .A3(n5369), .A4(data[34]), 
        .Y(n351) );
  AO22X1_HVT U2864 ( .A1(\ram[13][120] ), .A2(n5377), .A3(n5378), .A4(
        data[120]), .Y(n3509) );
  AO22X1_HVT U2865 ( .A1(\ram[13][119] ), .A2(n5377), .A3(n5378), .A4(
        data[119]), .Y(n3508) );
  AO22X1_HVT U2866 ( .A1(\ram[13][118] ), .A2(n5377), .A3(n5378), .A4(
        data[118]), .Y(n3507) );
  AO22X1_HVT U2867 ( .A1(\ram[13][117] ), .A2(n5377), .A3(n5378), .A4(
        data[117]), .Y(n3506) );
  AO22X1_HVT U2868 ( .A1(\ram[13][116] ), .A2(n5377), .A3(n5378), .A4(
        data[116]), .Y(n3505) );
  AO22X1_HVT U2869 ( .A1(\ram[13][115] ), .A2(n5377), .A3(n5378), .A4(
        data[115]), .Y(n3504) );
  AO22X1_HVT U2870 ( .A1(\ram[13][114] ), .A2(n5377), .A3(n5378), .A4(
        data[114]), .Y(n3503) );
  AO22X1_HVT U2871 ( .A1(\ram[13][113] ), .A2(n5377), .A3(n5378), .A4(
        data[113]), .Y(n3502) );
  AO22X1_HVT U2872 ( .A1(\ram[13][112] ), .A2(n5377), .A3(n5378), .A4(
        data[112]), .Y(n3501) );
  AO22X1_HVT U2873 ( .A1(\ram[13][111] ), .A2(n5377), .A3(n5378), .A4(
        data[111]), .Y(n3500) );
  AO22X1_HVT U2874 ( .A1(\ram[1][33] ), .A2(n5368), .A3(n5369), .A4(data[33]), 
        .Y(n350) );
  AO22X1_HVT U2875 ( .A1(\ram[13][110] ), .A2(n5377), .A3(n5378), .A4(
        data[110]), .Y(n3499) );
  AO22X1_HVT U2876 ( .A1(\ram[13][109] ), .A2(n5377), .A3(n5378), .A4(
        data[109]), .Y(n3498) );
  AO22X1_HVT U2877 ( .A1(\ram[13][108] ), .A2(n5377), .A3(n5378), .A4(
        data[108]), .Y(n3497) );
  AO22X1_HVT U2878 ( .A1(\ram[13][107] ), .A2(n5377), .A3(n5378), .A4(
        data[107]), .Y(n3496) );
  AO22X1_HVT U2879 ( .A1(\ram[13][106] ), .A2(n5377), .A3(n5378), .A4(
        data[106]), .Y(n3495) );
  AO22X1_HVT U2880 ( .A1(\ram[13][105] ), .A2(n5377), .A3(n5378), .A4(
        data[105]), .Y(n3494) );
  AO22X1_HVT U2881 ( .A1(\ram[13][104] ), .A2(n5377), .A3(n5378), .A4(
        data[104]), .Y(n3493) );
  AO22X1_HVT U2882 ( .A1(\ram[13][103] ), .A2(n5377), .A3(n5378), .A4(
        data[103]), .Y(n3492) );
  AO22X1_HVT U2883 ( .A1(\ram[13][102] ), .A2(n5377), .A3(n5378), .A4(
        data[102]), .Y(n3491) );
  AO22X1_HVT U2884 ( .A1(\ram[13][101] ), .A2(n5377), .A3(n5378), .A4(
        data[101]), .Y(n3490) );
  AO22X1_HVT U2885 ( .A1(\ram[1][32] ), .A2(n5368), .A3(n5369), .A4(data[32]), 
        .Y(n349) );
  AO22X1_HVT U2886 ( .A1(\ram[13][100] ), .A2(n5377), .A3(n5378), .A4(
        data[100]), .Y(n3489) );
  AO22X1_HVT U2887 ( .A1(\ram[13][99] ), .A2(n5377), .A3(n5378), .A4(data[99]), 
        .Y(n3488) );
  AO22X1_HVT U2888 ( .A1(\ram[13][98] ), .A2(n5377), .A3(n5378), .A4(data[98]), 
        .Y(n3487) );
  AO22X1_HVT U2889 ( .A1(\ram[13][97] ), .A2(n5377), .A3(n5378), .A4(data[97]), 
        .Y(n3486) );
  AO22X1_HVT U2890 ( .A1(\ram[13][96] ), .A2(n5377), .A3(n5378), .A4(data[96]), 
        .Y(n3485) );
  AO22X1_HVT U2891 ( .A1(\ram[13][95] ), .A2(n5377), .A3(n5378), .A4(data[95]), 
        .Y(n3484) );
  AO22X1_HVT U2892 ( .A1(\ram[13][94] ), .A2(n5377), .A3(n5378), .A4(data[94]), 
        .Y(n3483) );
  AO22X1_HVT U2893 ( .A1(\ram[13][93] ), .A2(n5377), .A3(n5378), .A4(data[93]), 
        .Y(n3482) );
  AO22X1_HVT U2894 ( .A1(\ram[13][92] ), .A2(n5377), .A3(n5378), .A4(data[92]), 
        .Y(n3481) );
  AO22X1_HVT U2895 ( .A1(\ram[13][91] ), .A2(n5377), .A3(n5378), .A4(data[91]), 
        .Y(n3480) );
  AO22X1_HVT U2896 ( .A1(\ram[1][31] ), .A2(n5368), .A3(n5369), .A4(data[31]), 
        .Y(n348) );
  AO22X1_HVT U2897 ( .A1(\ram[13][90] ), .A2(n5377), .A3(n5378), .A4(data[90]), 
        .Y(n3479) );
  AO22X1_HVT U2898 ( .A1(\ram[13][89] ), .A2(n5377), .A3(n5378), .A4(data[89]), 
        .Y(n3478) );
  AO22X1_HVT U2899 ( .A1(\ram[13][88] ), .A2(n5377), .A3(n5378), .A4(data[88]), 
        .Y(n3477) );
  AO22X1_HVT U2900 ( .A1(\ram[13][87] ), .A2(n5377), .A3(n5378), .A4(data[87]), 
        .Y(n3476) );
  AO22X1_HVT U2901 ( .A1(\ram[13][86] ), .A2(n5377), .A3(n5378), .A4(data[86]), 
        .Y(n3475) );
  AO22X1_HVT U2902 ( .A1(\ram[13][85] ), .A2(n5377), .A3(n5378), .A4(data[85]), 
        .Y(n3474) );
  AO22X1_HVT U2903 ( .A1(\ram[13][84] ), .A2(n5377), .A3(n5378), .A4(data[84]), 
        .Y(n3473) );
  AO22X1_HVT U2904 ( .A1(\ram[13][83] ), .A2(n5377), .A3(n5378), .A4(data[83]), 
        .Y(n3472) );
  AO22X1_HVT U2905 ( .A1(\ram[13][82] ), .A2(n5377), .A3(n5378), .A4(data[82]), 
        .Y(n3471) );
  AO22X1_HVT U2906 ( .A1(\ram[13][81] ), .A2(n5377), .A3(n5378), .A4(data[81]), 
        .Y(n3470) );
  AO22X1_HVT U2907 ( .A1(\ram[1][30] ), .A2(n5368), .A3(n5369), .A4(data[30]), 
        .Y(n347) );
  AO22X1_HVT U2908 ( .A1(\ram[13][80] ), .A2(n5377), .A3(n5378), .A4(data[80]), 
        .Y(n3469) );
  AO22X1_HVT U2909 ( .A1(\ram[13][79] ), .A2(n5377), .A3(n5378), .A4(data[79]), 
        .Y(n3468) );
  AO22X1_HVT U2910 ( .A1(\ram[13][78] ), .A2(n5377), .A3(n5378), .A4(data[78]), 
        .Y(n3467) );
  AO22X1_HVT U2911 ( .A1(\ram[13][77] ), .A2(n5377), .A3(n5378), .A4(data[77]), 
        .Y(n3466) );
  AO22X1_HVT U2912 ( .A1(\ram[13][76] ), .A2(n5377), .A3(n5378), .A4(data[76]), 
        .Y(n3465) );
  AO22X1_HVT U2913 ( .A1(\ram[13][75] ), .A2(n5377), .A3(n5378), .A4(data[75]), 
        .Y(n3464) );
  AO22X1_HVT U2914 ( .A1(\ram[13][74] ), .A2(n5377), .A3(n5378), .A4(data[74]), 
        .Y(n3463) );
  AO22X1_HVT U2915 ( .A1(\ram[13][73] ), .A2(n5377), .A3(n5378), .A4(data[73]), 
        .Y(n3462) );
  AO22X1_HVT U2916 ( .A1(\ram[13][72] ), .A2(n5377), .A3(n5378), .A4(data[72]), 
        .Y(n3461) );
  AO22X1_HVT U2917 ( .A1(\ram[13][71] ), .A2(n5377), .A3(n5378), .A4(data[71]), 
        .Y(n3460) );
  AO22X1_HVT U2918 ( .A1(\ram[1][29] ), .A2(n5368), .A3(n5369), .A4(data[29]), 
        .Y(n346) );
  AO22X1_HVT U2919 ( .A1(\ram[13][70] ), .A2(n5377), .A3(n5378), .A4(data[70]), 
        .Y(n3459) );
  AO22X1_HVT U2920 ( .A1(\ram[13][69] ), .A2(n5377), .A3(n5378), .A4(data[69]), 
        .Y(n3458) );
  AO22X1_HVT U2921 ( .A1(\ram[13][68] ), .A2(n5377), .A3(n5378), .A4(data[68]), 
        .Y(n3457) );
  AO22X1_HVT U2922 ( .A1(\ram[13][67] ), .A2(n5377), .A3(n5378), .A4(data[67]), 
        .Y(n3456) );
  AO22X1_HVT U2923 ( .A1(\ram[13][66] ), .A2(n5377), .A3(n5378), .A4(data[66]), 
        .Y(n3455) );
  AO22X1_HVT U2924 ( .A1(\ram[13][65] ), .A2(n5377), .A3(n5378), .A4(data[65]), 
        .Y(n3454) );
  AO22X1_HVT U2925 ( .A1(\ram[13][64] ), .A2(n5377), .A3(n5378), .A4(data[64]), 
        .Y(n3453) );
  AO22X1_HVT U2926 ( .A1(\ram[13][63] ), .A2(n5377), .A3(n5378), .A4(data[63]), 
        .Y(n3452) );
  AO22X1_HVT U2927 ( .A1(\ram[13][62] ), .A2(n5377), .A3(n5378), .A4(data[62]), 
        .Y(n3451) );
  AO22X1_HVT U2928 ( .A1(\ram[13][61] ), .A2(n5377), .A3(n5378), .A4(data[61]), 
        .Y(n3450) );
  AO22X1_HVT U2929 ( .A1(\ram[1][28] ), .A2(n5368), .A3(n5369), .A4(data[28]), 
        .Y(n345) );
  AO22X1_HVT U2930 ( .A1(\ram[13][60] ), .A2(n5377), .A3(n5378), .A4(data[60]), 
        .Y(n3449) );
  AO22X1_HVT U2931 ( .A1(\ram[13][59] ), .A2(n5377), .A3(n5378), .A4(data[59]), 
        .Y(n3448) );
  AO22X1_HVT U2932 ( .A1(\ram[13][58] ), .A2(n5377), .A3(n5378), .A4(data[58]), 
        .Y(n3447) );
  AO22X1_HVT U2933 ( .A1(\ram[13][57] ), .A2(n5377), .A3(n5378), .A4(data[57]), 
        .Y(n3446) );
  AO22X1_HVT U2934 ( .A1(\ram[13][56] ), .A2(n5377), .A3(n5378), .A4(data[56]), 
        .Y(n3445) );
  AO22X1_HVT U2935 ( .A1(\ram[13][55] ), .A2(n5377), .A3(n5378), .A4(data[55]), 
        .Y(n3444) );
  AO22X1_HVT U2936 ( .A1(\ram[13][54] ), .A2(n5377), .A3(n5378), .A4(data[54]), 
        .Y(n3443) );
  AO22X1_HVT U2937 ( .A1(\ram[13][53] ), .A2(n5377), .A3(n5378), .A4(data[53]), 
        .Y(n3442) );
  AO22X1_HVT U2938 ( .A1(\ram[13][52] ), .A2(n5377), .A3(n5378), .A4(data[52]), 
        .Y(n3441) );
  AO22X1_HVT U2939 ( .A1(\ram[13][51] ), .A2(n5377), .A3(n5378), .A4(data[51]), 
        .Y(n3440) );
  AO22X1_HVT U2940 ( .A1(\ram[1][27] ), .A2(n5368), .A3(n5369), .A4(data[27]), 
        .Y(n344) );
  AO22X1_HVT U2941 ( .A1(\ram[13][50] ), .A2(n5377), .A3(n5378), .A4(data[50]), 
        .Y(n3439) );
  AO22X1_HVT U2942 ( .A1(\ram[13][49] ), .A2(n5377), .A3(n5378), .A4(data[49]), 
        .Y(n3438) );
  AO22X1_HVT U2943 ( .A1(\ram[13][48] ), .A2(n5377), .A3(n5378), .A4(data[48]), 
        .Y(n3437) );
  AO22X1_HVT U2944 ( .A1(\ram[13][47] ), .A2(n5377), .A3(n5378), .A4(data[47]), 
        .Y(n3436) );
  AO22X1_HVT U2945 ( .A1(\ram[13][46] ), .A2(n5377), .A3(n5378), .A4(data[46]), 
        .Y(n3435) );
  AO22X1_HVT U2946 ( .A1(\ram[13][45] ), .A2(n5377), .A3(n5378), .A4(data[45]), 
        .Y(n3434) );
  AO22X1_HVT U2947 ( .A1(\ram[13][44] ), .A2(n5377), .A3(n5378), .A4(data[44]), 
        .Y(n3433) );
  AO22X1_HVT U2948 ( .A1(\ram[13][43] ), .A2(n5377), .A3(n5378), .A4(data[43]), 
        .Y(n3432) );
  AO22X1_HVT U2949 ( .A1(\ram[13][42] ), .A2(n5377), .A3(n5378), .A4(data[42]), 
        .Y(n3431) );
  AO22X1_HVT U2950 ( .A1(\ram[13][41] ), .A2(n5377), .A3(n5378), .A4(data[41]), 
        .Y(n3430) );
  AO22X1_HVT U2951 ( .A1(\ram[1][26] ), .A2(n5368), .A3(n5369), .A4(data[26]), 
        .Y(n343) );
  AO22X1_HVT U2952 ( .A1(\ram[13][40] ), .A2(n5377), .A3(n5378), .A4(data[40]), 
        .Y(n3429) );
  AO22X1_HVT U2953 ( .A1(\ram[13][39] ), .A2(n5377), .A3(n5378), .A4(data[39]), 
        .Y(n3428) );
  AO22X1_HVT U2954 ( .A1(\ram[13][38] ), .A2(n5377), .A3(n5378), .A4(data[38]), 
        .Y(n3427) );
  AO22X1_HVT U2955 ( .A1(\ram[13][37] ), .A2(n5377), .A3(n5378), .A4(data[37]), 
        .Y(n3426) );
  AO22X1_HVT U2956 ( .A1(\ram[13][36] ), .A2(n5377), .A3(n5378), .A4(data[36]), 
        .Y(n3425) );
  AO22X1_HVT U2957 ( .A1(\ram[13][35] ), .A2(n5377), .A3(n5378), .A4(data[35]), 
        .Y(n3424) );
  AO22X1_HVT U2958 ( .A1(\ram[13][34] ), .A2(n5377), .A3(n5378), .A4(data[34]), 
        .Y(n3423) );
  AO22X1_HVT U2959 ( .A1(\ram[13][33] ), .A2(n5377), .A3(n5378), .A4(data[33]), 
        .Y(n3422) );
  AO22X1_HVT U2960 ( .A1(\ram[13][32] ), .A2(n5377), .A3(n5378), .A4(data[32]), 
        .Y(n3421) );
  AO22X1_HVT U2961 ( .A1(\ram[13][31] ), .A2(n5377), .A3(n5378), .A4(data[31]), 
        .Y(n3420) );
  AO22X1_HVT U2962 ( .A1(\ram[1][25] ), .A2(n5368), .A3(n5369), .A4(data[25]), 
        .Y(n342) );
  AO22X1_HVT U2963 ( .A1(\ram[13][30] ), .A2(n5377), .A3(n5378), .A4(data[30]), 
        .Y(n3419) );
  AO22X1_HVT U2964 ( .A1(\ram[13][29] ), .A2(n5377), .A3(n5378), .A4(data[29]), 
        .Y(n3418) );
  AO22X1_HVT U2965 ( .A1(\ram[13][28] ), .A2(n5377), .A3(n5378), .A4(data[28]), 
        .Y(n3417) );
  AO22X1_HVT U2966 ( .A1(\ram[13][27] ), .A2(n5377), .A3(n5378), .A4(data[27]), 
        .Y(n3416) );
  AO22X1_HVT U2967 ( .A1(\ram[13][26] ), .A2(n5377), .A3(n5378), .A4(data[26]), 
        .Y(n3415) );
  AO22X1_HVT U2968 ( .A1(\ram[13][25] ), .A2(n5377), .A3(n5378), .A4(data[25]), 
        .Y(n3414) );
  AO22X1_HVT U2969 ( .A1(\ram[13][24] ), .A2(n5377), .A3(n5378), .A4(data[24]), 
        .Y(n3413) );
  AO22X1_HVT U2970 ( .A1(\ram[13][23] ), .A2(n5377), .A3(n5378), .A4(data[23]), 
        .Y(n3412) );
  AO22X1_HVT U2971 ( .A1(\ram[13][22] ), .A2(n5377), .A3(n5378), .A4(data[22]), 
        .Y(n3411) );
  AO22X1_HVT U2972 ( .A1(\ram[13][21] ), .A2(n5377), .A3(n5378), .A4(data[21]), 
        .Y(n3410) );
  AO22X1_HVT U2973 ( .A1(\ram[1][24] ), .A2(n5368), .A3(n5369), .A4(data[24]), 
        .Y(n341) );
  AO22X1_HVT U2974 ( .A1(\ram[13][20] ), .A2(n5377), .A3(n5378), .A4(data[20]), 
        .Y(n3409) );
  AO22X1_HVT U2975 ( .A1(\ram[13][19] ), .A2(n5377), .A3(n5378), .A4(data[19]), 
        .Y(n3408) );
  AO22X1_HVT U2976 ( .A1(\ram[13][18] ), .A2(n5377), .A3(n5378), .A4(data[18]), 
        .Y(n3407) );
  AO22X1_HVT U2977 ( .A1(\ram[13][17] ), .A2(n5377), .A3(n5378), .A4(data[17]), 
        .Y(n3406) );
  AO22X1_HVT U2978 ( .A1(\ram[13][16] ), .A2(n5377), .A3(n5378), .A4(data[16]), 
        .Y(n3405) );
  AO22X1_HVT U2979 ( .A1(\ram[13][15] ), .A2(n5377), .A3(n5378), .A4(data[15]), 
        .Y(n3404) );
  AO22X1_HVT U2980 ( .A1(\ram[13][14] ), .A2(n5377), .A3(n5378), .A4(data[14]), 
        .Y(n3403) );
  AO22X1_HVT U2981 ( .A1(\ram[13][13] ), .A2(n5377), .A3(n5378), .A4(data[13]), 
        .Y(n3402) );
  AO22X1_HVT U2982 ( .A1(\ram[13][12] ), .A2(n5377), .A3(n5378), .A4(data[12]), 
        .Y(n3401) );
  AO22X1_HVT U2983 ( .A1(\ram[13][11] ), .A2(n5377), .A3(n5378), .A4(data[11]), 
        .Y(n3400) );
  AO22X1_HVT U2984 ( .A1(\ram[1][23] ), .A2(n5368), .A3(n5369), .A4(data[23]), 
        .Y(n340) );
  AO22X1_HVT U2985 ( .A1(\ram[13][10] ), .A2(n5377), .A3(n5378), .A4(data[10]), 
        .Y(n3399) );
  AO22X1_HVT U2986 ( .A1(\ram[13][9] ), .A2(n5377), .A3(n5378), .A4(data[9]), 
        .Y(n3398) );
  AO22X1_HVT U2987 ( .A1(\ram[13][8] ), .A2(n5377), .A3(n5378), .A4(data[8]), 
        .Y(n3397) );
  AO22X1_HVT U2988 ( .A1(\ram[13][7] ), .A2(n5377), .A3(n5378), .A4(data[7]), 
        .Y(n3396) );
  AO22X1_HVT U2989 ( .A1(\ram[13][6] ), .A2(n5377), .A3(n5378), .A4(data[6]), 
        .Y(n3395) );
  AO22X1_HVT U2990 ( .A1(\ram[13][5] ), .A2(n5377), .A3(n5378), .A4(data[5]), 
        .Y(n3394) );
  AO22X1_HVT U2991 ( .A1(\ram[13][4] ), .A2(n5377), .A3(n5378), .A4(data[4]), 
        .Y(n3393) );
  AO22X1_HVT U2992 ( .A1(\ram[13][3] ), .A2(n5377), .A3(n5378), .A4(data[3]), 
        .Y(n3392) );
  AO22X1_HVT U2993 ( .A1(\ram[13][2] ), .A2(n5377), .A3(n5378), .A4(data[2]), 
        .Y(n3391) );
  AO22X1_HVT U2994 ( .A1(\ram[13][1] ), .A2(n5377), .A3(n5378), .A4(data[1]), 
        .Y(n3390) );
  AO22X1_HVT U2995 ( .A1(\ram[1][22] ), .A2(n5368), .A3(n5369), .A4(data[22]), 
        .Y(n339) );
  AO22X1_HVT U2996 ( .A1(\ram[13][0] ), .A2(n5377), .A3(n5378), .A4(data[0]), 
        .Y(n3389) );
  INVX0_HVT U2997 ( .A(n5379), .Y(n5378) );
  AND2X1_HVT U2998 ( .A1(n5379), .A2(n5365), .Y(n5377) );
  NAND3X0_HVT U2999 ( .A1(n4182), .A2(n4280), .A3(n5373), .Y(n5379) );
  AO22X1_HVT U3000 ( .A1(\ram[12][255] ), .A2(n5380), .A3(n5381), .A4(
        data[255]), .Y(n3388) );
  AO22X1_HVT U3001 ( .A1(\ram[12][254] ), .A2(n5380), .A3(n5381), .A4(
        data[254]), .Y(n3387) );
  AO22X1_HVT U3002 ( .A1(\ram[12][253] ), .A2(n5380), .A3(n5381), .A4(
        data[253]), .Y(n3386) );
  AO22X1_HVT U3003 ( .A1(\ram[12][252] ), .A2(n5380), .A3(n5381), .A4(
        data[252]), .Y(n3385) );
  AO22X1_HVT U3004 ( .A1(\ram[12][251] ), .A2(n5380), .A3(n5381), .A4(
        data[251]), .Y(n3384) );
  AO22X1_HVT U3005 ( .A1(\ram[12][250] ), .A2(n5380), .A3(n5381), .A4(
        data[250]), .Y(n3383) );
  AO22X1_HVT U3006 ( .A1(\ram[12][249] ), .A2(n5380), .A3(n5381), .A4(
        data[249]), .Y(n3382) );
  AO22X1_HVT U3007 ( .A1(\ram[12][248] ), .A2(n5380), .A3(n5381), .A4(
        data[248]), .Y(n3381) );
  AO22X1_HVT U3008 ( .A1(\ram[12][247] ), .A2(n5380), .A3(n5381), .A4(
        data[247]), .Y(n3380) );
  AO22X1_HVT U3009 ( .A1(\ram[1][21] ), .A2(n5368), .A3(n5369), .A4(data[21]), 
        .Y(n338) );
  AO22X1_HVT U3010 ( .A1(\ram[12][246] ), .A2(n5380), .A3(n5381), .A4(
        data[246]), .Y(n3379) );
  AO22X1_HVT U3011 ( .A1(\ram[12][245] ), .A2(n5380), .A3(n5381), .A4(
        data[245]), .Y(n3378) );
  AO22X1_HVT U3012 ( .A1(\ram[12][244] ), .A2(n5380), .A3(n5381), .A4(
        data[244]), .Y(n3377) );
  AO22X1_HVT U3013 ( .A1(\ram[12][243] ), .A2(n5380), .A3(n5381), .A4(
        data[243]), .Y(n3376) );
  AO22X1_HVT U3014 ( .A1(\ram[12][242] ), .A2(n5380), .A3(n5381), .A4(
        data[242]), .Y(n3375) );
  AO22X1_HVT U3015 ( .A1(\ram[12][241] ), .A2(n5380), .A3(n5381), .A4(
        data[241]), .Y(n3374) );
  AO22X1_HVT U3016 ( .A1(\ram[12][240] ), .A2(n5380), .A3(n5381), .A4(
        data[240]), .Y(n3373) );
  AO22X1_HVT U3017 ( .A1(\ram[12][239] ), .A2(n5380), .A3(n5381), .A4(
        data[239]), .Y(n3372) );
  AO22X1_HVT U3018 ( .A1(\ram[12][238] ), .A2(n5380), .A3(n5381), .A4(
        data[238]), .Y(n3371) );
  AO22X1_HVT U3019 ( .A1(\ram[12][237] ), .A2(n5380), .A3(n5381), .A4(
        data[237]), .Y(n3370) );
  AO22X1_HVT U3020 ( .A1(\ram[1][20] ), .A2(n5368), .A3(n5369), .A4(data[20]), 
        .Y(n337) );
  AO22X1_HVT U3021 ( .A1(\ram[12][236] ), .A2(n5380), .A3(n5381), .A4(
        data[236]), .Y(n3369) );
  AO22X1_HVT U3022 ( .A1(\ram[12][235] ), .A2(n5380), .A3(n5381), .A4(
        data[235]), .Y(n3368) );
  AO22X1_HVT U3023 ( .A1(\ram[12][234] ), .A2(n5380), .A3(n5381), .A4(
        data[234]), .Y(n3367) );
  AO22X1_HVT U3024 ( .A1(\ram[12][233] ), .A2(n5380), .A3(n5381), .A4(
        data[233]), .Y(n3366) );
  AO22X1_HVT U3025 ( .A1(\ram[12][232] ), .A2(n5380), .A3(n5381), .A4(
        data[232]), .Y(n3365) );
  AO22X1_HVT U3026 ( .A1(\ram[12][231] ), .A2(n5380), .A3(n5381), .A4(
        data[231]), .Y(n3364) );
  AO22X1_HVT U3027 ( .A1(\ram[12][230] ), .A2(n5380), .A3(n5381), .A4(
        data[230]), .Y(n3363) );
  AO22X1_HVT U3028 ( .A1(\ram[12][229] ), .A2(n5380), .A3(n5381), .A4(
        data[229]), .Y(n3362) );
  AO22X1_HVT U3029 ( .A1(\ram[12][228] ), .A2(n5380), .A3(n5381), .A4(
        data[228]), .Y(n3361) );
  AO22X1_HVT U3030 ( .A1(\ram[12][227] ), .A2(n5380), .A3(n5381), .A4(
        data[227]), .Y(n3360) );
  AO22X1_HVT U3031 ( .A1(\ram[1][19] ), .A2(n5368), .A3(n5369), .A4(data[19]), 
        .Y(n336) );
  AO22X1_HVT U3032 ( .A1(\ram[12][226] ), .A2(n5380), .A3(n5381), .A4(
        data[226]), .Y(n3359) );
  AO22X1_HVT U3033 ( .A1(\ram[12][225] ), .A2(n5380), .A3(n5381), .A4(
        data[225]), .Y(n3358) );
  AO22X1_HVT U3034 ( .A1(\ram[12][224] ), .A2(n5380), .A3(n5381), .A4(
        data[224]), .Y(n3357) );
  AO22X1_HVT U3035 ( .A1(\ram[12][223] ), .A2(n5380), .A3(n5381), .A4(
        data[223]), .Y(n3356) );
  AO22X1_HVT U3036 ( .A1(\ram[12][222] ), .A2(n5380), .A3(n5381), .A4(
        data[222]), .Y(n3355) );
  AO22X1_HVT U3037 ( .A1(\ram[12][221] ), .A2(n5380), .A3(n5381), .A4(
        data[221]), .Y(n3354) );
  AO22X1_HVT U3038 ( .A1(\ram[12][220] ), .A2(n5380), .A3(n5381), .A4(
        data[220]), .Y(n3353) );
  AO22X1_HVT U3039 ( .A1(\ram[12][219] ), .A2(n5380), .A3(n5381), .A4(
        data[219]), .Y(n3352) );
  AO22X1_HVT U3040 ( .A1(\ram[12][218] ), .A2(n5380), .A3(n5381), .A4(
        data[218]), .Y(n3351) );
  AO22X1_HVT U3041 ( .A1(\ram[12][217] ), .A2(n5380), .A3(n5381), .A4(
        data[217]), .Y(n3350) );
  AO22X1_HVT U3042 ( .A1(\ram[1][18] ), .A2(n5368), .A3(n5369), .A4(data[18]), 
        .Y(n335) );
  AO22X1_HVT U3043 ( .A1(\ram[12][216] ), .A2(n5380), .A3(n5381), .A4(
        data[216]), .Y(n3349) );
  AO22X1_HVT U3044 ( .A1(\ram[12][215] ), .A2(n5380), .A3(n5381), .A4(
        data[215]), .Y(n3348) );
  AO22X1_HVT U3045 ( .A1(\ram[12][214] ), .A2(n5380), .A3(n5381), .A4(
        data[214]), .Y(n3347) );
  AO22X1_HVT U3046 ( .A1(\ram[12][213] ), .A2(n5380), .A3(n5381), .A4(
        data[213]), .Y(n3346) );
  AO22X1_HVT U3047 ( .A1(\ram[12][212] ), .A2(n5380), .A3(n5381), .A4(
        data[212]), .Y(n3345) );
  AO22X1_HVT U3048 ( .A1(\ram[12][211] ), .A2(n5380), .A3(n5381), .A4(
        data[211]), .Y(n3344) );
  AO22X1_HVT U3049 ( .A1(\ram[12][210] ), .A2(n5380), .A3(n5381), .A4(
        data[210]), .Y(n3343) );
  AO22X1_HVT U3050 ( .A1(\ram[12][209] ), .A2(n5380), .A3(n5381), .A4(
        data[209]), .Y(n3342) );
  AO22X1_HVT U3051 ( .A1(\ram[12][208] ), .A2(n5380), .A3(n5381), .A4(
        data[208]), .Y(n3341) );
  AO22X1_HVT U3052 ( .A1(\ram[12][207] ), .A2(n5380), .A3(n5381), .A4(
        data[207]), .Y(n3340) );
  AO22X1_HVT U3053 ( .A1(\ram[1][17] ), .A2(n5368), .A3(n5369), .A4(data[17]), 
        .Y(n334) );
  AO22X1_HVT U3054 ( .A1(\ram[12][206] ), .A2(n5380), .A3(n5381), .A4(
        data[206]), .Y(n3339) );
  AO22X1_HVT U3055 ( .A1(\ram[12][205] ), .A2(n5380), .A3(n5381), .A4(
        data[205]), .Y(n3338) );
  AO22X1_HVT U3056 ( .A1(\ram[12][204] ), .A2(n5380), .A3(n5381), .A4(
        data[204]), .Y(n3337) );
  AO22X1_HVT U3057 ( .A1(\ram[12][203] ), .A2(n5380), .A3(n5381), .A4(
        data[203]), .Y(n3336) );
  AO22X1_HVT U3058 ( .A1(\ram[12][202] ), .A2(n5380), .A3(n5381), .A4(
        data[202]), .Y(n3335) );
  AO22X1_HVT U3059 ( .A1(\ram[12][201] ), .A2(n5380), .A3(n5381), .A4(
        data[201]), .Y(n3334) );
  AO22X1_HVT U3060 ( .A1(\ram[12][200] ), .A2(n5380), .A3(n5381), .A4(
        data[200]), .Y(n3333) );
  AO22X1_HVT U3061 ( .A1(\ram[12][199] ), .A2(n5380), .A3(n5381), .A4(
        data[199]), .Y(n3332) );
  AO22X1_HVT U3062 ( .A1(\ram[12][198] ), .A2(n5380), .A3(n5381), .A4(
        data[198]), .Y(n3331) );
  AO22X1_HVT U3063 ( .A1(\ram[12][197] ), .A2(n5380), .A3(n5381), .A4(
        data[197]), .Y(n3330) );
  AO22X1_HVT U3064 ( .A1(\ram[1][16] ), .A2(n5368), .A3(n5369), .A4(data[16]), 
        .Y(n333) );
  AO22X1_HVT U3065 ( .A1(\ram[12][196] ), .A2(n5380), .A3(n5381), .A4(
        data[196]), .Y(n3329) );
  AO22X1_HVT U3066 ( .A1(\ram[12][195] ), .A2(n5380), .A3(n5381), .A4(
        data[195]), .Y(n3328) );
  AO22X1_HVT U3067 ( .A1(\ram[12][194] ), .A2(n5380), .A3(n5381), .A4(
        data[194]), .Y(n3327) );
  AO22X1_HVT U3068 ( .A1(\ram[12][193] ), .A2(n5380), .A3(n5381), .A4(
        data[193]), .Y(n3326) );
  AO22X1_HVT U3069 ( .A1(\ram[12][192] ), .A2(n5380), .A3(n5381), .A4(
        data[192]), .Y(n3325) );
  AO22X1_HVT U3070 ( .A1(\ram[12][191] ), .A2(n5380), .A3(n5381), .A4(
        data[191]), .Y(n3324) );
  AO22X1_HVT U3071 ( .A1(\ram[12][190] ), .A2(n5380), .A3(n5381), .A4(
        data[190]), .Y(n3323) );
  AO22X1_HVT U3072 ( .A1(\ram[12][189] ), .A2(n5380), .A3(n5381), .A4(
        data[189]), .Y(n3322) );
  AO22X1_HVT U3073 ( .A1(\ram[12][188] ), .A2(n5380), .A3(n5381), .A4(
        data[188]), .Y(n3321) );
  AO22X1_HVT U3074 ( .A1(\ram[12][187] ), .A2(n5380), .A3(n5381), .A4(
        data[187]), .Y(n3320) );
  AO22X1_HVT U3075 ( .A1(\ram[1][15] ), .A2(n5368), .A3(n5369), .A4(data[15]), 
        .Y(n332) );
  AO22X1_HVT U3076 ( .A1(\ram[12][186] ), .A2(n5380), .A3(n5381), .A4(
        data[186]), .Y(n3319) );
  AO22X1_HVT U3077 ( .A1(\ram[12][185] ), .A2(n5380), .A3(n5381), .A4(
        data[185]), .Y(n3318) );
  AO22X1_HVT U3078 ( .A1(\ram[12][184] ), .A2(n5380), .A3(n5381), .A4(
        data[184]), .Y(n3317) );
  AO22X1_HVT U3079 ( .A1(\ram[12][183] ), .A2(n5380), .A3(n5381), .A4(
        data[183]), .Y(n3316) );
  AO22X1_HVT U3080 ( .A1(\ram[12][182] ), .A2(n5380), .A3(n5381), .A4(
        data[182]), .Y(n3315) );
  AO22X1_HVT U3081 ( .A1(\ram[12][181] ), .A2(n5380), .A3(n5381), .A4(
        data[181]), .Y(n3314) );
  AO22X1_HVT U3082 ( .A1(\ram[12][180] ), .A2(n5380), .A3(n5381), .A4(
        data[180]), .Y(n3313) );
  AO22X1_HVT U3083 ( .A1(\ram[12][179] ), .A2(n5380), .A3(n5381), .A4(
        data[179]), .Y(n3312) );
  AO22X1_HVT U3084 ( .A1(\ram[12][178] ), .A2(n5380), .A3(n5381), .A4(
        data[178]), .Y(n3311) );
  AO22X1_HVT U3085 ( .A1(\ram[12][177] ), .A2(n5380), .A3(n5381), .A4(
        data[177]), .Y(n3310) );
  AO22X1_HVT U3086 ( .A1(\ram[1][14] ), .A2(n5368), .A3(n5369), .A4(data[14]), 
        .Y(n331) );
  AO22X1_HVT U3087 ( .A1(\ram[12][176] ), .A2(n5380), .A3(n5381), .A4(
        data[176]), .Y(n3309) );
  AO22X1_HVT U3088 ( .A1(\ram[12][175] ), .A2(n5380), .A3(n5381), .A4(
        data[175]), .Y(n3308) );
  AO22X1_HVT U3089 ( .A1(\ram[12][174] ), .A2(n5380), .A3(n5381), .A4(
        data[174]), .Y(n3307) );
  AO22X1_HVT U3090 ( .A1(\ram[12][173] ), .A2(n5380), .A3(n5381), .A4(
        data[173]), .Y(n3306) );
  AO22X1_HVT U3091 ( .A1(\ram[12][172] ), .A2(n5380), .A3(n5381), .A4(
        data[172]), .Y(n3305) );
  AO22X1_HVT U3092 ( .A1(\ram[12][171] ), .A2(n5380), .A3(n5381), .A4(
        data[171]), .Y(n3304) );
  AO22X1_HVT U3093 ( .A1(\ram[12][170] ), .A2(n5380), .A3(n5381), .A4(
        data[170]), .Y(n3303) );
  AO22X1_HVT U3094 ( .A1(\ram[12][169] ), .A2(n5380), .A3(n5381), .A4(
        data[169]), .Y(n3302) );
  AO22X1_HVT U3095 ( .A1(\ram[12][168] ), .A2(n5380), .A3(n5381), .A4(
        data[168]), .Y(n3301) );
  AO22X1_HVT U3096 ( .A1(\ram[12][167] ), .A2(n5380), .A3(n5381), .A4(
        data[167]), .Y(n3300) );
  AO22X1_HVT U3097 ( .A1(\ram[1][13] ), .A2(n5368), .A3(n5369), .A4(data[13]), 
        .Y(n330) );
  AO22X1_HVT U3098 ( .A1(\ram[12][166] ), .A2(n5380), .A3(n5381), .A4(
        data[166]), .Y(n3299) );
  AO22X1_HVT U3099 ( .A1(\ram[12][165] ), .A2(n5380), .A3(n5381), .A4(
        data[165]), .Y(n3298) );
  AO22X1_HVT U3100 ( .A1(\ram[12][164] ), .A2(n5380), .A3(n5381), .A4(
        data[164]), .Y(n3297) );
  AO22X1_HVT U3101 ( .A1(\ram[12][163] ), .A2(n5380), .A3(n5381), .A4(
        data[163]), .Y(n3296) );
  AO22X1_HVT U3102 ( .A1(\ram[12][162] ), .A2(n5380), .A3(n5381), .A4(
        data[162]), .Y(n3295) );
  AO22X1_HVT U3103 ( .A1(\ram[12][161] ), .A2(n5380), .A3(n5381), .A4(
        data[161]), .Y(n3294) );
  AO22X1_HVT U3104 ( .A1(\ram[12][160] ), .A2(n5380), .A3(n5381), .A4(
        data[160]), .Y(n3293) );
  AO22X1_HVT U3105 ( .A1(\ram[12][159] ), .A2(n5380), .A3(n5381), .A4(
        data[159]), .Y(n3292) );
  AO22X1_HVT U3106 ( .A1(\ram[12][158] ), .A2(n5380), .A3(n5381), .A4(
        data[158]), .Y(n3291) );
  AO22X1_HVT U3107 ( .A1(\ram[12][157] ), .A2(n5380), .A3(n5381), .A4(
        data[157]), .Y(n3290) );
  AO22X1_HVT U3108 ( .A1(\ram[1][12] ), .A2(n5368), .A3(n5369), .A4(data[12]), 
        .Y(n329) );
  AO22X1_HVT U3109 ( .A1(\ram[12][156] ), .A2(n5380), .A3(n5381), .A4(
        data[156]), .Y(n3289) );
  AO22X1_HVT U3110 ( .A1(\ram[12][155] ), .A2(n5380), .A3(n5381), .A4(
        data[155]), .Y(n3288) );
  AO22X1_HVT U3111 ( .A1(\ram[12][154] ), .A2(n5380), .A3(n5381), .A4(
        data[154]), .Y(n3287) );
  AO22X1_HVT U3112 ( .A1(\ram[12][153] ), .A2(n5380), .A3(n5381), .A4(
        data[153]), .Y(n3286) );
  AO22X1_HVT U3113 ( .A1(\ram[12][152] ), .A2(n5380), .A3(n5381), .A4(
        data[152]), .Y(n3285) );
  AO22X1_HVT U3114 ( .A1(\ram[12][151] ), .A2(n5380), .A3(n5381), .A4(
        data[151]), .Y(n3284) );
  AO22X1_HVT U3115 ( .A1(\ram[12][150] ), .A2(n5380), .A3(n5381), .A4(
        data[150]), .Y(n3283) );
  AO22X1_HVT U3116 ( .A1(\ram[12][149] ), .A2(n5380), .A3(n5381), .A4(
        data[149]), .Y(n3282) );
  AO22X1_HVT U3117 ( .A1(\ram[12][148] ), .A2(n5380), .A3(n5381), .A4(
        data[148]), .Y(n3281) );
  AO22X1_HVT U3118 ( .A1(\ram[12][147] ), .A2(n5380), .A3(n5381), .A4(
        data[147]), .Y(n3280) );
  AO22X1_HVT U3119 ( .A1(\ram[1][11] ), .A2(n5368), .A3(n5369), .A4(data[11]), 
        .Y(n328) );
  AO22X1_HVT U3120 ( .A1(\ram[12][146] ), .A2(n5380), .A3(n5381), .A4(
        data[146]), .Y(n3279) );
  AO22X1_HVT U3121 ( .A1(\ram[12][145] ), .A2(n5380), .A3(n5381), .A4(
        data[145]), .Y(n3278) );
  AO22X1_HVT U3122 ( .A1(\ram[12][144] ), .A2(n5380), .A3(n5381), .A4(
        data[144]), .Y(n3277) );
  AO22X1_HVT U3123 ( .A1(\ram[12][143] ), .A2(n5380), .A3(n5381), .A4(
        data[143]), .Y(n3276) );
  AO22X1_HVT U3124 ( .A1(\ram[12][142] ), .A2(n5380), .A3(n5381), .A4(
        data[142]), .Y(n3275) );
  AO22X1_HVT U3125 ( .A1(\ram[12][141] ), .A2(n5380), .A3(n5381), .A4(
        data[141]), .Y(n3274) );
  AO22X1_HVT U3126 ( .A1(\ram[12][140] ), .A2(n5380), .A3(n5381), .A4(
        data[140]), .Y(n3273) );
  AO22X1_HVT U3127 ( .A1(\ram[12][139] ), .A2(n5380), .A3(n5381), .A4(
        data[139]), .Y(n3272) );
  AO22X1_HVT U3128 ( .A1(\ram[12][138] ), .A2(n5380), .A3(n5381), .A4(
        data[138]), .Y(n3271) );
  AO22X1_HVT U3129 ( .A1(\ram[12][137] ), .A2(n5380), .A3(n5381), .A4(
        data[137]), .Y(n3270) );
  AO22X1_HVT U3130 ( .A1(\ram[1][10] ), .A2(n5368), .A3(n5369), .A4(data[10]), 
        .Y(n327) );
  AO22X1_HVT U3131 ( .A1(\ram[12][136] ), .A2(n5380), .A3(n5381), .A4(
        data[136]), .Y(n3269) );
  AO22X1_HVT U3132 ( .A1(\ram[12][135] ), .A2(n5380), .A3(n5381), .A4(
        data[135]), .Y(n3268) );
  AO22X1_HVT U3133 ( .A1(\ram[12][134] ), .A2(n5380), .A3(n5381), .A4(
        data[134]), .Y(n3267) );
  AO22X1_HVT U3134 ( .A1(\ram[12][133] ), .A2(n5380), .A3(n5381), .A4(
        data[133]), .Y(n3266) );
  AO22X1_HVT U3135 ( .A1(\ram[12][132] ), .A2(n5380), .A3(n5381), .A4(
        data[132]), .Y(n3265) );
  AO22X1_HVT U3136 ( .A1(\ram[12][131] ), .A2(n5380), .A3(n5381), .A4(
        data[131]), .Y(n3264) );
  AO22X1_HVT U3137 ( .A1(\ram[12][130] ), .A2(n5380), .A3(n5381), .A4(
        data[130]), .Y(n3263) );
  AO22X1_HVT U3138 ( .A1(\ram[12][129] ), .A2(n5380), .A3(n5381), .A4(
        data[129]), .Y(n3262) );
  AO22X1_HVT U3139 ( .A1(\ram[12][128] ), .A2(n5380), .A3(n5381), .A4(
        data[128]), .Y(n3261) );
  AO22X1_HVT U3140 ( .A1(\ram[12][127] ), .A2(n5380), .A3(n5381), .A4(
        data[127]), .Y(n3260) );
  AO22X1_HVT U3141 ( .A1(\ram[1][9] ), .A2(n5368), .A3(n5369), .A4(data[9]), 
        .Y(n326) );
  AO22X1_HVT U3142 ( .A1(\ram[12][126] ), .A2(n5380), .A3(n5381), .A4(
        data[126]), .Y(n3259) );
  AO22X1_HVT U3143 ( .A1(\ram[12][125] ), .A2(n5380), .A3(n5381), .A4(
        data[125]), .Y(n3258) );
  AO22X1_HVT U3144 ( .A1(\ram[12][124] ), .A2(n5380), .A3(n5381), .A4(
        data[124]), .Y(n3257) );
  AO22X1_HVT U3145 ( .A1(\ram[12][123] ), .A2(n5380), .A3(n5381), .A4(
        data[123]), .Y(n3256) );
  AO22X1_HVT U3146 ( .A1(\ram[12][122] ), .A2(n5380), .A3(n5381), .A4(
        data[122]), .Y(n3255) );
  AO22X1_HVT U3147 ( .A1(\ram[12][121] ), .A2(n5380), .A3(n5381), .A4(
        data[121]), .Y(n3254) );
  AO22X1_HVT U3148 ( .A1(\ram[12][120] ), .A2(n5380), .A3(n5381), .A4(
        data[120]), .Y(n3253) );
  AO22X1_HVT U3149 ( .A1(\ram[12][119] ), .A2(n5380), .A3(n5381), .A4(
        data[119]), .Y(n3252) );
  AO22X1_HVT U3150 ( .A1(\ram[12][118] ), .A2(n5380), .A3(n5381), .A4(
        data[118]), .Y(n3251) );
  AO22X1_HVT U3151 ( .A1(\ram[12][117] ), .A2(n5380), .A3(n5381), .A4(
        data[117]), .Y(n3250) );
  AO22X1_HVT U3152 ( .A1(\ram[1][8] ), .A2(n5368), .A3(n5369), .A4(data[8]), 
        .Y(n325) );
  AO22X1_HVT U3153 ( .A1(\ram[12][116] ), .A2(n5380), .A3(n5381), .A4(
        data[116]), .Y(n3249) );
  AO22X1_HVT U3154 ( .A1(\ram[12][115] ), .A2(n5380), .A3(n5381), .A4(
        data[115]), .Y(n3248) );
  AO22X1_HVT U3155 ( .A1(\ram[12][114] ), .A2(n5380), .A3(n5381), .A4(
        data[114]), .Y(n3247) );
  AO22X1_HVT U3156 ( .A1(\ram[12][113] ), .A2(n5380), .A3(n5381), .A4(
        data[113]), .Y(n3246) );
  AO22X1_HVT U3157 ( .A1(\ram[12][112] ), .A2(n5380), .A3(n5381), .A4(
        data[112]), .Y(n3245) );
  AO22X1_HVT U3158 ( .A1(\ram[12][111] ), .A2(n5380), .A3(n5381), .A4(
        data[111]), .Y(n3244) );
  AO22X1_HVT U3159 ( .A1(\ram[12][110] ), .A2(n5380), .A3(n5381), .A4(
        data[110]), .Y(n3243) );
  AO22X1_HVT U3160 ( .A1(\ram[12][109] ), .A2(n5380), .A3(n5381), .A4(
        data[109]), .Y(n3242) );
  AO22X1_HVT U3161 ( .A1(\ram[12][108] ), .A2(n5380), .A3(n5381), .A4(
        data[108]), .Y(n3241) );
  AO22X1_HVT U3162 ( .A1(\ram[12][107] ), .A2(n5380), .A3(n5381), .A4(
        data[107]), .Y(n3240) );
  AO22X1_HVT U3163 ( .A1(\ram[1][7] ), .A2(n5368), .A3(n5369), .A4(data[7]), 
        .Y(n324) );
  AO22X1_HVT U3164 ( .A1(\ram[12][106] ), .A2(n5380), .A3(n5381), .A4(
        data[106]), .Y(n3239) );
  AO22X1_HVT U3165 ( .A1(\ram[12][105] ), .A2(n5380), .A3(n5381), .A4(
        data[105]), .Y(n3238) );
  AO22X1_HVT U3166 ( .A1(\ram[12][104] ), .A2(n5380), .A3(n5381), .A4(
        data[104]), .Y(n3237) );
  AO22X1_HVT U3167 ( .A1(\ram[12][103] ), .A2(n5380), .A3(n5381), .A4(
        data[103]), .Y(n3236) );
  AO22X1_HVT U3168 ( .A1(\ram[12][102] ), .A2(n5380), .A3(n5381), .A4(
        data[102]), .Y(n3235) );
  AO22X1_HVT U3169 ( .A1(\ram[12][101] ), .A2(n5380), .A3(n5381), .A4(
        data[101]), .Y(n3234) );
  AO22X1_HVT U3170 ( .A1(\ram[12][100] ), .A2(n5380), .A3(n5381), .A4(
        data[100]), .Y(n3233) );
  AO22X1_HVT U3171 ( .A1(\ram[12][99] ), .A2(n5380), .A3(n5381), .A4(data[99]), 
        .Y(n3232) );
  AO22X1_HVT U3172 ( .A1(\ram[12][98] ), .A2(n5380), .A3(n5381), .A4(data[98]), 
        .Y(n3231) );
  AO22X1_HVT U3173 ( .A1(\ram[12][97] ), .A2(n5380), .A3(n5381), .A4(data[97]), 
        .Y(n3230) );
  AO22X1_HVT U3174 ( .A1(\ram[1][6] ), .A2(n5368), .A3(n5369), .A4(data[6]), 
        .Y(n323) );
  AO22X1_HVT U3175 ( .A1(\ram[12][96] ), .A2(n5380), .A3(n5381), .A4(data[96]), 
        .Y(n3229) );
  AO22X1_HVT U3176 ( .A1(\ram[12][95] ), .A2(n5380), .A3(n5381), .A4(data[95]), 
        .Y(n3228) );
  AO22X1_HVT U3177 ( .A1(\ram[12][94] ), .A2(n5380), .A3(n5381), .A4(data[94]), 
        .Y(n3227) );
  AO22X1_HVT U3178 ( .A1(\ram[12][93] ), .A2(n5380), .A3(n5381), .A4(data[93]), 
        .Y(n3226) );
  AO22X1_HVT U3179 ( .A1(\ram[12][92] ), .A2(n5380), .A3(n5381), .A4(data[92]), 
        .Y(n3225) );
  AO22X1_HVT U3180 ( .A1(\ram[12][91] ), .A2(n5380), .A3(n5381), .A4(data[91]), 
        .Y(n3224) );
  AO22X1_HVT U3181 ( .A1(\ram[12][90] ), .A2(n5380), .A3(n5381), .A4(data[90]), 
        .Y(n3223) );
  AO22X1_HVT U3182 ( .A1(\ram[12][89] ), .A2(n5380), .A3(n5381), .A4(data[89]), 
        .Y(n3222) );
  AO22X1_HVT U3183 ( .A1(\ram[12][88] ), .A2(n5380), .A3(n5381), .A4(data[88]), 
        .Y(n3221) );
  AO22X1_HVT U3184 ( .A1(\ram[12][87] ), .A2(n5380), .A3(n5381), .A4(data[87]), 
        .Y(n3220) );
  AO22X1_HVT U3185 ( .A1(\ram[1][5] ), .A2(n5368), .A3(n5369), .A4(data[5]), 
        .Y(n322) );
  AO22X1_HVT U3186 ( .A1(\ram[12][86] ), .A2(n5380), .A3(n5381), .A4(data[86]), 
        .Y(n3219) );
  AO22X1_HVT U3187 ( .A1(\ram[12][85] ), .A2(n5380), .A3(n5381), .A4(data[85]), 
        .Y(n3218) );
  AO22X1_HVT U3188 ( .A1(\ram[12][84] ), .A2(n5380), .A3(n5381), .A4(data[84]), 
        .Y(n3217) );
  AO22X1_HVT U3189 ( .A1(\ram[12][83] ), .A2(n5380), .A3(n5381), .A4(data[83]), 
        .Y(n3216) );
  AO22X1_HVT U3190 ( .A1(\ram[12][82] ), .A2(n5380), .A3(n5381), .A4(data[82]), 
        .Y(n3215) );
  AO22X1_HVT U3191 ( .A1(\ram[12][81] ), .A2(n5380), .A3(n5381), .A4(data[81]), 
        .Y(n3214) );
  AO22X1_HVT U3192 ( .A1(\ram[12][80] ), .A2(n5380), .A3(n5381), .A4(data[80]), 
        .Y(n3213) );
  AO22X1_HVT U3193 ( .A1(\ram[12][79] ), .A2(n5380), .A3(n5381), .A4(data[79]), 
        .Y(n3212) );
  AO22X1_HVT U3194 ( .A1(\ram[12][78] ), .A2(n5380), .A3(n5381), .A4(data[78]), 
        .Y(n3211) );
  AO22X1_HVT U3195 ( .A1(\ram[12][77] ), .A2(n5380), .A3(n5381), .A4(data[77]), 
        .Y(n3210) );
  AO22X1_HVT U3196 ( .A1(\ram[1][4] ), .A2(n5368), .A3(n5369), .A4(data[4]), 
        .Y(n321) );
  AO22X1_HVT U3197 ( .A1(\ram[12][76] ), .A2(n5380), .A3(n5381), .A4(data[76]), 
        .Y(n3209) );
  AO22X1_HVT U3198 ( .A1(\ram[12][75] ), .A2(n5380), .A3(n5381), .A4(data[75]), 
        .Y(n3208) );
  AO22X1_HVT U3199 ( .A1(\ram[12][74] ), .A2(n5380), .A3(n5381), .A4(data[74]), 
        .Y(n3207) );
  AO22X1_HVT U3200 ( .A1(\ram[12][73] ), .A2(n5380), .A3(n5381), .A4(data[73]), 
        .Y(n3206) );
  AO22X1_HVT U3201 ( .A1(\ram[12][72] ), .A2(n5380), .A3(n5381), .A4(data[72]), 
        .Y(n3205) );
  AO22X1_HVT U3202 ( .A1(\ram[12][71] ), .A2(n5380), .A3(n5381), .A4(data[71]), 
        .Y(n3204) );
  AO22X1_HVT U3203 ( .A1(\ram[12][70] ), .A2(n5380), .A3(n5381), .A4(data[70]), 
        .Y(n3203) );
  AO22X1_HVT U3204 ( .A1(\ram[12][69] ), .A2(n5380), .A3(n5381), .A4(data[69]), 
        .Y(n3202) );
  AO22X1_HVT U3205 ( .A1(\ram[12][68] ), .A2(n5380), .A3(n5381), .A4(data[68]), 
        .Y(n3201) );
  AO22X1_HVT U3206 ( .A1(\ram[12][67] ), .A2(n5380), .A3(n5381), .A4(data[67]), 
        .Y(n3200) );
  AO22X1_HVT U3207 ( .A1(\ram[1][3] ), .A2(n5368), .A3(n5369), .A4(data[3]), 
        .Y(n320) );
  AO22X1_HVT U3208 ( .A1(\ram[12][66] ), .A2(n5380), .A3(n5381), .A4(data[66]), 
        .Y(n3199) );
  AO22X1_HVT U3209 ( .A1(\ram[12][65] ), .A2(n5380), .A3(n5381), .A4(data[65]), 
        .Y(n3198) );
  AO22X1_HVT U3210 ( .A1(\ram[12][64] ), .A2(n5380), .A3(n5381), .A4(data[64]), 
        .Y(n3197) );
  AO22X1_HVT U3211 ( .A1(\ram[12][63] ), .A2(n5380), .A3(n5381), .A4(data[63]), 
        .Y(n3196) );
  AO22X1_HVT U3212 ( .A1(\ram[12][62] ), .A2(n5380), .A3(n5381), .A4(data[62]), 
        .Y(n3195) );
  AO22X1_HVT U3213 ( .A1(\ram[12][61] ), .A2(n5380), .A3(n5381), .A4(data[61]), 
        .Y(n3194) );
  AO22X1_HVT U3214 ( .A1(\ram[12][60] ), .A2(n5380), .A3(n5381), .A4(data[60]), 
        .Y(n3193) );
  AO22X1_HVT U3215 ( .A1(\ram[12][59] ), .A2(n5380), .A3(n5381), .A4(data[59]), 
        .Y(n3192) );
  AO22X1_HVT U3216 ( .A1(\ram[12][58] ), .A2(n5380), .A3(n5381), .A4(data[58]), 
        .Y(n3191) );
  AO22X1_HVT U3217 ( .A1(\ram[12][57] ), .A2(n5380), .A3(n5381), .A4(data[57]), 
        .Y(n3190) );
  AO22X1_HVT U3218 ( .A1(\ram[1][2] ), .A2(n5368), .A3(n5369), .A4(data[2]), 
        .Y(n319) );
  AO22X1_HVT U3219 ( .A1(\ram[12][56] ), .A2(n5380), .A3(n5381), .A4(data[56]), 
        .Y(n3189) );
  AO22X1_HVT U3220 ( .A1(\ram[12][55] ), .A2(n5380), .A3(n5381), .A4(data[55]), 
        .Y(n3188) );
  AO22X1_HVT U3221 ( .A1(\ram[12][54] ), .A2(n5380), .A3(n5381), .A4(data[54]), 
        .Y(n3187) );
  AO22X1_HVT U3222 ( .A1(\ram[12][53] ), .A2(n5380), .A3(n5381), .A4(data[53]), 
        .Y(n3186) );
  AO22X1_HVT U3223 ( .A1(\ram[12][52] ), .A2(n5380), .A3(n5381), .A4(data[52]), 
        .Y(n3185) );
  AO22X1_HVT U3224 ( .A1(\ram[12][51] ), .A2(n5380), .A3(n5381), .A4(data[51]), 
        .Y(n3184) );
  AO22X1_HVT U3225 ( .A1(\ram[12][50] ), .A2(n5380), .A3(n5381), .A4(data[50]), 
        .Y(n3183) );
  AO22X1_HVT U3226 ( .A1(\ram[12][49] ), .A2(n5380), .A3(n5381), .A4(data[49]), 
        .Y(n3182) );
  AO22X1_HVT U3227 ( .A1(\ram[12][48] ), .A2(n5380), .A3(n5381), .A4(data[48]), 
        .Y(n3181) );
  AO22X1_HVT U3228 ( .A1(\ram[12][47] ), .A2(n5380), .A3(n5381), .A4(data[47]), 
        .Y(n3180) );
  AO22X1_HVT U3229 ( .A1(\ram[1][1] ), .A2(n5368), .A3(n5369), .A4(data[1]), 
        .Y(n318) );
  AO22X1_HVT U3230 ( .A1(\ram[12][46] ), .A2(n5380), .A3(n5381), .A4(data[46]), 
        .Y(n3179) );
  AO22X1_HVT U3231 ( .A1(\ram[12][45] ), .A2(n5380), .A3(n5381), .A4(data[45]), 
        .Y(n3178) );
  AO22X1_HVT U3232 ( .A1(\ram[12][44] ), .A2(n5380), .A3(n5381), .A4(data[44]), 
        .Y(n3177) );
  AO22X1_HVT U3233 ( .A1(\ram[12][43] ), .A2(n5380), .A3(n5381), .A4(data[43]), 
        .Y(n3176) );
  AO22X1_HVT U3234 ( .A1(\ram[12][42] ), .A2(n5380), .A3(n5381), .A4(data[42]), 
        .Y(n3175) );
  AO22X1_HVT U3235 ( .A1(\ram[12][41] ), .A2(n5380), .A3(n5381), .A4(data[41]), 
        .Y(n3174) );
  AO22X1_HVT U3236 ( .A1(\ram[12][40] ), .A2(n5380), .A3(n5381), .A4(data[40]), 
        .Y(n3173) );
  AO22X1_HVT U3237 ( .A1(\ram[12][39] ), .A2(n5380), .A3(n5381), .A4(data[39]), 
        .Y(n3172) );
  AO22X1_HVT U3238 ( .A1(\ram[12][38] ), .A2(n5380), .A3(n5381), .A4(data[38]), 
        .Y(n3171) );
  AO22X1_HVT U3239 ( .A1(\ram[12][37] ), .A2(n5380), .A3(n5381), .A4(data[37]), 
        .Y(n3170) );
  AO22X1_HVT U3240 ( .A1(\ram[1][0] ), .A2(n5368), .A3(n5369), .A4(data[0]), 
        .Y(n317) );
  INVX0_HVT U3241 ( .A(n5382), .Y(n5369) );
  AND2X1_HVT U3242 ( .A1(n5382), .A2(n5365), .Y(n5368) );
  NAND3X0_HVT U3243 ( .A1(n4182), .A2(n5367), .A3(n5383), .Y(n5382) );
  AO22X1_HVT U3244 ( .A1(\ram[12][36] ), .A2(n5380), .A3(n5381), .A4(data[36]), 
        .Y(n3169) );
  AO22X1_HVT U3245 ( .A1(\ram[12][35] ), .A2(n5380), .A3(n5381), .A4(data[35]), 
        .Y(n3168) );
  AO22X1_HVT U3246 ( .A1(\ram[12][34] ), .A2(n5380), .A3(n5381), .A4(data[34]), 
        .Y(n3167) );
  AO22X1_HVT U3247 ( .A1(\ram[12][33] ), .A2(n5380), .A3(n5381), .A4(data[33]), 
        .Y(n3166) );
  AO22X1_HVT U3248 ( .A1(\ram[12][32] ), .A2(n5380), .A3(n5381), .A4(data[32]), 
        .Y(n3165) );
  AO22X1_HVT U3249 ( .A1(\ram[12][31] ), .A2(n5380), .A3(n5381), .A4(data[31]), 
        .Y(n3164) );
  AO22X1_HVT U3250 ( .A1(\ram[12][30] ), .A2(n5380), .A3(n5381), .A4(data[30]), 
        .Y(n3163) );
  AO22X1_HVT U3251 ( .A1(\ram[12][29] ), .A2(n5380), .A3(n5381), .A4(data[29]), 
        .Y(n3162) );
  AO22X1_HVT U3252 ( .A1(\ram[12][28] ), .A2(n5380), .A3(n5381), .A4(data[28]), 
        .Y(n3161) );
  AO22X1_HVT U3253 ( .A1(\ram[12][27] ), .A2(n5380), .A3(n5381), .A4(data[27]), 
        .Y(n3160) );
  AO22X1_HVT U3254 ( .A1(\ram[0][255] ), .A2(n5360), .A3(data[255]), .A4(n5361), .Y(n316) );
  AO22X1_HVT U3255 ( .A1(\ram[12][26] ), .A2(n5380), .A3(n5381), .A4(data[26]), 
        .Y(n3159) );
  AO22X1_HVT U3256 ( .A1(\ram[12][25] ), .A2(n5380), .A3(n5381), .A4(data[25]), 
        .Y(n3158) );
  AO22X1_HVT U3257 ( .A1(\ram[12][24] ), .A2(n5380), .A3(n5381), .A4(data[24]), 
        .Y(n3157) );
  AO22X1_HVT U3258 ( .A1(\ram[12][23] ), .A2(n5380), .A3(n5381), .A4(data[23]), 
        .Y(n3156) );
  AO22X1_HVT U3259 ( .A1(\ram[12][22] ), .A2(n5380), .A3(n5381), .A4(data[22]), 
        .Y(n3155) );
  AO22X1_HVT U3260 ( .A1(\ram[12][21] ), .A2(n5380), .A3(n5381), .A4(data[21]), 
        .Y(n3154) );
  AO22X1_HVT U3261 ( .A1(\ram[12][20] ), .A2(n5380), .A3(n5381), .A4(data[20]), 
        .Y(n3153) );
  AO22X1_HVT U3262 ( .A1(\ram[12][19] ), .A2(n5380), .A3(n5381), .A4(data[19]), 
        .Y(n3152) );
  AO22X1_HVT U3263 ( .A1(\ram[12][18] ), .A2(n5380), .A3(n5381), .A4(data[18]), 
        .Y(n3151) );
  AO22X1_HVT U3264 ( .A1(\ram[12][17] ), .A2(n5380), .A3(n5381), .A4(data[17]), 
        .Y(n3150) );
  AO22X1_HVT U3265 ( .A1(\ram[0][254] ), .A2(n5360), .A3(data[254]), .A4(n5361), .Y(n315) );
  AO22X1_HVT U3266 ( .A1(\ram[12][16] ), .A2(n5380), .A3(n5381), .A4(data[16]), 
        .Y(n3149) );
  AO22X1_HVT U3267 ( .A1(\ram[12][15] ), .A2(n5380), .A3(n5381), .A4(data[15]), 
        .Y(n3148) );
  AO22X1_HVT U3268 ( .A1(\ram[12][14] ), .A2(n5380), .A3(n5381), .A4(data[14]), 
        .Y(n3147) );
  AO22X1_HVT U3269 ( .A1(\ram[12][13] ), .A2(n5380), .A3(n5381), .A4(data[13]), 
        .Y(n3146) );
  AO22X1_HVT U3270 ( .A1(\ram[12][12] ), .A2(n5380), .A3(n5381), .A4(data[12]), 
        .Y(n3145) );
  AO22X1_HVT U3271 ( .A1(\ram[12][11] ), .A2(n5380), .A3(n5381), .A4(data[11]), 
        .Y(n3144) );
  AO22X1_HVT U3272 ( .A1(\ram[12][10] ), .A2(n5380), .A3(n5381), .A4(data[10]), 
        .Y(n3143) );
  AO22X1_HVT U3273 ( .A1(\ram[12][9] ), .A2(n5380), .A3(n5381), .A4(data[9]), 
        .Y(n3142) );
  AO22X1_HVT U3274 ( .A1(\ram[12][8] ), .A2(n5380), .A3(n5381), .A4(data[8]), 
        .Y(n3141) );
  AO22X1_HVT U3275 ( .A1(\ram[12][7] ), .A2(n5380), .A3(n5381), .A4(data[7]), 
        .Y(n3140) );
  AO22X1_HVT U3276 ( .A1(\ram[0][253] ), .A2(n5360), .A3(data[253]), .A4(n5361), .Y(n314) );
  AO22X1_HVT U3277 ( .A1(\ram[12][6] ), .A2(n5380), .A3(n5381), .A4(data[6]), 
        .Y(n3139) );
  AO22X1_HVT U3278 ( .A1(\ram[12][5] ), .A2(n5380), .A3(n5381), .A4(data[5]), 
        .Y(n3138) );
  AO22X1_HVT U3279 ( .A1(\ram[12][4] ), .A2(n5380), .A3(n5381), .A4(data[4]), 
        .Y(n3137) );
  AO22X1_HVT U3280 ( .A1(\ram[12][3] ), .A2(n5380), .A3(n5381), .A4(data[3]), 
        .Y(n3136) );
  AO22X1_HVT U3281 ( .A1(\ram[12][2] ), .A2(n5380), .A3(n5381), .A4(data[2]), 
        .Y(n3135) );
  AO22X1_HVT U3282 ( .A1(\ram[12][1] ), .A2(n5380), .A3(n5381), .A4(data[1]), 
        .Y(n3134) );
  AO22X1_HVT U3283 ( .A1(\ram[12][0] ), .A2(n5380), .A3(n5381), .A4(data[0]), 
        .Y(n3133) );
  INVX0_HVT U3284 ( .A(n5384), .Y(n5381) );
  AND2X1_HVT U3285 ( .A1(n5384), .A2(n5365), .Y(n5380) );
  NAND3X0_HVT U3286 ( .A1(n4183), .A2(n4279), .A3(n5373), .Y(n5384) );
  AND2X1_HVT U3287 ( .A1(N28), .A2(n5385), .Y(n5373) );
  AO22X1_HVT U3288 ( .A1(\ram[11][255] ), .A2(n5386), .A3(n5387), .A4(
        data[255]), .Y(n3132) );
  AO22X1_HVT U3289 ( .A1(\ram[11][254] ), .A2(n5386), .A3(n5387), .A4(
        data[254]), .Y(n3131) );
  AO22X1_HVT U3290 ( .A1(\ram[11][253] ), .A2(n5386), .A3(n5387), .A4(
        data[253]), .Y(n3130) );
  AO22X1_HVT U3291 ( .A1(\ram[0][252] ), .A2(n5360), .A3(data[252]), .A4(n5361), .Y(n313) );
  AO22X1_HVT U3292 ( .A1(\ram[11][252] ), .A2(n5386), .A3(n5387), .A4(
        data[252]), .Y(n3129) );
  AO22X1_HVT U3293 ( .A1(\ram[11][251] ), .A2(n5386), .A3(n5387), .A4(
        data[251]), .Y(n3128) );
  AO22X1_HVT U3294 ( .A1(\ram[11][250] ), .A2(n5386), .A3(n5387), .A4(
        data[250]), .Y(n3127) );
  AO22X1_HVT U3295 ( .A1(\ram[11][249] ), .A2(n5386), .A3(n5387), .A4(
        data[249]), .Y(n3126) );
  AO22X1_HVT U3296 ( .A1(\ram[11][248] ), .A2(n5386), .A3(n5387), .A4(
        data[248]), .Y(n3125) );
  AO22X1_HVT U3297 ( .A1(\ram[11][247] ), .A2(n5386), .A3(n5387), .A4(
        data[247]), .Y(n3124) );
  AO22X1_HVT U3298 ( .A1(\ram[11][246] ), .A2(n5386), .A3(n5387), .A4(
        data[246]), .Y(n3123) );
  AO22X1_HVT U3299 ( .A1(\ram[11][245] ), .A2(n5386), .A3(n5387), .A4(
        data[245]), .Y(n3122) );
  AO22X1_HVT U3300 ( .A1(\ram[11][244] ), .A2(n5386), .A3(n5387), .A4(
        data[244]), .Y(n3121) );
  AO22X1_HVT U3301 ( .A1(\ram[11][243] ), .A2(n5386), .A3(n5387), .A4(
        data[243]), .Y(n3120) );
  AO22X1_HVT U3302 ( .A1(\ram[0][251] ), .A2(n5360), .A3(data[251]), .A4(n5361), .Y(n312) );
  AO22X1_HVT U3303 ( .A1(\ram[11][242] ), .A2(n5386), .A3(n5387), .A4(
        data[242]), .Y(n3119) );
  AO22X1_HVT U3304 ( .A1(\ram[11][241] ), .A2(n5386), .A3(n5387), .A4(
        data[241]), .Y(n3118) );
  AO22X1_HVT U3305 ( .A1(\ram[11][240] ), .A2(n5386), .A3(n5387), .A4(
        data[240]), .Y(n3117) );
  AO22X1_HVT U3306 ( .A1(\ram[11][239] ), .A2(n5386), .A3(n5387), .A4(
        data[239]), .Y(n3116) );
  AO22X1_HVT U3307 ( .A1(\ram[11][238] ), .A2(n5386), .A3(n5387), .A4(
        data[238]), .Y(n3115) );
  AO22X1_HVT U3308 ( .A1(\ram[11][237] ), .A2(n5386), .A3(n5387), .A4(
        data[237]), .Y(n3114) );
  AO22X1_HVT U3309 ( .A1(\ram[11][236] ), .A2(n5386), .A3(n5387), .A4(
        data[236]), .Y(n3113) );
  AO22X1_HVT U3310 ( .A1(\ram[11][235] ), .A2(n5386), .A3(n5387), .A4(
        data[235]), .Y(n3112) );
  AO22X1_HVT U3311 ( .A1(\ram[11][234] ), .A2(n5386), .A3(n5387), .A4(
        data[234]), .Y(n3111) );
  AO22X1_HVT U3312 ( .A1(\ram[11][233] ), .A2(n5386), .A3(n5387), .A4(
        data[233]), .Y(n3110) );
  AO22X1_HVT U3313 ( .A1(\ram[0][250] ), .A2(n5360), .A3(data[250]), .A4(n5361), .Y(n311) );
  AO22X1_HVT U3314 ( .A1(\ram[11][232] ), .A2(n5386), .A3(n5387), .A4(
        data[232]), .Y(n3109) );
  AO22X1_HVT U3315 ( .A1(\ram[11][231] ), .A2(n5386), .A3(n5387), .A4(
        data[231]), .Y(n3108) );
  AO22X1_HVT U3316 ( .A1(\ram[11][230] ), .A2(n5386), .A3(n5387), .A4(
        data[230]), .Y(n3107) );
  AO22X1_HVT U3317 ( .A1(\ram[11][229] ), .A2(n5386), .A3(n5387), .A4(
        data[229]), .Y(n3106) );
  AO22X1_HVT U3318 ( .A1(\ram[11][228] ), .A2(n5386), .A3(n5387), .A4(
        data[228]), .Y(n3105) );
  AO22X1_HVT U3319 ( .A1(\ram[11][227] ), .A2(n5386), .A3(n5387), .A4(
        data[227]), .Y(n3104) );
  AO22X1_HVT U3320 ( .A1(\ram[11][226] ), .A2(n5386), .A3(n5387), .A4(
        data[226]), .Y(n3103) );
  AO22X1_HVT U3321 ( .A1(\ram[11][225] ), .A2(n5386), .A3(n5387), .A4(
        data[225]), .Y(n3102) );
  AO22X1_HVT U3322 ( .A1(\ram[11][224] ), .A2(n5386), .A3(n5387), .A4(
        data[224]), .Y(n3101) );
  AO22X1_HVT U3323 ( .A1(\ram[11][223] ), .A2(n5386), .A3(n5387), .A4(
        data[223]), .Y(n3100) );
  AO22X1_HVT U3324 ( .A1(\ram[0][249] ), .A2(n5360), .A3(data[249]), .A4(n5361), .Y(n310) );
  AO22X1_HVT U3325 ( .A1(\ram[11][222] ), .A2(n5386), .A3(n5387), .A4(
        data[222]), .Y(n3099) );
  AO22X1_HVT U3326 ( .A1(\ram[11][221] ), .A2(n5386), .A3(n5387), .A4(
        data[221]), .Y(n3098) );
  AO22X1_HVT U3327 ( .A1(\ram[11][220] ), .A2(n5386), .A3(n5387), .A4(
        data[220]), .Y(n3097) );
  AO22X1_HVT U3328 ( .A1(\ram[11][219] ), .A2(n5386), .A3(n5387), .A4(
        data[219]), .Y(n3096) );
  AO22X1_HVT U3329 ( .A1(\ram[11][218] ), .A2(n5386), .A3(n5387), .A4(
        data[218]), .Y(n3095) );
  AO22X1_HVT U3330 ( .A1(\ram[11][217] ), .A2(n5386), .A3(n5387), .A4(
        data[217]), .Y(n3094) );
  AO22X1_HVT U3331 ( .A1(\ram[11][216] ), .A2(n5386), .A3(n5387), .A4(
        data[216]), .Y(n3093) );
  AO22X1_HVT U3332 ( .A1(\ram[11][215] ), .A2(n5386), .A3(n5387), .A4(
        data[215]), .Y(n3092) );
  AO22X1_HVT U3333 ( .A1(\ram[11][214] ), .A2(n5386), .A3(n5387), .A4(
        data[214]), .Y(n3091) );
  AO22X1_HVT U3334 ( .A1(\ram[11][213] ), .A2(n5386), .A3(n5387), .A4(
        data[213]), .Y(n3090) );
  AO22X1_HVT U3335 ( .A1(\ram[0][248] ), .A2(n5360), .A3(data[248]), .A4(n5361), .Y(n309) );
  AO22X1_HVT U3336 ( .A1(\ram[11][212] ), .A2(n5386), .A3(n5387), .A4(
        data[212]), .Y(n3089) );
  AO22X1_HVT U3337 ( .A1(\ram[11][211] ), .A2(n5386), .A3(n5387), .A4(
        data[211]), .Y(n3088) );
  AO22X1_HVT U3338 ( .A1(\ram[11][210] ), .A2(n5386), .A3(n5387), .A4(
        data[210]), .Y(n3087) );
  AO22X1_HVT U3339 ( .A1(\ram[11][209] ), .A2(n5386), .A3(n5387), .A4(
        data[209]), .Y(n3086) );
  AO22X1_HVT U3340 ( .A1(\ram[11][208] ), .A2(n5386), .A3(n5387), .A4(
        data[208]), .Y(n3085) );
  AO22X1_HVT U3341 ( .A1(\ram[11][207] ), .A2(n5386), .A3(n5387), .A4(
        data[207]), .Y(n3084) );
  AO22X1_HVT U3342 ( .A1(\ram[11][206] ), .A2(n5386), .A3(n5387), .A4(
        data[206]), .Y(n3083) );
  AO22X1_HVT U3343 ( .A1(\ram[11][205] ), .A2(n5386), .A3(n5387), .A4(
        data[205]), .Y(n3082) );
  AO22X1_HVT U3344 ( .A1(\ram[11][204] ), .A2(n5386), .A3(n5387), .A4(
        data[204]), .Y(n3081) );
  AO22X1_HVT U3345 ( .A1(\ram[11][203] ), .A2(n5386), .A3(n5387), .A4(
        data[203]), .Y(n3080) );
  AO22X1_HVT U3346 ( .A1(\ram[0][247] ), .A2(n5360), .A3(data[247]), .A4(n5361), .Y(n308) );
  AO22X1_HVT U3347 ( .A1(\ram[11][202] ), .A2(n5386), .A3(n5387), .A4(
        data[202]), .Y(n3079) );
  AO22X1_HVT U3348 ( .A1(\ram[11][201] ), .A2(n5386), .A3(n5387), .A4(
        data[201]), .Y(n3078) );
  AO22X1_HVT U3349 ( .A1(\ram[11][200] ), .A2(n5386), .A3(n5387), .A4(
        data[200]), .Y(n3077) );
  AO22X1_HVT U3350 ( .A1(\ram[11][199] ), .A2(n5386), .A3(n5387), .A4(
        data[199]), .Y(n3076) );
  AO22X1_HVT U3351 ( .A1(\ram[11][198] ), .A2(n5386), .A3(n5387), .A4(
        data[198]), .Y(n3075) );
  AO22X1_HVT U3352 ( .A1(\ram[11][197] ), .A2(n5386), .A3(n5387), .A4(
        data[197]), .Y(n3074) );
  AO22X1_HVT U3353 ( .A1(\ram[11][196] ), .A2(n5386), .A3(n5387), .A4(
        data[196]), .Y(n3073) );
  AO22X1_HVT U3354 ( .A1(\ram[11][195] ), .A2(n5386), .A3(n5387), .A4(
        data[195]), .Y(n3072) );
  AO22X1_HVT U3355 ( .A1(\ram[11][194] ), .A2(n5386), .A3(n5387), .A4(
        data[194]), .Y(n3071) );
  AO22X1_HVT U3356 ( .A1(\ram[11][193] ), .A2(n5386), .A3(n5387), .A4(
        data[193]), .Y(n3070) );
  AO22X1_HVT U3357 ( .A1(\ram[0][246] ), .A2(n5360), .A3(data[246]), .A4(n5361), .Y(n307) );
  AO22X1_HVT U3358 ( .A1(\ram[11][192] ), .A2(n5386), .A3(n5387), .A4(
        data[192]), .Y(n3069) );
  AO22X1_HVT U3359 ( .A1(\ram[11][191] ), .A2(n5386), .A3(n5387), .A4(
        data[191]), .Y(n3068) );
  AO22X1_HVT U3360 ( .A1(\ram[11][190] ), .A2(n5386), .A3(n5387), .A4(
        data[190]), .Y(n3067) );
  AO22X1_HVT U3361 ( .A1(\ram[11][189] ), .A2(n5386), .A3(n5387), .A4(
        data[189]), .Y(n3066) );
  AO22X1_HVT U3362 ( .A1(\ram[11][188] ), .A2(n5386), .A3(n5387), .A4(
        data[188]), .Y(n3065) );
  AO22X1_HVT U3363 ( .A1(\ram[11][187] ), .A2(n5386), .A3(n5387), .A4(
        data[187]), .Y(n3064) );
  AO22X1_HVT U3364 ( .A1(\ram[11][186] ), .A2(n5386), .A3(n5387), .A4(
        data[186]), .Y(n3063) );
  AO22X1_HVT U3365 ( .A1(\ram[11][185] ), .A2(n5386), .A3(n5387), .A4(
        data[185]), .Y(n3062) );
  AO22X1_HVT U3366 ( .A1(\ram[11][184] ), .A2(n5386), .A3(n5387), .A4(
        data[184]), .Y(n3061) );
  AO22X1_HVT U3367 ( .A1(\ram[11][183] ), .A2(n5386), .A3(n5387), .A4(
        data[183]), .Y(n3060) );
  AO22X1_HVT U3368 ( .A1(\ram[0][245] ), .A2(n5360), .A3(data[245]), .A4(n5361), .Y(n306) );
  AO22X1_HVT U3369 ( .A1(\ram[11][182] ), .A2(n5386), .A3(n5387), .A4(
        data[182]), .Y(n3059) );
  AO22X1_HVT U3370 ( .A1(\ram[11][181] ), .A2(n5386), .A3(n5387), .A4(
        data[181]), .Y(n3058) );
  AO22X1_HVT U3371 ( .A1(\ram[11][180] ), .A2(n5386), .A3(n5387), .A4(
        data[180]), .Y(n3057) );
  AO22X1_HVT U3372 ( .A1(\ram[11][179] ), .A2(n5386), .A3(n5387), .A4(
        data[179]), .Y(n3056) );
  AO22X1_HVT U3373 ( .A1(\ram[11][178] ), .A2(n5386), .A3(n5387), .A4(
        data[178]), .Y(n3055) );
  AO22X1_HVT U3374 ( .A1(\ram[11][177] ), .A2(n5386), .A3(n5387), .A4(
        data[177]), .Y(n3054) );
  AO22X1_HVT U3375 ( .A1(\ram[11][176] ), .A2(n5386), .A3(n5387), .A4(
        data[176]), .Y(n3053) );
  AO22X1_HVT U3376 ( .A1(\ram[11][175] ), .A2(n5386), .A3(n5387), .A4(
        data[175]), .Y(n3052) );
  AO22X1_HVT U3377 ( .A1(\ram[11][174] ), .A2(n5386), .A3(n5387), .A4(
        data[174]), .Y(n3051) );
  AO22X1_HVT U3378 ( .A1(\ram[11][173] ), .A2(n5386), .A3(n5387), .A4(
        data[173]), .Y(n3050) );
  AO22X1_HVT U3379 ( .A1(\ram[0][244] ), .A2(n5360), .A3(data[244]), .A4(n5361), .Y(n305) );
  AO22X1_HVT U3380 ( .A1(\ram[11][172] ), .A2(n5386), .A3(n5387), .A4(
        data[172]), .Y(n3049) );
  AO22X1_HVT U3381 ( .A1(\ram[11][171] ), .A2(n5386), .A3(n5387), .A4(
        data[171]), .Y(n3048) );
  AO22X1_HVT U3382 ( .A1(\ram[11][170] ), .A2(n5386), .A3(n5387), .A4(
        data[170]), .Y(n3047) );
  AO22X1_HVT U3383 ( .A1(\ram[11][169] ), .A2(n5386), .A3(n5387), .A4(
        data[169]), .Y(n3046) );
  AO22X1_HVT U3384 ( .A1(\ram[11][168] ), .A2(n5386), .A3(n5387), .A4(
        data[168]), .Y(n3045) );
  AO22X1_HVT U3385 ( .A1(\ram[11][167] ), .A2(n5386), .A3(n5387), .A4(
        data[167]), .Y(n3044) );
  AO22X1_HVT U3386 ( .A1(\ram[11][166] ), .A2(n5386), .A3(n5387), .A4(
        data[166]), .Y(n3043) );
  AO22X1_HVT U3387 ( .A1(\ram[11][165] ), .A2(n5386), .A3(n5387), .A4(
        data[165]), .Y(n3042) );
  AO22X1_HVT U3388 ( .A1(\ram[11][164] ), .A2(n5386), .A3(n5387), .A4(
        data[164]), .Y(n3041) );
  AO22X1_HVT U3389 ( .A1(\ram[11][163] ), .A2(n5386), .A3(n5387), .A4(
        data[163]), .Y(n3040) );
  AO22X1_HVT U3390 ( .A1(\ram[0][243] ), .A2(n5360), .A3(data[243]), .A4(n5361), .Y(n304) );
  AO22X1_HVT U3391 ( .A1(\ram[11][162] ), .A2(n5386), .A3(n5387), .A4(
        data[162]), .Y(n3039) );
  AO22X1_HVT U3392 ( .A1(\ram[11][161] ), .A2(n5386), .A3(n5387), .A4(
        data[161]), .Y(n3038) );
  AO22X1_HVT U3393 ( .A1(\ram[11][160] ), .A2(n5386), .A3(n5387), .A4(
        data[160]), .Y(n3037) );
  AO22X1_HVT U3394 ( .A1(\ram[11][159] ), .A2(n5386), .A3(n5387), .A4(
        data[159]), .Y(n3036) );
  AO22X1_HVT U3395 ( .A1(\ram[11][158] ), .A2(n5386), .A3(n5387), .A4(
        data[158]), .Y(n3035) );
  AO22X1_HVT U3396 ( .A1(\ram[11][157] ), .A2(n5386), .A3(n5387), .A4(
        data[157]), .Y(n3034) );
  AO22X1_HVT U3397 ( .A1(\ram[11][156] ), .A2(n5386), .A3(n5387), .A4(
        data[156]), .Y(n3033) );
  AO22X1_HVT U3398 ( .A1(\ram[11][155] ), .A2(n5386), .A3(n5387), .A4(
        data[155]), .Y(n3032) );
  AO22X1_HVT U3399 ( .A1(\ram[11][154] ), .A2(n5386), .A3(n5387), .A4(
        data[154]), .Y(n3031) );
  AO22X1_HVT U3400 ( .A1(\ram[11][153] ), .A2(n5386), .A3(n5387), .A4(
        data[153]), .Y(n3030) );
  AO22X1_HVT U3401 ( .A1(\ram[0][242] ), .A2(n5360), .A3(data[242]), .A4(n5361), .Y(n303) );
  AO22X1_HVT U3402 ( .A1(\ram[11][152] ), .A2(n5386), .A3(n5387), .A4(
        data[152]), .Y(n3029) );
  AO22X1_HVT U3403 ( .A1(\ram[11][151] ), .A2(n5386), .A3(n5387), .A4(
        data[151]), .Y(n3028) );
  AO22X1_HVT U3404 ( .A1(\ram[11][150] ), .A2(n5386), .A3(n5387), .A4(
        data[150]), .Y(n3027) );
  AO22X1_HVT U3405 ( .A1(\ram[11][149] ), .A2(n5386), .A3(n5387), .A4(
        data[149]), .Y(n3026) );
  AO22X1_HVT U3406 ( .A1(\ram[11][148] ), .A2(n5386), .A3(n5387), .A4(
        data[148]), .Y(n3025) );
  AO22X1_HVT U3407 ( .A1(\ram[11][147] ), .A2(n5386), .A3(n5387), .A4(
        data[147]), .Y(n3024) );
  AO22X1_HVT U3408 ( .A1(\ram[11][146] ), .A2(n5386), .A3(n5387), .A4(
        data[146]), .Y(n3023) );
  AO22X1_HVT U3409 ( .A1(\ram[11][145] ), .A2(n5386), .A3(n5387), .A4(
        data[145]), .Y(n3022) );
  AO22X1_HVT U3410 ( .A1(\ram[11][144] ), .A2(n5386), .A3(n5387), .A4(
        data[144]), .Y(n3021) );
  AO22X1_HVT U3411 ( .A1(\ram[11][143] ), .A2(n5386), .A3(n5387), .A4(
        data[143]), .Y(n3020) );
  AO22X1_HVT U3412 ( .A1(\ram[0][241] ), .A2(n5360), .A3(data[241]), .A4(n5361), .Y(n302) );
  AO22X1_HVT U3413 ( .A1(\ram[11][142] ), .A2(n5386), .A3(n5387), .A4(
        data[142]), .Y(n3019) );
  AO22X1_HVT U3414 ( .A1(\ram[11][141] ), .A2(n5386), .A3(n5387), .A4(
        data[141]), .Y(n3018) );
  AO22X1_HVT U3415 ( .A1(\ram[11][140] ), .A2(n5386), .A3(n5387), .A4(
        data[140]), .Y(n3017) );
  AO22X1_HVT U3416 ( .A1(\ram[11][139] ), .A2(n5386), .A3(n5387), .A4(
        data[139]), .Y(n3016) );
  AO22X1_HVT U3417 ( .A1(\ram[11][138] ), .A2(n5386), .A3(n5387), .A4(
        data[138]), .Y(n3015) );
  AO22X1_HVT U3418 ( .A1(\ram[11][137] ), .A2(n5386), .A3(n5387), .A4(
        data[137]), .Y(n3014) );
  AO22X1_HVT U3419 ( .A1(\ram[11][136] ), .A2(n5386), .A3(n5387), .A4(
        data[136]), .Y(n3013) );
  AO22X1_HVT U3420 ( .A1(\ram[11][135] ), .A2(n5386), .A3(n5387), .A4(
        data[135]), .Y(n3012) );
  AO22X1_HVT U3421 ( .A1(\ram[11][134] ), .A2(n5386), .A3(n5387), .A4(
        data[134]), .Y(n3011) );
  AO22X1_HVT U3422 ( .A1(\ram[11][133] ), .A2(n5386), .A3(n5387), .A4(
        data[133]), .Y(n3010) );
  AO22X1_HVT U3423 ( .A1(\ram[0][240] ), .A2(n5360), .A3(data[240]), .A4(n5361), .Y(n301) );
  AO22X1_HVT U3424 ( .A1(\ram[11][132] ), .A2(n5386), .A3(n5387), .A4(
        data[132]), .Y(n3009) );
  AO22X1_HVT U3425 ( .A1(\ram[11][131] ), .A2(n5386), .A3(n5387), .A4(
        data[131]), .Y(n3008) );
  AO22X1_HVT U3426 ( .A1(\ram[11][130] ), .A2(n5386), .A3(n5387), .A4(
        data[130]), .Y(n3007) );
  AO22X1_HVT U3427 ( .A1(\ram[11][129] ), .A2(n5386), .A3(n5387), .A4(
        data[129]), .Y(n3006) );
  AO22X1_HVT U3428 ( .A1(\ram[11][128] ), .A2(n5386), .A3(n5387), .A4(
        data[128]), .Y(n3005) );
  AO22X1_HVT U3429 ( .A1(\ram[11][127] ), .A2(n5386), .A3(n5387), .A4(
        data[127]), .Y(n3004) );
  AO22X1_HVT U3430 ( .A1(\ram[11][126] ), .A2(n5386), .A3(n5387), .A4(
        data[126]), .Y(n3003) );
  AO22X1_HVT U3431 ( .A1(\ram[11][125] ), .A2(n5386), .A3(n5387), .A4(
        data[125]), .Y(n3002) );
  AO22X1_HVT U3432 ( .A1(\ram[11][124] ), .A2(n5386), .A3(n5387), .A4(
        data[124]), .Y(n3001) );
  AO22X1_HVT U3433 ( .A1(\ram[11][123] ), .A2(n5386), .A3(n5387), .A4(
        data[123]), .Y(n3000) );
  AO22X1_HVT U3434 ( .A1(\ram[0][239] ), .A2(n5360), .A3(data[239]), .A4(n5361), .Y(n300) );
  AO22X1_HVT U3435 ( .A1(\ram[11][122] ), .A2(n5386), .A3(n5387), .A4(
        data[122]), .Y(n2999) );
  AO22X1_HVT U3436 ( .A1(\ram[11][121] ), .A2(n5386), .A3(n5387), .A4(
        data[121]), .Y(n2998) );
  AO22X1_HVT U3437 ( .A1(\ram[11][120] ), .A2(n5386), .A3(n5387), .A4(
        data[120]), .Y(n2997) );
  AO22X1_HVT U3438 ( .A1(\ram[11][119] ), .A2(n5386), .A3(n5387), .A4(
        data[119]), .Y(n2996) );
  AO22X1_HVT U3439 ( .A1(\ram[11][118] ), .A2(n5386), .A3(n5387), .A4(
        data[118]), .Y(n2995) );
  AO22X1_HVT U3440 ( .A1(\ram[11][117] ), .A2(n5386), .A3(n5387), .A4(
        data[117]), .Y(n2994) );
  AO22X1_HVT U3441 ( .A1(\ram[11][116] ), .A2(n5386), .A3(n5387), .A4(
        data[116]), .Y(n2993) );
  AO22X1_HVT U3442 ( .A1(\ram[11][115] ), .A2(n5386), .A3(n5387), .A4(
        data[115]), .Y(n2992) );
  AO22X1_HVT U3443 ( .A1(\ram[11][114] ), .A2(n5386), .A3(n5387), .A4(
        data[114]), .Y(n2991) );
  AO22X1_HVT U3444 ( .A1(\ram[11][113] ), .A2(n5386), .A3(n5387), .A4(
        data[113]), .Y(n2990) );
  AO22X1_HVT U3445 ( .A1(\ram[0][238] ), .A2(n5360), .A3(data[238]), .A4(n5361), .Y(n299) );
  AO22X1_HVT U3446 ( .A1(\ram[11][112] ), .A2(n5386), .A3(n5387), .A4(
        data[112]), .Y(n2989) );
  AO22X1_HVT U3447 ( .A1(\ram[11][111] ), .A2(n5386), .A3(n5387), .A4(
        data[111]), .Y(n2988) );
  AO22X1_HVT U3448 ( .A1(\ram[11][110] ), .A2(n5386), .A3(n5387), .A4(
        data[110]), .Y(n2987) );
  AO22X1_HVT U3449 ( .A1(\ram[11][109] ), .A2(n5386), .A3(n5387), .A4(
        data[109]), .Y(n2986) );
  AO22X1_HVT U3450 ( .A1(\ram[11][108] ), .A2(n5386), .A3(n5387), .A4(
        data[108]), .Y(n2985) );
  AO22X1_HVT U3451 ( .A1(\ram[11][107] ), .A2(n5386), .A3(n5387), .A4(
        data[107]), .Y(n2984) );
  AO22X1_HVT U3452 ( .A1(\ram[11][106] ), .A2(n5386), .A3(n5387), .A4(
        data[106]), .Y(n2983) );
  AO22X1_HVT U3453 ( .A1(\ram[11][105] ), .A2(n5386), .A3(n5387), .A4(
        data[105]), .Y(n2982) );
  AO22X1_HVT U3454 ( .A1(\ram[11][104] ), .A2(n5386), .A3(n5387), .A4(
        data[104]), .Y(n2981) );
  AO22X1_HVT U3455 ( .A1(\ram[11][103] ), .A2(n5386), .A3(n5387), .A4(
        data[103]), .Y(n2980) );
  AO22X1_HVT U3456 ( .A1(\ram[0][237] ), .A2(n5360), .A3(data[237]), .A4(n5361), .Y(n298) );
  AO22X1_HVT U3457 ( .A1(\ram[11][102] ), .A2(n5386), .A3(n5387), .A4(
        data[102]), .Y(n2979) );
  AO22X1_HVT U3458 ( .A1(\ram[11][101] ), .A2(n5386), .A3(n5387), .A4(
        data[101]), .Y(n2978) );
  AO22X1_HVT U3459 ( .A1(\ram[11][100] ), .A2(n5386), .A3(n5387), .A4(
        data[100]), .Y(n2977) );
  AO22X1_HVT U3460 ( .A1(\ram[11][99] ), .A2(n5386), .A3(n5387), .A4(data[99]), 
        .Y(n2976) );
  AO22X1_HVT U3461 ( .A1(\ram[11][98] ), .A2(n5386), .A3(n5387), .A4(data[98]), 
        .Y(n2975) );
  AO22X1_HVT U3462 ( .A1(\ram[11][97] ), .A2(n5386), .A3(n5387), .A4(data[97]), 
        .Y(n2974) );
  AO22X1_HVT U3463 ( .A1(\ram[11][96] ), .A2(n5386), .A3(n5387), .A4(data[96]), 
        .Y(n2973) );
  AO22X1_HVT U3464 ( .A1(\ram[11][95] ), .A2(n5386), .A3(n5387), .A4(data[95]), 
        .Y(n2972) );
  AO22X1_HVT U3465 ( .A1(\ram[11][94] ), .A2(n5386), .A3(n5387), .A4(data[94]), 
        .Y(n2971) );
  AO22X1_HVT U3466 ( .A1(\ram[11][93] ), .A2(n5386), .A3(n5387), .A4(data[93]), 
        .Y(n2970) );
  AO22X1_HVT U3467 ( .A1(\ram[0][236] ), .A2(n5360), .A3(data[236]), .A4(n5361), .Y(n297) );
  AO22X1_HVT U3468 ( .A1(\ram[11][92] ), .A2(n5386), .A3(n5387), .A4(data[92]), 
        .Y(n2969) );
  AO22X1_HVT U3469 ( .A1(\ram[11][91] ), .A2(n5386), .A3(n5387), .A4(data[91]), 
        .Y(n2968) );
  AO22X1_HVT U3470 ( .A1(\ram[11][90] ), .A2(n5386), .A3(n5387), .A4(data[90]), 
        .Y(n2967) );
  AO22X1_HVT U3471 ( .A1(\ram[11][89] ), .A2(n5386), .A3(n5387), .A4(data[89]), 
        .Y(n2966) );
  AO22X1_HVT U3472 ( .A1(\ram[11][88] ), .A2(n5386), .A3(n5387), .A4(data[88]), 
        .Y(n2965) );
  AO22X1_HVT U3473 ( .A1(\ram[11][87] ), .A2(n5386), .A3(n5387), .A4(data[87]), 
        .Y(n2964) );
  AO22X1_HVT U3474 ( .A1(\ram[11][86] ), .A2(n5386), .A3(n5387), .A4(data[86]), 
        .Y(n2963) );
  AO22X1_HVT U3475 ( .A1(\ram[11][85] ), .A2(n5386), .A3(n5387), .A4(data[85]), 
        .Y(n2962) );
  AO22X1_HVT U3476 ( .A1(\ram[11][84] ), .A2(n5386), .A3(n5387), .A4(data[84]), 
        .Y(n2961) );
  AO22X1_HVT U3477 ( .A1(\ram[11][83] ), .A2(n5386), .A3(n5387), .A4(data[83]), 
        .Y(n2960) );
  AO22X1_HVT U3478 ( .A1(\ram[0][235] ), .A2(n5360), .A3(data[235]), .A4(n5361), .Y(n296) );
  AO22X1_HVT U3479 ( .A1(\ram[11][82] ), .A2(n5386), .A3(n5387), .A4(data[82]), 
        .Y(n2959) );
  AO22X1_HVT U3480 ( .A1(\ram[11][81] ), .A2(n5386), .A3(n5387), .A4(data[81]), 
        .Y(n2958) );
  AO22X1_HVT U3481 ( .A1(\ram[11][80] ), .A2(n5386), .A3(n5387), .A4(data[80]), 
        .Y(n2957) );
  AO22X1_HVT U3482 ( .A1(\ram[11][79] ), .A2(n5386), .A3(n5387), .A4(data[79]), 
        .Y(n2956) );
  AO22X1_HVT U3483 ( .A1(\ram[11][78] ), .A2(n5386), .A3(n5387), .A4(data[78]), 
        .Y(n2955) );
  AO22X1_HVT U3484 ( .A1(\ram[11][77] ), .A2(n5386), .A3(n5387), .A4(data[77]), 
        .Y(n2954) );
  AO22X1_HVT U3485 ( .A1(\ram[11][76] ), .A2(n5386), .A3(n5387), .A4(data[76]), 
        .Y(n2953) );
  AO22X1_HVT U3486 ( .A1(\ram[11][75] ), .A2(n5386), .A3(n5387), .A4(data[75]), 
        .Y(n2952) );
  AO22X1_HVT U3487 ( .A1(\ram[11][74] ), .A2(n5386), .A3(n5387), .A4(data[74]), 
        .Y(n2951) );
  AO22X1_HVT U3488 ( .A1(\ram[11][73] ), .A2(n5386), .A3(n5387), .A4(data[73]), 
        .Y(n2950) );
  AO22X1_HVT U3489 ( .A1(\ram[0][234] ), .A2(n5360), .A3(data[234]), .A4(n5361), .Y(n295) );
  AO22X1_HVT U3490 ( .A1(\ram[11][72] ), .A2(n5386), .A3(n5387), .A4(data[72]), 
        .Y(n2949) );
  AO22X1_HVT U3491 ( .A1(\ram[11][71] ), .A2(n5386), .A3(n5387), .A4(data[71]), 
        .Y(n2948) );
  AO22X1_HVT U3492 ( .A1(\ram[11][70] ), .A2(n5386), .A3(n5387), .A4(data[70]), 
        .Y(n2947) );
  AO22X1_HVT U3493 ( .A1(\ram[11][69] ), .A2(n5386), .A3(n5387), .A4(data[69]), 
        .Y(n2946) );
  AO22X1_HVT U3494 ( .A1(\ram[11][68] ), .A2(n5386), .A3(n5387), .A4(data[68]), 
        .Y(n2945) );
  AO22X1_HVT U3495 ( .A1(\ram[11][67] ), .A2(n5386), .A3(n5387), .A4(data[67]), 
        .Y(n2944) );
  AO22X1_HVT U3496 ( .A1(\ram[11][66] ), .A2(n5386), .A3(n5387), .A4(data[66]), 
        .Y(n2943) );
  AO22X1_HVT U3497 ( .A1(\ram[11][65] ), .A2(n5386), .A3(n5387), .A4(data[65]), 
        .Y(n2942) );
  AO22X1_HVT U3498 ( .A1(\ram[11][64] ), .A2(n5386), .A3(n5387), .A4(data[64]), 
        .Y(n2941) );
  AO22X1_HVT U3499 ( .A1(\ram[11][63] ), .A2(n5386), .A3(n5387), .A4(data[63]), 
        .Y(n2940) );
  AO22X1_HVT U3500 ( .A1(\ram[0][233] ), .A2(n5360), .A3(data[233]), .A4(n5361), .Y(n294) );
  AO22X1_HVT U3501 ( .A1(\ram[11][62] ), .A2(n5386), .A3(n5387), .A4(data[62]), 
        .Y(n2939) );
  AO22X1_HVT U3502 ( .A1(\ram[11][61] ), .A2(n5386), .A3(n5387), .A4(data[61]), 
        .Y(n2938) );
  AO22X1_HVT U3503 ( .A1(\ram[11][60] ), .A2(n5386), .A3(n5387), .A4(data[60]), 
        .Y(n2937) );
  AO22X1_HVT U3504 ( .A1(\ram[11][59] ), .A2(n5386), .A3(n5387), .A4(data[59]), 
        .Y(n2936) );
  AO22X1_HVT U3505 ( .A1(\ram[11][58] ), .A2(n5386), .A3(n5387), .A4(data[58]), 
        .Y(n2935) );
  AO22X1_HVT U3506 ( .A1(\ram[11][57] ), .A2(n5386), .A3(n5387), .A4(data[57]), 
        .Y(n2934) );
  AO22X1_HVT U3507 ( .A1(\ram[11][56] ), .A2(n5386), .A3(n5387), .A4(data[56]), 
        .Y(n2933) );
  AO22X1_HVT U3508 ( .A1(\ram[11][55] ), .A2(n5386), .A3(n5387), .A4(data[55]), 
        .Y(n2932) );
  AO22X1_HVT U3509 ( .A1(\ram[11][54] ), .A2(n5386), .A3(n5387), .A4(data[54]), 
        .Y(n2931) );
  AO22X1_HVT U3510 ( .A1(\ram[11][53] ), .A2(n5386), .A3(n5387), .A4(data[53]), 
        .Y(n2930) );
  AO22X1_HVT U3511 ( .A1(\ram[0][232] ), .A2(n5360), .A3(data[232]), .A4(n5361), .Y(n293) );
  AO22X1_HVT U3512 ( .A1(\ram[11][52] ), .A2(n5386), .A3(n5387), .A4(data[52]), 
        .Y(n2929) );
  AO22X1_HVT U3513 ( .A1(\ram[11][51] ), .A2(n5386), .A3(n5387), .A4(data[51]), 
        .Y(n2928) );
  AO22X1_HVT U3514 ( .A1(\ram[11][50] ), .A2(n5386), .A3(n5387), .A4(data[50]), 
        .Y(n2927) );
  AO22X1_HVT U3515 ( .A1(\ram[11][49] ), .A2(n5386), .A3(n5387), .A4(data[49]), 
        .Y(n2926) );
  AO22X1_HVT U3516 ( .A1(\ram[11][48] ), .A2(n5386), .A3(n5387), .A4(data[48]), 
        .Y(n2925) );
  AO22X1_HVT U3517 ( .A1(\ram[11][47] ), .A2(n5386), .A3(n5387), .A4(data[47]), 
        .Y(n2924) );
  AO22X1_HVT U3518 ( .A1(\ram[11][46] ), .A2(n5386), .A3(n5387), .A4(data[46]), 
        .Y(n2923) );
  AO22X1_HVT U3519 ( .A1(\ram[11][45] ), .A2(n5386), .A3(n5387), .A4(data[45]), 
        .Y(n2922) );
  AO22X1_HVT U3520 ( .A1(\ram[11][44] ), .A2(n5386), .A3(n5387), .A4(data[44]), 
        .Y(n2921) );
  AO22X1_HVT U3521 ( .A1(\ram[11][43] ), .A2(n5386), .A3(n5387), .A4(data[43]), 
        .Y(n2920) );
  AO22X1_HVT U3522 ( .A1(\ram[0][231] ), .A2(n5360), .A3(data[231]), .A4(n5361), .Y(n292) );
  AO22X1_HVT U3523 ( .A1(\ram[11][42] ), .A2(n5386), .A3(n5387), .A4(data[42]), 
        .Y(n2919) );
  AO22X1_HVT U3524 ( .A1(\ram[11][41] ), .A2(n5386), .A3(n5387), .A4(data[41]), 
        .Y(n2918) );
  AO22X1_HVT U3525 ( .A1(\ram[11][40] ), .A2(n5386), .A3(n5387), .A4(data[40]), 
        .Y(n2917) );
  AO22X1_HVT U3526 ( .A1(\ram[11][39] ), .A2(n5386), .A3(n5387), .A4(data[39]), 
        .Y(n2916) );
  AO22X1_HVT U3527 ( .A1(\ram[11][38] ), .A2(n5386), .A3(n5387), .A4(data[38]), 
        .Y(n2915) );
  AO22X1_HVT U3528 ( .A1(\ram[11][37] ), .A2(n5386), .A3(n5387), .A4(data[37]), 
        .Y(n2914) );
  AO22X1_HVT U3529 ( .A1(\ram[11][36] ), .A2(n5386), .A3(n5387), .A4(data[36]), 
        .Y(n2913) );
  AO22X1_HVT U3530 ( .A1(\ram[11][35] ), .A2(n5386), .A3(n5387), .A4(data[35]), 
        .Y(n2912) );
  AO22X1_HVT U3531 ( .A1(\ram[11][34] ), .A2(n5386), .A3(n5387), .A4(data[34]), 
        .Y(n2911) );
  AO22X1_HVT U3532 ( .A1(\ram[11][33] ), .A2(n5386), .A3(n5387), .A4(data[33]), 
        .Y(n2910) );
  AO22X1_HVT U3533 ( .A1(\ram[0][230] ), .A2(n5360), .A3(data[230]), .A4(n5361), .Y(n291) );
  AO22X1_HVT U3534 ( .A1(\ram[11][32] ), .A2(n5386), .A3(n5387), .A4(data[32]), 
        .Y(n2909) );
  AO22X1_HVT U3535 ( .A1(\ram[11][31] ), .A2(n5386), .A3(n5387), .A4(data[31]), 
        .Y(n2908) );
  AO22X1_HVT U3536 ( .A1(\ram[11][30] ), .A2(n5386), .A3(n5387), .A4(data[30]), 
        .Y(n2907) );
  AO22X1_HVT U3537 ( .A1(\ram[11][29] ), .A2(n5386), .A3(n5387), .A4(data[29]), 
        .Y(n2906) );
  AO22X1_HVT U3538 ( .A1(\ram[11][28] ), .A2(n5386), .A3(n5387), .A4(data[28]), 
        .Y(n2905) );
  AO22X1_HVT U3539 ( .A1(\ram[11][27] ), .A2(n5386), .A3(n5387), .A4(data[27]), 
        .Y(n2904) );
  AO22X1_HVT U3540 ( .A1(\ram[11][26] ), .A2(n5386), .A3(n5387), .A4(data[26]), 
        .Y(n2903) );
  AO22X1_HVT U3541 ( .A1(\ram[11][25] ), .A2(n5386), .A3(n5387), .A4(data[25]), 
        .Y(n2902) );
  AO22X1_HVT U3542 ( .A1(\ram[11][24] ), .A2(n5386), .A3(n5387), .A4(data[24]), 
        .Y(n2901) );
  AO22X1_HVT U3543 ( .A1(\ram[11][23] ), .A2(n5386), .A3(n5387), .A4(data[23]), 
        .Y(n2900) );
  AO22X1_HVT U3544 ( .A1(\ram[0][229] ), .A2(n5360), .A3(data[229]), .A4(n5361), .Y(n290) );
  AO22X1_HVT U3545 ( .A1(\ram[11][22] ), .A2(n5386), .A3(n5387), .A4(data[22]), 
        .Y(n2899) );
  AO22X1_HVT U3546 ( .A1(\ram[11][21] ), .A2(n5386), .A3(n5387), .A4(data[21]), 
        .Y(n2898) );
  AO22X1_HVT U3547 ( .A1(\ram[11][20] ), .A2(n5386), .A3(n5387), .A4(data[20]), 
        .Y(n2897) );
  AO22X1_HVT U3548 ( .A1(\ram[11][19] ), .A2(n5386), .A3(n5387), .A4(data[19]), 
        .Y(n2896) );
  AO22X1_HVT U3549 ( .A1(\ram[11][18] ), .A2(n5386), .A3(n5387), .A4(data[18]), 
        .Y(n2895) );
  AO22X1_HVT U3550 ( .A1(\ram[11][17] ), .A2(n5386), .A3(n5387), .A4(data[17]), 
        .Y(n2894) );
  AO22X1_HVT U3551 ( .A1(\ram[11][16] ), .A2(n5386), .A3(n5387), .A4(data[16]), 
        .Y(n2893) );
  AO22X1_HVT U3552 ( .A1(\ram[11][15] ), .A2(n5386), .A3(n5387), .A4(data[15]), 
        .Y(n2892) );
  AO22X1_HVT U3553 ( .A1(\ram[11][14] ), .A2(n5386), .A3(n5387), .A4(data[14]), 
        .Y(n2891) );
  AO22X1_HVT U3554 ( .A1(\ram[11][13] ), .A2(n5386), .A3(n5387), .A4(data[13]), 
        .Y(n2890) );
  AO22X1_HVT U3555 ( .A1(\ram[0][228] ), .A2(n5360), .A3(data[228]), .A4(n5361), .Y(n289) );
  AO22X1_HVT U3556 ( .A1(\ram[11][12] ), .A2(n5386), .A3(n5387), .A4(data[12]), 
        .Y(n2889) );
  AO22X1_HVT U3557 ( .A1(\ram[11][11] ), .A2(n5386), .A3(n5387), .A4(data[11]), 
        .Y(n2888) );
  AO22X1_HVT U3558 ( .A1(\ram[11][10] ), .A2(n5386), .A3(n5387), .A4(data[10]), 
        .Y(n2887) );
  AO22X1_HVT U3559 ( .A1(\ram[11][9] ), .A2(n5386), .A3(n5387), .A4(data[9]), 
        .Y(n2886) );
  AO22X1_HVT U3560 ( .A1(\ram[11][8] ), .A2(n5386), .A3(n5387), .A4(data[8]), 
        .Y(n2885) );
  AO22X1_HVT U3561 ( .A1(\ram[11][7] ), .A2(n5386), .A3(n5387), .A4(data[7]), 
        .Y(n2884) );
  AO22X1_HVT U3562 ( .A1(\ram[11][6] ), .A2(n5386), .A3(n5387), .A4(data[6]), 
        .Y(n2883) );
  AO22X1_HVT U3563 ( .A1(\ram[11][5] ), .A2(n5386), .A3(n5387), .A4(data[5]), 
        .Y(n2882) );
  AO22X1_HVT U3564 ( .A1(\ram[11][4] ), .A2(n5386), .A3(n5387), .A4(data[4]), 
        .Y(n2881) );
  AO22X1_HVT U3565 ( .A1(\ram[11][3] ), .A2(n5386), .A3(n5387), .A4(data[3]), 
        .Y(n2880) );
  AO22X1_HVT U3566 ( .A1(\ram[0][227] ), .A2(n5360), .A3(data[227]), .A4(n5361), .Y(n288) );
  AO22X1_HVT U3567 ( .A1(\ram[11][2] ), .A2(n5386), .A3(n5387), .A4(data[2]), 
        .Y(n2879) );
  AO22X1_HVT U3568 ( .A1(\ram[11][1] ), .A2(n5386), .A3(n5387), .A4(data[1]), 
        .Y(n2878) );
  AO22X1_HVT U3569 ( .A1(\ram[11][0] ), .A2(n5386), .A3(n5387), .A4(data[0]), 
        .Y(n2877) );
  INVX0_HVT U3570 ( .A(n5388), .Y(n5387) );
  AND2X1_HVT U3571 ( .A1(n5388), .A2(n5365), .Y(n5386) );
  NAND3X0_HVT U3572 ( .A1(n4182), .A2(n5366), .A3(n5385), .Y(n5388) );
  AO22X1_HVT U3573 ( .A1(\ram[10][255] ), .A2(n5389), .A3(n5390), .A4(
        data[255]), .Y(n2876) );
  AO22X1_HVT U3574 ( .A1(\ram[10][254] ), .A2(n5389), .A3(n5390), .A4(
        data[254]), .Y(n2875) );
  AO22X1_HVT U3575 ( .A1(\ram[10][253] ), .A2(n5389), .A3(n5390), .A4(
        data[253]), .Y(n2874) );
  AO22X1_HVT U3576 ( .A1(\ram[10][252] ), .A2(n5389), .A3(n5390), .A4(
        data[252]), .Y(n2873) );
  AO22X1_HVT U3577 ( .A1(\ram[10][251] ), .A2(n5389), .A3(n5390), .A4(
        data[251]), .Y(n2872) );
  AO22X1_HVT U3578 ( .A1(\ram[10][250] ), .A2(n5389), .A3(n5390), .A4(
        data[250]), .Y(n2871) );
  AO22X1_HVT U3579 ( .A1(\ram[10][249] ), .A2(n5389), .A3(n5390), .A4(
        data[249]), .Y(n2870) );
  AO22X1_HVT U3580 ( .A1(\ram[0][226] ), .A2(n5360), .A3(data[226]), .A4(n5361), .Y(n287) );
  AO22X1_HVT U3581 ( .A1(\ram[10][248] ), .A2(n5389), .A3(n5390), .A4(
        data[248]), .Y(n2869) );
  AO22X1_HVT U3582 ( .A1(\ram[10][247] ), .A2(n5389), .A3(n5390), .A4(
        data[247]), .Y(n2868) );
  AO22X1_HVT U3583 ( .A1(\ram[10][246] ), .A2(n5389), .A3(n5390), .A4(
        data[246]), .Y(n2867) );
  AO22X1_HVT U3584 ( .A1(\ram[10][245] ), .A2(n5389), .A3(n5390), .A4(
        data[245]), .Y(n2866) );
  AO22X1_HVT U3585 ( .A1(\ram[10][244] ), .A2(n5389), .A3(n5390), .A4(
        data[244]), .Y(n2865) );
  AO22X1_HVT U3586 ( .A1(\ram[10][243] ), .A2(n5389), .A3(n5390), .A4(
        data[243]), .Y(n2864) );
  AO22X1_HVT U3587 ( .A1(\ram[10][242] ), .A2(n5389), .A3(n5390), .A4(
        data[242]), .Y(n2863) );
  AO22X1_HVT U3588 ( .A1(\ram[10][241] ), .A2(n5389), .A3(n5390), .A4(
        data[241]), .Y(n2862) );
  AO22X1_HVT U3589 ( .A1(\ram[10][240] ), .A2(n5389), .A3(n5390), .A4(
        data[240]), .Y(n2861) );
  AO22X1_HVT U3590 ( .A1(\ram[10][239] ), .A2(n5389), .A3(n5390), .A4(
        data[239]), .Y(n2860) );
  AO22X1_HVT U3591 ( .A1(\ram[0][225] ), .A2(n5360), .A3(data[225]), .A4(n5361), .Y(n286) );
  AO22X1_HVT U3592 ( .A1(\ram[10][238] ), .A2(n5389), .A3(n5390), .A4(
        data[238]), .Y(n2859) );
  AO22X1_HVT U3593 ( .A1(\ram[10][237] ), .A2(n5389), .A3(n5390), .A4(
        data[237]), .Y(n2858) );
  AO22X1_HVT U3594 ( .A1(\ram[10][236] ), .A2(n5389), .A3(n5390), .A4(
        data[236]), .Y(n2857) );
  AO22X1_HVT U3595 ( .A1(\ram[10][235] ), .A2(n5389), .A3(n5390), .A4(
        data[235]), .Y(n2856) );
  AO22X1_HVT U3596 ( .A1(\ram[10][234] ), .A2(n5389), .A3(n5390), .A4(
        data[234]), .Y(n2855) );
  AO22X1_HVT U3597 ( .A1(\ram[10][233] ), .A2(n5389), .A3(n5390), .A4(
        data[233]), .Y(n2854) );
  AO22X1_HVT U3598 ( .A1(\ram[10][232] ), .A2(n5389), .A3(n5390), .A4(
        data[232]), .Y(n2853) );
  AO22X1_HVT U3599 ( .A1(\ram[10][231] ), .A2(n5389), .A3(n5390), .A4(
        data[231]), .Y(n2852) );
  AO22X1_HVT U3600 ( .A1(\ram[10][230] ), .A2(n5389), .A3(n5390), .A4(
        data[230]), .Y(n2851) );
  AO22X1_HVT U3601 ( .A1(\ram[10][229] ), .A2(n5389), .A3(n5390), .A4(
        data[229]), .Y(n2850) );
  AO22X1_HVT U3602 ( .A1(\ram[0][224] ), .A2(n5360), .A3(data[224]), .A4(n5361), .Y(n285) );
  AO22X1_HVT U3603 ( .A1(\ram[10][228] ), .A2(n5389), .A3(n5390), .A4(
        data[228]), .Y(n2849) );
  AO22X1_HVT U3604 ( .A1(\ram[10][227] ), .A2(n5389), .A3(n5390), .A4(
        data[227]), .Y(n2848) );
  AO22X1_HVT U3605 ( .A1(\ram[10][226] ), .A2(n5389), .A3(n5390), .A4(
        data[226]), .Y(n2847) );
  AO22X1_HVT U3606 ( .A1(\ram[10][225] ), .A2(n5389), .A3(n5390), .A4(
        data[225]), .Y(n2846) );
  AO22X1_HVT U3607 ( .A1(\ram[10][224] ), .A2(n5389), .A3(n5390), .A4(
        data[224]), .Y(n2845) );
  AO22X1_HVT U3608 ( .A1(\ram[10][223] ), .A2(n5389), .A3(n5390), .A4(
        data[223]), .Y(n2844) );
  AO22X1_HVT U3609 ( .A1(\ram[10][222] ), .A2(n5389), .A3(n5390), .A4(
        data[222]), .Y(n2843) );
  AO22X1_HVT U3610 ( .A1(\ram[10][221] ), .A2(n5389), .A3(n5390), .A4(
        data[221]), .Y(n2842) );
  AO22X1_HVT U3611 ( .A1(\ram[10][220] ), .A2(n5389), .A3(n5390), .A4(
        data[220]), .Y(n2841) );
  AO22X1_HVT U3612 ( .A1(\ram[10][219] ), .A2(n5389), .A3(n5390), .A4(
        data[219]), .Y(n2840) );
  AO22X1_HVT U3613 ( .A1(\ram[0][223] ), .A2(n5360), .A3(data[223]), .A4(n5361), .Y(n284) );
  AO22X1_HVT U3614 ( .A1(\ram[10][218] ), .A2(n5389), .A3(n5390), .A4(
        data[218]), .Y(n2839) );
  AO22X1_HVT U3615 ( .A1(\ram[10][217] ), .A2(n5389), .A3(n5390), .A4(
        data[217]), .Y(n2838) );
  AO22X1_HVT U3616 ( .A1(\ram[10][216] ), .A2(n5389), .A3(n5390), .A4(
        data[216]), .Y(n2837) );
  AO22X1_HVT U3617 ( .A1(\ram[10][215] ), .A2(n5389), .A3(n5390), .A4(
        data[215]), .Y(n2836) );
  AO22X1_HVT U3618 ( .A1(\ram[10][214] ), .A2(n5389), .A3(n5390), .A4(
        data[214]), .Y(n2835) );
  AO22X1_HVT U3619 ( .A1(\ram[10][213] ), .A2(n5389), .A3(n5390), .A4(
        data[213]), .Y(n2834) );
  AO22X1_HVT U3620 ( .A1(\ram[10][212] ), .A2(n5389), .A3(n5390), .A4(
        data[212]), .Y(n2833) );
  AO22X1_HVT U3621 ( .A1(\ram[10][211] ), .A2(n5389), .A3(n5390), .A4(
        data[211]), .Y(n2832) );
  AO22X1_HVT U3622 ( .A1(\ram[10][210] ), .A2(n5389), .A3(n5390), .A4(
        data[210]), .Y(n2831) );
  AO22X1_HVT U3623 ( .A1(\ram[10][209] ), .A2(n5389), .A3(n5390), .A4(
        data[209]), .Y(n2830) );
  AO22X1_HVT U3624 ( .A1(\ram[0][222] ), .A2(n5360), .A3(data[222]), .A4(n5361), .Y(n283) );
  AO22X1_HVT U3625 ( .A1(\ram[10][208] ), .A2(n5389), .A3(n5390), .A4(
        data[208]), .Y(n2829) );
  AO22X1_HVT U3626 ( .A1(\ram[10][207] ), .A2(n5389), .A3(n5390), .A4(
        data[207]), .Y(n2828) );
  AO22X1_HVT U3627 ( .A1(\ram[10][206] ), .A2(n5389), .A3(n5390), .A4(
        data[206]), .Y(n2827) );
  AO22X1_HVT U3628 ( .A1(\ram[10][205] ), .A2(n5389), .A3(n5390), .A4(
        data[205]), .Y(n2826) );
  AO22X1_HVT U3629 ( .A1(\ram[10][204] ), .A2(n5389), .A3(n5390), .A4(
        data[204]), .Y(n2825) );
  AO22X1_HVT U3630 ( .A1(\ram[10][203] ), .A2(n5389), .A3(n5390), .A4(
        data[203]), .Y(n2824) );
  AO22X1_HVT U3631 ( .A1(\ram[10][202] ), .A2(n5389), .A3(n5390), .A4(
        data[202]), .Y(n2823) );
  AO22X1_HVT U3632 ( .A1(\ram[10][201] ), .A2(n5389), .A3(n5390), .A4(
        data[201]), .Y(n2822) );
  AO22X1_HVT U3633 ( .A1(\ram[10][200] ), .A2(n5389), .A3(n5390), .A4(
        data[200]), .Y(n2821) );
  AO22X1_HVT U3634 ( .A1(\ram[10][199] ), .A2(n5389), .A3(n5390), .A4(
        data[199]), .Y(n2820) );
  AO22X1_HVT U3635 ( .A1(\ram[0][221] ), .A2(n5360), .A3(data[221]), .A4(n5361), .Y(n282) );
  AO22X1_HVT U3636 ( .A1(\ram[10][198] ), .A2(n5389), .A3(n5390), .A4(
        data[198]), .Y(n2819) );
  AO22X1_HVT U3637 ( .A1(\ram[10][197] ), .A2(n5389), .A3(n5390), .A4(
        data[197]), .Y(n2818) );
  AO22X1_HVT U3638 ( .A1(\ram[10][196] ), .A2(n5389), .A3(n5390), .A4(
        data[196]), .Y(n2817) );
  AO22X1_HVT U3639 ( .A1(\ram[10][195] ), .A2(n5389), .A3(n5390), .A4(
        data[195]), .Y(n2816) );
  AO22X1_HVT U3640 ( .A1(\ram[10][194] ), .A2(n5389), .A3(n5390), .A4(
        data[194]), .Y(n2815) );
  AO22X1_HVT U3641 ( .A1(\ram[10][193] ), .A2(n5389), .A3(n5390), .A4(
        data[193]), .Y(n2814) );
  AO22X1_HVT U3642 ( .A1(\ram[10][192] ), .A2(n5389), .A3(n5390), .A4(
        data[192]), .Y(n2813) );
  AO22X1_HVT U3643 ( .A1(\ram[10][191] ), .A2(n5389), .A3(n5390), .A4(
        data[191]), .Y(n2812) );
  AO22X1_HVT U3644 ( .A1(\ram[10][190] ), .A2(n5389), .A3(n5390), .A4(
        data[190]), .Y(n2811) );
  AO22X1_HVT U3645 ( .A1(\ram[10][189] ), .A2(n5389), .A3(n5390), .A4(
        data[189]), .Y(n2810) );
  AO22X1_HVT U3646 ( .A1(\ram[0][220] ), .A2(n5360), .A3(data[220]), .A4(n5361), .Y(n281) );
  AO22X1_HVT U3647 ( .A1(\ram[10][188] ), .A2(n5389), .A3(n5390), .A4(
        data[188]), .Y(n2809) );
  AO22X1_HVT U3648 ( .A1(\ram[10][187] ), .A2(n5389), .A3(n5390), .A4(
        data[187]), .Y(n2808) );
  AO22X1_HVT U3649 ( .A1(\ram[10][186] ), .A2(n5389), .A3(n5390), .A4(
        data[186]), .Y(n2807) );
  AO22X1_HVT U3650 ( .A1(\ram[10][185] ), .A2(n5389), .A3(n5390), .A4(
        data[185]), .Y(n2806) );
  AO22X1_HVT U3651 ( .A1(\ram[10][184] ), .A2(n5389), .A3(n5390), .A4(
        data[184]), .Y(n2805) );
  AO22X1_HVT U3652 ( .A1(\ram[10][183] ), .A2(n5389), .A3(n5390), .A4(
        data[183]), .Y(n2804) );
  AO22X1_HVT U3653 ( .A1(\ram[10][182] ), .A2(n5389), .A3(n5390), .A4(
        data[182]), .Y(n2803) );
  AO22X1_HVT U3654 ( .A1(\ram[10][181] ), .A2(n5389), .A3(n5390), .A4(
        data[181]), .Y(n2802) );
  AO22X1_HVT U3655 ( .A1(\ram[10][180] ), .A2(n5389), .A3(n5390), .A4(
        data[180]), .Y(n2801) );
  AO22X1_HVT U3656 ( .A1(\ram[10][179] ), .A2(n5389), .A3(n5390), .A4(
        data[179]), .Y(n2800) );
  AO22X1_HVT U3657 ( .A1(\ram[0][219] ), .A2(n5360), .A3(data[219]), .A4(n5361), .Y(n280) );
  AO22X1_HVT U3658 ( .A1(\ram[10][178] ), .A2(n5389), .A3(n5390), .A4(
        data[178]), .Y(n2799) );
  AO22X1_HVT U3659 ( .A1(\ram[10][177] ), .A2(n5389), .A3(n5390), .A4(
        data[177]), .Y(n2798) );
  AO22X1_HVT U3660 ( .A1(\ram[10][176] ), .A2(n5389), .A3(n5390), .A4(
        data[176]), .Y(n2797) );
  AO22X1_HVT U3661 ( .A1(\ram[10][175] ), .A2(n5389), .A3(n5390), .A4(
        data[175]), .Y(n2796) );
  AO22X1_HVT U3662 ( .A1(\ram[10][174] ), .A2(n5389), .A3(n5390), .A4(
        data[174]), .Y(n2795) );
  AO22X1_HVT U3663 ( .A1(\ram[10][173] ), .A2(n5389), .A3(n5390), .A4(
        data[173]), .Y(n2794) );
  AO22X1_HVT U3664 ( .A1(\ram[10][172] ), .A2(n5389), .A3(n5390), .A4(
        data[172]), .Y(n2793) );
  AO22X1_HVT U3665 ( .A1(\ram[10][171] ), .A2(n5389), .A3(n5390), .A4(
        data[171]), .Y(n2792) );
  AO22X1_HVT U3666 ( .A1(\ram[10][170] ), .A2(n5389), .A3(n5390), .A4(
        data[170]), .Y(n2791) );
  AO22X1_HVT U3667 ( .A1(\ram[10][169] ), .A2(n5389), .A3(n5390), .A4(
        data[169]), .Y(n2790) );
  AO22X1_HVT U3668 ( .A1(\ram[0][218] ), .A2(n5360), .A3(data[218]), .A4(n5361), .Y(n279) );
  AO22X1_HVT U3669 ( .A1(\ram[10][168] ), .A2(n5389), .A3(n5390), .A4(
        data[168]), .Y(n2789) );
  AO22X1_HVT U3670 ( .A1(\ram[10][167] ), .A2(n5389), .A3(n5390), .A4(
        data[167]), .Y(n2788) );
  AO22X1_HVT U3671 ( .A1(\ram[10][166] ), .A2(n5389), .A3(n5390), .A4(
        data[166]), .Y(n2787) );
  AO22X1_HVT U3672 ( .A1(\ram[10][165] ), .A2(n5389), .A3(n5390), .A4(
        data[165]), .Y(n2786) );
  AO22X1_HVT U3673 ( .A1(\ram[10][164] ), .A2(n5389), .A3(n5390), .A4(
        data[164]), .Y(n2785) );
  AO22X1_HVT U3674 ( .A1(\ram[10][163] ), .A2(n5389), .A3(n5390), .A4(
        data[163]), .Y(n2784) );
  AO22X1_HVT U3675 ( .A1(\ram[10][162] ), .A2(n5389), .A3(n5390), .A4(
        data[162]), .Y(n2783) );
  AO22X1_HVT U3676 ( .A1(\ram[10][161] ), .A2(n5389), .A3(n5390), .A4(
        data[161]), .Y(n2782) );
  AO22X1_HVT U3677 ( .A1(\ram[10][160] ), .A2(n5389), .A3(n5390), .A4(
        data[160]), .Y(n2781) );
  AO22X1_HVT U3678 ( .A1(\ram[10][159] ), .A2(n5389), .A3(n5390), .A4(
        data[159]), .Y(n2780) );
  AO22X1_HVT U3679 ( .A1(\ram[0][217] ), .A2(n5360), .A3(data[217]), .A4(n5361), .Y(n278) );
  AO22X1_HVT U3680 ( .A1(\ram[10][158] ), .A2(n5389), .A3(n5390), .A4(
        data[158]), .Y(n2779) );
  AO22X1_HVT U3681 ( .A1(\ram[10][157] ), .A2(n5389), .A3(n5390), .A4(
        data[157]), .Y(n2778) );
  AO22X1_HVT U3682 ( .A1(\ram[10][156] ), .A2(n5389), .A3(n5390), .A4(
        data[156]), .Y(n2777) );
  AO22X1_HVT U3683 ( .A1(\ram[10][155] ), .A2(n5389), .A3(n5390), .A4(
        data[155]), .Y(n2776) );
  AO22X1_HVT U3684 ( .A1(\ram[10][154] ), .A2(n5389), .A3(n5390), .A4(
        data[154]), .Y(n2775) );
  AO22X1_HVT U3685 ( .A1(\ram[10][153] ), .A2(n5389), .A3(n5390), .A4(
        data[153]), .Y(n2774) );
  AO22X1_HVT U3686 ( .A1(\ram[10][152] ), .A2(n5389), .A3(n5390), .A4(
        data[152]), .Y(n2773) );
  AO22X1_HVT U3687 ( .A1(\ram[10][151] ), .A2(n5389), .A3(n5390), .A4(
        data[151]), .Y(n2772) );
  AO22X1_HVT U3688 ( .A1(\ram[10][150] ), .A2(n5389), .A3(n5390), .A4(
        data[150]), .Y(n2771) );
  AO22X1_HVT U3689 ( .A1(\ram[10][149] ), .A2(n5389), .A3(n5390), .A4(
        data[149]), .Y(n2770) );
  AO22X1_HVT U3690 ( .A1(\ram[0][216] ), .A2(n5360), .A3(data[216]), .A4(n5361), .Y(n277) );
  AO22X1_HVT U3691 ( .A1(\ram[10][148] ), .A2(n5389), .A3(n5390), .A4(
        data[148]), .Y(n2769) );
  AO22X1_HVT U3692 ( .A1(\ram[10][147] ), .A2(n5389), .A3(n5390), .A4(
        data[147]), .Y(n2768) );
  AO22X1_HVT U3693 ( .A1(\ram[10][146] ), .A2(n5389), .A3(n5390), .A4(
        data[146]), .Y(n2767) );
  AO22X1_HVT U3694 ( .A1(\ram[10][145] ), .A2(n5389), .A3(n5390), .A4(
        data[145]), .Y(n2766) );
  AO22X1_HVT U3695 ( .A1(\ram[10][144] ), .A2(n5389), .A3(n5390), .A4(
        data[144]), .Y(n2765) );
  AO22X1_HVT U3696 ( .A1(\ram[10][143] ), .A2(n5389), .A3(n5390), .A4(
        data[143]), .Y(n2764) );
  AO22X1_HVT U3697 ( .A1(\ram[10][142] ), .A2(n5389), .A3(n5390), .A4(
        data[142]), .Y(n2763) );
  AO22X1_HVT U3698 ( .A1(\ram[10][141] ), .A2(n5389), .A3(n5390), .A4(
        data[141]), .Y(n2762) );
  AO22X1_HVT U3699 ( .A1(\ram[10][140] ), .A2(n5389), .A3(n5390), .A4(
        data[140]), .Y(n2761) );
  AO22X1_HVT U3700 ( .A1(\ram[10][139] ), .A2(n5389), .A3(n5390), .A4(
        data[139]), .Y(n2760) );
  AO22X1_HVT U3701 ( .A1(\ram[0][215] ), .A2(n5360), .A3(data[215]), .A4(n5361), .Y(n276) );
  AO22X1_HVT U3702 ( .A1(\ram[10][138] ), .A2(n5389), .A3(n5390), .A4(
        data[138]), .Y(n2759) );
  AO22X1_HVT U3703 ( .A1(\ram[10][137] ), .A2(n5389), .A3(n5390), .A4(
        data[137]), .Y(n2758) );
  AO22X1_HVT U3704 ( .A1(\ram[10][136] ), .A2(n5389), .A3(n5390), .A4(
        data[136]), .Y(n2757) );
  AO22X1_HVT U3705 ( .A1(\ram[10][135] ), .A2(n5389), .A3(n5390), .A4(
        data[135]), .Y(n2756) );
  AO22X1_HVT U3706 ( .A1(\ram[10][134] ), .A2(n5389), .A3(n5390), .A4(
        data[134]), .Y(n2755) );
  AO22X1_HVT U3707 ( .A1(\ram[10][133] ), .A2(n5389), .A3(n5390), .A4(
        data[133]), .Y(n2754) );
  AO22X1_HVT U3708 ( .A1(\ram[10][132] ), .A2(n5389), .A3(n5390), .A4(
        data[132]), .Y(n2753) );
  AO22X1_HVT U3709 ( .A1(\ram[10][131] ), .A2(n5389), .A3(n5390), .A4(
        data[131]), .Y(n2752) );
  AO22X1_HVT U3710 ( .A1(\ram[10][130] ), .A2(n5389), .A3(n5390), .A4(
        data[130]), .Y(n2751) );
  AO22X1_HVT U3711 ( .A1(\ram[10][129] ), .A2(n5389), .A3(n5390), .A4(
        data[129]), .Y(n2750) );
  AO22X1_HVT U3712 ( .A1(\ram[0][214] ), .A2(n5360), .A3(data[214]), .A4(n5361), .Y(n275) );
  AO22X1_HVT U3713 ( .A1(\ram[10][128] ), .A2(n5389), .A3(n5390), .A4(
        data[128]), .Y(n2749) );
  AO22X1_HVT U3714 ( .A1(\ram[10][127] ), .A2(n5389), .A3(n5390), .A4(
        data[127]), .Y(n2748) );
  AO22X1_HVT U3715 ( .A1(\ram[10][126] ), .A2(n5389), .A3(n5390), .A4(
        data[126]), .Y(n2747) );
  AO22X1_HVT U3716 ( .A1(\ram[10][125] ), .A2(n5389), .A3(n5390), .A4(
        data[125]), .Y(n2746) );
  AO22X1_HVT U3717 ( .A1(\ram[10][124] ), .A2(n5389), .A3(n5390), .A4(
        data[124]), .Y(n2745) );
  AO22X1_HVT U3718 ( .A1(\ram[10][123] ), .A2(n5389), .A3(n5390), .A4(
        data[123]), .Y(n2744) );
  AO22X1_HVT U3719 ( .A1(\ram[10][122] ), .A2(n5389), .A3(n5390), .A4(
        data[122]), .Y(n2743) );
  AO22X1_HVT U3720 ( .A1(\ram[10][121] ), .A2(n5389), .A3(n5390), .A4(
        data[121]), .Y(n2742) );
  AO22X1_HVT U3721 ( .A1(\ram[10][120] ), .A2(n5389), .A3(n5390), .A4(
        data[120]), .Y(n2741) );
  AO22X1_HVT U3722 ( .A1(\ram[10][119] ), .A2(n5389), .A3(n5390), .A4(
        data[119]), .Y(n2740) );
  AO22X1_HVT U3723 ( .A1(\ram[0][213] ), .A2(n5360), .A3(data[213]), .A4(n5361), .Y(n274) );
  AO22X1_HVT U3724 ( .A1(\ram[10][118] ), .A2(n5389), .A3(n5390), .A4(
        data[118]), .Y(n2739) );
  AO22X1_HVT U3725 ( .A1(\ram[10][117] ), .A2(n5389), .A3(n5390), .A4(
        data[117]), .Y(n2738) );
  AO22X1_HVT U3726 ( .A1(\ram[10][116] ), .A2(n5389), .A3(n5390), .A4(
        data[116]), .Y(n2737) );
  AO22X1_HVT U3727 ( .A1(\ram[10][115] ), .A2(n5389), .A3(n5390), .A4(
        data[115]), .Y(n2736) );
  AO22X1_HVT U3728 ( .A1(\ram[10][114] ), .A2(n5389), .A3(n5390), .A4(
        data[114]), .Y(n2735) );
  AO22X1_HVT U3729 ( .A1(\ram[10][113] ), .A2(n5389), .A3(n5390), .A4(
        data[113]), .Y(n2734) );
  AO22X1_HVT U3730 ( .A1(\ram[10][112] ), .A2(n5389), .A3(n5390), .A4(
        data[112]), .Y(n2733) );
  AO22X1_HVT U3731 ( .A1(\ram[10][111] ), .A2(n5389), .A3(n5390), .A4(
        data[111]), .Y(n2732) );
  AO22X1_HVT U3732 ( .A1(\ram[10][110] ), .A2(n5389), .A3(n5390), .A4(
        data[110]), .Y(n2731) );
  AO22X1_HVT U3733 ( .A1(\ram[10][109] ), .A2(n5389), .A3(n5390), .A4(
        data[109]), .Y(n2730) );
  AO22X1_HVT U3734 ( .A1(\ram[0][212] ), .A2(n5360), .A3(data[212]), .A4(n5361), .Y(n273) );
  AO22X1_HVT U3735 ( .A1(\ram[10][108] ), .A2(n5389), .A3(n5390), .A4(
        data[108]), .Y(n2729) );
  AO22X1_HVT U3736 ( .A1(\ram[10][107] ), .A2(n5389), .A3(n5390), .A4(
        data[107]), .Y(n2728) );
  AO22X1_HVT U3737 ( .A1(\ram[10][106] ), .A2(n5389), .A3(n5390), .A4(
        data[106]), .Y(n2727) );
  AO22X1_HVT U3738 ( .A1(\ram[10][105] ), .A2(n5389), .A3(n5390), .A4(
        data[105]), .Y(n2726) );
  AO22X1_HVT U3739 ( .A1(\ram[10][104] ), .A2(n5389), .A3(n5390), .A4(
        data[104]), .Y(n2725) );
  AO22X1_HVT U3740 ( .A1(\ram[10][103] ), .A2(n5389), .A3(n5390), .A4(
        data[103]), .Y(n2724) );
  AO22X1_HVT U3741 ( .A1(\ram[10][102] ), .A2(n5389), .A3(n5390), .A4(
        data[102]), .Y(n2723) );
  AO22X1_HVT U3742 ( .A1(\ram[10][101] ), .A2(n5389), .A3(n5390), .A4(
        data[101]), .Y(n2722) );
  AO22X1_HVT U3743 ( .A1(\ram[10][100] ), .A2(n5389), .A3(n5390), .A4(
        data[100]), .Y(n2721) );
  AO22X1_HVT U3744 ( .A1(\ram[10][99] ), .A2(n5389), .A3(n5390), .A4(data[99]), 
        .Y(n2720) );
  AO22X1_HVT U3745 ( .A1(\ram[0][211] ), .A2(n5360), .A3(data[211]), .A4(n5361), .Y(n272) );
  AO22X1_HVT U3746 ( .A1(\ram[10][98] ), .A2(n5389), .A3(n5390), .A4(data[98]), 
        .Y(n2719) );
  AO22X1_HVT U3747 ( .A1(\ram[10][97] ), .A2(n5389), .A3(n5390), .A4(data[97]), 
        .Y(n2718) );
  AO22X1_HVT U3748 ( .A1(\ram[10][96] ), .A2(n5389), .A3(n5390), .A4(data[96]), 
        .Y(n2717) );
  AO22X1_HVT U3749 ( .A1(\ram[10][95] ), .A2(n5389), .A3(n5390), .A4(data[95]), 
        .Y(n2716) );
  AO22X1_HVT U3750 ( .A1(\ram[10][94] ), .A2(n5389), .A3(n5390), .A4(data[94]), 
        .Y(n2715) );
  AO22X1_HVT U3751 ( .A1(\ram[10][93] ), .A2(n5389), .A3(n5390), .A4(data[93]), 
        .Y(n2714) );
  AO22X1_HVT U3752 ( .A1(\ram[10][92] ), .A2(n5389), .A3(n5390), .A4(data[92]), 
        .Y(n2713) );
  AO22X1_HVT U3753 ( .A1(\ram[10][91] ), .A2(n5389), .A3(n5390), .A4(data[91]), 
        .Y(n2712) );
  AO22X1_HVT U3754 ( .A1(\ram[10][90] ), .A2(n5389), .A3(n5390), .A4(data[90]), 
        .Y(n2711) );
  AO22X1_HVT U3755 ( .A1(\ram[10][89] ), .A2(n5389), .A3(n5390), .A4(data[89]), 
        .Y(n2710) );
  AO22X1_HVT U3756 ( .A1(\ram[0][210] ), .A2(n5360), .A3(data[210]), .A4(n5361), .Y(n271) );
  AO22X1_HVT U3757 ( .A1(\ram[10][88] ), .A2(n5389), .A3(n5390), .A4(data[88]), 
        .Y(n2709) );
  AO22X1_HVT U3758 ( .A1(\ram[10][87] ), .A2(n5389), .A3(n5390), .A4(data[87]), 
        .Y(n2708) );
  AO22X1_HVT U3759 ( .A1(\ram[10][86] ), .A2(n5389), .A3(n5390), .A4(data[86]), 
        .Y(n2707) );
  AO22X1_HVT U3760 ( .A1(\ram[10][85] ), .A2(n5389), .A3(n5390), .A4(data[85]), 
        .Y(n2706) );
  AO22X1_HVT U3761 ( .A1(\ram[10][84] ), .A2(n5389), .A3(n5390), .A4(data[84]), 
        .Y(n2705) );
  AO22X1_HVT U3762 ( .A1(\ram[10][83] ), .A2(n5389), .A3(n5390), .A4(data[83]), 
        .Y(n2704) );
  AO22X1_HVT U3763 ( .A1(\ram[10][82] ), .A2(n5389), .A3(n5390), .A4(data[82]), 
        .Y(n2703) );
  AO22X1_HVT U3764 ( .A1(\ram[10][81] ), .A2(n5389), .A3(n5390), .A4(data[81]), 
        .Y(n2702) );
  AO22X1_HVT U3765 ( .A1(\ram[10][80] ), .A2(n5389), .A3(n5390), .A4(data[80]), 
        .Y(n2701) );
  AO22X1_HVT U3766 ( .A1(\ram[10][79] ), .A2(n5389), .A3(n5390), .A4(data[79]), 
        .Y(n2700) );
  AO22X1_HVT U3767 ( .A1(\ram[0][209] ), .A2(n5360), .A3(data[209]), .A4(n5361), .Y(n270) );
  AO22X1_HVT U3768 ( .A1(\ram[10][78] ), .A2(n5389), .A3(n5390), .A4(data[78]), 
        .Y(n2699) );
  AO22X1_HVT U3769 ( .A1(\ram[10][77] ), .A2(n5389), .A3(n5390), .A4(data[77]), 
        .Y(n2698) );
  AO22X1_HVT U3770 ( .A1(\ram[10][76] ), .A2(n5389), .A3(n5390), .A4(data[76]), 
        .Y(n2697) );
  AO22X1_HVT U3771 ( .A1(\ram[10][75] ), .A2(n5389), .A3(n5390), .A4(data[75]), 
        .Y(n2696) );
  AO22X1_HVT U3772 ( .A1(\ram[10][74] ), .A2(n5389), .A3(n5390), .A4(data[74]), 
        .Y(n2695) );
  AO22X1_HVT U3773 ( .A1(\ram[10][73] ), .A2(n5389), .A3(n5390), .A4(data[73]), 
        .Y(n2694) );
  AO22X1_HVT U3774 ( .A1(\ram[10][72] ), .A2(n5389), .A3(n5390), .A4(data[72]), 
        .Y(n2693) );
  AO22X1_HVT U3775 ( .A1(\ram[10][71] ), .A2(n5389), .A3(n5390), .A4(data[71]), 
        .Y(n2692) );
  AO22X1_HVT U3776 ( .A1(\ram[10][70] ), .A2(n5389), .A3(n5390), .A4(data[70]), 
        .Y(n2691) );
  AO22X1_HVT U3777 ( .A1(\ram[10][69] ), .A2(n5389), .A3(n5390), .A4(data[69]), 
        .Y(n2690) );
  AO22X1_HVT U3778 ( .A1(\ram[0][208] ), .A2(n5360), .A3(data[208]), .A4(n5361), .Y(n269) );
  AO22X1_HVT U3779 ( .A1(\ram[10][68] ), .A2(n5389), .A3(n5390), .A4(data[68]), 
        .Y(n2689) );
  AO22X1_HVT U3780 ( .A1(\ram[10][67] ), .A2(n5389), .A3(n5390), .A4(data[67]), 
        .Y(n2688) );
  AO22X1_HVT U3781 ( .A1(\ram[10][66] ), .A2(n5389), .A3(n5390), .A4(data[66]), 
        .Y(n2687) );
  AO22X1_HVT U3782 ( .A1(\ram[10][65] ), .A2(n5389), .A3(n5390), .A4(data[65]), 
        .Y(n2686) );
  AO22X1_HVT U3783 ( .A1(\ram[10][64] ), .A2(n5389), .A3(n5390), .A4(data[64]), 
        .Y(n2685) );
  AO22X1_HVT U3784 ( .A1(\ram[10][63] ), .A2(n5389), .A3(n5390), .A4(data[63]), 
        .Y(n2684) );
  AO22X1_HVT U3785 ( .A1(\ram[10][62] ), .A2(n5389), .A3(n5390), .A4(data[62]), 
        .Y(n2683) );
  AO22X1_HVT U3786 ( .A1(\ram[10][61] ), .A2(n5389), .A3(n5390), .A4(data[61]), 
        .Y(n2682) );
  AO22X1_HVT U3787 ( .A1(\ram[10][60] ), .A2(n5389), .A3(n5390), .A4(data[60]), 
        .Y(n2681) );
  AO22X1_HVT U3788 ( .A1(\ram[10][59] ), .A2(n5389), .A3(n5390), .A4(data[59]), 
        .Y(n2680) );
  AO22X1_HVT U3789 ( .A1(\ram[0][207] ), .A2(n5360), .A3(data[207]), .A4(n5361), .Y(n268) );
  AO22X1_HVT U3790 ( .A1(\ram[10][58] ), .A2(n5389), .A3(n5390), .A4(data[58]), 
        .Y(n2679) );
  AO22X1_HVT U3791 ( .A1(\ram[10][57] ), .A2(n5389), .A3(n5390), .A4(data[57]), 
        .Y(n2678) );
  AO22X1_HVT U3792 ( .A1(\ram[10][56] ), .A2(n5389), .A3(n5390), .A4(data[56]), 
        .Y(n2677) );
  AO22X1_HVT U3793 ( .A1(\ram[10][55] ), .A2(n5389), .A3(n5390), .A4(data[55]), 
        .Y(n2676) );
  AO22X1_HVT U3794 ( .A1(\ram[10][54] ), .A2(n5389), .A3(n5390), .A4(data[54]), 
        .Y(n2675) );
  AO22X1_HVT U3795 ( .A1(\ram[10][53] ), .A2(n5389), .A3(n5390), .A4(data[53]), 
        .Y(n2674) );
  AO22X1_HVT U3796 ( .A1(\ram[10][52] ), .A2(n5389), .A3(n5390), .A4(data[52]), 
        .Y(n2673) );
  AO22X1_HVT U3797 ( .A1(\ram[10][51] ), .A2(n5389), .A3(n5390), .A4(data[51]), 
        .Y(n2672) );
  AO22X1_HVT U3798 ( .A1(\ram[10][50] ), .A2(n5389), .A3(n5390), .A4(data[50]), 
        .Y(n2671) );
  AO22X1_HVT U3799 ( .A1(\ram[10][49] ), .A2(n5389), .A3(n5390), .A4(data[49]), 
        .Y(n2670) );
  AO22X1_HVT U3800 ( .A1(\ram[0][206] ), .A2(n5360), .A3(data[206]), .A4(n5361), .Y(n267) );
  AO22X1_HVT U3801 ( .A1(\ram[10][48] ), .A2(n5389), .A3(n5390), .A4(data[48]), 
        .Y(n2669) );
  AO22X1_HVT U3802 ( .A1(\ram[10][47] ), .A2(n5389), .A3(n5390), .A4(data[47]), 
        .Y(n2668) );
  AO22X1_HVT U3803 ( .A1(\ram[10][46] ), .A2(n5389), .A3(n5390), .A4(data[46]), 
        .Y(n2667) );
  AO22X1_HVT U3804 ( .A1(\ram[10][45] ), .A2(n5389), .A3(n5390), .A4(data[45]), 
        .Y(n2666) );
  AO22X1_HVT U3805 ( .A1(\ram[10][44] ), .A2(n5389), .A3(n5390), .A4(data[44]), 
        .Y(n2665) );
  AO22X1_HVT U3806 ( .A1(\ram[10][43] ), .A2(n5389), .A3(n5390), .A4(data[43]), 
        .Y(n2664) );
  AO22X1_HVT U3807 ( .A1(\ram[10][42] ), .A2(n5389), .A3(n5390), .A4(data[42]), 
        .Y(n2663) );
  AO22X1_HVT U3808 ( .A1(\ram[10][41] ), .A2(n5389), .A3(n5390), .A4(data[41]), 
        .Y(n2662) );
  AO22X1_HVT U3809 ( .A1(\ram[10][40] ), .A2(n5389), .A3(n5390), .A4(data[40]), 
        .Y(n2661) );
  AO22X1_HVT U3810 ( .A1(\ram[10][39] ), .A2(n5389), .A3(n5390), .A4(data[39]), 
        .Y(n2660) );
  AO22X1_HVT U3811 ( .A1(\ram[0][205] ), .A2(n5360), .A3(data[205]), .A4(n5361), .Y(n266) );
  AO22X1_HVT U3812 ( .A1(\ram[10][38] ), .A2(n5389), .A3(n5390), .A4(data[38]), 
        .Y(n2659) );
  AO22X1_HVT U3813 ( .A1(\ram[10][37] ), .A2(n5389), .A3(n5390), .A4(data[37]), 
        .Y(n2658) );
  AO22X1_HVT U3814 ( .A1(\ram[10][36] ), .A2(n5389), .A3(n5390), .A4(data[36]), 
        .Y(n2657) );
  AO22X1_HVT U3815 ( .A1(\ram[10][35] ), .A2(n5389), .A3(n5390), .A4(data[35]), 
        .Y(n2656) );
  AO22X1_HVT U3816 ( .A1(\ram[10][34] ), .A2(n5389), .A3(n5390), .A4(data[34]), 
        .Y(n2655) );
  AO22X1_HVT U3817 ( .A1(\ram[10][33] ), .A2(n5389), .A3(n5390), .A4(data[33]), 
        .Y(n2654) );
  AO22X1_HVT U3818 ( .A1(\ram[10][32] ), .A2(n5389), .A3(n5390), .A4(data[32]), 
        .Y(n2653) );
  AO22X1_HVT U3819 ( .A1(\ram[10][31] ), .A2(n5389), .A3(n5390), .A4(data[31]), 
        .Y(n2652) );
  AO22X1_HVT U3820 ( .A1(\ram[10][30] ), .A2(n5389), .A3(n5390), .A4(data[30]), 
        .Y(n2651) );
  AO22X1_HVT U3821 ( .A1(\ram[10][29] ), .A2(n5389), .A3(n5390), .A4(data[29]), 
        .Y(n2650) );
  AO22X1_HVT U3822 ( .A1(\ram[0][204] ), .A2(n5360), .A3(data[204]), .A4(n5361), .Y(n265) );
  AO22X1_HVT U3823 ( .A1(\ram[10][28] ), .A2(n5389), .A3(n5390), .A4(data[28]), 
        .Y(n2649) );
  AO22X1_HVT U3824 ( .A1(\ram[10][27] ), .A2(n5389), .A3(n5390), .A4(data[27]), 
        .Y(n2648) );
  AO22X1_HVT U3825 ( .A1(\ram[10][26] ), .A2(n5389), .A3(n5390), .A4(data[26]), 
        .Y(n2647) );
  AO22X1_HVT U3826 ( .A1(\ram[10][25] ), .A2(n5389), .A3(n5390), .A4(data[25]), 
        .Y(n2646) );
  AO22X1_HVT U3827 ( .A1(\ram[10][24] ), .A2(n5389), .A3(n5390), .A4(data[24]), 
        .Y(n2645) );
  AO22X1_HVT U3828 ( .A1(\ram[10][23] ), .A2(n5389), .A3(n5390), .A4(data[23]), 
        .Y(n2644) );
  AO22X1_HVT U3829 ( .A1(\ram[10][22] ), .A2(n5389), .A3(n5390), .A4(data[22]), 
        .Y(n2643) );
  AO22X1_HVT U3830 ( .A1(\ram[10][21] ), .A2(n5389), .A3(n5390), .A4(data[21]), 
        .Y(n2642) );
  AO22X1_HVT U3831 ( .A1(\ram[10][20] ), .A2(n5389), .A3(n5390), .A4(data[20]), 
        .Y(n2641) );
  AO22X1_HVT U3832 ( .A1(\ram[10][19] ), .A2(n5389), .A3(n5390), .A4(data[19]), 
        .Y(n2640) );
  AO22X1_HVT U3833 ( .A1(\ram[0][203] ), .A2(n5360), .A3(data[203]), .A4(n5361), .Y(n264) );
  AO22X1_HVT U3834 ( .A1(\ram[10][18] ), .A2(n5389), .A3(n5390), .A4(data[18]), 
        .Y(n2639) );
  AO22X1_HVT U3835 ( .A1(\ram[10][17] ), .A2(n5389), .A3(n5390), .A4(data[17]), 
        .Y(n2638) );
  AO22X1_HVT U3836 ( .A1(\ram[10][16] ), .A2(n5389), .A3(n5390), .A4(data[16]), 
        .Y(n2637) );
  AO22X1_HVT U3837 ( .A1(\ram[10][15] ), .A2(n5389), .A3(n5390), .A4(data[15]), 
        .Y(n2636) );
  AO22X1_HVT U3838 ( .A1(\ram[10][14] ), .A2(n5389), .A3(n5390), .A4(data[14]), 
        .Y(n2635) );
  AO22X1_HVT U3839 ( .A1(\ram[10][13] ), .A2(n5389), .A3(n5390), .A4(data[13]), 
        .Y(n2634) );
  AO22X1_HVT U3840 ( .A1(\ram[10][12] ), .A2(n5389), .A3(n5390), .A4(data[12]), 
        .Y(n2633) );
  AO22X1_HVT U3841 ( .A1(\ram[10][11] ), .A2(n5389), .A3(n5390), .A4(data[11]), 
        .Y(n2632) );
  AO22X1_HVT U3842 ( .A1(\ram[10][10] ), .A2(n5389), .A3(n5390), .A4(data[10]), 
        .Y(n2631) );
  AO22X1_HVT U3843 ( .A1(\ram[10][9] ), .A2(n5389), .A3(n5390), .A4(data[9]), 
        .Y(n2630) );
  AO22X1_HVT U3844 ( .A1(\ram[0][202] ), .A2(n5360), .A3(data[202]), .A4(n5361), .Y(n263) );
  AO22X1_HVT U3845 ( .A1(\ram[10][8] ), .A2(n5389), .A3(n5390), .A4(data[8]), 
        .Y(n2629) );
  AO22X1_HVT U3846 ( .A1(\ram[10][7] ), .A2(n5389), .A3(n5390), .A4(data[7]), 
        .Y(n2628) );
  AO22X1_HVT U3847 ( .A1(\ram[10][6] ), .A2(n5389), .A3(n5390), .A4(data[6]), 
        .Y(n2627) );
  AO22X1_HVT U3848 ( .A1(\ram[10][5] ), .A2(n5389), .A3(n5390), .A4(data[5]), 
        .Y(n2626) );
  AO22X1_HVT U3849 ( .A1(\ram[10][4] ), .A2(n5389), .A3(n5390), .A4(data[4]), 
        .Y(n2625) );
  AO22X1_HVT U3850 ( .A1(\ram[10][3] ), .A2(n5389), .A3(n5390), .A4(data[3]), 
        .Y(n2624) );
  AO22X1_HVT U3851 ( .A1(\ram[10][2] ), .A2(n5389), .A3(n5390), .A4(data[2]), 
        .Y(n2623) );
  AO22X1_HVT U3852 ( .A1(\ram[10][1] ), .A2(n5389), .A3(n5390), .A4(data[1]), 
        .Y(n2622) );
  AO22X1_HVT U3853 ( .A1(\ram[10][0] ), .A2(n5389), .A3(n5390), .A4(data[0]), 
        .Y(n2621) );
  INVX0_HVT U3854 ( .A(n5391), .Y(n5390) );
  AND2X1_HVT U3855 ( .A1(n5391), .A2(n5365), .Y(n5389) );
  NAND3X0_HVT U3856 ( .A1(n5366), .A2(n4183), .A3(n5385), .Y(n5391) );
  AO22X1_HVT U3857 ( .A1(\ram[9][255] ), .A2(n5392), .A3(n5393), .A4(data[255]), .Y(n2620) );
  AO22X1_HVT U3858 ( .A1(\ram[0][201] ), .A2(n5360), .A3(data[201]), .A4(n5361), .Y(n262) );
  AO22X1_HVT U3859 ( .A1(\ram[9][254] ), .A2(n5392), .A3(n5393), .A4(data[254]), .Y(n2619) );
  AO22X1_HVT U3860 ( .A1(\ram[9][253] ), .A2(n5392), .A3(n5393), .A4(data[253]), .Y(n2618) );
  AO22X1_HVT U3861 ( .A1(\ram[9][252] ), .A2(n5392), .A3(n5393), .A4(data[252]), .Y(n2617) );
  AO22X1_HVT U3862 ( .A1(\ram[9][251] ), .A2(n5392), .A3(n5393), .A4(data[251]), .Y(n2616) );
  AO22X1_HVT U3863 ( .A1(\ram[9][250] ), .A2(n5392), .A3(n5393), .A4(data[250]), .Y(n2615) );
  AO22X1_HVT U3864 ( .A1(\ram[9][249] ), .A2(n5392), .A3(n5393), .A4(data[249]), .Y(n2614) );
  AO22X1_HVT U3865 ( .A1(\ram[9][248] ), .A2(n5392), .A3(n5393), .A4(data[248]), .Y(n2613) );
  AO22X1_HVT U3866 ( .A1(\ram[9][247] ), .A2(n5392), .A3(n5393), .A4(data[247]), .Y(n2612) );
  AO22X1_HVT U3867 ( .A1(\ram[9][246] ), .A2(n5392), .A3(n5393), .A4(data[246]), .Y(n2611) );
  AO22X1_HVT U3868 ( .A1(\ram[9][245] ), .A2(n5392), .A3(n5393), .A4(data[245]), .Y(n2610) );
  AO22X1_HVT U3869 ( .A1(\ram[0][200] ), .A2(n5360), .A3(data[200]), .A4(n5361), .Y(n261) );
  AO22X1_HVT U3870 ( .A1(\ram[9][244] ), .A2(n5392), .A3(n5393), .A4(data[244]), .Y(n2609) );
  AO22X1_HVT U3871 ( .A1(\ram[9][243] ), .A2(n5392), .A3(n5393), .A4(data[243]), .Y(n2608) );
  AO22X1_HVT U3872 ( .A1(\ram[9][242] ), .A2(n5392), .A3(n5393), .A4(data[242]), .Y(n2607) );
  AO22X1_HVT U3873 ( .A1(\ram[9][241] ), .A2(n5392), .A3(n5393), .A4(data[241]), .Y(n2606) );
  AO22X1_HVT U3874 ( .A1(\ram[9][240] ), .A2(n5392), .A3(n5393), .A4(data[240]), .Y(n2605) );
  AO22X1_HVT U3875 ( .A1(\ram[9][239] ), .A2(n5392), .A3(n5393), .A4(data[239]), .Y(n2604) );
  AO22X1_HVT U3876 ( .A1(\ram[9][238] ), .A2(n5392), .A3(n5393), .A4(data[238]), .Y(n2603) );
  AO22X1_HVT U3877 ( .A1(\ram[9][237] ), .A2(n5392), .A3(n5393), .A4(data[237]), .Y(n2602) );
  AO22X1_HVT U3878 ( .A1(\ram[9][236] ), .A2(n5392), .A3(n5393), .A4(data[236]), .Y(n2601) );
  AO22X1_HVT U3879 ( .A1(\ram[9][235] ), .A2(n5392), .A3(n5393), .A4(data[235]), .Y(n2600) );
  AO22X1_HVT U3880 ( .A1(\ram[0][199] ), .A2(n5360), .A3(data[199]), .A4(n5361), .Y(n260) );
  AO22X1_HVT U3881 ( .A1(\ram[9][234] ), .A2(n5392), .A3(n5393), .A4(data[234]), .Y(n2599) );
  AO22X1_HVT U3882 ( .A1(\ram[9][233] ), .A2(n5392), .A3(n5393), .A4(data[233]), .Y(n2598) );
  AO22X1_HVT U3883 ( .A1(\ram[9][232] ), .A2(n5392), .A3(n5393), .A4(data[232]), .Y(n2597) );
  AO22X1_HVT U3884 ( .A1(\ram[9][231] ), .A2(n5392), .A3(n5393), .A4(data[231]), .Y(n2596) );
  AO22X1_HVT U3885 ( .A1(\ram[9][230] ), .A2(n5392), .A3(n5393), .A4(data[230]), .Y(n2595) );
  AO22X1_HVT U3886 ( .A1(\ram[9][229] ), .A2(n5392), .A3(n5393), .A4(data[229]), .Y(n2594) );
  AO22X1_HVT U3887 ( .A1(\ram[9][228] ), .A2(n5392), .A3(n5393), .A4(data[228]), .Y(n2593) );
  AO22X1_HVT U3888 ( .A1(\ram[9][227] ), .A2(n5392), .A3(n5393), .A4(data[227]), .Y(n2592) );
  AO22X1_HVT U3889 ( .A1(\ram[9][226] ), .A2(n5392), .A3(n5393), .A4(data[226]), .Y(n2591) );
  AO22X1_HVT U3890 ( .A1(\ram[9][225] ), .A2(n5392), .A3(n5393), .A4(data[225]), .Y(n2590) );
  AO22X1_HVT U3891 ( .A1(\ram[0][198] ), .A2(n5360), .A3(data[198]), .A4(n5361), .Y(n259) );
  AO22X1_HVT U3892 ( .A1(\ram[9][224] ), .A2(n5392), .A3(n5393), .A4(data[224]), .Y(n2589) );
  AO22X1_HVT U3893 ( .A1(\ram[9][223] ), .A2(n5392), .A3(n5393), .A4(data[223]), .Y(n2588) );
  AO22X1_HVT U3894 ( .A1(\ram[9][222] ), .A2(n5392), .A3(n5393), .A4(data[222]), .Y(n2587) );
  AO22X1_HVT U3895 ( .A1(\ram[9][221] ), .A2(n5392), .A3(n5393), .A4(data[221]), .Y(n2586) );
  AO22X1_HVT U3896 ( .A1(\ram[9][220] ), .A2(n5392), .A3(n5393), .A4(data[220]), .Y(n2585) );
  AO22X1_HVT U3897 ( .A1(\ram[9][219] ), .A2(n5392), .A3(n5393), .A4(data[219]), .Y(n2584) );
  AO22X1_HVT U3898 ( .A1(\ram[9][218] ), .A2(n5392), .A3(n5393), .A4(data[218]), .Y(n2583) );
  AO22X1_HVT U3899 ( .A1(\ram[9][217] ), .A2(n5392), .A3(n5393), .A4(data[217]), .Y(n2582) );
  AO22X1_HVT U3900 ( .A1(\ram[9][216] ), .A2(n5392), .A3(n5393), .A4(data[216]), .Y(n2581) );
  AO22X1_HVT U3901 ( .A1(\ram[9][215] ), .A2(n5392), .A3(n5393), .A4(data[215]), .Y(n2580) );
  AO22X1_HVT U3902 ( .A1(\ram[0][197] ), .A2(n5360), .A3(data[197]), .A4(n5361), .Y(n258) );
  AO22X1_HVT U3903 ( .A1(\ram[9][214] ), .A2(n5392), .A3(n5393), .A4(data[214]), .Y(n2579) );
  AO22X1_HVT U3904 ( .A1(\ram[9][213] ), .A2(n5392), .A3(n5393), .A4(data[213]), .Y(n2578) );
  AO22X1_HVT U3905 ( .A1(\ram[9][212] ), .A2(n5392), .A3(n5393), .A4(data[212]), .Y(n2577) );
  AO22X1_HVT U3906 ( .A1(\ram[9][211] ), .A2(n5392), .A3(n5393), .A4(data[211]), .Y(n2576) );
  AO22X1_HVT U3907 ( .A1(\ram[9][210] ), .A2(n5392), .A3(n5393), .A4(data[210]), .Y(n2575) );
  AO22X1_HVT U3908 ( .A1(\ram[9][209] ), .A2(n5392), .A3(n5393), .A4(data[209]), .Y(n2574) );
  AO22X1_HVT U3909 ( .A1(\ram[9][208] ), .A2(n5392), .A3(n5393), .A4(data[208]), .Y(n2573) );
  AO22X1_HVT U3910 ( .A1(\ram[9][207] ), .A2(n5392), .A3(n5393), .A4(data[207]), .Y(n2572) );
  AO22X1_HVT U3911 ( .A1(\ram[9][206] ), .A2(n5392), .A3(n5393), .A4(data[206]), .Y(n2571) );
  AO22X1_HVT U3912 ( .A1(\ram[9][205] ), .A2(n5392), .A3(n5393), .A4(data[205]), .Y(n2570) );
  AO22X1_HVT U3913 ( .A1(\ram[0][196] ), .A2(n5360), .A3(data[196]), .A4(n5361), .Y(n257) );
  AO22X1_HVT U3914 ( .A1(\ram[9][204] ), .A2(n5392), .A3(n5393), .A4(data[204]), .Y(n2569) );
  AO22X1_HVT U3915 ( .A1(\ram[9][203] ), .A2(n5392), .A3(n5393), .A4(data[203]), .Y(n2568) );
  AO22X1_HVT U3916 ( .A1(\ram[9][202] ), .A2(n5392), .A3(n5393), .A4(data[202]), .Y(n2567) );
  AO22X1_HVT U3917 ( .A1(\ram[9][201] ), .A2(n5392), .A3(n5393), .A4(data[201]), .Y(n2566) );
  AO22X1_HVT U3918 ( .A1(\ram[9][200] ), .A2(n5392), .A3(n5393), .A4(data[200]), .Y(n2565) );
  AO22X1_HVT U3919 ( .A1(\ram[9][199] ), .A2(n5392), .A3(n5393), .A4(data[199]), .Y(n2564) );
  AO22X1_HVT U3920 ( .A1(\ram[9][198] ), .A2(n5392), .A3(n5393), .A4(data[198]), .Y(n2563) );
  AO22X1_HVT U3921 ( .A1(\ram[9][197] ), .A2(n5392), .A3(n5393), .A4(data[197]), .Y(n2562) );
  AO22X1_HVT U3922 ( .A1(\ram[9][196] ), .A2(n5392), .A3(n5393), .A4(data[196]), .Y(n2561) );
  AO22X1_HVT U3923 ( .A1(\ram[9][195] ), .A2(n5392), .A3(n5393), .A4(data[195]), .Y(n2560) );
  AO22X1_HVT U3924 ( .A1(\ram[0][195] ), .A2(n5360), .A3(data[195]), .A4(n5361), .Y(n256) );
  AO22X1_HVT U3925 ( .A1(\ram[9][194] ), .A2(n5392), .A3(n5393), .A4(data[194]), .Y(n2559) );
  AO22X1_HVT U3926 ( .A1(\ram[9][193] ), .A2(n5392), .A3(n5393), .A4(data[193]), .Y(n2558) );
  AO22X1_HVT U3927 ( .A1(\ram[9][192] ), .A2(n5392), .A3(n5393), .A4(data[192]), .Y(n2557) );
  AO22X1_HVT U3928 ( .A1(\ram[9][191] ), .A2(n5392), .A3(n5393), .A4(data[191]), .Y(n2556) );
  AO22X1_HVT U3929 ( .A1(\ram[9][190] ), .A2(n5392), .A3(n5393), .A4(data[190]), .Y(n2555) );
  AO22X1_HVT U3930 ( .A1(\ram[9][189] ), .A2(n5392), .A3(n5393), .A4(data[189]), .Y(n2554) );
  AO22X1_HVT U3931 ( .A1(\ram[9][188] ), .A2(n5392), .A3(n5393), .A4(data[188]), .Y(n2553) );
  AO22X1_HVT U3932 ( .A1(\ram[9][187] ), .A2(n5392), .A3(n5393), .A4(data[187]), .Y(n2552) );
  AO22X1_HVT U3933 ( .A1(\ram[9][186] ), .A2(n5392), .A3(n5393), .A4(data[186]), .Y(n2551) );
  AO22X1_HVT U3934 ( .A1(\ram[9][185] ), .A2(n5392), .A3(n5393), .A4(data[185]), .Y(n2550) );
  AO22X1_HVT U3935 ( .A1(\ram[0][194] ), .A2(n5360), .A3(data[194]), .A4(n5361), .Y(n255) );
  AO22X1_HVT U3936 ( .A1(\ram[9][184] ), .A2(n5392), .A3(n5393), .A4(data[184]), .Y(n2549) );
  AO22X1_HVT U3937 ( .A1(\ram[9][183] ), .A2(n5392), .A3(n5393), .A4(data[183]), .Y(n2548) );
  AO22X1_HVT U3938 ( .A1(\ram[9][182] ), .A2(n5392), .A3(n5393), .A4(data[182]), .Y(n2547) );
  AO22X1_HVT U3939 ( .A1(\ram[9][181] ), .A2(n5392), .A3(n5393), .A4(data[181]), .Y(n2546) );
  AO22X1_HVT U3940 ( .A1(\ram[9][180] ), .A2(n5392), .A3(n5393), .A4(data[180]), .Y(n2545) );
  AO22X1_HVT U3941 ( .A1(\ram[9][179] ), .A2(n5392), .A3(n5393), .A4(data[179]), .Y(n2544) );
  AO22X1_HVT U3942 ( .A1(\ram[9][178] ), .A2(n5392), .A3(n5393), .A4(data[178]), .Y(n2543) );
  AO22X1_HVT U3943 ( .A1(\ram[9][177] ), .A2(n5392), .A3(n5393), .A4(data[177]), .Y(n2542) );
  AO22X1_HVT U3944 ( .A1(\ram[9][176] ), .A2(n5392), .A3(n5393), .A4(data[176]), .Y(n2541) );
  AO22X1_HVT U3945 ( .A1(\ram[9][175] ), .A2(n5392), .A3(n5393), .A4(data[175]), .Y(n2540) );
  AO22X1_HVT U3946 ( .A1(\ram[0][193] ), .A2(n5360), .A3(data[193]), .A4(n5361), .Y(n254) );
  AO22X1_HVT U3947 ( .A1(\ram[9][174] ), .A2(n5392), .A3(n5393), .A4(data[174]), .Y(n2539) );
  AO22X1_HVT U3948 ( .A1(\ram[9][173] ), .A2(n5392), .A3(n5393), .A4(data[173]), .Y(n2538) );
  AO22X1_HVT U3949 ( .A1(\ram[9][172] ), .A2(n5392), .A3(n5393), .A4(data[172]), .Y(n2537) );
  AO22X1_HVT U3950 ( .A1(\ram[9][171] ), .A2(n5392), .A3(n5393), .A4(data[171]), .Y(n2536) );
  AO22X1_HVT U3951 ( .A1(\ram[9][170] ), .A2(n5392), .A3(n5393), .A4(data[170]), .Y(n2535) );
  AO22X1_HVT U3952 ( .A1(\ram[9][169] ), .A2(n5392), .A3(n5393), .A4(data[169]), .Y(n2534) );
  AO22X1_HVT U3953 ( .A1(\ram[9][168] ), .A2(n5392), .A3(n5393), .A4(data[168]), .Y(n2533) );
  AO22X1_HVT U3954 ( .A1(\ram[9][167] ), .A2(n5392), .A3(n5393), .A4(data[167]), .Y(n2532) );
  AO22X1_HVT U3955 ( .A1(\ram[9][166] ), .A2(n5392), .A3(n5393), .A4(data[166]), .Y(n2531) );
  AO22X1_HVT U3956 ( .A1(\ram[9][165] ), .A2(n5392), .A3(n5393), .A4(data[165]), .Y(n2530) );
  AO22X1_HVT U3957 ( .A1(\ram[0][192] ), .A2(n5360), .A3(data[192]), .A4(n5361), .Y(n253) );
  AO22X1_HVT U3958 ( .A1(\ram[9][164] ), .A2(n5392), .A3(n5393), .A4(data[164]), .Y(n2529) );
  AO22X1_HVT U3959 ( .A1(\ram[9][163] ), .A2(n5392), .A3(n5393), .A4(data[163]), .Y(n2528) );
  AO22X1_HVT U3960 ( .A1(\ram[9][162] ), .A2(n5392), .A3(n5393), .A4(data[162]), .Y(n2527) );
  AO22X1_HVT U3961 ( .A1(\ram[9][161] ), .A2(n5392), .A3(n5393), .A4(data[161]), .Y(n2526) );
  AO22X1_HVT U3962 ( .A1(\ram[9][160] ), .A2(n5392), .A3(n5393), .A4(data[160]), .Y(n2525) );
  AO22X1_HVT U3963 ( .A1(\ram[9][159] ), .A2(n5392), .A3(n5393), .A4(data[159]), .Y(n2524) );
  AO22X1_HVT U3964 ( .A1(\ram[9][158] ), .A2(n5392), .A3(n5393), .A4(data[158]), .Y(n2523) );
  AO22X1_HVT U3965 ( .A1(\ram[9][157] ), .A2(n5392), .A3(n5393), .A4(data[157]), .Y(n2522) );
  AO22X1_HVT U3966 ( .A1(\ram[9][156] ), .A2(n5392), .A3(n5393), .A4(data[156]), .Y(n2521) );
  AO22X1_HVT U3967 ( .A1(\ram[9][155] ), .A2(n5392), .A3(n5393), .A4(data[155]), .Y(n2520) );
  AO22X1_HVT U3968 ( .A1(\ram[0][191] ), .A2(n5360), .A3(data[191]), .A4(n5361), .Y(n252) );
  AO22X1_HVT U3969 ( .A1(\ram[9][154] ), .A2(n5392), .A3(n5393), .A4(data[154]), .Y(n2519) );
  AO22X1_HVT U3970 ( .A1(\ram[9][153] ), .A2(n5392), .A3(n5393), .A4(data[153]), .Y(n2518) );
  AO22X1_HVT U3971 ( .A1(\ram[9][152] ), .A2(n5392), .A3(n5393), .A4(data[152]), .Y(n2517) );
  AO22X1_HVT U3972 ( .A1(\ram[9][151] ), .A2(n5392), .A3(n5393), .A4(data[151]), .Y(n2516) );
  AO22X1_HVT U3973 ( .A1(\ram[9][150] ), .A2(n5392), .A3(n5393), .A4(data[150]), .Y(n2515) );
  AO22X1_HVT U3974 ( .A1(\ram[9][149] ), .A2(n5392), .A3(n5393), .A4(data[149]), .Y(n2514) );
  AO22X1_HVT U3975 ( .A1(\ram[9][148] ), .A2(n5392), .A3(n5393), .A4(data[148]), .Y(n2513) );
  AO22X1_HVT U3976 ( .A1(\ram[9][147] ), .A2(n5392), .A3(n5393), .A4(data[147]), .Y(n2512) );
  AO22X1_HVT U3977 ( .A1(\ram[9][146] ), .A2(n5392), .A3(n5393), .A4(data[146]), .Y(n2511) );
  AO22X1_HVT U3978 ( .A1(\ram[9][145] ), .A2(n5392), .A3(n5393), .A4(data[145]), .Y(n2510) );
  AO22X1_HVT U3979 ( .A1(\ram[0][190] ), .A2(n5360), .A3(data[190]), .A4(n5361), .Y(n251) );
  AO22X1_HVT U3980 ( .A1(\ram[9][144] ), .A2(n5392), .A3(n5393), .A4(data[144]), .Y(n2509) );
  AO22X1_HVT U3981 ( .A1(\ram[9][143] ), .A2(n5392), .A3(n5393), .A4(data[143]), .Y(n2508) );
  AO22X1_HVT U3982 ( .A1(\ram[9][142] ), .A2(n5392), .A3(n5393), .A4(data[142]), .Y(n2507) );
  AO22X1_HVT U3983 ( .A1(\ram[9][141] ), .A2(n5392), .A3(n5393), .A4(data[141]), .Y(n2506) );
  AO22X1_HVT U3984 ( .A1(\ram[9][140] ), .A2(n5392), .A3(n5393), .A4(data[140]), .Y(n2505) );
  AO22X1_HVT U3985 ( .A1(\ram[9][139] ), .A2(n5392), .A3(n5393), .A4(data[139]), .Y(n2504) );
  AO22X1_HVT U3986 ( .A1(\ram[9][138] ), .A2(n5392), .A3(n5393), .A4(data[138]), .Y(n2503) );
  AO22X1_HVT U3987 ( .A1(\ram[9][137] ), .A2(n5392), .A3(n5393), .A4(data[137]), .Y(n2502) );
  AO22X1_HVT U3988 ( .A1(\ram[9][136] ), .A2(n5392), .A3(n5393), .A4(data[136]), .Y(n2501) );
  AO22X1_HVT U3989 ( .A1(\ram[9][135] ), .A2(n5392), .A3(n5393), .A4(data[135]), .Y(n2500) );
  AO22X1_HVT U3990 ( .A1(\ram[0][189] ), .A2(n5360), .A3(data[189]), .A4(n5361), .Y(n250) );
  AO22X1_HVT U3991 ( .A1(\ram[9][134] ), .A2(n5392), .A3(n5393), .A4(data[134]), .Y(n2499) );
  AO22X1_HVT U3992 ( .A1(\ram[9][133] ), .A2(n5392), .A3(n5393), .A4(data[133]), .Y(n2498) );
  AO22X1_HVT U3993 ( .A1(\ram[9][132] ), .A2(n5392), .A3(n5393), .A4(data[132]), .Y(n2497) );
  AO22X1_HVT U3994 ( .A1(\ram[9][131] ), .A2(n5392), .A3(n5393), .A4(data[131]), .Y(n2496) );
  AO22X1_HVT U3995 ( .A1(\ram[9][130] ), .A2(n5392), .A3(n5393), .A4(data[130]), .Y(n2495) );
  AO22X1_HVT U3996 ( .A1(\ram[9][129] ), .A2(n5392), .A3(n5393), .A4(data[129]), .Y(n2494) );
  AO22X1_HVT U3997 ( .A1(\ram[9][128] ), .A2(n5392), .A3(n5393), .A4(data[128]), .Y(n2493) );
  AO22X1_HVT U3998 ( .A1(\ram[9][127] ), .A2(n5392), .A3(n5393), .A4(data[127]), .Y(n2492) );
  AO22X1_HVT U3999 ( .A1(\ram[9][126] ), .A2(n5392), .A3(n5393), .A4(data[126]), .Y(n2491) );
  AO22X1_HVT U4000 ( .A1(\ram[9][125] ), .A2(n5392), .A3(n5393), .A4(data[125]), .Y(n2490) );
  AO22X1_HVT U4001 ( .A1(\ram[0][188] ), .A2(n5360), .A3(data[188]), .A4(n5361), .Y(n249) );
  AO22X1_HVT U4002 ( .A1(\ram[9][124] ), .A2(n5392), .A3(n5393), .A4(data[124]), .Y(n2489) );
  AO22X1_HVT U4003 ( .A1(\ram[9][123] ), .A2(n5392), .A3(n5393), .A4(data[123]), .Y(n2488) );
  AO22X1_HVT U4004 ( .A1(\ram[9][122] ), .A2(n5392), .A3(n5393), .A4(data[122]), .Y(n2487) );
  AO22X1_HVT U4005 ( .A1(\ram[9][121] ), .A2(n5392), .A3(n5393), .A4(data[121]), .Y(n2486) );
  AO22X1_HVT U4006 ( .A1(\ram[9][120] ), .A2(n5392), .A3(n5393), .A4(data[120]), .Y(n2485) );
  AO22X1_HVT U4007 ( .A1(\ram[9][119] ), .A2(n5392), .A3(n5393), .A4(data[119]), .Y(n2484) );
  AO22X1_HVT U4008 ( .A1(\ram[9][118] ), .A2(n5392), .A3(n5393), .A4(data[118]), .Y(n2483) );
  AO22X1_HVT U4009 ( .A1(\ram[9][117] ), .A2(n5392), .A3(n5393), .A4(data[117]), .Y(n2482) );
  AO22X1_HVT U4010 ( .A1(\ram[9][116] ), .A2(n5392), .A3(n5393), .A4(data[116]), .Y(n2481) );
  AO22X1_HVT U4011 ( .A1(\ram[9][115] ), .A2(n5392), .A3(n5393), .A4(data[115]), .Y(n2480) );
  AO22X1_HVT U4012 ( .A1(\ram[0][187] ), .A2(n5360), .A3(data[187]), .A4(n5361), .Y(n248) );
  AO22X1_HVT U4013 ( .A1(\ram[9][114] ), .A2(n5392), .A3(n5393), .A4(data[114]), .Y(n2479) );
  AO22X1_HVT U4014 ( .A1(\ram[9][113] ), .A2(n5392), .A3(n5393), .A4(data[113]), .Y(n2478) );
  AO22X1_HVT U4015 ( .A1(\ram[9][112] ), .A2(n5392), .A3(n5393), .A4(data[112]), .Y(n2477) );
  AO22X1_HVT U4016 ( .A1(\ram[9][111] ), .A2(n5392), .A3(n5393), .A4(data[111]), .Y(n2476) );
  AO22X1_HVT U4017 ( .A1(\ram[9][110] ), .A2(n5392), .A3(n5393), .A4(data[110]), .Y(n2475) );
  AO22X1_HVT U4018 ( .A1(\ram[9][109] ), .A2(n5392), .A3(n5393), .A4(data[109]), .Y(n2474) );
  AO22X1_HVT U4019 ( .A1(\ram[9][108] ), .A2(n5392), .A3(n5393), .A4(data[108]), .Y(n2473) );
  AO22X1_HVT U4020 ( .A1(\ram[9][107] ), .A2(n5392), .A3(n5393), .A4(data[107]), .Y(n2472) );
  AO22X1_HVT U4021 ( .A1(\ram[9][106] ), .A2(n5392), .A3(n5393), .A4(data[106]), .Y(n2471) );
  AO22X1_HVT U4022 ( .A1(\ram[9][105] ), .A2(n5392), .A3(n5393), .A4(data[105]), .Y(n2470) );
  AO22X1_HVT U4023 ( .A1(\ram[0][186] ), .A2(n5360), .A3(data[186]), .A4(n5361), .Y(n247) );
  AO22X1_HVT U4024 ( .A1(\ram[9][104] ), .A2(n5392), .A3(n5393), .A4(data[104]), .Y(n2469) );
  AO22X1_HVT U4025 ( .A1(\ram[9][103] ), .A2(n5392), .A3(n5393), .A4(data[103]), .Y(n2468) );
  AO22X1_HVT U4026 ( .A1(\ram[9][102] ), .A2(n5392), .A3(n5393), .A4(data[102]), .Y(n2467) );
  AO22X1_HVT U4027 ( .A1(\ram[9][101] ), .A2(n5392), .A3(n5393), .A4(data[101]), .Y(n2466) );
  AO22X1_HVT U4028 ( .A1(\ram[9][100] ), .A2(n5392), .A3(n5393), .A4(data[100]), .Y(n2465) );
  AO22X1_HVT U4029 ( .A1(\ram[9][99] ), .A2(n5392), .A3(n5393), .A4(data[99]), 
        .Y(n2464) );
  AO22X1_HVT U4030 ( .A1(\ram[9][98] ), .A2(n5392), .A3(n5393), .A4(data[98]), 
        .Y(n2463) );
  AO22X1_HVT U4031 ( .A1(\ram[9][97] ), .A2(n5392), .A3(n5393), .A4(data[97]), 
        .Y(n2462) );
  AO22X1_HVT U4032 ( .A1(\ram[9][96] ), .A2(n5392), .A3(n5393), .A4(data[96]), 
        .Y(n2461) );
  AO22X1_HVT U4033 ( .A1(\ram[9][95] ), .A2(n5392), .A3(n5393), .A4(data[95]), 
        .Y(n2460) );
  AO22X1_HVT U4034 ( .A1(\ram[0][185] ), .A2(n5360), .A3(data[185]), .A4(n5361), .Y(n246) );
  AO22X1_HVT U4035 ( .A1(\ram[9][94] ), .A2(n5392), .A3(n5393), .A4(data[94]), 
        .Y(n2459) );
  AO22X1_HVT U4036 ( .A1(\ram[9][93] ), .A2(n5392), .A3(n5393), .A4(data[93]), 
        .Y(n2458) );
  AO22X1_HVT U4037 ( .A1(\ram[9][92] ), .A2(n5392), .A3(n5393), .A4(data[92]), 
        .Y(n2457) );
  AO22X1_HVT U4038 ( .A1(\ram[9][91] ), .A2(n5392), .A3(n5393), .A4(data[91]), 
        .Y(n2456) );
  AO22X1_HVT U4039 ( .A1(\ram[9][90] ), .A2(n5392), .A3(n5393), .A4(data[90]), 
        .Y(n2455) );
  AO22X1_HVT U4040 ( .A1(\ram[9][89] ), .A2(n5392), .A3(n5393), .A4(data[89]), 
        .Y(n2454) );
  AO22X1_HVT U4041 ( .A1(\ram[9][88] ), .A2(n5392), .A3(n5393), .A4(data[88]), 
        .Y(n2453) );
  AO22X1_HVT U4042 ( .A1(\ram[9][87] ), .A2(n5392), .A3(n5393), .A4(data[87]), 
        .Y(n2452) );
  AO22X1_HVT U4043 ( .A1(\ram[9][86] ), .A2(n5392), .A3(n5393), .A4(data[86]), 
        .Y(n2451) );
  AO22X1_HVT U4044 ( .A1(\ram[9][85] ), .A2(n5392), .A3(n5393), .A4(data[85]), 
        .Y(n2450) );
  AO22X1_HVT U4045 ( .A1(\ram[0][184] ), .A2(n5360), .A3(data[184]), .A4(n5361), .Y(n245) );
  AO22X1_HVT U4046 ( .A1(\ram[9][84] ), .A2(n5392), .A3(n5393), .A4(data[84]), 
        .Y(n2449) );
  AO22X1_HVT U4047 ( .A1(\ram[9][83] ), .A2(n5392), .A3(n5393), .A4(data[83]), 
        .Y(n2448) );
  AO22X1_HVT U4048 ( .A1(\ram[9][82] ), .A2(n5392), .A3(n5393), .A4(data[82]), 
        .Y(n2447) );
  AO22X1_HVT U4049 ( .A1(\ram[9][81] ), .A2(n5392), .A3(n5393), .A4(data[81]), 
        .Y(n2446) );
  AO22X1_HVT U4050 ( .A1(\ram[9][80] ), .A2(n5392), .A3(n5393), .A4(data[80]), 
        .Y(n2445) );
  AO22X1_HVT U4051 ( .A1(\ram[9][79] ), .A2(n5392), .A3(n5393), .A4(data[79]), 
        .Y(n2444) );
  AO22X1_HVT U4052 ( .A1(\ram[9][78] ), .A2(n5392), .A3(n5393), .A4(data[78]), 
        .Y(n2443) );
  AO22X1_HVT U4053 ( .A1(\ram[9][77] ), .A2(n5392), .A3(n5393), .A4(data[77]), 
        .Y(n2442) );
  AO22X1_HVT U4054 ( .A1(\ram[9][76] ), .A2(n5392), .A3(n5393), .A4(data[76]), 
        .Y(n2441) );
  AO22X1_HVT U4055 ( .A1(\ram[9][75] ), .A2(n5392), .A3(n5393), .A4(data[75]), 
        .Y(n2440) );
  AO22X1_HVT U4056 ( .A1(\ram[0][183] ), .A2(n5360), .A3(data[183]), .A4(n5361), .Y(n244) );
  AO22X1_HVT U4057 ( .A1(\ram[9][74] ), .A2(n5392), .A3(n5393), .A4(data[74]), 
        .Y(n2439) );
  AO22X1_HVT U4058 ( .A1(\ram[9][73] ), .A2(n5392), .A3(n5393), .A4(data[73]), 
        .Y(n2438) );
  AO22X1_HVT U4059 ( .A1(\ram[9][72] ), .A2(n5392), .A3(n5393), .A4(data[72]), 
        .Y(n2437) );
  AO22X1_HVT U4060 ( .A1(\ram[9][71] ), .A2(n5392), .A3(n5393), .A4(data[71]), 
        .Y(n2436) );
  AO22X1_HVT U4061 ( .A1(\ram[9][70] ), .A2(n5392), .A3(n5393), .A4(data[70]), 
        .Y(n2435) );
  AO22X1_HVT U4062 ( .A1(\ram[9][69] ), .A2(n5392), .A3(n5393), .A4(data[69]), 
        .Y(n2434) );
  AO22X1_HVT U4063 ( .A1(\ram[9][68] ), .A2(n5392), .A3(n5393), .A4(data[68]), 
        .Y(n2433) );
  AO22X1_HVT U4064 ( .A1(\ram[9][67] ), .A2(n5392), .A3(n5393), .A4(data[67]), 
        .Y(n2432) );
  AO22X1_HVT U4065 ( .A1(\ram[9][66] ), .A2(n5392), .A3(n5393), .A4(data[66]), 
        .Y(n2431) );
  AO22X1_HVT U4066 ( .A1(\ram[9][65] ), .A2(n5392), .A3(n5393), .A4(data[65]), 
        .Y(n2430) );
  AO22X1_HVT U4067 ( .A1(\ram[0][182] ), .A2(n5360), .A3(data[182]), .A4(n5361), .Y(n243) );
  AO22X1_HVT U4068 ( .A1(\ram[9][64] ), .A2(n5392), .A3(n5393), .A4(data[64]), 
        .Y(n2429) );
  AO22X1_HVT U4069 ( .A1(\ram[9][63] ), .A2(n5392), .A3(n5393), .A4(data[63]), 
        .Y(n2428) );
  AO22X1_HVT U4070 ( .A1(\ram[9][62] ), .A2(n5392), .A3(n5393), .A4(data[62]), 
        .Y(n2427) );
  AO22X1_HVT U4071 ( .A1(\ram[9][61] ), .A2(n5392), .A3(n5393), .A4(data[61]), 
        .Y(n2426) );
  AO22X1_HVT U4072 ( .A1(\ram[9][60] ), .A2(n5392), .A3(n5393), .A4(data[60]), 
        .Y(n2425) );
  AO22X1_HVT U4073 ( .A1(\ram[9][59] ), .A2(n5392), .A3(n5393), .A4(data[59]), 
        .Y(n2424) );
  AO22X1_HVT U4074 ( .A1(\ram[9][58] ), .A2(n5392), .A3(n5393), .A4(data[58]), 
        .Y(n2423) );
  AO22X1_HVT U4075 ( .A1(\ram[9][57] ), .A2(n5392), .A3(n5393), .A4(data[57]), 
        .Y(n2422) );
  AO22X1_HVT U4076 ( .A1(\ram[9][56] ), .A2(n5392), .A3(n5393), .A4(data[56]), 
        .Y(n2421) );
  AO22X1_HVT U4077 ( .A1(\ram[9][55] ), .A2(n5392), .A3(n5393), .A4(data[55]), 
        .Y(n2420) );
  AO22X1_HVT U4078 ( .A1(\ram[0][181] ), .A2(n5360), .A3(data[181]), .A4(n5361), .Y(n242) );
  AO22X1_HVT U4079 ( .A1(\ram[9][54] ), .A2(n5392), .A3(n5393), .A4(data[54]), 
        .Y(n2419) );
  AO22X1_HVT U4080 ( .A1(\ram[9][53] ), .A2(n5392), .A3(n5393), .A4(data[53]), 
        .Y(n2418) );
  AO22X1_HVT U4081 ( .A1(\ram[9][52] ), .A2(n5392), .A3(n5393), .A4(data[52]), 
        .Y(n2417) );
  AO22X1_HVT U4082 ( .A1(\ram[9][51] ), .A2(n5392), .A3(n5393), .A4(data[51]), 
        .Y(n2416) );
  AO22X1_HVT U4083 ( .A1(\ram[9][50] ), .A2(n5392), .A3(n5393), .A4(data[50]), 
        .Y(n2415) );
  AO22X1_HVT U4084 ( .A1(\ram[9][49] ), .A2(n5392), .A3(n5393), .A4(data[49]), 
        .Y(n2414) );
  AO22X1_HVT U4085 ( .A1(\ram[9][48] ), .A2(n5392), .A3(n5393), .A4(data[48]), 
        .Y(n2413) );
  AO22X1_HVT U4086 ( .A1(\ram[9][47] ), .A2(n5392), .A3(n5393), .A4(data[47]), 
        .Y(n2412) );
  AO22X1_HVT U4087 ( .A1(\ram[9][46] ), .A2(n5392), .A3(n5393), .A4(data[46]), 
        .Y(n2411) );
  AO22X1_HVT U4088 ( .A1(\ram[9][45] ), .A2(n5392), .A3(n5393), .A4(data[45]), 
        .Y(n2410) );
  AO22X1_HVT U4089 ( .A1(\ram[0][180] ), .A2(n5360), .A3(data[180]), .A4(n5361), .Y(n241) );
  AO22X1_HVT U4090 ( .A1(\ram[9][44] ), .A2(n5392), .A3(n5393), .A4(data[44]), 
        .Y(n2409) );
  AO22X1_HVT U4091 ( .A1(\ram[9][43] ), .A2(n5392), .A3(n5393), .A4(data[43]), 
        .Y(n2408) );
  AO22X1_HVT U4092 ( .A1(\ram[9][42] ), .A2(n5392), .A3(n5393), .A4(data[42]), 
        .Y(n2407) );
  AO22X1_HVT U4093 ( .A1(\ram[9][41] ), .A2(n5392), .A3(n5393), .A4(data[41]), 
        .Y(n2406) );
  AO22X1_HVT U4094 ( .A1(\ram[9][40] ), .A2(n5392), .A3(n5393), .A4(data[40]), 
        .Y(n2405) );
  AO22X1_HVT U4095 ( .A1(\ram[9][39] ), .A2(n5392), .A3(n5393), .A4(data[39]), 
        .Y(n2404) );
  AO22X1_HVT U4096 ( .A1(\ram[9][38] ), .A2(n5392), .A3(n5393), .A4(data[38]), 
        .Y(n2403) );
  AO22X1_HVT U4097 ( .A1(\ram[9][37] ), .A2(n5392), .A3(n5393), .A4(data[37]), 
        .Y(n2402) );
  AO22X1_HVT U4098 ( .A1(\ram[9][36] ), .A2(n5392), .A3(n5393), .A4(data[36]), 
        .Y(n2401) );
  AO22X1_HVT U4099 ( .A1(\ram[9][35] ), .A2(n5392), .A3(n5393), .A4(data[35]), 
        .Y(n2400) );
  AO22X1_HVT U4100 ( .A1(\ram[0][179] ), .A2(n5360), .A3(data[179]), .A4(n5361), .Y(n240) );
  AO22X1_HVT U4101 ( .A1(\ram[9][34] ), .A2(n5392), .A3(n5393), .A4(data[34]), 
        .Y(n2399) );
  AO22X1_HVT U4102 ( .A1(\ram[9][33] ), .A2(n5392), .A3(n5393), .A4(data[33]), 
        .Y(n2398) );
  AO22X1_HVT U4103 ( .A1(\ram[9][32] ), .A2(n5392), .A3(n5393), .A4(data[32]), 
        .Y(n2397) );
  AO22X1_HVT U4104 ( .A1(\ram[9][31] ), .A2(n5392), .A3(n5393), .A4(data[31]), 
        .Y(n2396) );
  AO22X1_HVT U4105 ( .A1(\ram[9][30] ), .A2(n5392), .A3(n5393), .A4(data[30]), 
        .Y(n2395) );
  AO22X1_HVT U4106 ( .A1(\ram[9][29] ), .A2(n5392), .A3(n5393), .A4(data[29]), 
        .Y(n2394) );
  AO22X1_HVT U4107 ( .A1(\ram[9][28] ), .A2(n5392), .A3(n5393), .A4(data[28]), 
        .Y(n2393) );
  AO22X1_HVT U4108 ( .A1(\ram[9][27] ), .A2(n5392), .A3(n5393), .A4(data[27]), 
        .Y(n2392) );
  AO22X1_HVT U4109 ( .A1(\ram[9][26] ), .A2(n5392), .A3(n5393), .A4(data[26]), 
        .Y(n2391) );
  AO22X1_HVT U4110 ( .A1(\ram[9][25] ), .A2(n5392), .A3(n5393), .A4(data[25]), 
        .Y(n2390) );
  AO22X1_HVT U4111 ( .A1(\ram[0][178] ), .A2(n5360), .A3(data[178]), .A4(n5361), .Y(n239) );
  AO22X1_HVT U4112 ( .A1(\ram[9][24] ), .A2(n5392), .A3(n5393), .A4(data[24]), 
        .Y(n2389) );
  AO22X1_HVT U4113 ( .A1(\ram[9][23] ), .A2(n5392), .A3(n5393), .A4(data[23]), 
        .Y(n2388) );
  AO22X1_HVT U4114 ( .A1(\ram[9][22] ), .A2(n5392), .A3(n5393), .A4(data[22]), 
        .Y(n2387) );
  AO22X1_HVT U4115 ( .A1(\ram[9][21] ), .A2(n5392), .A3(n5393), .A4(data[21]), 
        .Y(n2386) );
  AO22X1_HVT U4116 ( .A1(\ram[9][20] ), .A2(n5392), .A3(n5393), .A4(data[20]), 
        .Y(n2385) );
  AO22X1_HVT U4117 ( .A1(\ram[9][19] ), .A2(n5392), .A3(n5393), .A4(data[19]), 
        .Y(n2384) );
  AO22X1_HVT U4118 ( .A1(\ram[9][18] ), .A2(n5392), .A3(n5393), .A4(data[18]), 
        .Y(n2383) );
  AO22X1_HVT U4119 ( .A1(\ram[9][17] ), .A2(n5392), .A3(n5393), .A4(data[17]), 
        .Y(n2382) );
  AO22X1_HVT U4120 ( .A1(\ram[9][16] ), .A2(n5392), .A3(n5393), .A4(data[16]), 
        .Y(n2381) );
  AO22X1_HVT U4121 ( .A1(\ram[9][15] ), .A2(n5392), .A3(n5393), .A4(data[15]), 
        .Y(n2380) );
  AO22X1_HVT U4122 ( .A1(\ram[0][177] ), .A2(n5360), .A3(data[177]), .A4(n5361), .Y(n238) );
  AO22X1_HVT U4123 ( .A1(\ram[9][14] ), .A2(n5392), .A3(n5393), .A4(data[14]), 
        .Y(n2379) );
  AO22X1_HVT U4124 ( .A1(\ram[9][13] ), .A2(n5392), .A3(n5393), .A4(data[13]), 
        .Y(n2378) );
  AO22X1_HVT U4125 ( .A1(\ram[9][12] ), .A2(n5392), .A3(n5393), .A4(data[12]), 
        .Y(n2377) );
  AO22X1_HVT U4126 ( .A1(\ram[9][11] ), .A2(n5392), .A3(n5393), .A4(data[11]), 
        .Y(n2376) );
  AO22X1_HVT U4127 ( .A1(\ram[9][10] ), .A2(n5392), .A3(n5393), .A4(data[10]), 
        .Y(n2375) );
  AO22X1_HVT U4128 ( .A1(\ram[9][9] ), .A2(n5392), .A3(n5393), .A4(data[9]), 
        .Y(n2374) );
  AO22X1_HVT U4129 ( .A1(\ram[9][8] ), .A2(n5392), .A3(n5393), .A4(data[8]), 
        .Y(n2373) );
  AO22X1_HVT U4130 ( .A1(\ram[9][7] ), .A2(n5392), .A3(n5393), .A4(data[7]), 
        .Y(n2372) );
  AO22X1_HVT U4131 ( .A1(\ram[9][6] ), .A2(n5392), .A3(n5393), .A4(data[6]), 
        .Y(n2371) );
  AO22X1_HVT U4132 ( .A1(\ram[9][5] ), .A2(n5392), .A3(n5393), .A4(data[5]), 
        .Y(n2370) );
  AO22X1_HVT U4133 ( .A1(\ram[0][176] ), .A2(n5360), .A3(data[176]), .A4(n5361), .Y(n237) );
  AO22X1_HVT U4134 ( .A1(\ram[9][4] ), .A2(n5392), .A3(n5393), .A4(data[4]), 
        .Y(n2369) );
  AO22X1_HVT U4135 ( .A1(\ram[9][3] ), .A2(n5392), .A3(n5393), .A4(data[3]), 
        .Y(n2368) );
  AO22X1_HVT U4136 ( .A1(\ram[9][2] ), .A2(n5392), .A3(n5393), .A4(data[2]), 
        .Y(n2367) );
  AO22X1_HVT U4137 ( .A1(\ram[9][1] ), .A2(n5392), .A3(n5393), .A4(data[1]), 
        .Y(n2366) );
  AO22X1_HVT U4138 ( .A1(\ram[9][0] ), .A2(n5392), .A3(n5393), .A4(data[0]), 
        .Y(n2365) );
  INVX0_HVT U4139 ( .A(n5394), .Y(n5393) );
  AND2X1_HVT U4140 ( .A1(n5394), .A2(n5365), .Y(n5392) );
  NAND3X0_HVT U4141 ( .A1(n5383), .A2(n4182), .A3(n5385), .Y(n5394) );
  AO22X1_HVT U4142 ( .A1(\ram[8][255] ), .A2(n5395), .A3(n5396), .A4(data[255]), .Y(n2364) );
  AO22X1_HVT U4143 ( .A1(\ram[8][254] ), .A2(n5395), .A3(n5396), .A4(data[254]), .Y(n2363) );
  AO22X1_HVT U4144 ( .A1(\ram[8][253] ), .A2(n5395), .A3(n5396), .A4(data[253]), .Y(n2362) );
  AO22X1_HVT U4145 ( .A1(\ram[8][252] ), .A2(n5395), .A3(n5396), .A4(data[252]), .Y(n2361) );
  AO22X1_HVT U4146 ( .A1(\ram[8][251] ), .A2(n5395), .A3(n5396), .A4(data[251]), .Y(n2360) );
  AO22X1_HVT U4147 ( .A1(\ram[0][175] ), .A2(n5360), .A3(data[175]), .A4(n5361), .Y(n236) );
  AO22X1_HVT U4148 ( .A1(\ram[8][250] ), .A2(n5395), .A3(n5396), .A4(data[250]), .Y(n2359) );
  AO22X1_HVT U4149 ( .A1(\ram[8][249] ), .A2(n5395), .A3(n5396), .A4(data[249]), .Y(n2358) );
  AO22X1_HVT U4150 ( .A1(\ram[8][248] ), .A2(n5395), .A3(n5396), .A4(data[248]), .Y(n2357) );
  AO22X1_HVT U4151 ( .A1(\ram[8][247] ), .A2(n5395), .A3(n5396), .A4(data[247]), .Y(n2356) );
  AO22X1_HVT U4152 ( .A1(\ram[8][246] ), .A2(n5395), .A3(n5396), .A4(data[246]), .Y(n2355) );
  AO22X1_HVT U4153 ( .A1(\ram[8][245] ), .A2(n5395), .A3(n5396), .A4(data[245]), .Y(n2354) );
  AO22X1_HVT U4154 ( .A1(\ram[8][244] ), .A2(n5395), .A3(n5396), .A4(data[244]), .Y(n2353) );
  AO22X1_HVT U4155 ( .A1(\ram[8][243] ), .A2(n5395), .A3(n5396), .A4(data[243]), .Y(n2352) );
  AO22X1_HVT U4156 ( .A1(\ram[8][242] ), .A2(n5395), .A3(n5396), .A4(data[242]), .Y(n2351) );
  AO22X1_HVT U4157 ( .A1(\ram[8][241] ), .A2(n5395), .A3(n5396), .A4(data[241]), .Y(n2350) );
  AO22X1_HVT U4158 ( .A1(\ram[0][174] ), .A2(n5360), .A3(data[174]), .A4(n5361), .Y(n235) );
  AO22X1_HVT U4159 ( .A1(\ram[8][240] ), .A2(n5395), .A3(n5396), .A4(data[240]), .Y(n2349) );
  AO22X1_HVT U4160 ( .A1(\ram[8][239] ), .A2(n5395), .A3(n5396), .A4(data[239]), .Y(n2348) );
  AO22X1_HVT U4161 ( .A1(\ram[8][238] ), .A2(n5395), .A3(n5396), .A4(data[238]), .Y(n2347) );
  AO22X1_HVT U4162 ( .A1(\ram[8][237] ), .A2(n5395), .A3(n5396), .A4(data[237]), .Y(n2346) );
  AO22X1_HVT U4163 ( .A1(\ram[8][236] ), .A2(n5395), .A3(n5396), .A4(data[236]), .Y(n2345) );
  AO22X1_HVT U4164 ( .A1(\ram[8][235] ), .A2(n5395), .A3(n5396), .A4(data[235]), .Y(n2344) );
  AO22X1_HVT U4165 ( .A1(\ram[8][234] ), .A2(n5395), .A3(n5396), .A4(data[234]), .Y(n2343) );
  AO22X1_HVT U4166 ( .A1(\ram[8][233] ), .A2(n5395), .A3(n5396), .A4(data[233]), .Y(n2342) );
  AO22X1_HVT U4167 ( .A1(\ram[8][232] ), .A2(n5395), .A3(n5396), .A4(data[232]), .Y(n2341) );
  AO22X1_HVT U4168 ( .A1(\ram[8][231] ), .A2(n5395), .A3(n5396), .A4(data[231]), .Y(n2340) );
  AO22X1_HVT U4169 ( .A1(\ram[0][173] ), .A2(n5360), .A3(data[173]), .A4(n5361), .Y(n234) );
  AO22X1_HVT U4170 ( .A1(\ram[8][230] ), .A2(n5395), .A3(n5396), .A4(data[230]), .Y(n2339) );
  AO22X1_HVT U4171 ( .A1(\ram[8][229] ), .A2(n5395), .A3(n5396), .A4(data[229]), .Y(n2338) );
  AO22X1_HVT U4172 ( .A1(\ram[8][228] ), .A2(n5395), .A3(n5396), .A4(data[228]), .Y(n2337) );
  AO22X1_HVT U4173 ( .A1(\ram[8][227] ), .A2(n5395), .A3(n5396), .A4(data[227]), .Y(n2336) );
  AO22X1_HVT U4174 ( .A1(\ram[8][226] ), .A2(n5395), .A3(n5396), .A4(data[226]), .Y(n2335) );
  AO22X1_HVT U4175 ( .A1(\ram[8][225] ), .A2(n5395), .A3(n5396), .A4(data[225]), .Y(n2334) );
  AO22X1_HVT U4176 ( .A1(\ram[8][224] ), .A2(n5395), .A3(n5396), .A4(data[224]), .Y(n2333) );
  AO22X1_HVT U4177 ( .A1(\ram[8][223] ), .A2(n5395), .A3(n5396), .A4(data[223]), .Y(n2332) );
  AO22X1_HVT U4178 ( .A1(\ram[8][222] ), .A2(n5395), .A3(n5396), .A4(data[222]), .Y(n2331) );
  AO22X1_HVT U4179 ( .A1(\ram[8][221] ), .A2(n5395), .A3(n5396), .A4(data[221]), .Y(n2330) );
  AO22X1_HVT U4180 ( .A1(\ram[0][172] ), .A2(n5360), .A3(data[172]), .A4(n5361), .Y(n233) );
  AO22X1_HVT U4181 ( .A1(\ram[8][220] ), .A2(n5395), .A3(n5396), .A4(data[220]), .Y(n2329) );
  AO22X1_HVT U4182 ( .A1(\ram[8][219] ), .A2(n5395), .A3(n5396), .A4(data[219]), .Y(n2328) );
  AO22X1_HVT U4183 ( .A1(\ram[8][218] ), .A2(n5395), .A3(n5396), .A4(data[218]), .Y(n2327) );
  AO22X1_HVT U4184 ( .A1(\ram[8][217] ), .A2(n5395), .A3(n5396), .A4(data[217]), .Y(n2326) );
  AO22X1_HVT U4185 ( .A1(\ram[8][216] ), .A2(n5395), .A3(n5396), .A4(data[216]), .Y(n2325) );
  AO22X1_HVT U4186 ( .A1(\ram[8][215] ), .A2(n5395), .A3(n5396), .A4(data[215]), .Y(n2324) );
  AO22X1_HVT U4187 ( .A1(\ram[8][214] ), .A2(n5395), .A3(n5396), .A4(data[214]), .Y(n2323) );
  AO22X1_HVT U4188 ( .A1(\ram[8][213] ), .A2(n5395), .A3(n5396), .A4(data[213]), .Y(n2322) );
  AO22X1_HVT U4189 ( .A1(\ram[8][212] ), .A2(n5395), .A3(n5396), .A4(data[212]), .Y(n2321) );
  AO22X1_HVT U4190 ( .A1(\ram[8][211] ), .A2(n5395), .A3(n5396), .A4(data[211]), .Y(n2320) );
  AO22X1_HVT U4191 ( .A1(\ram[0][171] ), .A2(n5360), .A3(data[171]), .A4(n5361), .Y(n232) );
  AO22X1_HVT U4192 ( .A1(\ram[8][210] ), .A2(n5395), .A3(n5396), .A4(data[210]), .Y(n2319) );
  AO22X1_HVT U4193 ( .A1(\ram[8][209] ), .A2(n5395), .A3(n5396), .A4(data[209]), .Y(n2318) );
  AO22X1_HVT U4194 ( .A1(\ram[8][208] ), .A2(n5395), .A3(n5396), .A4(data[208]), .Y(n2317) );
  AO22X1_HVT U4195 ( .A1(\ram[8][207] ), .A2(n5395), .A3(n5396), .A4(data[207]), .Y(n2316) );
  AO22X1_HVT U4196 ( .A1(\ram[8][206] ), .A2(n5395), .A3(n5396), .A4(data[206]), .Y(n2315) );
  AO22X1_HVT U4197 ( .A1(\ram[8][205] ), .A2(n5395), .A3(n5396), .A4(data[205]), .Y(n2314) );
  AO22X1_HVT U4198 ( .A1(\ram[8][204] ), .A2(n5395), .A3(n5396), .A4(data[204]), .Y(n2313) );
  AO22X1_HVT U4199 ( .A1(\ram[8][203] ), .A2(n5395), .A3(n5396), .A4(data[203]), .Y(n2312) );
  AO22X1_HVT U4200 ( .A1(\ram[8][202] ), .A2(n5395), .A3(n5396), .A4(data[202]), .Y(n2311) );
  AO22X1_HVT U4201 ( .A1(\ram[8][201] ), .A2(n5395), .A3(n5396), .A4(data[201]), .Y(n2310) );
  AO22X1_HVT U4202 ( .A1(\ram[0][170] ), .A2(n5360), .A3(n5361), .A4(data[170]), .Y(n231) );
  AO22X1_HVT U4203 ( .A1(\ram[8][200] ), .A2(n5395), .A3(n5396), .A4(data[200]), .Y(n2309) );
  AO22X1_HVT U4204 ( .A1(\ram[8][199] ), .A2(n5395), .A3(n5396), .A4(data[199]), .Y(n2308) );
  AO22X1_HVT U4205 ( .A1(\ram[8][198] ), .A2(n5395), .A3(n5396), .A4(data[198]), .Y(n2307) );
  AO22X1_HVT U4206 ( .A1(\ram[8][197] ), .A2(n5395), .A3(n5396), .A4(data[197]), .Y(n2306) );
  AO22X1_HVT U4207 ( .A1(\ram[8][196] ), .A2(n5395), .A3(n5396), .A4(data[196]), .Y(n2305) );
  AO22X1_HVT U4208 ( .A1(\ram[8][195] ), .A2(n5395), .A3(n5396), .A4(data[195]), .Y(n2304) );
  AO22X1_HVT U4209 ( .A1(\ram[8][194] ), .A2(n5395), .A3(n5396), .A4(data[194]), .Y(n2303) );
  AO22X1_HVT U4210 ( .A1(\ram[8][193] ), .A2(n5395), .A3(n5396), .A4(data[193]), .Y(n2302) );
  AO22X1_HVT U4211 ( .A1(\ram[8][192] ), .A2(n5395), .A3(n5396), .A4(data[192]), .Y(n2301) );
  AO22X1_HVT U4212 ( .A1(\ram[8][191] ), .A2(n5395), .A3(n5396), .A4(data[191]), .Y(n2300) );
  AO22X1_HVT U4213 ( .A1(\ram[0][169] ), .A2(n5360), .A3(n5361), .A4(data[169]), .Y(n230) );
  AO22X1_HVT U4214 ( .A1(\ram[8][190] ), .A2(n5395), .A3(n5396), .A4(data[190]), .Y(n2299) );
  AO22X1_HVT U4215 ( .A1(\ram[8][189] ), .A2(n5395), .A3(n5396), .A4(data[189]), .Y(n2298) );
  AO22X1_HVT U4216 ( .A1(\ram[8][188] ), .A2(n5395), .A3(n5396), .A4(data[188]), .Y(n2297) );
  AO22X1_HVT U4217 ( .A1(\ram[8][187] ), .A2(n5395), .A3(n5396), .A4(data[187]), .Y(n2296) );
  AO22X1_HVT U4218 ( .A1(\ram[8][186] ), .A2(n5395), .A3(n5396), .A4(data[186]), .Y(n2295) );
  AO22X1_HVT U4219 ( .A1(\ram[8][185] ), .A2(n5395), .A3(n5396), .A4(data[185]), .Y(n2294) );
  AO22X1_HVT U4220 ( .A1(\ram[8][184] ), .A2(n5395), .A3(n5396), .A4(data[184]), .Y(n2293) );
  AO22X1_HVT U4221 ( .A1(\ram[8][183] ), .A2(n5395), .A3(n5396), .A4(data[183]), .Y(n2292) );
  AO22X1_HVT U4222 ( .A1(\ram[8][182] ), .A2(n5395), .A3(n5396), .A4(data[182]), .Y(n2291) );
  AO22X1_HVT U4223 ( .A1(\ram[8][181] ), .A2(n5395), .A3(n5396), .A4(data[181]), .Y(n2290) );
  AO22X1_HVT U4224 ( .A1(\ram[0][168] ), .A2(n5360), .A3(n5361), .A4(data[168]), .Y(n229) );
  AO22X1_HVT U4225 ( .A1(\ram[8][180] ), .A2(n5395), .A3(n5396), .A4(data[180]), .Y(n2289) );
  AO22X1_HVT U4226 ( .A1(\ram[8][179] ), .A2(n5395), .A3(n5396), .A4(data[179]), .Y(n2288) );
  AO22X1_HVT U4227 ( .A1(\ram[8][178] ), .A2(n5395), .A3(n5396), .A4(data[178]), .Y(n2287) );
  AO22X1_HVT U4228 ( .A1(\ram[8][177] ), .A2(n5395), .A3(n5396), .A4(data[177]), .Y(n2286) );
  AO22X1_HVT U4229 ( .A1(\ram[8][176] ), .A2(n5395), .A3(n5396), .A4(data[176]), .Y(n2285) );
  AO22X1_HVT U4230 ( .A1(\ram[8][175] ), .A2(n5395), .A3(n5396), .A4(data[175]), .Y(n2284) );
  AO22X1_HVT U4231 ( .A1(\ram[8][174] ), .A2(n5395), .A3(n5396), .A4(data[174]), .Y(n2283) );
  AO22X1_HVT U4232 ( .A1(\ram[8][173] ), .A2(n5395), .A3(n5396), .A4(data[173]), .Y(n2282) );
  AO22X1_HVT U4233 ( .A1(\ram[8][172] ), .A2(n5395), .A3(n5396), .A4(data[172]), .Y(n2281) );
  AO22X1_HVT U4234 ( .A1(\ram[8][171] ), .A2(n5395), .A3(n5396), .A4(data[171]), .Y(n2280) );
  AO22X1_HVT U4235 ( .A1(\ram[0][167] ), .A2(n5360), .A3(n5361), .A4(data[167]), .Y(n228) );
  AO22X1_HVT U4236 ( .A1(\ram[8][170] ), .A2(n5395), .A3(n5396), .A4(data[170]), .Y(n2279) );
  AO22X1_HVT U4237 ( .A1(\ram[8][169] ), .A2(n5395), .A3(n5396), .A4(data[169]), .Y(n2278) );
  AO22X1_HVT U4238 ( .A1(\ram[8][168] ), .A2(n5395), .A3(n5396), .A4(data[168]), .Y(n2277) );
  AO22X1_HVT U4239 ( .A1(\ram[8][167] ), .A2(n5395), .A3(n5396), .A4(data[167]), .Y(n2276) );
  AO22X1_HVT U4240 ( .A1(\ram[8][166] ), .A2(n5395), .A3(n5396), .A4(data[166]), .Y(n2275) );
  AO22X1_HVT U4241 ( .A1(\ram[8][165] ), .A2(n5395), .A3(n5396), .A4(data[165]), .Y(n2274) );
  AO22X1_HVT U4242 ( .A1(\ram[8][164] ), .A2(n5395), .A3(n5396), .A4(data[164]), .Y(n2273) );
  AO22X1_HVT U4243 ( .A1(\ram[8][163] ), .A2(n5395), .A3(n5396), .A4(data[163]), .Y(n2272) );
  AO22X1_HVT U4244 ( .A1(\ram[8][162] ), .A2(n5395), .A3(n5396), .A4(data[162]), .Y(n2271) );
  AO22X1_HVT U4245 ( .A1(\ram[8][161] ), .A2(n5395), .A3(n5396), .A4(data[161]), .Y(n2270) );
  AO22X1_HVT U4246 ( .A1(\ram[0][166] ), .A2(n5360), .A3(n5361), .A4(data[166]), .Y(n227) );
  AO22X1_HVT U4247 ( .A1(\ram[8][160] ), .A2(n5395), .A3(n5396), .A4(data[160]), .Y(n2269) );
  AO22X1_HVT U4248 ( .A1(\ram[8][159] ), .A2(n5395), .A3(n5396), .A4(data[159]), .Y(n2268) );
  AO22X1_HVT U4249 ( .A1(\ram[8][158] ), .A2(n5395), .A3(n5396), .A4(data[158]), .Y(n2267) );
  AO22X1_HVT U4250 ( .A1(\ram[8][157] ), .A2(n5395), .A3(n5396), .A4(data[157]), .Y(n2266) );
  AO22X1_HVT U4251 ( .A1(\ram[8][156] ), .A2(n5395), .A3(n5396), .A4(data[156]), .Y(n2265) );
  AO22X1_HVT U4252 ( .A1(\ram[8][155] ), .A2(n5395), .A3(n5396), .A4(data[155]), .Y(n2264) );
  AO22X1_HVT U4253 ( .A1(\ram[8][154] ), .A2(n5395), .A3(n5396), .A4(data[154]), .Y(n2263) );
  AO22X1_HVT U4254 ( .A1(\ram[8][153] ), .A2(n5395), .A3(n5396), .A4(data[153]), .Y(n2262) );
  AO22X1_HVT U4255 ( .A1(\ram[8][152] ), .A2(n5395), .A3(n5396), .A4(data[152]), .Y(n2261) );
  AO22X1_HVT U4256 ( .A1(\ram[8][151] ), .A2(n5395), .A3(n5396), .A4(data[151]), .Y(n2260) );
  AO22X1_HVT U4257 ( .A1(\ram[0][165] ), .A2(n5360), .A3(n5361), .A4(data[165]), .Y(n226) );
  AO22X1_HVT U4258 ( .A1(\ram[8][150] ), .A2(n5395), .A3(n5396), .A4(data[150]), .Y(n2259) );
  AO22X1_HVT U4259 ( .A1(\ram[8][149] ), .A2(n5395), .A3(n5396), .A4(data[149]), .Y(n2258) );
  AO22X1_HVT U4260 ( .A1(\ram[8][148] ), .A2(n5395), .A3(n5396), .A4(data[148]), .Y(n2257) );
  AO22X1_HVT U4261 ( .A1(\ram[8][147] ), .A2(n5395), .A3(n5396), .A4(data[147]), .Y(n2256) );
  AO22X1_HVT U4262 ( .A1(\ram[8][146] ), .A2(n5395), .A3(n5396), .A4(data[146]), .Y(n2255) );
  AO22X1_HVT U4263 ( .A1(\ram[8][145] ), .A2(n5395), .A3(n5396), .A4(data[145]), .Y(n2254) );
  AO22X1_HVT U4264 ( .A1(\ram[8][144] ), .A2(n5395), .A3(n5396), .A4(data[144]), .Y(n2253) );
  AO22X1_HVT U4265 ( .A1(\ram[8][143] ), .A2(n5395), .A3(n5396), .A4(data[143]), .Y(n2252) );
  AO22X1_HVT U4266 ( .A1(\ram[8][142] ), .A2(n5395), .A3(n5396), .A4(data[142]), .Y(n2251) );
  AO22X1_HVT U4267 ( .A1(\ram[8][141] ), .A2(n5395), .A3(n5396), .A4(data[141]), .Y(n2250) );
  AO22X1_HVT U4268 ( .A1(\ram[0][164] ), .A2(n5360), .A3(n5361), .A4(data[164]), .Y(n225) );
  AO22X1_HVT U4269 ( .A1(\ram[8][140] ), .A2(n5395), .A3(n5396), .A4(data[140]), .Y(n2249) );
  AO22X1_HVT U4270 ( .A1(\ram[8][139] ), .A2(n5395), .A3(n5396), .A4(data[139]), .Y(n2248) );
  AO22X1_HVT U4271 ( .A1(\ram[8][138] ), .A2(n5395), .A3(n5396), .A4(data[138]), .Y(n2247) );
  AO22X1_HVT U4272 ( .A1(\ram[8][137] ), .A2(n5395), .A3(n5396), .A4(data[137]), .Y(n2246) );
  AO22X1_HVT U4273 ( .A1(\ram[8][136] ), .A2(n5395), .A3(n5396), .A4(data[136]), .Y(n2245) );
  AO22X1_HVT U4274 ( .A1(\ram[8][135] ), .A2(n5395), .A3(n5396), .A4(data[135]), .Y(n2244) );
  AO22X1_HVT U4275 ( .A1(\ram[8][134] ), .A2(n5395), .A3(n5396), .A4(data[134]), .Y(n2243) );
  AO22X1_HVT U4276 ( .A1(\ram[8][133] ), .A2(n5395), .A3(n5396), .A4(data[133]), .Y(n2242) );
  AO22X1_HVT U4277 ( .A1(\ram[8][132] ), .A2(n5395), .A3(n5396), .A4(data[132]), .Y(n2241) );
  AO22X1_HVT U4278 ( .A1(\ram[8][131] ), .A2(n5395), .A3(n5396), .A4(data[131]), .Y(n2240) );
  AO22X1_HVT U4279 ( .A1(\ram[0][163] ), .A2(n5360), .A3(n5361), .A4(data[163]), .Y(n224) );
  AO22X1_HVT U4280 ( .A1(\ram[8][130] ), .A2(n5395), .A3(n5396), .A4(data[130]), .Y(n2239) );
  AO22X1_HVT U4281 ( .A1(\ram[8][129] ), .A2(n5395), .A3(n5396), .A4(data[129]), .Y(n2238) );
  AO22X1_HVT U4282 ( .A1(\ram[8][128] ), .A2(n5395), .A3(n5396), .A4(data[128]), .Y(n2237) );
  AO22X1_HVT U4283 ( .A1(\ram[8][127] ), .A2(n5395), .A3(n5396), .A4(data[127]), .Y(n2236) );
  AO22X1_HVT U4284 ( .A1(\ram[8][126] ), .A2(n5395), .A3(n5396), .A4(data[126]), .Y(n2235) );
  AO22X1_HVT U4285 ( .A1(\ram[8][125] ), .A2(n5395), .A3(n5396), .A4(data[125]), .Y(n2234) );
  AO22X1_HVT U4286 ( .A1(\ram[8][124] ), .A2(n5395), .A3(n5396), .A4(data[124]), .Y(n2233) );
  AO22X1_HVT U4287 ( .A1(\ram[8][123] ), .A2(n5395), .A3(n5396), .A4(data[123]), .Y(n2232) );
  AO22X1_HVT U4288 ( .A1(\ram[8][122] ), .A2(n5395), .A3(n5396), .A4(data[122]), .Y(n2231) );
  AO22X1_HVT U4289 ( .A1(\ram[8][121] ), .A2(n5395), .A3(n5396), .A4(data[121]), .Y(n2230) );
  AO22X1_HVT U4290 ( .A1(\ram[0][162] ), .A2(n5360), .A3(n5361), .A4(data[162]), .Y(n223) );
  AO22X1_HVT U4291 ( .A1(\ram[8][120] ), .A2(n5395), .A3(n5396), .A4(data[120]), .Y(n2229) );
  AO22X1_HVT U4292 ( .A1(\ram[8][119] ), .A2(n5395), .A3(n5396), .A4(data[119]), .Y(n2228) );
  AO22X1_HVT U4293 ( .A1(\ram[8][118] ), .A2(n5395), .A3(n5396), .A4(data[118]), .Y(n2227) );
  AO22X1_HVT U4294 ( .A1(\ram[8][117] ), .A2(n5395), .A3(n5396), .A4(data[117]), .Y(n2226) );
  AO22X1_HVT U4295 ( .A1(\ram[8][116] ), .A2(n5395), .A3(n5396), .A4(data[116]), .Y(n2225) );
  AO22X1_HVT U4296 ( .A1(\ram[8][115] ), .A2(n5395), .A3(n5396), .A4(data[115]), .Y(n2224) );
  AO22X1_HVT U4297 ( .A1(\ram[8][114] ), .A2(n5395), .A3(n5396), .A4(data[114]), .Y(n2223) );
  AO22X1_HVT U4298 ( .A1(\ram[8][113] ), .A2(n5395), .A3(n5396), .A4(data[113]), .Y(n2222) );
  AO22X1_HVT U4299 ( .A1(\ram[8][112] ), .A2(n5395), .A3(n5396), .A4(data[112]), .Y(n2221) );
  AO22X1_HVT U4300 ( .A1(\ram[8][111] ), .A2(n5395), .A3(n5396), .A4(data[111]), .Y(n2220) );
  AO22X1_HVT U4301 ( .A1(\ram[0][161] ), .A2(n5360), .A3(n5361), .A4(data[161]), .Y(n222) );
  AO22X1_HVT U4302 ( .A1(\ram[8][110] ), .A2(n5395), .A3(n5396), .A4(data[110]), .Y(n2219) );
  AO22X1_HVT U4303 ( .A1(\ram[8][109] ), .A2(n5395), .A3(n5396), .A4(data[109]), .Y(n2218) );
  AO22X1_HVT U4304 ( .A1(\ram[8][108] ), .A2(n5395), .A3(n5396), .A4(data[108]), .Y(n2217) );
  AO22X1_HVT U4305 ( .A1(\ram[8][107] ), .A2(n5395), .A3(n5396), .A4(data[107]), .Y(n2216) );
  AO22X1_HVT U4306 ( .A1(\ram[8][106] ), .A2(n5395), .A3(n5396), .A4(data[106]), .Y(n2215) );
  AO22X1_HVT U4307 ( .A1(\ram[8][105] ), .A2(n5395), .A3(n5396), .A4(data[105]), .Y(n2214) );
  AO22X1_HVT U4308 ( .A1(\ram[8][104] ), .A2(n5395), .A3(n5396), .A4(data[104]), .Y(n2213) );
  AO22X1_HVT U4309 ( .A1(\ram[8][103] ), .A2(n5395), .A3(n5396), .A4(data[103]), .Y(n2212) );
  AO22X1_HVT U4310 ( .A1(\ram[8][102] ), .A2(n5395), .A3(n5396), .A4(data[102]), .Y(n2211) );
  AO22X1_HVT U4311 ( .A1(\ram[8][101] ), .A2(n5395), .A3(n5396), .A4(data[101]), .Y(n2210) );
  AO22X1_HVT U4312 ( .A1(\ram[0][160] ), .A2(n5360), .A3(data[160]), .A4(n5361), .Y(n221) );
  AO22X1_HVT U4313 ( .A1(\ram[8][100] ), .A2(n5395), .A3(n5396), .A4(data[100]), .Y(n2209) );
  AO22X1_HVT U4314 ( .A1(\ram[8][99] ), .A2(n5395), .A3(n5396), .A4(data[99]), 
        .Y(n2208) );
  AO22X1_HVT U4315 ( .A1(\ram[8][98] ), .A2(n5395), .A3(n5396), .A4(data[98]), 
        .Y(n2207) );
  AO22X1_HVT U4316 ( .A1(\ram[8][97] ), .A2(n5395), .A3(n5396), .A4(data[97]), 
        .Y(n2206) );
  AO22X1_HVT U4317 ( .A1(\ram[8][96] ), .A2(n5395), .A3(n5396), .A4(data[96]), 
        .Y(n2205) );
  AO22X1_HVT U4318 ( .A1(\ram[8][95] ), .A2(n5395), .A3(n5396), .A4(data[95]), 
        .Y(n2204) );
  AO22X1_HVT U4319 ( .A1(\ram[8][94] ), .A2(n5395), .A3(n5396), .A4(data[94]), 
        .Y(n2203) );
  AO22X1_HVT U4320 ( .A1(\ram[8][93] ), .A2(n5395), .A3(n5396), .A4(data[93]), 
        .Y(n2202) );
  AO22X1_HVT U4321 ( .A1(\ram[8][92] ), .A2(n5395), .A3(n5396), .A4(data[92]), 
        .Y(n2201) );
  AO22X1_HVT U4322 ( .A1(\ram[8][91] ), .A2(n5395), .A3(n5396), .A4(data[91]), 
        .Y(n2200) );
  AO22X1_HVT U4323 ( .A1(\ram[0][159] ), .A2(n5360), .A3(data[159]), .A4(n5361), .Y(n220) );
  AO22X1_HVT U4324 ( .A1(\ram[8][90] ), .A2(n5395), .A3(n5396), .A4(data[90]), 
        .Y(n2199) );
  AO22X1_HVT U4325 ( .A1(\ram[8][89] ), .A2(n5395), .A3(n5396), .A4(data[89]), 
        .Y(n2198) );
  AO22X1_HVT U4326 ( .A1(\ram[8][88] ), .A2(n5395), .A3(n5396), .A4(data[88]), 
        .Y(n2197) );
  AO22X1_HVT U4327 ( .A1(\ram[8][87] ), .A2(n5395), .A3(n5396), .A4(data[87]), 
        .Y(n2196) );
  AO22X1_HVT U4328 ( .A1(\ram[8][86] ), .A2(n5395), .A3(n5396), .A4(data[86]), 
        .Y(n2195) );
  AO22X1_HVT U4329 ( .A1(\ram[8][85] ), .A2(n5395), .A3(n5396), .A4(data[85]), 
        .Y(n2194) );
  AO22X1_HVT U4330 ( .A1(\ram[8][84] ), .A2(n5395), .A3(n5396), .A4(data[84]), 
        .Y(n2193) );
  AO22X1_HVT U4331 ( .A1(\ram[8][83] ), .A2(n5395), .A3(n5396), .A4(data[83]), 
        .Y(n2192) );
  AO22X1_HVT U4332 ( .A1(\ram[8][82] ), .A2(n5395), .A3(n5396), .A4(data[82]), 
        .Y(n2191) );
  AO22X1_HVT U4333 ( .A1(\ram[8][81] ), .A2(n5395), .A3(n5396), .A4(data[81]), 
        .Y(n2190) );
  AO22X1_HVT U4334 ( .A1(\ram[0][158] ), .A2(n5360), .A3(data[158]), .A4(n5361), .Y(n219) );
  AO22X1_HVT U4335 ( .A1(\ram[8][80] ), .A2(n5395), .A3(n5396), .A4(data[80]), 
        .Y(n2189) );
  AO22X1_HVT U4336 ( .A1(\ram[8][79] ), .A2(n5395), .A3(n5396), .A4(data[79]), 
        .Y(n2188) );
  AO22X1_HVT U4337 ( .A1(\ram[8][78] ), .A2(n5395), .A3(n5396), .A4(data[78]), 
        .Y(n2187) );
  AO22X1_HVT U4338 ( .A1(\ram[8][77] ), .A2(n5395), .A3(n5396), .A4(data[77]), 
        .Y(n2186) );
  AO22X1_HVT U4339 ( .A1(\ram[8][76] ), .A2(n5395), .A3(n5396), .A4(data[76]), 
        .Y(n2185) );
  AO22X1_HVT U4340 ( .A1(\ram[8][75] ), .A2(n5395), .A3(n5396), .A4(data[75]), 
        .Y(n2184) );
  AO22X1_HVT U4341 ( .A1(\ram[8][74] ), .A2(n5395), .A3(n5396), .A4(data[74]), 
        .Y(n2183) );
  AO22X1_HVT U4342 ( .A1(\ram[8][73] ), .A2(n5395), .A3(n5396), .A4(data[73]), 
        .Y(n2182) );
  AO22X1_HVT U4343 ( .A1(\ram[8][72] ), .A2(n5395), .A3(n5396), .A4(data[72]), 
        .Y(n2181) );
  AO22X1_HVT U4344 ( .A1(\ram[8][71] ), .A2(n5395), .A3(n5396), .A4(data[71]), 
        .Y(n2180) );
  AO22X1_HVT U4345 ( .A1(\ram[0][157] ), .A2(n5360), .A3(data[157]), .A4(n5361), .Y(n218) );
  AO22X1_HVT U4346 ( .A1(\ram[8][70] ), .A2(n5395), .A3(n5396), .A4(data[70]), 
        .Y(n2179) );
  AO22X1_HVT U4347 ( .A1(\ram[8][69] ), .A2(n5395), .A3(n5396), .A4(data[69]), 
        .Y(n2178) );
  AO22X1_HVT U4348 ( .A1(\ram[8][68] ), .A2(n5395), .A3(n5396), .A4(data[68]), 
        .Y(n2177) );
  AO22X1_HVT U4349 ( .A1(\ram[8][67] ), .A2(n5395), .A3(n5396), .A4(data[67]), 
        .Y(n2176) );
  AO22X1_HVT U4350 ( .A1(\ram[8][66] ), .A2(n5395), .A3(n5396), .A4(data[66]), 
        .Y(n2175) );
  AO22X1_HVT U4351 ( .A1(\ram[8][65] ), .A2(n5395), .A3(n5396), .A4(data[65]), 
        .Y(n2174) );
  AO22X1_HVT U4352 ( .A1(\ram[8][64] ), .A2(n5395), .A3(n5396), .A4(data[64]), 
        .Y(n2173) );
  AO22X1_HVT U4353 ( .A1(\ram[8][63] ), .A2(n5395), .A3(n5396), .A4(data[63]), 
        .Y(n2172) );
  AO22X1_HVT U4354 ( .A1(\ram[8][62] ), .A2(n5395), .A3(n5396), .A4(data[62]), 
        .Y(n2171) );
  AO22X1_HVT U4355 ( .A1(\ram[8][61] ), .A2(n5395), .A3(n5396), .A4(data[61]), 
        .Y(n2170) );
  AO22X1_HVT U4356 ( .A1(\ram[0][156] ), .A2(n5360), .A3(data[156]), .A4(n5361), .Y(n217) );
  AO22X1_HVT U4357 ( .A1(\ram[8][60] ), .A2(n5395), .A3(n5396), .A4(data[60]), 
        .Y(n2169) );
  AO22X1_HVT U4358 ( .A1(\ram[8][59] ), .A2(n5395), .A3(n5396), .A4(data[59]), 
        .Y(n2168) );
  AO22X1_HVT U4359 ( .A1(\ram[8][58] ), .A2(n5395), .A3(n5396), .A4(data[58]), 
        .Y(n2167) );
  AO22X1_HVT U4360 ( .A1(\ram[8][57] ), .A2(n5395), .A3(n5396), .A4(data[57]), 
        .Y(n2166) );
  AO22X1_HVT U4361 ( .A1(\ram[8][56] ), .A2(n5395), .A3(n5396), .A4(data[56]), 
        .Y(n2165) );
  AO22X1_HVT U4362 ( .A1(\ram[8][55] ), .A2(n5395), .A3(n5396), .A4(data[55]), 
        .Y(n2164) );
  AO22X1_HVT U4363 ( .A1(\ram[8][54] ), .A2(n5395), .A3(n5396), .A4(data[54]), 
        .Y(n2163) );
  AO22X1_HVT U4364 ( .A1(\ram[8][53] ), .A2(n5395), .A3(n5396), .A4(data[53]), 
        .Y(n2162) );
  AO22X1_HVT U4365 ( .A1(\ram[8][52] ), .A2(n5395), .A3(n5396), .A4(data[52]), 
        .Y(n2161) );
  AO22X1_HVT U4366 ( .A1(\ram[8][51] ), .A2(n5395), .A3(n5396), .A4(data[51]), 
        .Y(n2160) );
  AO22X1_HVT U4367 ( .A1(\ram[0][155] ), .A2(n5360), .A3(data[155]), .A4(n5361), .Y(n216) );
  AO22X1_HVT U4368 ( .A1(\ram[8][50] ), .A2(n5395), .A3(n5396), .A4(data[50]), 
        .Y(n2159) );
  AO22X1_HVT U4369 ( .A1(\ram[8][49] ), .A2(n5395), .A3(n5396), .A4(data[49]), 
        .Y(n2158) );
  AO22X1_HVT U4370 ( .A1(\ram[8][48] ), .A2(n5395), .A3(n5396), .A4(data[48]), 
        .Y(n2157) );
  AO22X1_HVT U4371 ( .A1(\ram[8][47] ), .A2(n5395), .A3(n5396), .A4(data[47]), 
        .Y(n2156) );
  AO22X1_HVT U4372 ( .A1(\ram[8][46] ), .A2(n5395), .A3(n5396), .A4(data[46]), 
        .Y(n2155) );
  AO22X1_HVT U4373 ( .A1(\ram[8][45] ), .A2(n5395), .A3(n5396), .A4(data[45]), 
        .Y(n2154) );
  AO22X1_HVT U4374 ( .A1(\ram[8][44] ), .A2(n5395), .A3(n5396), .A4(data[44]), 
        .Y(n2153) );
  AO22X1_HVT U4375 ( .A1(\ram[8][43] ), .A2(n5395), .A3(n5396), .A4(data[43]), 
        .Y(n2152) );
  AO22X1_HVT U4376 ( .A1(\ram[8][42] ), .A2(n5395), .A3(n5396), .A4(data[42]), 
        .Y(n2151) );
  AO22X1_HVT U4377 ( .A1(\ram[8][41] ), .A2(n5395), .A3(n5396), .A4(data[41]), 
        .Y(n2150) );
  AO22X1_HVT U4378 ( .A1(\ram[0][154] ), .A2(n5360), .A3(data[154]), .A4(n5361), .Y(n215) );
  AO22X1_HVT U4379 ( .A1(\ram[8][40] ), .A2(n5395), .A3(n5396), .A4(data[40]), 
        .Y(n2149) );
  AO22X1_HVT U4380 ( .A1(\ram[8][39] ), .A2(n5395), .A3(n5396), .A4(data[39]), 
        .Y(n2148) );
  AO22X1_HVT U4381 ( .A1(\ram[8][38] ), .A2(n5395), .A3(n5396), .A4(data[38]), 
        .Y(n2147) );
  AO22X1_HVT U4382 ( .A1(\ram[8][37] ), .A2(n5395), .A3(n5396), .A4(data[37]), 
        .Y(n2146) );
  AO22X1_HVT U4383 ( .A1(\ram[8][36] ), .A2(n5395), .A3(n5396), .A4(data[36]), 
        .Y(n2145) );
  AO22X1_HVT U4384 ( .A1(\ram[8][35] ), .A2(n5395), .A3(n5396), .A4(data[35]), 
        .Y(n2144) );
  AO22X1_HVT U4385 ( .A1(\ram[8][34] ), .A2(n5395), .A3(n5396), .A4(data[34]), 
        .Y(n2143) );
  AO22X1_HVT U4386 ( .A1(\ram[8][33] ), .A2(n5395), .A3(n5396), .A4(data[33]), 
        .Y(n2142) );
  AO22X1_HVT U4387 ( .A1(\ram[8][32] ), .A2(n5395), .A3(n5396), .A4(data[32]), 
        .Y(n2141) );
  AO22X1_HVT U4388 ( .A1(\ram[8][31] ), .A2(n5395), .A3(n5396), .A4(data[31]), 
        .Y(n2140) );
  AO22X1_HVT U4389 ( .A1(\ram[0][153] ), .A2(n5360), .A3(data[153]), .A4(n5361), .Y(n214) );
  AO22X1_HVT U4390 ( .A1(\ram[8][30] ), .A2(n5395), .A3(n5396), .A4(data[30]), 
        .Y(n2139) );
  AO22X1_HVT U4391 ( .A1(\ram[8][29] ), .A2(n5395), .A3(n5396), .A4(data[29]), 
        .Y(n2138) );
  AO22X1_HVT U4392 ( .A1(\ram[8][28] ), .A2(n5395), .A3(n5396), .A4(data[28]), 
        .Y(n2137) );
  AO22X1_HVT U4393 ( .A1(\ram[8][27] ), .A2(n5395), .A3(n5396), .A4(data[27]), 
        .Y(n2136) );
  AO22X1_HVT U4394 ( .A1(\ram[8][26] ), .A2(n5395), .A3(n5396), .A4(data[26]), 
        .Y(n2135) );
  AO22X1_HVT U4395 ( .A1(\ram[8][25] ), .A2(n5395), .A3(n5396), .A4(data[25]), 
        .Y(n2134) );
  AO22X1_HVT U4396 ( .A1(\ram[8][24] ), .A2(n5395), .A3(n5396), .A4(data[24]), 
        .Y(n2133) );
  AO22X1_HVT U4397 ( .A1(\ram[8][23] ), .A2(n5395), .A3(n5396), .A4(data[23]), 
        .Y(n2132) );
  AO22X1_HVT U4398 ( .A1(\ram[8][22] ), .A2(n5395), .A3(n5396), .A4(data[22]), 
        .Y(n2131) );
  AO22X1_HVT U4399 ( .A1(\ram[8][21] ), .A2(n5395), .A3(n5396), .A4(data[21]), 
        .Y(n2130) );
  AO22X1_HVT U4400 ( .A1(\ram[0][152] ), .A2(n5360), .A3(data[152]), .A4(n5361), .Y(n213) );
  AO22X1_HVT U4401 ( .A1(\ram[8][20] ), .A2(n5395), .A3(n5396), .A4(data[20]), 
        .Y(n2129) );
  AO22X1_HVT U4402 ( .A1(\ram[8][19] ), .A2(n5395), .A3(n5396), .A4(data[19]), 
        .Y(n2128) );
  AO22X1_HVT U4403 ( .A1(\ram[8][18] ), .A2(n5395), .A3(n5396), .A4(data[18]), 
        .Y(n2127) );
  AO22X1_HVT U4404 ( .A1(\ram[8][17] ), .A2(n5395), .A3(n5396), .A4(data[17]), 
        .Y(n2126) );
  AO22X1_HVT U4405 ( .A1(\ram[8][16] ), .A2(n5395), .A3(n5396), .A4(data[16]), 
        .Y(n2125) );
  AO22X1_HVT U4406 ( .A1(\ram[8][15] ), .A2(n5395), .A3(n5396), .A4(data[15]), 
        .Y(n2124) );
  AO22X1_HVT U4407 ( .A1(\ram[8][14] ), .A2(n5395), .A3(n5396), .A4(data[14]), 
        .Y(n2123) );
  AO22X1_HVT U4408 ( .A1(\ram[8][13] ), .A2(n5395), .A3(n5396), .A4(data[13]), 
        .Y(n2122) );
  AO22X1_HVT U4409 ( .A1(\ram[8][12] ), .A2(n5395), .A3(n5396), .A4(data[12]), 
        .Y(n2121) );
  AO22X1_HVT U4410 ( .A1(\ram[8][11] ), .A2(n5395), .A3(n5396), .A4(data[11]), 
        .Y(n2120) );
  AO22X1_HVT U4411 ( .A1(\ram[0][151] ), .A2(n5360), .A3(data[151]), .A4(n5361), .Y(n212) );
  AO22X1_HVT U4412 ( .A1(\ram[8][10] ), .A2(n5395), .A3(n5396), .A4(data[10]), 
        .Y(n2119) );
  AO22X1_HVT U4413 ( .A1(\ram[8][9] ), .A2(n5395), .A3(n5396), .A4(data[9]), 
        .Y(n2118) );
  AO22X1_HVT U4414 ( .A1(\ram[8][8] ), .A2(n5395), .A3(n5396), .A4(data[8]), 
        .Y(n2117) );
  AO22X1_HVT U4415 ( .A1(\ram[8][7] ), .A2(n5395), .A3(n5396), .A4(data[7]), 
        .Y(n2116) );
  AO22X1_HVT U4416 ( .A1(\ram[8][6] ), .A2(n5395), .A3(n5396), .A4(data[6]), 
        .Y(n2115) );
  AO22X1_HVT U4417 ( .A1(\ram[8][5] ), .A2(n5395), .A3(n5396), .A4(data[5]), 
        .Y(n2114) );
  AO22X1_HVT U4418 ( .A1(\ram[8][4] ), .A2(n5395), .A3(n5396), .A4(data[4]), 
        .Y(n2113) );
  AO22X1_HVT U4419 ( .A1(\ram[8][3] ), .A2(n5395), .A3(n5396), .A4(data[3]), 
        .Y(n2112) );
  AO22X1_HVT U4420 ( .A1(\ram[8][2] ), .A2(n5395), .A3(n5396), .A4(data[2]), 
        .Y(n2111) );
  AO22X1_HVT U4421 ( .A1(\ram[8][1] ), .A2(n5395), .A3(n5396), .A4(data[1]), 
        .Y(n2110) );
  AO22X1_HVT U4422 ( .A1(\ram[0][150] ), .A2(n5360), .A3(data[150]), .A4(n5361), .Y(n211) );
  AO22X1_HVT U4423 ( .A1(\ram[8][0] ), .A2(n5395), .A3(n5396), .A4(data[0]), 
        .Y(n2109) );
  INVX0_HVT U4424 ( .A(n5397), .Y(n5396) );
  AND2X1_HVT U4425 ( .A1(n5397), .A2(n5365), .Y(n5395) );
  NAND3X0_HVT U4426 ( .A1(n5383), .A2(n4183), .A3(n5385), .Y(n5397) );
  AND2X1_HVT U4427 ( .A1(N29), .A2(we), .Y(n5385) );
  AO22X1_HVT U4428 ( .A1(\ram[7][255] ), .A2(n5398), .A3(n5399), .A4(data[255]), .Y(n2108) );
  AO22X1_HVT U4429 ( .A1(\ram[7][254] ), .A2(n5398), .A3(n5399), .A4(data[254]), .Y(n2107) );
  AO22X1_HVT U4430 ( .A1(\ram[7][253] ), .A2(n5398), .A3(n5399), .A4(data[253]), .Y(n2106) );
  AO22X1_HVT U4431 ( .A1(\ram[7][252] ), .A2(n5398), .A3(n5399), .A4(data[252]), .Y(n2105) );
  AO22X1_HVT U4432 ( .A1(\ram[7][251] ), .A2(n5398), .A3(n5399), .A4(data[251]), .Y(n2104) );
  AO22X1_HVT U4433 ( .A1(\ram[7][250] ), .A2(n5398), .A3(n5399), .A4(data[250]), .Y(n2103) );
  AO22X1_HVT U4434 ( .A1(\ram[7][249] ), .A2(n5398), .A3(n5399), .A4(data[249]), .Y(n2102) );
  AO22X1_HVT U4435 ( .A1(\ram[7][248] ), .A2(n5398), .A3(n5399), .A4(data[248]), .Y(n2101) );
  AO22X1_HVT U4436 ( .A1(\ram[7][247] ), .A2(n5398), .A3(n5399), .A4(data[247]), .Y(n2100) );
  AO22X1_HVT U4437 ( .A1(\ram[0][149] ), .A2(n5360), .A3(data[149]), .A4(n5361), .Y(n210) );
  AO22X1_HVT U4438 ( .A1(\ram[7][246] ), .A2(n5398), .A3(n5399), .A4(data[246]), .Y(n2099) );
  AO22X1_HVT U4439 ( .A1(\ram[7][245] ), .A2(n5398), .A3(n5399), .A4(data[245]), .Y(n2098) );
  AO22X1_HVT U4440 ( .A1(\ram[7][244] ), .A2(n5398), .A3(n5399), .A4(data[244]), .Y(n2097) );
  AO22X1_HVT U4441 ( .A1(\ram[7][243] ), .A2(n5398), .A3(n5399), .A4(data[243]), .Y(n2096) );
  AO22X1_HVT U4442 ( .A1(\ram[7][242] ), .A2(n5398), .A3(n5399), .A4(data[242]), .Y(n2095) );
  AO22X1_HVT U4443 ( .A1(\ram[7][241] ), .A2(n5398), .A3(n5399), .A4(data[241]), .Y(n2094) );
  AO22X1_HVT U4444 ( .A1(\ram[7][240] ), .A2(n5398), .A3(n5399), .A4(data[240]), .Y(n2093) );
  AO22X1_HVT U4445 ( .A1(\ram[7][239] ), .A2(n5398), .A3(n5399), .A4(data[239]), .Y(n2092) );
  AO22X1_HVT U4446 ( .A1(\ram[7][238] ), .A2(n5398), .A3(n5399), .A4(data[238]), .Y(n2091) );
  AO22X1_HVT U4447 ( .A1(\ram[7][237] ), .A2(n5398), .A3(n5399), .A4(data[237]), .Y(n2090) );
  AO22X1_HVT U4448 ( .A1(\ram[0][148] ), .A2(n5360), .A3(data[148]), .A4(n5361), .Y(n209) );
  AO22X1_HVT U4449 ( .A1(\ram[7][236] ), .A2(n5398), .A3(n5399), .A4(data[236]), .Y(n2089) );
  AO22X1_HVT U4450 ( .A1(\ram[7][235] ), .A2(n5398), .A3(n5399), .A4(data[235]), .Y(n2088) );
  AO22X1_HVT U4451 ( .A1(\ram[7][234] ), .A2(n5398), .A3(n5399), .A4(data[234]), .Y(n2087) );
  AO22X1_HVT U4452 ( .A1(\ram[7][233] ), .A2(n5398), .A3(n5399), .A4(data[233]), .Y(n2086) );
  AO22X1_HVT U4453 ( .A1(\ram[7][232] ), .A2(n5398), .A3(n5399), .A4(data[232]), .Y(n2085) );
  AO22X1_HVT U4454 ( .A1(\ram[7][231] ), .A2(n5398), .A3(n5399), .A4(data[231]), .Y(n2084) );
  AO22X1_HVT U4455 ( .A1(\ram[7][230] ), .A2(n5398), .A3(n5399), .A4(data[230]), .Y(n2083) );
  AO22X1_HVT U4456 ( .A1(\ram[7][229] ), .A2(n5398), .A3(n5399), .A4(data[229]), .Y(n2082) );
  AO22X1_HVT U4457 ( .A1(\ram[7][228] ), .A2(n5398), .A3(n5399), .A4(data[228]), .Y(n2081) );
  AO22X1_HVT U4458 ( .A1(\ram[7][227] ), .A2(n5398), .A3(n5399), .A4(data[227]), .Y(n2080) );
  AO22X1_HVT U4459 ( .A1(\ram[0][147] ), .A2(n5360), .A3(data[147]), .A4(n5361), .Y(n208) );
  AO22X1_HVT U4460 ( .A1(\ram[7][226] ), .A2(n5398), .A3(n5399), .A4(data[226]), .Y(n2079) );
  AO22X1_HVT U4461 ( .A1(\ram[7][225] ), .A2(n5398), .A3(n5399), .A4(data[225]), .Y(n2078) );
  AO22X1_HVT U4462 ( .A1(\ram[7][224] ), .A2(n5398), .A3(n5399), .A4(data[224]), .Y(n2077) );
  AO22X1_HVT U4463 ( .A1(\ram[7][223] ), .A2(n5398), .A3(n5399), .A4(data[223]), .Y(n2076) );
  AO22X1_HVT U4464 ( .A1(\ram[7][222] ), .A2(n5398), .A3(n5399), .A4(data[222]), .Y(n2075) );
  AO22X1_HVT U4465 ( .A1(\ram[7][221] ), .A2(n5398), .A3(n5399), .A4(data[221]), .Y(n2074) );
  AO22X1_HVT U4466 ( .A1(\ram[7][220] ), .A2(n5398), .A3(n5399), .A4(data[220]), .Y(n2073) );
  AO22X1_HVT U4467 ( .A1(\ram[7][219] ), .A2(n5398), .A3(n5399), .A4(data[219]), .Y(n2072) );
  AO22X1_HVT U4468 ( .A1(\ram[7][218] ), .A2(n5398), .A3(n5399), .A4(data[218]), .Y(n2071) );
  AO22X1_HVT U4469 ( .A1(\ram[7][217] ), .A2(n5398), .A3(n5399), .A4(data[217]), .Y(n2070) );
  AO22X1_HVT U4470 ( .A1(\ram[0][146] ), .A2(n5360), .A3(data[146]), .A4(n5361), .Y(n207) );
  AO22X1_HVT U4471 ( .A1(\ram[7][216] ), .A2(n5398), .A3(n5399), .A4(data[216]), .Y(n2069) );
  AO22X1_HVT U4472 ( .A1(\ram[7][215] ), .A2(n5398), .A3(n5399), .A4(data[215]), .Y(n2068) );
  AO22X1_HVT U4473 ( .A1(\ram[7][214] ), .A2(n5398), .A3(n5399), .A4(data[214]), .Y(n2067) );
  AO22X1_HVT U4474 ( .A1(\ram[7][213] ), .A2(n5398), .A3(n5399), .A4(data[213]), .Y(n2066) );
  AO22X1_HVT U4475 ( .A1(\ram[7][212] ), .A2(n5398), .A3(n5399), .A4(data[212]), .Y(n2065) );
  AO22X1_HVT U4476 ( .A1(\ram[7][211] ), .A2(n5398), .A3(n5399), .A4(data[211]), .Y(n2064) );
  AO22X1_HVT U4477 ( .A1(\ram[7][210] ), .A2(n5398), .A3(n5399), .A4(data[210]), .Y(n2063) );
  AO22X1_HVT U4478 ( .A1(\ram[7][209] ), .A2(n5398), .A3(n5399), .A4(data[209]), .Y(n2062) );
  AO22X1_HVT U4479 ( .A1(\ram[7][208] ), .A2(n5398), .A3(n5399), .A4(data[208]), .Y(n2061) );
  AO22X1_HVT U4480 ( .A1(\ram[7][207] ), .A2(n5398), .A3(n5399), .A4(data[207]), .Y(n2060) );
  AO22X1_HVT U4481 ( .A1(\ram[0][145] ), .A2(n5360), .A3(data[145]), .A4(n5361), .Y(n206) );
  AO22X1_HVT U4482 ( .A1(\ram[7][206] ), .A2(n5398), .A3(n5399), .A4(data[206]), .Y(n2059) );
  AO22X1_HVT U4483 ( .A1(\ram[7][205] ), .A2(n5398), .A3(n5399), .A4(data[205]), .Y(n2058) );
  AO22X1_HVT U4484 ( .A1(\ram[7][204] ), .A2(n5398), .A3(n5399), .A4(data[204]), .Y(n2057) );
  AO22X1_HVT U4485 ( .A1(\ram[7][203] ), .A2(n5398), .A3(n5399), .A4(data[203]), .Y(n2056) );
  AO22X1_HVT U4486 ( .A1(\ram[7][202] ), .A2(n5398), .A3(n5399), .A4(data[202]), .Y(n2055) );
  AO22X1_HVT U4487 ( .A1(\ram[7][201] ), .A2(n5398), .A3(n5399), .A4(data[201]), .Y(n2054) );
  AO22X1_HVT U4488 ( .A1(\ram[7][200] ), .A2(n5398), .A3(n5399), .A4(data[200]), .Y(n2053) );
  AO22X1_HVT U4489 ( .A1(\ram[7][199] ), .A2(n5398), .A3(n5399), .A4(data[199]), .Y(n2052) );
  AO22X1_HVT U4490 ( .A1(\ram[7][198] ), .A2(n5398), .A3(n5399), .A4(data[198]), .Y(n2051) );
  AO22X1_HVT U4491 ( .A1(\ram[7][197] ), .A2(n5398), .A3(n5399), .A4(data[197]), .Y(n2050) );
  AO22X1_HVT U4492 ( .A1(\ram[0][144] ), .A2(n5360), .A3(data[144]), .A4(n5361), .Y(n205) );
  AO22X1_HVT U4493 ( .A1(\ram[7][196] ), .A2(n5398), .A3(n5399), .A4(data[196]), .Y(n2049) );
  AO22X1_HVT U4494 ( .A1(\ram[7][195] ), .A2(n5398), .A3(n5399), .A4(data[195]), .Y(n2048) );
  AO22X1_HVT U4495 ( .A1(\ram[7][194] ), .A2(n5398), .A3(n5399), .A4(data[194]), .Y(n2047) );
  AO22X1_HVT U4496 ( .A1(\ram[7][193] ), .A2(n5398), .A3(n5399), .A4(data[193]), .Y(n2046) );
  AO22X1_HVT U4497 ( .A1(\ram[7][192] ), .A2(n5398), .A3(n5399), .A4(data[192]), .Y(n2045) );
  AO22X1_HVT U4498 ( .A1(\ram[7][191] ), .A2(n5398), .A3(n5399), .A4(data[191]), .Y(n2044) );
  AO22X1_HVT U4499 ( .A1(\ram[7][190] ), .A2(n5398), .A3(n5399), .A4(data[190]), .Y(n2043) );
  AO22X1_HVT U4500 ( .A1(\ram[7][189] ), .A2(n5398), .A3(n5399), .A4(data[189]), .Y(n2042) );
  AO22X1_HVT U4501 ( .A1(\ram[7][188] ), .A2(n5398), .A3(n5399), .A4(data[188]), .Y(n2041) );
  AO22X1_HVT U4502 ( .A1(\ram[7][187] ), .A2(n5398), .A3(n5399), .A4(data[187]), .Y(n2040) );
  AO22X1_HVT U4503 ( .A1(\ram[0][143] ), .A2(n5360), .A3(data[143]), .A4(n5361), .Y(n204) );
  AO22X1_HVT U4504 ( .A1(\ram[7][186] ), .A2(n5398), .A3(n5399), .A4(data[186]), .Y(n2039) );
  AO22X1_HVT U4505 ( .A1(\ram[7][185] ), .A2(n5398), .A3(n5399), .A4(data[185]), .Y(n2038) );
  AO22X1_HVT U4506 ( .A1(\ram[7][184] ), .A2(n5398), .A3(n5399), .A4(data[184]), .Y(n2037) );
  AO22X1_HVT U4507 ( .A1(\ram[7][183] ), .A2(n5398), .A3(n5399), .A4(data[183]), .Y(n2036) );
  AO22X1_HVT U4508 ( .A1(\ram[7][182] ), .A2(n5398), .A3(n5399), .A4(data[182]), .Y(n2035) );
  AO22X1_HVT U4509 ( .A1(\ram[7][181] ), .A2(n5398), .A3(n5399), .A4(data[181]), .Y(n2034) );
  AO22X1_HVT U4510 ( .A1(\ram[7][180] ), .A2(n5398), .A3(n5399), .A4(data[180]), .Y(n2033) );
  AO22X1_HVT U4511 ( .A1(\ram[7][179] ), .A2(n5398), .A3(n5399), .A4(data[179]), .Y(n2032) );
  AO22X1_HVT U4512 ( .A1(\ram[7][178] ), .A2(n5398), .A3(n5399), .A4(data[178]), .Y(n2031) );
  AO22X1_HVT U4513 ( .A1(\ram[7][177] ), .A2(n5398), .A3(n5399), .A4(data[177]), .Y(n2030) );
  AO22X1_HVT U4514 ( .A1(\ram[0][142] ), .A2(n5360), .A3(data[142]), .A4(n5361), .Y(n203) );
  AO22X1_HVT U4515 ( .A1(\ram[7][176] ), .A2(n5398), .A3(n5399), .A4(data[176]), .Y(n2029) );
  AO22X1_HVT U4516 ( .A1(\ram[7][175] ), .A2(n5398), .A3(n5399), .A4(data[175]), .Y(n2028) );
  AO22X1_HVT U4517 ( .A1(\ram[7][174] ), .A2(n5398), .A3(n5399), .A4(data[174]), .Y(n2027) );
  AO22X1_HVT U4518 ( .A1(\ram[7][173] ), .A2(n5398), .A3(n5399), .A4(data[173]), .Y(n2026) );
  AO22X1_HVT U4519 ( .A1(\ram[7][172] ), .A2(n5398), .A3(n5399), .A4(data[172]), .Y(n2025) );
  AO22X1_HVT U4520 ( .A1(\ram[7][171] ), .A2(n5398), .A3(n5399), .A4(data[171]), .Y(n2024) );
  AO22X1_HVT U4521 ( .A1(\ram[7][170] ), .A2(n5398), .A3(n5399), .A4(data[170]), .Y(n2023) );
  AO22X1_HVT U4522 ( .A1(\ram[7][169] ), .A2(n5398), .A3(n5399), .A4(data[169]), .Y(n2022) );
  AO22X1_HVT U4523 ( .A1(\ram[7][168] ), .A2(n5398), .A3(n5399), .A4(data[168]), .Y(n2021) );
  AO22X1_HVT U4524 ( .A1(\ram[7][167] ), .A2(n5398), .A3(n5399), .A4(data[167]), .Y(n2020) );
  AO22X1_HVT U4525 ( .A1(\ram[0][141] ), .A2(n5360), .A3(data[141]), .A4(n5361), .Y(n202) );
  AO22X1_HVT U4526 ( .A1(\ram[7][166] ), .A2(n5398), .A3(n5399), .A4(data[166]), .Y(n2019) );
  AO22X1_HVT U4527 ( .A1(\ram[7][165] ), .A2(n5398), .A3(n5399), .A4(data[165]), .Y(n2018) );
  AO22X1_HVT U4528 ( .A1(\ram[7][164] ), .A2(n5398), .A3(n5399), .A4(data[164]), .Y(n2017) );
  AO22X1_HVT U4529 ( .A1(\ram[7][163] ), .A2(n5398), .A3(n5399), .A4(data[163]), .Y(n2016) );
  AO22X1_HVT U4530 ( .A1(\ram[7][162] ), .A2(n5398), .A3(n5399), .A4(data[162]), .Y(n2015) );
  AO22X1_HVT U4531 ( .A1(\ram[7][161] ), .A2(n5398), .A3(n5399), .A4(data[161]), .Y(n2014) );
  AO22X1_HVT U4532 ( .A1(\ram[7][160] ), .A2(n5398), .A3(n5399), .A4(data[160]), .Y(n2013) );
  AO22X1_HVT U4533 ( .A1(\ram[7][159] ), .A2(n5398), .A3(n5399), .A4(data[159]), .Y(n2012) );
  AO22X1_HVT U4534 ( .A1(\ram[7][158] ), .A2(n5398), .A3(n5399), .A4(data[158]), .Y(n2011) );
  AO22X1_HVT U4535 ( .A1(\ram[7][157] ), .A2(n5398), .A3(n5399), .A4(data[157]), .Y(n2010) );
  AO22X1_HVT U4536 ( .A1(\ram[0][140] ), .A2(n5360), .A3(data[140]), .A4(n5361), .Y(n201) );
  AO22X1_HVT U4537 ( .A1(\ram[7][156] ), .A2(n5398), .A3(n5399), .A4(data[156]), .Y(n2009) );
  AO22X1_HVT U4538 ( .A1(\ram[7][155] ), .A2(n5398), .A3(n5399), .A4(data[155]), .Y(n2008) );
  AO22X1_HVT U4539 ( .A1(\ram[7][154] ), .A2(n5398), .A3(n5399), .A4(data[154]), .Y(n2007) );
  AO22X1_HVT U4540 ( .A1(\ram[7][153] ), .A2(n5398), .A3(n5399), .A4(data[153]), .Y(n2006) );
  AO22X1_HVT U4541 ( .A1(\ram[7][152] ), .A2(n5398), .A3(n5399), .A4(data[152]), .Y(n2005) );
  AO22X1_HVT U4542 ( .A1(\ram[7][151] ), .A2(n5398), .A3(n5399), .A4(data[151]), .Y(n2004) );
  AO22X1_HVT U4543 ( .A1(\ram[7][150] ), .A2(n5398), .A3(n5399), .A4(data[150]), .Y(n2003) );
  AO22X1_HVT U4544 ( .A1(\ram[7][149] ), .A2(n5398), .A3(n5399), .A4(data[149]), .Y(n2002) );
  AO22X1_HVT U4545 ( .A1(\ram[7][148] ), .A2(n5398), .A3(n5399), .A4(data[148]), .Y(n2001) );
  AO22X1_HVT U4546 ( .A1(\ram[7][147] ), .A2(n5398), .A3(n5399), .A4(data[147]), .Y(n2000) );
  AO22X1_HVT U4547 ( .A1(\ram[0][139] ), .A2(n5360), .A3(data[139]), .A4(n5361), .Y(n200) );
  AO22X1_HVT U4548 ( .A1(\ram[7][146] ), .A2(n5398), .A3(n5399), .A4(data[146]), .Y(n1999) );
  AO22X1_HVT U4549 ( .A1(\ram[7][145] ), .A2(n5398), .A3(n5399), .A4(data[145]), .Y(n1998) );
  AO22X1_HVT U4550 ( .A1(\ram[7][144] ), .A2(n5398), .A3(n5399), .A4(data[144]), .Y(n1997) );
  AO22X1_HVT U4551 ( .A1(\ram[7][143] ), .A2(n5398), .A3(n5399), .A4(data[143]), .Y(n1996) );
  AO22X1_HVT U4552 ( .A1(\ram[7][142] ), .A2(n5398), .A3(n5399), .A4(data[142]), .Y(n1995) );
  AO22X1_HVT U4553 ( .A1(\ram[7][141] ), .A2(n5398), .A3(n5399), .A4(data[141]), .Y(n1994) );
  AO22X1_HVT U4554 ( .A1(\ram[7][140] ), .A2(n5398), .A3(n5399), .A4(data[140]), .Y(n1993) );
  AO22X1_HVT U4555 ( .A1(\ram[7][139] ), .A2(n5398), .A3(n5399), .A4(data[139]), .Y(n1992) );
  AO22X1_HVT U4556 ( .A1(\ram[7][138] ), .A2(n5398), .A3(n5399), .A4(data[138]), .Y(n1991) );
  AO22X1_HVT U4557 ( .A1(\ram[7][137] ), .A2(n5398), .A3(n5399), .A4(data[137]), .Y(n1990) );
  AO22X1_HVT U4558 ( .A1(\ram[0][138] ), .A2(n5360), .A3(data[138]), .A4(n5361), .Y(n199) );
  AO22X1_HVT U4559 ( .A1(\ram[7][136] ), .A2(n5398), .A3(n5399), .A4(data[136]), .Y(n1989) );
  AO22X1_HVT U4560 ( .A1(\ram[7][135] ), .A2(n5398), .A3(n5399), .A4(data[135]), .Y(n1988) );
  AO22X1_HVT U4561 ( .A1(\ram[7][134] ), .A2(n5398), .A3(n5399), .A4(data[134]), .Y(n1987) );
  AO22X1_HVT U4562 ( .A1(\ram[7][133] ), .A2(n5398), .A3(n5399), .A4(data[133]), .Y(n1986) );
  AO22X1_HVT U4563 ( .A1(\ram[7][132] ), .A2(n5398), .A3(n5399), .A4(data[132]), .Y(n1985) );
  AO22X1_HVT U4564 ( .A1(\ram[7][131] ), .A2(n5398), .A3(n5399), .A4(data[131]), .Y(n1984) );
  AO22X1_HVT U4565 ( .A1(\ram[7][130] ), .A2(n5398), .A3(n5399), .A4(data[130]), .Y(n1983) );
  AO22X1_HVT U4566 ( .A1(\ram[7][129] ), .A2(n5398), .A3(n5399), .A4(data[129]), .Y(n1982) );
  AO22X1_HVT U4567 ( .A1(\ram[7][128] ), .A2(n5398), .A3(n5399), .A4(data[128]), .Y(n1981) );
  AO22X1_HVT U4568 ( .A1(\ram[7][127] ), .A2(n5398), .A3(n5399), .A4(data[127]), .Y(n1980) );
  AO22X1_HVT U4569 ( .A1(\ram[0][137] ), .A2(n5360), .A3(data[137]), .A4(n5361), .Y(n198) );
  AO22X1_HVT U4570 ( .A1(\ram[7][126] ), .A2(n5398), .A3(n5399), .A4(data[126]), .Y(n1979) );
  AO22X1_HVT U4571 ( .A1(\ram[7][125] ), .A2(n5398), .A3(n5399), .A4(data[125]), .Y(n1978) );
  AO22X1_HVT U4572 ( .A1(\ram[7][124] ), .A2(n5398), .A3(n5399), .A4(data[124]), .Y(n1977) );
  AO22X1_HVT U4573 ( .A1(\ram[7][123] ), .A2(n5398), .A3(n5399), .A4(data[123]), .Y(n1976) );
  AO22X1_HVT U4574 ( .A1(\ram[7][122] ), .A2(n5398), .A3(n5399), .A4(data[122]), .Y(n1975) );
  AO22X1_HVT U4575 ( .A1(\ram[7][121] ), .A2(n5398), .A3(n5399), .A4(data[121]), .Y(n1974) );
  AO22X1_HVT U4576 ( .A1(\ram[7][120] ), .A2(n5398), .A3(n5399), .A4(data[120]), .Y(n1973) );
  AO22X1_HVT U4577 ( .A1(\ram[7][119] ), .A2(n5398), .A3(n5399), .A4(data[119]), .Y(n1972) );
  AO22X1_HVT U4578 ( .A1(\ram[7][118] ), .A2(n5398), .A3(n5399), .A4(data[118]), .Y(n1971) );
  AO22X1_HVT U4579 ( .A1(\ram[7][117] ), .A2(n5398), .A3(n5399), .A4(data[117]), .Y(n1970) );
  AO22X1_HVT U4580 ( .A1(\ram[0][136] ), .A2(n5360), .A3(data[136]), .A4(n5361), .Y(n197) );
  AO22X1_HVT U4581 ( .A1(\ram[7][116] ), .A2(n5398), .A3(n5399), .A4(data[116]), .Y(n1969) );
  AO22X1_HVT U4582 ( .A1(\ram[7][115] ), .A2(n5398), .A3(n5399), .A4(data[115]), .Y(n1968) );
  AO22X1_HVT U4583 ( .A1(\ram[7][114] ), .A2(n5398), .A3(n5399), .A4(data[114]), .Y(n1967) );
  AO22X1_HVT U4584 ( .A1(\ram[7][113] ), .A2(n5398), .A3(n5399), .A4(data[113]), .Y(n1966) );
  AO22X1_HVT U4585 ( .A1(\ram[7][112] ), .A2(n5398), .A3(n5399), .A4(data[112]), .Y(n1965) );
  AO22X1_HVT U4586 ( .A1(\ram[7][111] ), .A2(n5398), .A3(n5399), .A4(data[111]), .Y(n1964) );
  AO22X1_HVT U4587 ( .A1(\ram[7][110] ), .A2(n5398), .A3(n5399), .A4(data[110]), .Y(n1963) );
  AO22X1_HVT U4588 ( .A1(\ram[7][109] ), .A2(n5398), .A3(n5399), .A4(data[109]), .Y(n1962) );
  AO22X1_HVT U4589 ( .A1(\ram[7][108] ), .A2(n5398), .A3(n5399), .A4(data[108]), .Y(n1961) );
  AO22X1_HVT U4590 ( .A1(\ram[7][107] ), .A2(n5398), .A3(n5399), .A4(data[107]), .Y(n1960) );
  AO22X1_HVT U4591 ( .A1(\ram[0][135] ), .A2(n5360), .A3(data[135]), .A4(n5361), .Y(n196) );
  AO22X1_HVT U4592 ( .A1(\ram[7][106] ), .A2(n5398), .A3(n5399), .A4(data[106]), .Y(n1959) );
  AO22X1_HVT U4593 ( .A1(\ram[7][105] ), .A2(n5398), .A3(n5399), .A4(data[105]), .Y(n1958) );
  AO22X1_HVT U4594 ( .A1(\ram[7][104] ), .A2(n5398), .A3(n5399), .A4(data[104]), .Y(n1957) );
  AO22X1_HVT U4595 ( .A1(\ram[7][103] ), .A2(n5398), .A3(n5399), .A4(data[103]), .Y(n1956) );
  AO22X1_HVT U4596 ( .A1(\ram[7][102] ), .A2(n5398), .A3(n5399), .A4(data[102]), .Y(n1955) );
  AO22X1_HVT U4597 ( .A1(\ram[7][101] ), .A2(n5398), .A3(n5399), .A4(data[101]), .Y(n1954) );
  AO22X1_HVT U4598 ( .A1(\ram[7][100] ), .A2(n5398), .A3(n5399), .A4(data[100]), .Y(n1953) );
  AO22X1_HVT U4599 ( .A1(\ram[7][99] ), .A2(n5398), .A3(n5399), .A4(data[99]), 
        .Y(n1952) );
  AO22X1_HVT U4600 ( .A1(\ram[7][98] ), .A2(n5398), .A3(n5399), .A4(data[98]), 
        .Y(n1951) );
  AO22X1_HVT U4601 ( .A1(\ram[7][97] ), .A2(n5398), .A3(n5399), .A4(data[97]), 
        .Y(n1950) );
  AO22X1_HVT U4602 ( .A1(\ram[0][134] ), .A2(n5360), .A3(data[134]), .A4(n5361), .Y(n195) );
  AO22X1_HVT U4603 ( .A1(\ram[7][96] ), .A2(n5398), .A3(n5399), .A4(data[96]), 
        .Y(n1949) );
  AO22X1_HVT U4604 ( .A1(\ram[7][95] ), .A2(n5398), .A3(n5399), .A4(data[95]), 
        .Y(n1948) );
  AO22X1_HVT U4605 ( .A1(\ram[7][94] ), .A2(n5398), .A3(n5399), .A4(data[94]), 
        .Y(n1947) );
  AO22X1_HVT U4606 ( .A1(\ram[7][93] ), .A2(n5398), .A3(n5399), .A4(data[93]), 
        .Y(n1946) );
  AO22X1_HVT U4607 ( .A1(\ram[7][92] ), .A2(n5398), .A3(n5399), .A4(data[92]), 
        .Y(n1945) );
  AO22X1_HVT U4608 ( .A1(\ram[7][91] ), .A2(n5398), .A3(n5399), .A4(data[91]), 
        .Y(n1944) );
  AO22X1_HVT U4609 ( .A1(\ram[7][90] ), .A2(n5398), .A3(n5399), .A4(data[90]), 
        .Y(n1943) );
  AO22X1_HVT U4610 ( .A1(\ram[7][89] ), .A2(n5398), .A3(n5399), .A4(data[89]), 
        .Y(n1942) );
  AO22X1_HVT U4611 ( .A1(\ram[7][88] ), .A2(n5398), .A3(n5399), .A4(data[88]), 
        .Y(n1941) );
  AO22X1_HVT U4612 ( .A1(\ram[7][87] ), .A2(n5398), .A3(n5399), .A4(data[87]), 
        .Y(n1940) );
  AO22X1_HVT U4613 ( .A1(\ram[0][133] ), .A2(n5360), .A3(data[133]), .A4(n5361), .Y(n194) );
  AO22X1_HVT U4614 ( .A1(\ram[7][86] ), .A2(n5398), .A3(n5399), .A4(data[86]), 
        .Y(n1939) );
  AO22X1_HVT U4615 ( .A1(\ram[7][85] ), .A2(n5398), .A3(n5399), .A4(data[85]), 
        .Y(n1938) );
  AO22X1_HVT U4616 ( .A1(\ram[7][84] ), .A2(n5398), .A3(n5399), .A4(data[84]), 
        .Y(n1937) );
  AO22X1_HVT U4617 ( .A1(\ram[7][83] ), .A2(n5398), .A3(n5399), .A4(data[83]), 
        .Y(n1936) );
  AO22X1_HVT U4618 ( .A1(\ram[7][82] ), .A2(n5398), .A3(n5399), .A4(data[82]), 
        .Y(n1935) );
  AO22X1_HVT U4619 ( .A1(\ram[7][81] ), .A2(n5398), .A3(n5399), .A4(data[81]), 
        .Y(n1934) );
  AO22X1_HVT U4620 ( .A1(\ram[7][80] ), .A2(n5398), .A3(n5399), .A4(data[80]), 
        .Y(n1933) );
  AO22X1_HVT U4621 ( .A1(\ram[7][79] ), .A2(n5398), .A3(n5399), .A4(data[79]), 
        .Y(n1932) );
  AO22X1_HVT U4622 ( .A1(\ram[7][78] ), .A2(n5398), .A3(n5399), .A4(data[78]), 
        .Y(n1931) );
  AO22X1_HVT U4623 ( .A1(\ram[7][77] ), .A2(n5398), .A3(n5399), .A4(data[77]), 
        .Y(n1930) );
  AO22X1_HVT U4624 ( .A1(\ram[0][132] ), .A2(n5360), .A3(data[132]), .A4(n5361), .Y(n193) );
  AO22X1_HVT U4625 ( .A1(\ram[7][76] ), .A2(n5398), .A3(n5399), .A4(data[76]), 
        .Y(n1929) );
  AO22X1_HVT U4626 ( .A1(\ram[7][75] ), .A2(n5398), .A3(n5399), .A4(data[75]), 
        .Y(n1928) );
  AO22X1_HVT U4627 ( .A1(\ram[7][74] ), .A2(n5398), .A3(n5399), .A4(data[74]), 
        .Y(n1927) );
  AO22X1_HVT U4628 ( .A1(\ram[7][73] ), .A2(n5398), .A3(n5399), .A4(data[73]), 
        .Y(n1926) );
  AO22X1_HVT U4629 ( .A1(\ram[7][72] ), .A2(n5398), .A3(n5399), .A4(data[72]), 
        .Y(n1925) );
  AO22X1_HVT U4630 ( .A1(\ram[7][71] ), .A2(n5398), .A3(n5399), .A4(data[71]), 
        .Y(n1924) );
  AO22X1_HVT U4631 ( .A1(\ram[7][70] ), .A2(n5398), .A3(n5399), .A4(data[70]), 
        .Y(n1923) );
  AO22X1_HVT U4632 ( .A1(\ram[7][69] ), .A2(n5398), .A3(n5399), .A4(data[69]), 
        .Y(n1922) );
  AO22X1_HVT U4633 ( .A1(\ram[7][68] ), .A2(n5398), .A3(n5399), .A4(data[68]), 
        .Y(n1921) );
  AO22X1_HVT U4634 ( .A1(\ram[7][67] ), .A2(n5398), .A3(n5399), .A4(data[67]), 
        .Y(n1920) );
  AO22X1_HVT U4635 ( .A1(\ram[0][131] ), .A2(n5360), .A3(data[131]), .A4(n5361), .Y(n192) );
  AO22X1_HVT U4636 ( .A1(\ram[7][66] ), .A2(n5398), .A3(n5399), .A4(data[66]), 
        .Y(n1919) );
  AO22X1_HVT U4637 ( .A1(\ram[7][65] ), .A2(n5398), .A3(n5399), .A4(data[65]), 
        .Y(n1918) );
  AO22X1_HVT U4638 ( .A1(\ram[7][64] ), .A2(n5398), .A3(n5399), .A4(data[64]), 
        .Y(n1917) );
  AO22X1_HVT U4639 ( .A1(\ram[7][63] ), .A2(n5398), .A3(n5399), .A4(data[63]), 
        .Y(n1916) );
  AO22X1_HVT U4640 ( .A1(\ram[7][62] ), .A2(n5398), .A3(n5399), .A4(data[62]), 
        .Y(n1915) );
  AO22X1_HVT U4641 ( .A1(\ram[7][61] ), .A2(n5398), .A3(n5399), .A4(data[61]), 
        .Y(n1914) );
  AO22X1_HVT U4642 ( .A1(\ram[7][60] ), .A2(n5398), .A3(n5399), .A4(data[60]), 
        .Y(n1913) );
  AO22X1_HVT U4643 ( .A1(\ram[7][59] ), .A2(n5398), .A3(n5399), .A4(data[59]), 
        .Y(n1912) );
  AO22X1_HVT U4644 ( .A1(\ram[7][58] ), .A2(n5398), .A3(n5399), .A4(data[58]), 
        .Y(n1911) );
  AO22X1_HVT U4645 ( .A1(\ram[7][57] ), .A2(n5398), .A3(n5399), .A4(data[57]), 
        .Y(n1910) );
  AO22X1_HVT U4646 ( .A1(\ram[0][130] ), .A2(n5360), .A3(data[130]), .A4(n5361), .Y(n191) );
  AO22X1_HVT U4647 ( .A1(\ram[7][56] ), .A2(n5398), .A3(n5399), .A4(data[56]), 
        .Y(n1909) );
  AO22X1_HVT U4648 ( .A1(\ram[7][55] ), .A2(n5398), .A3(n5399), .A4(data[55]), 
        .Y(n1908) );
  AO22X1_HVT U4649 ( .A1(\ram[7][54] ), .A2(n5398), .A3(n5399), .A4(data[54]), 
        .Y(n1907) );
  AO22X1_HVT U4650 ( .A1(\ram[7][53] ), .A2(n5398), .A3(n5399), .A4(data[53]), 
        .Y(n1906) );
  AO22X1_HVT U4651 ( .A1(\ram[7][52] ), .A2(n5398), .A3(n5399), .A4(data[52]), 
        .Y(n1905) );
  AO22X1_HVT U4652 ( .A1(\ram[7][51] ), .A2(n5398), .A3(n5399), .A4(data[51]), 
        .Y(n1904) );
  AO22X1_HVT U4653 ( .A1(\ram[7][50] ), .A2(n5398), .A3(n5399), .A4(data[50]), 
        .Y(n1903) );
  AO22X1_HVT U4654 ( .A1(\ram[7][49] ), .A2(n5398), .A3(n5399), .A4(data[49]), 
        .Y(n1902) );
  AO22X1_HVT U4655 ( .A1(\ram[7][48] ), .A2(n5398), .A3(n5399), .A4(data[48]), 
        .Y(n1901) );
  AO22X1_HVT U4656 ( .A1(\ram[7][47] ), .A2(n5398), .A3(n5399), .A4(data[47]), 
        .Y(n1900) );
  AO22X1_HVT U4657 ( .A1(\ram[0][129] ), .A2(n5360), .A3(data[129]), .A4(n5361), .Y(n190) );
  AO22X1_HVT U4658 ( .A1(\ram[7][46] ), .A2(n5398), .A3(n5399), .A4(data[46]), 
        .Y(n1899) );
  AO22X1_HVT U4659 ( .A1(\ram[7][45] ), .A2(n5398), .A3(n5399), .A4(data[45]), 
        .Y(n1898) );
  AO22X1_HVT U4660 ( .A1(\ram[7][44] ), .A2(n5398), .A3(n5399), .A4(data[44]), 
        .Y(n1897) );
  AO22X1_HVT U4661 ( .A1(\ram[7][43] ), .A2(n5398), .A3(n5399), .A4(data[43]), 
        .Y(n1896) );
  AO22X1_HVT U4662 ( .A1(\ram[7][42] ), .A2(n5398), .A3(n5399), .A4(data[42]), 
        .Y(n1895) );
  AO22X1_HVT U4663 ( .A1(\ram[7][41] ), .A2(n5398), .A3(n5399), .A4(data[41]), 
        .Y(n1894) );
  AO22X1_HVT U4664 ( .A1(\ram[7][40] ), .A2(n5398), .A3(n5399), .A4(data[40]), 
        .Y(n1893) );
  AO22X1_HVT U4665 ( .A1(\ram[7][39] ), .A2(n5398), .A3(n5399), .A4(data[39]), 
        .Y(n1892) );
  AO22X1_HVT U4666 ( .A1(\ram[7][38] ), .A2(n5398), .A3(n5399), .A4(data[38]), 
        .Y(n1891) );
  AO22X1_HVT U4667 ( .A1(\ram[7][37] ), .A2(n5398), .A3(n5399), .A4(data[37]), 
        .Y(n1890) );
  AO22X1_HVT U4668 ( .A1(\ram[0][128] ), .A2(n5360), .A3(data[128]), .A4(n5361), .Y(n189) );
  AO22X1_HVT U4669 ( .A1(\ram[7][36] ), .A2(n5398), .A3(n5399), .A4(data[36]), 
        .Y(n1889) );
  AO22X1_HVT U4670 ( .A1(\ram[7][35] ), .A2(n5398), .A3(n5399), .A4(data[35]), 
        .Y(n1888) );
  AO22X1_HVT U4671 ( .A1(\ram[7][34] ), .A2(n5398), .A3(n5399), .A4(data[34]), 
        .Y(n1887) );
  AO22X1_HVT U4672 ( .A1(\ram[7][33] ), .A2(n5398), .A3(n5399), .A4(data[33]), 
        .Y(n1886) );
  AO22X1_HVT U4673 ( .A1(\ram[7][32] ), .A2(n5398), .A3(n5399), .A4(data[32]), 
        .Y(n1885) );
  AO22X1_HVT U4674 ( .A1(\ram[7][31] ), .A2(n5398), .A3(n5399), .A4(data[31]), 
        .Y(n1884) );
  AO22X1_HVT U4675 ( .A1(\ram[7][30] ), .A2(n5398), .A3(n5399), .A4(data[30]), 
        .Y(n1883) );
  AO22X1_HVT U4676 ( .A1(\ram[7][29] ), .A2(n5398), .A3(n5399), .A4(data[29]), 
        .Y(n1882) );
  AO22X1_HVT U4677 ( .A1(\ram[7][28] ), .A2(n5398), .A3(n5399), .A4(data[28]), 
        .Y(n1881) );
  AO22X1_HVT U4678 ( .A1(\ram[7][27] ), .A2(n5398), .A3(n5399), .A4(data[27]), 
        .Y(n1880) );
  AO22X1_HVT U4679 ( .A1(\ram[0][127] ), .A2(n5360), .A3(data[127]), .A4(n5361), .Y(n188) );
  AO22X1_HVT U4680 ( .A1(\ram[7][26] ), .A2(n5398), .A3(n5399), .A4(data[26]), 
        .Y(n1879) );
  AO22X1_HVT U4681 ( .A1(\ram[7][25] ), .A2(n5398), .A3(n5399), .A4(data[25]), 
        .Y(n1878) );
  AO22X1_HVT U4682 ( .A1(\ram[7][24] ), .A2(n5398), .A3(n5399), .A4(data[24]), 
        .Y(n1877) );
  AO22X1_HVT U4683 ( .A1(\ram[7][23] ), .A2(n5398), .A3(n5399), .A4(data[23]), 
        .Y(n1876) );
  AO22X1_HVT U4684 ( .A1(\ram[7][22] ), .A2(n5398), .A3(n5399), .A4(data[22]), 
        .Y(n1875) );
  AO22X1_HVT U4685 ( .A1(\ram[7][21] ), .A2(n5398), .A3(n5399), .A4(data[21]), 
        .Y(n1874) );
  AO22X1_HVT U4686 ( .A1(\ram[7][20] ), .A2(n5398), .A3(n5399), .A4(data[20]), 
        .Y(n1873) );
  AO22X1_HVT U4687 ( .A1(\ram[7][19] ), .A2(n5398), .A3(n5399), .A4(data[19]), 
        .Y(n1872) );
  AO22X1_HVT U4688 ( .A1(\ram[7][18] ), .A2(n5398), .A3(n5399), .A4(data[18]), 
        .Y(n1871) );
  AO22X1_HVT U4689 ( .A1(\ram[7][17] ), .A2(n5398), .A3(n5399), .A4(data[17]), 
        .Y(n1870) );
  AO22X1_HVT U4690 ( .A1(\ram[0][126] ), .A2(n5360), .A3(data[126]), .A4(n5361), .Y(n187) );
  AO22X1_HVT U4691 ( .A1(\ram[7][16] ), .A2(n5398), .A3(n5399), .A4(data[16]), 
        .Y(n1869) );
  AO22X1_HVT U4692 ( .A1(\ram[7][15] ), .A2(n5398), .A3(n5399), .A4(data[15]), 
        .Y(n1868) );
  AO22X1_HVT U4693 ( .A1(\ram[7][14] ), .A2(n5398), .A3(n5399), .A4(data[14]), 
        .Y(n1867) );
  AO22X1_HVT U4694 ( .A1(\ram[7][13] ), .A2(n5398), .A3(n5399), .A4(data[13]), 
        .Y(n1866) );
  AO22X1_HVT U4695 ( .A1(\ram[7][12] ), .A2(n5398), .A3(n5399), .A4(data[12]), 
        .Y(n1865) );
  AO22X1_HVT U4696 ( .A1(\ram[7][11] ), .A2(n5398), .A3(n5399), .A4(data[11]), 
        .Y(n1864) );
  AO22X1_HVT U4697 ( .A1(\ram[7][10] ), .A2(n5398), .A3(n5399), .A4(data[10]), 
        .Y(n1863) );
  AO22X1_HVT U4698 ( .A1(\ram[7][9] ), .A2(n5398), .A3(n5399), .A4(data[9]), 
        .Y(n1862) );
  AO22X1_HVT U4699 ( .A1(\ram[7][8] ), .A2(n5398), .A3(n5399), .A4(data[8]), 
        .Y(n1861) );
  AO22X1_HVT U4700 ( .A1(\ram[7][7] ), .A2(n5398), .A3(n5399), .A4(data[7]), 
        .Y(n1860) );
  AO22X1_HVT U4701 ( .A1(\ram[0][125] ), .A2(n5360), .A3(data[125]), .A4(n5361), .Y(n186) );
  AO22X1_HVT U4702 ( .A1(\ram[7][6] ), .A2(n5398), .A3(n5399), .A4(data[6]), 
        .Y(n1859) );
  AO22X1_HVT U4703 ( .A1(\ram[7][5] ), .A2(n5398), .A3(n5399), .A4(data[5]), 
        .Y(n1858) );
  AO22X1_HVT U4704 ( .A1(\ram[7][4] ), .A2(n5398), .A3(n5399), .A4(data[4]), 
        .Y(n1857) );
  AO22X1_HVT U4705 ( .A1(\ram[7][3] ), .A2(n5398), .A3(n5399), .A4(data[3]), 
        .Y(n1856) );
  AO22X1_HVT U4706 ( .A1(\ram[7][2] ), .A2(n5398), .A3(n5399), .A4(data[2]), 
        .Y(n1855) );
  AO22X1_HVT U4707 ( .A1(\ram[7][1] ), .A2(n5398), .A3(n5399), .A4(data[1]), 
        .Y(n1854) );
  AO22X1_HVT U4708 ( .A1(\ram[7][0] ), .A2(n5398), .A3(n5399), .A4(data[0]), 
        .Y(n1853) );
  INVX0_HVT U4709 ( .A(n5400), .Y(n5399) );
  AND2X1_HVT U4710 ( .A1(n5400), .A2(n5365), .Y(n5398) );
  NAND3X0_HVT U4711 ( .A1(n4182), .A2(n4276), .A3(n5401), .Y(n5400) );
  AO22X1_HVT U4712 ( .A1(\ram[6][255] ), .A2(n5402), .A3(n5403), .A4(data[255]), .Y(n1852) );
  AO22X1_HVT U4713 ( .A1(\ram[6][254] ), .A2(n5402), .A3(n5403), .A4(data[254]), .Y(n1851) );
  AO22X1_HVT U4714 ( .A1(\ram[6][253] ), .A2(n5402), .A3(n5403), .A4(data[253]), .Y(n1850) );
  AO22X1_HVT U4715 ( .A1(\ram[0][124] ), .A2(n5360), .A3(data[124]), .A4(n5361), .Y(n185) );
  AO22X1_HVT U4716 ( .A1(\ram[6][252] ), .A2(n5402), .A3(n5403), .A4(data[252]), .Y(n1849) );
  AO22X1_HVT U4717 ( .A1(\ram[6][251] ), .A2(n5402), .A3(n5403), .A4(data[251]), .Y(n1848) );
  AO22X1_HVT U4718 ( .A1(\ram[6][250] ), .A2(n5402), .A3(n5403), .A4(data[250]), .Y(n1847) );
  AO22X1_HVT U4719 ( .A1(\ram[6][249] ), .A2(n5402), .A3(n5403), .A4(data[249]), .Y(n1846) );
  AO22X1_HVT U4720 ( .A1(\ram[6][248] ), .A2(n5402), .A3(n5403), .A4(data[248]), .Y(n1845) );
  AO22X1_HVT U4721 ( .A1(\ram[6][247] ), .A2(n5402), .A3(n5403), .A4(data[247]), .Y(n1844) );
  AO22X1_HVT U4722 ( .A1(\ram[6][246] ), .A2(n5402), .A3(n5403), .A4(data[246]), .Y(n1843) );
  AO22X1_HVT U4723 ( .A1(\ram[6][245] ), .A2(n5402), .A3(n5403), .A4(data[245]), .Y(n1842) );
  AO22X1_HVT U4724 ( .A1(\ram[6][244] ), .A2(n5402), .A3(n5403), .A4(data[244]), .Y(n1841) );
  AO22X1_HVT U4725 ( .A1(\ram[6][243] ), .A2(n5402), .A3(n5403), .A4(data[243]), .Y(n1840) );
  AO22X1_HVT U4726 ( .A1(\ram[0][123] ), .A2(n5360), .A3(data[123]), .A4(n5361), .Y(n184) );
  AO22X1_HVT U4727 ( .A1(\ram[6][242] ), .A2(n5402), .A3(n5403), .A4(data[242]), .Y(n1839) );
  AO22X1_HVT U4728 ( .A1(\ram[6][241] ), .A2(n5402), .A3(n5403), .A4(data[241]), .Y(n1838) );
  AO22X1_HVT U4729 ( .A1(\ram[6][240] ), .A2(n5402), .A3(n5403), .A4(data[240]), .Y(n1837) );
  AO22X1_HVT U4730 ( .A1(\ram[6][239] ), .A2(n5402), .A3(n5403), .A4(data[239]), .Y(n1836) );
  AO22X1_HVT U4731 ( .A1(\ram[6][238] ), .A2(n5402), .A3(n5403), .A4(data[238]), .Y(n1835) );
  AO22X1_HVT U4732 ( .A1(\ram[6][237] ), .A2(n5402), .A3(n5403), .A4(data[237]), .Y(n1834) );
  AO22X1_HVT U4733 ( .A1(\ram[6][236] ), .A2(n5402), .A3(n5403), .A4(data[236]), .Y(n1833) );
  AO22X1_HVT U4734 ( .A1(\ram[6][235] ), .A2(n5402), .A3(n5403), .A4(data[235]), .Y(n1832) );
  AO22X1_HVT U4735 ( .A1(\ram[6][234] ), .A2(n5402), .A3(n5403), .A4(data[234]), .Y(n1831) );
  AO22X1_HVT U4736 ( .A1(\ram[6][233] ), .A2(n5402), .A3(n5403), .A4(data[233]), .Y(n1830) );
  AO22X1_HVT U4737 ( .A1(\ram[0][122] ), .A2(n5360), .A3(data[122]), .A4(n5361), .Y(n183) );
  AO22X1_HVT U4738 ( .A1(\ram[6][232] ), .A2(n5402), .A3(n5403), .A4(data[232]), .Y(n1829) );
  AO22X1_HVT U4739 ( .A1(\ram[6][231] ), .A2(n5402), .A3(n5403), .A4(data[231]), .Y(n1828) );
  AO22X1_HVT U4740 ( .A1(\ram[6][230] ), .A2(n5402), .A3(n5403), .A4(data[230]), .Y(n1827) );
  AO22X1_HVT U4741 ( .A1(\ram[6][229] ), .A2(n5402), .A3(n5403), .A4(data[229]), .Y(n1826) );
  AO22X1_HVT U4742 ( .A1(\ram[6][228] ), .A2(n5402), .A3(n5403), .A4(data[228]), .Y(n1825) );
  AO22X1_HVT U4743 ( .A1(\ram[6][227] ), .A2(n5402), .A3(n5403), .A4(data[227]), .Y(n1824) );
  AO22X1_HVT U4744 ( .A1(\ram[6][226] ), .A2(n5402), .A3(n5403), .A4(data[226]), .Y(n1823) );
  AO22X1_HVT U4745 ( .A1(\ram[6][225] ), .A2(n5402), .A3(n5403), .A4(data[225]), .Y(n1822) );
  AO22X1_HVT U4746 ( .A1(\ram[6][224] ), .A2(n5402), .A3(n5403), .A4(data[224]), .Y(n1821) );
  AO22X1_HVT U4747 ( .A1(\ram[6][223] ), .A2(n5402), .A3(n5403), .A4(data[223]), .Y(n1820) );
  AO22X1_HVT U4748 ( .A1(\ram[0][121] ), .A2(n5360), .A3(data[121]), .A4(n5361), .Y(n182) );
  AO22X1_HVT U4749 ( .A1(\ram[6][222] ), .A2(n5402), .A3(n5403), .A4(data[222]), .Y(n1819) );
  AO22X1_HVT U4750 ( .A1(\ram[6][221] ), .A2(n5402), .A3(n5403), .A4(data[221]), .Y(n1818) );
  AO22X1_HVT U4751 ( .A1(\ram[6][220] ), .A2(n5402), .A3(n5403), .A4(data[220]), .Y(n1817) );
  AO22X1_HVT U4752 ( .A1(\ram[6][219] ), .A2(n5402), .A3(n5403), .A4(data[219]), .Y(n1816) );
  AO22X1_HVT U4753 ( .A1(\ram[6][218] ), .A2(n5402), .A3(n5403), .A4(data[218]), .Y(n1815) );
  AO22X1_HVT U4754 ( .A1(\ram[6][217] ), .A2(n5402), .A3(n5403), .A4(data[217]), .Y(n1814) );
  AO22X1_HVT U4755 ( .A1(\ram[6][216] ), .A2(n5402), .A3(n5403), .A4(data[216]), .Y(n1813) );
  AO22X1_HVT U4756 ( .A1(\ram[6][215] ), .A2(n5402), .A3(n5403), .A4(data[215]), .Y(n1812) );
  AO22X1_HVT U4757 ( .A1(\ram[6][214] ), .A2(n5402), .A3(n5403), .A4(data[214]), .Y(n1811) );
  AO22X1_HVT U4758 ( .A1(\ram[6][213] ), .A2(n5402), .A3(n5403), .A4(data[213]), .Y(n1810) );
  AO22X1_HVT U4759 ( .A1(\ram[0][120] ), .A2(n5360), .A3(data[120]), .A4(n5361), .Y(n181) );
  AO22X1_HVT U4760 ( .A1(\ram[6][212] ), .A2(n5402), .A3(n5403), .A4(data[212]), .Y(n1809) );
  AO22X1_HVT U4761 ( .A1(\ram[6][211] ), .A2(n5402), .A3(n5403), .A4(data[211]), .Y(n1808) );
  AO22X1_HVT U4762 ( .A1(\ram[6][210] ), .A2(n5402), .A3(n5403), .A4(data[210]), .Y(n1807) );
  AO22X1_HVT U4763 ( .A1(\ram[6][209] ), .A2(n5402), .A3(n5403), .A4(data[209]), .Y(n1806) );
  AO22X1_HVT U4764 ( .A1(\ram[6][208] ), .A2(n5402), .A3(n5403), .A4(data[208]), .Y(n1805) );
  AO22X1_HVT U4765 ( .A1(\ram[6][207] ), .A2(n5402), .A3(n5403), .A4(data[207]), .Y(n1804) );
  AO22X1_HVT U4766 ( .A1(\ram[6][206] ), .A2(n5402), .A3(n5403), .A4(data[206]), .Y(n1803) );
  AO22X1_HVT U4767 ( .A1(\ram[6][205] ), .A2(n5402), .A3(n5403), .A4(data[205]), .Y(n1802) );
  AO22X1_HVT U4768 ( .A1(\ram[6][204] ), .A2(n5402), .A3(n5403), .A4(data[204]), .Y(n1801) );
  AO22X1_HVT U4769 ( .A1(\ram[6][203] ), .A2(n5402), .A3(n5403), .A4(data[203]), .Y(n1800) );
  AO22X1_HVT U4770 ( .A1(\ram[0][119] ), .A2(n5360), .A3(data[119]), .A4(n5361), .Y(n180) );
  AO22X1_HVT U4771 ( .A1(\ram[6][202] ), .A2(n5402), .A3(n5403), .A4(data[202]), .Y(n1799) );
  AO22X1_HVT U4772 ( .A1(\ram[6][201] ), .A2(n5402), .A3(n5403), .A4(data[201]), .Y(n1798) );
  AO22X1_HVT U4773 ( .A1(\ram[6][200] ), .A2(n5402), .A3(n5403), .A4(data[200]), .Y(n1797) );
  AO22X1_HVT U4774 ( .A1(\ram[6][199] ), .A2(n5402), .A3(n5403), .A4(data[199]), .Y(n1796) );
  AO22X1_HVT U4775 ( .A1(\ram[6][198] ), .A2(n5402), .A3(n5403), .A4(data[198]), .Y(n1795) );
  AO22X1_HVT U4776 ( .A1(\ram[6][197] ), .A2(n5402), .A3(n5403), .A4(data[197]), .Y(n1794) );
  AO22X1_HVT U4777 ( .A1(\ram[6][196] ), .A2(n5402), .A3(n5403), .A4(data[196]), .Y(n1793) );
  AO22X1_HVT U4778 ( .A1(\ram[6][195] ), .A2(n5402), .A3(n5403), .A4(data[195]), .Y(n1792) );
  AO22X1_HVT U4779 ( .A1(\ram[6][194] ), .A2(n5402), .A3(n5403), .A4(data[194]), .Y(n1791) );
  AO22X1_HVT U4780 ( .A1(\ram[6][193] ), .A2(n5402), .A3(n5403), .A4(data[193]), .Y(n1790) );
  AO22X1_HVT U4781 ( .A1(\ram[0][118] ), .A2(n5360), .A3(data[118]), .A4(n5361), .Y(n179) );
  AO22X1_HVT U4782 ( .A1(\ram[6][192] ), .A2(n5402), .A3(n5403), .A4(data[192]), .Y(n1789) );
  AO22X1_HVT U4783 ( .A1(\ram[6][191] ), .A2(n5402), .A3(n5403), .A4(data[191]), .Y(n1788) );
  AO22X1_HVT U4784 ( .A1(\ram[6][190] ), .A2(n5402), .A3(n5403), .A4(data[190]), .Y(n1787) );
  AO22X1_HVT U4785 ( .A1(\ram[6][189] ), .A2(n5402), .A3(n5403), .A4(data[189]), .Y(n1786) );
  AO22X1_HVT U4786 ( .A1(\ram[6][188] ), .A2(n5402), .A3(n5403), .A4(data[188]), .Y(n1785) );
  AO22X1_HVT U4787 ( .A1(\ram[6][187] ), .A2(n5402), .A3(n5403), .A4(data[187]), .Y(n1784) );
  AO22X1_HVT U4788 ( .A1(\ram[6][186] ), .A2(n5402), .A3(n5403), .A4(data[186]), .Y(n1783) );
  AO22X1_HVT U4789 ( .A1(\ram[6][185] ), .A2(n5402), .A3(n5403), .A4(data[185]), .Y(n1782) );
  AO22X1_HVT U4790 ( .A1(\ram[6][184] ), .A2(n5402), .A3(n5403), .A4(data[184]), .Y(n1781) );
  AO22X1_HVT U4791 ( .A1(\ram[6][183] ), .A2(n5402), .A3(n5403), .A4(data[183]), .Y(n1780) );
  AO22X1_HVT U4792 ( .A1(\ram[0][117] ), .A2(n5360), .A3(data[117]), .A4(n5361), .Y(n178) );
  AO22X1_HVT U4793 ( .A1(\ram[6][182] ), .A2(n5402), .A3(n5403), .A4(data[182]), .Y(n1779) );
  AO22X1_HVT U4794 ( .A1(\ram[6][181] ), .A2(n5402), .A3(n5403), .A4(data[181]), .Y(n1778) );
  AO22X1_HVT U4795 ( .A1(\ram[6][180] ), .A2(n5402), .A3(n5403), .A4(data[180]), .Y(n1777) );
  AO22X1_HVT U4796 ( .A1(\ram[6][179] ), .A2(n5402), .A3(n5403), .A4(data[179]), .Y(n1776) );
  AO22X1_HVT U4797 ( .A1(\ram[6][178] ), .A2(n5402), .A3(n5403), .A4(data[178]), .Y(n1775) );
  AO22X1_HVT U4798 ( .A1(\ram[6][177] ), .A2(n5402), .A3(n5403), .A4(data[177]), .Y(n1774) );
  AO22X1_HVT U4799 ( .A1(\ram[6][176] ), .A2(n5402), .A3(n5403), .A4(data[176]), .Y(n1773) );
  AO22X1_HVT U4800 ( .A1(\ram[6][175] ), .A2(n5402), .A3(n5403), .A4(data[175]), .Y(n1772) );
  AO22X1_HVT U4801 ( .A1(\ram[6][174] ), .A2(n5402), .A3(n5403), .A4(data[174]), .Y(n1771) );
  AO22X1_HVT U4802 ( .A1(\ram[6][173] ), .A2(n5402), .A3(n5403), .A4(data[173]), .Y(n1770) );
  AO22X1_HVT U4803 ( .A1(\ram[0][116] ), .A2(n5360), .A3(data[116]), .A4(n5361), .Y(n177) );
  AO22X1_HVT U4804 ( .A1(\ram[6][172] ), .A2(n5402), .A3(n5403), .A4(data[172]), .Y(n1769) );
  AO22X1_HVT U4805 ( .A1(\ram[6][171] ), .A2(n5402), .A3(n5403), .A4(data[171]), .Y(n1768) );
  AO22X1_HVT U4806 ( .A1(\ram[6][170] ), .A2(n5402), .A3(n5403), .A4(data[170]), .Y(n1767) );
  AO22X1_HVT U4807 ( .A1(\ram[6][169] ), .A2(n5402), .A3(n5403), .A4(data[169]), .Y(n1766) );
  AO22X1_HVT U4808 ( .A1(\ram[6][168] ), .A2(n5402), .A3(n5403), .A4(data[168]), .Y(n1765) );
  AO22X1_HVT U4809 ( .A1(\ram[6][167] ), .A2(n5402), .A3(n5403), .A4(data[167]), .Y(n1764) );
  AO22X1_HVT U4810 ( .A1(\ram[6][166] ), .A2(n5402), .A3(n5403), .A4(data[166]), .Y(n1763) );
  AO22X1_HVT U4811 ( .A1(\ram[6][165] ), .A2(n5402), .A3(n5403), .A4(data[165]), .Y(n1762) );
  AO22X1_HVT U4812 ( .A1(\ram[6][164] ), .A2(n5402), .A3(n5403), .A4(data[164]), .Y(n1761) );
  AO22X1_HVT U4813 ( .A1(\ram[6][163] ), .A2(n5402), .A3(n5403), .A4(data[163]), .Y(n1760) );
  AO22X1_HVT U4814 ( .A1(\ram[0][115] ), .A2(n5360), .A3(data[115]), .A4(n5361), .Y(n176) );
  AO22X1_HVT U4815 ( .A1(\ram[6][162] ), .A2(n5402), .A3(n5403), .A4(data[162]), .Y(n1759) );
  AO22X1_HVT U4816 ( .A1(\ram[6][161] ), .A2(n5402), .A3(n5403), .A4(data[161]), .Y(n1758) );
  AO22X1_HVT U4817 ( .A1(\ram[6][160] ), .A2(n5402), .A3(n5403), .A4(data[160]), .Y(n1757) );
  AO22X1_HVT U4818 ( .A1(\ram[6][159] ), .A2(n5402), .A3(n5403), .A4(data[159]), .Y(n1756) );
  AO22X1_HVT U4819 ( .A1(\ram[6][158] ), .A2(n5402), .A3(n5403), .A4(data[158]), .Y(n1755) );
  AO22X1_HVT U4820 ( .A1(\ram[6][157] ), .A2(n5402), .A3(n5403), .A4(data[157]), .Y(n1754) );
  AO22X1_HVT U4821 ( .A1(\ram[6][156] ), .A2(n5402), .A3(n5403), .A4(data[156]), .Y(n1753) );
  AO22X1_HVT U4822 ( .A1(\ram[6][155] ), .A2(n5402), .A3(n5403), .A4(data[155]), .Y(n1752) );
  AO22X1_HVT U4823 ( .A1(\ram[6][154] ), .A2(n5402), .A3(n5403), .A4(data[154]), .Y(n1751) );
  AO22X1_HVT U4824 ( .A1(\ram[6][153] ), .A2(n5402), .A3(n5403), .A4(data[153]), .Y(n1750) );
  AO22X1_HVT U4825 ( .A1(\ram[0][114] ), .A2(n5360), .A3(data[114]), .A4(n5361), .Y(n175) );
  AO22X1_HVT U4826 ( .A1(\ram[6][152] ), .A2(n5402), .A3(n5403), .A4(data[152]), .Y(n1749) );
  AO22X1_HVT U4827 ( .A1(\ram[6][151] ), .A2(n5402), .A3(n5403), .A4(data[151]), .Y(n1748) );
  AO22X1_HVT U4828 ( .A1(\ram[6][150] ), .A2(n5402), .A3(n5403), .A4(data[150]), .Y(n1747) );
  AO22X1_HVT U4829 ( .A1(\ram[6][149] ), .A2(n5402), .A3(n5403), .A4(data[149]), .Y(n1746) );
  AO22X1_HVT U4830 ( .A1(\ram[6][148] ), .A2(n5402), .A3(n5403), .A4(data[148]), .Y(n1745) );
  AO22X1_HVT U4831 ( .A1(\ram[6][147] ), .A2(n5402), .A3(n5403), .A4(data[147]), .Y(n1744) );
  AO22X1_HVT U4832 ( .A1(\ram[6][146] ), .A2(n5402), .A3(n5403), .A4(data[146]), .Y(n1743) );
  AO22X1_HVT U4833 ( .A1(\ram[6][145] ), .A2(n5402), .A3(n5403), .A4(data[145]), .Y(n1742) );
  AO22X1_HVT U4834 ( .A1(\ram[6][144] ), .A2(n5402), .A3(n5403), .A4(data[144]), .Y(n1741) );
  AO22X1_HVT U4835 ( .A1(\ram[6][143] ), .A2(n5402), .A3(n5403), .A4(data[143]), .Y(n1740) );
  AO22X1_HVT U4836 ( .A1(\ram[0][113] ), .A2(n5360), .A3(data[113]), .A4(n5361), .Y(n174) );
  AO22X1_HVT U4837 ( .A1(\ram[6][142] ), .A2(n5402), .A3(n5403), .A4(data[142]), .Y(n1739) );
  AO22X1_HVT U4838 ( .A1(\ram[6][141] ), .A2(n5402), .A3(n5403), .A4(data[141]), .Y(n1738) );
  AO22X1_HVT U4839 ( .A1(\ram[6][140] ), .A2(n5402), .A3(n5403), .A4(data[140]), .Y(n1737) );
  AO22X1_HVT U4840 ( .A1(\ram[6][139] ), .A2(n5402), .A3(n5403), .A4(data[139]), .Y(n1736) );
  AO22X1_HVT U4841 ( .A1(\ram[6][138] ), .A2(n5402), .A3(n5403), .A4(data[138]), .Y(n1735) );
  AO22X1_HVT U4842 ( .A1(\ram[6][137] ), .A2(n5402), .A3(n5403), .A4(data[137]), .Y(n1734) );
  AO22X1_HVT U4843 ( .A1(\ram[6][136] ), .A2(n5402), .A3(n5403), .A4(data[136]), .Y(n1733) );
  AO22X1_HVT U4844 ( .A1(\ram[6][135] ), .A2(n5402), .A3(n5403), .A4(data[135]), .Y(n1732) );
  AO22X1_HVT U4845 ( .A1(\ram[6][134] ), .A2(n5402), .A3(n5403), .A4(data[134]), .Y(n1731) );
  AO22X1_HVT U4846 ( .A1(\ram[6][133] ), .A2(n5402), .A3(n5403), .A4(data[133]), .Y(n1730) );
  AO22X1_HVT U4847 ( .A1(\ram[0][112] ), .A2(n5360), .A3(data[112]), .A4(n5361), .Y(n173) );
  AO22X1_HVT U4848 ( .A1(\ram[6][132] ), .A2(n5402), .A3(n5403), .A4(data[132]), .Y(n1729) );
  AO22X1_HVT U4849 ( .A1(\ram[6][131] ), .A2(n5402), .A3(n5403), .A4(data[131]), .Y(n1728) );
  AO22X1_HVT U4850 ( .A1(\ram[6][130] ), .A2(n5402), .A3(n5403), .A4(data[130]), .Y(n1727) );
  AO22X1_HVT U4851 ( .A1(\ram[6][129] ), .A2(n5402), .A3(n5403), .A4(data[129]), .Y(n1726) );
  AO22X1_HVT U4852 ( .A1(\ram[6][128] ), .A2(n5402), .A3(n5403), .A4(data[128]), .Y(n1725) );
  AO22X1_HVT U4853 ( .A1(\ram[6][127] ), .A2(n5402), .A3(n5403), .A4(data[127]), .Y(n1724) );
  AO22X1_HVT U4854 ( .A1(\ram[6][126] ), .A2(n5402), .A3(n5403), .A4(data[126]), .Y(n1723) );
  AO22X1_HVT U4855 ( .A1(\ram[6][125] ), .A2(n5402), .A3(n5403), .A4(data[125]), .Y(n1722) );
  AO22X1_HVT U4856 ( .A1(\ram[6][124] ), .A2(n5402), .A3(n5403), .A4(data[124]), .Y(n1721) );
  AO22X1_HVT U4857 ( .A1(\ram[6][123] ), .A2(n5402), .A3(n5403), .A4(data[123]), .Y(n1720) );
  AO22X1_HVT U4858 ( .A1(\ram[0][111] ), .A2(n5360), .A3(data[111]), .A4(n5361), .Y(n172) );
  AO22X1_HVT U4859 ( .A1(\ram[6][122] ), .A2(n5402), .A3(n5403), .A4(data[122]), .Y(n1719) );
  AO22X1_HVT U4860 ( .A1(\ram[6][121] ), .A2(n5402), .A3(n5403), .A4(data[121]), .Y(n1718) );
  AO22X1_HVT U4861 ( .A1(\ram[6][120] ), .A2(n5402), .A3(n5403), .A4(data[120]), .Y(n1717) );
  AO22X1_HVT U4862 ( .A1(\ram[6][119] ), .A2(n5402), .A3(n5403), .A4(data[119]), .Y(n1716) );
  AO22X1_HVT U4863 ( .A1(\ram[6][118] ), .A2(n5402), .A3(n5403), .A4(data[118]), .Y(n1715) );
  AO22X1_HVT U4864 ( .A1(\ram[6][117] ), .A2(n5402), .A3(n5403), .A4(data[117]), .Y(n1714) );
  AO22X1_HVT U4865 ( .A1(\ram[6][116] ), .A2(n5402), .A3(n5403), .A4(data[116]), .Y(n1713) );
  AO22X1_HVT U4866 ( .A1(\ram[6][115] ), .A2(n5402), .A3(n5403), .A4(data[115]), .Y(n1712) );
  AO22X1_HVT U4867 ( .A1(\ram[6][114] ), .A2(n5402), .A3(n5403), .A4(data[114]), .Y(n1711) );
  AO22X1_HVT U4868 ( .A1(\ram[6][113] ), .A2(n5402), .A3(n5403), .A4(data[113]), .Y(n1710) );
  AO22X1_HVT U4869 ( .A1(\ram[0][110] ), .A2(n5360), .A3(data[110]), .A4(n5361), .Y(n171) );
  AO22X1_HVT U4870 ( .A1(\ram[6][112] ), .A2(n5402), .A3(n5403), .A4(data[112]), .Y(n1709) );
  AO22X1_HVT U4871 ( .A1(\ram[6][111] ), .A2(n5402), .A3(n5403), .A4(data[111]), .Y(n1708) );
  AO22X1_HVT U4872 ( .A1(\ram[6][110] ), .A2(n5402), .A3(n5403), .A4(data[110]), .Y(n1707) );
  AO22X1_HVT U4873 ( .A1(\ram[6][109] ), .A2(n5402), .A3(n5403), .A4(data[109]), .Y(n1706) );
  AO22X1_HVT U4874 ( .A1(\ram[6][108] ), .A2(n5402), .A3(n5403), .A4(data[108]), .Y(n1705) );
  AO22X1_HVT U4875 ( .A1(\ram[6][107] ), .A2(n5402), .A3(n5403), .A4(data[107]), .Y(n1704) );
  AO22X1_HVT U4876 ( .A1(\ram[6][106] ), .A2(n5402), .A3(n5403), .A4(data[106]), .Y(n1703) );
  AO22X1_HVT U4877 ( .A1(\ram[6][105] ), .A2(n5402), .A3(n5403), .A4(data[105]), .Y(n1702) );
  AO22X1_HVT U4878 ( .A1(\ram[6][104] ), .A2(n5402), .A3(n5403), .A4(data[104]), .Y(n1701) );
  AO22X1_HVT U4879 ( .A1(\ram[6][103] ), .A2(n5402), .A3(n5403), .A4(data[103]), .Y(n1700) );
  AO22X1_HVT U4880 ( .A1(\ram[0][109] ), .A2(n5360), .A3(data[109]), .A4(n5361), .Y(n170) );
  AO22X1_HVT U4881 ( .A1(\ram[6][102] ), .A2(n5402), .A3(n5403), .A4(data[102]), .Y(n1699) );
  AO22X1_HVT U4882 ( .A1(\ram[6][101] ), .A2(n5402), .A3(n5403), .A4(data[101]), .Y(n1698) );
  AO22X1_HVT U4883 ( .A1(\ram[6][100] ), .A2(n5402), .A3(n5403), .A4(data[100]), .Y(n1697) );
  AO22X1_HVT U4884 ( .A1(\ram[6][99] ), .A2(n5402), .A3(n5403), .A4(data[99]), 
        .Y(n1696) );
  AO22X1_HVT U4885 ( .A1(\ram[6][98] ), .A2(n5402), .A3(n5403), .A4(data[98]), 
        .Y(n1695) );
  AO22X1_HVT U4886 ( .A1(\ram[6][97] ), .A2(n5402), .A3(n5403), .A4(data[97]), 
        .Y(n1694) );
  AO22X1_HVT U4887 ( .A1(\ram[6][96] ), .A2(n5402), .A3(n5403), .A4(data[96]), 
        .Y(n1693) );
  AO22X1_HVT U4888 ( .A1(\ram[6][95] ), .A2(n5402), .A3(n5403), .A4(data[95]), 
        .Y(n1692) );
  AO22X1_HVT U4889 ( .A1(\ram[6][94] ), .A2(n5402), .A3(n5403), .A4(data[94]), 
        .Y(n1691) );
  AO22X1_HVT U4890 ( .A1(\ram[6][93] ), .A2(n5402), .A3(n5403), .A4(data[93]), 
        .Y(n1690) );
  AO22X1_HVT U4891 ( .A1(\ram[0][108] ), .A2(n5360), .A3(data[108]), .A4(n5361), .Y(n169) );
  AO22X1_HVT U4892 ( .A1(\ram[6][92] ), .A2(n5402), .A3(n5403), .A4(data[92]), 
        .Y(n1689) );
  AO22X1_HVT U4893 ( .A1(\ram[6][91] ), .A2(n5402), .A3(n5403), .A4(data[91]), 
        .Y(n1688) );
  AO22X1_HVT U4894 ( .A1(\ram[6][90] ), .A2(n5402), .A3(n5403), .A4(data[90]), 
        .Y(n1687) );
  AO22X1_HVT U4895 ( .A1(\ram[6][89] ), .A2(n5402), .A3(n5403), .A4(data[89]), 
        .Y(n1686) );
  AO22X1_HVT U4896 ( .A1(\ram[6][88] ), .A2(n5402), .A3(n5403), .A4(data[88]), 
        .Y(n1685) );
  AO22X1_HVT U4897 ( .A1(\ram[6][87] ), .A2(n5402), .A3(n5403), .A4(data[87]), 
        .Y(n1684) );
  AO22X1_HVT U4898 ( .A1(\ram[6][86] ), .A2(n5402), .A3(n5403), .A4(data[86]), 
        .Y(n1683) );
  AO22X1_HVT U4899 ( .A1(\ram[6][85] ), .A2(n5402), .A3(n5403), .A4(data[85]), 
        .Y(n1682) );
  AO22X1_HVT U4900 ( .A1(\ram[6][84] ), .A2(n5402), .A3(n5403), .A4(data[84]), 
        .Y(n1681) );
  AO22X1_HVT U4901 ( .A1(\ram[6][83] ), .A2(n5402), .A3(n5403), .A4(data[83]), 
        .Y(n1680) );
  AO22X1_HVT U4902 ( .A1(\ram[0][107] ), .A2(n5360), .A3(data[107]), .A4(n5361), .Y(n168) );
  AO22X1_HVT U4903 ( .A1(\ram[6][82] ), .A2(n5402), .A3(n5403), .A4(data[82]), 
        .Y(n1679) );
  AO22X1_HVT U4904 ( .A1(\ram[6][81] ), .A2(n5402), .A3(n5403), .A4(data[81]), 
        .Y(n1678) );
  AO22X1_HVT U4905 ( .A1(\ram[6][80] ), .A2(n5402), .A3(n5403), .A4(data[80]), 
        .Y(n1677) );
  AO22X1_HVT U4906 ( .A1(\ram[6][79] ), .A2(n5402), .A3(n5403), .A4(data[79]), 
        .Y(n1676) );
  AO22X1_HVT U4907 ( .A1(\ram[6][78] ), .A2(n5402), .A3(n5403), .A4(data[78]), 
        .Y(n1675) );
  AO22X1_HVT U4908 ( .A1(\ram[6][77] ), .A2(n5402), .A3(n5403), .A4(data[77]), 
        .Y(n1674) );
  AO22X1_HVT U4909 ( .A1(\ram[6][76] ), .A2(n5402), .A3(n5403), .A4(data[76]), 
        .Y(n1673) );
  AO22X1_HVT U4910 ( .A1(\ram[6][75] ), .A2(n5402), .A3(n5403), .A4(data[75]), 
        .Y(n1672) );
  AO22X1_HVT U4911 ( .A1(\ram[6][74] ), .A2(n5402), .A3(n5403), .A4(data[74]), 
        .Y(n1671) );
  AO22X1_HVT U4912 ( .A1(\ram[6][73] ), .A2(n5402), .A3(n5403), .A4(data[73]), 
        .Y(n1670) );
  AO22X1_HVT U4913 ( .A1(\ram[0][106] ), .A2(n5360), .A3(data[106]), .A4(n5361), .Y(n167) );
  AO22X1_HVT U4914 ( .A1(\ram[6][72] ), .A2(n5402), .A3(n5403), .A4(data[72]), 
        .Y(n1669) );
  AO22X1_HVT U4915 ( .A1(\ram[6][71] ), .A2(n5402), .A3(n5403), .A4(data[71]), 
        .Y(n1668) );
  AO22X1_HVT U4916 ( .A1(\ram[6][70] ), .A2(n5402), .A3(n5403), .A4(data[70]), 
        .Y(n1667) );
  AO22X1_HVT U4917 ( .A1(\ram[6][69] ), .A2(n5402), .A3(n5403), .A4(data[69]), 
        .Y(n1666) );
  AO22X1_HVT U4918 ( .A1(\ram[6][68] ), .A2(n5402), .A3(n5403), .A4(data[68]), 
        .Y(n1665) );
  AO22X1_HVT U4919 ( .A1(\ram[6][67] ), .A2(n5402), .A3(n5403), .A4(data[67]), 
        .Y(n1664) );
  AO22X1_HVT U4920 ( .A1(\ram[6][66] ), .A2(n5402), .A3(n5403), .A4(data[66]), 
        .Y(n1663) );
  AO22X1_HVT U4921 ( .A1(\ram[6][65] ), .A2(n5402), .A3(n5403), .A4(data[65]), 
        .Y(n1662) );
  AO22X1_HVT U4922 ( .A1(\ram[6][64] ), .A2(n5402), .A3(n5403), .A4(data[64]), 
        .Y(n1661) );
  AO22X1_HVT U4923 ( .A1(\ram[6][63] ), .A2(n5402), .A3(n5403), .A4(data[63]), 
        .Y(n1660) );
  AO22X1_HVT U4924 ( .A1(\ram[0][105] ), .A2(n5360), .A3(data[105]), .A4(n5361), .Y(n166) );
  AO22X1_HVT U4925 ( .A1(\ram[6][62] ), .A2(n5402), .A3(n5403), .A4(data[62]), 
        .Y(n1659) );
  AO22X1_HVT U4926 ( .A1(\ram[6][61] ), .A2(n5402), .A3(n5403), .A4(data[61]), 
        .Y(n1658) );
  AO22X1_HVT U4927 ( .A1(\ram[6][60] ), .A2(n5402), .A3(n5403), .A4(data[60]), 
        .Y(n1657) );
  AO22X1_HVT U4928 ( .A1(\ram[6][59] ), .A2(n5402), .A3(n5403), .A4(data[59]), 
        .Y(n1656) );
  AO22X1_HVT U4929 ( .A1(\ram[6][58] ), .A2(n5402), .A3(n5403), .A4(data[58]), 
        .Y(n1655) );
  AO22X1_HVT U4930 ( .A1(\ram[6][57] ), .A2(n5402), .A3(n5403), .A4(data[57]), 
        .Y(n1654) );
  AO22X1_HVT U4931 ( .A1(\ram[6][56] ), .A2(n5402), .A3(n5403), .A4(data[56]), 
        .Y(n1653) );
  AO22X1_HVT U4932 ( .A1(\ram[6][55] ), .A2(n5402), .A3(n5403), .A4(data[55]), 
        .Y(n1652) );
  AO22X1_HVT U4933 ( .A1(\ram[6][54] ), .A2(n5402), .A3(n5403), .A4(data[54]), 
        .Y(n1651) );
  AO22X1_HVT U4934 ( .A1(\ram[6][53] ), .A2(n5402), .A3(n5403), .A4(data[53]), 
        .Y(n1650) );
  AO22X1_HVT U4935 ( .A1(\ram[0][104] ), .A2(n5360), .A3(data[104]), .A4(n5361), .Y(n165) );
  AO22X1_HVT U4936 ( .A1(\ram[6][52] ), .A2(n5402), .A3(n5403), .A4(data[52]), 
        .Y(n1649) );
  AO22X1_HVT U4937 ( .A1(\ram[6][51] ), .A2(n5402), .A3(n5403), .A4(data[51]), 
        .Y(n1648) );
  AO22X1_HVT U4938 ( .A1(\ram[6][50] ), .A2(n5402), .A3(n5403), .A4(data[50]), 
        .Y(n1647) );
  AO22X1_HVT U4939 ( .A1(\ram[6][49] ), .A2(n5402), .A3(n5403), .A4(data[49]), 
        .Y(n1646) );
  AO22X1_HVT U4940 ( .A1(\ram[6][48] ), .A2(n5402), .A3(n5403), .A4(data[48]), 
        .Y(n1645) );
  AO22X1_HVT U4941 ( .A1(\ram[6][47] ), .A2(n5402), .A3(n5403), .A4(data[47]), 
        .Y(n1644) );
  AO22X1_HVT U4942 ( .A1(\ram[6][46] ), .A2(n5402), .A3(n5403), .A4(data[46]), 
        .Y(n1643) );
  AO22X1_HVT U4943 ( .A1(\ram[6][45] ), .A2(n5402), .A3(n5403), .A4(data[45]), 
        .Y(n1642) );
  AO22X1_HVT U4944 ( .A1(\ram[6][44] ), .A2(n5402), .A3(n5403), .A4(data[44]), 
        .Y(n1641) );
  AO22X1_HVT U4945 ( .A1(\ram[6][43] ), .A2(n5402), .A3(n5403), .A4(data[43]), 
        .Y(n1640) );
  AO22X1_HVT U4946 ( .A1(\ram[0][103] ), .A2(n5360), .A3(data[103]), .A4(n5361), .Y(n164) );
  AO22X1_HVT U4947 ( .A1(\ram[6][42] ), .A2(n5402), .A3(n5403), .A4(data[42]), 
        .Y(n1639) );
  AO22X1_HVT U4948 ( .A1(\ram[6][41] ), .A2(n5402), .A3(n5403), .A4(data[41]), 
        .Y(n1638) );
  AO22X1_HVT U4949 ( .A1(\ram[6][40] ), .A2(n5402), .A3(n5403), .A4(data[40]), 
        .Y(n1637) );
  AO22X1_HVT U4950 ( .A1(\ram[6][39] ), .A2(n5402), .A3(n5403), .A4(data[39]), 
        .Y(n1636) );
  AO22X1_HVT U4951 ( .A1(\ram[6][38] ), .A2(n5402), .A3(n5403), .A4(data[38]), 
        .Y(n1635) );
  AO22X1_HVT U4952 ( .A1(\ram[6][37] ), .A2(n5402), .A3(n5403), .A4(data[37]), 
        .Y(n1634) );
  AO22X1_HVT U4953 ( .A1(\ram[6][36] ), .A2(n5402), .A3(n5403), .A4(data[36]), 
        .Y(n1633) );
  AO22X1_HVT U4954 ( .A1(\ram[6][35] ), .A2(n5402), .A3(n5403), .A4(data[35]), 
        .Y(n1632) );
  AO22X1_HVT U4955 ( .A1(\ram[6][34] ), .A2(n5402), .A3(n5403), .A4(data[34]), 
        .Y(n1631) );
  AO22X1_HVT U4956 ( .A1(\ram[6][33] ), .A2(n5402), .A3(n5403), .A4(data[33]), 
        .Y(n1630) );
  AO22X1_HVT U4957 ( .A1(\ram[0][102] ), .A2(n5360), .A3(data[102]), .A4(n5361), .Y(n163) );
  AO22X1_HVT U4958 ( .A1(\ram[6][32] ), .A2(n5402), .A3(n5403), .A4(data[32]), 
        .Y(n1629) );
  AO22X1_HVT U4959 ( .A1(\ram[6][31] ), .A2(n5402), .A3(n5403), .A4(data[31]), 
        .Y(n1628) );
  AO22X1_HVT U4960 ( .A1(\ram[6][30] ), .A2(n5402), .A3(n5403), .A4(data[30]), 
        .Y(n1627) );
  AO22X1_HVT U4961 ( .A1(\ram[6][29] ), .A2(n5402), .A3(n5403), .A4(data[29]), 
        .Y(n1626) );
  AO22X1_HVT U4962 ( .A1(\ram[6][28] ), .A2(n5402), .A3(n5403), .A4(data[28]), 
        .Y(n1625) );
  AO22X1_HVT U4963 ( .A1(\ram[6][27] ), .A2(n5402), .A3(n5403), .A4(data[27]), 
        .Y(n1624) );
  AO22X1_HVT U4964 ( .A1(\ram[6][26] ), .A2(n5402), .A3(n5403), .A4(data[26]), 
        .Y(n1623) );
  AO22X1_HVT U4965 ( .A1(\ram[6][25] ), .A2(n5402), .A3(n5403), .A4(data[25]), 
        .Y(n1622) );
  AO22X1_HVT U4966 ( .A1(\ram[6][24] ), .A2(n5402), .A3(n5403), .A4(data[24]), 
        .Y(n1621) );
  AO22X1_HVT U4967 ( .A1(\ram[6][23] ), .A2(n5402), .A3(n5403), .A4(data[23]), 
        .Y(n1620) );
  AO22X1_HVT U4968 ( .A1(\ram[0][101] ), .A2(n5360), .A3(data[101]), .A4(n5361), .Y(n162) );
  AO22X1_HVT U4969 ( .A1(\ram[6][22] ), .A2(n5402), .A3(n5403), .A4(data[22]), 
        .Y(n1619) );
  AO22X1_HVT U4970 ( .A1(\ram[6][21] ), .A2(n5402), .A3(n5403), .A4(data[21]), 
        .Y(n1618) );
  AO22X1_HVT U4971 ( .A1(\ram[6][20] ), .A2(n5402), .A3(n5403), .A4(data[20]), 
        .Y(n1617) );
  AO22X1_HVT U4972 ( .A1(\ram[6][19] ), .A2(n5402), .A3(n5403), .A4(data[19]), 
        .Y(n1616) );
  AO22X1_HVT U4973 ( .A1(\ram[6][18] ), .A2(n5402), .A3(n5403), .A4(data[18]), 
        .Y(n1615) );
  AO22X1_HVT U4974 ( .A1(\ram[6][17] ), .A2(n5402), .A3(n5403), .A4(data[17]), 
        .Y(n1614) );
  AO22X1_HVT U4975 ( .A1(\ram[6][16] ), .A2(n5402), .A3(n5403), .A4(data[16]), 
        .Y(n1613) );
  AO22X1_HVT U4976 ( .A1(\ram[6][15] ), .A2(n5402), .A3(n5403), .A4(data[15]), 
        .Y(n1612) );
  AO22X1_HVT U4977 ( .A1(\ram[6][14] ), .A2(n5402), .A3(n5403), .A4(data[14]), 
        .Y(n1611) );
  AO22X1_HVT U4978 ( .A1(\ram[6][13] ), .A2(n5402), .A3(n5403), .A4(data[13]), 
        .Y(n1610) );
  AO22X1_HVT U4979 ( .A1(\ram[0][100] ), .A2(n5360), .A3(data[100]), .A4(n5361), .Y(n161) );
  AO22X1_HVT U4980 ( .A1(\ram[6][12] ), .A2(n5402), .A3(n5403), .A4(data[12]), 
        .Y(n1609) );
  AO22X1_HVT U4981 ( .A1(\ram[6][11] ), .A2(n5402), .A3(n5403), .A4(data[11]), 
        .Y(n1608) );
  AO22X1_HVT U4982 ( .A1(\ram[6][10] ), .A2(n5402), .A3(n5403), .A4(data[10]), 
        .Y(n1607) );
  AO22X1_HVT U4983 ( .A1(\ram[6][9] ), .A2(n5402), .A3(n5403), .A4(data[9]), 
        .Y(n1606) );
  AO22X1_HVT U4984 ( .A1(\ram[6][8] ), .A2(n5402), .A3(n5403), .A4(data[8]), 
        .Y(n1605) );
  AO22X1_HVT U4985 ( .A1(\ram[6][7] ), .A2(n5402), .A3(n5403), .A4(data[7]), 
        .Y(n1604) );
  AO22X1_HVT U4986 ( .A1(\ram[6][6] ), .A2(n5402), .A3(n5403), .A4(data[6]), 
        .Y(n1603) );
  AO22X1_HVT U4987 ( .A1(\ram[6][5] ), .A2(n5402), .A3(n5403), .A4(data[5]), 
        .Y(n1602) );
  AO22X1_HVT U4988 ( .A1(\ram[6][4] ), .A2(n5402), .A3(n5403), .A4(data[4]), 
        .Y(n1601) );
  AO22X1_HVT U4989 ( .A1(\ram[6][3] ), .A2(n5402), .A3(n5403), .A4(data[3]), 
        .Y(n1600) );
  AO22X1_HVT U4990 ( .A1(\ram[0][99] ), .A2(n5360), .A3(data[99]), .A4(n5361), 
        .Y(n160) );
  AO22X1_HVT U4991 ( .A1(\ram[6][2] ), .A2(n5402), .A3(n5403), .A4(data[2]), 
        .Y(n1599) );
  AO22X1_HVT U4992 ( .A1(\ram[6][1] ), .A2(n5402), .A3(n5403), .A4(data[1]), 
        .Y(n1598) );
  AO22X1_HVT U4993 ( .A1(\ram[6][0] ), .A2(n5402), .A3(n5403), .A4(data[0]), 
        .Y(n1597) );
  INVX0_HVT U4994 ( .A(n5404), .Y(n5403) );
  AND2X1_HVT U4995 ( .A1(n5404), .A2(n5365), .Y(n5402) );
  NAND3X0_HVT U4996 ( .A1(n4276), .A2(n4183), .A3(n5401), .Y(n5404) );
  AO22X1_HVT U4997 ( .A1(\ram[5][255] ), .A2(n5405), .A3(n5406), .A4(data[255]), .Y(n1596) );
  AO22X1_HVT U4998 ( .A1(\ram[5][254] ), .A2(n5405), .A3(n5406), .A4(data[254]), .Y(n1595) );
  AO22X1_HVT U4999 ( .A1(\ram[5][253] ), .A2(n5405), .A3(n5406), .A4(data[253]), .Y(n1594) );
  AO22X1_HVT U5000 ( .A1(\ram[5][252] ), .A2(n5405), .A3(n5406), .A4(data[252]), .Y(n1593) );
  AO22X1_HVT U5001 ( .A1(\ram[5][251] ), .A2(n5405), .A3(n5406), .A4(data[251]), .Y(n1592) );
  AO22X1_HVT U5002 ( .A1(\ram[5][250] ), .A2(n5405), .A3(n5406), .A4(data[250]), .Y(n1591) );
  AO22X1_HVT U5003 ( .A1(\ram[5][249] ), .A2(n5405), .A3(n5406), .A4(data[249]), .Y(n1590) );
  AO22X1_HVT U5004 ( .A1(\ram[0][98] ), .A2(n5360), .A3(data[98]), .A4(n5361), 
        .Y(n159) );
  AO22X1_HVT U5005 ( .A1(\ram[5][248] ), .A2(n5405), .A3(n5406), .A4(data[248]), .Y(n1589) );
  AO22X1_HVT U5006 ( .A1(\ram[5][247] ), .A2(n5405), .A3(n5406), .A4(data[247]), .Y(n1588) );
  AO22X1_HVT U5007 ( .A1(\ram[5][246] ), .A2(n5405), .A3(n5406), .A4(data[246]), .Y(n1587) );
  AO22X1_HVT U5008 ( .A1(\ram[5][245] ), .A2(n5405), .A3(n5406), .A4(data[245]), .Y(n1586) );
  AO22X1_HVT U5009 ( .A1(\ram[5][244] ), .A2(n5405), .A3(n5406), .A4(data[244]), .Y(n1585) );
  AO22X1_HVT U5010 ( .A1(\ram[5][243] ), .A2(n5405), .A3(n5406), .A4(data[243]), .Y(n1584) );
  AO22X1_HVT U5011 ( .A1(\ram[5][242] ), .A2(n5405), .A3(n5406), .A4(data[242]), .Y(n1583) );
  AO22X1_HVT U5012 ( .A1(\ram[5][241] ), .A2(n5405), .A3(n5406), .A4(data[241]), .Y(n1582) );
  AO22X1_HVT U5013 ( .A1(\ram[5][240] ), .A2(n5405), .A3(n5406), .A4(data[240]), .Y(n1581) );
  AO22X1_HVT U5014 ( .A1(\ram[5][239] ), .A2(n5405), .A3(n5406), .A4(data[239]), .Y(n1580) );
  AO22X1_HVT U5015 ( .A1(\ram[0][97] ), .A2(n5360), .A3(data[97]), .A4(n5361), 
        .Y(n158) );
  AO22X1_HVT U5016 ( .A1(\ram[5][238] ), .A2(n5405), .A3(n5406), .A4(data[238]), .Y(n1579) );
  AO22X1_HVT U5017 ( .A1(\ram[5][237] ), .A2(n5405), .A3(n5406), .A4(data[237]), .Y(n1578) );
  AO22X1_HVT U5018 ( .A1(\ram[5][236] ), .A2(n5405), .A3(n5406), .A4(data[236]), .Y(n1577) );
  AO22X1_HVT U5019 ( .A1(\ram[5][235] ), .A2(n5405), .A3(n5406), .A4(data[235]), .Y(n1576) );
  AO22X1_HVT U5020 ( .A1(\ram[5][234] ), .A2(n5405), .A3(n5406), .A4(data[234]), .Y(n1575) );
  AO22X1_HVT U5021 ( .A1(\ram[5][233] ), .A2(n5405), .A3(n5406), .A4(data[233]), .Y(n1574) );
  AO22X1_HVT U5022 ( .A1(\ram[5][232] ), .A2(n5405), .A3(n5406), .A4(data[232]), .Y(n1573) );
  AO22X1_HVT U5023 ( .A1(\ram[5][231] ), .A2(n5405), .A3(n5406), .A4(data[231]), .Y(n1572) );
  AO22X1_HVT U5024 ( .A1(\ram[5][230] ), .A2(n5405), .A3(n5406), .A4(data[230]), .Y(n1571) );
  AO22X1_HVT U5025 ( .A1(\ram[5][229] ), .A2(n5405), .A3(n5406), .A4(data[229]), .Y(n1570) );
  AO22X1_HVT U5026 ( .A1(\ram[0][96] ), .A2(n5360), .A3(data[96]), .A4(n5361), 
        .Y(n157) );
  AO22X1_HVT U5027 ( .A1(\ram[5][228] ), .A2(n5405), .A3(n5406), .A4(data[228]), .Y(n1569) );
  AO22X1_HVT U5028 ( .A1(\ram[5][227] ), .A2(n5405), .A3(n5406), .A4(data[227]), .Y(n1568) );
  AO22X1_HVT U5029 ( .A1(\ram[5][226] ), .A2(n5405), .A3(n5406), .A4(data[226]), .Y(n1567) );
  AO22X1_HVT U5030 ( .A1(\ram[5][225] ), .A2(n5405), .A3(n5406), .A4(data[225]), .Y(n1566) );
  AO22X1_HVT U5031 ( .A1(\ram[5][224] ), .A2(n5405), .A3(n5406), .A4(data[224]), .Y(n1565) );
  AO22X1_HVT U5032 ( .A1(\ram[5][223] ), .A2(n5405), .A3(n5406), .A4(data[223]), .Y(n1564) );
  AO22X1_HVT U5033 ( .A1(\ram[5][222] ), .A2(n5405), .A3(n5406), .A4(data[222]), .Y(n1563) );
  AO22X1_HVT U5034 ( .A1(\ram[5][221] ), .A2(n5405), .A3(n5406), .A4(data[221]), .Y(n1562) );
  AO22X1_HVT U5035 ( .A1(\ram[5][220] ), .A2(n5405), .A3(n5406), .A4(data[220]), .Y(n1561) );
  AO22X1_HVT U5036 ( .A1(\ram[5][219] ), .A2(n5405), .A3(n5406), .A4(data[219]), .Y(n1560) );
  AO22X1_HVT U5037 ( .A1(\ram[0][95] ), .A2(n5360), .A3(data[95]), .A4(n5361), 
        .Y(n156) );
  AO22X1_HVT U5038 ( .A1(\ram[5][218] ), .A2(n5405), .A3(n5406), .A4(data[218]), .Y(n1559) );
  AO22X1_HVT U5039 ( .A1(\ram[5][217] ), .A2(n5405), .A3(n5406), .A4(data[217]), .Y(n1558) );
  AO22X1_HVT U5040 ( .A1(\ram[5][216] ), .A2(n5405), .A3(n5406), .A4(data[216]), .Y(n1557) );
  AO22X1_HVT U5041 ( .A1(\ram[5][215] ), .A2(n5405), .A3(n5406), .A4(data[215]), .Y(n1556) );
  AO22X1_HVT U5042 ( .A1(\ram[5][214] ), .A2(n5405), .A3(n5406), .A4(data[214]), .Y(n1555) );
  AO22X1_HVT U5043 ( .A1(\ram[5][213] ), .A2(n5405), .A3(n5406), .A4(data[213]), .Y(n1554) );
  AO22X1_HVT U5044 ( .A1(\ram[5][212] ), .A2(n5405), .A3(n5406), .A4(data[212]), .Y(n1553) );
  AO22X1_HVT U5045 ( .A1(\ram[5][211] ), .A2(n5405), .A3(n5406), .A4(data[211]), .Y(n1552) );
  AO22X1_HVT U5046 ( .A1(\ram[5][210] ), .A2(n5405), .A3(n5406), .A4(data[210]), .Y(n1551) );
  AO22X1_HVT U5047 ( .A1(\ram[5][209] ), .A2(n5405), .A3(n5406), .A4(data[209]), .Y(n1550) );
  AO22X1_HVT U5048 ( .A1(\ram[0][94] ), .A2(n5360), .A3(data[94]), .A4(n5361), 
        .Y(n155) );
  AO22X1_HVT U5049 ( .A1(\ram[5][208] ), .A2(n5405), .A3(n5406), .A4(data[208]), .Y(n1549) );
  AO22X1_HVT U5050 ( .A1(\ram[5][207] ), .A2(n5405), .A3(n5406), .A4(data[207]), .Y(n1548) );
  AO22X1_HVT U5051 ( .A1(\ram[5][206] ), .A2(n5405), .A3(n5406), .A4(data[206]), .Y(n1547) );
  AO22X1_HVT U5052 ( .A1(\ram[5][205] ), .A2(n5405), .A3(n5406), .A4(data[205]), .Y(n1546) );
  AO22X1_HVT U5053 ( .A1(\ram[5][204] ), .A2(n5405), .A3(n5406), .A4(data[204]), .Y(n1545) );
  AO22X1_HVT U5054 ( .A1(\ram[5][203] ), .A2(n5405), .A3(n5406), .A4(data[203]), .Y(n1544) );
  AO22X1_HVT U5055 ( .A1(\ram[5][202] ), .A2(n5405), .A3(n5406), .A4(data[202]), .Y(n1543) );
  AO22X1_HVT U5056 ( .A1(\ram[5][201] ), .A2(n5405), .A3(n5406), .A4(data[201]), .Y(n1542) );
  AO22X1_HVT U5057 ( .A1(\ram[5][200] ), .A2(n5405), .A3(n5406), .A4(data[200]), .Y(n1541) );
  AO22X1_HVT U5058 ( .A1(\ram[5][199] ), .A2(n5405), .A3(n5406), .A4(data[199]), .Y(n1540) );
  AO22X1_HVT U5059 ( .A1(\ram[0][93] ), .A2(n5360), .A3(data[93]), .A4(n5361), 
        .Y(n154) );
  AO22X1_HVT U5060 ( .A1(\ram[5][198] ), .A2(n5405), .A3(n5406), .A4(data[198]), .Y(n1539) );
  AO22X1_HVT U5061 ( .A1(\ram[5][197] ), .A2(n5405), .A3(n5406), .A4(data[197]), .Y(n1538) );
  AO22X1_HVT U5062 ( .A1(\ram[5][196] ), .A2(n5405), .A3(n5406), .A4(data[196]), .Y(n1537) );
  AO22X1_HVT U5063 ( .A1(\ram[5][195] ), .A2(n5405), .A3(n5406), .A4(data[195]), .Y(n1536) );
  AO22X1_HVT U5064 ( .A1(\ram[5][194] ), .A2(n5405), .A3(n5406), .A4(data[194]), .Y(n1535) );
  AO22X1_HVT U5065 ( .A1(\ram[5][193] ), .A2(n5405), .A3(n5406), .A4(data[193]), .Y(n1534) );
  AO22X1_HVT U5066 ( .A1(\ram[5][192] ), .A2(n5405), .A3(n5406), .A4(data[192]), .Y(n1533) );
  AO22X1_HVT U5067 ( .A1(\ram[5][191] ), .A2(n5405), .A3(n5406), .A4(data[191]), .Y(n1532) );
  AO22X1_HVT U5068 ( .A1(\ram[5][190] ), .A2(n5405), .A3(n5406), .A4(data[190]), .Y(n1531) );
  AO22X1_HVT U5069 ( .A1(\ram[5][189] ), .A2(n5405), .A3(n5406), .A4(data[189]), .Y(n1530) );
  AO22X1_HVT U5070 ( .A1(\ram[0][92] ), .A2(n5360), .A3(data[92]), .A4(n5361), 
        .Y(n153) );
  AO22X1_HVT U5071 ( .A1(\ram[5][188] ), .A2(n5405), .A3(n5406), .A4(data[188]), .Y(n1529) );
  AO22X1_HVT U5072 ( .A1(\ram[5][187] ), .A2(n5405), .A3(n5406), .A4(data[187]), .Y(n1528) );
  AO22X1_HVT U5073 ( .A1(\ram[5][186] ), .A2(n5405), .A3(n5406), .A4(data[186]), .Y(n1527) );
  AO22X1_HVT U5074 ( .A1(\ram[5][185] ), .A2(n5405), .A3(n5406), .A4(data[185]), .Y(n1526) );
  AO22X1_HVT U5075 ( .A1(\ram[5][184] ), .A2(n5405), .A3(n5406), .A4(data[184]), .Y(n1525) );
  AO22X1_HVT U5076 ( .A1(\ram[5][183] ), .A2(n5405), .A3(n5406), .A4(data[183]), .Y(n1524) );
  AO22X1_HVT U5077 ( .A1(\ram[5][182] ), .A2(n5405), .A3(n5406), .A4(data[182]), .Y(n1523) );
  AO22X1_HVT U5078 ( .A1(\ram[5][181] ), .A2(n5405), .A3(n5406), .A4(data[181]), .Y(n1522) );
  AO22X1_HVT U5079 ( .A1(\ram[5][180] ), .A2(n5405), .A3(n5406), .A4(data[180]), .Y(n1521) );
  AO22X1_HVT U5080 ( .A1(\ram[5][179] ), .A2(n5405), .A3(n5406), .A4(data[179]), .Y(n1520) );
  AO22X1_HVT U5081 ( .A1(\ram[0][91] ), .A2(n5360), .A3(data[91]), .A4(n5361), 
        .Y(n152) );
  AO22X1_HVT U5082 ( .A1(\ram[5][178] ), .A2(n5405), .A3(n5406), .A4(data[178]), .Y(n1519) );
  AO22X1_HVT U5083 ( .A1(\ram[5][177] ), .A2(n5405), .A3(n5406), .A4(data[177]), .Y(n1518) );
  AO22X1_HVT U5084 ( .A1(\ram[5][176] ), .A2(n5405), .A3(n5406), .A4(data[176]), .Y(n1517) );
  AO22X1_HVT U5085 ( .A1(\ram[5][175] ), .A2(n5405), .A3(n5406), .A4(data[175]), .Y(n1516) );
  AO22X1_HVT U5086 ( .A1(\ram[5][174] ), .A2(n5405), .A3(n5406), .A4(data[174]), .Y(n1515) );
  AO22X1_HVT U5087 ( .A1(\ram[5][173] ), .A2(n5405), .A3(n5406), .A4(data[173]), .Y(n1514) );
  AO22X1_HVT U5088 ( .A1(\ram[5][172] ), .A2(n5405), .A3(n5406), .A4(data[172]), .Y(n1513) );
  AO22X1_HVT U5089 ( .A1(\ram[5][171] ), .A2(n5405), .A3(n5406), .A4(data[171]), .Y(n1512) );
  AO22X1_HVT U5090 ( .A1(\ram[5][170] ), .A2(n5405), .A3(n5406), .A4(data[170]), .Y(n1511) );
  AO22X1_HVT U5091 ( .A1(\ram[5][169] ), .A2(n5405), .A3(n5406), .A4(data[169]), .Y(n1510) );
  AO22X1_HVT U5092 ( .A1(\ram[0][90] ), .A2(n5360), .A3(data[90]), .A4(n5361), 
        .Y(n151) );
  AO22X1_HVT U5093 ( .A1(\ram[5][168] ), .A2(n5405), .A3(n5406), .A4(data[168]), .Y(n1509) );
  AO22X1_HVT U5094 ( .A1(\ram[5][167] ), .A2(n5405), .A3(n5406), .A4(data[167]), .Y(n1508) );
  AO22X1_HVT U5095 ( .A1(\ram[5][166] ), .A2(n5405), .A3(n5406), .A4(data[166]), .Y(n1507) );
  AO22X1_HVT U5096 ( .A1(\ram[5][165] ), .A2(n5405), .A3(n5406), .A4(data[165]), .Y(n1506) );
  AO22X1_HVT U5097 ( .A1(\ram[5][164] ), .A2(n5405), .A3(n5406), .A4(data[164]), .Y(n1505) );
  AO22X1_HVT U5098 ( .A1(\ram[5][163] ), .A2(n5405), .A3(n5406), .A4(data[163]), .Y(n1504) );
  AO22X1_HVT U5099 ( .A1(\ram[5][162] ), .A2(n5405), .A3(n5406), .A4(data[162]), .Y(n1503) );
  AO22X1_HVT U5100 ( .A1(\ram[5][161] ), .A2(n5405), .A3(n5406), .A4(data[161]), .Y(n1502) );
  AO22X1_HVT U5101 ( .A1(\ram[5][160] ), .A2(n5405), .A3(n5406), .A4(data[160]), .Y(n1501) );
  AO22X1_HVT U5102 ( .A1(\ram[5][159] ), .A2(n5405), .A3(n5406), .A4(data[159]), .Y(n1500) );
  AO22X1_HVT U5103 ( .A1(\ram[0][89] ), .A2(n5360), .A3(data[89]), .A4(n5361), 
        .Y(n150) );
  AO22X1_HVT U5104 ( .A1(\ram[5][158] ), .A2(n5405), .A3(n5406), .A4(data[158]), .Y(n1499) );
  AO22X1_HVT U5105 ( .A1(\ram[5][157] ), .A2(n5405), .A3(n5406), .A4(data[157]), .Y(n1498) );
  AO22X1_HVT U5106 ( .A1(\ram[5][156] ), .A2(n5405), .A3(n5406), .A4(data[156]), .Y(n1497) );
  AO22X1_HVT U5107 ( .A1(\ram[5][155] ), .A2(n5405), .A3(n5406), .A4(data[155]), .Y(n1496) );
  AO22X1_HVT U5108 ( .A1(\ram[5][154] ), .A2(n5405), .A3(n5406), .A4(data[154]), .Y(n1495) );
  AO22X1_HVT U5109 ( .A1(\ram[5][153] ), .A2(n5405), .A3(n5406), .A4(data[153]), .Y(n1494) );
  AO22X1_HVT U5110 ( .A1(\ram[5][152] ), .A2(n5405), .A3(n5406), .A4(data[152]), .Y(n1493) );
  AO22X1_HVT U5111 ( .A1(\ram[5][151] ), .A2(n5405), .A3(n5406), .A4(data[151]), .Y(n1492) );
  AO22X1_HVT U5112 ( .A1(\ram[5][150] ), .A2(n5405), .A3(n5406), .A4(data[150]), .Y(n1491) );
  AO22X1_HVT U5113 ( .A1(\ram[5][149] ), .A2(n5405), .A3(n5406), .A4(data[149]), .Y(n1490) );
  AO22X1_HVT U5114 ( .A1(\ram[0][88] ), .A2(n5360), .A3(data[88]), .A4(n5361), 
        .Y(n149) );
  AO22X1_HVT U5115 ( .A1(\ram[5][148] ), .A2(n5405), .A3(n5406), .A4(data[148]), .Y(n1489) );
  AO22X1_HVT U5116 ( .A1(\ram[5][147] ), .A2(n5405), .A3(n5406), .A4(data[147]), .Y(n1488) );
  AO22X1_HVT U5117 ( .A1(\ram[5][146] ), .A2(n5405), .A3(n5406), .A4(data[146]), .Y(n1487) );
  AO22X1_HVT U5118 ( .A1(\ram[5][145] ), .A2(n5405), .A3(n5406), .A4(data[145]), .Y(n1486) );
  AO22X1_HVT U5119 ( .A1(\ram[5][144] ), .A2(n5405), .A3(n5406), .A4(data[144]), .Y(n1485) );
  AO22X1_HVT U5120 ( .A1(\ram[5][143] ), .A2(n5405), .A3(n5406), .A4(data[143]), .Y(n1484) );
  AO22X1_HVT U5121 ( .A1(\ram[5][142] ), .A2(n5405), .A3(n5406), .A4(data[142]), .Y(n1483) );
  AO22X1_HVT U5122 ( .A1(\ram[5][141] ), .A2(n5405), .A3(n5406), .A4(data[141]), .Y(n1482) );
  AO22X1_HVT U5123 ( .A1(\ram[5][140] ), .A2(n5405), .A3(n5406), .A4(data[140]), .Y(n1481) );
  AO22X1_HVT U5124 ( .A1(\ram[5][139] ), .A2(n5405), .A3(n5406), .A4(data[139]), .Y(n1480) );
  AO22X1_HVT U5125 ( .A1(\ram[0][87] ), .A2(n5360), .A3(data[87]), .A4(n5361), 
        .Y(n148) );
  AO22X1_HVT U5126 ( .A1(\ram[5][138] ), .A2(n5405), .A3(n5406), .A4(data[138]), .Y(n1479) );
  AO22X1_HVT U5127 ( .A1(\ram[5][137] ), .A2(n5405), .A3(n5406), .A4(data[137]), .Y(n1478) );
  AO22X1_HVT U5128 ( .A1(\ram[5][136] ), .A2(n5405), .A3(n5406), .A4(data[136]), .Y(n1477) );
  AO22X1_HVT U5129 ( .A1(\ram[5][135] ), .A2(n5405), .A3(n5406), .A4(data[135]), .Y(n1476) );
  AO22X1_HVT U5130 ( .A1(\ram[5][134] ), .A2(n5405), .A3(n5406), .A4(data[134]), .Y(n1475) );
  AO22X1_HVT U5131 ( .A1(\ram[5][133] ), .A2(n5405), .A3(n5406), .A4(data[133]), .Y(n1474) );
  AO22X1_HVT U5132 ( .A1(\ram[5][132] ), .A2(n5405), .A3(n5406), .A4(data[132]), .Y(n1473) );
  AO22X1_HVT U5133 ( .A1(\ram[5][131] ), .A2(n5405), .A3(n5406), .A4(data[131]), .Y(n1472) );
  AO22X1_HVT U5134 ( .A1(\ram[5][130] ), .A2(n5405), .A3(n5406), .A4(data[130]), .Y(n1471) );
  AO22X1_HVT U5135 ( .A1(\ram[5][129] ), .A2(n5405), .A3(n5406), .A4(data[129]), .Y(n1470) );
  AO22X1_HVT U5136 ( .A1(\ram[0][86] ), .A2(n5360), .A3(data[86]), .A4(n5361), 
        .Y(n147) );
  AO22X1_HVT U5137 ( .A1(\ram[5][128] ), .A2(n5405), .A3(n5406), .A4(data[128]), .Y(n1469) );
  AO22X1_HVT U5138 ( .A1(\ram[5][127] ), .A2(n5405), .A3(n5406), .A4(data[127]), .Y(n1468) );
  AO22X1_HVT U5139 ( .A1(\ram[5][126] ), .A2(n5405), .A3(n5406), .A4(data[126]), .Y(n1467) );
  AO22X1_HVT U5140 ( .A1(\ram[5][125] ), .A2(n5405), .A3(n5406), .A4(data[125]), .Y(n1466) );
  AO22X1_HVT U5141 ( .A1(\ram[5][124] ), .A2(n5405), .A3(n5406), .A4(data[124]), .Y(n1465) );
  AO22X1_HVT U5142 ( .A1(\ram[5][123] ), .A2(n5405), .A3(n5406), .A4(data[123]), .Y(n1464) );
  AO22X1_HVT U5143 ( .A1(\ram[5][122] ), .A2(n5405), .A3(n5406), .A4(data[122]), .Y(n1463) );
  AO22X1_HVT U5144 ( .A1(\ram[5][121] ), .A2(n5405), .A3(n5406), .A4(data[121]), .Y(n1462) );
  AO22X1_HVT U5145 ( .A1(\ram[5][120] ), .A2(n5405), .A3(n5406), .A4(data[120]), .Y(n1461) );
  AO22X1_HVT U5146 ( .A1(\ram[5][119] ), .A2(n5405), .A3(n5406), .A4(data[119]), .Y(n1460) );
  AO22X1_HVT U5147 ( .A1(\ram[0][85] ), .A2(n5360), .A3(data[85]), .A4(n5361), 
        .Y(n146) );
  AO22X1_HVT U5148 ( .A1(\ram[5][118] ), .A2(n5405), .A3(n5406), .A4(data[118]), .Y(n1459) );
  AO22X1_HVT U5149 ( .A1(\ram[5][117] ), .A2(n5405), .A3(n5406), .A4(data[117]), .Y(n1458) );
  AO22X1_HVT U5150 ( .A1(\ram[5][116] ), .A2(n5405), .A3(n5406), .A4(data[116]), .Y(n1457) );
  AO22X1_HVT U5151 ( .A1(\ram[5][115] ), .A2(n5405), .A3(n5406), .A4(data[115]), .Y(n1456) );
  AO22X1_HVT U5152 ( .A1(\ram[5][114] ), .A2(n5405), .A3(n5406), .A4(data[114]), .Y(n1455) );
  AO22X1_HVT U5153 ( .A1(\ram[5][113] ), .A2(n5405), .A3(n5406), .A4(data[113]), .Y(n1454) );
  AO22X1_HVT U5154 ( .A1(\ram[5][112] ), .A2(n5405), .A3(n5406), .A4(data[112]), .Y(n1453) );
  AO22X1_HVT U5155 ( .A1(\ram[5][111] ), .A2(n5405), .A3(n5406), .A4(data[111]), .Y(n1452) );
  AO22X1_HVT U5156 ( .A1(\ram[5][110] ), .A2(n5405), .A3(n5406), .A4(data[110]), .Y(n1451) );
  AO22X1_HVT U5157 ( .A1(\ram[5][109] ), .A2(n5405), .A3(n5406), .A4(data[109]), .Y(n1450) );
  AO22X1_HVT U5158 ( .A1(\ram[0][84] ), .A2(n5360), .A3(data[84]), .A4(n5361), 
        .Y(n145) );
  AO22X1_HVT U5159 ( .A1(\ram[5][108] ), .A2(n5405), .A3(n5406), .A4(data[108]), .Y(n1449) );
  AO22X1_HVT U5160 ( .A1(\ram[5][107] ), .A2(n5405), .A3(n5406), .A4(data[107]), .Y(n1448) );
  AO22X1_HVT U5161 ( .A1(\ram[5][106] ), .A2(n5405), .A3(n5406), .A4(data[106]), .Y(n1447) );
  AO22X1_HVT U5162 ( .A1(\ram[5][105] ), .A2(n5405), .A3(n5406), .A4(data[105]), .Y(n1446) );
  AO22X1_HVT U5163 ( .A1(\ram[5][104] ), .A2(n5405), .A3(n5406), .A4(data[104]), .Y(n1445) );
  AO22X1_HVT U5164 ( .A1(\ram[5][103] ), .A2(n5405), .A3(n5406), .A4(data[103]), .Y(n1444) );
  AO22X1_HVT U5165 ( .A1(\ram[5][102] ), .A2(n5405), .A3(n5406), .A4(data[102]), .Y(n1443) );
  AO22X1_HVT U5166 ( .A1(\ram[5][101] ), .A2(n5405), .A3(n5406), .A4(data[101]), .Y(n1442) );
  AO22X1_HVT U5167 ( .A1(\ram[5][100] ), .A2(n5405), .A3(n5406), .A4(data[100]), .Y(n1441) );
  AO22X1_HVT U5168 ( .A1(\ram[5][99] ), .A2(n5405), .A3(n5406), .A4(data[99]), 
        .Y(n1440) );
  AO22X1_HVT U5169 ( .A1(\ram[0][83] ), .A2(n5360), .A3(data[83]), .A4(n5361), 
        .Y(n144) );
  AO22X1_HVT U5170 ( .A1(\ram[5][98] ), .A2(n5405), .A3(n5406), .A4(data[98]), 
        .Y(n1439) );
  AO22X1_HVT U5171 ( .A1(\ram[5][97] ), .A2(n5405), .A3(n5406), .A4(data[97]), 
        .Y(n1438) );
  AO22X1_HVT U5172 ( .A1(\ram[5][96] ), .A2(n5405), .A3(n5406), .A4(data[96]), 
        .Y(n1437) );
  AO22X1_HVT U5173 ( .A1(\ram[5][95] ), .A2(n5405), .A3(n5406), .A4(data[95]), 
        .Y(n1436) );
  AO22X1_HVT U5174 ( .A1(\ram[5][94] ), .A2(n5405), .A3(n5406), .A4(data[94]), 
        .Y(n1435) );
  AO22X1_HVT U5175 ( .A1(\ram[5][93] ), .A2(n5405), .A3(n5406), .A4(data[93]), 
        .Y(n1434) );
  AO22X1_HVT U5176 ( .A1(\ram[5][92] ), .A2(n5405), .A3(n5406), .A4(data[92]), 
        .Y(n1433) );
  AO22X1_HVT U5177 ( .A1(\ram[5][91] ), .A2(n5405), .A3(n5406), .A4(data[91]), 
        .Y(n1432) );
  AO22X1_HVT U5178 ( .A1(\ram[5][90] ), .A2(n5405), .A3(n5406), .A4(data[90]), 
        .Y(n1431) );
  AO22X1_HVT U5179 ( .A1(\ram[5][89] ), .A2(n5405), .A3(n5406), .A4(data[89]), 
        .Y(n1430) );
  AO22X1_HVT U5180 ( .A1(\ram[0][82] ), .A2(n5360), .A3(data[82]), .A4(n5361), 
        .Y(n143) );
  AO22X1_HVT U5181 ( .A1(\ram[5][88] ), .A2(n5405), .A3(n5406), .A4(data[88]), 
        .Y(n1429) );
  AO22X1_HVT U5182 ( .A1(\ram[5][87] ), .A2(n5405), .A3(n5406), .A4(data[87]), 
        .Y(n1428) );
  AO22X1_HVT U5183 ( .A1(\ram[5][86] ), .A2(n5405), .A3(n5406), .A4(data[86]), 
        .Y(n1427) );
  AO22X1_HVT U5184 ( .A1(\ram[5][85] ), .A2(n5405), .A3(n5406), .A4(data[85]), 
        .Y(n1426) );
  AO22X1_HVT U5185 ( .A1(\ram[5][84] ), .A2(n5405), .A3(n5406), .A4(data[84]), 
        .Y(n1425) );
  AO22X1_HVT U5186 ( .A1(\ram[5][83] ), .A2(n5405), .A3(n5406), .A4(data[83]), 
        .Y(n1424) );
  AO22X1_HVT U5187 ( .A1(\ram[5][82] ), .A2(n5405), .A3(n5406), .A4(data[82]), 
        .Y(n1423) );
  AO22X1_HVT U5188 ( .A1(\ram[5][81] ), .A2(n5405), .A3(n5406), .A4(data[81]), 
        .Y(n1422) );
  AO22X1_HVT U5189 ( .A1(\ram[5][80] ), .A2(n5405), .A3(n5406), .A4(data[80]), 
        .Y(n1421) );
  AO22X1_HVT U5190 ( .A1(\ram[5][79] ), .A2(n5405), .A3(n5406), .A4(data[79]), 
        .Y(n1420) );
  AO22X1_HVT U5191 ( .A1(\ram[0][81] ), .A2(n5360), .A3(data[81]), .A4(n5361), 
        .Y(n142) );
  AO22X1_HVT U5192 ( .A1(\ram[5][78] ), .A2(n5405), .A3(n5406), .A4(data[78]), 
        .Y(n1419) );
  AO22X1_HVT U5193 ( .A1(\ram[5][77] ), .A2(n5405), .A3(n5406), .A4(data[77]), 
        .Y(n1418) );
  AO22X1_HVT U5194 ( .A1(\ram[5][76] ), .A2(n5405), .A3(n5406), .A4(data[76]), 
        .Y(n1417) );
  AO22X1_HVT U5195 ( .A1(\ram[5][75] ), .A2(n5405), .A3(n5406), .A4(data[75]), 
        .Y(n1416) );
  AO22X1_HVT U5196 ( .A1(\ram[5][74] ), .A2(n5405), .A3(n5406), .A4(data[74]), 
        .Y(n1415) );
  AO22X1_HVT U5197 ( .A1(\ram[5][73] ), .A2(n5405), .A3(n5406), .A4(data[73]), 
        .Y(n1414) );
  AO22X1_HVT U5198 ( .A1(\ram[5][72] ), .A2(n5405), .A3(n5406), .A4(data[72]), 
        .Y(n1413) );
  AO22X1_HVT U5199 ( .A1(\ram[5][71] ), .A2(n5405), .A3(n5406), .A4(data[71]), 
        .Y(n1412) );
  AO22X1_HVT U5200 ( .A1(\ram[5][70] ), .A2(n5405), .A3(n5406), .A4(data[70]), 
        .Y(n1411) );
  AO22X1_HVT U5201 ( .A1(\ram[5][69] ), .A2(n5405), .A3(n5406), .A4(data[69]), 
        .Y(n1410) );
  AO22X1_HVT U5202 ( .A1(\ram[0][80] ), .A2(n5360), .A3(data[80]), .A4(n5361), 
        .Y(n141) );
  AO22X1_HVT U5203 ( .A1(\ram[5][68] ), .A2(n5405), .A3(n5406), .A4(data[68]), 
        .Y(n1409) );
  AO22X1_HVT U5204 ( .A1(\ram[5][67] ), .A2(n5405), .A3(n5406), .A4(data[67]), 
        .Y(n1408) );
  AO22X1_HVT U5205 ( .A1(\ram[5][66] ), .A2(n5405), .A3(n5406), .A4(data[66]), 
        .Y(n1407) );
  AO22X1_HVT U5206 ( .A1(\ram[5][65] ), .A2(n5405), .A3(n5406), .A4(data[65]), 
        .Y(n1406) );
  AO22X1_HVT U5207 ( .A1(\ram[5][64] ), .A2(n5405), .A3(n5406), .A4(data[64]), 
        .Y(n1405) );
  AO22X1_HVT U5208 ( .A1(\ram[5][63] ), .A2(n5405), .A3(n5406), .A4(data[63]), 
        .Y(n1404) );
  AO22X1_HVT U5209 ( .A1(\ram[5][62] ), .A2(n5405), .A3(n5406), .A4(data[62]), 
        .Y(n1403) );
  AO22X1_HVT U5210 ( .A1(\ram[5][61] ), .A2(n5405), .A3(n5406), .A4(data[61]), 
        .Y(n1402) );
  AO22X1_HVT U5211 ( .A1(\ram[5][60] ), .A2(n5405), .A3(n5406), .A4(data[60]), 
        .Y(n1401) );
  AO22X1_HVT U5212 ( .A1(\ram[5][59] ), .A2(n5405), .A3(n5406), .A4(data[59]), 
        .Y(n1400) );
  AO22X1_HVT U5213 ( .A1(\ram[0][79] ), .A2(n5360), .A3(data[79]), .A4(n5361), 
        .Y(n140) );
  AO22X1_HVT U5214 ( .A1(\ram[5][58] ), .A2(n5405), .A3(n5406), .A4(data[58]), 
        .Y(n1399) );
  AO22X1_HVT U5215 ( .A1(\ram[5][57] ), .A2(n5405), .A3(n5406), .A4(data[57]), 
        .Y(n1398) );
  AO22X1_HVT U5216 ( .A1(\ram[5][56] ), .A2(n5405), .A3(n5406), .A4(data[56]), 
        .Y(n1397) );
  AO22X1_HVT U5217 ( .A1(\ram[5][55] ), .A2(n5405), .A3(n5406), .A4(data[55]), 
        .Y(n1396) );
  AO22X1_HVT U5218 ( .A1(\ram[5][54] ), .A2(n5405), .A3(n5406), .A4(data[54]), 
        .Y(n1395) );
  AO22X1_HVT U5219 ( .A1(\ram[5][53] ), .A2(n5405), .A3(n5406), .A4(data[53]), 
        .Y(n1394) );
  AO22X1_HVT U5220 ( .A1(\ram[5][52] ), .A2(n5405), .A3(n5406), .A4(data[52]), 
        .Y(n1393) );
  AO22X1_HVT U5221 ( .A1(\ram[5][51] ), .A2(n5405), .A3(n5406), .A4(data[51]), 
        .Y(n1392) );
  AO22X1_HVT U5222 ( .A1(\ram[5][50] ), .A2(n5405), .A3(n5406), .A4(data[50]), 
        .Y(n1391) );
  AO22X1_HVT U5223 ( .A1(\ram[5][49] ), .A2(n5405), .A3(n5406), .A4(data[49]), 
        .Y(n1390) );
  AO22X1_HVT U5224 ( .A1(\ram[0][78] ), .A2(n5360), .A3(data[78]), .A4(n5361), 
        .Y(n139) );
  AO22X1_HVT U5225 ( .A1(\ram[5][48] ), .A2(n5405), .A3(n5406), .A4(data[48]), 
        .Y(n1389) );
  AO22X1_HVT U5226 ( .A1(\ram[5][47] ), .A2(n5405), .A3(n5406), .A4(data[47]), 
        .Y(n1388) );
  AO22X1_HVT U5227 ( .A1(\ram[5][46] ), .A2(n5405), .A3(n5406), .A4(data[46]), 
        .Y(n1387) );
  AO22X1_HVT U5228 ( .A1(\ram[5][45] ), .A2(n5405), .A3(n5406), .A4(data[45]), 
        .Y(n1386) );
  AO22X1_HVT U5229 ( .A1(\ram[5][44] ), .A2(n5405), .A3(n5406), .A4(data[44]), 
        .Y(n1385) );
  AO22X1_HVT U5230 ( .A1(\ram[5][43] ), .A2(n5405), .A3(n5406), .A4(data[43]), 
        .Y(n1384) );
  AO22X1_HVT U5231 ( .A1(\ram[5][42] ), .A2(n5405), .A3(n5406), .A4(data[42]), 
        .Y(n1383) );
  AO22X1_HVT U5232 ( .A1(\ram[5][41] ), .A2(n5405), .A3(n5406), .A4(data[41]), 
        .Y(n1382) );
  AO22X1_HVT U5233 ( .A1(\ram[5][40] ), .A2(n5405), .A3(n5406), .A4(data[40]), 
        .Y(n1381) );
  AO22X1_HVT U5234 ( .A1(\ram[5][39] ), .A2(n5405), .A3(n5406), .A4(data[39]), 
        .Y(n1380) );
  AO22X1_HVT U5235 ( .A1(\ram[0][77] ), .A2(n5360), .A3(data[77]), .A4(n5361), 
        .Y(n138) );
  AO22X1_HVT U5236 ( .A1(\ram[5][38] ), .A2(n5405), .A3(n5406), .A4(data[38]), 
        .Y(n1379) );
  AO22X1_HVT U5237 ( .A1(\ram[5][37] ), .A2(n5405), .A3(n5406), .A4(data[37]), 
        .Y(n1378) );
  AO22X1_HVT U5238 ( .A1(\ram[5][36] ), .A2(n5405), .A3(n5406), .A4(data[36]), 
        .Y(n1377) );
  AO22X1_HVT U5239 ( .A1(\ram[5][35] ), .A2(n5405), .A3(n5406), .A4(data[35]), 
        .Y(n1376) );
  AO22X1_HVT U5240 ( .A1(\ram[5][34] ), .A2(n5405), .A3(n5406), .A4(data[34]), 
        .Y(n1375) );
  AO22X1_HVT U5241 ( .A1(\ram[5][33] ), .A2(n5405), .A3(n5406), .A4(data[33]), 
        .Y(n1374) );
  AO22X1_HVT U5242 ( .A1(\ram[5][32] ), .A2(n5405), .A3(n5406), .A4(data[32]), 
        .Y(n1373) );
  AO22X1_HVT U5243 ( .A1(\ram[5][31] ), .A2(n5405), .A3(n5406), .A4(data[31]), 
        .Y(n1372) );
  AO22X1_HVT U5244 ( .A1(\ram[5][30] ), .A2(n5405), .A3(n5406), .A4(data[30]), 
        .Y(n1371) );
  AO22X1_HVT U5245 ( .A1(\ram[5][29] ), .A2(n5405), .A3(n5406), .A4(data[29]), 
        .Y(n1370) );
  AO22X1_HVT U5246 ( .A1(\ram[0][76] ), .A2(n5360), .A3(data[76]), .A4(n5361), 
        .Y(n137) );
  AO22X1_HVT U5247 ( .A1(\ram[5][28] ), .A2(n5405), .A3(n5406), .A4(data[28]), 
        .Y(n1369) );
  AO22X1_HVT U5248 ( .A1(\ram[5][27] ), .A2(n5405), .A3(n5406), .A4(data[27]), 
        .Y(n1368) );
  AO22X1_HVT U5249 ( .A1(\ram[5][26] ), .A2(n5405), .A3(n5406), .A4(data[26]), 
        .Y(n1367) );
  AO22X1_HVT U5250 ( .A1(\ram[5][25] ), .A2(n5405), .A3(n5406), .A4(data[25]), 
        .Y(n1366) );
  AO22X1_HVT U5251 ( .A1(\ram[5][24] ), .A2(n5405), .A3(n5406), .A4(data[24]), 
        .Y(n1365) );
  AO22X1_HVT U5252 ( .A1(\ram[5][23] ), .A2(n5405), .A3(n5406), .A4(data[23]), 
        .Y(n1364) );
  AO22X1_HVT U5253 ( .A1(\ram[5][22] ), .A2(n5405), .A3(n5406), .A4(data[22]), 
        .Y(n1363) );
  AO22X1_HVT U5254 ( .A1(\ram[5][21] ), .A2(n5405), .A3(n5406), .A4(data[21]), 
        .Y(n1362) );
  AO22X1_HVT U5255 ( .A1(\ram[5][20] ), .A2(n5405), .A3(n5406), .A4(data[20]), 
        .Y(n1361) );
  AO22X1_HVT U5256 ( .A1(\ram[5][19] ), .A2(n5405), .A3(n5406), .A4(data[19]), 
        .Y(n1360) );
  AO22X1_HVT U5257 ( .A1(\ram[0][75] ), .A2(n5360), .A3(data[75]), .A4(n5361), 
        .Y(n136) );
  AO22X1_HVT U5258 ( .A1(\ram[5][18] ), .A2(n5405), .A3(n5406), .A4(data[18]), 
        .Y(n1359) );
  AO22X1_HVT U5259 ( .A1(\ram[5][17] ), .A2(n5405), .A3(n5406), .A4(data[17]), 
        .Y(n1358) );
  AO22X1_HVT U5260 ( .A1(\ram[5][16] ), .A2(n5405), .A3(n5406), .A4(data[16]), 
        .Y(n1357) );
  AO22X1_HVT U5261 ( .A1(\ram[5][15] ), .A2(n5405), .A3(n5406), .A4(data[15]), 
        .Y(n1356) );
  AO22X1_HVT U5262 ( .A1(\ram[5][14] ), .A2(n5405), .A3(n5406), .A4(data[14]), 
        .Y(n1355) );
  AO22X1_HVT U5263 ( .A1(\ram[5][13] ), .A2(n5405), .A3(n5406), .A4(data[13]), 
        .Y(n1354) );
  AO22X1_HVT U5264 ( .A1(\ram[5][12] ), .A2(n5405), .A3(n5406), .A4(data[12]), 
        .Y(n1353) );
  AO22X1_HVT U5265 ( .A1(\ram[5][11] ), .A2(n5405), .A3(n5406), .A4(data[11]), 
        .Y(n1352) );
  AO22X1_HVT U5266 ( .A1(\ram[5][10] ), .A2(n5405), .A3(n5406), .A4(data[10]), 
        .Y(n1351) );
  AO22X1_HVT U5267 ( .A1(\ram[5][9] ), .A2(n5405), .A3(n5406), .A4(data[9]), 
        .Y(n1350) );
  AO22X1_HVT U5268 ( .A1(\ram[0][74] ), .A2(n5360), .A3(data[74]), .A4(n5361), 
        .Y(n135) );
  AO22X1_HVT U5269 ( .A1(\ram[5][8] ), .A2(n5405), .A3(n5406), .A4(data[8]), 
        .Y(n1349) );
  AO22X1_HVT U5270 ( .A1(\ram[5][7] ), .A2(n5405), .A3(n5406), .A4(data[7]), 
        .Y(n1348) );
  AO22X1_HVT U5271 ( .A1(\ram[5][6] ), .A2(n5405), .A3(n5406), .A4(data[6]), 
        .Y(n1347) );
  AO22X1_HVT U5272 ( .A1(\ram[5][5] ), .A2(n5405), .A3(n5406), .A4(data[5]), 
        .Y(n1346) );
  AO22X1_HVT U5273 ( .A1(\ram[5][4] ), .A2(n5405), .A3(n5406), .A4(data[4]), 
        .Y(n1345) );
  AO22X1_HVT U5274 ( .A1(\ram[5][3] ), .A2(n5405), .A3(n5406), .A4(data[3]), 
        .Y(n1344) );
  AO22X1_HVT U5275 ( .A1(\ram[5][2] ), .A2(n5405), .A3(n5406), .A4(data[2]), 
        .Y(n1343) );
  AO22X1_HVT U5276 ( .A1(\ram[5][1] ), .A2(n5405), .A3(n5406), .A4(data[1]), 
        .Y(n1342) );
  AO22X1_HVT U5277 ( .A1(\ram[5][0] ), .A2(n5405), .A3(n5406), .A4(data[0]), 
        .Y(n1341) );
  INVX0_HVT U5278 ( .A(n5407), .Y(n5406) );
  AND2X1_HVT U5279 ( .A1(n5407), .A2(n5365), .Y(n5405) );
  NAND3X0_HVT U5280 ( .A1(n4182), .A2(n4278), .A3(n5401), .Y(n5407) );
  AO22X1_HVT U5281 ( .A1(\ram[4][255] ), .A2(n5408), .A3(n5409), .A4(data[255]), .Y(n1340) );
  AO22X1_HVT U5282 ( .A1(\ram[0][73] ), .A2(n5360), .A3(data[73]), .A4(n5361), 
        .Y(n134) );
  AO22X1_HVT U5283 ( .A1(\ram[4][254] ), .A2(n5408), .A3(n5409), .A4(data[254]), .Y(n1339) );
  AO22X1_HVT U5284 ( .A1(\ram[4][253] ), .A2(n5408), .A3(n5409), .A4(data[253]), .Y(n1338) );
  AO22X1_HVT U5285 ( .A1(\ram[4][252] ), .A2(n5408), .A3(n5409), .A4(data[252]), .Y(n1337) );
  AO22X1_HVT U5286 ( .A1(\ram[4][251] ), .A2(n5408), .A3(n5409), .A4(data[251]), .Y(n1336) );
  AO22X1_HVT U5287 ( .A1(\ram[4][250] ), .A2(n5408), .A3(n5409), .A4(data[250]), .Y(n1335) );
  AO22X1_HVT U5288 ( .A1(\ram[4][249] ), .A2(n5408), .A3(n5409), .A4(data[249]), .Y(n1334) );
  AO22X1_HVT U5289 ( .A1(\ram[4][248] ), .A2(n5408), .A3(n5409), .A4(data[248]), .Y(n1333) );
  AO22X1_HVT U5290 ( .A1(\ram[4][247] ), .A2(n5408), .A3(n5409), .A4(data[247]), .Y(n1332) );
  AO22X1_HVT U5291 ( .A1(\ram[4][246] ), .A2(n5408), .A3(n5409), .A4(data[246]), .Y(n1331) );
  AO22X1_HVT U5292 ( .A1(\ram[4][245] ), .A2(n5408), .A3(n5409), .A4(data[245]), .Y(n1330) );
  AO22X1_HVT U5293 ( .A1(\ram[0][72] ), .A2(n5360), .A3(data[72]), .A4(n5361), 
        .Y(n133) );
  AO22X1_HVT U5294 ( .A1(\ram[4][244] ), .A2(n5408), .A3(n5409), .A4(data[244]), .Y(n1329) );
  AO22X1_HVT U5295 ( .A1(\ram[4][243] ), .A2(n5408), .A3(n5409), .A4(data[243]), .Y(n1328) );
  AO22X1_HVT U5296 ( .A1(\ram[4][242] ), .A2(n5408), .A3(n5409), .A4(data[242]), .Y(n1327) );
  AO22X1_HVT U5297 ( .A1(\ram[4][241] ), .A2(n5408), .A3(n5409), .A4(data[241]), .Y(n1326) );
  AO22X1_HVT U5298 ( .A1(\ram[4][240] ), .A2(n5408), .A3(n5409), .A4(data[240]), .Y(n1325) );
  AO22X1_HVT U5299 ( .A1(\ram[4][239] ), .A2(n5408), .A3(n5409), .A4(data[239]), .Y(n1324) );
  AO22X1_HVT U5300 ( .A1(\ram[4][238] ), .A2(n5408), .A3(n5409), .A4(data[238]), .Y(n1323) );
  AO22X1_HVT U5301 ( .A1(\ram[4][237] ), .A2(n5408), .A3(n5409), .A4(data[237]), .Y(n1322) );
  AO22X1_HVT U5302 ( .A1(\ram[4][236] ), .A2(n5408), .A3(n5409), .A4(data[236]), .Y(n1321) );
  AO22X1_HVT U5303 ( .A1(\ram[4][235] ), .A2(n5408), .A3(n5409), .A4(data[235]), .Y(n1320) );
  AO22X1_HVT U5304 ( .A1(\ram[0][71] ), .A2(n5360), .A3(data[71]), .A4(n5361), 
        .Y(n132) );
  AO22X1_HVT U5305 ( .A1(\ram[4][234] ), .A2(n5408), .A3(n5409), .A4(data[234]), .Y(n1319) );
  AO22X1_HVT U5306 ( .A1(\ram[4][233] ), .A2(n5408), .A3(n5409), .A4(data[233]), .Y(n1318) );
  AO22X1_HVT U5307 ( .A1(\ram[4][232] ), .A2(n5408), .A3(n5409), .A4(data[232]), .Y(n1317) );
  AO22X1_HVT U5308 ( .A1(\ram[4][231] ), .A2(n5408), .A3(n5409), .A4(data[231]), .Y(n1316) );
  AO22X1_HVT U5309 ( .A1(\ram[4][230] ), .A2(n5408), .A3(n5409), .A4(data[230]), .Y(n1315) );
  AO22X1_HVT U5310 ( .A1(\ram[4][229] ), .A2(n5408), .A3(n5409), .A4(data[229]), .Y(n1314) );
  AO22X1_HVT U5311 ( .A1(\ram[4][228] ), .A2(n5408), .A3(n5409), .A4(data[228]), .Y(n1313) );
  AO22X1_HVT U5312 ( .A1(\ram[4][227] ), .A2(n5408), .A3(n5409), .A4(data[227]), .Y(n1312) );
  AO22X1_HVT U5313 ( .A1(\ram[4][226] ), .A2(n5408), .A3(n5409), .A4(data[226]), .Y(n1311) );
  AO22X1_HVT U5314 ( .A1(\ram[4][225] ), .A2(n5408), .A3(n5409), .A4(data[225]), .Y(n1310) );
  AO22X1_HVT U5315 ( .A1(\ram[0][70] ), .A2(n5360), .A3(data[70]), .A4(n5361), 
        .Y(n131) );
  AO22X1_HVT U5316 ( .A1(\ram[4][224] ), .A2(n5408), .A3(n5409), .A4(data[224]), .Y(n1309) );
  AO22X1_HVT U5317 ( .A1(\ram[4][223] ), .A2(n5408), .A3(n5409), .A4(data[223]), .Y(n1308) );
  AO22X1_HVT U5318 ( .A1(\ram[4][222] ), .A2(n5408), .A3(n5409), .A4(data[222]), .Y(n1307) );
  AO22X1_HVT U5319 ( .A1(\ram[4][221] ), .A2(n5408), .A3(n5409), .A4(data[221]), .Y(n1306) );
  AO22X1_HVT U5320 ( .A1(\ram[4][220] ), .A2(n5408), .A3(n5409), .A4(data[220]), .Y(n1305) );
  AO22X1_HVT U5321 ( .A1(\ram[4][219] ), .A2(n5408), .A3(n5409), .A4(data[219]), .Y(n1304) );
  AO22X1_HVT U5322 ( .A1(\ram[4][218] ), .A2(n5408), .A3(n5409), .A4(data[218]), .Y(n1303) );
  AO22X1_HVT U5323 ( .A1(\ram[4][217] ), .A2(n5408), .A3(n5409), .A4(data[217]), .Y(n1302) );
  AO22X1_HVT U5324 ( .A1(\ram[4][216] ), .A2(n5408), .A3(n5409), .A4(data[216]), .Y(n1301) );
  AO22X1_HVT U5325 ( .A1(\ram[4][215] ), .A2(n5408), .A3(n5409), .A4(data[215]), .Y(n1300) );
  AO22X1_HVT U5326 ( .A1(\ram[0][69] ), .A2(n5360), .A3(data[69]), .A4(n5361), 
        .Y(n130) );
  AO22X1_HVT U5327 ( .A1(\ram[4][214] ), .A2(n5408), .A3(n5409), .A4(data[214]), .Y(n1299) );
  AO22X1_HVT U5328 ( .A1(\ram[4][213] ), .A2(n5408), .A3(n5409), .A4(data[213]), .Y(n1298) );
  AO22X1_HVT U5329 ( .A1(\ram[4][212] ), .A2(n5408), .A3(n5409), .A4(data[212]), .Y(n1297) );
  AO22X1_HVT U5330 ( .A1(\ram[4][211] ), .A2(n5408), .A3(n5409), .A4(data[211]), .Y(n1296) );
  AO22X1_HVT U5331 ( .A1(\ram[4][210] ), .A2(n5408), .A3(n5409), .A4(data[210]), .Y(n1295) );
  AO22X1_HVT U5332 ( .A1(\ram[4][209] ), .A2(n5408), .A3(n5409), .A4(data[209]), .Y(n1294) );
  AO22X1_HVT U5333 ( .A1(\ram[4][208] ), .A2(n5408), .A3(n5409), .A4(data[208]), .Y(n1293) );
  AO22X1_HVT U5334 ( .A1(\ram[4][207] ), .A2(n5408), .A3(n5409), .A4(data[207]), .Y(n1292) );
  AO22X1_HVT U5335 ( .A1(\ram[4][206] ), .A2(n5408), .A3(n5409), .A4(data[206]), .Y(n1291) );
  AO22X1_HVT U5336 ( .A1(\ram[4][205] ), .A2(n5408), .A3(n5409), .A4(data[205]), .Y(n1290) );
  AO22X1_HVT U5337 ( .A1(\ram[0][68] ), .A2(n5360), .A3(data[68]), .A4(n5361), 
        .Y(n129) );
  AO22X1_HVT U5338 ( .A1(\ram[4][204] ), .A2(n5408), .A3(n5409), .A4(data[204]), .Y(n1289) );
  AO22X1_HVT U5339 ( .A1(\ram[4][203] ), .A2(n5408), .A3(n5409), .A4(data[203]), .Y(n1288) );
  AO22X1_HVT U5340 ( .A1(\ram[4][202] ), .A2(n5408), .A3(n5409), .A4(data[202]), .Y(n1287) );
  AO22X1_HVT U5341 ( .A1(\ram[4][201] ), .A2(n5408), .A3(n5409), .A4(data[201]), .Y(n1286) );
  AO22X1_HVT U5342 ( .A1(\ram[4][200] ), .A2(n5408), .A3(n5409), .A4(data[200]), .Y(n1285) );
  AO22X1_HVT U5343 ( .A1(\ram[4][199] ), .A2(n5408), .A3(n5409), .A4(data[199]), .Y(n1284) );
  AO22X1_HVT U5344 ( .A1(\ram[4][198] ), .A2(n5408), .A3(n5409), .A4(data[198]), .Y(n1283) );
  AO22X1_HVT U5345 ( .A1(\ram[4][197] ), .A2(n5408), .A3(n5409), .A4(data[197]), .Y(n1282) );
  AO22X1_HVT U5346 ( .A1(\ram[4][196] ), .A2(n5408), .A3(n5409), .A4(data[196]), .Y(n1281) );
  AO22X1_HVT U5347 ( .A1(\ram[4][195] ), .A2(n5408), .A3(n5409), .A4(data[195]), .Y(n1280) );
  AO22X1_HVT U5348 ( .A1(\ram[0][67] ), .A2(n5360), .A3(data[67]), .A4(n5361), 
        .Y(n128) );
  AO22X1_HVT U5349 ( .A1(\ram[4][194] ), .A2(n5408), .A3(n5409), .A4(data[194]), .Y(n1279) );
  AO22X1_HVT U5350 ( .A1(\ram[4][193] ), .A2(n5408), .A3(n5409), .A4(data[193]), .Y(n1278) );
  AO22X1_HVT U5351 ( .A1(\ram[4][192] ), .A2(n5408), .A3(n5409), .A4(data[192]), .Y(n1277) );
  AO22X1_HVT U5352 ( .A1(\ram[4][191] ), .A2(n5408), .A3(n5409), .A4(data[191]), .Y(n1276) );
  AO22X1_HVT U5353 ( .A1(\ram[4][190] ), .A2(n5408), .A3(n5409), .A4(data[190]), .Y(n1275) );
  AO22X1_HVT U5354 ( .A1(\ram[4][189] ), .A2(n5408), .A3(n5409), .A4(data[189]), .Y(n1274) );
  AO22X1_HVT U5355 ( .A1(\ram[4][188] ), .A2(n5408), .A3(n5409), .A4(data[188]), .Y(n1273) );
  AO22X1_HVT U5356 ( .A1(\ram[4][187] ), .A2(n5408), .A3(n5409), .A4(data[187]), .Y(n1272) );
  AO22X1_HVT U5357 ( .A1(\ram[4][186] ), .A2(n5408), .A3(n5409), .A4(data[186]), .Y(n1271) );
  AO22X1_HVT U5358 ( .A1(\ram[4][185] ), .A2(n5408), .A3(n5409), .A4(data[185]), .Y(n1270) );
  AO22X1_HVT U5359 ( .A1(\ram[0][66] ), .A2(n5360), .A3(data[66]), .A4(n5361), 
        .Y(n127) );
  AO22X1_HVT U5360 ( .A1(\ram[4][184] ), .A2(n5408), .A3(n5409), .A4(data[184]), .Y(n1269) );
  AO22X1_HVT U5361 ( .A1(\ram[4][183] ), .A2(n5408), .A3(n5409), .A4(data[183]), .Y(n1268) );
  AO22X1_HVT U5362 ( .A1(\ram[4][182] ), .A2(n5408), .A3(n5409), .A4(data[182]), .Y(n1267) );
  AO22X1_HVT U5363 ( .A1(\ram[4][181] ), .A2(n5408), .A3(n5409), .A4(data[181]), .Y(n1266) );
  AO22X1_HVT U5364 ( .A1(\ram[4][180] ), .A2(n5408), .A3(n5409), .A4(data[180]), .Y(n1265) );
  AO22X1_HVT U5365 ( .A1(\ram[4][179] ), .A2(n5408), .A3(n5409), .A4(data[179]), .Y(n1264) );
  AO22X1_HVT U5366 ( .A1(\ram[4][178] ), .A2(n5408), .A3(n5409), .A4(data[178]), .Y(n1263) );
  AO22X1_HVT U5367 ( .A1(\ram[4][177] ), .A2(n5408), .A3(n5409), .A4(data[177]), .Y(n1262) );
  AO22X1_HVT U5368 ( .A1(\ram[4][176] ), .A2(n5408), .A3(n5409), .A4(data[176]), .Y(n1261) );
  AO22X1_HVT U5369 ( .A1(\ram[4][175] ), .A2(n5408), .A3(n5409), .A4(data[175]), .Y(n1260) );
  AO22X1_HVT U5370 ( .A1(\ram[0][65] ), .A2(n5360), .A3(data[65]), .A4(n5361), 
        .Y(n126) );
  AO22X1_HVT U5371 ( .A1(\ram[4][174] ), .A2(n5408), .A3(n5409), .A4(data[174]), .Y(n1259) );
  AO22X1_HVT U5372 ( .A1(\ram[4][173] ), .A2(n5408), .A3(n5409), .A4(data[173]), .Y(n1258) );
  AO22X1_HVT U5373 ( .A1(\ram[4][172] ), .A2(n5408), .A3(n5409), .A4(data[172]), .Y(n1257) );
  AO22X1_HVT U5374 ( .A1(\ram[4][171] ), .A2(n5408), .A3(n5409), .A4(data[171]), .Y(n1256) );
  AO22X1_HVT U5375 ( .A1(\ram[4][170] ), .A2(n5408), .A3(n5409), .A4(data[170]), .Y(n1255) );
  AO22X1_HVT U5376 ( .A1(\ram[4][169] ), .A2(n5408), .A3(n5409), .A4(data[169]), .Y(n1254) );
  AO22X1_HVT U5377 ( .A1(\ram[4][168] ), .A2(n5408), .A3(n5409), .A4(data[168]), .Y(n1253) );
  AO22X1_HVT U5378 ( .A1(\ram[4][167] ), .A2(n5408), .A3(n5409), .A4(data[167]), .Y(n1252) );
  AO22X1_HVT U5379 ( .A1(\ram[4][166] ), .A2(n5408), .A3(n5409), .A4(data[166]), .Y(n1251) );
  AO22X1_HVT U5380 ( .A1(\ram[4][165] ), .A2(n5408), .A3(n5409), .A4(data[165]), .Y(n1250) );
  AO22X1_HVT U5381 ( .A1(\ram[0][64] ), .A2(n5360), .A3(data[64]), .A4(n5361), 
        .Y(n125) );
  AO22X1_HVT U5382 ( .A1(\ram[4][164] ), .A2(n5408), .A3(n5409), .A4(data[164]), .Y(n1249) );
  AO22X1_HVT U5383 ( .A1(\ram[4][163] ), .A2(n5408), .A3(n5409), .A4(data[163]), .Y(n1248) );
  AO22X1_HVT U5384 ( .A1(\ram[4][162] ), .A2(n5408), .A3(n5409), .A4(data[162]), .Y(n1247) );
  AO22X1_HVT U5385 ( .A1(\ram[4][161] ), .A2(n5408), .A3(n5409), .A4(data[161]), .Y(n1246) );
  AO22X1_HVT U5386 ( .A1(\ram[4][160] ), .A2(n5408), .A3(n5409), .A4(data[160]), .Y(n1245) );
  AO22X1_HVT U5387 ( .A1(\ram[4][159] ), .A2(n5408), .A3(n5409), .A4(data[159]), .Y(n1244) );
  AO22X1_HVT U5388 ( .A1(\ram[4][158] ), .A2(n5408), .A3(n5409), .A4(data[158]), .Y(n1243) );
  AO22X1_HVT U5389 ( .A1(\ram[4][157] ), .A2(n5408), .A3(n5409), .A4(data[157]), .Y(n1242) );
  AO22X1_HVT U5390 ( .A1(\ram[4][156] ), .A2(n5408), .A3(n5409), .A4(data[156]), .Y(n1241) );
  AO22X1_HVT U5391 ( .A1(\ram[4][155] ), .A2(n5408), .A3(n5409), .A4(data[155]), .Y(n1240) );
  AO22X1_HVT U5392 ( .A1(\ram[0][63] ), .A2(n5360), .A3(data[63]), .A4(n5361), 
        .Y(n124) );
  AO22X1_HVT U5393 ( .A1(\ram[4][154] ), .A2(n5408), .A3(n5409), .A4(data[154]), .Y(n1239) );
  AO22X1_HVT U5394 ( .A1(\ram[4][153] ), .A2(n5408), .A3(n5409), .A4(data[153]), .Y(n1238) );
  AO22X1_HVT U5395 ( .A1(\ram[4][152] ), .A2(n5408), .A3(n5409), .A4(data[152]), .Y(n1237) );
  AO22X1_HVT U5396 ( .A1(\ram[4][151] ), .A2(n5408), .A3(n5409), .A4(data[151]), .Y(n1236) );
  AO22X1_HVT U5397 ( .A1(\ram[4][150] ), .A2(n5408), .A3(n5409), .A4(data[150]), .Y(n1235) );
  AO22X1_HVT U5398 ( .A1(\ram[4][149] ), .A2(n5408), .A3(n5409), .A4(data[149]), .Y(n1234) );
  AO22X1_HVT U5399 ( .A1(\ram[4][148] ), .A2(n5408), .A3(n5409), .A4(data[148]), .Y(n1233) );
  AO22X1_HVT U5400 ( .A1(\ram[4][147] ), .A2(n5408), .A3(n5409), .A4(data[147]), .Y(n1232) );
  AO22X1_HVT U5401 ( .A1(\ram[4][146] ), .A2(n5408), .A3(n5409), .A4(data[146]), .Y(n1231) );
  AO22X1_HVT U5402 ( .A1(\ram[4][145] ), .A2(n5408), .A3(n5409), .A4(data[145]), .Y(n1230) );
  AO22X1_HVT U5403 ( .A1(\ram[0][62] ), .A2(n5360), .A3(data[62]), .A4(n5361), 
        .Y(n123) );
  AO22X1_HVT U5404 ( .A1(\ram[4][144] ), .A2(n5408), .A3(n5409), .A4(data[144]), .Y(n1229) );
  AO22X1_HVT U5405 ( .A1(\ram[4][143] ), .A2(n5408), .A3(n5409), .A4(data[143]), .Y(n1228) );
  AO22X1_HVT U5406 ( .A1(\ram[4][142] ), .A2(n5408), .A3(n5409), .A4(data[142]), .Y(n1227) );
  AO22X1_HVT U5407 ( .A1(\ram[4][141] ), .A2(n5408), .A3(n5409), .A4(data[141]), .Y(n1226) );
  AO22X1_HVT U5408 ( .A1(\ram[4][140] ), .A2(n5408), .A3(n5409), .A4(data[140]), .Y(n1225) );
  AO22X1_HVT U5409 ( .A1(\ram[4][139] ), .A2(n5408), .A3(n5409), .A4(data[139]), .Y(n1224) );
  AO22X1_HVT U5410 ( .A1(\ram[4][138] ), .A2(n5408), .A3(n5409), .A4(data[138]), .Y(n1223) );
  AO22X1_HVT U5411 ( .A1(\ram[4][137] ), .A2(n5408), .A3(n5409), .A4(data[137]), .Y(n1222) );
  AO22X1_HVT U5412 ( .A1(\ram[4][136] ), .A2(n5408), .A3(n5409), .A4(data[136]), .Y(n1221) );
  AO22X1_HVT U5413 ( .A1(\ram[4][135] ), .A2(n5408), .A3(n5409), .A4(data[135]), .Y(n1220) );
  AO22X1_HVT U5414 ( .A1(\ram[0][61] ), .A2(n5360), .A3(data[61]), .A4(n5361), 
        .Y(n122) );
  AO22X1_HVT U5415 ( .A1(\ram[4][134] ), .A2(n5408), .A3(n5409), .A4(data[134]), .Y(n1219) );
  AO22X1_HVT U5416 ( .A1(\ram[4][133] ), .A2(n5408), .A3(n5409), .A4(data[133]), .Y(n1218) );
  AO22X1_HVT U5417 ( .A1(\ram[4][132] ), .A2(n5408), .A3(n5409), .A4(data[132]), .Y(n1217) );
  AO22X1_HVT U5418 ( .A1(\ram[4][131] ), .A2(n5408), .A3(n5409), .A4(data[131]), .Y(n1216) );
  AO22X1_HVT U5419 ( .A1(\ram[4][130] ), .A2(n5408), .A3(n5409), .A4(data[130]), .Y(n1215) );
  AO22X1_HVT U5420 ( .A1(\ram[4][129] ), .A2(n5408), .A3(n5409), .A4(data[129]), .Y(n1214) );
  AO22X1_HVT U5421 ( .A1(\ram[4][128] ), .A2(n5408), .A3(n5409), .A4(data[128]), .Y(n1213) );
  AO22X1_HVT U5422 ( .A1(\ram[4][127] ), .A2(n5408), .A3(n5409), .A4(data[127]), .Y(n1212) );
  AO22X1_HVT U5423 ( .A1(\ram[4][126] ), .A2(n5408), .A3(n5409), .A4(data[126]), .Y(n1211) );
  AO22X1_HVT U5424 ( .A1(\ram[4][125] ), .A2(n5408), .A3(n5409), .A4(data[125]), .Y(n1210) );
  AO22X1_HVT U5425 ( .A1(\ram[0][60] ), .A2(n5360), .A3(data[60]), .A4(n5361), 
        .Y(n121) );
  AO22X1_HVT U5426 ( .A1(\ram[4][124] ), .A2(n5408), .A3(n5409), .A4(data[124]), .Y(n1209) );
  AO22X1_HVT U5427 ( .A1(\ram[4][123] ), .A2(n5408), .A3(n5409), .A4(data[123]), .Y(n1208) );
  AO22X1_HVT U5428 ( .A1(\ram[4][122] ), .A2(n5408), .A3(n5409), .A4(data[122]), .Y(n1207) );
  AO22X1_HVT U5429 ( .A1(\ram[4][121] ), .A2(n5408), .A3(n5409), .A4(data[121]), .Y(n1206) );
  AO22X1_HVT U5430 ( .A1(\ram[4][120] ), .A2(n5408), .A3(n5409), .A4(data[120]), .Y(n1205) );
  AO22X1_HVT U5431 ( .A1(\ram[4][119] ), .A2(n5408), .A3(n5409), .A4(data[119]), .Y(n1204) );
  AO22X1_HVT U5432 ( .A1(\ram[4][118] ), .A2(n5408), .A3(n5409), .A4(data[118]), .Y(n1203) );
  AO22X1_HVT U5433 ( .A1(\ram[4][117] ), .A2(n5408), .A3(n5409), .A4(data[117]), .Y(n1202) );
  AO22X1_HVT U5434 ( .A1(\ram[4][116] ), .A2(n5408), .A3(n5409), .A4(data[116]), .Y(n1201) );
  AO22X1_HVT U5435 ( .A1(\ram[4][115] ), .A2(n5408), .A3(n5409), .A4(data[115]), .Y(n1200) );
  AO22X1_HVT U5436 ( .A1(\ram[0][59] ), .A2(n5360), .A3(data[59]), .A4(n5361), 
        .Y(n120) );
  AO22X1_HVT U5437 ( .A1(\ram[4][114] ), .A2(n5408), .A3(n5409), .A4(data[114]), .Y(n1199) );
  AO22X1_HVT U5438 ( .A1(\ram[4][113] ), .A2(n5408), .A3(n5409), .A4(data[113]), .Y(n1198) );
  AO22X1_HVT U5439 ( .A1(\ram[4][112] ), .A2(n5408), .A3(n5409), .A4(data[112]), .Y(n1197) );
  AO22X1_HVT U5440 ( .A1(\ram[4][111] ), .A2(n5408), .A3(n5409), .A4(data[111]), .Y(n1196) );
  AO22X1_HVT U5441 ( .A1(\ram[4][110] ), .A2(n5408), .A3(n5409), .A4(data[110]), .Y(n1195) );
  AO22X1_HVT U5442 ( .A1(\ram[4][109] ), .A2(n5408), .A3(n5409), .A4(data[109]), .Y(n1194) );
  AO22X1_HVT U5443 ( .A1(\ram[4][108] ), .A2(n5408), .A3(n5409), .A4(data[108]), .Y(n1193) );
  AO22X1_HVT U5444 ( .A1(\ram[4][107] ), .A2(n5408), .A3(n5409), .A4(data[107]), .Y(n1192) );
  AO22X1_HVT U5445 ( .A1(\ram[4][106] ), .A2(n5408), .A3(n5409), .A4(data[106]), .Y(n1191) );
  AO22X1_HVT U5446 ( .A1(\ram[4][105] ), .A2(n5408), .A3(n5409), .A4(data[105]), .Y(n1190) );
  AO22X1_HVT U5447 ( .A1(\ram[0][58] ), .A2(n5360), .A3(data[58]), .A4(n5361), 
        .Y(n119) );
  AO22X1_HVT U5448 ( .A1(\ram[4][104] ), .A2(n5408), .A3(n5409), .A4(data[104]), .Y(n1189) );
  AO22X1_HVT U5449 ( .A1(\ram[4][103] ), .A2(n5408), .A3(n5409), .A4(data[103]), .Y(n1188) );
  AO22X1_HVT U5450 ( .A1(\ram[4][102] ), .A2(n5408), .A3(n5409), .A4(data[102]), .Y(n1187) );
  AO22X1_HVT U5451 ( .A1(\ram[4][101] ), .A2(n5408), .A3(n5409), .A4(data[101]), .Y(n1186) );
  AO22X1_HVT U5452 ( .A1(\ram[4][100] ), .A2(n5408), .A3(n5409), .A4(data[100]), .Y(n1185) );
  AO22X1_HVT U5453 ( .A1(\ram[4][99] ), .A2(n5408), .A3(n5409), .A4(data[99]), 
        .Y(n1184) );
  AO22X1_HVT U5454 ( .A1(\ram[4][98] ), .A2(n5408), .A3(n5409), .A4(data[98]), 
        .Y(n1183) );
  AO22X1_HVT U5455 ( .A1(\ram[4][97] ), .A2(n5408), .A3(n5409), .A4(data[97]), 
        .Y(n1182) );
  AO22X1_HVT U5456 ( .A1(\ram[4][96] ), .A2(n5408), .A3(n5409), .A4(data[96]), 
        .Y(n1181) );
  AO22X1_HVT U5457 ( .A1(\ram[4][95] ), .A2(n5408), .A3(n5409), .A4(data[95]), 
        .Y(n1180) );
  AO22X1_HVT U5458 ( .A1(\ram[0][57] ), .A2(n5360), .A3(data[57]), .A4(n5361), 
        .Y(n118) );
  AO22X1_HVT U5459 ( .A1(\ram[4][94] ), .A2(n5408), .A3(n5409), .A4(data[94]), 
        .Y(n1179) );
  AO22X1_HVT U5460 ( .A1(\ram[4][93] ), .A2(n5408), .A3(n5409), .A4(data[93]), 
        .Y(n1178) );
  AO22X1_HVT U5461 ( .A1(\ram[4][92] ), .A2(n5408), .A3(n5409), .A4(data[92]), 
        .Y(n1177) );
  AO22X1_HVT U5462 ( .A1(\ram[4][91] ), .A2(n5408), .A3(n5409), .A4(data[91]), 
        .Y(n1176) );
  AO22X1_HVT U5463 ( .A1(\ram[4][90] ), .A2(n5408), .A3(n5409), .A4(data[90]), 
        .Y(n1175) );
  AO22X1_HVT U5464 ( .A1(\ram[4][89] ), .A2(n5408), .A3(n5409), .A4(data[89]), 
        .Y(n1174) );
  AO22X1_HVT U5465 ( .A1(\ram[4][88] ), .A2(n5408), .A3(n5409), .A4(data[88]), 
        .Y(n1173) );
  AO22X1_HVT U5466 ( .A1(\ram[4][87] ), .A2(n5408), .A3(n5409), .A4(data[87]), 
        .Y(n1172) );
  AO22X1_HVT U5467 ( .A1(\ram[4][86] ), .A2(n5408), .A3(n5409), .A4(data[86]), 
        .Y(n1171) );
  AO22X1_HVT U5468 ( .A1(\ram[4][85] ), .A2(n5408), .A3(n5409), .A4(data[85]), 
        .Y(n1170) );
  AO22X1_HVT U5469 ( .A1(\ram[0][56] ), .A2(n5360), .A3(data[56]), .A4(n5361), 
        .Y(n117) );
  AO22X1_HVT U5470 ( .A1(\ram[4][84] ), .A2(n5408), .A3(n5409), .A4(data[84]), 
        .Y(n1169) );
  AO22X1_HVT U5471 ( .A1(\ram[4][83] ), .A2(n5408), .A3(n5409), .A4(data[83]), 
        .Y(n1168) );
  AO22X1_HVT U5472 ( .A1(\ram[4][82] ), .A2(n5408), .A3(n5409), .A4(data[82]), 
        .Y(n1167) );
  AO22X1_HVT U5473 ( .A1(\ram[4][81] ), .A2(n5408), .A3(n5409), .A4(data[81]), 
        .Y(n1166) );
  AO22X1_HVT U5474 ( .A1(\ram[4][80] ), .A2(n5408), .A3(n5409), .A4(data[80]), 
        .Y(n1165) );
  AO22X1_HVT U5475 ( .A1(\ram[4][79] ), .A2(n5408), .A3(n5409), .A4(data[79]), 
        .Y(n1164) );
  AO22X1_HVT U5476 ( .A1(\ram[4][78] ), .A2(n5408), .A3(n5409), .A4(data[78]), 
        .Y(n1163) );
  AO22X1_HVT U5477 ( .A1(\ram[4][77] ), .A2(n5408), .A3(n5409), .A4(data[77]), 
        .Y(n1162) );
  AO22X1_HVT U5478 ( .A1(\ram[4][76] ), .A2(n5408), .A3(n5409), .A4(data[76]), 
        .Y(n1161) );
  AO22X1_HVT U5479 ( .A1(\ram[4][75] ), .A2(n5408), .A3(n5409), .A4(data[75]), 
        .Y(n1160) );
  AO22X1_HVT U5480 ( .A1(\ram[0][55] ), .A2(n5360), .A3(data[55]), .A4(n5361), 
        .Y(n116) );
  AO22X1_HVT U5481 ( .A1(\ram[4][74] ), .A2(n5408), .A3(n5409), .A4(data[74]), 
        .Y(n1159) );
  AO22X1_HVT U5482 ( .A1(\ram[4][73] ), .A2(n5408), .A3(n5409), .A4(data[73]), 
        .Y(n1158) );
  AO22X1_HVT U5483 ( .A1(\ram[4][72] ), .A2(n5408), .A3(n5409), .A4(data[72]), 
        .Y(n1157) );
  AO22X1_HVT U5484 ( .A1(\ram[4][71] ), .A2(n5408), .A3(n5409), .A4(data[71]), 
        .Y(n1156) );
  AO22X1_HVT U5485 ( .A1(\ram[4][70] ), .A2(n5408), .A3(n5409), .A4(data[70]), 
        .Y(n1155) );
  AO22X1_HVT U5486 ( .A1(\ram[4][69] ), .A2(n5408), .A3(n5409), .A4(data[69]), 
        .Y(n1154) );
  AO22X1_HVT U5487 ( .A1(\ram[4][68] ), .A2(n5408), .A3(n5409), .A4(data[68]), 
        .Y(n1153) );
  AO22X1_HVT U5488 ( .A1(\ram[4][67] ), .A2(n5408), .A3(n5409), .A4(data[67]), 
        .Y(n1152) );
  AO22X1_HVT U5489 ( .A1(\ram[4][66] ), .A2(n5408), .A3(n5409), .A4(data[66]), 
        .Y(n1151) );
  AO22X1_HVT U5490 ( .A1(\ram[4][65] ), .A2(n5408), .A3(n5409), .A4(data[65]), 
        .Y(n1150) );
  AO22X1_HVT U5491 ( .A1(\ram[0][54] ), .A2(n5360), .A3(data[54]), .A4(n5361), 
        .Y(n115) );
  AO22X1_HVT U5492 ( .A1(\ram[4][64] ), .A2(n5408), .A3(n5409), .A4(data[64]), 
        .Y(n1149) );
  AO22X1_HVT U5493 ( .A1(\ram[4][63] ), .A2(n5408), .A3(n5409), .A4(data[63]), 
        .Y(n1148) );
  AO22X1_HVT U5494 ( .A1(\ram[4][62] ), .A2(n5408), .A3(n5409), .A4(data[62]), 
        .Y(n1147) );
  AO22X1_HVT U5495 ( .A1(\ram[4][61] ), .A2(n5408), .A3(n5409), .A4(data[61]), 
        .Y(n1146) );
  AO22X1_HVT U5496 ( .A1(\ram[4][60] ), .A2(n5408), .A3(n5409), .A4(data[60]), 
        .Y(n1145) );
  AO22X1_HVT U5497 ( .A1(\ram[4][59] ), .A2(n5408), .A3(n5409), .A4(data[59]), 
        .Y(n1144) );
  AO22X1_HVT U5498 ( .A1(\ram[4][58] ), .A2(n5408), .A3(n5409), .A4(data[58]), 
        .Y(n1143) );
  AO22X1_HVT U5499 ( .A1(\ram[4][57] ), .A2(n5408), .A3(n5409), .A4(data[57]), 
        .Y(n1142) );
  AO22X1_HVT U5500 ( .A1(\ram[4][56] ), .A2(n5408), .A3(n5409), .A4(data[56]), 
        .Y(n1141) );
  AO22X1_HVT U5501 ( .A1(\ram[4][55] ), .A2(n5408), .A3(n5409), .A4(data[55]), 
        .Y(n1140) );
  AO22X1_HVT U5502 ( .A1(\ram[0][53] ), .A2(n5360), .A3(data[53]), .A4(n5361), 
        .Y(n114) );
  AO22X1_HVT U5503 ( .A1(\ram[4][54] ), .A2(n5408), .A3(n5409), .A4(data[54]), 
        .Y(n1139) );
  AO22X1_HVT U5504 ( .A1(\ram[4][53] ), .A2(n5408), .A3(n5409), .A4(data[53]), 
        .Y(n1138) );
  AO22X1_HVT U5505 ( .A1(\ram[4][52] ), .A2(n5408), .A3(n5409), .A4(data[52]), 
        .Y(n1137) );
  AO22X1_HVT U5506 ( .A1(\ram[4][51] ), .A2(n5408), .A3(n5409), .A4(data[51]), 
        .Y(n1136) );
  AO22X1_HVT U5507 ( .A1(\ram[4][50] ), .A2(n5408), .A3(n5409), .A4(data[50]), 
        .Y(n1135) );
  AO22X1_HVT U5508 ( .A1(\ram[4][49] ), .A2(n5408), .A3(n5409), .A4(data[49]), 
        .Y(n1134) );
  AO22X1_HVT U5509 ( .A1(\ram[4][48] ), .A2(n5408), .A3(n5409), .A4(data[48]), 
        .Y(n1133) );
  AO22X1_HVT U5510 ( .A1(\ram[4][47] ), .A2(n5408), .A3(n5409), .A4(data[47]), 
        .Y(n1132) );
  AO22X1_HVT U5511 ( .A1(\ram[4][46] ), .A2(n5408), .A3(n5409), .A4(data[46]), 
        .Y(n1131) );
  AO22X1_HVT U5512 ( .A1(\ram[4][45] ), .A2(n5408), .A3(n5409), .A4(data[45]), 
        .Y(n1130) );
  AO22X1_HVT U5513 ( .A1(\ram[0][52] ), .A2(n5360), .A3(data[52]), .A4(n5361), 
        .Y(n113) );
  AO22X1_HVT U5514 ( .A1(\ram[4][44] ), .A2(n5408), .A3(n5409), .A4(data[44]), 
        .Y(n1129) );
  AO22X1_HVT U5515 ( .A1(\ram[4][43] ), .A2(n5408), .A3(n5409), .A4(data[43]), 
        .Y(n1128) );
  AO22X1_HVT U5516 ( .A1(\ram[4][42] ), .A2(n5408), .A3(n5409), .A4(data[42]), 
        .Y(n1127) );
  AO22X1_HVT U5517 ( .A1(\ram[4][41] ), .A2(n5408), .A3(n5409), .A4(data[41]), 
        .Y(n1126) );
  AO22X1_HVT U5518 ( .A1(\ram[4][40] ), .A2(n5408), .A3(n5409), .A4(data[40]), 
        .Y(n1125) );
  AO22X1_HVT U5519 ( .A1(\ram[4][39] ), .A2(n5408), .A3(n5409), .A4(data[39]), 
        .Y(n1124) );
  AO22X1_HVT U5520 ( .A1(\ram[4][38] ), .A2(n5408), .A3(n5409), .A4(data[38]), 
        .Y(n1123) );
  AO22X1_HVT U5521 ( .A1(\ram[4][37] ), .A2(n5408), .A3(n5409), .A4(data[37]), 
        .Y(n1122) );
  AO22X1_HVT U5522 ( .A1(\ram[4][36] ), .A2(n5408), .A3(n5409), .A4(data[36]), 
        .Y(n1121) );
  AO22X1_HVT U5523 ( .A1(\ram[4][35] ), .A2(n5408), .A3(n5409), .A4(data[35]), 
        .Y(n1120) );
  AO22X1_HVT U5524 ( .A1(\ram[0][51] ), .A2(n5360), .A3(data[51]), .A4(n5361), 
        .Y(n112) );
  AO22X1_HVT U5525 ( .A1(\ram[4][34] ), .A2(n5408), .A3(n5409), .A4(data[34]), 
        .Y(n1119) );
  AO22X1_HVT U5526 ( .A1(\ram[4][33] ), .A2(n5408), .A3(n5409), .A4(data[33]), 
        .Y(n1118) );
  AO22X1_HVT U5527 ( .A1(\ram[4][32] ), .A2(n5408), .A3(n5409), .A4(data[32]), 
        .Y(n1117) );
  AO22X1_HVT U5528 ( .A1(\ram[4][31] ), .A2(n5408), .A3(n5409), .A4(data[31]), 
        .Y(n1116) );
  AO22X1_HVT U5529 ( .A1(\ram[4][30] ), .A2(n5408), .A3(n5409), .A4(data[30]), 
        .Y(n1115) );
  AO22X1_HVT U5530 ( .A1(\ram[4][29] ), .A2(n5408), .A3(n5409), .A4(data[29]), 
        .Y(n1114) );
  AO22X1_HVT U5531 ( .A1(\ram[4][28] ), .A2(n5408), .A3(n5409), .A4(data[28]), 
        .Y(n1113) );
  AO22X1_HVT U5532 ( .A1(\ram[4][27] ), .A2(n5408), .A3(n5409), .A4(data[27]), 
        .Y(n1112) );
  AO22X1_HVT U5533 ( .A1(\ram[4][26] ), .A2(n5408), .A3(n5409), .A4(data[26]), 
        .Y(n1111) );
  AO22X1_HVT U5534 ( .A1(\ram[4][25] ), .A2(n5408), .A3(n5409), .A4(data[25]), 
        .Y(n1110) );
  AO22X1_HVT U5535 ( .A1(\ram[0][50] ), .A2(n5360), .A3(data[50]), .A4(n5361), 
        .Y(n111) );
  AO22X1_HVT U5536 ( .A1(\ram[4][24] ), .A2(n5408), .A3(n5409), .A4(data[24]), 
        .Y(n1109) );
  AO22X1_HVT U5537 ( .A1(\ram[4][23] ), .A2(n5408), .A3(n5409), .A4(data[23]), 
        .Y(n1108) );
  AO22X1_HVT U5538 ( .A1(\ram[4][22] ), .A2(n5408), .A3(n5409), .A4(data[22]), 
        .Y(n1107) );
  AO22X1_HVT U5539 ( .A1(\ram[4][21] ), .A2(n5408), .A3(n5409), .A4(data[21]), 
        .Y(n1106) );
  AO22X1_HVT U5540 ( .A1(\ram[4][20] ), .A2(n5408), .A3(n5409), .A4(data[20]), 
        .Y(n1105) );
  AO22X1_HVT U5541 ( .A1(\ram[4][19] ), .A2(n5408), .A3(n5409), .A4(data[19]), 
        .Y(n1104) );
  AO22X1_HVT U5542 ( .A1(\ram[4][18] ), .A2(n5408), .A3(n5409), .A4(data[18]), 
        .Y(n1103) );
  AO22X1_HVT U5543 ( .A1(\ram[4][17] ), .A2(n5408), .A3(n5409), .A4(data[17]), 
        .Y(n1102) );
  AO22X1_HVT U5544 ( .A1(\ram[4][16] ), .A2(n5408), .A3(n5409), .A4(data[16]), 
        .Y(n1101) );
  AO22X1_HVT U5545 ( .A1(\ram[4][15] ), .A2(n5408), .A3(n5409), .A4(data[15]), 
        .Y(n1100) );
  AO22X1_HVT U5546 ( .A1(\ram[0][49] ), .A2(n5360), .A3(data[49]), .A4(n5361), 
        .Y(n110) );
  AO22X1_HVT U5547 ( .A1(\ram[4][14] ), .A2(n5408), .A3(n5409), .A4(data[14]), 
        .Y(n1099) );
  AO22X1_HVT U5548 ( .A1(\ram[4][13] ), .A2(n5408), .A3(n5409), .A4(data[13]), 
        .Y(n1098) );
  AO22X1_HVT U5549 ( .A1(\ram[4][12] ), .A2(n5408), .A3(n5409), .A4(data[12]), 
        .Y(n1097) );
  AO22X1_HVT U5550 ( .A1(\ram[4][11] ), .A2(n5408), .A3(n5409), .A4(data[11]), 
        .Y(n1096) );
  AO22X1_HVT U5551 ( .A1(\ram[4][10] ), .A2(n5408), .A3(n5409), .A4(data[10]), 
        .Y(n1095) );
  AO22X1_HVT U5552 ( .A1(\ram[4][9] ), .A2(n5408), .A3(n5409), .A4(data[9]), 
        .Y(n1094) );
  AO22X1_HVT U5553 ( .A1(\ram[4][8] ), .A2(n5408), .A3(n5409), .A4(data[8]), 
        .Y(n1093) );
  AO22X1_HVT U5554 ( .A1(\ram[4][7] ), .A2(n5408), .A3(n5409), .A4(data[7]), 
        .Y(n1092) );
  AO22X1_HVT U5555 ( .A1(\ram[4][6] ), .A2(n5408), .A3(n5409), .A4(data[6]), 
        .Y(n1091) );
  AO22X1_HVT U5556 ( .A1(\ram[4][5] ), .A2(n5408), .A3(n5409), .A4(data[5]), 
        .Y(n1090) );
  AO22X1_HVT U5557 ( .A1(\ram[0][48] ), .A2(n5360), .A3(data[48]), .A4(n5361), 
        .Y(n109) );
  AO22X1_HVT U5558 ( .A1(\ram[4][4] ), .A2(n5408), .A3(n5409), .A4(data[4]), 
        .Y(n1089) );
  AO22X1_HVT U5559 ( .A1(\ram[4][3] ), .A2(n5408), .A3(n5409), .A4(data[3]), 
        .Y(n1088) );
  AO22X1_HVT U5560 ( .A1(\ram[4][2] ), .A2(n5408), .A3(n5409), .A4(data[2]), 
        .Y(n1087) );
  AO22X1_HVT U5561 ( .A1(\ram[4][1] ), .A2(n5408), .A3(n5409), .A4(data[1]), 
        .Y(n1086) );
  AO22X1_HVT U5562 ( .A1(\ram[4][0] ), .A2(n5408), .A3(n5409), .A4(data[0]), 
        .Y(n1085) );
  INVX0_HVT U5563 ( .A(n5410), .Y(n5409) );
  AND2X1_HVT U5564 ( .A1(n5410), .A2(n5365), .Y(n5408) );
  NAND3X0_HVT U5565 ( .A1(n4183), .A2(n4280), .A3(n5401), .Y(n5410) );
  AND2X1_HVT U5566 ( .A1(N28), .A2(n5367), .Y(n5401) );
  AO22X1_HVT U5567 ( .A1(\ram[3][255] ), .A2(n5358), .A3(data[255]), .A4(n5359), .Y(n1084) );
  AO22X1_HVT U5568 ( .A1(\ram[3][254] ), .A2(n5358), .A3(data[254]), .A4(n5359), .Y(n1083) );
  AO22X1_HVT U5569 ( .A1(\ram[3][253] ), .A2(n5358), .A3(data[253]), .A4(n5359), .Y(n1082) );
  AO22X1_HVT U5570 ( .A1(\ram[3][252] ), .A2(n5358), .A3(data[252]), .A4(n5359), .Y(n1081) );
  AO22X1_HVT U5571 ( .A1(\ram[3][251] ), .A2(n5358), .A3(data[251]), .A4(n5359), .Y(n1080) );
  AO22X1_HVT U5572 ( .A1(\ram[0][47] ), .A2(n5360), .A3(data[47]), .A4(n5361), 
        .Y(n108) );
  AO22X1_HVT U5573 ( .A1(\ram[3][250] ), .A2(n5358), .A3(data[250]), .A4(n5359), .Y(n1079) );
  AO22X1_HVT U5574 ( .A1(\ram[3][249] ), .A2(n5358), .A3(data[249]), .A4(n5359), .Y(n1078) );
  AO22X1_HVT U5575 ( .A1(\ram[3][248] ), .A2(n5358), .A3(data[248]), .A4(n5359), .Y(n1077) );
  AO22X1_HVT U5576 ( .A1(\ram[3][247] ), .A2(n5358), .A3(data[247]), .A4(n5359), .Y(n1076) );
  AO22X1_HVT U5577 ( .A1(\ram[3][246] ), .A2(n5358), .A3(data[246]), .A4(n5359), .Y(n1075) );
  AO22X1_HVT U5578 ( .A1(\ram[3][245] ), .A2(n5358), .A3(data[245]), .A4(n5359), .Y(n1074) );
  AO22X1_HVT U5579 ( .A1(\ram[3][244] ), .A2(n5358), .A3(data[244]), .A4(n5359), .Y(n1073) );
  AO22X1_HVT U5580 ( .A1(\ram[3][243] ), .A2(n5358), .A3(data[243]), .A4(n5359), .Y(n1072) );
  AO22X1_HVT U5581 ( .A1(\ram[3][242] ), .A2(n5358), .A3(data[242]), .A4(n5359), .Y(n1071) );
  AO22X1_HVT U5582 ( .A1(\ram[3][241] ), .A2(n5358), .A3(data[241]), .A4(n5359), .Y(n1070) );
  AO22X1_HVT U5583 ( .A1(\ram[0][46] ), .A2(n5360), .A3(data[46]), .A4(n5361), 
        .Y(n107) );
  AO22X1_HVT U5584 ( .A1(\ram[3][240] ), .A2(n5358), .A3(data[240]), .A4(n5359), .Y(n1069) );
  AO22X1_HVT U5585 ( .A1(\ram[3][239] ), .A2(n5358), .A3(data[239]), .A4(n5359), .Y(n1068) );
  AO22X1_HVT U5586 ( .A1(\ram[3][238] ), .A2(n5358), .A3(data[238]), .A4(n5359), .Y(n1067) );
  AO22X1_HVT U5587 ( .A1(\ram[3][237] ), .A2(n5358), .A3(data[237]), .A4(n5359), .Y(n1066) );
  AO22X1_HVT U5588 ( .A1(\ram[3][236] ), .A2(n5358), .A3(data[236]), .A4(n5359), .Y(n1065) );
  AO22X1_HVT U5589 ( .A1(\ram[3][235] ), .A2(n5358), .A3(data[235]), .A4(n5359), .Y(n1064) );
  AO22X1_HVT U5590 ( .A1(\ram[3][234] ), .A2(n5358), .A3(data[234]), .A4(n5359), .Y(n1063) );
  AO22X1_HVT U5591 ( .A1(\ram[3][233] ), .A2(n5358), .A3(data[233]), .A4(n5359), .Y(n1062) );
  AO22X1_HVT U5592 ( .A1(\ram[3][232] ), .A2(n5358), .A3(data[232]), .A4(n5359), .Y(n1061) );
  AO22X1_HVT U5593 ( .A1(\ram[3][231] ), .A2(n5358), .A3(data[231]), .A4(n5359), .Y(n1060) );
  AO22X1_HVT U5594 ( .A1(\ram[0][45] ), .A2(n5360), .A3(data[45]), .A4(n5361), 
        .Y(n106) );
  AO22X1_HVT U5595 ( .A1(\ram[3][230] ), .A2(n5358), .A3(data[230]), .A4(n5359), .Y(n1059) );
  AO22X1_HVT U5596 ( .A1(\ram[3][229] ), .A2(n5358), .A3(data[229]), .A4(n5359), .Y(n1058) );
  AO22X1_HVT U5597 ( .A1(\ram[3][228] ), .A2(n5358), .A3(data[228]), .A4(n5359), .Y(n1057) );
  AO22X1_HVT U5598 ( .A1(\ram[3][227] ), .A2(n5358), .A3(data[227]), .A4(n5359), .Y(n1056) );
  AO22X1_HVT U5599 ( .A1(\ram[3][226] ), .A2(n5358), .A3(data[226]), .A4(n5359), .Y(n1055) );
  AO22X1_HVT U5600 ( .A1(\ram[3][225] ), .A2(n5358), .A3(data[225]), .A4(n5359), .Y(n1054) );
  AO22X1_HVT U5601 ( .A1(\ram[3][224] ), .A2(n5358), .A3(data[224]), .A4(n5359), .Y(n1053) );
  AO22X1_HVT U5602 ( .A1(\ram[3][223] ), .A2(n5358), .A3(data[223]), .A4(n5359), .Y(n1052) );
  AO22X1_HVT U5603 ( .A1(\ram[3][222] ), .A2(n5358), .A3(data[222]), .A4(n5359), .Y(n1051) );
  AO22X1_HVT U5604 ( .A1(\ram[3][221] ), .A2(n5358), .A3(data[221]), .A4(n5359), .Y(n1050) );
  AO22X1_HVT U5605 ( .A1(\ram[0][44] ), .A2(n5360), .A3(data[44]), .A4(n5361), 
        .Y(n105) );
  AO22X1_HVT U5606 ( .A1(\ram[3][220] ), .A2(n5358), .A3(data[220]), .A4(n5359), .Y(n1049) );
  AO22X1_HVT U5607 ( .A1(\ram[3][219] ), .A2(n5358), .A3(data[219]), .A4(n5359), .Y(n1048) );
  AO22X1_HVT U5608 ( .A1(\ram[3][218] ), .A2(n5358), .A3(data[218]), .A4(n5359), .Y(n1047) );
  AO22X1_HVT U5609 ( .A1(\ram[3][217] ), .A2(n5358), .A3(data[217]), .A4(n5359), .Y(n1046) );
  AO22X1_HVT U5610 ( .A1(\ram[3][216] ), .A2(n5358), .A3(data[216]), .A4(n5359), .Y(n1045) );
  AO22X1_HVT U5611 ( .A1(\ram[3][215] ), .A2(n5358), .A3(data[215]), .A4(n5359), .Y(n1044) );
  AO22X1_HVT U5612 ( .A1(\ram[3][214] ), .A2(n5358), .A3(data[214]), .A4(n5359), .Y(n1043) );
  AO22X1_HVT U5613 ( .A1(\ram[3][213] ), .A2(n5358), .A3(data[213]), .A4(n5359), .Y(n1042) );
  AO22X1_HVT U5614 ( .A1(\ram[3][212] ), .A2(n5358), .A3(data[212]), .A4(n5359), .Y(n1041) );
  AO22X1_HVT U5615 ( .A1(\ram[3][211] ), .A2(n5358), .A3(data[211]), .A4(n5359), .Y(n1040) );
  AO22X1_HVT U5616 ( .A1(\ram[0][43] ), .A2(n5360), .A3(data[43]), .A4(n5361), 
        .Y(n104) );
  AO22X1_HVT U5617 ( .A1(\ram[3][210] ), .A2(n5358), .A3(data[210]), .A4(n5359), .Y(n1039) );
  AO22X1_HVT U5618 ( .A1(\ram[3][209] ), .A2(n5358), .A3(data[209]), .A4(n5359), .Y(n1038) );
  AO22X1_HVT U5619 ( .A1(\ram[3][208] ), .A2(n5358), .A3(data[208]), .A4(n5359), .Y(n1037) );
  AO22X1_HVT U5620 ( .A1(\ram[3][207] ), .A2(n5358), .A3(data[207]), .A4(n5359), .Y(n1036) );
  AO22X1_HVT U5621 ( .A1(\ram[3][206] ), .A2(n5358), .A3(data[206]), .A4(n5359), .Y(n1035) );
  AO22X1_HVT U5622 ( .A1(\ram[3][205] ), .A2(n5358), .A3(data[205]), .A4(n5359), .Y(n1034) );
  AO22X1_HVT U5623 ( .A1(\ram[3][204] ), .A2(n5358), .A3(data[204]), .A4(n5359), .Y(n1033) );
  AO22X1_HVT U5624 ( .A1(\ram[3][203] ), .A2(n5358), .A3(data[203]), .A4(n5359), .Y(n1032) );
  AO22X1_HVT U5625 ( .A1(\ram[3][202] ), .A2(n5358), .A3(data[202]), .A4(n5359), .Y(n1031) );
  AO22X1_HVT U5626 ( .A1(\ram[3][201] ), .A2(n5358), .A3(data[201]), .A4(n5359), .Y(n1030) );
  AO22X1_HVT U5627 ( .A1(\ram[0][42] ), .A2(n5360), .A3(data[42]), .A4(n5361), 
        .Y(n103) );
  AO22X1_HVT U5628 ( .A1(\ram[3][200] ), .A2(n5358), .A3(data[200]), .A4(n5359), .Y(n1029) );
  AO22X1_HVT U5629 ( .A1(\ram[3][199] ), .A2(n5358), .A3(data[199]), .A4(n5359), .Y(n1028) );
  AO22X1_HVT U5630 ( .A1(\ram[3][198] ), .A2(n5358), .A3(data[198]), .A4(n5359), .Y(n1027) );
  AO22X1_HVT U5631 ( .A1(\ram[3][197] ), .A2(n5358), .A3(data[197]), .A4(n5359), .Y(n1026) );
  AO22X1_HVT U5632 ( .A1(\ram[3][196] ), .A2(n5358), .A3(data[196]), .A4(n5359), .Y(n1025) );
  AO22X1_HVT U5633 ( .A1(\ram[3][195] ), .A2(n5358), .A3(data[195]), .A4(n5359), .Y(n1024) );
  AO22X1_HVT U5634 ( .A1(\ram[3][194] ), .A2(n5358), .A3(data[194]), .A4(n5359), .Y(n1023) );
  AO22X1_HVT U5635 ( .A1(\ram[3][193] ), .A2(n5358), .A3(data[193]), .A4(n5359), .Y(n1022) );
  AO22X1_HVT U5636 ( .A1(\ram[3][192] ), .A2(n5358), .A3(data[192]), .A4(n5359), .Y(n1021) );
  AO22X1_HVT U5637 ( .A1(\ram[3][191] ), .A2(n5358), .A3(data[191]), .A4(n5359), .Y(n1020) );
  AO22X1_HVT U5638 ( .A1(\ram[0][41] ), .A2(n5360), .A3(data[41]), .A4(n5361), 
        .Y(n102) );
  AO22X1_HVT U5639 ( .A1(\ram[3][190] ), .A2(n5358), .A3(data[190]), .A4(n5359), .Y(n1019) );
  AO22X1_HVT U5640 ( .A1(\ram[3][189] ), .A2(n5358), .A3(data[189]), .A4(n5359), .Y(n1018) );
  AO22X1_HVT U5641 ( .A1(\ram[3][188] ), .A2(n5358), .A3(data[188]), .A4(n5359), .Y(n1017) );
  AO22X1_HVT U5642 ( .A1(\ram[3][187] ), .A2(n5358), .A3(data[187]), .A4(n5359), .Y(n1016) );
  AO22X1_HVT U5643 ( .A1(\ram[3][186] ), .A2(n5358), .A3(data[186]), .A4(n5359), .Y(n1015) );
  AO22X1_HVT U5644 ( .A1(\ram[3][185] ), .A2(n5358), .A3(data[185]), .A4(n5359), .Y(n1014) );
  AO22X1_HVT U5645 ( .A1(\ram[3][184] ), .A2(n5358), .A3(data[184]), .A4(n5359), .Y(n1013) );
  AO22X1_HVT U5646 ( .A1(\ram[3][183] ), .A2(n5358), .A3(data[183]), .A4(n5359), .Y(n1012) );
  AO22X1_HVT U5647 ( .A1(\ram[3][182] ), .A2(n5358), .A3(data[182]), .A4(n5359), .Y(n1011) );
  AO22X1_HVT U5648 ( .A1(\ram[3][181] ), .A2(n5358), .A3(data[181]), .A4(n5359), .Y(n1010) );
  AO22X1_HVT U5649 ( .A1(\ram[0][40] ), .A2(n5360), .A3(data[40]), .A4(n5361), 
        .Y(n101) );
  AO22X1_HVT U5650 ( .A1(\ram[3][180] ), .A2(n5358), .A3(data[180]), .A4(n5359), .Y(n1009) );
  AO22X1_HVT U5651 ( .A1(\ram[3][179] ), .A2(n5358), .A3(data[179]), .A4(n5359), .Y(n1008) );
  AO22X1_HVT U5652 ( .A1(\ram[3][178] ), .A2(n5358), .A3(data[178]), .A4(n5359), .Y(n1007) );
  AO22X1_HVT U5653 ( .A1(\ram[3][177] ), .A2(n5358), .A3(data[177]), .A4(n5359), .Y(n1006) );
  AO22X1_HVT U5654 ( .A1(\ram[3][176] ), .A2(n5358), .A3(data[176]), .A4(n5359), .Y(n1005) );
  AO22X1_HVT U5655 ( .A1(\ram[3][175] ), .A2(n5358), .A3(data[175]), .A4(n5359), .Y(n1004) );
  AO22X1_HVT U5656 ( .A1(\ram[3][174] ), .A2(n5358), .A3(data[174]), .A4(n5359), .Y(n1003) );
  AO22X1_HVT U5657 ( .A1(\ram[3][173] ), .A2(n5358), .A3(data[173]), .A4(n5359), .Y(n1002) );
  AO22X1_HVT U5658 ( .A1(\ram[3][172] ), .A2(n5358), .A3(data[172]), .A4(n5359), .Y(n1001) );
  AO22X1_HVT U5659 ( .A1(\ram[3][171] ), .A2(n5358), .A3(data[171]), .A4(n5359), .Y(n1000) );
  INVX0_HVT U5660 ( .A(n5411), .Y(n5359) );
  AND2X1_HVT U5661 ( .A1(n5411), .A2(n5365), .Y(n5358) );
  NAND3X0_HVT U5662 ( .A1(n5367), .A2(n5366), .A3(n4182), .Y(n5411) );
  AND2X1_HVT U5663 ( .A1(n4276), .A2(n4308), .Y(n5366) );
  AO22X1_HVT U5664 ( .A1(\ram[0][39] ), .A2(n5360), .A3(data[39]), .A4(n5361), 
        .Y(n100) );
  INVX0_HVT U5665 ( .A(n5412), .Y(n5361) );
  AND2X1_HVT U5666 ( .A1(n5412), .A2(n5365), .Y(n5360) );
  INVX0_HVT U5667 ( .A(rst), .Y(n5365) );
  NAND3X0_HVT U5668 ( .A1(n5367), .A2(n4183), .A3(n5383), .Y(n5412) );
  AND2X1_HVT U5669 ( .A1(n4277), .A2(n4308), .Y(n5383) );
  AND2X1_HVT U5670 ( .A1(we), .A2(n4331), .Y(n5367) );
endmodule

