
module sbox_5 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n3, n19, n23, n34, n35, n38, n50, n82, n118, n119, n147, n148, n210,
         n211, n212, n213, n216, n217, n218, n219, n220, n227, n230, n231,
         n232, n236, n238, n241, n252, n254, n255, n257, n261, n264, n266,
         n269, n272, n273, n275, n279, n280, n282, n283, n284, n285, n289,
         n290, n292, n293, n294, n297, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771;

  NAND2X0_HVT U4 ( .A1(n400), .A2(n429), .Y(n769) );
  NAND2X0_HVT U5 ( .A1(n511), .A2(n504), .Y(n767) );
  NAND2X0_HVT U13 ( .A1(n759), .A2(n319), .Y(n760) );
  NAND2X0_HVT U15 ( .A1(n429), .A2(n473), .Y(n757) );
  NAND2X0_HVT U21 ( .A1(n400), .A2(n326), .Y(n752) );
  NAND2X0_HVT U24 ( .A1(n406), .A2(n355), .Y(n750) );
  NAND2X0_HVT U35 ( .A1(n501), .A2(n326), .Y(n741) );
  NAND2X0_HVT U42 ( .A1(n272), .A2(n500), .Y(n735) );
  NAND2X0_HVT U53 ( .A1(n724), .A2(n734), .Y(n725) );
  NAND2X0_HVT U56 ( .A1(n400), .A2(n720), .Y(n721) );
  MUX41X1_HVT U57 ( .A1(n534), .A3(n754), .A2(n721), .A4(n762), .S0(n517), 
        .S1(n494), .Y(n719) );
  NAND2X0_HVT U58 ( .A1(n319), .A2(n232), .Y(n718) );
  MUX41X1_HVT U59 ( .A1(n483), .A3(n718), .A2(n482), .A4(n410), .S0(n254), 
        .S1(n494), .Y(n717) );
  MUX41X1_HVT U61 ( .A1(n480), .A3(n551), .A2(n352), .A4(n473), .S0(n518), 
        .S1(n494), .Y(n715) );
  NAND2X0_HVT U62 ( .A1(n355), .A2(n461), .Y(n714) );
  MUX41X1_HVT U63 ( .A1(n714), .A3(n529), .A2(n418), .A4(n407), .S0(n519), 
        .S1(n494), .Y(n713) );
  AO21X1_HVT U66 ( .A1(n558), .A2(n493), .A3(n560), .Y(n710) );
  MUX41X1_HVT U69 ( .A1(n708), .A3(n716), .A2(n712), .A4(n722), .S0(n327), 
        .S1(n499), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n241), .A2(n703), .Y(n704) );
  MUX41X1_HVT U74 ( .A1(n705), .A3(n748), .A2(n704), .A4(n750), .S0(n210), 
        .S1(n517), .Y(n702) );
  AND2X1_HVT U83 ( .A1(n388), .A2(n453), .Y(n693) );
  MUX41X1_HVT U84 ( .A1(n356), .A3(n283), .A2(n756), .A4(n693), .S0(n488), 
        .S1(n332), .Y(n692) );
  NAND2X0_HVT U85 ( .A1(n326), .A2(n559), .Y(n691) );
  MUX41X1_HVT U90 ( .A1(n731), .A3(n735), .A2(n218), .A4(n688), .S0(n489), 
        .S1(n332), .Y(n687) );
  MUX41X1_HVT U97 ( .A1(n556), .A3(n479), .A2(n511), .A4(n757), .S0(n488), 
        .S1(n332), .Y(n679) );
  NAND2X0_HVT U101 ( .A1(n674), .A2(n673), .Y(n675) );
  MUX41X1_HVT U103 ( .A1(n429), .A3(n546), .A2(n452), .A4(n741), .S0(n488), 
        .S1(n518), .Y(n671) );
  MUX41X1_HVT U105 ( .A1(n550), .A3(n729), .A2(n670), .A4(n543), .S0(n488), 
        .S1(n518), .Y(n669) );
  NAND2X0_HVT U110 ( .A1(n460), .A2(n664), .Y(n665) );
  AND2X1_HVT U115 ( .A1(n511), .A2(n357), .Y(n661) );
  NAND2X0_HVT U123 ( .A1(n651), .A2(n652), .Y(n653) );
  MUX41X1_HVT U125 ( .A1(n752), .A3(n483), .A2(n531), .A4(n540), .S0(n489), 
        .S1(n519), .Y(n649) );
  AND2X1_HVT U154 ( .A1(n496), .A2(n500), .Y(n624) );
  NAND2X0_HVT U158 ( .A1(n344), .A2(n315), .Y(n620) );
  MUX41X1_HVT U159 ( .A1(n341), .A3(n471), .A2(n620), .A4(n561), .S0(n395), 
        .S1(n465), .Y(n619) );
  AND2X1_HVT U162 ( .A1(n366), .A2(n330), .Y(n616) );
  MUX41X1_HVT U165 ( .A1(n752), .A3(n549), .A2(n731), .A4(n614), .S0(n518), 
        .S1(n485), .Y(n613) );
  NAND2X0_HVT U166 ( .A1(n319), .A2(n720), .Y(n612) );
  NAND2X0_HVT U167 ( .A1(n464), .A2(n326), .Y(n611) );
  MUX41X1_HVT U168 ( .A1(n534), .A3(n257), .A2(n611), .A4(n612), .S0(n491), 
        .S1(n519), .Y(n610) );
  NAND2X0_HVT U174 ( .A1(n510), .A2(n470), .Y(n759) );
  NAND2X0_HVT U177 ( .A1(n511), .A2(n501), .Y(n603) );
  MUX41X1_HVT U179 ( .A1(n746), .A3(n3), .A2(n535), .A4(n548), .S0(n395), .S1(
        n332), .Y(n601) );
  MUX41X1_HVT U182 ( .A1(n539), .A3(n399), .A2(n363), .A4(n440), .S0(n519), 
        .S1(n485), .Y(n598) );
  AO21X1_HVT U197 ( .A1(n481), .A2(n498), .A3(n552), .Y(n584) );
  MUX41X1_HVT U204 ( .A1(n721), .A3(n760), .A2(n405), .A4(n751), .S0(n210), 
        .S1(n466), .Y(n577) );
  NAND2X0_HVT U208 ( .A1(n509), .A2(n289), .Y(n664) );
  NAND2X0_HVT U214 ( .A1(n283), .A2(n428), .Y(n574) );
  NAND2X0_HVT U215 ( .A1(n664), .A2(n257), .Y(n573) );
  NAND2X0_HVT U218 ( .A1(n255), .A2(n358), .Y(n627) );
  NAND2X0_HVT U220 ( .A1(n497), .A2(n574), .Y(n696) );
  INVX0_HVT U241 ( .A(n750), .Y(n564) );
  INVX0_HVT U242 ( .A(n735), .Y(n563) );
  INVX0_HVT U245 ( .A(n767), .Y(n561) );
  INVX0_HVT U256 ( .A(n627), .Y(n552) );
  INVX0_HVT U268 ( .A(n752), .Y(n544) );
  INVX0_HVT U270 ( .A(n573), .Y(n543) );
  INVX0_HVT U284 ( .A(n574), .Y(n535) );
  INVX0_HVT U289 ( .A(n673), .Y(n532) );
  INVX0_HVT U295 ( .A(n769), .Y(n530) );
  INVX0_HVT U296 ( .A(n757), .Y(n529) );
  INVX0_HVT U306 ( .A(n611), .Y(n525) );
  INVX0_HVT U309 ( .A(n754), .Y(n522) );
  MUX21X1_HVT U1 ( .A1(n453), .A2(n554), .S0(n451), .Y(n755) );
  OA21X1_HVT U2 ( .A1(n261), .A2(n324), .A3(n356), .Y(n596) );
  INVX1_HVT U3 ( .A(n316), .Y(n318) );
  INVX0_HVT U6 ( .A(n502), .Y(n441) );
  AND3X1_HVT U7 ( .A1(n491), .A2(n428), .A3(n453), .Y(n646) );
  MUX21X1_HVT U8 ( .A1(n628), .A2(n629), .S0(n492), .Y(n626) );
  INVX1_HVT U9 ( .A(n514), .Y(n484) );
  AND2X1_HVT U10 ( .A1(n231), .A2(n365), .Y(n3) );
  INVX1_HVT U11 ( .A(n499), .Y(n118) );
  AND2X1_HVT U12 ( .A1(n241), .A2(n355), .Y(n19) );
  IBUFFX2_HVT U14 ( .A(n720), .Y(n556) );
  INVX0_HVT U16 ( .A(n506), .Y(n526) );
  AND2X1_HVT U17 ( .A1(n371), .A2(n370), .Y(n23) );
  MUX41X1_HVT U18 ( .A1(n524), .A3(n742), .A2(n740), .A4(n761), .S0(n465), 
        .S1(n459), .Y(n578) );
  INVX0_HVT U19 ( .A(n376), .Y(n377) );
  INVX0_HVT U20 ( .A(n375), .Y(n359) );
  INVX1_HVT U22 ( .A(n374), .Y(n358) );
  INVX1_HVT U23 ( .A(n486), .Y(n460) );
  MUX41X1_HVT U25 ( .A1(n533), .A3(n700), .A2(n541), .A4(n764), .S0(n474), 
        .S1(n484), .Y(n699) );
  INVX1_HVT U26 ( .A(n360), .Y(n34) );
  INVX1_HVT U27 ( .A(n34), .Y(n35) );
  INVX0_HVT U28 ( .A(n771), .Y(n316) );
  INVX0_HVT U29 ( .A(n562), .Y(n406) );
  INVX1_HVT U30 ( .A(n380), .Y(n468) );
  MUX21X1_HVT U31 ( .A1(n501), .A2(n473), .S0(n428), .Y(n673) );
  MUX41X1_HVT U32 ( .A1(n501), .A3(n605), .A2(n532), .A4(n342), .S0(n517), 
        .S1(n485), .Y(n604) );
  OR2X1_HVT U33 ( .A1(n119), .A2(n38), .Y(n348) );
  NAND2X0_HVT U34 ( .A1(n453), .A2(n38), .Y(n50) );
  NAND2X0_HVT U36 ( .A1(n398), .A2(n386), .Y(n82) );
  NAND2X0_HVT U37 ( .A1(n50), .A2(n82), .Y(n742) );
  INVX0_HVT U38 ( .A(n386), .Y(n38) );
  INVX1_HVT U39 ( .A(n502), .Y(n453) );
  MUX41X1_HVT U40 ( .A1(n553), .A3(n556), .A2(n523), .A4(n463), .S0(n484), 
        .S1(n332), .Y(n701) );
  INVX1_HVT U41 ( .A(n749), .Y(n523) );
  MUX41X1_HVT U43 ( .A1(n625), .A3(n619), .A2(n626), .A4(n621), .S0(n118), 
        .S1(n495), .Y(n618) );
  OR2X1_HVT U44 ( .A1(n377), .A2(n359), .Y(n213) );
  NBUFFX2_HVT U45 ( .A(n763), .Y(n364) );
  MUX21X2_HVT U46 ( .A1(n476), .A2(n756), .S0(n367), .Y(n581) );
  INVX0_HVT U47 ( .A(n766), .Y(n467) );
  MUX41X1_HVT U48 ( .A1(n679), .A3(n680), .A2(n682), .A4(n687), .S0(n493), 
        .S1(n499), .Y(n678) );
  INVX1_HVT U49 ( .A(n506), .Y(n463) );
  INVX0_HVT U50 ( .A(n469), .Y(n119) );
  NAND2X0_HVT U51 ( .A1(n753), .A2(n211), .Y(n147) );
  AND2X1_HVT U52 ( .A1(n147), .A2(n148), .Y(n336) );
  OR2X1_HVT U54 ( .A1(n210), .A2(n457), .Y(n148) );
  INVX0_HVT U55 ( .A(n459), .Y(n210) );
  AND2X1_HVT U60 ( .A1(n324), .A2(n459), .Y(n211) );
  MUX41X1_HVT U64 ( .A1(n481), .A3(n477), .A2(n553), .A4(n691), .S0(n488), 
        .S1(n435), .Y(n690) );
  NAND2X0_HVT U65 ( .A1(n311), .A2(n312), .Y(n212) );
  INVX1_HVT U67 ( .A(n766), .Y(n380) );
  IBUFFX2_HVT U68 ( .A(n212), .Y(n536) );
  NAND2X0_HVT U70 ( .A1(n504), .A2(n216), .Y(n217) );
  NAND2X0_HVT U71 ( .A1(n217), .A2(n349), .Y(n589) );
  INVX0_HVT U72 ( .A(n451), .Y(n216) );
  MUX41X1_HVT U75 ( .A1(n578), .A3(n576), .A2(n579), .A4(n577), .S0(n118), 
        .S1(n495), .Y(n575) );
  INVX1_HVT U76 ( .A(n565), .Y(n273) );
  INVX1_HVT U77 ( .A(n417), .Y(n241) );
  AO21X1_HVT U78 ( .A1(n492), .A2(n241), .A3(n283), .Y(n658) );
  XNOR2X1_HVT U79 ( .A1(n433), .A2(n238), .Y(n236) );
  NBUFFX2_HVT U80 ( .A(n219), .Y(n419) );
  INVX1_HVT U81 ( .A(n515), .Y(n514) );
  NAND2X0_HVT U82 ( .A1(n697), .A2(n395), .Y(n335) );
  INVX1_HVT U86 ( .A(n746), .Y(n550) );
  INVX1_HVT U87 ( .A(n492), .Y(n338) );
  MUX21X1_HVT U88 ( .A1(n763), .A2(n399), .S0(n355), .Y(n688) );
  MUX21X1_HVT U89 ( .A1(n213), .A2(n399), .S0(n344), .Y(n410) );
  INVX1_HVT U91 ( .A(n492), .Y(n475) );
  INVX0_HVT U92 ( .A(n470), .Y(n471) );
  INVX1_HVT U93 ( .A(n419), .Y(n386) );
  INVX1_HVT U94 ( .A(n520), .Y(n465) );
  MUX21X1_HVT U95 ( .A1(n329), .A2(n315), .S0(n238), .Y(n765) );
  INVX1_HVT U96 ( .A(n490), .Y(n454) );
  INVX1_HVT U98 ( .A(n762), .Y(n558) );
  INVX1_HVT U99 ( .A(n488), .Y(n320) );
  NAND2X0_HVT U100 ( .A1(n725), .A2(n297), .Y(n415) );
  NAND2X0_HVT U102 ( .A1(n658), .A2(n297), .Y(n401) );
  INVX1_HVT U104 ( .A(n744), .Y(n549) );
  INVX0_HVT U106 ( .A(n492), .Y(n459) );
  INVX1_HVT U107 ( .A(in[7]), .Y(n520) );
  INVX1_HVT U108 ( .A(n520), .Y(n517) );
  INVX1_HVT U109 ( .A(n520), .Y(n332) );
  NBUFFX2_HVT U111 ( .A(n514), .Y(n489) );
  INVX1_HVT U112 ( .A(n517), .Y(n324) );
  INVX1_HVT U113 ( .A(n494), .Y(n325) );
  INVX1_HVT U114 ( .A(n314), .Y(n512) );
  NBUFFX2_HVT U116 ( .A(n514), .Y(n492) );
  INVX1_HVT U117 ( .A(n510), .Y(n347) );
  INVX1_HVT U118 ( .A(n496), .Y(n474) );
  INVX1_HVT U119 ( .A(n386), .Y(n328) );
  INVX1_HVT U120 ( .A(n374), .Y(n510) );
  INVX1_HVT U121 ( .A(n495), .Y(n252) );
  INVX0_HVT U122 ( .A(n520), .Y(n519) );
  INVX0_HVT U124 ( .A(n419), .Y(n326) );
  INVX0_HVT U126 ( .A(n512), .Y(n238) );
  INVX1_HVT U127 ( .A(n491), .Y(n444) );
  INVX1_HVT U128 ( .A(n499), .Y(n414) );
  INVX0_HVT U129 ( .A(n512), .Y(n508) );
  INVX1_HVT U130 ( .A(n398), .Y(n400) );
  INVX0_HVT U131 ( .A(n441), .Y(n354) );
  AND2X1_HVT U132 ( .A1(n321), .A2(n349), .Y(n218) );
  INVX1_HVT U133 ( .A(n743), .Y(n557) );
  INVX1_HVT U134 ( .A(n418), .Y(n341) );
  NBUFFX2_HVT U135 ( .A(n368), .Y(n498) );
  INVX0_HVT U136 ( .A(n313), .Y(n219) );
  INVX1_HVT U137 ( .A(n374), .Y(n344) );
  INVX1_HVT U138 ( .A(n526), .Y(n462) );
  MUX41X1_HVT U139 ( .A1(n662), .A3(n648), .A2(n656), .A4(n643), .S0(n391), 
        .S1(n414), .Y(out[3]) );
  XNOR2X2_HVT U140 ( .A1(n526), .A2(n272), .Y(n728) );
  AO21X1_HVT U141 ( .A1(n428), .A2(n417), .A3(n324), .Y(n674) );
  OA21X1_HVT U142 ( .A1(n482), .A2(n324), .A3(n220), .Y(n608) );
  INVX1_HVT U143 ( .A(n352), .Y(n756) );
  INVX1_HVT U144 ( .A(n316), .Y(n319) );
  INVX0_HVT U145 ( .A(n557), .Y(n220) );
  INVX0_HVT U146 ( .A(n742), .Y(n537) );
  INVX1_HVT U147 ( .A(n755), .Y(n551) );
  NAND2X0_HVT U148 ( .A1(n354), .A2(n227), .Y(n230) );
  NAND2X0_HVT U149 ( .A1(n317), .A2(n508), .Y(n231) );
  NAND2X0_HVT U150 ( .A1(n230), .A2(n231), .Y(n411) );
  INVX0_HVT U151 ( .A(n508), .Y(n227) );
  INVX0_HVT U152 ( .A(n316), .Y(n317) );
  MUX21X1_HVT U153 ( .A1(n411), .A2(n232), .S0(n490), .Y(n667) );
  NAND2X0_HVT U155 ( .A1(n509), .A2(n462), .Y(n232) );
  MUX41X1_HVT U156 ( .A1(n330), .A3(n731), .A2(n527), .A4(n556), .S0(n254), 
        .S1(n320), .Y(n631) );
  INVX1_HVT U157 ( .A(n768), .Y(n398) );
  INVX0_HVT U160 ( .A(n506), .Y(n486) );
  MUX21X2_HVT U161 ( .A1(n453), .A2(n460), .S0(n388), .Y(n753) );
  INVX0_HVT U163 ( .A(n363), .Y(n736) );
  INVX0_HVT U164 ( .A(n467), .Y(n472) );
  NBUFFX2_HVT U169 ( .A(n368), .Y(n497) );
  NBUFFX2_HVT U170 ( .A(n368), .Y(n496) );
  XNOR2X2_HVT U171 ( .A1(n318), .A2(n328), .Y(n481) );
  AND3X1_HVT U172 ( .A1(n460), .A2(n720), .A3(n696), .Y(n697) );
  XNOR2X1_HVT U173 ( .A1(n498), .A2(n747), .Y(n733) );
  INVX0_HVT U175 ( .A(n737), .Y(n524) );
  INVX1_HVT U176 ( .A(n505), .Y(n255) );
  INVX0_HVT U178 ( .A(n411), .Y(n740) );
  MUX41X1_HVT U180 ( .A1(n615), .A3(n610), .A2(n613), .A4(n607), .S0(n118), 
        .S1(n252), .Y(n606) );
  INVX1_HVT U181 ( .A(n261), .Y(n405) );
  MUX41X1_HVT U183 ( .A1(n542), .A3(n241), .A2(n356), .A4(n473), .S0(n489), 
        .S1(n433), .Y(n635) );
  MUX41X1_HVT U184 ( .A1(n632), .A3(n631), .A2(n409), .A4(n635), .S0(n252), 
        .S1(n499), .Y(n630) );
  XOR2X1_HVT U185 ( .A1(n511), .A2(n484), .Y(n487) );
  INVX1_HVT U186 ( .A(n703), .Y(n560) );
  MUX21X1_HVT U187 ( .A1(n213), .A2(n501), .S0(n361), .Y(n705) );
  MUX21X1_HVT U188 ( .A1(n538), .A2(n655), .S0(n491), .Y(n654) );
  NBUFFX2_HVT U189 ( .A(n465), .Y(n254) );
  MUX21X1_HVT U190 ( .A1(n503), .A2(n464), .S0(n388), .Y(n737) );
  MUX41X1_HVT U191 ( .A1(n690), .A3(n692), .A2(n694), .A4(n695), .S0(n493), 
        .S1(n499), .Y(n689) );
  INVX0_HVT U192 ( .A(n766), .Y(n329) );
  MUX41X1_HVT U193 ( .A1(n587), .A3(n583), .A2(n588), .A4(n586), .S0(n118), 
        .S1(n495), .Y(n582) );
  INVX1_HVT U194 ( .A(n255), .Y(n257) );
  INVX1_HVT U195 ( .A(n367), .Y(n368) );
  MUX21X1_HVT U196 ( .A1(n364), .A2(n471), .S0(n508), .Y(n670) );
  MUX21X1_HVT U198 ( .A1(n559), .A2(n504), .S0(n272), .Y(n261) );
  INVX1_HVT U199 ( .A(in[3]), .Y(n376) );
  MUX21X1_HVT U200 ( .A1(n468), .A2(n500), .S0(n38), .Y(n352) );
  INVX0_HVT U201 ( .A(n520), .Y(n466) );
  INVX1_HVT U202 ( .A(n364), .Y(n417) );
  NAND2X0_HVT U203 ( .A1(n289), .A2(n347), .Y(n264) );
  NAND2X0_HVT U205 ( .A1(n503), .A2(n508), .Y(n266) );
  NAND2X0_HVT U206 ( .A1(n264), .A2(n266), .Y(n761) );
  NAND2X0_HVT U207 ( .A1(n471), .A2(n355), .Y(n269) );
  MUX21X2_HVT U209 ( .A1(n743), .A2(n665), .S0(n489), .Y(n663) );
  NAND2X0_HVT U210 ( .A1(n238), .A2(n763), .Y(n720) );
  INVX1_HVT U211 ( .A(n219), .Y(n374) );
  INVX1_HVT U212 ( .A(n213), .Y(n554) );
  NBUFFX2_HVT U213 ( .A(n314), .Y(n272) );
  XNOR2X1_HVT U216 ( .A1(n400), .A2(n508), .Y(n478) );
  XNOR2X2_HVT U217 ( .A1(n227), .A2(n554), .Y(n732) );
  INVX0_HVT U219 ( .A(n565), .Y(n548) );
  INVX0_HVT U221 ( .A(n386), .Y(n361) );
  MUX21X2_HVT U222 ( .A1(n317), .A2(n213), .S0(n510), .Y(n743) );
  MUX41X1_HVT U223 ( .A1(n23), .A3(n667), .A2(n663), .A4(n666), .S0(n493), 
        .S1(n254), .Y(n662) );
  MUX41X1_HVT U224 ( .A1(n736), .A3(n337), .A2(n434), .A4(n257), .S0(n496), 
        .S1(n485), .Y(n587) );
  NAND2X0_HVT U225 ( .A1(n329), .A2(n347), .Y(n275) );
  NAND2X0_HVT U226 ( .A1(n364), .A2(n361), .Y(n279) );
  NAND2X0_HVT U227 ( .A1(n269), .A2(n279), .Y(n434) );
  INVX1_HVT U228 ( .A(n484), .Y(n485) );
  INVX0_HVT U229 ( .A(n761), .Y(n545) );
  MUX41X1_HVT U230 ( .A1(n232), .A3(n441), .A2(n557), .A4(n3), .S0(n454), .S1(
        n465), .Y(n576) );
  MUX21X2_HVT U231 ( .A1(n563), .A2(n273), .S0(n497), .Y(n585) );
  XNOR2X2_HVT U232 ( .A1(n375), .A2(n360), .Y(n766) );
  MUX41X1_HVT U233 ( .A1(n601), .A3(n604), .A2(n600), .A4(n602), .S0(n499), 
        .S1(n252), .Y(n599) );
  NAND2X0_HVT U234 ( .A1(n550), .A2(n338), .Y(n280) );
  NAND2X0_HVT U235 ( .A1(n744), .A2(n513), .Y(n282) );
  NAND2X0_HVT U236 ( .A1(n280), .A2(n282), .Y(n647) );
  MUX41X1_HVT U237 ( .A1(n647), .A3(n646), .A2(n645), .A4(n644), .S0(n297), 
        .S1(n325), .Y(n643) );
  MUX21X1_HVT U238 ( .A1(n331), .A2(n357), .S0(n326), .Y(n681) );
  INVX1_HVT U239 ( .A(n466), .Y(n433) );
  MUX41X1_HVT U240 ( .A1(n711), .A3(n710), .A2(n709), .A4(n531), .S0(n297), 
        .S1(n320), .Y(n708) );
  INVX0_HVT U243 ( .A(n357), .Y(n283) );
  INVX1_HVT U244 ( .A(in[1]), .Y(n313) );
  NBUFFX2_HVT U246 ( .A(n770), .Y(n506) );
  INVX1_HVT U247 ( .A(n419), .Y(n428) );
  NBUFFX2_HVT U248 ( .A(n430), .Y(n501) );
  INVX1_HVT U249 ( .A(n501), .Y(n306) );
  MUX21X1_HVT U250 ( .A1(n634), .A2(n633), .S0(n491), .Y(n632) );
  NAND2X0_HVT U251 ( .A1(n713), .A2(n444), .Y(n284) );
  NAND2X0_HVT U252 ( .A1(n715), .A2(n395), .Y(n285) );
  NAND2X0_HVT U253 ( .A1(n284), .A2(n285), .Y(n712) );
  INVX0_HVT U254 ( .A(n765), .Y(n531) );
  INVX1_HVT U255 ( .A(n512), .Y(n511) );
  NAND2X0_HVT U257 ( .A1(n502), .A2(n562), .Y(n289) );
  MUX41X1_HVT U258 ( .A1(n528), .A3(n732), .A2(n758), .A4(n564), .S0(n320), 
        .S1(n518), .Y(n694) );
  INVX1_HVT U259 ( .A(n515), .Y(n513) );
  INVX1_HVT U260 ( .A(n487), .Y(n369) );
  INVX0_HVT U261 ( .A(n498), .Y(n297) );
  INVX1_HVT U262 ( .A(in[4]), .Y(n430) );
  NAND2X0_HVT U263 ( .A1(n668), .A2(n391), .Y(n290) );
  NAND2X0_HVT U264 ( .A1(n678), .A2(n327), .Y(n292) );
  NAND2X0_HVT U265 ( .A1(n290), .A2(n292), .Y(out[2]) );
  MUX41X1_HVT U266 ( .A1(n676), .A3(n672), .A2(n671), .A4(n669), .S0(n325), 
        .S1(n118), .Y(n668) );
  NAND2X0_HVT U267 ( .A1(n480), .A2(n394), .Y(n293) );
  NAND2X0_HVT U269 ( .A1(n677), .A2(n730), .Y(n294) );
  NAND2X0_HVT U271 ( .A1(n293), .A2(n294), .Y(n676) );
  INVX1_HVT U272 ( .A(n394), .Y(n730) );
  INVX0_HVT U273 ( .A(n497), .Y(n435) );
  INVX0_HVT U274 ( .A(n741), .Y(n547) );
  OA21X1_HVT U275 ( .A1(n737), .A2(n435), .A3(n627), .Y(n628) );
  INVX0_HVT U276 ( .A(n305), .Y(n686) );
  NAND2X0_HVT U277 ( .A1(n297), .A2(n533), .Y(n303) );
  NAND2X0_HVT U278 ( .A1(n417), .A2(n496), .Y(n304) );
  NAND2X0_HVT U279 ( .A1(n303), .A2(n304), .Y(n629) );
  MUX41X1_HVT U280 ( .A1(n480), .A3(n547), .A2(n665), .A4(n461), .S0(n254), 
        .S1(n320), .Y(n625) );
  MUX21X1_HVT U281 ( .A1(n503), .A2(n306), .S0(n498), .Y(n305) );
  NAND2X0_HVT U282 ( .A1(n608), .A2(n210), .Y(n307) );
  NAND2X0_HVT U283 ( .A1(n609), .A2(n444), .Y(n308) );
  NAND2X0_HVT U285 ( .A1(n307), .A2(n308), .Y(n607) );
  NAND2X0_HVT U286 ( .A1(n727), .A2(n490), .Y(n309) );
  NAND2X0_HVT U287 ( .A1(n723), .A2(n444), .Y(n310) );
  NAND2X0_HVT U288 ( .A1(n309), .A2(n310), .Y(n722) );
  INVX1_HVT U290 ( .A(n572), .Y(n534) );
  OA21X1_HVT U291 ( .A1(n525), .A2(n324), .A3(n743), .Y(n633) );
  NAND2X0_HVT U292 ( .A1(n289), .A2(n355), .Y(n311) );
  NAND2X0_HVT U293 ( .A1(n472), .A2(n510), .Y(n312) );
  INVX1_HVT U294 ( .A(n313), .Y(n314) );
  XOR2X1_HVT U297 ( .A1(n238), .A2(n500), .Y(n729) );
  MUX21X1_HVT U298 ( .A1(n317), .A2(n399), .S0(n512), .Y(n683) );
  INVX0_HVT U299 ( .A(n419), .Y(n355) );
  INVX1_HVT U300 ( .A(n428), .Y(n509) );
  INVX1_HVT U301 ( .A(n430), .Y(n375) );
  INVX1_HVT U302 ( .A(n507), .Y(n315) );
  NAND2X0_HVT U303 ( .A1(n461), .A2(n227), .Y(n321) );
  INVX0_HVT U304 ( .A(n486), .Y(n461) );
  INVX1_HVT U305 ( .A(n520), .Y(n518) );
  INVX1_HVT U307 ( .A(n472), .Y(n473) );
  AO21X1_HVT U308 ( .A1(n496), .A2(n683), .A3(n552), .Y(n684) );
  INVX1_HVT U310 ( .A(n683), .Y(n541) );
  NAND2X0_HVT U311 ( .A1(n463), .A2(n347), .Y(n322) );
  NAND2X0_HVT U312 ( .A1(n500), .A2(n38), .Y(n323) );
  NAND2X0_HVT U313 ( .A1(n322), .A2(n323), .Y(n754) );
  NBUFFX2_HVT U314 ( .A(n35), .Y(n500) );
  MUX41X1_HVT U315 ( .A1(n528), .A3(n522), .A2(n544), .A4(n218), .S0(n324), 
        .S1(n325), .Y(n727) );
  OA21X1_HVT U316 ( .A1(n435), .A2(n765), .A3(n408), .Y(n580) );
  INVX1_HVT U317 ( .A(n571), .Y(n555) );
  INVX0_HVT U318 ( .A(in[7]), .Y(n367) );
  INVX1_HVT U319 ( .A(n376), .Y(n360) );
  MUX21X1_HVT U320 ( .A1(n504), .A2(n453), .S0(n388), .Y(n744) );
  MUX21X1_HVT U321 ( .A1(n751), .A2(n539), .S0(n466), .Y(n638) );
  NAND2X0_HVT U322 ( .A1(n582), .A2(in[6]), .Y(n431) );
  INVX0_HVT U323 ( .A(n512), .Y(n451) );
  INVX0_HVT U324 ( .A(n374), .Y(n388) );
  INVX1_HVT U325 ( .A(n391), .Y(n327) );
  INVX1_HVT U326 ( .A(in[6]), .Y(n391) );
  INVX1_HVT U327 ( .A(n343), .Y(n731) );
  MUX41X1_HVT U328 ( .A1(n641), .A3(n640), .A2(n639), .A4(n637), .S0(n325), 
        .S1(n414), .Y(n636) );
  INVX0_HVT U329 ( .A(n452), .Y(n745) );
  INVX1_HVT U330 ( .A(n560), .Y(n330) );
  MUX41X1_HVT U331 ( .A1(n749), .A3(n19), .A2(n408), .A4(n537), .S0(n254), 
        .S1(n513), .Y(n409) );
  INVX1_HVT U332 ( .A(n768), .Y(n331) );
  INVX1_HVT U333 ( .A(n440), .Y(n748) );
  NAND2X0_HVT U334 ( .A1(n289), .A2(n347), .Y(n333) );
  NAND2X0_HVT U335 ( .A1(n500), .A2(n358), .Y(n334) );
  NAND2X0_HVT U336 ( .A1(n333), .A2(n334), .Y(n764) );
  INVX1_HVT U337 ( .A(n764), .Y(n546) );
  NAND2X0_HVT U338 ( .A1(n335), .A2(n336), .Y(n695) );
  INVX1_HVT U339 ( .A(n753), .Y(n528) );
  NAND2X0_HVT U340 ( .A1(n322), .A2(n387), .Y(n337) );
  NAND2X0_HVT U341 ( .A1(n557), .A2(n338), .Y(n339) );
  NAND2X0_HVT U342 ( .A1(n758), .A2(n492), .Y(n340) );
  NAND2X0_HVT U343 ( .A1(n339), .A2(n340), .Y(n677) );
  NAND2X0_HVT U344 ( .A1(n511), .A2(n317), .Y(n703) );
  MUX21X1_HVT U345 ( .A1(n486), .A2(n255), .S0(n508), .Y(n407) );
  INVX1_HVT U346 ( .A(n738), .Y(n539) );
  MUX41X1_HVT U347 ( .A1(n417), .A3(n434), .A2(n337), .A4(n767), .S0(n475), 
        .S1(n517), .Y(n640) );
  INVX0_HVT U348 ( .A(n770), .Y(n464) );
  NBUFFX2_HVT U349 ( .A(n759), .Y(n342) );
  XOR2X1_HVT U350 ( .A1(n329), .A2(n344), .Y(n343) );
  MUX41X1_HVT U351 ( .A1(n738), .A3(n479), .A2(n731), .A4(n330), .S0(n338), 
        .S1(n519), .Y(n594) );
  NAND2X0_HVT U352 ( .A1(n653), .A2(n254), .Y(n345) );
  NAND2X0_HVT U353 ( .A1(n654), .A2(n324), .Y(n346) );
  NAND2X0_HVT U354 ( .A1(n345), .A2(n346), .Y(n650) );
  MUX21X1_HVT U355 ( .A1(n501), .A2(n504), .S0(n451), .Y(n655) );
  MUX21X1_HVT U356 ( .A1(n469), .A2(n463), .S0(n38), .Y(n749) );
  NAND2X0_HVT U357 ( .A1(n501), .A2(n344), .Y(n349) );
  NAND2X0_HVT U358 ( .A1(n348), .A2(n349), .Y(n700) );
  INVX1_HVT U359 ( .A(n398), .Y(n399) );
  NAND2X0_HVT U360 ( .A1(n490), .A2(n352), .Y(n350) );
  NAND2X0_HVT U361 ( .A1(n478), .A2(n338), .Y(n351) );
  NAND2X0_HVT U362 ( .A1(n350), .A2(n351), .Y(n645) );
  INVX0_HVT U363 ( .A(n82), .Y(n538) );
  OA21X1_HVT U364 ( .A1(n536), .A2(n454), .A3(n410), .Y(n666) );
  MUX21X1_HVT U365 ( .A1(n504), .A2(n354), .S0(n489), .Y(n353) );
  INVX1_HVT U366 ( .A(n570), .Y(n553) );
  AND2X1_HVT U367 ( .A1(n362), .A2(n275), .Y(n356) );
  INVX0_HVT U368 ( .A(n469), .Y(n357) );
  INVX0_HVT U369 ( .A(n467), .Y(n469) );
  OR2X1_HVT U370 ( .A1(n35), .A2(n359), .Y(n763) );
  NAND2X0_HVT U371 ( .A1(n406), .A2(n361), .Y(n362) );
  NAND2X0_HVT U372 ( .A1(n275), .A2(n362), .Y(n751) );
  MUX21X1_HVT U373 ( .A1(n464), .A2(n472), .S0(n358), .Y(n363) );
  MUX41X1_HVT U374 ( .A1(n728), .A3(n589), .A2(n735), .A4(n741), .S0(n489), 
        .S1(n433), .Y(n588) );
  MUX41X1_HVT U375 ( .A1(n479), .A3(n564), .A2(n681), .A4(n555), .S0(n444), 
        .S1(n465), .Y(n680) );
  NAND2X0_HVT U376 ( .A1(n441), .A2(n347), .Y(n365) );
  NBUFFX2_HVT U377 ( .A(n470), .Y(n366) );
  NAND2X0_HVT U378 ( .A1(n405), .A2(n210), .Y(n403) );
  NAND2X0_HVT U379 ( .A1(n464), .A2(n369), .Y(n370) );
  NAND2X0_HVT U380 ( .A1(n353), .A2(n487), .Y(n371) );
  INVX1_HVT U381 ( .A(n407), .Y(n758) );
  NAND2X0_HVT U382 ( .A1(n537), .A2(n491), .Y(n372) );
  NAND2X0_HVT U383 ( .A1(n755), .A2(n454), .Y(n373) );
  NAND2X0_HVT U384 ( .A1(n373), .A2(n372), .Y(n644) );
  NBUFFX2_HVT U385 ( .A(n514), .Y(n491) );
  MUX41X1_HVT U386 ( .A1(n527), .A3(n477), .A2(n740), .A4(n82), .S0(n474), 
        .S1(n489), .Y(n639) );
  NAND2X0_HVT U387 ( .A1(n717), .A2(n444), .Y(n378) );
  NAND2X0_HVT U388 ( .A1(n719), .A2(n490), .Y(n379) );
  NAND2X0_HVT U389 ( .A1(n378), .A2(n379), .Y(n716) );
  MUX21X1_HVT U390 ( .A1(n503), .A2(n315), .S0(n509), .Y(n762) );
  NBUFFX2_HVT U391 ( .A(n430), .Y(n502) );
  NAND2X0_HVT U392 ( .A1(n745), .A2(n435), .Y(n436) );
  MUX41X1_HVT U393 ( .A1(n555), .A3(n366), .A2(n212), .A4(n318), .S0(n338), 
        .S1(n466), .Y(n586) );
  INVX1_HVT U394 ( .A(n507), .Y(n559) );
  NAND2X0_HVT U395 ( .A1(n624), .A2(n381), .Y(n382) );
  NAND2X0_HVT U396 ( .A1(n461), .A2(n236), .Y(n383) );
  NAND2X0_HVT U397 ( .A1(n382), .A2(n383), .Y(n623) );
  INVX0_HVT U398 ( .A(n236), .Y(n381) );
  MUX21X1_HVT U399 ( .A1(n500), .A2(n741), .S0(n493), .Y(n726) );
  NAND2X0_HVT U400 ( .A1(n707), .A2(n395), .Y(n384) );
  NAND2X0_HVT U401 ( .A1(n733), .A2(n444), .Y(n385) );
  NAND2X0_HVT U402 ( .A1(n384), .A2(n385), .Y(n706) );
  NAND2X0_HVT U403 ( .A1(n315), .A2(n272), .Y(n387) );
  NAND2X0_HVT U404 ( .A1(n322), .A2(n387), .Y(n747) );
  NAND2X0_HVT U405 ( .A1(n596), .A2(n444), .Y(n389) );
  NAND2X0_HVT U406 ( .A1(n597), .A2(n490), .Y(n390) );
  NAND2X0_HVT U407 ( .A1(n389), .A2(n390), .Y(n595) );
  NAND2X0_HVT U408 ( .A1(n590), .A2(n391), .Y(n392) );
  NAND2X0_HVT U409 ( .A1(n599), .A2(n327), .Y(n393) );
  NAND2X0_HVT U410 ( .A1(n392), .A2(n393), .Y(out[6]) );
  MUX21X1_HVT U411 ( .A1(n691), .A2(n406), .S0(n496), .Y(n597) );
  NBUFFX2_HVT U412 ( .A(n514), .Y(n490) );
  XNOR2X1_HVT U413 ( .A1(n395), .A2(n368), .Y(n394) );
  NAND2X0_HVT U414 ( .A1(n769), .A2(n395), .Y(n396) );
  NAND2X0_HVT U415 ( .A1(n638), .A2(n475), .Y(n397) );
  NAND2X0_HVT U416 ( .A1(n397), .A2(n396), .Y(n637) );
  INVX0_HVT U417 ( .A(n475), .Y(n395) );
  NAND2X0_HVT U418 ( .A1(n502), .A2(n562), .Y(n768) );
  NAND2X0_HVT U419 ( .A1(n659), .A2(n496), .Y(n402) );
  NAND2X0_HVT U420 ( .A1(n401), .A2(n402), .Y(n657) );
  NAND2X0_HVT U421 ( .A1(n547), .A2(n338), .Y(n404) );
  NAND2X0_HVT U422 ( .A1(n403), .A2(n404), .Y(n659) );
  INVX0_HVT U423 ( .A(n664), .Y(n542) );
  INVX0_HVT U424 ( .A(n408), .Y(n739) );
  INVX1_HVT U425 ( .A(n569), .Y(n533) );
  MUX21X1_HVT U426 ( .A1(n317), .A2(n289), .S0(n272), .Y(n408) );
  MUX41X1_HVT U427 ( .A1(n603), .A3(n755), .A2(n739), .A4(n548), .S0(n338), 
        .S1(n518), .Y(n602) );
  NAND2X0_HVT U428 ( .A1(n649), .A2(n252), .Y(n412) );
  NAND2X0_HVT U429 ( .A1(n650), .A2(n495), .Y(n413) );
  NAND2X0_HVT U430 ( .A1(n412), .A2(n413), .Y(n648) );
  MUX41X1_HVT U431 ( .A1(n595), .A3(n598), .A2(n591), .A4(n594), .S0(n495), 
        .S1(n414), .Y(n590) );
  NAND2X0_HVT U432 ( .A1(n726), .A2(n498), .Y(n416) );
  NAND2X0_HVT U433 ( .A1(n415), .A2(n416), .Y(n723) );
  AND2X1_HVT U434 ( .A1(n342), .A2(n319), .Y(n418) );
  MUX41X1_HVT U435 ( .A1(n341), .A3(n476), .A2(n530), .A4(n764), .S0(n498), 
        .S1(n454), .Y(n600) );
  MUX41X1_HVT U436 ( .A1(n593), .A3(n543), .A2(n592), .A4(n342), .S0(n496), 
        .S1(n475), .Y(n591) );
  NAND2X0_HVT U437 ( .A1(n657), .A2(n252), .Y(n420) );
  NAND2X0_HVT U438 ( .A1(n660), .A2(n516), .Y(n421) );
  NAND2X0_HVT U439 ( .A1(n420), .A2(n421), .Y(n656) );
  NAND2X0_HVT U440 ( .A1(n689), .A2(n391), .Y(n422) );
  NAND2X0_HVT U441 ( .A1(n698), .A2(n327), .Y(n423) );
  NAND2X0_HVT U442 ( .A1(n423), .A2(n422), .Y(out[1]) );
  MUX41X1_HVT U443 ( .A1(n706), .A3(n702), .A2(n701), .A4(n699), .S0(n252), 
        .S1(n414), .Y(n698) );
  NAND2X0_HVT U444 ( .A1(n622), .A2(n444), .Y(n424) );
  NAND2X0_HVT U445 ( .A1(n623), .A2(n492), .Y(n425) );
  NAND2X0_HVT U446 ( .A1(n425), .A2(n424), .Y(n621) );
  NAND2X0_HVT U447 ( .A1(n606), .A2(n391), .Y(n426) );
  NAND2X0_HVT U448 ( .A1(n618), .A2(n327), .Y(n427) );
  NAND2X0_HVT U449 ( .A1(n427), .A2(n426), .Y(out[5]) );
  MUX21X1_HVT U450 ( .A1(n739), .A2(n541), .S0(n498), .Y(n622) );
  INVX1_HVT U451 ( .A(n566), .Y(n527) );
  MUX41X1_HVT U452 ( .A1(n617), .A3(n478), .A2(n616), .A4(n551), .S0(n484), 
        .S1(n435), .Y(n615) );
  INVX1_HVT U453 ( .A(n458), .Y(n429) );
  MUX41X1_HVT U454 ( .A1(n523), .A3(n220), .A2(n341), .A4(n661), .S0(n513), 
        .S1(n474), .Y(n660) );
  NAND2X0_HVT U455 ( .A1(n575), .A2(n391), .Y(n432) );
  NAND2X0_HVT U456 ( .A1(n432), .A2(n431), .Y(out[7]) );
  NAND2X0_HVT U457 ( .A1(n458), .A2(n498), .Y(n437) );
  NAND2X0_HVT U458 ( .A1(n436), .A2(n437), .Y(n634) );
  NAND2X0_HVT U459 ( .A1(n630), .A2(n391), .Y(n438) );
  NAND2X0_HVT U460 ( .A1(n636), .A2(n327), .Y(n439) );
  NAND2X0_HVT U461 ( .A1(n438), .A2(n439), .Y(out[4]) );
  XNOR2X1_HVT U462 ( .A1(n441), .A2(n216), .Y(n440) );
  NAND2X0_HVT U463 ( .A1(n585), .A2(n459), .Y(n442) );
  NAND2X0_HVT U464 ( .A1(n584), .A2(n490), .Y(n443) );
  NAND2X0_HVT U465 ( .A1(n442), .A2(n443), .Y(n583) );
  NAND2X0_HVT U466 ( .A1(n521), .A2(n444), .Y(n445) );
  NAND2X0_HVT U467 ( .A1(n642), .A2(n491), .Y(n446) );
  NAND2X0_HVT U468 ( .A1(n445), .A2(n446), .Y(n641) );
  MUX21X1_HVT U469 ( .A1(n540), .A2(n257), .S0(n496), .Y(n642) );
  INVX1_HVT U470 ( .A(n568), .Y(n521) );
  INVX1_HVT U471 ( .A(n567), .Y(n540) );
  NAND2X0_HVT U472 ( .A1(n461), .A2(n381), .Y(n447) );
  NAND2X0_HVT U473 ( .A1(n686), .A2(n236), .Y(n448) );
  NAND2X0_HVT U474 ( .A1(n447), .A2(n448), .Y(n685) );
  NAND2X0_HVT U475 ( .A1(n684), .A2(n444), .Y(n449) );
  NAND2X0_HVT U476 ( .A1(n685), .A2(n492), .Y(n450) );
  NAND2X0_HVT U477 ( .A1(n449), .A2(n450), .Y(n682) );
  MUX21X1_HVT U478 ( .A1(n453), .A2(n400), .S0(n388), .Y(n452) );
  NAND2X0_HVT U479 ( .A1(n580), .A2(n454), .Y(n455) );
  NAND2X0_HVT U480 ( .A1(n581), .A2(n490), .Y(n456) );
  NAND2X0_HVT U481 ( .A1(n456), .A2(n455), .Y(n579) );
  NAND2X0_HVT U482 ( .A1(n364), .A2(n519), .Y(n457) );
  AND2X1_HVT U483 ( .A1(n509), .A2(n462), .Y(n458) );
  INVX1_HVT U484 ( .A(n380), .Y(n470) );
  AND2X1_HVT U485 ( .A1(n357), .A2(n720), .Y(n476) );
  MUX21X1_HVT U486 ( .A1(n331), .A2(n315), .S0(n493), .Y(n724) );
  AND2X1_HVT U487 ( .A1(n462), .A2(n703), .Y(n477) );
  MUX21X1_HVT U488 ( .A1(n546), .A2(n417), .S0(n493), .Y(n709) );
  MUX21X1_HVT U489 ( .A1(n331), .A2(n464), .S0(n328), .Y(n605) );
  MUX21X1_HVT U490 ( .A1(n315), .A2(n119), .S0(n328), .Y(n617) );
  MUX21X1_HVT U491 ( .A1(n331), .A2(n501), .S0(n511), .Y(n567) );
  MUX21X1_HVT U492 ( .A1(n503), .A2(n468), .S0(n344), .Y(n569) );
  MUX21X1_HVT U493 ( .A1(n504), .A2(n318), .S0(n358), .Y(n592) );
  MUX21X1_HVT U494 ( .A1(n318), .A2(n461), .S0(n358), .Y(n593) );
  MUX21X1_HVT U495 ( .A1(n462), .A2(n400), .S0(n238), .Y(n566) );
  AND2X1_HVT U496 ( .A1(n511), .A2(n463), .Y(n479) );
  MUX21X1_HVT U497 ( .A1(n213), .A2(n503), .S0(n510), .Y(n571) );
  AND2X1_HVT U498 ( .A1(n319), .A2(n664), .Y(n480) );
  MUX21X1_HVT U499 ( .A1(n257), .A2(n319), .S0(n491), .Y(n652) );
  NBUFFX2_HVT U500 ( .A(n562), .Y(n503) );
  NBUFFX2_HVT U501 ( .A(n562), .Y(n504) );
  NBUFFX2_HVT U502 ( .A(n516), .Y(n495) );
  NBUFFX2_HVT U503 ( .A(n516), .Y(n494) );
  NBUFFX2_HVT U504 ( .A(n513), .Y(n488) );
  NBUFFX2_HVT U505 ( .A(n516), .Y(n493) );
  MUX21X1_HVT U506 ( .A1(n675), .A2(n521), .S0(n491), .Y(n672) );
  MUX21X1_HVT U507 ( .A1(n406), .A2(n398), .S0(n451), .Y(n738) );
  MUX21X1_HVT U508 ( .A1(n241), .A2(n555), .S0(n497), .Y(n609) );
  NAND2X0_HVT U509 ( .A1(n35), .A2(n502), .Y(n770) );
  AND2X1_HVT U510 ( .A1(n471), .A2(n355), .Y(n482) );
  MUX21X1_HVT U511 ( .A1(n559), .A2(n555), .S0(n497), .Y(n707) );
  MUX21X1_HVT U512 ( .A1(n554), .A2(n464), .S0(n272), .Y(n614) );
  NBUFFX2_HVT U513 ( .A(n771), .Y(n507) );
  MUX21X1_HVT U514 ( .A1(n429), .A2(n326), .S0(n490), .Y(n651) );
  MUX21X1_HVT U515 ( .A1(n744), .A2(n573), .S0(n497), .Y(n568) );
  MUX21X1_HVT U516 ( .A1(n406), .A2(n554), .S0(n272), .Y(n570) );
  XOR2X1_HVT U517 ( .A1(n361), .A2(n495), .Y(n734) );
  NBUFFX2_HVT U518 ( .A(n763), .Y(n505) );
  MUX21X1_HVT U519 ( .A1(n545), .A2(n326), .S0(n493), .Y(n711) );
  INVX1_HVT U520 ( .A(n377), .Y(n562) );
  AND2X1_HVT U521 ( .A1(n503), .A2(n428), .Y(n483) );
  NBUFFX2_HVT U522 ( .A(in[5]), .Y(n516) );
  NAND2X0_HVT U523 ( .A1(n377), .A2(n375), .Y(n771) );
  MUX21X1_HVT U524 ( .A1(n441), .A2(n366), .S0(n344), .Y(n572) );
  MUX21X1_HVT U525 ( .A1(n318), .A2(n441), .S0(n344), .Y(n746) );
  MUX21X1_HVT U526 ( .A1(n453), .A2(n505), .S0(n328), .Y(n565) );
  NBUFFX2_HVT U527 ( .A(in[0]), .Y(n499) );
  INVX1_HVT U528 ( .A(in[2]), .Y(n515) );
endmodule

