
module inv_sbox_2 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n6, n58, n196, n197, n198, n199, n200, n201, n202, n206, n208, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598;

  NAND2X0_HVT U1 ( .A1(n258), .A2(n392), .Y(n598) );
  NAND2X0_HVT U5 ( .A1(n265), .A2(n269), .Y(n594) );
  NAND2X0_HVT U6 ( .A1(n326), .A2(n305), .Y(n593) );
  NAND2X0_HVT U7 ( .A1(n252), .A2(n322), .Y(n592) );
  NAND2X0_HVT U8 ( .A1(n251), .A2(n268), .Y(n591) );
  NAND2X0_HVT U9 ( .A1(n301), .A2(n591), .Y(n590) );
  NAND2X0_HVT U10 ( .A1(n305), .A2(n588), .Y(n589) );
  NAND2X0_HVT U11 ( .A1(n330), .A2(n263), .Y(n587) );
  NAND2X0_HVT U12 ( .A1(n326), .A2(n317), .Y(n586) );
  NAND2X0_HVT U13 ( .A1(n323), .A2(n591), .Y(n585) );
  NAND2X0_HVT U15 ( .A1(n284), .A2(n328), .Y(n583) );
  NAND2X0_HVT U19 ( .A1(n325), .A2(n391), .Y(n578) );
  NAND2X0_HVT U32 ( .A1(n318), .A2(n330), .Y(n566) );
  NAND2X0_HVT U35 ( .A1(n591), .A2(n291), .Y(n563) );
  NAND2X0_HVT U38 ( .A1(n317), .A2(n330), .Y(n560) );
  NAND2X0_HVT U42 ( .A1(n593), .A2(n286), .Y(n556) );
  NAND2X0_HVT U55 ( .A1(n323), .A2(n595), .Y(n544) );
  AO21X1_HVT U60 ( .A1(n539), .A2(n314), .A3(n577), .Y(n540) );
  MUX41X1_HVT U62 ( .A1(n538), .A3(n543), .A2(n542), .A4(n545), .S0(n321), 
        .S1(n248), .Y(n537) );
  MUX41X1_HVT U65 ( .A1(n356), .A3(n358), .A2(n357), .A4(n560), .S0(n312), 
        .S1(n245), .Y(n534) );
  NAND2X0_HVT U66 ( .A1(n252), .A2(n273), .Y(n533) );
  MUX41X1_HVT U67 ( .A1(n353), .A3(n377), .A2(n355), .A4(n533), .S0(n316), 
        .S1(n309), .Y(n532) );
  MUX41X1_HVT U71 ( .A1(n593), .A3(n303), .A2(n587), .A4(n349), .S0(n311), 
        .S1(n244), .Y(n529) );
  NAND2X0_HVT U72 ( .A1(n285), .A2(n592), .Y(n528) );
  MUX41X1_HVT U73 ( .A1(n571), .A3(n528), .A2(n378), .A4(n257), .S0(n315), 
        .S1(n308), .Y(n527) );
  MUX41X1_HVT U74 ( .A1(n589), .A3(n369), .A2(n368), .A4(n359), .S0(n312), 
        .S1(n245), .Y(n526) );
  MUX41X1_HVT U80 ( .A1(n379), .A3(n376), .A2(n590), .A4(n594), .S0(n311), 
        .S1(n244), .Y(n520) );
  NAND2X0_HVT U81 ( .A1(n597), .A2(n592), .Y(n519) );
  AND2X1_HVT U82 ( .A1(n593), .A2(n596), .Y(n518) );
  MUX41X1_HVT U83 ( .A1(n518), .A3(n366), .A2(n292), .A4(n519), .S0(n311), 
        .S1(n245), .Y(n517) );
  MUX41X1_HVT U84 ( .A1(n299), .A3(n365), .A2(n380), .A4(n241), .S0(n312), 
        .S1(n333), .Y(n516) );
  MUX41X1_HVT U85 ( .A1(n516), .A3(n520), .A2(n517), .A4(n521), .S0(n321), 
        .S1(n248), .Y(n515) );
  MUX41X1_HVT U88 ( .A1(n355), .A3(n340), .A2(n568), .A4(n552), .S0(n311), 
        .S1(n334), .Y(n513) );
  NAND2X0_HVT U89 ( .A1(n330), .A2(n270), .Y(n512) );
  MUX41X1_HVT U95 ( .A1(n507), .A3(n513), .A2(n511), .A4(n514), .S0(n321), 
        .S1(n319), .Y(n506) );
  MUX41X1_HVT U96 ( .A1(n377), .A3(n585), .A2(n223), .A4(n382), .S0(n312), 
        .S1(n333), .Y(n505) );
  MUX41X1_HVT U98 ( .A1(n504), .A3(n383), .A2(n370), .A4(n570), .S0(n312), 
        .S1(n244), .Y(n503) );
  MUX41X1_HVT U99 ( .A1(n566), .A3(n357), .A2(n550), .A4(n284), .S0(n334), 
        .S1(n309), .Y(n502) );
  NAND2X0_HVT U100 ( .A1(n330), .A2(n262), .Y(n501) );
  MUX41X1_HVT U101 ( .A1(n384), .A3(n586), .A2(n264), .A4(n501), .S0(n334), 
        .S1(n307), .Y(n500) );
  MUX41X1_HVT U102 ( .A1(n500), .A3(n503), .A2(n502), .A4(n505), .S0(n321), 
        .S1(n248), .Y(n499) );
  AND2X1_HVT U104 ( .A1(n592), .A2(n269), .Y(n498) );
  MUX41X1_HVT U105 ( .A1(n584), .A3(n385), .A2(n519), .A4(n498), .S0(n312), 
        .S1(n244), .Y(n497) );
  MUX41X1_HVT U107 ( .A1(n384), .A3(n596), .A2(n496), .A4(n346), .S0(n311), 
        .S1(n334), .Y(n495) );
  MUX41X1_HVT U108 ( .A1(n359), .A3(n288), .A2(n362), .A4(n597), .S0(n312), 
        .S1(n333), .Y(n494) );
  MUX41X1_HVT U109 ( .A1(n383), .A3(n340), .A2(n380), .A4(n374), .S0(n311), 
        .S1(n238), .Y(n493) );
  MUX41X1_HVT U110 ( .A1(n493), .A3(n495), .A2(n494), .A4(n497), .S0(n321), 
        .S1(n319), .Y(n492) );
  AO21X1_HVT U112 ( .A1(n371), .A2(n315), .A3(n574), .Y(n490) );
  NAND2X0_HVT U114 ( .A1(n301), .A2(n592), .Y(n488) );
  MUX41X1_HVT U115 ( .A1(n488), .A3(n587), .A2(n371), .A4(n596), .S0(n334), 
        .S1(n309), .Y(n487) );
  MUX41X1_HVT U116 ( .A1(n282), .A3(n365), .A2(n340), .A4(n583), .S0(n310), 
        .S1(n334), .Y(n486) );
  NAND2X0_HVT U118 ( .A1(n330), .A2(n258), .Y(n484) );
  MUX41X1_HVT U119 ( .A1(n386), .A3(n485), .A2(n561), .A4(n484), .S0(n310), 
        .S1(n333), .Y(n483) );
  MUX41X1_HVT U120 ( .A1(n483), .A3(n487), .A2(n486), .A4(n489), .S0(in[5]), 
        .S1(n319), .Y(n482) );
  MUX41X1_HVT U122 ( .A1(n375), .A3(n295), .A2(n552), .A4(n261), .S0(n310), 
        .S1(n333), .Y(n481) );
  MUX41X1_HVT U124 ( .A1(n297), .A3(n480), .A2(n575), .A4(n287), .S0(n314), 
        .S1(n310), .Y(n479) );
  AOI21X1_HVT U127 ( .A1(n313), .A2(n475), .A3(n347), .Y(n476) );
  NAND2X0_HVT U129 ( .A1(n313), .A2(n305), .Y(n473) );
  MUX41X1_HVT U130 ( .A1(n473), .A3(n474), .A2(n477), .A4(n476), .S0(n316), 
        .S1(n319), .Y(n472) );
  AND2X1_HVT U131 ( .A1(n273), .A2(n230), .Y(n471) );
  MUX41X1_HVT U132 ( .A1(n344), .A3(n471), .A2(n388), .A4(n353), .S0(n315), 
        .S1(n308), .Y(n470) );
  MUX41X1_HVT U133 ( .A1(n389), .A3(n346), .A2(n544), .A4(n345), .S0(n314), 
        .S1(n307), .Y(n469) );
  MUX41X1_HVT U136 ( .A1(n549), .A3(n501), .A2(n467), .A4(n351), .S0(n331), 
        .S1(n334), .Y(n466) );
  MUX41X1_HVT U137 ( .A1(n591), .A3(n569), .A2(n241), .A4(n382), .S0(n316), 
        .S1(n307), .Y(n465) );
  MUX41X1_HVT U139 ( .A1(n464), .A3(n468), .A2(n472), .A4(n478), .S0(n321), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n368), .A3(n296), .A2(n361), .A4(n587), .S0(n315), 
        .S1(n309), .Y(n463) );
  NAND2X0_HVT U141 ( .A1(n285), .A2(n330), .Y(n462) );
  MUX41X1_HVT U142 ( .A1(n462), .A3(n559), .A2(n387), .A4(n361), .S0(n313), 
        .S1(n245), .Y(n461) );
  MUX41X1_HVT U145 ( .A1(n567), .A3(n385), .A2(n459), .A4(n519), .S0(n313), 
        .S1(n245), .Y(n458) );
  MUX41X1_HVT U146 ( .A1(n458), .A3(n460), .A2(n461), .A4(n463), .S0(n248), 
        .S1(n321), .Y(n457) );
  AO21X1_HVT U148 ( .A1(n316), .A2(n348), .A3(n262), .Y(n455) );
  MUX41X1_HVT U151 ( .A1(n292), .A3(n370), .A2(n360), .A4(n453), .S0(n314), 
        .S1(n307), .Y(n452) );
  MUX41X1_HVT U155 ( .A1(n361), .A3(n587), .A2(n579), .A4(n223), .S0(n309), 
        .S1(n333), .Y(n448) );
  MUX41X1_HVT U156 ( .A1(n448), .A3(n452), .A2(n449), .A4(n454), .S0(in[5]), 
        .S1(n319), .Y(n447) );
  NAND2X0_HVT U159 ( .A1(n444), .A2(n443), .Y(n445) );
  MUX41X1_HVT U162 ( .A1(n372), .A3(n358), .A2(n563), .A4(n441), .S0(n309), 
        .S1(n244), .Y(n440) );
  NAND2X0_HVT U163 ( .A1(n252), .A2(n270), .Y(n439) );
  MUX41X1_HVT U164 ( .A1(n590), .A3(n439), .A2(n561), .A4(n359), .S0(n310), 
        .S1(n244), .Y(n438) );
  NAND2X0_HVT U166 ( .A1(n588), .A2(n435), .Y(n436) );
  MUX41X1_HVT U168 ( .A1(n434), .A3(n440), .A2(n438), .A4(n442), .S0(n321), 
        .S1(n319), .Y(n433) );
  NAND2X0_HVT U177 ( .A1(n326), .A2(n258), .Y(n425) );
  AND2X1_HVT U179 ( .A1(n593), .A2(n268), .Y(n423) );
  MUX41X1_HVT U182 ( .A1(n346), .A3(n265), .A2(n343), .A4(n292), .S0(n310), 
        .S1(n333), .Y(n420) );
  MUX41X1_HVT U183 ( .A1(n232), .A3(n376), .A2(n359), .A4(n556), .S0(n314), 
        .S1(n308), .Y(n419) );
  AND2X1_HVT U185 ( .A1(n286), .A2(n230), .Y(n417) );
  NAND2X0_HVT U191 ( .A1(n337), .A2(n352), .Y(n411) );
  AND2X1_HVT U192 ( .A1(n369), .A2(n409), .Y(n410) );
  NAND2X0_HVT U194 ( .A1(n556), .A2(n409), .Y(n407) );
  MUX41X1_HVT U195 ( .A1(n408), .A3(n407), .A2(n410), .A4(n411), .S0(n311), 
        .S1(n248), .Y(n406) );
  NAND2X0_HVT U198 ( .A1(n229), .A2(n291), .Y(n588) );
  NAND2X0_HVT U200 ( .A1(n267), .A2(n330), .Y(n475) );
  NAND2X0_HVT U207 ( .A1(n330), .A2(n303), .Y(n539) );
  OA21X2_HVT U2 ( .A1(n337), .A2(n548), .A3(n364), .Y(n546) );
  NAND2X0_HVT U3 ( .A1(n417), .A2(n6), .Y(n58) );
  NAND2X0_HVT U4 ( .A1(n379), .A2(n314), .Y(n196) );
  NAND2X0_HVT U14 ( .A1(n58), .A2(n196), .Y(n416) );
  IBUFFX2_HVT U16 ( .A(n314), .Y(n6) );
  INVX0_HVT U17 ( .A(n577), .Y(n359) );
  INVX1_HVT U18 ( .A(n336), .Y(n335) );
  IBUFFX2_HVT U20 ( .A(n336), .Y(n244) );
  MUX21X1_HVT U21 ( .A1(n303), .A2(n318), .S0(n251), .Y(n430) );
  MUX21X1_HVT U22 ( .A1(n261), .A2(n339), .S0(n316), .Y(n525) );
  INVX1_HVT U23 ( .A(n286), .Y(n284) );
  AO21X2_HVT U24 ( .A1(n327), .A2(n262), .A3(n336), .Y(n409) );
  AO21X2_HVT U25 ( .A1(n230), .A2(n306), .A3(n336), .Y(n443) );
  MUX41X1_HVT U26 ( .A1(n430), .A3(n512), .A2(n576), .A4(n294), .S0(n197), 
        .S1(n245), .Y(n429) );
  IBUFFX16_HVT U27 ( .A(n308), .Y(n197) );
  MUX21X1_HVT U28 ( .A1(n490), .A2(n491), .S0(n313), .Y(n489) );
  INVX1_HVT U29 ( .A(in[3]), .Y(n257) );
  INVX2_HVT U30 ( .A(n306), .Y(n302) );
  IBUFFX2_HVT U31 ( .A(n336), .Y(n245) );
  IBUFFX2_HVT U33 ( .A(n336), .Y(n333) );
  INVX1_HVT U34 ( .A(n393), .Y(n389) );
  INVX0_HVT U36 ( .A(n277), .Y(n263) );
  INVX1_HVT U37 ( .A(n277), .Y(n266) );
  NAND2X1_HVT U39 ( .A1(n257), .A2(n392), .Y(n597) );
  MUX21X2_HVT U40 ( .A1(n546), .A2(n547), .S0(n198), .Y(n545) );
  IBUFFX16_HVT U41 ( .A(n308), .Y(n198) );
  MUX21X2_HVT U43 ( .A1(n322), .A2(n510), .S0(n199), .Y(n509) );
  IBUFFX16_HVT U44 ( .A(n327), .Y(n199) );
  MUX21X2_HVT U45 ( .A1(n426), .A2(n433), .S0(n200), .Y(out[6]) );
  IBUFFX16_HVT U46 ( .A(n254), .Y(n200) );
  MUX41X1_HVT U47 ( .A1(n412), .A3(n406), .A2(n421), .A4(n418), .S0(n320), 
        .S1(n201), .Y(out[7]) );
  IBUFFX16_HVT U48 ( .A(n254), .Y(n201) );
  MUX21X2_HVT U49 ( .A1(n363), .A2(n354), .S0(n316), .Y(n547) );
  MUX21X1_HVT U50 ( .A1(n277), .A2(n318), .S0(n202), .Y(n572) );
  IBUFFX16_HVT U51 ( .A(n325), .Y(n202) );
  MUX41X1_HVT U52 ( .A1(n413), .A3(n416), .A2(n414), .A4(n415), .S0(n248), 
        .S1(n206), .Y(n412) );
  IBUFFX16_HVT U53 ( .A(n308), .Y(n206) );
  MUX21X2_HVT U54 ( .A1(n522), .A2(n515), .S0(n208), .Y(out[1]) );
  IBUFFX16_HVT U56 ( .A(in[7]), .Y(n208) );
  MUX21X1_HVT U57 ( .A1(n557), .A2(n378), .S0(n283), .Y(n414) );
  IBUFFX16_HVT U58 ( .A(n249), .Y(n319) );
  NBUFFX4_HVT U59 ( .A(n392), .Y(n318) );
  NAND2X0_HVT U61 ( .A1(n373), .A2(n218), .Y(n219) );
  NAND2X0_HVT U63 ( .A1(n297), .A2(n314), .Y(n220) );
  NAND2X0_HVT U64 ( .A1(n219), .A2(n220), .Y(n408) );
  IBUFFX2_HVT U68 ( .A(n314), .Y(n218) );
  MUX21X1_HVT U69 ( .A1(n318), .A2(n317), .S0(n221), .Y(n553) );
  IBUFFX16_HVT U70 ( .A(n324), .Y(n221) );
  INVX2_HVT U75 ( .A(in[6]), .Y(n392) );
  MUX21X2_HVT U76 ( .A1(n436), .A2(n437), .S0(n313), .Y(n434) );
  IBUFFX2_HVT U77 ( .A(n572), .Y(n362) );
  INVX0_HVT U78 ( .A(n363), .Y(n222) );
  INVX0_HVT U79 ( .A(n222), .Y(n223) );
  NAND2X0_HVT U86 ( .A1(n258), .A2(n224), .Y(n225) );
  NAND2X0_HVT U87 ( .A1(n318), .A2(n227), .Y(n226) );
  NAND2X0_HVT U90 ( .A1(n225), .A2(n226), .Y(n571) );
  INVX0_HVT U91 ( .A(n227), .Y(n224) );
  IBUFFX2_HVT U92 ( .A(n328), .Y(n227) );
  INVX0_HVT U93 ( .A(n571), .Y(n363) );
  INVX2_HVT U94 ( .A(n249), .Y(n248) );
  INVX2_HVT U97 ( .A(n336), .Y(n334) );
  INVX1_HVT U103 ( .A(in[4]), .Y(n336) );
  MUX21X1_HVT U106 ( .A1(n481), .A2(n479), .S0(n249), .Y(n478) );
  IBUFFX16_HVT U111 ( .A(in[1]), .Y(n249) );
  INVX0_HVT U113 ( .A(n392), .Y(n272) );
  NBUFFX2_HVT U117 ( .A(n337), .Y(n228) );
  INVX1_HVT U121 ( .A(in[4]), .Y(n337) );
  MUX21X2_HVT U123 ( .A1(n469), .A2(n470), .S0(n319), .Y(n468) );
  AO21X1_HVT U125 ( .A1(n285), .A2(n595), .A3(n337), .Y(n435) );
  OA21X1_HVT U126 ( .A1(n341), .A2(n228), .A3(n350), .Y(n450) );
  INVX1_HVT U128 ( .A(n293), .Y(n229) );
  INVX1_HVT U134 ( .A(n253), .Y(n230) );
  INVX1_HVT U135 ( .A(n325), .Y(n293) );
  NBUFFX2_HVT U138 ( .A(in[0]), .Y(n253) );
  MUX21X2_HVT U143 ( .A1(n347), .A2(n557), .S0(n316), .Y(n491) );
  OA21X1_HVT U144 ( .A1(n365), .A2(n337), .A3(n539), .Y(n413) );
  MUX41X1_HVT U147 ( .A1(n294), .A3(n298), .A2(n432), .A4(n297), .S0(n231), 
        .S1(n334), .Y(n431) );
  IBUFFX16_HVT U149 ( .A(n307), .Y(n231) );
  MUX21X2_HVT U150 ( .A1(n349), .A2(n582), .S0(n316), .Y(n508) );
  OA21X1_HVT U152 ( .A1(n342), .A2(n337), .A3(n577), .Y(n524) );
  MUX21X1_HVT U153 ( .A1(n299), .A2(n241), .S0(n283), .Y(n451) );
  MUX21X1_HVT U154 ( .A1(n287), .A2(n544), .S0(n315), .Y(n541) );
  INVX1_HVT U157 ( .A(n235), .Y(n542) );
  MUX21X1_HVT U158 ( .A1(n574), .A2(n234), .S0(n300), .Y(n235) );
  MUX21X1_HVT U160 ( .A1(n359), .A2(n536), .S0(n300), .Y(n535) );
  MUX21X1_HVT U161 ( .A1(n360), .A2(n265), .S0(n331), .Y(n536) );
  INVX1_HVT U165 ( .A(n331), .Y(n250) );
  INVX0_HVT U167 ( .A(n267), .Y(n270) );
  INVX1_HVT U169 ( .A(n312), .Y(n247) );
  INVX1_HVT U170 ( .A(in[5]), .Y(n320) );
  INVX1_HVT U171 ( .A(in[7]), .Y(n254) );
  INVX0_HVT U172 ( .A(n317), .Y(n233) );
  INVX1_HVT U173 ( .A(n301), .Y(n303) );
  INVX1_HVT U174 ( .A(n304), .Y(n306) );
  INVX1_HVT U175 ( .A(n598), .Y(n304) );
  INVX0_HVT U176 ( .A(n288), .Y(n291) );
  INVX1_HVT U178 ( .A(n582), .Y(n286) );
  INVX1_HVT U180 ( .A(n263), .Y(n262) );
  INVX0_HVT U181 ( .A(n316), .Y(n246) );
  MUX21X2_HVT U184 ( .A1(n508), .A2(n509), .S0(n307), .Y(n507) );
  INVX1_HVT U186 ( .A(n569), .Y(n365) );
  INVX0_HVT U187 ( .A(n232), .Y(n555) );
  MUX21X1_HVT U188 ( .A1(n233), .A2(n323), .S0(n326), .Y(n232) );
  INVX1_HVT U189 ( .A(n329), .Y(n251) );
  IBUFFX2_HVT U190 ( .A(n329), .Y(n324) );
  IBUFFX2_HVT U193 ( .A(n230), .Y(n325) );
  IBUFFX2_HVT U196 ( .A(n329), .Y(n327) );
  INVX1_HVT U197 ( .A(in[0]), .Y(n329) );
  INVX2_HVT U199 ( .A(n253), .Y(n330) );
  MUX21X2_HVT U201 ( .A1(n450), .A2(n451), .S0(n313), .Y(n449) );
  MUX21X1_HVT U202 ( .A1(n344), .A2(n573), .S0(n250), .Y(n234) );
  INVX0_HVT U203 ( .A(n573), .Y(n361) );
  NAND2X0_HVT U204 ( .A1(n422), .A2(n249), .Y(n236) );
  NAND2X0_HVT U205 ( .A1(n424), .A2(n248), .Y(n237) );
  NAND2X0_HVT U206 ( .A1(n236), .A2(n237), .Y(n421) );
  MUX21X1_HVT U208 ( .A1(n272), .A2(n582), .S0(n253), .Y(n264) );
  MUX21X2_HVT U209 ( .A1(n506), .A2(n499), .S0(n254), .Y(out[2]) );
  MUX21X2_HVT U210 ( .A1(n524), .A2(n525), .S0(n250), .Y(n523) );
  NAND2X0_HVT U211 ( .A1(n550), .A2(n238), .Y(n239) );
  NAND2X0_HVT U212 ( .A1(n299), .A2(n246), .Y(n240) );
  NAND2X0_HVT U213 ( .A1(n239), .A2(n240), .Y(n415) );
  INVX1_HVT U214 ( .A(n246), .Y(n238) );
  XOR2X1_HVT U215 ( .A1(n269), .A2(n251), .Y(n550) );
  MUX41X1_HVT U216 ( .A1(n562), .A3(n266), .A2(n302), .A4(n305), .S0(n247), 
        .S1(n246), .Y(n428) );
  INVX0_HVT U217 ( .A(n264), .Y(n562) );
  MUX41X1_HVT U218 ( .A1(n338), .A3(n566), .A2(n553), .A4(n423), .S0(n247), 
        .S1(n245), .Y(n422) );
  NAND2X0_HVT U219 ( .A1(n274), .A2(n275), .Y(n241) );
  NAND2X0_HVT U220 ( .A1(n419), .A2(n249), .Y(n242) );
  NAND2X0_HVT U221 ( .A1(n420), .A2(in[1]), .Y(n243) );
  NAND2X0_HVT U222 ( .A1(n242), .A2(n243), .Y(n418) );
  MUX41X1_HVT U223 ( .A1(n544), .A3(n362), .A2(n284), .A4(n376), .S0(n247), 
        .S1(n283), .Y(n543) );
  INVX1_HVT U224 ( .A(n315), .Y(n283) );
  MUX41X1_HVT U225 ( .A1(n580), .A3(n365), .A2(n581), .A4(n367), .S0(n247), 
        .S1(n244), .Y(n521) );
  MUX41X1_HVT U226 ( .A1(n529), .A3(n526), .A2(n527), .A4(n523), .S0(n320), 
        .S1(n249), .Y(n522) );
  MUX21X1_HVT U227 ( .A1(n597), .A2(n257), .S0(n253), .Y(n287) );
  MUX21X2_HVT U228 ( .A1(n540), .A2(n541), .S0(n250), .Y(n538) );
  INVX0_HVT U229 ( .A(n287), .Y(n575) );
  MUX41X1_HVT U230 ( .A1(n512), .A3(n551), .A2(n592), .A4(n304), .S0(n247), 
        .S1(n228), .Y(n511) );
  INVX0_HVT U231 ( .A(n329), .Y(n252) );
  IBUFFX2_HVT U232 ( .A(n329), .Y(n328) );
  INVX1_HVT U233 ( .A(n402), .Y(n379) );
  MUX41X1_HVT U234 ( .A1(n431), .A3(n428), .A2(n429), .A4(n427), .S0(n320), 
        .S1(n249), .Y(n426) );
  MUX21X1_HVT U235 ( .A1(n286), .A2(n262), .S0(n328), .Y(n576) );
  MUX21X1_HVT U236 ( .A1(n270), .A2(n302), .S0(n327), .Y(n554) );
  INVX0_HVT U237 ( .A(n282), .Y(n559) );
  MUX21X1_HVT U238 ( .A1(n273), .A2(n391), .S0(n326), .Y(n557) );
  INVX0_HVT U239 ( .A(n392), .Y(n273) );
  MUX21X1_HVT U240 ( .A1(n582), .A2(n318), .S0(n315), .Y(n510) );
  INVX1_HVT U241 ( .A(n320), .Y(n321) );
  INVX0_HVT U242 ( .A(n255), .Y(n531) );
  INVX0_HVT U243 ( .A(n354), .Y(n256) );
  INVX0_HVT U244 ( .A(n268), .Y(n271) );
  INVX1_HVT U245 ( .A(n291), .Y(n285) );
  MUX41X1_HVT U246 ( .A1(n256), .A3(n303), .A2(n584), .A4(n257), .S0(n311), 
        .S1(n228), .Y(n255) );
  MUX21X2_HVT U247 ( .A1(n530), .A2(n537), .S0(in[7]), .Y(out[0]) );
  MUX21X2_HVT U248 ( .A1(n482), .A2(n492), .S0(in[7]), .Y(out[3]) );
  MUX41X1_HVT U249 ( .A1(n362), .A3(n381), .A2(n299), .A4(n343), .S0(n250), 
        .S1(n337), .Y(n514) );
  INVX1_HVT U250 ( .A(n257), .Y(n258) );
  MUX21X2_HVT U251 ( .A1(n445), .A2(n446), .S0(n313), .Y(n442) );
  NAND2X0_HVT U252 ( .A1(n261), .A2(n335), .Y(n259) );
  NAND2X0_HVT U253 ( .A1(n555), .A2(n283), .Y(n260) );
  NAND2X0_HVT U254 ( .A1(n259), .A2(n260), .Y(n446) );
  INVX0_HVT U255 ( .A(in[3]), .Y(n390) );
  MUX21X1_HVT U256 ( .A1(n233), .A2(n596), .S0(n230), .Y(n261) );
  INVX1_HVT U257 ( .A(n596), .Y(n391) );
  OR2X1_HVT U258 ( .A1(n390), .A2(n392), .Y(n596) );
  INVX1_HVT U259 ( .A(n597), .Y(n277) );
  INVX1_HVT U260 ( .A(n343), .Y(n265) );
  INVX1_HVT U261 ( .A(n595), .Y(n343) );
  NAND2X0_HVT U262 ( .A1(n328), .A2(n266), .Y(n595) );
  MUX41X1_HVT U263 ( .A1(n544), .A3(n381), .A2(n286), .A4(n389), .S0(n250), 
        .S1(n335), .Y(n427) );
  XNOR2X1_HVT U264 ( .A1(n392), .A2(n390), .Y(n582) );
  INVX0_HVT U265 ( .A(n576), .Y(n360) );
  NAND2X0_HVT U266 ( .A1(n272), .A2(n317), .Y(n267) );
  NAND2X0_HVT U267 ( .A1(n272), .A2(n317), .Y(n268) );
  INVX0_HVT U268 ( .A(n271), .Y(n269) );
  MUX41X1_HVT U269 ( .A1(n554), .A3(n425), .A2(n303), .A4(n298), .S0(n283), 
        .S1(n247), .Y(n424) );
  INVX1_HVT U270 ( .A(n554), .Y(n372) );
  INVX1_HVT U271 ( .A(n276), .Y(n292) );
  MUX41X1_HVT U272 ( .A1(n535), .A3(n532), .A2(n534), .A4(n531), .S0(n320), 
        .S1(n249), .Y(n530) );
  MUX21X1_HVT U273 ( .A1(n284), .A2(n317), .S0(n324), .Y(n577) );
  NAND2X0_HVT U274 ( .A1(n318), .A2(n251), .Y(n274) );
  NAND2X0_HVT U275 ( .A1(n284), .A2(n330), .Y(n275) );
  NAND2X0_HVT U276 ( .A1(n274), .A2(n275), .Y(n573) );
  MUX21X1_HVT U277 ( .A1(n291), .A2(n257), .S0(n293), .Y(n276) );
  NAND2X0_HVT U278 ( .A1(n455), .A2(n307), .Y(n278) );
  NAND2X0_HVT U279 ( .A1(n456), .A2(n250), .Y(n279) );
  NAND2X0_HVT U280 ( .A1(n278), .A2(n279), .Y(n454) );
  NAND2X0_HVT U281 ( .A1(n447), .A2(n254), .Y(n280) );
  NAND2X0_HVT U282 ( .A1(n457), .A2(in[7]), .Y(n281) );
  NAND2X0_HVT U283 ( .A1(n280), .A2(n281), .Y(out[5]) );
  MUX21X1_HVT U284 ( .A1(n388), .A2(n344), .S0(n314), .Y(n456) );
  MUX21X1_HVT U285 ( .A1(n233), .A2(n288), .S0(n330), .Y(n282) );
  INVX0_HVT U286 ( .A(n286), .Y(n288) );
  NAND2X0_HVT U287 ( .A1(n572), .A2(n283), .Y(n289) );
  NAND2X0_HVT U288 ( .A1(n575), .A2(n314), .Y(n290) );
  NAND2X0_HVT U289 ( .A1(n289), .A2(n290), .Y(n437) );
  MUX41X1_HVT U290 ( .A1(n575), .A3(n578), .A2(n232), .A4(n270), .S0(n250), 
        .S1(n228), .Y(n460) );
  AND2X1_HVT U291 ( .A1(n593), .A2(n266), .Y(n294) );
  AND2X1_HVT U292 ( .A1(n266), .A2(n583), .Y(n295) );
  MUX21X1_HVT U293 ( .A1(n262), .A2(n286), .S0(n326), .Y(n565) );
  MUX21X1_HVT U294 ( .A1(n318), .A2(n271), .S0(n324), .Y(n453) );
  MUX21X1_HVT U295 ( .A1(n286), .A2(n318), .S0(n326), .Y(n395) );
  MUX21X1_HVT U296 ( .A1(n277), .A2(n318), .S0(n325), .Y(n403) );
  MUX21X1_HVT U297 ( .A1(n267), .A2(n322), .S0(n327), .Y(n441) );
  MUX21X1_HVT U298 ( .A1(n285), .A2(n302), .S0(n324), .Y(n567) );
  MUX21X1_HVT U299 ( .A1(n317), .A2(n277), .S0(n251), .Y(n568) );
  MUX21X1_HVT U300 ( .A1(n262), .A2(n391), .S0(n324), .Y(n548) );
  MUX21X1_HVT U301 ( .A1(n288), .A2(n270), .S0(n251), .Y(n564) );
  MUX21X1_HVT U302 ( .A1(n302), .A2(n288), .S0(n252), .Y(n400) );
  MUX21X1_HVT U303 ( .A1(n269), .A2(n263), .S0(n251), .Y(n394) );
  MUX21X1_HVT U304 ( .A1(n317), .A2(n266), .S0(n325), .Y(n402) );
  MUX21X1_HVT U305 ( .A1(n565), .A2(n295), .S0(n313), .Y(n474) );
  MUX21X1_HVT U306 ( .A1(n303), .A2(n391), .S0(n252), .Y(n432) );
  MUX21X1_HVT U307 ( .A1(n318), .A2(n597), .S0(n327), .Y(n496) );
  MUX21X1_HVT U308 ( .A1(n387), .A2(n296), .S0(n311), .Y(n477) );
  XOR2X1_HVT U309 ( .A1(n306), .A2(n326), .Y(n561) );
  XOR2X1_HVT U310 ( .A1(n284), .A2(n327), .Y(n552) );
  XNOR2X1_HVT U311 ( .A1(n597), .A2(n328), .Y(n296) );
  MUX21X1_HVT U312 ( .A1(n302), .A2(n270), .S0(n326), .Y(n570) );
  MUX21X1_HVT U313 ( .A1(n323), .A2(n266), .S0(n327), .Y(n580) );
  MUX21X1_HVT U314 ( .A1(n318), .A2(n285), .S0(n328), .Y(n558) );
  MUX21X1_HVT U315 ( .A1(n306), .A2(n263), .S0(n252), .Y(n584) );
  MUX21X1_HVT U316 ( .A1(n322), .A2(n257), .S0(n251), .Y(n579) );
  XOR2X1_HVT U317 ( .A1(n323), .A2(n252), .Y(n551) );
  AND2X1_HVT U318 ( .A1(n251), .A2(n318), .Y(n297) );
  MUX21X1_HVT U319 ( .A1(n323), .A2(n318), .S0(n229), .Y(n480) );
  MUX21X1_HVT U320 ( .A1(n317), .A2(n322), .S0(n324), .Y(n397) );
  NBUFFX2_HVT U321 ( .A(n335), .Y(n315) );
  NBUFFX2_HVT U322 ( .A(n335), .Y(n314) );
  NBUFFX2_HVT U323 ( .A(n335), .Y(n316) );
  AND2X1_HVT U324 ( .A1(n391), .A2(n330), .Y(n298) );
  MUX21X1_HVT U325 ( .A1(n263), .A2(n268), .S0(n229), .Y(n459) );
  AND2X1_HVT U326 ( .A1(n323), .A2(n330), .Y(n299) );
  NBUFFX2_HVT U327 ( .A(n596), .Y(n323) );
  NBUFFX2_HVT U328 ( .A(n596), .Y(n322) );
  NBUFFX2_HVT U329 ( .A(n390), .Y(n317) );
  INVX1_HVT U330 ( .A(n329), .Y(n326) );
  NBUFFX2_HVT U331 ( .A(n332), .Y(n313) );
  XNOR2X1_HVT U332 ( .A1(n337), .A2(n310), .Y(n300) );
  NBUFFX2_HVT U333 ( .A(n332), .Y(n310) );
  NBUFFX2_HVT U334 ( .A(n332), .Y(n311) );
  NBUFFX2_HVT U335 ( .A(n332), .Y(n312) );
  NBUFFX2_HVT U336 ( .A(n331), .Y(n308) );
  NBUFFX2_HVT U337 ( .A(n331), .Y(n309) );
  NBUFFX2_HVT U338 ( .A(n331), .Y(n307) );
  MUX21X1_HVT U339 ( .A1(n465), .A2(n466), .S0(in[1]), .Y(n464) );
  MUX21X1_HVT U340 ( .A1(n273), .A2(n270), .S0(n325), .Y(n405) );
  MUX21X1_HVT U341 ( .A1(n273), .A2(n301), .S0(n327), .Y(n581) );
  MUX21X1_HVT U342 ( .A1(n305), .A2(n258), .S0(n252), .Y(n444) );
  MUX21X1_HVT U343 ( .A1(n267), .A2(n258), .S0(n324), .Y(n504) );
  XOR2X1_HVT U344 ( .A1(n328), .A2(n273), .Y(n549) );
  MUX21X1_HVT U345 ( .A1(n262), .A2(n273), .S0(n252), .Y(n467) );
  MUX21X1_HVT U346 ( .A1(n258), .A2(n306), .S0(n327), .Y(n399) );
  MUX21X1_HVT U347 ( .A1(n302), .A2(n258), .S0(n328), .Y(n393) );
  MUX21X1_HVT U348 ( .A1(n268), .A2(n273), .S0(n252), .Y(n569) );
  MUX21X1_HVT U349 ( .A1(n273), .A2(n302), .S0(n324), .Y(n574) );
  MUX21X1_HVT U350 ( .A1(n391), .A2(n271), .S0(n326), .Y(n485) );
  MUX21X1_HVT U351 ( .A1(n258), .A2(n267), .S0(n229), .Y(n398) );
  MUX21X1_HVT U352 ( .A1(n273), .A2(n323), .S0(n328), .Y(n404) );
  MUX21X1_HVT U353 ( .A1(n322), .A2(n273), .S0(n251), .Y(n401) );
  MUX21X1_HVT U354 ( .A1(n317), .A2(n273), .S0(n324), .Y(n396) );
  NBUFFX2_HVT U355 ( .A(in[2]), .Y(n332) );
  NBUFFX2_HVT U356 ( .A(in[2]), .Y(n331) );
  INVX0_HVT U357 ( .A(n304), .Y(n301) );
  INVX0_HVT U358 ( .A(n304), .Y(n305) );
  INVX0_HVT U359 ( .A(n587), .Y(n338) );
  INVX0_HVT U360 ( .A(n566), .Y(n339) );
  INVX0_HVT U361 ( .A(n560), .Y(n340) );
  INVX0_HVT U362 ( .A(n501), .Y(n341) );
  INVX0_HVT U363 ( .A(n462), .Y(n342) );
  INVX0_HVT U364 ( .A(n594), .Y(n344) );
  INVX0_HVT U365 ( .A(n593), .Y(n345) );
  INVX0_HVT U366 ( .A(n556), .Y(n346) );
  INVX0_HVT U367 ( .A(n592), .Y(n347) );
  INVX0_HVT U368 ( .A(n591), .Y(n348) );
  INVX0_HVT U369 ( .A(n563), .Y(n349) );
  INVX0_HVT U370 ( .A(n585), .Y(n350) );
  INVX0_HVT U371 ( .A(n590), .Y(n351) );
  INVX0_HVT U372 ( .A(n586), .Y(n352) );
  INVX0_HVT U373 ( .A(n584), .Y(n353) );
  INVX0_HVT U374 ( .A(n583), .Y(n354) );
  INVX0_HVT U375 ( .A(n581), .Y(n355) );
  INVX0_HVT U376 ( .A(n580), .Y(n356) );
  INVX0_HVT U377 ( .A(n579), .Y(n357) );
  INVX0_HVT U378 ( .A(n578), .Y(n358) );
  INVX0_HVT U379 ( .A(n570), .Y(n364) );
  INVX0_HVT U380 ( .A(n568), .Y(n366) );
  INVX0_HVT U381 ( .A(n567), .Y(n367) );
  INVX0_HVT U382 ( .A(n565), .Y(n368) );
  INVX0_HVT U383 ( .A(n564), .Y(n369) );
  INVX0_HVT U384 ( .A(n561), .Y(n370) );
  INVX0_HVT U385 ( .A(n558), .Y(n371) );
  INVX0_HVT U386 ( .A(n553), .Y(n373) );
  INVX0_HVT U387 ( .A(n552), .Y(n374) );
  INVX0_HVT U388 ( .A(n589), .Y(n375) );
  INVX0_HVT U389 ( .A(n405), .Y(n376) );
  INVX0_HVT U390 ( .A(n404), .Y(n377) );
  INVX0_HVT U391 ( .A(n403), .Y(n378) );
  INVX0_HVT U392 ( .A(n401), .Y(n380) );
  INVX0_HVT U393 ( .A(n400), .Y(n381) );
  INVX0_HVT U394 ( .A(n399), .Y(n382) );
  INVX0_HVT U395 ( .A(n398), .Y(n383) );
  INVX0_HVT U396 ( .A(n397), .Y(n384) );
  INVX0_HVT U397 ( .A(n396), .Y(n385) );
  INVX0_HVT U398 ( .A(n444), .Y(n386) );
  INVX0_HVT U399 ( .A(n395), .Y(n387) );
  INVX0_HVT U400 ( .A(n394), .Y(n388) );
endmodule

