
module add_round_keys_0 ( state, subkey, out );
  input [127:0] state;
  input [127:0] subkey;
  output [127:0] out;


  XOR2X1_HVT U1 ( .A1(subkey[60]), .A2(state[60]), .Y(out[60]) );
  XOR2X1_HVT U2 ( .A1(subkey[113]), .A2(state[113]), .Y(out[113]) );
  XOR2X1_HVT U3 ( .A1(subkey[111]), .A2(state[111]), .Y(out[111]) );
  XOR2X1_HVT U4 ( .A1(subkey[121]), .A2(state[121]), .Y(out[121]) );
  XOR2X1_HVT U5 ( .A1(subkey[100]), .A2(state[100]), .Y(out[100]) );
  XOR2X1_HVT U6 ( .A1(subkey[116]), .A2(state[116]), .Y(out[116]) );
  XOR2X1_HVT U7 ( .A1(subkey[20]), .A2(state[20]), .Y(out[20]) );
  XOR2X1_HVT U8 ( .A1(subkey[19]), .A2(state[19]), .Y(out[19]) );
  XOR2X1_HVT U9 ( .A1(subkey[36]), .A2(state[36]), .Y(out[36]) );
  XOR2X1_HVT U10 ( .A1(subkey[67]), .A2(state[67]), .Y(out[67]) );
  XOR2X1_HVT U11 ( .A1(subkey[68]), .A2(state[68]), .Y(out[68]) );
  XOR2X1_HVT U12 ( .A1(subkey[51]), .A2(state[51]), .Y(out[51]) );
  XOR2X1_HVT U13 ( .A1(subkey[17]), .A2(state[17]), .Y(out[17]) );
  XOR2X1_HVT U14 ( .A1(subkey[43]), .A2(state[43]), .Y(out[43]) );
  XOR2X1_HVT U15 ( .A1(subkey[59]), .A2(state[59]), .Y(out[59]) );
  XOR2X1_HVT U16 ( .A1(subkey[73]), .A2(state[73]), .Y(out[73]) );
  XOR2X1_HVT U17 ( .A1(subkey[105]), .A2(state[105]), .Y(out[105]) );
  XOR2X1_HVT U18 ( .A1(subkey[65]), .A2(state[65]), .Y(out[65]) );
  XOR2X1_HVT U19 ( .A1(subkey[33]), .A2(state[33]), .Y(out[33]) );
  XOR2X1_HVT U20 ( .A1(subkey[41]), .A2(state[41]), .Y(out[41]) );
  XOR2X1_HVT U21 ( .A1(subkey[57]), .A2(state[57]), .Y(out[57]) );
  XOR2X1_HVT U22 ( .A1(subkey[89]), .A2(state[89]), .Y(out[89]) );
  XOR2X1_HVT U23 ( .A1(subkey[99]), .A2(state[99]), .Y(out[99]) );
  XOR2X1_HVT U24 ( .A1(subkey[16]), .A2(state[16]), .Y(out[16]) );
  XOR2X1_HVT U25 ( .A1(subkey[81]), .A2(state[81]), .Y(out[81]) );
  XOR2X1_HVT U26 ( .A1(subkey[4]), .A2(state[4]), .Y(out[4]) );
  XOR2X1_HVT U27 ( .A1(subkey[49]), .A2(state[49]), .Y(out[49]) );
  XOR2X1_HVT U28 ( .A1(subkey[9]), .A2(state[9]), .Y(out[9]) );
  XOR2X1_HVT U29 ( .A1(subkey[1]), .A2(state[1]), .Y(out[1]) );
  XOR2X1_HVT U30 ( .A1(subkey[103]), .A2(state[103]), .Y(out[103]) );
  XOR2X1_HVT U31 ( .A1(subkey[97]), .A2(state[97]), .Y(out[97]) );
  XOR2X1_HVT U32 ( .A1(subkey[12]), .A2(state[12]), .Y(out[12]) );
  XOR2X1_HVT U33 ( .A1(subkey[28]), .A2(state[28]), .Y(out[28]) );
  XOR2X1_HVT U34 ( .A1(subkey[79]), .A2(state[79]), .Y(out[79]) );
  XOR2X1_HVT U35 ( .A1(subkey[47]), .A2(state[47]), .Y(out[47]) );
  XOR2X1_HVT U36 ( .A1(subkey[31]), .A2(state[31]), .Y(out[31]) );
  XOR2X1_HVT U37 ( .A1(subkey[25]), .A2(state[25]), .Y(out[25]) );
  XOR2X1_HVT U38 ( .A1(subkey[123]), .A2(state[123]), .Y(out[123]) );
  XOR2X1_HVT U39 ( .A1(subkey[3]), .A2(state[3]), .Y(out[3]) );
  XOR2X1_HVT U40 ( .A1(subkey[71]), .A2(state[71]), .Y(out[71]) );
  XOR2X1_HVT U41 ( .A1(subkey[24]), .A2(state[24]), .Y(out[24]) );
  XOR2X1_HVT U42 ( .A1(subkey[75]), .A2(state[75]), .Y(out[75]) );
  XOR2X1_HVT U43 ( .A1(subkey[124]), .A2(state[124]), .Y(out[124]) );
  XOR2X1_HVT U44 ( .A1(subkey[84]), .A2(state[84]), .Y(out[84]) );
  XOR2X1_HVT U45 ( .A1(subkey[39]), .A2(state[39]), .Y(out[39]) );
  XOR2X1_HVT U46 ( .A1(subkey[27]), .A2(state[27]), .Y(out[27]) );
  XOR2X1_HVT U47 ( .A1(subkey[76]), .A2(state[76]), .Y(out[76]) );
  XOR2X1_HVT U48 ( .A1(subkey[48]), .A2(state[48]), .Y(out[48]) );
  XOR2X1_HVT U49 ( .A1(subkey[52]), .A2(state[52]), .Y(out[52]) );
  XOR2X1_HVT U50 ( .A1(subkey[92]), .A2(state[92]), .Y(out[92]) );
  XOR2X1_HVT U51 ( .A1(subkey[112]), .A2(state[112]), .Y(out[112]) );
  XOR2X1_HVT U52 ( .A1(subkey[127]), .A2(state[127]), .Y(out[127]) );
  XOR2X1_HVT U53 ( .A1(subkey[119]), .A2(state[119]), .Y(out[119]) );
  XOR2X1_HVT U54 ( .A1(subkey[55]), .A2(state[55]), .Y(out[55]) );
  XOR2X1_HVT U55 ( .A1(subkey[87]), .A2(state[87]), .Y(out[87]) );
  XOR2X1_HVT U56 ( .A1(subkey[56]), .A2(state[56]), .Y(out[56]) );
  XOR2X1_HVT U57 ( .A1(subkey[88]), .A2(state[88]), .Y(out[88]) );
  XOR2X1_HVT U58 ( .A1(subkey[108]), .A2(state[108]), .Y(out[108]) );
  XOR2X1_HVT U59 ( .A1(subkey[35]), .A2(state[35]), .Y(out[35]) );
  XOR2X1_HVT U60 ( .A1(subkey[44]), .A2(state[44]), .Y(out[44]) );
  XOR2X1_HVT U61 ( .A1(subkey[83]), .A2(state[83]), .Y(out[83]) );
  XOR2X1_HVT U62 ( .A1(subkey[115]), .A2(state[115]), .Y(out[115]) );
  XOR2X1_HVT U63 ( .A1(subkey[11]), .A2(state[11]), .Y(out[11]) );
  XOR2X1_HVT U64 ( .A1(subkey[120]), .A2(state[120]), .Y(out[120]) );
  XOR2X1_HVT U65 ( .A1(subkey[91]), .A2(state[91]), .Y(out[91]) );
  XOR2X1_HVT U66 ( .A1(subkey[63]), .A2(state[63]), .Y(out[63]) );
  XOR2X1_HVT U67 ( .A1(subkey[95]), .A2(state[95]), .Y(out[95]) );
  XOR2X1_HVT U68 ( .A1(subkey[45]), .A2(state[45]), .Y(out[45]) );
  XOR2X1_HVT U69 ( .A1(subkey[107]), .A2(state[107]), .Y(out[107]) );
  XOR2X1_HVT U70 ( .A1(subkey[0]), .A2(state[0]), .Y(out[0]) );
  XOR2X1_HVT U71 ( .A1(subkey[62]), .A2(state[62]), .Y(out[62]) );
  XOR2X1_HVT U72 ( .A1(subkey[94]), .A2(state[94]), .Y(out[94]) );
  XOR2X1_HVT U73 ( .A1(subkey[30]), .A2(state[30]), .Y(out[30]) );
  XOR2X1_HVT U74 ( .A1(subkey[15]), .A2(state[15]), .Y(out[15]) );
  XOR2X1_HVT U75 ( .A1(subkey[23]), .A2(state[23]), .Y(out[23]) );
  XOR2X1_HVT U76 ( .A1(subkey[104]), .A2(state[104]), .Y(out[104]) );
  XOR2X1_HVT U77 ( .A1(subkey[13]), .A2(state[13]), .Y(out[13]) );
  XOR2X1_HVT U78 ( .A1(subkey[98]), .A2(state[98]), .Y(out[98]) );
  XOR2X1_HVT U79 ( .A1(subkey[109]), .A2(state[109]), .Y(out[109]) );
  XOR2X1_HVT U80 ( .A1(subkey[53]), .A2(state[53]), .Y(out[53]) );
  XOR2X1_HVT U81 ( .A1(subkey[18]), .A2(state[18]), .Y(out[18]) );
  XOR2X1_HVT U82 ( .A1(subkey[69]), .A2(state[69]), .Y(out[69]) );
  XOR2X1_HVT U83 ( .A1(subkey[117]), .A2(state[117]), .Y(out[117]) );
  XOR2X1_HVT U84 ( .A1(subkey[101]), .A2(state[101]), .Y(out[101]) );
  XOR2X1_HVT U85 ( .A1(subkey[64]), .A2(state[64]), .Y(out[64]) );
  XOR2X1_HVT U86 ( .A1(subkey[32]), .A2(state[32]), .Y(out[32]) );
  XOR2X1_HVT U87 ( .A1(subkey[50]), .A2(state[50]), .Y(out[50]) );
  XOR2X1_HVT U88 ( .A1(subkey[37]), .A2(state[37]), .Y(out[37]) );
  XOR2X1_HVT U89 ( .A1(subkey[7]), .A2(state[7]), .Y(out[7]) );
  XOR2X1_HVT U90 ( .A1(subkey[102]), .A2(state[102]), .Y(out[102]) );
  XOR2X1_HVT U91 ( .A1(subkey[70]), .A2(state[70]), .Y(out[70]) );
  XOR2X1_HVT U92 ( .A1(subkey[38]), .A2(state[38]), .Y(out[38]) );
  XOR2X1_HVT U93 ( .A1(subkey[96]), .A2(state[96]), .Y(out[96]) );
  XOR2X1_HVT U94 ( .A1(subkey[77]), .A2(state[77]), .Y(out[77]) );
  XOR2X1_HVT U95 ( .A1(subkey[74]), .A2(state[74]), .Y(out[74]) );
  XOR2X1_HVT U96 ( .A1(subkey[106]), .A2(state[106]), .Y(out[106]) );
  XOR2X1_HVT U97 ( .A1(subkey[10]), .A2(state[10]), .Y(out[10]) );
  XOR2X1_HVT U98 ( .A1(subkey[2]), .A2(state[2]), .Y(out[2]) );
  XOR2X1_HVT U99 ( .A1(subkey[80]), .A2(state[80]), .Y(out[80]) );
  XOR2X1_HVT U100 ( .A1(subkey[82]), .A2(state[82]), .Y(out[82]) );
  XOR2X1_HVT U101 ( .A1(subkey[42]), .A2(state[42]), .Y(out[42]) );
  XOR2X1_HVT U102 ( .A1(subkey[61]), .A2(state[61]), .Y(out[61]) );
  XOR2X1_HVT U103 ( .A1(subkey[46]), .A2(state[46]), .Y(out[46]) );
  XOR2X1_HVT U104 ( .A1(subkey[5]), .A2(state[5]), .Y(out[5]) );
  XOR2X1_HVT U105 ( .A1(subkey[78]), .A2(state[78]), .Y(out[78]) );
  XOR2X1_HVT U106 ( .A1(subkey[93]), .A2(state[93]), .Y(out[93]) );
  XOR2X1_HVT U107 ( .A1(subkey[118]), .A2(state[118]), .Y(out[118]) );
  XOR2X1_HVT U108 ( .A1(subkey[85]), .A2(state[85]), .Y(out[85]) );
  XOR2X1_HVT U109 ( .A1(subkey[125]), .A2(state[125]), .Y(out[125]) );
  XOR2X1_HVT U110 ( .A1(subkey[110]), .A2(state[110]), .Y(out[110]) );
  XOR2X1_HVT U111 ( .A1(subkey[58]), .A2(state[58]), .Y(out[58]) );
  XOR2X1_HVT U112 ( .A1(subkey[14]), .A2(state[14]), .Y(out[14]) );
  XOR2X1_HVT U113 ( .A1(subkey[122]), .A2(state[122]), .Y(out[122]) );
  XOR2X1_HVT U114 ( .A1(subkey[114]), .A2(state[114]), .Y(out[114]) );
  XOR2X1_HVT U115 ( .A1(subkey[126]), .A2(state[126]), .Y(out[126]) );
  XOR2X1_HVT U116 ( .A1(subkey[8]), .A2(state[8]), .Y(out[8]) );
  XOR2X1_HVT U117 ( .A1(subkey[40]), .A2(state[40]), .Y(out[40]) );
  XOR2X1_HVT U118 ( .A1(subkey[72]), .A2(state[72]), .Y(out[72]) );
  XOR2X1_HVT U119 ( .A1(subkey[6]), .A2(state[6]), .Y(out[6]) );
  XOR2X1_HVT U120 ( .A1(subkey[90]), .A2(state[90]), .Y(out[90]) );
  XOR2X1_HVT U121 ( .A1(subkey[26]), .A2(state[26]), .Y(out[26]) );
  XOR2X1_HVT U122 ( .A1(subkey[66]), .A2(state[66]), .Y(out[66]) );
  XOR2X1_HVT U123 ( .A1(subkey[34]), .A2(state[34]), .Y(out[34]) );
  XOR2X1_HVT U124 ( .A1(subkey[22]), .A2(state[22]), .Y(out[22]) );
  XOR2X1_HVT U125 ( .A1(subkey[86]), .A2(state[86]), .Y(out[86]) );
  XOR2X1_HVT U126 ( .A1(subkey[54]), .A2(state[54]), .Y(out[54]) );
  XOR2X1_HVT U127 ( .A1(subkey[29]), .A2(state[29]), .Y(out[29]) );
  XOR2X1_HVT U128 ( .A1(subkey[21]), .A2(state[21]), .Y(out[21]) );
endmodule

