
module sbox_1 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n7, n10, n17, n18, n19, n23, n24, n48, n50, n118, n160, n170, n210,
         n211, n212, n213, n216, n217, n218, n219, n224, n225, n231, n232,
         n236, n238, n241, n242, n246, n249, n252, n261, n264, n269, n273,
         n274, n278, n280, n282, n283, n284, n285, n293, n296, n297, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781;

  NAND2X0_HVT U4 ( .A1(n348), .A2(n779), .Y(n778) );
  NAND2X0_HVT U5 ( .A1(n460), .A2(n344), .Y(n776) );
  NAND2X0_HVT U15 ( .A1(n779), .A2(n238), .Y(n768) );
  NAND2X0_HVT U21 ( .A1(n348), .A2(n367), .Y(n765) );
  NAND2X0_HVT U24 ( .A1(n466), .A2(n396), .Y(n764) );
  NAND2X0_HVT U33 ( .A1(n549), .A2(n464), .Y(n755) );
  NAND2X0_HVT U35 ( .A1(n280), .A2(n464), .Y(n753) );
  NAND2X0_HVT U42 ( .A1(n397), .A2(n443), .Y(n746) );
  NAND2X0_HVT U53 ( .A1(n736), .A2(n745), .Y(n737) );
  NAND2X0_HVT U56 ( .A1(n348), .A2(n732), .Y(n733) );
  NAND2X0_HVT U58 ( .A1(n510), .A2(n779), .Y(n730) );
  MUX41X1_HVT U61 ( .A1(n486), .A3(n432), .A2(n384), .A4(n238), .S0(n523), 
        .S1(n519), .Y(n727) );
  NAND2X0_HVT U62 ( .A1(n367), .A2(n370), .Y(n726) );
  MUX41X1_HVT U68 ( .A1(n538), .A3(n722), .A2(n721), .A4(n723), .S0(n497), 
        .S1(n522), .Y(n720) );
  NAND2X0_HVT U73 ( .A1(n416), .A2(n715), .Y(n716) );
  MUX41X1_HVT U75 ( .A1(n566), .A3(n564), .A2(n494), .A4(n527), .S0(n496), 
        .S1(n467), .Y(n713) );
  AND2X1_HVT U83 ( .A1(n343), .A2(n394), .Y(n704) );
  MUX41X1_HVT U90 ( .A1(n742), .A3(n746), .A2(n531), .A4(n699), .S0(n420), 
        .S1(n522), .Y(n698) );
  NAND2X0_HVT U101 ( .A1(n685), .A2(n684), .Y(n686) );
  MUX41X1_HVT U103 ( .A1(n303), .A3(n555), .A2(n544), .A4(n753), .S0(n497), 
        .S1(n468), .Y(n682) );
  MUX41X1_HVT U105 ( .A1(n562), .A3(n741), .A2(n681), .A4(n552), .S0(n420), 
        .S1(n521), .Y(n680) );
  NAND2X0_HVT U110 ( .A1(n507), .A2(n675), .Y(n676) );
  AND2X1_HVT U115 ( .A1(n308), .A2(n405), .Y(n671) );
  MUX41X1_HVT U116 ( .A1(n304), .A3(n671), .A2(n527), .A4(n757), .S0(n496), 
        .S1(n333), .Y(n670) );
  NAND2X0_HVT U123 ( .A1(n662), .A2(n661), .Y(n663) );
  MUX41X1_HVT U125 ( .A1(n765), .A3(n490), .A2(n538), .A4(n548), .S0(n496), 
        .S1(n297), .Y(n659) );
  MUX41X1_HVT U131 ( .A1(n654), .A3(n656), .A2(n655), .A4(n657), .S0(n499), 
        .S1(n297), .Y(n653) );
  MUX41X1_HVT U135 ( .A1(n540), .A3(n414), .A2(n776), .A4(n761), .S0(n497), 
        .S1(n523), .Y(n650) );
  AND2X1_HVT U140 ( .A1(n417), .A2(n391), .Y(n645) );
  NAND2X0_HVT U158 ( .A1(n318), .A2(n568), .Y(n629) );
  MUX41X1_HVT U159 ( .A1(n304), .A3(n238), .A2(n629), .A4(n570), .S0(n376), 
        .S1(n333), .Y(n628) );
  AND2X1_HVT U162 ( .A1(n372), .A2(n252), .Y(n625) );
  MUX41X1_HVT U165 ( .A1(n765), .A3(n561), .A2(n742), .A4(n19), .S0(n523), 
        .S1(n492), .Y(n623) );
  NAND2X0_HVT U167 ( .A1(n494), .A2(n367), .Y(n621) );
  MUX41X1_HVT U176 ( .A1(n217), .A3(n615), .A2(n539), .A4(n218), .S0(n467), 
        .S1(n492), .Y(n614) );
  NAND2X0_HVT U177 ( .A1(n435), .A2(n505), .Y(n613) );
  MUX41X1_HVT U178 ( .A1(n305), .A3(n613), .A2(n560), .A4(n750), .S0(n497), 
        .S1(n521), .Y(n612) );
  MUX41X1_HVT U179 ( .A1(n760), .A3(n559), .A2(n542), .A4(n560), .S0(n330), 
        .S1(n333), .Y(n611) );
  MUX41X1_HVT U180 ( .A1(n537), .A3(n284), .A2(n304), .A4(n482), .S0(n501), 
        .S1(n376), .Y(n610) );
  MUX41X1_HVT U182 ( .A1(n547), .A3(n348), .A2(n532), .A4(n556), .S0(n501), 
        .S1(n492), .Y(n608) );
  MUX41X1_HVT U189 ( .A1(n602), .A3(n218), .A2(n603), .A4(n552), .S0(n502), 
        .S1(n439), .Y(n601) );
  MUX41X1_HVT U194 ( .A1(n747), .A3(n406), .A2(n540), .A4(n417), .S0(n501), 
        .S1(n516), .Y(n597) );
  MUX41X1_HVT U195 ( .A1(n387), .A3(n565), .A2(n216), .A4(n751), .S0(n439), 
        .S1(n521), .Y(n596) );
  AO21X1_HVT U197 ( .A1(n487), .A2(n501), .A3(n563), .Y(n594) );
  MUX41X1_HVT U205 ( .A1(n394), .A3(n303), .A2(n559), .A4(n567), .S0(n376), 
        .S1(n522), .Y(n586) );
  NAND2X0_HVT U208 ( .A1(n397), .A2(n345), .Y(n675) );
  NAND2X0_HVT U212 ( .A1(n249), .A2(n415), .Y(n732) );
  NAND2X0_HVT U214 ( .A1(n372), .A2(n464), .Y(n584) );
  NAND2X0_HVT U215 ( .A1(n675), .A2(n416), .Y(n583) );
  NAND2X0_HVT U218 ( .A1(n414), .A2(n460), .Y(n635) );
  NAND2X0_HVT U220 ( .A1(n502), .A2(n584), .Y(n707) );
  INVX0_HVT U241 ( .A(n764), .Y(n573) );
  INVX0_HVT U242 ( .A(n746), .Y(n572) );
  INVX0_HVT U245 ( .A(n776), .Y(n570) );
  INVX0_HVT U256 ( .A(n635), .Y(n563) );
  INVX0_HVT U264 ( .A(n753), .Y(n557) );
  INVX0_HVT U265 ( .A(n762), .Y(n556) );
  INVX0_HVT U268 ( .A(n765), .Y(n553) );
  INVX0_HVT U270 ( .A(n583), .Y(n552) );
  INVX0_HVT U287 ( .A(n577), .Y(n540) );
  INVX0_HVT U289 ( .A(n684), .Y(n539) );
  INVX0_HVT U295 ( .A(n778), .Y(n537) );
  INVX0_HVT U296 ( .A(n768), .Y(n536) );
  INVX0_HVT U300 ( .A(n747), .Y(n532) );
  INVX0_HVT U303 ( .A(n576), .Y(n530) );
  INVX0_HVT U306 ( .A(n621), .Y(n529) );
  INVX1_HVT U1 ( .A(n769), .Y(n534) );
  INVX0_HVT U2 ( .A(n395), .Y(n754) );
  INVX1_HVT U3 ( .A(n10), .Y(n742) );
  INVX1_HVT U6 ( .A(n777), .Y(n347) );
  INVX1_HVT U7 ( .A(n518), .Y(n516) );
  INVX0_HVT U8 ( .A(n339), .Y(n280) );
  INVX1_HVT U9 ( .A(n775), .Y(n538) );
  AND2X1_HVT U10 ( .A1(n350), .A2(n571), .Y(n7) );
  INVX1_HVT U11 ( .A(n525), .Y(n476) );
  INVX1_HVT U12 ( .A(n473), .Y(n404) );
  XOR2X1_HVT U13 ( .A1(n473), .A2(n379), .Y(n10) );
  MUX41X1_HVT U14 ( .A1(n640), .A3(n639), .A2(n644), .A4(n643), .S0(n307), 
        .S1(n503), .Y(n638) );
  INVX0_HVT U16 ( .A(n338), .Y(n371) );
  MUX21X2_HVT U17 ( .A1(n484), .A2(n384), .S0(n495), .Y(n655) );
  MUX41X1_HVT U18 ( .A1(n672), .A3(n666), .A2(n658), .A4(n653), .S0(n311), 
        .S1(n451), .Y(out[3]) );
  INVX0_HVT U19 ( .A(n558), .Y(n350) );
  MUX41X1_HVT U20 ( .A1(n763), .A3(n434), .A2(n645), .A4(n545), .S0(n496), 
        .S1(n500), .Y(n644) );
  INVX0_HVT U22 ( .A(n500), .Y(n477) );
  INVX0_HVT U23 ( .A(n341), .Y(n369) );
  INVX1_HVT U25 ( .A(n524), .Y(n467) );
  XNOR2X1_HVT U26 ( .A1(n345), .A2(n318), .Y(n484) );
  NBUFFX2_HVT U27 ( .A(n461), .Y(n308) );
  MUX21X1_HVT U28 ( .A1(n347), .A2(n463), .S0(n460), .Y(n756) );
  INVX1_HVT U29 ( .A(n504), .Y(n463) );
  INVX1_HVT U30 ( .A(n371), .Y(n372) );
  INVX1_HVT U31 ( .A(n349), .Y(n343) );
  INVX1_HVT U32 ( .A(n525), .Y(n523) );
  INVX1_HVT U34 ( .A(n524), .Y(n333) );
  MUX21X1_HVT U36 ( .A1(n466), .A2(n753), .S0(n499), .Y(n738) );
  MUX21X1_HVT U37 ( .A1(n405), .A2(n568), .S0(n343), .Y(n775) );
  INVX1_HVT U38 ( .A(n497), .Y(n388) );
  INVX1_HVT U39 ( .A(n344), .Y(n443) );
  INVX1_HVT U40 ( .A(n489), .Y(n455) );
  MUX21X1_HVT U41 ( .A1(n415), .A2(n346), .S0(n461), .Y(n433) );
  INVX1_HVT U43 ( .A(n496), .Y(n383) );
  INVX1_HVT U44 ( .A(n755), .Y(n546) );
  INVX1_HVT U45 ( .A(n420), .Y(n444) );
  AO21X1_HVT U46 ( .A1(n497), .A2(n316), .A3(n338), .Y(n668) );
  INVX1_HVT U47 ( .A(n412), .Y(n413) );
  XOR2X1_HVT U48 ( .A1(n280), .A2(n460), .Y(n762) );
  INVX1_HVT U49 ( .A(n748), .Y(n528) );
  XNOR2X1_HVT U50 ( .A1(n518), .A2(n477), .Y(n454) );
  AO21X1_HVT U51 ( .A1(n464), .A2(n413), .A3(n246), .Y(n685) );
  MUX21X1_HVT U52 ( .A1(n549), .A2(n317), .S0(n391), .Y(n692) );
  MUX21X1_HVT U54 ( .A1(n676), .A2(n757), .S0(n436), .Y(n674) );
  AND3X1_HVT U55 ( .A1(n439), .A2(n396), .A3(n394), .Y(n656) );
  NAND2X0_HVT U57 ( .A1(n547), .A2(n297), .Y(n285) );
  NAND2X0_HVT U59 ( .A1(n535), .A2(n297), .Y(n336) );
  INVX1_HVT U60 ( .A(n675), .Y(n551) );
  MUX21X1_HVT U63 ( .A1(n631), .A2(n632), .S0(n373), .Y(n630) );
  MUX21X1_HVT U64 ( .A1(n619), .A2(n618), .S0(n376), .Y(n617) );
  OA21X1_HVT U65 ( .A1(n754), .A2(n50), .A3(n17), .Y(n606) );
  INVX1_HVT U66 ( .A(n491), .Y(n492) );
  MUX21X1_HVT U67 ( .A1(n417), .A2(n317), .S0(n435), .Y(n681) );
  INVX1_HVT U69 ( .A(n383), .Y(n330) );
  INVX1_HVT U70 ( .A(n584), .Y(n542) );
  INVX0_HVT U71 ( .A(n524), .Y(n468) );
  INVX1_HVT U72 ( .A(n467), .Y(n324) );
  INVX1_HVT U74 ( .A(n380), .Y(n511) );
  INVX1_HVT U76 ( .A(n424), .Y(n170) );
  INVX0_HVT U77 ( .A(n380), .Y(n460) );
  INVX1_HVT U78 ( .A(n512), .Y(n431) );
  INVX1_HVT U79 ( .A(n515), .Y(n379) );
  INVX1_HVT U80 ( .A(n379), .Y(n212) );
  INVX1_HVT U81 ( .A(n513), .Y(n396) );
  NBUFFX2_HVT U82 ( .A(n520), .Y(n499) );
  NBUFFX2_HVT U84 ( .A(n476), .Y(n500) );
  INVX0_HVT U85 ( .A(n380), .Y(n435) );
  INVX1_HVT U86 ( .A(n461), .Y(n391) );
  INVX0_HVT U87 ( .A(n7), .Y(n415) );
  INVX0_HVT U88 ( .A(n280), .Y(n394) );
  INVX0_HVT U89 ( .A(n568), .Y(n216) );
  AND2X1_HVT U91 ( .A1(n210), .A2(n211), .Y(n17) );
  AND2X1_HVT U92 ( .A1(n355), .A2(n356), .Y(n18) );
  AND2X1_HVT U93 ( .A1(n381), .A2(n382), .Y(n19) );
  INVX0_HVT U94 ( .A(n715), .Y(n569) );
  NAND2X0_HVT U95 ( .A1(n737), .A2(n324), .Y(n309) );
  INVX1_HVT U96 ( .A(n524), .Y(n297) );
  MUX21X1_HVT U97 ( .A1(n494), .A2(n421), .S0(n331), .Y(n493) );
  INVX0_HVT U98 ( .A(n365), .Y(n344) );
  AND3X1_HVT U99 ( .A1(n507), .A2(n118), .A3(n707), .Y(n708) );
  NAND2X0_HVT U100 ( .A1(n210), .A2(n211), .Y(n23) );
  MUX41X1_HVT U102 ( .A1(n772), .A3(n752), .A2(n756), .A4(n528), .S0(n324), 
        .S1(n492), .Y(n588) );
  MUX21X2_HVT U104 ( .A1(n507), .A2(n371), .S0(n511), .Y(n747) );
  INVX0_HVT U106 ( .A(n347), .Y(n346) );
  AND2X1_HVT U107 ( .A1(n328), .A2(n329), .Y(n24) );
  MUX41X1_HVT U108 ( .A1(n541), .A3(n733), .A2(n767), .A4(n773), .S0(n519), 
        .S1(n523), .Y(n731) );
  INVX1_HVT U109 ( .A(n772), .Y(n554) );
  INVX1_HVT U111 ( .A(n340), .Y(n320) );
  NBUFFX2_HVT U112 ( .A(n476), .Y(n502) );
  INVX1_HVT U113 ( .A(n502), .Y(n50) );
  INVX0_HVT U114 ( .A(n454), .Y(n428) );
  INVX0_HVT U117 ( .A(n7), .Y(n416) );
  MUX21X2_HVT U118 ( .A1(n345), .A2(n466), .S0(n514), .Y(n774) );
  INVX1_HVT U119 ( .A(n694), .Y(n550) );
  INVX1_HVT U120 ( .A(in[0]), .Y(n311) );
  NAND2X0_HVT U121 ( .A1(n316), .A2(n48), .Y(n770) );
  AND2X1_HVT U122 ( .A1(n315), .A2(n514), .Y(n48) );
  MUX41X1_HVT U124 ( .A1(n550), .A3(n774), .A2(n465), .A4(n712), .S0(n50), 
        .S1(n516), .Y(n711) );
  INVX1_HVT U126 ( .A(n516), .Y(n491) );
  OA21X1_HVT U127 ( .A1(n518), .A2(n423), .A3(n433), .Y(n677) );
  INVX0_HVT U128 ( .A(n368), .Y(n426) );
  NBUFFX2_HVT U129 ( .A(n781), .Y(n508) );
  INVX0_HVT U130 ( .A(n566), .Y(n118) );
  INVX0_HVT U132 ( .A(n342), .Y(n160) );
  MUX21X1_HVT U133 ( .A1(n415), .A2(n508), .S0(n396), .Y(n757) );
  MUX41X1_HVT U134 ( .A1(n526), .A3(n533), .A2(n531), .A4(n553), .S0(n297), 
        .S1(n409), .Y(n739) );
  NAND2X0_HVT U136 ( .A1(n443), .A2(n170), .Y(n210) );
  NAND2X0_HVT U137 ( .A1(n354), .A2(n424), .Y(n211) );
  MUX21X1_HVT U138 ( .A1(n345), .A2(n506), .S0(n514), .Y(n772) );
  INVX1_HVT U139 ( .A(n498), .Y(n307) );
  MUX41X1_HVT U141 ( .A1(n698), .A3(n691), .A2(n693), .A4(n690), .S0(n311), 
        .S1(n307), .Y(n689) );
  INVX1_HVT U142 ( .A(n353), .Y(n752) );
  MUX41X1_HVT U143 ( .A1(n252), .A3(n530), .A2(n742), .A4(n566), .S0(n388), 
        .S1(n333), .Y(n639) );
  INVX1_HVT U144 ( .A(n213), .Y(n719) );
  INVX0_HVT U145 ( .A(n379), .Y(n380) );
  INVX0_HVT U146 ( .A(n766), .Y(n533) );
  MUX21X1_HVT U147 ( .A1(n216), .A2(n580), .S0(n500), .Y(n213) );
  INVX0_HVT U148 ( .A(n580), .Y(n565) );
  INVX1_HVT U149 ( .A(n369), .Y(n370) );
  INVX1_HVT U150 ( .A(n463), .Y(n217) );
  INVX0_HVT U151 ( .A(n442), .Y(n773) );
  INVX0_HVT U152 ( .A(n763), .Y(n527) );
  NBUFFX2_HVT U153 ( .A(n770), .Y(n218) );
  NAND2X0_HVT U154 ( .A1(n314), .A2(n422), .Y(n219) );
  INVX0_HVT U155 ( .A(n759), .Y(n544) );
  NAND2X0_HVT U156 ( .A1(n406), .A2(n501), .Y(n225) );
  NAND2X0_HVT U157 ( .A1(n224), .A2(n477), .Y(n231) );
  NAND2X0_HVT U160 ( .A1(n225), .A2(n231), .Y(n744) );
  INVX0_HVT U161 ( .A(n761), .Y(n224) );
  MUX41X1_HVT U163 ( .A1(n651), .A3(n650), .A2(n649), .A4(n647), .S0(n307), 
        .S1(n311), .Y(n646) );
  NAND2X0_HVT U164 ( .A1(n372), .A2(n367), .Y(n232) );
  NAND2X0_HVT U166 ( .A1(n217), .A2(n511), .Y(n236) );
  NAND2X0_HVT U168 ( .A1(n232), .A2(n236), .Y(n712) );
  NAND2X0_HVT U169 ( .A1(n219), .A2(n315), .Y(n238) );
  INVX0_HVT U170 ( .A(n771), .Y(n543) );
  INVX1_HVT U171 ( .A(n522), .Y(n246) );
  INVX0_HVT U172 ( .A(n524), .Y(n522) );
  MUX21X2_HVT U173 ( .A1(n466), .A2(n405), .S0(n460), .Y(n465) );
  INVX1_HVT U174 ( .A(n404), .Y(n405) );
  INVX0_HVT U175 ( .A(n524), .Y(n521) );
  MUX21X1_HVT U181 ( .A1(n305), .A2(n545), .S0(n495), .Y(n654) );
  INVX0_HVT U183 ( .A(n305), .Y(n432) );
  INVX1_HVT U184 ( .A(n212), .Y(n461) );
  NAND2X0_HVT U185 ( .A1(n241), .A2(n500), .Y(n242) );
  AND2X1_HVT U186 ( .A1(n242), .A2(n757), .Y(n618) );
  INVX0_HVT U187 ( .A(n488), .Y(n241) );
  MUX41X1_HVT U188 ( .A1(n674), .A3(n677), .A2(n673), .A4(n678), .S0(n499), 
        .S1(n246), .Y(n672) );
  MUX41X1_HVT U190 ( .A1(n610), .A3(n612), .A2(n611), .A4(n614), .S0(n503), 
        .S1(n498), .Y(n609) );
  INVX1_HVT U191 ( .A(n212), .Y(n249) );
  INVX1_HVT U192 ( .A(n569), .Y(n252) );
  NAND2X0_HVT U193 ( .A1(n170), .A2(n510), .Y(n715) );
  NAND2X0_HVT U196 ( .A1(n466), .A2(n170), .Y(n261) );
  NAND2X0_HVT U198 ( .A1(n426), .A2(n396), .Y(n264) );
  NAND2X0_HVT U199 ( .A1(n261), .A2(n264), .Y(n767) );
  INVX1_HVT U200 ( .A(n344), .Y(n466) );
  INVX0_HVT U201 ( .A(n756), .Y(n545) );
  NAND2X0_HVT U202 ( .A1(n413), .A2(n498), .Y(n269) );
  NAND2X0_HVT U203 ( .A1(n555), .A2(n409), .Y(n273) );
  NAND2X0_HVT U204 ( .A1(n269), .A2(n273), .Y(n721) );
  INVX0_HVT U206 ( .A(n767), .Y(n526) );
  NBUFFX2_HVT U207 ( .A(n280), .Y(n505) );
  MUX21X2_HVT U209 ( .A1(n508), .A2(n443), .S0(n512), .Y(n395) );
  INVX1_HVT U210 ( .A(n212), .Y(n318) );
  INVX0_HVT U211 ( .A(n513), .Y(n367) );
  INVX0_HVT U213 ( .A(n513), .Y(n464) );
  INVX0_HVT U216 ( .A(n366), .Y(n339) );
  NAND2X0_HVT U217 ( .A1(n414), .A2(n523), .Y(n274) );
  NAND2X0_HVT U219 ( .A1(n462), .A2(n465), .Y(n278) );
  NAND2X0_HVT U221 ( .A1(n274), .A2(n278), .Y(n637) );
  XNOR2X2_HVT U222 ( .A1(n504), .A2(n320), .Y(n317) );
  MUX21X1_HVT U223 ( .A1(n568), .A2(n317), .S0(n249), .Y(n626) );
  MUX41X1_HVT U224 ( .A1(n586), .A3(n588), .A2(n587), .A4(n589), .S0(n503), 
        .S1(n498), .Y(n585) );
  INVX1_HVT U225 ( .A(n571), .Y(n323) );
  NAND2X0_HVT U226 ( .A1(n554), .A2(n409), .Y(n282) );
  NAND2X0_HVT U227 ( .A1(n396), .A2(n499), .Y(n283) );
  NAND2X0_HVT U228 ( .A1(n282), .A2(n283), .Y(n723) );
  INVX0_HVT U229 ( .A(n555), .Y(n284) );
  INVX1_HVT U230 ( .A(n574), .Y(n559) );
  NAND2X0_HVT U231 ( .A1(n50), .A2(n23), .Y(n293) );
  NAND2X0_HVT U232 ( .A1(n285), .A2(n293), .Y(n648) );
  MUX21X1_HVT U233 ( .A1(n346), .A2(n508), .S0(n424), .Y(n434) );
  INVX1_HVT U234 ( .A(n319), .Y(n296) );
  INVX1_HVT U235 ( .A(n370), .Y(n319) );
  MUX41X1_HVT U236 ( .A1(n701), .A3(n703), .A2(n705), .A4(n706), .S0(n520), 
        .S1(n503), .Y(n700) );
  INVX1_HVT U237 ( .A(n582), .Y(n531) );
  NAND2X0_HVT U238 ( .A1(n538), .A2(n297), .Y(n302) );
  AND2X1_HVT U239 ( .A1(n302), .A2(n434), .Y(n590) );
  INVX1_HVT U240 ( .A(n535), .Y(n303) );
  INVX0_HVT U243 ( .A(n779), .Y(n535) );
  INVX0_HVT U244 ( .A(n543), .Y(n304) );
  INVX1_HVT U246 ( .A(n504), .Y(n314) );
  MUX21X1_HVT U247 ( .A1(n314), .A2(n160), .S0(n461), .Y(n305) );
  MUX41X1_HVT U248 ( .A1(n17), .A3(n238), .A2(n551), .A4(n416), .S0(n420), 
        .S1(n523), .Y(n643) );
  NBUFFX2_HVT U249 ( .A(n517), .Y(n420) );
  NAND2X0_HVT U250 ( .A1(n571), .A2(n558), .Y(n777) );
  INVX0_HVT U251 ( .A(n571), .Y(n365) );
  INVX1_HVT U252 ( .A(in[3]), .Y(n571) );
  NBUFFX2_HVT U253 ( .A(n541), .Y(n306) );
  INVX0_HVT U254 ( .A(n518), .Y(n517) );
  MUX41X1_HVT U255 ( .A1(n682), .A3(n687), .A2(n680), .A4(n683), .S0(in[0]), 
        .S1(n307), .Y(n679) );
  NAND2X0_HVT U257 ( .A1(n738), .A2(n501), .Y(n310) );
  NAND2X0_HVT U258 ( .A1(n309), .A2(n310), .Y(n735) );
  MUX41X1_HVT U259 ( .A1(n624), .A3(n623), .A2(n620), .A4(n617), .S0(n409), 
        .S1(n311), .Y(n616) );
  NAND2X0_HVT U260 ( .A1(n708), .A2(n373), .Y(n312) );
  NAND2X0_HVT U261 ( .A1(n709), .A2(n436), .Y(n313) );
  NAND2X0_HVT U262 ( .A1(n312), .A2(n313), .Y(n706) );
  NAND2X0_HVT U263 ( .A1(n504), .A2(n320), .Y(n315) );
  NAND2X0_HVT U266 ( .A1(n314), .A2(n422), .Y(n316) );
  NAND2X0_HVT U267 ( .A1(n316), .A2(n315), .Y(n354) );
  INVX1_HVT U269 ( .A(n380), .Y(n514) );
  INVX0_HVT U271 ( .A(n749), .Y(n547) );
  MUX21X1_HVT U272 ( .A1(n417), .A2(n548), .S0(n477), .Y(n652) );
  INVX0_HVT U273 ( .A(n513), .Y(n424) );
  MUX41X1_HVT U274 ( .A1(n536), .A3(n726), .A2(n534), .A4(n543), .S0(n50), 
        .S1(n519), .Y(n725) );
  NBUFFX2_HVT U275 ( .A(n517), .Y(n495) );
  NBUFFX2_HVT U276 ( .A(n517), .Y(n496) );
  NBUFFX2_HVT U277 ( .A(n517), .Y(n497) );
  INVX0_HVT U278 ( .A(n760), .Y(n562) );
  INVX1_HVT U279 ( .A(n774), .Y(n555) );
  XOR2X2_HVT U280 ( .A1(n318), .A2(n413), .Y(n743) );
  MUX21X2_HVT U281 ( .A1(n557), .A2(n395), .S0(n495), .Y(n669) );
  NAND2X0_HVT U282 ( .A1(n394), .A2(n431), .Y(n321) );
  NAND2X0_HVT U283 ( .A1(n338), .A2(n435), .Y(n322) );
  NAND2X0_HVT U284 ( .A1(n322), .A2(n321), .Y(n581) );
  INVX0_HVT U285 ( .A(n581), .Y(n541) );
  INVX1_HVT U286 ( .A(in[7]), .Y(n525) );
  MUX41X1_HVT U288 ( .A1(n487), .A3(n564), .A2(n483), .A4(n702), .S0(n324), 
        .S1(n420), .Y(n701) );
  INVX1_HVT U290 ( .A(n476), .Y(n524) );
  MUX41X1_HVT U291 ( .A1(n598), .A3(n597), .A2(n596), .A4(n593), .S0(n307), 
        .S1(n311), .Y(n592) );
  NAND2X0_HVT U292 ( .A1(n638), .A2(n451), .Y(n478) );
  MUX21X1_HVT U293 ( .A1(n404), .A2(n494), .S0(n249), .Y(n763) );
  INVX0_HVT U294 ( .A(in[4]), .Y(n558) );
  INVX0_HVT U297 ( .A(n323), .Y(n422) );
  NAND2X0_HVT U298 ( .A1(n339), .A2(n340), .Y(n325) );
  INVX1_HVT U299 ( .A(n365), .Y(n340) );
  NAND2X0_HVT U301 ( .A1(n443), .A2(n431), .Y(n326) );
  NAND2X0_HVT U302 ( .A1(n509), .A2(n511), .Y(n327) );
  NAND2X0_HVT U304 ( .A1(n326), .A2(n327), .Y(n442) );
  INVX1_HVT U305 ( .A(n515), .Y(n513) );
  NAND2X0_HVT U307 ( .A1(n466), .A2(n170), .Y(n328) );
  NAND2X0_HVT U308 ( .A1(n338), .A2(n391), .Y(n329) );
  NAND2X0_HVT U309 ( .A1(n328), .A2(n329), .Y(n384) );
  MUX41X1_HVT U310 ( .A1(n605), .A3(n608), .A2(n601), .A4(n604), .S0(n520), 
        .S1(n311), .Y(n600) );
  INVX1_HVT U311 ( .A(in[2]), .Y(n518) );
  NAND2X0_HVT U312 ( .A1(n770), .A2(n510), .Y(n771) );
  MUX41X1_HVT U313 ( .A1(n483), .A3(n755), .A2(n530), .A4(n752), .S0(n330), 
        .S1(n523), .Y(n649) );
  INVX0_HVT U314 ( .A(n757), .Y(n567) );
  XNOR2X1_HVT U315 ( .A1(n510), .A2(n249), .Y(n487) );
  MUX41X1_HVT U316 ( .A1(n17), .A3(n387), .A2(n24), .A4(n704), .S0(n496), .S1(
        n467), .Y(n703) );
  XNOR2X1_HVT U317 ( .A1(n391), .A2(n491), .Y(n331) );
  INVX0_HVT U318 ( .A(n508), .Y(n568) );
  INVX1_HVT U319 ( .A(n493), .Y(n673) );
  INVX1_HVT U320 ( .A(in[1]), .Y(n515) );
  NAND2X0_HVT U321 ( .A1(n695), .A2(n436), .Y(n458) );
  NAND2X0_HVT U322 ( .A1(n442), .A2(n499), .Y(n332) );
  NAND2X0_HVT U323 ( .A1(n332), .A2(n252), .Y(n722) );
  NAND2X0_HVT U324 ( .A1(n750), .A2(n477), .Y(n334) );
  NAND2X0_HVT U325 ( .A1(n550), .A2(n500), .Y(n335) );
  NAND2X0_HVT U326 ( .A1(n334), .A2(n335), .Y(n631) );
  INVX0_HVT U327 ( .A(n434), .Y(n750) );
  MUX41X1_HVT U328 ( .A1(n743), .A3(n533), .A2(n573), .A4(n769), .S0(n420), 
        .S1(n467), .Y(n705) );
  MUX21X1_HVT U329 ( .A1(n217), .A2(n317), .S0(n431), .Y(n684) );
  MUX21X1_HVT U330 ( .A1(n567), .A2(n769), .S0(n516), .Y(n688) );
  NAND2X0_HVT U331 ( .A1(n479), .A2(n478), .Y(out[4]) );
  NAND2X0_HVT U332 ( .A1(n759), .A2(n462), .Y(n337) );
  NAND2X0_HVT U333 ( .A1(n336), .A2(n337), .Y(n642) );
  AND2X1_HVT U334 ( .A1(n342), .A2(n780), .Y(n338) );
  NAND2X0_HVT U335 ( .A1(n323), .A2(n366), .Y(n341) );
  NAND2X0_HVT U336 ( .A1(n339), .A2(n340), .Y(n342) );
  NAND2X0_HVT U337 ( .A1(n325), .A2(n341), .Y(n473) );
  OR2X1_HVT U338 ( .A1(n509), .A2(n396), .Y(n418) );
  MUX21X2_HVT U339 ( .A1(n368), .A2(n415), .S0(n514), .Y(n769) );
  INVX1_HVT U340 ( .A(n379), .Y(n349) );
  OA21X1_HVT U341 ( .A1(n529), .A2(n324), .A3(n352), .Y(n641) );
  INVX0_HVT U342 ( .A(n567), .Y(n352) );
  NBUFFX2_HVT U343 ( .A(n558), .Y(n504) );
  MUX21X1_HVT U344 ( .A1(n217), .A2(n549), .S0(n308), .Y(n759) );
  INVX1_HVT U345 ( .A(n349), .Y(n512) );
  NBUFFX2_HVT U346 ( .A(n777), .Y(n345) );
  INVX1_HVT U347 ( .A(n347), .Y(n348) );
  INVX1_HVT U348 ( .A(n346), .Y(n549) );
  INVX0_HVT U349 ( .A(in[4]), .Y(n366) );
  INVX1_HVT U350 ( .A(n451), .Y(n351) );
  INVX1_HVT U351 ( .A(in[6]), .Y(n451) );
  MUX21X1_HVT U352 ( .A1(n510), .A2(n280), .S0(n367), .Y(n353) );
  XNOR2X1_HVT U353 ( .A1(n296), .A2(n464), .Y(n740) );
  MUX41X1_HVT U354 ( .A1(n740), .A3(n599), .A2(n746), .A4(n753), .S0(n330), 
        .S1(n462), .Y(n598) );
  NAND2X0_HVT U355 ( .A1(n367), .A2(n568), .Y(n702) );
  MUX41X1_HVT U356 ( .A1(n720), .A3(n728), .A2(n724), .A4(n734), .S0(n351), 
        .S1(n503), .Y(out[0]) );
  INVX1_HVT U357 ( .A(n758), .Y(n561) );
  MUX21X1_HVT U358 ( .A1(n344), .A2(n463), .S0(n318), .Y(n758) );
  NAND2X0_HVT U359 ( .A1(n583), .A2(n297), .Y(n355) );
  NAND2X0_HVT U360 ( .A1(n758), .A2(n462), .Y(n356) );
  NAND2X0_HVT U361 ( .A1(n739), .A2(n439), .Y(n357) );
  NAND2X0_HVT U362 ( .A1(n735), .A2(n383), .Y(n358) );
  NAND2X0_HVT U363 ( .A1(n357), .A2(n358), .Y(n734) );
  MUX41X1_HVT U364 ( .A1(n485), .A3(n566), .A2(n768), .A4(n343), .S0(n388), 
        .S1(n522), .Y(n690) );
  NAND2X0_HVT U365 ( .A1(n641), .A2(n439), .Y(n359) );
  NAND2X0_HVT U366 ( .A1(n642), .A2(n383), .Y(n360) );
  NAND2X0_HVT U367 ( .A1(n359), .A2(n360), .Y(n640) );
  MUX41X1_HVT U368 ( .A1(n711), .A3(n713), .A2(n714), .A4(n718), .S0(n520), 
        .S1(n503), .Y(n710) );
  NAND2X0_HVT U369 ( .A1(n731), .A2(n376), .Y(n361) );
  NAND2X0_HVT U370 ( .A1(n729), .A2(n444), .Y(n362) );
  NAND2X0_HVT U371 ( .A1(n362), .A2(n361), .Y(n728) );
  INVX0_HVT U372 ( .A(n732), .Y(n566) );
  MUX41X1_HVT U373 ( .A1(n485), .A3(n573), .A2(n692), .A4(n565), .S0(n444), 
        .S1(n468), .Y(n691) );
  NAND2X0_HVT U374 ( .A1(n778), .A2(n439), .Y(n363) );
  NAND2X0_HVT U375 ( .A1(n648), .A2(n436), .Y(n364) );
  NAND2X0_HVT U376 ( .A1(n364), .A2(n363), .Y(n647) );
  XNOR2X1_HVT U377 ( .A1(n476), .A2(n424), .Y(n489) );
  MUX41X1_HVT U378 ( .A1(n630), .A3(n628), .A2(n634), .A4(n633), .S0(n307), 
        .S1(n503), .Y(n627) );
  MUX41X1_HVT U379 ( .A1(n304), .A3(n733), .A2(n23), .A4(n395), .S0(n491), 
        .S1(n468), .Y(n587) );
  XNOR2X1_HVT U380 ( .A1(n343), .A2(n422), .Y(n741) );
  INVX1_HVT U381 ( .A(n369), .Y(n368) );
  NAND2X0_HVT U382 ( .A1(n303), .A2(n373), .Y(n374) );
  NAND2X0_HVT U383 ( .A1(n353), .A2(n383), .Y(n375) );
  NAND2X0_HVT U384 ( .A1(n374), .A2(n375), .Y(n678) );
  INVX0_HVT U385 ( .A(n383), .Y(n373) );
  NAND2X0_HVT U386 ( .A1(n719), .A2(n376), .Y(n377) );
  NAND2X0_HVT U387 ( .A1(n744), .A2(n436), .Y(n378) );
  NAND2X0_HVT U388 ( .A1(n377), .A2(n378), .Y(n718) );
  INVX0_HVT U389 ( .A(n436), .Y(n376) );
  INVX1_HVT U390 ( .A(n517), .Y(n436) );
  INVX0_HVT U391 ( .A(n425), .Y(n632) );
  NAND2X0_HVT U392 ( .A1(n18), .A2(n388), .Y(n437) );
  NAND2X0_HVT U393 ( .A1(n296), .A2(n170), .Y(n381) );
  NAND2X0_HVT U394 ( .A1(n417), .A2(n431), .Y(n382) );
  INVX0_HVT U395 ( .A(n423), .Y(n751) );
  MUX21X2_HVT U396 ( .A1(n668), .A2(n669), .S0(n502), .Y(n667) );
  NAND2X0_HVT U397 ( .A1(n416), .A2(n50), .Y(n385) );
  NAND2X0_HVT U398 ( .A1(n565), .A2(n500), .Y(n386) );
  NAND2X0_HVT U399 ( .A1(n385), .A2(n386), .Y(n619) );
  NBUFFX2_HVT U400 ( .A(n372), .Y(n387) );
  MUX41X1_HVT U401 ( .A1(n762), .A3(n717), .A2(n764), .A4(n716), .S0(n388), 
        .S1(n333), .Y(n714) );
  NAND2X0_HVT U402 ( .A1(n727), .A2(n373), .Y(n389) );
  NAND2X0_HVT U403 ( .A1(n725), .A2(n444), .Y(n390) );
  NAND2X0_HVT U404 ( .A1(n390), .A2(n389), .Y(n724) );
  MUX41X1_HVT U405 ( .A1(n625), .A3(n432), .A2(n626), .A4(n484), .S0(n491), 
        .S1(n468), .Y(n624) );
  OA21X1_HVT U406 ( .A1(n748), .A2(n324), .A3(n635), .Y(n636) );
  MUX21X1_HVT U407 ( .A1(n506), .A2(n494), .S0(n512), .Y(n748) );
  NAND2X0_HVT U408 ( .A1(n600), .A2(n451), .Y(n392) );
  NAND2X0_HVT U409 ( .A1(n609), .A2(n351), .Y(n393) );
  NAND2X0_HVT U410 ( .A1(n392), .A2(n393), .Y(out[6]) );
  MUX21X1_HVT U411 ( .A1(n607), .A2(n606), .S0(n436), .Y(n605) );
  INVX1_HVT U412 ( .A(n368), .Y(n494) );
  AO21X1_HVT U413 ( .A1(n502), .A2(n694), .A3(n563), .Y(n695) );
  INVX1_HVT U414 ( .A(n349), .Y(n397) );
  INVX1_HVT U415 ( .A(n519), .Y(n409) );
  NAND2X0_HVT U416 ( .A1(n416), .A2(n467), .Y(n398) );
  NAND2X0_HVT U417 ( .A1(n766), .A2(n50), .Y(n399) );
  NAND2X0_HVT U418 ( .A1(n398), .A2(n399), .Y(n709) );
  MUX21X1_HVT U419 ( .A1(n463), .A2(n370), .S0(n512), .Y(n766) );
  NAND2X0_HVT U420 ( .A1(n562), .A2(n444), .Y(n400) );
  NAND2X0_HVT U421 ( .A1(n758), .A2(n496), .Y(n401) );
  NAND2X0_HVT U422 ( .A1(n401), .A2(n400), .Y(n657) );
  NAND2X0_HVT U423 ( .A1(n686), .A2(n388), .Y(n402) );
  NAND2X0_HVT U424 ( .A1(n18), .A2(n330), .Y(n403) );
  NAND2X0_HVT U425 ( .A1(n403), .A2(n402), .Y(n683) );
  NAND2X0_HVT U426 ( .A1(n418), .A2(n419), .Y(n406) );
  NAND2X0_HVT U427 ( .A1(n594), .A2(n330), .Y(n407) );
  NAND2X0_HVT U428 ( .A1(n595), .A2(n388), .Y(n408) );
  NAND2X0_HVT U429 ( .A1(n407), .A2(n408), .Y(n593) );
  MUX21X1_HVT U430 ( .A1(n572), .A2(n560), .S0(n500), .Y(n595) );
  NAND2X0_HVT U431 ( .A1(n636), .A2(n388), .Y(n410) );
  NAND2X0_HVT U432 ( .A1(n637), .A2(n330), .Y(n411) );
  NAND2X0_HVT U433 ( .A1(n410), .A2(n411), .Y(n634) );
  MUX41X1_HVT U434 ( .A1(n306), .A3(n417), .A2(n621), .A4(n622), .S0(n330), 
        .S1(n521), .Y(n620) );
  NAND2X0_HVT U435 ( .A1(n216), .A2(n732), .Y(n622) );
  INVX1_HVT U436 ( .A(n160), .Y(n412) );
  INVX1_HVT U437 ( .A(n412), .Y(n414) );
  INVX1_HVT U438 ( .A(n7), .Y(n417) );
  NAND2X0_HVT U439 ( .A1(n426), .A2(n464), .Y(n419) );
  NAND2X0_HVT U440 ( .A1(n418), .A2(n419), .Y(n761) );
  MUX21X1_HVT U441 ( .A1(n422), .A2(n505), .S0(n495), .Y(n421) );
  NBUFFX2_HVT U442 ( .A(n476), .Y(n501) );
  INVX0_HVT U443 ( .A(n500), .Y(n462) );
  MUX21X1_HVT U444 ( .A1(n405), .A2(n549), .S0(n464), .Y(n423) );
  INVX1_HVT U445 ( .A(n575), .Y(n560) );
  MUX21X1_HVT U446 ( .A1(n427), .A2(n426), .S0(n489), .Y(n425) );
  NAND2X0_HVT U447 ( .A1(n501), .A2(n443), .Y(n427) );
  INVX1_HVT U448 ( .A(n579), .Y(n564) );
  NAND2X0_HVT U449 ( .A1(n688), .A2(n428), .Y(n429) );
  NAND2X0_HVT U450 ( .A1(n486), .A2(n454), .Y(n430) );
  NAND2X0_HVT U451 ( .A1(n429), .A2(n430), .Y(n687) );
  NAND2X0_HVT U452 ( .A1(n453), .A2(n452), .Y(out[1]) );
  NAND2X0_HVT U453 ( .A1(n689), .A2(n351), .Y(n449) );
  NAND2X0_HVT U454 ( .A1(n480), .A2(n481), .Y(n666) );
  NAND2X0_HVT U455 ( .A1(n652), .A2(n373), .Y(n438) );
  NAND2X0_HVT U456 ( .A1(n437), .A2(n438), .Y(n651) );
  NAND2X0_HVT U457 ( .A1(n472), .A2(n471), .Y(out[5]) );
  OR2X1_HVT U458 ( .A1(n424), .A2(n319), .Y(n779) );
  NAND2X0_HVT U459 ( .A1(n591), .A2(n439), .Y(n440) );
  NAND2X0_HVT U460 ( .A1(n590), .A2(n388), .Y(n441) );
  NAND2X0_HVT U461 ( .A1(n441), .A2(n440), .Y(n589) );
  INVX0_HVT U462 ( .A(n436), .Y(n439) );
  NAND2X0_HVT U463 ( .A1(n546), .A2(n444), .Y(n445) );
  NAND2X0_HVT U464 ( .A1(n665), .A2(n420), .Y(n446) );
  NAND2X0_HVT U465 ( .A1(n445), .A2(n446), .Y(n664) );
  NAND2X0_HVT U466 ( .A1(n659), .A2(n307), .Y(n447) );
  NAND2X0_HVT U467 ( .A1(n660), .A2(n498), .Y(n448) );
  NAND2X0_HVT U468 ( .A1(n447), .A2(n448), .Y(n658) );
  MUX21X1_HVT U469 ( .A1(n664), .A2(n663), .S0(n501), .Y(n660) );
  MUX41X1_HVT U470 ( .A1(n730), .A3(n490), .A2(n433), .A4(n488), .S0(n50), 
        .S1(n519), .Y(n729) );
  NAND2X0_HVT U471 ( .A1(n679), .A2(n451), .Y(n450) );
  NAND2X0_HVT U472 ( .A1(n449), .A2(n450), .Y(out[2]) );
  NAND2X0_HVT U473 ( .A1(n700), .A2(n451), .Y(n452) );
  NAND2X0_HVT U474 ( .A1(n710), .A2(n351), .Y(n453) );
  INVX1_HVT U475 ( .A(n578), .Y(n548) );
  NAND2X0_HVT U476 ( .A1(n296), .A2(n455), .Y(n456) );
  NAND2X0_HVT U477 ( .A1(n697), .A2(n489), .Y(n457) );
  NAND2X0_HVT U478 ( .A1(n457), .A2(n456), .Y(n696) );
  NAND2X0_HVT U479 ( .A1(n696), .A2(n373), .Y(n459) );
  NAND2X0_HVT U480 ( .A1(n458), .A2(n459), .Y(n693) );
  MUX41X1_HVT U481 ( .A1(n749), .A3(n485), .A2(n742), .A4(n252), .S0(n491), 
        .S1(n521), .Y(n604) );
  NAND2X0_HVT U482 ( .A1(n585), .A2(n451), .Y(n469) );
  NAND2X0_HVT U483 ( .A1(n592), .A2(n351), .Y(n470) );
  NAND2X0_HVT U484 ( .A1(n469), .A2(n470), .Y(out[7]) );
  MUX41X1_HVT U485 ( .A1(n676), .A3(n296), .A2(n486), .A4(n557), .S0(n468), 
        .S1(n497), .Y(n633) );
  NAND2X0_HVT U486 ( .A1(n627), .A2(in[6]), .Y(n471) );
  NAND2X0_HVT U487 ( .A1(n616), .A2(n451), .Y(n472) );
  NAND2X0_HVT U488 ( .A1(n482), .A2(n297), .Y(n474) );
  NAND2X0_HVT U489 ( .A1(n24), .A2(n50), .Y(n475) );
  NAND2X0_HVT U490 ( .A1(n474), .A2(n475), .Y(n591) );
  NAND2X0_HVT U491 ( .A1(n646), .A2(n351), .Y(n479) );
  NAND2X0_HVT U492 ( .A1(n667), .A2(n409), .Y(n480) );
  NAND2X0_HVT U493 ( .A1(n670), .A2(n499), .Y(n481) );
  AND2X1_HVT U494 ( .A1(n238), .A2(n732), .Y(n482) );
  MUX21X1_HVT U495 ( .A1(n347), .A2(n568), .S0(n499), .Y(n736) );
  AND2X1_HVT U496 ( .A1(n507), .A2(n715), .Y(n483) );
  MUX21X1_HVT U497 ( .A1(n549), .A2(n426), .S0(n511), .Y(n615) );
  MUX21X1_HVT U498 ( .A1(n338), .A2(n413), .S0(n308), .Y(n577) );
  MUX21X1_HVT U499 ( .A1(n549), .A2(n505), .S0(n343), .Y(n578) );
  NBUFFX2_HVT U500 ( .A(n780), .Y(n507) );
  MUX21X1_HVT U501 ( .A1(n348), .A2(n417), .S0(n435), .Y(n699) );
  MUX21X1_HVT U502 ( .A1(n507), .A2(n348), .S0(n511), .Y(n576) );
  MUX21X1_HVT U503 ( .A1(n348), .A2(n509), .S0(n513), .Y(n694) );
  MUX21X1_HVT U504 ( .A1(n217), .A2(n506), .S0(n397), .Y(n665) );
  MUX21X1_HVT U505 ( .A1(n506), .A2(n216), .S0(n318), .Y(n602) );
  MUX21X1_HVT U506 ( .A1(n509), .A2(n507), .S0(n170), .Y(n603) );
  MUX21X1_HVT U507 ( .A1(n344), .A2(n505), .S0(n435), .Y(n599) );
  MUX21X1_HVT U508 ( .A1(n370), .A2(n280), .S0(n511), .Y(n582) );
  AND2X1_HVT U509 ( .A1(n308), .A2(n426), .Y(n485) );
  MUX21X1_HVT U510 ( .A1(n219), .A2(n506), .S0(n249), .Y(n580) );
  AND2X1_HVT U511 ( .A1(n509), .A2(n675), .Y(n486) );
  MUX21X1_HVT U512 ( .A1(n415), .A2(n366), .S0(n343), .Y(n717) );
  MUX21X1_HVT U513 ( .A1(n416), .A2(n216), .S0(n495), .Y(n662) );
  NBUFFX2_HVT U514 ( .A(n422), .Y(n506) );
  NBUFFX2_HVT U515 ( .A(n520), .Y(n498) );
  MUX21X1_HVT U516 ( .A1(n702), .A2(n466), .S0(n501), .Y(n607) );
  MUX21X1_HVT U517 ( .A1(n443), .A2(n549), .S0(n397), .Y(n749) );
  NAND2X0_HVT U518 ( .A1(n323), .A2(n366), .Y(n780) );
  AND2X1_HVT U519 ( .A1(n317), .A2(n396), .Y(n488) );
  XOR2X1_HVT U520 ( .A1(n308), .A2(n498), .Y(n745) );
  MUX21X1_HVT U521 ( .A1(n466), .A2(n414), .S0(n397), .Y(n579) );
  MUX21X1_HVT U522 ( .A1(n779), .A2(n391), .S0(n495), .Y(n661) );
  NBUFFX2_HVT U523 ( .A(n781), .Y(n510) );
  MUX21X1_HVT U524 ( .A1(n443), .A2(n217), .S0(n502), .Y(n697) );
  NBUFFX2_HVT U525 ( .A(n781), .Y(n509) );
  AND2X1_HVT U526 ( .A1(n506), .A2(n367), .Y(n490) );
  NBUFFX2_HVT U527 ( .A(in[5]), .Y(n520) );
  NBUFFX2_HVT U528 ( .A(in[5]), .Y(n519) );
  NAND2X0_HVT U529 ( .A1(n350), .A2(n323), .Y(n781) );
  MUX21X1_HVT U530 ( .A1(n463), .A2(n416), .S0(n435), .Y(n575) );
  MUX21X1_HVT U531 ( .A1(n509), .A2(n394), .S0(n397), .Y(n760) );
  MUX21X1_HVT U532 ( .A1(n394), .A2(n510), .S0(n512), .Y(n574) );
  NBUFFX2_HVT U533 ( .A(in[0]), .Y(n503) );
endmodule

