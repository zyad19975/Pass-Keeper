
module sbox_12 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n50, n210, n211, n212, n213, n216, n217, n218, n219, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604;

  NAND2X0_HVT U4 ( .A1(n307), .A2(n602), .Y(n601) );
  NAND2X0_HVT U5 ( .A1(n311), .A2(n296), .Y(n599) );
  NAND2X0_HVT U13 ( .A1(n591), .A2(n309), .Y(n592) );
  NAND2X0_HVT U15 ( .A1(n602), .A2(n298), .Y(n589) );
  NAND2X0_HVT U21 ( .A1(n307), .A2(n316), .Y(n583) );
  NAND2X0_HVT U24 ( .A1(n304), .A2(n316), .Y(n581) );
  NAND2X0_HVT U33 ( .A1(n380), .A2(n316), .Y(n572) );
  NAND2X0_HVT U35 ( .A1(n301), .A2(n316), .Y(n570) );
  NAND2X0_HVT U42 ( .A1(n246), .A2(n304), .Y(n563) );
  MUX41X1_HVT U51 ( .A1(n368), .A3(n326), .A2(n344), .A4(n345), .S0(n324), 
        .S1(n289), .Y(n556) );
  NAND2X0_HVT U53 ( .A1(n553), .A2(n562), .Y(n554) );
  NAND2X0_HVT U56 ( .A1(n307), .A2(n549), .Y(n550) );
  MUX41X1_HVT U57 ( .A1(n369), .A3(n585), .A2(n550), .A4(n594), .S0(n324), 
        .S1(n289), .Y(n548) );
  NAND2X0_HVT U58 ( .A1(n309), .A2(n602), .Y(n547) );
  MUX41X1_HVT U59 ( .A1(n284), .A3(n547), .A2(n282), .A4(n343), .S0(n324), 
        .S1(n289), .Y(n546) );
  MUX41X1_HVT U61 ( .A1(n280), .A3(n342), .A2(n341), .A4(n297), .S0(n324), 
        .S1(n289), .Y(n544) );
  NAND2X0_HVT U62 ( .A1(n316), .A2(n237), .Y(n543) );
  MUX41X1_HVT U63 ( .A1(n543), .A3(n333), .A2(n363), .A4(n340), .S0(n324), 
        .S1(n289), .Y(n542) );
  AO21X1_HVT U66 ( .A1(n338), .A2(n291), .A3(n362), .Y(n539) );
  MUX41X1_HVT U68 ( .A1(n336), .A3(n539), .A2(n538), .A4(n540), .S0(n285), 
        .S1(n273), .Y(n537) );
  MUX41X1_HVT U69 ( .A1(n537), .A3(n545), .A2(n541), .A4(n551), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n305), .A2(n532), .Y(n533) );
  MUX41X1_HVT U74 ( .A1(n534), .A3(n579), .A2(n533), .A4(n581), .S0(n287), 
        .S1(n322), .Y(n531) );
  MUX41X1_HVT U75 ( .A1(n366), .A3(n371), .A2(n232), .A4(n347), .S0(n285), 
        .S1(n322), .Y(n530) );
  MUX41X1_HVT U77 ( .A1(n596), .A3(n373), .A2(n529), .A4(n372), .S0(n292), 
        .S1(n317), .Y(n528) );
  MUX41X1_HVT U78 ( .A1(n528), .A3(n531), .A2(n530), .A4(n535), .S0(in[0]), 
        .S1(n289), .Y(n527) );
  MUX41X1_HVT U82 ( .A1(n560), .A3(n345), .A2(n327), .A4(n590), .S0(n285), 
        .S1(n273), .Y(n522) );
  AND2X1_HVT U83 ( .A1(n314), .A2(n274), .Y(n521) );
  MUX41X1_HVT U84 ( .A1(n346), .A3(n598), .A2(n588), .A4(n521), .S0(n285), 
        .S1(n321), .Y(n520) );
  NAND2X0_HVT U85 ( .A1(n316), .A2(n383), .Y(n519) );
  MUX41X1_HVT U86 ( .A1(n371), .A3(n519), .A2(n281), .A4(n277), .S0(n285), 
        .S1(n273), .Y(n518) );
  MUX41X1_HVT U87 ( .A1(n518), .A3(n522), .A2(n520), .A4(n523), .S0(n303), 
        .S1(in[5]), .Y(n517) );
  AO21X1_HVT U93 ( .A1(n294), .A2(n511), .A3(n367), .Y(n512) );
  MUX41X1_HVT U96 ( .A1(n327), .A3(n279), .A2(n370), .A4(n509), .S0(n285), 
        .S1(n273), .Y(n508) );
  MUX41X1_HVT U97 ( .A1(n366), .A3(n279), .A2(n310), .A4(n589), .S0(n285), 
        .S1(n321), .Y(n507) );
  NAND2X0_HVT U101 ( .A1(n502), .A2(n501), .Y(n503) );
  MUX41X1_HVT U103 ( .A1(n602), .A3(n337), .A2(n255), .A4(n570), .S0(n285), 
        .S1(n273), .Y(n499) );
  MUX41X1_HVT U105 ( .A1(n349), .A3(n558), .A2(n498), .A4(n365), .S0(n285), 
        .S1(n322), .Y(n497) );
  OA21X1_HVT U109 ( .A1(n356), .A2(n319), .A3(n343), .Y(n494) );
  NAND2X0_HVT U110 ( .A1(n236), .A2(n492), .Y(n493) );
  MUX41X1_HVT U114 ( .A1(n489), .A3(n495), .A2(n491), .A4(n494), .S0(n291), 
        .S1(n273), .Y(n488) );
  AND2X1_HVT U115 ( .A1(n246), .A2(n297), .Y(n487) );
  NAND2X0_HVT U123 ( .A1(n478), .A2(n477), .Y(n479) );
  MUX41X1_HVT U125 ( .A1(n583), .A3(n284), .A2(n336), .A4(n375), .S0(n286), 
        .S1(n324), .Y(n475) );
  AND3X1_HVT U128 ( .A1(n288), .A2(n316), .A3(n274), .Y(n472) );
  MUX41X1_HVT U131 ( .A1(n470), .A3(n472), .A2(n471), .A4(n473), .S0(n291), 
        .S1(n324), .Y(n469) );
  MUX41X1_HVT U135 ( .A1(n376), .A3(n381), .A2(n599), .A4(n578), .S0(n285), 
        .S1(n323), .Y(n466) );
  MUX41X1_HVT U136 ( .A1(n277), .A3(n572), .A2(n377), .A4(n569), .S0(n286), 
        .S1(n324), .Y(n465) );
  MUX41X1_HVT U139 ( .A1(n463), .A3(n466), .A2(n465), .A4(n467), .S0(n302), 
        .S1(n320), .Y(n462) );
  AND2X1_HVT U140 ( .A1(n595), .A2(n315), .Y(n461) );
  MUX41X1_HVT U141 ( .A1(n580), .A3(n357), .A2(n461), .A4(n353), .S0(n287), 
        .S1(n323), .Y(n460) );
  MUX41X1_HVT U142 ( .A1(n346), .A3(n297), .A2(n364), .A4(n595), .S0(n286), 
        .S1(n323), .Y(n459) );
  NAND2X0_HVT U146 ( .A1(n247), .A2(n309), .Y(n532) );
  MUX41X1_HVT U147 ( .A1(n377), .A3(n532), .A2(n366), .A4(n559), .S0(n259), 
        .S1(n324), .Y(n455) );
  OA21X1_HVT U151 ( .A1(n565), .A2(n267), .A3(n451), .Y(n452) );
  MUX41X1_HVT U153 ( .A1(n493), .A3(n280), .A2(n235), .A4(n329), .S0(n286), 
        .S1(n321), .Y(n449) );
  AND2X1_HVT U154 ( .A1(n294), .A2(n304), .Y(n448) );
  NAND2X0_HVT U158 ( .A1(n314), .A2(n383), .Y(n444) );
  MUX41X1_HVT U159 ( .A1(n50), .A3(n297), .A2(n444), .A4(n335), .S0(n317), 
        .S1(n322), .Y(n443) );
  MUX41X1_HVT U160 ( .A1(n443), .A3(n449), .A2(n445), .A4(n450), .S0(n302), 
        .S1(n290), .Y(n442) );
  AND2X1_HVT U162 ( .A1(n598), .A2(n532), .Y(n440) );
  MUX41X1_HVT U163 ( .A1(n342), .A3(n440), .A2(n278), .A4(n441), .S0(n317), 
        .S1(n321), .Y(n439) );
  MUX41X1_HVT U165 ( .A1(n583), .A3(n350), .A2(n559), .A4(n438), .S0(n324), 
        .S1(n318), .Y(n437) );
  NAND2X0_HVT U166 ( .A1(n309), .A2(n549), .Y(n436) );
  NAND2X0_HVT U167 ( .A1(n233), .A2(n316), .Y(n435) );
  MUX41X1_HVT U168 ( .A1(n369), .A3(n595), .A2(n435), .A4(n436), .S0(n318), 
        .S1(n322), .Y(n434) );
  MUX41X1_HVT U172 ( .A1(n431), .A3(n437), .A2(n434), .A4(n439), .S0(n303), 
        .S1(n320), .Y(n430) );
  NAND2X0_HVT U174 ( .A1(n310), .A2(n598), .Y(n591) );
  MUX41X1_HVT U176 ( .A1(n300), .A3(n429), .A2(n374), .A4(n591), .S0(n324), 
        .S1(n318), .Y(n428) );
  NAND2X0_HVT U177 ( .A1(n247), .A2(n301), .Y(n427) );
  MUX41X1_HVT U178 ( .A1(n587), .A3(n427), .A2(n378), .A4(n567), .S0(n259), 
        .S1(n321), .Y(n426) );
  MUX41X1_HVT U179 ( .A1(n577), .A3(n379), .A2(n331), .A4(n378), .S0(n318), 
        .S1(n321), .Y(n425) );
  MUX41X1_HVT U180 ( .A1(n334), .A3(n596), .A2(n50), .A4(n276), .S0(n292), 
        .S1(n318), .Y(n424) );
  MUX41X1_HVT U181 ( .A1(n424), .A3(n426), .A2(n425), .A4(n428), .S0(n302), 
        .S1(n290), .Y(n423) );
  OA21X1_HVT U184 ( .A1(n571), .A2(n258), .A3(n346), .Y(n420) );
  MUX41X1_HVT U186 ( .A1(n279), .A3(n566), .A2(n532), .A4(n559), .S0(n318), 
        .S1(n321), .Y(n418) );
  MUX41X1_HVT U189 ( .A1(n416), .A3(n591), .A2(n417), .A4(n365), .S0(n292), 
        .S1(n318), .Y(n415) );
  MUX41X1_HVT U190 ( .A1(n415), .A3(n418), .A2(n419), .A4(n422), .S0(n290), 
        .S1(n303), .Y(n414) );
  MUX41X1_HVT U195 ( .A1(n598), .A3(n370), .A2(n604), .A4(n568), .S0(n317), 
        .S1(n273), .Y(n410) );
  AO21X1_HVT U197 ( .A1(n281), .A2(n293), .A3(n367), .Y(n408) );
  NAND2X0_HVT U208 ( .A1(n310), .A2(n307), .Y(n492) );
  NAND2X0_HVT U212 ( .A1(n314), .A2(n305), .Y(n549) );
  NAND2X0_HVT U214 ( .A1(n598), .A2(n316), .Y(n398) );
  NAND2X0_HVT U215 ( .A1(n492), .A2(n305), .Y(n397) );
  AO21X1_HVT U216 ( .A1(n315), .A2(n381), .A3(n258), .Y(n502) );
  NAND2X0_HVT U218 ( .A1(n381), .A2(n313), .Y(n451) );
  NAND2X0_HVT U220 ( .A1(n293), .A2(n398), .Y(n524) );
  MUX21X2_HVT U1 ( .A1(n236), .A2(n298), .S0(n310), .Y(n564) );
  XOR2X1_HVT U2 ( .A1(n267), .A2(n578), .Y(n561) );
  MUX41X1_HVT U3 ( .A1(n510), .A3(n507), .A2(n515), .A4(n508), .S0(n23), .S1(
        n320), .Y(n506) );
  IBUFFX16_HVT U6 ( .A(n302), .Y(n23) );
  INVX0_HVT U7 ( .A(n592), .Y(n48) );
  INVX1_HVT U8 ( .A(n48), .Y(n50) );
  NAND2X0_HVT U9 ( .A1(n408), .A2(n210), .Y(n211) );
  NAND2X0_HVT U10 ( .A1(n409), .A2(n218), .Y(n212) );
  NAND2X0_HVT U11 ( .A1(n211), .A2(n212), .Y(n407) );
  INVX0_HVT U12 ( .A(n218), .Y(n210) );
  MUX21X1_HVT U14 ( .A1(n361), .A2(n378), .S0(n293), .Y(n409) );
  IBUFFX2_HVT U16 ( .A(n287), .Y(n218) );
  IBUFFX2_HVT U17 ( .A(n50), .Y(n363) );
  MUX21X1_HVT U18 ( .A1(n235), .A2(n514), .S0(n283), .Y(n513) );
  XNOR2X2_HVT U19 ( .A1(n272), .A2(n246), .Y(n283) );
  MUX21X1_HVT U20 ( .A1(n512), .A2(n513), .S0(n285), .Y(n510) );
  XOR2X2_HVT U22 ( .A1(n598), .A2(n314), .Y(n559) );
  MUX41X1_HVT U23 ( .A1(n410), .A3(n412), .A2(n407), .A4(n411), .S0(n213), 
        .S1(n216), .Y(n406) );
  IBUFFX16_HVT U25 ( .A(n244), .Y(n213) );
  IBUFFX16_HVT U26 ( .A(n290), .Y(n216) );
  IBUFFX2_HVT U27 ( .A(n315), .Y(n313) );
  MUX41X1_HVT U28 ( .A1(n354), .A3(n582), .A2(n550), .A4(n592), .S0(n217), 
        .S1(n268), .Y(n401) );
  IBUFFX16_HVT U29 ( .A(n250), .Y(n217) );
  IBUFFX2_HVT U30 ( .A(n568), .Y(n356) );
  IBUFFX2_HVT U31 ( .A(n549), .Y(n366) );
  AND3X2_HVT U32 ( .A1(n236), .A2(n549), .A3(n524), .Y(n525) );
  INVX2_HVT U34 ( .A(n242), .Y(n598) );
  DELLN1X2_HVT U36 ( .A(in[2]), .Y(n285) );
  MUX21X1_HVT U37 ( .A1(n561), .A2(n536), .S0(n287), .Y(n535) );
  MUX21X1_HVT U38 ( .A1(n420), .A2(n421), .S0(n287), .Y(n419) );
  MUX21X1_HVT U39 ( .A1(n278), .A2(n341), .S0(n286), .Y(n471) );
  IBUFFX2_HVT U40 ( .A(n315), .Y(n311) );
  IBUFFX16_HVT U41 ( .A(n325), .Y(n324) );
  INVX2_HVT U43 ( .A(n325), .Y(n323) );
  INVX2_HVT U44 ( .A(in[7]), .Y(n325) );
  INVX1_HVT U45 ( .A(n315), .Y(n246) );
  MUX21X1_HVT U46 ( .A1(n454), .A2(n462), .S0(in[6]), .Y(out[4]) );
  INVX1_HVT U47 ( .A(n384), .Y(n219) );
  INVX1_HVT U48 ( .A(n384), .Y(n231) );
  INVX1_HVT U49 ( .A(n219), .Y(n232) );
  INVX1_HVT U50 ( .A(n231), .Y(n233) );
  IBUFFX2_HVT U52 ( .A(n603), .Y(n234) );
  INVX1_HVT U54 ( .A(n234), .Y(n235) );
  INVX0_HVT U55 ( .A(n234), .Y(n236) );
  INVX0_HVT U60 ( .A(n234), .Y(n237) );
  NAND2X0_HVT U64 ( .A1(n496), .A2(n238), .Y(n239) );
  NAND2X0_HVT U65 ( .A1(n506), .A2(in[6]), .Y(n240) );
  NAND2X2_HVT U67 ( .A1(n239), .A2(n240), .Y(out[2]) );
  IBUFFX2_HVT U70 ( .A(in[6]), .Y(n238) );
  INVX1_HVT U71 ( .A(n308), .Y(n384) );
  INVX0_HVT U72 ( .A(n595), .Y(n381) );
  AO21X1_HVT U76 ( .A1(n287), .A2(n595), .A3(n598), .Y(n484) );
  NAND2X2_HVT U79 ( .A1(in[4]), .A2(n295), .Y(n595) );
  MUX41X1_HVT U80 ( .A1(n368), .A3(n516), .A2(n559), .A4(n563), .S0(n286), 
        .S1(n241), .Y(n515) );
  IBUFFX16_HVT U81 ( .A(n322), .Y(n241) );
  INVX0_HVT U88 ( .A(n312), .Y(n243) );
  IBUFFX2_HVT U89 ( .A(n315), .Y(n247) );
  XNOR2X1_HVT U90 ( .A1(n300), .A2(in[3]), .Y(n242) );
  INVX0_HVT U91 ( .A(n588), .Y(n341) );
  NBUFFX4_HVT U92 ( .A(n242), .Y(n299) );
  MUX21X2_HVT U94 ( .A1(n383), .A2(n299), .S0(n243), .Y(n597) );
  IBUFFX16_HVT U95 ( .A(n303), .Y(n244) );
  MUX41X1_HVT U98 ( .A1(n403), .A3(n401), .A2(n402), .A4(n400), .S0(n269), 
        .S1(n245), .Y(n399) );
  IBUFFX16_HVT U99 ( .A(n290), .Y(n245) );
  INVX0_HVT U100 ( .A(n597), .Y(n336) );
  MUX21X2_HVT U102 ( .A1(n298), .A2(n296), .S0(n247), .Y(n588) );
  NAND2X2_HVT U104 ( .A1(n246), .A2(n235), .Y(n602) );
  MUX21X2_HVT U106 ( .A1(n232), .A2(n383), .S0(n311), .Y(n578) );
  MUX21X1_HVT U107 ( .A1(n235), .A2(n490), .S0(n275), .Y(n489) );
  NBUFFX16_HVT U108 ( .A(n385), .Y(n300) );
  IBUFFX2_HVT U111 ( .A(n315), .Y(n314) );
  MUX21X1_HVT U112 ( .A1(n373), .A2(n567), .S0(n272), .Y(n446) );
  MUX21X1_HVT U113 ( .A1(n358), .A2(n582), .S0(n272), .Y(n464) );
  NAND2X0_HVT U116 ( .A1(n479), .A2(n252), .Y(n253) );
  MUX21X1_HVT U117 ( .A1(n601), .A2(n464), .S0(n250), .Y(n463) );
  MUX21X1_HVT U118 ( .A1(n475), .A2(n476), .S0(n291), .Y(n474) );
  INVX1_HVT U119 ( .A(n273), .Y(n268) );
  OA21X1_HVT U120 ( .A1(n597), .A2(n267), .A3(n357), .Y(n404) );
  INVX1_HVT U121 ( .A(n292), .Y(n272) );
  INVX0_HVT U122 ( .A(n321), .Y(n258) );
  INVX1_HVT U124 ( .A(n322), .Y(n267) );
  INVX1_HVT U126 ( .A(in[2]), .Y(n319) );
  NAND2X0_HVT U127 ( .A1(n265), .A2(n266), .Y(out[6]) );
  INVX1_HVT U129 ( .A(in[4]), .Y(n385) );
  INVX1_HVT U130 ( .A(n267), .Y(n252) );
  INVX1_HVT U132 ( .A(n320), .Y(n251) );
  INVX1_HVT U133 ( .A(n302), .Y(n269) );
  INVX0_HVT U134 ( .A(n287), .Y(n250) );
  INVX1_HVT U137 ( .A(n319), .Y(n259) );
  INVX0_HVT U138 ( .A(in[6]), .Y(n264) );
  INVX1_HVT U143 ( .A(n300), .Y(n274) );
  IBUFFX2_HVT U144 ( .A(n315), .Y(n312) );
  NAND2X0_HVT U145 ( .A1(n458), .A2(n250), .Y(n248) );
  NAND2X0_HVT U148 ( .A1(n457), .A2(n288), .Y(n249) );
  NAND2X0_HVT U149 ( .A1(n248), .A2(n249), .Y(n456) );
  MUX21X1_HVT U150 ( .A1(n332), .A2(n576), .S0(n267), .Y(n458) );
  OA21X2_HVT U152 ( .A1(n330), .A2(n258), .A3(n574), .Y(n457) );
  INVX1_HVT U155 ( .A(n255), .Y(n576) );
  OA21X1_HVT U156 ( .A1(n282), .A2(n258), .A3(n574), .Y(n432) );
  MUX21X2_HVT U157 ( .A1(n526), .A2(n525), .S0(n259), .Y(n523) );
  IBUFFX2_HVT U161 ( .A(n584), .Y(n345) );
  MUX21X2_HVT U164 ( .A1(n447), .A2(n446), .S0(n250), .Y(n445) );
  MUX41X1_HVT U169 ( .A1(n456), .A3(n460), .A2(n455), .A4(n459), .S0(n303), 
        .S1(n251), .Y(n454) );
  NAND2X0_HVT U170 ( .A1(n480), .A2(n267), .Y(n254) );
  NAND2X0_HVT U171 ( .A1(n253), .A2(n254), .Y(n476) );
  MUX21X2_HVT U173 ( .A1(n453), .A2(n452), .S0(n250), .Y(n450) );
  MUX21X1_HVT U175 ( .A1(n574), .A2(n493), .S0(n286), .Y(n491) );
  MUX21X1_HVT U182 ( .A1(n274), .A2(n306), .S0(n314), .Y(n255) );
  INVX0_HVT U183 ( .A(n567), .Y(n357) );
  IBUFFX2_HVT U185 ( .A(n582), .Y(n346) );
  INVX0_HVT U187 ( .A(n573), .Y(n353) );
  NAND2X0_HVT U188 ( .A1(n399), .A2(n264), .Y(n256) );
  NAND2X0_HVT U191 ( .A1(n406), .A2(in[6]), .Y(n257) );
  NAND2X0_HVT U192 ( .A1(n256), .A2(n257), .Y(out[7]) );
  MUX41X1_HVT U193 ( .A1(n593), .A3(n573), .A2(n569), .A4(n359), .S0(n317), 
        .S1(n258), .Y(n402) );
  MUX41X1_HVT U194 ( .A1(n352), .A3(n379), .A2(n602), .A4(n274), .S0(n250), 
        .S1(n272), .Y(n400) );
  INVX1_HVT U196 ( .A(n387), .Y(n378) );
  MUX21X2_HVT U198 ( .A1(n305), .A2(n584), .S0(n272), .Y(n526) );
  MUX41X1_HVT U199 ( .A1(n488), .A3(n474), .A2(n482), .A4(n469), .S0(n264), 
        .S1(n269), .Y(out[3]) );
  MUX41X1_HVT U200 ( .A1(n564), .A3(n578), .A2(n376), .A4(n595), .S0(n252), 
        .S1(n259), .Y(n411) );
  MUX21X1_HVT U201 ( .A1(n483), .A2(n486), .S0(n291), .Y(n482) );
  NAND2X0_HVT U202 ( .A1(n280), .A2(n260), .Y(n261) );
  NAND2X0_HVT U203 ( .A1(n505), .A2(n263), .Y(n262) );
  NAND2X0_HVT U204 ( .A1(n261), .A2(n262), .Y(n504) );
  INVX0_HVT U205 ( .A(n263), .Y(n260) );
  IBUFFX2_HVT U206 ( .A(n564), .Y(n360) );
  XOR2X1_HVT U207 ( .A1(n317), .A2(n323), .Y(n263) );
  INVX0_HVT U209 ( .A(n574), .Y(n352) );
  NAND2X0_HVT U210 ( .A1(n414), .A2(n264), .Y(n265) );
  NAND2X0_HVT U211 ( .A1(n423), .A2(in[6]), .Y(n266) );
  MUX41X1_HVT U213 ( .A1(n413), .A3(n557), .A2(n570), .A4(n563), .S0(n250), 
        .S1(n267), .Y(n412) );
  NAND2X0_HVT U217 ( .A1(n276), .A2(n252), .Y(n270) );
  NAND2X0_HVT U219 ( .A1(n588), .A2(n272), .Y(n271) );
  NAND2X0_HVT U221 ( .A1(n270), .A2(n271), .Y(n405) );
  MUX21X2_HVT U222 ( .A1(n405), .A2(n404), .S0(n250), .Y(n403) );
  MUX41X1_HVT U223 ( .A1(n574), .A3(n347), .A2(n487), .A4(n50), .S0(n319), 
        .S1(n267), .Y(n486) );
  MUX21X2_HVT U224 ( .A1(n328), .A2(n481), .S0(n259), .Y(n480) );
  IBUFFX2_HVT U225 ( .A(in[1]), .Y(n316) );
  MUX21X2_HVT U226 ( .A1(n517), .A2(n527), .S0(in[6]), .Y(out[1]) );
  INVX2_HVT U227 ( .A(in[1]), .Y(n315) );
  NBUFFX2_HVT U228 ( .A(in[2]), .Y(n286) );
  IBUFFX2_HVT U229 ( .A(n325), .Y(n321) );
  IBUFFX2_HVT U230 ( .A(n325), .Y(n322) );
  IBUFFX2_HVT U231 ( .A(n325), .Y(n273) );
  INVX1_HVT U232 ( .A(n319), .Y(n317) );
  IBUFFX2_HVT U233 ( .A(n319), .Y(n318) );
  MUX41X1_HVT U234 ( .A1(n348), .A3(n360), .A2(n306), .A4(n358), .S0(n325), 
        .S1(n319), .Y(n422) );
  MUX41X1_HVT U235 ( .A1(n504), .A3(n499), .A2(n500), .A4(n497), .S0(n269), 
        .S1(n251), .Y(n496) );
  XNOR2X1_HVT U236 ( .A1(n315), .A2(n319), .Y(n275) );
  IBUFFX2_HVT U237 ( .A(n315), .Y(n310) );
  MUX21X2_HVT U238 ( .A1(n430), .A2(n442), .S0(in[6]), .Y(out[5]) );
  INVX0_HVT U239 ( .A(in[3]), .Y(n382) );
  INVX1_HVT U240 ( .A(n306), .Y(n380) );
  NBUFFX2_HVT U241 ( .A(n242), .Y(n298) );
  NBUFFX2_HVT U242 ( .A(n242), .Y(n297) );
  AND2X1_HVT U243 ( .A1(n299), .A2(n549), .Y(n276) );
  NBUFFX2_HVT U244 ( .A(n600), .Y(n306) );
  MUX21X1_HVT U245 ( .A1(n380), .A2(n383), .S0(n291), .Y(n553) );
  NBUFFX2_HVT U246 ( .A(n600), .Y(n307) );
  MUX21X1_HVT U247 ( .A1(n337), .A2(n381), .S0(n291), .Y(n538) );
  AND2X1_HVT U248 ( .A1(n235), .A2(n532), .Y(n277) );
  MUX21X1_HVT U249 ( .A1(n297), .A2(n301), .S0(n314), .Y(n501) );
  MUX21X1_HVT U250 ( .A1(n380), .A2(n233), .S0(n311), .Y(n429) );
  MUX21X1_HVT U251 ( .A1(n307), .A2(n598), .S0(n313), .Y(n568) );
  MUX21X1_HVT U252 ( .A1(n383), .A2(n298), .S0(n313), .Y(n441) );
  MUX21X1_HVT U253 ( .A1(n298), .A2(n380), .S0(n247), .Y(n509) );
  MUX21X1_HVT U254 ( .A1(n598), .A2(n381), .S0(n246), .Y(n389) );
  MUX21X1_HVT U255 ( .A1(n598), .A2(n233), .S0(n311), .Y(n580) );
  MUX21X1_HVT U256 ( .A1(n307), .A2(n305), .S0(n314), .Y(n516) );
  MUX21X1_HVT U257 ( .A1(n598), .A2(n301), .S0(n246), .Y(n529) );
  MUX21X1_HVT U258 ( .A1(n383), .A2(n380), .S0(n313), .Y(n567) );
  MUX21X1_HVT U259 ( .A1(n296), .A2(n232), .S0(n314), .Y(n565) );
  MUX21X1_HVT U260 ( .A1(n484), .A2(n485), .S0(n293), .Y(n483) );
  MUX21X1_HVT U261 ( .A1(n329), .A2(n354), .S0(n286), .Y(n485) );
  MUX21X1_HVT U262 ( .A1(n351), .A2(n468), .S0(n288), .Y(n467) );
  MUX21X1_HVT U263 ( .A1(n375), .A2(n305), .S0(n293), .Y(n468) );
  NAND2X0_HVT U264 ( .A1(n300), .A2(n295), .Y(n600) );
  MUX21X1_HVT U265 ( .A1(n380), .A2(n301), .S0(n314), .Y(n390) );
  MUX21X1_HVT U266 ( .A1(n295), .A2(n598), .S0(n310), .Y(n392) );
  NBUFFX2_HVT U267 ( .A(n603), .Y(n308) );
  MUX21X1_HVT U268 ( .A1(n383), .A2(n296), .S0(n246), .Y(n571) );
  MUX21X1_HVT U269 ( .A1(n381), .A2(n380), .S0(n247), .Y(n586) );
  MUX21X1_HVT U270 ( .A1(n301), .A2(n296), .S0(n312), .Y(n481) );
  MUX21X1_HVT U271 ( .A1(n295), .A2(n309), .S0(n313), .Y(n416) );
  MUX21X1_HVT U272 ( .A1(n604), .A2(n236), .S0(n310), .Y(n417) );
  INVX1_HVT U273 ( .A(n604), .Y(n383) );
  MUX21X1_HVT U274 ( .A1(n237), .A2(n305), .S0(n246), .Y(n590) );
  MUX21X1_HVT U275 ( .A1(n306), .A2(n309), .S0(n313), .Y(n511) );
  MUX21X1_HVT U276 ( .A1(n296), .A2(n383), .S0(n247), .Y(n594) );
  MUX21X1_HVT U277 ( .A1(n352), .A2(n590), .S0(n287), .Y(n505) );
  MUX21X1_HVT U278 ( .A1(n295), .A2(n301), .S0(n310), .Y(n413) );
  XOR2X1_HVT U279 ( .A1(n235), .A2(n311), .Y(n557) );
  XOR2X1_HVT U280 ( .A1(n246), .A2(n381), .Y(n560) );
  XNOR2X1_HVT U281 ( .A1(n306), .A2(n311), .Y(n278) );
  AND2X1_HVT U282 ( .A1(n312), .A2(n233), .Y(n279) );
  MUX21X1_HVT U283 ( .A1(n604), .A2(n305), .S0(n311), .Y(n574) );
  MUX21X1_HVT U284 ( .A1(n307), .A2(n296), .S0(n247), .Y(n593) );
  MUX21X1_HVT U285 ( .A1(n237), .A2(n301), .S0(n311), .Y(n396) );
  MUX21X1_HVT U286 ( .A1(n237), .A2(n307), .S0(n313), .Y(n388) );
  MUX21X1_HVT U287 ( .A1(n305), .A2(n296), .S0(n247), .Y(n394) );
  AND2X1_HVT U288 ( .A1(n309), .A2(n492), .Y(n280) );
  XNOR2X1_HVT U289 ( .A1(n604), .A2(n313), .Y(n281) );
  MUX21X1_HVT U290 ( .A1(n305), .A2(n301), .S0(n312), .Y(n534) );
  MUX21X1_HVT U291 ( .A1(n595), .A2(n309), .S0(n288), .Y(n478) );
  XOR2X1_HVT U292 ( .A1(n300), .A2(n246), .Y(n579) );
  NBUFFX2_HVT U293 ( .A(n382), .Y(n295) );
  NBUFFX2_HVT U294 ( .A(n323), .Y(n294) );
  NBUFFX2_HVT U295 ( .A(n323), .Y(n292) );
  NBUFFX2_HVT U296 ( .A(n323), .Y(n293) );
  NBUFFX2_HVT U297 ( .A(n382), .Y(n296) );
  NBUFFX2_HVT U298 ( .A(in[5]), .Y(n291) );
  NBUFFX2_HVT U299 ( .A(in[5]), .Y(n290) );
  NBUFFX2_HVT U300 ( .A(n317), .Y(n288) );
  NBUFFX2_HVT U301 ( .A(in[2]), .Y(n287) );
  NBUFFX2_HVT U302 ( .A(n320), .Y(n289) );
  MUX21X1_HVT U303 ( .A1(n299), .A2(n304), .S0(n312), .Y(n582) );
  MUX21X1_HVT U304 ( .A1(n503), .A2(n351), .S0(n288), .Y(n500) );
  MUX21X1_HVT U305 ( .A1(n519), .A2(n304), .S0(n293), .Y(n421) );
  MUX21X1_HVT U306 ( .A1(n542), .A2(n544), .S0(n287), .Y(n541) );
  XOR2X1_HVT U307 ( .A1(n312), .A2(in[3]), .Y(n558) );
  MUX21X1_HVT U308 ( .A1(n305), .A2(n299), .S0(n313), .Y(n498) );
  AND2X1_HVT U309 ( .A1(n299), .A2(n316), .Y(n282) );
  MUX21X1_HVT U310 ( .A1(n304), .A2(n380), .S0(n312), .Y(n566) );
  MUX21X1_HVT U311 ( .A1(n383), .A2(n370), .S0(n294), .Y(n536) );
  MUX21X1_HVT U312 ( .A1(n433), .A2(n432), .S0(n288), .Y(n431) );
  MUX21X1_HVT U313 ( .A1(n595), .A2(n370), .S0(n294), .Y(n433) );
  MUX21X1_HVT U314 ( .A1(n372), .A2(n381), .S0(n293), .Y(n453) );
  MUX21X1_HVT U315 ( .A1(n381), .A2(n232), .S0(n310), .Y(n438) );
  NAND2X0_HVT U316 ( .A1(n304), .A2(n301), .Y(n603) );
  NBUFFX2_HVT U317 ( .A(n385), .Y(n301) );
  MUX21X1_HVT U318 ( .A1(n232), .A2(n304), .S0(n314), .Y(n585) );
  MUX21X1_HVT U319 ( .A1(n355), .A2(n602), .S0(n259), .Y(n495) );
  MUX21X1_HVT U320 ( .A1(n448), .A2(n237), .S0(n283), .Y(n447) );
  MUX21X1_HVT U321 ( .A1(n587), .A2(n353), .S0(n259), .Y(n470) );
  MUX21X1_HVT U322 ( .A1(n602), .A2(n315), .S0(n287), .Y(n477) );
  MUX21X1_HVT U323 ( .A1(n554), .A2(n555), .S0(n292), .Y(n552) );
  MUX21X1_HVT U324 ( .A1(n304), .A2(n570), .S0(n291), .Y(n555) );
  XOR2X1_HVT U325 ( .A1(n312), .A2(n290), .Y(n562) );
  MUX21X1_HVT U326 ( .A1(n304), .A2(n381), .S0(n311), .Y(n393) );
  MUX21X1_HVT U327 ( .A1(n307), .A2(n304), .S0(n247), .Y(n596) );
  NBUFFX2_HVT U328 ( .A(n595), .Y(n305) );
  MUX21X1_HVT U329 ( .A1(n575), .A2(n397), .S0(n292), .Y(n391) );
  MUX21X1_HVT U330 ( .A1(n349), .A2(n575), .S0(n259), .Y(n473) );
  MUX21X1_HVT U331 ( .A1(n339), .A2(n316), .S0(n291), .Y(n540) );
  MUX21X1_HVT U332 ( .A1(n304), .A2(n301), .S0(n294), .Y(n514) );
  NBUFFX2_HVT U333 ( .A(n604), .Y(n309) );
  AND2X1_HVT U334 ( .A1(n296), .A2(n316), .Y(n284) );
  NBUFFX2_HVT U335 ( .A(in[5]), .Y(n320) );
  MUX21X1_HVT U336 ( .A1(n552), .A2(n556), .S0(n288), .Y(n551) );
  MUX21X1_HVT U337 ( .A1(n546), .A2(n548), .S0(n287), .Y(n545) );
  MUX21X1_HVT U338 ( .A1(n380), .A2(n274), .S0(n311), .Y(n573) );
  MUX21X1_HVT U339 ( .A1(n274), .A2(n598), .S0(n310), .Y(n395) );
  MUX21X1_HVT U340 ( .A1(n274), .A2(n383), .S0(n312), .Y(n569) );
  MUX21X1_HVT U341 ( .A1(n274), .A2(n381), .S0(n310), .Y(n587) );
  NAND2X0_HVT U342 ( .A1(in[3]), .A2(in[4]), .Y(n604) );
  MUX21X1_HVT U343 ( .A1(n274), .A2(n236), .S0(n310), .Y(n584) );
  MUX21X1_HVT U344 ( .A1(n309), .A2(n274), .S0(n312), .Y(n577) );
  MUX21X1_HVT U345 ( .A1(n304), .A2(n274), .S0(n286), .Y(n490) );
  MUX21X1_HVT U346 ( .A1(n274), .A2(n305), .S0(n314), .Y(n387) );
  MUX21X1_HVT U347 ( .A1(n274), .A2(n309), .S0(n313), .Y(n386) );
  MUX21X1_HVT U348 ( .A1(n296), .A2(n274), .S0(n247), .Y(n575) );
  NBUFFX2_HVT U349 ( .A(in[3]), .Y(n304) );
  NBUFFX2_HVT U350 ( .A(in[0]), .Y(n302) );
  NBUFFX2_HVT U351 ( .A(in[0]), .Y(n303) );
  INVX0_HVT U352 ( .A(n583), .Y(n326) );
  INVX0_HVT U353 ( .A(n581), .Y(n327) );
  INVX0_HVT U354 ( .A(n572), .Y(n328) );
  INVX0_HVT U355 ( .A(n570), .Y(n329) );
  INVX0_HVT U356 ( .A(n435), .Y(n330) );
  INVX0_HVT U357 ( .A(n398), .Y(n331) );
  INVX0_HVT U358 ( .A(n602), .Y(n332) );
  INVX0_HVT U359 ( .A(n589), .Y(n333) );
  INVX0_HVT U360 ( .A(n601), .Y(n334) );
  INVX0_HVT U361 ( .A(n599), .Y(n335) );
  INVX0_HVT U362 ( .A(n596), .Y(n337) );
  INVX0_HVT U363 ( .A(n594), .Y(n338) );
  INVX0_HVT U364 ( .A(n593), .Y(n339) );
  INVX0_HVT U365 ( .A(n590), .Y(n340) );
  INVX0_HVT U366 ( .A(n587), .Y(n342) );
  INVX0_HVT U367 ( .A(n586), .Y(n343) );
  INVX0_HVT U368 ( .A(n585), .Y(n344) );
  INVX0_HVT U369 ( .A(n580), .Y(n347) );
  INVX0_HVT U370 ( .A(n579), .Y(n348) );
  INVX0_HVT U371 ( .A(n577), .Y(n349) );
  INVX0_HVT U372 ( .A(n575), .Y(n350) );
  INVX0_HVT U373 ( .A(n391), .Y(n351) );
  INVX0_HVT U374 ( .A(n571), .Y(n354) );
  INVX0_HVT U375 ( .A(n569), .Y(n355) );
  INVX0_HVT U376 ( .A(n566), .Y(n358) );
  INVX0_HVT U377 ( .A(n565), .Y(n359) );
  INVX0_HVT U378 ( .A(n563), .Y(n361) );
  INVX0_HVT U379 ( .A(n532), .Y(n362) );
  INVX0_HVT U380 ( .A(n492), .Y(n364) );
  INVX0_HVT U381 ( .A(n397), .Y(n365) );
  INVX0_HVT U382 ( .A(n451), .Y(n367) );
  INVX0_HVT U383 ( .A(n396), .Y(n368) );
  INVX0_HVT U384 ( .A(n395), .Y(n369) );
  INVX0_HVT U385 ( .A(n394), .Y(n370) );
  INVX0_HVT U386 ( .A(n393), .Y(n371) );
  INVX0_HVT U387 ( .A(n392), .Y(n372) );
  INVX0_HVT U388 ( .A(n511), .Y(n373) );
  INVX0_HVT U389 ( .A(n501), .Y(n374) );
  INVX0_HVT U390 ( .A(n390), .Y(n375) );
  INVX0_HVT U391 ( .A(n389), .Y(n376) );
  INVX0_HVT U392 ( .A(n388), .Y(n377) );
  INVX0_HVT U393 ( .A(n386), .Y(n379) );
endmodule

