
module aes ( plaintext, key, clk, reset, start, cipher_text, ready );
  input [127:0] plaintext;
  input [127:0] key;
  output [127:0] cipher_text;
  input clk, reset, start;
  output ready;
  wire   n12, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305;
  wire   [127:0] adk_out0;
  wire   [127:0] adk_in;
  wire   [3:0] round_number;
  wire   [127:0] key_round;
  wire   [127:0] keyout;

  DFFASX1_HVT d_reg ( .D(n287), .CLK(clk), .SETB(n25), .Q(n2), .QN(n12) );
  DFFARX1_HVT \round_number_reg[3]  ( .D(n286), .CLK(clk), .RSTB(n14), .Q(
        round_number[3]) );
  DFFARX1_HVT \round_number_reg[0]  ( .D(n285), .CLK(clk), .RSTB(n15), .Q(
        round_number[0]), .QN(n3) );
  DFFARX1_HVT \round_number_reg[1]  ( .D(n284), .CLK(clk), .RSTB(n15), .Q(
        round_number[1]), .QN(n4) );
  DFFARX1_HVT \round_number_reg[2]  ( .D(n283), .CLK(clk), .RSTB(n14), .Q(
        round_number[2]), .QN(n1) );
  DFFARX1_HVT \key_round_reg[0]  ( .D(n282), .CLK(clk), .RSTB(n11), .Q(
        key_round[0]) );
  DFFARX1_HVT \adk_in_reg[0]  ( .D(n281), .CLK(clk), .RSTB(n24), .Q(adk_in[0])
         );
  DFFARX1_HVT \adk_in_reg[1]  ( .D(n280), .CLK(clk), .RSTB(n20), .Q(adk_in[1])
         );
  DFFARX1_HVT \adk_in_reg[2]  ( .D(n279), .CLK(clk), .RSTB(n20), .Q(adk_in[2])
         );
  DFFARX1_HVT \adk_in_reg[3]  ( .D(n278), .CLK(clk), .RSTB(n19), .Q(adk_in[3])
         );
  DFFARX1_HVT \adk_in_reg[4]  ( .D(n277), .CLK(clk), .RSTB(n20), .Q(adk_in[4])
         );
  DFFARX1_HVT \adk_in_reg[5]  ( .D(n276), .CLK(clk), .RSTB(n19), .Q(adk_in[5])
         );
  DFFARX1_HVT \adk_in_reg[6]  ( .D(n275), .CLK(clk), .RSTB(n21), .Q(adk_in[6])
         );
  DFFARX1_HVT \adk_in_reg[7]  ( .D(n274), .CLK(clk), .RSTB(n21), .Q(adk_in[7])
         );
  DFFARX1_HVT \adk_in_reg[8]  ( .D(n273), .CLK(clk), .RSTB(n17), .Q(adk_in[8])
         );
  DFFARX1_HVT \adk_in_reg[9]  ( .D(n272), .CLK(clk), .RSTB(n17), .Q(adk_in[9])
         );
  DFFARX1_HVT \adk_in_reg[10]  ( .D(n271), .CLK(clk), .RSTB(n17), .Q(
        adk_in[10]) );
  DFFARX1_HVT \adk_in_reg[11]  ( .D(n270), .CLK(clk), .RSTB(n18), .Q(
        adk_in[11]) );
  DFFARX1_HVT \adk_in_reg[12]  ( .D(n269), .CLK(clk), .RSTB(n17), .Q(
        adk_in[12]) );
  DFFARX1_HVT \adk_in_reg[13]  ( .D(n268), .CLK(clk), .RSTB(n17), .Q(
        adk_in[13]) );
  DFFARX1_HVT \adk_in_reg[14]  ( .D(n267), .CLK(clk), .RSTB(n17), .Q(
        adk_in[14]) );
  DFFARX1_HVT \adk_in_reg[15]  ( .D(n266), .CLK(clk), .RSTB(n18), .Q(
        adk_in[15]) );
  DFFARX1_HVT \adk_in_reg[16]  ( .D(n265), .CLK(clk), .RSTB(n24), .Q(
        adk_in[16]) );
  DFFARX1_HVT \adk_in_reg[17]  ( .D(n264), .CLK(clk), .RSTB(n23), .Q(
        adk_in[17]) );
  DFFARX1_HVT \adk_in_reg[18]  ( .D(n263), .CLK(clk), .RSTB(n22), .Q(
        adk_in[18]) );
  DFFARX1_HVT \adk_in_reg[19]  ( .D(n262), .CLK(clk), .RSTB(n9), .Q(adk_in[19]) );
  DFFARX1_HVT \adk_in_reg[20]  ( .D(n261), .CLK(clk), .RSTB(n22), .Q(
        adk_in[20]) );
  DFFARX1_HVT \adk_in_reg[21]  ( .D(n260), .CLK(clk), .RSTB(n23), .Q(
        adk_in[21]) );
  DFFARX1_HVT \adk_in_reg[22]  ( .D(n259), .CLK(clk), .RSTB(n23), .Q(
        adk_in[22]) );
  DFFARX1_HVT \adk_in_reg[23]  ( .D(n258), .CLK(clk), .RSTB(n24), .Q(
        adk_in[23]) );
  DFFARX1_HVT \adk_in_reg[24]  ( .D(n257), .CLK(clk), .RSTB(n15), .Q(
        adk_in[24]) );
  DFFARX1_HVT \adk_in_reg[25]  ( .D(n256), .CLK(clk), .RSTB(n15), .Q(
        adk_in[25]) );
  DFFARX1_HVT \adk_in_reg[26]  ( .D(n255), .CLK(clk), .RSTB(n20), .Q(
        adk_in[26]) );
  DFFARX1_HVT \adk_in_reg[27]  ( .D(n254), .CLK(clk), .RSTB(n15), .Q(
        adk_in[27]) );
  DFFARX1_HVT \adk_in_reg[28]  ( .D(n253), .CLK(clk), .RSTB(n15), .Q(
        adk_in[28]) );
  DFFARX1_HVT \adk_in_reg[29]  ( .D(n252), .CLK(clk), .RSTB(n15), .Q(
        adk_in[29]) );
  DFFARX1_HVT \adk_in_reg[30]  ( .D(n251), .CLK(clk), .RSTB(n15), .Q(
        adk_in[30]) );
  DFFARX1_HVT \adk_in_reg[31]  ( .D(n250), .CLK(clk), .RSTB(n15), .Q(
        adk_in[31]) );
  DFFARX1_HVT \adk_in_reg[32]  ( .D(n249), .CLK(clk), .RSTB(n24), .Q(
        adk_in[32]) );
  DFFARX1_HVT \adk_in_reg[33]  ( .D(n248), .CLK(clk), .RSTB(n20), .Q(
        adk_in[33]) );
  DFFARX1_HVT \adk_in_reg[34]  ( .D(n247), .CLK(clk), .RSTB(n21), .Q(
        adk_in[34]) );
  DFFARX1_HVT \adk_in_reg[35]  ( .D(n246), .CLK(clk), .RSTB(n19), .Q(
        adk_in[35]) );
  DFFARX1_HVT \adk_in_reg[36]  ( .D(n245), .CLK(clk), .RSTB(n20), .Q(
        adk_in[36]) );
  DFFARX1_HVT \adk_in_reg[37]  ( .D(n244), .CLK(clk), .RSTB(n19), .Q(
        adk_in[37]) );
  DFFARX1_HVT \adk_in_reg[38]  ( .D(n243), .CLK(clk), .RSTB(n20), .Q(
        adk_in[38]) );
  DFFARX1_HVT \adk_in_reg[39]  ( .D(n242), .CLK(clk), .RSTB(n21), .Q(
        adk_in[39]) );
  DFFARX1_HVT \adk_in_reg[40]  ( .D(n241), .CLK(clk), .RSTB(n22), .Q(
        adk_in[40]) );
  DFFARX1_HVT \adk_in_reg[41]  ( .D(n240), .CLK(clk), .RSTB(n15), .Q(
        adk_in[41]) );
  DFFARX1_HVT \adk_in_reg[42]  ( .D(n239), .CLK(clk), .RSTB(n22), .Q(
        adk_in[42]) );
  DFFARX1_HVT \adk_in_reg[43]  ( .D(n238), .CLK(clk), .RSTB(n19), .Q(
        adk_in[43]) );
  DFFARX1_HVT \adk_in_reg[44]  ( .D(n237), .CLK(clk), .RSTB(n21), .Q(
        adk_in[44]) );
  DFFARX1_HVT \adk_in_reg[45]  ( .D(n236), .CLK(clk), .RSTB(n21), .Q(
        adk_in[45]) );
  DFFARX1_HVT \adk_in_reg[46]  ( .D(n235), .CLK(clk), .RSTB(n21), .Q(
        adk_in[46]) );
  DFFARX1_HVT \adk_in_reg[47]  ( .D(n234), .CLK(clk), .RSTB(n22), .Q(
        adk_in[47]) );
  DFFARX1_HVT \adk_in_reg[48]  ( .D(n233), .CLK(clk), .RSTB(n23), .Q(
        adk_in[48]) );
  DFFARX1_HVT \adk_in_reg[49]  ( .D(n232), .CLK(clk), .RSTB(n23), .Q(
        adk_in[49]) );
  DFFARX1_HVT \adk_in_reg[50]  ( .D(n231), .CLK(clk), .RSTB(n24), .Q(
        adk_in[50]) );
  DFFARX1_HVT \adk_in_reg[51]  ( .D(n230), .CLK(clk), .RSTB(n18), .Q(
        adk_in[51]) );
  DFFARX1_HVT \adk_in_reg[52]  ( .D(n229), .CLK(clk), .RSTB(n23), .Q(
        adk_in[52]) );
  DFFARX1_HVT \adk_in_reg[53]  ( .D(n228), .CLK(clk), .RSTB(n22), .Q(
        adk_in[53]) );
  DFFARX1_HVT \adk_in_reg[54]  ( .D(n227), .CLK(clk), .RSTB(n23), .Q(
        adk_in[54]) );
  DFFARX1_HVT \adk_in_reg[55]  ( .D(n226), .CLK(clk), .RSTB(n24), .Q(
        adk_in[55]) );
  DFFARX1_HVT \adk_in_reg[56]  ( .D(n225), .CLK(clk), .RSTB(n18), .Q(
        adk_in[56]) );
  DFFARX1_HVT \adk_in_reg[57]  ( .D(n224), .CLK(clk), .RSTB(n18), .Q(
        adk_in[57]) );
  DFFARX1_HVT \adk_in_reg[58]  ( .D(n223), .CLK(clk), .RSTB(n18), .Q(
        adk_in[58]) );
  DFFARX1_HVT \adk_in_reg[59]  ( .D(n222), .CLK(clk), .RSTB(n19), .Q(
        adk_in[59]) );
  DFFARX1_HVT \adk_in_reg[60]  ( .D(n221), .CLK(clk), .RSTB(n18), .Q(
        adk_in[60]) );
  DFFARX1_HVT \adk_in_reg[61]  ( .D(n220), .CLK(clk), .RSTB(n18), .Q(
        adk_in[61]) );
  DFFARX1_HVT \adk_in_reg[62]  ( .D(n219), .CLK(clk), .RSTB(n18), .Q(
        adk_in[62]) );
  DFFARX1_HVT \adk_in_reg[63]  ( .D(n218), .CLK(clk), .RSTB(n19), .Q(
        adk_in[63]) );
  DFFARX1_HVT \adk_in_reg[64]  ( .D(n217), .CLK(clk), .RSTB(n24), .Q(
        adk_in[64]) );
  DFFARX1_HVT \adk_in_reg[65]  ( .D(n216), .CLK(clk), .RSTB(n20), .Q(
        adk_in[65]) );
  DFFARX1_HVT \adk_in_reg[66]  ( .D(n215), .CLK(clk), .RSTB(n19), .Q(
        adk_in[66]) );
  DFFARX1_HVT \adk_in_reg[67]  ( .D(n214), .CLK(clk), .RSTB(n19), .Q(
        adk_in[67]) );
  DFFARX1_HVT \adk_in_reg[68]  ( .D(n213), .CLK(clk), .RSTB(n20), .Q(
        adk_in[68]) );
  DFFARX1_HVT \adk_in_reg[69]  ( .D(n212), .CLK(clk), .RSTB(n19), .Q(
        adk_in[69]) );
  DFFARX1_HVT \adk_in_reg[70]  ( .D(n211), .CLK(clk), .RSTB(n20), .Q(
        adk_in[70]) );
  DFFARX1_HVT \adk_in_reg[71]  ( .D(n210), .CLK(clk), .RSTB(n21), .Q(
        adk_in[71]) );
  DFFARX1_HVT \adk_in_reg[72]  ( .D(n209), .CLK(clk), .RSTB(n17), .Q(
        adk_in[72]) );
  DFFARX1_HVT \adk_in_reg[73]  ( .D(n208), .CLK(clk), .RSTB(n17), .Q(
        adk_in[73]) );
  DFFARX1_HVT \adk_in_reg[74]  ( .D(n207), .CLK(clk), .RSTB(n15), .Q(
        adk_in[74]) );
  DFFARX1_HVT \adk_in_reg[75]  ( .D(n206), .CLK(clk), .RSTB(n17), .Q(
        adk_in[75]) );
  DFFARX1_HVT \adk_in_reg[76]  ( .D(n205), .CLK(clk), .RSTB(n17), .Q(
        adk_in[76]) );
  DFFARX1_HVT \adk_in_reg[77]  ( .D(n204), .CLK(clk), .RSTB(n18), .Q(
        adk_in[77]) );
  DFFARX1_HVT \adk_in_reg[78]  ( .D(n203), .CLK(clk), .RSTB(n17), .Q(
        adk_in[78]) );
  DFFARX1_HVT \adk_in_reg[79]  ( .D(n202), .CLK(clk), .RSTB(n18), .Q(
        adk_in[79]) );
  DFFARX1_HVT \adk_in_reg[80]  ( .D(n201), .CLK(clk), .RSTB(n23), .Q(
        adk_in[80]) );
  DFFARX1_HVT \adk_in_reg[81]  ( .D(n200), .CLK(clk), .RSTB(n22), .Q(
        adk_in[81]) );
  DFFARX1_HVT \adk_in_reg[82]  ( .D(n199), .CLK(clk), .RSTB(n23), .Q(
        adk_in[82]) );
  DFFARX1_HVT \adk_in_reg[83]  ( .D(n198), .CLK(clk), .RSTB(n18), .Q(
        adk_in[83]) );
  DFFARX1_HVT \adk_in_reg[84]  ( .D(n197), .CLK(clk), .RSTB(n23), .Q(
        adk_in[84]) );
  DFFARX1_HVT \adk_in_reg[85]  ( .D(n196), .CLK(clk), .RSTB(n22), .Q(
        adk_in[85]) );
  DFFARX1_HVT \adk_in_reg[86]  ( .D(n195), .CLK(clk), .RSTB(n24), .Q(
        adk_in[86]) );
  DFFARX1_HVT \adk_in_reg[87]  ( .D(n194), .CLK(clk), .RSTB(n24), .Q(
        adk_in[87]) );
  DFFARX1_HVT \adk_in_reg[88]  ( .D(n193), .CLK(clk), .RSTB(n16), .Q(
        adk_in[88]) );
  DFFARX1_HVT \adk_in_reg[89]  ( .D(n192), .CLK(clk), .RSTB(n15), .Q(
        adk_in[89]) );
  DFFARX1_HVT \adk_in_reg[90]  ( .D(n191), .CLK(clk), .RSTB(n17), .Q(
        adk_in[90]) );
  DFFARX1_HVT \adk_in_reg[91]  ( .D(n190), .CLK(clk), .RSTB(n16), .Q(
        adk_in[91]) );
  DFFARX1_HVT \adk_in_reg[92]  ( .D(n189), .CLK(clk), .RSTB(n16), .Q(
        adk_in[92]) );
  DFFARX1_HVT \adk_in_reg[93]  ( .D(n188), .CLK(clk), .RSTB(n16), .Q(
        adk_in[93]) );
  DFFARX1_HVT \adk_in_reg[94]  ( .D(n187), .CLK(clk), .RSTB(n16), .Q(
        adk_in[94]) );
  DFFARX1_HVT \adk_in_reg[95]  ( .D(n186), .CLK(clk), .RSTB(n17), .Q(
        adk_in[95]) );
  DFFARX1_HVT \adk_in_reg[96]  ( .D(n185), .CLK(clk), .RSTB(n24), .Q(
        adk_in[96]) );
  DFFARX1_HVT \adk_in_reg[97]  ( .D(n184), .CLK(clk), .RSTB(n21), .Q(
        adk_in[97]) );
  DFFARX1_HVT \adk_in_reg[98]  ( .D(n183), .CLK(clk), .RSTB(n19), .Q(
        adk_in[98]) );
  DFFARX1_HVT \adk_in_reg[99]  ( .D(n182), .CLK(clk), .RSTB(n19), .Q(
        adk_in[99]) );
  DFFARX1_HVT \adk_in_reg[100]  ( .D(n181), .CLK(clk), .RSTB(n20), .Q(
        adk_in[100]) );
  DFFARX1_HVT \adk_in_reg[101]  ( .D(n180), .CLK(clk), .RSTB(n20), .Q(
        adk_in[101]) );
  DFFARX1_HVT \adk_in_reg[102]  ( .D(n179), .CLK(clk), .RSTB(n20), .Q(
        adk_in[102]) );
  DFFARX1_HVT \adk_in_reg[103]  ( .D(n178), .CLK(clk), .RSTB(n21), .Q(
        adk_in[103]) );
  DFFARX1_HVT \adk_in_reg[104]  ( .D(n177), .CLK(clk), .RSTB(n22), .Q(
        adk_in[104]) );
  DFFARX1_HVT \adk_in_reg[105]  ( .D(n176), .CLK(clk), .RSTB(n21), .Q(
        adk_in[105]) );
  DFFARX1_HVT \adk_in_reg[106]  ( .D(n175), .CLK(clk), .RSTB(n21), .Q(
        adk_in[106]) );
  DFFARX1_HVT \adk_in_reg[107]  ( .D(n174), .CLK(clk), .RSTB(n15), .Q(
        adk_in[107]) );
  DFFARX1_HVT \adk_in_reg[108]  ( .D(n173), .CLK(clk), .RSTB(n19), .Q(
        adk_in[108]) );
  DFFARX1_HVT \adk_in_reg[109]  ( .D(n172), .CLK(clk), .RSTB(n21), .Q(
        adk_in[109]) );
  DFFARX1_HVT \adk_in_reg[110]  ( .D(n171), .CLK(clk), .RSTB(n22), .Q(
        adk_in[110]) );
  DFFARX1_HVT \adk_in_reg[111]  ( .D(n170), .CLK(clk), .RSTB(n22), .Q(
        adk_in[111]) );
  DFFARX1_HVT \adk_in_reg[112]  ( .D(n169), .CLK(clk), .RSTB(n24), .Q(
        adk_in[112]) );
  DFFARX1_HVT \adk_in_reg[113]  ( .D(n168), .CLK(clk), .RSTB(n22), .Q(
        adk_in[113]) );
  DFFARX1_HVT \adk_in_reg[114]  ( .D(n167), .CLK(clk), .RSTB(n23), .Q(
        adk_in[114]) );
  DFFARX1_HVT \adk_in_reg[115]  ( .D(n166), .CLK(clk), .RSTB(n18), .Q(
        adk_in[115]) );
  DFFARX1_HVT \adk_in_reg[116]  ( .D(n165), .CLK(clk), .RSTB(n22), .Q(
        adk_in[116]) );
  DFFARX1_HVT \adk_in_reg[117]  ( .D(n164), .CLK(clk), .RSTB(n23), .Q(
        adk_in[117]) );
  DFFARX1_HVT \adk_in_reg[118]  ( .D(n163), .CLK(clk), .RSTB(n23), .Q(
        adk_in[118]) );
  DFFARX1_HVT \adk_in_reg[119]  ( .D(n162), .CLK(clk), .RSTB(n24), .Q(
        adk_in[119]) );
  DFFARX1_HVT \adk_in_reg[120]  ( .D(n161), .CLK(clk), .RSTB(n16), .Q(
        adk_in[120]) );
  DFFARX1_HVT \adk_in_reg[121]  ( .D(n160), .CLK(clk), .RSTB(n16), .Q(
        adk_in[121]) );
  DFFARX1_HVT \adk_in_reg[122]  ( .D(n159), .CLK(clk), .RSTB(n16), .Q(
        adk_in[122]) );
  DFFARX1_HVT \adk_in_reg[123]  ( .D(n158), .CLK(clk), .RSTB(n16), .Q(
        adk_in[123]) );
  DFFARX1_HVT \adk_in_reg[124]  ( .D(n157), .CLK(clk), .RSTB(n16), .Q(
        adk_in[124]) );
  DFFARX1_HVT \adk_in_reg[125]  ( .D(n156), .CLK(clk), .RSTB(n16), .Q(
        adk_in[125]) );
  DFFARX1_HVT \adk_in_reg[126]  ( .D(n155), .CLK(clk), .RSTB(n16), .Q(
        adk_in[126]) );
  DFFARX1_HVT \adk_in_reg[127]  ( .D(n154), .CLK(clk), .RSTB(n16), .Q(
        adk_in[127]) );
  DFFARX1_HVT \key_round_reg[1]  ( .D(n153), .CLK(clk), .RSTB(n10), .Q(
        key_round[1]) );
  DFFARX1_HVT \key_round_reg[2]  ( .D(n152), .CLK(clk), .RSTB(n13), .Q(
        key_round[2]) );
  DFFARX1_HVT \key_round_reg[3]  ( .D(n151), .CLK(clk), .RSTB(n8), .Q(
        key_round[3]) );
  DFFARX1_HVT \key_round_reg[4]  ( .D(n150), .CLK(clk), .RSTB(n5), .Q(
        key_round[4]) );
  DFFARX1_HVT \key_round_reg[5]  ( .D(n149), .CLK(clk), .RSTB(n7), .Q(
        key_round[5]) );
  DFFARX1_HVT \key_round_reg[6]  ( .D(n148), .CLK(clk), .RSTB(n25), .Q(
        key_round[6]) );
  DFFARX1_HVT \key_round_reg[7]  ( .D(n147), .CLK(clk), .RSTB(n9), .Q(
        key_round[7]) );
  DFFARX1_HVT \key_round_reg[8]  ( .D(n146), .CLK(clk), .RSTB(n14), .Q(
        key_round[8]) );
  DFFARX1_HVT \key_round_reg[9]  ( .D(n145), .CLK(clk), .RSTB(n11), .Q(
        key_round[9]) );
  DFFARX1_HVT \key_round_reg[10]  ( .D(n144), .CLK(clk), .RSTB(n13), .Q(
        key_round[10]) );
  DFFARX1_HVT \key_round_reg[11]  ( .D(n143), .CLK(clk), .RSTB(n10), .Q(
        key_round[11]) );
  DFFARX1_HVT \key_round_reg[12]  ( .D(n142), .CLK(clk), .RSTB(n9), .Q(
        key_round[12]) );
  DFFARX1_HVT \key_round_reg[13]  ( .D(n141), .CLK(clk), .RSTB(n7), .Q(
        key_round[13]) );
  DFFARX1_HVT \key_round_reg[14]  ( .D(n140), .CLK(clk), .RSTB(n6), .Q(
        key_round[14]) );
  DFFARX1_HVT \key_round_reg[15]  ( .D(n139), .CLK(clk), .RSTB(n5), .Q(
        key_round[15]) );
  DFFARX1_HVT \key_round_reg[16]  ( .D(n138), .CLK(clk), .RSTB(n11), .Q(
        key_round[16]) );
  DFFARX1_HVT \key_round_reg[17]  ( .D(n137), .CLK(clk), .RSTB(n14), .Q(
        key_round[17]) );
  DFFARX1_HVT \key_round_reg[18]  ( .D(n136), .CLK(clk), .RSTB(n13), .Q(
        key_round[18]) );
  DFFARX1_HVT \key_round_reg[19]  ( .D(n135), .CLK(clk), .RSTB(n8), .Q(
        key_round[19]) );
  DFFARX1_HVT \key_round_reg[20]  ( .D(n134), .CLK(clk), .RSTB(n7), .Q(
        key_round[20]) );
  DFFARX1_HVT \key_round_reg[21]  ( .D(n133), .CLK(clk), .RSTB(n9), .Q(
        key_round[21]) );
  DFFARX1_HVT \key_round_reg[22]  ( .D(n132), .CLK(clk), .RSTB(n6), .Q(
        key_round[22]) );
  DFFARX1_HVT \key_round_reg[23]  ( .D(n131), .CLK(clk), .RSTB(n5), .Q(
        key_round[23]) );
  DFFARX1_HVT \key_round_reg[24]  ( .D(n130), .CLK(clk), .RSTB(n8), .Q(
        key_round[24]) );
  DFFARX1_HVT \key_round_reg[25]  ( .D(n129), .CLK(clk), .RSTB(n6), .Q(
        key_round[25]) );
  DFFARX1_HVT \key_round_reg[26]  ( .D(n128), .CLK(clk), .RSTB(n13), .Q(
        key_round[26]) );
  DFFARX1_HVT \key_round_reg[27]  ( .D(n127), .CLK(clk), .RSTB(n7), .Q(
        key_round[27]) );
  DFFARX1_HVT \key_round_reg[28]  ( .D(n126), .CLK(clk), .RSTB(n14), .Q(
        key_round[28]) );
  DFFARX1_HVT \key_round_reg[29]  ( .D(n125), .CLK(clk), .RSTB(n10), .Q(
        key_round[29]) );
  DFFARX1_HVT \key_round_reg[30]  ( .D(n124), .CLK(clk), .RSTB(n9), .Q(
        key_round[30]) );
  DFFARX1_HVT \key_round_reg[31]  ( .D(n123), .CLK(clk), .RSTB(n25), .Q(
        key_round[31]) );
  DFFARX1_HVT \key_round_reg[32]  ( .D(n122), .CLK(clk), .RSTB(n11), .Q(
        key_round[32]) );
  DFFARX1_HVT \key_round_reg[33]  ( .D(n121), .CLK(clk), .RSTB(n10), .Q(
        key_round[33]) );
  DFFARX1_HVT \key_round_reg[34]  ( .D(n120), .CLK(clk), .RSTB(n13), .Q(
        key_round[34]) );
  DFFARX1_HVT \key_round_reg[35]  ( .D(n119), .CLK(clk), .RSTB(n8), .Q(
        key_round[35]) );
  DFFARX1_HVT \key_round_reg[36]  ( .D(n118), .CLK(clk), .RSTB(n5), .Q(
        key_round[36]) );
  DFFARX1_HVT \key_round_reg[37]  ( .D(n117), .CLK(clk), .RSTB(n7), .Q(
        key_round[37]) );
  DFFARX1_HVT \key_round_reg[38]  ( .D(n116), .CLK(clk), .RSTB(n25), .Q(
        key_round[38]) );
  DFFARX1_HVT \key_round_reg[39]  ( .D(n115), .CLK(clk), .RSTB(n9), .Q(
        key_round[39]) );
  DFFARX1_HVT \key_round_reg[40]  ( .D(n114), .CLK(clk), .RSTB(n6), .Q(
        key_round[40]) );
  DFFARX1_HVT \key_round_reg[41]  ( .D(n113), .CLK(clk), .RSTB(n11), .Q(
        key_round[41]) );
  DFFARX1_HVT \key_round_reg[42]  ( .D(n112), .CLK(clk), .RSTB(n13), .Q(
        key_round[42]) );
  DFFARX1_HVT \key_round_reg[43]  ( .D(n111), .CLK(clk), .RSTB(n10), .Q(
        key_round[43]) );
  DFFARX1_HVT \key_round_reg[44]  ( .D(n110), .CLK(clk), .RSTB(n25), .Q(
        key_round[44]) );
  DFFARX1_HVT \key_round_reg[45]  ( .D(n109), .CLK(clk), .RSTB(n7), .Q(
        key_round[45]) );
  DFFARX1_HVT \key_round_reg[46]  ( .D(n108), .CLK(clk), .RSTB(n6), .Q(
        key_round[46]) );
  DFFARX1_HVT \key_round_reg[47]  ( .D(n107), .CLK(clk), .RSTB(n5), .Q(
        key_round[47]) );
  DFFARX1_HVT \key_round_reg[48]  ( .D(n106), .CLK(clk), .RSTB(n11), .Q(
        key_round[48]) );
  DFFARX1_HVT \key_round_reg[49]  ( .D(n105), .CLK(clk), .RSTB(n14), .Q(
        key_round[49]) );
  DFFARX1_HVT \key_round_reg[50]  ( .D(n104), .CLK(clk), .RSTB(n13), .Q(
        key_round[50]) );
  DFFARX1_HVT \key_round_reg[51]  ( .D(n103), .CLK(clk), .RSTB(n8), .Q(
        key_round[51]) );
  DFFARX1_HVT \key_round_reg[52]  ( .D(n102), .CLK(clk), .RSTB(n25), .Q(
        key_round[52]) );
  DFFARX1_HVT \key_round_reg[53]  ( .D(n101), .CLK(clk), .RSTB(n10), .Q(
        key_round[53]) );
  DFFARX1_HVT \key_round_reg[54]  ( .D(n100), .CLK(clk), .RSTB(n6), .Q(
        key_round[54]) );
  DFFARX1_HVT \key_round_reg[55]  ( .D(n99), .CLK(clk), .RSTB(n5), .Q(
        key_round[55]) );
  DFFARX1_HVT \key_round_reg[56]  ( .D(n98), .CLK(clk), .RSTB(n8), .Q(
        key_round[56]) );
  DFFARX1_HVT \key_round_reg[57]  ( .D(n97), .CLK(clk), .RSTB(n6), .Q(
        key_round[57]) );
  DFFARX1_HVT \key_round_reg[58]  ( .D(n96), .CLK(clk), .RSTB(n13), .Q(
        key_round[58]) );
  DFFARX1_HVT \key_round_reg[59]  ( .D(n95), .CLK(clk), .RSTB(n7), .Q(
        key_round[59]) );
  DFFARX1_HVT \key_round_reg[60]  ( .D(n94), .CLK(clk), .RSTB(n14), .Q(
        key_round[60]) );
  DFFARX1_HVT \key_round_reg[61]  ( .D(n93), .CLK(clk), .RSTB(n10), .Q(
        key_round[61]) );
  DFFARX1_HVT \key_round_reg[62]  ( .D(n92), .CLK(clk), .RSTB(n9), .Q(
        key_round[62]) );
  DFFARX1_HVT \key_round_reg[63]  ( .D(n91), .CLK(clk), .RSTB(n5), .Q(
        key_round[63]) );
  DFFARX1_HVT \key_round_reg[64]  ( .D(n90), .CLK(clk), .RSTB(n11), .Q(
        key_round[64]) );
  DFFARX1_HVT \key_round_reg[65]  ( .D(n89), .CLK(clk), .RSTB(n10), .Q(
        key_round[65]) );
  DFFARX1_HVT \key_round_reg[66]  ( .D(n88), .CLK(clk), .RSTB(n14), .Q(
        key_round[66]) );
  DFFARX1_HVT \key_round_reg[67]  ( .D(n87), .CLK(clk), .RSTB(n8), .Q(
        key_round[67]) );
  DFFARX1_HVT \key_round_reg[68]  ( .D(n86), .CLK(clk), .RSTB(n6), .Q(
        key_round[68]) );
  DFFARX1_HVT \key_round_reg[69]  ( .D(n85), .CLK(clk), .RSTB(n7), .Q(
        key_round[69]) );
  DFFARX1_HVT \key_round_reg[70]  ( .D(n84), .CLK(clk), .RSTB(n25), .Q(
        key_round[70]) );
  DFFARX1_HVT \key_round_reg[71]  ( .D(n83), .CLK(clk), .RSTB(n9), .Q(
        key_round[71]) );
  DFFARX1_HVT \key_round_reg[72]  ( .D(n82), .CLK(clk), .RSTB(n25), .Q(
        key_round[72]) );
  DFFARX1_HVT \key_round_reg[73]  ( .D(n81), .CLK(clk), .RSTB(n11), .Q(
        key_round[73]) );
  DFFARX1_HVT \key_round_reg[74]  ( .D(n80), .CLK(clk), .RSTB(n13), .Q(
        key_round[74]) );
  DFFARX1_HVT \key_round_reg[75]  ( .D(n79), .CLK(clk), .RSTB(n10), .Q(
        key_round[75]) );
  DFFARX1_HVT \key_round_reg[76]  ( .D(n78), .CLK(clk), .RSTB(n9), .Q(
        key_round[76]) );
  DFFARX1_HVT \key_round_reg[77]  ( .D(n77), .CLK(clk), .RSTB(n7), .Q(
        key_round[77]) );
  DFFARX1_HVT \key_round_reg[78]  ( .D(n76), .CLK(clk), .RSTB(n6), .Q(
        key_round[78]) );
  DFFARX1_HVT \key_round_reg[79]  ( .D(n75), .CLK(clk), .RSTB(n5), .Q(
        key_round[79]) );
  DFFARX1_HVT \key_round_reg[80]  ( .D(n74), .CLK(clk), .RSTB(n11), .Q(
        key_round[80]) );
  DFFARX1_HVT \key_round_reg[81]  ( .D(n73), .CLK(clk), .RSTB(n14), .Q(
        key_round[81]) );
  DFFARX1_HVT \key_round_reg[82]  ( .D(n72), .CLK(clk), .RSTB(n13), .Q(
        key_round[82]) );
  DFFARX1_HVT \key_round_reg[83]  ( .D(n71), .CLK(clk), .RSTB(n8), .Q(
        key_round[83]) );
  DFFARX1_HVT \key_round_reg[84]  ( .D(n70), .CLK(clk), .RSTB(n7), .Q(
        key_round[84]) );
  DFFARX1_HVT \key_round_reg[85]  ( .D(n69), .CLK(clk), .RSTB(n10), .Q(
        key_round[85]) );
  DFFARX1_HVT \key_round_reg[86]  ( .D(n68), .CLK(clk), .RSTB(n6), .Q(
        key_round[86]) );
  DFFARX1_HVT \key_round_reg[87]  ( .D(n67), .CLK(clk), .RSTB(n5), .Q(
        key_round[87]) );
  DFFARX1_HVT \key_round_reg[88]  ( .D(n66), .CLK(clk), .RSTB(n8), .Q(
        key_round[88]) );
  DFFARX1_HVT \key_round_reg[89]  ( .D(n65), .CLK(clk), .RSTB(n6), .Q(
        key_round[89]) );
  DFFARX1_HVT \key_round_reg[90]  ( .D(n64), .CLK(clk), .RSTB(n13), .Q(
        key_round[90]) );
  DFFARX1_HVT \key_round_reg[91]  ( .D(n63), .CLK(clk), .RSTB(n7), .Q(
        key_round[91]) );
  DFFARX1_HVT \key_round_reg[92]  ( .D(n62), .CLK(clk), .RSTB(n14), .Q(
        key_round[92]) );
  DFFARX1_HVT \key_round_reg[93]  ( .D(n61), .CLK(clk), .RSTB(n11), .Q(
        key_round[93]) );
  DFFARX1_HVT \key_round_reg[94]  ( .D(n60), .CLK(clk), .RSTB(n9), .Q(
        key_round[94]) );
  DFFARX1_HVT \key_round_reg[95]  ( .D(n59), .CLK(clk), .RSTB(n5), .Q(
        key_round[95]) );
  DFFARX1_HVT \key_round_reg[96]  ( .D(n58), .CLK(clk), .RSTB(n11), .Q(
        key_round[96]) );
  DFFARX1_HVT \key_round_reg[97]  ( .D(n57), .CLK(clk), .RSTB(n10), .Q(
        key_round[97]) );
  DFFARX1_HVT \key_round_reg[98]  ( .D(n56), .CLK(clk), .RSTB(n14), .Q(
        key_round[98]) );
  DFFARX1_HVT \key_round_reg[99]  ( .D(n55), .CLK(clk), .RSTB(n8), .Q(
        key_round[99]) );
  DFFARX1_HVT \key_round_reg[100]  ( .D(n54), .CLK(clk), .RSTB(n6), .Q(
        key_round[100]) );
  DFFARX1_HVT \key_round_reg[101]  ( .D(n53), .CLK(clk), .RSTB(n7), .Q(
        key_round[101]) );
  DFFARX1_HVT \key_round_reg[102]  ( .D(n52), .CLK(clk), .RSTB(n25), .Q(
        key_round[102]) );
  DFFARX1_HVT \key_round_reg[103]  ( .D(n51), .CLK(clk), .RSTB(n9), .Q(
        key_round[103]) );
  DFFARX1_HVT \key_round_reg[104]  ( .D(n50), .CLK(clk), .RSTB(n9), .Q(
        key_round[104]) );
  DFFARX1_HVT \key_round_reg[105]  ( .D(n49), .CLK(clk), .RSTB(n11), .Q(
        key_round[105]) );
  DFFARX1_HVT \key_round_reg[106]  ( .D(n48), .CLK(clk), .RSTB(n13), .Q(
        key_round[106]) );
  DFFARX1_HVT \key_round_reg[107]  ( .D(n47), .CLK(clk), .RSTB(n10), .Q(
        key_round[107]) );
  DFFARX1_HVT \key_round_reg[108]  ( .D(n46), .CLK(clk), .RSTB(n9), .Q(
        key_round[108]) );
  DFFARX1_HVT \key_round_reg[109]  ( .D(n45), .CLK(clk), .RSTB(n8), .Q(
        key_round[109]) );
  DFFARX1_HVT \key_round_reg[110]  ( .D(n44), .CLK(clk), .RSTB(n6), .Q(
        key_round[110]) );
  DFFARX1_HVT \key_round_reg[111]  ( .D(n43), .CLK(clk), .RSTB(n5), .Q(
        key_round[111]) );
  DFFARX1_HVT \key_round_reg[112]  ( .D(n42), .CLK(clk), .RSTB(n25), .Q(
        key_round[112]) );
  DFFARX1_HVT \key_round_reg[113]  ( .D(n41), .CLK(clk), .RSTB(n14), .Q(
        key_round[113]) );
  DFFARX1_HVT \key_round_reg[114]  ( .D(n40), .CLK(clk), .RSTB(n13), .Q(
        key_round[114]) );
  DFFARX1_HVT \key_round_reg[115]  ( .D(n39), .CLK(clk), .RSTB(n8), .Q(
        key_round[115]) );
  DFFARX1_HVT \key_round_reg[116]  ( .D(n38), .CLK(clk), .RSTB(n7), .Q(
        key_round[116]) );
  DFFARX1_HVT \key_round_reg[117]  ( .D(n37), .CLK(clk), .RSTB(n10), .Q(
        key_round[117]) );
  DFFARX1_HVT \key_round_reg[118]  ( .D(n36), .CLK(clk), .RSTB(n6), .Q(
        key_round[118]) );
  DFFARX1_HVT \key_round_reg[119]  ( .D(n35), .CLK(clk), .RSTB(n5), .Q(
        key_round[119]) );
  DFFARX1_HVT \key_round_reg[120]  ( .D(n34), .CLK(clk), .RSTB(n8), .Q(
        key_round[120]) );
  DFFARX1_HVT \key_round_reg[121]  ( .D(n33), .CLK(clk), .RSTB(n25), .Q(
        key_round[121]) );
  DFFARX1_HVT \key_round_reg[122]  ( .D(n32), .CLK(clk), .RSTB(n25), .Q(
        key_round[122]) );
  DFFARX1_HVT \key_round_reg[123]  ( .D(n31), .CLK(clk), .RSTB(n25), .Q(
        key_round[123]) );
  DFFARX1_HVT \key_round_reg[124]  ( .D(n30), .CLK(clk), .RSTB(n24), .Q(
        key_round[124]) );
  DFFARX1_HVT \key_round_reg[125]  ( .D(n29), .CLK(clk), .RSTB(n11), .Q(
        key_round[125]) );
  DFFARX1_HVT \key_round_reg[126]  ( .D(n28), .CLK(clk), .RSTB(n9), .Q(
        key_round[126]) );
  DFFARX1_HVT \key_round_reg[127]  ( .D(n27), .CLK(clk), .RSTB(n5), .Q(
        key_round[127]) );
  DFFARX1_HVT ready_reg ( .D(n26), .CLK(clk), .RSTB(n14), .Q(ready), .QN(n304)
         );
  add_round_keys_0 adk_0 ( .state(plaintext), .subkey(key), .out(adk_out0) );
  round r1 ( .in(adk_in), .round_num(round_number), .keyin(key_round), 
        .keyout(keyout), .out(cipher_text) );
  NBUFFX2_HVT U3 ( .A(n305), .Y(n25) );
  NBUFFX2_HVT U4 ( .A(n305), .Y(n6) );
  NBUFFX2_HVT U5 ( .A(n305), .Y(n9) );
  NBUFFX2_HVT U6 ( .A(n305), .Y(n7) );
  NBUFFX2_HVT U7 ( .A(n305), .Y(n5) );
  NBUFFX2_HVT U8 ( .A(n305), .Y(n8) );
  NBUFFX2_HVT U9 ( .A(n305), .Y(n13) );
  NBUFFX2_HVT U10 ( .A(n305), .Y(n10) );
  NBUFFX2_HVT U11 ( .A(n305), .Y(n16) );
  NBUFFX2_HVT U12 ( .A(n305), .Y(n22) );
  NBUFFX2_HVT U13 ( .A(n305), .Y(n23) );
  NBUFFX2_HVT U14 ( .A(n305), .Y(n18) );
  NBUFFX2_HVT U15 ( .A(n305), .Y(n17) );
  NBUFFX2_HVT U16 ( .A(n305), .Y(n21) );
  NBUFFX2_HVT U17 ( .A(n305), .Y(n19) );
  NBUFFX2_HVT U18 ( .A(n305), .Y(n20) );
  NBUFFX2_HVT U19 ( .A(n305), .Y(n24) );
  NBUFFX2_HVT U20 ( .A(n305), .Y(n11) );
  NBUFFX2_HVT U21 ( .A(n305), .Y(n15) );
  NBUFFX2_HVT U22 ( .A(n305), .Y(n14) );
  INVX0_HVT U23 ( .A(reset), .Y(n305) );
  AO222X1_HVT U24 ( .A1(n288), .A2(key_round[55]), .A3(keyout[55]), .A4(n289), 
        .A5(key[55]), .A6(n290), .Y(n99) );
  AO222X1_HVT U25 ( .A1(n288), .A2(key_round[56]), .A3(keyout[56]), .A4(n289), 
        .A5(key[56]), .A6(n290), .Y(n98) );
  AO222X1_HVT U26 ( .A1(n288), .A2(key_round[57]), .A3(keyout[57]), .A4(n289), 
        .A5(key[57]), .A6(n290), .Y(n97) );
  AO222X1_HVT U27 ( .A1(n288), .A2(key_round[58]), .A3(keyout[58]), .A4(n289), 
        .A5(key[58]), .A6(n290), .Y(n96) );
  AO222X1_HVT U28 ( .A1(n288), .A2(key_round[59]), .A3(keyout[59]), .A4(n289), 
        .A5(key[59]), .A6(n290), .Y(n95) );
  AO222X1_HVT U29 ( .A1(n288), .A2(key_round[60]), .A3(keyout[60]), .A4(n289), 
        .A5(key[60]), .A6(n290), .Y(n94) );
  AO222X1_HVT U30 ( .A1(n288), .A2(key_round[61]), .A3(keyout[61]), .A4(n289), 
        .A5(key[61]), .A6(n290), .Y(n93) );
  AO222X1_HVT U31 ( .A1(n288), .A2(key_round[62]), .A3(keyout[62]), .A4(n289), 
        .A5(key[62]), .A6(n290), .Y(n92) );
  AO222X1_HVT U32 ( .A1(n288), .A2(key_round[63]), .A3(keyout[63]), .A4(n289), 
        .A5(key[63]), .A6(n290), .Y(n91) );
  AO222X1_HVT U33 ( .A1(n288), .A2(key_round[64]), .A3(keyout[64]), .A4(n289), 
        .A5(key[64]), .A6(n290), .Y(n90) );
  AO222X1_HVT U34 ( .A1(n288), .A2(key_round[65]), .A3(keyout[65]), .A4(n289), 
        .A5(key[65]), .A6(n290), .Y(n89) );
  AO222X1_HVT U35 ( .A1(n288), .A2(key_round[66]), .A3(keyout[66]), .A4(n289), 
        .A5(key[66]), .A6(n290), .Y(n88) );
  AO222X1_HVT U36 ( .A1(n288), .A2(key_round[67]), .A3(keyout[67]), .A4(n289), 
        .A5(key[67]), .A6(n290), .Y(n87) );
  AO222X1_HVT U37 ( .A1(n288), .A2(key_round[68]), .A3(keyout[68]), .A4(n289), 
        .A5(key[68]), .A6(n290), .Y(n86) );
  AO222X1_HVT U38 ( .A1(n288), .A2(key_round[69]), .A3(keyout[69]), .A4(n289), 
        .A5(key[69]), .A6(n290), .Y(n85) );
  AO222X1_HVT U39 ( .A1(n288), .A2(key_round[70]), .A3(keyout[70]), .A4(n289), 
        .A5(key[70]), .A6(n290), .Y(n84) );
  AO222X1_HVT U40 ( .A1(n288), .A2(key_round[71]), .A3(keyout[71]), .A4(n289), 
        .A5(key[71]), .A6(n290), .Y(n83) );
  AO222X1_HVT U41 ( .A1(n288), .A2(key_round[72]), .A3(keyout[72]), .A4(n289), 
        .A5(key[72]), .A6(n290), .Y(n82) );
  AO222X1_HVT U42 ( .A1(n288), .A2(key_round[73]), .A3(keyout[73]), .A4(n289), 
        .A5(key[73]), .A6(n290), .Y(n81) );
  AO222X1_HVT U43 ( .A1(n288), .A2(key_round[74]), .A3(keyout[74]), .A4(n289), 
        .A5(key[74]), .A6(n290), .Y(n80) );
  AO222X1_HVT U44 ( .A1(n288), .A2(key_round[75]), .A3(keyout[75]), .A4(n289), 
        .A5(key[75]), .A6(n290), .Y(n79) );
  AO222X1_HVT U45 ( .A1(n288), .A2(key_round[76]), .A3(keyout[76]), .A4(n289), 
        .A5(key[76]), .A6(n290), .Y(n78) );
  AO222X1_HVT U46 ( .A1(n288), .A2(key_round[77]), .A3(keyout[77]), .A4(n289), 
        .A5(key[77]), .A6(n290), .Y(n77) );
  AO222X1_HVT U47 ( .A1(n288), .A2(key_round[78]), .A3(keyout[78]), .A4(n289), 
        .A5(key[78]), .A6(n290), .Y(n76) );
  AO222X1_HVT U48 ( .A1(n288), .A2(key_round[79]), .A3(keyout[79]), .A4(n289), 
        .A5(key[79]), .A6(n290), .Y(n75) );
  AO222X1_HVT U49 ( .A1(n288), .A2(key_round[80]), .A3(keyout[80]), .A4(n289), 
        .A5(key[80]), .A6(n290), .Y(n74) );
  AO222X1_HVT U50 ( .A1(n288), .A2(key_round[81]), .A3(keyout[81]), .A4(n289), 
        .A5(key[81]), .A6(n290), .Y(n73) );
  AO222X1_HVT U51 ( .A1(n288), .A2(key_round[82]), .A3(keyout[82]), .A4(n289), 
        .A5(key[82]), .A6(n290), .Y(n72) );
  AO222X1_HVT U52 ( .A1(n288), .A2(key_round[83]), .A3(keyout[83]), .A4(n289), 
        .A5(key[83]), .A6(n290), .Y(n71) );
  AO222X1_HVT U53 ( .A1(n288), .A2(key_round[84]), .A3(keyout[84]), .A4(n289), 
        .A5(key[84]), .A6(n290), .Y(n70) );
  AO222X1_HVT U54 ( .A1(n288), .A2(key_round[85]), .A3(keyout[85]), .A4(n289), 
        .A5(key[85]), .A6(n290), .Y(n69) );
  AO222X1_HVT U55 ( .A1(n288), .A2(key_round[86]), .A3(keyout[86]), .A4(n289), 
        .A5(key[86]), .A6(n290), .Y(n68) );
  AO222X1_HVT U56 ( .A1(n288), .A2(key_round[87]), .A3(keyout[87]), .A4(n289), 
        .A5(key[87]), .A6(n290), .Y(n67) );
  AO222X1_HVT U57 ( .A1(n288), .A2(key_round[88]), .A3(keyout[88]), .A4(n289), 
        .A5(key[88]), .A6(n290), .Y(n66) );
  AO222X1_HVT U58 ( .A1(n288), .A2(key_round[89]), .A3(keyout[89]), .A4(n289), 
        .A5(key[89]), .A6(n290), .Y(n65) );
  AO222X1_HVT U59 ( .A1(n288), .A2(key_round[90]), .A3(keyout[90]), .A4(n289), 
        .A5(key[90]), .A6(n290), .Y(n64) );
  AO222X1_HVT U60 ( .A1(n288), .A2(key_round[91]), .A3(keyout[91]), .A4(n289), 
        .A5(key[91]), .A6(n290), .Y(n63) );
  AO222X1_HVT U61 ( .A1(n288), .A2(key_round[92]), .A3(keyout[92]), .A4(n289), 
        .A5(key[92]), .A6(n290), .Y(n62) );
  AO222X1_HVT U62 ( .A1(n288), .A2(key_round[93]), .A3(keyout[93]), .A4(n289), 
        .A5(key[93]), .A6(n290), .Y(n61) );
  AO222X1_HVT U63 ( .A1(n288), .A2(key_round[94]), .A3(keyout[94]), .A4(n289), 
        .A5(key[94]), .A6(n290), .Y(n60) );
  AO222X1_HVT U64 ( .A1(n288), .A2(key_round[95]), .A3(keyout[95]), .A4(n289), 
        .A5(key[95]), .A6(n290), .Y(n59) );
  AO222X1_HVT U65 ( .A1(n288), .A2(key_round[96]), .A3(keyout[96]), .A4(n289), 
        .A5(key[96]), .A6(n290), .Y(n58) );
  AO222X1_HVT U66 ( .A1(n288), .A2(key_round[97]), .A3(keyout[97]), .A4(n289), 
        .A5(key[97]), .A6(n290), .Y(n57) );
  AO222X1_HVT U67 ( .A1(n288), .A2(key_round[98]), .A3(keyout[98]), .A4(n289), 
        .A5(key[98]), .A6(n290), .Y(n56) );
  AO222X1_HVT U68 ( .A1(n288), .A2(key_round[99]), .A3(keyout[99]), .A4(n289), 
        .A5(key[99]), .A6(n290), .Y(n55) );
  AO222X1_HVT U69 ( .A1(n288), .A2(key_round[100]), .A3(keyout[100]), .A4(n289), .A5(key[100]), .A6(n290), .Y(n54) );
  AO222X1_HVT U70 ( .A1(n288), .A2(key_round[101]), .A3(keyout[101]), .A4(n289), .A5(key[101]), .A6(n290), .Y(n53) );
  AO222X1_HVT U71 ( .A1(n288), .A2(key_round[102]), .A3(keyout[102]), .A4(n289), .A5(key[102]), .A6(n290), .Y(n52) );
  AO222X1_HVT U72 ( .A1(n288), .A2(key_round[103]), .A3(keyout[103]), .A4(n289), .A5(key[103]), .A6(n290), .Y(n51) );
  AO222X1_HVT U73 ( .A1(n288), .A2(key_round[104]), .A3(keyout[104]), .A4(n289), .A5(key[104]), .A6(n290), .Y(n50) );
  AO222X1_HVT U74 ( .A1(n288), .A2(key_round[105]), .A3(keyout[105]), .A4(n289), .A5(key[105]), .A6(n290), .Y(n49) );
  AO222X1_HVT U75 ( .A1(n288), .A2(key_round[106]), .A3(keyout[106]), .A4(n289), .A5(key[106]), .A6(n290), .Y(n48) );
  AO222X1_HVT U76 ( .A1(n288), .A2(key_round[107]), .A3(keyout[107]), .A4(n289), .A5(key[107]), .A6(n290), .Y(n47) );
  AO222X1_HVT U77 ( .A1(n288), .A2(key_round[108]), .A3(keyout[108]), .A4(n289), .A5(key[108]), .A6(n290), .Y(n46) );
  AO222X1_HVT U78 ( .A1(n288), .A2(key_round[109]), .A3(keyout[109]), .A4(n289), .A5(key[109]), .A6(n290), .Y(n45) );
  AO222X1_HVT U79 ( .A1(n288), .A2(key_round[110]), .A3(keyout[110]), .A4(n289), .A5(key[110]), .A6(n290), .Y(n44) );
  AO222X1_HVT U80 ( .A1(n288), .A2(key_round[111]), .A3(keyout[111]), .A4(n289), .A5(key[111]), .A6(n290), .Y(n43) );
  AO222X1_HVT U81 ( .A1(n288), .A2(key_round[112]), .A3(keyout[112]), .A4(n289), .A5(key[112]), .A6(n290), .Y(n42) );
  AO222X1_HVT U82 ( .A1(n288), .A2(key_round[113]), .A3(keyout[113]), .A4(n289), .A5(key[113]), .A6(n290), .Y(n41) );
  AO222X1_HVT U83 ( .A1(n288), .A2(key_round[114]), .A3(keyout[114]), .A4(n289), .A5(key[114]), .A6(n290), .Y(n40) );
  AO222X1_HVT U84 ( .A1(n288), .A2(key_round[115]), .A3(keyout[115]), .A4(n289), .A5(key[115]), .A6(n290), .Y(n39) );
  AO222X1_HVT U85 ( .A1(n288), .A2(key_round[116]), .A3(keyout[116]), .A4(n289), .A5(key[116]), .A6(n290), .Y(n38) );
  AO222X1_HVT U86 ( .A1(n288), .A2(key_round[117]), .A3(keyout[117]), .A4(n289), .A5(key[117]), .A6(n290), .Y(n37) );
  AO222X1_HVT U87 ( .A1(n288), .A2(key_round[118]), .A3(keyout[118]), .A4(n289), .A5(key[118]), .A6(n290), .Y(n36) );
  AO222X1_HVT U88 ( .A1(n288), .A2(key_round[119]), .A3(keyout[119]), .A4(n289), .A5(key[119]), .A6(n290), .Y(n35) );
  AO222X1_HVT U89 ( .A1(n288), .A2(key_round[120]), .A3(keyout[120]), .A4(n289), .A5(key[120]), .A6(n290), .Y(n34) );
  AO222X1_HVT U90 ( .A1(n288), .A2(key_round[121]), .A3(keyout[121]), .A4(n289), .A5(key[121]), .A6(n290), .Y(n33) );
  AO222X1_HVT U91 ( .A1(n288), .A2(key_round[122]), .A3(keyout[122]), .A4(n289), .A5(key[122]), .A6(n290), .Y(n32) );
  AO222X1_HVT U92 ( .A1(n288), .A2(key_round[123]), .A3(keyout[123]), .A4(n289), .A5(key[123]), .A6(n290), .Y(n31) );
  AO222X1_HVT U93 ( .A1(n288), .A2(key_round[124]), .A3(keyout[124]), .A4(n289), .A5(key[124]), .A6(n290), .Y(n30) );
  AO222X1_HVT U94 ( .A1(n288), .A2(key_round[125]), .A3(keyout[125]), .A4(n289), .A5(key[125]), .A6(n290), .Y(n29) );
  NAND2X0_HVT U95 ( .A1(n291), .A2(n292), .Y(n287) );
  AO21X1_HVT U96 ( .A1(start), .A2(n288), .A3(n12), .Y(n292) );
  AO22X1_HVT U97 ( .A1(round_number[3]), .A2(n293), .A3(round_number[2]), .A4(
        n294), .Y(n286) );
  MUX21X1_HVT U98 ( .A1(n295), .A2(n296), .S0(n3), .Y(n285) );
  AND2X1_HVT U99 ( .A1(n288), .A2(n297), .Y(n295) );
  MUX21X1_HVT U100 ( .A1(n298), .A2(n299), .S0(n4), .Y(n284) );
  AND2X1_HVT U101 ( .A1(round_number[0]), .A2(n296), .Y(n299) );
  MUX21X1_HVT U102 ( .A1(n293), .A2(n294), .S0(n1), .Y(n283) );
  AND3X1_HVT U103 ( .A1(round_number[1]), .A2(n296), .A3(round_number[0]), .Y(
        n294) );
  AO21X1_HVT U104 ( .A1(n296), .A2(n4), .A3(n298), .Y(n293) );
  MUX21X1_HVT U105 ( .A1(n3), .A2(n297), .S0(n288), .Y(n298) );
  NAND2X0_HVT U106 ( .A1(start), .A2(n2), .Y(n297) );
  AO222X1_HVT U107 ( .A1(n288), .A2(key_round[0]), .A3(keyout[0]), .A4(n289), 
        .A5(key[0]), .A6(n290), .Y(n282) );
  AO222X1_HVT U108 ( .A1(n288), .A2(adk_in[0]), .A3(cipher_text[0]), .A4(n289), 
        .A5(adk_out0[0]), .A6(n290), .Y(n281) );
  AO222X1_HVT U109 ( .A1(n288), .A2(adk_in[1]), .A3(cipher_text[1]), .A4(n289), 
        .A5(adk_out0[1]), .A6(n290), .Y(n280) );
  AO222X1_HVT U110 ( .A1(n288), .A2(key_round[126]), .A3(keyout[126]), .A4(
        n289), .A5(key[126]), .A6(n290), .Y(n28) );
  AO222X1_HVT U111 ( .A1(n288), .A2(adk_in[2]), .A3(cipher_text[2]), .A4(n289), 
        .A5(adk_out0[2]), .A6(n290), .Y(n279) );
  AO222X1_HVT U112 ( .A1(n288), .A2(adk_in[3]), .A3(cipher_text[3]), .A4(n289), 
        .A5(adk_out0[3]), .A6(n290), .Y(n278) );
  AO222X1_HVT U113 ( .A1(n288), .A2(adk_in[4]), .A3(cipher_text[4]), .A4(n289), 
        .A5(adk_out0[4]), .A6(n290), .Y(n277) );
  AO222X1_HVT U114 ( .A1(n288), .A2(adk_in[5]), .A3(cipher_text[5]), .A4(n289), 
        .A5(adk_out0[5]), .A6(n290), .Y(n276) );
  AO222X1_HVT U115 ( .A1(n288), .A2(adk_in[6]), .A3(cipher_text[6]), .A4(n289), 
        .A5(adk_out0[6]), .A6(n290), .Y(n275) );
  AO222X1_HVT U116 ( .A1(n288), .A2(adk_in[7]), .A3(cipher_text[7]), .A4(n289), 
        .A5(adk_out0[7]), .A6(n290), .Y(n274) );
  AO222X1_HVT U117 ( .A1(n288), .A2(adk_in[8]), .A3(cipher_text[8]), .A4(n289), 
        .A5(adk_out0[8]), .A6(n290), .Y(n273) );
  AO222X1_HVT U118 ( .A1(n288), .A2(adk_in[9]), .A3(cipher_text[9]), .A4(n289), 
        .A5(adk_out0[9]), .A6(n290), .Y(n272) );
  AO222X1_HVT U119 ( .A1(n288), .A2(adk_in[10]), .A3(cipher_text[10]), .A4(
        n289), .A5(adk_out0[10]), .A6(n290), .Y(n271) );
  AO222X1_HVT U120 ( .A1(n288), .A2(adk_in[11]), .A3(cipher_text[11]), .A4(
        n289), .A5(adk_out0[11]), .A6(n290), .Y(n270) );
  AO222X1_HVT U121 ( .A1(n288), .A2(key_round[127]), .A3(keyout[127]), .A4(
        n289), .A5(key[127]), .A6(n290), .Y(n27) );
  AO222X1_HVT U122 ( .A1(n288), .A2(adk_in[12]), .A3(cipher_text[12]), .A4(
        n289), .A5(adk_out0[12]), .A6(n290), .Y(n269) );
  AO222X1_HVT U123 ( .A1(n288), .A2(adk_in[13]), .A3(cipher_text[13]), .A4(
        n289), .A5(adk_out0[13]), .A6(n290), .Y(n268) );
  AO222X1_HVT U124 ( .A1(n288), .A2(adk_in[14]), .A3(cipher_text[14]), .A4(
        n289), .A5(adk_out0[14]), .A6(n290), .Y(n267) );
  AO222X1_HVT U125 ( .A1(n288), .A2(adk_in[15]), .A3(cipher_text[15]), .A4(
        n289), .A5(adk_out0[15]), .A6(n290), .Y(n266) );
  AO222X1_HVT U126 ( .A1(n288), .A2(adk_in[16]), .A3(cipher_text[16]), .A4(
        n289), .A5(adk_out0[16]), .A6(n290), .Y(n265) );
  AO222X1_HVT U127 ( .A1(n288), .A2(adk_in[17]), .A3(cipher_text[17]), .A4(
        n289), .A5(adk_out0[17]), .A6(n290), .Y(n264) );
  AO222X1_HVT U128 ( .A1(n288), .A2(adk_in[18]), .A3(cipher_text[18]), .A4(
        n289), .A5(adk_out0[18]), .A6(n290), .Y(n263) );
  AO222X1_HVT U129 ( .A1(n288), .A2(adk_in[19]), .A3(cipher_text[19]), .A4(
        n289), .A5(adk_out0[19]), .A6(n290), .Y(n262) );
  AO222X1_HVT U130 ( .A1(n288), .A2(adk_in[20]), .A3(cipher_text[20]), .A4(
        n289), .A5(adk_out0[20]), .A6(n290), .Y(n261) );
  AO222X1_HVT U131 ( .A1(n288), .A2(adk_in[21]), .A3(cipher_text[21]), .A4(
        n289), .A5(adk_out0[21]), .A6(n290), .Y(n260) );
  NAND2X0_HVT U132 ( .A1(n291), .A2(n300), .Y(n26) );
  AO21X1_HVT U133 ( .A1(n288), .A2(n2), .A3(n304), .Y(n300) );
  NAND4X0_HVT U134 ( .A1(n3), .A2(n1), .A3(round_number[3]), .A4(n301), .Y(
        n291) );
  AND2X1_HVT U135 ( .A1(round_number[1]), .A2(n12), .Y(n301) );
  AO222X1_HVT U136 ( .A1(n288), .A2(adk_in[22]), .A3(cipher_text[22]), .A4(
        n289), .A5(adk_out0[22]), .A6(n290), .Y(n259) );
  AO222X1_HVT U137 ( .A1(n288), .A2(adk_in[23]), .A3(cipher_text[23]), .A4(
        n289), .A5(adk_out0[23]), .A6(n290), .Y(n258) );
  AO222X1_HVT U138 ( .A1(n288), .A2(adk_in[24]), .A3(cipher_text[24]), .A4(
        n289), .A5(adk_out0[24]), .A6(n290), .Y(n257) );
  AO222X1_HVT U139 ( .A1(n288), .A2(adk_in[25]), .A3(cipher_text[25]), .A4(
        n289), .A5(adk_out0[25]), .A6(n290), .Y(n256) );
  AO222X1_HVT U140 ( .A1(n288), .A2(adk_in[26]), .A3(cipher_text[26]), .A4(
        n289), .A5(adk_out0[26]), .A6(n290), .Y(n255) );
  AO222X1_HVT U141 ( .A1(n288), .A2(adk_in[27]), .A3(cipher_text[27]), .A4(
        n289), .A5(adk_out0[27]), .A6(n290), .Y(n254) );
  AO222X1_HVT U142 ( .A1(n288), .A2(adk_in[28]), .A3(cipher_text[28]), .A4(
        n289), .A5(adk_out0[28]), .A6(n290), .Y(n253) );
  AO222X1_HVT U143 ( .A1(n288), .A2(adk_in[29]), .A3(cipher_text[29]), .A4(
        n289), .A5(adk_out0[29]), .A6(n290), .Y(n252) );
  AO222X1_HVT U144 ( .A1(n288), .A2(adk_in[30]), .A3(cipher_text[30]), .A4(
        n289), .A5(adk_out0[30]), .A6(n290), .Y(n251) );
  AO222X1_HVT U145 ( .A1(n288), .A2(adk_in[31]), .A3(cipher_text[31]), .A4(
        n289), .A5(adk_out0[31]), .A6(n290), .Y(n250) );
  AO222X1_HVT U146 ( .A1(n288), .A2(adk_in[32]), .A3(cipher_text[32]), .A4(
        n289), .A5(adk_out0[32]), .A6(n290), .Y(n249) );
  AO222X1_HVT U147 ( .A1(n288), .A2(adk_in[33]), .A3(cipher_text[33]), .A4(
        n289), .A5(adk_out0[33]), .A6(n290), .Y(n248) );
  AO222X1_HVT U148 ( .A1(n288), .A2(adk_in[34]), .A3(cipher_text[34]), .A4(
        n289), .A5(adk_out0[34]), .A6(n290), .Y(n247) );
  AO222X1_HVT U149 ( .A1(n288), .A2(adk_in[35]), .A3(cipher_text[35]), .A4(
        n289), .A5(adk_out0[35]), .A6(n290), .Y(n246) );
  AO222X1_HVT U150 ( .A1(n288), .A2(adk_in[36]), .A3(cipher_text[36]), .A4(
        n289), .A5(adk_out0[36]), .A6(n290), .Y(n245) );
  AO222X1_HVT U151 ( .A1(n288), .A2(adk_in[37]), .A3(cipher_text[37]), .A4(
        n289), .A5(adk_out0[37]), .A6(n290), .Y(n244) );
  AO222X1_HVT U152 ( .A1(n288), .A2(adk_in[38]), .A3(cipher_text[38]), .A4(
        n289), .A5(adk_out0[38]), .A6(n290), .Y(n243) );
  AO222X1_HVT U153 ( .A1(n288), .A2(adk_in[39]), .A3(cipher_text[39]), .A4(
        n289), .A5(adk_out0[39]), .A6(n290), .Y(n242) );
  AO222X1_HVT U154 ( .A1(n288), .A2(adk_in[40]), .A3(cipher_text[40]), .A4(
        n289), .A5(adk_out0[40]), .A6(n290), .Y(n241) );
  AO222X1_HVT U155 ( .A1(n288), .A2(adk_in[41]), .A3(cipher_text[41]), .A4(
        n289), .A5(adk_out0[41]), .A6(n290), .Y(n240) );
  AO222X1_HVT U156 ( .A1(n288), .A2(adk_in[42]), .A3(cipher_text[42]), .A4(
        n289), .A5(adk_out0[42]), .A6(n290), .Y(n239) );
  AO222X1_HVT U157 ( .A1(n288), .A2(adk_in[43]), .A3(cipher_text[43]), .A4(
        n289), .A5(adk_out0[43]), .A6(n290), .Y(n238) );
  AO222X1_HVT U158 ( .A1(n288), .A2(adk_in[44]), .A3(cipher_text[44]), .A4(
        n289), .A5(adk_out0[44]), .A6(n290), .Y(n237) );
  AO222X1_HVT U159 ( .A1(n288), .A2(adk_in[45]), .A3(cipher_text[45]), .A4(
        n289), .A5(adk_out0[45]), .A6(n290), .Y(n236) );
  AO222X1_HVT U160 ( .A1(n288), .A2(adk_in[46]), .A3(cipher_text[46]), .A4(
        n289), .A5(adk_out0[46]), .A6(n290), .Y(n235) );
  AO222X1_HVT U161 ( .A1(n288), .A2(adk_in[47]), .A3(cipher_text[47]), .A4(
        n289), .A5(adk_out0[47]), .A6(n290), .Y(n234) );
  AO222X1_HVT U162 ( .A1(n288), .A2(adk_in[48]), .A3(cipher_text[48]), .A4(
        n289), .A5(adk_out0[48]), .A6(n290), .Y(n233) );
  AO222X1_HVT U163 ( .A1(n288), .A2(adk_in[49]), .A3(cipher_text[49]), .A4(
        n289), .A5(adk_out0[49]), .A6(n290), .Y(n232) );
  AO222X1_HVT U164 ( .A1(n288), .A2(adk_in[50]), .A3(cipher_text[50]), .A4(
        n289), .A5(adk_out0[50]), .A6(n290), .Y(n231) );
  AO222X1_HVT U165 ( .A1(n288), .A2(adk_in[51]), .A3(cipher_text[51]), .A4(
        n289), .A5(adk_out0[51]), .A6(n290), .Y(n230) );
  AO222X1_HVT U166 ( .A1(n288), .A2(adk_in[52]), .A3(cipher_text[52]), .A4(
        n289), .A5(adk_out0[52]), .A6(n290), .Y(n229) );
  AO222X1_HVT U167 ( .A1(n288), .A2(adk_in[53]), .A3(cipher_text[53]), .A4(
        n289), .A5(adk_out0[53]), .A6(n290), .Y(n228) );
  AO222X1_HVT U168 ( .A1(n288), .A2(adk_in[54]), .A3(cipher_text[54]), .A4(
        n289), .A5(adk_out0[54]), .A6(n290), .Y(n227) );
  AO222X1_HVT U169 ( .A1(n288), .A2(adk_in[55]), .A3(cipher_text[55]), .A4(
        n289), .A5(adk_out0[55]), .A6(n290), .Y(n226) );
  AO222X1_HVT U170 ( .A1(n288), .A2(adk_in[56]), .A3(cipher_text[56]), .A4(
        n289), .A5(adk_out0[56]), .A6(n290), .Y(n225) );
  AO222X1_HVT U171 ( .A1(n288), .A2(adk_in[57]), .A3(cipher_text[57]), .A4(
        n289), .A5(adk_out0[57]), .A6(n290), .Y(n224) );
  AO222X1_HVT U172 ( .A1(n288), .A2(adk_in[58]), .A3(cipher_text[58]), .A4(
        n289), .A5(adk_out0[58]), .A6(n290), .Y(n223) );
  AO222X1_HVT U173 ( .A1(n288), .A2(adk_in[59]), .A3(cipher_text[59]), .A4(
        n289), .A5(adk_out0[59]), .A6(n290), .Y(n222) );
  AO222X1_HVT U174 ( .A1(n288), .A2(adk_in[60]), .A3(cipher_text[60]), .A4(
        n289), .A5(adk_out0[60]), .A6(n290), .Y(n221) );
  AO222X1_HVT U175 ( .A1(n288), .A2(adk_in[61]), .A3(cipher_text[61]), .A4(
        n289), .A5(adk_out0[61]), .A6(n290), .Y(n220) );
  AO222X1_HVT U176 ( .A1(n288), .A2(adk_in[62]), .A3(cipher_text[62]), .A4(
        n289), .A5(adk_out0[62]), .A6(n290), .Y(n219) );
  AO222X1_HVT U177 ( .A1(n288), .A2(adk_in[63]), .A3(cipher_text[63]), .A4(
        n289), .A5(adk_out0[63]), .A6(n290), .Y(n218) );
  AO222X1_HVT U178 ( .A1(n288), .A2(adk_in[64]), .A3(cipher_text[64]), .A4(
        n289), .A5(adk_out0[64]), .A6(n290), .Y(n217) );
  AO222X1_HVT U179 ( .A1(n288), .A2(adk_in[65]), .A3(cipher_text[65]), .A4(
        n289), .A5(adk_out0[65]), .A6(n290), .Y(n216) );
  AO222X1_HVT U180 ( .A1(n288), .A2(adk_in[66]), .A3(cipher_text[66]), .A4(
        n289), .A5(adk_out0[66]), .A6(n290), .Y(n215) );
  AO222X1_HVT U181 ( .A1(n288), .A2(adk_in[67]), .A3(cipher_text[67]), .A4(
        n289), .A5(adk_out0[67]), .A6(n290), .Y(n214) );
  AO222X1_HVT U182 ( .A1(n288), .A2(adk_in[68]), .A3(cipher_text[68]), .A4(
        n289), .A5(adk_out0[68]), .A6(n290), .Y(n213) );
  AO222X1_HVT U183 ( .A1(n288), .A2(adk_in[69]), .A3(cipher_text[69]), .A4(
        n289), .A5(adk_out0[69]), .A6(n290), .Y(n212) );
  AO222X1_HVT U184 ( .A1(n288), .A2(adk_in[70]), .A3(cipher_text[70]), .A4(
        n289), .A5(adk_out0[70]), .A6(n290), .Y(n211) );
  AO222X1_HVT U185 ( .A1(n288), .A2(adk_in[71]), .A3(cipher_text[71]), .A4(
        n289), .A5(adk_out0[71]), .A6(n290), .Y(n210) );
  AO222X1_HVT U186 ( .A1(n288), .A2(adk_in[72]), .A3(cipher_text[72]), .A4(
        n289), .A5(adk_out0[72]), .A6(n290), .Y(n209) );
  AO222X1_HVT U187 ( .A1(n288), .A2(adk_in[73]), .A3(cipher_text[73]), .A4(
        n289), .A5(adk_out0[73]), .A6(n290), .Y(n208) );
  AO222X1_HVT U188 ( .A1(n288), .A2(adk_in[74]), .A3(cipher_text[74]), .A4(
        n289), .A5(adk_out0[74]), .A6(n290), .Y(n207) );
  AO222X1_HVT U189 ( .A1(n288), .A2(adk_in[75]), .A3(cipher_text[75]), .A4(
        n289), .A5(adk_out0[75]), .A6(n290), .Y(n206) );
  AO222X1_HVT U190 ( .A1(n288), .A2(adk_in[76]), .A3(cipher_text[76]), .A4(
        n289), .A5(adk_out0[76]), .A6(n290), .Y(n205) );
  AO222X1_HVT U191 ( .A1(n288), .A2(adk_in[77]), .A3(cipher_text[77]), .A4(
        n289), .A5(adk_out0[77]), .A6(n290), .Y(n204) );
  AO222X1_HVT U192 ( .A1(n288), .A2(adk_in[78]), .A3(cipher_text[78]), .A4(
        n289), .A5(adk_out0[78]), .A6(n290), .Y(n203) );
  AO222X1_HVT U193 ( .A1(n288), .A2(adk_in[79]), .A3(cipher_text[79]), .A4(
        n289), .A5(adk_out0[79]), .A6(n290), .Y(n202) );
  AO222X1_HVT U194 ( .A1(n288), .A2(adk_in[80]), .A3(cipher_text[80]), .A4(
        n289), .A5(adk_out0[80]), .A6(n290), .Y(n201) );
  AO222X1_HVT U195 ( .A1(n288), .A2(adk_in[81]), .A3(cipher_text[81]), .A4(
        n289), .A5(adk_out0[81]), .A6(n290), .Y(n200) );
  AO222X1_HVT U196 ( .A1(n288), .A2(adk_in[82]), .A3(cipher_text[82]), .A4(
        n289), .A5(adk_out0[82]), .A6(n290), .Y(n199) );
  AO222X1_HVT U197 ( .A1(n288), .A2(adk_in[83]), .A3(cipher_text[83]), .A4(
        n289), .A5(adk_out0[83]), .A6(n290), .Y(n198) );
  AO222X1_HVT U198 ( .A1(n288), .A2(adk_in[84]), .A3(cipher_text[84]), .A4(
        n289), .A5(adk_out0[84]), .A6(n290), .Y(n197) );
  AO222X1_HVT U199 ( .A1(n288), .A2(adk_in[85]), .A3(cipher_text[85]), .A4(
        n289), .A5(adk_out0[85]), .A6(n290), .Y(n196) );
  AO222X1_HVT U200 ( .A1(n288), .A2(adk_in[86]), .A3(cipher_text[86]), .A4(
        n289), .A5(adk_out0[86]), .A6(n290), .Y(n195) );
  AO222X1_HVT U201 ( .A1(n288), .A2(adk_in[87]), .A3(cipher_text[87]), .A4(
        n289), .A5(adk_out0[87]), .A6(n290), .Y(n194) );
  AO222X1_HVT U202 ( .A1(n288), .A2(adk_in[88]), .A3(cipher_text[88]), .A4(
        n289), .A5(adk_out0[88]), .A6(n290), .Y(n193) );
  AO222X1_HVT U203 ( .A1(n288), .A2(adk_in[89]), .A3(cipher_text[89]), .A4(
        n289), .A5(adk_out0[89]), .A6(n290), .Y(n192) );
  AO222X1_HVT U204 ( .A1(n288), .A2(adk_in[90]), .A3(cipher_text[90]), .A4(
        n289), .A5(adk_out0[90]), .A6(n290), .Y(n191) );
  AO222X1_HVT U205 ( .A1(n288), .A2(adk_in[91]), .A3(cipher_text[91]), .A4(
        n289), .A5(adk_out0[91]), .A6(n290), .Y(n190) );
  AO222X1_HVT U206 ( .A1(n288), .A2(adk_in[92]), .A3(cipher_text[92]), .A4(
        n289), .A5(adk_out0[92]), .A6(n290), .Y(n189) );
  AO222X1_HVT U207 ( .A1(n288), .A2(adk_in[93]), .A3(cipher_text[93]), .A4(
        n289), .A5(adk_out0[93]), .A6(n290), .Y(n188) );
  AO222X1_HVT U208 ( .A1(n288), .A2(adk_in[94]), .A3(cipher_text[94]), .A4(
        n289), .A5(adk_out0[94]), .A6(n290), .Y(n187) );
  AO222X1_HVT U209 ( .A1(n288), .A2(adk_in[95]), .A3(cipher_text[95]), .A4(
        n289), .A5(adk_out0[95]), .A6(n290), .Y(n186) );
  AO222X1_HVT U210 ( .A1(n288), .A2(adk_in[96]), .A3(cipher_text[96]), .A4(
        n289), .A5(adk_out0[96]), .A6(n290), .Y(n185) );
  AO222X1_HVT U211 ( .A1(n288), .A2(adk_in[97]), .A3(cipher_text[97]), .A4(
        n289), .A5(adk_out0[97]), .A6(n290), .Y(n184) );
  AO222X1_HVT U212 ( .A1(n288), .A2(adk_in[98]), .A3(cipher_text[98]), .A4(
        n289), .A5(adk_out0[98]), .A6(n290), .Y(n183) );
  AO222X1_HVT U213 ( .A1(n288), .A2(adk_in[99]), .A3(cipher_text[99]), .A4(
        n289), .A5(adk_out0[99]), .A6(n290), .Y(n182) );
  AO222X1_HVT U214 ( .A1(n288), .A2(adk_in[100]), .A3(cipher_text[100]), .A4(
        n289), .A5(adk_out0[100]), .A6(n290), .Y(n181) );
  AO222X1_HVT U215 ( .A1(n288), .A2(adk_in[101]), .A3(cipher_text[101]), .A4(
        n289), .A5(adk_out0[101]), .A6(n290), .Y(n180) );
  AO222X1_HVT U216 ( .A1(n288), .A2(adk_in[102]), .A3(cipher_text[102]), .A4(
        n289), .A5(adk_out0[102]), .A6(n290), .Y(n179) );
  AO222X1_HVT U217 ( .A1(n288), .A2(adk_in[103]), .A3(cipher_text[103]), .A4(
        n289), .A5(adk_out0[103]), .A6(n290), .Y(n178) );
  AO222X1_HVT U218 ( .A1(n288), .A2(adk_in[104]), .A3(cipher_text[104]), .A4(
        n289), .A5(adk_out0[104]), .A6(n290), .Y(n177) );
  AO222X1_HVT U219 ( .A1(n288), .A2(adk_in[105]), .A3(cipher_text[105]), .A4(
        n289), .A5(adk_out0[105]), .A6(n290), .Y(n176) );
  AO222X1_HVT U220 ( .A1(n288), .A2(adk_in[106]), .A3(cipher_text[106]), .A4(
        n289), .A5(adk_out0[106]), .A6(n290), .Y(n175) );
  AO222X1_HVT U221 ( .A1(n288), .A2(adk_in[107]), .A3(cipher_text[107]), .A4(
        n289), .A5(adk_out0[107]), .A6(n290), .Y(n174) );
  AO222X1_HVT U222 ( .A1(n288), .A2(adk_in[108]), .A3(cipher_text[108]), .A4(
        n289), .A5(adk_out0[108]), .A6(n290), .Y(n173) );
  AO222X1_HVT U223 ( .A1(n288), .A2(adk_in[109]), .A3(cipher_text[109]), .A4(
        n289), .A5(adk_out0[109]), .A6(n290), .Y(n172) );
  AO222X1_HVT U224 ( .A1(n288), .A2(adk_in[110]), .A3(cipher_text[110]), .A4(
        n289), .A5(adk_out0[110]), .A6(n290), .Y(n171) );
  AO222X1_HVT U225 ( .A1(n288), .A2(adk_in[111]), .A3(cipher_text[111]), .A4(
        n289), .A5(adk_out0[111]), .A6(n290), .Y(n170) );
  AO222X1_HVT U226 ( .A1(n288), .A2(adk_in[112]), .A3(cipher_text[112]), .A4(
        n289), .A5(adk_out0[112]), .A6(n290), .Y(n169) );
  AO222X1_HVT U227 ( .A1(n288), .A2(adk_in[113]), .A3(cipher_text[113]), .A4(
        n289), .A5(adk_out0[113]), .A6(n290), .Y(n168) );
  AO222X1_HVT U228 ( .A1(n288), .A2(adk_in[114]), .A3(cipher_text[114]), .A4(
        n289), .A5(adk_out0[114]), .A6(n290), .Y(n167) );
  AO222X1_HVT U229 ( .A1(n288), .A2(adk_in[115]), .A3(cipher_text[115]), .A4(
        n289), .A5(adk_out0[115]), .A6(n290), .Y(n166) );
  AO222X1_HVT U230 ( .A1(n288), .A2(adk_in[116]), .A3(cipher_text[116]), .A4(
        n289), .A5(adk_out0[116]), .A6(n290), .Y(n165) );
  AO222X1_HVT U231 ( .A1(n288), .A2(adk_in[117]), .A3(cipher_text[117]), .A4(
        n289), .A5(adk_out0[117]), .A6(n290), .Y(n164) );
  AO222X1_HVT U232 ( .A1(n288), .A2(adk_in[118]), .A3(cipher_text[118]), .A4(
        n289), .A5(adk_out0[118]), .A6(n290), .Y(n163) );
  AO222X1_HVT U233 ( .A1(n288), .A2(adk_in[119]), .A3(cipher_text[119]), .A4(
        n289), .A5(adk_out0[119]), .A6(n290), .Y(n162) );
  AO222X1_HVT U234 ( .A1(n288), .A2(adk_in[120]), .A3(cipher_text[120]), .A4(
        n289), .A5(adk_out0[120]), .A6(n290), .Y(n161) );
  AO222X1_HVT U235 ( .A1(n288), .A2(adk_in[121]), .A3(cipher_text[121]), .A4(
        n289), .A5(adk_out0[121]), .A6(n290), .Y(n160) );
  AO222X1_HVT U236 ( .A1(n288), .A2(adk_in[122]), .A3(cipher_text[122]), .A4(
        n289), .A5(adk_out0[122]), .A6(n290), .Y(n159) );
  AO222X1_HVT U237 ( .A1(n288), .A2(adk_in[123]), .A3(cipher_text[123]), .A4(
        n289), .A5(adk_out0[123]), .A6(n290), .Y(n158) );
  AO222X1_HVT U238 ( .A1(n288), .A2(adk_in[124]), .A3(cipher_text[124]), .A4(
        n289), .A5(adk_out0[124]), .A6(n290), .Y(n157) );
  AO222X1_HVT U239 ( .A1(n288), .A2(adk_in[125]), .A3(cipher_text[125]), .A4(
        n289), .A5(adk_out0[125]), .A6(n290), .Y(n156) );
  AO222X1_HVT U240 ( .A1(n288), .A2(adk_in[126]), .A3(cipher_text[126]), .A4(
        n289), .A5(adk_out0[126]), .A6(n290), .Y(n155) );
  AO222X1_HVT U241 ( .A1(n288), .A2(adk_in[127]), .A3(cipher_text[127]), .A4(
        n289), .A5(adk_out0[127]), .A6(n290), .Y(n154) );
  AO222X1_HVT U242 ( .A1(n288), .A2(key_round[1]), .A3(keyout[1]), .A4(n289), 
        .A5(key[1]), .A6(n290), .Y(n153) );
  AO222X1_HVT U243 ( .A1(n288), .A2(key_round[2]), .A3(keyout[2]), .A4(n289), 
        .A5(key[2]), .A6(n290), .Y(n152) );
  AO222X1_HVT U244 ( .A1(n288), .A2(key_round[3]), .A3(keyout[3]), .A4(n289), 
        .A5(key[3]), .A6(n290), .Y(n151) );
  AO222X1_HVT U245 ( .A1(n288), .A2(key_round[4]), .A3(keyout[4]), .A4(n289), 
        .A5(key[4]), .A6(n290), .Y(n150) );
  AO222X1_HVT U246 ( .A1(n288), .A2(key_round[5]), .A3(keyout[5]), .A4(n289), 
        .A5(key[5]), .A6(n290), .Y(n149) );
  AO222X1_HVT U247 ( .A1(n288), .A2(key_round[6]), .A3(keyout[6]), .A4(n289), 
        .A5(key[6]), .A6(n290), .Y(n148) );
  AO222X1_HVT U248 ( .A1(n288), .A2(key_round[7]), .A3(keyout[7]), .A4(n289), 
        .A5(key[7]), .A6(n290), .Y(n147) );
  AO222X1_HVT U249 ( .A1(n288), .A2(key_round[8]), .A3(keyout[8]), .A4(n289), 
        .A5(key[8]), .A6(n290), .Y(n146) );
  AO222X1_HVT U250 ( .A1(n288), .A2(key_round[9]), .A3(keyout[9]), .A4(n289), 
        .A5(key[9]), .A6(n290), .Y(n145) );
  AO222X1_HVT U251 ( .A1(n288), .A2(key_round[10]), .A3(keyout[10]), .A4(n289), 
        .A5(key[10]), .A6(n290), .Y(n144) );
  AO222X1_HVT U252 ( .A1(n288), .A2(key_round[11]), .A3(keyout[11]), .A4(n289), 
        .A5(key[11]), .A6(n290), .Y(n143) );
  AO222X1_HVT U253 ( .A1(n288), .A2(key_round[12]), .A3(keyout[12]), .A4(n289), 
        .A5(key[12]), .A6(n290), .Y(n142) );
  AO222X1_HVT U254 ( .A1(n288), .A2(key_round[13]), .A3(keyout[13]), .A4(n289), 
        .A5(key[13]), .A6(n290), .Y(n141) );
  AO222X1_HVT U255 ( .A1(n288), .A2(key_round[14]), .A3(keyout[14]), .A4(n289), 
        .A5(key[14]), .A6(n290), .Y(n140) );
  AO222X1_HVT U256 ( .A1(n288), .A2(key_round[15]), .A3(keyout[15]), .A4(n289), 
        .A5(key[15]), .A6(n290), .Y(n139) );
  AO222X1_HVT U257 ( .A1(n288), .A2(key_round[16]), .A3(keyout[16]), .A4(n289), 
        .A5(key[16]), .A6(n290), .Y(n138) );
  AO222X1_HVT U258 ( .A1(n288), .A2(key_round[17]), .A3(keyout[17]), .A4(n289), 
        .A5(key[17]), .A6(n290), .Y(n137) );
  AO222X1_HVT U259 ( .A1(n288), .A2(key_round[18]), .A3(keyout[18]), .A4(n289), 
        .A5(key[18]), .A6(n290), .Y(n136) );
  AO222X1_HVT U260 ( .A1(n288), .A2(key_round[19]), .A3(keyout[19]), .A4(n289), 
        .A5(key[19]), .A6(n290), .Y(n135) );
  AO222X1_HVT U261 ( .A1(n288), .A2(key_round[20]), .A3(keyout[20]), .A4(n289), 
        .A5(key[20]), .A6(n290), .Y(n134) );
  AO222X1_HVT U262 ( .A1(n288), .A2(key_round[21]), .A3(keyout[21]), .A4(n289), 
        .A5(key[21]), .A6(n290), .Y(n133) );
  AO222X1_HVT U263 ( .A1(n288), .A2(key_round[22]), .A3(keyout[22]), .A4(n289), 
        .A5(key[22]), .A6(n290), .Y(n132) );
  AO222X1_HVT U264 ( .A1(n288), .A2(key_round[23]), .A3(keyout[23]), .A4(n289), 
        .A5(key[23]), .A6(n290), .Y(n131) );
  AO222X1_HVT U265 ( .A1(n288), .A2(key_round[24]), .A3(keyout[24]), .A4(n289), 
        .A5(key[24]), .A6(n290), .Y(n130) );
  AO222X1_HVT U266 ( .A1(n288), .A2(key_round[25]), .A3(keyout[25]), .A4(n289), 
        .A5(key[25]), .A6(n290), .Y(n129) );
  AO222X1_HVT U267 ( .A1(n288), .A2(key_round[26]), .A3(keyout[26]), .A4(n289), 
        .A5(key[26]), .A6(n290), .Y(n128) );
  AO222X1_HVT U268 ( .A1(n288), .A2(key_round[27]), .A3(keyout[27]), .A4(n289), 
        .A5(key[27]), .A6(n290), .Y(n127) );
  AO222X1_HVT U269 ( .A1(n288), .A2(key_round[28]), .A3(keyout[28]), .A4(n289), 
        .A5(key[28]), .A6(n290), .Y(n126) );
  AO222X1_HVT U270 ( .A1(n288), .A2(key_round[29]), .A3(keyout[29]), .A4(n289), 
        .A5(key[29]), .A6(n290), .Y(n125) );
  AO222X1_HVT U271 ( .A1(n288), .A2(key_round[30]), .A3(keyout[30]), .A4(n289), 
        .A5(key[30]), .A6(n290), .Y(n124) );
  AO222X1_HVT U272 ( .A1(n288), .A2(key_round[31]), .A3(keyout[31]), .A4(n289), 
        .A5(key[31]), .A6(n290), .Y(n123) );
  AO222X1_HVT U273 ( .A1(n288), .A2(key_round[32]), .A3(keyout[32]), .A4(n289), 
        .A5(key[32]), .A6(n290), .Y(n122) );
  AO222X1_HVT U274 ( .A1(n288), .A2(key_round[33]), .A3(keyout[33]), .A4(n289), 
        .A5(key[33]), .A6(n290), .Y(n121) );
  AO222X1_HVT U275 ( .A1(n288), .A2(key_round[34]), .A3(keyout[34]), .A4(n289), 
        .A5(key[34]), .A6(n290), .Y(n120) );
  AO222X1_HVT U276 ( .A1(n288), .A2(key_round[35]), .A3(keyout[35]), .A4(n289), 
        .A5(key[35]), .A6(n290), .Y(n119) );
  AO222X1_HVT U277 ( .A1(n288), .A2(key_round[36]), .A3(keyout[36]), .A4(n289), 
        .A5(key[36]), .A6(n290), .Y(n118) );
  AO222X1_HVT U278 ( .A1(n288), .A2(key_round[37]), .A3(keyout[37]), .A4(n289), 
        .A5(key[37]), .A6(n290), .Y(n117) );
  AO222X1_HVT U279 ( .A1(n288), .A2(key_round[38]), .A3(keyout[38]), .A4(n289), 
        .A5(key[38]), .A6(n290), .Y(n116) );
  AO222X1_HVT U280 ( .A1(n288), .A2(key_round[39]), .A3(keyout[39]), .A4(n289), 
        .A5(key[39]), .A6(n290), .Y(n115) );
  AO222X1_HVT U281 ( .A1(n288), .A2(key_round[40]), .A3(keyout[40]), .A4(n289), 
        .A5(key[40]), .A6(n290), .Y(n114) );
  AO222X1_HVT U282 ( .A1(n288), .A2(key_round[41]), .A3(keyout[41]), .A4(n289), 
        .A5(key[41]), .A6(n290), .Y(n113) );
  AO222X1_HVT U283 ( .A1(n288), .A2(key_round[42]), .A3(keyout[42]), .A4(n289), 
        .A5(key[42]), .A6(n290), .Y(n112) );
  AO222X1_HVT U284 ( .A1(n288), .A2(key_round[43]), .A3(keyout[43]), .A4(n289), 
        .A5(key[43]), .A6(n290), .Y(n111) );
  AO222X1_HVT U285 ( .A1(n288), .A2(key_round[44]), .A3(keyout[44]), .A4(n289), 
        .A5(key[44]), .A6(n290), .Y(n110) );
  AO222X1_HVT U286 ( .A1(n288), .A2(key_round[45]), .A3(keyout[45]), .A4(n289), 
        .A5(key[45]), .A6(n290), .Y(n109) );
  AO222X1_HVT U287 ( .A1(n288), .A2(key_round[46]), .A3(keyout[46]), .A4(n289), 
        .A5(key[46]), .A6(n290), .Y(n108) );
  AO222X1_HVT U288 ( .A1(n288), .A2(key_round[47]), .A3(keyout[47]), .A4(n289), 
        .A5(key[47]), .A6(n290), .Y(n107) );
  AO222X1_HVT U289 ( .A1(n288), .A2(key_round[48]), .A3(keyout[48]), .A4(n289), 
        .A5(key[48]), .A6(n290), .Y(n106) );
  AO222X1_HVT U290 ( .A1(n288), .A2(key_round[49]), .A3(keyout[49]), .A4(n289), 
        .A5(key[49]), .A6(n290), .Y(n105) );
  AO222X1_HVT U291 ( .A1(n288), .A2(key_round[50]), .A3(keyout[50]), .A4(n289), 
        .A5(key[50]), .A6(n290), .Y(n104) );
  AO222X1_HVT U292 ( .A1(n288), .A2(key_round[51]), .A3(keyout[51]), .A4(n289), 
        .A5(key[51]), .A6(n290), .Y(n103) );
  AO222X1_HVT U293 ( .A1(n288), .A2(key_round[52]), .A3(keyout[52]), .A4(n289), 
        .A5(key[52]), .A6(n290), .Y(n102) );
  AO222X1_HVT U294 ( .A1(n288), .A2(key_round[53]), .A3(keyout[53]), .A4(n289), 
        .A5(key[53]), .A6(n290), .Y(n101) );
  AO222X1_HVT U295 ( .A1(n288), .A2(key_round[54]), .A3(keyout[54]), .A4(n289), 
        .A5(key[54]), .A6(n290), .Y(n100) );
  INVX0_HVT U296 ( .A(n302), .Y(n290) );
  AND2X1_HVT U297 ( .A1(n302), .A2(n296), .Y(n289) );
  OR3X1_HVT U298 ( .A1(round_number[0]), .A2(round_number[3]), .A3(n303), .Y(
        n302) );
  INVX0_HVT U299 ( .A(n296), .Y(n288) );
  NAND2X0_HVT U300 ( .A1(round_number[3]), .A2(n303), .Y(n296) );
  NAND2X0_HVT U301 ( .A1(n1), .A2(n4), .Y(n303) );
endmodule

