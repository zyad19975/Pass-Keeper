
module inv_sbox_5 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n196, n197, n198, n199, n200, n201, n202, n203, n208, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629;

  NAND2X0_HVT U1 ( .A1(n297), .A2(n335), .Y(n629) );
  NAND2X0_HVT U4 ( .A1(n355), .A2(n349), .Y(n626) );
  NAND2X0_HVT U5 ( .A1(n626), .A2(n345), .Y(n625) );
  NAND2X0_HVT U7 ( .A1(n353), .A2(n346), .Y(n622) );
  NAND2X0_HVT U8 ( .A1(n354), .A2(n344), .Y(n621) );
  NAND2X0_HVT U9 ( .A1(n352), .A2(n621), .Y(n620) );
  NAND2X0_HVT U10 ( .A1(n351), .A2(n618), .Y(n619) );
  NAND2X0_HVT U11 ( .A1(n239), .A2(n350), .Y(n617) );
  NAND2X0_HVT U12 ( .A1(n354), .A2(n244), .Y(n616) );
  NAND2X0_HVT U13 ( .A1(n347), .A2(n621), .Y(n615) );
  NAND2X0_HVT U15 ( .A1(n342), .A2(n354), .Y(n613) );
  NAND2X0_HVT U19 ( .A1(n353), .A2(n421), .Y(n608) );
  NAND2X0_HVT U25 ( .A1(n307), .A2(n419), .Y(n624) );
  NAND2X0_HVT U32 ( .A1(n335), .A2(n239), .Y(n596) );
  NAND2X0_HVT U35 ( .A1(n208), .A2(n263), .Y(n593) );
  NAND2X0_HVT U38 ( .A1(n244), .A2(n258), .Y(n590) );
  NAND2X0_HVT U42 ( .A1(n623), .A2(n278), .Y(n586) );
  OA21X1_HVT U53 ( .A1(n283), .A2(n578), .A3(n390), .Y(n576) );
  NAND2X0_HVT U55 ( .A1(n347), .A2(n626), .Y(n574) );
  MUX41X1_HVT U56 ( .A1(n304), .A3(n341), .A2(n388), .A4(n231), .S0(n326), 
        .S1(n361), .Y(n573) );
  MUX41X1_HVT U65 ( .A1(n382), .A3(n384), .A2(n383), .A4(n590), .S0(n326), 
        .S1(n282), .Y(n563) );
  NAND2X0_HVT U66 ( .A1(n254), .A2(n198), .Y(n562) );
  MUX41X1_HVT U67 ( .A1(n379), .A3(n403), .A2(n381), .A4(n562), .S0(n332), 
        .S1(n324), .Y(n561) );
  NAND2X0_HVT U72 ( .A1(n343), .A2(n622), .Y(n557) );
  MUX41X1_HVT U73 ( .A1(n601), .A3(n557), .A2(n404), .A4(n333), .S0(n331), 
        .S1(n323), .Y(n556) );
  MUX41X1_HVT U74 ( .A1(n619), .A3(n395), .A2(n394), .A4(n196), .S0(n326), 
        .S1(n281), .Y(n555) );
  MUX41X1_HVT U80 ( .A1(n406), .A3(n304), .A2(n203), .A4(n625), .S0(n326), 
        .S1(n274), .Y(n549) );
  NAND2X0_HVT U81 ( .A1(n350), .A2(n622), .Y(n548) );
  AND2X1_HVT U82 ( .A1(n623), .A2(n348), .Y(n547) );
  MUX41X1_HVT U83 ( .A1(n547), .A3(n392), .A2(n312), .A4(n548), .S0(n324), 
        .S1(n361), .Y(n546) );
  MUX41X1_HVT U88 ( .A1(n381), .A3(n366), .A2(n598), .A4(n582), .S0(n256), 
        .S1(n361), .Y(n542) );
  NAND2X0_HVT U89 ( .A1(n258), .A2(n418), .Y(n541) );
  MUX41X1_HVT U90 ( .A1(n420), .A3(n622), .A2(n581), .A4(n541), .S0(n324), 
        .S1(n281), .Y(n540) );
  MUX41X1_HVT U96 ( .A1(n403), .A3(n615), .A2(n389), .A4(n409), .S0(n326), 
        .S1(n361), .Y(n534) );
  MUX41X1_HVT U99 ( .A1(n596), .A3(n383), .A2(n580), .A4(n341), .S0(n361), 
        .S1(n324), .Y(n531) );
  NAND2X0_HVT U100 ( .A1(n242), .A2(n310), .Y(n530) );
  AND2X1_HVT U104 ( .A1(n622), .A2(n345), .Y(n527) );
  MUX41X1_HVT U105 ( .A1(n614), .A3(n412), .A2(n548), .A4(n527), .S0(n326), 
        .S1(n281), .Y(n526) );
  MUX41X1_HVT U107 ( .A1(n411), .A3(n347), .A2(n525), .A4(n372), .S0(n326), 
        .S1(n281), .Y(n524) );
  MUX41X1_HVT U108 ( .A1(n196), .A3(n341), .A2(n388), .A4(n299), .S0(n326), 
        .S1(n282), .Y(n523) );
  MUX41X1_HVT U109 ( .A1(n410), .A3(n366), .A2(n407), .A4(n401), .S0(n256), 
        .S1(n282), .Y(n522) );
  MUX41X1_HVT U110 ( .A1(n522), .A3(n524), .A2(n523), .A4(n526), .S0(n340), 
        .S1(n338), .Y(n521) );
  AO21X1_HVT U112 ( .A1(n398), .A2(n331), .A3(n604), .Y(n519) );
  NAND2X0_HVT U114 ( .A1(n629), .A2(n622), .Y(n517) );
  MUX41X1_HVT U115 ( .A1(n517), .A3(n617), .A2(n398), .A4(n348), .S0(n281), 
        .S1(n324), .Y(n516) );
  MUX41X1_HVT U116 ( .A1(n397), .A3(n391), .A2(n366), .A4(n613), .S0(n325), 
        .S1(n281), .Y(n515) );
  NAND2X0_HVT U118 ( .A1(n258), .A2(n297), .Y(n513) );
  MUX41X1_HVT U119 ( .A1(n413), .A3(n514), .A2(n591), .A4(n513), .S0(n325), 
        .S1(n274), .Y(n512) );
  MUX41X1_HVT U120 ( .A1(n512), .A3(n516), .A2(n515), .A4(n518), .S0(n340), 
        .S1(n338), .Y(n511) );
  MUX41X1_HVT U122 ( .A1(n402), .A3(n314), .A2(n582), .A4(n405), .S0(n325), 
        .S1(n282), .Y(n510) );
  MUX41X1_HVT U124 ( .A1(n317), .A3(n509), .A2(n605), .A4(n284), .S0(n330), 
        .S1(n325), .Y(n508) );
  AOI21X1_HVT U127 ( .A1(n329), .A2(n504), .A3(n373), .Y(n505) );
  NAND2X0_HVT U129 ( .A1(n328), .A2(n351), .Y(n502) );
  MUX41X1_HVT U130 ( .A1(n502), .A3(n503), .A2(n506), .A4(n505), .S0(n332), 
        .S1(n338), .Y(n501) );
  AND2X1_HVT U131 ( .A1(n198), .A2(n258), .Y(n500) );
  MUX41X1_HVT U132 ( .A1(n370), .A3(n500), .A2(n415), .A4(n379), .S0(n331), 
        .S1(n323), .Y(n499) );
  MUX41X1_HVT U133 ( .A1(n416), .A3(n372), .A2(n231), .A4(n371), .S0(n330), 
        .S1(n322), .Y(n498) );
  MUX41X1_HVT U136 ( .A1(n579), .A3(n530), .A2(n496), .A4(n377), .S0(n328), 
        .S1(n361), .Y(n495) );
  MUX41X1_HVT U137 ( .A1(n208), .A3(n235), .A2(n603), .A4(n409), .S0(n332), 
        .S1(n322), .Y(n494) );
  MUX41X1_HVT U139 ( .A1(n493), .A3(n497), .A2(n501), .A4(n507), .S0(n340), 
        .S1(n261), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n394), .A3(n315), .A2(n387), .A4(n617), .S0(n331), 
        .S1(n324), .Y(n492) );
  NAND2X0_HVT U141 ( .A1(n342), .A2(n258), .Y(n491) );
  MUX41X1_HVT U142 ( .A1(n491), .A3(n589), .A2(n414), .A4(n387), .S0(n329), 
        .S1(n282), .Y(n490) );
  MUX41X1_HVT U143 ( .A1(n418), .A3(n399), .A2(n608), .A4(n605), .S0(n327), 
        .S1(n360), .Y(n489) );
  MUX41X1_HVT U145 ( .A1(n597), .A3(n412), .A2(n488), .A4(n548), .S0(n329), 
        .S1(n361), .Y(n487) );
  OA21X1_HVT U153 ( .A1(n367), .A2(n283), .A3(n376), .Y(n479) );
  MUX41X1_HVT U155 ( .A1(n387), .A3(n617), .A2(n609), .A4(n389), .S0(n327), 
        .S1(n360), .Y(n477) );
  NAND2X0_HVT U159 ( .A1(n473), .A2(n472), .Y(n474) );
  NAND2X0_HVT U163 ( .A1(n253), .A2(n418), .Y(n468) );
  NAND2X0_HVT U166 ( .A1(n618), .A2(n464), .Y(n465) );
  MUX41X1_HVT U170 ( .A1(n319), .A3(n316), .A2(n317), .A4(n461), .S0(n327), 
        .S1(n282), .Y(n460) );
  MUX41X1_HVT U173 ( .A1(n352), .A3(n420), .A2(n299), .A4(n592), .S0(n327), 
        .S1(n360), .Y(n457) );
  NAND2X0_HVT U177 ( .A1(n353), .A2(n297), .Y(n454) );
  AND2X1_HVT U179 ( .A1(n623), .A2(n345), .Y(n452) );
  MUX41X1_HVT U180 ( .A1(n596), .A3(n364), .A2(n452), .A4(n583), .S0(n327), 
        .S1(n360), .Y(n451) );
  MUX41X1_HVT U182 ( .A1(n372), .A3(n232), .A2(n369), .A4(n312), .S0(n325), 
        .S1(n360), .Y(n449) );
  AND2X1_HVT U185 ( .A1(n278), .A2(n242), .Y(n446) );
  NAND2X0_HVT U191 ( .A1(n283), .A2(n378), .Y(n440) );
  AND2X1_HVT U192 ( .A1(n395), .A2(n438), .Y(n439) );
  NAND2X0_HVT U194 ( .A1(n586), .A2(n438), .Y(n436) );
  MUX41X1_HVT U195 ( .A1(n437), .A3(n436), .A2(n439), .A4(n440), .S0(n324), 
        .S1(n291), .Y(n435) );
  NAND2X0_HVT U198 ( .A1(n356), .A2(n278), .Y(n618) );
  NAND2X0_HVT U200 ( .A1(n345), .A2(n258), .Y(n504) );
  NAND2X0_HVT U207 ( .A1(n258), .A2(n420), .Y(n568) );
  OR2X1_HVT U2 ( .A1(n419), .A2(n306), .Y(n627) );
  INVX0_HVT U3 ( .A(n358), .Y(n357) );
  IBUFFX2_HVT U6 ( .A(n358), .Y(n356) );
  INVX1_HVT U14 ( .A(n358), .Y(n253) );
  INVX0_HVT U16 ( .A(n607), .Y(n196) );
  INVX0_HVT U17 ( .A(n607), .Y(n385) );
  MUX21X1_HVT U18 ( .A1(n342), .A2(n244), .S0(n257), .Y(n607) );
  MUX21X2_HVT U20 ( .A1(n344), .A2(n306), .S0(n305), .Y(n304) );
  IBUFFX2_HVT U21 ( .A(in[3]), .Y(n244) );
  MUX41X1_HVT U22 ( .A1(n304), .A3(n586), .A2(n399), .A4(n385), .S0(n199), 
        .S1(n224), .Y(n448) );
  INVX0_HVT U23 ( .A(n585), .Y(n399) );
  IBUFFX2_HVT U24 ( .A(n330), .Y(n224) );
  INVX1_HVT U26 ( .A(n225), .Y(n199) );
  MUX21X2_HVT U27 ( .A1(n350), .A2(n352), .S0(n197), .Y(n614) );
  IBUFFX16_HVT U28 ( .A(n353), .Y(n197) );
  MUX21X2_HVT U29 ( .A1(n343), .A2(n336), .S0(n357), .Y(n603) );
  XNOR2X2_HVT U30 ( .A1(n344), .A2(n305), .Y(n580) );
  OA21X1_HVT U31 ( .A1(n368), .A2(n303), .A3(n607), .Y(n553) );
  AO21X1_HVT U33 ( .A1(n568), .A2(n330), .A3(n607), .Y(n569) );
  INVX0_HVT U34 ( .A(n336), .Y(n198) );
  NBUFFX2_HVT U36 ( .A(n306), .Y(n336) );
  IBUFFX2_HVT U37 ( .A(n306), .Y(n307) );
  INVX1_HVT U39 ( .A(n419), .Y(n297) );
  MUX21X2_HVT U40 ( .A1(n391), .A2(n318), .S0(n255), .Y(n285) );
  INVX0_HVT U41 ( .A(n356), .Y(n239) );
  INVX0_HVT U43 ( .A(n254), .Y(n242) );
  NAND2X0_HVT U44 ( .A1(n585), .A2(n200), .Y(n201) );
  NAND2X0_HVT U45 ( .A1(n405), .A2(n331), .Y(n202) );
  NAND2X0_HVT U46 ( .A1(n201), .A2(n202), .Y(n475) );
  IBUFFX2_HVT U47 ( .A(n331), .Y(n200) );
  MUX21X1_HVT U48 ( .A1(n244), .A2(n421), .S0(n353), .Y(n585) );
  MUX21X1_HVT U49 ( .A1(n474), .A2(n475), .S0(n329), .Y(n471) );
  INVX1_HVT U50 ( .A(n243), .Y(n228) );
  IBUFFX2_HVT U51 ( .A(n339), .Y(n229) );
  INVX0_HVT U52 ( .A(n377), .Y(n203) );
  INVX1_HVT U54 ( .A(n374), .Y(n208) );
  INVX1_HVT U57 ( .A(n620), .Y(n377) );
  INVX1_HVT U58 ( .A(n621), .Y(n374) );
  INVX1_HVT U59 ( .A(n599), .Y(n391) );
  IBUFFX2_HVT U60 ( .A(n600), .Y(n390) );
  MUX21X2_HVT U61 ( .A1(n407), .A2(n603), .S0(n218), .Y(n286) );
  IBUFFX16_HVT U62 ( .A(n255), .Y(n218) );
  INVX1_HVT U63 ( .A(n358), .Y(n254) );
  INVX0_HVT U64 ( .A(n628), .Y(n219) );
  INVX1_HVT U68 ( .A(n219), .Y(n220) );
  MUX21X1_HVT U69 ( .A1(n299), .A2(n244), .S0(n357), .Y(n284) );
  NAND2X0_HVT U70 ( .A1(n297), .A2(n221), .Y(n222) );
  NAND2X0_HVT U71 ( .A1(n345), .A2(n239), .Y(n223) );
  NAND2X0_HVT U75 ( .A1(n222), .A2(n223), .Y(n533) );
  INVX0_HVT U76 ( .A(n239), .Y(n221) );
  MUX21X1_HVT U77 ( .A1(n284), .A2(n574), .S0(n331), .Y(n570) );
  MUX21X2_HVT U78 ( .A1(n351), .A2(n345), .S0(n239), .Y(n313) );
  MUX21X2_HVT U79 ( .A1(n334), .A2(n418), .S0(n254), .Y(n482) );
  INVX0_HVT U84 ( .A(n313), .Y(n584) );
  IBUFFX16_HVT U85 ( .A(n323), .Y(n225) );
  MUX41X1_HVT U86 ( .A1(n420), .A3(n623), .A2(n375), .A4(n617), .S0(n226), 
        .S1(n281), .Y(n558) );
  IBUFFX16_HVT U87 ( .A(n256), .Y(n226) );
  MUX21X2_HVT U91 ( .A1(n286), .A2(n285), .S0(n227), .Y(n545) );
  IBUFFX16_HVT U92 ( .A(n281), .Y(n227) );
  MUX41X1_HVT U93 ( .A1(n463), .A3(n467), .A2(n469), .A4(n471), .S0(n228), 
        .S1(n229), .Y(n462) );
  INVX0_HVT U94 ( .A(n574), .Y(n230) );
  INVX0_HVT U95 ( .A(n230), .Y(n231) );
  INVX1_HVT U97 ( .A(n369), .Y(n232) );
  INVX1_HVT U98 ( .A(n626), .Y(n369) );
  INVX1_HVT U101 ( .A(n292), .Y(n560) );
  IBUFFX2_HVT U102 ( .A(n337), .Y(n233) );
  OA21X1_HVT U103 ( .A1(n391), .A2(n287), .A3(n568), .Y(n442) );
  MUX41X1_HVT U106 ( .A1(n532), .A3(n529), .A2(n534), .A4(n531), .S0(n339), 
        .S1(n233), .Y(n528) );
  MUX41X1_HVT U111 ( .A1(n555), .A3(n558), .A2(n552), .A4(n556), .S0(n234), 
        .S1(n337), .Y(n551) );
  IBUFFX16_HVT U113 ( .A(n237), .Y(n234) );
  MUX41X1_HVT U117 ( .A1(n441), .A3(n435), .A2(n450), .A4(n447), .S0(n339), 
        .S1(n261), .Y(out[7]) );
  NBUFFX2_HVT U121 ( .A(n599), .Y(n235) );
  MUX21X2_HVT U123 ( .A1(n486), .A2(n476), .S0(n236), .Y(out[5]) );
  IBUFFX16_HVT U125 ( .A(n261), .Y(n236) );
  INVX1_HVT U126 ( .A(n594), .Y(n395) );
  IBUFFX16_HVT U128 ( .A(n340), .Y(n237) );
  MUX41X1_HVT U134 ( .A1(n458), .A3(n460), .A2(n456), .A4(n457), .S0(n238), 
        .S1(n339), .Y(n455) );
  IBUFFX16_HVT U135 ( .A(n337), .Y(n238) );
  IBUFFX2_HVT U138 ( .A(n220), .Y(n310) );
  MUX21X2_HVT U144 ( .A1(n420), .A2(n418), .S0(n253), .Y(n600) );
  MUX21X1_HVT U146 ( .A1(n466), .A2(n465), .S0(n290), .Y(n463) );
  NBUFFX2_HVT U147 ( .A(n362), .Y(n332) );
  INVX1_HVT U148 ( .A(n363), .Y(n362) );
  MUX41X1_HVT U149 ( .A1(n545), .A3(n549), .A2(n546), .A4(n550), .S0(in[5]), 
        .S1(n291), .Y(n544) );
  MUX21X2_HVT U150 ( .A1(n569), .A2(n570), .S0(n240), .Y(n567) );
  IBUFFX16_HVT U151 ( .A(n328), .Y(n240) );
  MUX21X1_HVT U152 ( .A1(n386), .A2(n572), .S0(n320), .Y(n571) );
  AO21X1_HVT U154 ( .A1(n254), .A2(n310), .A3(n287), .Y(n438) );
  INVX2_HVT U156 ( .A(n330), .Y(n287) );
  MUX21X2_HVT U157 ( .A1(n508), .A2(n510), .S0(n291), .Y(n507) );
  MUX41X1_HVT U158 ( .A1(n263), .A3(n416), .A2(n574), .A4(n408), .S0(n241), 
        .S1(n363), .Y(n456) );
  IBUFFX16_HVT U160 ( .A(n327), .Y(n241) );
  IBUFFX2_HVT U161 ( .A(n363), .Y(n360) );
  MUX21X2_HVT U162 ( .A1(n404), .A2(n587), .S0(n331), .Y(n443) );
  INVX1_HVT U164 ( .A(n344), .Y(n418) );
  MUX21X1_HVT U165 ( .A1(n405), .A2(n365), .S0(n332), .Y(n554) );
  MUX21X1_HVT U167 ( .A1(n333), .A2(n421), .S0(n242), .Y(n432) );
  INVX1_HVT U168 ( .A(n432), .Y(n405) );
  IBUFFX16_HVT U169 ( .A(n338), .Y(n243) );
  INVX1_HVT U171 ( .A(in[4]), .Y(n363) );
  INVX1_HVT U172 ( .A(n586), .Y(n372) );
  NAND2X0_HVT U174 ( .A1(n347), .A2(n354), .Y(n265) );
  NAND2X0_HVT U175 ( .A1(n253), .A2(n321), .Y(n623) );
  AO21X1_HVT U176 ( .A1(n343), .A2(n626), .A3(n303), .Y(n464) );
  NAND2X0_HVT U178 ( .A1(n519), .A2(n290), .Y(n247) );
  MUX21X1_HVT U181 ( .A1(n342), .A2(n264), .S0(n305), .Y(n311) );
  INVX0_HVT U183 ( .A(n352), .Y(n294) );
  INVX0_HVT U184 ( .A(n380), .Y(n293) );
  NAND2X0_HVT U186 ( .A1(n260), .A2(n259), .Y(n447) );
  MUX41X1_HVT U187 ( .A1(n369), .A3(n318), .A2(n408), .A4(n388), .S0(n325), 
        .S1(n282), .Y(n543) );
  INVX1_HVT U188 ( .A(in[1]), .Y(n337) );
  INVX1_HVT U189 ( .A(n328), .Y(n290) );
  INVX0_HVT U190 ( .A(n358), .Y(n353) );
  INVX1_HVT U193 ( .A(n341), .Y(n278) );
  INVX1_HVT U196 ( .A(n342), .Y(n263) );
  INVX1_HVT U197 ( .A(n336), .Y(n264) );
  INVX1_HVT U199 ( .A(n302), .Y(n261) );
  INVX0_HVT U201 ( .A(in[7]), .Y(n302) );
  INVX1_HVT U202 ( .A(n283), .Y(n274) );
  INVX0_HVT U203 ( .A(n331), .Y(n283) );
  INVX1_HVT U204 ( .A(n322), .Y(n255) );
  INVX0_HVT U205 ( .A(n309), .Y(n256) );
  INVX1_HVT U206 ( .A(n327), .Y(n309) );
  INVX1_HVT U208 ( .A(n337), .Y(n338) );
  INVX1_HVT U209 ( .A(n337), .Y(n291) );
  INVX1_HVT U210 ( .A(in[6]), .Y(n306) );
  MUX41X1_HVT U211 ( .A1(n575), .A3(n571), .A2(n573), .A4(n567), .S0(n339), 
        .S1(n337), .Y(n566) );
  MUX21X2_HVT U212 ( .A1(n554), .A2(n553), .S0(n329), .Y(n552) );
  MUX21X2_HVT U213 ( .A1(n577), .A2(n576), .S0(n328), .Y(n575) );
  NAND2X0_HVT U214 ( .A1(n484), .A2(n326), .Y(n245) );
  NAND2X0_HVT U215 ( .A1(n485), .A2(n309), .Y(n246) );
  NAND2X0_HVT U216 ( .A1(n245), .A2(n246), .Y(n483) );
  AO21X2_HVT U217 ( .A1(n332), .A2(n374), .A3(n310), .Y(n484) );
  NAND2X0_HVT U218 ( .A1(n520), .A2(n329), .Y(n248) );
  NAND2X0_HVT U219 ( .A1(n247), .A2(n248), .Y(n518) );
  NAND2X2_HVT U220 ( .A1(n521), .A2(n261), .Y(n249) );
  NAND2X0_HVT U221 ( .A1(n511), .A2(n302), .Y(n250) );
  NAND2X0_HVT U222 ( .A1(n249), .A2(n250), .Y(out[3]) );
  MUX41X1_HVT U223 ( .A1(n536), .A3(n540), .A2(n542), .A4(n543), .S0(n338), 
        .S1(n340), .Y(n535) );
  NAND2X0_HVT U224 ( .A1(n538), .A2(n326), .Y(n251) );
  NAND2X0_HVT U225 ( .A1(n537), .A2(n290), .Y(n252) );
  NAND2X0_HVT U226 ( .A1(n251), .A2(n252), .Y(n536) );
  INVX1_HVT U227 ( .A(n339), .Y(n340) );
  INVX0_HVT U228 ( .A(n332), .Y(n303) );
  MUX21X1_HVT U229 ( .A1(n318), .A2(n580), .S0(n332), .Y(n444) );
  NBUFFX4_HVT U230 ( .A(n362), .Y(n330) );
  MUX21X1_HVT U231 ( .A1(n344), .A2(n348), .S0(n253), .Y(n470) );
  INVX1_HVT U232 ( .A(n358), .Y(n354) );
  INVX1_HVT U233 ( .A(n358), .Y(n355) );
  MUX41X1_HVT U234 ( .A1(n311), .A3(n530), .A2(n411), .A4(n616), .S0(n282), 
        .S1(n255), .Y(n529) );
  IBUFFX2_HVT U235 ( .A(n623), .Y(n371) );
  MUX41X1_HVT U236 ( .A1(n444), .A3(n443), .A2(n445), .A4(n442), .S0(n337), 
        .S1(n256), .Y(n441) );
  INVX0_HVT U237 ( .A(n358), .Y(n257) );
  INVX1_HVT U238 ( .A(n354), .Y(n258) );
  MUX41X1_HVT U239 ( .A1(n298), .A3(n482), .A2(n312), .A4(n396), .S0(n330), 
        .S1(n255), .Y(n481) );
  MUX41X1_HVT U240 ( .A1(n454), .A3(n319), .A2(n584), .A4(n420), .S0(n290), 
        .S1(n360), .Y(n453) );
  INVX1_HVT U241 ( .A(n262), .Y(n539) );
  INVX1_HVT U242 ( .A(n298), .Y(n606) );
  MUX41X1_HVT U243 ( .A1(n313), .A3(n384), .A2(n593), .A4(n470), .S0(n327), 
        .S1(n361), .Y(n469) );
  NAND2X0_HVT U244 ( .A1(n449), .A2(n338), .Y(n259) );
  NAND2X0_HVT U245 ( .A1(n448), .A2(n337), .Y(n260) );
  MUX41X1_HVT U246 ( .A1(n481), .A3(n477), .A2(n483), .A4(n478), .S0(n339), 
        .S1(n291), .Y(n476) );
  AO21X2_HVT U247 ( .A1(n258), .A2(n352), .A3(n283), .Y(n472) );
  MUX21X1_HVT U248 ( .A1(n263), .A2(n264), .S0(n331), .Y(n262) );
  INVX1_HVT U249 ( .A(n277), .Y(n312) );
  INVX1_HVT U250 ( .A(n433), .Y(n404) );
  NAND2X0_HVT U251 ( .A1(n539), .A2(n258), .Y(n266) );
  NAND2X0_HVT U252 ( .A1(n265), .A2(n266), .Y(n538) );
  NAND2X0_HVT U253 ( .A1(n196), .A2(n267), .Y(n268) );
  NAND2X0_HVT U254 ( .A1(n565), .A2(n320), .Y(n269) );
  NAND2X0_HVT U255 ( .A1(n268), .A2(n269), .Y(n564) );
  INVX0_HVT U256 ( .A(n320), .Y(n267) );
  NAND2X0_HVT U257 ( .A1(n566), .A2(in[7]), .Y(n270) );
  NAND2X0_HVT U258 ( .A1(n559), .A2(n302), .Y(n271) );
  NAND2X0_HVT U259 ( .A1(n270), .A2(n271), .Y(out[0]) );
  MUX21X1_HVT U260 ( .A1(n232), .A2(n298), .S0(n309), .Y(n565) );
  NAND2X0_HVT U261 ( .A1(n451), .A2(n337), .Y(n272) );
  NAND2X0_HVT U262 ( .A1(n453), .A2(n338), .Y(n273) );
  NAND2X0_HVT U263 ( .A1(n273), .A2(n272), .Y(n450) );
  NAND2X0_HVT U264 ( .A1(n318), .A2(n274), .Y(n275) );
  NAND2X0_HVT U265 ( .A1(n603), .A2(n283), .Y(n276) );
  NAND2X0_HVT U266 ( .A1(n275), .A2(n276), .Y(n480) );
  MUX21X1_HVT U267 ( .A1(n278), .A2(n333), .S0(n305), .Y(n277) );
  NAND2X0_HVT U268 ( .A1(n462), .A2(n261), .Y(n279) );
  NAND2X0_HVT U269 ( .A1(n455), .A2(n302), .Y(n280) );
  NAND2X0_HVT U270 ( .A1(n279), .A2(n280), .Y(out[6]) );
  INVX1_HVT U271 ( .A(n363), .Y(n281) );
  INVX1_HVT U272 ( .A(n363), .Y(n282) );
  IBUFFX2_HVT U273 ( .A(n603), .Y(n387) );
  INVX0_HVT U274 ( .A(n284), .Y(n605) );
  MUX41X1_HVT U275 ( .A1(n468), .A3(n620), .A2(n385), .A4(n591), .S0(n255), 
        .S1(n360), .Y(n467) );
  INVX2_HVT U276 ( .A(n363), .Y(n361) );
  NAND2X0_HVT U277 ( .A1(n602), .A2(n287), .Y(n288) );
  NAND2X0_HVT U278 ( .A1(n605), .A2(n330), .Y(n289) );
  NAND2X0_HVT U279 ( .A1(n288), .A2(n289), .Y(n466) );
  MUX41X1_HVT U280 ( .A1(n490), .A3(n492), .A2(n487), .A4(n489), .S0(n291), 
        .S1(n339), .Y(n486) );
  MUX41X1_HVT U281 ( .A1(n294), .A3(n293), .A2(n244), .A4(n614), .S0(n255), 
        .S1(n303), .Y(n292) );
  NAND2X0_HVT U282 ( .A1(n544), .A2(n302), .Y(n295) );
  NAND2X0_HVT U283 ( .A1(n551), .A2(in[7]), .Y(n296) );
  NAND2X0_HVT U284 ( .A1(n295), .A2(n296), .Y(out[1]) );
  NBUFFX2_HVT U285 ( .A(n419), .Y(n333) );
  INVX0_HVT U286 ( .A(n311), .Y(n592) );
  INVX0_HVT U287 ( .A(n308), .Y(n461) );
  MUX21X1_HVT U288 ( .A1(n415), .A2(n370), .S0(n330), .Y(n485) );
  INVX1_HVT U289 ( .A(n355), .Y(n305) );
  INVX1_HVT U290 ( .A(n417), .Y(n299) );
  MUX21X2_HVT U291 ( .A1(n479), .A2(n480), .S0(n329), .Y(n478) );
  INVX1_HVT U292 ( .A(in[0]), .Y(n358) );
  MUX41X1_HVT U293 ( .A1(n611), .A3(n393), .A2(n610), .A4(n391), .S0(n309), 
        .S1(n287), .Y(n550) );
  INVX0_HVT U294 ( .A(in[3]), .Y(n419) );
  MUX21X1_HVT U295 ( .A1(n350), .A2(n342), .S0(n239), .Y(n298) );
  INVX0_HVT U296 ( .A(n628), .Y(n417) );
  NAND2X0_HVT U297 ( .A1(n535), .A2(n261), .Y(n300) );
  NAND2X0_HVT U298 ( .A1(n528), .A2(n302), .Y(n301) );
  NAND2X0_HVT U299 ( .A1(n301), .A2(n300), .Y(out[2]) );
  MUX41X1_HVT U300 ( .A1(n600), .A3(n396), .A2(n410), .A4(n533), .S0(n309), 
        .S1(n303), .Y(n532) );
  XOR2X1_HVT U301 ( .A1(n334), .A2(in[3]), .Y(n612) );
  MUX21X1_HVT U302 ( .A1(n348), .A2(n321), .S0(n242), .Y(n308) );
  INVX1_HVT U303 ( .A(n346), .Y(n421) );
  INVX1_HVT U304 ( .A(n321), .Y(n420) );
  MUX41X1_HVT U305 ( .A1(n606), .A3(n316), .A2(n459), .A4(n541), .S0(n309), 
        .S1(n287), .Y(n458) );
  NBUFFX2_HVT U306 ( .A(n629), .Y(n351) );
  MUX41X1_HVT U307 ( .A1(n564), .A3(n561), .A2(n563), .A4(n560), .S0(n339), 
        .S1(n337), .Y(n559) );
  INVX1_HVT U308 ( .A(in[5]), .Y(n339) );
  INVX1_HVT U309 ( .A(n595), .Y(n394) );
  INVX1_HVT U310 ( .A(n422), .Y(n416) );
  NBUFFX2_HVT U311 ( .A(n220), .Y(n349) );
  NBUFFX2_HVT U312 ( .A(n220), .Y(n350) );
  AND2X1_HVT U313 ( .A1(n349), .A2(n613), .Y(n314) );
  MUX21X1_HVT U314 ( .A1(n400), .A2(n317), .S0(n330), .Y(n437) );
  MUX21X1_HVT U315 ( .A1(n310), .A2(n263), .S0(n357), .Y(n595) );
  NAND2X0_HVT U316 ( .A1(n333), .A2(n334), .Y(n628) );
  MUX21X1_HVT U317 ( .A1(n263), .A2(n244), .S0(n257), .Y(n589) );
  MUX21X1_HVT U318 ( .A1(n342), .A2(n420), .S0(n253), .Y(n597) );
  MUX21X1_HVT U319 ( .A1(n335), .A2(n417), .S0(n254), .Y(n602) );
  MUX21X1_HVT U320 ( .A1(n420), .A2(n336), .S0(n354), .Y(n459) );
  MUX21X1_HVT U321 ( .A1(n420), .A2(n343), .S0(n355), .Y(n429) );
  MUX21X1_HVT U322 ( .A1(n263), .A2(n336), .S0(n257), .Y(n424) );
  MUX21X1_HVT U323 ( .A1(n417), .A2(n335), .S0(n357), .Y(n433) );
  MUX21X1_HVT U324 ( .A1(n244), .A2(n310), .S0(n356), .Y(n598) );
  MUX21X1_HVT U325 ( .A1(n414), .A2(n315), .S0(n328), .Y(n506) );
  MUX21X1_HVT U326 ( .A1(n375), .A2(n342), .S0(n332), .Y(n537) );
  MUX21X1_HVT U327 ( .A1(n595), .A2(n314), .S0(n329), .Y(n503) );
  MUX21X1_HVT U328 ( .A1(n345), .A2(n350), .S0(n354), .Y(n423) );
  XNOR2X1_HVT U329 ( .A1(n299), .A2(n253), .Y(n315) );
  MUX21X1_HVT U330 ( .A1(n334), .A2(n350), .S0(n257), .Y(n525) );
  XOR2X1_HVT U331 ( .A1(n341), .A2(n355), .Y(n582) );
  MUX21X1_HVT U332 ( .A1(n343), .A2(n418), .S0(n354), .Y(n594) );
  MUX21X1_HVT U333 ( .A1(n334), .A2(n343), .S0(n355), .Y(n588) );
  MUX21X1_HVT U334 ( .A1(n333), .A2(n349), .S0(n253), .Y(n431) );
  MUX21X1_HVT U335 ( .A1(n347), .A2(n349), .S0(n356), .Y(n610) );
  XOR2X1_HVT U336 ( .A1(n347), .A2(n357), .Y(n581) );
  MUX21X1_HVT U337 ( .A1(n348), .A2(n244), .S0(n254), .Y(n609) );
  MUX21X1_HVT U338 ( .A1(n244), .A2(n335), .S0(n257), .Y(n583) );
  AND2X1_HVT U339 ( .A1(n623), .A2(n349), .Y(n316) );
  MUX21X1_HVT U340 ( .A1(n346), .A2(n335), .S0(n357), .Y(n509) );
  MUX21X1_HVT U341 ( .A1(n333), .A2(n348), .S0(n257), .Y(n426) );
  AND2X1_HVT U342 ( .A1(n353), .A2(n336), .Y(n317) );
  NBUFFX2_HVT U343 ( .A(n362), .Y(n331) );
  NBUFFX2_HVT U344 ( .A(n306), .Y(n334) );
  NBUFFX2_HVT U345 ( .A(n612), .Y(n341) );
  MUX21X1_HVT U346 ( .A1(n446), .A2(n406), .S0(n330), .Y(n445) );
  NBUFFX2_HVT U347 ( .A(n306), .Y(n335) );
  NBUFFX2_HVT U348 ( .A(n612), .Y(n343) );
  MUX21X1_HVT U349 ( .A1(n389), .A2(n380), .S0(n332), .Y(n577) );
  MUX21X1_HVT U350 ( .A1(n310), .A2(n421), .S0(n354), .Y(n578) );
  MUX21X1_HVT U351 ( .A1(n299), .A2(n345), .S0(n356), .Y(n488) );
  NBUFFX2_HVT U352 ( .A(n629), .Y(n352) );
  NBUFFX2_HVT U353 ( .A(n612), .Y(n342) );
  MUX21X1_HVT U354 ( .A1(n387), .A2(n625), .S0(n329), .Y(n572) );
  NBUFFX2_HVT U355 ( .A(n624), .Y(n344) );
  AND2X1_HVT U356 ( .A1(n347), .A2(n242), .Y(n318) );
  AND2X1_HVT U357 ( .A1(n421), .A2(n258), .Y(n319) );
  MUX21X1_HVT U358 ( .A1(n373), .A2(n587), .S0(n332), .Y(n520) );
  XOR2X1_HVT U359 ( .A1(n629), .A2(n257), .Y(n591) );
  NBUFFX2_HVT U360 ( .A(n624), .Y(n345) );
  NBUFFX2_HVT U361 ( .A(n627), .Y(n346) );
  NBUFFX2_HVT U362 ( .A(n627), .Y(n348) );
  NBUFFX2_HVT U363 ( .A(n627), .Y(n347) );
  NBUFFX2_HVT U364 ( .A(in[2]), .Y(n327) );
  NBUFFX2_HVT U365 ( .A(n359), .Y(n329) );
  NBUFFX2_HVT U366 ( .A(n323), .Y(n328) );
  XNOR2X1_HVT U367 ( .A1(n283), .A2(n325), .Y(n320) );
  NBUFFX2_HVT U368 ( .A(n359), .Y(n325) );
  NBUFFX2_HVT U369 ( .A(n359), .Y(n326) );
  NBUFFX2_HVT U370 ( .A(n359), .Y(n324) );
  NBUFFX2_HVT U371 ( .A(n359), .Y(n322) );
  NBUFFX2_HVT U372 ( .A(n359), .Y(n323) );
  MUX21X1_HVT U373 ( .A1(n420), .A2(n297), .S0(n355), .Y(n422) );
  MUX21X1_HVT U374 ( .A1(n352), .A2(n297), .S0(n254), .Y(n473) );
  MUX21X1_HVT U375 ( .A1(n498), .A2(n499), .S0(n338), .Y(n497) );
  MUX21X1_HVT U376 ( .A1(n494), .A2(n495), .S0(n291), .Y(n493) );
  MUX21X1_HVT U377 ( .A1(n198), .A2(n420), .S0(n357), .Y(n604) );
  XOR2X1_HVT U378 ( .A1(n357), .A2(n307), .Y(n579) );
  MUX21X1_HVT U379 ( .A1(n310), .A2(n198), .S0(n253), .Y(n496) );
  MUX21X1_HVT U380 ( .A1(n421), .A2(n418), .S0(n355), .Y(n514) );
  MUX21X1_HVT U381 ( .A1(n344), .A2(n307), .S0(n356), .Y(n599) );
  MUX21X1_HVT U382 ( .A1(n307), .A2(n421), .S0(n257), .Y(n587) );
  MUX21X1_HVT U383 ( .A1(n307), .A2(n321), .S0(n356), .Y(n611) );
  MUX21X1_HVT U384 ( .A1(n297), .A2(n345), .S0(n356), .Y(n427) );
  MUX21X1_HVT U385 ( .A1(n297), .A2(n351), .S0(n355), .Y(n428) );
  MUX21X1_HVT U386 ( .A1(n336), .A2(n297), .S0(n254), .Y(n601) );
  MUX21X1_HVT U387 ( .A1(n333), .A2(n307), .S0(n353), .Y(n425) );
  MUX21X1_HVT U388 ( .A1(n198), .A2(n348), .S0(n353), .Y(n434) );
  MUX21X1_HVT U389 ( .A1(n348), .A2(n307), .S0(n353), .Y(n430) );
  NBUFFX2_HVT U390 ( .A(in[2]), .Y(n359) );
  NAND2X0_HVT U391 ( .A1(in[3]), .A2(n335), .Y(n321) );
  INVX0_HVT U392 ( .A(n617), .Y(n364) );
  INVX0_HVT U393 ( .A(n596), .Y(n365) );
  INVX0_HVT U394 ( .A(n590), .Y(n366) );
  INVX0_HVT U395 ( .A(n530), .Y(n367) );
  INVX0_HVT U396 ( .A(n491), .Y(n368) );
  INVX0_HVT U397 ( .A(n625), .Y(n370) );
  INVX0_HVT U398 ( .A(n622), .Y(n373) );
  INVX0_HVT U399 ( .A(n593), .Y(n375) );
  INVX0_HVT U400 ( .A(n615), .Y(n376) );
  INVX0_HVT U401 ( .A(n616), .Y(n378) );
  INVX0_HVT U402 ( .A(n614), .Y(n379) );
  INVX0_HVT U403 ( .A(n613), .Y(n380) );
  INVX0_HVT U404 ( .A(n611), .Y(n381) );
  INVX0_HVT U405 ( .A(n610), .Y(n382) );
  INVX0_HVT U406 ( .A(n609), .Y(n383) );
  INVX0_HVT U407 ( .A(n608), .Y(n384) );
  INVX0_HVT U408 ( .A(n604), .Y(n386) );
  INVX0_HVT U409 ( .A(n602), .Y(n388) );
  INVX0_HVT U410 ( .A(n601), .Y(n389) );
  INVX0_HVT U411 ( .A(n598), .Y(n392) );
  INVX0_HVT U412 ( .A(n597), .Y(n393) );
  INVX0_HVT U413 ( .A(n591), .Y(n396) );
  INVX0_HVT U414 ( .A(n589), .Y(n397) );
  INVX0_HVT U415 ( .A(n588), .Y(n398) );
  INVX0_HVT U416 ( .A(n583), .Y(n400) );
  INVX0_HVT U417 ( .A(n582), .Y(n401) );
  INVX0_HVT U418 ( .A(n619), .Y(n402) );
  INVX0_HVT U419 ( .A(n434), .Y(n403) );
  INVX0_HVT U420 ( .A(n431), .Y(n406) );
  INVX0_HVT U421 ( .A(n430), .Y(n407) );
  INVX0_HVT U422 ( .A(n429), .Y(n408) );
  INVX0_HVT U423 ( .A(n428), .Y(n409) );
  INVX0_HVT U424 ( .A(n427), .Y(n410) );
  INVX0_HVT U425 ( .A(n426), .Y(n411) );
  INVX0_HVT U426 ( .A(n425), .Y(n412) );
  INVX0_HVT U427 ( .A(n473), .Y(n413) );
  INVX0_HVT U428 ( .A(n424), .Y(n414) );
  INVX0_HVT U429 ( .A(n423), .Y(n415) );
endmodule

