
module RAM_memory ( data, addr, we, clk, rst, q );
  input [255:0] data;
  input [3:0] addr;
  output [255:0] q;
  input we, clk, rst;
  wire   N26, N27, N28, N29, \ram[15][255] , \ram[15][254] , \ram[15][253] ,
         \ram[15][252] , \ram[15][251] , \ram[15][250] , \ram[15][249] ,
         \ram[15][248] , \ram[15][247] , \ram[15][246] , \ram[15][245] ,
         \ram[15][244] , \ram[15][243] , \ram[15][242] , \ram[15][241] ,
         \ram[15][240] , \ram[15][239] , \ram[15][238] , \ram[15][237] ,
         \ram[15][236] , \ram[15][235] , \ram[15][234] , \ram[15][233] ,
         \ram[15][232] , \ram[15][231] , \ram[15][230] , \ram[15][229] ,
         \ram[15][228] , \ram[15][227] , \ram[15][226] , \ram[15][225] ,
         \ram[15][224] , \ram[15][223] , \ram[15][222] , \ram[15][221] ,
         \ram[15][220] , \ram[15][219] , \ram[15][218] , \ram[15][217] ,
         \ram[15][216] , \ram[15][215] , \ram[15][214] , \ram[15][213] ,
         \ram[15][212] , \ram[15][211] , \ram[15][210] , \ram[15][209] ,
         \ram[15][208] , \ram[15][207] , \ram[15][206] , \ram[15][205] ,
         \ram[15][204] , \ram[15][203] , \ram[15][202] , \ram[15][201] ,
         \ram[15][200] , \ram[15][199] , \ram[15][198] , \ram[15][197] ,
         \ram[15][196] , \ram[15][195] , \ram[15][194] , \ram[15][193] ,
         \ram[15][192] , \ram[15][191] , \ram[15][190] , \ram[15][189] ,
         \ram[15][188] , \ram[15][187] , \ram[15][186] , \ram[15][185] ,
         \ram[15][184] , \ram[15][183] , \ram[15][182] , \ram[15][181] ,
         \ram[15][180] , \ram[15][179] , \ram[15][178] , \ram[15][177] ,
         \ram[15][176] , \ram[15][175] , \ram[15][174] , \ram[15][173] ,
         \ram[15][172] , \ram[15][171] , \ram[15][170] , \ram[15][169] ,
         \ram[15][168] , \ram[15][167] , \ram[15][166] , \ram[15][165] ,
         \ram[15][164] , \ram[15][163] , \ram[15][162] , \ram[15][161] ,
         \ram[15][160] , \ram[15][159] , \ram[15][158] , \ram[15][157] ,
         \ram[15][156] , \ram[15][155] , \ram[15][154] , \ram[15][153] ,
         \ram[15][152] , \ram[15][151] , \ram[15][150] , \ram[15][149] ,
         \ram[15][148] , \ram[15][147] , \ram[15][146] , \ram[15][145] ,
         \ram[15][144] , \ram[15][143] , \ram[15][142] , \ram[15][141] ,
         \ram[15][140] , \ram[15][139] , \ram[15][138] , \ram[15][137] ,
         \ram[15][136] , \ram[15][135] , \ram[15][134] , \ram[15][133] ,
         \ram[15][132] , \ram[15][131] , \ram[15][130] , \ram[15][129] ,
         \ram[15][128] , \ram[15][127] , \ram[15][126] , \ram[15][125] ,
         \ram[15][124] , \ram[15][123] , \ram[15][122] , \ram[15][121] ,
         \ram[15][120] , \ram[15][119] , \ram[15][118] , \ram[15][117] ,
         \ram[15][116] , \ram[15][115] , \ram[15][114] , \ram[15][113] ,
         \ram[15][112] , \ram[15][111] , \ram[15][110] , \ram[15][109] ,
         \ram[15][108] , \ram[15][107] , \ram[15][106] , \ram[15][105] ,
         \ram[15][104] , \ram[15][102] , \ram[15][101] , \ram[15][100] ,
         \ram[15][99] , \ram[15][98] , \ram[15][97] , \ram[15][96] ,
         \ram[15][95] , \ram[15][94] , \ram[15][93] , \ram[15][92] ,
         \ram[15][91] , \ram[15][90] , \ram[15][89] , \ram[15][88] ,
         \ram[15][87] , \ram[15][86] , \ram[15][85] , \ram[15][84] ,
         \ram[15][83] , \ram[15][82] , \ram[15][81] , \ram[15][80] ,
         \ram[15][79] , \ram[15][78] , \ram[15][77] , \ram[15][76] ,
         \ram[15][75] , \ram[15][74] , \ram[15][73] , \ram[15][72] ,
         \ram[15][71] , \ram[15][70] , \ram[15][69] , \ram[15][68] ,
         \ram[15][67] , \ram[15][66] , \ram[15][65] , \ram[15][64] ,
         \ram[15][63] , \ram[15][62] , \ram[15][61] , \ram[15][60] ,
         \ram[15][59] , \ram[15][58] , \ram[15][57] , \ram[15][56] ,
         \ram[15][55] , \ram[15][54] , \ram[15][53] , \ram[15][52] ,
         \ram[15][51] , \ram[15][50] , \ram[15][49] , \ram[15][48] ,
         \ram[15][47] , \ram[15][46] , \ram[15][45] , \ram[15][44] ,
         \ram[15][43] , \ram[15][42] , \ram[15][41] , \ram[15][40] ,
         \ram[15][39] , \ram[15][38] , \ram[15][37] , \ram[15][36] ,
         \ram[15][35] , \ram[15][34] , \ram[15][33] , \ram[15][32] ,
         \ram[15][31] , \ram[15][30] , \ram[15][29] , \ram[15][28] ,
         \ram[15][27] , \ram[15][26] , \ram[15][25] , \ram[15][24] ,
         \ram[15][23] , \ram[15][22] , \ram[15][21] , \ram[15][20] ,
         \ram[15][19] , \ram[15][18] , \ram[15][17] , \ram[15][16] ,
         \ram[15][15] , \ram[15][14] , \ram[15][13] , \ram[15][12] ,
         \ram[15][11] , \ram[15][10] , \ram[15][9] , \ram[15][8] ,
         \ram[15][7] , \ram[15][6] , \ram[15][5] , \ram[15][4] , \ram[15][3] ,
         \ram[15][2] , \ram[15][1] , \ram[15][0] , \ram[14][255] ,
         \ram[14][254] , \ram[14][253] , \ram[14][252] , \ram[14][251] ,
         \ram[14][250] , \ram[14][249] , \ram[14][248] , \ram[14][247] ,
         \ram[14][246] , \ram[14][245] , \ram[14][244] , \ram[14][243] ,
         \ram[14][242] , \ram[14][241] , \ram[14][240] , \ram[14][239] ,
         \ram[14][238] , \ram[14][237] , \ram[14][236] , \ram[14][235] ,
         \ram[14][234] , \ram[14][233] , \ram[14][232] , \ram[14][231] ,
         \ram[14][230] , \ram[14][229] , \ram[14][228] , \ram[14][227] ,
         \ram[14][226] , \ram[14][225] , \ram[14][224] , \ram[14][223] ,
         \ram[14][222] , \ram[14][221] , \ram[14][220] , \ram[14][219] ,
         \ram[14][218] , \ram[14][217] , \ram[14][216] , \ram[14][215] ,
         \ram[14][214] , \ram[14][213] , \ram[14][212] , \ram[14][211] ,
         \ram[14][210] , \ram[14][209] , \ram[14][208] , \ram[14][207] ,
         \ram[14][206] , \ram[14][205] , \ram[14][204] , \ram[14][203] ,
         \ram[14][202] , \ram[14][201] , \ram[14][200] , \ram[14][199] ,
         \ram[14][198] , \ram[14][197] , \ram[14][196] , \ram[14][195] ,
         \ram[14][194] , \ram[14][193] , \ram[14][192] , \ram[14][191] ,
         \ram[14][190] , \ram[14][189] , \ram[14][188] , \ram[14][187] ,
         \ram[14][186] , \ram[14][185] , \ram[14][184] , \ram[14][183] ,
         \ram[14][182] , \ram[14][181] , \ram[14][180] , \ram[14][179] ,
         \ram[14][178] , \ram[14][177] , \ram[14][176] , \ram[14][175] ,
         \ram[14][174] , \ram[14][173] , \ram[14][172] , \ram[14][171] ,
         \ram[14][170] , \ram[14][169] , \ram[14][168] , \ram[14][167] ,
         \ram[14][166] , \ram[14][165] , \ram[14][164] , \ram[14][163] ,
         \ram[14][162] , \ram[14][161] , \ram[14][160] , \ram[14][159] ,
         \ram[14][158] , \ram[14][157] , \ram[14][156] , \ram[14][155] ,
         \ram[14][154] , \ram[14][153] , \ram[14][152] , \ram[14][151] ,
         \ram[14][150] , \ram[14][149] , \ram[14][148] , \ram[14][147] ,
         \ram[14][146] , \ram[14][145] , \ram[14][144] , \ram[14][143] ,
         \ram[14][142] , \ram[14][141] , \ram[14][140] , \ram[14][139] ,
         \ram[14][138] , \ram[14][137] , \ram[14][136] , \ram[14][135] ,
         \ram[14][134] , \ram[14][133] , \ram[14][132] , \ram[14][131] ,
         \ram[14][130] , \ram[14][129] , \ram[14][128] , \ram[14][127] ,
         \ram[14][126] , \ram[14][125] , \ram[14][124] , \ram[14][123] ,
         \ram[14][122] , \ram[14][121] , \ram[14][120] , \ram[14][119] ,
         \ram[14][118] , \ram[14][117] , \ram[14][116] , \ram[14][115] ,
         \ram[14][114] , \ram[14][113] , \ram[14][112] , \ram[14][111] ,
         \ram[14][110] , \ram[14][109] , \ram[14][108] , \ram[14][107] ,
         \ram[14][106] , \ram[14][105] , \ram[14][104] , \ram[14][103] ,
         \ram[14][102] , \ram[14][101] , \ram[14][100] , \ram[14][99] ,
         \ram[14][98] , \ram[14][97] , \ram[14][96] , \ram[14][95] ,
         \ram[14][94] , \ram[14][93] , \ram[14][92] , \ram[14][91] ,
         \ram[14][90] , \ram[14][89] , \ram[14][88] , \ram[14][87] ,
         \ram[14][86] , \ram[14][85] , \ram[14][84] , \ram[14][83] ,
         \ram[14][82] , \ram[14][81] , \ram[14][80] , \ram[14][79] ,
         \ram[14][78] , \ram[14][77] , \ram[14][76] , \ram[14][75] ,
         \ram[14][74] , \ram[14][73] , \ram[14][72] , \ram[14][71] ,
         \ram[14][70] , \ram[14][69] , \ram[14][68] , \ram[14][67] ,
         \ram[14][66] , \ram[14][65] , \ram[14][64] , \ram[14][63] ,
         \ram[14][62] , \ram[14][61] , \ram[14][60] , \ram[14][59] ,
         \ram[14][58] , \ram[14][57] , \ram[14][56] , \ram[14][55] ,
         \ram[14][54] , \ram[14][53] , \ram[14][52] , \ram[14][51] ,
         \ram[14][50] , \ram[14][49] , \ram[14][48] , \ram[14][47] ,
         \ram[14][46] , \ram[14][45] , \ram[14][44] , \ram[14][43] ,
         \ram[14][42] , \ram[14][41] , \ram[14][40] , \ram[14][39] ,
         \ram[14][38] , \ram[14][37] , \ram[14][36] , \ram[14][35] ,
         \ram[14][34] , \ram[14][33] , \ram[14][32] , \ram[14][31] ,
         \ram[14][30] , \ram[14][29] , \ram[14][28] , \ram[14][27] ,
         \ram[14][26] , \ram[14][25] , \ram[14][24] , \ram[14][23] ,
         \ram[14][22] , \ram[14][21] , \ram[14][20] , \ram[14][19] ,
         \ram[14][18] , \ram[14][17] , \ram[14][16] , \ram[14][15] ,
         \ram[14][14] , \ram[14][13] , \ram[14][12] , \ram[14][11] ,
         \ram[14][10] , \ram[14][9] , \ram[14][8] , \ram[14][7] , \ram[14][6] ,
         \ram[14][5] , \ram[14][4] , \ram[14][3] , \ram[14][2] , \ram[14][1] ,
         \ram[14][0] , \ram[13][255] , \ram[13][254] , \ram[13][253] ,
         \ram[13][252] , \ram[13][251] , \ram[13][250] , \ram[13][249] ,
         \ram[13][248] , \ram[13][247] , \ram[13][246] , \ram[13][245] ,
         \ram[13][244] , \ram[13][243] , \ram[13][242] , \ram[13][241] ,
         \ram[13][240] , \ram[13][239] , \ram[13][238] , \ram[13][237] ,
         \ram[13][236] , \ram[13][235] , \ram[13][234] , \ram[13][233] ,
         \ram[13][232] , \ram[13][231] , \ram[13][230] , \ram[13][229] ,
         \ram[13][228] , \ram[13][227] , \ram[13][226] , \ram[13][225] ,
         \ram[13][224] , \ram[13][223] , \ram[13][222] , \ram[13][221] ,
         \ram[13][220] , \ram[13][219] , \ram[13][218] , \ram[13][217] ,
         \ram[13][216] , \ram[13][215] , \ram[13][214] , \ram[13][213] ,
         \ram[13][212] , \ram[13][211] , \ram[13][210] , \ram[13][209] ,
         \ram[13][208] , \ram[13][207] , \ram[13][206] , \ram[13][205] ,
         \ram[13][204] , \ram[13][203] , \ram[13][202] , \ram[13][201] ,
         \ram[13][200] , \ram[13][199] , \ram[13][198] , \ram[13][197] ,
         \ram[13][196] , \ram[13][195] , \ram[13][194] , \ram[13][193] ,
         \ram[13][192] , \ram[13][191] , \ram[13][190] , \ram[13][189] ,
         \ram[13][188] , \ram[13][187] , \ram[13][186] , \ram[13][185] ,
         \ram[13][184] , \ram[13][183] , \ram[13][182] , \ram[13][181] ,
         \ram[13][180] , \ram[13][179] , \ram[13][178] , \ram[13][177] ,
         \ram[13][176] , \ram[13][175] , \ram[13][174] , \ram[13][173] ,
         \ram[13][172] , \ram[13][171] , \ram[13][170] , \ram[13][169] ,
         \ram[13][168] , \ram[13][167] , \ram[13][166] , \ram[13][165] ,
         \ram[13][164] , \ram[13][163] , \ram[13][162] , \ram[13][161] ,
         \ram[13][160] , \ram[13][159] , \ram[13][158] , \ram[13][157] ,
         \ram[13][156] , \ram[13][155] , \ram[13][154] , \ram[13][153] ,
         \ram[13][152] , \ram[13][151] , \ram[13][150] , \ram[13][149] ,
         \ram[13][148] , \ram[13][147] , \ram[13][146] , \ram[13][145] ,
         \ram[13][144] , \ram[13][143] , \ram[13][142] , \ram[13][141] ,
         \ram[13][140] , \ram[13][139] , \ram[13][138] , \ram[13][137] ,
         \ram[13][136] , \ram[13][135] , \ram[13][134] , \ram[13][133] ,
         \ram[13][132] , \ram[13][131] , \ram[13][130] , \ram[13][129] ,
         \ram[13][128] , \ram[13][127] , \ram[13][126] , \ram[13][125] ,
         \ram[13][124] , \ram[13][123] , \ram[13][122] , \ram[13][121] ,
         \ram[13][120] , \ram[13][119] , \ram[13][118] , \ram[13][117] ,
         \ram[13][116] , \ram[13][115] , \ram[13][114] , \ram[13][113] ,
         \ram[13][112] , \ram[13][111] , \ram[13][110] , \ram[13][109] ,
         \ram[13][108] , \ram[13][107] , \ram[13][106] , \ram[13][105] ,
         \ram[13][104] , \ram[13][103] , \ram[13][102] , \ram[13][100] ,
         \ram[13][99] , \ram[13][98] , \ram[13][97] , \ram[13][96] ,
         \ram[13][95] , \ram[13][94] , \ram[13][93] , \ram[13][92] ,
         \ram[13][91] , \ram[13][90] , \ram[13][89] , \ram[13][88] ,
         \ram[13][87] , \ram[13][86] , \ram[13][85] , \ram[13][84] ,
         \ram[13][83] , \ram[13][82] , \ram[13][81] , \ram[13][80] ,
         \ram[13][79] , \ram[13][78] , \ram[13][77] , \ram[13][76] ,
         \ram[13][75] , \ram[13][74] , \ram[13][73] , \ram[13][72] ,
         \ram[13][71] , \ram[13][70] , \ram[13][69] , \ram[13][68] ,
         \ram[13][67] , \ram[13][66] , \ram[13][65] , \ram[13][64] ,
         \ram[13][63] , \ram[13][62] , \ram[13][61] , \ram[13][60] ,
         \ram[13][59] , \ram[13][58] , \ram[13][57] , \ram[13][56] ,
         \ram[13][55] , \ram[13][54] , \ram[13][53] , \ram[13][52] ,
         \ram[13][51] , \ram[13][50] , \ram[13][49] , \ram[13][48] ,
         \ram[13][47] , \ram[13][46] , \ram[13][45] , \ram[13][44] ,
         \ram[13][43] , \ram[13][42] , \ram[13][41] , \ram[13][40] ,
         \ram[13][39] , \ram[13][38] , \ram[13][37] , \ram[13][36] ,
         \ram[13][35] , \ram[13][34] , \ram[13][33] , \ram[13][32] ,
         \ram[13][31] , \ram[13][30] , \ram[13][29] , \ram[13][28] ,
         \ram[13][27] , \ram[13][26] , \ram[13][25] , \ram[13][24] ,
         \ram[13][23] , \ram[13][22] , \ram[13][21] , \ram[13][20] ,
         \ram[13][19] , \ram[13][18] , \ram[13][17] , \ram[13][16] ,
         \ram[13][15] , \ram[13][14] , \ram[13][13] , \ram[13][12] ,
         \ram[13][11] , \ram[13][10] , \ram[13][9] , \ram[13][8] ,
         \ram[13][7] , \ram[13][6] , \ram[13][5] , \ram[13][4] , \ram[13][3] ,
         \ram[13][2] , \ram[13][1] , \ram[13][0] , \ram[12][255] ,
         \ram[12][254] , \ram[12][253] , \ram[12][252] , \ram[12][251] ,
         \ram[12][250] , \ram[12][249] , \ram[12][248] , \ram[12][247] ,
         \ram[12][246] , \ram[12][245] , \ram[12][244] , \ram[12][243] ,
         \ram[12][242] , \ram[12][241] , \ram[12][240] , \ram[12][239] ,
         \ram[12][238] , \ram[12][237] , \ram[12][236] , \ram[12][235] ,
         \ram[12][234] , \ram[12][233] , \ram[12][232] , \ram[12][231] ,
         \ram[12][230] , \ram[12][229] , \ram[12][228] , \ram[12][227] ,
         \ram[12][226] , \ram[12][225] , \ram[12][224] , \ram[12][223] ,
         \ram[12][222] , \ram[12][221] , \ram[12][220] , \ram[12][219] ,
         \ram[12][218] , \ram[12][217] , \ram[12][216] , \ram[12][215] ,
         \ram[12][214] , \ram[12][213] , \ram[12][212] , \ram[12][211] ,
         \ram[12][210] , \ram[12][209] , \ram[12][208] , \ram[12][207] ,
         \ram[12][206] , \ram[12][205] , \ram[12][204] , \ram[12][203] ,
         \ram[12][202] , \ram[12][201] , \ram[12][200] , \ram[12][199] ,
         \ram[12][198] , \ram[12][197] , \ram[12][196] , \ram[12][195] ,
         \ram[12][194] , \ram[12][193] , \ram[12][192] , \ram[12][191] ,
         \ram[12][190] , \ram[12][189] , \ram[12][188] , \ram[12][187] ,
         \ram[12][186] , \ram[12][185] , \ram[12][184] , \ram[12][183] ,
         \ram[12][182] , \ram[12][181] , \ram[12][180] , \ram[12][179] ,
         \ram[12][178] , \ram[12][177] , \ram[12][176] , \ram[12][175] ,
         \ram[12][174] , \ram[12][173] , \ram[12][172] , \ram[12][171] ,
         \ram[12][170] , \ram[12][169] , \ram[12][168] , \ram[12][167] ,
         \ram[12][166] , \ram[12][165] , \ram[12][164] , \ram[12][163] ,
         \ram[12][162] , \ram[12][161] , \ram[12][160] , \ram[12][159] ,
         \ram[12][158] , \ram[12][157] , \ram[12][156] , \ram[12][155] ,
         \ram[12][154] , \ram[12][153] , \ram[12][152] , \ram[12][151] ,
         \ram[12][150] , \ram[12][149] , \ram[12][148] , \ram[12][147] ,
         \ram[12][146] , \ram[12][145] , \ram[12][144] , \ram[12][143] ,
         \ram[12][142] , \ram[12][141] , \ram[12][140] , \ram[12][139] ,
         \ram[12][138] , \ram[12][137] , \ram[12][136] , \ram[12][135] ,
         \ram[12][134] , \ram[12][133] , \ram[12][132] , \ram[12][131] ,
         \ram[12][130] , \ram[12][129] , \ram[12][128] , \ram[12][127] ,
         \ram[12][126] , \ram[12][125] , \ram[12][124] , \ram[12][123] ,
         \ram[12][122] , \ram[12][121] , \ram[12][120] , \ram[12][119] ,
         \ram[12][118] , \ram[12][117] , \ram[12][116] , \ram[12][115] ,
         \ram[12][114] , \ram[12][113] , \ram[12][112] , \ram[12][111] ,
         \ram[12][110] , \ram[12][109] , \ram[12][108] , \ram[12][107] ,
         \ram[12][106] , \ram[12][105] , \ram[12][104] , \ram[12][103] ,
         \ram[12][102] , \ram[12][101] , \ram[12][100] , \ram[12][99] ,
         \ram[12][98] , \ram[12][97] , \ram[12][96] , \ram[12][95] ,
         \ram[12][94] , \ram[12][93] , \ram[12][92] , \ram[12][91] ,
         \ram[12][90] , \ram[12][89] , \ram[12][88] , \ram[12][87] ,
         \ram[12][86] , \ram[12][85] , \ram[12][84] , \ram[12][83] ,
         \ram[12][82] , \ram[12][81] , \ram[12][80] , \ram[12][79] ,
         \ram[12][78] , \ram[12][77] , \ram[12][76] , \ram[12][75] ,
         \ram[12][74] , \ram[12][73] , \ram[12][72] , \ram[12][71] ,
         \ram[12][70] , \ram[12][69] , \ram[12][68] , \ram[12][67] ,
         \ram[12][66] , \ram[12][65] , \ram[12][64] , \ram[12][63] ,
         \ram[12][62] , \ram[12][61] , \ram[12][60] , \ram[12][59] ,
         \ram[12][58] , \ram[12][57] , \ram[12][56] , \ram[12][55] ,
         \ram[12][54] , \ram[12][53] , \ram[12][52] , \ram[12][51] ,
         \ram[12][50] , \ram[12][49] , \ram[12][48] , \ram[12][47] ,
         \ram[12][46] , \ram[12][45] , \ram[12][44] , \ram[12][43] ,
         \ram[12][42] , \ram[12][41] , \ram[12][40] , \ram[12][39] ,
         \ram[12][38] , \ram[12][37] , \ram[12][36] , \ram[12][35] ,
         \ram[12][34] , \ram[12][33] , \ram[12][32] , \ram[12][31] ,
         \ram[12][30] , \ram[12][29] , \ram[12][28] , \ram[12][27] ,
         \ram[12][26] , \ram[12][25] , \ram[12][24] , \ram[12][23] ,
         \ram[12][22] , \ram[12][21] , \ram[12][20] , \ram[12][19] ,
         \ram[12][18] , \ram[12][17] , \ram[12][16] , \ram[12][15] ,
         \ram[12][14] , \ram[12][13] , \ram[12][12] , \ram[12][11] ,
         \ram[12][10] , \ram[12][9] , \ram[12][8] , \ram[12][7] , \ram[12][6] ,
         \ram[12][5] , \ram[12][4] , \ram[12][3] , \ram[12][2] , \ram[12][1] ,
         \ram[12][0] , \ram[11][255] , \ram[11][254] , \ram[11][253] ,
         \ram[11][252] , \ram[11][251] , \ram[11][250] , \ram[11][249] ,
         \ram[11][248] , \ram[11][247] , \ram[11][246] , \ram[11][245] ,
         \ram[11][244] , \ram[11][243] , \ram[11][242] , \ram[11][241] ,
         \ram[11][240] , \ram[11][239] , \ram[11][238] , \ram[11][237] ,
         \ram[11][236] , \ram[11][235] , \ram[11][234] , \ram[11][233] ,
         \ram[11][232] , \ram[11][231] , \ram[11][230] , \ram[11][229] ,
         \ram[11][228] , \ram[11][227] , \ram[11][226] , \ram[11][225] ,
         \ram[11][224] , \ram[11][223] , \ram[11][222] , \ram[11][221] ,
         \ram[11][220] , \ram[11][219] , \ram[11][218] , \ram[11][217] ,
         \ram[11][216] , \ram[11][215] , \ram[11][214] , \ram[11][213] ,
         \ram[11][212] , \ram[11][211] , \ram[11][210] , \ram[11][209] ,
         \ram[11][208] , \ram[11][207] , \ram[11][206] , \ram[11][205] ,
         \ram[11][204] , \ram[11][203] , \ram[11][202] , \ram[11][201] ,
         \ram[11][200] , \ram[11][199] , \ram[11][198] , \ram[11][197] ,
         \ram[11][196] , \ram[11][195] , \ram[11][194] , \ram[11][193] ,
         \ram[11][192] , \ram[11][191] , \ram[11][190] , \ram[11][189] ,
         \ram[11][188] , \ram[11][187] , \ram[11][186] , \ram[11][185] ,
         \ram[11][184] , \ram[11][183] , \ram[11][182] , \ram[11][181] ,
         \ram[11][180] , \ram[11][179] , \ram[11][178] , \ram[11][177] ,
         \ram[11][176] , \ram[11][175] , \ram[11][174] , \ram[11][173] ,
         \ram[11][172] , \ram[11][171] , \ram[11][170] , \ram[11][169] ,
         \ram[11][168] , \ram[11][167] , \ram[11][166] , \ram[11][165] ,
         \ram[11][164] , \ram[11][163] , \ram[11][162] , \ram[11][161] ,
         \ram[11][160] , \ram[11][159] , \ram[11][158] , \ram[11][157] ,
         \ram[11][156] , \ram[11][155] , \ram[11][154] , \ram[11][153] ,
         \ram[11][152] , \ram[11][151] , \ram[11][150] , \ram[11][149] ,
         \ram[11][148] , \ram[11][147] , \ram[11][146] , \ram[11][145] ,
         \ram[11][144] , \ram[11][143] , \ram[11][142] , \ram[11][141] ,
         \ram[11][140] , \ram[11][139] , \ram[11][138] , \ram[11][137] ,
         \ram[11][136] , \ram[11][135] , \ram[11][134] , \ram[11][133] ,
         \ram[11][132] , \ram[11][131] , \ram[11][130] , \ram[11][129] ,
         \ram[11][128] , \ram[11][127] , \ram[11][126] , \ram[11][125] ,
         \ram[11][124] , \ram[11][123] , \ram[11][122] , \ram[11][121] ,
         \ram[11][120] , \ram[11][119] , \ram[11][118] , \ram[11][117] ,
         \ram[11][116] , \ram[11][115] , \ram[11][114] , \ram[11][113] ,
         \ram[11][112] , \ram[11][111] , \ram[11][110] , \ram[11][109] ,
         \ram[11][108] , \ram[11][107] , \ram[11][106] , \ram[11][105] ,
         \ram[11][104] , \ram[11][103] , \ram[11][102] , \ram[11][101] ,
         \ram[11][100] , \ram[11][99] , \ram[11][98] , \ram[11][97] ,
         \ram[11][96] , \ram[11][95] , \ram[11][94] , \ram[11][93] ,
         \ram[11][92] , \ram[11][91] , \ram[11][90] , \ram[11][89] ,
         \ram[11][88] , \ram[11][87] , \ram[11][86] , \ram[11][85] ,
         \ram[11][84] , \ram[11][83] , \ram[11][82] , \ram[11][81] ,
         \ram[11][80] , \ram[11][79] , \ram[11][78] , \ram[11][77] ,
         \ram[11][76] , \ram[11][75] , \ram[11][74] , \ram[11][73] ,
         \ram[11][72] , \ram[11][71] , \ram[11][70] , \ram[11][69] ,
         \ram[11][68] , \ram[11][67] , \ram[11][66] , \ram[11][65] ,
         \ram[11][64] , \ram[11][63] , \ram[11][62] , \ram[11][61] ,
         \ram[11][60] , \ram[11][59] , \ram[11][58] , \ram[11][57] ,
         \ram[11][56] , \ram[11][55] , \ram[11][54] , \ram[11][53] ,
         \ram[11][52] , \ram[11][51] , \ram[11][50] , \ram[11][49] ,
         \ram[11][48] , \ram[11][47] , \ram[11][46] , \ram[11][45] ,
         \ram[11][44] , \ram[11][43] , \ram[11][42] , \ram[11][41] ,
         \ram[11][40] , \ram[11][39] , \ram[11][38] , \ram[11][37] ,
         \ram[11][36] , \ram[11][35] , \ram[11][34] , \ram[11][33] ,
         \ram[11][32] , \ram[11][31] , \ram[11][30] , \ram[11][29] ,
         \ram[11][28] , \ram[11][27] , \ram[11][26] , \ram[11][25] ,
         \ram[11][24] , \ram[11][23] , \ram[11][22] , \ram[11][21] ,
         \ram[11][20] , \ram[11][19] , \ram[11][18] , \ram[11][17] ,
         \ram[11][16] , \ram[11][15] , \ram[11][14] , \ram[11][13] ,
         \ram[11][12] , \ram[11][11] , \ram[11][10] , \ram[11][9] ,
         \ram[11][8] , \ram[11][7] , \ram[11][6] , \ram[11][5] , \ram[11][4] ,
         \ram[11][3] , \ram[11][2] , \ram[11][1] , \ram[11][0] ,
         \ram[10][255] , \ram[10][254] , \ram[10][253] , \ram[10][252] ,
         \ram[10][251] , \ram[10][250] , \ram[10][249] , \ram[10][248] ,
         \ram[10][247] , \ram[10][246] , \ram[10][245] , \ram[10][244] ,
         \ram[10][243] , \ram[10][242] , \ram[10][241] , \ram[10][240] ,
         \ram[10][239] , \ram[10][238] , \ram[10][237] , \ram[10][236] ,
         \ram[10][235] , \ram[10][234] , \ram[10][233] , \ram[10][232] ,
         \ram[10][231] , \ram[10][230] , \ram[10][229] , \ram[10][228] ,
         \ram[10][227] , \ram[10][226] , \ram[10][225] , \ram[10][224] ,
         \ram[10][223] , \ram[10][222] , \ram[10][221] , \ram[10][220] ,
         \ram[10][219] , \ram[10][218] , \ram[10][217] , \ram[10][216] ,
         \ram[10][215] , \ram[10][214] , \ram[10][213] , \ram[10][212] ,
         \ram[10][211] , \ram[10][210] , \ram[10][209] , \ram[10][208] ,
         \ram[10][207] , \ram[10][206] , \ram[10][205] , \ram[10][204] ,
         \ram[10][203] , \ram[10][202] , \ram[10][201] , \ram[10][200] ,
         \ram[10][199] , \ram[10][198] , \ram[10][197] , \ram[10][196] ,
         \ram[10][195] , \ram[10][194] , \ram[10][193] , \ram[10][192] ,
         \ram[10][191] , \ram[10][190] , \ram[10][189] , \ram[10][188] ,
         \ram[10][187] , \ram[10][186] , \ram[10][185] , \ram[10][184] ,
         \ram[10][183] , \ram[10][182] , \ram[10][181] , \ram[10][180] ,
         \ram[10][179] , \ram[10][178] , \ram[10][177] , \ram[10][176] ,
         \ram[10][175] , \ram[10][174] , \ram[10][173] , \ram[10][172] ,
         \ram[10][171] , \ram[10][170] , \ram[10][169] , \ram[10][168] ,
         \ram[10][167] , \ram[10][166] , \ram[10][165] , \ram[10][164] ,
         \ram[10][163] , \ram[10][162] , \ram[10][161] , \ram[10][160] ,
         \ram[10][159] , \ram[10][158] , \ram[10][157] , \ram[10][156] ,
         \ram[10][155] , \ram[10][154] , \ram[10][153] , \ram[10][152] ,
         \ram[10][151] , \ram[10][150] , \ram[10][149] , \ram[10][148] ,
         \ram[10][147] , \ram[10][146] , \ram[10][145] , \ram[10][144] ,
         \ram[10][143] , \ram[10][142] , \ram[10][141] , \ram[10][140] ,
         \ram[10][139] , \ram[10][138] , \ram[10][137] , \ram[10][136] ,
         \ram[10][135] , \ram[10][134] , \ram[10][133] , \ram[10][132] ,
         \ram[10][131] , \ram[10][130] , \ram[10][129] , \ram[10][128] ,
         \ram[10][127] , \ram[10][126] , \ram[10][125] , \ram[10][124] ,
         \ram[10][123] , \ram[10][122] , \ram[10][121] , \ram[10][120] ,
         \ram[10][119] , \ram[10][118] , \ram[10][117] , \ram[10][116] ,
         \ram[10][115] , \ram[10][114] , \ram[10][113] , \ram[10][112] ,
         \ram[10][111] , \ram[10][110] , \ram[10][109] , \ram[10][108] ,
         \ram[10][107] , \ram[10][106] , \ram[10][105] , \ram[10][104] ,
         \ram[10][103] , \ram[10][102] , \ram[10][101] , \ram[10][100] ,
         \ram[10][99] , \ram[10][98] , \ram[10][97] , \ram[10][96] ,
         \ram[10][95] , \ram[10][94] , \ram[10][93] , \ram[10][92] ,
         \ram[10][91] , \ram[10][90] , \ram[10][89] , \ram[10][88] ,
         \ram[10][87] , \ram[10][86] , \ram[10][85] , \ram[10][84] ,
         \ram[10][83] , \ram[10][82] , \ram[10][81] , \ram[10][80] ,
         \ram[10][79] , \ram[10][78] , \ram[10][77] , \ram[10][76] ,
         \ram[10][75] , \ram[10][74] , \ram[10][73] , \ram[10][72] ,
         \ram[10][71] , \ram[10][70] , \ram[10][69] , \ram[10][68] ,
         \ram[10][67] , \ram[10][66] , \ram[10][65] , \ram[10][64] ,
         \ram[10][63] , \ram[10][62] , \ram[10][61] , \ram[10][60] ,
         \ram[10][59] , \ram[10][58] , \ram[10][57] , \ram[10][56] ,
         \ram[10][55] , \ram[10][54] , \ram[10][53] , \ram[10][52] ,
         \ram[10][51] , \ram[10][50] , \ram[10][49] , \ram[10][48] ,
         \ram[10][47] , \ram[10][46] , \ram[10][45] , \ram[10][44] ,
         \ram[10][43] , \ram[10][42] , \ram[10][41] , \ram[10][40] ,
         \ram[10][39] , \ram[10][38] , \ram[10][37] , \ram[10][36] ,
         \ram[10][35] , \ram[10][34] , \ram[10][33] , \ram[10][32] ,
         \ram[10][31] , \ram[10][30] , \ram[10][29] , \ram[10][28] ,
         \ram[10][27] , \ram[10][26] , \ram[10][25] , \ram[10][24] ,
         \ram[10][23] , \ram[10][22] , \ram[10][21] , \ram[10][20] ,
         \ram[10][19] , \ram[10][18] , \ram[10][17] , \ram[10][16] ,
         \ram[10][15] , \ram[10][14] , \ram[10][13] , \ram[10][12] ,
         \ram[10][11] , \ram[10][10] , \ram[10][9] , \ram[10][8] ,
         \ram[10][7] , \ram[10][6] , \ram[10][5] , \ram[10][4] , \ram[10][3] ,
         \ram[10][2] , \ram[10][1] , \ram[10][0] , \ram[9][255] ,
         \ram[9][254] , \ram[9][253] , \ram[9][252] , \ram[9][251] ,
         \ram[9][250] , \ram[9][249] , \ram[9][248] , \ram[9][247] ,
         \ram[9][246] , \ram[9][245] , \ram[9][244] , \ram[9][243] ,
         \ram[9][242] , \ram[9][241] , \ram[9][240] , \ram[9][239] ,
         \ram[9][238] , \ram[9][237] , \ram[9][236] , \ram[9][235] ,
         \ram[9][234] , \ram[9][233] , \ram[9][232] , \ram[9][231] ,
         \ram[9][230] , \ram[9][229] , \ram[9][228] , \ram[9][227] ,
         \ram[9][226] , \ram[9][225] , \ram[9][224] , \ram[9][223] ,
         \ram[9][222] , \ram[9][221] , \ram[9][220] , \ram[9][219] ,
         \ram[9][218] , \ram[9][217] , \ram[9][216] , \ram[9][215] ,
         \ram[9][214] , \ram[9][213] , \ram[9][212] , \ram[9][211] ,
         \ram[9][210] , \ram[9][209] , \ram[9][208] , \ram[9][207] ,
         \ram[9][206] , \ram[9][205] , \ram[9][204] , \ram[9][203] ,
         \ram[9][202] , \ram[9][201] , \ram[9][200] , \ram[9][199] ,
         \ram[9][198] , \ram[9][197] , \ram[9][196] , \ram[9][195] ,
         \ram[9][194] , \ram[9][193] , \ram[9][192] , \ram[9][191] ,
         \ram[9][190] , \ram[9][189] , \ram[9][188] , \ram[9][187] ,
         \ram[9][186] , \ram[9][185] , \ram[9][184] , \ram[9][183] ,
         \ram[9][182] , \ram[9][181] , \ram[9][180] , \ram[9][179] ,
         \ram[9][178] , \ram[9][177] , \ram[9][176] , \ram[9][175] ,
         \ram[9][174] , \ram[9][173] , \ram[9][172] , \ram[9][171] ,
         \ram[9][170] , \ram[9][169] , \ram[9][168] , \ram[9][167] ,
         \ram[9][166] , \ram[9][165] , \ram[9][164] , \ram[9][163] ,
         \ram[9][162] , \ram[9][161] , \ram[9][160] , \ram[9][159] ,
         \ram[9][158] , \ram[9][157] , \ram[9][156] , \ram[9][155] ,
         \ram[9][154] , \ram[9][153] , \ram[9][152] , \ram[9][151] ,
         \ram[9][150] , \ram[9][149] , \ram[9][148] , \ram[9][147] ,
         \ram[9][146] , \ram[9][145] , \ram[9][144] , \ram[9][143] ,
         \ram[9][142] , \ram[9][141] , \ram[9][140] , \ram[9][139] ,
         \ram[9][138] , \ram[9][137] , \ram[9][136] , \ram[9][135] ,
         \ram[9][134] , \ram[9][133] , \ram[9][132] , \ram[9][131] ,
         \ram[9][130] , \ram[9][129] , \ram[9][128] , \ram[9][127] ,
         \ram[9][126] , \ram[9][125] , \ram[9][124] , \ram[9][123] ,
         \ram[9][122] , \ram[9][121] , \ram[9][120] , \ram[9][119] ,
         \ram[9][118] , \ram[9][117] , \ram[9][116] , \ram[9][115] ,
         \ram[9][114] , \ram[9][113] , \ram[9][112] , \ram[9][111] ,
         \ram[9][110] , \ram[9][109] , \ram[9][108] , \ram[9][107] ,
         \ram[9][106] , \ram[9][105] , \ram[9][104] , \ram[9][103] ,
         \ram[9][102] , \ram[9][101] , \ram[9][100] , \ram[9][99] ,
         \ram[9][98] , \ram[9][97] , \ram[9][96] , \ram[9][95] , \ram[9][94] ,
         \ram[9][93] , \ram[9][92] , \ram[9][91] , \ram[9][90] , \ram[9][89] ,
         \ram[9][88] , \ram[9][87] , \ram[9][86] , \ram[9][85] , \ram[9][84] ,
         \ram[9][83] , \ram[9][82] , \ram[9][81] , \ram[9][80] , \ram[9][79] ,
         \ram[9][78] , \ram[9][77] , \ram[9][76] , \ram[9][75] , \ram[9][74] ,
         \ram[9][73] , \ram[9][72] , \ram[9][71] , \ram[9][70] , \ram[9][69] ,
         \ram[9][68] , \ram[9][67] , \ram[9][66] , \ram[9][65] , \ram[9][64] ,
         \ram[9][63] , \ram[9][62] , \ram[9][61] , \ram[9][60] , \ram[9][59] ,
         \ram[9][58] , \ram[9][57] , \ram[9][56] , \ram[9][55] , \ram[9][54] ,
         \ram[9][53] , \ram[9][52] , \ram[9][51] , \ram[9][50] , \ram[9][49] ,
         \ram[9][48] , \ram[9][47] , \ram[9][46] , \ram[9][45] , \ram[9][44] ,
         \ram[9][43] , \ram[9][42] , \ram[9][41] , \ram[9][40] , \ram[9][39] ,
         \ram[9][38] , \ram[9][37] , \ram[9][36] , \ram[9][35] , \ram[9][34] ,
         \ram[9][33] , \ram[9][32] , \ram[9][31] , \ram[9][30] , \ram[9][29] ,
         \ram[9][28] , \ram[9][27] , \ram[9][26] , \ram[9][25] , \ram[9][24] ,
         \ram[9][23] , \ram[9][22] , \ram[9][21] , \ram[9][20] , \ram[9][19] ,
         \ram[9][18] , \ram[9][17] , \ram[9][16] , \ram[9][15] , \ram[9][14] ,
         \ram[9][13] , \ram[9][12] , \ram[9][11] , \ram[9][10] , \ram[9][9] ,
         \ram[9][8] , \ram[9][7] , \ram[9][6] , \ram[9][5] , \ram[9][4] ,
         \ram[9][3] , \ram[9][2] , \ram[9][1] , \ram[9][0] , \ram[8][255] ,
         \ram[8][254] , \ram[8][253] , \ram[8][252] , \ram[8][251] ,
         \ram[8][250] , \ram[8][249] , \ram[8][248] , \ram[8][247] ,
         \ram[8][246] , \ram[8][245] , \ram[8][244] , \ram[8][243] ,
         \ram[8][242] , \ram[8][241] , \ram[8][240] , \ram[8][239] ,
         \ram[8][238] , \ram[8][237] , \ram[8][236] , \ram[8][235] ,
         \ram[8][234] , \ram[8][233] , \ram[8][232] , \ram[8][231] ,
         \ram[8][230] , \ram[8][229] , \ram[8][228] , \ram[8][227] ,
         \ram[8][226] , \ram[8][225] , \ram[8][224] , \ram[8][223] ,
         \ram[8][222] , \ram[8][221] , \ram[8][220] , \ram[8][219] ,
         \ram[8][218] , \ram[8][217] , \ram[8][216] , \ram[8][215] ,
         \ram[8][214] , \ram[8][213] , \ram[8][212] , \ram[8][211] ,
         \ram[8][210] , \ram[8][209] , \ram[8][208] , \ram[8][207] ,
         \ram[8][206] , \ram[8][205] , \ram[8][204] , \ram[8][203] ,
         \ram[8][202] , \ram[8][201] , \ram[8][200] , \ram[8][199] ,
         \ram[8][198] , \ram[8][197] , \ram[8][196] , \ram[8][195] ,
         \ram[8][194] , \ram[8][193] , \ram[8][192] , \ram[8][191] ,
         \ram[8][190] , \ram[8][189] , \ram[8][188] , \ram[8][187] ,
         \ram[8][186] , \ram[8][185] , \ram[8][184] , \ram[8][183] ,
         \ram[8][182] , \ram[8][181] , \ram[8][180] , \ram[8][179] ,
         \ram[8][178] , \ram[8][177] , \ram[8][176] , \ram[8][175] ,
         \ram[8][174] , \ram[8][173] , \ram[8][172] , \ram[8][171] ,
         \ram[8][170] , \ram[8][169] , \ram[8][168] , \ram[8][167] ,
         \ram[8][166] , \ram[8][165] , \ram[8][164] , \ram[8][163] ,
         \ram[8][162] , \ram[8][161] , \ram[8][160] , \ram[8][159] ,
         \ram[8][158] , \ram[8][157] , \ram[8][156] , \ram[8][155] ,
         \ram[8][154] , \ram[8][153] , \ram[8][152] , \ram[8][151] ,
         \ram[8][150] , \ram[8][149] , \ram[8][148] , \ram[8][147] ,
         \ram[8][146] , \ram[8][145] , \ram[8][144] , \ram[8][143] ,
         \ram[8][142] , \ram[8][141] , \ram[8][140] , \ram[8][139] ,
         \ram[8][138] , \ram[8][137] , \ram[8][136] , \ram[8][135] ,
         \ram[8][134] , \ram[8][133] , \ram[8][132] , \ram[8][131] ,
         \ram[8][130] , \ram[8][129] , \ram[8][128] , \ram[8][127] ,
         \ram[8][126] , \ram[8][125] , \ram[8][124] , \ram[8][123] ,
         \ram[8][122] , \ram[8][121] , \ram[8][120] , \ram[8][119] ,
         \ram[8][118] , \ram[8][117] , \ram[8][116] , \ram[8][115] ,
         \ram[8][114] , \ram[8][113] , \ram[8][112] , \ram[8][111] ,
         \ram[8][110] , \ram[8][109] , \ram[8][108] , \ram[8][107] ,
         \ram[8][106] , \ram[8][105] , \ram[8][104] , \ram[8][103] ,
         \ram[8][102] , \ram[8][101] , \ram[8][100] , \ram[8][99] ,
         \ram[8][98] , \ram[8][97] , \ram[8][96] , \ram[8][95] , \ram[8][94] ,
         \ram[8][93] , \ram[8][92] , \ram[8][91] , \ram[8][90] , \ram[8][89] ,
         \ram[8][88] , \ram[8][87] , \ram[8][86] , \ram[8][85] , \ram[8][84] ,
         \ram[8][83] , \ram[8][82] , \ram[8][81] , \ram[8][80] , \ram[8][79] ,
         \ram[8][78] , \ram[8][77] , \ram[8][76] , \ram[8][75] , \ram[8][74] ,
         \ram[8][73] , \ram[8][72] , \ram[8][71] , \ram[8][70] , \ram[8][69] ,
         \ram[8][68] , \ram[8][67] , \ram[8][66] , \ram[8][65] , \ram[8][64] ,
         \ram[8][63] , \ram[8][62] , \ram[8][61] , \ram[8][60] , \ram[8][59] ,
         \ram[8][57] , \ram[8][56] , \ram[8][55] , \ram[8][54] , \ram[8][53] ,
         \ram[8][52] , \ram[8][51] , \ram[8][50] , \ram[8][49] , \ram[8][48] ,
         \ram[8][47] , \ram[8][46] , \ram[8][45] , \ram[8][44] , \ram[8][43] ,
         \ram[8][42] , \ram[8][41] , \ram[8][40] , \ram[8][39] , \ram[8][38] ,
         \ram[8][37] , \ram[8][36] , \ram[8][35] , \ram[8][34] , \ram[8][33] ,
         \ram[8][32] , \ram[8][31] , \ram[8][30] , \ram[8][29] , \ram[8][28] ,
         \ram[8][27] , \ram[8][26] , \ram[8][25] , \ram[8][24] , \ram[8][23] ,
         \ram[8][22] , \ram[8][21] , \ram[8][20] , \ram[8][19] , \ram[8][18] ,
         \ram[8][17] , \ram[8][16] , \ram[8][15] , \ram[8][14] , \ram[8][13] ,
         \ram[8][12] , \ram[8][11] , \ram[8][10] , \ram[8][9] , \ram[8][8] ,
         \ram[8][7] , \ram[8][6] , \ram[8][5] , \ram[8][4] , \ram[8][3] ,
         \ram[8][2] , \ram[8][1] , \ram[8][0] , \ram[7][255] , \ram[7][254] ,
         \ram[7][253] , \ram[7][252] , \ram[7][251] , \ram[7][250] ,
         \ram[7][249] , \ram[7][248] , \ram[7][247] , \ram[7][246] ,
         \ram[7][245] , \ram[7][244] , \ram[7][243] , \ram[7][242] ,
         \ram[7][241] , \ram[7][240] , \ram[7][239] , \ram[7][238] ,
         \ram[7][237] , \ram[7][236] , \ram[7][235] , \ram[7][234] ,
         \ram[7][233] , \ram[7][232] , \ram[7][231] , \ram[7][230] ,
         \ram[7][229] , \ram[7][228] , \ram[7][227] , \ram[7][226] ,
         \ram[7][225] , \ram[7][224] , \ram[7][223] , \ram[7][222] ,
         \ram[7][221] , \ram[7][220] , \ram[7][219] , \ram[7][218] ,
         \ram[7][217] , \ram[7][216] , \ram[7][215] , \ram[7][214] ,
         \ram[7][213] , \ram[7][212] , \ram[7][211] , \ram[7][210] ,
         \ram[7][209] , \ram[7][208] , \ram[7][207] , \ram[7][206] ,
         \ram[7][205] , \ram[7][204] , \ram[7][203] , \ram[7][202] ,
         \ram[7][201] , \ram[7][200] , \ram[7][199] , \ram[7][198] ,
         \ram[7][197] , \ram[7][196] , \ram[7][195] , \ram[7][194] ,
         \ram[7][193] , \ram[7][192] , \ram[7][191] , \ram[7][190] ,
         \ram[7][189] , \ram[7][188] , \ram[7][187] , \ram[7][186] ,
         \ram[7][185] , \ram[7][184] , \ram[7][183] , \ram[7][182] ,
         \ram[7][181] , \ram[7][180] , \ram[7][179] , \ram[7][178] ,
         \ram[7][177] , \ram[7][176] , \ram[7][175] , \ram[7][174] ,
         \ram[7][173] , \ram[7][172] , \ram[7][171] , \ram[7][170] ,
         \ram[7][169] , \ram[7][168] , \ram[7][167] , \ram[7][166] ,
         \ram[7][165] , \ram[7][164] , \ram[7][163] , \ram[7][162] ,
         \ram[7][161] , \ram[7][160] , \ram[7][159] , \ram[7][158] ,
         \ram[7][157] , \ram[7][156] , \ram[7][155] , \ram[7][154] ,
         \ram[7][153] , \ram[7][152] , \ram[7][151] , \ram[7][150] ,
         \ram[7][149] , \ram[7][148] , \ram[7][147] , \ram[7][146] ,
         \ram[7][145] , \ram[7][144] , \ram[7][143] , \ram[7][142] ,
         \ram[7][141] , \ram[7][140] , \ram[7][139] , \ram[7][138] ,
         \ram[7][137] , \ram[7][136] , \ram[7][135] , \ram[7][134] ,
         \ram[7][133] , \ram[7][132] , \ram[7][131] , \ram[7][130] ,
         \ram[7][129] , \ram[7][128] , \ram[7][127] , \ram[7][126] ,
         \ram[7][125] , \ram[7][124] , \ram[7][123] , \ram[7][122] ,
         \ram[7][121] , \ram[7][120] , \ram[7][119] , \ram[7][118] ,
         \ram[7][117] , \ram[7][116] , \ram[7][115] , \ram[7][114] ,
         \ram[7][113] , \ram[7][112] , \ram[7][111] , \ram[7][110] ,
         \ram[7][109] , \ram[7][108] , \ram[7][107] , \ram[7][106] ,
         \ram[7][105] , \ram[7][104] , \ram[7][103] , \ram[7][102] ,
         \ram[7][101] , \ram[7][100] , \ram[7][99] , \ram[7][98] ,
         \ram[7][97] , \ram[7][96] , \ram[7][95] , \ram[7][94] , \ram[7][93] ,
         \ram[7][92] , \ram[7][91] , \ram[7][90] , \ram[7][89] , \ram[7][88] ,
         \ram[7][87] , \ram[7][86] , \ram[7][85] , \ram[7][84] , \ram[7][83] ,
         \ram[7][82] , \ram[7][81] , \ram[7][80] , \ram[7][79] , \ram[7][78] ,
         \ram[7][77] , \ram[7][76] , \ram[7][75] , \ram[7][74] , \ram[7][73] ,
         \ram[7][72] , \ram[7][71] , \ram[7][70] , \ram[7][69] , \ram[7][68] ,
         \ram[7][67] , \ram[7][66] , \ram[7][65] , \ram[7][64] , \ram[7][63] ,
         \ram[7][62] , \ram[7][61] , \ram[7][60] , \ram[7][59] , \ram[7][58] ,
         \ram[7][57] , \ram[7][56] , \ram[7][55] , \ram[7][54] , \ram[7][53] ,
         \ram[7][52] , \ram[7][51] , \ram[7][50] , \ram[7][49] , \ram[7][48] ,
         \ram[7][47] , \ram[7][46] , \ram[7][45] , \ram[7][44] , \ram[7][43] ,
         \ram[7][42] , \ram[7][41] , \ram[7][40] , \ram[7][39] , \ram[7][38] ,
         \ram[7][37] , \ram[7][36] , \ram[7][35] , \ram[7][34] , \ram[7][33] ,
         \ram[7][32] , \ram[7][31] , \ram[7][30] , \ram[7][29] , \ram[7][28] ,
         \ram[7][27] , \ram[7][26] , \ram[7][25] , \ram[7][24] , \ram[7][23] ,
         \ram[7][22] , \ram[7][21] , \ram[7][20] , \ram[7][19] , \ram[7][18] ,
         \ram[7][17] , \ram[7][16] , \ram[7][15] , \ram[7][14] , \ram[7][13] ,
         \ram[7][12] , \ram[7][11] , \ram[7][10] , \ram[7][9] , \ram[7][8] ,
         \ram[7][7] , \ram[7][6] , \ram[7][5] , \ram[7][4] , \ram[7][3] ,
         \ram[7][2] , \ram[7][1] , \ram[7][0] , \ram[6][255] , \ram[6][254] ,
         \ram[6][253] , \ram[6][252] , \ram[6][251] , \ram[6][250] ,
         \ram[6][249] , \ram[6][248] , \ram[6][247] , \ram[6][246] ,
         \ram[6][245] , \ram[6][244] , \ram[6][243] , \ram[6][242] ,
         \ram[6][241] , \ram[6][240] , \ram[6][239] , \ram[6][238] ,
         \ram[6][237] , \ram[6][236] , \ram[6][235] , \ram[6][234] ,
         \ram[6][233] , \ram[6][232] , \ram[6][231] , \ram[6][230] ,
         \ram[6][229] , \ram[6][228] , \ram[6][227] , \ram[6][226] ,
         \ram[6][225] , \ram[6][224] , \ram[6][223] , \ram[6][222] ,
         \ram[6][221] , \ram[6][220] , \ram[6][219] , \ram[6][218] ,
         \ram[6][217] , \ram[6][216] , \ram[6][215] , \ram[6][214] ,
         \ram[6][213] , \ram[6][212] , \ram[6][211] , \ram[6][210] ,
         \ram[6][209] , \ram[6][208] , \ram[6][207] , \ram[6][206] ,
         \ram[6][205] , \ram[6][204] , \ram[6][203] , \ram[6][202] ,
         \ram[6][201] , \ram[6][200] , \ram[6][199] , \ram[6][198] ,
         \ram[6][197] , \ram[6][196] , \ram[6][195] , \ram[6][194] ,
         \ram[6][193] , \ram[6][192] , \ram[6][191] , \ram[6][190] ,
         \ram[6][189] , \ram[6][188] , \ram[6][187] , \ram[6][186] ,
         \ram[6][185] , \ram[6][184] , \ram[6][183] , \ram[6][182] ,
         \ram[6][181] , \ram[6][180] , \ram[6][179] , \ram[6][178] ,
         \ram[6][177] , \ram[6][176] , \ram[6][175] , \ram[6][174] ,
         \ram[6][173] , \ram[6][172] , \ram[6][171] , \ram[6][170] ,
         \ram[6][169] , \ram[6][168] , \ram[6][167] , \ram[6][166] ,
         \ram[6][165] , \ram[6][164] , \ram[6][163] , \ram[6][162] ,
         \ram[6][161] , \ram[6][160] , \ram[6][159] , \ram[6][158] ,
         \ram[6][157] , \ram[6][156] , \ram[6][155] , \ram[6][154] ,
         \ram[6][153] , \ram[6][152] , \ram[6][151] , \ram[6][150] ,
         \ram[6][149] , \ram[6][148] , \ram[6][147] , \ram[6][146] ,
         \ram[6][145] , \ram[6][144] , \ram[6][143] , \ram[6][142] ,
         \ram[6][141] , \ram[6][140] , \ram[6][139] , \ram[6][138] ,
         \ram[6][137] , \ram[6][136] , \ram[6][135] , \ram[6][134] ,
         \ram[6][133] , \ram[6][132] , \ram[6][131] , \ram[6][130] ,
         \ram[6][129] , \ram[6][128] , \ram[6][127] , \ram[6][126] ,
         \ram[6][125] , \ram[6][124] , \ram[6][123] , \ram[6][122] ,
         \ram[6][121] , \ram[6][120] , \ram[6][119] , \ram[6][118] ,
         \ram[6][117] , \ram[6][116] , \ram[6][115] , \ram[6][114] ,
         \ram[6][113] , \ram[6][112] , \ram[6][111] , \ram[6][110] ,
         \ram[6][109] , \ram[6][108] , \ram[6][107] , \ram[6][106] ,
         \ram[6][105] , \ram[6][104] , \ram[6][103] , \ram[6][102] ,
         \ram[6][101] , \ram[6][100] , \ram[6][99] , \ram[6][98] ,
         \ram[6][97] , \ram[6][96] , \ram[6][95] , \ram[6][94] , \ram[6][93] ,
         \ram[6][92] , \ram[6][91] , \ram[6][90] , \ram[6][89] , \ram[6][88] ,
         \ram[6][87] , \ram[6][86] , \ram[6][85] , \ram[6][84] , \ram[6][83] ,
         \ram[6][82] , \ram[6][81] , \ram[6][80] , \ram[6][79] , \ram[6][78] ,
         \ram[6][77] , \ram[6][76] , \ram[6][75] , \ram[6][74] , \ram[6][73] ,
         \ram[6][72] , \ram[6][71] , \ram[6][70] , \ram[6][69] , \ram[6][68] ,
         \ram[6][67] , \ram[6][66] , \ram[6][65] , \ram[6][64] , \ram[6][63] ,
         \ram[6][62] , \ram[6][61] , \ram[6][60] , \ram[6][59] , \ram[6][58] ,
         \ram[6][57] , \ram[6][56] , \ram[6][55] , \ram[6][53] , \ram[6][52] ,
         \ram[6][51] , \ram[6][50] , \ram[6][49] , \ram[6][48] , \ram[6][47] ,
         \ram[6][46] , \ram[6][45] , \ram[6][44] , \ram[6][43] , \ram[6][42] ,
         \ram[6][41] , \ram[6][40] , \ram[6][39] , \ram[6][38] , \ram[6][37] ,
         \ram[6][36] , \ram[6][35] , \ram[6][34] , \ram[6][33] , \ram[6][32] ,
         \ram[6][31] , \ram[6][30] , \ram[6][29] , \ram[6][28] , \ram[6][27] ,
         \ram[6][26] , \ram[6][25] , \ram[6][24] , \ram[6][23] , \ram[6][22] ,
         \ram[6][21] , \ram[6][19] , \ram[6][18] , \ram[6][17] , \ram[6][16] ,
         \ram[6][15] , \ram[6][14] , \ram[6][13] , \ram[6][12] , \ram[6][11] ,
         \ram[6][10] , \ram[6][9] , \ram[6][8] , \ram[6][7] , \ram[6][6] ,
         \ram[6][5] , \ram[6][4] , \ram[6][3] , \ram[6][2] , \ram[6][1] ,
         \ram[6][0] , \ram[5][255] , \ram[5][254] , \ram[5][253] ,
         \ram[5][252] , \ram[5][251] , \ram[5][250] , \ram[5][249] ,
         \ram[5][248] , \ram[5][247] , \ram[5][246] , \ram[5][245] ,
         \ram[5][244] , \ram[5][243] , \ram[5][242] , \ram[5][241] ,
         \ram[5][240] , \ram[5][239] , \ram[5][238] , \ram[5][237] ,
         \ram[5][236] , \ram[5][235] , \ram[5][234] , \ram[5][233] ,
         \ram[5][232] , \ram[5][231] , \ram[5][230] , \ram[5][229] ,
         \ram[5][228] , \ram[5][227] , \ram[5][226] , \ram[5][225] ,
         \ram[5][224] , \ram[5][223] , \ram[5][222] , \ram[5][221] ,
         \ram[5][220] , \ram[5][219] , \ram[5][218] , \ram[5][217] ,
         \ram[5][216] , \ram[5][215] , \ram[5][214] , \ram[5][213] ,
         \ram[5][212] , \ram[5][211] , \ram[5][210] , \ram[5][209] ,
         \ram[5][208] , \ram[5][207] , \ram[5][206] , \ram[5][205] ,
         \ram[5][204] , \ram[5][203] , \ram[5][202] , \ram[5][201] ,
         \ram[5][200] , \ram[5][199] , \ram[5][198] , \ram[5][197] ,
         \ram[5][196] , \ram[5][195] , \ram[5][194] , \ram[5][193] ,
         \ram[5][192] , \ram[5][191] , \ram[5][190] , \ram[5][189] ,
         \ram[5][188] , \ram[5][187] , \ram[5][186] , \ram[5][185] ,
         \ram[5][184] , \ram[5][183] , \ram[5][182] , \ram[5][181] ,
         \ram[5][180] , \ram[5][179] , \ram[5][178] , \ram[5][177] ,
         \ram[5][176] , \ram[5][175] , \ram[5][174] , \ram[5][173] ,
         \ram[5][172] , \ram[5][171] , \ram[5][170] , \ram[5][169] ,
         \ram[5][168] , \ram[5][167] , \ram[5][166] , \ram[5][165] ,
         \ram[5][164] , \ram[5][163] , \ram[5][162] , \ram[5][161] ,
         \ram[5][160] , \ram[5][159] , \ram[5][158] , \ram[5][157] ,
         \ram[5][156] , \ram[5][155] , \ram[5][154] , \ram[5][153] ,
         \ram[5][152] , \ram[5][151] , \ram[5][150] , \ram[5][149] ,
         \ram[5][148] , \ram[5][147] , \ram[5][146] , \ram[5][145] ,
         \ram[5][144] , \ram[5][143] , \ram[5][142] , \ram[5][141] ,
         \ram[5][140] , \ram[5][139] , \ram[5][138] , \ram[5][137] ,
         \ram[5][136] , \ram[5][135] , \ram[5][134] , \ram[5][133] ,
         \ram[5][132] , \ram[5][131] , \ram[5][130] , \ram[5][129] ,
         \ram[5][128] , \ram[5][127] , \ram[5][126] , \ram[5][125] ,
         \ram[5][124] , \ram[5][123] , \ram[5][122] , \ram[5][121] ,
         \ram[5][120] , \ram[5][119] , \ram[5][118] , \ram[5][117] ,
         \ram[5][116] , \ram[5][115] , \ram[5][114] , \ram[5][113] ,
         \ram[5][112] , \ram[5][111] , \ram[5][110] , \ram[5][109] ,
         \ram[5][108] , \ram[5][107] , \ram[5][106] , \ram[5][105] ,
         \ram[5][104] , \ram[5][103] , \ram[5][102] , \ram[5][101] ,
         \ram[5][100] , \ram[5][99] , \ram[5][98] , \ram[5][97] , \ram[5][96] ,
         \ram[5][95] , \ram[5][94] , \ram[5][93] , \ram[5][92] , \ram[5][91] ,
         \ram[5][90] , \ram[5][89] , \ram[5][88] , \ram[5][87] , \ram[5][86] ,
         \ram[5][85] , \ram[5][84] , \ram[5][83] , \ram[5][82] , \ram[5][81] ,
         \ram[5][80] , \ram[5][79] , \ram[5][78] , \ram[5][77] , \ram[5][76] ,
         \ram[5][75] , \ram[5][74] , \ram[5][73] , \ram[5][72] , \ram[5][71] ,
         \ram[5][70] , \ram[5][69] , \ram[5][68] , \ram[5][67] , \ram[5][66] ,
         \ram[5][65] , \ram[5][64] , \ram[5][63] , \ram[5][62] , \ram[5][61] ,
         \ram[5][60] , \ram[5][59] , \ram[5][58] , \ram[5][57] , \ram[5][56] ,
         \ram[5][55] , \ram[5][54] , \ram[5][53] , \ram[5][52] , \ram[5][51] ,
         \ram[5][50] , \ram[5][49] , \ram[5][48] , \ram[5][47] , \ram[5][46] ,
         \ram[5][45] , \ram[5][44] , \ram[5][43] , \ram[5][42] , \ram[5][41] ,
         \ram[5][40] , \ram[5][39] , \ram[5][38] , \ram[5][37] , \ram[5][36] ,
         \ram[5][35] , \ram[5][34] , \ram[5][33] , \ram[5][32] , \ram[5][31] ,
         \ram[5][30] , \ram[5][29] , \ram[5][28] , \ram[5][27] , \ram[5][26] ,
         \ram[5][25] , \ram[5][24] , \ram[5][23] , \ram[5][22] , \ram[5][21] ,
         \ram[5][19] , \ram[5][18] , \ram[5][17] , \ram[5][16] , \ram[5][15] ,
         \ram[5][14] , \ram[5][13] , \ram[5][12] , \ram[5][11] , \ram[5][10] ,
         \ram[5][9] , \ram[5][8] , \ram[5][7] , \ram[5][6] , \ram[5][5] ,
         \ram[5][4] , \ram[5][3] , \ram[5][2] , \ram[5][1] , \ram[5][0] ,
         \ram[4][255] , \ram[4][254] , \ram[4][253] , \ram[4][252] ,
         \ram[4][251] , \ram[4][250] , \ram[4][249] , \ram[4][248] ,
         \ram[4][247] , \ram[4][246] , \ram[4][245] , \ram[4][244] ,
         \ram[4][243] , \ram[4][242] , \ram[4][241] , \ram[4][240] ,
         \ram[4][239] , \ram[4][238] , \ram[4][237] , \ram[4][236] ,
         \ram[4][235] , \ram[4][234] , \ram[4][233] , \ram[4][232] ,
         \ram[4][231] , \ram[4][230] , \ram[4][229] , \ram[4][228] ,
         \ram[4][227] , \ram[4][226] , \ram[4][225] , \ram[4][224] ,
         \ram[4][223] , \ram[4][222] , \ram[4][221] , \ram[4][220] ,
         \ram[4][219] , \ram[4][218] , \ram[4][217] , \ram[4][216] ,
         \ram[4][215] , \ram[4][214] , \ram[4][213] , \ram[4][212] ,
         \ram[4][211] , \ram[4][210] , \ram[4][209] , \ram[4][208] ,
         \ram[4][207] , \ram[4][206] , \ram[4][205] , \ram[4][204] ,
         \ram[4][203] , \ram[4][202] , \ram[4][201] , \ram[4][200] ,
         \ram[4][199] , \ram[4][198] , \ram[4][197] , \ram[4][196] ,
         \ram[4][195] , \ram[4][194] , \ram[4][193] , \ram[4][192] ,
         \ram[4][191] , \ram[4][190] , \ram[4][189] , \ram[4][188] ,
         \ram[4][187] , \ram[4][186] , \ram[4][185] , \ram[4][184] ,
         \ram[4][183] , \ram[4][182] , \ram[4][181] , \ram[4][180] ,
         \ram[4][179] , \ram[4][178] , \ram[4][177] , \ram[4][176] ,
         \ram[4][175] , \ram[4][174] , \ram[4][173] , \ram[4][172] ,
         \ram[4][171] , \ram[4][170] , \ram[4][169] , \ram[4][168] ,
         \ram[4][167] , \ram[4][166] , \ram[4][165] , \ram[4][164] ,
         \ram[4][163] , \ram[4][162] , \ram[4][161] , \ram[4][160] ,
         \ram[4][159] , \ram[4][158] , \ram[4][157] , \ram[4][156] ,
         \ram[4][155] , \ram[4][154] , \ram[4][153] , \ram[4][152] ,
         \ram[4][151] , \ram[4][150] , \ram[4][149] , \ram[4][148] ,
         \ram[4][147] , \ram[4][146] , \ram[4][145] , \ram[4][144] ,
         \ram[4][143] , \ram[4][142] , \ram[4][141] , \ram[4][140] ,
         \ram[4][139] , \ram[4][138] , \ram[4][137] , \ram[4][136] ,
         \ram[4][135] , \ram[4][134] , \ram[4][133] , \ram[4][132] ,
         \ram[4][131] , \ram[4][130] , \ram[4][129] , \ram[4][128] ,
         \ram[4][127] , \ram[4][126] , \ram[4][125] , \ram[4][124] ,
         \ram[4][123] , \ram[4][122] , \ram[4][121] , \ram[4][120] ,
         \ram[4][119] , \ram[4][118] , \ram[4][117] , \ram[4][116] ,
         \ram[4][115] , \ram[4][114] , \ram[4][113] , \ram[4][112] ,
         \ram[4][111] , \ram[4][110] , \ram[4][109] , \ram[4][108] ,
         \ram[4][107] , \ram[4][106] , \ram[4][105] , \ram[4][104] ,
         \ram[4][103] , \ram[4][102] , \ram[4][101] , \ram[4][100] ,
         \ram[4][99] , \ram[4][98] , \ram[4][97] , \ram[4][96] , \ram[4][95] ,
         \ram[4][94] , \ram[4][93] , \ram[4][92] , \ram[4][91] , \ram[4][90] ,
         \ram[4][89] , \ram[4][88] , \ram[4][87] , \ram[4][86] , \ram[4][85] ,
         \ram[4][84] , \ram[4][83] , \ram[4][82] , \ram[4][81] , \ram[4][80] ,
         \ram[4][79] , \ram[4][78] , \ram[4][77] , \ram[4][76] , \ram[4][75] ,
         \ram[4][74] , \ram[4][73] , \ram[4][72] , \ram[4][71] , \ram[4][70] ,
         \ram[4][69] , \ram[4][68] , \ram[4][67] , \ram[4][66] , \ram[4][65] ,
         \ram[4][64] , \ram[4][63] , \ram[4][62] , \ram[4][61] , \ram[4][60] ,
         \ram[4][59] , \ram[4][58] , \ram[4][57] , \ram[4][56] , \ram[4][55] ,
         \ram[4][54] , \ram[4][53] , \ram[4][52] , \ram[4][51] , \ram[4][50] ,
         \ram[4][49] , \ram[4][48] , \ram[4][47] , \ram[4][46] , \ram[4][45] ,
         \ram[4][44] , \ram[4][43] , \ram[4][42] , \ram[4][41] , \ram[4][40] ,
         \ram[4][39] , \ram[4][38] , \ram[4][37] , \ram[4][36] , \ram[4][35] ,
         \ram[4][34] , \ram[4][33] , \ram[4][32] , \ram[4][31] , \ram[4][30] ,
         \ram[4][29] , \ram[4][28] , \ram[4][27] , \ram[4][26] , \ram[4][25] ,
         \ram[4][24] , \ram[4][23] , \ram[4][22] , \ram[4][21] , \ram[4][19] ,
         \ram[4][18] , \ram[4][17] , \ram[4][16] , \ram[4][15] , \ram[4][14] ,
         \ram[4][13] , \ram[4][12] , \ram[4][11] , \ram[4][10] , \ram[4][9] ,
         \ram[4][8] , \ram[4][7] , \ram[4][6] , \ram[4][5] , \ram[4][4] ,
         \ram[4][3] , \ram[4][2] , \ram[4][1] , \ram[4][0] , \ram[3][255] ,
         \ram[3][254] , \ram[3][253] , \ram[3][252] , \ram[3][251] ,
         \ram[3][250] , \ram[3][249] , \ram[3][248] , \ram[3][247] ,
         \ram[3][246] , \ram[3][245] , \ram[3][244] , \ram[3][243] ,
         \ram[3][242] , \ram[3][241] , \ram[3][240] , \ram[3][239] ,
         \ram[3][238] , \ram[3][237] , \ram[3][236] , \ram[3][235] ,
         \ram[3][234] , \ram[3][233] , \ram[3][232] , \ram[3][231] ,
         \ram[3][230] , \ram[3][229] , \ram[3][228] , \ram[3][227] ,
         \ram[3][226] , \ram[3][225] , \ram[3][224] , \ram[3][223] ,
         \ram[3][222] , \ram[3][221] , \ram[3][220] , \ram[3][219] ,
         \ram[3][218] , \ram[3][217] , \ram[3][216] , \ram[3][215] ,
         \ram[3][214] , \ram[3][213] , \ram[3][212] , \ram[3][211] ,
         \ram[3][210] , \ram[3][209] , \ram[3][208] , \ram[3][207] ,
         \ram[3][206] , \ram[3][205] , \ram[3][204] , \ram[3][203] ,
         \ram[3][202] , \ram[3][201] , \ram[3][200] , \ram[3][199] ,
         \ram[3][198] , \ram[3][197] , \ram[3][196] , \ram[3][195] ,
         \ram[3][194] , \ram[3][193] , \ram[3][192] , \ram[3][191] ,
         \ram[3][190] , \ram[3][189] , \ram[3][188] , \ram[3][187] ,
         \ram[3][186] , \ram[3][185] , \ram[3][184] , \ram[3][183] ,
         \ram[3][182] , \ram[3][181] , \ram[3][180] , \ram[3][179] ,
         \ram[3][178] , \ram[3][177] , \ram[3][176] , \ram[3][175] ,
         \ram[3][174] , \ram[3][173] , \ram[3][172] , \ram[3][171] ,
         \ram[3][170] , \ram[3][169] , \ram[3][168] , \ram[3][167] ,
         \ram[3][166] , \ram[3][165] , \ram[3][164] , \ram[3][163] ,
         \ram[3][162] , \ram[3][161] , \ram[3][160] , \ram[3][159] ,
         \ram[3][158] , \ram[3][157] , \ram[3][156] , \ram[3][155] ,
         \ram[3][154] , \ram[3][153] , \ram[3][152] , \ram[3][151] ,
         \ram[3][150] , \ram[3][149] , \ram[3][148] , \ram[3][147] ,
         \ram[3][146] , \ram[3][145] , \ram[3][144] , \ram[3][143] ,
         \ram[3][142] , \ram[3][141] , \ram[3][140] , \ram[3][139] ,
         \ram[3][138] , \ram[3][137] , \ram[3][136] , \ram[3][135] ,
         \ram[3][134] , \ram[3][133] , \ram[3][132] , \ram[3][131] ,
         \ram[3][130] , \ram[3][129] , \ram[3][128] , \ram[3][127] ,
         \ram[3][126] , \ram[3][125] , \ram[3][124] , \ram[3][123] ,
         \ram[3][122] , \ram[3][121] , \ram[3][120] , \ram[3][119] ,
         \ram[3][118] , \ram[3][117] , \ram[3][116] , \ram[3][115] ,
         \ram[3][114] , \ram[3][113] , \ram[3][112] , \ram[3][111] ,
         \ram[3][110] , \ram[3][109] , \ram[3][108] , \ram[3][107] ,
         \ram[3][106] , \ram[3][105] , \ram[3][104] , \ram[3][103] ,
         \ram[3][102] , \ram[3][101] , \ram[3][100] , \ram[3][99] ,
         \ram[3][98] , \ram[3][97] , \ram[3][96] , \ram[3][95] , \ram[3][94] ,
         \ram[3][93] , \ram[3][92] , \ram[3][91] , \ram[3][90] , \ram[3][89] ,
         \ram[3][88] , \ram[3][87] , \ram[3][86] , \ram[3][85] , \ram[3][84] ,
         \ram[3][83] , \ram[3][82] , \ram[3][81] , \ram[3][80] , \ram[3][79] ,
         \ram[3][78] , \ram[3][77] , \ram[3][76] , \ram[3][75] , \ram[3][74] ,
         \ram[3][73] , \ram[3][72] , \ram[3][71] , \ram[3][70] , \ram[3][69] ,
         \ram[3][68] , \ram[3][67] , \ram[3][66] , \ram[3][65] , \ram[3][64] ,
         \ram[3][63] , \ram[3][62] , \ram[3][61] , \ram[3][60] , \ram[3][59] ,
         \ram[3][58] , \ram[3][57] , \ram[3][56] , \ram[3][55] , \ram[3][54] ,
         \ram[3][53] , \ram[3][52] , \ram[3][51] , \ram[3][50] , \ram[3][49] ,
         \ram[3][48] , \ram[3][47] , \ram[3][46] , \ram[3][45] , \ram[3][44] ,
         \ram[3][43] , \ram[3][42] , \ram[3][41] , \ram[3][40] , \ram[3][39] ,
         \ram[3][38] , \ram[3][37] , \ram[3][36] , \ram[3][35] , \ram[3][34] ,
         \ram[3][33] , \ram[3][32] , \ram[3][31] , \ram[3][30] , \ram[3][29] ,
         \ram[3][28] , \ram[3][27] , \ram[3][26] , \ram[3][25] , \ram[3][24] ,
         \ram[3][23] , \ram[3][22] , \ram[3][21] , \ram[3][20] , \ram[3][19] ,
         \ram[3][18] , \ram[3][17] , \ram[3][16] , \ram[3][15] , \ram[3][14] ,
         \ram[3][13] , \ram[3][12] , \ram[3][11] , \ram[3][10] , \ram[3][9] ,
         \ram[3][8] , \ram[3][7] , \ram[3][6] , \ram[3][5] , \ram[3][4] ,
         \ram[3][3] , \ram[3][2] , \ram[3][1] , \ram[3][0] , \ram[2][255] ,
         \ram[2][254] , \ram[2][253] , \ram[2][252] , \ram[2][251] ,
         \ram[2][250] , \ram[2][249] , \ram[2][248] , \ram[2][247] ,
         \ram[2][246] , \ram[2][245] , \ram[2][244] , \ram[2][243] ,
         \ram[2][242] , \ram[2][241] , \ram[2][240] , \ram[2][239] ,
         \ram[2][238] , \ram[2][237] , \ram[2][236] , \ram[2][235] ,
         \ram[2][234] , \ram[2][233] , \ram[2][232] , \ram[2][231] ,
         \ram[2][230] , \ram[2][229] , \ram[2][228] , \ram[2][227] ,
         \ram[2][226] , \ram[2][225] , \ram[2][224] , \ram[2][223] ,
         \ram[2][222] , \ram[2][221] , \ram[2][220] , \ram[2][219] ,
         \ram[2][218] , \ram[2][217] , \ram[2][216] , \ram[2][215] ,
         \ram[2][214] , \ram[2][213] , \ram[2][212] , \ram[2][211] ,
         \ram[2][210] , \ram[2][209] , \ram[2][208] , \ram[2][207] ,
         \ram[2][206] , \ram[2][205] , \ram[2][204] , \ram[2][203] ,
         \ram[2][202] , \ram[2][201] , \ram[2][200] , \ram[2][199] ,
         \ram[2][198] , \ram[2][197] , \ram[2][196] , \ram[2][195] ,
         \ram[2][194] , \ram[2][193] , \ram[2][192] , \ram[2][191] ,
         \ram[2][190] , \ram[2][189] , \ram[2][188] , \ram[2][187] ,
         \ram[2][186] , \ram[2][185] , \ram[2][184] , \ram[2][183] ,
         \ram[2][182] , \ram[2][181] , \ram[2][180] , \ram[2][179] ,
         \ram[2][178] , \ram[2][177] , \ram[2][176] , \ram[2][175] ,
         \ram[2][174] , \ram[2][173] , \ram[2][172] , \ram[2][171] ,
         \ram[2][170] , \ram[2][169] , \ram[2][168] , \ram[2][167] ,
         \ram[2][166] , \ram[2][165] , \ram[2][164] , \ram[2][163] ,
         \ram[2][162] , \ram[2][161] , \ram[2][160] , \ram[2][159] ,
         \ram[2][158] , \ram[2][157] , \ram[2][156] , \ram[2][155] ,
         \ram[2][154] , \ram[2][153] , \ram[2][152] , \ram[2][151] ,
         \ram[2][150] , \ram[2][149] , \ram[2][148] , \ram[2][147] ,
         \ram[2][146] , \ram[2][145] , \ram[2][144] , \ram[2][143] ,
         \ram[2][142] , \ram[2][141] , \ram[2][140] , \ram[2][139] ,
         \ram[2][138] , \ram[2][137] , \ram[2][136] , \ram[2][135] ,
         \ram[2][134] , \ram[2][133] , \ram[2][132] , \ram[2][131] ,
         \ram[2][130] , \ram[2][129] , \ram[2][128] , \ram[2][127] ,
         \ram[2][126] , \ram[2][125] , \ram[2][124] , \ram[2][123] ,
         \ram[2][122] , \ram[2][121] , \ram[2][120] , \ram[2][119] ,
         \ram[2][118] , \ram[2][117] , \ram[2][116] , \ram[2][115] ,
         \ram[2][114] , \ram[2][113] , \ram[2][112] , \ram[2][111] ,
         \ram[2][110] , \ram[2][109] , \ram[2][108] , \ram[2][107] ,
         \ram[2][106] , \ram[2][105] , \ram[2][104] , \ram[2][103] ,
         \ram[2][102] , \ram[2][101] , \ram[2][100] , \ram[2][99] ,
         \ram[2][98] , \ram[2][97] , \ram[2][96] , \ram[2][95] , \ram[2][94] ,
         \ram[2][93] , \ram[2][92] , \ram[2][91] , \ram[2][90] , \ram[2][89] ,
         \ram[2][88] , \ram[2][87] , \ram[2][86] , \ram[2][85] , \ram[2][84] ,
         \ram[2][83] , \ram[2][82] , \ram[2][81] , \ram[2][80] , \ram[2][79] ,
         \ram[2][78] , \ram[2][77] , \ram[2][76] , \ram[2][75] , \ram[2][74] ,
         \ram[2][73] , \ram[2][72] , \ram[2][71] , \ram[2][70] , \ram[2][69] ,
         \ram[2][68] , \ram[2][67] , \ram[2][66] , \ram[2][65] , \ram[2][64] ,
         \ram[2][63] , \ram[2][62] , \ram[2][61] , \ram[2][60] , \ram[2][59] ,
         \ram[2][58] , \ram[2][57] , \ram[2][56] , \ram[2][55] , \ram[2][54] ,
         \ram[2][53] , \ram[2][52] , \ram[2][51] , \ram[2][50] , \ram[2][49] ,
         \ram[2][48] , \ram[2][47] , \ram[2][46] , \ram[2][45] , \ram[2][44] ,
         \ram[2][43] , \ram[2][42] , \ram[2][41] , \ram[2][40] , \ram[2][39] ,
         \ram[2][38] , \ram[2][37] , \ram[2][36] , \ram[2][35] , \ram[2][34] ,
         \ram[2][33] , \ram[2][32] , \ram[2][31] , \ram[2][30] , \ram[2][29] ,
         \ram[2][28] , \ram[2][27] , \ram[2][26] , \ram[2][25] , \ram[2][24] ,
         \ram[2][23] , \ram[2][22] , \ram[2][21] , \ram[2][20] , \ram[2][19] ,
         \ram[2][18] , \ram[2][17] , \ram[2][16] , \ram[2][15] , \ram[2][14] ,
         \ram[2][13] , \ram[2][12] , \ram[2][11] , \ram[2][10] , \ram[2][9] ,
         \ram[2][8] , \ram[2][7] , \ram[2][6] , \ram[2][5] , \ram[2][4] ,
         \ram[2][3] , \ram[2][2] , \ram[2][1] , \ram[2][0] , \ram[1][255] ,
         \ram[1][254] , \ram[1][253] , \ram[1][252] , \ram[1][251] ,
         \ram[1][250] , \ram[1][249] , \ram[1][248] , \ram[1][247] ,
         \ram[1][246] , \ram[1][245] , \ram[1][244] , \ram[1][243] ,
         \ram[1][242] , \ram[1][241] , \ram[1][240] , \ram[1][239] ,
         \ram[1][238] , \ram[1][237] , \ram[1][236] , \ram[1][235] ,
         \ram[1][234] , \ram[1][233] , \ram[1][232] , \ram[1][231] ,
         \ram[1][230] , \ram[1][229] , \ram[1][228] , \ram[1][227] ,
         \ram[1][226] , \ram[1][225] , \ram[1][224] , \ram[1][223] ,
         \ram[1][222] , \ram[1][221] , \ram[1][220] , \ram[1][219] ,
         \ram[1][218] , \ram[1][217] , \ram[1][216] , \ram[1][215] ,
         \ram[1][214] , \ram[1][213] , \ram[1][212] , \ram[1][211] ,
         \ram[1][210] , \ram[1][209] , \ram[1][208] , \ram[1][207] ,
         \ram[1][206] , \ram[1][205] , \ram[1][204] , \ram[1][203] ,
         \ram[1][202] , \ram[1][201] , \ram[1][200] , \ram[1][199] ,
         \ram[1][198] , \ram[1][197] , \ram[1][196] , \ram[1][195] ,
         \ram[1][194] , \ram[1][193] , \ram[1][192] , \ram[1][191] ,
         \ram[1][190] , \ram[1][189] , \ram[1][188] , \ram[1][187] ,
         \ram[1][186] , \ram[1][185] , \ram[1][184] , \ram[1][183] ,
         \ram[1][182] , \ram[1][181] , \ram[1][180] , \ram[1][179] ,
         \ram[1][178] , \ram[1][177] , \ram[1][176] , \ram[1][175] ,
         \ram[1][174] , \ram[1][173] , \ram[1][172] , \ram[1][171] ,
         \ram[1][170] , \ram[1][169] , \ram[1][168] , \ram[1][167] ,
         \ram[1][166] , \ram[1][165] , \ram[1][164] , \ram[1][163] ,
         \ram[1][162] , \ram[1][161] , \ram[1][160] , \ram[1][159] ,
         \ram[1][158] , \ram[1][157] , \ram[1][156] , \ram[1][155] ,
         \ram[1][154] , \ram[1][153] , \ram[1][152] , \ram[1][151] ,
         \ram[1][150] , \ram[1][149] , \ram[1][148] , \ram[1][147] ,
         \ram[1][146] , \ram[1][145] , \ram[1][144] , \ram[1][143] ,
         \ram[1][142] , \ram[1][141] , \ram[1][140] , \ram[1][139] ,
         \ram[1][138] , \ram[1][137] , \ram[1][136] , \ram[1][135] ,
         \ram[1][134] , \ram[1][133] , \ram[1][132] , \ram[1][131] ,
         \ram[1][130] , \ram[1][129] , \ram[1][128] , \ram[1][127] ,
         \ram[1][126] , \ram[1][125] , \ram[1][124] , \ram[1][123] ,
         \ram[1][122] , \ram[1][121] , \ram[1][120] , \ram[1][119] ,
         \ram[1][118] , \ram[1][117] , \ram[1][116] , \ram[1][115] ,
         \ram[1][114] , \ram[1][113] , \ram[1][112] , \ram[1][111] ,
         \ram[1][110] , \ram[1][109] , \ram[1][108] , \ram[1][107] ,
         \ram[1][106] , \ram[1][105] , \ram[1][104] , \ram[1][103] ,
         \ram[1][102] , \ram[1][101] , \ram[1][100] , \ram[1][99] ,
         \ram[1][98] , \ram[1][97] , \ram[1][96] , \ram[1][95] , \ram[1][94] ,
         \ram[1][93] , \ram[1][92] , \ram[1][91] , \ram[1][90] , \ram[1][89] ,
         \ram[1][88] , \ram[1][87] , \ram[1][86] , \ram[1][85] , \ram[1][84] ,
         \ram[1][83] , \ram[1][82] , \ram[1][81] , \ram[1][80] , \ram[1][79] ,
         \ram[1][78] , \ram[1][77] , \ram[1][76] , \ram[1][75] , \ram[1][74] ,
         \ram[1][73] , \ram[1][72] , \ram[1][71] , \ram[1][70] , \ram[1][69] ,
         \ram[1][68] , \ram[1][67] , \ram[1][66] , \ram[1][65] , \ram[1][64] ,
         \ram[1][63] , \ram[1][62] , \ram[1][61] , \ram[1][60] , \ram[1][59] ,
         \ram[1][58] , \ram[1][57] , \ram[1][56] , \ram[1][55] , \ram[1][54] ,
         \ram[1][53] , \ram[1][52] , \ram[1][51] , \ram[1][50] , \ram[1][49] ,
         \ram[1][48] , \ram[1][47] , \ram[1][46] , \ram[1][45] , \ram[1][44] ,
         \ram[1][43] , \ram[1][42] , \ram[1][41] , \ram[1][40] , \ram[1][39] ,
         \ram[1][38] , \ram[1][37] , \ram[1][36] , \ram[1][35] , \ram[1][34] ,
         \ram[1][33] , \ram[1][32] , \ram[1][31] , \ram[1][30] , \ram[1][29] ,
         \ram[1][28] , \ram[1][27] , \ram[1][26] , \ram[1][25] , \ram[1][24] ,
         \ram[1][23] , \ram[1][22] , \ram[1][21] , \ram[1][20] , \ram[1][19] ,
         \ram[1][18] , \ram[1][17] , \ram[1][16] , \ram[1][15] , \ram[1][14] ,
         \ram[1][13] , \ram[1][12] , \ram[1][11] , \ram[1][10] , \ram[1][9] ,
         \ram[1][8] , \ram[1][7] , \ram[1][6] , \ram[1][5] , \ram[1][4] ,
         \ram[1][3] , \ram[1][2] , \ram[1][1] , \ram[1][0] , \ram[0][255] ,
         \ram[0][254] , \ram[0][253] , \ram[0][252] , \ram[0][251] ,
         \ram[0][250] , \ram[0][249] , \ram[0][248] , \ram[0][247] ,
         \ram[0][246] , \ram[0][245] , \ram[0][244] , \ram[0][243] ,
         \ram[0][242] , \ram[0][241] , \ram[0][240] , \ram[0][239] ,
         \ram[0][238] , \ram[0][237] , \ram[0][236] , \ram[0][235] ,
         \ram[0][234] , \ram[0][233] , \ram[0][232] , \ram[0][231] ,
         \ram[0][230] , \ram[0][229] , \ram[0][228] , \ram[0][227] ,
         \ram[0][226] , \ram[0][225] , \ram[0][224] , \ram[0][223] ,
         \ram[0][222] , \ram[0][221] , \ram[0][220] , \ram[0][219] ,
         \ram[0][218] , \ram[0][217] , \ram[0][216] , \ram[0][215] ,
         \ram[0][214] , \ram[0][213] , \ram[0][212] , \ram[0][211] ,
         \ram[0][210] , \ram[0][209] , \ram[0][208] , \ram[0][207] ,
         \ram[0][206] , \ram[0][205] , \ram[0][204] , \ram[0][203] ,
         \ram[0][202] , \ram[0][201] , \ram[0][200] , \ram[0][199] ,
         \ram[0][198] , \ram[0][197] , \ram[0][196] , \ram[0][195] ,
         \ram[0][194] , \ram[0][193] , \ram[0][192] , \ram[0][191] ,
         \ram[0][190] , \ram[0][189] , \ram[0][188] , \ram[0][187] ,
         \ram[0][186] , \ram[0][185] , \ram[0][184] , \ram[0][183] ,
         \ram[0][182] , \ram[0][181] , \ram[0][180] , \ram[0][179] ,
         \ram[0][178] , \ram[0][177] , \ram[0][176] , \ram[0][175] ,
         \ram[0][174] , \ram[0][173] , \ram[0][172] , \ram[0][171] ,
         \ram[0][170] , \ram[0][169] , \ram[0][168] , \ram[0][167] ,
         \ram[0][166] , \ram[0][165] , \ram[0][164] , \ram[0][163] ,
         \ram[0][162] , \ram[0][161] , \ram[0][160] , \ram[0][159] ,
         \ram[0][158] , \ram[0][157] , \ram[0][156] , \ram[0][155] ,
         \ram[0][154] , \ram[0][153] , \ram[0][152] , \ram[0][151] ,
         \ram[0][150] , \ram[0][149] , \ram[0][148] , \ram[0][147] ,
         \ram[0][146] , \ram[0][145] , \ram[0][143] , \ram[0][142] ,
         \ram[0][141] , \ram[0][140] , \ram[0][139] , \ram[0][138] ,
         \ram[0][137] , \ram[0][136] , \ram[0][135] , \ram[0][134] ,
         \ram[0][133] , \ram[0][132] , \ram[0][131] , \ram[0][130] ,
         \ram[0][129] , \ram[0][128] , \ram[0][127] , \ram[0][126] ,
         \ram[0][125] , \ram[0][124] , \ram[0][123] , \ram[0][122] ,
         \ram[0][121] , \ram[0][120] , \ram[0][119] , \ram[0][118] ,
         \ram[0][117] , \ram[0][116] , \ram[0][115] , \ram[0][114] ,
         \ram[0][113] , \ram[0][112] , \ram[0][111] , \ram[0][110] ,
         \ram[0][109] , \ram[0][108] , \ram[0][107] , \ram[0][106] ,
         \ram[0][105] , \ram[0][104] , \ram[0][103] , \ram[0][102] ,
         \ram[0][101] , \ram[0][100] , \ram[0][99] , \ram[0][98] ,
         \ram[0][97] , \ram[0][96] , \ram[0][95] , \ram[0][94] , \ram[0][93] ,
         \ram[0][92] , \ram[0][91] , \ram[0][90] , \ram[0][89] , \ram[0][88] ,
         \ram[0][87] , \ram[0][86] , \ram[0][85] , \ram[0][84] , \ram[0][83] ,
         \ram[0][82] , \ram[0][81] , \ram[0][80] , \ram[0][79] , \ram[0][78] ,
         \ram[0][77] , \ram[0][76] , \ram[0][75] , \ram[0][74] , \ram[0][73] ,
         \ram[0][72] , \ram[0][71] , \ram[0][70] , \ram[0][69] , \ram[0][68] ,
         \ram[0][67] , \ram[0][66] , \ram[0][65] , \ram[0][64] , \ram[0][63] ,
         \ram[0][62] , \ram[0][61] , \ram[0][60] , \ram[0][59] , \ram[0][58] ,
         \ram[0][57] , \ram[0][56] , \ram[0][55] , \ram[0][54] , \ram[0][53] ,
         \ram[0][52] , \ram[0][51] , \ram[0][50] , \ram[0][49] , \ram[0][48] ,
         \ram[0][47] , \ram[0][46] , \ram[0][45] , \ram[0][44] , \ram[0][43] ,
         \ram[0][42] , \ram[0][41] , \ram[0][40] , \ram[0][39] , \ram[0][38] ,
         \ram[0][37] , \ram[0][36] , \ram[0][35] , \ram[0][34] , \ram[0][33] ,
         \ram[0][32] , \ram[0][31] , \ram[0][30] , \ram[0][29] , \ram[0][28] ,
         \ram[0][27] , \ram[0][26] , \ram[0][25] , \ram[0][24] , \ram[0][23] ,
         \ram[0][22] , \ram[0][21] , \ram[0][20] , \ram[0][19] , \ram[0][18] ,
         \ram[0][17] , \ram[0][16] , \ram[0][15] , \ram[0][14] , \ram[0][13] ,
         \ram[0][12] , \ram[0][11] , \ram[0][10] , \ram[0][9] , \ram[0][8] ,
         \ram[0][7] , \ram[0][6] , \ram[0][5] , \ram[0][4] , \ram[0][3] ,
         \ram[0][2] , \ram[0][1] , \ram[0][0] , n7, n8, n9, n10, n12, n13, n16,
         n17, n18, n20, n21, n22, n24, n25, n28, n30, n33, n34, n37, n38, n40,
         n41, n44, n47, n49, n50, n51, n52, n53, n54, n55, n56, n57, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n830, n831, n832, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1138, n1139, n1140,
         n1141, n1142, n1143, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1358, n1360, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1390, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1462, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1799, n1800, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n1, n2,
         n3, n4, n5, n6, n11, n14, n15, n19, n23, n26, n27, n29, n31, n32, n35,
         n36, n39, n42, n43, n45, n46, n48, n58, n829, n833, n866, n877, n917,
         n1023, n1078, n1137, n1144, n1344, n1357, n1359, n1361, n1389, n1391,
         n1461, n1463, n1597, n1633, n1651, n1798, n1801, n3929, n3949, n4105,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381;
  assign N26 = addr[0];
  assign N27 = addr[1];
  assign N28 = addr[2];
  assign N29 = addr[3];

  DFFX1_HVT \ram_reg[15][255]  ( .D(n4156), .CLK(clk), .Q(\ram[15][255] ) );
  DFFX1_HVT \ram_reg[15][254]  ( .D(n4155), .CLK(clk), .Q(\ram[15][254] ) );
  DFFX1_HVT \ram_reg[15][253]  ( .D(n4154), .CLK(clk), .Q(\ram[15][253] ) );
  DFFX1_HVT \ram_reg[15][252]  ( .D(n4153), .CLK(clk), .Q(\ram[15][252] ) );
  DFFX1_HVT \ram_reg[15][251]  ( .D(n4152), .CLK(clk), .Q(\ram[15][251] ) );
  DFFX1_HVT \ram_reg[15][250]  ( .D(n4151), .CLK(clk), .Q(\ram[15][250] ) );
  DFFX1_HVT \ram_reg[15][249]  ( .D(n4150), .CLK(clk), .Q(\ram[15][249] ) );
  DFFX1_HVT \ram_reg[15][248]  ( .D(n4149), .CLK(clk), .Q(\ram[15][248] ) );
  DFFX1_HVT \ram_reg[15][247]  ( .D(n4148), .CLK(clk), .Q(\ram[15][247] ), 
        .QN(n5597) );
  DFFX1_HVT \ram_reg[15][246]  ( .D(n4147), .CLK(clk), .Q(\ram[15][246] ) );
  DFFX1_HVT \ram_reg[15][245]  ( .D(n4146), .CLK(clk), .Q(\ram[15][245] ) );
  DFFX1_HVT \ram_reg[15][244]  ( .D(n4145), .CLK(clk), .Q(\ram[15][244] ) );
  DFFX1_HVT \ram_reg[15][243]  ( .D(n4144), .CLK(clk), .Q(\ram[15][243] ) );
  DFFX1_HVT \ram_reg[15][242]  ( .D(n4143), .CLK(clk), .Q(\ram[15][242] ) );
  DFFX1_HVT \ram_reg[15][241]  ( .D(n4142), .CLK(clk), .Q(\ram[15][241] ) );
  DFFX1_HVT \ram_reg[15][240]  ( .D(n4141), .CLK(clk), .Q(\ram[15][240] ), 
        .QN(n5598) );
  DFFX1_HVT \ram_reg[15][239]  ( .D(n4140), .CLK(clk), .Q(\ram[15][239] ) );
  DFFX1_HVT \ram_reg[15][238]  ( .D(n4139), .CLK(clk), .Q(\ram[15][238] ) );
  DFFX1_HVT \ram_reg[15][237]  ( .D(n4138), .CLK(clk), .Q(\ram[15][237] ) );
  DFFX1_HVT \ram_reg[15][236]  ( .D(n4137), .CLK(clk), .Q(\ram[15][236] ) );
  DFFX1_HVT \ram_reg[15][235]  ( .D(n4136), .CLK(clk), .Q(\ram[15][235] ) );
  DFFX1_HVT \ram_reg[15][234]  ( .D(n4135), .CLK(clk), .Q(\ram[15][234] ) );
  DFFX1_HVT \ram_reg[15][233]  ( .D(n4134), .CLK(clk), .Q(\ram[15][233] ) );
  DFFX1_HVT \ram_reg[15][232]  ( .D(n4133), .CLK(clk), .Q(\ram[15][232] ) );
  DFFX1_HVT \ram_reg[15][231]  ( .D(n4132), .CLK(clk), .Q(\ram[15][231] ) );
  DFFX1_HVT \ram_reg[15][230]  ( .D(n4131), .CLK(clk), .Q(\ram[15][230] ) );
  DFFX1_HVT \ram_reg[15][229]  ( .D(n4130), .CLK(clk), .Q(\ram[15][229] ) );
  DFFX1_HVT \ram_reg[15][228]  ( .D(n4129), .CLK(clk), .Q(\ram[15][228] ) );
  DFFX1_HVT \ram_reg[15][227]  ( .D(n4128), .CLK(clk), .Q(\ram[15][227] ) );
  DFFX1_HVT \ram_reg[15][226]  ( .D(n4127), .CLK(clk), .Q(\ram[15][226] ) );
  DFFX1_HVT \ram_reg[15][225]  ( .D(n4126), .CLK(clk), .Q(\ram[15][225] ) );
  DFFX1_HVT \ram_reg[15][224]  ( .D(n4125), .CLK(clk), .Q(\ram[15][224] ) );
  DFFX1_HVT \ram_reg[15][223]  ( .D(n4124), .CLK(clk), .Q(\ram[15][223] ) );
  DFFX1_HVT \ram_reg[15][222]  ( .D(n4123), .CLK(clk), .Q(\ram[15][222] ) );
  DFFX1_HVT \ram_reg[15][221]  ( .D(n4122), .CLK(clk), .Q(\ram[15][221] ) );
  DFFX1_HVT \ram_reg[15][220]  ( .D(n4121), .CLK(clk), .Q(\ram[15][220] ) );
  DFFX1_HVT \ram_reg[15][219]  ( .D(n4120), .CLK(clk), .Q(\ram[15][219] ) );
  DFFX1_HVT \ram_reg[15][218]  ( .D(n4119), .CLK(clk), .Q(\ram[15][218] ) );
  DFFX1_HVT \ram_reg[15][217]  ( .D(n4118), .CLK(clk), .Q(\ram[15][217] ) );
  DFFX1_HVT \ram_reg[15][216]  ( .D(n4117), .CLK(clk), .Q(\ram[15][216] ) );
  DFFX1_HVT \ram_reg[15][215]  ( .D(n4116), .CLK(clk), .Q(\ram[15][215] ) );
  DFFX1_HVT \ram_reg[15][214]  ( .D(n4115), .CLK(clk), .Q(\ram[15][214] ) );
  DFFX1_HVT \ram_reg[15][213]  ( .D(n4114), .CLK(clk), .Q(\ram[15][213] ) );
  DFFX1_HVT \ram_reg[15][212]  ( .D(n4113), .CLK(clk), .Q(\ram[15][212] ) );
  DFFX1_HVT \ram_reg[15][211]  ( .D(n4112), .CLK(clk), .Q(\ram[15][211] ) );
  DFFX1_HVT \ram_reg[15][210]  ( .D(n4111), .CLK(clk), .Q(\ram[15][210] ) );
  DFFX1_HVT \ram_reg[15][209]  ( .D(n4110), .CLK(clk), .Q(\ram[15][209] ) );
  DFFX1_HVT \ram_reg[15][208]  ( .D(n4109), .CLK(clk), .Q(\ram[15][208] ) );
  DFFX1_HVT \ram_reg[15][207]  ( .D(n4108), .CLK(clk), .Q(\ram[15][207] ) );
  DFFX1_HVT \ram_reg[15][206]  ( .D(n4107), .CLK(clk), .Q(\ram[15][206] ) );
  DFFX1_HVT \ram_reg[15][205]  ( .D(n4106), .CLK(clk), .Q(\ram[15][205] ) );
  DFFX1_HVT \ram_reg[15][204]  ( .D(n5024), .CLK(clk), .Q(\ram[15][204] ), 
        .QN(n5897) );
  DFFX1_HVT \ram_reg[15][203]  ( .D(n4104), .CLK(clk), .Q(\ram[15][203] ) );
  DFFX1_HVT \ram_reg[15][202]  ( .D(n4103), .CLK(clk), .Q(\ram[15][202] ) );
  DFFX1_HVT \ram_reg[15][201]  ( .D(n4102), .CLK(clk), .Q(\ram[15][201] ) );
  DFFX1_HVT \ram_reg[15][200]  ( .D(n4101), .CLK(clk), .Q(\ram[15][200] ) );
  DFFX1_HVT \ram_reg[15][199]  ( .D(n4100), .CLK(clk), .Q(\ram[15][199] ) );
  DFFX1_HVT \ram_reg[15][198]  ( .D(n4099), .CLK(clk), .Q(\ram[15][198] ) );
  DFFX1_HVT \ram_reg[15][197]  ( .D(n4098), .CLK(clk), .Q(\ram[15][197] ) );
  DFFX1_HVT \ram_reg[15][196]  ( .D(n4097), .CLK(clk), .Q(\ram[15][196] ) );
  DFFX1_HVT \ram_reg[15][195]  ( .D(n4096), .CLK(clk), .Q(\ram[15][195] ) );
  DFFX1_HVT \ram_reg[15][194]  ( .D(n4095), .CLK(clk), .Q(\ram[15][194] ) );
  DFFX1_HVT \ram_reg[15][193]  ( .D(n4094), .CLK(clk), .Q(\ram[15][193] ) );
  DFFX1_HVT \ram_reg[15][192]  ( .D(n4093), .CLK(clk), .Q(\ram[15][192] ) );
  DFFX1_HVT \ram_reg[15][191]  ( .D(n4092), .CLK(clk), .Q(\ram[15][191] ) );
  DFFX1_HVT \ram_reg[15][190]  ( .D(n4091), .CLK(clk), .Q(\ram[15][190] ) );
  DFFX1_HVT \ram_reg[15][189]  ( .D(n4090), .CLK(clk), .Q(\ram[15][189] ) );
  DFFX1_HVT \ram_reg[15][188]  ( .D(n4089), .CLK(clk), .Q(\ram[15][188] ) );
  DFFX1_HVT \ram_reg[15][187]  ( .D(n4088), .CLK(clk), .Q(\ram[15][187] ) );
  DFFX1_HVT \ram_reg[15][186]  ( .D(n4087), .CLK(clk), .Q(\ram[15][186] ) );
  DFFX1_HVT \ram_reg[15][185]  ( .D(n4086), .CLK(clk), .Q(\ram[15][185] ) );
  DFFX1_HVT \ram_reg[15][184]  ( .D(n4085), .CLK(clk), .Q(\ram[15][184] ) );
  DFFX1_HVT \ram_reg[15][183]  ( .D(n4084), .CLK(clk), .Q(\ram[15][183] ) );
  DFFX1_HVT \ram_reg[15][182]  ( .D(n4083), .CLK(clk), .Q(\ram[15][182] ) );
  DFFX1_HVT \ram_reg[15][181]  ( .D(n4082), .CLK(clk), .Q(\ram[15][181] ) );
  DFFX1_HVT \ram_reg[15][180]  ( .D(n4081), .CLK(clk), .Q(\ram[15][180] ) );
  DFFX1_HVT \ram_reg[15][179]  ( .D(n4080), .CLK(clk), .Q(\ram[15][179] ) );
  DFFX1_HVT \ram_reg[15][178]  ( .D(n4079), .CLK(clk), .Q(\ram[15][178] ) );
  DFFX1_HVT \ram_reg[15][177]  ( .D(n4078), .CLK(clk), .Q(\ram[15][177] ) );
  DFFX1_HVT \ram_reg[15][176]  ( .D(n4077), .CLK(clk), .Q(\ram[15][176] ) );
  DFFX1_HVT \ram_reg[15][175]  ( .D(n4076), .CLK(clk), .Q(\ram[15][175] ) );
  DFFX1_HVT \ram_reg[15][174]  ( .D(n4075), .CLK(clk), .Q(\ram[15][174] ) );
  DFFX1_HVT \ram_reg[15][173]  ( .D(n4074), .CLK(clk), .Q(\ram[15][173] ) );
  DFFX1_HVT \ram_reg[15][172]  ( .D(n4073), .CLK(clk), .Q(\ram[15][172] ) );
  DFFX1_HVT \ram_reg[15][171]  ( .D(n4072), .CLK(clk), .Q(\ram[15][171] ) );
  DFFX1_HVT \ram_reg[15][170]  ( .D(n4071), .CLK(clk), .Q(\ram[15][170] ) );
  DFFX1_HVT \ram_reg[15][169]  ( .D(n4070), .CLK(clk), .Q(\ram[15][169] ) );
  DFFX1_HVT \ram_reg[15][168]  ( .D(n4069), .CLK(clk), .Q(\ram[15][168] ) );
  DFFX1_HVT \ram_reg[15][167]  ( .D(n4068), .CLK(clk), .Q(\ram[15][167] ) );
  DFFX1_HVT \ram_reg[15][166]  ( .D(n4067), .CLK(clk), .Q(\ram[15][166] ) );
  DFFX1_HVT \ram_reg[15][165]  ( .D(n4066), .CLK(clk), .Q(\ram[15][165] ) );
  DFFX1_HVT \ram_reg[15][164]  ( .D(n4065), .CLK(clk), .Q(\ram[15][164] ) );
  DFFX1_HVT \ram_reg[15][163]  ( .D(n4064), .CLK(clk), .Q(\ram[15][163] ) );
  DFFX1_HVT \ram_reg[15][162]  ( .D(n4063), .CLK(clk), .Q(\ram[15][162] ) );
  DFFX1_HVT \ram_reg[15][161]  ( .D(n4062), .CLK(clk), .Q(\ram[15][161] ) );
  DFFX1_HVT \ram_reg[15][160]  ( .D(n4061), .CLK(clk), .Q(\ram[15][160] ) );
  DFFX1_HVT \ram_reg[15][159]  ( .D(n4060), .CLK(clk), .Q(\ram[15][159] ) );
  DFFX1_HVT \ram_reg[15][158]  ( .D(n4059), .CLK(clk), .Q(\ram[15][158] ) );
  DFFX1_HVT \ram_reg[15][157]  ( .D(n4058), .CLK(clk), .Q(\ram[15][157] ) );
  DFFX1_HVT \ram_reg[15][156]  ( .D(n4057), .CLK(clk), .Q(\ram[15][156] ) );
  DFFX1_HVT \ram_reg[15][155]  ( .D(n4056), .CLK(clk), .Q(\ram[15][155] ) );
  DFFX1_HVT \ram_reg[15][154]  ( .D(n4055), .CLK(clk), .Q(\ram[15][154] ) );
  DFFX1_HVT \ram_reg[15][153]  ( .D(n4054), .CLK(clk), .Q(\ram[15][153] ) );
  DFFX1_HVT \ram_reg[15][152]  ( .D(n4053), .CLK(clk), .Q(\ram[15][152] ), 
        .QN(n5530) );
  DFFX1_HVT \ram_reg[15][151]  ( .D(n4052), .CLK(clk), .Q(\ram[15][151] ) );
  DFFX1_HVT \ram_reg[15][150]  ( .D(n4051), .CLK(clk), .Q(\ram[15][150] ) );
  DFFX1_HVT \ram_reg[15][149]  ( .D(n4050), .CLK(clk), .Q(\ram[15][149] ) );
  DFFX1_HVT \ram_reg[15][148]  ( .D(n4049), .CLK(clk), .Q(\ram[15][148] ), 
        .QN(n5599) );
  DFFX1_HVT \ram_reg[15][147]  ( .D(n4048), .CLK(clk), .Q(\ram[15][147] ) );
  DFFX1_HVT \ram_reg[15][146]  ( .D(n4047), .CLK(clk), .Q(\ram[15][146] ) );
  DFFX1_HVT \ram_reg[15][145]  ( .D(n4046), .CLK(clk), .Q(\ram[15][145] ) );
  DFFX1_HVT \ram_reg[15][144]  ( .D(n4045), .CLK(clk), .Q(\ram[15][144] ) );
  DFFX1_HVT \ram_reg[15][143]  ( .D(n4044), .CLK(clk), .Q(\ram[15][143] ) );
  DFFX1_HVT \ram_reg[15][142]  ( .D(n4043), .CLK(clk), .Q(\ram[15][142] ) );
  DFFX1_HVT \ram_reg[15][141]  ( .D(n4042), .CLK(clk), .Q(\ram[15][141] ) );
  DFFX1_HVT \ram_reg[15][140]  ( .D(n4041), .CLK(clk), .Q(\ram[15][140] ) );
  DFFX1_HVT \ram_reg[15][139]  ( .D(n4040), .CLK(clk), .Q(\ram[15][139] ) );
  DFFX1_HVT \ram_reg[15][138]  ( .D(n4039), .CLK(clk), .Q(\ram[15][138] ) );
  DFFX1_HVT \ram_reg[15][137]  ( .D(n4038), .CLK(clk), .Q(\ram[15][137] ) );
  DFFX1_HVT \ram_reg[15][136]  ( .D(n4037), .CLK(clk), .Q(\ram[15][136] ) );
  DFFX1_HVT \ram_reg[15][135]  ( .D(n4036), .CLK(clk), .Q(\ram[15][135] ) );
  DFFX1_HVT \ram_reg[15][134]  ( .D(n4035), .CLK(clk), .Q(\ram[15][134] ) );
  DFFX1_HVT \ram_reg[15][133]  ( .D(n4034), .CLK(clk), .Q(\ram[15][133] ) );
  DFFX1_HVT \ram_reg[15][132]  ( .D(n4033), .CLK(clk), .Q(\ram[15][132] ) );
  DFFX1_HVT \ram_reg[15][131]  ( .D(n4032), .CLK(clk), .Q(\ram[15][131] ) );
  DFFX1_HVT \ram_reg[15][130]  ( .D(n4031), .CLK(clk), .Q(\ram[15][130] ) );
  DFFX1_HVT \ram_reg[15][129]  ( .D(n4030), .CLK(clk), .Q(\ram[15][129] ) );
  DFFX1_HVT \ram_reg[15][128]  ( .D(n4029), .CLK(clk), .Q(\ram[15][128] ) );
  DFFX1_HVT \ram_reg[15][127]  ( .D(n4028), .CLK(clk), .Q(\ram[15][127] ) );
  DFFX1_HVT \ram_reg[15][126]  ( .D(n4027), .CLK(clk), .Q(\ram[15][126] ) );
  DFFX1_HVT \ram_reg[15][125]  ( .D(n4026), .CLK(clk), .Q(\ram[15][125] ) );
  DFFX1_HVT \ram_reg[15][124]  ( .D(n4025), .CLK(clk), .Q(\ram[15][124] ) );
  DFFX1_HVT \ram_reg[15][123]  ( .D(n4024), .CLK(clk), .Q(\ram[15][123] ) );
  DFFX1_HVT \ram_reg[15][122]  ( .D(n4023), .CLK(clk), .Q(\ram[15][122] ) );
  DFFX1_HVT \ram_reg[15][121]  ( .D(n4022), .CLK(clk), .Q(\ram[15][121] ) );
  DFFX1_HVT \ram_reg[15][120]  ( .D(n4021), .CLK(clk), .Q(\ram[15][120] ) );
  DFFX1_HVT \ram_reg[15][119]  ( .D(n4020), .CLK(clk), .Q(\ram[15][119] ) );
  DFFX1_HVT \ram_reg[15][118]  ( .D(n4019), .CLK(clk), .Q(\ram[15][118] ) );
  DFFX1_HVT \ram_reg[15][117]  ( .D(n4018), .CLK(clk), .Q(\ram[15][117] ) );
  DFFX1_HVT \ram_reg[15][116]  ( .D(n4017), .CLK(clk), .Q(\ram[15][116] ) );
  DFFX1_HVT \ram_reg[15][115]  ( .D(n4016), .CLK(clk), .Q(\ram[15][115] ) );
  DFFX1_HVT \ram_reg[15][114]  ( .D(n4015), .CLK(clk), .Q(\ram[15][114] ) );
  DFFX1_HVT \ram_reg[15][113]  ( .D(n4014), .CLK(clk), .Q(\ram[15][113] ) );
  DFFX1_HVT \ram_reg[15][112]  ( .D(n4013), .CLK(clk), .Q(\ram[15][112] ) );
  DFFX1_HVT \ram_reg[15][111]  ( .D(n4012), .CLK(clk), .Q(\ram[15][111] ) );
  DFFX1_HVT \ram_reg[15][110]  ( .D(n4011), .CLK(clk), .Q(\ram[15][110] ) );
  DFFX1_HVT \ram_reg[15][109]  ( .D(n4010), .CLK(clk), .Q(\ram[15][109] ) );
  DFFX1_HVT \ram_reg[15][108]  ( .D(n4009), .CLK(clk), .Q(\ram[15][108] ) );
  DFFX1_HVT \ram_reg[15][107]  ( .D(n4008), .CLK(clk), .Q(\ram[15][107] ) );
  DFFX1_HVT \ram_reg[15][106]  ( .D(n4007), .CLK(clk), .Q(\ram[15][106] ) );
  DFFX1_HVT \ram_reg[15][105]  ( .D(n4006), .CLK(clk), .Q(\ram[15][105] ) );
  DFFX1_HVT \ram_reg[15][104]  ( .D(n4005), .CLK(clk), .Q(\ram[15][104] ) );
  DFFX1_HVT \ram_reg[15][103]  ( .D(n4004), .CLK(clk), .QN(n5856) );
  DFFX1_HVT \ram_reg[15][102]  ( .D(n4003), .CLK(clk), .Q(\ram[15][102] ) );
  DFFX1_HVT \ram_reg[15][101]  ( .D(n4002), .CLK(clk), .Q(\ram[15][101] ), 
        .QN(n4809) );
  DFFX1_HVT \ram_reg[15][100]  ( .D(n4001), .CLK(clk), .Q(\ram[15][100] ) );
  DFFX1_HVT \ram_reg[15][99]  ( .D(n4000), .CLK(clk), .Q(\ram[15][99] ) );
  DFFX1_HVT \ram_reg[15][98]  ( .D(n3999), .CLK(clk), .Q(\ram[15][98] ) );
  DFFX1_HVT \ram_reg[15][97]  ( .D(n3998), .CLK(clk), .Q(\ram[15][97] ) );
  DFFX1_HVT \ram_reg[15][96]  ( .D(n3997), .CLK(clk), .Q(\ram[15][96] ) );
  DFFX1_HVT \ram_reg[15][95]  ( .D(n3996), .CLK(clk), .Q(\ram[15][95] ) );
  DFFX1_HVT \ram_reg[15][94]  ( .D(n3995), .CLK(clk), .Q(\ram[15][94] ) );
  DFFX1_HVT \ram_reg[15][93]  ( .D(n3994), .CLK(clk), .Q(\ram[15][93] ) );
  DFFX1_HVT \ram_reg[15][92]  ( .D(n3993), .CLK(clk), .Q(\ram[15][92] ) );
  DFFX1_HVT \ram_reg[15][91]  ( .D(n3992), .CLK(clk), .Q(\ram[15][91] ) );
  DFFX1_HVT \ram_reg[15][90]  ( .D(n3991), .CLK(clk), .Q(\ram[15][90] ) );
  DFFX1_HVT \ram_reg[15][89]  ( .D(n3990), .CLK(clk), .Q(\ram[15][89] ) );
  DFFX1_HVT \ram_reg[15][88]  ( .D(n3989), .CLK(clk), .Q(\ram[15][88] ) );
  DFFX1_HVT \ram_reg[15][87]  ( .D(n3988), .CLK(clk), .Q(\ram[15][87] ) );
  DFFX1_HVT \ram_reg[15][86]  ( .D(n3987), .CLK(clk), .Q(\ram[15][86] ) );
  DFFX1_HVT \ram_reg[15][85]  ( .D(n3986), .CLK(clk), .Q(\ram[15][85] ) );
  DFFX1_HVT \ram_reg[15][84]  ( .D(n3985), .CLK(clk), .Q(\ram[15][84] ) );
  DFFX1_HVT \ram_reg[15][83]  ( .D(n3984), .CLK(clk), .Q(\ram[15][83] ), .QN(
        n5522) );
  DFFX1_HVT \ram_reg[15][82]  ( .D(n3983), .CLK(clk), .Q(\ram[15][82] ) );
  DFFX1_HVT \ram_reg[15][81]  ( .D(n3982), .CLK(clk), .Q(\ram[15][81] ) );
  DFFX1_HVT \ram_reg[15][80]  ( .D(n3981), .CLK(clk), .Q(\ram[15][80] ) );
  DFFX1_HVT \ram_reg[15][79]  ( .D(n3980), .CLK(clk), .Q(\ram[15][79] ) );
  DFFX1_HVT \ram_reg[15][78]  ( .D(n3979), .CLK(clk), .Q(\ram[15][78] ) );
  DFFX1_HVT \ram_reg[15][77]  ( .D(n3978), .CLK(clk), .Q(\ram[15][77] ) );
  DFFX1_HVT \ram_reg[15][76]  ( .D(n3977), .CLK(clk), .Q(\ram[15][76] ) );
  DFFX1_HVT \ram_reg[15][75]  ( .D(n3976), .CLK(clk), .Q(\ram[15][75] ), .QN(
        n5498) );
  DFFX1_HVT \ram_reg[15][74]  ( .D(n3975), .CLK(clk), .Q(\ram[15][74] ) );
  DFFX1_HVT \ram_reg[15][73]  ( .D(n3974), .CLK(clk), .Q(\ram[15][73] ) );
  DFFX1_HVT \ram_reg[15][72]  ( .D(n3973), .CLK(clk), .Q(\ram[15][72] ) );
  DFFX1_HVT \ram_reg[15][71]  ( .D(n3972), .CLK(clk), .Q(\ram[15][71] ) );
  DFFX1_HVT \ram_reg[15][70]  ( .D(n3971), .CLK(clk), .Q(\ram[15][70] ) );
  DFFX1_HVT \ram_reg[15][69]  ( .D(n3970), .CLK(clk), .Q(\ram[15][69] ) );
  DFFX1_HVT \ram_reg[15][68]  ( .D(n3969), .CLK(clk), .Q(\ram[15][68] ) );
  DFFX1_HVT \ram_reg[15][67]  ( .D(n3968), .CLK(clk), .Q(\ram[15][67] ) );
  DFFX1_HVT \ram_reg[15][66]  ( .D(n3967), .CLK(clk), .Q(\ram[15][66] ) );
  DFFX1_HVT \ram_reg[15][65]  ( .D(n3966), .CLK(clk), .Q(\ram[15][65] ), .QN(
        n4882) );
  DFFX1_HVT \ram_reg[15][64]  ( .D(n3965), .CLK(clk), .Q(\ram[15][64] ) );
  DFFX1_HVT \ram_reg[15][63]  ( .D(n3964), .CLK(clk), .Q(\ram[15][63] ) );
  DFFX1_HVT \ram_reg[15][62]  ( .D(n3963), .CLK(clk), .Q(\ram[15][62] ) );
  DFFX1_HVT \ram_reg[15][61]  ( .D(n3962), .CLK(clk), .Q(\ram[15][61] ) );
  DFFX1_HVT \ram_reg[15][60]  ( .D(n3961), .CLK(clk), .Q(\ram[15][60] ) );
  DFFX1_HVT \ram_reg[15][59]  ( .D(n3960), .CLK(clk), .Q(\ram[15][59] ) );
  DFFX1_HVT \ram_reg[15][58]  ( .D(n3959), .CLK(clk), .Q(\ram[15][58] ) );
  DFFX1_HVT \ram_reg[15][57]  ( .D(n3958), .CLK(clk), .Q(\ram[15][57] ) );
  DFFX1_HVT \ram_reg[15][56]  ( .D(n3957), .CLK(clk), .Q(\ram[15][56] ) );
  DFFX1_HVT \ram_reg[15][55]  ( .D(n3956), .CLK(clk), .Q(\ram[15][55] ) );
  DFFX1_HVT \ram_reg[15][54]  ( .D(n3955), .CLK(clk), .Q(\ram[15][54] ) );
  DFFX1_HVT \ram_reg[15][53]  ( .D(n3954), .CLK(clk), .Q(\ram[15][53] ) );
  DFFX1_HVT \ram_reg[15][52]  ( .D(n3953), .CLK(clk), .Q(\ram[15][52] ) );
  DFFX1_HVT \ram_reg[15][51]  ( .D(n3952), .CLK(clk), .Q(\ram[15][51] ) );
  DFFX1_HVT \ram_reg[15][50]  ( .D(n3951), .CLK(clk), .Q(\ram[15][50] ) );
  DFFX1_HVT \ram_reg[15][49]  ( .D(n3950), .CLK(clk), .Q(\ram[15][49] ) );
  DFFX1_HVT \ram_reg[15][48]  ( .D(n5035), .CLK(clk), .Q(\ram[15][48] ), .QN(
        n6016) );
  DFFX1_HVT \ram_reg[15][47]  ( .D(n3948), .CLK(clk), .Q(\ram[15][47] ) );
  DFFX1_HVT \ram_reg[15][46]  ( .D(n3947), .CLK(clk), .Q(\ram[15][46] ) );
  DFFX1_HVT \ram_reg[15][45]  ( .D(n3946), .CLK(clk), .Q(\ram[15][45] ) );
  DFFX1_HVT \ram_reg[15][44]  ( .D(n3945), .CLK(clk), .Q(\ram[15][44] ) );
  DFFX1_HVT \ram_reg[15][43]  ( .D(n3944), .CLK(clk), .Q(\ram[15][43] ) );
  DFFX1_HVT \ram_reg[15][42]  ( .D(n3943), .CLK(clk), .Q(\ram[15][42] ) );
  DFFX1_HVT \ram_reg[15][41]  ( .D(n3942), .CLK(clk), .Q(\ram[15][41] ) );
  DFFX1_HVT \ram_reg[15][40]  ( .D(n3941), .CLK(clk), .Q(\ram[15][40] ) );
  DFFX1_HVT \ram_reg[15][39]  ( .D(n3940), .CLK(clk), .Q(\ram[15][39] ) );
  DFFX1_HVT \ram_reg[15][38]  ( .D(n3939), .CLK(clk), .Q(\ram[15][38] ) );
  DFFX1_HVT \ram_reg[15][37]  ( .D(n3938), .CLK(clk), .Q(\ram[15][37] ) );
  DFFX1_HVT \ram_reg[15][36]  ( .D(n3937), .CLK(clk), .Q(\ram[15][36] ) );
  DFFX1_HVT \ram_reg[15][35]  ( .D(n3936), .CLK(clk), .Q(\ram[15][35] ) );
  DFFX1_HVT \ram_reg[15][34]  ( .D(n3935), .CLK(clk), .Q(\ram[15][34] ) );
  DFFX1_HVT \ram_reg[15][33]  ( .D(n3934), .CLK(clk), .Q(\ram[15][33] ) );
  DFFX1_HVT \ram_reg[15][32]  ( .D(n3933), .CLK(clk), .Q(\ram[15][32] ) );
  DFFX1_HVT \ram_reg[15][31]  ( .D(n3932), .CLK(clk), .Q(\ram[15][31] ) );
  DFFX1_HVT \ram_reg[15][30]  ( .D(n3931), .CLK(clk), .Q(\ram[15][30] ), .QN(
        n5521) );
  DFFX1_HVT \ram_reg[15][29]  ( .D(n3930), .CLK(clk), .Q(\ram[15][29] ) );
  DFFX1_HVT \ram_reg[15][28]  ( .D(n5036), .CLK(clk), .Q(\ram[15][28] ), .QN(
        n5604) );
  DFFX1_HVT \ram_reg[15][27]  ( .D(n3928), .CLK(clk), .Q(\ram[15][27] ), .QN(
        n5524) );
  DFFX1_HVT \ram_reg[15][26]  ( .D(n3927), .CLK(clk), .Q(\ram[15][26] ), .QN(
        n4196) );
  DFFX1_HVT \ram_reg[15][25]  ( .D(n3926), .CLK(clk), .Q(\ram[15][25] ) );
  DFFX1_HVT \ram_reg[15][24]  ( .D(n3925), .CLK(clk), .Q(\ram[15][24] ) );
  DFFX1_HVT \ram_reg[15][23]  ( .D(n3924), .CLK(clk), .Q(\ram[15][23] ) );
  DFFX1_HVT \ram_reg[15][22]  ( .D(n3923), .CLK(clk), .Q(\ram[15][22] ) );
  DFFX1_HVT \ram_reg[15][21]  ( .D(n3922), .CLK(clk), .Q(\ram[15][21] ) );
  DFFX1_HVT \ram_reg[15][20]  ( .D(n3921), .CLK(clk), .Q(\ram[15][20] ) );
  DFFX1_HVT \ram_reg[15][19]  ( .D(n3920), .CLK(clk), .Q(\ram[15][19] ) );
  DFFX1_HVT \ram_reg[15][18]  ( .D(n3919), .CLK(clk), .Q(\ram[15][18] ) );
  DFFX1_HVT \ram_reg[15][17]  ( .D(n3918), .CLK(clk), .Q(\ram[15][17] ) );
  DFFX1_HVT \ram_reg[15][16]  ( .D(n3917), .CLK(clk), .Q(\ram[15][16] ) );
  DFFX1_HVT \ram_reg[15][15]  ( .D(n3916), .CLK(clk), .Q(\ram[15][15] ) );
  DFFX1_HVT \ram_reg[15][14]  ( .D(n3915), .CLK(clk), .Q(\ram[15][14] ) );
  DFFX1_HVT \ram_reg[15][13]  ( .D(n3914), .CLK(clk), .Q(\ram[15][13] ) );
  DFFX1_HVT \ram_reg[15][12]  ( .D(n3913), .CLK(clk), .Q(\ram[15][12] ), .QN(
        n5529) );
  DFFX1_HVT \ram_reg[15][11]  ( .D(n3912), .CLK(clk), .Q(\ram[15][11] ) );
  DFFX1_HVT \ram_reg[15][10]  ( .D(n3911), .CLK(clk), .Q(\ram[15][10] ) );
  DFFX1_HVT \ram_reg[15][9]  ( .D(n3910), .CLK(clk), .Q(\ram[15][9] ) );
  DFFX1_HVT \ram_reg[15][8]  ( .D(n3909), .CLK(clk), .Q(\ram[15][8] ) );
  DFFX1_HVT \ram_reg[15][7]  ( .D(n3908), .CLK(clk), .Q(\ram[15][7] ) );
  DFFX1_HVT \ram_reg[15][6]  ( .D(n3907), .CLK(clk), .Q(\ram[15][6] ) );
  DFFX1_HVT \ram_reg[15][5]  ( .D(n3906), .CLK(clk), .Q(\ram[15][5] ) );
  DFFX1_HVT \ram_reg[15][4]  ( .D(n3905), .CLK(clk), .Q(\ram[15][4] ) );
  DFFX1_HVT \ram_reg[15][3]  ( .D(n3904), .CLK(clk), .Q(\ram[15][3] ) );
  DFFX1_HVT \ram_reg[15][2]  ( .D(n3903), .CLK(clk), .Q(\ram[15][2] ) );
  DFFX1_HVT \ram_reg[15][1]  ( .D(n3902), .CLK(clk), .Q(\ram[15][1] ) );
  DFFX1_HVT \ram_reg[15][0]  ( .D(n3901), .CLK(clk), .Q(\ram[15][0] ) );
  DFFX1_HVT \ram_reg[14][255]  ( .D(n3900), .CLK(clk), .Q(\ram[14][255] ) );
  DFFX1_HVT \ram_reg[14][254]  ( .D(n3899), .CLK(clk), .Q(\ram[14][254] ) );
  DFFX1_HVT \ram_reg[14][253]  ( .D(n3898), .CLK(clk), .Q(\ram[14][253] ) );
  DFFX1_HVT \ram_reg[14][252]  ( .D(n3897), .CLK(clk), .Q(\ram[14][252] ) );
  DFFX1_HVT \ram_reg[14][251]  ( .D(n3896), .CLK(clk), .Q(\ram[14][251] ) );
  DFFX1_HVT \ram_reg[14][250]  ( .D(n3895), .CLK(clk), .Q(\ram[14][250] ) );
  DFFX1_HVT \ram_reg[14][249]  ( .D(n3894), .CLK(clk), .Q(\ram[14][249] ) );
  DFFX1_HVT \ram_reg[14][248]  ( .D(n3893), .CLK(clk), .Q(\ram[14][248] ) );
  DFFX1_HVT \ram_reg[14][247]  ( .D(n3892), .CLK(clk), .Q(\ram[14][247] ) );
  DFFX1_HVT \ram_reg[14][246]  ( .D(n3891), .CLK(clk), .Q(\ram[14][246] ) );
  DFFX1_HVT \ram_reg[14][245]  ( .D(n3890), .CLK(clk), .Q(\ram[14][245] ) );
  DFFX1_HVT \ram_reg[14][244]  ( .D(n3889), .CLK(clk), .Q(\ram[14][244] ) );
  DFFX1_HVT \ram_reg[14][243]  ( .D(n3888), .CLK(clk), .Q(\ram[14][243] ) );
  DFFX1_HVT \ram_reg[14][242]  ( .D(n3887), .CLK(clk), .Q(\ram[14][242] ) );
  DFFX1_HVT \ram_reg[14][241]  ( .D(n3886), .CLK(clk), .Q(\ram[14][241] ) );
  DFFX1_HVT \ram_reg[14][240]  ( .D(n3885), .CLK(clk), .Q(\ram[14][240] ) );
  DFFX1_HVT \ram_reg[14][239]  ( .D(n3884), .CLK(clk), .Q(\ram[14][239] ) );
  DFFX1_HVT \ram_reg[14][238]  ( .D(n3883), .CLK(clk), .Q(\ram[14][238] ) );
  DFFX1_HVT \ram_reg[14][237]  ( .D(n3882), .CLK(clk), .Q(\ram[14][237] ) );
  DFFX1_HVT \ram_reg[14][236]  ( .D(n3881), .CLK(clk), .Q(\ram[14][236] ) );
  DFFX1_HVT \ram_reg[14][235]  ( .D(n3880), .CLK(clk), .Q(\ram[14][235] ) );
  DFFX1_HVT \ram_reg[14][234]  ( .D(n3879), .CLK(clk), .Q(\ram[14][234] ) );
  DFFX1_HVT \ram_reg[14][233]  ( .D(n3878), .CLK(clk), .Q(\ram[14][233] ) );
  DFFX1_HVT \ram_reg[14][232]  ( .D(n3877), .CLK(clk), .Q(\ram[14][232] ) );
  DFFX1_HVT \ram_reg[14][231]  ( .D(n3876), .CLK(clk), .Q(\ram[14][231] ) );
  DFFX1_HVT \ram_reg[14][230]  ( .D(n3875), .CLK(clk), .Q(\ram[14][230] ) );
  DFFX1_HVT \ram_reg[14][229]  ( .D(n3874), .CLK(clk), .Q(\ram[14][229] ) );
  DFFX1_HVT \ram_reg[14][228]  ( .D(n3873), .CLK(clk), .Q(\ram[14][228] ) );
  DFFX1_HVT \ram_reg[14][227]  ( .D(n3872), .CLK(clk), .Q(\ram[14][227] ) );
  DFFX1_HVT \ram_reg[14][226]  ( .D(n3871), .CLK(clk), .Q(\ram[14][226] ) );
  DFFX1_HVT \ram_reg[14][225]  ( .D(n3870), .CLK(clk), .Q(\ram[14][225] ) );
  DFFX1_HVT \ram_reg[14][224]  ( .D(n3869), .CLK(clk), .Q(\ram[14][224] ) );
  DFFX1_HVT \ram_reg[14][223]  ( .D(n3868), .CLK(clk), .Q(\ram[14][223] ) );
  DFFX1_HVT \ram_reg[14][222]  ( .D(n3867), .CLK(clk), .Q(\ram[14][222] ) );
  DFFX1_HVT \ram_reg[14][221]  ( .D(n3866), .CLK(clk), .Q(\ram[14][221] ) );
  DFFX1_HVT \ram_reg[14][220]  ( .D(n3865), .CLK(clk), .Q(\ram[14][220] ) );
  DFFX1_HVT \ram_reg[14][219]  ( .D(n3864), .CLK(clk), .Q(\ram[14][219] ) );
  DFFX1_HVT \ram_reg[14][218]  ( .D(n3863), .CLK(clk), .Q(\ram[14][218] ) );
  DFFX1_HVT \ram_reg[14][217]  ( .D(n3862), .CLK(clk), .Q(\ram[14][217] ) );
  DFFX1_HVT \ram_reg[14][216]  ( .D(n3861), .CLK(clk), .Q(\ram[14][216] ) );
  DFFX1_HVT \ram_reg[14][215]  ( .D(n3860), .CLK(clk), .Q(\ram[14][215] ) );
  DFFX1_HVT \ram_reg[14][214]  ( .D(n3859), .CLK(clk), .Q(\ram[14][214] ) );
  DFFX1_HVT \ram_reg[14][213]  ( .D(n3858), .CLK(clk), .Q(\ram[14][213] ) );
  DFFX1_HVT \ram_reg[14][212]  ( .D(n3857), .CLK(clk), .Q(\ram[14][212] ) );
  DFFX1_HVT \ram_reg[14][211]  ( .D(n3856), .CLK(clk), .Q(\ram[14][211] ) );
  DFFX1_HVT \ram_reg[14][210]  ( .D(n3855), .CLK(clk), .Q(\ram[14][210] ) );
  DFFX1_HVT \ram_reg[14][209]  ( .D(n3854), .CLK(clk), .Q(\ram[14][209] ) );
  DFFX1_HVT \ram_reg[14][208]  ( .D(n3853), .CLK(clk), .Q(\ram[14][208] ) );
  DFFX1_HVT \ram_reg[14][207]  ( .D(n3852), .CLK(clk), .Q(\ram[14][207] ) );
  DFFX1_HVT \ram_reg[14][206]  ( .D(n3851), .CLK(clk), .Q(\ram[14][206] ) );
  DFFX1_HVT \ram_reg[14][205]  ( .D(n3850), .CLK(clk), .Q(\ram[14][205] ) );
  DFFX1_HVT \ram_reg[14][204]  ( .D(n3849), .CLK(clk), .Q(\ram[14][204] ) );
  DFFX1_HVT \ram_reg[14][203]  ( .D(n3848), .CLK(clk), .Q(\ram[14][203] ) );
  DFFX1_HVT \ram_reg[14][202]  ( .D(n3847), .CLK(clk), .Q(\ram[14][202] ) );
  DFFX1_HVT \ram_reg[14][201]  ( .D(n3846), .CLK(clk), .Q(\ram[14][201] ) );
  DFFX1_HVT \ram_reg[14][200]  ( .D(n3845), .CLK(clk), .Q(\ram[14][200] ) );
  DFFX1_HVT \ram_reg[14][199]  ( .D(n3844), .CLK(clk), .Q(\ram[14][199] ) );
  DFFX1_HVT \ram_reg[14][198]  ( .D(n3843), .CLK(clk), .Q(\ram[14][198] ) );
  DFFX1_HVT \ram_reg[14][197]  ( .D(n3842), .CLK(clk), .Q(\ram[14][197] ) );
  DFFX1_HVT \ram_reg[14][196]  ( .D(n3841), .CLK(clk), .Q(\ram[14][196] ) );
  DFFX1_HVT \ram_reg[14][195]  ( .D(n3840), .CLK(clk), .Q(\ram[14][195] ) );
  DFFX1_HVT \ram_reg[14][194]  ( .D(n3839), .CLK(clk), .Q(\ram[14][194] ) );
  DFFX1_HVT \ram_reg[14][193]  ( .D(n3838), .CLK(clk), .Q(\ram[14][193] ) );
  DFFX1_HVT \ram_reg[14][192]  ( .D(n3837), .CLK(clk), .Q(\ram[14][192] ) );
  DFFX1_HVT \ram_reg[14][191]  ( .D(n3836), .CLK(clk), .Q(\ram[14][191] ) );
  DFFX1_HVT \ram_reg[14][190]  ( .D(n3835), .CLK(clk), .Q(\ram[14][190] ) );
  DFFX1_HVT \ram_reg[14][189]  ( .D(n3834), .CLK(clk), .Q(\ram[14][189] ) );
  DFFX1_HVT \ram_reg[14][188]  ( .D(n3833), .CLK(clk), .Q(\ram[14][188] ) );
  DFFX1_HVT \ram_reg[14][187]  ( .D(n3832), .CLK(clk), .Q(\ram[14][187] ) );
  DFFX1_HVT \ram_reg[14][186]  ( .D(n3831), .CLK(clk), .Q(\ram[14][186] ) );
  DFFX1_HVT \ram_reg[14][185]  ( .D(n3830), .CLK(clk), .Q(\ram[14][185] ) );
  DFFX1_HVT \ram_reg[14][184]  ( .D(n3829), .CLK(clk), .Q(\ram[14][184] ) );
  DFFX1_HVT \ram_reg[14][183]  ( .D(n3828), .CLK(clk), .Q(\ram[14][183] ) );
  DFFX1_HVT \ram_reg[14][182]  ( .D(n3827), .CLK(clk), .Q(\ram[14][182] ) );
  DFFX1_HVT \ram_reg[14][181]  ( .D(n3826), .CLK(clk), .Q(\ram[14][181] ) );
  DFFX1_HVT \ram_reg[14][180]  ( .D(n3825), .CLK(clk), .Q(\ram[14][180] ) );
  DFFX1_HVT \ram_reg[14][179]  ( .D(n3824), .CLK(clk), .Q(\ram[14][179] ) );
  DFFX1_HVT \ram_reg[14][178]  ( .D(n3823), .CLK(clk), .Q(\ram[14][178] ) );
  DFFX1_HVT \ram_reg[14][177]  ( .D(n3822), .CLK(clk), .Q(\ram[14][177] ) );
  DFFX1_HVT \ram_reg[14][176]  ( .D(n3821), .CLK(clk), .Q(\ram[14][176] ) );
  DFFX1_HVT \ram_reg[14][175]  ( .D(n3820), .CLK(clk), .Q(\ram[14][175] ) );
  DFFX1_HVT \ram_reg[14][174]  ( .D(n3819), .CLK(clk), .Q(\ram[14][174] ) );
  DFFX1_HVT \ram_reg[14][173]  ( .D(n3818), .CLK(clk), .Q(\ram[14][173] ) );
  DFFX1_HVT \ram_reg[14][172]  ( .D(n3817), .CLK(clk), .Q(\ram[14][172] ) );
  DFFX1_HVT \ram_reg[14][171]  ( .D(n3816), .CLK(clk), .Q(\ram[14][171] ) );
  DFFX1_HVT \ram_reg[14][170]  ( .D(n3815), .CLK(clk), .Q(\ram[14][170] ) );
  DFFX1_HVT \ram_reg[14][169]  ( .D(n3814), .CLK(clk), .Q(\ram[14][169] ) );
  DFFX1_HVT \ram_reg[14][168]  ( .D(n3813), .CLK(clk), .Q(\ram[14][168] ) );
  DFFX1_HVT \ram_reg[14][167]  ( .D(n3812), .CLK(clk), .Q(\ram[14][167] ) );
  DFFX1_HVT \ram_reg[14][166]  ( .D(n3811), .CLK(clk), .Q(\ram[14][166] ) );
  DFFX1_HVT \ram_reg[14][165]  ( .D(n3810), .CLK(clk), .Q(\ram[14][165] ) );
  DFFX1_HVT \ram_reg[14][164]  ( .D(n3809), .CLK(clk), .Q(\ram[14][164] ) );
  DFFX1_HVT \ram_reg[14][163]  ( .D(n3808), .CLK(clk), .Q(\ram[14][163] ) );
  DFFX1_HVT \ram_reg[14][162]  ( .D(n3807), .CLK(clk), .Q(\ram[14][162] ) );
  DFFX1_HVT \ram_reg[14][161]  ( .D(n3806), .CLK(clk), .Q(\ram[14][161] ) );
  DFFX1_HVT \ram_reg[14][160]  ( .D(n3805), .CLK(clk), .Q(\ram[14][160] ) );
  DFFX1_HVT \ram_reg[14][159]  ( .D(n3804), .CLK(clk), .Q(\ram[14][159] ) );
  DFFX1_HVT \ram_reg[14][158]  ( .D(n3803), .CLK(clk), .Q(\ram[14][158] ) );
  DFFX1_HVT \ram_reg[14][157]  ( .D(n3802), .CLK(clk), .Q(\ram[14][157] ) );
  DFFX1_HVT \ram_reg[14][156]  ( .D(n3801), .CLK(clk), .Q(\ram[14][156] ) );
  DFFX1_HVT \ram_reg[14][155]  ( .D(n3800), .CLK(clk), .Q(\ram[14][155] ) );
  DFFX1_HVT \ram_reg[14][154]  ( .D(n3799), .CLK(clk), .Q(\ram[14][154] ) );
  DFFX1_HVT \ram_reg[14][153]  ( .D(n3798), .CLK(clk), .Q(\ram[14][153] ) );
  DFFX1_HVT \ram_reg[14][152]  ( .D(n3797), .CLK(clk), .Q(\ram[14][152] ) );
  DFFX1_HVT \ram_reg[14][151]  ( .D(n3796), .CLK(clk), .Q(\ram[14][151] ) );
  DFFX1_HVT \ram_reg[14][150]  ( .D(n3795), .CLK(clk), .Q(\ram[14][150] ) );
  DFFX1_HVT \ram_reg[14][149]  ( .D(n3794), .CLK(clk), .Q(\ram[14][149] ) );
  DFFX1_HVT \ram_reg[14][148]  ( .D(n3793), .CLK(clk), .Q(\ram[14][148] ) );
  DFFX1_HVT \ram_reg[14][147]  ( .D(n3792), .CLK(clk), .Q(\ram[14][147] ) );
  DFFX1_HVT \ram_reg[14][146]  ( .D(n3791), .CLK(clk), .Q(\ram[14][146] ) );
  DFFX1_HVT \ram_reg[14][145]  ( .D(n3790), .CLK(clk), .Q(\ram[14][145] ) );
  DFFX1_HVT \ram_reg[14][144]  ( .D(n3789), .CLK(clk), .Q(\ram[14][144] ) );
  DFFX1_HVT \ram_reg[14][143]  ( .D(n3788), .CLK(clk), .Q(\ram[14][143] ) );
  DFFX1_HVT \ram_reg[14][142]  ( .D(n3787), .CLK(clk), .Q(\ram[14][142] ) );
  DFFX1_HVT \ram_reg[14][141]  ( .D(n3786), .CLK(clk), .Q(\ram[14][141] ) );
  DFFX1_HVT \ram_reg[14][140]  ( .D(n3785), .CLK(clk), .Q(\ram[14][140] ) );
  DFFX1_HVT \ram_reg[14][139]  ( .D(n3784), .CLK(clk), .Q(\ram[14][139] ) );
  DFFX1_HVT \ram_reg[14][138]  ( .D(n3783), .CLK(clk), .Q(\ram[14][138] ) );
  DFFX1_HVT \ram_reg[14][137]  ( .D(n3782), .CLK(clk), .Q(\ram[14][137] ) );
  DFFX1_HVT \ram_reg[14][136]  ( .D(n3781), .CLK(clk), .Q(\ram[14][136] ) );
  DFFX1_HVT \ram_reg[14][135]  ( .D(n3780), .CLK(clk), .Q(\ram[14][135] ) );
  DFFX1_HVT \ram_reg[14][134]  ( .D(n3779), .CLK(clk), .Q(\ram[14][134] ) );
  DFFX1_HVT \ram_reg[14][133]  ( .D(n3778), .CLK(clk), .Q(\ram[14][133] ) );
  DFFX1_HVT \ram_reg[14][132]  ( .D(n3777), .CLK(clk), .Q(\ram[14][132] ) );
  DFFX1_HVT \ram_reg[14][131]  ( .D(n3776), .CLK(clk), .Q(\ram[14][131] ) );
  DFFX1_HVT \ram_reg[14][130]  ( .D(n3775), .CLK(clk), .Q(\ram[14][130] ) );
  DFFX1_HVT \ram_reg[14][129]  ( .D(n3774), .CLK(clk), .Q(\ram[14][129] ) );
  DFFX1_HVT \ram_reg[14][128]  ( .D(n3773), .CLK(clk), .Q(\ram[14][128] ) );
  DFFX1_HVT \ram_reg[14][127]  ( .D(n3772), .CLK(clk), .Q(\ram[14][127] ) );
  DFFX1_HVT \ram_reg[14][126]  ( .D(n3771), .CLK(clk), .Q(\ram[14][126] ) );
  DFFX1_HVT \ram_reg[14][125]  ( .D(n3770), .CLK(clk), .Q(\ram[14][125] ) );
  DFFX1_HVT \ram_reg[14][124]  ( .D(n3769), .CLK(clk), .Q(\ram[14][124] ) );
  DFFX1_HVT \ram_reg[14][123]  ( .D(n3768), .CLK(clk), .Q(\ram[14][123] ) );
  DFFX1_HVT \ram_reg[14][122]  ( .D(n3767), .CLK(clk), .Q(\ram[14][122] ) );
  DFFX1_HVT \ram_reg[14][121]  ( .D(n3766), .CLK(clk), .Q(\ram[14][121] ) );
  DFFX1_HVT \ram_reg[14][120]  ( .D(n3765), .CLK(clk), .Q(\ram[14][120] ) );
  DFFX1_HVT \ram_reg[14][119]  ( .D(n3764), .CLK(clk), .Q(\ram[14][119] ) );
  DFFX1_HVT \ram_reg[14][118]  ( .D(n3763), .CLK(clk), .Q(\ram[14][118] ) );
  DFFX1_HVT \ram_reg[14][117]  ( .D(n3762), .CLK(clk), .Q(\ram[14][117] ) );
  DFFX1_HVT \ram_reg[14][116]  ( .D(n3761), .CLK(clk), .Q(\ram[14][116] ) );
  DFFX1_HVT \ram_reg[14][115]  ( .D(n3760), .CLK(clk), .Q(\ram[14][115] ) );
  DFFX1_HVT \ram_reg[14][114]  ( .D(n3759), .CLK(clk), .Q(\ram[14][114] ) );
  DFFX1_HVT \ram_reg[14][113]  ( .D(n3758), .CLK(clk), .Q(\ram[14][113] ) );
  DFFX1_HVT \ram_reg[14][112]  ( .D(n3757), .CLK(clk), .Q(\ram[14][112] ) );
  DFFX1_HVT \ram_reg[14][111]  ( .D(n3756), .CLK(clk), .Q(\ram[14][111] ) );
  DFFX1_HVT \ram_reg[14][110]  ( .D(n3755), .CLK(clk), .Q(\ram[14][110] ) );
  DFFX1_HVT \ram_reg[14][109]  ( .D(n3754), .CLK(clk), .Q(\ram[14][109] ) );
  DFFX1_HVT \ram_reg[14][108]  ( .D(n3753), .CLK(clk), .Q(\ram[14][108] ) );
  DFFX1_HVT \ram_reg[14][107]  ( .D(n3752), .CLK(clk), .Q(\ram[14][107] ) );
  DFFX1_HVT \ram_reg[14][106]  ( .D(n3751), .CLK(clk), .Q(\ram[14][106] ) );
  DFFX1_HVT \ram_reg[14][105]  ( .D(n3750), .CLK(clk), .Q(\ram[14][105] ) );
  DFFX1_HVT \ram_reg[14][104]  ( .D(n3749), .CLK(clk), .Q(\ram[14][104] ) );
  DFFX1_HVT \ram_reg[14][103]  ( .D(n3748), .CLK(clk), .Q(\ram[14][103] ), 
        .QN(n5857) );
  DFFX1_HVT \ram_reg[14][102]  ( .D(n3747), .CLK(clk), .Q(\ram[14][102] ), 
        .QN(n4479) );
  DFFX1_HVT \ram_reg[14][101]  ( .D(n3746), .CLK(clk), .Q(\ram[14][101] ), 
        .QN(n4811) );
  DFFX1_HVT \ram_reg[14][100]  ( .D(n3745), .CLK(clk), .Q(\ram[14][100] ) );
  DFFX1_HVT \ram_reg[14][99]  ( .D(n3744), .CLK(clk), .Q(\ram[14][99] ) );
  DFFX1_HVT \ram_reg[14][98]  ( .D(n3743), .CLK(clk), .Q(\ram[14][98] ) );
  DFFX1_HVT \ram_reg[14][97]  ( .D(n3742), .CLK(clk), .Q(\ram[14][97] ) );
  DFFX1_HVT \ram_reg[14][96]  ( .D(n3741), .CLK(clk), .Q(\ram[14][96] ) );
  DFFX1_HVT \ram_reg[14][95]  ( .D(n3740), .CLK(clk), .Q(\ram[14][95] ) );
  DFFX1_HVT \ram_reg[14][94]  ( .D(n3739), .CLK(clk), .Q(\ram[14][94] ) );
  DFFX1_HVT \ram_reg[14][93]  ( .D(n3738), .CLK(clk), .Q(\ram[14][93] ) );
  DFFX1_HVT \ram_reg[14][92]  ( .D(n3737), .CLK(clk), .Q(\ram[14][92] ) );
  DFFX1_HVT \ram_reg[14][91]  ( .D(n3736), .CLK(clk), .Q(\ram[14][91] ) );
  DFFX1_HVT \ram_reg[14][90]  ( .D(n3735), .CLK(clk), .Q(\ram[14][90] ) );
  DFFX1_HVT \ram_reg[14][89]  ( .D(n3734), .CLK(clk), .Q(\ram[14][89] ) );
  DFFX1_HVT \ram_reg[14][88]  ( .D(n3733), .CLK(clk), .Q(\ram[14][88] ) );
  DFFX1_HVT \ram_reg[14][87]  ( .D(n3732), .CLK(clk), .Q(\ram[14][87] ) );
  DFFX1_HVT \ram_reg[14][86]  ( .D(n3731), .CLK(clk), .Q(\ram[14][86] ) );
  DFFX1_HVT \ram_reg[14][85]  ( .D(n3730), .CLK(clk), .Q(\ram[14][85] ) );
  DFFX1_HVT \ram_reg[14][84]  ( .D(n3729), .CLK(clk), .Q(\ram[14][84] ) );
  DFFX1_HVT \ram_reg[14][83]  ( .D(n3728), .CLK(clk), .Q(\ram[14][83] ) );
  DFFX1_HVT \ram_reg[14][82]  ( .D(n3727), .CLK(clk), .Q(\ram[14][82] ) );
  DFFX1_HVT \ram_reg[14][81]  ( .D(n3726), .CLK(clk), .Q(\ram[14][81] ) );
  DFFX1_HVT \ram_reg[14][80]  ( .D(n3725), .CLK(clk), .Q(\ram[14][80] ) );
  DFFX1_HVT \ram_reg[14][79]  ( .D(n3724), .CLK(clk), .Q(\ram[14][79] ) );
  DFFX1_HVT \ram_reg[14][78]  ( .D(n3723), .CLK(clk), .Q(\ram[14][78] ) );
  DFFX1_HVT \ram_reg[14][77]  ( .D(n3722), .CLK(clk), .Q(\ram[14][77] ) );
  DFFX1_HVT \ram_reg[14][76]  ( .D(n3721), .CLK(clk), .Q(\ram[14][76] ) );
  DFFX1_HVT \ram_reg[14][75]  ( .D(n3720), .CLK(clk), .Q(\ram[14][75] ) );
  DFFX1_HVT \ram_reg[14][74]  ( .D(n3719), .CLK(clk), .Q(\ram[14][74] ) );
  DFFX1_HVT \ram_reg[14][73]  ( .D(n3718), .CLK(clk), .Q(\ram[14][73] ) );
  DFFX1_HVT \ram_reg[14][72]  ( .D(n3717), .CLK(clk), .Q(\ram[14][72] ) );
  DFFX1_HVT \ram_reg[14][71]  ( .D(n3716), .CLK(clk), .Q(\ram[14][71] ) );
  DFFX1_HVT \ram_reg[14][70]  ( .D(n3715), .CLK(clk), .Q(\ram[14][70] ) );
  DFFX1_HVT \ram_reg[14][69]  ( .D(n3714), .CLK(clk), .Q(\ram[14][69] ) );
  DFFX1_HVT \ram_reg[14][68]  ( .D(n3713), .CLK(clk), .Q(\ram[14][68] ) );
  DFFX1_HVT \ram_reg[14][67]  ( .D(n3712), .CLK(clk), .Q(\ram[14][67] ), .QN(
        n4618) );
  DFFX1_HVT \ram_reg[14][66]  ( .D(n3711), .CLK(clk), .Q(\ram[14][66] ) );
  DFFX1_HVT \ram_reg[14][65]  ( .D(n3710), .CLK(clk), .Q(\ram[14][65] ) );
  DFFX1_HVT \ram_reg[14][64]  ( .D(n3709), .CLK(clk), .Q(\ram[14][64] ) );
  DFFX1_HVT \ram_reg[14][63]  ( .D(n3708), .CLK(clk), .Q(\ram[14][63] ) );
  DFFX1_HVT \ram_reg[14][62]  ( .D(n3707), .CLK(clk), .Q(\ram[14][62] ) );
  DFFX1_HVT \ram_reg[14][61]  ( .D(n3706), .CLK(clk), .Q(\ram[14][61] ) );
  DFFX1_HVT \ram_reg[14][60]  ( .D(n3705), .CLK(clk), .Q(\ram[14][60] ) );
  DFFX1_HVT \ram_reg[14][59]  ( .D(n3704), .CLK(clk), .Q(\ram[14][59] ) );
  DFFX1_HVT \ram_reg[14][58]  ( .D(n3703), .CLK(clk), .Q(\ram[14][58] ) );
  DFFX1_HVT \ram_reg[14][57]  ( .D(n3702), .CLK(clk), .Q(\ram[14][57] ) );
  DFFX1_HVT \ram_reg[14][56]  ( .D(n3701), .CLK(clk), .Q(\ram[14][56] ) );
  DFFX1_HVT \ram_reg[14][55]  ( .D(n3700), .CLK(clk), .Q(\ram[14][55] ), .QN(
        n4290) );
  DFFX1_HVT \ram_reg[14][54]  ( .D(n3699), .CLK(clk), .Q(\ram[14][54] ) );
  DFFX1_HVT \ram_reg[14][53]  ( .D(n3698), .CLK(clk), .Q(\ram[14][53] ) );
  DFFX1_HVT \ram_reg[14][52]  ( .D(n3697), .CLK(clk), .Q(\ram[14][52] ) );
  DFFX1_HVT \ram_reg[14][51]  ( .D(n3696), .CLK(clk), .Q(\ram[14][51] ) );
  DFFX1_HVT \ram_reg[14][50]  ( .D(n3695), .CLK(clk), .Q(\ram[14][50] ) );
  DFFX1_HVT \ram_reg[14][49]  ( .D(n3694), .CLK(clk), .Q(\ram[14][49] ) );
  DFFX1_HVT \ram_reg[14][48]  ( .D(n3693), .CLK(clk), .Q(\ram[14][48] ), .QN(
        n4288) );
  DFFX1_HVT \ram_reg[14][47]  ( .D(n3692), .CLK(clk), .Q(\ram[14][47] ) );
  DFFX1_HVT \ram_reg[14][46]  ( .D(n3691), .CLK(clk), .Q(\ram[14][46] ) );
  DFFX1_HVT \ram_reg[14][45]  ( .D(n3690), .CLK(clk), .Q(\ram[14][45] ) );
  DFFX1_HVT \ram_reg[14][44]  ( .D(n3689), .CLK(clk), .Q(\ram[14][44] ) );
  DFFX1_HVT \ram_reg[14][43]  ( .D(n3688), .CLK(clk), .Q(\ram[14][43] ) );
  DFFX1_HVT \ram_reg[14][42]  ( .D(n3687), .CLK(clk), .Q(\ram[14][42] ) );
  DFFX1_HVT \ram_reg[14][41]  ( .D(n3686), .CLK(clk), .Q(\ram[14][41] ) );
  DFFX1_HVT \ram_reg[14][40]  ( .D(n3685), .CLK(clk), .Q(\ram[14][40] ) );
  DFFX1_HVT \ram_reg[14][39]  ( .D(n3684), .CLK(clk), .Q(\ram[14][39] ) );
  DFFX1_HVT \ram_reg[14][38]  ( .D(n3683), .CLK(clk), .Q(\ram[14][38] ) );
  DFFX1_HVT \ram_reg[14][37]  ( .D(n3682), .CLK(clk), .Q(\ram[14][37] ) );
  DFFX1_HVT \ram_reg[14][36]  ( .D(n3681), .CLK(clk), .Q(\ram[14][36] ) );
  DFFX1_HVT \ram_reg[14][35]  ( .D(n3680), .CLK(clk), .Q(\ram[14][35] ) );
  DFFX1_HVT \ram_reg[14][34]  ( .D(n3679), .CLK(clk), .Q(\ram[14][34] ) );
  DFFX1_HVT \ram_reg[14][33]  ( .D(n3678), .CLK(clk), .Q(\ram[14][33] ) );
  DFFX1_HVT \ram_reg[14][32]  ( .D(n3677), .CLK(clk), .Q(\ram[14][32] ) );
  DFFX1_HVT \ram_reg[14][31]  ( .D(n3676), .CLK(clk), .Q(\ram[14][31] ) );
  DFFX1_HVT \ram_reg[14][30]  ( .D(n3675), .CLK(clk), .Q(\ram[14][30] ) );
  DFFX1_HVT \ram_reg[14][29]  ( .D(n3674), .CLK(clk), .Q(\ram[14][29] ) );
  DFFX1_HVT \ram_reg[14][28]  ( .D(n3673), .CLK(clk), .Q(\ram[14][28] ) );
  DFFX1_HVT \ram_reg[14][27]  ( .D(n3672), .CLK(clk), .Q(\ram[14][27] ) );
  DFFX1_HVT \ram_reg[14][26]  ( .D(n3671), .CLK(clk), .Q(\ram[14][26] ) );
  DFFX1_HVT \ram_reg[14][25]  ( .D(n3670), .CLK(clk), .Q(\ram[14][25] ) );
  DFFX1_HVT \ram_reg[14][24]  ( .D(n3669), .CLK(clk), .Q(\ram[14][24] ) );
  DFFX1_HVT \ram_reg[14][23]  ( .D(n3668), .CLK(clk), .Q(\ram[14][23] ) );
  DFFX1_HVT \ram_reg[14][22]  ( .D(n3667), .CLK(clk), .Q(\ram[14][22] ) );
  DFFX1_HVT \ram_reg[14][21]  ( .D(n3666), .CLK(clk), .Q(\ram[14][21] ) );
  DFFX1_HVT \ram_reg[14][20]  ( .D(n3665), .CLK(clk), .Q(\ram[14][20] ) );
  DFFX1_HVT \ram_reg[14][19]  ( .D(n3664), .CLK(clk), .Q(\ram[14][19] ) );
  DFFX1_HVT \ram_reg[14][18]  ( .D(n3663), .CLK(clk), .Q(\ram[14][18] ) );
  DFFX1_HVT \ram_reg[14][17]  ( .D(n3662), .CLK(clk), .Q(\ram[14][17] ) );
  DFFX1_HVT \ram_reg[14][16]  ( .D(n3661), .CLK(clk), .Q(\ram[14][16] ) );
  DFFX1_HVT \ram_reg[14][15]  ( .D(n3660), .CLK(clk), .Q(\ram[14][15] ) );
  DFFX1_HVT \ram_reg[14][14]  ( .D(n3659), .CLK(clk), .Q(\ram[14][14] ) );
  DFFX1_HVT \ram_reg[14][13]  ( .D(n3658), .CLK(clk), .Q(\ram[14][13] ) );
  DFFX1_HVT \ram_reg[14][12]  ( .D(n3657), .CLK(clk), .Q(\ram[14][12] ) );
  DFFX1_HVT \ram_reg[14][11]  ( .D(n3656), .CLK(clk), .Q(\ram[14][11] ) );
  DFFX1_HVT \ram_reg[14][10]  ( .D(n3655), .CLK(clk), .Q(\ram[14][10] ) );
  DFFX1_HVT \ram_reg[14][9]  ( .D(n3654), .CLK(clk), .Q(\ram[14][9] ), .QN(
        n4598) );
  DFFX1_HVT \ram_reg[14][8]  ( .D(n3653), .CLK(clk), .Q(\ram[14][8] ) );
  DFFX1_HVT \ram_reg[14][7]  ( .D(n3652), .CLK(clk), .Q(\ram[14][7] ) );
  DFFX1_HVT \ram_reg[14][6]  ( .D(n3651), .CLK(clk), .Q(\ram[14][6] ) );
  DFFX1_HVT \ram_reg[14][5]  ( .D(n3650), .CLK(clk), .Q(\ram[14][5] ) );
  DFFX1_HVT \ram_reg[14][4]  ( .D(n3649), .CLK(clk), .Q(\ram[14][4] ) );
  DFFX1_HVT \ram_reg[14][3]  ( .D(n3648), .CLK(clk), .Q(\ram[14][3] ) );
  DFFX1_HVT \ram_reg[14][2]  ( .D(n3647), .CLK(clk), .Q(\ram[14][2] ) );
  DFFX1_HVT \ram_reg[14][1]  ( .D(n3646), .CLK(clk), .Q(\ram[14][1] ) );
  DFFX1_HVT \ram_reg[14][0]  ( .D(n3645), .CLK(clk), .Q(\ram[14][0] ) );
  DFFX1_HVT \ram_reg[13][255]  ( .D(n3644), .CLK(clk), .Q(\ram[13][255] ) );
  DFFX1_HVT \ram_reg[13][254]  ( .D(n3643), .CLK(clk), .Q(\ram[13][254] ) );
  DFFX1_HVT \ram_reg[13][253]  ( .D(n3642), .CLK(clk), .Q(\ram[13][253] ) );
  DFFX1_HVT \ram_reg[13][252]  ( .D(n3641), .CLK(clk), .Q(\ram[13][252] ), 
        .QN(n4577) );
  DFFX1_HVT \ram_reg[13][251]  ( .D(n3640), .CLK(clk), .Q(\ram[13][251] ) );
  DFFX1_HVT \ram_reg[13][250]  ( .D(n3639), .CLK(clk), .Q(\ram[13][250] ) );
  DFFX1_HVT \ram_reg[13][249]  ( .D(n3638), .CLK(clk), .Q(\ram[13][249] ) );
  DFFX1_HVT \ram_reg[13][248]  ( .D(n3637), .CLK(clk), .Q(\ram[13][248] ) );
  DFFX1_HVT \ram_reg[13][247]  ( .D(n3636), .CLK(clk), .Q(\ram[13][247] ) );
  DFFX1_HVT \ram_reg[13][246]  ( .D(n3635), .CLK(clk), .Q(\ram[13][246] ) );
  DFFX1_HVT \ram_reg[13][245]  ( .D(n3634), .CLK(clk), .Q(\ram[13][245] ) );
  DFFX1_HVT \ram_reg[13][244]  ( .D(n3633), .CLK(clk), .Q(\ram[13][244] ) );
  DFFX1_HVT \ram_reg[13][243]  ( .D(n3632), .CLK(clk), .Q(\ram[13][243] ) );
  DFFX1_HVT \ram_reg[13][242]  ( .D(n3631), .CLK(clk), .Q(\ram[13][242] ) );
  DFFX1_HVT \ram_reg[13][241]  ( .D(n3630), .CLK(clk), .Q(\ram[13][241] ) );
  DFFX1_HVT \ram_reg[13][240]  ( .D(n3629), .CLK(clk), .Q(\ram[13][240] ) );
  DFFX1_HVT \ram_reg[13][239]  ( .D(n3628), .CLK(clk), .Q(\ram[13][239] ) );
  DFFX1_HVT \ram_reg[13][238]  ( .D(n3627), .CLK(clk), .Q(\ram[13][238] ) );
  DFFX1_HVT \ram_reg[13][237]  ( .D(n3626), .CLK(clk), .Q(\ram[13][237] ) );
  DFFX1_HVT \ram_reg[13][236]  ( .D(n3625), .CLK(clk), .Q(\ram[13][236] ) );
  DFFX1_HVT \ram_reg[13][235]  ( .D(n3624), .CLK(clk), .Q(\ram[13][235] ) );
  DFFX1_HVT \ram_reg[13][234]  ( .D(n3623), .CLK(clk), .Q(\ram[13][234] ) );
  DFFX1_HVT \ram_reg[13][233]  ( .D(n3622), .CLK(clk), .Q(\ram[13][233] ) );
  DFFX1_HVT \ram_reg[13][232]  ( .D(n3621), .CLK(clk), .Q(\ram[13][232] ) );
  DFFX1_HVT \ram_reg[13][231]  ( .D(n3620), .CLK(clk), .Q(\ram[13][231] ) );
  DFFX1_HVT \ram_reg[13][230]  ( .D(n3619), .CLK(clk), .Q(\ram[13][230] ) );
  DFFX1_HVT \ram_reg[13][229]  ( .D(n3618), .CLK(clk), .Q(\ram[13][229] ) );
  DFFX1_HVT \ram_reg[13][228]  ( .D(n3617), .CLK(clk), .Q(\ram[13][228] ) );
  DFFX1_HVT \ram_reg[13][227]  ( .D(n3616), .CLK(clk), .Q(\ram[13][227] ) );
  DFFX1_HVT \ram_reg[13][226]  ( .D(n3615), .CLK(clk), .Q(\ram[13][226] ) );
  DFFX1_HVT \ram_reg[13][225]  ( .D(n3614), .CLK(clk), .Q(\ram[13][225] ) );
  DFFX1_HVT \ram_reg[13][224]  ( .D(n3613), .CLK(clk), .Q(\ram[13][224] ) );
  DFFX1_HVT \ram_reg[13][223]  ( .D(n3612), .CLK(clk), .Q(\ram[13][223] ) );
  DFFX1_HVT \ram_reg[13][222]  ( .D(n3611), .CLK(clk), .Q(\ram[13][222] ) );
  DFFX1_HVT \ram_reg[13][221]  ( .D(n3610), .CLK(clk), .Q(\ram[13][221] ) );
  DFFX1_HVT \ram_reg[13][220]  ( .D(n3609), .CLK(clk), .Q(\ram[13][220] ) );
  DFFX1_HVT \ram_reg[13][219]  ( .D(n3608), .CLK(clk), .Q(\ram[13][219] ) );
  DFFX1_HVT \ram_reg[13][218]  ( .D(n3607), .CLK(clk), .Q(\ram[13][218] ), 
        .QN(n4539) );
  DFFX1_HVT \ram_reg[13][217]  ( .D(n3606), .CLK(clk), .Q(\ram[13][217] ) );
  DFFX1_HVT \ram_reg[13][216]  ( .D(n3605), .CLK(clk), .Q(\ram[13][216] ) );
  DFFX1_HVT \ram_reg[13][215]  ( .D(n3604), .CLK(clk), .Q(\ram[13][215] ) );
  DFFX1_HVT \ram_reg[13][214]  ( .D(n3603), .CLK(clk), .Q(\ram[13][214] ) );
  DFFX1_HVT \ram_reg[13][213]  ( .D(n3602), .CLK(clk), .Q(\ram[13][213] ) );
  DFFX1_HVT \ram_reg[13][212]  ( .D(n3601), .CLK(clk), .Q(\ram[13][212] ) );
  DFFX1_HVT \ram_reg[13][211]  ( .D(n3600), .CLK(clk), .Q(\ram[13][211] ) );
  DFFX1_HVT \ram_reg[13][210]  ( .D(n3599), .CLK(clk), .Q(\ram[13][210] ) );
  DFFX1_HVT \ram_reg[13][209]  ( .D(n3598), .CLK(clk), .Q(\ram[13][209] ) );
  DFFX1_HVT \ram_reg[13][208]  ( .D(n3597), .CLK(clk), .Q(\ram[13][208] ) );
  DFFX1_HVT \ram_reg[13][207]  ( .D(n3596), .CLK(clk), .Q(\ram[13][207] ) );
  DFFX1_HVT \ram_reg[13][206]  ( .D(n3595), .CLK(clk), .Q(\ram[13][206] ) );
  DFFX1_HVT \ram_reg[13][205]  ( .D(n3594), .CLK(clk), .Q(\ram[13][205] ) );
  DFFX1_HVT \ram_reg[13][204]  ( .D(n3593), .CLK(clk), .Q(\ram[13][204] ) );
  DFFX1_HVT \ram_reg[13][203]  ( .D(n3592), .CLK(clk), .Q(\ram[13][203] ) );
  DFFX1_HVT \ram_reg[13][202]  ( .D(n3591), .CLK(clk), .Q(\ram[13][202] ) );
  DFFX1_HVT \ram_reg[13][201]  ( .D(n3590), .CLK(clk), .Q(\ram[13][201] ) );
  DFFX1_HVT \ram_reg[13][200]  ( .D(n3589), .CLK(clk), .Q(\ram[13][200] ) );
  DFFX1_HVT \ram_reg[13][199]  ( .D(n3588), .CLK(clk), .Q(\ram[13][199] ) );
  DFFX1_HVT \ram_reg[13][198]  ( .D(n3587), .CLK(clk), .Q(\ram[13][198] ) );
  DFFX1_HVT \ram_reg[13][197]  ( .D(n3586), .CLK(clk), .Q(\ram[13][197] ) );
  DFFX1_HVT \ram_reg[13][196]  ( .D(n3585), .CLK(clk), .Q(\ram[13][196] ) );
  DFFX1_HVT \ram_reg[13][195]  ( .D(n3584), .CLK(clk), .Q(\ram[13][195] ) );
  DFFX1_HVT \ram_reg[13][194]  ( .D(n3583), .CLK(clk), .Q(\ram[13][194] ) );
  DFFX1_HVT \ram_reg[13][193]  ( .D(n3582), .CLK(clk), .Q(\ram[13][193] ) );
  DFFX1_HVT \ram_reg[13][192]  ( .D(n3581), .CLK(clk), .Q(\ram[13][192] ) );
  DFFX1_HVT \ram_reg[13][191]  ( .D(n3580), .CLK(clk), .Q(\ram[13][191] ) );
  DFFX1_HVT \ram_reg[13][190]  ( .D(n3579), .CLK(clk), .Q(\ram[13][190] ) );
  DFFX1_HVT \ram_reg[13][189]  ( .D(n3578), .CLK(clk), .Q(\ram[13][189] ), 
        .QN(n4565) );
  DFFX1_HVT \ram_reg[13][188]  ( .D(n3577), .CLK(clk), .Q(\ram[13][188] ) );
  DFFX1_HVT \ram_reg[13][187]  ( .D(n3576), .CLK(clk), .Q(\ram[13][187] ) );
  DFFX1_HVT \ram_reg[13][186]  ( .D(n3575), .CLK(clk), .Q(\ram[13][186] ) );
  DFFX1_HVT \ram_reg[13][185]  ( .D(n3574), .CLK(clk), .Q(\ram[13][185] ) );
  DFFX1_HVT \ram_reg[13][184]  ( .D(n3573), .CLK(clk), .Q(\ram[13][184] ) );
  DFFX1_HVT \ram_reg[13][183]  ( .D(n3572), .CLK(clk), .Q(\ram[13][183] ) );
  DFFX1_HVT \ram_reg[13][182]  ( .D(n3571), .CLK(clk), .Q(\ram[13][182] ) );
  DFFX1_HVT \ram_reg[13][181]  ( .D(n3570), .CLK(clk), .Q(\ram[13][181] ) );
  DFFX1_HVT \ram_reg[13][180]  ( .D(n3569), .CLK(clk), .Q(\ram[13][180] ) );
  DFFX1_HVT \ram_reg[13][179]  ( .D(n3568), .CLK(clk), .Q(\ram[13][179] ) );
  DFFX1_HVT \ram_reg[13][178]  ( .D(n3567), .CLK(clk), .Q(\ram[13][178] ) );
  DFFX1_HVT \ram_reg[13][177]  ( .D(n3566), .CLK(clk), .Q(\ram[13][177] ) );
  DFFX1_HVT \ram_reg[13][176]  ( .D(n3565), .CLK(clk), .Q(\ram[13][176] ) );
  DFFX1_HVT \ram_reg[13][175]  ( .D(n3564), .CLK(clk), .Q(\ram[13][175] ) );
  DFFX1_HVT \ram_reg[13][174]  ( .D(n3563), .CLK(clk), .Q(\ram[13][174] ) );
  DFFX1_HVT \ram_reg[13][173]  ( .D(n3562), .CLK(clk), .Q(\ram[13][173] ) );
  DFFX1_HVT \ram_reg[13][172]  ( .D(n3561), .CLK(clk), .Q(\ram[13][172] ) );
  DFFX1_HVT \ram_reg[13][171]  ( .D(n3560), .CLK(clk), .Q(\ram[13][171] ) );
  DFFX1_HVT \ram_reg[13][170]  ( .D(n3559), .CLK(clk), .Q(\ram[13][170] ) );
  DFFX1_HVT \ram_reg[13][169]  ( .D(n3558), .CLK(clk), .Q(\ram[13][169] ) );
  DFFX1_HVT \ram_reg[13][168]  ( .D(n3557), .CLK(clk), .Q(\ram[13][168] ) );
  DFFX1_HVT \ram_reg[13][167]  ( .D(n3556), .CLK(clk), .Q(\ram[13][167] ) );
  DFFX1_HVT \ram_reg[13][166]  ( .D(n3555), .CLK(clk), .Q(\ram[13][166] ) );
  DFFX1_HVT \ram_reg[13][165]  ( .D(n3554), .CLK(clk), .Q(\ram[13][165] ) );
  DFFX1_HVT \ram_reg[13][164]  ( .D(n3553), .CLK(clk), .Q(\ram[13][164] ) );
  DFFX1_HVT \ram_reg[13][163]  ( .D(n3552), .CLK(clk), .Q(\ram[13][163] ) );
  DFFX1_HVT \ram_reg[13][162]  ( .D(n3551), .CLK(clk), .Q(\ram[13][162] ) );
  DFFX1_HVT \ram_reg[13][161]  ( .D(n3550), .CLK(clk), .Q(\ram[13][161] ), 
        .QN(n4456) );
  DFFX1_HVT \ram_reg[13][160]  ( .D(n3549), .CLK(clk), .Q(\ram[13][160] ) );
  DFFX1_HVT \ram_reg[13][159]  ( .D(n3548), .CLK(clk), .Q(\ram[13][159] ) );
  DFFX1_HVT \ram_reg[13][158]  ( .D(n3547), .CLK(clk), .Q(\ram[13][158] ) );
  DFFX1_HVT \ram_reg[13][157]  ( .D(n3546), .CLK(clk), .Q(\ram[13][157] ) );
  DFFX1_HVT \ram_reg[13][156]  ( .D(n3545), .CLK(clk), .Q(\ram[13][156] ) );
  DFFX1_HVT \ram_reg[13][155]  ( .D(n3544), .CLK(clk), .Q(\ram[13][155] ) );
  DFFX1_HVT \ram_reg[13][154]  ( .D(n3543), .CLK(clk), .Q(\ram[13][154] ) );
  DFFX1_HVT \ram_reg[13][153]  ( .D(n3542), .CLK(clk), .Q(\ram[13][153] ) );
  DFFX1_HVT \ram_reg[13][152]  ( .D(n3541), .CLK(clk), .Q(\ram[13][152] ) );
  DFFX1_HVT \ram_reg[13][151]  ( .D(n3540), .CLK(clk), .Q(\ram[13][151] ) );
  DFFX1_HVT \ram_reg[13][150]  ( .D(n3539), .CLK(clk), .Q(\ram[13][150] ) );
  DFFX1_HVT \ram_reg[13][149]  ( .D(n3538), .CLK(clk), .Q(\ram[13][149] ) );
  DFFX1_HVT \ram_reg[13][148]  ( .D(n3537), .CLK(clk), .Q(\ram[13][148] ) );
  DFFX1_HVT \ram_reg[13][147]  ( .D(n3536), .CLK(clk), .Q(\ram[13][147] ) );
  DFFX1_HVT \ram_reg[13][146]  ( .D(n3535), .CLK(clk), .Q(\ram[13][146] ) );
  DFFX1_HVT \ram_reg[13][145]  ( .D(n3534), .CLK(clk), .Q(\ram[13][145] ) );
  DFFX1_HVT \ram_reg[13][144]  ( .D(n3533), .CLK(clk), .Q(\ram[13][144] ) );
  DFFX1_HVT \ram_reg[13][143]  ( .D(n3532), .CLK(clk), .Q(\ram[13][143] ) );
  DFFX1_HVT \ram_reg[13][142]  ( .D(n3531), .CLK(clk), .Q(\ram[13][142] ), 
        .QN(n4458) );
  DFFX1_HVT \ram_reg[13][141]  ( .D(n3530), .CLK(clk), .Q(\ram[13][141] ) );
  DFFX1_HVT \ram_reg[13][140]  ( .D(n3529), .CLK(clk), .Q(\ram[13][140] ) );
  DFFX1_HVT \ram_reg[13][139]  ( .D(n3528), .CLK(clk), .Q(\ram[13][139] ) );
  DFFX1_HVT \ram_reg[13][138]  ( .D(n3527), .CLK(clk), .Q(\ram[13][138] ) );
  DFFX1_HVT \ram_reg[13][137]  ( .D(n3526), .CLK(clk), .Q(\ram[13][137] ) );
  DFFX1_HVT \ram_reg[13][136]  ( .D(n3525), .CLK(clk), .Q(\ram[13][136] ), 
        .QN(n5495) );
  DFFX1_HVT \ram_reg[13][135]  ( .D(n3524), .CLK(clk), .Q(\ram[13][135] ) );
  DFFX1_HVT \ram_reg[13][134]  ( .D(n3523), .CLK(clk), .Q(\ram[13][134] ) );
  DFFX1_HVT \ram_reg[13][133]  ( .D(n3522), .CLK(clk), .Q(\ram[13][133] ) );
  DFFX1_HVT \ram_reg[13][132]  ( .D(n3521), .CLK(clk), .Q(\ram[13][132] ) );
  DFFX1_HVT \ram_reg[13][131]  ( .D(n3520), .CLK(clk), .Q(\ram[13][131] ) );
  DFFX1_HVT \ram_reg[13][130]  ( .D(n3519), .CLK(clk), .Q(\ram[13][130] ) );
  DFFX1_HVT \ram_reg[13][129]  ( .D(n3518), .CLK(clk), .Q(\ram[13][129] ) );
  DFFX1_HVT \ram_reg[13][128]  ( .D(n3517), .CLK(clk), .Q(\ram[13][128] ) );
  DFFX1_HVT \ram_reg[13][127]  ( .D(n3516), .CLK(clk), .Q(\ram[13][127] ) );
  DFFX1_HVT \ram_reg[13][126]  ( .D(n3515), .CLK(clk), .Q(\ram[13][126] ) );
  DFFX1_HVT \ram_reg[13][125]  ( .D(n3514), .CLK(clk), .Q(\ram[13][125] ) );
  DFFX1_HVT \ram_reg[13][124]  ( .D(n3513), .CLK(clk), .Q(\ram[13][124] ) );
  DFFX1_HVT \ram_reg[13][123]  ( .D(n3512), .CLK(clk), .Q(\ram[13][123] ) );
  DFFX1_HVT \ram_reg[13][122]  ( .D(n3511), .CLK(clk), .Q(\ram[13][122] ) );
  DFFX1_HVT \ram_reg[13][121]  ( .D(n3510), .CLK(clk), .Q(\ram[13][121] ), 
        .QN(n4421) );
  DFFX1_HVT \ram_reg[13][120]  ( .D(n3509), .CLK(clk), .Q(\ram[13][120] ) );
  DFFX1_HVT \ram_reg[13][119]  ( .D(n3508), .CLK(clk), .Q(\ram[13][119] ) );
  DFFX1_HVT \ram_reg[13][118]  ( .D(n3507), .CLK(clk), .Q(\ram[13][118] ) );
  DFFX1_HVT \ram_reg[13][117]  ( .D(n3506), .CLK(clk), .Q(\ram[13][117] ) );
  DFFX1_HVT \ram_reg[13][116]  ( .D(n3505), .CLK(clk), .Q(\ram[13][116] ) );
  DFFX1_HVT \ram_reg[13][115]  ( .D(n3504), .CLK(clk), .Q(\ram[13][115] ) );
  DFFX1_HVT \ram_reg[13][114]  ( .D(n3503), .CLK(clk), .Q(\ram[13][114] ) );
  DFFX1_HVT \ram_reg[13][113]  ( .D(n3502), .CLK(clk), .Q(\ram[13][113] ) );
  DFFX1_HVT \ram_reg[13][112]  ( .D(n3501), .CLK(clk), .Q(\ram[13][112] ) );
  DFFX1_HVT \ram_reg[13][111]  ( .D(n3500), .CLK(clk), .Q(\ram[13][111] ) );
  DFFX1_HVT \ram_reg[13][110]  ( .D(n3499), .CLK(clk), .Q(\ram[13][110] ) );
  DFFX1_HVT \ram_reg[13][109]  ( .D(n3498), .CLK(clk), .Q(\ram[13][109] ) );
  DFFX1_HVT \ram_reg[13][108]  ( .D(n3497), .CLK(clk), .Q(\ram[13][108] ) );
  DFFX1_HVT \ram_reg[13][107]  ( .D(n3496), .CLK(clk), .Q(\ram[13][107] ) );
  DFFX1_HVT \ram_reg[13][106]  ( .D(n3495), .CLK(clk), .Q(\ram[13][106] ) );
  DFFX1_HVT \ram_reg[13][105]  ( .D(n3494), .CLK(clk), .Q(\ram[13][105] ) );
  DFFX1_HVT \ram_reg[13][104]  ( .D(n3493), .CLK(clk), .Q(\ram[13][104] ) );
  DFFX1_HVT \ram_reg[13][103]  ( .D(n3492), .CLK(clk), .Q(\ram[13][103] ), 
        .QN(n5437) );
  DFFX1_HVT \ram_reg[13][102]  ( .D(n3491), .CLK(clk), .Q(\ram[13][102] ) );
  DFFX1_HVT \ram_reg[13][101]  ( .D(n3490), .CLK(clk), .QN(n4810) );
  DFFX1_HVT \ram_reg[13][100]  ( .D(n3489), .CLK(clk), .Q(\ram[13][100] ) );
  DFFX1_HVT \ram_reg[13][99]  ( .D(n3488), .CLK(clk), .Q(\ram[13][99] ) );
  DFFX1_HVT \ram_reg[13][98]  ( .D(n3487), .CLK(clk), .Q(\ram[13][98] ) );
  DFFX1_HVT \ram_reg[13][97]  ( .D(n3486), .CLK(clk), .Q(\ram[13][97] ) );
  DFFX1_HVT \ram_reg[13][96]  ( .D(n3485), .CLK(clk), .Q(\ram[13][96] ) );
  DFFX1_HVT \ram_reg[13][95]  ( .D(n3484), .CLK(clk), .Q(\ram[13][95] ) );
  DFFX1_HVT \ram_reg[13][94]  ( .D(n3483), .CLK(clk), .Q(\ram[13][94] ) );
  DFFX1_HVT \ram_reg[13][93]  ( .D(n3482), .CLK(clk), .Q(\ram[13][93] ) );
  DFFX1_HVT \ram_reg[13][92]  ( .D(n3481), .CLK(clk), .Q(\ram[13][92] ) );
  DFFX1_HVT \ram_reg[13][91]  ( .D(n3480), .CLK(clk), .Q(\ram[13][91] ) );
  DFFX1_HVT \ram_reg[13][90]  ( .D(n3479), .CLK(clk), .Q(\ram[13][90] ) );
  DFFX1_HVT \ram_reg[13][89]  ( .D(n3478), .CLK(clk), .Q(\ram[13][89] ) );
  DFFX1_HVT \ram_reg[13][88]  ( .D(n3477), .CLK(clk), .Q(\ram[13][88] ) );
  DFFX1_HVT \ram_reg[13][87]  ( .D(n3476), .CLK(clk), .Q(\ram[13][87] ) );
  DFFX1_HVT \ram_reg[13][86]  ( .D(n3475), .CLK(clk), .Q(\ram[13][86] ) );
  DFFX1_HVT \ram_reg[13][85]  ( .D(n3474), .CLK(clk), .Q(\ram[13][85] ) );
  DFFX1_HVT \ram_reg[13][84]  ( .D(n3473), .CLK(clk), .Q(\ram[13][84] ) );
  DFFX1_HVT \ram_reg[13][83]  ( .D(n3472), .CLK(clk), .Q(\ram[13][83] ), .QN(
        n4771) );
  DFFX1_HVT \ram_reg[13][82]  ( .D(n3471), .CLK(clk), .Q(\ram[13][82] ) );
  DFFX1_HVT \ram_reg[13][81]  ( .D(n3470), .CLK(clk), .Q(\ram[13][81] ) );
  DFFX1_HVT \ram_reg[13][80]  ( .D(n3469), .CLK(clk), .Q(\ram[13][80] ) );
  DFFX1_HVT \ram_reg[13][79]  ( .D(n3468), .CLK(clk), .Q(\ram[13][79] ) );
  DFFX1_HVT \ram_reg[13][78]  ( .D(n3467), .CLK(clk), .Q(\ram[13][78] ) );
  DFFX1_HVT \ram_reg[13][77]  ( .D(n3466), .CLK(clk), .Q(\ram[13][77] ), .QN(
        n4679) );
  DFFX1_HVT \ram_reg[13][76]  ( .D(n3465), .CLK(clk), .Q(\ram[13][76] ) );
  DFFX1_HVT \ram_reg[13][75]  ( .D(n3464), .CLK(clk), .Q(\ram[13][75] ), .QN(
        n4827) );
  DFFX1_HVT \ram_reg[13][74]  ( .D(n3463), .CLK(clk), .Q(\ram[13][74] ) );
  DFFX1_HVT \ram_reg[13][73]  ( .D(n3462), .CLK(clk), .Q(\ram[13][73] ) );
  DFFX1_HVT \ram_reg[13][72]  ( .D(n3461), .CLK(clk), .Q(\ram[13][72] ) );
  DFFX1_HVT \ram_reg[13][71]  ( .D(n3460), .CLK(clk), .Q(\ram[13][71] ), .QN(
        n4460) );
  DFFX1_HVT \ram_reg[13][70]  ( .D(n3459), .CLK(clk), .Q(\ram[13][70] ) );
  DFFX1_HVT \ram_reg[13][69]  ( .D(n3458), .CLK(clk), .Q(\ram[13][69] ) );
  DFFX1_HVT \ram_reg[13][68]  ( .D(n3457), .CLK(clk), .Q(\ram[13][68] ), .QN(
        n4769) );
  DFFX1_HVT \ram_reg[13][67]  ( .D(n3456), .CLK(clk), .Q(\ram[13][67] ) );
  DFFX1_HVT \ram_reg[13][66]  ( .D(n3455), .CLK(clk), .Q(\ram[13][66] ) );
  DFFX1_HVT \ram_reg[13][65]  ( .D(n3454), .CLK(clk), .Q(\ram[13][65] ), .QN(
        n4881) );
  DFFX1_HVT \ram_reg[13][64]  ( .D(n3453), .CLK(clk), .Q(\ram[13][64] ) );
  DFFX1_HVT \ram_reg[13][63]  ( .D(n3452), .CLK(clk), .Q(\ram[13][63] ) );
  DFFX1_HVT \ram_reg[13][62]  ( .D(n3451), .CLK(clk), .Q(\ram[13][62] ) );
  DFFX1_HVT \ram_reg[13][61]  ( .D(n3450), .CLK(clk), .Q(\ram[13][61] ), .QN(
        n4486) );
  DFFX1_HVT \ram_reg[13][60]  ( .D(n3449), .CLK(clk), .Q(\ram[13][60] ), .QN(
        n4642) );
  DFFX1_HVT \ram_reg[13][59]  ( .D(n3448), .CLK(clk), .Q(\ram[13][59] ), .QN(
        n4644) );
  DFFX1_HVT \ram_reg[13][58]  ( .D(n3447), .CLK(clk), .Q(\ram[13][58] ) );
  DFFX1_HVT \ram_reg[13][57]  ( .D(n3446), .CLK(clk), .Q(\ram[13][57] ) );
  DFFX1_HVT \ram_reg[13][56]  ( .D(n3445), .CLK(clk), .Q(\ram[13][56] ) );
  DFFX1_HVT \ram_reg[13][55]  ( .D(n3444), .CLK(clk), .Q(\ram[13][55] ) );
  DFFX1_HVT \ram_reg[13][54]  ( .D(n3443), .CLK(clk), .Q(\ram[13][54] ) );
  DFFX1_HVT \ram_reg[13][53]  ( .D(n3442), .CLK(clk), .Q(\ram[13][53] ) );
  DFFX1_HVT \ram_reg[13][52]  ( .D(n3441), .CLK(clk), .Q(\ram[13][52] ) );
  DFFX1_HVT \ram_reg[13][51]  ( .D(n3440), .CLK(clk), .Q(\ram[13][51] ) );
  DFFX1_HVT \ram_reg[13][50]  ( .D(n3439), .CLK(clk), .Q(\ram[13][50] ) );
  DFFX1_HVT \ram_reg[13][49]  ( .D(n3438), .CLK(clk), .Q(\ram[13][49] ) );
  DFFX1_HVT \ram_reg[13][48]  ( .D(n3437), .CLK(clk), .Q(\ram[13][48] ) );
  DFFX1_HVT \ram_reg[13][47]  ( .D(n3436), .CLK(clk), .Q(\ram[13][47] ) );
  DFFX1_HVT \ram_reg[13][46]  ( .D(n3435), .CLK(clk), .Q(\ram[13][46] ) );
  DFFX1_HVT \ram_reg[13][45]  ( .D(n3434), .CLK(clk), .Q(\ram[13][45] ) );
  DFFX1_HVT \ram_reg[13][44]  ( .D(n3433), .CLK(clk), .Q(\ram[13][44] ) );
  DFFX1_HVT \ram_reg[13][43]  ( .D(n3432), .CLK(clk), .Q(\ram[13][43] ) );
  DFFX1_HVT \ram_reg[13][42]  ( .D(n3431), .CLK(clk), .Q(\ram[13][42] ) );
  DFFX1_HVT \ram_reg[13][41]  ( .D(n3430), .CLK(clk), .Q(\ram[13][41] ) );
  DFFX1_HVT \ram_reg[13][40]  ( .D(n3429), .CLK(clk), .Q(\ram[13][40] ) );
  DFFX1_HVT \ram_reg[13][39]  ( .D(n3428), .CLK(clk), .Q(\ram[13][39] ) );
  DFFX1_HVT \ram_reg[13][38]  ( .D(n3427), .CLK(clk), .Q(\ram[13][38] ) );
  DFFX1_HVT \ram_reg[13][37]  ( .D(n3426), .CLK(clk), .Q(\ram[13][37] ) );
  DFFX1_HVT \ram_reg[13][36]  ( .D(n3425), .CLK(clk), .Q(\ram[13][36] ) );
  DFFX1_HVT \ram_reg[13][35]  ( .D(n3424), .CLK(clk), .Q(\ram[13][35] ) );
  DFFX1_HVT \ram_reg[13][34]  ( .D(n3423), .CLK(clk), .Q(\ram[13][34] ) );
  DFFX1_HVT \ram_reg[13][33]  ( .D(n3422), .CLK(clk), .Q(\ram[13][33] ) );
  DFFX1_HVT \ram_reg[13][32]  ( .D(n3421), .CLK(clk), .Q(\ram[13][32] ) );
  DFFX1_HVT \ram_reg[13][31]  ( .D(n3420), .CLK(clk), .Q(\ram[13][31] ) );
  DFFX1_HVT \ram_reg[13][30]  ( .D(n3419), .CLK(clk), .Q(\ram[13][30] ), .QN(
        n4856) );
  DFFX1_HVT \ram_reg[13][29]  ( .D(n3418), .CLK(clk), .Q(\ram[13][29] ) );
  DFFX1_HVT \ram_reg[13][28]  ( .D(n3417), .CLK(clk), .Q(\ram[13][28] ), .QN(
        n4846) );
  DFFX1_HVT \ram_reg[13][27]  ( .D(n3416), .CLK(clk), .Q(\ram[13][27] ), .QN(
        n4784) );
  DFFX1_HVT \ram_reg[13][26]  ( .D(n3415), .CLK(clk), .Q(\ram[13][26] ) );
  DFFX1_HVT \ram_reg[13][25]  ( .D(n3414), .CLK(clk), .Q(\ram[13][25] ) );
  DFFX1_HVT \ram_reg[13][24]  ( .D(n3413), .CLK(clk), .Q(\ram[13][24] ) );
  DFFX1_HVT \ram_reg[13][23]  ( .D(n3412), .CLK(clk), .Q(\ram[13][23] ) );
  DFFX1_HVT \ram_reg[13][22]  ( .D(n3411), .CLK(clk), .Q(\ram[13][22] ) );
  DFFX1_HVT \ram_reg[13][21]  ( .D(n3410), .CLK(clk), .Q(\ram[13][21] ) );
  DFFX1_HVT \ram_reg[13][20]  ( .D(n3409), .CLK(clk), .Q(\ram[13][20] ) );
  DFFX1_HVT \ram_reg[13][19]  ( .D(n3408), .CLK(clk), .Q(\ram[13][19] ) );
  DFFX1_HVT \ram_reg[13][18]  ( .D(n3407), .CLK(clk), .Q(\ram[13][18] ) );
  DFFX1_HVT \ram_reg[13][17]  ( .D(n3406), .CLK(clk), .Q(\ram[13][17] ) );
  DFFX1_HVT \ram_reg[13][16]  ( .D(n3405), .CLK(clk), .Q(\ram[13][16] ) );
  DFFX1_HVT \ram_reg[13][15]  ( .D(n3404), .CLK(clk), .Q(\ram[13][15] ) );
  DFFX1_HVT \ram_reg[13][14]  ( .D(n3403), .CLK(clk), .Q(\ram[13][14] ) );
  DFFX1_HVT \ram_reg[13][13]  ( .D(n3402), .CLK(clk), .Q(\ram[13][13] ) );
  DFFX1_HVT \ram_reg[13][12]  ( .D(n3401), .CLK(clk), .Q(\ram[13][12] ) );
  DFFX1_HVT \ram_reg[13][11]  ( .D(n3400), .CLK(clk), .Q(\ram[13][11] ), .QN(
        n4757) );
  DFFX1_HVT \ram_reg[13][10]  ( .D(n3399), .CLK(clk), .Q(\ram[13][10] ) );
  DFFX1_HVT \ram_reg[13][9]  ( .D(n3398), .CLK(clk), .Q(\ram[13][9] ) );
  DFFX1_HVT \ram_reg[13][8]  ( .D(n3397), .CLK(clk), .Q(\ram[13][8] ) );
  DFFX1_HVT \ram_reg[13][7]  ( .D(n3396), .CLK(clk), .Q(\ram[13][7] ) );
  DFFX1_HVT \ram_reg[13][6]  ( .D(n3395), .CLK(clk), .Q(\ram[13][6] ) );
  DFFX1_HVT \ram_reg[13][5]  ( .D(n3394), .CLK(clk), .Q(\ram[13][5] ) );
  DFFX1_HVT \ram_reg[13][4]  ( .D(n3393), .CLK(clk), .Q(\ram[13][4] ) );
  DFFX1_HVT \ram_reg[13][3]  ( .D(n3392), .CLK(clk), .Q(\ram[13][3] ), .QN(
        n4721) );
  DFFX1_HVT \ram_reg[13][2]  ( .D(n3391), .CLK(clk), .Q(\ram[13][2] ) );
  DFFX1_HVT \ram_reg[13][1]  ( .D(n3390), .CLK(clk), .Q(\ram[13][1] ) );
  DFFX1_HVT \ram_reg[13][0]  ( .D(n3389), .CLK(clk), .Q(\ram[13][0] ) );
  DFFX1_HVT \ram_reg[12][255]  ( .D(n3388), .CLK(clk), .Q(\ram[12][255] ) );
  DFFX1_HVT \ram_reg[12][254]  ( .D(n3387), .CLK(clk), .Q(\ram[12][254] ) );
  DFFX1_HVT \ram_reg[12][253]  ( .D(n3386), .CLK(clk), .Q(\ram[12][253] ) );
  DFFX1_HVT \ram_reg[12][252]  ( .D(n3385), .CLK(clk), .Q(\ram[12][252] ) );
  DFFX1_HVT \ram_reg[12][251]  ( .D(n3384), .CLK(clk), .Q(\ram[12][251] ) );
  DFFX1_HVT \ram_reg[12][250]  ( .D(n3383), .CLK(clk), .Q(\ram[12][250] ) );
  DFFX1_HVT \ram_reg[12][249]  ( .D(n3382), .CLK(clk), .Q(\ram[12][249] ) );
  DFFX1_HVT \ram_reg[12][248]  ( .D(n3381), .CLK(clk), .Q(\ram[12][248] ) );
  DFFX1_HVT \ram_reg[12][247]  ( .D(n3380), .CLK(clk), .Q(\ram[12][247] ) );
  DFFX1_HVT \ram_reg[12][246]  ( .D(n3379), .CLK(clk), .Q(\ram[12][246] ) );
  DFFX1_HVT \ram_reg[12][245]  ( .D(n3378), .CLK(clk), .Q(\ram[12][245] ) );
  DFFX1_HVT \ram_reg[12][244]  ( .D(n3377), .CLK(clk), .Q(\ram[12][244] ) );
  DFFX1_HVT \ram_reg[12][243]  ( .D(n3376), .CLK(clk), .Q(\ram[12][243] ) );
  DFFX1_HVT \ram_reg[12][242]  ( .D(n3375), .CLK(clk), .Q(\ram[12][242] ) );
  DFFX1_HVT \ram_reg[12][241]  ( .D(n3374), .CLK(clk), .Q(\ram[12][241] ) );
  DFFX1_HVT \ram_reg[12][240]  ( .D(n3373), .CLK(clk), .Q(\ram[12][240] ) );
  DFFX1_HVT \ram_reg[12][239]  ( .D(n3372), .CLK(clk), .Q(\ram[12][239] ) );
  DFFX1_HVT \ram_reg[12][238]  ( .D(n3371), .CLK(clk), .Q(\ram[12][238] ) );
  DFFX1_HVT \ram_reg[12][237]  ( .D(n3370), .CLK(clk), .Q(\ram[12][237] ) );
  DFFX1_HVT \ram_reg[12][236]  ( .D(n3369), .CLK(clk), .Q(\ram[12][236] ) );
  DFFX1_HVT \ram_reg[12][235]  ( .D(n3368), .CLK(clk), .Q(\ram[12][235] ) );
  DFFX1_HVT \ram_reg[12][234]  ( .D(n3367), .CLK(clk), .Q(\ram[12][234] ) );
  DFFX1_HVT \ram_reg[12][233]  ( .D(n3366), .CLK(clk), .Q(\ram[12][233] ) );
  DFFX1_HVT \ram_reg[12][232]  ( .D(n3365), .CLK(clk), .Q(\ram[12][232] ) );
  DFFX1_HVT \ram_reg[12][231]  ( .D(n3364), .CLK(clk), .Q(\ram[12][231] ) );
  DFFX1_HVT \ram_reg[12][230]  ( .D(n3363), .CLK(clk), .Q(\ram[12][230] ) );
  DFFX1_HVT \ram_reg[12][229]  ( .D(n3362), .CLK(clk), .Q(\ram[12][229] ) );
  DFFX1_HVT \ram_reg[12][228]  ( .D(n3361), .CLK(clk), .Q(\ram[12][228] ) );
  DFFX1_HVT \ram_reg[12][227]  ( .D(n3360), .CLK(clk), .Q(\ram[12][227] ) );
  DFFX1_HVT \ram_reg[12][226]  ( .D(n3359), .CLK(clk), .Q(\ram[12][226] ) );
  DFFX1_HVT \ram_reg[12][225]  ( .D(n3358), .CLK(clk), .Q(\ram[12][225] ) );
  DFFX1_HVT \ram_reg[12][224]  ( .D(n3357), .CLK(clk), .Q(\ram[12][224] ) );
  DFFX1_HVT \ram_reg[12][223]  ( .D(n3356), .CLK(clk), .Q(\ram[12][223] ) );
  DFFX1_HVT \ram_reg[12][222]  ( .D(n3355), .CLK(clk), .Q(\ram[12][222] ) );
  DFFX1_HVT \ram_reg[12][221]  ( .D(n3354), .CLK(clk), .Q(\ram[12][221] ) );
  DFFX1_HVT \ram_reg[12][220]  ( .D(n3353), .CLK(clk), .Q(\ram[12][220] ) );
  DFFX1_HVT \ram_reg[12][219]  ( .D(n3352), .CLK(clk), .Q(\ram[12][219] ) );
  DFFX1_HVT \ram_reg[12][218]  ( .D(n3351), .CLK(clk), .Q(\ram[12][218] ) );
  DFFX1_HVT \ram_reg[12][217]  ( .D(n3350), .CLK(clk), .Q(\ram[12][217] ) );
  DFFX1_HVT \ram_reg[12][216]  ( .D(n3349), .CLK(clk), .Q(\ram[12][216] ) );
  DFFX1_HVT \ram_reg[12][215]  ( .D(n3348), .CLK(clk), .Q(\ram[12][215] ) );
  DFFX1_HVT \ram_reg[12][214]  ( .D(n3347), .CLK(clk), .Q(\ram[12][214] ) );
  DFFX1_HVT \ram_reg[12][213]  ( .D(n3346), .CLK(clk), .Q(\ram[12][213] ) );
  DFFX1_HVT \ram_reg[12][212]  ( .D(n3345), .CLK(clk), .Q(\ram[12][212] ) );
  DFFX1_HVT \ram_reg[12][211]  ( .D(n3344), .CLK(clk), .Q(\ram[12][211] ) );
  DFFX1_HVT \ram_reg[12][210]  ( .D(n3343), .CLK(clk), .Q(\ram[12][210] ) );
  DFFX1_HVT \ram_reg[12][209]  ( .D(n3342), .CLK(clk), .Q(\ram[12][209] ) );
  DFFX1_HVT \ram_reg[12][208]  ( .D(n3341), .CLK(clk), .Q(\ram[12][208] ) );
  DFFX1_HVT \ram_reg[12][207]  ( .D(n3340), .CLK(clk), .Q(\ram[12][207] ) );
  DFFX1_HVT \ram_reg[12][206]  ( .D(n3339), .CLK(clk), .Q(\ram[12][206] ), 
        .QN(n4620) );
  DFFX1_HVT \ram_reg[12][205]  ( .D(n3338), .CLK(clk), .Q(\ram[12][205] ) );
  DFFX1_HVT \ram_reg[12][204]  ( .D(n3337), .CLK(clk), .Q(\ram[12][204] ) );
  DFFX1_HVT \ram_reg[12][203]  ( .D(n3336), .CLK(clk), .Q(\ram[12][203] ) );
  DFFX1_HVT \ram_reg[12][202]  ( .D(n3335), .CLK(clk), .Q(\ram[12][202] ) );
  DFFX1_HVT \ram_reg[12][201]  ( .D(n3334), .CLK(clk), .Q(\ram[12][201] ) );
  DFFX1_HVT \ram_reg[12][200]  ( .D(n3333), .CLK(clk), .Q(\ram[12][200] ) );
  DFFX1_HVT \ram_reg[12][199]  ( .D(n3332), .CLK(clk), .Q(\ram[12][199] ) );
  DFFX1_HVT \ram_reg[12][198]  ( .D(n3331), .CLK(clk), .Q(\ram[12][198] ) );
  DFFX1_HVT \ram_reg[12][197]  ( .D(n3330), .CLK(clk), .Q(\ram[12][197] ) );
  DFFX1_HVT \ram_reg[12][196]  ( .D(n3329), .CLK(clk), .Q(\ram[12][196] ) );
  DFFX1_HVT \ram_reg[12][195]  ( .D(n3328), .CLK(clk), .Q(\ram[12][195] ) );
  DFFX1_HVT \ram_reg[12][194]  ( .D(n3327), .CLK(clk), .Q(\ram[12][194] ) );
  DFFX1_HVT \ram_reg[12][193]  ( .D(n3326), .CLK(clk), .Q(\ram[12][193] ) );
  DFFX1_HVT \ram_reg[12][192]  ( .D(n3325), .CLK(clk), .Q(\ram[12][192] ) );
  DFFX1_HVT \ram_reg[12][191]  ( .D(n3324), .CLK(clk), .Q(\ram[12][191] ) );
  DFFX1_HVT \ram_reg[12][190]  ( .D(n3323), .CLK(clk), .Q(\ram[12][190] ) );
  DFFX1_HVT \ram_reg[12][189]  ( .D(n3322), .CLK(clk), .Q(\ram[12][189] ) );
  DFFX1_HVT \ram_reg[12][188]  ( .D(n3321), .CLK(clk), .Q(\ram[12][188] ) );
  DFFX1_HVT \ram_reg[12][187]  ( .D(n3320), .CLK(clk), .Q(\ram[12][187] ) );
  DFFX1_HVT \ram_reg[12][186]  ( .D(n3319), .CLK(clk), .Q(\ram[12][186] ) );
  DFFX1_HVT \ram_reg[12][185]  ( .D(n3318), .CLK(clk), .Q(\ram[12][185] ) );
  DFFX1_HVT \ram_reg[12][184]  ( .D(n3317), .CLK(clk), .Q(\ram[12][184] ) );
  DFFX1_HVT \ram_reg[12][183]  ( .D(n3316), .CLK(clk), .Q(\ram[12][183] ) );
  DFFX1_HVT \ram_reg[12][182]  ( .D(n3315), .CLK(clk), .Q(\ram[12][182] ) );
  DFFX1_HVT \ram_reg[12][181]  ( .D(n3314), .CLK(clk), .Q(\ram[12][181] ) );
  DFFX1_HVT \ram_reg[12][180]  ( .D(n3313), .CLK(clk), .Q(\ram[12][180] ) );
  DFFX1_HVT \ram_reg[12][179]  ( .D(n3312), .CLK(clk), .Q(\ram[12][179] ) );
  DFFX1_HVT \ram_reg[12][178]  ( .D(n3311), .CLK(clk), .Q(\ram[12][178] ) );
  DFFX1_HVT \ram_reg[12][177]  ( .D(n3310), .CLK(clk), .Q(\ram[12][177] ) );
  DFFX1_HVT \ram_reg[12][176]  ( .D(n3309), .CLK(clk), .Q(\ram[12][176] ) );
  DFFX1_HVT \ram_reg[12][175]  ( .D(n3308), .CLK(clk), .Q(\ram[12][175] ) );
  DFFX1_HVT \ram_reg[12][174]  ( .D(n3307), .CLK(clk), .Q(\ram[12][174] ) );
  DFFX1_HVT \ram_reg[12][173]  ( .D(n3306), .CLK(clk), .Q(\ram[12][173] ) );
  DFFX1_HVT \ram_reg[12][172]  ( .D(n3305), .CLK(clk), .Q(\ram[12][172] ) );
  DFFX1_HVT \ram_reg[12][171]  ( .D(n3304), .CLK(clk), .Q(\ram[12][171] ), 
        .QN(n4609) );
  DFFX1_HVT \ram_reg[12][170]  ( .D(n3303), .CLK(clk), .Q(\ram[12][170] ) );
  DFFX1_HVT \ram_reg[12][169]  ( .D(n3302), .CLK(clk), .Q(\ram[12][169] ) );
  DFFX1_HVT \ram_reg[12][168]  ( .D(n3301), .CLK(clk), .Q(\ram[12][168] ) );
  DFFX1_HVT \ram_reg[12][167]  ( .D(n3300), .CLK(clk), .Q(\ram[12][167] ) );
  DFFX1_HVT \ram_reg[12][166]  ( .D(n3299), .CLK(clk), .Q(\ram[12][166] ) );
  DFFX1_HVT \ram_reg[12][165]  ( .D(n3298), .CLK(clk), .Q(\ram[12][165] ) );
  DFFX1_HVT \ram_reg[12][164]  ( .D(n3297), .CLK(clk), .Q(\ram[12][164] ) );
  DFFX1_HVT \ram_reg[12][163]  ( .D(n3296), .CLK(clk), .Q(\ram[12][163] ) );
  DFFX1_HVT \ram_reg[12][162]  ( .D(n3295), .CLK(clk), .Q(\ram[12][162] ) );
  DFFX1_HVT \ram_reg[12][161]  ( .D(n3294), .CLK(clk), .Q(\ram[12][161] ) );
  DFFX1_HVT \ram_reg[12][160]  ( .D(n3293), .CLK(clk), .Q(\ram[12][160] ) );
  DFFX1_HVT \ram_reg[12][159]  ( .D(n3292), .CLK(clk), .Q(\ram[12][159] ) );
  DFFX1_HVT \ram_reg[12][158]  ( .D(n3291), .CLK(clk), .Q(\ram[12][158] ) );
  DFFX1_HVT \ram_reg[12][157]  ( .D(n3290), .CLK(clk), .Q(\ram[12][157] ) );
  DFFX1_HVT \ram_reg[12][156]  ( .D(n3289), .CLK(clk), .Q(\ram[12][156] ) );
  DFFX1_HVT \ram_reg[12][155]  ( .D(n3288), .CLK(clk), .Q(\ram[12][155] ) );
  DFFX1_HVT \ram_reg[12][154]  ( .D(n3287), .CLK(clk), .Q(\ram[12][154] ) );
  DFFX1_HVT \ram_reg[12][153]  ( .D(n3286), .CLK(clk), .Q(\ram[12][153] ) );
  DFFX1_HVT \ram_reg[12][152]  ( .D(n3285), .CLK(clk), .Q(\ram[12][152] ) );
  DFFX1_HVT \ram_reg[12][151]  ( .D(n3284), .CLK(clk), .Q(\ram[12][151] ) );
  DFFX1_HVT \ram_reg[12][150]  ( .D(n3283), .CLK(clk), .Q(\ram[12][150] ) );
  DFFX1_HVT \ram_reg[12][149]  ( .D(n3282), .CLK(clk), .Q(\ram[12][149] ) );
  DFFX1_HVT \ram_reg[12][148]  ( .D(n3281), .CLK(clk), .Q(\ram[12][148] ) );
  DFFX1_HVT \ram_reg[12][147]  ( .D(n3280), .CLK(clk), .Q(\ram[12][147] ) );
  DFFX1_HVT \ram_reg[12][146]  ( .D(n3279), .CLK(clk), .Q(\ram[12][146] ) );
  DFFX1_HVT \ram_reg[12][145]  ( .D(n3278), .CLK(clk), .Q(\ram[12][145] ) );
  DFFX1_HVT \ram_reg[12][144]  ( .D(n3277), .CLK(clk), .Q(\ram[12][144] ) );
  DFFX1_HVT \ram_reg[12][143]  ( .D(n3276), .CLK(clk), .Q(\ram[12][143] ), 
        .QN(n4548) );
  DFFX1_HVT \ram_reg[12][142]  ( .D(n3275), .CLK(clk), .Q(\ram[12][142] ) );
  DFFX1_HVT \ram_reg[12][141]  ( .D(n3274), .CLK(clk), .Q(\ram[12][141] ) );
  DFFX1_HVT \ram_reg[12][140]  ( .D(n3273), .CLK(clk), .Q(\ram[12][140] ), 
        .QN(n4284) );
  DFFX1_HVT \ram_reg[12][139]  ( .D(n3272), .CLK(clk), .Q(\ram[12][139] ) );
  DFFX1_HVT \ram_reg[12][138]  ( .D(n3271), .CLK(clk), .Q(\ram[12][138] ) );
  DFFX1_HVT \ram_reg[12][137]  ( .D(n3270), .CLK(clk), .Q(\ram[12][137] ) );
  DFFX1_HVT \ram_reg[12][136]  ( .D(n3269), .CLK(clk), .Q(\ram[12][136] ) );
  DFFX1_HVT \ram_reg[12][135]  ( .D(n3268), .CLK(clk), .Q(\ram[12][135] ) );
  DFFX1_HVT \ram_reg[12][134]  ( .D(n3267), .CLK(clk), .Q(\ram[12][134] ) );
  DFFX1_HVT \ram_reg[12][133]  ( .D(n3266), .CLK(clk), .Q(\ram[12][133] ) );
  DFFX1_HVT \ram_reg[12][132]  ( .D(n3265), .CLK(clk), .Q(\ram[12][132] ) );
  DFFX1_HVT \ram_reg[12][131]  ( .D(n3264), .CLK(clk), .Q(\ram[12][131] ) );
  DFFX1_HVT \ram_reg[12][130]  ( .D(n3263), .CLK(clk), .Q(\ram[12][130] ) );
  DFFX1_HVT \ram_reg[12][129]  ( .D(n3262), .CLK(clk), .Q(\ram[12][129] ) );
  DFFX1_HVT \ram_reg[12][128]  ( .D(n3261), .CLK(clk), .Q(\ram[12][128] ) );
  DFFX1_HVT \ram_reg[12][127]  ( .D(n3260), .CLK(clk), .Q(\ram[12][127] ) );
  DFFX1_HVT \ram_reg[12][126]  ( .D(n3259), .CLK(clk), .Q(\ram[12][126] ) );
  DFFX1_HVT \ram_reg[12][125]  ( .D(n3258), .CLK(clk), .Q(\ram[12][125] ) );
  DFFX1_HVT \ram_reg[12][124]  ( .D(n3257), .CLK(clk), .Q(\ram[12][124] ) );
  DFFX1_HVT \ram_reg[12][123]  ( .D(n3256), .CLK(clk), .Q(\ram[12][123] ) );
  DFFX1_HVT \ram_reg[12][122]  ( .D(n3255), .CLK(clk), .Q(\ram[12][122] ) );
  DFFX1_HVT \ram_reg[12][121]  ( .D(n3254), .CLK(clk), .Q(\ram[12][121] ) );
  DFFX1_HVT \ram_reg[12][120]  ( .D(n3253), .CLK(clk), .Q(\ram[12][120] ) );
  DFFX1_HVT \ram_reg[12][119]  ( .D(n3252), .CLK(clk), .Q(\ram[12][119] ) );
  DFFX1_HVT \ram_reg[12][118]  ( .D(n3251), .CLK(clk), .Q(\ram[12][118] ) );
  DFFX1_HVT \ram_reg[12][117]  ( .D(n3250), .CLK(clk), .Q(\ram[12][117] ) );
  DFFX1_HVT \ram_reg[12][116]  ( .D(n3249), .CLK(clk), .Q(\ram[12][116] ) );
  DFFX1_HVT \ram_reg[12][115]  ( .D(n3248), .CLK(clk), .Q(\ram[12][115] ) );
  DFFX1_HVT \ram_reg[12][114]  ( .D(n3247), .CLK(clk), .Q(\ram[12][114] ) );
  DFFX1_HVT \ram_reg[12][113]  ( .D(n3246), .CLK(clk), .Q(\ram[12][113] ) );
  DFFX1_HVT \ram_reg[12][112]  ( .D(n3245), .CLK(clk), .Q(\ram[12][112] ) );
  DFFX1_HVT \ram_reg[12][111]  ( .D(n3244), .CLK(clk), .Q(\ram[12][111] ) );
  DFFX1_HVT \ram_reg[12][110]  ( .D(n3243), .CLK(clk), .Q(\ram[12][110] ) );
  DFFX1_HVT \ram_reg[12][109]  ( .D(n3242), .CLK(clk), .Q(\ram[12][109] ) );
  DFFX1_HVT \ram_reg[12][108]  ( .D(n3241), .CLK(clk), .Q(\ram[12][108] ) );
  DFFX1_HVT \ram_reg[12][107]  ( .D(n3240), .CLK(clk), .Q(\ram[12][107] ) );
  DFFX1_HVT \ram_reg[12][106]  ( .D(n3239), .CLK(clk), .Q(\ram[12][106] ) );
  DFFX1_HVT \ram_reg[12][105]  ( .D(n3238), .CLK(clk), .Q(\ram[12][105] ) );
  DFFX1_HVT \ram_reg[12][104]  ( .D(n3237), .CLK(clk), .Q(\ram[12][104] ) );
  DFFX1_HVT \ram_reg[12][103]  ( .D(n3236), .CLK(clk), .Q(\ram[12][103] ), 
        .QN(n5858) );
  DFFX1_HVT \ram_reg[12][102]  ( .D(n3235), .CLK(clk), .Q(\ram[12][102] ) );
  DFFX1_HVT \ram_reg[12][101]  ( .D(n3234), .CLK(clk), .Q(\ram[12][101] ), 
        .QN(n4812) );
  DFFX1_HVT \ram_reg[12][100]  ( .D(n3233), .CLK(clk), .Q(\ram[12][100] ) );
  DFFX1_HVT \ram_reg[12][99]  ( .D(n3232), .CLK(clk), .Q(\ram[12][99] ) );
  DFFX1_HVT \ram_reg[12][98]  ( .D(n3231), .CLK(clk), .Q(\ram[12][98] ), .QN(
        n4369) );
  DFFX1_HVT \ram_reg[12][97]  ( .D(n3230), .CLK(clk), .Q(\ram[12][97] ) );
  DFFX1_HVT \ram_reg[12][96]  ( .D(n3229), .CLK(clk), .Q(\ram[12][96] ) );
  DFFX1_HVT \ram_reg[12][95]  ( .D(n3228), .CLK(clk), .Q(\ram[12][95] ) );
  DFFX1_HVT \ram_reg[12][94]  ( .D(n3227), .CLK(clk), .Q(\ram[12][94] ) );
  DFFX1_HVT \ram_reg[12][93]  ( .D(n3226), .CLK(clk), .Q(\ram[12][93] ) );
  DFFX1_HVT \ram_reg[12][92]  ( .D(n3225), .CLK(clk), .Q(\ram[12][92] ) );
  DFFX1_HVT \ram_reg[12][91]  ( .D(n3224), .CLK(clk), .Q(\ram[12][91] ) );
  DFFX1_HVT \ram_reg[12][90]  ( .D(n3223), .CLK(clk), .Q(\ram[12][90] ) );
  DFFX1_HVT \ram_reg[12][89]  ( .D(n3222), .CLK(clk), .Q(\ram[12][89] ) );
  DFFX1_HVT \ram_reg[12][88]  ( .D(n3221), .CLK(clk), .Q(\ram[12][88] ) );
  DFFX1_HVT \ram_reg[12][87]  ( .D(n3220), .CLK(clk), .Q(\ram[12][87] ) );
  DFFX1_HVT \ram_reg[12][86]  ( .D(n3219), .CLK(clk), .Q(\ram[12][86] ) );
  DFFX1_HVT \ram_reg[12][85]  ( .D(n3218), .CLK(clk), .Q(\ram[12][85] ), .QN(
        n4276) );
  DFFX1_HVT \ram_reg[12][84]  ( .D(n3217), .CLK(clk), .Q(\ram[12][84] ) );
  DFFX1_HVT \ram_reg[12][83]  ( .D(n3216), .CLK(clk), .Q(\ram[12][83] ), .QN(
        n4501) );
  DFFX1_HVT \ram_reg[12][82]  ( .D(n3215), .CLK(clk), .Q(\ram[12][82] ) );
  DFFX1_HVT \ram_reg[12][81]  ( .D(n3214), .CLK(clk), .Q(\ram[12][81] ) );
  DFFX1_HVT \ram_reg[12][80]  ( .D(n3213), .CLK(clk), .Q(\ram[12][80] ) );
  DFFX1_HVT \ram_reg[12][79]  ( .D(n3212), .CLK(clk), .Q(\ram[12][79] ) );
  DFFX1_HVT \ram_reg[12][78]  ( .D(n3211), .CLK(clk), .Q(\ram[12][78] ) );
  DFFX1_HVT \ram_reg[12][77]  ( .D(n3210), .CLK(clk), .Q(\ram[12][77] ) );
  DFFX1_HVT \ram_reg[12][76]  ( .D(n3209), .CLK(clk), .Q(\ram[12][76] ) );
  DFFX1_HVT \ram_reg[12][75]  ( .D(n3208), .CLK(clk), .Q(\ram[12][75] ) );
  DFFX1_HVT \ram_reg[12][74]  ( .D(n3207), .CLK(clk), .Q(\ram[12][74] ) );
  DFFX1_HVT \ram_reg[12][73]  ( .D(n3206), .CLK(clk), .Q(\ram[12][73] ) );
  DFFX1_HVT \ram_reg[12][72]  ( .D(n3205), .CLK(clk), .Q(\ram[12][72] ) );
  DFFX1_HVT \ram_reg[12][71]  ( .D(n3204), .CLK(clk), .Q(\ram[12][71] ) );
  DFFX1_HVT \ram_reg[12][70]  ( .D(n3203), .CLK(clk), .Q(\ram[12][70] ) );
  DFFX1_HVT \ram_reg[12][69]  ( .D(n3202), .CLK(clk), .Q(\ram[12][69] ), .QN(
        n4687) );
  DFFX1_HVT \ram_reg[12][68]  ( .D(n3201), .CLK(clk), .Q(\ram[12][68] ) );
  DFFX1_HVT \ram_reg[12][67]  ( .D(n3200), .CLK(clk), .Q(\ram[12][67] ) );
  DFFX1_HVT \ram_reg[12][66]  ( .D(n3199), .CLK(clk), .Q(\ram[12][66] ) );
  DFFX1_HVT \ram_reg[12][65]  ( .D(n3198), .CLK(clk), .Q(\ram[12][65] ), .QN(
        n4880) );
  DFFX1_HVT \ram_reg[12][64]  ( .D(n3197), .CLK(clk), .Q(\ram[12][64] ) );
  DFFX1_HVT \ram_reg[12][63]  ( .D(n3196), .CLK(clk), .Q(\ram[12][63] ) );
  DFFX1_HVT \ram_reg[12][62]  ( .D(n3195), .CLK(clk), .Q(\ram[12][62] ) );
  DFFX1_HVT \ram_reg[12][61]  ( .D(n3194), .CLK(clk), .Q(\ram[12][61] ) );
  DFFX1_HVT \ram_reg[12][60]  ( .D(n3193), .CLK(clk), .Q(\ram[12][60] ) );
  DFFX1_HVT \ram_reg[12][59]  ( .D(n3192), .CLK(clk), .Q(\ram[12][59] ) );
  DFFX1_HVT \ram_reg[12][58]  ( .D(n3191), .CLK(clk), .Q(\ram[12][58] ) );
  DFFX1_HVT \ram_reg[12][57]  ( .D(n3190), .CLK(clk), .Q(\ram[12][57] ) );
  DFFX1_HVT \ram_reg[12][56]  ( .D(n3189), .CLK(clk), .Q(\ram[12][56] ) );
  DFFX1_HVT \ram_reg[12][55]  ( .D(n3188), .CLK(clk), .Q(\ram[12][55] ) );
  DFFX1_HVT \ram_reg[12][54]  ( .D(n3187), .CLK(clk), .Q(\ram[12][54] ) );
  DFFX1_HVT \ram_reg[12][53]  ( .D(n3186), .CLK(clk), .Q(\ram[12][53] ) );
  DFFX1_HVT \ram_reg[12][52]  ( .D(n3185), .CLK(clk), .Q(\ram[12][52] ) );
  DFFX1_HVT \ram_reg[12][51]  ( .D(n3184), .CLK(clk), .Q(\ram[12][51] ) );
  DFFX1_HVT \ram_reg[12][50]  ( .D(n3183), .CLK(clk), .Q(\ram[12][50] ) );
  DFFX1_HVT \ram_reg[12][49]  ( .D(n3182), .CLK(clk), .Q(\ram[12][49] ), .QN(
        n4554) );
  DFFX1_HVT \ram_reg[12][48]  ( .D(n3181), .CLK(clk), .Q(\ram[12][48] ) );
  DFFX1_HVT \ram_reg[12][47]  ( .D(n3180), .CLK(clk), .Q(\ram[12][47] ) );
  DFFX1_HVT \ram_reg[12][46]  ( .D(n3179), .CLK(clk), .Q(\ram[12][46] ) );
  DFFX1_HVT \ram_reg[12][45]  ( .D(n3178), .CLK(clk), .Q(\ram[12][45] ) );
  DFFX1_HVT \ram_reg[12][44]  ( .D(n3177), .CLK(clk), .Q(\ram[12][44] ) );
  DFFX1_HVT \ram_reg[12][43]  ( .D(n3176), .CLK(clk), .Q(\ram[12][43] ) );
  DFFX1_HVT \ram_reg[12][42]  ( .D(n3175), .CLK(clk), .Q(\ram[12][42] ) );
  DFFX1_HVT \ram_reg[12][41]  ( .D(n3174), .CLK(clk), .Q(\ram[12][41] ) );
  DFFX1_HVT \ram_reg[12][40]  ( .D(n3173), .CLK(clk), .Q(\ram[12][40] ) );
  DFFX1_HVT \ram_reg[12][39]  ( .D(n3172), .CLK(clk), .Q(\ram[12][39] ) );
  DFFX1_HVT \ram_reg[12][38]  ( .D(n3171), .CLK(clk), .Q(\ram[12][38] ) );
  DFFX1_HVT \ram_reg[12][37]  ( .D(n3170), .CLK(clk), .Q(\ram[12][37] ) );
  DFFX1_HVT \ram_reg[12][36]  ( .D(n3169), .CLK(clk), .Q(\ram[12][36] ) );
  DFFX1_HVT \ram_reg[12][35]  ( .D(n3168), .CLK(clk), .Q(\ram[12][35] ), .QN(
        n4555) );
  DFFX1_HVT \ram_reg[12][34]  ( .D(n3167), .CLK(clk), .Q(\ram[12][34] ), .QN(
        n4746) );
  DFFX1_HVT \ram_reg[12][33]  ( .D(n3166), .CLK(clk), .Q(\ram[12][33] ) );
  DFFX1_HVT \ram_reg[12][32]  ( .D(n3165), .CLK(clk), .Q(\ram[12][32] ), .QN(
        n4401) );
  DFFX1_HVT \ram_reg[12][31]  ( .D(n3164), .CLK(clk), .Q(\ram[12][31] ) );
  DFFX1_HVT \ram_reg[12][30]  ( .D(n3163), .CLK(clk), .Q(\ram[12][30] ) );
  DFFX1_HVT \ram_reg[12][29]  ( .D(n3162), .CLK(clk), .Q(\ram[12][29] ) );
  DFFX1_HVT \ram_reg[12][28]  ( .D(n3161), .CLK(clk), .Q(\ram[12][28] ), .QN(
        n4404) );
  DFFX1_HVT \ram_reg[12][27]  ( .D(n3160), .CLK(clk), .Q(\ram[12][27] ) );
  DFFX1_HVT \ram_reg[12][26]  ( .D(n3159), .CLK(clk), .Q(\ram[12][26] ) );
  DFFX1_HVT \ram_reg[12][25]  ( .D(n3158), .CLK(clk), .Q(\ram[12][25] ) );
  DFFX1_HVT \ram_reg[12][24]  ( .D(n3157), .CLK(clk), .Q(\ram[12][24] ) );
  DFFX1_HVT \ram_reg[12][23]  ( .D(n3156), .CLK(clk), .Q(\ram[12][23] ) );
  DFFX1_HVT \ram_reg[12][22]  ( .D(n3155), .CLK(clk), .Q(\ram[12][22] ) );
  DFFX1_HVT \ram_reg[12][21]  ( .D(n3154), .CLK(clk), .Q(\ram[12][21] ) );
  DFFX1_HVT \ram_reg[12][20]  ( .D(n3153), .CLK(clk), .Q(\ram[12][20] ) );
  DFFX1_HVT \ram_reg[12][19]  ( .D(n3152), .CLK(clk), .Q(\ram[12][19] ) );
  DFFX1_HVT \ram_reg[12][18]  ( .D(n3151), .CLK(clk), .Q(\ram[12][18] ) );
  DFFX1_HVT \ram_reg[12][17]  ( .D(n3150), .CLK(clk), .Q(\ram[12][17] ) );
  DFFX1_HVT \ram_reg[12][16]  ( .D(n3149), .CLK(clk), .Q(\ram[12][16] ) );
  DFFX1_HVT \ram_reg[12][15]  ( .D(n3148), .CLK(clk), .Q(\ram[12][15] ) );
  DFFX1_HVT \ram_reg[12][14]  ( .D(n3147), .CLK(clk), .Q(\ram[12][14] ), .QN(
        n4277) );
  DFFX1_HVT \ram_reg[12][13]  ( .D(n3146), .CLK(clk), .Q(\ram[12][13] ) );
  DFFX1_HVT \ram_reg[12][12]  ( .D(n3145), .CLK(clk), .Q(\ram[12][12] ) );
  DFFX1_HVT \ram_reg[12][11]  ( .D(n3144), .CLK(clk), .Q(\ram[12][11] ) );
  DFFX1_HVT \ram_reg[12][10]  ( .D(n3143), .CLK(clk), .Q(\ram[12][10] ) );
  DFFX1_HVT \ram_reg[12][9]  ( .D(n3142), .CLK(clk), .Q(\ram[12][9] ) );
  DFFX1_HVT \ram_reg[12][8]  ( .D(n3141), .CLK(clk), .Q(\ram[12][8] ) );
  DFFX1_HVT \ram_reg[12][7]  ( .D(n3140), .CLK(clk), .Q(\ram[12][7] ) );
  DFFX1_HVT \ram_reg[12][6]  ( .D(n3139), .CLK(clk), .Q(\ram[12][6] ) );
  DFFX1_HVT \ram_reg[12][5]  ( .D(n3138), .CLK(clk), .Q(\ram[12][5] ) );
  DFFX1_HVT \ram_reg[12][4]  ( .D(n3137), .CLK(clk), .Q(\ram[12][4] ) );
  DFFX1_HVT \ram_reg[12][3]  ( .D(n3136), .CLK(clk), .Q(\ram[12][3] ) );
  DFFX1_HVT \ram_reg[12][2]  ( .D(n3135), .CLK(clk), .Q(\ram[12][2] ) );
  DFFX1_HVT \ram_reg[12][1]  ( .D(n3134), .CLK(clk), .Q(\ram[12][1] ) );
  DFFX1_HVT \ram_reg[12][0]  ( .D(n3133), .CLK(clk), .Q(\ram[12][0] ) );
  DFFX1_HVT \ram_reg[11][255]  ( .D(n3132), .CLK(clk), .Q(\ram[11][255] ) );
  DFFX1_HVT \ram_reg[11][254]  ( .D(n3131), .CLK(clk), .Q(\ram[11][254] ) );
  DFFX1_HVT \ram_reg[11][253]  ( .D(n3130), .CLK(clk), .Q(\ram[11][253] ) );
  DFFX1_HVT \ram_reg[11][252]  ( .D(n3129), .CLK(clk), .Q(\ram[11][252] ) );
  DFFX1_HVT \ram_reg[11][251]  ( .D(n3128), .CLK(clk), .Q(\ram[11][251] ) );
  DFFX1_HVT \ram_reg[11][250]  ( .D(n3127), .CLK(clk), .Q(\ram[11][250] ) );
  DFFX1_HVT \ram_reg[11][249]  ( .D(n3126), .CLK(clk), .Q(\ram[11][249] ) );
  DFFX1_HVT \ram_reg[11][248]  ( .D(n3125), .CLK(clk), .Q(\ram[11][248] ) );
  DFFX1_HVT \ram_reg[11][247]  ( .D(n3124), .CLK(clk), .Q(\ram[11][247] ) );
  DFFX1_HVT \ram_reg[11][246]  ( .D(n3123), .CLK(clk), .Q(\ram[11][246] ) );
  DFFX1_HVT \ram_reg[11][245]  ( .D(n3122), .CLK(clk), .Q(\ram[11][245] ) );
  DFFX1_HVT \ram_reg[11][244]  ( .D(n3121), .CLK(clk), .Q(\ram[11][244] ) );
  DFFX1_HVT \ram_reg[11][243]  ( .D(n3120), .CLK(clk), .Q(\ram[11][243] ) );
  DFFX1_HVT \ram_reg[11][242]  ( .D(n3119), .CLK(clk), .Q(\ram[11][242] ) );
  DFFX1_HVT \ram_reg[11][241]  ( .D(n3118), .CLK(clk), .Q(\ram[11][241] ) );
  DFFX1_HVT \ram_reg[11][240]  ( .D(n3117), .CLK(clk), .Q(\ram[11][240] ) );
  DFFX1_HVT \ram_reg[11][239]  ( .D(n3116), .CLK(clk), .Q(\ram[11][239] ) );
  DFFX1_HVT \ram_reg[11][238]  ( .D(n3115), .CLK(clk), .Q(\ram[11][238] ) );
  DFFX1_HVT \ram_reg[11][237]  ( .D(n3114), .CLK(clk), .Q(\ram[11][237] ) );
  DFFX1_HVT \ram_reg[11][236]  ( .D(n3113), .CLK(clk), .Q(\ram[11][236] ) );
  DFFX1_HVT \ram_reg[11][235]  ( .D(n3112), .CLK(clk), .Q(\ram[11][235] ) );
  DFFX1_HVT \ram_reg[11][234]  ( .D(n3111), .CLK(clk), .Q(\ram[11][234] ) );
  DFFX1_HVT \ram_reg[11][233]  ( .D(n3110), .CLK(clk), .Q(\ram[11][233] ) );
  DFFX1_HVT \ram_reg[11][232]  ( .D(n3109), .CLK(clk), .Q(\ram[11][232] ) );
  DFFX1_HVT \ram_reg[11][231]  ( .D(n3108), .CLK(clk), .Q(\ram[11][231] ) );
  DFFX1_HVT \ram_reg[11][230]  ( .D(n3107), .CLK(clk), .Q(\ram[11][230] ) );
  DFFX1_HVT \ram_reg[11][229]  ( .D(n3106), .CLK(clk), .Q(\ram[11][229] ) );
  DFFX1_HVT \ram_reg[11][228]  ( .D(n3105), .CLK(clk), .Q(\ram[11][228] ) );
  DFFX1_HVT \ram_reg[11][227]  ( .D(n3104), .CLK(clk), .Q(\ram[11][227] ) );
  DFFX1_HVT \ram_reg[11][226]  ( .D(n3103), .CLK(clk), .Q(\ram[11][226] ) );
  DFFX1_HVT \ram_reg[11][225]  ( .D(n3102), .CLK(clk), .Q(\ram[11][225] ) );
  DFFX1_HVT \ram_reg[11][224]  ( .D(n3101), .CLK(clk), .Q(\ram[11][224] ) );
  DFFX1_HVT \ram_reg[11][223]  ( .D(n3100), .CLK(clk), .Q(\ram[11][223] ) );
  DFFX1_HVT \ram_reg[11][222]  ( .D(n3099), .CLK(clk), .Q(\ram[11][222] ) );
  DFFX1_HVT \ram_reg[11][221]  ( .D(n3098), .CLK(clk), .Q(\ram[11][221] ) );
  DFFX1_HVT \ram_reg[11][220]  ( .D(n3097), .CLK(clk), .Q(\ram[11][220] ), 
        .QN(n5930) );
  DFFX1_HVT \ram_reg[11][219]  ( .D(n3096), .CLK(clk), .Q(\ram[11][219] ) );
  DFFX1_HVT \ram_reg[11][218]  ( .D(n3095), .CLK(clk), .Q(\ram[11][218] ) );
  DFFX1_HVT \ram_reg[11][217]  ( .D(n3094), .CLK(clk), .Q(\ram[11][217] ) );
  DFFX1_HVT \ram_reg[11][216]  ( .D(n3093), .CLK(clk), .Q(\ram[11][216] ) );
  DFFX1_HVT \ram_reg[11][215]  ( .D(n3092), .CLK(clk), .Q(\ram[11][215] ) );
  DFFX1_HVT \ram_reg[11][214]  ( .D(n3091), .CLK(clk), .Q(\ram[11][214] ) );
  DFFX1_HVT \ram_reg[11][213]  ( .D(n3090), .CLK(clk), .Q(\ram[11][213] ) );
  DFFX1_HVT \ram_reg[11][212]  ( .D(n3089), .CLK(clk), .Q(\ram[11][212] ) );
  DFFX1_HVT \ram_reg[11][211]  ( .D(n3088), .CLK(clk), .Q(\ram[11][211] ) );
  DFFX1_HVT \ram_reg[11][210]  ( .D(n3087), .CLK(clk), .Q(\ram[11][210] ) );
  DFFX1_HVT \ram_reg[11][209]  ( .D(n3086), .CLK(clk), .Q(\ram[11][209] ) );
  DFFX1_HVT \ram_reg[11][208]  ( .D(n3085), .CLK(clk), .Q(\ram[11][208] ) );
  DFFX1_HVT \ram_reg[11][207]  ( .D(n3084), .CLK(clk), .Q(\ram[11][207] ) );
  DFFX1_HVT \ram_reg[11][206]  ( .D(n3083), .CLK(clk), .Q(\ram[11][206] ) );
  DFFX1_HVT \ram_reg[11][205]  ( .D(n3082), .CLK(clk), .Q(\ram[11][205] ) );
  DFFX1_HVT \ram_reg[11][204]  ( .D(n3081), .CLK(clk), .Q(\ram[11][204] ) );
  DFFX1_HVT \ram_reg[11][203]  ( .D(n3080), .CLK(clk), .Q(\ram[11][203] ) );
  DFFX1_HVT \ram_reg[11][202]  ( .D(n3079), .CLK(clk), .Q(\ram[11][202] ) );
  DFFX1_HVT \ram_reg[11][201]  ( .D(n3078), .CLK(clk), .Q(\ram[11][201] ) );
  DFFX1_HVT \ram_reg[11][200]  ( .D(n3077), .CLK(clk), .Q(\ram[11][200] ) );
  DFFX1_HVT \ram_reg[11][199]  ( .D(n3076), .CLK(clk), .Q(\ram[11][199] ) );
  DFFX1_HVT \ram_reg[11][198]  ( .D(n3075), .CLK(clk), .Q(\ram[11][198] ) );
  DFFX1_HVT \ram_reg[11][197]  ( .D(n3074), .CLK(clk), .Q(\ram[11][197] ) );
  DFFX1_HVT \ram_reg[11][196]  ( .D(n3073), .CLK(clk), .Q(\ram[11][196] ) );
  DFFX1_HVT \ram_reg[11][195]  ( .D(n3072), .CLK(clk), .Q(\ram[11][195] ) );
  DFFX1_HVT \ram_reg[11][194]  ( .D(n3071), .CLK(clk), .Q(\ram[11][194] ) );
  DFFX1_HVT \ram_reg[11][193]  ( .D(n3070), .CLK(clk), .Q(\ram[11][193] ) );
  DFFX1_HVT \ram_reg[11][192]  ( .D(n3069), .CLK(clk), .Q(\ram[11][192] ) );
  DFFX1_HVT \ram_reg[11][191]  ( .D(n3068), .CLK(clk), .Q(\ram[11][191] ) );
  DFFX1_HVT \ram_reg[11][190]  ( .D(n3067), .CLK(clk), .Q(\ram[11][190] ) );
  DFFX1_HVT \ram_reg[11][189]  ( .D(n3066), .CLK(clk), .Q(\ram[11][189] ) );
  DFFX1_HVT \ram_reg[11][188]  ( .D(n3065), .CLK(clk), .Q(\ram[11][188] ) );
  DFFX1_HVT \ram_reg[11][187]  ( .D(n3064), .CLK(clk), .Q(\ram[11][187] ) );
  DFFX1_HVT \ram_reg[11][186]  ( .D(n3063), .CLK(clk), .Q(\ram[11][186] ) );
  DFFX1_HVT \ram_reg[11][185]  ( .D(n3062), .CLK(clk), .Q(\ram[11][185] ) );
  DFFX1_HVT \ram_reg[11][184]  ( .D(n3061), .CLK(clk), .Q(\ram[11][184] ) );
  DFFX1_HVT \ram_reg[11][183]  ( .D(n3060), .CLK(clk), .Q(\ram[11][183] ) );
  DFFX1_HVT \ram_reg[11][182]  ( .D(n3059), .CLK(clk), .Q(\ram[11][182] ) );
  DFFX1_HVT \ram_reg[11][181]  ( .D(n3058), .CLK(clk), .Q(\ram[11][181] ) );
  DFFX1_HVT \ram_reg[11][180]  ( .D(n3057), .CLK(clk), .Q(\ram[11][180] ) );
  DFFX1_HVT \ram_reg[11][179]  ( .D(n3056), .CLK(clk), .Q(\ram[11][179] ) );
  DFFX1_HVT \ram_reg[11][178]  ( .D(n3055), .CLK(clk), .Q(\ram[11][178] ) );
  DFFX1_HVT \ram_reg[11][177]  ( .D(n3054), .CLK(clk), .Q(\ram[11][177] ) );
  DFFX1_HVT \ram_reg[11][176]  ( .D(n3053), .CLK(clk), .Q(\ram[11][176] ) );
  DFFX1_HVT \ram_reg[11][175]  ( .D(n3052), .CLK(clk), .Q(\ram[11][175] ) );
  DFFX1_HVT \ram_reg[11][174]  ( .D(n3051), .CLK(clk), .Q(\ram[11][174] ) );
  DFFX1_HVT \ram_reg[11][173]  ( .D(n3050), .CLK(clk), .Q(\ram[11][173] ) );
  DFFX1_HVT \ram_reg[11][172]  ( .D(n3049), .CLK(clk), .Q(\ram[11][172] ) );
  DFFX1_HVT \ram_reg[11][171]  ( .D(n3048), .CLK(clk), .Q(\ram[11][171] ) );
  DFFX1_HVT \ram_reg[11][170]  ( .D(n3047), .CLK(clk), .Q(\ram[11][170] ) );
  DFFX1_HVT \ram_reg[11][169]  ( .D(n3046), .CLK(clk), .Q(\ram[11][169] ) );
  DFFX1_HVT \ram_reg[11][168]  ( .D(n3045), .CLK(clk), .Q(\ram[11][168] ) );
  DFFX1_HVT \ram_reg[11][167]  ( .D(n3044), .CLK(clk), .Q(\ram[11][167] ) );
  DFFX1_HVT \ram_reg[11][166]  ( .D(n3043), .CLK(clk), .Q(\ram[11][166] ) );
  DFFX1_HVT \ram_reg[11][165]  ( .D(n3042), .CLK(clk), .Q(\ram[11][165] ) );
  DFFX1_HVT \ram_reg[11][164]  ( .D(n3041), .CLK(clk), .Q(\ram[11][164] ) );
  DFFX1_HVT \ram_reg[11][163]  ( .D(n3040), .CLK(clk), .Q(\ram[11][163] ) );
  DFFX1_HVT \ram_reg[11][162]  ( .D(n3039), .CLK(clk), .Q(\ram[11][162] ), 
        .QN(n4105) );
  DFFX1_HVT \ram_reg[11][161]  ( .D(n3038), .CLK(clk), .Q(\ram[11][161] ) );
  DFFX1_HVT \ram_reg[11][160]  ( .D(n3037), .CLK(clk), .Q(\ram[11][160] ) );
  DFFX1_HVT \ram_reg[11][159]  ( .D(n3036), .CLK(clk), .Q(\ram[11][159] ) );
  DFFX1_HVT \ram_reg[11][158]  ( .D(n3035), .CLK(clk), .Q(\ram[11][158] ) );
  DFFX1_HVT \ram_reg[11][157]  ( .D(n3034), .CLK(clk), .Q(\ram[11][157] ) );
  DFFX1_HVT \ram_reg[11][156]  ( .D(n3033), .CLK(clk), .Q(\ram[11][156] ) );
  DFFX1_HVT \ram_reg[11][155]  ( .D(n3032), .CLK(clk), .Q(\ram[11][155] ) );
  DFFX1_HVT \ram_reg[11][154]  ( .D(n3031), .CLK(clk), .Q(\ram[11][154] ) );
  DFFX1_HVT \ram_reg[11][153]  ( .D(n3030), .CLK(clk), .Q(\ram[11][153] ) );
  DFFX1_HVT \ram_reg[11][152]  ( .D(n3029), .CLK(clk), .Q(\ram[11][152] ) );
  DFFX1_HVT \ram_reg[11][151]  ( .D(n3028), .CLK(clk), .Q(\ram[11][151] ) );
  DFFX1_HVT \ram_reg[11][150]  ( .D(n3027), .CLK(clk), .Q(\ram[11][150] ) );
  DFFX1_HVT \ram_reg[11][149]  ( .D(n3026), .CLK(clk), .Q(\ram[11][149] ) );
  DFFX1_HVT \ram_reg[11][148]  ( .D(n3025), .CLK(clk), .Q(\ram[11][148] ) );
  DFFX1_HVT \ram_reg[11][147]  ( .D(n3024), .CLK(clk), .Q(\ram[11][147] ) );
  DFFX1_HVT \ram_reg[11][146]  ( .D(n3023), .CLK(clk), .Q(\ram[11][146] ) );
  DFFX1_HVT \ram_reg[11][145]  ( .D(n3022), .CLK(clk), .Q(\ram[11][145] ) );
  DFFX1_HVT \ram_reg[11][144]  ( .D(n3021), .CLK(clk), .Q(\ram[11][144] ) );
  DFFX1_HVT \ram_reg[11][143]  ( .D(n3020), .CLK(clk), .Q(\ram[11][143] ) );
  DFFX1_HVT \ram_reg[11][142]  ( .D(n3019), .CLK(clk), .Q(\ram[11][142] ) );
  DFFX1_HVT \ram_reg[11][141]  ( .D(n3018), .CLK(clk), .Q(\ram[11][141] ) );
  DFFX1_HVT \ram_reg[11][140]  ( .D(n3017), .CLK(clk), .Q(\ram[11][140] ) );
  DFFX1_HVT \ram_reg[11][139]  ( .D(n3016), .CLK(clk), .Q(\ram[11][139] ) );
  DFFX1_HVT \ram_reg[11][138]  ( .D(n3015), .CLK(clk), .Q(\ram[11][138] ) );
  DFFX1_HVT \ram_reg[11][137]  ( .D(n3014), .CLK(clk), .Q(\ram[11][137] ) );
  DFFX1_HVT \ram_reg[11][136]  ( .D(n3013), .CLK(clk), .Q(\ram[11][136] ) );
  DFFX1_HVT \ram_reg[11][135]  ( .D(n3012), .CLK(clk), .Q(\ram[11][135] ) );
  DFFX1_HVT \ram_reg[11][134]  ( .D(n3011), .CLK(clk), .Q(\ram[11][134] ) );
  DFFX1_HVT \ram_reg[11][133]  ( .D(n3010), .CLK(clk), .Q(\ram[11][133] ) );
  DFFX1_HVT \ram_reg[11][132]  ( .D(n3009), .CLK(clk), .Q(\ram[11][132] ) );
  DFFX1_HVT \ram_reg[11][131]  ( .D(n3008), .CLK(clk), .Q(\ram[11][131] ) );
  DFFX1_HVT \ram_reg[11][130]  ( .D(n3007), .CLK(clk), .Q(\ram[11][130] ) );
  DFFX1_HVT \ram_reg[11][129]  ( .D(n3006), .CLK(clk), .Q(\ram[11][129] ) );
  DFFX1_HVT \ram_reg[11][128]  ( .D(n3005), .CLK(clk), .Q(\ram[11][128] ) );
  DFFX1_HVT \ram_reg[11][127]  ( .D(n3004), .CLK(clk), .Q(\ram[11][127] ) );
  DFFX1_HVT \ram_reg[11][126]  ( .D(n3003), .CLK(clk), .Q(\ram[11][126] ) );
  DFFX1_HVT \ram_reg[11][125]  ( .D(n3002), .CLK(clk), .Q(\ram[11][125] ) );
  DFFX1_HVT \ram_reg[11][124]  ( .D(n3001), .CLK(clk), .Q(\ram[11][124] ) );
  DFFX1_HVT \ram_reg[11][123]  ( .D(n3000), .CLK(clk), .Q(\ram[11][123] ) );
  DFFX1_HVT \ram_reg[11][122]  ( .D(n2999), .CLK(clk), .Q(\ram[11][122] ) );
  DFFX1_HVT \ram_reg[11][121]  ( .D(n2998), .CLK(clk), .Q(\ram[11][121] ) );
  DFFX1_HVT \ram_reg[11][120]  ( .D(n2997), .CLK(clk), .Q(\ram[11][120] ) );
  DFFX1_HVT \ram_reg[11][119]  ( .D(n2996), .CLK(clk), .Q(\ram[11][119] ) );
  DFFX1_HVT \ram_reg[11][118]  ( .D(n2995), .CLK(clk), .Q(\ram[11][118] ) );
  DFFX1_HVT \ram_reg[11][117]  ( .D(n2994), .CLK(clk), .Q(\ram[11][117] ) );
  DFFX1_HVT \ram_reg[11][116]  ( .D(n2993), .CLK(clk), .Q(\ram[11][116] ) );
  DFFX1_HVT \ram_reg[11][115]  ( .D(n2992), .CLK(clk), .Q(\ram[11][115] ) );
  DFFX1_HVT \ram_reg[11][114]  ( .D(n2991), .CLK(clk), .Q(\ram[11][114] ) );
  DFFX1_HVT \ram_reg[11][113]  ( .D(n2990), .CLK(clk), .Q(\ram[11][113] ) );
  DFFX1_HVT \ram_reg[11][112]  ( .D(n2989), .CLK(clk), .Q(\ram[11][112] ) );
  DFFX1_HVT \ram_reg[11][111]  ( .D(n2988), .CLK(clk), .Q(\ram[11][111] ) );
  DFFX1_HVT \ram_reg[11][110]  ( .D(n2987), .CLK(clk), .Q(\ram[11][110] ) );
  DFFX1_HVT \ram_reg[11][109]  ( .D(n2986), .CLK(clk), .Q(\ram[11][109] ) );
  DFFX1_HVT \ram_reg[11][108]  ( .D(n2985), .CLK(clk), .Q(\ram[11][108] ) );
  DFFX1_HVT \ram_reg[11][107]  ( .D(n2984), .CLK(clk), .Q(\ram[11][107] ) );
  DFFX1_HVT \ram_reg[11][106]  ( .D(n2983), .CLK(clk), .Q(\ram[11][106] ) );
  DFFX1_HVT \ram_reg[11][105]  ( .D(n2982), .CLK(clk), .Q(\ram[11][105] ) );
  DFFX1_HVT \ram_reg[11][104]  ( .D(n2981), .CLK(clk), .Q(\ram[11][104] ) );
  DFFX1_HVT \ram_reg[11][103]  ( .D(n2980), .CLK(clk), .Q(\ram[11][103] ) );
  DFFX1_HVT \ram_reg[11][102]  ( .D(n2979), .CLK(clk), .Q(\ram[11][102] ) );
  DFFX1_HVT \ram_reg[11][101]  ( .D(n2978), .CLK(clk), .Q(\ram[11][101] ) );
  DFFX1_HVT \ram_reg[11][100]  ( .D(n2977), .CLK(clk), .Q(\ram[11][100] ) );
  DFFX1_HVT \ram_reg[11][99]  ( .D(n2976), .CLK(clk), .Q(\ram[11][99] ) );
  DFFX1_HVT \ram_reg[11][98]  ( .D(n2975), .CLK(clk), .Q(\ram[11][98] ) );
  DFFX1_HVT \ram_reg[11][97]  ( .D(n2974), .CLK(clk), .Q(\ram[11][97] ) );
  DFFX1_HVT \ram_reg[11][96]  ( .D(n2973), .CLK(clk), .Q(\ram[11][96] ) );
  DFFX1_HVT \ram_reg[11][95]  ( .D(n2972), .CLK(clk), .Q(\ram[11][95] ) );
  DFFX1_HVT \ram_reg[11][94]  ( .D(n2971), .CLK(clk), .Q(\ram[11][94] ) );
  DFFX1_HVT \ram_reg[11][93]  ( .D(n2970), .CLK(clk), .Q(\ram[11][93] ) );
  DFFX1_HVT \ram_reg[11][92]  ( .D(n2969), .CLK(clk), .Q(\ram[11][92] ) );
  DFFX1_HVT \ram_reg[11][91]  ( .D(n2968), .CLK(clk), .Q(\ram[11][91] ) );
  DFFX1_HVT \ram_reg[11][90]  ( .D(n2967), .CLK(clk), .Q(\ram[11][90] ) );
  DFFX1_HVT \ram_reg[11][89]  ( .D(n2966), .CLK(clk), .Q(\ram[11][89] ) );
  DFFX1_HVT \ram_reg[11][88]  ( .D(n2965), .CLK(clk), .Q(\ram[11][88] ) );
  DFFX1_HVT \ram_reg[11][87]  ( .D(n2964), .CLK(clk), .Q(\ram[11][87] ) );
  DFFX1_HVT \ram_reg[11][86]  ( .D(n2963), .CLK(clk), .Q(\ram[11][86] ) );
  DFFX1_HVT \ram_reg[11][85]  ( .D(n2962), .CLK(clk), .Q(\ram[11][85] ) );
  DFFX1_HVT \ram_reg[11][84]  ( .D(n2961), .CLK(clk), .Q(\ram[11][84] ) );
  DFFX1_HVT \ram_reg[11][83]  ( .D(n2960), .CLK(clk), .Q(\ram[11][83] ) );
  DFFX1_HVT \ram_reg[11][82]  ( .D(n2959), .CLK(clk), .Q(\ram[11][82] ) );
  DFFX1_HVT \ram_reg[11][81]  ( .D(n2958), .CLK(clk), .Q(\ram[11][81] ) );
  DFFX1_HVT \ram_reg[11][80]  ( .D(n2957), .CLK(clk), .Q(\ram[11][80] ) );
  DFFX1_HVT \ram_reg[11][79]  ( .D(n2956), .CLK(clk), .Q(\ram[11][79] ) );
  DFFX1_HVT \ram_reg[11][78]  ( .D(n2955), .CLK(clk), .Q(\ram[11][78] ) );
  DFFX1_HVT \ram_reg[11][77]  ( .D(n2954), .CLK(clk), .Q(\ram[11][77] ) );
  DFFX1_HVT \ram_reg[11][76]  ( .D(n2953), .CLK(clk), .Q(\ram[11][76] ) );
  DFFX1_HVT \ram_reg[11][75]  ( .D(n2952), .CLK(clk), .Q(\ram[11][75] ) );
  DFFX1_HVT \ram_reg[11][74]  ( .D(n2951), .CLK(clk), .Q(\ram[11][74] ) );
  DFFX1_HVT \ram_reg[11][73]  ( .D(n2950), .CLK(clk), .Q(\ram[11][73] ) );
  DFFX1_HVT \ram_reg[11][72]  ( .D(n2949), .CLK(clk), .Q(\ram[11][72] ) );
  DFFX1_HVT \ram_reg[11][71]  ( .D(n2948), .CLK(clk), .Q(\ram[11][71] ) );
  DFFX1_HVT \ram_reg[11][70]  ( .D(n2947), .CLK(clk), .Q(\ram[11][70] ) );
  DFFX1_HVT \ram_reg[11][69]  ( .D(n2946), .CLK(clk), .Q(\ram[11][69] ) );
  DFFX1_HVT \ram_reg[11][68]  ( .D(n2945), .CLK(clk), .Q(\ram[11][68] ) );
  DFFX1_HVT \ram_reg[11][67]  ( .D(n2944), .CLK(clk), .Q(\ram[11][67] ) );
  DFFX1_HVT \ram_reg[11][66]  ( .D(n2943), .CLK(clk), .Q(\ram[11][66] ) );
  DFFX1_HVT \ram_reg[11][65]  ( .D(n2942), .CLK(clk), .Q(\ram[11][65] ) );
  DFFX1_HVT \ram_reg[11][64]  ( .D(n2941), .CLK(clk), .Q(\ram[11][64] ) );
  DFFX1_HVT \ram_reg[11][63]  ( .D(n2940), .CLK(clk), .Q(\ram[11][63] ) );
  DFFX1_HVT \ram_reg[11][62]  ( .D(n2939), .CLK(clk), .Q(\ram[11][62] ) );
  DFFX1_HVT \ram_reg[11][61]  ( .D(n2938), .CLK(clk), .Q(\ram[11][61] ) );
  DFFX1_HVT \ram_reg[11][60]  ( .D(n2937), .CLK(clk), .Q(\ram[11][60] ) );
  DFFX1_HVT \ram_reg[11][59]  ( .D(n2936), .CLK(clk), .Q(\ram[11][59] ) );
  DFFX1_HVT \ram_reg[11][58]  ( .D(n2935), .CLK(clk), .Q(\ram[11][58] ), .QN(
        n4815) );
  DFFX1_HVT \ram_reg[11][57]  ( .D(n2934), .CLK(clk), .Q(\ram[11][57] ) );
  DFFX1_HVT \ram_reg[11][56]  ( .D(n2933), .CLK(clk), .Q(\ram[11][56] ) );
  DFFX1_HVT \ram_reg[11][55]  ( .D(n2932), .CLK(clk), .Q(\ram[11][55] ) );
  DFFX1_HVT \ram_reg[11][54]  ( .D(n2931), .CLK(clk), .Q(\ram[11][54] ) );
  DFFX1_HVT \ram_reg[11][53]  ( .D(n2930), .CLK(clk), .Q(\ram[11][53] ) );
  DFFX1_HVT \ram_reg[11][52]  ( .D(n2929), .CLK(clk), .Q(\ram[11][52] ) );
  DFFX1_HVT \ram_reg[11][51]  ( .D(n2928), .CLK(clk), .Q(\ram[11][51] ) );
  DFFX1_HVT \ram_reg[11][50]  ( .D(n2927), .CLK(clk), .Q(\ram[11][50] ) );
  DFFX1_HVT \ram_reg[11][49]  ( .D(n2926), .CLK(clk), .Q(\ram[11][49] ) );
  DFFX1_HVT \ram_reg[11][48]  ( .D(n2925), .CLK(clk), .Q(\ram[11][48] ) );
  DFFX1_HVT \ram_reg[11][47]  ( .D(n2924), .CLK(clk), .Q(\ram[11][47] ) );
  DFFX1_HVT \ram_reg[11][46]  ( .D(n2923), .CLK(clk), .Q(\ram[11][46] ) );
  DFFX1_HVT \ram_reg[11][45]  ( .D(n2922), .CLK(clk), .Q(\ram[11][45] ) );
  DFFX1_HVT \ram_reg[11][44]  ( .D(n2921), .CLK(clk), .Q(\ram[11][44] ) );
  DFFX1_HVT \ram_reg[11][43]  ( .D(n2920), .CLK(clk), .Q(\ram[11][43] ) );
  DFFX1_HVT \ram_reg[11][42]  ( .D(n2919), .CLK(clk), .Q(\ram[11][42] ) );
  DFFX1_HVT \ram_reg[11][41]  ( .D(n2918), .CLK(clk), .Q(\ram[11][41] ) );
  DFFX1_HVT \ram_reg[11][40]  ( .D(n2917), .CLK(clk), .Q(\ram[11][40] ) );
  DFFX1_HVT \ram_reg[11][39]  ( .D(n2916), .CLK(clk), .Q(\ram[11][39] ) );
  DFFX1_HVT \ram_reg[11][38]  ( .D(n2915), .CLK(clk), .Q(\ram[11][38] ), .QN(
        n1359) );
  DFFX1_HVT \ram_reg[11][37]  ( .D(n2914), .CLK(clk), .Q(\ram[11][37] ) );
  DFFX1_HVT \ram_reg[11][36]  ( .D(n2913), .CLK(clk), .Q(\ram[11][36] ) );
  DFFX1_HVT \ram_reg[11][35]  ( .D(n2912), .CLK(clk), .Q(\ram[11][35] ) );
  DFFX1_HVT \ram_reg[11][34]  ( .D(n2911), .CLK(clk), .Q(\ram[11][34] ) );
  DFFX1_HVT \ram_reg[11][33]  ( .D(n2910), .CLK(clk), .Q(\ram[11][33] ), .QN(
        n4388) );
  DFFX1_HVT \ram_reg[11][32]  ( .D(n2909), .CLK(clk), .Q(\ram[11][32] ), .QN(
        n4391) );
  DFFX1_HVT \ram_reg[11][31]  ( .D(n2908), .CLK(clk), .Q(\ram[11][31] ), .QN(
        n4394) );
  DFFX1_HVT \ram_reg[11][30]  ( .D(n2907), .CLK(clk), .Q(\ram[11][30] ) );
  DFFX1_HVT \ram_reg[11][29]  ( .D(n2906), .CLK(clk), .Q(\ram[11][29] ), .QN(
        n4904) );
  DFFX1_HVT \ram_reg[11][28]  ( .D(n2905), .CLK(clk), .Q(\ram[11][28] ) );
  DFFX1_HVT \ram_reg[11][27]  ( .D(n2904), .CLK(clk), .Q(\ram[11][27] ) );
  DFFX1_HVT \ram_reg[11][26]  ( .D(n2903), .CLK(clk), .Q(\ram[11][26] ) );
  DFFX1_HVT \ram_reg[11][25]  ( .D(n2902), .CLK(clk), .Q(\ram[11][25] ) );
  DFFX1_HVT \ram_reg[11][24]  ( .D(n2901), .CLK(clk), .Q(\ram[11][24] ) );
  DFFX1_HVT \ram_reg[11][23]  ( .D(n2900), .CLK(clk), .Q(\ram[11][23] ) );
  DFFX1_HVT \ram_reg[11][22]  ( .D(n2899), .CLK(clk), .Q(\ram[11][22] ) );
  DFFX1_HVT \ram_reg[11][21]  ( .D(n2898), .CLK(clk), .Q(\ram[11][21] ) );
  DFFX1_HVT \ram_reg[11][20]  ( .D(n2897), .CLK(clk), .Q(\ram[11][20] ), .QN(
        n6481) );
  DFFX1_HVT \ram_reg[11][19]  ( .D(n2896), .CLK(clk), .Q(\ram[11][19] ) );
  DFFX1_HVT \ram_reg[11][18]  ( .D(n2895), .CLK(clk), .Q(\ram[11][18] ) );
  DFFX1_HVT \ram_reg[11][17]  ( .D(n2894), .CLK(clk), .Q(\ram[11][17] ) );
  DFFX1_HVT \ram_reg[11][16]  ( .D(n2893), .CLK(clk), .Q(\ram[11][16] ) );
  DFFX1_HVT \ram_reg[11][15]  ( .D(n2892), .CLK(clk), .Q(\ram[11][15] ) );
  DFFX1_HVT \ram_reg[11][14]  ( .D(n2891), .CLK(clk), .Q(\ram[11][14] ) );
  DFFX1_HVT \ram_reg[11][13]  ( .D(n2890), .CLK(clk), .Q(\ram[11][13] ) );
  DFFX1_HVT \ram_reg[11][12]  ( .D(n2889), .CLK(clk), .Q(\ram[11][12] ) );
  DFFX1_HVT \ram_reg[11][11]  ( .D(n2888), .CLK(clk), .Q(\ram[11][11] ) );
  DFFX1_HVT \ram_reg[11][10]  ( .D(n2887), .CLK(clk), .Q(\ram[11][10] ) );
  DFFX1_HVT \ram_reg[11][9]  ( .D(n2886), .CLK(clk), .Q(\ram[11][9] ) );
  DFFX1_HVT \ram_reg[11][8]  ( .D(n2885), .CLK(clk), .Q(\ram[11][8] ) );
  DFFX1_HVT \ram_reg[11][7]  ( .D(n2884), .CLK(clk), .Q(\ram[11][7] ), .QN(
        n4429) );
  DFFX1_HVT \ram_reg[11][6]  ( .D(n2883), .CLK(clk), .Q(\ram[11][6] ) );
  DFFX1_HVT \ram_reg[11][5]  ( .D(n2882), .CLK(clk), .Q(\ram[11][5] ) );
  DFFX1_HVT \ram_reg[11][4]  ( .D(n2881), .CLK(clk), .Q(\ram[11][4] ) );
  DFFX1_HVT \ram_reg[11][3]  ( .D(n2880), .CLK(clk), .Q(\ram[11][3] ) );
  DFFX1_HVT \ram_reg[11][2]  ( .D(n2879), .CLK(clk), .Q(\ram[11][2] ) );
  DFFX1_HVT \ram_reg[11][1]  ( .D(n2878), .CLK(clk), .Q(\ram[11][1] ) );
  DFFX1_HVT \ram_reg[11][0]  ( .D(n2877), .CLK(clk), .Q(\ram[11][0] ) );
  DFFX1_HVT \ram_reg[10][255]  ( .D(n2876), .CLK(clk), .Q(\ram[10][255] ) );
  DFFX1_HVT \ram_reg[10][254]  ( .D(n2875), .CLK(clk), .Q(\ram[10][254] ) );
  DFFX1_HVT \ram_reg[10][253]  ( .D(n2874), .CLK(clk), .Q(\ram[10][253] ) );
  DFFX1_HVT \ram_reg[10][252]  ( .D(n2873), .CLK(clk), .Q(\ram[10][252] ) );
  DFFX1_HVT \ram_reg[10][251]  ( .D(n2872), .CLK(clk), .Q(\ram[10][251] ) );
  DFFX1_HVT \ram_reg[10][250]  ( .D(n2871), .CLK(clk), .Q(\ram[10][250] ) );
  DFFX1_HVT \ram_reg[10][249]  ( .D(n2870), .CLK(clk), .Q(\ram[10][249] ) );
  DFFX1_HVT \ram_reg[10][248]  ( .D(n2869), .CLK(clk), .Q(\ram[10][248] ) );
  DFFX1_HVT \ram_reg[10][247]  ( .D(n2868), .CLK(clk), .Q(\ram[10][247] ) );
  DFFX1_HVT \ram_reg[10][246]  ( .D(n2867), .CLK(clk), .Q(\ram[10][246] ) );
  DFFX1_HVT \ram_reg[10][245]  ( .D(n2866), .CLK(clk), .Q(\ram[10][245] ) );
  DFFX1_HVT \ram_reg[10][244]  ( .D(n2865), .CLK(clk), .Q(\ram[10][244] ) );
  DFFX1_HVT \ram_reg[10][243]  ( .D(n2864), .CLK(clk), .Q(\ram[10][243] ) );
  DFFX1_HVT \ram_reg[10][242]  ( .D(n2863), .CLK(clk), .Q(\ram[10][242] ) );
  DFFX1_HVT \ram_reg[10][241]  ( .D(n2862), .CLK(clk), .Q(\ram[10][241] ) );
  DFFX1_HVT \ram_reg[10][240]  ( .D(n2861), .CLK(clk), .Q(\ram[10][240] ) );
  DFFX1_HVT \ram_reg[10][239]  ( .D(n2860), .CLK(clk), .Q(\ram[10][239] ) );
  DFFX1_HVT \ram_reg[10][238]  ( .D(n2859), .CLK(clk), .Q(\ram[10][238] ) );
  DFFX1_HVT \ram_reg[10][237]  ( .D(n2858), .CLK(clk), .Q(\ram[10][237] ) );
  DFFX1_HVT \ram_reg[10][236]  ( .D(n2857), .CLK(clk), .Q(\ram[10][236] ) );
  DFFX1_HVT \ram_reg[10][235]  ( .D(n2856), .CLK(clk), .Q(\ram[10][235] ) );
  DFFX1_HVT \ram_reg[10][234]  ( .D(n2855), .CLK(clk), .Q(\ram[10][234] ) );
  DFFX1_HVT \ram_reg[10][233]  ( .D(n2854), .CLK(clk), .Q(\ram[10][233] ) );
  DFFX1_HVT \ram_reg[10][232]  ( .D(n2853), .CLK(clk), .Q(\ram[10][232] ) );
  DFFX1_HVT \ram_reg[10][231]  ( .D(n2852), .CLK(clk), .Q(\ram[10][231] ) );
  DFFX1_HVT \ram_reg[10][230]  ( .D(n2851), .CLK(clk), .Q(\ram[10][230] ) );
  DFFX1_HVT \ram_reg[10][229]  ( .D(n2850), .CLK(clk), .Q(\ram[10][229] ) );
  DFFX1_HVT \ram_reg[10][228]  ( .D(n2849), .CLK(clk), .Q(\ram[10][228] ) );
  DFFX1_HVT \ram_reg[10][227]  ( .D(n2848), .CLK(clk), .Q(\ram[10][227] ) );
  DFFX1_HVT \ram_reg[10][226]  ( .D(n2847), .CLK(clk), .Q(\ram[10][226] ) );
  DFFX1_HVT \ram_reg[10][225]  ( .D(n2846), .CLK(clk), .Q(\ram[10][225] ) );
  DFFX1_HVT \ram_reg[10][224]  ( .D(n2845), .CLK(clk), .Q(\ram[10][224] ) );
  DFFX1_HVT \ram_reg[10][223]  ( .D(n2844), .CLK(clk), .Q(\ram[10][223] ) );
  DFFX1_HVT \ram_reg[10][222]  ( .D(n2843), .CLK(clk), .Q(\ram[10][222] ) );
  DFFX1_HVT \ram_reg[10][221]  ( .D(n2842), .CLK(clk), .Q(\ram[10][221] ) );
  DFFX1_HVT \ram_reg[10][220]  ( .D(n2841), .CLK(clk), .Q(\ram[10][220] ), 
        .QN(n5438) );
  DFFX1_HVT \ram_reg[10][219]  ( .D(n2840), .CLK(clk), .Q(\ram[10][219] ) );
  DFFX1_HVT \ram_reg[10][218]  ( .D(n2839), .CLK(clk), .Q(\ram[10][218] ) );
  DFFX1_HVT \ram_reg[10][217]  ( .D(n2838), .CLK(clk), .Q(\ram[10][217] ) );
  DFFX1_HVT \ram_reg[10][216]  ( .D(n2837), .CLK(clk), .Q(\ram[10][216] ) );
  DFFX1_HVT \ram_reg[10][215]  ( .D(n2836), .CLK(clk), .Q(\ram[10][215] ) );
  DFFX1_HVT \ram_reg[10][214]  ( .D(n2835), .CLK(clk), .Q(\ram[10][214] ) );
  DFFX1_HVT \ram_reg[10][213]  ( .D(n2834), .CLK(clk), .Q(\ram[10][213] ) );
  DFFX1_HVT \ram_reg[10][212]  ( .D(n2833), .CLK(clk), .Q(\ram[10][212] ) );
  DFFX1_HVT \ram_reg[10][211]  ( .D(n2832), .CLK(clk), .Q(\ram[10][211] ) );
  DFFX1_HVT \ram_reg[10][210]  ( .D(n2831), .CLK(clk), .Q(\ram[10][210] ) );
  DFFX1_HVT \ram_reg[10][209]  ( .D(n2830), .CLK(clk), .Q(\ram[10][209] ) );
  DFFX1_HVT \ram_reg[10][208]  ( .D(n2829), .CLK(clk), .Q(\ram[10][208] ) );
  DFFX1_HVT \ram_reg[10][207]  ( .D(n2828), .CLK(clk), .Q(\ram[10][207] ) );
  DFFX1_HVT \ram_reg[10][206]  ( .D(n2827), .CLK(clk), .Q(\ram[10][206] ) );
  DFFX1_HVT \ram_reg[10][205]  ( .D(n2826), .CLK(clk), .Q(\ram[10][205] ) );
  DFFX1_HVT \ram_reg[10][204]  ( .D(n2825), .CLK(clk), .Q(\ram[10][204] ) );
  DFFX1_HVT \ram_reg[10][203]  ( .D(n2824), .CLK(clk), .Q(\ram[10][203] ) );
  DFFX1_HVT \ram_reg[10][202]  ( .D(n2823), .CLK(clk), .Q(\ram[10][202] ) );
  DFFX1_HVT \ram_reg[10][201]  ( .D(n2822), .CLK(clk), .Q(\ram[10][201] ) );
  DFFX1_HVT \ram_reg[10][200]  ( .D(n2821), .CLK(clk), .Q(\ram[10][200] ) );
  DFFX1_HVT \ram_reg[10][199]  ( .D(n2820), .CLK(clk), .Q(\ram[10][199] ) );
  DFFX1_HVT \ram_reg[10][198]  ( .D(n2819), .CLK(clk), .Q(\ram[10][198] ) );
  DFFX1_HVT \ram_reg[10][197]  ( .D(n2818), .CLK(clk), .Q(\ram[10][197] ) );
  DFFX1_HVT \ram_reg[10][196]  ( .D(n2817), .CLK(clk), .Q(\ram[10][196] ) );
  DFFX1_HVT \ram_reg[10][195]  ( .D(n2816), .CLK(clk), .Q(\ram[10][195] ) );
  DFFX1_HVT \ram_reg[10][194]  ( .D(n2815), .CLK(clk), .Q(\ram[10][194] ) );
  DFFX1_HVT \ram_reg[10][193]  ( .D(n2814), .CLK(clk), .Q(\ram[10][193] ) );
  DFFX1_HVT \ram_reg[10][192]  ( .D(n2813), .CLK(clk), .Q(\ram[10][192] ) );
  DFFX1_HVT \ram_reg[10][191]  ( .D(n2812), .CLK(clk), .Q(\ram[10][191] ) );
  DFFX1_HVT \ram_reg[10][190]  ( .D(n2811), .CLK(clk), .Q(\ram[10][190] ) );
  DFFX1_HVT \ram_reg[10][189]  ( .D(n2810), .CLK(clk), .Q(\ram[10][189] ) );
  DFFX1_HVT \ram_reg[10][188]  ( .D(n2809), .CLK(clk), .Q(\ram[10][188] ) );
  DFFX1_HVT \ram_reg[10][187]  ( .D(n2808), .CLK(clk), .Q(\ram[10][187] ) );
  DFFX1_HVT \ram_reg[10][186]  ( .D(n2807), .CLK(clk), .Q(\ram[10][186] ) );
  DFFX1_HVT \ram_reg[10][185]  ( .D(n2806), .CLK(clk), .Q(\ram[10][185] ) );
  DFFX1_HVT \ram_reg[10][184]  ( .D(n2805), .CLK(clk), .Q(\ram[10][184] ) );
  DFFX1_HVT \ram_reg[10][183]  ( .D(n2804), .CLK(clk), .Q(\ram[10][183] ) );
  DFFX1_HVT \ram_reg[10][182]  ( .D(n2803), .CLK(clk), .Q(\ram[10][182] ) );
  DFFX1_HVT \ram_reg[10][181]  ( .D(n2802), .CLK(clk), .Q(\ram[10][181] ) );
  DFFX1_HVT \ram_reg[10][180]  ( .D(n2801), .CLK(clk), .Q(\ram[10][180] ) );
  DFFX1_HVT \ram_reg[10][179]  ( .D(n2800), .CLK(clk), .Q(\ram[10][179] ) );
  DFFX1_HVT \ram_reg[10][178]  ( .D(n2799), .CLK(clk), .Q(\ram[10][178] ) );
  DFFX1_HVT \ram_reg[10][177]  ( .D(n2798), .CLK(clk), .Q(\ram[10][177] ) );
  DFFX1_HVT \ram_reg[10][176]  ( .D(n2797), .CLK(clk), .Q(\ram[10][176] ) );
  DFFX1_HVT \ram_reg[10][175]  ( .D(n2796), .CLK(clk), .Q(\ram[10][175] ) );
  DFFX1_HVT \ram_reg[10][174]  ( .D(n2795), .CLK(clk), .Q(\ram[10][174] ) );
  DFFX1_HVT \ram_reg[10][173]  ( .D(n2794), .CLK(clk), .Q(\ram[10][173] ) );
  DFFX1_HVT \ram_reg[10][172]  ( .D(n2793), .CLK(clk), .Q(\ram[10][172] ) );
  DFFX1_HVT \ram_reg[10][171]  ( .D(n2792), .CLK(clk), .Q(\ram[10][171] ) );
  DFFX1_HVT \ram_reg[10][170]  ( .D(n2791), .CLK(clk), .Q(\ram[10][170] ) );
  DFFX1_HVT \ram_reg[10][169]  ( .D(n2790), .CLK(clk), .Q(\ram[10][169] ) );
  DFFX1_HVT \ram_reg[10][168]  ( .D(n2789), .CLK(clk), .Q(\ram[10][168] ) );
  DFFX1_HVT \ram_reg[10][167]  ( .D(n2788), .CLK(clk), .Q(\ram[10][167] ) );
  DFFX1_HVT \ram_reg[10][166]  ( .D(n2787), .CLK(clk), .Q(\ram[10][166] ) );
  DFFX1_HVT \ram_reg[10][165]  ( .D(n2786), .CLK(clk), .Q(\ram[10][165] ) );
  DFFX1_HVT \ram_reg[10][164]  ( .D(n2785), .CLK(clk), .Q(\ram[10][164] ) );
  DFFX1_HVT \ram_reg[10][163]  ( .D(n2784), .CLK(clk), .Q(\ram[10][163] ) );
  DFFX1_HVT \ram_reg[10][162]  ( .D(n2783), .CLK(clk), .Q(\ram[10][162] ), 
        .QN(n3949) );
  DFFX1_HVT \ram_reg[10][161]  ( .D(n2782), .CLK(clk), .Q(\ram[10][161] ) );
  DFFX1_HVT \ram_reg[10][160]  ( .D(n2781), .CLK(clk), .Q(\ram[10][160] ) );
  DFFX1_HVT \ram_reg[10][159]  ( .D(n2780), .CLK(clk), .Q(\ram[10][159] ) );
  DFFX1_HVT \ram_reg[10][158]  ( .D(n2779), .CLK(clk), .Q(\ram[10][158] ) );
  DFFX1_HVT \ram_reg[10][157]  ( .D(n2778), .CLK(clk), .Q(\ram[10][157] ) );
  DFFX1_HVT \ram_reg[10][156]  ( .D(n2777), .CLK(clk), .Q(\ram[10][156] ) );
  DFFX1_HVT \ram_reg[10][155]  ( .D(n2776), .CLK(clk), .Q(\ram[10][155] ) );
  DFFX1_HVT \ram_reg[10][154]  ( .D(n2775), .CLK(clk), .Q(\ram[10][154] ) );
  DFFX1_HVT \ram_reg[10][153]  ( .D(n2774), .CLK(clk), .Q(\ram[10][153] ) );
  DFFX1_HVT \ram_reg[10][152]  ( .D(n2773), .CLK(clk), .Q(\ram[10][152] ) );
  DFFX1_HVT \ram_reg[10][151]  ( .D(n2772), .CLK(clk), .Q(\ram[10][151] ) );
  DFFX1_HVT \ram_reg[10][150]  ( .D(n2771), .CLK(clk), .Q(\ram[10][150] ) );
  DFFX1_HVT \ram_reg[10][149]  ( .D(n2770), .CLK(clk), .Q(\ram[10][149] ) );
  DFFX1_HVT \ram_reg[10][148]  ( .D(n2769), .CLK(clk), .Q(\ram[10][148] ) );
  DFFX1_HVT \ram_reg[10][147]  ( .D(n2768), .CLK(clk), .Q(\ram[10][147] ) );
  DFFX1_HVT \ram_reg[10][146]  ( .D(n2767), .CLK(clk), .Q(\ram[10][146] ) );
  DFFX1_HVT \ram_reg[10][145]  ( .D(n2766), .CLK(clk), .Q(\ram[10][145] ) );
  DFFX1_HVT \ram_reg[10][144]  ( .D(n2765), .CLK(clk), .Q(\ram[10][144] ) );
  DFFX1_HVT \ram_reg[10][143]  ( .D(n2764), .CLK(clk), .Q(\ram[10][143] ) );
  DFFX1_HVT \ram_reg[10][142]  ( .D(n2763), .CLK(clk), .Q(\ram[10][142] ) );
  DFFX1_HVT \ram_reg[10][141]  ( .D(n2762), .CLK(clk), .Q(\ram[10][141] ) );
  DFFX1_HVT \ram_reg[10][140]  ( .D(n2761), .CLK(clk), .Q(\ram[10][140] ) );
  DFFX1_HVT \ram_reg[10][139]  ( .D(n2760), .CLK(clk), .Q(\ram[10][139] ) );
  DFFX1_HVT \ram_reg[10][138]  ( .D(n2759), .CLK(clk), .Q(\ram[10][138] ) );
  DFFX1_HVT \ram_reg[10][137]  ( .D(n2758), .CLK(clk), .Q(\ram[10][137] ) );
  DFFX1_HVT \ram_reg[10][136]  ( .D(n2757), .CLK(clk), .Q(\ram[10][136] ), 
        .QN(n4172) );
  DFFX1_HVT \ram_reg[10][135]  ( .D(n2756), .CLK(clk), .Q(\ram[10][135] ) );
  DFFX1_HVT \ram_reg[10][134]  ( .D(n2755), .CLK(clk), .Q(\ram[10][134] ) );
  DFFX1_HVT \ram_reg[10][133]  ( .D(n2754), .CLK(clk), .Q(\ram[10][133] ) );
  DFFX1_HVT \ram_reg[10][132]  ( .D(n2753), .CLK(clk), .Q(\ram[10][132] ) );
  DFFX1_HVT \ram_reg[10][131]  ( .D(n2752), .CLK(clk), .Q(\ram[10][131] ) );
  DFFX1_HVT \ram_reg[10][130]  ( .D(n2751), .CLK(clk), .Q(\ram[10][130] ) );
  DFFX1_HVT \ram_reg[10][129]  ( .D(n2750), .CLK(clk), .Q(\ram[10][129] ) );
  DFFX1_HVT \ram_reg[10][128]  ( .D(n2749), .CLK(clk), .Q(\ram[10][128] ) );
  DFFX1_HVT \ram_reg[10][127]  ( .D(n2748), .CLK(clk), .Q(\ram[10][127] ) );
  DFFX1_HVT \ram_reg[10][126]  ( .D(n2747), .CLK(clk), .Q(\ram[10][126] ) );
  DFFX1_HVT \ram_reg[10][125]  ( .D(n2746), .CLK(clk), .Q(\ram[10][125] ) );
  DFFX1_HVT \ram_reg[10][124]  ( .D(n2745), .CLK(clk), .Q(\ram[10][124] ) );
  DFFX1_HVT \ram_reg[10][123]  ( .D(n2744), .CLK(clk), .Q(\ram[10][123] ) );
  DFFX1_HVT \ram_reg[10][122]  ( .D(n2743), .CLK(clk), .Q(\ram[10][122] ) );
  DFFX1_HVT \ram_reg[10][121]  ( .D(n2742), .CLK(clk), .Q(\ram[10][121] ) );
  DFFX1_HVT \ram_reg[10][120]  ( .D(n2741), .CLK(clk), .Q(\ram[10][120] ) );
  DFFX1_HVT \ram_reg[10][119]  ( .D(n2740), .CLK(clk), .Q(\ram[10][119] ) );
  DFFX1_HVT \ram_reg[10][118]  ( .D(n2739), .CLK(clk), .Q(\ram[10][118] ) );
  DFFX1_HVT \ram_reg[10][117]  ( .D(n2738), .CLK(clk), .Q(\ram[10][117] ) );
  DFFX1_HVT \ram_reg[10][116]  ( .D(n2737), .CLK(clk), .Q(\ram[10][116] ) );
  DFFX1_HVT \ram_reg[10][115]  ( .D(n2736), .CLK(clk), .Q(\ram[10][115] ) );
  DFFX1_HVT \ram_reg[10][114]  ( .D(n2735), .CLK(clk), .Q(\ram[10][114] ) );
  DFFX1_HVT \ram_reg[10][113]  ( .D(n2734), .CLK(clk), .Q(\ram[10][113] ) );
  DFFX1_HVT \ram_reg[10][112]  ( .D(n2733), .CLK(clk), .Q(\ram[10][112] ) );
  DFFX1_HVT \ram_reg[10][111]  ( .D(n2732), .CLK(clk), .Q(\ram[10][111] ) );
  DFFX1_HVT \ram_reg[10][110]  ( .D(n2731), .CLK(clk), .Q(\ram[10][110] ) );
  DFFX1_HVT \ram_reg[10][109]  ( .D(n2730), .CLK(clk), .Q(\ram[10][109] ) );
  DFFX1_HVT \ram_reg[10][108]  ( .D(n2729), .CLK(clk), .Q(\ram[10][108] ) );
  DFFX1_HVT \ram_reg[10][107]  ( .D(n2728), .CLK(clk), .Q(\ram[10][107] ) );
  DFFX1_HVT \ram_reg[10][106]  ( .D(n2727), .CLK(clk), .Q(\ram[10][106] ) );
  DFFX1_HVT \ram_reg[10][105]  ( .D(n2726), .CLK(clk), .Q(\ram[10][105] ) );
  DFFX1_HVT \ram_reg[10][104]  ( .D(n2725), .CLK(clk), .Q(\ram[10][104] ) );
  DFFX1_HVT \ram_reg[10][103]  ( .D(n2724), .CLK(clk), .Q(\ram[10][103] ) );
  DFFX1_HVT \ram_reg[10][102]  ( .D(n2723), .CLK(clk), .Q(\ram[10][102] ) );
  DFFX1_HVT \ram_reg[10][101]  ( .D(n2722), .CLK(clk), .Q(\ram[10][101] ) );
  DFFX1_HVT \ram_reg[10][100]  ( .D(n2721), .CLK(clk), .Q(\ram[10][100] ) );
  DFFX1_HVT \ram_reg[10][99]  ( .D(n2720), .CLK(clk), .Q(\ram[10][99] ) );
  DFFX1_HVT \ram_reg[10][98]  ( .D(n2719), .CLK(clk), .Q(\ram[10][98] ) );
  DFFX1_HVT \ram_reg[10][97]  ( .D(n2718), .CLK(clk), .Q(\ram[10][97] ) );
  DFFX1_HVT \ram_reg[10][96]  ( .D(n2717), .CLK(clk), .Q(\ram[10][96] ) );
  DFFX1_HVT \ram_reg[10][95]  ( .D(n2716), .CLK(clk), .Q(\ram[10][95] ) );
  DFFX1_HVT \ram_reg[10][94]  ( .D(n2715), .CLK(clk), .Q(\ram[10][94] ) );
  DFFX1_HVT \ram_reg[10][93]  ( .D(n2714), .CLK(clk), .Q(\ram[10][93] ) );
  DFFX1_HVT \ram_reg[10][92]  ( .D(n2713), .CLK(clk), .Q(\ram[10][92] ) );
  DFFX1_HVT \ram_reg[10][91]  ( .D(n2712), .CLK(clk), .Q(\ram[10][91] ) );
  DFFX1_HVT \ram_reg[10][90]  ( .D(n2711), .CLK(clk), .Q(\ram[10][90] ) );
  DFFX1_HVT \ram_reg[10][89]  ( .D(n2710), .CLK(clk), .Q(\ram[10][89] ) );
  DFFX1_HVT \ram_reg[10][88]  ( .D(n2709), .CLK(clk), .Q(\ram[10][88] ) );
  DFFX1_HVT \ram_reg[10][87]  ( .D(n2708), .CLK(clk), .Q(\ram[10][87] ) );
  DFFX1_HVT \ram_reg[10][86]  ( .D(n2707), .CLK(clk), .Q(\ram[10][86] ) );
  DFFX1_HVT \ram_reg[10][85]  ( .D(n2706), .CLK(clk), .Q(\ram[10][85] ) );
  DFFX1_HVT \ram_reg[10][84]  ( .D(n2705), .CLK(clk), .Q(\ram[10][84] ) );
  DFFX1_HVT \ram_reg[10][83]  ( .D(n2704), .CLK(clk), .Q(\ram[10][83] ) );
  DFFX1_HVT \ram_reg[10][82]  ( .D(n2703), .CLK(clk), .Q(\ram[10][82] ) );
  DFFX1_HVT \ram_reg[10][81]  ( .D(n2702), .CLK(clk), .Q(\ram[10][81] ) );
  DFFX1_HVT \ram_reg[10][80]  ( .D(n2701), .CLK(clk), .Q(\ram[10][80] ) );
  DFFX1_HVT \ram_reg[10][79]  ( .D(n2700), .CLK(clk), .Q(\ram[10][79] ) );
  DFFX1_HVT \ram_reg[10][78]  ( .D(n2699), .CLK(clk), .Q(\ram[10][78] ) );
  DFFX1_HVT \ram_reg[10][77]  ( .D(n2698), .CLK(clk), .Q(\ram[10][77] ) );
  DFFX1_HVT \ram_reg[10][76]  ( .D(n2697), .CLK(clk), .Q(\ram[10][76] ) );
  DFFX1_HVT \ram_reg[10][75]  ( .D(n2696), .CLK(clk), .Q(\ram[10][75] ) );
  DFFX1_HVT \ram_reg[10][74]  ( .D(n2695), .CLK(clk), .Q(\ram[10][74] ) );
  DFFX1_HVT \ram_reg[10][73]  ( .D(n2694), .CLK(clk), .Q(\ram[10][73] ) );
  DFFX1_HVT \ram_reg[10][72]  ( .D(n2693), .CLK(clk), .Q(\ram[10][72] ) );
  DFFX1_HVT \ram_reg[10][71]  ( .D(n2692), .CLK(clk), .Q(\ram[10][71] ) );
  DFFX1_HVT \ram_reg[10][70]  ( .D(n2691), .CLK(clk), .Q(\ram[10][70] ) );
  DFFX1_HVT \ram_reg[10][69]  ( .D(n2690), .CLK(clk), .Q(\ram[10][69] ) );
  DFFX1_HVT \ram_reg[10][68]  ( .D(n2689), .CLK(clk), .Q(\ram[10][68] ) );
  DFFX1_HVT \ram_reg[10][67]  ( .D(n2688), .CLK(clk), .Q(\ram[10][67] ) );
  DFFX1_HVT \ram_reg[10][66]  ( .D(n2687), .CLK(clk), .Q(\ram[10][66] ) );
  DFFX1_HVT \ram_reg[10][65]  ( .D(n2686), .CLK(clk), .Q(\ram[10][65] ) );
  DFFX1_HVT \ram_reg[10][64]  ( .D(n2685), .CLK(clk), .Q(\ram[10][64] ) );
  DFFX1_HVT \ram_reg[10][63]  ( .D(n2684), .CLK(clk), .Q(\ram[10][63] ) );
  DFFX1_HVT \ram_reg[10][62]  ( .D(n2683), .CLK(clk), .Q(\ram[10][62] ) );
  DFFX1_HVT \ram_reg[10][61]  ( .D(n2682), .CLK(clk), .Q(\ram[10][61] ) );
  DFFX1_HVT \ram_reg[10][60]  ( .D(n2681), .CLK(clk), .Q(\ram[10][60] ) );
  DFFX1_HVT \ram_reg[10][59]  ( .D(n2680), .CLK(clk), .Q(\ram[10][59] ) );
  DFFX1_HVT \ram_reg[10][58]  ( .D(n2679), .CLK(clk), .Q(\ram[10][58] ), .QN(
        n4817) );
  DFFX1_HVT \ram_reg[10][57]  ( .D(n2678), .CLK(clk), .Q(\ram[10][57] ) );
  DFFX1_HVT \ram_reg[10][56]  ( .D(n2677), .CLK(clk), .Q(\ram[10][56] ) );
  DFFX1_HVT \ram_reg[10][55]  ( .D(n2676), .CLK(clk), .Q(\ram[10][55] ) );
  DFFX1_HVT \ram_reg[10][54]  ( .D(n2675), .CLK(clk), .Q(\ram[10][54] ) );
  DFFX1_HVT \ram_reg[10][53]  ( .D(n2674), .CLK(clk), .Q(\ram[10][53] ) );
  DFFX1_HVT \ram_reg[10][52]  ( .D(n2673), .CLK(clk), .Q(\ram[10][52] ) );
  DFFX1_HVT \ram_reg[10][51]  ( .D(n2672), .CLK(clk), .Q(\ram[10][51] ) );
  DFFX1_HVT \ram_reg[10][50]  ( .D(n2671), .CLK(clk), .Q(\ram[10][50] ) );
  DFFX1_HVT \ram_reg[10][49]  ( .D(n2670), .CLK(clk), .Q(\ram[10][49] ) );
  DFFX1_HVT \ram_reg[10][48]  ( .D(n2669), .CLK(clk), .Q(\ram[10][48] ) );
  DFFX1_HVT \ram_reg[10][47]  ( .D(n2668), .CLK(clk), .Q(\ram[10][47] ) );
  DFFX1_HVT \ram_reg[10][46]  ( .D(n2667), .CLK(clk), .Q(\ram[10][46] ) );
  DFFX1_HVT \ram_reg[10][45]  ( .D(n2666), .CLK(clk), .Q(\ram[10][45] ) );
  DFFX1_HVT \ram_reg[10][44]  ( .D(n2665), .CLK(clk), .Q(\ram[10][44] ) );
  DFFX1_HVT \ram_reg[10][43]  ( .D(n2664), .CLK(clk), .Q(\ram[10][43] ) );
  DFFX1_HVT \ram_reg[10][42]  ( .D(n2663), .CLK(clk), .Q(\ram[10][42] ) );
  DFFX1_HVT \ram_reg[10][41]  ( .D(n2662), .CLK(clk), .Q(\ram[10][41] ) );
  DFFX1_HVT \ram_reg[10][40]  ( .D(n2661), .CLK(clk), .Q(\ram[10][40] ) );
  DFFX1_HVT \ram_reg[10][39]  ( .D(n2660), .CLK(clk), .Q(\ram[10][39] ) );
  DFFX1_HVT \ram_reg[10][38]  ( .D(n2659), .CLK(clk), .Q(\ram[10][38] ), .QN(
        n1357) );
  DFFX1_HVT \ram_reg[10][37]  ( .D(n2658), .CLK(clk), .Q(\ram[10][37] ) );
  DFFX1_HVT \ram_reg[10][36]  ( .D(n2657), .CLK(clk), .Q(\ram[10][36] ) );
  DFFX1_HVT \ram_reg[10][35]  ( .D(n2656), .CLK(clk), .Q(\ram[10][35] ) );
  DFFX1_HVT \ram_reg[10][34]  ( .D(n2655), .CLK(clk), .Q(\ram[10][34] ) );
  DFFX1_HVT \ram_reg[10][33]  ( .D(n2654), .CLK(clk), .Q(\ram[10][33] ) );
  DFFX1_HVT \ram_reg[10][32]  ( .D(n2653), .CLK(clk), .Q(\ram[10][32] ) );
  DFFX1_HVT \ram_reg[10][31]  ( .D(n2652), .CLK(clk), .Q(\ram[10][31] ) );
  DFFX1_HVT \ram_reg[10][30]  ( .D(n2651), .CLK(clk), .Q(\ram[10][30] ) );
  DFFX1_HVT \ram_reg[10][29]  ( .D(n2650), .CLK(clk), .Q(\ram[10][29] ) );
  DFFX1_HVT \ram_reg[10][28]  ( .D(n2649), .CLK(clk), .Q(\ram[10][28] ) );
  DFFX1_HVT \ram_reg[10][27]  ( .D(n2648), .CLK(clk), .Q(\ram[10][27] ) );
  DFFX1_HVT \ram_reg[10][26]  ( .D(n2647), .CLK(clk), .Q(\ram[10][26] ) );
  DFFX1_HVT \ram_reg[10][25]  ( .D(n2646), .CLK(clk), .Q(\ram[10][25] ) );
  DFFX1_HVT \ram_reg[10][24]  ( .D(n2645), .CLK(clk), .Q(\ram[10][24] ) );
  DFFX1_HVT \ram_reg[10][23]  ( .D(n2644), .CLK(clk), .Q(\ram[10][23] ) );
  DFFX1_HVT \ram_reg[10][22]  ( .D(n2643), .CLK(clk), .Q(\ram[10][22] ) );
  DFFX1_HVT \ram_reg[10][21]  ( .D(n2642), .CLK(clk), .Q(\ram[10][21] ) );
  DFFX1_HVT \ram_reg[10][20]  ( .D(n2641), .CLK(clk), .Q(\ram[10][20] ), .QN(
        n6483) );
  DFFX1_HVT \ram_reg[10][19]  ( .D(n2640), .CLK(clk), .Q(\ram[10][19] ) );
  DFFX1_HVT \ram_reg[10][18]  ( .D(n2639), .CLK(clk), .Q(\ram[10][18] ) );
  DFFX1_HVT \ram_reg[10][17]  ( .D(n2638), .CLK(clk), .Q(\ram[10][17] ) );
  DFFX1_HVT \ram_reg[10][16]  ( .D(n2637), .CLK(clk), .Q(\ram[10][16] ) );
  DFFX1_HVT \ram_reg[10][15]  ( .D(n2636), .CLK(clk), .Q(\ram[10][15] ) );
  DFFX1_HVT \ram_reg[10][14]  ( .D(n2635), .CLK(clk), .Q(\ram[10][14] ) );
  DFFX1_HVT \ram_reg[10][13]  ( .D(n2634), .CLK(clk), .Q(\ram[10][13] ) );
  DFFX1_HVT \ram_reg[10][12]  ( .D(n2633), .CLK(clk), .Q(\ram[10][12] ) );
  DFFX1_HVT \ram_reg[10][11]  ( .D(n2632), .CLK(clk), .Q(\ram[10][11] ) );
  DFFX1_HVT \ram_reg[10][10]  ( .D(n2631), .CLK(clk), .Q(\ram[10][10] ) );
  DFFX1_HVT \ram_reg[10][9]  ( .D(n2630), .CLK(clk), .Q(\ram[10][9] ) );
  DFFX1_HVT \ram_reg[10][8]  ( .D(n2629), .CLK(clk), .Q(\ram[10][8] ) );
  DFFX1_HVT \ram_reg[10][7]  ( .D(n2628), .CLK(clk), .Q(\ram[10][7] ) );
  DFFX1_HVT \ram_reg[10][6]  ( .D(n2627), .CLK(clk), .Q(\ram[10][6] ) );
  DFFX1_HVT \ram_reg[10][5]  ( .D(n2626), .CLK(clk), .Q(\ram[10][5] ) );
  DFFX1_HVT \ram_reg[10][4]  ( .D(n2625), .CLK(clk), .Q(\ram[10][4] ) );
  DFFX1_HVT \ram_reg[10][3]  ( .D(n2624), .CLK(clk), .Q(\ram[10][3] ) );
  DFFX1_HVT \ram_reg[10][2]  ( .D(n2623), .CLK(clk), .Q(\ram[10][2] ) );
  DFFX1_HVT \ram_reg[10][1]  ( .D(n2622), .CLK(clk), .Q(\ram[10][1] ) );
  DFFX1_HVT \ram_reg[10][0]  ( .D(n2621), .CLK(clk), .Q(\ram[10][0] ) );
  DFFX1_HVT \ram_reg[9][255]  ( .D(n2620), .CLK(clk), .Q(\ram[9][255] ) );
  DFFX1_HVT \ram_reg[9][254]  ( .D(n2619), .CLK(clk), .Q(\ram[9][254] ) );
  DFFX1_HVT \ram_reg[9][253]  ( .D(n2618), .CLK(clk), .Q(\ram[9][253] ) );
  DFFX1_HVT \ram_reg[9][252]  ( .D(n2617), .CLK(clk), .Q(\ram[9][252] ) );
  DFFX1_HVT \ram_reg[9][251]  ( .D(n2616), .CLK(clk), .Q(\ram[9][251] ) );
  DFFX1_HVT \ram_reg[9][250]  ( .D(n2615), .CLK(clk), .Q(\ram[9][250] ) );
  DFFX1_HVT \ram_reg[9][249]  ( .D(n2614), .CLK(clk), .Q(\ram[9][249] ) );
  DFFX1_HVT \ram_reg[9][248]  ( .D(n2613), .CLK(clk), .Q(\ram[9][248] ) );
  DFFX1_HVT \ram_reg[9][247]  ( .D(n2612), .CLK(clk), .Q(\ram[9][247] ) );
  DFFX1_HVT \ram_reg[9][246]  ( .D(n2611), .CLK(clk), .Q(\ram[9][246] ) );
  DFFX1_HVT \ram_reg[9][245]  ( .D(n2610), .CLK(clk), .Q(\ram[9][245] ) );
  DFFX1_HVT \ram_reg[9][244]  ( .D(n2609), .CLK(clk), .Q(\ram[9][244] ) );
  DFFX1_HVT \ram_reg[9][243]  ( .D(n2608), .CLK(clk), .Q(\ram[9][243] ) );
  DFFX1_HVT \ram_reg[9][242]  ( .D(n2607), .CLK(clk), .Q(\ram[9][242] ) );
  DFFX1_HVT \ram_reg[9][241]  ( .D(n2606), .CLK(clk), .Q(\ram[9][241] ) );
  DFFX1_HVT \ram_reg[9][240]  ( .D(n2605), .CLK(clk), .Q(\ram[9][240] ) );
  DFFX1_HVT \ram_reg[9][239]  ( .D(n2604), .CLK(clk), .Q(\ram[9][239] ) );
  DFFX1_HVT \ram_reg[9][238]  ( .D(n2603), .CLK(clk), .Q(\ram[9][238] ) );
  DFFX1_HVT \ram_reg[9][237]  ( .D(n2602), .CLK(clk), .Q(\ram[9][237] ) );
  DFFX1_HVT \ram_reg[9][236]  ( .D(n2601), .CLK(clk), .Q(\ram[9][236] ) );
  DFFX1_HVT \ram_reg[9][235]  ( .D(n2600), .CLK(clk), .Q(\ram[9][235] ) );
  DFFX1_HVT \ram_reg[9][234]  ( .D(n2599), .CLK(clk), .Q(\ram[9][234] ) );
  DFFX1_HVT \ram_reg[9][233]  ( .D(n2598), .CLK(clk), .Q(\ram[9][233] ) );
  DFFX1_HVT \ram_reg[9][232]  ( .D(n2597), .CLK(clk), .Q(\ram[9][232] ) );
  DFFX1_HVT \ram_reg[9][231]  ( .D(n2596), .CLK(clk), .Q(\ram[9][231] ) );
  DFFX1_HVT \ram_reg[9][230]  ( .D(n2595), .CLK(clk), .Q(\ram[9][230] ) );
  DFFX1_HVT \ram_reg[9][229]  ( .D(n2594), .CLK(clk), .Q(\ram[9][229] ) );
  DFFX1_HVT \ram_reg[9][228]  ( .D(n2593), .CLK(clk), .Q(\ram[9][228] ) );
  DFFX1_HVT \ram_reg[9][227]  ( .D(n2592), .CLK(clk), .Q(\ram[9][227] ) );
  DFFX1_HVT \ram_reg[9][226]  ( .D(n2591), .CLK(clk), .Q(\ram[9][226] ), .QN(
        n4235) );
  DFFX1_HVT \ram_reg[9][225]  ( .D(n2590), .CLK(clk), .Q(\ram[9][225] ), .QN(
        n4226) );
  DFFX1_HVT \ram_reg[9][224]  ( .D(n2589), .CLK(clk), .Q(\ram[9][224] ) );
  DFFX1_HVT \ram_reg[9][223]  ( .D(n2588), .CLK(clk), .Q(\ram[9][223] ) );
  DFFX1_HVT \ram_reg[9][222]  ( .D(n2587), .CLK(clk), .Q(\ram[9][222] ) );
  DFFX1_HVT \ram_reg[9][221]  ( .D(n2586), .CLK(clk), .Q(\ram[9][221] ) );
  DFFX1_HVT \ram_reg[9][220]  ( .D(n2585), .CLK(clk), .Q(\ram[9][220] ), .QN(
        n5929) );
  DFFX1_HVT \ram_reg[9][219]  ( .D(n2584), .CLK(clk), .Q(\ram[9][219] ) );
  DFFX1_HVT \ram_reg[9][218]  ( .D(n2583), .CLK(clk), .Q(\ram[9][218] ) );
  DFFX1_HVT \ram_reg[9][217]  ( .D(n2582), .CLK(clk), .Q(\ram[9][217] ) );
  DFFX1_HVT \ram_reg[9][216]  ( .D(n2581), .CLK(clk), .Q(\ram[9][216] ) );
  DFFX1_HVT \ram_reg[9][215]  ( .D(n2580), .CLK(clk), .Q(\ram[9][215] ) );
  DFFX1_HVT \ram_reg[9][214]  ( .D(n2579), .CLK(clk), .Q(\ram[9][214] ) );
  DFFX1_HVT \ram_reg[9][213]  ( .D(n2578), .CLK(clk), .Q(\ram[9][213] ) );
  DFFX1_HVT \ram_reg[9][212]  ( .D(n2577), .CLK(clk), .Q(\ram[9][212] ) );
  DFFX1_HVT \ram_reg[9][211]  ( .D(n2576), .CLK(clk), .Q(\ram[9][211] ) );
  DFFX1_HVT \ram_reg[9][210]  ( .D(n2575), .CLK(clk), .Q(\ram[9][210] ) );
  DFFX1_HVT \ram_reg[9][209]  ( .D(n2574), .CLK(clk), .Q(\ram[9][209] ) );
  DFFX1_HVT \ram_reg[9][208]  ( .D(n2573), .CLK(clk), .Q(\ram[9][208] ) );
  DFFX1_HVT \ram_reg[9][207]  ( .D(n2572), .CLK(clk), .Q(\ram[9][207] ) );
  DFFX1_HVT \ram_reg[9][206]  ( .D(n2571), .CLK(clk), .Q(\ram[9][206] ) );
  DFFX1_HVT \ram_reg[9][205]  ( .D(n2570), .CLK(clk), .Q(\ram[9][205] ) );
  DFFX1_HVT \ram_reg[9][204]  ( .D(n2569), .CLK(clk), .Q(\ram[9][204] ) );
  DFFX1_HVT \ram_reg[9][203]  ( .D(n2568), .CLK(clk), .Q(\ram[9][203] ) );
  DFFX1_HVT \ram_reg[9][202]  ( .D(n2567), .CLK(clk), .Q(\ram[9][202] ) );
  DFFX1_HVT \ram_reg[9][201]  ( .D(n2566), .CLK(clk), .Q(\ram[9][201] ) );
  DFFX1_HVT \ram_reg[9][200]  ( .D(n2565), .CLK(clk), .Q(\ram[9][200] ) );
  DFFX1_HVT \ram_reg[9][199]  ( .D(n2564), .CLK(clk), .Q(\ram[9][199] ) );
  DFFX1_HVT \ram_reg[9][198]  ( .D(n2563), .CLK(clk), .Q(\ram[9][198] ) );
  DFFX1_HVT \ram_reg[9][197]  ( .D(n2562), .CLK(clk), .Q(\ram[9][197] ) );
  DFFX1_HVT \ram_reg[9][196]  ( .D(n2561), .CLK(clk), .Q(\ram[9][196] ) );
  DFFX1_HVT \ram_reg[9][195]  ( .D(n2560), .CLK(clk), .Q(\ram[9][195] ) );
  DFFX1_HVT \ram_reg[9][194]  ( .D(n2559), .CLK(clk), .Q(\ram[9][194] ) );
  DFFX1_HVT \ram_reg[9][193]  ( .D(n2558), .CLK(clk), .Q(\ram[9][193] ) );
  DFFX1_HVT \ram_reg[9][192]  ( .D(n2557), .CLK(clk), .Q(\ram[9][192] ) );
  DFFX1_HVT \ram_reg[9][191]  ( .D(n2556), .CLK(clk), .Q(\ram[9][191] ) );
  DFFX1_HVT \ram_reg[9][190]  ( .D(n2555), .CLK(clk), .Q(\ram[9][190] ) );
  DFFX1_HVT \ram_reg[9][189]  ( .D(n2554), .CLK(clk), .Q(\ram[9][189] ) );
  DFFX1_HVT \ram_reg[9][188]  ( .D(n2553), .CLK(clk), .Q(\ram[9][188] ) );
  DFFX1_HVT \ram_reg[9][187]  ( .D(n2552), .CLK(clk), .Q(\ram[9][187] ) );
  DFFX1_HVT \ram_reg[9][186]  ( .D(n2551), .CLK(clk), .Q(\ram[9][186] ) );
  DFFX1_HVT \ram_reg[9][185]  ( .D(n2550), .CLK(clk), .Q(\ram[9][185] ) );
  DFFX1_HVT \ram_reg[9][184]  ( .D(n2549), .CLK(clk), .Q(\ram[9][184] ) );
  DFFX1_HVT \ram_reg[9][183]  ( .D(n2548), .CLK(clk), .Q(\ram[9][183] ) );
  DFFX1_HVT \ram_reg[9][182]  ( .D(n2547), .CLK(clk), .Q(\ram[9][182] ) );
  DFFX1_HVT \ram_reg[9][181]  ( .D(n2546), .CLK(clk), .Q(\ram[9][181] ) );
  DFFX1_HVT \ram_reg[9][180]  ( .D(n2545), .CLK(clk), .Q(\ram[9][180] ) );
  DFFX1_HVT \ram_reg[9][179]  ( .D(n2544), .CLK(clk), .Q(\ram[9][179] ) );
  DFFX1_HVT \ram_reg[9][178]  ( .D(n2543), .CLK(clk), .Q(\ram[9][178] ) );
  DFFX1_HVT \ram_reg[9][177]  ( .D(n2542), .CLK(clk), .Q(\ram[9][177] ) );
  DFFX1_HVT \ram_reg[9][176]  ( .D(n2541), .CLK(clk), .Q(\ram[9][176] ) );
  DFFX1_HVT \ram_reg[9][175]  ( .D(n2540), .CLK(clk), .Q(\ram[9][175] ) );
  DFFX1_HVT \ram_reg[9][174]  ( .D(n2539), .CLK(clk), .Q(\ram[9][174] ) );
  DFFX1_HVT \ram_reg[9][173]  ( .D(n2538), .CLK(clk), .Q(\ram[9][173] ) );
  DFFX1_HVT \ram_reg[9][172]  ( .D(n2537), .CLK(clk), .Q(\ram[9][172] ) );
  DFFX1_HVT \ram_reg[9][171]  ( .D(n2536), .CLK(clk), .Q(\ram[9][171] ), .QN(
        n4351) );
  DFFX1_HVT \ram_reg[9][170]  ( .D(n2535), .CLK(clk), .Q(\ram[9][170] ) );
  DFFX1_HVT \ram_reg[9][169]  ( .D(n2534), .CLK(clk), .Q(\ram[9][169] ) );
  DFFX1_HVT \ram_reg[9][168]  ( .D(n2533), .CLK(clk), .Q(\ram[9][168] ) );
  DFFX1_HVT \ram_reg[9][167]  ( .D(n2532), .CLK(clk), .Q(\ram[9][167] ) );
  DFFX1_HVT \ram_reg[9][166]  ( .D(n2531), .CLK(clk), .Q(\ram[9][166] ) );
  DFFX1_HVT \ram_reg[9][165]  ( .D(n2530), .CLK(clk), .Q(\ram[9][165] ) );
  DFFX1_HVT \ram_reg[9][164]  ( .D(n2529), .CLK(clk), .Q(\ram[9][164] ) );
  DFFX1_HVT \ram_reg[9][163]  ( .D(n2528), .CLK(clk), .Q(\ram[9][163] ) );
  DFFX1_HVT \ram_reg[9][162]  ( .D(n2527), .CLK(clk), .Q(\ram[9][162] ), .QN(
        n4157) );
  DFFX1_HVT \ram_reg[9][161]  ( .D(n2526), .CLK(clk), .Q(\ram[9][161] ) );
  DFFX1_HVT \ram_reg[9][160]  ( .D(n2525), .CLK(clk), .Q(\ram[9][160] ) );
  DFFX1_HVT \ram_reg[9][159]  ( .D(n2524), .CLK(clk), .Q(\ram[9][159] ) );
  DFFX1_HVT \ram_reg[9][158]  ( .D(n2523), .CLK(clk), .Q(\ram[9][158] ) );
  DFFX1_HVT \ram_reg[9][157]  ( .D(n2522), .CLK(clk), .Q(\ram[9][157] ), .QN(
        n4505) );
  DFFX1_HVT \ram_reg[9][156]  ( .D(n2521), .CLK(clk), .Q(\ram[9][156] ) );
  DFFX1_HVT \ram_reg[9][155]  ( .D(n2520), .CLK(clk), .Q(\ram[9][155] ) );
  DFFX1_HVT \ram_reg[9][154]  ( .D(n2519), .CLK(clk), .Q(\ram[9][154] ) );
  DFFX1_HVT \ram_reg[9][153]  ( .D(n2518), .CLK(clk), .Q(\ram[9][153] ) );
  DFFX1_HVT \ram_reg[9][152]  ( .D(n2517), .CLK(clk), .Q(\ram[9][152] ) );
  DFFX1_HVT \ram_reg[9][151]  ( .D(n2516), .CLK(clk), .Q(\ram[9][151] ) );
  DFFX1_HVT \ram_reg[9][150]  ( .D(n2515), .CLK(clk), .Q(\ram[9][150] ) );
  DFFX1_HVT \ram_reg[9][149]  ( .D(n2514), .CLK(clk), .Q(\ram[9][149] ) );
  DFFX1_HVT \ram_reg[9][148]  ( .D(n2513), .CLK(clk), .Q(\ram[9][148] ) );
  DFFX1_HVT \ram_reg[9][147]  ( .D(n2512), .CLK(clk), .Q(\ram[9][147] ) );
  DFFX1_HVT \ram_reg[9][146]  ( .D(n2511), .CLK(clk), .Q(\ram[9][146] ) );
  DFFX1_HVT \ram_reg[9][145]  ( .D(n2510), .CLK(clk), .Q(\ram[9][145] ) );
  DFFX1_HVT \ram_reg[9][144]  ( .D(n2509), .CLK(clk), .Q(\ram[9][144] ) );
  DFFX1_HVT \ram_reg[9][143]  ( .D(n2508), .CLK(clk), .Q(\ram[9][143] ) );
  DFFX1_HVT \ram_reg[9][142]  ( .D(n2507), .CLK(clk), .Q(\ram[9][142] ) );
  DFFX1_HVT \ram_reg[9][141]  ( .D(n2506), .CLK(clk), .Q(\ram[9][141] ) );
  DFFX1_HVT \ram_reg[9][140]  ( .D(n2505), .CLK(clk), .Q(\ram[9][140] ) );
  DFFX1_HVT \ram_reg[9][139]  ( .D(n2504), .CLK(clk), .Q(\ram[9][139] ) );
  DFFX1_HVT \ram_reg[9][138]  ( .D(n2503), .CLK(clk), .Q(\ram[9][138] ) );
  DFFX1_HVT \ram_reg[9][137]  ( .D(n2502), .CLK(clk), .Q(\ram[9][137] ) );
  DFFX1_HVT \ram_reg[9][136]  ( .D(n2501), .CLK(clk), .Q(\ram[9][136] ), .QN(
        n4170) );
  DFFX1_HVT \ram_reg[9][135]  ( .D(n2500), .CLK(clk), .Q(\ram[9][135] ) );
  DFFX1_HVT \ram_reg[9][134]  ( .D(n2499), .CLK(clk), .Q(\ram[9][134] ) );
  DFFX1_HVT \ram_reg[9][133]  ( .D(n2498), .CLK(clk), .Q(\ram[9][133] ) );
  DFFX1_HVT \ram_reg[9][132]  ( .D(n2497), .CLK(clk), .Q(\ram[9][132] ) );
  DFFX1_HVT \ram_reg[9][131]  ( .D(n2496), .CLK(clk), .Q(\ram[9][131] ) );
  DFFX1_HVT \ram_reg[9][130]  ( .D(n2495), .CLK(clk), .Q(\ram[9][130] ) );
  DFFX1_HVT \ram_reg[9][129]  ( .D(n2494), .CLK(clk), .Q(\ram[9][129] ) );
  DFFX1_HVT \ram_reg[9][128]  ( .D(n2493), .CLK(clk), .Q(\ram[9][128] ) );
  DFFX1_HVT \ram_reg[9][127]  ( .D(n2492), .CLK(clk), .Q(\ram[9][127] ) );
  DFFX1_HVT \ram_reg[9][126]  ( .D(n2491), .CLK(clk), .Q(\ram[9][126] ), .QN(
        n4381) );
  DFFX1_HVT \ram_reg[9][125]  ( .D(n2490), .CLK(clk), .Q(\ram[9][125] ) );
  DFFX1_HVT \ram_reg[9][124]  ( .D(n2489), .CLK(clk), .Q(\ram[9][124] ) );
  DFFX1_HVT \ram_reg[9][123]  ( .D(n2488), .CLK(clk), .Q(\ram[9][123] ) );
  DFFX1_HVT \ram_reg[9][122]  ( .D(n2487), .CLK(clk), .Q(\ram[9][122] ) );
  DFFX1_HVT \ram_reg[9][121]  ( .D(n2486), .CLK(clk), .Q(\ram[9][121] ) );
  DFFX1_HVT \ram_reg[9][120]  ( .D(n2485), .CLK(clk), .Q(\ram[9][120] ) );
  DFFX1_HVT \ram_reg[9][119]  ( .D(n2484), .CLK(clk), .Q(\ram[9][119] ) );
  DFFX1_HVT \ram_reg[9][118]  ( .D(n2483), .CLK(clk), .Q(\ram[9][118] ) );
  DFFX1_HVT \ram_reg[9][117]  ( .D(n2482), .CLK(clk), .Q(\ram[9][117] ) );
  DFFX1_HVT \ram_reg[9][116]  ( .D(n2481), .CLK(clk), .Q(\ram[9][116] ) );
  DFFX1_HVT \ram_reg[9][115]  ( .D(n2480), .CLK(clk), .Q(\ram[9][115] ) );
  DFFX1_HVT \ram_reg[9][114]  ( .D(n2479), .CLK(clk), .Q(\ram[9][114] ) );
  DFFX1_HVT \ram_reg[9][113]  ( .D(n2478), .CLK(clk), .Q(\ram[9][113] ) );
  DFFX1_HVT \ram_reg[9][112]  ( .D(n2477), .CLK(clk), .Q(\ram[9][112] ) );
  DFFX1_HVT \ram_reg[9][111]  ( .D(n2476), .CLK(clk), .Q(\ram[9][111] ) );
  DFFX1_HVT \ram_reg[9][110]  ( .D(n2475), .CLK(clk), .Q(\ram[9][110] ) );
  DFFX1_HVT \ram_reg[9][109]  ( .D(n2474), .CLK(clk), .Q(\ram[9][109] ) );
  DFFX1_HVT \ram_reg[9][108]  ( .D(n2473), .CLK(clk), .Q(\ram[9][108] ) );
  DFFX1_HVT \ram_reg[9][107]  ( .D(n2472), .CLK(clk), .Q(\ram[9][107] ), .QN(
        n4468) );
  DFFX1_HVT \ram_reg[9][106]  ( .D(n2471), .CLK(clk), .Q(\ram[9][106] ) );
  DFFX1_HVT \ram_reg[9][105]  ( .D(n2470), .CLK(clk), .Q(\ram[9][105] ) );
  DFFX1_HVT \ram_reg[9][104]  ( .D(n2469), .CLK(clk), .Q(\ram[9][104] ) );
  DFFX1_HVT \ram_reg[9][103]  ( .D(n2468), .CLK(clk), .Q(\ram[9][103] ) );
  DFFX1_HVT \ram_reg[9][102]  ( .D(n2467), .CLK(clk), .Q(\ram[9][102] ) );
  DFFX1_HVT \ram_reg[9][101]  ( .D(n2466), .CLK(clk), .Q(\ram[9][101] ) );
  DFFX1_HVT \ram_reg[9][100]  ( .D(n2465), .CLK(clk), .Q(\ram[9][100] ) );
  DFFX1_HVT \ram_reg[9][99]  ( .D(n2464), .CLK(clk), .Q(\ram[9][99] ) );
  DFFX1_HVT \ram_reg[9][98]  ( .D(n2463), .CLK(clk), .Q(\ram[9][98] ) );
  DFFX1_HVT \ram_reg[9][97]  ( .D(n2462), .CLK(clk), .Q(\ram[9][97] ) );
  DFFX1_HVT \ram_reg[9][96]  ( .D(n2461), .CLK(clk), .Q(\ram[9][96] ) );
  DFFX1_HVT \ram_reg[9][95]  ( .D(n2460), .CLK(clk), .Q(\ram[9][95] ) );
  DFFX1_HVT \ram_reg[9][94]  ( .D(n2459), .CLK(clk), .Q(\ram[9][94] ) );
  DFFX1_HVT \ram_reg[9][93]  ( .D(n2458), .CLK(clk), .Q(\ram[9][93] ) );
  DFFX1_HVT \ram_reg[9][92]  ( .D(n2457), .CLK(clk), .Q(\ram[9][92] ) );
  DFFX1_HVT \ram_reg[9][91]  ( .D(n2456), .CLK(clk), .Q(\ram[9][91] ) );
  DFFX1_HVT \ram_reg[9][90]  ( .D(n2455), .CLK(clk), .Q(\ram[9][90] ) );
  DFFX1_HVT \ram_reg[9][89]  ( .D(n2454), .CLK(clk), .Q(\ram[9][89] ) );
  DFFX1_HVT \ram_reg[9][88]  ( .D(n2453), .CLK(clk), .Q(\ram[9][88] ) );
  DFFX1_HVT \ram_reg[9][87]  ( .D(n2452), .CLK(clk), .Q(\ram[9][87] ) );
  DFFX1_HVT \ram_reg[9][86]  ( .D(n2451), .CLK(clk), .Q(\ram[9][86] ) );
  DFFX1_HVT \ram_reg[9][85]  ( .D(n2450), .CLK(clk), .Q(\ram[9][85] ) );
  DFFX1_HVT \ram_reg[9][84]  ( .D(n2449), .CLK(clk), .Q(\ram[9][84] ) );
  DFFX1_HVT \ram_reg[9][83]  ( .D(n2448), .CLK(clk), .Q(\ram[9][83] ) );
  DFFX1_HVT \ram_reg[9][82]  ( .D(n2447), .CLK(clk), .Q(\ram[9][82] ), .QN(
        n4654) );
  DFFX1_HVT \ram_reg[9][81]  ( .D(n2446), .CLK(clk), .Q(\ram[9][81] ) );
  DFFX1_HVT \ram_reg[9][80]  ( .D(n2445), .CLK(clk), .Q(\ram[9][80] ) );
  DFFX1_HVT \ram_reg[9][79]  ( .D(n2444), .CLK(clk), .Q(\ram[9][79] ) );
  DFFX1_HVT \ram_reg[9][78]  ( .D(n2443), .CLK(clk), .Q(\ram[9][78] ) );
  DFFX1_HVT \ram_reg[9][77]  ( .D(n2442), .CLK(clk), .Q(\ram[9][77] ) );
  DFFX1_HVT \ram_reg[9][76]  ( .D(n2441), .CLK(clk), .Q(\ram[9][76] ) );
  DFFX1_HVT \ram_reg[9][75]  ( .D(n2440), .CLK(clk), .Q(\ram[9][75] ) );
  DFFX1_HVT \ram_reg[9][74]  ( .D(n2439), .CLK(clk), .Q(\ram[9][74] ) );
  DFFX1_HVT \ram_reg[9][73]  ( .D(n2438), .CLK(clk), .Q(\ram[9][73] ) );
  DFFX1_HVT \ram_reg[9][72]  ( .D(n2437), .CLK(clk), .Q(\ram[9][72] ) );
  DFFX1_HVT \ram_reg[9][71]  ( .D(n2436), .CLK(clk), .Q(\ram[9][71] ) );
  DFFX1_HVT \ram_reg[9][70]  ( .D(n2435), .CLK(clk), .Q(\ram[9][70] ) );
  DFFX1_HVT \ram_reg[9][69]  ( .D(n2434), .CLK(clk), .Q(\ram[9][69] ) );
  DFFX1_HVT \ram_reg[9][68]  ( .D(n2433), .CLK(clk), .Q(\ram[9][68] ) );
  DFFX1_HVT \ram_reg[9][67]  ( .D(n2432), .CLK(clk), .Q(\ram[9][67] ) );
  DFFX1_HVT \ram_reg[9][66]  ( .D(n2431), .CLK(clk), .Q(\ram[9][66] ) );
  DFFX1_HVT \ram_reg[9][65]  ( .D(n2430), .CLK(clk), .Q(\ram[9][65] ) );
  DFFX1_HVT \ram_reg[9][64]  ( .D(n2429), .CLK(clk), .Q(\ram[9][64] ) );
  DFFX1_HVT \ram_reg[9][63]  ( .D(n2428), .CLK(clk), .Q(\ram[9][63] ) );
  DFFX1_HVT \ram_reg[9][62]  ( .D(n2427), .CLK(clk), .Q(\ram[9][62] ), .QN(
        n4488) );
  DFFX1_HVT \ram_reg[9][61]  ( .D(n2426), .CLK(clk), .Q(\ram[9][61] ) );
  DFFX1_HVT \ram_reg[9][60]  ( .D(n2425), .CLK(clk), .Q(\ram[9][60] ) );
  DFFX1_HVT \ram_reg[9][59]  ( .D(n2424), .CLK(clk), .Q(\ram[9][59] ) );
  DFFX1_HVT \ram_reg[9][58]  ( .D(n2423), .CLK(clk), .Q(\ram[9][58] ), .QN(
        n4816) );
  DFFX1_HVT \ram_reg[9][57]  ( .D(n2422), .CLK(clk), .Q(\ram[9][57] ) );
  DFFX1_HVT \ram_reg[9][56]  ( .D(n2421), .CLK(clk), .Q(\ram[9][56] ) );
  DFFX1_HVT \ram_reg[9][55]  ( .D(n2420), .CLK(clk), .Q(\ram[9][55] ), .QN(
        n4490) );
  DFFX1_HVT \ram_reg[9][54]  ( .D(n2419), .CLK(clk), .Q(\ram[9][54] ) );
  DFFX1_HVT \ram_reg[9][53]  ( .D(n2418), .CLK(clk), .Q(\ram[9][53] ) );
  DFFX1_HVT \ram_reg[9][52]  ( .D(n2417), .CLK(clk), .Q(\ram[9][52] ) );
  DFFX1_HVT \ram_reg[9][51]  ( .D(n2416), .CLK(clk), .Q(\ram[9][51] ) );
  DFFX1_HVT \ram_reg[9][50]  ( .D(n2415), .CLK(clk), .Q(\ram[9][50] ) );
  DFFX1_HVT \ram_reg[9][49]  ( .D(n2414), .CLK(clk), .Q(\ram[9][49] ) );
  DFFX1_HVT \ram_reg[9][48]  ( .D(n2413), .CLK(clk), .Q(\ram[9][48] ), .QN(
        n4450) );
  DFFX1_HVT \ram_reg[9][47]  ( .D(n2412), .CLK(clk), .Q(\ram[9][47] ), .QN(
        n4452) );
  DFFX1_HVT \ram_reg[9][46]  ( .D(n2411), .CLK(clk), .Q(\ram[9][46] ), .QN(
        n4454) );
  DFFX1_HVT \ram_reg[9][45]  ( .D(n2410), .CLK(clk), .Q(\ram[9][45] ), .QN(
        n4491) );
  DFFX1_HVT \ram_reg[9][44]  ( .D(n2409), .CLK(clk), .Q(\ram[9][44] ) );
  DFFX1_HVT \ram_reg[9][43]  ( .D(n2408), .CLK(clk), .Q(\ram[9][43] ) );
  DFFX1_HVT \ram_reg[9][42]  ( .D(n2407), .CLK(clk), .Q(\ram[9][42] ) );
  DFFX1_HVT \ram_reg[9][41]  ( .D(n2406), .CLK(clk), .Q(\ram[9][41] ) );
  DFFX1_HVT \ram_reg[9][40]  ( .D(n2405), .CLK(clk), .Q(\ram[9][40] ) );
  DFFX1_HVT \ram_reg[9][39]  ( .D(n2404), .CLK(clk), .Q(\ram[9][39] ) );
  DFFX1_HVT \ram_reg[9][38]  ( .D(n2403), .CLK(clk), .Q(\ram[9][38] ), .QN(
        n1361) );
  DFFX1_HVT \ram_reg[9][37]  ( .D(n2402), .CLK(clk), .Q(\ram[9][37] ), .QN(
        n4751) );
  DFFX1_HVT \ram_reg[9][36]  ( .D(n2401), .CLK(clk), .Q(\ram[9][36] ), .QN(
        n4753) );
  DFFX1_HVT \ram_reg[9][35]  ( .D(n2400), .CLK(clk), .Q(\ram[9][35] ) );
  DFFX1_HVT \ram_reg[9][34]  ( .D(n2399), .CLK(clk), .Q(\ram[9][34] ) );
  DFFX1_HVT \ram_reg[9][33]  ( .D(n2398), .CLK(clk), .Q(\ram[9][33] ) );
  DFFX1_HVT \ram_reg[9][32]  ( .D(n2397), .CLK(clk), .Q(\ram[9][32] ) );
  DFFX1_HVT \ram_reg[9][31]  ( .D(n2396), .CLK(clk), .Q(\ram[9][31] ) );
  DFFX1_HVT \ram_reg[9][30]  ( .D(n2395), .CLK(clk), .Q(\ram[9][30] ) );
  DFFX1_HVT \ram_reg[9][29]  ( .D(n2394), .CLK(clk), .Q(\ram[9][29] ) );
  DFFX1_HVT \ram_reg[9][28]  ( .D(n2393), .CLK(clk), .Q(\ram[9][28] ) );
  DFFX1_HVT \ram_reg[9][27]  ( .D(n2392), .CLK(clk), .Q(\ram[9][27] ) );
  DFFX1_HVT \ram_reg[9][26]  ( .D(n2391), .CLK(clk), .Q(\ram[9][26] ), .QN(
        n4660) );
  DFFX1_HVT \ram_reg[9][25]  ( .D(n2390), .CLK(clk), .Q(\ram[9][25] ) );
  DFFX1_HVT \ram_reg[9][24]  ( .D(n2389), .CLK(clk), .Q(\ram[9][24] ), .QN(
        n4661) );
  DFFX1_HVT \ram_reg[9][23]  ( .D(n2388), .CLK(clk), .Q(\ram[9][23] ) );
  DFFX1_HVT \ram_reg[9][22]  ( .D(n2387), .CLK(clk), .Q(\ram[9][22] ) );
  DFFX1_HVT \ram_reg[9][21]  ( .D(n2386), .CLK(clk), .Q(\ram[9][21] ) );
  DFFX1_HVT \ram_reg[9][20]  ( .D(n2385), .CLK(clk), .Q(\ram[9][20] ), .QN(
        n6482) );
  DFFX1_HVT \ram_reg[9][19]  ( .D(n2384), .CLK(clk), .Q(\ram[9][19] ) );
  DFFX1_HVT \ram_reg[9][18]  ( .D(n2383), .CLK(clk), .Q(\ram[9][18] ) );
  DFFX1_HVT \ram_reg[9][17]  ( .D(n2382), .CLK(clk), .Q(\ram[9][17] ) );
  DFFX1_HVT \ram_reg[9][16]  ( .D(n2381), .CLK(clk), .Q(\ram[9][16] ) );
  DFFX1_HVT \ram_reg[9][15]  ( .D(n2380), .CLK(clk), .Q(\ram[9][15] ) );
  DFFX1_HVT \ram_reg[9][14]  ( .D(n2379), .CLK(clk), .Q(\ram[9][14] ) );
  DFFX1_HVT \ram_reg[9][13]  ( .D(n2378), .CLK(clk), .Q(\ram[9][13] ) );
  DFFX1_HVT \ram_reg[9][12]  ( .D(n2377), .CLK(clk), .Q(\ram[9][12] ) );
  DFFX1_HVT \ram_reg[9][11]  ( .D(n2376), .CLK(clk), .Q(\ram[9][11] ) );
  DFFX1_HVT \ram_reg[9][10]  ( .D(n2375), .CLK(clk), .Q(\ram[9][10] ), .QN(
        n4383) );
  DFFX1_HVT \ram_reg[9][9]  ( .D(n2374), .CLK(clk), .Q(\ram[9][9] ) );
  DFFX1_HVT \ram_reg[9][8]  ( .D(n2373), .CLK(clk), .Q(\ram[9][8] ) );
  DFFX1_HVT \ram_reg[9][7]  ( .D(n2372), .CLK(clk), .Q(\ram[9][7] ) );
  DFFX1_HVT \ram_reg[9][6]  ( .D(n2371), .CLK(clk), .Q(\ram[9][6] ) );
  DFFX1_HVT \ram_reg[9][5]  ( .D(n2370), .CLK(clk), .Q(\ram[9][5] ) );
  DFFX1_HVT \ram_reg[9][4]  ( .D(n2369), .CLK(clk), .Q(\ram[9][4] ) );
  DFFX1_HVT \ram_reg[9][3]  ( .D(n2368), .CLK(clk), .Q(\ram[9][3] ) );
  DFFX1_HVT \ram_reg[9][2]  ( .D(n2367), .CLK(clk), .Q(\ram[9][2] ) );
  DFFX1_HVT \ram_reg[9][1]  ( .D(n2366), .CLK(clk), .Q(\ram[9][1] ) );
  DFFX1_HVT \ram_reg[9][0]  ( .D(n2365), .CLK(clk), .Q(\ram[9][0] ) );
  DFFX1_HVT \ram_reg[8][255]  ( .D(n2364), .CLK(clk), .Q(\ram[8][255] ) );
  DFFX1_HVT \ram_reg[8][254]  ( .D(n2363), .CLK(clk), .Q(\ram[8][254] ) );
  DFFX1_HVT \ram_reg[8][253]  ( .D(n2362), .CLK(clk), .Q(\ram[8][253] ) );
  DFFX1_HVT \ram_reg[8][252]  ( .D(n2361), .CLK(clk), .Q(\ram[8][252] ) );
  DFFX1_HVT \ram_reg[8][251]  ( .D(n2360), .CLK(clk), .Q(\ram[8][251] ) );
  DFFX1_HVT \ram_reg[8][250]  ( .D(n2359), .CLK(clk), .Q(\ram[8][250] ) );
  DFFX1_HVT \ram_reg[8][249]  ( .D(n2358), .CLK(clk), .Q(\ram[8][249] ) );
  DFFX1_HVT \ram_reg[8][248]  ( .D(n2357), .CLK(clk), .Q(\ram[8][248] ) );
  DFFX1_HVT \ram_reg[8][247]  ( .D(n2356), .CLK(clk), .Q(\ram[8][247] ) );
  DFFX1_HVT \ram_reg[8][246]  ( .D(n2355), .CLK(clk), .Q(\ram[8][246] ) );
  DFFX1_HVT \ram_reg[8][245]  ( .D(n2354), .CLK(clk), .Q(\ram[8][245] ) );
  DFFX1_HVT \ram_reg[8][244]  ( .D(n2353), .CLK(clk), .Q(\ram[8][244] ) );
  DFFX1_HVT \ram_reg[8][243]  ( .D(n2352), .CLK(clk), .Q(\ram[8][243] ) );
  DFFX1_HVT \ram_reg[8][242]  ( .D(n2351), .CLK(clk), .Q(\ram[8][242] ) );
  DFFX1_HVT \ram_reg[8][241]  ( .D(n2350), .CLK(clk), .Q(\ram[8][241] ) );
  DFFX1_HVT \ram_reg[8][240]  ( .D(n2349), .CLK(clk), .Q(\ram[8][240] ) );
  DFFX1_HVT \ram_reg[8][239]  ( .D(n2348), .CLK(clk), .Q(\ram[8][239] ) );
  DFFX1_HVT \ram_reg[8][238]  ( .D(n2347), .CLK(clk), .Q(\ram[8][238] ) );
  DFFX1_HVT \ram_reg[8][237]  ( .D(n2346), .CLK(clk), .Q(\ram[8][237] ) );
  DFFX1_HVT \ram_reg[8][236]  ( .D(n2345), .CLK(clk), .Q(\ram[8][236] ) );
  DFFX1_HVT \ram_reg[8][235]  ( .D(n2344), .CLK(clk), .Q(\ram[8][235] ) );
  DFFX1_HVT \ram_reg[8][234]  ( .D(n2343), .CLK(clk), .Q(\ram[8][234] ) );
  DFFX1_HVT \ram_reg[8][233]  ( .D(n2342), .CLK(clk), .Q(\ram[8][233] ) );
  DFFX1_HVT \ram_reg[8][232]  ( .D(n2341), .CLK(clk), .Q(\ram[8][232] ) );
  DFFX1_HVT \ram_reg[8][231]  ( .D(n2340), .CLK(clk), .Q(\ram[8][231] ) );
  DFFX1_HVT \ram_reg[8][230]  ( .D(n2339), .CLK(clk), .Q(\ram[8][230] ) );
  DFFX1_HVT \ram_reg[8][229]  ( .D(n2338), .CLK(clk), .Q(\ram[8][229] ) );
  DFFX1_HVT \ram_reg[8][228]  ( .D(n2337), .CLK(clk), .Q(\ram[8][228] ) );
  DFFX1_HVT \ram_reg[8][227]  ( .D(n2336), .CLK(clk), .Q(\ram[8][227] ) );
  DFFX1_HVT \ram_reg[8][226]  ( .D(n2335), .CLK(clk), .Q(\ram[8][226] ) );
  DFFX1_HVT \ram_reg[8][225]  ( .D(n2334), .CLK(clk), .Q(\ram[8][225] ) );
  DFFX1_HVT \ram_reg[8][224]  ( .D(n2333), .CLK(clk), .Q(\ram[8][224] ) );
  DFFX1_HVT \ram_reg[8][223]  ( .D(n2332), .CLK(clk), .Q(\ram[8][223] ) );
  DFFX1_HVT \ram_reg[8][222]  ( .D(n2331), .CLK(clk), .Q(\ram[8][222] ) );
  DFFX1_HVT \ram_reg[8][221]  ( .D(n2330), .CLK(clk), .Q(\ram[8][221] ) );
  DFFX1_HVT \ram_reg[8][220]  ( .D(n2329), .CLK(clk), .Q(\ram[8][220] ), .QN(
        n5928) );
  DFFX1_HVT \ram_reg[8][219]  ( .D(n2328), .CLK(clk), .Q(\ram[8][219] ) );
  DFFX1_HVT \ram_reg[8][218]  ( .D(n2327), .CLK(clk), .Q(\ram[8][218] ) );
  DFFX1_HVT \ram_reg[8][217]  ( .D(n2326), .CLK(clk), .Q(\ram[8][217] ) );
  DFFX1_HVT \ram_reg[8][216]  ( .D(n2325), .CLK(clk), .Q(\ram[8][216] ) );
  DFFX1_HVT \ram_reg[8][215]  ( .D(n2324), .CLK(clk), .Q(\ram[8][215] ) );
  DFFX1_HVT \ram_reg[8][214]  ( .D(n2323), .CLK(clk), .Q(\ram[8][214] ) );
  DFFX1_HVT \ram_reg[8][213]  ( .D(n2322), .CLK(clk), .Q(\ram[8][213] ) );
  DFFX1_HVT \ram_reg[8][212]  ( .D(n2321), .CLK(clk), .Q(\ram[8][212] ) );
  DFFX1_HVT \ram_reg[8][211]  ( .D(n2320), .CLK(clk), .Q(\ram[8][211] ) );
  DFFX1_HVT \ram_reg[8][210]  ( .D(n2319), .CLK(clk), .Q(\ram[8][210] ) );
  DFFX1_HVT \ram_reg[8][209]  ( .D(n2318), .CLK(clk), .Q(\ram[8][209] ) );
  DFFX1_HVT \ram_reg[8][208]  ( .D(n2317), .CLK(clk), .Q(\ram[8][208] ) );
  DFFX1_HVT \ram_reg[8][207]  ( .D(n2316), .CLK(clk), .Q(\ram[8][207] ) );
  DFFX1_HVT \ram_reg[8][206]  ( .D(n2315), .CLK(clk), .Q(\ram[8][206] ) );
  DFFX1_HVT \ram_reg[8][205]  ( .D(n2314), .CLK(clk), .Q(\ram[8][205] ) );
  DFFX1_HVT \ram_reg[8][204]  ( .D(n2313), .CLK(clk), .Q(\ram[8][204] ) );
  DFFX1_HVT \ram_reg[8][203]  ( .D(n2312), .CLK(clk), .Q(\ram[8][203] ) );
  DFFX1_HVT \ram_reg[8][202]  ( .D(n2311), .CLK(clk), .Q(\ram[8][202] ) );
  DFFX1_HVT \ram_reg[8][201]  ( .D(n2310), .CLK(clk), .Q(\ram[8][201] ) );
  DFFX1_HVT \ram_reg[8][200]  ( .D(n2309), .CLK(clk), .Q(\ram[8][200] ) );
  DFFX1_HVT \ram_reg[8][199]  ( .D(n2308), .CLK(clk), .Q(\ram[8][199] ) );
  DFFX1_HVT \ram_reg[8][198]  ( .D(n2307), .CLK(clk), .Q(\ram[8][198] ) );
  DFFX1_HVT \ram_reg[8][197]  ( .D(n2306), .CLK(clk), .Q(\ram[8][197] ) );
  DFFX1_HVT \ram_reg[8][196]  ( .D(n2305), .CLK(clk), .Q(\ram[8][196] ) );
  DFFX1_HVT \ram_reg[8][195]  ( .D(n2304), .CLK(clk), .Q(\ram[8][195] ) );
  DFFX1_HVT \ram_reg[8][194]  ( .D(n2303), .CLK(clk), .Q(\ram[8][194] ) );
  DFFX1_HVT \ram_reg[8][193]  ( .D(n2302), .CLK(clk), .Q(\ram[8][193] ) );
  DFFX1_HVT \ram_reg[8][192]  ( .D(n2301), .CLK(clk), .Q(\ram[8][192] ) );
  DFFX1_HVT \ram_reg[8][191]  ( .D(n2300), .CLK(clk), .Q(\ram[8][191] ) );
  DFFX1_HVT \ram_reg[8][190]  ( .D(n2299), .CLK(clk), .Q(\ram[8][190] ) );
  DFFX1_HVT \ram_reg[8][189]  ( .D(n2298), .CLK(clk), .Q(\ram[8][189] ) );
  DFFX1_HVT \ram_reg[8][188]  ( .D(n2297), .CLK(clk), .Q(\ram[8][188] ) );
  DFFX1_HVT \ram_reg[8][187]  ( .D(n2296), .CLK(clk), .Q(\ram[8][187] ) );
  DFFX1_HVT \ram_reg[8][186]  ( .D(n2295), .CLK(clk), .Q(\ram[8][186] ) );
  DFFX1_HVT \ram_reg[8][185]  ( .D(n2294), .CLK(clk), .Q(\ram[8][185] ) );
  DFFX1_HVT \ram_reg[8][184]  ( .D(n2293), .CLK(clk), .Q(\ram[8][184] ) );
  DFFX1_HVT \ram_reg[8][183]  ( .D(n2292), .CLK(clk), .Q(\ram[8][183] ) );
  DFFX1_HVT \ram_reg[8][182]  ( .D(n2291), .CLK(clk), .Q(\ram[8][182] ) );
  DFFX1_HVT \ram_reg[8][181]  ( .D(n2290), .CLK(clk), .Q(\ram[8][181] ) );
  DFFX1_HVT \ram_reg[8][180]  ( .D(n2289), .CLK(clk), .Q(\ram[8][180] ) );
  DFFX1_HVT \ram_reg[8][179]  ( .D(n2288), .CLK(clk), .Q(\ram[8][179] ) );
  DFFX1_HVT \ram_reg[8][178]  ( .D(n2287), .CLK(clk), .Q(\ram[8][178] ) );
  DFFX1_HVT \ram_reg[8][177]  ( .D(n2286), .CLK(clk), .Q(\ram[8][177] ) );
  DFFX1_HVT \ram_reg[8][176]  ( .D(n2285), .CLK(clk), .Q(\ram[8][176] ) );
  DFFX1_HVT \ram_reg[8][175]  ( .D(n2284), .CLK(clk), .Q(\ram[8][175] ) );
  DFFX1_HVT \ram_reg[8][174]  ( .D(n2283), .CLK(clk), .Q(\ram[8][174] ) );
  DFFX1_HVT \ram_reg[8][173]  ( .D(n2282), .CLK(clk), .Q(\ram[8][173] ) );
  DFFX1_HVT \ram_reg[8][172]  ( .D(n2281), .CLK(clk), .Q(\ram[8][172] ) );
  DFFX1_HVT \ram_reg[8][171]  ( .D(n2280), .CLK(clk), .Q(\ram[8][171] ) );
  DFFX1_HVT \ram_reg[8][170]  ( .D(n2279), .CLK(clk), .Q(\ram[8][170] ) );
  DFFX1_HVT \ram_reg[8][169]  ( .D(n2278), .CLK(clk), .Q(\ram[8][169] ) );
  DFFX1_HVT \ram_reg[8][168]  ( .D(n2277), .CLK(clk), .Q(\ram[8][168] ) );
  DFFX1_HVT \ram_reg[8][167]  ( .D(n2276), .CLK(clk), .Q(\ram[8][167] ) );
  DFFX1_HVT \ram_reg[8][166]  ( .D(n2275), .CLK(clk), .Q(\ram[8][166] ) );
  DFFX1_HVT \ram_reg[8][165]  ( .D(n2274), .CLK(clk), .Q(\ram[8][165] ) );
  DFFX1_HVT \ram_reg[8][164]  ( .D(n2273), .CLK(clk), .Q(\ram[8][164] ) );
  DFFX1_HVT \ram_reg[8][163]  ( .D(n2272), .CLK(clk), .Q(\ram[8][163] ) );
  DFFX1_HVT \ram_reg[8][162]  ( .D(n2271), .CLK(clk), .Q(\ram[8][162] ) );
  DFFX1_HVT \ram_reg[8][161]  ( .D(n2270), .CLK(clk), .Q(\ram[8][161] ) );
  DFFX1_HVT \ram_reg[8][160]  ( .D(n2269), .CLK(clk), .Q(\ram[8][160] ) );
  DFFX1_HVT \ram_reg[8][159]  ( .D(n2268), .CLK(clk), .Q(\ram[8][159] ) );
  DFFX1_HVT \ram_reg[8][158]  ( .D(n2267), .CLK(clk), .Q(\ram[8][158] ) );
  DFFX1_HVT \ram_reg[8][157]  ( .D(n2266), .CLK(clk), .Q(\ram[8][157] ) );
  DFFX1_HVT \ram_reg[8][156]  ( .D(n2265), .CLK(clk), .Q(\ram[8][156] ) );
  DFFX1_HVT \ram_reg[8][155]  ( .D(n2264), .CLK(clk), .Q(\ram[8][155] ) );
  DFFX1_HVT \ram_reg[8][154]  ( .D(n2263), .CLK(clk), .Q(\ram[8][154] ) );
  DFFX1_HVT \ram_reg[8][153]  ( .D(n2262), .CLK(clk), .Q(\ram[8][153] ) );
  DFFX1_HVT \ram_reg[8][152]  ( .D(n2261), .CLK(clk), .Q(\ram[8][152] ) );
  DFFX1_HVT \ram_reg[8][151]  ( .D(n2260), .CLK(clk), .Q(\ram[8][151] ) );
  DFFX1_HVT \ram_reg[8][150]  ( .D(n2259), .CLK(clk), .Q(\ram[8][150] ) );
  DFFX1_HVT \ram_reg[8][149]  ( .D(n2258), .CLK(clk), .Q(\ram[8][149] ) );
  DFFX1_HVT \ram_reg[8][148]  ( .D(n2257), .CLK(clk), .Q(\ram[8][148] ) );
  DFFX1_HVT \ram_reg[8][147]  ( .D(n2256), .CLK(clk), .Q(\ram[8][147] ) );
  DFFX1_HVT \ram_reg[8][146]  ( .D(n2255), .CLK(clk), .Q(\ram[8][146] ) );
  DFFX1_HVT \ram_reg[8][145]  ( .D(n2254), .CLK(clk), .Q(\ram[8][145] ) );
  DFFX1_HVT \ram_reg[8][144]  ( .D(n2253), .CLK(clk), .Q(\ram[8][144] ) );
  DFFX1_HVT \ram_reg[8][143]  ( .D(n2252), .CLK(clk), .Q(\ram[8][143] ) );
  DFFX1_HVT \ram_reg[8][142]  ( .D(n2251), .CLK(clk), .Q(\ram[8][142] ) );
  DFFX1_HVT \ram_reg[8][141]  ( .D(n2250), .CLK(clk), .Q(\ram[8][141] ) );
  DFFX1_HVT \ram_reg[8][140]  ( .D(n2249), .CLK(clk), .Q(\ram[8][140] ) );
  DFFX1_HVT \ram_reg[8][139]  ( .D(n2248), .CLK(clk), .Q(\ram[8][139] ) );
  DFFX1_HVT \ram_reg[8][138]  ( .D(n2247), .CLK(clk), .Q(\ram[8][138] ) );
  DFFX1_HVT \ram_reg[8][137]  ( .D(n2246), .CLK(clk), .Q(\ram[8][137] ) );
  DFFX1_HVT \ram_reg[8][136]  ( .D(n2245), .CLK(clk), .Q(\ram[8][136] ), .QN(
        n4171) );
  DFFX1_HVT \ram_reg[8][135]  ( .D(n2244), .CLK(clk), .Q(\ram[8][135] ) );
  DFFX1_HVT \ram_reg[8][134]  ( .D(n2243), .CLK(clk), .Q(\ram[8][134] ) );
  DFFX1_HVT \ram_reg[8][133]  ( .D(n2242), .CLK(clk), .Q(\ram[8][133] ) );
  DFFX1_HVT \ram_reg[8][132]  ( .D(n2241), .CLK(clk), .Q(\ram[8][132] ) );
  DFFX1_HVT \ram_reg[8][131]  ( .D(n2240), .CLK(clk), .Q(\ram[8][131] ) );
  DFFX1_HVT \ram_reg[8][130]  ( .D(n2239), .CLK(clk), .Q(\ram[8][130] ) );
  DFFX1_HVT \ram_reg[8][129]  ( .D(n2238), .CLK(clk), .Q(\ram[8][129] ) );
  DFFX1_HVT \ram_reg[8][128]  ( .D(n2237), .CLK(clk), .Q(\ram[8][128] ) );
  DFFX1_HVT \ram_reg[8][127]  ( .D(n2236), .CLK(clk), .Q(\ram[8][127] ) );
  DFFX1_HVT \ram_reg[8][126]  ( .D(n2235), .CLK(clk), .Q(\ram[8][126] ) );
  DFFX1_HVT \ram_reg[8][125]  ( .D(n2234), .CLK(clk), .Q(\ram[8][125] ) );
  DFFX1_HVT \ram_reg[8][124]  ( .D(n2233), .CLK(clk), .Q(\ram[8][124] ) );
  DFFX1_HVT \ram_reg[8][123]  ( .D(n2232), .CLK(clk), .Q(\ram[8][123] ) );
  DFFX1_HVT \ram_reg[8][122]  ( .D(n2231), .CLK(clk), .Q(\ram[8][122] ) );
  DFFX1_HVT \ram_reg[8][121]  ( .D(n2230), .CLK(clk), .Q(\ram[8][121] ) );
  DFFX1_HVT \ram_reg[8][120]  ( .D(n2229), .CLK(clk), .Q(\ram[8][120] ) );
  DFFX1_HVT \ram_reg[8][119]  ( .D(n2228), .CLK(clk), .Q(\ram[8][119] ) );
  DFFX1_HVT \ram_reg[8][118]  ( .D(n2227), .CLK(clk), .Q(\ram[8][118] ) );
  DFFX1_HVT \ram_reg[8][117]  ( .D(n2226), .CLK(clk), .Q(\ram[8][117] ) );
  DFFX1_HVT \ram_reg[8][116]  ( .D(n2225), .CLK(clk), .Q(\ram[8][116] ) );
  DFFX1_HVT \ram_reg[8][115]  ( .D(n2224), .CLK(clk), .Q(\ram[8][115] ) );
  DFFX1_HVT \ram_reg[8][114]  ( .D(n2223), .CLK(clk), .Q(\ram[8][114] ) );
  DFFX1_HVT \ram_reg[8][113]  ( .D(n2222), .CLK(clk), .Q(\ram[8][113] ) );
  DFFX1_HVT \ram_reg[8][112]  ( .D(n2221), .CLK(clk), .Q(\ram[8][112] ) );
  DFFX1_HVT \ram_reg[8][111]  ( .D(n2220), .CLK(clk), .Q(\ram[8][111] ) );
  DFFX1_HVT \ram_reg[8][110]  ( .D(n2219), .CLK(clk), .Q(\ram[8][110] ) );
  DFFX1_HVT \ram_reg[8][109]  ( .D(n2218), .CLK(clk), .Q(\ram[8][109] ) );
  DFFX1_HVT \ram_reg[8][108]  ( .D(n2217), .CLK(clk), .Q(\ram[8][108] ) );
  DFFX1_HVT \ram_reg[8][107]  ( .D(n2216), .CLK(clk), .Q(\ram[8][107] ) );
  DFFX1_HVT \ram_reg[8][106]  ( .D(n2215), .CLK(clk), .Q(\ram[8][106] ) );
  DFFX1_HVT \ram_reg[8][105]  ( .D(n2214), .CLK(clk), .Q(\ram[8][105] ) );
  DFFX1_HVT \ram_reg[8][104]  ( .D(n2213), .CLK(clk), .Q(\ram[8][104] ) );
  DFFX1_HVT \ram_reg[8][103]  ( .D(n2212), .CLK(clk), .Q(\ram[8][103] ) );
  DFFX1_HVT \ram_reg[8][102]  ( .D(n2211), .CLK(clk), .Q(\ram[8][102] ) );
  DFFX1_HVT \ram_reg[8][101]  ( .D(n2210), .CLK(clk), .Q(\ram[8][101] ) );
  DFFX1_HVT \ram_reg[8][100]  ( .D(n2209), .CLK(clk), .Q(\ram[8][100] ) );
  DFFX1_HVT \ram_reg[8][99]  ( .D(n2208), .CLK(clk), .Q(\ram[8][99] ) );
  DFFX1_HVT \ram_reg[8][98]  ( .D(n2207), .CLK(clk), .Q(\ram[8][98] ) );
  DFFX1_HVT \ram_reg[8][97]  ( .D(n2206), .CLK(clk), .Q(\ram[8][97] ) );
  DFFX1_HVT \ram_reg[8][96]  ( .D(n2205), .CLK(clk), .Q(\ram[8][96] ) );
  DFFX1_HVT \ram_reg[8][95]  ( .D(n2204), .CLK(clk), .Q(\ram[8][95] ) );
  DFFX1_HVT \ram_reg[8][94]  ( .D(n2203), .CLK(clk), .Q(\ram[8][94] ) );
  DFFX1_HVT \ram_reg[8][93]  ( .D(n2202), .CLK(clk), .Q(\ram[8][93] ) );
  DFFX1_HVT \ram_reg[8][92]  ( .D(n2201), .CLK(clk), .Q(\ram[8][92] ) );
  DFFX1_HVT \ram_reg[8][91]  ( .D(n2200), .CLK(clk), .Q(\ram[8][91] ) );
  DFFX1_HVT \ram_reg[8][90]  ( .D(n2199), .CLK(clk), .Q(\ram[8][90] ) );
  DFFX1_HVT \ram_reg[8][89]  ( .D(n2198), .CLK(clk), .Q(\ram[8][89] ) );
  DFFX1_HVT \ram_reg[8][88]  ( .D(n2197), .CLK(clk), .Q(\ram[8][88] ) );
  DFFX1_HVT \ram_reg[8][87]  ( .D(n2196), .CLK(clk), .Q(\ram[8][87] ) );
  DFFX1_HVT \ram_reg[8][86]  ( .D(n2195), .CLK(clk), .Q(\ram[8][86] ) );
  DFFX1_HVT \ram_reg[8][85]  ( .D(n2194), .CLK(clk), .Q(\ram[8][85] ) );
  DFFX1_HVT \ram_reg[8][84]  ( .D(n2193), .CLK(clk), .Q(\ram[8][84] ) );
  DFFX1_HVT \ram_reg[8][83]  ( .D(n2192), .CLK(clk), .Q(\ram[8][83] ) );
  DFFX1_HVT \ram_reg[8][82]  ( .D(n2191), .CLK(clk), .Q(\ram[8][82] ) );
  DFFX1_HVT \ram_reg[8][81]  ( .D(n2190), .CLK(clk), .Q(\ram[8][81] ) );
  DFFX1_HVT \ram_reg[8][80]  ( .D(n2189), .CLK(clk), .Q(\ram[8][80] ) );
  DFFX1_HVT \ram_reg[8][79]  ( .D(n2188), .CLK(clk), .Q(\ram[8][79] ) );
  DFFX1_HVT \ram_reg[8][78]  ( .D(n2187), .CLK(clk), .Q(\ram[8][78] ) );
  DFFX1_HVT \ram_reg[8][77]  ( .D(n2186), .CLK(clk), .Q(\ram[8][77] ) );
  DFFX1_HVT \ram_reg[8][76]  ( .D(n2185), .CLK(clk), .Q(\ram[8][76] ) );
  DFFX1_HVT \ram_reg[8][75]  ( .D(n2184), .CLK(clk), .Q(\ram[8][75] ) );
  DFFX1_HVT \ram_reg[8][74]  ( .D(n2183), .CLK(clk), .Q(\ram[8][74] ) );
  DFFX1_HVT \ram_reg[8][73]  ( .D(n2182), .CLK(clk), .Q(\ram[8][73] ) );
  DFFX1_HVT \ram_reg[8][72]  ( .D(n2181), .CLK(clk), .Q(\ram[8][72] ) );
  DFFX1_HVT \ram_reg[8][71]  ( .D(n2180), .CLK(clk), .Q(\ram[8][71] ) );
  DFFX1_HVT \ram_reg[8][70]  ( .D(n2179), .CLK(clk), .Q(\ram[8][70] ) );
  DFFX1_HVT \ram_reg[8][69]  ( .D(n2178), .CLK(clk), .Q(\ram[8][69] ) );
  DFFX1_HVT \ram_reg[8][68]  ( .D(n2177), .CLK(clk), .Q(\ram[8][68] ) );
  DFFX1_HVT \ram_reg[8][67]  ( .D(n2176), .CLK(clk), .Q(\ram[8][67] ) );
  DFFX1_HVT \ram_reg[8][66]  ( .D(n2175), .CLK(clk), .Q(\ram[8][66] ) );
  DFFX1_HVT \ram_reg[8][65]  ( .D(n2174), .CLK(clk), .Q(\ram[8][65] ) );
  DFFX1_HVT \ram_reg[8][64]  ( .D(n2173), .CLK(clk), .Q(\ram[8][64] ) );
  DFFX1_HVT \ram_reg[8][63]  ( .D(n2172), .CLK(clk), .Q(\ram[8][63] ) );
  DFFX1_HVT \ram_reg[8][62]  ( .D(n2171), .CLK(clk), .Q(\ram[8][62] ) );
  DFFX1_HVT \ram_reg[8][61]  ( .D(n2170), .CLK(clk), .Q(\ram[8][61] ) );
  DFFX1_HVT \ram_reg[8][60]  ( .D(n2169), .CLK(clk), .Q(\ram[8][60] ) );
  DFFX1_HVT \ram_reg[8][59]  ( .D(n2168), .CLK(clk), .Q(\ram[8][59] ) );
  DFFX1_HVT \ram_reg[8][58]  ( .D(n2167), .CLK(clk), .QN(n4818) );
  DFFX1_HVT \ram_reg[8][57]  ( .D(n2166), .CLK(clk), .Q(\ram[8][57] ) );
  DFFX1_HVT \ram_reg[8][56]  ( .D(n2165), .CLK(clk), .Q(\ram[8][56] ) );
  DFFX1_HVT \ram_reg[8][55]  ( .D(n2164), .CLK(clk), .Q(\ram[8][55] ) );
  DFFX1_HVT \ram_reg[8][54]  ( .D(n2163), .CLK(clk), .Q(\ram[8][54] ) );
  DFFX1_HVT \ram_reg[8][53]  ( .D(n2162), .CLK(clk), .Q(\ram[8][53] ) );
  DFFX1_HVT \ram_reg[8][52]  ( .D(n2161), .CLK(clk), .Q(\ram[8][52] ) );
  DFFX1_HVT \ram_reg[8][51]  ( .D(n2160), .CLK(clk), .Q(\ram[8][51] ) );
  DFFX1_HVT \ram_reg[8][50]  ( .D(n2159), .CLK(clk), .Q(\ram[8][50] ) );
  DFFX1_HVT \ram_reg[8][49]  ( .D(n2158), .CLK(clk), .Q(\ram[8][49] ) );
  DFFX1_HVT \ram_reg[8][48]  ( .D(n2157), .CLK(clk), .Q(\ram[8][48] ) );
  DFFX1_HVT \ram_reg[8][47]  ( .D(n2156), .CLK(clk), .Q(\ram[8][47] ), .QN(
        n4221) );
  DFFX1_HVT \ram_reg[8][46]  ( .D(n2155), .CLK(clk), .Q(\ram[8][46] ) );
  DFFX1_HVT \ram_reg[8][45]  ( .D(n2154), .CLK(clk), .Q(\ram[8][45] ) );
  DFFX1_HVT \ram_reg[8][44]  ( .D(n2153), .CLK(clk), .Q(\ram[8][44] ) );
  DFFX1_HVT \ram_reg[8][43]  ( .D(n2152), .CLK(clk), .Q(\ram[8][43] ) );
  DFFX1_HVT \ram_reg[8][42]  ( .D(n2151), .CLK(clk), .Q(\ram[8][42] ) );
  DFFX1_HVT \ram_reg[8][41]  ( .D(n2150), .CLK(clk), .Q(\ram[8][41] ) );
  DFFX1_HVT \ram_reg[8][40]  ( .D(n2149), .CLK(clk), .Q(\ram[8][40] ) );
  DFFX1_HVT \ram_reg[8][39]  ( .D(n2148), .CLK(clk), .Q(\ram[8][39] ), .QN(
        n4224) );
  DFFX1_HVT \ram_reg[8][38]  ( .D(n2147), .CLK(clk), .Q(\ram[8][38] ) );
  DFFX1_HVT \ram_reg[8][37]  ( .D(n2146), .CLK(clk), .Q(\ram[8][37] ) );
  DFFX1_HVT \ram_reg[8][36]  ( .D(n2145), .CLK(clk), .Q(\ram[8][36] ) );
  DFFX1_HVT \ram_reg[8][35]  ( .D(n2144), .CLK(clk), .Q(\ram[8][35] ) );
  DFFX1_HVT \ram_reg[8][34]  ( .D(n2143), .CLK(clk), .Q(\ram[8][34] ) );
  DFFX1_HVT \ram_reg[8][33]  ( .D(n2142), .CLK(clk), .Q(\ram[8][33] ) );
  DFFX1_HVT \ram_reg[8][32]  ( .D(n2141), .CLK(clk), .Q(\ram[8][32] ), .QN(
        n4282) );
  DFFX1_HVT \ram_reg[8][31]  ( .D(n2140), .CLK(clk), .Q(\ram[8][31] ) );
  DFFX1_HVT \ram_reg[8][30]  ( .D(n2139), .CLK(clk), .Q(\ram[8][30] ) );
  DFFX1_HVT \ram_reg[8][29]  ( .D(n2138), .CLK(clk), .Q(\ram[8][29] ) );
  DFFX1_HVT \ram_reg[8][28]  ( .D(n2137), .CLK(clk), .Q(\ram[8][28] ) );
  DFFX1_HVT \ram_reg[8][27]  ( .D(n2136), .CLK(clk), .Q(\ram[8][27] ) );
  DFFX1_HVT \ram_reg[8][26]  ( .D(n2135), .CLK(clk), .Q(\ram[8][26] ), .QN(
        n4595) );
  DFFX1_HVT \ram_reg[8][25]  ( .D(n2134), .CLK(clk), .Q(\ram[8][25] ), .QN(
        n4471) );
  DFFX1_HVT \ram_reg[8][24]  ( .D(n2133), .CLK(clk), .Q(\ram[8][24] ) );
  DFFX1_HVT \ram_reg[8][23]  ( .D(n2132), .CLK(clk), .Q(\ram[8][23] ) );
  DFFX1_HVT \ram_reg[8][22]  ( .D(n2131), .CLK(clk), .Q(\ram[8][22] ) );
  DFFX1_HVT \ram_reg[8][21]  ( .D(n2130), .CLK(clk), .Q(\ram[8][21] ) );
  DFFX1_HVT \ram_reg[8][20]  ( .D(n2129), .CLK(clk), .Q(\ram[8][20] ), .QN(
        n6484) );
  DFFX1_HVT \ram_reg[8][19]  ( .D(n2128), .CLK(clk), .Q(\ram[8][19] ) );
  DFFX1_HVT \ram_reg[8][18]  ( .D(n2127), .CLK(clk), .Q(\ram[8][18] ), .QN(
        n4364) );
  DFFX1_HVT \ram_reg[8][17]  ( .D(n2126), .CLK(clk), .Q(\ram[8][17] ), .QN(
        n4366) );
  DFFX1_HVT \ram_reg[8][16]  ( .D(n2125), .CLK(clk), .Q(\ram[8][16] ) );
  DFFX1_HVT \ram_reg[8][15]  ( .D(n2124), .CLK(clk), .Q(\ram[8][15] ), .QN(
        n4437) );
  DFFX1_HVT \ram_reg[8][14]  ( .D(n2123), .CLK(clk), .Q(\ram[8][14] ) );
  DFFX1_HVT \ram_reg[8][13]  ( .D(n2122), .CLK(clk), .Q(\ram[8][13] ) );
  DFFX1_HVT \ram_reg[8][12]  ( .D(n2121), .CLK(clk), .Q(\ram[8][12] ) );
  DFFX1_HVT \ram_reg[8][11]  ( .D(n2120), .CLK(clk), .Q(\ram[8][11] ), .QN(
        n4213) );
  DFFX1_HVT \ram_reg[8][10]  ( .D(n2119), .CLK(clk), .Q(\ram[8][10] ) );
  DFFX1_HVT \ram_reg[8][9]  ( .D(n2118), .CLK(clk), .Q(\ram[8][9] ) );
  DFFX1_HVT \ram_reg[8][8]  ( .D(n2117), .CLK(clk), .Q(\ram[8][8] ) );
  DFFX1_HVT \ram_reg[8][7]  ( .D(n2116), .CLK(clk), .Q(\ram[8][7] ) );
  DFFX1_HVT \ram_reg[8][6]  ( .D(n2115), .CLK(clk), .Q(\ram[8][6] ) );
  DFFX1_HVT \ram_reg[8][5]  ( .D(n2114), .CLK(clk), .Q(\ram[8][5] ) );
  DFFX1_HVT \ram_reg[8][4]  ( .D(n2113), .CLK(clk), .Q(\ram[8][4] ) );
  DFFX1_HVT \ram_reg[8][3]  ( .D(n2112), .CLK(clk), .Q(\ram[8][3] ) );
  DFFX1_HVT \ram_reg[8][2]  ( .D(n2111), .CLK(clk), .Q(\ram[8][2] ) );
  DFFX1_HVT \ram_reg[8][1]  ( .D(n2110), .CLK(clk), .Q(\ram[8][1] ) );
  DFFX1_HVT \ram_reg[8][0]  ( .D(n2109), .CLK(clk), .Q(\ram[8][0] ) );
  DFFX1_HVT \ram_reg[7][255]  ( .D(n2108), .CLK(clk), .Q(\ram[7][255] ) );
  DFFX1_HVT \ram_reg[7][254]  ( .D(n2107), .CLK(clk), .Q(\ram[7][254] ) );
  DFFX1_HVT \ram_reg[7][253]  ( .D(n2106), .CLK(clk), .Q(\ram[7][253] ) );
  DFFX1_HVT \ram_reg[7][252]  ( .D(n2105), .CLK(clk), .Q(\ram[7][252] ) );
  DFFX1_HVT \ram_reg[7][251]  ( .D(n2104), .CLK(clk), .Q(\ram[7][251] ) );
  DFFX1_HVT \ram_reg[7][250]  ( .D(n2103), .CLK(clk), .Q(\ram[7][250] ) );
  DFFX1_HVT \ram_reg[7][249]  ( .D(n2102), .CLK(clk), .Q(\ram[7][249] ) );
  DFFX1_HVT \ram_reg[7][248]  ( .D(n2101), .CLK(clk), .Q(\ram[7][248] ) );
  DFFX1_HVT \ram_reg[7][247]  ( .D(n2100), .CLK(clk), .Q(\ram[7][247] ) );
  DFFX1_HVT \ram_reg[7][246]  ( .D(n2099), .CLK(clk), .Q(\ram[7][246] ) );
  DFFX1_HVT \ram_reg[7][245]  ( .D(n2098), .CLK(clk), .Q(\ram[7][245] ) );
  DFFX1_HVT \ram_reg[7][244]  ( .D(n2097), .CLK(clk), .Q(\ram[7][244] ) );
  DFFX1_HVT \ram_reg[7][243]  ( .D(n2096), .CLK(clk), .Q(\ram[7][243] ) );
  DFFX1_HVT \ram_reg[7][242]  ( .D(n2095), .CLK(clk), .Q(\ram[7][242] ) );
  DFFX1_HVT \ram_reg[7][241]  ( .D(n2094), .CLK(clk), .Q(\ram[7][241] ) );
  DFFX1_HVT \ram_reg[7][240]  ( .D(n2093), .CLK(clk), .Q(\ram[7][240] ) );
  DFFX1_HVT \ram_reg[7][239]  ( .D(n2092), .CLK(clk), .Q(\ram[7][239] ) );
  DFFX1_HVT \ram_reg[7][238]  ( .D(n2091), .CLK(clk), .Q(\ram[7][238] ) );
  DFFX1_HVT \ram_reg[7][237]  ( .D(n2090), .CLK(clk), .Q(\ram[7][237] ) );
  DFFX1_HVT \ram_reg[7][236]  ( .D(n2089), .CLK(clk), .Q(\ram[7][236] ) );
  DFFX1_HVT \ram_reg[7][235]  ( .D(n2088), .CLK(clk), .Q(\ram[7][235] ) );
  DFFX1_HVT \ram_reg[7][234]  ( .D(n2087), .CLK(clk), .Q(\ram[7][234] ), .QN(
        n5716) );
  DFFX1_HVT \ram_reg[7][233]  ( .D(n2086), .CLK(clk), .Q(\ram[7][233] ) );
  DFFX1_HVT \ram_reg[7][232]  ( .D(n2085), .CLK(clk), .Q(\ram[7][232] ) );
  DFFX1_HVT \ram_reg[7][231]  ( .D(n2084), .CLK(clk), .Q(\ram[7][231] ) );
  DFFX1_HVT \ram_reg[7][230]  ( .D(n2083), .CLK(clk), .Q(\ram[7][230] ) );
  DFFX1_HVT \ram_reg[7][229]  ( .D(n2082), .CLK(clk), .Q(\ram[7][229] ) );
  DFFX1_HVT \ram_reg[7][228]  ( .D(n2081), .CLK(clk), .Q(\ram[7][228] ) );
  DFFX1_HVT \ram_reg[7][227]  ( .D(n2080), .CLK(clk), .Q(\ram[7][227] ) );
  DFFX1_HVT \ram_reg[7][226]  ( .D(n2079), .CLK(clk), .Q(\ram[7][226] ) );
  DFFX1_HVT \ram_reg[7][225]  ( .D(n2078), .CLK(clk), .Q(\ram[7][225] ) );
  DFFX1_HVT \ram_reg[7][224]  ( .D(n2077), .CLK(clk), .Q(\ram[7][224] ) );
  DFFX1_HVT \ram_reg[7][223]  ( .D(n2076), .CLK(clk), .Q(\ram[7][223] ) );
  DFFX1_HVT \ram_reg[7][222]  ( .D(n2075), .CLK(clk), .Q(\ram[7][222] ) );
  DFFX1_HVT \ram_reg[7][221]  ( .D(n2074), .CLK(clk), .Q(\ram[7][221] ) );
  DFFX1_HVT \ram_reg[7][220]  ( .D(n2073), .CLK(clk), .Q(\ram[7][220] ) );
  DFFX1_HVT \ram_reg[7][219]  ( .D(n2072), .CLK(clk), .Q(\ram[7][219] ) );
  DFFX1_HVT \ram_reg[7][218]  ( .D(n2071), .CLK(clk), .Q(\ram[7][218] ) );
  DFFX1_HVT \ram_reg[7][217]  ( .D(n2070), .CLK(clk), .Q(\ram[7][217] ) );
  DFFX1_HVT \ram_reg[7][216]  ( .D(n2069), .CLK(clk), .Q(\ram[7][216] ) );
  DFFX1_HVT \ram_reg[7][215]  ( .D(n2068), .CLK(clk), .Q(\ram[7][215] ) );
  DFFX1_HVT \ram_reg[7][214]  ( .D(n2067), .CLK(clk), .Q(\ram[7][214] ) );
  DFFX1_HVT \ram_reg[7][213]  ( .D(n2066), .CLK(clk), .Q(\ram[7][213] ) );
  DFFX1_HVT \ram_reg[7][212]  ( .D(n2065), .CLK(clk), .Q(\ram[7][212] ) );
  DFFX1_HVT \ram_reg[7][211]  ( .D(n2064), .CLK(clk), .Q(\ram[7][211] ) );
  DFFX1_HVT \ram_reg[7][210]  ( .D(n2063), .CLK(clk), .Q(\ram[7][210] ) );
  DFFX1_HVT \ram_reg[7][209]  ( .D(n2062), .CLK(clk), .Q(\ram[7][209] ) );
  DFFX1_HVT \ram_reg[7][208]  ( .D(n2061), .CLK(clk), .Q(\ram[7][208] ) );
  DFFX1_HVT \ram_reg[7][207]  ( .D(n2060), .CLK(clk), .Q(\ram[7][207] ) );
  DFFX1_HVT \ram_reg[7][206]  ( .D(n2059), .CLK(clk), .Q(\ram[7][206] ), .QN(
        n39) );
  DFFX1_HVT \ram_reg[7][205]  ( .D(n2058), .CLK(clk), .Q(\ram[7][205] ) );
  DFFX1_HVT \ram_reg[7][204]  ( .D(n2057), .CLK(clk), .Q(\ram[7][204] ) );
  DFFX1_HVT \ram_reg[7][203]  ( .D(n2056), .CLK(clk), .Q(\ram[7][203] ) );
  DFFX1_HVT \ram_reg[7][202]  ( .D(n2055), .CLK(clk), .Q(\ram[7][202] ) );
  DFFX1_HVT \ram_reg[7][201]  ( .D(n2054), .CLK(clk), .Q(\ram[7][201] ) );
  DFFX1_HVT \ram_reg[7][200]  ( .D(n2053), .CLK(clk), .Q(\ram[7][200] ) );
  DFFX1_HVT \ram_reg[7][199]  ( .D(n2052), .CLK(clk), .Q(\ram[7][199] ) );
  DFFX1_HVT \ram_reg[7][198]  ( .D(n2051), .CLK(clk), .Q(\ram[7][198] ) );
  DFFX1_HVT \ram_reg[7][197]  ( .D(n2050), .CLK(clk), .Q(\ram[7][197] ) );
  DFFX1_HVT \ram_reg[7][196]  ( .D(n2049), .CLK(clk), .Q(\ram[7][196] ) );
  DFFX1_HVT \ram_reg[7][195]  ( .D(n2048), .CLK(clk), .Q(\ram[7][195] ) );
  DFFX1_HVT \ram_reg[7][194]  ( .D(n2047), .CLK(clk), .Q(\ram[7][194] ) );
  DFFX1_HVT \ram_reg[7][193]  ( .D(n2046), .CLK(clk), .Q(\ram[7][193] ) );
  DFFX1_HVT \ram_reg[7][192]  ( .D(n2045), .CLK(clk), .Q(\ram[7][192] ) );
  DFFX1_HVT \ram_reg[7][191]  ( .D(n2044), .CLK(clk), .Q(\ram[7][191] ) );
  DFFX1_HVT \ram_reg[7][190]  ( .D(n2043), .CLK(clk), .Q(\ram[7][190] ) );
  DFFX1_HVT \ram_reg[7][189]  ( .D(n2042), .CLK(clk), .Q(\ram[7][189] ) );
  DFFX1_HVT \ram_reg[7][188]  ( .D(n2041), .CLK(clk), .Q(\ram[7][188] ) );
  DFFX1_HVT \ram_reg[7][187]  ( .D(n2040), .CLK(clk), .Q(\ram[7][187] ) );
  DFFX1_HVT \ram_reg[7][186]  ( .D(n2039), .CLK(clk), .Q(\ram[7][186] ) );
  DFFX1_HVT \ram_reg[7][185]  ( .D(n2038), .CLK(clk), .Q(\ram[7][185] ) );
  DFFX1_HVT \ram_reg[7][184]  ( .D(n2037), .CLK(clk), .Q(\ram[7][184] ) );
  DFFX1_HVT \ram_reg[7][183]  ( .D(n2036), .CLK(clk), .Q(\ram[7][183] ) );
  DFFX1_HVT \ram_reg[7][182]  ( .D(n2035), .CLK(clk), .Q(\ram[7][182] ) );
  DFFX1_HVT \ram_reg[7][181]  ( .D(n2034), .CLK(clk), .Q(\ram[7][181] ) );
  DFFX1_HVT \ram_reg[7][180]  ( .D(n2033), .CLK(clk), .Q(\ram[7][180] ) );
  DFFX1_HVT \ram_reg[7][179]  ( .D(n2032), .CLK(clk), .Q(\ram[7][179] ) );
  DFFX1_HVT \ram_reg[7][178]  ( .D(n2031), .CLK(clk), .Q(\ram[7][178] ) );
  DFFX1_HVT \ram_reg[7][177]  ( .D(n2030), .CLK(clk), .Q(\ram[7][177] ) );
  DFFX1_HVT \ram_reg[7][176]  ( .D(n2029), .CLK(clk), .Q(\ram[7][176] ) );
  DFFX1_HVT \ram_reg[7][175]  ( .D(n2028), .CLK(clk), .Q(\ram[7][175] ) );
  DFFX1_HVT \ram_reg[7][174]  ( .D(n2027), .CLK(clk), .Q(\ram[7][174] ) );
  DFFX1_HVT \ram_reg[7][173]  ( .D(n2026), .CLK(clk), .Q(\ram[7][173] ) );
  DFFX1_HVT \ram_reg[7][172]  ( .D(n2025), .CLK(clk), .Q(\ram[7][172] ) );
  DFFX1_HVT \ram_reg[7][171]  ( .D(n2024), .CLK(clk), .Q(\ram[7][171] ) );
  DFFX1_HVT \ram_reg[7][170]  ( .D(n2023), .CLK(clk), .Q(\ram[7][170] ) );
  DFFX1_HVT \ram_reg[7][169]  ( .D(n2022), .CLK(clk), .Q(\ram[7][169] ) );
  DFFX1_HVT \ram_reg[7][168]  ( .D(n2021), .CLK(clk), .Q(\ram[7][168] ) );
  DFFX1_HVT \ram_reg[7][167]  ( .D(n2020), .CLK(clk), .Q(\ram[7][167] ) );
  DFFX1_HVT \ram_reg[7][166]  ( .D(n2019), .CLK(clk), .Q(\ram[7][166] ) );
  DFFX1_HVT \ram_reg[7][165]  ( .D(n2018), .CLK(clk), .Q(\ram[7][165] ) );
  DFFX1_HVT \ram_reg[7][164]  ( .D(n2017), .CLK(clk), .Q(\ram[7][164] ) );
  DFFX1_HVT \ram_reg[7][163]  ( .D(n2016), .CLK(clk), .Q(\ram[7][163] ) );
  DFFX1_HVT \ram_reg[7][162]  ( .D(n2015), .CLK(clk), .Q(\ram[7][162] ) );
  DFFX1_HVT \ram_reg[7][161]  ( .D(n2014), .CLK(clk), .Q(\ram[7][161] ) );
  DFFX1_HVT \ram_reg[7][160]  ( .D(n2013), .CLK(clk), .Q(\ram[7][160] ) );
  DFFX1_HVT \ram_reg[7][159]  ( .D(n2012), .CLK(clk), .Q(\ram[7][159] ) );
  DFFX1_HVT \ram_reg[7][158]  ( .D(n2011), .CLK(clk), .Q(\ram[7][158] ) );
  DFFX1_HVT \ram_reg[7][157]  ( .D(n2010), .CLK(clk), .Q(\ram[7][157] ) );
  DFFX1_HVT \ram_reg[7][156]  ( .D(n2009), .CLK(clk), .Q(\ram[7][156] ) );
  DFFX1_HVT \ram_reg[7][155]  ( .D(n2008), .CLK(clk), .Q(\ram[7][155] ) );
  DFFX1_HVT \ram_reg[7][154]  ( .D(n2007), .CLK(clk), .Q(\ram[7][154] ) );
  DFFX1_HVT \ram_reg[7][153]  ( .D(n2006), .CLK(clk), .Q(\ram[7][153] ) );
  DFFX1_HVT \ram_reg[7][152]  ( .D(n2005), .CLK(clk), .Q(\ram[7][152] ) );
  DFFX1_HVT \ram_reg[7][151]  ( .D(n2004), .CLK(clk), .Q(\ram[7][151] ) );
  DFFX1_HVT \ram_reg[7][150]  ( .D(n2003), .CLK(clk), .Q(\ram[7][150] ) );
  DFFX1_HVT \ram_reg[7][149]  ( .D(n2002), .CLK(clk), .Q(\ram[7][149] ) );
  DFFX1_HVT \ram_reg[7][148]  ( .D(n2001), .CLK(clk), .Q(\ram[7][148] ) );
  DFFX1_HVT \ram_reg[7][147]  ( .D(n2000), .CLK(clk), .Q(\ram[7][147] ) );
  DFFX1_HVT \ram_reg[7][146]  ( .D(n1999), .CLK(clk), .Q(\ram[7][146] ) );
  DFFX1_HVT \ram_reg[7][145]  ( .D(n1998), .CLK(clk), .Q(\ram[7][145] ) );
  DFFX1_HVT \ram_reg[7][144]  ( .D(n1997), .CLK(clk), .Q(\ram[7][144] ) );
  DFFX1_HVT \ram_reg[7][143]  ( .D(n1996), .CLK(clk), .Q(\ram[7][143] ) );
  DFFX1_HVT \ram_reg[7][142]  ( .D(n1995), .CLK(clk), .Q(\ram[7][142] ) );
  DFFX1_HVT \ram_reg[7][141]  ( .D(n1994), .CLK(clk), .Q(\ram[7][141] ) );
  DFFX1_HVT \ram_reg[7][140]  ( .D(n1993), .CLK(clk), .Q(\ram[7][140] ) );
  DFFX1_HVT \ram_reg[7][139]  ( .D(n1992), .CLK(clk), .Q(\ram[7][139] ) );
  DFFX1_HVT \ram_reg[7][138]  ( .D(n1991), .CLK(clk), .Q(\ram[7][138] ) );
  DFFX1_HVT \ram_reg[7][137]  ( .D(n1990), .CLK(clk), .Q(\ram[7][137] ) );
  DFFX1_HVT \ram_reg[7][136]  ( .D(n1989), .CLK(clk), .Q(\ram[7][136] ) );
  DFFX1_HVT \ram_reg[7][135]  ( .D(n1988), .CLK(clk), .Q(\ram[7][135] ) );
  DFFX1_HVT \ram_reg[7][134]  ( .D(n1987), .CLK(clk), .Q(\ram[7][134] ) );
  DFFX1_HVT \ram_reg[7][133]  ( .D(n1986), .CLK(clk), .Q(\ram[7][133] ) );
  DFFX1_HVT \ram_reg[7][132]  ( .D(n1985), .CLK(clk), .Q(\ram[7][132] ) );
  DFFX1_HVT \ram_reg[7][131]  ( .D(n1984), .CLK(clk), .Q(\ram[7][131] ) );
  DFFX1_HVT \ram_reg[7][130]  ( .D(n1983), .CLK(clk), .Q(\ram[7][130] ) );
  DFFX1_HVT \ram_reg[7][129]  ( .D(n1982), .CLK(clk), .Q(\ram[7][129] ) );
  DFFX1_HVT \ram_reg[7][128]  ( .D(n1981), .CLK(clk), .Q(\ram[7][128] ) );
  DFFX1_HVT \ram_reg[7][127]  ( .D(n1980), .CLK(clk), .Q(\ram[7][127] ) );
  DFFX1_HVT \ram_reg[7][126]  ( .D(n1979), .CLK(clk), .Q(\ram[7][126] ) );
  DFFX1_HVT \ram_reg[7][125]  ( .D(n1978), .CLK(clk), .Q(\ram[7][125] ) );
  DFFX1_HVT \ram_reg[7][124]  ( .D(n1977), .CLK(clk), .Q(\ram[7][124] ) );
  DFFX1_HVT \ram_reg[7][123]  ( .D(n1976), .CLK(clk), .Q(\ram[7][123] ) );
  DFFX1_HVT \ram_reg[7][122]  ( .D(n1975), .CLK(clk), .Q(\ram[7][122] ) );
  DFFX1_HVT \ram_reg[7][121]  ( .D(n1974), .CLK(clk), .Q(\ram[7][121] ) );
  DFFX1_HVT \ram_reg[7][120]  ( .D(n1973), .CLK(clk), .Q(\ram[7][120] ) );
  DFFX1_HVT \ram_reg[7][119]  ( .D(n1972), .CLK(clk), .Q(\ram[7][119] ) );
  DFFX1_HVT \ram_reg[7][118]  ( .D(n1971), .CLK(clk), .Q(\ram[7][118] ) );
  DFFX1_HVT \ram_reg[7][117]  ( .D(n1970), .CLK(clk), .Q(\ram[7][117] ) );
  DFFX1_HVT \ram_reg[7][116]  ( .D(n1969), .CLK(clk), .Q(\ram[7][116] ) );
  DFFX1_HVT \ram_reg[7][115]  ( .D(n1968), .CLK(clk), .Q(\ram[7][115] ) );
  DFFX1_HVT \ram_reg[7][114]  ( .D(n1967), .CLK(clk), .Q(\ram[7][114] ) );
  DFFX1_HVT \ram_reg[7][113]  ( .D(n1966), .CLK(clk), .Q(\ram[7][113] ) );
  DFFX1_HVT \ram_reg[7][112]  ( .D(n1965), .CLK(clk), .Q(\ram[7][112] ) );
  DFFX1_HVT \ram_reg[7][111]  ( .D(n1964), .CLK(clk), .Q(\ram[7][111] ) );
  DFFX1_HVT \ram_reg[7][110]  ( .D(n1963), .CLK(clk), .Q(\ram[7][110] ) );
  DFFX1_HVT \ram_reg[7][109]  ( .D(n1962), .CLK(clk), .Q(\ram[7][109] ) );
  DFFX1_HVT \ram_reg[7][108]  ( .D(n1961), .CLK(clk), .Q(\ram[7][108] ) );
  DFFX1_HVT \ram_reg[7][107]  ( .D(n1960), .CLK(clk), .Q(\ram[7][107] ) );
  DFFX1_HVT \ram_reg[7][106]  ( .D(n1959), .CLK(clk), .Q(\ram[7][106] ) );
  DFFX1_HVT \ram_reg[7][105]  ( .D(n1958), .CLK(clk), .Q(\ram[7][105] ) );
  DFFX1_HVT \ram_reg[7][104]  ( .D(n1957), .CLK(clk), .Q(\ram[7][104] ) );
  DFFX1_HVT \ram_reg[7][103]  ( .D(n1956), .CLK(clk), .Q(\ram[7][103] ) );
  DFFX1_HVT \ram_reg[7][102]  ( .D(n1955), .CLK(clk), .Q(\ram[7][102] ) );
  DFFX1_HVT \ram_reg[7][101]  ( .D(n1954), .CLK(clk), .Q(\ram[7][101] ) );
  DFFX1_HVT \ram_reg[7][100]  ( .D(n1953), .CLK(clk), .Q(\ram[7][100] ) );
  DFFX1_HVT \ram_reg[7][99]  ( .D(n1952), .CLK(clk), .Q(\ram[7][99] ) );
  DFFX1_HVT \ram_reg[7][98]  ( .D(n1951), .CLK(clk), .Q(\ram[7][98] ) );
  DFFX1_HVT \ram_reg[7][97]  ( .D(n1950), .CLK(clk), .Q(\ram[7][97] ) );
  DFFX1_HVT \ram_reg[7][96]  ( .D(n1949), .CLK(clk), .Q(\ram[7][96] ) );
  DFFX1_HVT \ram_reg[7][95]  ( .D(n1948), .CLK(clk), .Q(\ram[7][95] ) );
  DFFX1_HVT \ram_reg[7][94]  ( .D(n1947), .CLK(clk), .Q(\ram[7][94] ) );
  DFFX1_HVT \ram_reg[7][93]  ( .D(n1946), .CLK(clk), .Q(\ram[7][93] ) );
  DFFX1_HVT \ram_reg[7][92]  ( .D(n1945), .CLK(clk), .Q(\ram[7][92] ) );
  DFFX1_HVT \ram_reg[7][91]  ( .D(n1944), .CLK(clk), .Q(\ram[7][91] ) );
  DFFX1_HVT \ram_reg[7][90]  ( .D(n1943), .CLK(clk), .Q(\ram[7][90] ) );
  DFFX1_HVT \ram_reg[7][89]  ( .D(n1942), .CLK(clk), .Q(\ram[7][89] ) );
  DFFX1_HVT \ram_reg[7][88]  ( .D(n1941), .CLK(clk), .Q(\ram[7][88] ) );
  DFFX1_HVT \ram_reg[7][87]  ( .D(n1940), .CLK(clk), .Q(\ram[7][87] ) );
  DFFX1_HVT \ram_reg[7][86]  ( .D(n1939), .CLK(clk), .Q(\ram[7][86] ) );
  DFFX1_HVT \ram_reg[7][85]  ( .D(n1938), .CLK(clk), .Q(\ram[7][85] ) );
  DFFX1_HVT \ram_reg[7][84]  ( .D(n1937), .CLK(clk), .Q(\ram[7][84] ) );
  DFFX1_HVT \ram_reg[7][83]  ( .D(n1936), .CLK(clk), .Q(\ram[7][83] ) );
  DFFX1_HVT \ram_reg[7][82]  ( .D(n1935), .CLK(clk), .Q(\ram[7][82] ) );
  DFFX1_HVT \ram_reg[7][81]  ( .D(n1934), .CLK(clk), .Q(\ram[7][81] ) );
  DFFX1_HVT \ram_reg[7][80]  ( .D(n1933), .CLK(clk), .Q(\ram[7][80] ) );
  DFFX1_HVT \ram_reg[7][79]  ( .D(n1932), .CLK(clk), .Q(\ram[7][79] ) );
  DFFX1_HVT \ram_reg[7][78]  ( .D(n1931), .CLK(clk), .Q(\ram[7][78] ) );
  DFFX1_HVT \ram_reg[7][77]  ( .D(n1930), .CLK(clk), .Q(\ram[7][77] ) );
  DFFX1_HVT \ram_reg[7][76]  ( .D(n1929), .CLK(clk), .Q(\ram[7][76] ) );
  DFFX1_HVT \ram_reg[7][75]  ( .D(n1928), .CLK(clk), .Q(\ram[7][75] ) );
  DFFX1_HVT \ram_reg[7][74]  ( .D(n1927), .CLK(clk), .Q(\ram[7][74] ) );
  DFFX1_HVT \ram_reg[7][73]  ( .D(n1926), .CLK(clk), .Q(\ram[7][73] ) );
  DFFX1_HVT \ram_reg[7][72]  ( .D(n1925), .CLK(clk), .Q(\ram[7][72] ) );
  DFFX1_HVT \ram_reg[7][71]  ( .D(n1924), .CLK(clk), .Q(\ram[7][71] ) );
  DFFX1_HVT \ram_reg[7][70]  ( .D(n1923), .CLK(clk), .Q(\ram[7][70] ) );
  DFFX1_HVT \ram_reg[7][69]  ( .D(n1922), .CLK(clk), .Q(\ram[7][69] ) );
  DFFX1_HVT \ram_reg[7][68]  ( .D(n1921), .CLK(clk), .Q(\ram[7][68] ) );
  DFFX1_HVT \ram_reg[7][67]  ( .D(n1920), .CLK(clk), .Q(\ram[7][67] ) );
  DFFX1_HVT \ram_reg[7][66]  ( .D(n1919), .CLK(clk), .Q(\ram[7][66] ) );
  DFFX1_HVT \ram_reg[7][65]  ( .D(n1918), .CLK(clk), .Q(\ram[7][65] ) );
  DFFX1_HVT \ram_reg[7][64]  ( .D(n1917), .CLK(clk), .Q(\ram[7][64] ) );
  DFFX1_HVT \ram_reg[7][63]  ( .D(n1916), .CLK(clk), .Q(\ram[7][63] ) );
  DFFX1_HVT \ram_reg[7][62]  ( .D(n1915), .CLK(clk), .Q(\ram[7][62] ) );
  DFFX1_HVT \ram_reg[7][61]  ( .D(n1914), .CLK(clk), .Q(\ram[7][61] ) );
  DFFX1_HVT \ram_reg[7][60]  ( .D(n1913), .CLK(clk), .Q(\ram[7][60] ) );
  DFFX1_HVT \ram_reg[7][59]  ( .D(n1912), .CLK(clk), .Q(\ram[7][59] ) );
  DFFX1_HVT \ram_reg[7][58]  ( .D(n1911), .CLK(clk), .Q(\ram[7][58] ) );
  DFFX1_HVT \ram_reg[7][57]  ( .D(n1910), .CLK(clk), .Q(\ram[7][57] ) );
  DFFX1_HVT \ram_reg[7][56]  ( .D(n1909), .CLK(clk), .Q(\ram[7][56] ) );
  DFFX1_HVT \ram_reg[7][55]  ( .D(n1908), .CLK(clk), .Q(\ram[7][55] ) );
  DFFX1_HVT \ram_reg[7][54]  ( .D(n1907), .CLK(clk), .Q(\ram[7][54] ), .QN(
        n4804) );
  DFFX1_HVT \ram_reg[7][53]  ( .D(n1906), .CLK(clk), .Q(\ram[7][53] ) );
  DFFX1_HVT \ram_reg[7][52]  ( .D(n1905), .CLK(clk), .Q(\ram[7][52] ) );
  DFFX1_HVT \ram_reg[7][51]  ( .D(n1904), .CLK(clk), .Q(\ram[7][51] ) );
  DFFX1_HVT \ram_reg[7][50]  ( .D(n1903), .CLK(clk), .Q(\ram[7][50] ) );
  DFFX1_HVT \ram_reg[7][49]  ( .D(n1902), .CLK(clk), .Q(\ram[7][49] ) );
  DFFX1_HVT \ram_reg[7][48]  ( .D(n1901), .CLK(clk), .Q(\ram[7][48] ) );
  DFFX1_HVT \ram_reg[7][47]  ( .D(n1900), .CLK(clk), .Q(\ram[7][47] ) );
  DFFX1_HVT \ram_reg[7][46]  ( .D(n1899), .CLK(clk), .Q(\ram[7][46] ) );
  DFFX1_HVT \ram_reg[7][45]  ( .D(n1898), .CLK(clk), .Q(\ram[7][45] ) );
  DFFX1_HVT \ram_reg[7][44]  ( .D(n1897), .CLK(clk), .Q(\ram[7][44] ) );
  DFFX1_HVT \ram_reg[7][43]  ( .D(n1896), .CLK(clk), .Q(\ram[7][43] ) );
  DFFX1_HVT \ram_reg[7][42]  ( .D(n1895), .CLK(clk), .Q(\ram[7][42] ) );
  DFFX1_HVT \ram_reg[7][41]  ( .D(n1894), .CLK(clk), .Q(\ram[7][41] ) );
  DFFX1_HVT \ram_reg[7][40]  ( .D(n1893), .CLK(clk), .Q(\ram[7][40] ) );
  DFFX1_HVT \ram_reg[7][39]  ( .D(n1892), .CLK(clk), .Q(\ram[7][39] ) );
  DFFX1_HVT \ram_reg[7][38]  ( .D(n1891), .CLK(clk), .Q(\ram[7][38] ) );
  DFFX1_HVT \ram_reg[7][37]  ( .D(n1890), .CLK(clk), .Q(\ram[7][37] ) );
  DFFX1_HVT \ram_reg[7][36]  ( .D(n1889), .CLK(clk), .Q(\ram[7][36] ) );
  DFFX1_HVT \ram_reg[7][35]  ( .D(n1888), .CLK(clk), .Q(\ram[7][35] ) );
  DFFX1_HVT \ram_reg[7][34]  ( .D(n1887), .CLK(clk), .Q(\ram[7][34] ) );
  DFFX1_HVT \ram_reg[7][33]  ( .D(n1886), .CLK(clk), .Q(\ram[7][33] ) );
  DFFX1_HVT \ram_reg[7][32]  ( .D(n1885), .CLK(clk), .Q(\ram[7][32] ) );
  DFFX1_HVT \ram_reg[7][31]  ( .D(n1884), .CLK(clk), .Q(\ram[7][31] ) );
  DFFX1_HVT \ram_reg[7][30]  ( .D(n1883), .CLK(clk), .Q(\ram[7][30] ) );
  DFFX1_HVT \ram_reg[7][29]  ( .D(n1882), .CLK(clk), .Q(\ram[7][29] ) );
  DFFX1_HVT \ram_reg[7][28]  ( .D(n1881), .CLK(clk), .Q(\ram[7][28] ) );
  DFFX1_HVT \ram_reg[7][27]  ( .D(n1880), .CLK(clk), .Q(\ram[7][27] ) );
  DFFX1_HVT \ram_reg[7][26]  ( .D(n1879), .CLK(clk), .Q(\ram[7][26] ) );
  DFFX1_HVT \ram_reg[7][25]  ( .D(n1878), .CLK(clk), .Q(\ram[7][25] ) );
  DFFX1_HVT \ram_reg[7][24]  ( .D(n1877), .CLK(clk), .Q(\ram[7][24] ) );
  DFFX1_HVT \ram_reg[7][23]  ( .D(n1876), .CLK(clk), .Q(\ram[7][23] ) );
  DFFX1_HVT \ram_reg[7][22]  ( .D(n1875), .CLK(clk), .Q(\ram[7][22] ) );
  DFFX1_HVT \ram_reg[7][21]  ( .D(n1874), .CLK(clk), .Q(\ram[7][21] ) );
  DFFX1_HVT \ram_reg[7][20]  ( .D(n1873), .CLK(clk), .Q(\ram[7][20] ), .QN(
        n6552) );
  DFFX1_HVT \ram_reg[7][19]  ( .D(n1872), .CLK(clk), .Q(\ram[7][19] ) );
  DFFX1_HVT \ram_reg[7][18]  ( .D(n1871), .CLK(clk), .Q(\ram[7][18] ) );
  DFFX1_HVT \ram_reg[7][17]  ( .D(n1870), .CLK(clk), .Q(\ram[7][17] ) );
  DFFX1_HVT \ram_reg[7][16]  ( .D(n1869), .CLK(clk), .Q(\ram[7][16] ) );
  DFFX1_HVT \ram_reg[7][15]  ( .D(n1868), .CLK(clk), .Q(\ram[7][15] ) );
  DFFX1_HVT \ram_reg[7][14]  ( .D(n1867), .CLK(clk), .Q(\ram[7][14] ) );
  DFFX1_HVT \ram_reg[7][13]  ( .D(n1866), .CLK(clk), .Q(\ram[7][13] ) );
  DFFX1_HVT \ram_reg[7][12]  ( .D(n1865), .CLK(clk), .Q(\ram[7][12] ) );
  DFFX1_HVT \ram_reg[7][11]  ( .D(n1864), .CLK(clk), .Q(\ram[7][11] ) );
  DFFX1_HVT \ram_reg[7][10]  ( .D(n1863), .CLK(clk), .Q(\ram[7][10] ) );
  DFFX1_HVT \ram_reg[7][9]  ( .D(n1862), .CLK(clk), .Q(\ram[7][9] ) );
  DFFX1_HVT \ram_reg[7][8]  ( .D(n1861), .CLK(clk), .Q(\ram[7][8] ) );
  DFFX1_HVT \ram_reg[7][7]  ( .D(n1860), .CLK(clk), .Q(\ram[7][7] ) );
  DFFX1_HVT \ram_reg[7][6]  ( .D(n1859), .CLK(clk), .Q(\ram[7][6] ) );
  DFFX1_HVT \ram_reg[7][5]  ( .D(n1858), .CLK(clk), .Q(\ram[7][5] ) );
  DFFX1_HVT \ram_reg[7][4]  ( .D(n1857), .CLK(clk), .Q(\ram[7][4] ) );
  DFFX1_HVT \ram_reg[7][3]  ( .D(n1856), .CLK(clk), .Q(\ram[7][3] ) );
  DFFX1_HVT \ram_reg[7][2]  ( .D(n1855), .CLK(clk), .Q(\ram[7][2] ) );
  DFFX1_HVT \ram_reg[7][1]  ( .D(n1854), .CLK(clk), .Q(\ram[7][1] ) );
  DFFX1_HVT \ram_reg[7][0]  ( .D(n1853), .CLK(clk), .Q(\ram[7][0] ) );
  DFFX1_HVT \ram_reg[6][255]  ( .D(n1852), .CLK(clk), .Q(\ram[6][255] ) );
  DFFX1_HVT \ram_reg[6][254]  ( .D(n1851), .CLK(clk), .Q(\ram[6][254] ) );
  DFFX1_HVT \ram_reg[6][253]  ( .D(n1850), .CLK(clk), .Q(\ram[6][253] ) );
  DFFX1_HVT \ram_reg[6][252]  ( .D(n1849), .CLK(clk), .Q(\ram[6][252] ) );
  DFFX1_HVT \ram_reg[6][251]  ( .D(n1848), .CLK(clk), .Q(\ram[6][251] ) );
  DFFX1_HVT \ram_reg[6][250]  ( .D(n1847), .CLK(clk), .Q(\ram[6][250] ) );
  DFFX1_HVT \ram_reg[6][249]  ( .D(n1846), .CLK(clk), .Q(\ram[6][249] ) );
  DFFX1_HVT \ram_reg[6][248]  ( .D(n1845), .CLK(clk), .Q(\ram[6][248] ) );
  DFFX1_HVT \ram_reg[6][247]  ( .D(n1844), .CLK(clk), .Q(\ram[6][247] ) );
  DFFX1_HVT \ram_reg[6][246]  ( .D(n1843), .CLK(clk), .Q(\ram[6][246] ) );
  DFFX1_HVT \ram_reg[6][245]  ( .D(n1842), .CLK(clk), .Q(\ram[6][245] ) );
  DFFX1_HVT \ram_reg[6][244]  ( .D(n1841), .CLK(clk), .Q(\ram[6][244] ) );
  DFFX1_HVT \ram_reg[6][243]  ( .D(n1840), .CLK(clk), .Q(\ram[6][243] ) );
  DFFX1_HVT \ram_reg[6][242]  ( .D(n1839), .CLK(clk), .Q(\ram[6][242] ) );
  DFFX1_HVT \ram_reg[6][241]  ( .D(n1838), .CLK(clk), .Q(\ram[6][241] ) );
  DFFX1_HVT \ram_reg[6][240]  ( .D(n1837), .CLK(clk), .Q(\ram[6][240] ) );
  DFFX1_HVT \ram_reg[6][239]  ( .D(n1836), .CLK(clk), .Q(\ram[6][239] ) );
  DFFX1_HVT \ram_reg[6][238]  ( .D(n1835), .CLK(clk), .Q(\ram[6][238] ) );
  DFFX1_HVT \ram_reg[6][237]  ( .D(n1834), .CLK(clk), .Q(\ram[6][237] ) );
  DFFX1_HVT \ram_reg[6][236]  ( .D(n1833), .CLK(clk), .Q(\ram[6][236] ) );
  DFFX1_HVT \ram_reg[6][235]  ( .D(n1832), .CLK(clk), .Q(\ram[6][235] ) );
  DFFX1_HVT \ram_reg[6][234]  ( .D(n1831), .CLK(clk), .Q(\ram[6][234] ), .QN(
        n5717) );
  DFFX1_HVT \ram_reg[6][233]  ( .D(n1830), .CLK(clk), .Q(\ram[6][233] ) );
  DFFX1_HVT \ram_reg[6][232]  ( .D(n1829), .CLK(clk), .Q(\ram[6][232] ) );
  DFFX1_HVT \ram_reg[6][231]  ( .D(n1828), .CLK(clk), .Q(\ram[6][231] ) );
  DFFX1_HVT \ram_reg[6][230]  ( .D(n1827), .CLK(clk), .Q(\ram[6][230] ) );
  DFFX1_HVT \ram_reg[6][229]  ( .D(n1826), .CLK(clk), .Q(\ram[6][229] ) );
  DFFX1_HVT \ram_reg[6][228]  ( .D(n1825), .CLK(clk), .Q(\ram[6][228] ) );
  DFFX1_HVT \ram_reg[6][227]  ( .D(n1824), .CLK(clk), .Q(\ram[6][227] ) );
  DFFX1_HVT \ram_reg[6][226]  ( .D(n1823), .CLK(clk), .Q(\ram[6][226] ) );
  DFFX1_HVT \ram_reg[6][225]  ( .D(n1822), .CLK(clk), .Q(\ram[6][225] ) );
  DFFX1_HVT \ram_reg[6][224]  ( .D(n1821), .CLK(clk), .Q(\ram[6][224] ) );
  DFFX1_HVT \ram_reg[6][223]  ( .D(n1820), .CLK(clk), .Q(\ram[6][223] ) );
  DFFX1_HVT \ram_reg[6][222]  ( .D(n1819), .CLK(clk), .Q(\ram[6][222] ) );
  DFFX1_HVT \ram_reg[6][221]  ( .D(n1818), .CLK(clk), .Q(\ram[6][221] ) );
  DFFX1_HVT \ram_reg[6][220]  ( .D(n1817), .CLK(clk), .Q(\ram[6][220] ) );
  DFFX1_HVT \ram_reg[6][219]  ( .D(n1816), .CLK(clk), .Q(\ram[6][219] ) );
  DFFX1_HVT \ram_reg[6][218]  ( .D(n1815), .CLK(clk), .Q(\ram[6][218] ) );
  DFFX1_HVT \ram_reg[6][217]  ( .D(n1814), .CLK(clk), .Q(\ram[6][217] ), .QN(
        n5497) );
  DFFX1_HVT \ram_reg[6][216]  ( .D(n1813), .CLK(clk), .Q(\ram[6][216] ) );
  DFFX1_HVT \ram_reg[6][215]  ( .D(n1812), .CLK(clk), .Q(\ram[6][215] ) );
  DFFX1_HVT \ram_reg[6][214]  ( .D(n1811), .CLK(clk), .Q(\ram[6][214] ) );
  DFFX1_HVT \ram_reg[6][213]  ( .D(n1810), .CLK(clk), .Q(\ram[6][213] ) );
  DFFX1_HVT \ram_reg[6][212]  ( .D(n1809), .CLK(clk), .Q(\ram[6][212] ) );
  DFFX1_HVT \ram_reg[6][211]  ( .D(n1808), .CLK(clk), .Q(\ram[6][211] ) );
  DFFX1_HVT \ram_reg[6][210]  ( .D(n1807), .CLK(clk), .Q(\ram[6][210] ) );
  DFFX1_HVT \ram_reg[6][209]  ( .D(n1806), .CLK(clk), .Q(\ram[6][209] ) );
  DFFX1_HVT \ram_reg[6][208]  ( .D(n1805), .CLK(clk), .Q(\ram[6][208] ) );
  DFFX1_HVT \ram_reg[6][207]  ( .D(n1804), .CLK(clk), .Q(\ram[6][207] ) );
  DFFX1_HVT \ram_reg[6][206]  ( .D(n1803), .CLK(clk), .Q(\ram[6][206] ), .QN(
        n36) );
  DFFX1_HVT \ram_reg[6][205]  ( .D(n1802), .CLK(clk), .Q(\ram[6][205] ) );
  DFFX1_HVT \ram_reg[6][204]  ( .D(n5429), .CLK(clk), .Q(\ram[6][204] ), .QN(
        n6631) );
  DFFX1_HVT \ram_reg[6][203]  ( .D(n1800), .CLK(clk), .Q(\ram[6][203] ) );
  DFFX1_HVT \ram_reg[6][202]  ( .D(n1799), .CLK(clk), .Q(\ram[6][202] ) );
  DFFX1_HVT \ram_reg[6][201]  ( .D(n5023), .CLK(clk), .Q(\ram[6][201] ), .QN(
        n5526) );
  DFFX1_HVT \ram_reg[6][200]  ( .D(n1797), .CLK(clk), .Q(\ram[6][200] ) );
  DFFX1_HVT \ram_reg[6][199]  ( .D(n1796), .CLK(clk), .Q(\ram[6][199] ) );
  DFFX1_HVT \ram_reg[6][198]  ( .D(n1795), .CLK(clk), .Q(\ram[6][198] ) );
  DFFX1_HVT \ram_reg[6][197]  ( .D(n1794), .CLK(clk), .Q(\ram[6][197] ) );
  DFFX1_HVT \ram_reg[6][196]  ( .D(n1793), .CLK(clk), .Q(\ram[6][196] ) );
  DFFX1_HVT \ram_reg[6][195]  ( .D(n1792), .CLK(clk), .Q(\ram[6][195] ) );
  DFFX1_HVT \ram_reg[6][194]  ( .D(n1791), .CLK(clk), .Q(\ram[6][194] ) );
  DFFX1_HVT \ram_reg[6][193]  ( .D(n1790), .CLK(clk), .Q(\ram[6][193] ) );
  DFFX1_HVT \ram_reg[6][192]  ( .D(n1789), .CLK(clk), .Q(\ram[6][192] ) );
  DFFX1_HVT \ram_reg[6][191]  ( .D(n1788), .CLK(clk), .Q(\ram[6][191] ) );
  DFFX1_HVT \ram_reg[6][190]  ( .D(n1787), .CLK(clk), .Q(\ram[6][190] ) );
  DFFX1_HVT \ram_reg[6][189]  ( .D(n1786), .CLK(clk), .Q(\ram[6][189] ) );
  DFFX1_HVT \ram_reg[6][188]  ( .D(n1785), .CLK(clk), .Q(\ram[6][188] ) );
  DFFX1_HVT \ram_reg[6][187]  ( .D(n1784), .CLK(clk), .Q(\ram[6][187] ) );
  DFFX1_HVT \ram_reg[6][186]  ( .D(n1783), .CLK(clk), .Q(\ram[6][186] ) );
  DFFX1_HVT \ram_reg[6][185]  ( .D(n1782), .CLK(clk), .Q(\ram[6][185] ) );
  DFFX1_HVT \ram_reg[6][184]  ( .D(n1781), .CLK(clk), .Q(\ram[6][184] ) );
  DFFX1_HVT \ram_reg[6][183]  ( .D(n1780), .CLK(clk), .Q(\ram[6][183] ) );
  DFFX1_HVT \ram_reg[6][182]  ( .D(n1779), .CLK(clk), .Q(\ram[6][182] ) );
  DFFX1_HVT \ram_reg[6][181]  ( .D(n1778), .CLK(clk), .Q(\ram[6][181] ) );
  DFFX1_HVT \ram_reg[6][180]  ( .D(n1777), .CLK(clk), .Q(\ram[6][180] ) );
  DFFX1_HVT \ram_reg[6][179]  ( .D(n1776), .CLK(clk), .Q(\ram[6][179] ) );
  DFFX1_HVT \ram_reg[6][178]  ( .D(n1775), .CLK(clk), .Q(\ram[6][178] ) );
  DFFX1_HVT \ram_reg[6][177]  ( .D(n1774), .CLK(clk), .Q(\ram[6][177] ) );
  DFFX1_HVT \ram_reg[6][176]  ( .D(n1773), .CLK(clk), .Q(\ram[6][176] ) );
  DFFX1_HVT \ram_reg[6][175]  ( .D(n1772), .CLK(clk), .Q(\ram[6][175] ) );
  DFFX1_HVT \ram_reg[6][174]  ( .D(n1771), .CLK(clk), .Q(\ram[6][174] ) );
  DFFX1_HVT \ram_reg[6][173]  ( .D(n1770), .CLK(clk), .Q(\ram[6][173] ) );
  DFFX1_HVT \ram_reg[6][172]  ( .D(n1769), .CLK(clk), .Q(\ram[6][172] ) );
  DFFX1_HVT \ram_reg[6][171]  ( .D(n1768), .CLK(clk), .Q(\ram[6][171] ) );
  DFFX1_HVT \ram_reg[6][170]  ( .D(n1767), .CLK(clk), .Q(\ram[6][170] ) );
  DFFX1_HVT \ram_reg[6][169]  ( .D(n1766), .CLK(clk), .Q(\ram[6][169] ) );
  DFFX1_HVT \ram_reg[6][168]  ( .D(n1765), .CLK(clk), .Q(\ram[6][168] ) );
  DFFX1_HVT \ram_reg[6][167]  ( .D(n1764), .CLK(clk), .Q(\ram[6][167] ) );
  DFFX1_HVT \ram_reg[6][166]  ( .D(n1763), .CLK(clk), .Q(\ram[6][166] ) );
  DFFX1_HVT \ram_reg[6][165]  ( .D(n1762), .CLK(clk), .Q(\ram[6][165] ) );
  DFFX1_HVT \ram_reg[6][164]  ( .D(n1761), .CLK(clk), .Q(\ram[6][164] ) );
  DFFX1_HVT \ram_reg[6][163]  ( .D(n1760), .CLK(clk), .Q(\ram[6][163] ) );
  DFFX1_HVT \ram_reg[6][162]  ( .D(n1759), .CLK(clk), .Q(\ram[6][162] ) );
  DFFX1_HVT \ram_reg[6][161]  ( .D(n1758), .CLK(clk), .Q(\ram[6][161] ) );
  DFFX1_HVT \ram_reg[6][160]  ( .D(n1757), .CLK(clk), .Q(\ram[6][160] ) );
  DFFX1_HVT \ram_reg[6][159]  ( .D(n1756), .CLK(clk), .Q(\ram[6][159] ) );
  DFFX1_HVT \ram_reg[6][158]  ( .D(n1755), .CLK(clk), .Q(\ram[6][158] ) );
  DFFX1_HVT \ram_reg[6][157]  ( .D(n1754), .CLK(clk), .Q(\ram[6][157] ) );
  DFFX1_HVT \ram_reg[6][156]  ( .D(n1753), .CLK(clk), .Q(\ram[6][156] ) );
  DFFX1_HVT \ram_reg[6][155]  ( .D(n1752), .CLK(clk), .Q(\ram[6][155] ) );
  DFFX1_HVT \ram_reg[6][154]  ( .D(n1751), .CLK(clk), .Q(\ram[6][154] ) );
  DFFX1_HVT \ram_reg[6][153]  ( .D(n1750), .CLK(clk), .Q(\ram[6][153] ) );
  DFFX1_HVT \ram_reg[6][152]  ( .D(n1749), .CLK(clk), .Q(\ram[6][152] ) );
  DFFX1_HVT \ram_reg[6][151]  ( .D(n1748), .CLK(clk), .Q(\ram[6][151] ) );
  DFFX1_HVT \ram_reg[6][150]  ( .D(n1747), .CLK(clk), .Q(\ram[6][150] ) );
  DFFX1_HVT \ram_reg[6][149]  ( .D(n1746), .CLK(clk), .Q(\ram[6][149] ) );
  DFFX1_HVT \ram_reg[6][148]  ( .D(n1745), .CLK(clk), .Q(\ram[6][148] ) );
  DFFX1_HVT \ram_reg[6][147]  ( .D(n1744), .CLK(clk), .Q(\ram[6][147] ) );
  DFFX1_HVT \ram_reg[6][146]  ( .D(n1743), .CLK(clk), .Q(\ram[6][146] ) );
  DFFX1_HVT \ram_reg[6][145]  ( .D(n1742), .CLK(clk), .Q(\ram[6][145] ) );
  DFFX1_HVT \ram_reg[6][144]  ( .D(n1741), .CLK(clk), .Q(\ram[6][144] ) );
  DFFX1_HVT \ram_reg[6][143]  ( .D(n1740), .CLK(clk), .Q(\ram[6][143] ) );
  DFFX1_HVT \ram_reg[6][142]  ( .D(n1739), .CLK(clk), .Q(\ram[6][142] ) );
  DFFX1_HVT \ram_reg[6][141]  ( .D(n1738), .CLK(clk), .Q(\ram[6][141] ) );
  DFFX1_HVT \ram_reg[6][140]  ( .D(n1737), .CLK(clk), .Q(\ram[6][140] ) );
  DFFX1_HVT \ram_reg[6][139]  ( .D(n1736), .CLK(clk), .Q(\ram[6][139] ) );
  DFFX1_HVT \ram_reg[6][138]  ( .D(n1735), .CLK(clk), .Q(\ram[6][138] ) );
  DFFX1_HVT \ram_reg[6][137]  ( .D(n1734), .CLK(clk), .Q(\ram[6][137] ) );
  DFFX1_HVT \ram_reg[6][136]  ( .D(n1733), .CLK(clk), .Q(\ram[6][136] ) );
  DFFX1_HVT \ram_reg[6][135]  ( .D(n1732), .CLK(clk), .Q(\ram[6][135] ) );
  DFFX1_HVT \ram_reg[6][134]  ( .D(n1731), .CLK(clk), .Q(\ram[6][134] ) );
  DFFX1_HVT \ram_reg[6][133]  ( .D(n1730), .CLK(clk), .Q(\ram[6][133] ) );
  DFFX1_HVT \ram_reg[6][132]  ( .D(n1729), .CLK(clk), .Q(\ram[6][132] ) );
  DFFX1_HVT \ram_reg[6][131]  ( .D(n1728), .CLK(clk), .Q(\ram[6][131] ) );
  DFFX1_HVT \ram_reg[6][130]  ( .D(n1727), .CLK(clk), .Q(\ram[6][130] ) );
  DFFX1_HVT \ram_reg[6][129]  ( .D(n1726), .CLK(clk), .Q(\ram[6][129] ) );
  DFFX1_HVT \ram_reg[6][128]  ( .D(n1725), .CLK(clk), .Q(\ram[6][128] ) );
  DFFX1_HVT \ram_reg[6][127]  ( .D(n1724), .CLK(clk), .Q(\ram[6][127] ) );
  DFFX1_HVT \ram_reg[6][126]  ( .D(n1723), .CLK(clk), .Q(\ram[6][126] ) );
  DFFX1_HVT \ram_reg[6][125]  ( .D(n1722), .CLK(clk), .Q(\ram[6][125] ) );
  DFFX1_HVT \ram_reg[6][124]  ( .D(n1721), .CLK(clk), .Q(\ram[6][124] ) );
  DFFX1_HVT \ram_reg[6][123]  ( .D(n1720), .CLK(clk), .Q(\ram[6][123] ) );
  DFFX1_HVT \ram_reg[6][122]  ( .D(n1719), .CLK(clk), .Q(\ram[6][122] ) );
  DFFX1_HVT \ram_reg[6][121]  ( .D(n1718), .CLK(clk), .Q(\ram[6][121] ) );
  DFFX1_HVT \ram_reg[6][120]  ( .D(n1717), .CLK(clk), .Q(\ram[6][120] ) );
  DFFX1_HVT \ram_reg[6][119]  ( .D(n1716), .CLK(clk), .Q(\ram[6][119] ) );
  DFFX1_HVT \ram_reg[6][118]  ( .D(n1715), .CLK(clk), .Q(\ram[6][118] ), .QN(
        n5464) );
  DFFX1_HVT \ram_reg[6][117]  ( .D(n1714), .CLK(clk), .Q(\ram[6][117] ) );
  DFFX1_HVT \ram_reg[6][116]  ( .D(n1713), .CLK(clk), .Q(\ram[6][116] ) );
  DFFX1_HVT \ram_reg[6][115]  ( .D(n1712), .CLK(clk), .Q(\ram[6][115] ) );
  DFFX1_HVT \ram_reg[6][114]  ( .D(n1711), .CLK(clk), .Q(\ram[6][114] ) );
  DFFX1_HVT \ram_reg[6][113]  ( .D(n1710), .CLK(clk), .Q(\ram[6][113] ) );
  DFFX1_HVT \ram_reg[6][112]  ( .D(n1709), .CLK(clk), .Q(\ram[6][112] ) );
  DFFX1_HVT \ram_reg[6][111]  ( .D(n1708), .CLK(clk), .Q(\ram[6][111] ) );
  DFFX1_HVT \ram_reg[6][110]  ( .D(n1707), .CLK(clk), .Q(\ram[6][110] ) );
  DFFX1_HVT \ram_reg[6][109]  ( .D(n1706), .CLK(clk), .Q(\ram[6][109] ) );
  DFFX1_HVT \ram_reg[6][108]  ( .D(n1705), .CLK(clk), .Q(\ram[6][108] ) );
  DFFX1_HVT \ram_reg[6][107]  ( .D(n1704), .CLK(clk), .Q(\ram[6][107] ) );
  DFFX1_HVT \ram_reg[6][106]  ( .D(n1703), .CLK(clk), .Q(\ram[6][106] ) );
  DFFX1_HVT \ram_reg[6][105]  ( .D(n1702), .CLK(clk), .Q(\ram[6][105] ) );
  DFFX1_HVT \ram_reg[6][104]  ( .D(n1701), .CLK(clk), .Q(\ram[6][104] ) );
  DFFX1_HVT \ram_reg[6][103]  ( .D(n1700), .CLK(clk), .Q(\ram[6][103] ) );
  DFFX1_HVT \ram_reg[6][102]  ( .D(n1699), .CLK(clk), .Q(\ram[6][102] ) );
  DFFX1_HVT \ram_reg[6][101]  ( .D(n1698), .CLK(clk), .Q(\ram[6][101] ) );
  DFFX1_HVT \ram_reg[6][100]  ( .D(n1697), .CLK(clk), .Q(\ram[6][100] ) );
  DFFX1_HVT \ram_reg[6][99]  ( .D(n1696), .CLK(clk), .Q(\ram[6][99] ) );
  DFFX1_HVT \ram_reg[6][98]  ( .D(n1695), .CLK(clk), .Q(\ram[6][98] ) );
  DFFX1_HVT \ram_reg[6][97]  ( .D(n1694), .CLK(clk), .Q(\ram[6][97] ) );
  DFFX1_HVT \ram_reg[6][96]  ( .D(n1693), .CLK(clk), .Q(\ram[6][96] ) );
  DFFX1_HVT \ram_reg[6][95]  ( .D(n1692), .CLK(clk), .Q(\ram[6][95] ) );
  DFFX1_HVT \ram_reg[6][94]  ( .D(n1691), .CLK(clk), .Q(\ram[6][94] ) );
  DFFX1_HVT \ram_reg[6][93]  ( .D(n1690), .CLK(clk), .Q(\ram[6][93] ) );
  DFFX1_HVT \ram_reg[6][92]  ( .D(n1689), .CLK(clk), .Q(\ram[6][92] ) );
  DFFX1_HVT \ram_reg[6][91]  ( .D(n1688), .CLK(clk), .Q(\ram[6][91] ) );
  DFFX1_HVT \ram_reg[6][90]  ( .D(n1687), .CLK(clk), .Q(\ram[6][90] ) );
  DFFX1_HVT \ram_reg[6][89]  ( .D(n1686), .CLK(clk), .Q(\ram[6][89] ) );
  DFFX1_HVT \ram_reg[6][88]  ( .D(n1685), .CLK(clk), .Q(\ram[6][88] ) );
  DFFX1_HVT \ram_reg[6][87]  ( .D(n1684), .CLK(clk), .Q(\ram[6][87] ) );
  DFFX1_HVT \ram_reg[6][86]  ( .D(n1683), .CLK(clk), .Q(\ram[6][86] ) );
  DFFX1_HVT \ram_reg[6][85]  ( .D(n1682), .CLK(clk), .Q(\ram[6][85] ) );
  DFFX1_HVT \ram_reg[6][84]  ( .D(n1681), .CLK(clk), .Q(\ram[6][84] ) );
  DFFX1_HVT \ram_reg[6][83]  ( .D(n1680), .CLK(clk), .Q(\ram[6][83] ) );
  DFFX1_HVT \ram_reg[6][82]  ( .D(n1679), .CLK(clk), .Q(\ram[6][82] ) );
  DFFX1_HVT \ram_reg[6][81]  ( .D(n1678), .CLK(clk), .Q(\ram[6][81] ) );
  DFFX1_HVT \ram_reg[6][80]  ( .D(n1677), .CLK(clk), .Q(\ram[6][80] ) );
  DFFX1_HVT \ram_reg[6][79]  ( .D(n1676), .CLK(clk), .Q(\ram[6][79] ) );
  DFFX1_HVT \ram_reg[6][78]  ( .D(n1675), .CLK(clk), .Q(\ram[6][78] ) );
  DFFX1_HVT \ram_reg[6][77]  ( .D(n1674), .CLK(clk), .Q(\ram[6][77] ) );
  DFFX1_HVT \ram_reg[6][76]  ( .D(n1673), .CLK(clk), .Q(\ram[6][76] ) );
  DFFX1_HVT \ram_reg[6][75]  ( .D(n1672), .CLK(clk), .Q(\ram[6][75] ) );
  DFFX1_HVT \ram_reg[6][74]  ( .D(n1671), .CLK(clk), .Q(\ram[6][74] ) );
  DFFX1_HVT \ram_reg[6][73]  ( .D(n1670), .CLK(clk), .Q(\ram[6][73] ) );
  DFFX1_HVT \ram_reg[6][72]  ( .D(n1669), .CLK(clk), .Q(\ram[6][72] ) );
  DFFX1_HVT \ram_reg[6][71]  ( .D(n1668), .CLK(clk), .Q(\ram[6][71] ) );
  DFFX1_HVT \ram_reg[6][70]  ( .D(n1667), .CLK(clk), .Q(\ram[6][70] ) );
  DFFX1_HVT \ram_reg[6][69]  ( .D(n1666), .CLK(clk), .Q(\ram[6][69] ) );
  DFFX1_HVT \ram_reg[6][68]  ( .D(n1665), .CLK(clk), .Q(\ram[6][68] ), .QN(
        n4875) );
  DFFX1_HVT \ram_reg[6][67]  ( .D(n1664), .CLK(clk), .Q(\ram[6][67] ) );
  DFFX1_HVT \ram_reg[6][66]  ( .D(n1663), .CLK(clk), .Q(\ram[6][66] ) );
  DFFX1_HVT \ram_reg[6][65]  ( .D(n1662), .CLK(clk), .Q(\ram[6][65] ) );
  DFFX1_HVT \ram_reg[6][64]  ( .D(n1661), .CLK(clk), .Q(\ram[6][64] ) );
  DFFX1_HVT \ram_reg[6][63]  ( .D(n1660), .CLK(clk), .Q(\ram[6][63] ) );
  DFFX1_HVT \ram_reg[6][62]  ( .D(n1659), .CLK(clk), .Q(\ram[6][62] ) );
  DFFX1_HVT \ram_reg[6][61]  ( .D(n1658), .CLK(clk), .Q(\ram[6][61] ) );
  DFFX1_HVT \ram_reg[6][60]  ( .D(n1657), .CLK(clk), .Q(\ram[6][60] ) );
  DFFX1_HVT \ram_reg[6][59]  ( .D(n1656), .CLK(clk), .Q(\ram[6][59] ) );
  DFFX1_HVT \ram_reg[6][58]  ( .D(n1655), .CLK(clk), .Q(\ram[6][58] ) );
  DFFX1_HVT \ram_reg[6][57]  ( .D(n1654), .CLK(clk), .Q(\ram[6][57] ) );
  DFFX1_HVT \ram_reg[6][56]  ( .D(n1653), .CLK(clk), .Q(\ram[6][56] ) );
  DFFX1_HVT \ram_reg[6][55]  ( .D(n1652), .CLK(clk), .Q(\ram[6][55] ) );
  DFFX1_HVT \ram_reg[6][54]  ( .D(n4754), .CLK(clk), .QN(n5842) );
  DFFX1_HVT \ram_reg[6][53]  ( .D(n1650), .CLK(clk), .Q(\ram[6][53] ), .QN(
        n5844) );
  DFFX1_HVT \ram_reg[6][52]  ( .D(n1649), .CLK(clk), .Q(\ram[6][52] ) );
  DFFX1_HVT \ram_reg[6][51]  ( .D(n1648), .CLK(clk), .Q(\ram[6][51] ), .QN(
        n5847) );
  DFFX1_HVT \ram_reg[6][50]  ( .D(n1647), .CLK(clk), .Q(\ram[6][50] ) );
  DFFX1_HVT \ram_reg[6][49]  ( .D(n1646), .CLK(clk), .Q(\ram[6][49] ), .QN(
        n5850) );
  DFFX1_HVT \ram_reg[6][48]  ( .D(n1645), .CLK(clk), .Q(\ram[6][48] ) );
  DFFX1_HVT \ram_reg[6][47]  ( .D(n1644), .CLK(clk), .Q(\ram[6][47] ) );
  DFFX1_HVT \ram_reg[6][46]  ( .D(n1643), .CLK(clk), .Q(\ram[6][46] ) );
  DFFX1_HVT \ram_reg[6][45]  ( .D(n1642), .CLK(clk), .Q(\ram[6][45] ) );
  DFFX1_HVT \ram_reg[6][44]  ( .D(n1641), .CLK(clk), .Q(\ram[6][44] ) );
  DFFX1_HVT \ram_reg[6][43]  ( .D(n1640), .CLK(clk), .Q(\ram[6][43] ) );
  DFFX1_HVT \ram_reg[6][42]  ( .D(n1639), .CLK(clk), .Q(\ram[6][42] ) );
  DFFX1_HVT \ram_reg[6][41]  ( .D(n1638), .CLK(clk), .Q(\ram[6][41] ) );
  DFFX1_HVT \ram_reg[6][40]  ( .D(n1637), .CLK(clk), .Q(\ram[6][40] ) );
  DFFX1_HVT \ram_reg[6][39]  ( .D(n1636), .CLK(clk), .Q(\ram[6][39] ) );
  DFFX1_HVT \ram_reg[6][38]  ( .D(n1635), .CLK(clk), .Q(\ram[6][38] ) );
  DFFX1_HVT \ram_reg[6][37]  ( .D(n1634), .CLK(clk), .Q(\ram[6][37] ) );
  DFFX1_HVT \ram_reg[6][36]  ( .D(n5025), .CLK(clk), .Q(\ram[6][36] ), .QN(
        n6011) );
  DFFX1_HVT \ram_reg[6][35]  ( .D(n1632), .CLK(clk), .Q(\ram[6][35] ) );
  DFFX1_HVT \ram_reg[6][34]  ( .D(n1631), .CLK(clk), .Q(\ram[6][34] ) );
  DFFX1_HVT \ram_reg[6][33]  ( .D(n1630), .CLK(clk), .Q(\ram[6][33] ) );
  DFFX1_HVT \ram_reg[6][32]  ( .D(n1629), .CLK(clk), .Q(\ram[6][32] ) );
  DFFX1_HVT \ram_reg[6][31]  ( .D(n1628), .CLK(clk), .Q(\ram[6][31] ) );
  DFFX1_HVT \ram_reg[6][30]  ( .D(n1627), .CLK(clk), .Q(\ram[6][30] ), .QN(
        n5206) );
  DFFX1_HVT \ram_reg[6][29]  ( .D(n1626), .CLK(clk), .Q(\ram[6][29] ) );
  DFFX1_HVT \ram_reg[6][28]  ( .D(n1625), .CLK(clk), .Q(\ram[6][28] ) );
  DFFX1_HVT \ram_reg[6][27]  ( .D(n1624), .CLK(clk), .Q(\ram[6][27] ) );
  DFFX1_HVT \ram_reg[6][26]  ( .D(n1623), .CLK(clk), .Q(\ram[6][26] ) );
  DFFX1_HVT \ram_reg[6][25]  ( .D(n1622), .CLK(clk), .Q(\ram[6][25] ) );
  DFFX1_HVT \ram_reg[6][24]  ( .D(n1621), .CLK(clk), .Q(\ram[6][24] ) );
  DFFX1_HVT \ram_reg[6][23]  ( .D(n1620), .CLK(clk), .Q(\ram[6][23] ) );
  DFFX1_HVT \ram_reg[6][22]  ( .D(n1619), .CLK(clk), .Q(\ram[6][22] ) );
  DFFX1_HVT \ram_reg[6][21]  ( .D(n1618), .CLK(clk), .Q(\ram[6][21] ) );
  DFFX1_HVT \ram_reg[6][20]  ( .D(n1617), .CLK(clk), .QN(n6554) );
  DFFX1_HVT \ram_reg[6][19]  ( .D(n1616), .CLK(clk), .Q(\ram[6][19] ) );
  DFFX1_HVT \ram_reg[6][18]  ( .D(n1615), .CLK(clk), .Q(\ram[6][18] ) );
  DFFX1_HVT \ram_reg[6][17]  ( .D(n1614), .CLK(clk), .Q(\ram[6][17] ) );
  DFFX1_HVT \ram_reg[6][16]  ( .D(n1613), .CLK(clk), .Q(\ram[6][16] ), .QN(
        n5561) );
  DFFX1_HVT \ram_reg[6][15]  ( .D(n1612), .CLK(clk), .Q(\ram[6][15] ) );
  DFFX1_HVT \ram_reg[6][14]  ( .D(n1611), .CLK(clk), .Q(\ram[6][14] ) );
  DFFX1_HVT \ram_reg[6][13]  ( .D(n1610), .CLK(clk), .Q(\ram[6][13] ) );
  DFFX1_HVT \ram_reg[6][12]  ( .D(n1609), .CLK(clk), .Q(\ram[6][12] ) );
  DFFX1_HVT \ram_reg[6][11]  ( .D(n1608), .CLK(clk), .Q(\ram[6][11] ) );
  DFFX1_HVT \ram_reg[6][10]  ( .D(n1607), .CLK(clk), .Q(\ram[6][10] ) );
  DFFX1_HVT \ram_reg[6][9]  ( .D(n1606), .CLK(clk), .Q(\ram[6][9] ) );
  DFFX1_HVT \ram_reg[6][8]  ( .D(n1605), .CLK(clk), .Q(\ram[6][8] ) );
  DFFX1_HVT \ram_reg[6][7]  ( .D(n1604), .CLK(clk), .Q(\ram[6][7] ) );
  DFFX1_HVT \ram_reg[6][6]  ( .D(n1603), .CLK(clk), .Q(\ram[6][6] ) );
  DFFX1_HVT \ram_reg[6][5]  ( .D(n1602), .CLK(clk), .Q(\ram[6][5] ), .QN(n5534) );
  DFFX1_HVT \ram_reg[6][4]  ( .D(n1601), .CLK(clk), .Q(\ram[6][4] ) );
  DFFX1_HVT \ram_reg[6][3]  ( .D(n1600), .CLK(clk), .Q(\ram[6][3] ) );
  DFFX1_HVT \ram_reg[6][2]  ( .D(n1599), .CLK(clk), .Q(\ram[6][2] ), .QN(n4892) );
  DFFX1_HVT \ram_reg[6][1]  ( .D(n1598), .CLK(clk), .Q(\ram[6][1] ) );
  DFFX1_HVT \ram_reg[6][0]  ( .D(n5026), .CLK(clk), .Q(\ram[6][0] ), .QN(n5532) );
  DFFX1_HVT \ram_reg[5][255]  ( .D(n1596), .CLK(clk), .Q(\ram[5][255] ) );
  DFFX1_HVT \ram_reg[5][254]  ( .D(n1595), .CLK(clk), .Q(\ram[5][254] ) );
  DFFX1_HVT \ram_reg[5][253]  ( .D(n1594), .CLK(clk), .Q(\ram[5][253] ) );
  DFFX1_HVT \ram_reg[5][252]  ( .D(n1593), .CLK(clk), .Q(\ram[5][252] ) );
  DFFX1_HVT \ram_reg[5][251]  ( .D(n1592), .CLK(clk), .Q(\ram[5][251] ) );
  DFFX1_HVT \ram_reg[5][250]  ( .D(n1591), .CLK(clk), .Q(\ram[5][250] ) );
  DFFX1_HVT \ram_reg[5][249]  ( .D(n1590), .CLK(clk), .Q(\ram[5][249] ) );
  DFFX1_HVT \ram_reg[5][248]  ( .D(n1589), .CLK(clk), .Q(\ram[5][248] ) );
  DFFX1_HVT \ram_reg[5][247]  ( .D(n1588), .CLK(clk), .Q(\ram[5][247] ) );
  DFFX1_HVT \ram_reg[5][246]  ( .D(n1587), .CLK(clk), .Q(\ram[5][246] ) );
  DFFX1_HVT \ram_reg[5][245]  ( .D(n1586), .CLK(clk), .Q(\ram[5][245] ) );
  DFFX1_HVT \ram_reg[5][244]  ( .D(n1585), .CLK(clk), .Q(\ram[5][244] ) );
  DFFX1_HVT \ram_reg[5][243]  ( .D(n1584), .CLK(clk), .Q(\ram[5][243] ) );
  DFFX1_HVT \ram_reg[5][242]  ( .D(n1583), .CLK(clk), .Q(\ram[5][242] ) );
  DFFX1_HVT \ram_reg[5][241]  ( .D(n1582), .CLK(clk), .Q(\ram[5][241] ) );
  DFFX1_HVT \ram_reg[5][240]  ( .D(n1581), .CLK(clk), .Q(\ram[5][240] ) );
  DFFX1_HVT \ram_reg[5][239]  ( .D(n1580), .CLK(clk), .Q(\ram[5][239] ) );
  DFFX1_HVT \ram_reg[5][238]  ( .D(n1579), .CLK(clk), .Q(\ram[5][238] ) );
  DFFX1_HVT \ram_reg[5][237]  ( .D(n1578), .CLK(clk), .Q(\ram[5][237] ), .QN(
        n4329) );
  DFFX1_HVT \ram_reg[5][236]  ( .D(n1577), .CLK(clk), .Q(\ram[5][236] ) );
  DFFX1_HVT \ram_reg[5][235]  ( .D(n1576), .CLK(clk), .Q(\ram[5][235] ) );
  DFFX1_HVT \ram_reg[5][234]  ( .D(n1575), .CLK(clk), .Q(\ram[5][234] ), .QN(
        n5436) );
  DFFX1_HVT \ram_reg[5][233]  ( .D(n1574), .CLK(clk), .Q(\ram[5][233] ) );
  DFFX1_HVT \ram_reg[5][232]  ( .D(n1573), .CLK(clk), .Q(\ram[5][232] ) );
  DFFX1_HVT \ram_reg[5][231]  ( .D(n1572), .CLK(clk), .Q(\ram[5][231] ) );
  DFFX1_HVT \ram_reg[5][230]  ( .D(n1571), .CLK(clk), .Q(\ram[5][230] ), .QN(
        n4641) );
  DFFX1_HVT \ram_reg[5][229]  ( .D(n1570), .CLK(clk), .Q(\ram[5][229] ) );
  DFFX1_HVT \ram_reg[5][228]  ( .D(n1569), .CLK(clk), .Q(\ram[5][228] ) );
  DFFX1_HVT \ram_reg[5][227]  ( .D(n1568), .CLK(clk), .Q(\ram[5][227] ) );
  DFFX1_HVT \ram_reg[5][226]  ( .D(n1567), .CLK(clk), .Q(\ram[5][226] ) );
  DFFX1_HVT \ram_reg[5][225]  ( .D(n1566), .CLK(clk), .Q(\ram[5][225] ) );
  DFFX1_HVT \ram_reg[5][224]  ( .D(n1565), .CLK(clk), .Q(\ram[5][224] ) );
  DFFX1_HVT \ram_reg[5][223]  ( .D(n1564), .CLK(clk), .Q(\ram[5][223] ) );
  DFFX1_HVT \ram_reg[5][222]  ( .D(n1563), .CLK(clk), .Q(\ram[5][222] ) );
  DFFX1_HVT \ram_reg[5][221]  ( .D(n1562), .CLK(clk), .Q(\ram[5][221] ), .QN(
        n4587) );
  DFFX1_HVT \ram_reg[5][220]  ( .D(n1561), .CLK(clk), .Q(\ram[5][220] ), .QN(
        n4624) );
  DFFX1_HVT \ram_reg[5][219]  ( .D(n1560), .CLK(clk), .Q(\ram[5][219] ) );
  DFFX1_HVT \ram_reg[5][218]  ( .D(n1559), .CLK(clk), .Q(\ram[5][218] ) );
  DFFX1_HVT \ram_reg[5][217]  ( .D(n1558), .CLK(clk), .Q(\ram[5][217] ) );
  DFFX1_HVT \ram_reg[5][216]  ( .D(n1557), .CLK(clk), .Q(\ram[5][216] ) );
  DFFX1_HVT \ram_reg[5][215]  ( .D(n1556), .CLK(clk), .Q(\ram[5][215] ) );
  DFFX1_HVT \ram_reg[5][214]  ( .D(n1555), .CLK(clk), .Q(\ram[5][214] ) );
  DFFX1_HVT \ram_reg[5][213]  ( .D(n1554), .CLK(clk), .Q(\ram[5][213] ) );
  DFFX1_HVT \ram_reg[5][212]  ( .D(n1553), .CLK(clk), .Q(\ram[5][212] ), .QN(
        n4739) );
  DFFX1_HVT \ram_reg[5][211]  ( .D(n1552), .CLK(clk), .Q(\ram[5][211] ) );
  DFFX1_HVT \ram_reg[5][210]  ( .D(n1551), .CLK(clk), .Q(\ram[5][210] ) );
  DFFX1_HVT \ram_reg[5][209]  ( .D(n1550), .CLK(clk), .Q(\ram[5][209] ) );
  DFFX1_HVT \ram_reg[5][208]  ( .D(n1549), .CLK(clk), .Q(\ram[5][208] ) );
  DFFX1_HVT \ram_reg[5][207]  ( .D(n1548), .CLK(clk), .Q(\ram[5][207] ) );
  DFFX1_HVT \ram_reg[5][206]  ( .D(n1547), .CLK(clk), .Q(\ram[5][206] ), .QN(
        n42) );
  DFFX1_HVT \ram_reg[5][205]  ( .D(n1546), .CLK(clk), .Q(\ram[5][205] ) );
  DFFX1_HVT \ram_reg[5][204]  ( .D(n1545), .CLK(clk), .Q(\ram[5][204] ) );
  DFFX1_HVT \ram_reg[5][203]  ( .D(n1544), .CLK(clk), .Q(\ram[5][203] ) );
  DFFX1_HVT \ram_reg[5][202]  ( .D(n1543), .CLK(clk), .Q(\ram[5][202] ) );
  DFFX1_HVT \ram_reg[5][201]  ( .D(n1542), .CLK(clk), .Q(\ram[5][201] ) );
  DFFX1_HVT \ram_reg[5][200]  ( .D(n1541), .CLK(clk), .Q(\ram[5][200] ) );
  DFFX1_HVT \ram_reg[5][199]  ( .D(n1540), .CLK(clk), .Q(\ram[5][199] ) );
  DFFX1_HVT \ram_reg[5][198]  ( .D(n1539), .CLK(clk), .Q(\ram[5][198] ) );
  DFFX1_HVT \ram_reg[5][197]  ( .D(n1538), .CLK(clk), .Q(\ram[5][197] ) );
  DFFX1_HVT \ram_reg[5][196]  ( .D(n1537), .CLK(clk), .Q(\ram[5][196] ) );
  DFFX1_HVT \ram_reg[5][195]  ( .D(n1536), .CLK(clk), .Q(\ram[5][195] ) );
  DFFX1_HVT \ram_reg[5][194]  ( .D(n1535), .CLK(clk), .Q(\ram[5][194] ) );
  DFFX1_HVT \ram_reg[5][193]  ( .D(n1534), .CLK(clk), .Q(\ram[5][193] ) );
  DFFX1_HVT \ram_reg[5][192]  ( .D(n1533), .CLK(clk), .Q(\ram[5][192] ) );
  DFFX1_HVT \ram_reg[5][191]  ( .D(n1532), .CLK(clk), .Q(\ram[5][191] ) );
  DFFX1_HVT \ram_reg[5][190]  ( .D(n1531), .CLK(clk), .Q(\ram[5][190] ) );
  DFFX1_HVT \ram_reg[5][189]  ( .D(n1530), .CLK(clk), .Q(\ram[5][189] ) );
  DFFX1_HVT \ram_reg[5][188]  ( .D(n1529), .CLK(clk), .Q(\ram[5][188] ) );
  DFFX1_HVT \ram_reg[5][187]  ( .D(n1528), .CLK(clk), .Q(\ram[5][187] ) );
  DFFX1_HVT \ram_reg[5][186]  ( .D(n1527), .CLK(clk), .Q(\ram[5][186] ) );
  DFFX1_HVT \ram_reg[5][185]  ( .D(n1526), .CLK(clk), .Q(\ram[5][185] ) );
  DFFX1_HVT \ram_reg[5][184]  ( .D(n1525), .CLK(clk), .Q(\ram[5][184] ) );
  DFFX1_HVT \ram_reg[5][183]  ( .D(n1524), .CLK(clk), .Q(\ram[5][183] ) );
  DFFX1_HVT \ram_reg[5][182]  ( .D(n1523), .CLK(clk), .Q(\ram[5][182] ) );
  DFFX1_HVT \ram_reg[5][181]  ( .D(n1522), .CLK(clk), .Q(\ram[5][181] ) );
  DFFX1_HVT \ram_reg[5][180]  ( .D(n1521), .CLK(clk), .Q(\ram[5][180] ) );
  DFFX1_HVT \ram_reg[5][179]  ( .D(n1520), .CLK(clk), .Q(\ram[5][179] ) );
  DFFX1_HVT \ram_reg[5][178]  ( .D(n1519), .CLK(clk), .Q(\ram[5][178] ) );
  DFFX1_HVT \ram_reg[5][177]  ( .D(n1518), .CLK(clk), .Q(\ram[5][177] ) );
  DFFX1_HVT \ram_reg[5][176]  ( .D(n1517), .CLK(clk), .Q(\ram[5][176] ) );
  DFFX1_HVT \ram_reg[5][175]  ( .D(n1516), .CLK(clk), .Q(\ram[5][175] ) );
  DFFX1_HVT \ram_reg[5][174]  ( .D(n1515), .CLK(clk), .Q(\ram[5][174] ) );
  DFFX1_HVT \ram_reg[5][173]  ( .D(n1514), .CLK(clk), .Q(\ram[5][173] ) );
  DFFX1_HVT \ram_reg[5][172]  ( .D(n1513), .CLK(clk), .Q(\ram[5][172] ) );
  DFFX1_HVT \ram_reg[5][171]  ( .D(n1512), .CLK(clk), .Q(\ram[5][171] ) );
  DFFX1_HVT \ram_reg[5][170]  ( .D(n1511), .CLK(clk), .Q(\ram[5][170] ), .QN(
        n4267) );
  DFFX1_HVT \ram_reg[5][169]  ( .D(n1510), .CLK(clk), .Q(\ram[5][169] ) );
  DFFX1_HVT \ram_reg[5][168]  ( .D(n1509), .CLK(clk), .Q(\ram[5][168] ) );
  DFFX1_HVT \ram_reg[5][167]  ( .D(n1508), .CLK(clk), .Q(\ram[5][167] ) );
  DFFX1_HVT \ram_reg[5][166]  ( .D(n1507), .CLK(clk), .Q(\ram[5][166] ) );
  DFFX1_HVT \ram_reg[5][165]  ( .D(n1506), .CLK(clk), .Q(\ram[5][165] ) );
  DFFX1_HVT \ram_reg[5][164]  ( .D(n1505), .CLK(clk), .Q(\ram[5][164] ) );
  DFFX1_HVT \ram_reg[5][163]  ( .D(n1504), .CLK(clk), .Q(\ram[5][163] ) );
  DFFX1_HVT \ram_reg[5][162]  ( .D(n1503), .CLK(clk), .Q(\ram[5][162] ) );
  DFFX1_HVT \ram_reg[5][161]  ( .D(n1502), .CLK(clk), .Q(\ram[5][161] ) );
  DFFX1_HVT \ram_reg[5][160]  ( .D(n1501), .CLK(clk), .Q(\ram[5][160] ) );
  DFFX1_HVT \ram_reg[5][159]  ( .D(n1500), .CLK(clk), .Q(\ram[5][159] ) );
  DFFX1_HVT \ram_reg[5][158]  ( .D(n1499), .CLK(clk), .Q(\ram[5][158] ) );
  DFFX1_HVT \ram_reg[5][157]  ( .D(n1498), .CLK(clk), .Q(\ram[5][157] ) );
  DFFX1_HVT \ram_reg[5][156]  ( .D(n1497), .CLK(clk), .Q(\ram[5][156] ) );
  DFFX1_HVT \ram_reg[5][155]  ( .D(n1496), .CLK(clk), .Q(\ram[5][155] ) );
  DFFX1_HVT \ram_reg[5][154]  ( .D(n1495), .CLK(clk), .Q(\ram[5][154] ) );
  DFFX1_HVT \ram_reg[5][153]  ( .D(n1494), .CLK(clk), .Q(\ram[5][153] ) );
  DFFX1_HVT \ram_reg[5][152]  ( .D(n1493), .CLK(clk), .Q(\ram[5][152] ) );
  DFFX1_HVT \ram_reg[5][151]  ( .D(n1492), .CLK(clk), .Q(\ram[5][151] ) );
  DFFX1_HVT \ram_reg[5][150]  ( .D(n1491), .CLK(clk), .Q(\ram[5][150] ) );
  DFFX1_HVT \ram_reg[5][149]  ( .D(n1490), .CLK(clk), .Q(\ram[5][149] ) );
  DFFX1_HVT \ram_reg[5][148]  ( .D(n1489), .CLK(clk), .Q(\ram[5][148] ) );
  DFFX1_HVT \ram_reg[5][147]  ( .D(n1488), .CLK(clk), .Q(\ram[5][147] ) );
  DFFX1_HVT \ram_reg[5][146]  ( .D(n1487), .CLK(clk), .Q(\ram[5][146] ) );
  DFFX1_HVT \ram_reg[5][145]  ( .D(n1486), .CLK(clk), .Q(\ram[5][145] ) );
  DFFX1_HVT \ram_reg[5][144]  ( .D(n1485), .CLK(clk), .Q(\ram[5][144] ) );
  DFFX1_HVT \ram_reg[5][143]  ( .D(n1484), .CLK(clk), .Q(\ram[5][143] ) );
  DFFX1_HVT \ram_reg[5][142]  ( .D(n1483), .CLK(clk), .Q(\ram[5][142] ) );
  DFFX1_HVT \ram_reg[5][141]  ( .D(n1482), .CLK(clk), .Q(\ram[5][141] ) );
  DFFX1_HVT \ram_reg[5][140]  ( .D(n1481), .CLK(clk), .Q(\ram[5][140] ) );
  DFFX1_HVT \ram_reg[5][139]  ( .D(n1480), .CLK(clk), .Q(\ram[5][139] ) );
  DFFX1_HVT \ram_reg[5][138]  ( .D(n1479), .CLK(clk), .Q(\ram[5][138] ) );
  DFFX1_HVT \ram_reg[5][137]  ( .D(n1478), .CLK(clk), .Q(\ram[5][137] ) );
  DFFX1_HVT \ram_reg[5][136]  ( .D(n1477), .CLK(clk), .Q(\ram[5][136] ) );
  DFFX1_HVT \ram_reg[5][135]  ( .D(n1476), .CLK(clk), .Q(\ram[5][135] ) );
  DFFX1_HVT \ram_reg[5][134]  ( .D(n1475), .CLK(clk), .Q(\ram[5][134] ) );
  DFFX1_HVT \ram_reg[5][133]  ( .D(n1474), .CLK(clk), .Q(\ram[5][133] ) );
  DFFX1_HVT \ram_reg[5][132]  ( .D(n1473), .CLK(clk), .Q(\ram[5][132] ) );
  DFFX1_HVT \ram_reg[5][131]  ( .D(n1472), .CLK(clk), .Q(\ram[5][131] ) );
  DFFX1_HVT \ram_reg[5][130]  ( .D(n1471), .CLK(clk), .Q(\ram[5][130] ) );
  DFFX1_HVT \ram_reg[5][129]  ( .D(n1470), .CLK(clk), .Q(\ram[5][129] ) );
  DFFX1_HVT \ram_reg[5][128]  ( .D(n1469), .CLK(clk), .Q(\ram[5][128] ) );
  DFFX1_HVT \ram_reg[5][127]  ( .D(n1468), .CLK(clk), .Q(\ram[5][127] ) );
  DFFX1_HVT \ram_reg[5][126]  ( .D(n1467), .CLK(clk), .Q(\ram[5][126] ) );
  DFFX1_HVT \ram_reg[5][125]  ( .D(n1466), .CLK(clk), .Q(\ram[5][125] ) );
  DFFX1_HVT \ram_reg[5][124]  ( .D(n1465), .CLK(clk), .Q(\ram[5][124] ) );
  DFFX1_HVT \ram_reg[5][123]  ( .D(n1464), .CLK(clk), .Q(\ram[5][123] ) );
  DFFX1_HVT \ram_reg[5][122]  ( .D(n5435), .CLK(clk), .Q(\ram[5][122] ), .QN(
        n5952) );
  DFFX1_HVT \ram_reg[5][121]  ( .D(n1462), .CLK(clk), .Q(\ram[5][121] ) );
  DFFX1_HVT \ram_reg[5][120]  ( .D(n5430), .CLK(clk), .Q(\ram[5][120] ), .QN(
        n5963) );
  DFFX1_HVT \ram_reg[5][119]  ( .D(n1460), .CLK(clk), .Q(\ram[5][119] ) );
  DFFX1_HVT \ram_reg[5][118]  ( .D(n1459), .CLK(clk), .Q(\ram[5][118] ) );
  DFFX1_HVT \ram_reg[5][117]  ( .D(n1458), .CLK(clk), .Q(\ram[5][117] ) );
  DFFX1_HVT \ram_reg[5][116]  ( .D(n1457), .CLK(clk), .Q(\ram[5][116] ) );
  DFFX1_HVT \ram_reg[5][115]  ( .D(n1456), .CLK(clk), .Q(\ram[5][115] ) );
  DFFX1_HVT \ram_reg[5][114]  ( .D(n1455), .CLK(clk), .Q(\ram[5][114] ) );
  DFFX1_HVT \ram_reg[5][113]  ( .D(n1454), .CLK(clk), .Q(\ram[5][113] ) );
  DFFX1_HVT \ram_reg[5][112]  ( .D(n1453), .CLK(clk), .Q(\ram[5][112] ) );
  DFFX1_HVT \ram_reg[5][111]  ( .D(n1452), .CLK(clk), .Q(\ram[5][111] ) );
  DFFX1_HVT \ram_reg[5][110]  ( .D(n1451), .CLK(clk), .Q(\ram[5][110] ) );
  DFFX1_HVT \ram_reg[5][109]  ( .D(n1450), .CLK(clk), .Q(\ram[5][109] ), .QN(
        n4567) );
  DFFX1_HVT \ram_reg[5][108]  ( .D(n1449), .CLK(clk), .Q(\ram[5][108] ) );
  DFFX1_HVT \ram_reg[5][107]  ( .D(n1448), .CLK(clk), .Q(\ram[5][107] ) );
  DFFX1_HVT \ram_reg[5][106]  ( .D(n1447), .CLK(clk), .Q(\ram[5][106] ) );
  DFFX1_HVT \ram_reg[5][105]  ( .D(n1446), .CLK(clk), .Q(\ram[5][105] ) );
  DFFX1_HVT \ram_reg[5][104]  ( .D(n1445), .CLK(clk), .Q(\ram[5][104] ) );
  DFFX1_HVT \ram_reg[5][103]  ( .D(n1444), .CLK(clk), .Q(\ram[5][103] ) );
  DFFX1_HVT \ram_reg[5][102]  ( .D(n1443), .CLK(clk), .Q(\ram[5][102] ) );
  DFFX1_HVT \ram_reg[5][101]  ( .D(n1442), .CLK(clk), .Q(\ram[5][101] ) );
  DFFX1_HVT \ram_reg[5][100]  ( .D(n1441), .CLK(clk), .Q(\ram[5][100] ) );
  DFFX1_HVT \ram_reg[5][99]  ( .D(n1440), .CLK(clk), .Q(\ram[5][99] ) );
  DFFX1_HVT \ram_reg[5][98]  ( .D(n1439), .CLK(clk), .Q(\ram[5][98] ) );
  DFFX1_HVT \ram_reg[5][97]  ( .D(n1438), .CLK(clk), .Q(\ram[5][97] ), .QN(
        n4241) );
  DFFX1_HVT \ram_reg[5][96]  ( .D(n1437), .CLK(clk), .Q(\ram[5][96] ) );
  DFFX1_HVT \ram_reg[5][95]  ( .D(n1436), .CLK(clk), .Q(\ram[5][95] ) );
  DFFX1_HVT \ram_reg[5][94]  ( .D(n1435), .CLK(clk), .Q(\ram[5][94] ) );
  DFFX1_HVT \ram_reg[5][93]  ( .D(n1434), .CLK(clk), .Q(\ram[5][93] ) );
  DFFX1_HVT \ram_reg[5][92]  ( .D(n1433), .CLK(clk), .Q(\ram[5][92] ) );
  DFFX1_HVT \ram_reg[5][91]  ( .D(n1432), .CLK(clk), .Q(\ram[5][91] ), .QN(
        n4201) );
  DFFX1_HVT \ram_reg[5][90]  ( .D(n1431), .CLK(clk), .Q(\ram[5][90] ) );
  DFFX1_HVT \ram_reg[5][89]  ( .D(n1430), .CLK(clk), .Q(\ram[5][89] ) );
  DFFX1_HVT \ram_reg[5][88]  ( .D(n1429), .CLK(clk), .Q(\ram[5][88] ) );
  DFFX1_HVT \ram_reg[5][87]  ( .D(n1428), .CLK(clk), .Q(\ram[5][87] ) );
  DFFX1_HVT \ram_reg[5][86]  ( .D(n1427), .CLK(clk), .Q(\ram[5][86] ) );
  DFFX1_HVT \ram_reg[5][85]  ( .D(n1426), .CLK(clk), .Q(\ram[5][85] ) );
  DFFX1_HVT \ram_reg[5][84]  ( .D(n1425), .CLK(clk), .Q(\ram[5][84] ) );
  DFFX1_HVT \ram_reg[5][83]  ( .D(n1424), .CLK(clk), .Q(\ram[5][83] ) );
  DFFX1_HVT \ram_reg[5][82]  ( .D(n1423), .CLK(clk), .Q(\ram[5][82] ) );
  DFFX1_HVT \ram_reg[5][81]  ( .D(n1422), .CLK(clk), .Q(\ram[5][81] ) );
  DFFX1_HVT \ram_reg[5][80]  ( .D(n1421), .CLK(clk), .Q(\ram[5][80] ) );
  DFFX1_HVT \ram_reg[5][79]  ( .D(n1420), .CLK(clk), .Q(\ram[5][79] ) );
  DFFX1_HVT \ram_reg[5][78]  ( .D(n1419), .CLK(clk), .Q(\ram[5][78] ) );
  DFFX1_HVT \ram_reg[5][77]  ( .D(n1418), .CLK(clk), .Q(\ram[5][77] ) );
  DFFX1_HVT \ram_reg[5][76]  ( .D(n1417), .CLK(clk), .Q(\ram[5][76] ) );
  DFFX1_HVT \ram_reg[5][75]  ( .D(n1416), .CLK(clk), .Q(\ram[5][75] ) );
  DFFX1_HVT \ram_reg[5][74]  ( .D(n1415), .CLK(clk), .Q(\ram[5][74] ) );
  DFFX1_HVT \ram_reg[5][73]  ( .D(n1414), .CLK(clk), .Q(\ram[5][73] ) );
  DFFX1_HVT \ram_reg[5][72]  ( .D(n1413), .CLK(clk), .Q(\ram[5][72] ) );
  DFFX1_HVT \ram_reg[5][71]  ( .D(n1412), .CLK(clk), .Q(\ram[5][71] ) );
  DFFX1_HVT \ram_reg[5][70]  ( .D(n1411), .CLK(clk), .Q(\ram[5][70] ) );
  DFFX1_HVT \ram_reg[5][69]  ( .D(n1410), .CLK(clk), .Q(\ram[5][69] ) );
  DFFX1_HVT \ram_reg[5][68]  ( .D(n1409), .CLK(clk), .Q(\ram[5][68] ), .QN(
        n4204) );
  DFFX1_HVT \ram_reg[5][67]  ( .D(n1408), .CLK(clk), .Q(\ram[5][67] ) );
  DFFX1_HVT \ram_reg[5][66]  ( .D(n1407), .CLK(clk), .Q(\ram[5][66] ) );
  DFFX1_HVT \ram_reg[5][65]  ( .D(n1406), .CLK(clk), .Q(\ram[5][65] ), .QN(
        n4717) );
  DFFX1_HVT \ram_reg[5][64]  ( .D(n1405), .CLK(clk), .Q(\ram[5][64] ) );
  DFFX1_HVT \ram_reg[5][63]  ( .D(n1404), .CLK(clk), .Q(\ram[5][63] ) );
  DFFX1_HVT \ram_reg[5][62]  ( .D(n1403), .CLK(clk), .Q(\ram[5][62] ), .QN(
        n4944) );
  DFFX1_HVT \ram_reg[5][61]  ( .D(n1402), .CLK(clk), .Q(\ram[5][61] ) );
  DFFX1_HVT \ram_reg[5][60]  ( .D(n1401), .CLK(clk), .Q(\ram[5][60] ) );
  DFFX1_HVT \ram_reg[5][59]  ( .D(n1400), .CLK(clk), .Q(\ram[5][59] ) );
  DFFX1_HVT \ram_reg[5][58]  ( .D(n1399), .CLK(clk), .Q(\ram[5][58] ) );
  DFFX1_HVT \ram_reg[5][57]  ( .D(n1398), .CLK(clk), .Q(\ram[5][57] ) );
  DFFX1_HVT \ram_reg[5][56]  ( .D(n1397), .CLK(clk), .Q(\ram[5][56] ) );
  DFFX1_HVT \ram_reg[5][55]  ( .D(n1396), .CLK(clk), .Q(\ram[5][55] ) );
  DFFX1_HVT \ram_reg[5][54]  ( .D(n1395), .CLK(clk), .Q(\ram[5][54] ), .QN(
        n4805) );
  DFFX1_HVT \ram_reg[5][53]  ( .D(n1394), .CLK(clk), .Q(\ram[5][53] ) );
  DFFX1_HVT \ram_reg[5][52]  ( .D(n1393), .CLK(clk), .Q(\ram[5][52] ) );
  DFFX1_HVT \ram_reg[5][51]  ( .D(n1392), .CLK(clk), .Q(\ram[5][51] ), .QN(
        n4842) );
  DFFX1_HVT \ram_reg[5][50]  ( .D(n5428), .CLK(clk), .Q(\ram[5][50] ), .QN(
        n5876) );
  DFFX1_HVT \ram_reg[5][49]  ( .D(n1390), .CLK(clk), .Q(\ram[5][49] ), .QN(
        n5786) );
  DFFX1_HVT \ram_reg[5][48]  ( .D(n5427), .CLK(clk), .Q(\ram[5][48] ), .QN(
        n7270) );
  DFFX1_HVT \ram_reg[5][47]  ( .D(n1388), .CLK(clk), .Q(\ram[5][47] ), .QN(
        n4730) );
  DFFX1_HVT \ram_reg[5][46]  ( .D(n1387), .CLK(clk), .Q(\ram[5][46] ) );
  DFFX1_HVT \ram_reg[5][45]  ( .D(n1386), .CLK(clk), .Q(\ram[5][45] ) );
  DFFX1_HVT \ram_reg[5][44]  ( .D(n1385), .CLK(clk), .Q(\ram[5][44] ) );
  DFFX1_HVT \ram_reg[5][43]  ( .D(n1384), .CLK(clk), .Q(\ram[5][43] ) );
  DFFX1_HVT \ram_reg[5][42]  ( .D(n1383), .CLK(clk), .Q(\ram[5][42] ) );
  DFFX1_HVT \ram_reg[5][41]  ( .D(n1382), .CLK(clk), .Q(\ram[5][41] ) );
  DFFX1_HVT \ram_reg[5][40]  ( .D(n1381), .CLK(clk), .Q(\ram[5][40] ) );
  DFFX1_HVT \ram_reg[5][39]  ( .D(n1380), .CLK(clk), .Q(\ram[5][39] ) );
  DFFX1_HVT \ram_reg[5][38]  ( .D(n1379), .CLK(clk), .Q(\ram[5][38] ), .QN(
        n4740) );
  DFFX1_HVT \ram_reg[5][37]  ( .D(n1378), .CLK(clk), .Q(\ram[5][37] ) );
  DFFX1_HVT \ram_reg[5][36]  ( .D(n1377), .CLK(clk), .Q(\ram[5][36] ), .QN(
        n4895) );
  DFFX1_HVT \ram_reg[5][35]  ( .D(n1376), .CLK(clk), .Q(\ram[5][35] ) );
  DFFX1_HVT \ram_reg[5][34]  ( .D(n1375), .CLK(clk), .Q(\ram[5][34] ), .QN(
        n4843) );
  DFFX1_HVT \ram_reg[5][33]  ( .D(n1374), .CLK(clk), .Q(\ram[5][33] ) );
  DFFX1_HVT \ram_reg[5][32]  ( .D(n1373), .CLK(clk), .Q(\ram[5][32] ) );
  DFFX1_HVT \ram_reg[5][31]  ( .D(n1372), .CLK(clk), .Q(\ram[5][31] ) );
  DFFX1_HVT \ram_reg[5][30]  ( .D(n1371), .CLK(clk), .Q(\ram[5][30] ), .QN(
        n4963) );
  DFFX1_HVT \ram_reg[5][29]  ( .D(n1370), .CLK(clk), .Q(\ram[5][29] ), .QN(
        n4515) );
  DFFX1_HVT \ram_reg[5][28]  ( .D(n1369), .CLK(clk), .Q(\ram[5][28] ), .QN(
        n4946) );
  DFFX1_HVT \ram_reg[5][27]  ( .D(n1368), .CLK(clk), .Q(\ram[5][27] ) );
  DFFX1_HVT \ram_reg[5][26]  ( .D(n1367), .CLK(clk), .Q(\ram[5][26] ) );
  DFFX1_HVT \ram_reg[5][25]  ( .D(n1366), .CLK(clk), .Q(\ram[5][25] ) );
  DFFX1_HVT \ram_reg[5][24]  ( .D(n1365), .CLK(clk), .Q(\ram[5][24] ) );
  DFFX1_HVT \ram_reg[5][23]  ( .D(n1364), .CLK(clk), .Q(\ram[5][23] ) );
  DFFX1_HVT \ram_reg[5][22]  ( .D(n1363), .CLK(clk), .Q(\ram[5][22] ) );
  DFFX1_HVT \ram_reg[5][21]  ( .D(n1362), .CLK(clk), .Q(\ram[5][21] ) );
  DFFX1_HVT \ram_reg[5][20]  ( .D(n5431), .CLK(clk), .QN(n6553) );
  DFFX1_HVT \ram_reg[5][19]  ( .D(n1360), .CLK(clk), .Q(\ram[5][19] ) );
  DFFX1_HVT \ram_reg[5][18]  ( .D(n5434), .CLK(clk), .Q(\ram[5][18] ), .QN(
        n5781) );
  DFFX1_HVT \ram_reg[5][17]  ( .D(n1358), .CLK(clk), .Q(\ram[5][17] ), .QN(
        n4733) );
  DFFX1_HVT \ram_reg[5][16]  ( .D(n5433), .CLK(clk), .Q(\ram[5][16] ), .QN(
        n5783) );
  DFFX1_HVT \ram_reg[5][15]  ( .D(n1356), .CLK(clk), .Q(\ram[5][15] ), .QN(
        n4681) );
  DFFX1_HVT \ram_reg[5][14]  ( .D(n1355), .CLK(clk), .Q(\ram[5][14] ), .QN(
        n4840) );
  DFFX1_HVT \ram_reg[5][13]  ( .D(n1354), .CLK(clk), .Q(\ram[5][13] ), .QN(
        n4767) );
  DFFX1_HVT \ram_reg[5][12]  ( .D(n1353), .CLK(clk), .Q(\ram[5][12] ), .QN(
        n4287) );
  DFFX1_HVT \ram_reg[5][11]  ( .D(n1352), .CLK(clk), .Q(\ram[5][11] ) );
  DFFX1_HVT \ram_reg[5][10]  ( .D(n1351), .CLK(clk), .Q(\ram[5][10] ), .QN(
        n4694) );
  DFFX1_HVT \ram_reg[5][9]  ( .D(n1350), .CLK(clk), .Q(\ram[5][9] ) );
  DFFX1_HVT \ram_reg[5][8]  ( .D(n1349), .CLK(clk), .Q(\ram[5][8] ), .QN(n4712) );
  DFFX1_HVT \ram_reg[5][7]  ( .D(n1348), .CLK(clk), .Q(\ram[5][7] ) );
  DFFX1_HVT \ram_reg[5][6]  ( .D(n1347), .CLK(clk), .Q(\ram[5][6] ), .QN(n4951) );
  DFFX1_HVT \ram_reg[5][5]  ( .D(n1346), .CLK(clk), .Q(\ram[5][5] ) );
  DFFX1_HVT \ram_reg[5][4]  ( .D(n1345), .CLK(clk), .Q(\ram[5][4] ) );
  DFFX1_HVT \ram_reg[5][3]  ( .D(n5432), .CLK(clk), .Q(\ram[5][3] ), .QN(n5872) );
  DFFX1_HVT \ram_reg[5][2]  ( .D(n1343), .CLK(clk), .Q(\ram[5][2] ), .QN(n4713) );
  DFFX1_HVT \ram_reg[5][1]  ( .D(n1342), .CLK(clk), .Q(\ram[5][1] ) );
  DFFX1_HVT \ram_reg[5][0]  ( .D(n1341), .CLK(clk), .Q(\ram[5][0] ) );
  DFFX1_HVT \ram_reg[4][255]  ( .D(n1340), .CLK(clk), .Q(\ram[4][255] ) );
  DFFX1_HVT \ram_reg[4][254]  ( .D(n1339), .CLK(clk), .Q(\ram[4][254] ) );
  DFFX1_HVT \ram_reg[4][253]  ( .D(n1338), .CLK(clk), .Q(\ram[4][253] ) );
  DFFX1_HVT \ram_reg[4][252]  ( .D(n1337), .CLK(clk), .Q(\ram[4][252] ) );
  DFFX1_HVT \ram_reg[4][251]  ( .D(n1336), .CLK(clk), .Q(\ram[4][251] ) );
  DFFX1_HVT \ram_reg[4][250]  ( .D(n1335), .CLK(clk), .Q(\ram[4][250] ) );
  DFFX1_HVT \ram_reg[4][249]  ( .D(n1334), .CLK(clk), .Q(\ram[4][249] ) );
  DFFX1_HVT \ram_reg[4][248]  ( .D(n1333), .CLK(clk), .Q(\ram[4][248] ) );
  DFFX1_HVT \ram_reg[4][247]  ( .D(n1332), .CLK(clk), .Q(\ram[4][247] ) );
  DFFX1_HVT \ram_reg[4][246]  ( .D(n1331), .CLK(clk), .Q(\ram[4][246] ) );
  DFFX1_HVT \ram_reg[4][245]  ( .D(n1330), .CLK(clk), .Q(\ram[4][245] ) );
  DFFX1_HVT \ram_reg[4][244]  ( .D(n1329), .CLK(clk), .Q(\ram[4][244] ) );
  DFFX1_HVT \ram_reg[4][243]  ( .D(n1328), .CLK(clk), .Q(\ram[4][243] ) );
  DFFX1_HVT \ram_reg[4][242]  ( .D(n1327), .CLK(clk), .Q(\ram[4][242] ) );
  DFFX1_HVT \ram_reg[4][241]  ( .D(n1326), .CLK(clk), .Q(\ram[4][241] ) );
  DFFX1_HVT \ram_reg[4][240]  ( .D(n1325), .CLK(clk), .Q(\ram[4][240] ) );
  DFFX1_HVT \ram_reg[4][239]  ( .D(n1324), .CLK(clk), .Q(\ram[4][239] ) );
  DFFX1_HVT \ram_reg[4][238]  ( .D(n1323), .CLK(clk), .Q(\ram[4][238] ) );
  DFFX1_HVT \ram_reg[4][237]  ( .D(n1322), .CLK(clk), .Q(\ram[4][237] ) );
  DFFX1_HVT \ram_reg[4][236]  ( .D(n1321), .CLK(clk), .Q(\ram[4][236] ) );
  DFFX1_HVT \ram_reg[4][235]  ( .D(n1320), .CLK(clk), .Q(\ram[4][235] ) );
  DFFX1_HVT \ram_reg[4][234]  ( .D(n1319), .CLK(clk), .Q(\ram[4][234] ), .QN(
        n5718) );
  DFFX1_HVT \ram_reg[4][233]  ( .D(n1318), .CLK(clk), .Q(\ram[4][233] ) );
  DFFX1_HVT \ram_reg[4][232]  ( .D(n1317), .CLK(clk), .Q(\ram[4][232] ) );
  DFFX1_HVT \ram_reg[4][231]  ( .D(n1316), .CLK(clk), .Q(\ram[4][231] ) );
  DFFX1_HVT \ram_reg[4][230]  ( .D(n1315), .CLK(clk), .Q(\ram[4][230] ) );
  DFFX1_HVT \ram_reg[4][229]  ( .D(n1314), .CLK(clk), .Q(\ram[4][229] ) );
  DFFX1_HVT \ram_reg[4][228]  ( .D(n1313), .CLK(clk), .Q(\ram[4][228] ) );
  DFFX1_HVT \ram_reg[4][227]  ( .D(n1312), .CLK(clk), .Q(\ram[4][227] ) );
  DFFX1_HVT \ram_reg[4][226]  ( .D(n1311), .CLK(clk), .Q(\ram[4][226] ) );
  DFFX1_HVT \ram_reg[4][225]  ( .D(n1310), .CLK(clk), .Q(\ram[4][225] ) );
  DFFX1_HVT \ram_reg[4][224]  ( .D(n1309), .CLK(clk), .Q(\ram[4][224] ) );
  DFFX1_HVT \ram_reg[4][223]  ( .D(n1308), .CLK(clk), .Q(\ram[4][223] ) );
  DFFX1_HVT \ram_reg[4][222]  ( .D(n1307), .CLK(clk), .Q(\ram[4][222] ) );
  DFFX1_HVT \ram_reg[4][221]  ( .D(n1306), .CLK(clk), .Q(\ram[4][221] ) );
  DFFX1_HVT \ram_reg[4][220]  ( .D(n1305), .CLK(clk), .Q(\ram[4][220] ) );
  DFFX1_HVT \ram_reg[4][219]  ( .D(n1304), .CLK(clk), .Q(\ram[4][219] ) );
  DFFX1_HVT \ram_reg[4][218]  ( .D(n1303), .CLK(clk), .Q(\ram[4][218] ) );
  DFFX1_HVT \ram_reg[4][217]  ( .D(n1302), .CLK(clk), .Q(\ram[4][217] ) );
  DFFX1_HVT \ram_reg[4][216]  ( .D(n1301), .CLK(clk), .Q(\ram[4][216] ) );
  DFFX1_HVT \ram_reg[4][215]  ( .D(n1300), .CLK(clk), .Q(\ram[4][215] ) );
  DFFX1_HVT \ram_reg[4][214]  ( .D(n1299), .CLK(clk), .Q(\ram[4][214] ) );
  DFFX1_HVT \ram_reg[4][213]  ( .D(n1298), .CLK(clk), .Q(\ram[4][213] ), .QN(
        n5453) );
  DFFX1_HVT \ram_reg[4][212]  ( .D(n1297), .CLK(clk), .Q(\ram[4][212] ) );
  DFFX1_HVT \ram_reg[4][211]  ( .D(n1296), .CLK(clk), .Q(\ram[4][211] ) );
  DFFX1_HVT \ram_reg[4][210]  ( .D(n1295), .CLK(clk), .Q(\ram[4][210] ) );
  DFFX1_HVT \ram_reg[4][209]  ( .D(n1294), .CLK(clk), .Q(\ram[4][209] ) );
  DFFX1_HVT \ram_reg[4][208]  ( .D(n1293), .CLK(clk), .Q(\ram[4][208] ) );
  DFFX1_HVT \ram_reg[4][207]  ( .D(n1292), .CLK(clk), .Q(\ram[4][207] ) );
  DFFX1_HVT \ram_reg[4][206]  ( .D(n1291), .CLK(clk), .Q(\ram[4][206] ) );
  DFFX1_HVT \ram_reg[4][205]  ( .D(n1290), .CLK(clk), .Q(\ram[4][205] ) );
  DFFX1_HVT \ram_reg[4][204]  ( .D(n1289), .CLK(clk), .Q(\ram[4][204] ) );
  DFFX1_HVT \ram_reg[4][203]  ( .D(n1288), .CLK(clk), .Q(\ram[4][203] ) );
  DFFX1_HVT \ram_reg[4][202]  ( .D(n1287), .CLK(clk), .Q(\ram[4][202] ) );
  DFFX1_HVT \ram_reg[4][201]  ( .D(n1286), .CLK(clk), .Q(\ram[4][201] ) );
  DFFX1_HVT \ram_reg[4][200]  ( .D(n1285), .CLK(clk), .Q(\ram[4][200] ) );
  DFFX1_HVT \ram_reg[4][199]  ( .D(n1284), .CLK(clk), .Q(\ram[4][199] ) );
  DFFX1_HVT \ram_reg[4][198]  ( .D(n1283), .CLK(clk), .Q(\ram[4][198] ) );
  DFFX1_HVT \ram_reg[4][197]  ( .D(n1282), .CLK(clk), .Q(\ram[4][197] ) );
  DFFX1_HVT \ram_reg[4][196]  ( .D(n1281), .CLK(clk), .Q(\ram[4][196] ) );
  DFFX1_HVT \ram_reg[4][195]  ( .D(n1280), .CLK(clk), .Q(\ram[4][195] ), .QN(
        n4319) );
  DFFX1_HVT \ram_reg[4][194]  ( .D(n1279), .CLK(clk), .Q(\ram[4][194] ) );
  DFFX1_HVT \ram_reg[4][193]  ( .D(n1278), .CLK(clk), .Q(\ram[4][193] ) );
  DFFX1_HVT \ram_reg[4][192]  ( .D(n1277), .CLK(clk), .Q(\ram[4][192] ) );
  DFFX1_HVT \ram_reg[4][191]  ( .D(n1276), .CLK(clk), .Q(\ram[4][191] ) );
  DFFX1_HVT \ram_reg[4][190]  ( .D(n1275), .CLK(clk), .Q(\ram[4][190] ) );
  DFFX1_HVT \ram_reg[4][189]  ( .D(n1274), .CLK(clk), .Q(\ram[4][189] ) );
  DFFX1_HVT \ram_reg[4][188]  ( .D(n1273), .CLK(clk), .Q(\ram[4][188] ) );
  DFFX1_HVT \ram_reg[4][187]  ( .D(n1272), .CLK(clk), .Q(\ram[4][187] ) );
  DFFX1_HVT \ram_reg[4][186]  ( .D(n1271), .CLK(clk), .Q(\ram[4][186] ) );
  DFFX1_HVT \ram_reg[4][185]  ( .D(n1270), .CLK(clk), .Q(\ram[4][185] ) );
  DFFX1_HVT \ram_reg[4][184]  ( .D(n1269), .CLK(clk), .Q(\ram[4][184] ) );
  DFFX1_HVT \ram_reg[4][183]  ( .D(n1268), .CLK(clk), .Q(\ram[4][183] ) );
  DFFX1_HVT \ram_reg[4][182]  ( .D(n1267), .CLK(clk), .Q(\ram[4][182] ) );
  DFFX1_HVT \ram_reg[4][181]  ( .D(n1266), .CLK(clk), .Q(\ram[4][181] ) );
  DFFX1_HVT \ram_reg[4][180]  ( .D(n1265), .CLK(clk), .Q(\ram[4][180] ) );
  DFFX1_HVT \ram_reg[4][179]  ( .D(n1264), .CLK(clk), .Q(\ram[4][179] ) );
  DFFX1_HVT \ram_reg[4][178]  ( .D(n1263), .CLK(clk), .Q(\ram[4][178] ) );
  DFFX1_HVT \ram_reg[4][177]  ( .D(n1262), .CLK(clk), .Q(\ram[4][177] ) );
  DFFX1_HVT \ram_reg[4][176]  ( .D(n1261), .CLK(clk), .Q(\ram[4][176] ) );
  DFFX1_HVT \ram_reg[4][175]  ( .D(n1260), .CLK(clk), .Q(\ram[4][175] ) );
  DFFX1_HVT \ram_reg[4][174]  ( .D(n1259), .CLK(clk), .Q(\ram[4][174] ) );
  DFFX1_HVT \ram_reg[4][173]  ( .D(n1258), .CLK(clk), .Q(\ram[4][173] ) );
  DFFX1_HVT \ram_reg[4][172]  ( .D(n1257), .CLK(clk), .Q(\ram[4][172] ) );
  DFFX1_HVT \ram_reg[4][171]  ( .D(n1256), .CLK(clk), .Q(\ram[4][171] ) );
  DFFX1_HVT \ram_reg[4][170]  ( .D(n1255), .CLK(clk), .Q(\ram[4][170] ) );
  DFFX1_HVT \ram_reg[4][169]  ( .D(n1254), .CLK(clk), .Q(\ram[4][169] ) );
  DFFX1_HVT \ram_reg[4][168]  ( .D(n1253), .CLK(clk), .Q(\ram[4][168] ) );
  DFFX1_HVT \ram_reg[4][167]  ( .D(n1252), .CLK(clk), .Q(\ram[4][167] ) );
  DFFX1_HVT \ram_reg[4][166]  ( .D(n1251), .CLK(clk), .Q(\ram[4][166] ) );
  DFFX1_HVT \ram_reg[4][165]  ( .D(n1250), .CLK(clk), .Q(\ram[4][165] ) );
  DFFX1_HVT \ram_reg[4][164]  ( .D(n1249), .CLK(clk), .Q(\ram[4][164] ) );
  DFFX1_HVT \ram_reg[4][163]  ( .D(n1248), .CLK(clk), .Q(\ram[4][163] ) );
  DFFX1_HVT \ram_reg[4][162]  ( .D(n1247), .CLK(clk), .Q(\ram[4][162] ) );
  DFFX1_HVT \ram_reg[4][161]  ( .D(n1246), .CLK(clk), .Q(\ram[4][161] ) );
  DFFX1_HVT \ram_reg[4][160]  ( .D(n1245), .CLK(clk), .Q(\ram[4][160] ) );
  DFFX1_HVT \ram_reg[4][159]  ( .D(n1244), .CLK(clk), .Q(\ram[4][159] ) );
  DFFX1_HVT \ram_reg[4][158]  ( .D(n1243), .CLK(clk), .Q(\ram[4][158] ) );
  DFFX1_HVT \ram_reg[4][157]  ( .D(n1242), .CLK(clk), .Q(\ram[4][157] ) );
  DFFX1_HVT \ram_reg[4][156]  ( .D(n1241), .CLK(clk), .Q(\ram[4][156] ) );
  DFFX1_HVT \ram_reg[4][155]  ( .D(n1240), .CLK(clk), .Q(\ram[4][155] ) );
  DFFX1_HVT \ram_reg[4][154]  ( .D(n1239), .CLK(clk), .Q(\ram[4][154] ) );
  DFFX1_HVT \ram_reg[4][153]  ( .D(n1238), .CLK(clk), .Q(\ram[4][153] ) );
  DFFX1_HVT \ram_reg[4][152]  ( .D(n1237), .CLK(clk), .Q(\ram[4][152] ) );
  DFFX1_HVT \ram_reg[4][151]  ( .D(n1236), .CLK(clk), .Q(\ram[4][151] ) );
  DFFX1_HVT \ram_reg[4][150]  ( .D(n1235), .CLK(clk), .Q(\ram[4][150] ) );
  DFFX1_HVT \ram_reg[4][149]  ( .D(n1234), .CLK(clk), .Q(\ram[4][149] ) );
  DFFX1_HVT \ram_reg[4][148]  ( .D(n1233), .CLK(clk), .Q(\ram[4][148] ) );
  DFFX1_HVT \ram_reg[4][147]  ( .D(n1232), .CLK(clk), .Q(\ram[4][147] ) );
  DFFX1_HVT \ram_reg[4][146]  ( .D(n1231), .CLK(clk), .Q(\ram[4][146] ) );
  DFFX1_HVT \ram_reg[4][145]  ( .D(n1230), .CLK(clk), .Q(\ram[4][145] ) );
  DFFX1_HVT \ram_reg[4][144]  ( .D(n1229), .CLK(clk), .Q(\ram[4][144] ) );
  DFFX1_HVT \ram_reg[4][143]  ( .D(n1228), .CLK(clk), .Q(\ram[4][143] ) );
  DFFX1_HVT \ram_reg[4][142]  ( .D(n1227), .CLK(clk), .Q(\ram[4][142] ) );
  DFFX1_HVT \ram_reg[4][141]  ( .D(n1226), .CLK(clk), .Q(\ram[4][141] ), .QN(
        n4292) );
  DFFX1_HVT \ram_reg[4][140]  ( .D(n1225), .CLK(clk), .Q(\ram[4][140] ) );
  DFFX1_HVT \ram_reg[4][139]  ( .D(n1224), .CLK(clk), .Q(\ram[4][139] ), .QN(
        n4591) );
  DFFX1_HVT \ram_reg[4][138]  ( .D(n1223), .CLK(clk), .Q(\ram[4][138] ) );
  DFFX1_HVT \ram_reg[4][137]  ( .D(n1222), .CLK(clk), .Q(\ram[4][137] ) );
  DFFX1_HVT \ram_reg[4][136]  ( .D(n1221), .CLK(clk), .Q(\ram[4][136] ) );
  DFFX1_HVT \ram_reg[4][135]  ( .D(n1220), .CLK(clk), .Q(\ram[4][135] ) );
  DFFX1_HVT \ram_reg[4][134]  ( .D(n1219), .CLK(clk), .Q(\ram[4][134] ) );
  DFFX1_HVT \ram_reg[4][133]  ( .D(n1218), .CLK(clk), .Q(\ram[4][133] ) );
  DFFX1_HVT \ram_reg[4][132]  ( .D(n1217), .CLK(clk), .Q(\ram[4][132] ) );
  DFFX1_HVT \ram_reg[4][131]  ( .D(n1216), .CLK(clk), .Q(\ram[4][131] ), .QN(
        n4633) );
  DFFX1_HVT \ram_reg[4][130]  ( .D(n1215), .CLK(clk), .Q(\ram[4][130] ) );
  DFFX1_HVT \ram_reg[4][129]  ( .D(n1214), .CLK(clk), .Q(\ram[4][129] ) );
  DFFX1_HVT \ram_reg[4][128]  ( .D(n1213), .CLK(clk), .Q(\ram[4][128] ) );
  DFFX1_HVT \ram_reg[4][127]  ( .D(n1212), .CLK(clk), .Q(\ram[4][127] ) );
  DFFX1_HVT \ram_reg[4][126]  ( .D(n1211), .CLK(clk), .Q(\ram[4][126] ) );
  DFFX1_HVT \ram_reg[4][125]  ( .D(n1210), .CLK(clk), .Q(\ram[4][125] ) );
  DFFX1_HVT \ram_reg[4][124]  ( .D(n1209), .CLK(clk), .Q(\ram[4][124] ) );
  DFFX1_HVT \ram_reg[4][123]  ( .D(n1208), .CLK(clk), .Q(\ram[4][123] ) );
  DFFX1_HVT \ram_reg[4][122]  ( .D(n1207), .CLK(clk), .Q(\ram[4][122] ) );
  DFFX1_HVT \ram_reg[4][121]  ( .D(n1206), .CLK(clk), .Q(\ram[4][121] ), .QN(
        n5100) );
  DFFX1_HVT \ram_reg[4][120]  ( .D(n1205), .CLK(clk), .Q(\ram[4][120] ) );
  DFFX1_HVT \ram_reg[4][119]  ( .D(n1204), .CLK(clk), .Q(\ram[4][119] ) );
  DFFX1_HVT \ram_reg[4][118]  ( .D(n1203), .CLK(clk), .Q(\ram[4][118] ) );
  DFFX1_HVT \ram_reg[4][117]  ( .D(n1202), .CLK(clk), .Q(\ram[4][117] ) );
  DFFX1_HVT \ram_reg[4][116]  ( .D(n1201), .CLK(clk), .Q(\ram[4][116] ) );
  DFFX1_HVT \ram_reg[4][115]  ( .D(n1200), .CLK(clk), .Q(\ram[4][115] ) );
  DFFX1_HVT \ram_reg[4][114]  ( .D(n1199), .CLK(clk), .Q(\ram[4][114] ) );
  DFFX1_HVT \ram_reg[4][113]  ( .D(n1198), .CLK(clk), .Q(\ram[4][113] ) );
  DFFX1_HVT \ram_reg[4][112]  ( .D(n1197), .CLK(clk), .Q(\ram[4][112] ) );
  DFFX1_HVT \ram_reg[4][111]  ( .D(n1196), .CLK(clk), .Q(\ram[4][111] ) );
  DFFX1_HVT \ram_reg[4][110]  ( .D(n1195), .CLK(clk), .Q(\ram[4][110] ) );
  DFFX1_HVT \ram_reg[4][109]  ( .D(n1194), .CLK(clk), .Q(\ram[4][109] ) );
  DFFX1_HVT \ram_reg[4][108]  ( .D(n1193), .CLK(clk), .Q(\ram[4][108] ) );
  DFFX1_HVT \ram_reg[4][107]  ( .D(n1192), .CLK(clk), .Q(\ram[4][107] ) );
  DFFX1_HVT \ram_reg[4][106]  ( .D(n1191), .CLK(clk), .Q(\ram[4][106] ) );
  DFFX1_HVT \ram_reg[4][105]  ( .D(n1190), .CLK(clk), .Q(\ram[4][105] ) );
  DFFX1_HVT \ram_reg[4][104]  ( .D(n1189), .CLK(clk), .Q(\ram[4][104] ) );
  DFFX1_HVT \ram_reg[4][103]  ( .D(n1188), .CLK(clk), .Q(\ram[4][103] ) );
  DFFX1_HVT \ram_reg[4][102]  ( .D(n1187), .CLK(clk), .Q(\ram[4][102] ) );
  DFFX1_HVT \ram_reg[4][101]  ( .D(n1186), .CLK(clk), .Q(\ram[4][101] ) );
  DFFX1_HVT \ram_reg[4][100]  ( .D(n1185), .CLK(clk), .Q(\ram[4][100] ) );
  DFFX1_HVT \ram_reg[4][99]  ( .D(n1184), .CLK(clk), .Q(\ram[4][99] ) );
  DFFX1_HVT \ram_reg[4][98]  ( .D(n1183), .CLK(clk), .Q(\ram[4][98] ) );
  DFFX1_HVT \ram_reg[4][97]  ( .D(n1182), .CLK(clk), .Q(\ram[4][97] ) );
  DFFX1_HVT \ram_reg[4][96]  ( .D(n1181), .CLK(clk), .Q(\ram[4][96] ) );
  DFFX1_HVT \ram_reg[4][95]  ( .D(n1180), .CLK(clk), .Q(\ram[4][95] ) );
  DFFX1_HVT \ram_reg[4][94]  ( .D(n1179), .CLK(clk), .Q(\ram[4][94] ) );
  DFFX1_HVT \ram_reg[4][93]  ( .D(n1178), .CLK(clk), .Q(\ram[4][93] ) );
  DFFX1_HVT \ram_reg[4][92]  ( .D(n1177), .CLK(clk), .Q(\ram[4][92] ) );
  DFFX1_HVT \ram_reg[4][91]  ( .D(n1176), .CLK(clk), .Q(\ram[4][91] ) );
  DFFX1_HVT \ram_reg[4][90]  ( .D(n1175), .CLK(clk), .Q(\ram[4][90] ) );
  DFFX1_HVT \ram_reg[4][89]  ( .D(n1174), .CLK(clk), .Q(\ram[4][89] ) );
  DFFX1_HVT \ram_reg[4][88]  ( .D(n1173), .CLK(clk), .Q(\ram[4][88] ) );
  DFFX1_HVT \ram_reg[4][87]  ( .D(n1172), .CLK(clk), .Q(\ram[4][87] ) );
  DFFX1_HVT \ram_reg[4][86]  ( .D(n1171), .CLK(clk), .Q(\ram[4][86] ) );
  DFFX1_HVT \ram_reg[4][85]  ( .D(n1170), .CLK(clk), .Q(\ram[4][85] ) );
  DFFX1_HVT \ram_reg[4][84]  ( .D(n1169), .CLK(clk), .Q(\ram[4][84] ) );
  DFFX1_HVT \ram_reg[4][83]  ( .D(n1168), .CLK(clk), .Q(\ram[4][83] ) );
  DFFX1_HVT \ram_reg[4][82]  ( .D(n1167), .CLK(clk), .Q(\ram[4][82] ) );
  DFFX1_HVT \ram_reg[4][81]  ( .D(n1166), .CLK(clk), .Q(\ram[4][81] ) );
  DFFX1_HVT \ram_reg[4][80]  ( .D(n1165), .CLK(clk), .Q(\ram[4][80] ) );
  DFFX1_HVT \ram_reg[4][79]  ( .D(n1164), .CLK(clk), .Q(\ram[4][79] ) );
  DFFX1_HVT \ram_reg[4][78]  ( .D(n1163), .CLK(clk), .Q(\ram[4][78] ) );
  DFFX1_HVT \ram_reg[4][77]  ( .D(n1162), .CLK(clk), .Q(\ram[4][77] ) );
  DFFX1_HVT \ram_reg[4][76]  ( .D(n1161), .CLK(clk), .Q(\ram[4][76] ) );
  DFFX1_HVT \ram_reg[4][75]  ( .D(n1160), .CLK(clk), .Q(\ram[4][75] ) );
  DFFX1_HVT \ram_reg[4][74]  ( .D(n1159), .CLK(clk), .Q(\ram[4][74] ) );
  DFFX1_HVT \ram_reg[4][73]  ( .D(n1158), .CLK(clk), .Q(\ram[4][73] ) );
  DFFX1_HVT \ram_reg[4][72]  ( .D(n1157), .CLK(clk), .Q(\ram[4][72] ) );
  DFFX1_HVT \ram_reg[4][71]  ( .D(n1156), .CLK(clk), .Q(\ram[4][71] ) );
  DFFX1_HVT \ram_reg[4][70]  ( .D(n1155), .CLK(clk), .Q(\ram[4][70] ) );
  DFFX1_HVT \ram_reg[4][69]  ( .D(n1154), .CLK(clk), .Q(\ram[4][69] ) );
  DFFX1_HVT \ram_reg[4][68]  ( .D(n1153), .CLK(clk), .Q(\ram[4][68] ) );
  DFFX1_HVT \ram_reg[4][67]  ( .D(n1152), .CLK(clk), .Q(\ram[4][67] ), .QN(
        n4821) );
  DFFX1_HVT \ram_reg[4][66]  ( .D(n1151), .CLK(clk), .Q(\ram[4][66] ) );
  DFFX1_HVT \ram_reg[4][65]  ( .D(n1150), .CLK(clk), .Q(\ram[4][65] ) );
  DFFX1_HVT \ram_reg[4][64]  ( .D(n1149), .CLK(clk), .Q(\ram[4][64] ) );
  DFFX1_HVT \ram_reg[4][63]  ( .D(n1148), .CLK(clk), .Q(\ram[4][63] ) );
  DFFX1_HVT \ram_reg[4][62]  ( .D(n1147), .CLK(clk), .Q(\ram[4][62] ) );
  DFFX1_HVT \ram_reg[4][61]  ( .D(n1146), .CLK(clk), .Q(\ram[4][61] ) );
  DFFX1_HVT \ram_reg[4][60]  ( .D(n1145), .CLK(clk), .Q(\ram[4][60] ) );
  DFFX1_HVT \ram_reg[4][59]  ( .D(n5027), .CLK(clk), .Q(\ram[4][59] ) );
  DFFX1_HVT \ram_reg[4][58]  ( .D(n1143), .CLK(clk), .Q(\ram[4][58] ) );
  DFFX1_HVT \ram_reg[4][57]  ( .D(n1142), .CLK(clk), .Q(\ram[4][57] ) );
  DFFX1_HVT \ram_reg[4][56]  ( .D(n1141), .CLK(clk), .Q(\ram[4][56] ) );
  DFFX1_HVT \ram_reg[4][55]  ( .D(n1140), .CLK(clk), .Q(\ram[4][55] ) );
  DFFX1_HVT \ram_reg[4][54]  ( .D(n1139), .CLK(clk), .Q(\ram[4][54] ), .QN(
        n4806) );
  DFFX1_HVT \ram_reg[4][53]  ( .D(n1138), .CLK(clk), .Q(\ram[4][53] ) );
  DFFX1_HVT \ram_reg[4][52]  ( .D(n5028), .CLK(clk), .Q(\ram[4][52] ) );
  DFFX1_HVT \ram_reg[4][51]  ( .D(n1136), .CLK(clk), .Q(\ram[4][51] ) );
  DFFX1_HVT \ram_reg[4][50]  ( .D(n1135), .CLK(clk), .Q(\ram[4][50] ), .QN(
        n5065) );
  DFFX1_HVT \ram_reg[4][49]  ( .D(n1134), .CLK(clk), .Q(\ram[4][49] ) );
  DFFX1_HVT \ram_reg[4][48]  ( .D(n1133), .CLK(clk), .Q(\ram[4][48] ), .QN(
        n4960) );
  DFFX1_HVT \ram_reg[4][47]  ( .D(n1132), .CLK(clk), .Q(\ram[4][47] ) );
  DFFX1_HVT \ram_reg[4][46]  ( .D(n1131), .CLK(clk), .Q(\ram[4][46] ) );
  DFFX1_HVT \ram_reg[4][45]  ( .D(n1130), .CLK(clk), .Q(\ram[4][45] ) );
  DFFX1_HVT \ram_reg[4][44]  ( .D(n1129), .CLK(clk), .Q(\ram[4][44] ) );
  DFFX1_HVT \ram_reg[4][43]  ( .D(n1128), .CLK(clk), .Q(\ram[4][43] ) );
  DFFX1_HVT \ram_reg[4][42]  ( .D(n1127), .CLK(clk), .Q(\ram[4][42] ), .QN(
        n5547) );
  DFFX1_HVT \ram_reg[4][41]  ( .D(n1126), .CLK(clk), .Q(\ram[4][41] ) );
  DFFX1_HVT \ram_reg[4][40]  ( .D(n1125), .CLK(clk), .Q(\ram[4][40] ) );
  DFFX1_HVT \ram_reg[4][39]  ( .D(n1124), .CLK(clk), .Q(\ram[4][39] ), .QN(
        n4967) );
  DFFX1_HVT \ram_reg[4][38]  ( .D(n1123), .CLK(clk), .Q(\ram[4][38] ) );
  DFFX1_HVT \ram_reg[4][37]  ( .D(n1122), .CLK(clk), .Q(\ram[4][37] ) );
  DFFX1_HVT \ram_reg[4][36]  ( .D(n1121), .CLK(clk), .Q(\ram[4][36] ), .QN(
        n5548) );
  DFFX1_HVT \ram_reg[4][35]  ( .D(n1120), .CLK(clk), .Q(\ram[4][35] ) );
  DFFX1_HVT \ram_reg[4][34]  ( .D(n1119), .CLK(clk), .Q(\ram[4][34] ) );
  DFFX1_HVT \ram_reg[4][33]  ( .D(n1118), .CLK(clk), .Q(\ram[4][33] ) );
  DFFX1_HVT \ram_reg[4][32]  ( .D(n1117), .CLK(clk), .Q(\ram[4][32] ) );
  DFFX1_HVT \ram_reg[4][31]  ( .D(n1116), .CLK(clk), .Q(\ram[4][31] ) );
  DFFX1_HVT \ram_reg[4][30]  ( .D(n1115), .CLK(clk), .Q(\ram[4][30] ) );
  DFFX1_HVT \ram_reg[4][29]  ( .D(n1114), .CLK(clk), .Q(\ram[4][29] ), .QN(
        n5452) );
  DFFX1_HVT \ram_reg[4][28]  ( .D(n1113), .CLK(clk), .Q(\ram[4][28] ) );
  DFFX1_HVT \ram_reg[4][27]  ( .D(n1112), .CLK(clk), .Q(\ram[4][27] ), .QN(
        n5549) );
  DFFX1_HVT \ram_reg[4][26]  ( .D(n1111), .CLK(clk), .Q(\ram[4][26] ) );
  DFFX1_HVT \ram_reg[4][25]  ( .D(n1110), .CLK(clk), .Q(\ram[4][25] ), .QN(
        n5550) );
  DFFX1_HVT \ram_reg[4][24]  ( .D(n1109), .CLK(clk), .Q(\ram[4][24] ) );
  DFFX1_HVT \ram_reg[4][23]  ( .D(n1108), .CLK(clk), .Q(\ram[4][23] ) );
  DFFX1_HVT \ram_reg[4][22]  ( .D(n1107), .CLK(clk), .Q(\ram[4][22] ) );
  DFFX1_HVT \ram_reg[4][21]  ( .D(n1106), .CLK(clk), .Q(\ram[4][21] ), .QN(
        n5725) );
  DFFX1_HVT \ram_reg[4][20]  ( .D(n1105), .CLK(clk), .QN(n6555) );
  DFFX1_HVT \ram_reg[4][19]  ( .D(n1104), .CLK(clk), .Q(\ram[4][19] ) );
  DFFX1_HVT \ram_reg[4][18]  ( .D(n1103), .CLK(clk), .Q(\ram[4][18] ) );
  DFFX1_HVT \ram_reg[4][17]  ( .D(n1102), .CLK(clk), .Q(\ram[4][17] ) );
  DFFX1_HVT \ram_reg[4][16]  ( .D(n1101), .CLK(clk), .Q(\ram[4][16] ) );
  DFFX1_HVT \ram_reg[4][15]  ( .D(n1100), .CLK(clk), .Q(\ram[4][15] ) );
  DFFX1_HVT \ram_reg[4][14]  ( .D(n1099), .CLK(clk), .Q(\ram[4][14] ) );
  DFFX1_HVT \ram_reg[4][13]  ( .D(n1098), .CLK(clk), .Q(\ram[4][13] ) );
  DFFX1_HVT \ram_reg[4][12]  ( .D(n1097), .CLK(clk), .Q(\ram[4][12] ), .QN(
        n5198) );
  DFFX1_HVT \ram_reg[4][11]  ( .D(n1096), .CLK(clk), .Q(\ram[4][11] ) );
  DFFX1_HVT \ram_reg[4][10]  ( .D(n1095), .CLK(clk), .Q(\ram[4][10] ), .QN(
        n5068) );
  DFFX1_HVT \ram_reg[4][9]  ( .D(n1094), .CLK(clk), .Q(\ram[4][9] ), .QN(n5726) );
  DFFX1_HVT \ram_reg[4][8]  ( .D(n1093), .CLK(clk), .Q(\ram[4][8] ), .QN(n5727) );
  DFFX1_HVT \ram_reg[4][7]  ( .D(n1092), .CLK(clk), .Q(\ram[4][7] ), .QN(n5086) );
  DFFX1_HVT \ram_reg[4][6]  ( .D(n1091), .CLK(clk), .Q(\ram[4][6] ), .QN(n5146) );
  DFFX1_HVT \ram_reg[4][5]  ( .D(n1090), .CLK(clk), .Q(\ram[4][5] ) );
  DFFX1_HVT \ram_reg[4][4]  ( .D(n1089), .CLK(clk), .Q(\ram[4][4] ) );
  DFFX1_HVT \ram_reg[4][3]  ( .D(n1088), .CLK(clk), .Q(\ram[4][3] ) );
  DFFX1_HVT \ram_reg[4][2]  ( .D(n1087), .CLK(clk), .Q(\ram[4][2] ) );
  DFFX1_HVT \ram_reg[4][1]  ( .D(n1086), .CLK(clk), .Q(\ram[4][1] ) );
  DFFX1_HVT \ram_reg[4][0]  ( .D(n1085), .CLK(clk), .Q(\ram[4][0] ) );
  DFFX1_HVT \ram_reg[3][255]  ( .D(n1084), .CLK(clk), .Q(\ram[3][255] ) );
  DFFX1_HVT \ram_reg[3][254]  ( .D(n1083), .CLK(clk), .Q(\ram[3][254] ) );
  DFFX1_HVT \ram_reg[3][253]  ( .D(n1082), .CLK(clk), .Q(\ram[3][253] ) );
  DFFX1_HVT \ram_reg[3][252]  ( .D(n1081), .CLK(clk), .Q(\ram[3][252] ) );
  DFFX1_HVT \ram_reg[3][251]  ( .D(n1080), .CLK(clk), .Q(\ram[3][251] ) );
  DFFX1_HVT \ram_reg[3][250]  ( .D(n1079), .CLK(clk), .Q(\ram[3][250] ) );
  DFFX1_HVT \ram_reg[3][249]  ( .D(n5029), .CLK(clk), .Q(\ram[3][249] ), .QN(
        n5330) );
  DFFX1_HVT \ram_reg[3][248]  ( .D(n1077), .CLK(clk), .Q(\ram[3][248] ) );
  DFFX1_HVT \ram_reg[3][247]  ( .D(n1076), .CLK(clk), .Q(\ram[3][247] ) );
  DFFX1_HVT \ram_reg[3][246]  ( .D(n1075), .CLK(clk), .Q(\ram[3][246] ) );
  DFFX1_HVT \ram_reg[3][245]  ( .D(n1074), .CLK(clk), .Q(\ram[3][245] ) );
  DFFX1_HVT \ram_reg[3][244]  ( .D(n1073), .CLK(clk), .Q(\ram[3][244] ) );
  DFFX1_HVT \ram_reg[3][243]  ( .D(n1072), .CLK(clk), .Q(\ram[3][243] ) );
  DFFX1_HVT \ram_reg[3][242]  ( .D(n1071), .CLK(clk), .Q(\ram[3][242] ) );
  DFFX1_HVT \ram_reg[3][241]  ( .D(n1070), .CLK(clk), .Q(\ram[3][241] ) );
  DFFX1_HVT \ram_reg[3][240]  ( .D(n1069), .CLK(clk), .Q(\ram[3][240] ) );
  DFFX1_HVT \ram_reg[3][239]  ( .D(n1068), .CLK(clk), .Q(\ram[3][239] ) );
  DFFX1_HVT \ram_reg[3][238]  ( .D(n1067), .CLK(clk), .Q(\ram[3][238] ) );
  DFFX1_HVT \ram_reg[3][237]  ( .D(n1066), .CLK(clk), .Q(\ram[3][237] ) );
  DFFX1_HVT \ram_reg[3][236]  ( .D(n1065), .CLK(clk), .Q(\ram[3][236] ) );
  DFFX1_HVT \ram_reg[3][235]  ( .D(n1064), .CLK(clk), .Q(\ram[3][235] ) );
  DFFX1_HVT \ram_reg[3][234]  ( .D(n1063), .CLK(clk), .Q(\ram[3][234] ) );
  DFFX1_HVT \ram_reg[3][233]  ( .D(n1062), .CLK(clk), .Q(\ram[3][233] ) );
  DFFX1_HVT \ram_reg[3][232]  ( .D(n1061), .CLK(clk), .Q(\ram[3][232] ) );
  DFFX1_HVT \ram_reg[3][231]  ( .D(n1060), .CLK(clk), .Q(\ram[3][231] ) );
  DFFX1_HVT \ram_reg[3][230]  ( .D(n1059), .CLK(clk), .Q(\ram[3][230] ) );
  DFFX1_HVT \ram_reg[3][229]  ( .D(n1058), .CLK(clk), .Q(\ram[3][229] ) );
  DFFX1_HVT \ram_reg[3][228]  ( .D(n1057), .CLK(clk), .Q(\ram[3][228] ) );
  DFFX1_HVT \ram_reg[3][227]  ( .D(n1056), .CLK(clk), .Q(\ram[3][227] ) );
  DFFX1_HVT \ram_reg[3][226]  ( .D(n1055), .CLK(clk), .Q(\ram[3][226] ) );
  DFFX1_HVT \ram_reg[3][225]  ( .D(n1054), .CLK(clk), .Q(\ram[3][225] ) );
  DFFX1_HVT \ram_reg[3][224]  ( .D(n1053), .CLK(clk), .Q(\ram[3][224] ), .QN(
        n5033) );
  DFFX1_HVT \ram_reg[3][223]  ( .D(n1052), .CLK(clk), .Q(\ram[3][223] ), .QN(
        n4336) );
  DFFX1_HVT \ram_reg[3][222]  ( .D(n1051), .CLK(clk), .Q(\ram[3][222] ) );
  DFFX1_HVT \ram_reg[3][221]  ( .D(n1050), .CLK(clk), .Q(\ram[3][221] ) );
  DFFX1_HVT \ram_reg[3][220]  ( .D(n1049), .CLK(clk), .Q(\ram[3][220] ) );
  DFFX1_HVT \ram_reg[3][219]  ( .D(n1048), .CLK(clk), .Q(\ram[3][219] ) );
  DFFX1_HVT \ram_reg[3][218]  ( .D(n1047), .CLK(clk), .Q(\ram[3][218] ) );
  DFFX1_HVT \ram_reg[3][217]  ( .D(n1046), .CLK(clk), .Q(\ram[3][217] ) );
  DFFX1_HVT \ram_reg[3][216]  ( .D(n1045), .CLK(clk), .Q(\ram[3][216] ) );
  DFFX1_HVT \ram_reg[3][215]  ( .D(n1044), .CLK(clk), .Q(\ram[3][215] ) );
  DFFX1_HVT \ram_reg[3][214]  ( .D(n1043), .CLK(clk), .Q(\ram[3][214] ) );
  DFFX1_HVT \ram_reg[3][213]  ( .D(n1042), .CLK(clk), .Q(\ram[3][213] ) );
  DFFX1_HVT \ram_reg[3][212]  ( .D(n1041), .CLK(clk), .Q(\ram[3][212] ) );
  DFFX1_HVT \ram_reg[3][211]  ( .D(n1040), .CLK(clk), .Q(\ram[3][211] ) );
  DFFX1_HVT \ram_reg[3][210]  ( .D(n1039), .CLK(clk), .Q(\ram[3][210] ) );
  DFFX1_HVT \ram_reg[3][209]  ( .D(n1038), .CLK(clk), .Q(\ram[3][209] ) );
  DFFX1_HVT \ram_reg[3][208]  ( .D(n1037), .CLK(clk), .Q(\ram[3][208] ) );
  DFFX1_HVT \ram_reg[3][207]  ( .D(n1036), .CLK(clk), .Q(\ram[3][207] ) );
  DFFX1_HVT \ram_reg[3][206]  ( .D(n1035), .CLK(clk), .Q(\ram[3][206] ) );
  DFFX1_HVT \ram_reg[3][205]  ( .D(n1034), .CLK(clk), .Q(\ram[3][205] ) );
  DFFX1_HVT \ram_reg[3][204]  ( .D(n1033), .CLK(clk), .Q(\ram[3][204] ) );
  DFFX1_HVT \ram_reg[3][203]  ( .D(n1032), .CLK(clk), .Q(\ram[3][203] ) );
  DFFX1_HVT \ram_reg[3][202]  ( .D(n1031), .CLK(clk), .Q(\ram[3][202] ) );
  DFFX1_HVT \ram_reg[3][201]  ( .D(n1030), .CLK(clk), .Q(\ram[3][201] ) );
  DFFX1_HVT \ram_reg[3][200]  ( .D(n1029), .CLK(clk), .Q(\ram[3][200] ) );
  DFFX1_HVT \ram_reg[3][199]  ( .D(n1028), .CLK(clk), .Q(\ram[3][199] ) );
  DFFX1_HVT \ram_reg[3][198]  ( .D(n1027), .CLK(clk), .Q(\ram[3][198] ) );
  DFFX1_HVT \ram_reg[3][197]  ( .D(n1026), .CLK(clk), .Q(\ram[3][197] ) );
  DFFX1_HVT \ram_reg[3][196]  ( .D(n1025), .CLK(clk), .Q(\ram[3][196] ) );
  DFFX1_HVT \ram_reg[3][195]  ( .D(n1024), .CLK(clk), .Q(\ram[3][195] ) );
  DFFX1_HVT \ram_reg[3][194]  ( .D(n5462), .CLK(clk), .Q(\ram[3][194] ), .QN(
        n5861) );
  DFFX1_HVT \ram_reg[3][193]  ( .D(n1022), .CLK(clk), .Q(\ram[3][193] ) );
  DFFX1_HVT \ram_reg[3][192]  ( .D(n1021), .CLK(clk), .Q(\ram[3][192] ) );
  DFFX1_HVT \ram_reg[3][191]  ( .D(n1020), .CLK(clk), .Q(\ram[3][191] ) );
  DFFX1_HVT \ram_reg[3][190]  ( .D(n1019), .CLK(clk), .Q(\ram[3][190] ) );
  DFFX1_HVT \ram_reg[3][189]  ( .D(n1018), .CLK(clk), .Q(\ram[3][189] ) );
  DFFX1_HVT \ram_reg[3][188]  ( .D(n1017), .CLK(clk), .Q(\ram[3][188] ) );
  DFFX1_HVT \ram_reg[3][187]  ( .D(n1016), .CLK(clk), .Q(\ram[3][187] ) );
  DFFX1_HVT \ram_reg[3][186]  ( .D(n1015), .CLK(clk), .Q(\ram[3][186] ) );
  DFFX1_HVT \ram_reg[3][185]  ( .D(n1014), .CLK(clk), .Q(\ram[3][185] ) );
  DFFX1_HVT \ram_reg[3][184]  ( .D(n1013), .CLK(clk), .Q(\ram[3][184] ) );
  DFFX1_HVT \ram_reg[3][183]  ( .D(n1012), .CLK(clk), .Q(\ram[3][183] ) );
  DFFX1_HVT \ram_reg[3][182]  ( .D(n1011), .CLK(clk), .Q(\ram[3][182] ), .QN(
        n4384) );
  DFFX1_HVT \ram_reg[3][181]  ( .D(n1010), .CLK(clk), .Q(\ram[3][181] ) );
  DFFX1_HVT \ram_reg[3][180]  ( .D(n1009), .CLK(clk), .Q(\ram[3][180] ) );
  DFFX1_HVT \ram_reg[3][179]  ( .D(n1008), .CLK(clk), .Q(\ram[3][179] ) );
  DFFX1_HVT \ram_reg[3][178]  ( .D(n1007), .CLK(clk), .Q(\ram[3][178] ) );
  DFFX1_HVT \ram_reg[3][177]  ( .D(n1006), .CLK(clk), .Q(\ram[3][177] ) );
  DFFX1_HVT \ram_reg[3][176]  ( .D(n1005), .CLK(clk), .Q(\ram[3][176] ) );
  DFFX1_HVT \ram_reg[3][175]  ( .D(n1004), .CLK(clk), .Q(\ram[3][175] ), .QN(
        n4253) );
  DFFX1_HVT \ram_reg[3][174]  ( .D(n1003), .CLK(clk), .Q(\ram[3][174] ) );
  DFFX1_HVT \ram_reg[3][173]  ( .D(n1002), .CLK(clk), .Q(\ram[3][173] ) );
  DFFX1_HVT \ram_reg[3][172]  ( .D(n1001), .CLK(clk), .Q(\ram[3][172] ) );
  DFFX1_HVT \ram_reg[3][171]  ( .D(n1000), .CLK(clk), .Q(\ram[3][171] ) );
  DFFX1_HVT \ram_reg[3][170]  ( .D(n999), .CLK(clk), .Q(\ram[3][170] ) );
  DFFX1_HVT \ram_reg[3][169]  ( .D(n998), .CLK(clk), .Q(\ram[3][169] ) );
  DFFX1_HVT \ram_reg[3][168]  ( .D(n997), .CLK(clk), .Q(\ram[3][168] ) );
  DFFX1_HVT \ram_reg[3][167]  ( .D(n996), .CLK(clk), .Q(\ram[3][167] ) );
  DFFX1_HVT \ram_reg[3][166]  ( .D(n995), .CLK(clk), .Q(\ram[3][166] ) );
  DFFX1_HVT \ram_reg[3][165]  ( .D(n994), .CLK(clk), .Q(\ram[3][165] ) );
  DFFX1_HVT \ram_reg[3][164]  ( .D(n993), .CLK(clk), .Q(\ram[3][164] ), .QN(
        n4359) );
  DFFX1_HVT \ram_reg[3][163]  ( .D(n992), .CLK(clk), .Q(\ram[3][163] ) );
  DFFX1_HVT \ram_reg[3][162]  ( .D(n991), .CLK(clk), .Q(\ram[3][162] ) );
  DFFX1_HVT \ram_reg[3][161]  ( .D(n990), .CLK(clk), .Q(\ram[3][161] ) );
  DFFX1_HVT \ram_reg[3][160]  ( .D(n989), .CLK(clk), .Q(\ram[3][160] ) );
  DFFX1_HVT \ram_reg[3][159]  ( .D(n988), .CLK(clk), .Q(\ram[3][159] ) );
  DFFX1_HVT \ram_reg[3][158]  ( .D(n987), .CLK(clk), .Q(\ram[3][158] ) );
  DFFX1_HVT \ram_reg[3][157]  ( .D(n986), .CLK(clk), .Q(\ram[3][157] ) );
  DFFX1_HVT \ram_reg[3][156]  ( .D(n985), .CLK(clk), .Q(\ram[3][156] ) );
  DFFX1_HVT \ram_reg[3][155]  ( .D(n984), .CLK(clk), .Q(\ram[3][155] ) );
  DFFX1_HVT \ram_reg[3][154]  ( .D(n983), .CLK(clk), .Q(\ram[3][154] ) );
  DFFX1_HVT \ram_reg[3][153]  ( .D(n982), .CLK(clk), .Q(\ram[3][153] ) );
  DFFX1_HVT \ram_reg[3][152]  ( .D(n981), .CLK(clk), .Q(\ram[3][152] ) );
  DFFX1_HVT \ram_reg[3][151]  ( .D(n980), .CLK(clk), .Q(\ram[3][151] ) );
  DFFX1_HVT \ram_reg[3][150]  ( .D(n979), .CLK(clk), .Q(\ram[3][150] ) );
  DFFX1_HVT \ram_reg[3][149]  ( .D(n978), .CLK(clk), .Q(\ram[3][149] ) );
  DFFX1_HVT \ram_reg[3][148]  ( .D(n977), .CLK(clk), .Q(\ram[3][148] ) );
  DFFX1_HVT \ram_reg[3][147]  ( .D(n976), .CLK(clk), .Q(\ram[3][147] ) );
  DFFX1_HVT \ram_reg[3][146]  ( .D(n975), .CLK(clk), .Q(\ram[3][146] ) );
  DFFX1_HVT \ram_reg[3][145]  ( .D(n974), .CLK(clk), .Q(\ram[3][145] ) );
  DFFX1_HVT \ram_reg[3][144]  ( .D(n973), .CLK(clk), .Q(\ram[3][144] ) );
  DFFX1_HVT \ram_reg[3][143]  ( .D(n972), .CLK(clk), .Q(\ram[3][143] ) );
  DFFX1_HVT \ram_reg[3][142]  ( .D(n971), .CLK(clk), .Q(\ram[3][142] ) );
  DFFX1_HVT \ram_reg[3][141]  ( .D(n970), .CLK(clk), .Q(\ram[3][141] ) );
  DFFX1_HVT \ram_reg[3][140]  ( .D(n969), .CLK(clk), .Q(\ram[3][140] ) );
  DFFX1_HVT \ram_reg[3][139]  ( .D(n968), .CLK(clk), .Q(\ram[3][139] ) );
  DFFX1_HVT \ram_reg[3][138]  ( .D(n967), .CLK(clk), .Q(\ram[3][138] ) );
  DFFX1_HVT \ram_reg[3][137]  ( .D(n966), .CLK(clk), .Q(\ram[3][137] ) );
  DFFX1_HVT \ram_reg[3][136]  ( .D(n965), .CLK(clk), .Q(\ram[3][136] ) );
  DFFX1_HVT \ram_reg[3][135]  ( .D(n964), .CLK(clk), .Q(\ram[3][135] ) );
  DFFX1_HVT \ram_reg[3][134]  ( .D(n963), .CLK(clk), .Q(\ram[3][134] ) );
  DFFX1_HVT \ram_reg[3][133]  ( .D(n962), .CLK(clk), .Q(\ram[3][133] ) );
  DFFX1_HVT \ram_reg[3][132]  ( .D(n961), .CLK(clk), .Q(\ram[3][132] ) );
  DFFX1_HVT \ram_reg[3][131]  ( .D(n960), .CLK(clk), .Q(\ram[3][131] ) );
  DFFX1_HVT \ram_reg[3][130]  ( .D(n959), .CLK(clk), .Q(\ram[3][130] ) );
  DFFX1_HVT \ram_reg[3][129]  ( .D(n958), .CLK(clk), .Q(\ram[3][129] ) );
  DFFX1_HVT \ram_reg[3][128]  ( .D(n957), .CLK(clk), .Q(\ram[3][128] ) );
  DFFX1_HVT \ram_reg[3][127]  ( .D(n956), .CLK(clk), .Q(\ram[3][127] ) );
  DFFX1_HVT \ram_reg[3][126]  ( .D(n955), .CLK(clk), .Q(\ram[3][126] ) );
  DFFX1_HVT \ram_reg[3][125]  ( .D(n954), .CLK(clk), .Q(\ram[3][125] ) );
  DFFX1_HVT \ram_reg[3][124]  ( .D(n953), .CLK(clk), .Q(\ram[3][124] ) );
  DFFX1_HVT \ram_reg[3][123]  ( .D(n952), .CLK(clk), .Q(\ram[3][123] ) );
  DFFX1_HVT \ram_reg[3][122]  ( .D(n951), .CLK(clk), .Q(\ram[3][122] ) );
  DFFX1_HVT \ram_reg[3][121]  ( .D(n950), .CLK(clk), .Q(\ram[3][121] ) );
  DFFX1_HVT \ram_reg[3][120]  ( .D(n949), .CLK(clk), .Q(\ram[3][120] ) );
  DFFX1_HVT \ram_reg[3][119]  ( .D(n948), .CLK(clk), .Q(\ram[3][119] ) );
  DFFX1_HVT \ram_reg[3][118]  ( .D(n947), .CLK(clk), .Q(\ram[3][118] ), .QN(
        n4524) );
  DFFX1_HVT \ram_reg[3][117]  ( .D(n946), .CLK(clk), .Q(\ram[3][117] ) );
  DFFX1_HVT \ram_reg[3][116]  ( .D(n945), .CLK(clk), .Q(\ram[3][116] ) );
  DFFX1_HVT \ram_reg[3][115]  ( .D(n944), .CLK(clk), .Q(\ram[3][115] ) );
  DFFX1_HVT \ram_reg[3][114]  ( .D(n943), .CLK(clk), .Q(\ram[3][114] ), .QN(
        n4563) );
  DFFX1_HVT \ram_reg[3][113]  ( .D(n942), .CLK(clk), .Q(\ram[3][113] ) );
  DFFX1_HVT \ram_reg[3][112]  ( .D(n941), .CLK(clk), .Q(\ram[3][112] ), .QN(
        n5838) );
  DFFX1_HVT \ram_reg[3][111]  ( .D(n940), .CLK(clk), .Q(\ram[3][111] ) );
  DFFX1_HVT \ram_reg[3][110]  ( .D(n939), .CLK(clk), .Q(\ram[3][110] ) );
  DFFX1_HVT \ram_reg[3][109]  ( .D(n938), .CLK(clk), .Q(\ram[3][109] ) );
  DFFX1_HVT \ram_reg[3][108]  ( .D(n937), .CLK(clk), .Q(\ram[3][108] ) );
  DFFX1_HVT \ram_reg[3][107]  ( .D(n936), .CLK(clk), .Q(\ram[3][107] ) );
  DFFX1_HVT \ram_reg[3][106]  ( .D(n935), .CLK(clk), .Q(\ram[3][106] ) );
  DFFX1_HVT \ram_reg[3][105]  ( .D(n934), .CLK(clk), .Q(\ram[3][105] ), .QN(
        n4367) );
  DFFX1_HVT \ram_reg[3][104]  ( .D(n933), .CLK(clk), .Q(\ram[3][104] ) );
  DFFX1_HVT \ram_reg[3][103]  ( .D(n932), .CLK(clk), .Q(\ram[3][103] ) );
  DFFX1_HVT \ram_reg[3][102]  ( .D(n931), .CLK(clk), .Q(\ram[3][102] ) );
  DFFX1_HVT \ram_reg[3][101]  ( .D(n930), .CLK(clk), .Q(\ram[3][101] ) );
  DFFX1_HVT \ram_reg[3][100]  ( .D(n929), .CLK(clk), .Q(\ram[3][100] ) );
  DFFX1_HVT \ram_reg[3][99]  ( .D(n928), .CLK(clk), .Q(\ram[3][99] ) );
  DFFX1_HVT \ram_reg[3][98]  ( .D(n927), .CLK(clk), .Q(\ram[3][98] ) );
  DFFX1_HVT \ram_reg[3][97]  ( .D(n926), .CLK(clk), .Q(\ram[3][97] ), .QN(
        n4500) );
  DFFX1_HVT \ram_reg[3][96]  ( .D(n925), .CLK(clk), .Q(\ram[3][96] ) );
  DFFX1_HVT \ram_reg[3][95]  ( .D(n924), .CLK(clk), .Q(\ram[3][95] ) );
  DFFX1_HVT \ram_reg[3][94]  ( .D(n923), .CLK(clk), .Q(\ram[3][94] ) );
  DFFX1_HVT \ram_reg[3][93]  ( .D(n922), .CLK(clk), .Q(\ram[3][93] ) );
  DFFX1_HVT \ram_reg[3][92]  ( .D(n921), .CLK(clk), .Q(\ram[3][92] ) );
  DFFX1_HVT \ram_reg[3][91]  ( .D(n920), .CLK(clk), .Q(\ram[3][91] ) );
  DFFX1_HVT \ram_reg[3][90]  ( .D(n919), .CLK(clk), .Q(\ram[3][90] ) );
  DFFX1_HVT \ram_reg[3][89]  ( .D(n918), .CLK(clk), .Q(\ram[3][89] ) );
  DFFX1_HVT \ram_reg[3][88]  ( .D(n5034), .CLK(clk), .Q(\ram[3][88] ), .QN(
        n5286) );
  DFFX1_HVT \ram_reg[3][87]  ( .D(n916), .CLK(clk), .Q(\ram[3][87] ), .QN(
        n4376) );
  DFFX1_HVT \ram_reg[3][86]  ( .D(n915), .CLK(clk), .Q(\ram[3][86] ) );
  DFFX1_HVT \ram_reg[3][85]  ( .D(n914), .CLK(clk), .Q(\ram[3][85] ) );
  DFFX1_HVT \ram_reg[3][84]  ( .D(n913), .CLK(clk), .Q(\ram[3][84] ), .QN(
        n4519) );
  DFFX1_HVT \ram_reg[3][83]  ( .D(n912), .CLK(clk), .Q(\ram[3][83] ) );
  DFFX1_HVT \ram_reg[3][82]  ( .D(n911), .CLK(clk), .Q(\ram[3][82] ) );
  DFFX1_HVT \ram_reg[3][81]  ( .D(n910), .CLK(clk), .Q(\ram[3][81] ) );
  DFFX1_HVT \ram_reg[3][80]  ( .D(n909), .CLK(clk), .Q(\ram[3][80] ) );
  DFFX1_HVT \ram_reg[3][79]  ( .D(n908), .CLK(clk), .Q(\ram[3][79] ) );
  DFFX1_HVT \ram_reg[3][78]  ( .D(n907), .CLK(clk), .Q(\ram[3][78] ) );
  DFFX1_HVT \ram_reg[3][77]  ( .D(n906), .CLK(clk), .Q(\ram[3][77] ) );
  DFFX1_HVT \ram_reg[3][76]  ( .D(n905), .CLK(clk), .Q(\ram[3][76] ) );
  DFFX1_HVT \ram_reg[3][75]  ( .D(n904), .CLK(clk), .Q(\ram[3][75] ) );
  DFFX1_HVT \ram_reg[3][74]  ( .D(n903), .CLK(clk), .Q(\ram[3][74] ) );
  DFFX1_HVT \ram_reg[3][73]  ( .D(n902), .CLK(clk), .Q(\ram[3][73] ) );
  DFFX1_HVT \ram_reg[3][72]  ( .D(n901), .CLK(clk), .Q(\ram[3][72] ) );
  DFFX1_HVT \ram_reg[3][71]  ( .D(n900), .CLK(clk), .Q(\ram[3][71] ) );
  DFFX1_HVT \ram_reg[3][70]  ( .D(n899), .CLK(clk), .Q(\ram[3][70] ) );
  DFFX1_HVT \ram_reg[3][69]  ( .D(n898), .CLK(clk), .Q(\ram[3][69] ) );
  DFFX1_HVT \ram_reg[3][68]  ( .D(n897), .CLK(clk), .Q(\ram[3][68] ) );
  DFFX1_HVT \ram_reg[3][67]  ( .D(n896), .CLK(clk), .Q(\ram[3][67] ) );
  DFFX1_HVT \ram_reg[3][66]  ( .D(n895), .CLK(clk), .Q(\ram[3][66] ) );
  DFFX1_HVT \ram_reg[3][65]  ( .D(n894), .CLK(clk), .Q(\ram[3][65] ) );
  DFFX1_HVT \ram_reg[3][64]  ( .D(n893), .CLK(clk), .Q(\ram[3][64] ) );
  DFFX1_HVT \ram_reg[3][63]  ( .D(n892), .CLK(clk), .Q(\ram[3][63] ) );
  DFFX1_HVT \ram_reg[3][62]  ( .D(n891), .CLK(clk), .Q(\ram[3][62] ) );
  DFFX1_HVT \ram_reg[3][61]  ( .D(n890), .CLK(clk), .Q(\ram[3][61] ) );
  DFFX1_HVT \ram_reg[3][60]  ( .D(n889), .CLK(clk), .Q(\ram[3][60] ) );
  DFFX1_HVT \ram_reg[3][59]  ( .D(n888), .CLK(clk), .Q(\ram[3][59] ) );
  DFFX1_HVT \ram_reg[3][58]  ( .D(n887), .CLK(clk), .Q(\ram[3][58] ) );
  DFFX1_HVT \ram_reg[3][57]  ( .D(n886), .CLK(clk), .Q(\ram[3][57] ) );
  DFFX1_HVT \ram_reg[3][56]  ( .D(n885), .CLK(clk), .Q(\ram[3][56] ) );
  DFFX1_HVT \ram_reg[3][55]  ( .D(n884), .CLK(clk), .Q(\ram[3][55] ) );
  DFFX1_HVT \ram_reg[3][54]  ( .D(n883), .CLK(clk), .Q(\ram[3][54] ) );
  DFFX1_HVT \ram_reg[3][53]  ( .D(n882), .CLK(clk), .Q(\ram[3][53] ) );
  DFFX1_HVT \ram_reg[3][52]  ( .D(n881), .CLK(clk), .Q(\ram[3][52] ) );
  DFFX1_HVT \ram_reg[3][51]  ( .D(n880), .CLK(clk), .Q(\ram[3][51] ) );
  DFFX1_HVT \ram_reg[3][50]  ( .D(n879), .CLK(clk), .Q(\ram[3][50] ) );
  DFFX1_HVT \ram_reg[3][49]  ( .D(n878), .CLK(clk), .Q(\ram[3][49] ) );
  DFFX1_HVT \ram_reg[3][48]  ( .D(n5466), .CLK(clk), .Q(\ram[3][48] ) );
  DFFX1_HVT \ram_reg[3][47]  ( .D(n876), .CLK(clk), .Q(\ram[3][47] ) );
  DFFX1_HVT \ram_reg[3][46]  ( .D(n875), .CLK(clk), .Q(\ram[3][46] ) );
  DFFX1_HVT \ram_reg[3][45]  ( .D(n874), .CLK(clk), .Q(\ram[3][45] ) );
  DFFX1_HVT \ram_reg[3][44]  ( .D(n873), .CLK(clk), .Q(\ram[3][44] ) );
  DFFX1_HVT \ram_reg[3][43]  ( .D(n872), .CLK(clk), .Q(\ram[3][43] ) );
  DFFX1_HVT \ram_reg[3][42]  ( .D(n871), .CLK(clk), .Q(\ram[3][42] ) );
  DFFX1_HVT \ram_reg[3][41]  ( .D(n870), .CLK(clk), .Q(\ram[3][41] ) );
  DFFX1_HVT \ram_reg[3][40]  ( .D(n869), .CLK(clk), .Q(\ram[3][40] ) );
  DFFX1_HVT \ram_reg[3][39]  ( .D(n868), .CLK(clk), .Q(\ram[3][39] ) );
  DFFX1_HVT \ram_reg[3][38]  ( .D(n867), .CLK(clk), .Q(\ram[3][38] ) );
  DFFX1_HVT \ram_reg[3][37]  ( .D(n5030), .CLK(clk), .Q(\ram[3][37] ), .QN(
        n5350) );
  DFFX1_HVT \ram_reg[3][36]  ( .D(n865), .CLK(clk), .Q(\ram[3][36] ) );
  DFFX1_HVT \ram_reg[3][35]  ( .D(n864), .CLK(clk), .Q(\ram[3][35] ) );
  DFFX1_HVT \ram_reg[3][34]  ( .D(n863), .CLK(clk), .Q(\ram[3][34] ) );
  DFFX1_HVT \ram_reg[3][33]  ( .D(n862), .CLK(clk), .Q(\ram[3][33] ) );
  DFFX1_HVT \ram_reg[3][32]  ( .D(n861), .CLK(clk), .Q(\ram[3][32] ) );
  DFFX1_HVT \ram_reg[3][31]  ( .D(n860), .CLK(clk), .Q(\ram[3][31] ) );
  DFFX1_HVT \ram_reg[3][30]  ( .D(n859), .CLK(clk), .Q(\ram[3][30] ) );
  DFFX1_HVT \ram_reg[3][29]  ( .D(n858), .CLK(clk), .Q(\ram[3][29] ) );
  DFFX1_HVT \ram_reg[3][28]  ( .D(n857), .CLK(clk), .Q(\ram[3][28] ) );
  DFFX1_HVT \ram_reg[3][27]  ( .D(n856), .CLK(clk), .Q(\ram[3][27] ) );
  DFFX1_HVT \ram_reg[3][26]  ( .D(n855), .CLK(clk), .Q(\ram[3][26] ), .QN(
        n4522) );
  DFFX1_HVT \ram_reg[3][25]  ( .D(n854), .CLK(clk), .Q(\ram[3][25] ) );
  DFFX1_HVT \ram_reg[3][24]  ( .D(n853), .CLK(clk), .Q(\ram[3][24] ) );
  DFFX1_HVT \ram_reg[3][23]  ( .D(n852), .CLK(clk), .Q(\ram[3][23] ) );
  DFFX1_HVT \ram_reg[3][22]  ( .D(n851), .CLK(clk), .Q(\ram[3][22] ) );
  DFFX1_HVT \ram_reg[3][21]  ( .D(n850), .CLK(clk), .Q(\ram[3][21] ) );
  DFFX1_HVT \ram_reg[3][20]  ( .D(n849), .CLK(clk), .Q(\ram[3][20] ) );
  DFFX1_HVT \ram_reg[3][19]  ( .D(n848), .CLK(clk), .Q(\ram[3][19] ) );
  DFFX1_HVT \ram_reg[3][18]  ( .D(n847), .CLK(clk), .Q(\ram[3][18] ), .QN(
        n4244) );
  DFFX1_HVT \ram_reg[3][17]  ( .D(n846), .CLK(clk), .Q(\ram[3][17] ), .QN(
        n4247) );
  DFFX1_HVT \ram_reg[3][16]  ( .D(n845), .CLK(clk), .Q(\ram[3][16] ), .QN(
        n4373) );
  DFFX1_HVT \ram_reg[3][15]  ( .D(n844), .CLK(clk), .Q(\ram[3][15] ) );
  DFFX1_HVT \ram_reg[3][14]  ( .D(n843), .CLK(clk), .Q(\ram[3][14] ) );
  DFFX1_HVT \ram_reg[3][13]  ( .D(n842), .CLK(clk), .Q(\ram[3][13] ) );
  DFFX1_HVT \ram_reg[3][12]  ( .D(n841), .CLK(clk), .Q(\ram[3][12] ) );
  DFFX1_HVT \ram_reg[3][11]  ( .D(n840), .CLK(clk), .Q(\ram[3][11] ) );
  DFFX1_HVT \ram_reg[3][10]  ( .D(n839), .CLK(clk), .Q(\ram[3][10] ) );
  DFFX1_HVT \ram_reg[3][9]  ( .D(n838), .CLK(clk), .Q(\ram[3][9] ) );
  DFFX1_HVT \ram_reg[3][8]  ( .D(n837), .CLK(clk), .Q(\ram[3][8] ), .QN(n4250)
         );
  DFFX1_HVT \ram_reg[3][7]  ( .D(n836), .CLK(clk), .Q(\ram[3][7] ), .QN(n6402)
         );
  DFFX1_HVT \ram_reg[3][6]  ( .D(n835), .CLK(clk), .Q(\ram[3][6] ) );
  DFFX1_HVT \ram_reg[3][5]  ( .D(n834), .CLK(clk), .Q(\ram[3][5] ) );
  DFFX1_HVT \ram_reg[3][4]  ( .D(n5031), .CLK(clk), .Q(\ram[3][4] ), .QN(n6256) );
  DFFX1_HVT \ram_reg[3][3]  ( .D(n832), .CLK(clk), .Q(\ram[3][3] ), .QN(n4252)
         );
  DFFX1_HVT \ram_reg[3][2]  ( .D(n831), .CLK(clk), .Q(\ram[3][2] ), .QN(n4473)
         );
  DFFX1_HVT \ram_reg[3][1]  ( .D(n830), .CLK(clk), .Q(\ram[3][1] ) );
  DFFX1_HVT \ram_reg[3][0]  ( .D(n5032), .CLK(clk), .Q(\ram[3][0] ), .QN(n5375) );
  DFFX1_HVT \ram_reg[2][255]  ( .D(n828), .CLK(clk), .Q(\ram[2][255] ) );
  DFFX1_HVT \ram_reg[2][254]  ( .D(n827), .CLK(clk), .Q(\ram[2][254] ) );
  DFFX1_HVT \ram_reg[2][253]  ( .D(n826), .CLK(clk), .Q(\ram[2][253] ) );
  DFFX1_HVT \ram_reg[2][252]  ( .D(n825), .CLK(clk), .Q(\ram[2][252] ), .QN(
        n5443) );
  DFFX1_HVT \ram_reg[2][251]  ( .D(n824), .CLK(clk), .Q(\ram[2][251] ) );
  DFFX1_HVT \ram_reg[2][250]  ( .D(n823), .CLK(clk), .Q(\ram[2][250] ) );
  DFFX1_HVT \ram_reg[2][249]  ( .D(n822), .CLK(clk), .Q(\ram[2][249] ) );
  DFFX1_HVT \ram_reg[2][248]  ( .D(n821), .CLK(clk), .Q(\ram[2][248] ) );
  DFFX1_HVT \ram_reg[2][247]  ( .D(n820), .CLK(clk), .Q(\ram[2][247] ) );
  DFFX1_HVT \ram_reg[2][246]  ( .D(n819), .CLK(clk), .Q(\ram[2][246] ) );
  DFFX1_HVT \ram_reg[2][245]  ( .D(n818), .CLK(clk), .Q(\ram[2][245] ) );
  DFFX1_HVT \ram_reg[2][244]  ( .D(n817), .CLK(clk), .Q(\ram[2][244] ) );
  DFFX1_HVT \ram_reg[2][243]  ( .D(n816), .CLK(clk), .Q(\ram[2][243] ) );
  DFFX1_HVT \ram_reg[2][242]  ( .D(n815), .CLK(clk), .Q(\ram[2][242] ) );
  DFFX1_HVT \ram_reg[2][241]  ( .D(n814), .CLK(clk), .Q(\ram[2][241] ) );
  DFFX1_HVT \ram_reg[2][240]  ( .D(n813), .CLK(clk), .Q(\ram[2][240] ) );
  DFFX1_HVT \ram_reg[2][239]  ( .D(n812), .CLK(clk), .Q(\ram[2][239] ) );
  DFFX1_HVT \ram_reg[2][238]  ( .D(n811), .CLK(clk), .Q(\ram[2][238] ) );
  DFFX1_HVT \ram_reg[2][237]  ( .D(n810), .CLK(clk), .Q(\ram[2][237] ) );
  DFFX1_HVT \ram_reg[2][236]  ( .D(n809), .CLK(clk), .Q(\ram[2][236] ) );
  DFFX1_HVT \ram_reg[2][235]  ( .D(n808), .CLK(clk), .Q(\ram[2][235] ) );
  DFFX1_HVT \ram_reg[2][234]  ( .D(n807), .CLK(clk), .Q(\ram[2][234] ) );
  DFFX1_HVT \ram_reg[2][233]  ( .D(n806), .CLK(clk), .Q(\ram[2][233] ) );
  DFFX1_HVT \ram_reg[2][232]  ( .D(n805), .CLK(clk), .Q(\ram[2][232] ) );
  DFFX1_HVT \ram_reg[2][231]  ( .D(n804), .CLK(clk), .Q(\ram[2][231] ) );
  DFFX1_HVT \ram_reg[2][230]  ( .D(n803), .CLK(clk), .Q(\ram[2][230] ) );
  DFFX1_HVT \ram_reg[2][229]  ( .D(n802), .CLK(clk), .Q(\ram[2][229] ) );
  DFFX1_HVT \ram_reg[2][228]  ( .D(n801), .CLK(clk), .Q(\ram[2][228] ) );
  DFFX1_HVT \ram_reg[2][227]  ( .D(n800), .CLK(clk), .Q(\ram[2][227] ) );
  DFFX1_HVT \ram_reg[2][226]  ( .D(n799), .CLK(clk), .Q(\ram[2][226] ) );
  DFFX1_HVT \ram_reg[2][225]  ( .D(n798), .CLK(clk), .Q(\ram[2][225] ) );
  DFFX1_HVT \ram_reg[2][224]  ( .D(n797), .CLK(clk), .Q(\ram[2][224] ), .QN(
        n5169) );
  DFFX1_HVT \ram_reg[2][223]  ( .D(n796), .CLK(clk), .Q(\ram[2][223] ) );
  DFFX1_HVT \ram_reg[2][222]  ( .D(n795), .CLK(clk), .Q(\ram[2][222] ) );
  DFFX1_HVT \ram_reg[2][221]  ( .D(n794), .CLK(clk), .Q(\ram[2][221] ) );
  DFFX1_HVT \ram_reg[2][220]  ( .D(n793), .CLK(clk), .Q(\ram[2][220] ) );
  DFFX1_HVT \ram_reg[2][219]  ( .D(n792), .CLK(clk), .Q(\ram[2][219] ) );
  DFFX1_HVT \ram_reg[2][218]  ( .D(n791), .CLK(clk), .Q(\ram[2][218] ) );
  DFFX1_HVT \ram_reg[2][217]  ( .D(n790), .CLK(clk), .Q(\ram[2][217] ) );
  DFFX1_HVT \ram_reg[2][216]  ( .D(n789), .CLK(clk), .Q(\ram[2][216] ) );
  DFFX1_HVT \ram_reg[2][215]  ( .D(n788), .CLK(clk), .Q(\ram[2][215] ) );
  DFFX1_HVT \ram_reg[2][214]  ( .D(n787), .CLK(clk), .Q(\ram[2][214] ) );
  DFFX1_HVT \ram_reg[2][213]  ( .D(n786), .CLK(clk), .Q(\ram[2][213] ) );
  DFFX1_HVT \ram_reg[2][212]  ( .D(n785), .CLK(clk), .Q(\ram[2][212] ) );
  DFFX1_HVT \ram_reg[2][211]  ( .D(n784), .CLK(clk), .Q(\ram[2][211] ) );
  DFFX1_HVT \ram_reg[2][210]  ( .D(n783), .CLK(clk), .Q(\ram[2][210] ) );
  DFFX1_HVT \ram_reg[2][209]  ( .D(n782), .CLK(clk), .Q(\ram[2][209] ) );
  DFFX1_HVT \ram_reg[2][208]  ( .D(n781), .CLK(clk), .Q(\ram[2][208] ) );
  DFFX1_HVT \ram_reg[2][207]  ( .D(n780), .CLK(clk), .Q(\ram[2][207] ) );
  DFFX1_HVT \ram_reg[2][206]  ( .D(n779), .CLK(clk), .Q(\ram[2][206] ) );
  DFFX1_HVT \ram_reg[2][205]  ( .D(n778), .CLK(clk), .Q(\ram[2][205] ) );
  DFFX1_HVT \ram_reg[2][204]  ( .D(n777), .CLK(clk), .Q(\ram[2][204] ) );
  DFFX1_HVT \ram_reg[2][203]  ( .D(n776), .CLK(clk), .Q(\ram[2][203] ) );
  DFFX1_HVT \ram_reg[2][202]  ( .D(n775), .CLK(clk), .Q(\ram[2][202] ) );
  DFFX1_HVT \ram_reg[2][201]  ( .D(n774), .CLK(clk), .Q(\ram[2][201] ) );
  DFFX1_HVT \ram_reg[2][200]  ( .D(n773), .CLK(clk), .Q(\ram[2][200] ) );
  DFFX1_HVT \ram_reg[2][199]  ( .D(n772), .CLK(clk), .Q(\ram[2][199] ) );
  DFFX1_HVT \ram_reg[2][198]  ( .D(n771), .CLK(clk), .Q(\ram[2][198] ) );
  DFFX1_HVT \ram_reg[2][197]  ( .D(n770), .CLK(clk), .Q(\ram[2][197] ) );
  DFFX1_HVT \ram_reg[2][196]  ( .D(n769), .CLK(clk), .Q(\ram[2][196] ) );
  DFFX1_HVT \ram_reg[2][195]  ( .D(n768), .CLK(clk), .Q(\ram[2][195] ) );
  DFFX1_HVT \ram_reg[2][194]  ( .D(n767), .CLK(clk), .Q(\ram[2][194] ) );
  DFFX1_HVT \ram_reg[2][193]  ( .D(n766), .CLK(clk), .Q(\ram[2][193] ) );
  DFFX1_HVT \ram_reg[2][192]  ( .D(n765), .CLK(clk), .Q(\ram[2][192] ) );
  DFFX1_HVT \ram_reg[2][191]  ( .D(n764), .CLK(clk), .Q(\ram[2][191] ) );
  DFFX1_HVT \ram_reg[2][190]  ( .D(n763), .CLK(clk), .Q(\ram[2][190] ) );
  DFFX1_HVT \ram_reg[2][189]  ( .D(n762), .CLK(clk), .Q(\ram[2][189] ) );
  DFFX1_HVT \ram_reg[2][188]  ( .D(n761), .CLK(clk), .Q(\ram[2][188] ) );
  DFFX1_HVT \ram_reg[2][187]  ( .D(n760), .CLK(clk), .Q(\ram[2][187] ) );
  DFFX1_HVT \ram_reg[2][186]  ( .D(n759), .CLK(clk), .Q(\ram[2][186] ) );
  DFFX1_HVT \ram_reg[2][185]  ( .D(n758), .CLK(clk), .Q(\ram[2][185] ) );
  DFFX1_HVT \ram_reg[2][184]  ( .D(n757), .CLK(clk), .Q(\ram[2][184] ) );
  DFFX1_HVT \ram_reg[2][183]  ( .D(n756), .CLK(clk), .Q(\ram[2][183] ) );
  DFFX1_HVT \ram_reg[2][182]  ( .D(n755), .CLK(clk), .Q(\ram[2][182] ) );
  DFFX1_HVT \ram_reg[2][181]  ( .D(n754), .CLK(clk), .Q(\ram[2][181] ) );
  DFFX1_HVT \ram_reg[2][180]  ( .D(n753), .CLK(clk), .Q(\ram[2][180] ) );
  DFFX1_HVT \ram_reg[2][179]  ( .D(n752), .CLK(clk), .Q(\ram[2][179] ) );
  DFFX1_HVT \ram_reg[2][178]  ( .D(n751), .CLK(clk), .Q(\ram[2][178] ) );
  DFFX1_HVT \ram_reg[2][177]  ( .D(n750), .CLK(clk), .Q(\ram[2][177] ) );
  DFFX1_HVT \ram_reg[2][176]  ( .D(n749), .CLK(clk), .Q(\ram[2][176] ) );
  DFFX1_HVT \ram_reg[2][175]  ( .D(n748), .CLK(clk), .Q(\ram[2][175] ) );
  DFFX1_HVT \ram_reg[2][174]  ( .D(n747), .CLK(clk), .Q(\ram[2][174] ) );
  DFFX1_HVT \ram_reg[2][173]  ( .D(n746), .CLK(clk), .Q(\ram[2][173] ) );
  DFFX1_HVT \ram_reg[2][172]  ( .D(n745), .CLK(clk), .Q(\ram[2][172] ) );
  DFFX1_HVT \ram_reg[2][171]  ( .D(n744), .CLK(clk), .Q(\ram[2][171] ) );
  DFFX1_HVT \ram_reg[2][170]  ( .D(n743), .CLK(clk), .Q(\ram[2][170] ) );
  DFFX1_HVT \ram_reg[2][169]  ( .D(n742), .CLK(clk), .Q(\ram[2][169] ) );
  DFFX1_HVT \ram_reg[2][168]  ( .D(n741), .CLK(clk), .Q(\ram[2][168] ) );
  DFFX1_HVT \ram_reg[2][167]  ( .D(n740), .CLK(clk), .Q(\ram[2][167] ) );
  DFFX1_HVT \ram_reg[2][166]  ( .D(n739), .CLK(clk), .Q(\ram[2][166] ) );
  DFFX1_HVT \ram_reg[2][165]  ( .D(n738), .CLK(clk), .Q(\ram[2][165] ) );
  DFFX1_HVT \ram_reg[2][164]  ( .D(n737), .CLK(clk), .Q(\ram[2][164] ) );
  DFFX1_HVT \ram_reg[2][163]  ( .D(n736), .CLK(clk), .Q(\ram[2][163] ) );
  DFFX1_HVT \ram_reg[2][162]  ( .D(n735), .CLK(clk), .Q(\ram[2][162] ) );
  DFFX1_HVT \ram_reg[2][161]  ( .D(n734), .CLK(clk), .Q(\ram[2][161] ) );
  DFFX1_HVT \ram_reg[2][160]  ( .D(n733), .CLK(clk), .Q(\ram[2][160] ) );
  DFFX1_HVT \ram_reg[2][159]  ( .D(n732), .CLK(clk), .Q(\ram[2][159] ) );
  DFFX1_HVT \ram_reg[2][158]  ( .D(n731), .CLK(clk), .Q(\ram[2][158] ) );
  DFFX1_HVT \ram_reg[2][157]  ( .D(n730), .CLK(clk), .Q(\ram[2][157] ) );
  DFFX1_HVT \ram_reg[2][156]  ( .D(n729), .CLK(clk), .Q(\ram[2][156] ) );
  DFFX1_HVT \ram_reg[2][155]  ( .D(n728), .CLK(clk), .Q(\ram[2][155] ) );
  DFFX1_HVT \ram_reg[2][154]  ( .D(n727), .CLK(clk), .Q(\ram[2][154] ) );
  DFFX1_HVT \ram_reg[2][153]  ( .D(n726), .CLK(clk), .Q(\ram[2][153] ) );
  DFFX1_HVT \ram_reg[2][152]  ( .D(n725), .CLK(clk), .Q(\ram[2][152] ) );
  DFFX1_HVT \ram_reg[2][151]  ( .D(n724), .CLK(clk), .Q(\ram[2][151] ) );
  DFFX1_HVT \ram_reg[2][150]  ( .D(n723), .CLK(clk), .Q(\ram[2][150] ) );
  DFFX1_HVT \ram_reg[2][149]  ( .D(n722), .CLK(clk), .Q(\ram[2][149] ) );
  DFFX1_HVT \ram_reg[2][148]  ( .D(n721), .CLK(clk), .Q(\ram[2][148] ) );
  DFFX1_HVT \ram_reg[2][147]  ( .D(n720), .CLK(clk), .Q(\ram[2][147] ), .QN(
        n917) );
  DFFX1_HVT \ram_reg[2][146]  ( .D(n719), .CLK(clk), .Q(\ram[2][146] ) );
  DFFX1_HVT \ram_reg[2][145]  ( .D(n718), .CLK(clk), .Q(\ram[2][145] ) );
  DFFX1_HVT \ram_reg[2][144]  ( .D(n717), .CLK(clk), .Q(\ram[2][144] ) );
  DFFX1_HVT \ram_reg[2][143]  ( .D(n716), .CLK(clk), .Q(\ram[2][143] ) );
  DFFX1_HVT \ram_reg[2][142]  ( .D(n715), .CLK(clk), .Q(\ram[2][142] ) );
  DFFX1_HVT \ram_reg[2][141]  ( .D(n714), .CLK(clk), .Q(\ram[2][141] ) );
  DFFX1_HVT \ram_reg[2][140]  ( .D(n713), .CLK(clk), .Q(\ram[2][140] ) );
  DFFX1_HVT \ram_reg[2][139]  ( .D(n712), .CLK(clk), .Q(\ram[2][139] ) );
  DFFX1_HVT \ram_reg[2][138]  ( .D(n711), .CLK(clk), .Q(\ram[2][138] ) );
  DFFX1_HVT \ram_reg[2][137]  ( .D(n710), .CLK(clk), .Q(\ram[2][137] ) );
  DFFX1_HVT \ram_reg[2][136]  ( .D(n709), .CLK(clk), .Q(\ram[2][136] ) );
  DFFX1_HVT \ram_reg[2][135]  ( .D(n708), .CLK(clk), .Q(\ram[2][135] ) );
  DFFX1_HVT \ram_reg[2][134]  ( .D(n707), .CLK(clk), .Q(\ram[2][134] ) );
  DFFX1_HVT \ram_reg[2][133]  ( .D(n706), .CLK(clk), .Q(\ram[2][133] ) );
  DFFX1_HVT \ram_reg[2][132]  ( .D(n705), .CLK(clk), .Q(\ram[2][132] ) );
  DFFX1_HVT \ram_reg[2][131]  ( .D(n704), .CLK(clk), .Q(\ram[2][131] ) );
  DFFX1_HVT \ram_reg[2][130]  ( .D(n703), .CLK(clk), .Q(\ram[2][130] ) );
  DFFX1_HVT \ram_reg[2][129]  ( .D(n702), .CLK(clk), .Q(\ram[2][129] ) );
  DFFX1_HVT \ram_reg[2][128]  ( .D(n701), .CLK(clk), .Q(\ram[2][128] ) );
  DFFX1_HVT \ram_reg[2][127]  ( .D(n700), .CLK(clk), .Q(\ram[2][127] ) );
  DFFX1_HVT \ram_reg[2][126]  ( .D(n699), .CLK(clk), .Q(\ram[2][126] ) );
  DFFX1_HVT \ram_reg[2][125]  ( .D(n698), .CLK(clk), .Q(\ram[2][125] ) );
  DFFX1_HVT \ram_reg[2][124]  ( .D(n697), .CLK(clk), .Q(\ram[2][124] ) );
  DFFX1_HVT \ram_reg[2][123]  ( .D(n696), .CLK(clk), .Q(\ram[2][123] ) );
  DFFX1_HVT \ram_reg[2][122]  ( .D(n695), .CLK(clk), .Q(\ram[2][122] ) );
  DFFX1_HVT \ram_reg[2][121]  ( .D(n694), .CLK(clk), .Q(\ram[2][121] ) );
  DFFX1_HVT \ram_reg[2][120]  ( .D(n693), .CLK(clk), .Q(\ram[2][120] ) );
  DFFX1_HVT \ram_reg[2][119]  ( .D(n692), .CLK(clk), .Q(\ram[2][119] ) );
  DFFX1_HVT \ram_reg[2][118]  ( .D(n691), .CLK(clk), .Q(\ram[2][118] ) );
  DFFX1_HVT \ram_reg[2][117]  ( .D(n690), .CLK(clk), .Q(\ram[2][117] ) );
  DFFX1_HVT \ram_reg[2][116]  ( .D(n689), .CLK(clk), .Q(\ram[2][116] ) );
  DFFX1_HVT \ram_reg[2][115]  ( .D(n688), .CLK(clk), .Q(\ram[2][115] ) );
  DFFX1_HVT \ram_reg[2][114]  ( .D(n687), .CLK(clk), .Q(\ram[2][114] ) );
  DFFX1_HVT \ram_reg[2][113]  ( .D(n686), .CLK(clk), .Q(\ram[2][113] ) );
  DFFX1_HVT \ram_reg[2][112]  ( .D(n685), .CLK(clk), .Q(\ram[2][112] ), .QN(
        n5839) );
  DFFX1_HVT \ram_reg[2][111]  ( .D(n684), .CLK(clk), .Q(\ram[2][111] ) );
  DFFX1_HVT \ram_reg[2][110]  ( .D(n683), .CLK(clk), .Q(\ram[2][110] ) );
  DFFX1_HVT \ram_reg[2][109]  ( .D(n682), .CLK(clk), .Q(\ram[2][109] ) );
  DFFX1_HVT \ram_reg[2][108]  ( .D(n681), .CLK(clk), .Q(\ram[2][108] ) );
  DFFX1_HVT \ram_reg[2][107]  ( .D(n680), .CLK(clk), .Q(\ram[2][107] ) );
  DFFX1_HVT \ram_reg[2][106]  ( .D(n679), .CLK(clk), .Q(\ram[2][106] ) );
  DFFX1_HVT \ram_reg[2][105]  ( .D(n678), .CLK(clk), .Q(\ram[2][105] ) );
  DFFX1_HVT \ram_reg[2][104]  ( .D(n677), .CLK(clk), .Q(\ram[2][104] ) );
  DFFX1_HVT \ram_reg[2][103]  ( .D(n676), .CLK(clk), .Q(\ram[2][103] ) );
  DFFX1_HVT \ram_reg[2][102]  ( .D(n675), .CLK(clk), .Q(\ram[2][102] ) );
  DFFX1_HVT \ram_reg[2][101]  ( .D(n674), .CLK(clk), .Q(\ram[2][101] ) );
  DFFX1_HVT \ram_reg[2][100]  ( .D(n673), .CLK(clk), .Q(\ram[2][100] ) );
  DFFX1_HVT \ram_reg[2][99]  ( .D(n672), .CLK(clk), .Q(\ram[2][99] ) );
  DFFX1_HVT \ram_reg[2][98]  ( .D(n671), .CLK(clk), .Q(\ram[2][98] ) );
  DFFX1_HVT \ram_reg[2][97]  ( .D(n670), .CLK(clk), .Q(\ram[2][97] ) );
  DFFX1_HVT \ram_reg[2][96]  ( .D(n669), .CLK(clk), .Q(\ram[2][96] ) );
  DFFX1_HVT \ram_reg[2][95]  ( .D(n668), .CLK(clk), .Q(\ram[2][95] ) );
  DFFX1_HVT \ram_reg[2][94]  ( .D(n667), .CLK(clk), .Q(\ram[2][94] ) );
  DFFX1_HVT \ram_reg[2][93]  ( .D(n666), .CLK(clk), .Q(\ram[2][93] ) );
  DFFX1_HVT \ram_reg[2][92]  ( .D(n665), .CLK(clk), .Q(\ram[2][92] ) );
  DFFX1_HVT \ram_reg[2][91]  ( .D(n664), .CLK(clk), .Q(\ram[2][91] ) );
  DFFX1_HVT \ram_reg[2][90]  ( .D(n663), .CLK(clk), .Q(\ram[2][90] ) );
  DFFX1_HVT \ram_reg[2][89]  ( .D(n662), .CLK(clk), .Q(\ram[2][89] ) );
  DFFX1_HVT \ram_reg[2][88]  ( .D(n661), .CLK(clk), .Q(\ram[2][88] ) );
  DFFX1_HVT \ram_reg[2][87]  ( .D(n660), .CLK(clk), .Q(\ram[2][87] ) );
  DFFX1_HVT \ram_reg[2][86]  ( .D(n659), .CLK(clk), .Q(\ram[2][86] ) );
  DFFX1_HVT \ram_reg[2][85]  ( .D(n658), .CLK(clk), .Q(\ram[2][85] ) );
  DFFX1_HVT \ram_reg[2][84]  ( .D(n657), .CLK(clk), .Q(\ram[2][84] ) );
  DFFX1_HVT \ram_reg[2][83]  ( .D(n656), .CLK(clk), .Q(\ram[2][83] ) );
  DFFX1_HVT \ram_reg[2][82]  ( .D(n655), .CLK(clk), .Q(\ram[2][82] ) );
  DFFX1_HVT \ram_reg[2][81]  ( .D(n654), .CLK(clk), .Q(\ram[2][81] ) );
  DFFX1_HVT \ram_reg[2][80]  ( .D(n653), .CLK(clk), .Q(\ram[2][80] ) );
  DFFX1_HVT \ram_reg[2][79]  ( .D(n652), .CLK(clk), .Q(\ram[2][79] ) );
  DFFX1_HVT \ram_reg[2][78]  ( .D(n651), .CLK(clk), .Q(\ram[2][78] ) );
  DFFX1_HVT \ram_reg[2][77]  ( .D(n650), .CLK(clk), .Q(\ram[2][77] ) );
  DFFX1_HVT \ram_reg[2][76]  ( .D(n649), .CLK(clk), .Q(\ram[2][76] ) );
  DFFX1_HVT \ram_reg[2][75]  ( .D(n648), .CLK(clk), .Q(\ram[2][75] ) );
  DFFX1_HVT \ram_reg[2][74]  ( .D(n647), .CLK(clk), .Q(\ram[2][74] ) );
  DFFX1_HVT \ram_reg[2][73]  ( .D(n646), .CLK(clk), .Q(\ram[2][73] ) );
  DFFX1_HVT \ram_reg[2][72]  ( .D(n645), .CLK(clk), .Q(\ram[2][72] ), .QN(
        n5468) );
  DFFX1_HVT \ram_reg[2][71]  ( .D(n644), .CLK(clk), .Q(\ram[2][71] ) );
  DFFX1_HVT \ram_reg[2][70]  ( .D(n643), .CLK(clk), .Q(\ram[2][70] ) );
  DFFX1_HVT \ram_reg[2][69]  ( .D(n642), .CLK(clk), .Q(\ram[2][69] ) );
  DFFX1_HVT \ram_reg[2][68]  ( .D(n641), .CLK(clk), .Q(\ram[2][68] ) );
  DFFX1_HVT \ram_reg[2][67]  ( .D(n640), .CLK(clk), .Q(\ram[2][67] ), .QN(
        n4636) );
  DFFX1_HVT \ram_reg[2][66]  ( .D(n639), .CLK(clk), .Q(\ram[2][66] ) );
  DFFX1_HVT \ram_reg[2][65]  ( .D(n638), .CLK(clk), .Q(\ram[2][65] ) );
  DFFX1_HVT \ram_reg[2][64]  ( .D(n637), .CLK(clk), .Q(\ram[2][64] ) );
  DFFX1_HVT \ram_reg[2][63]  ( .D(n636), .CLK(clk), .Q(\ram[2][63] ) );
  DFFX1_HVT \ram_reg[2][62]  ( .D(n635), .CLK(clk), .Q(\ram[2][62] ) );
  DFFX1_HVT \ram_reg[2][61]  ( .D(n634), .CLK(clk), .Q(\ram[2][61] ) );
  DFFX1_HVT \ram_reg[2][60]  ( .D(n633), .CLK(clk), .Q(\ram[2][60] ) );
  DFFX1_HVT \ram_reg[2][59]  ( .D(n632), .CLK(clk), .Q(\ram[2][59] ) );
  DFFX1_HVT \ram_reg[2][58]  ( .D(n631), .CLK(clk), .Q(\ram[2][58] ) );
  DFFX1_HVT \ram_reg[2][57]  ( .D(n630), .CLK(clk), .Q(\ram[2][57] ) );
  DFFX1_HVT \ram_reg[2][56]  ( .D(n629), .CLK(clk), .Q(\ram[2][56] ) );
  DFFX1_HVT \ram_reg[2][55]  ( .D(n628), .CLK(clk), .Q(\ram[2][55] ) );
  DFFX1_HVT \ram_reg[2][54]  ( .D(n627), .CLK(clk), .Q(\ram[2][54] ) );
  DFFX1_HVT \ram_reg[2][53]  ( .D(n626), .CLK(clk), .Q(\ram[2][53] ) );
  DFFX1_HVT \ram_reg[2][52]  ( .D(n625), .CLK(clk), .Q(\ram[2][52] ) );
  DFFX1_HVT \ram_reg[2][51]  ( .D(n624), .CLK(clk), .Q(\ram[2][51] ) );
  DFFX1_HVT \ram_reg[2][50]  ( .D(n623), .CLK(clk), .Q(\ram[2][50] ) );
  DFFX1_HVT \ram_reg[2][49]  ( .D(n622), .CLK(clk), .Q(\ram[2][49] ) );
  DFFX1_HVT \ram_reg[2][48]  ( .D(n621), .CLK(clk), .Q(\ram[2][48] ) );
  DFFX1_HVT \ram_reg[2][47]  ( .D(n620), .CLK(clk), .Q(\ram[2][47] ) );
  DFFX1_HVT \ram_reg[2][46]  ( .D(n619), .CLK(clk), .Q(\ram[2][46] ) );
  DFFX1_HVT \ram_reg[2][45]  ( .D(n618), .CLK(clk), .Q(\ram[2][45] ) );
  DFFX1_HVT \ram_reg[2][44]  ( .D(n617), .CLK(clk), .Q(\ram[2][44] ) );
  DFFX1_HVT \ram_reg[2][43]  ( .D(n616), .CLK(clk), .Q(\ram[2][43] ) );
  DFFX1_HVT \ram_reg[2][42]  ( .D(n615), .CLK(clk), .Q(\ram[2][42] ) );
  DFFX1_HVT \ram_reg[2][41]  ( .D(n614), .CLK(clk), .Q(\ram[2][41] ) );
  DFFX1_HVT \ram_reg[2][40]  ( .D(n613), .CLK(clk), .Q(\ram[2][40] ) );
  DFFX1_HVT \ram_reg[2][39]  ( .D(n612), .CLK(clk), .Q(\ram[2][39] ) );
  DFFX1_HVT \ram_reg[2][38]  ( .D(n611), .CLK(clk), .Q(\ram[2][38] ) );
  DFFX1_HVT \ram_reg[2][37]  ( .D(n610), .CLK(clk), .Q(\ram[2][37] ) );
  DFFX1_HVT \ram_reg[2][36]  ( .D(n609), .CLK(clk), .Q(\ram[2][36] ) );
  DFFX1_HVT \ram_reg[2][35]  ( .D(n608), .CLK(clk), .Q(\ram[2][35] ) );
  DFFX1_HVT \ram_reg[2][34]  ( .D(n607), .CLK(clk), .Q(\ram[2][34] ) );
  DFFX1_HVT \ram_reg[2][33]  ( .D(n606), .CLK(clk), .Q(\ram[2][33] ) );
  DFFX1_HVT \ram_reg[2][32]  ( .D(n605), .CLK(clk), .Q(\ram[2][32] ) );
  DFFX1_HVT \ram_reg[2][31]  ( .D(n604), .CLK(clk), .Q(\ram[2][31] ) );
  DFFX1_HVT \ram_reg[2][30]  ( .D(n603), .CLK(clk), .Q(\ram[2][30] ) );
  DFFX1_HVT \ram_reg[2][29]  ( .D(n602), .CLK(clk), .Q(\ram[2][29] ) );
  DFFX1_HVT \ram_reg[2][28]  ( .D(n601), .CLK(clk), .Q(\ram[2][28] ) );
  DFFX1_HVT \ram_reg[2][27]  ( .D(n600), .CLK(clk), .Q(\ram[2][27] ) );
  DFFX1_HVT \ram_reg[2][26]  ( .D(n599), .CLK(clk), .Q(\ram[2][26] ) );
  DFFX1_HVT \ram_reg[2][25]  ( .D(n598), .CLK(clk), .Q(\ram[2][25] ) );
  DFFX1_HVT \ram_reg[2][24]  ( .D(n597), .CLK(clk), .Q(\ram[2][24] ) );
  DFFX1_HVT \ram_reg[2][23]  ( .D(n596), .CLK(clk), .Q(\ram[2][23] ) );
  DFFX1_HVT \ram_reg[2][22]  ( .D(n595), .CLK(clk), .Q(\ram[2][22] ) );
  DFFX1_HVT \ram_reg[2][21]  ( .D(n594), .CLK(clk), .Q(\ram[2][21] ) );
  DFFX1_HVT \ram_reg[2][20]  ( .D(n593), .CLK(clk), .Q(\ram[2][20] ) );
  DFFX1_HVT \ram_reg[2][19]  ( .D(n592), .CLK(clk), .Q(\ram[2][19] ) );
  DFFX1_HVT \ram_reg[2][18]  ( .D(n591), .CLK(clk), .Q(\ram[2][18] ) );
  DFFX1_HVT \ram_reg[2][17]  ( .D(n590), .CLK(clk), .Q(\ram[2][17] ) );
  DFFX1_HVT \ram_reg[2][16]  ( .D(n589), .CLK(clk), .Q(\ram[2][16] ) );
  DFFX1_HVT \ram_reg[2][15]  ( .D(n588), .CLK(clk), .Q(\ram[2][15] ) );
  DFFX1_HVT \ram_reg[2][14]  ( .D(n587), .CLK(clk), .Q(\ram[2][14] ) );
  DFFX1_HVT \ram_reg[2][13]  ( .D(n586), .CLK(clk), .Q(\ram[2][13] ) );
  DFFX1_HVT \ram_reg[2][12]  ( .D(n585), .CLK(clk), .Q(\ram[2][12] ) );
  DFFX1_HVT \ram_reg[2][11]  ( .D(n584), .CLK(clk), .Q(\ram[2][11] ) );
  DFFX1_HVT \ram_reg[2][10]  ( .D(n583), .CLK(clk), .Q(\ram[2][10] ) );
  DFFX1_HVT \ram_reg[2][9]  ( .D(n582), .CLK(clk), .Q(\ram[2][9] ) );
  DFFX1_HVT \ram_reg[2][8]  ( .D(n581), .CLK(clk), .Q(\ram[2][8] ) );
  DFFX1_HVT \ram_reg[2][7]  ( .D(n580), .CLK(clk), .Q(\ram[2][7] ), .QN(n6403)
         );
  DFFX1_HVT \ram_reg[2][6]  ( .D(n579), .CLK(clk), .Q(\ram[2][6] ) );
  DFFX1_HVT \ram_reg[2][5]  ( .D(n578), .CLK(clk), .Q(\ram[2][5] ) );
  DFFX1_HVT \ram_reg[2][4]  ( .D(n577), .CLK(clk), .Q(\ram[2][4] ) );
  DFFX1_HVT \ram_reg[2][3]  ( .D(n576), .CLK(clk), .Q(\ram[2][3] ) );
  DFFX1_HVT \ram_reg[2][2]  ( .D(n575), .CLK(clk), .Q(\ram[2][2] ) );
  DFFX1_HVT \ram_reg[2][1]  ( .D(n574), .CLK(clk), .Q(\ram[2][1] ) );
  DFFX1_HVT \ram_reg[2][0]  ( .D(n573), .CLK(clk), .Q(\ram[2][0] ) );
  DFFX1_HVT \ram_reg[1][255]  ( .D(n572), .CLK(clk), .Q(\ram[1][255] ) );
  DFFX1_HVT \ram_reg[1][254]  ( .D(n571), .CLK(clk), .Q(\ram[1][254] ) );
  DFFX1_HVT \ram_reg[1][253]  ( .D(n570), .CLK(clk), .Q(\ram[1][253] ) );
  DFFX1_HVT \ram_reg[1][252]  ( .D(n569), .CLK(clk), .Q(\ram[1][252] ), .QN(
        n4237) );
  DFFX1_HVT \ram_reg[1][251]  ( .D(n568), .CLK(clk), .Q(\ram[1][251] ) );
  DFFX1_HVT \ram_reg[1][250]  ( .D(n567), .CLK(clk), .Q(\ram[1][250] ) );
  DFFX1_HVT \ram_reg[1][249]  ( .D(n566), .CLK(clk), .Q(\ram[1][249] ) );
  DFFX1_HVT \ram_reg[1][248]  ( .D(n565), .CLK(clk), .Q(\ram[1][248] ) );
  DFFX1_HVT \ram_reg[1][247]  ( .D(n564), .CLK(clk), .Q(\ram[1][247] ) );
  DFFX1_HVT \ram_reg[1][246]  ( .D(n563), .CLK(clk), .Q(\ram[1][246] ) );
  DFFX1_HVT \ram_reg[1][245]  ( .D(n562), .CLK(clk), .Q(\ram[1][245] ) );
  DFFX1_HVT \ram_reg[1][244]  ( .D(n561), .CLK(clk), .Q(\ram[1][244] ), .QN(
        n4348) );
  DFFX1_HVT \ram_reg[1][243]  ( .D(n560), .CLK(clk), .Q(\ram[1][243] ) );
  DFFX1_HVT \ram_reg[1][242]  ( .D(n559), .CLK(clk), .Q(\ram[1][242] ) );
  DFFX1_HVT \ram_reg[1][241]  ( .D(n558), .CLK(clk), .Q(\ram[1][241] ) );
  DFFX1_HVT \ram_reg[1][240]  ( .D(n557), .CLK(clk), .Q(\ram[1][240] ) );
  DFFX1_HVT \ram_reg[1][239]  ( .D(n556), .CLK(clk), .Q(\ram[1][239] ) );
  DFFX1_HVT \ram_reg[1][238]  ( .D(n555), .CLK(clk), .Q(\ram[1][238] ) );
  DFFX1_HVT \ram_reg[1][237]  ( .D(n554), .CLK(clk), .Q(\ram[1][237] ) );
  DFFX1_HVT \ram_reg[1][236]  ( .D(n553), .CLK(clk), .Q(\ram[1][236] ) );
  DFFX1_HVT \ram_reg[1][235]  ( .D(n552), .CLK(clk), .Q(\ram[1][235] ) );
  DFFX1_HVT \ram_reg[1][234]  ( .D(n551), .CLK(clk), .Q(\ram[1][234] ) );
  DFFX1_HVT \ram_reg[1][233]  ( .D(n550), .CLK(clk), .Q(\ram[1][233] ) );
  DFFX1_HVT \ram_reg[1][232]  ( .D(n549), .CLK(clk), .Q(\ram[1][232] ) );
  DFFX1_HVT \ram_reg[1][231]  ( .D(n548), .CLK(clk), .Q(\ram[1][231] ) );
  DFFX1_HVT \ram_reg[1][230]  ( .D(n547), .CLK(clk), .Q(\ram[1][230] ) );
  DFFX1_HVT \ram_reg[1][229]  ( .D(n546), .CLK(clk), .Q(\ram[1][229] ) );
  DFFX1_HVT \ram_reg[1][228]  ( .D(n545), .CLK(clk), .Q(\ram[1][228] ) );
  DFFX1_HVT \ram_reg[1][227]  ( .D(n544), .CLK(clk), .Q(\ram[1][227] ) );
  DFFX1_HVT \ram_reg[1][226]  ( .D(n543), .CLK(clk), .Q(\ram[1][226] ) );
  DFFX1_HVT \ram_reg[1][225]  ( .D(n542), .CLK(clk), .Q(\ram[1][225] ) );
  DFFX1_HVT \ram_reg[1][224]  ( .D(n541), .CLK(clk), .Q(\ram[1][224] ), .QN(
        n5167) );
  DFFX1_HVT \ram_reg[1][223]  ( .D(n540), .CLK(clk), .Q(\ram[1][223] ) );
  DFFX1_HVT \ram_reg[1][222]  ( .D(n539), .CLK(clk), .Q(\ram[1][222] ) );
  DFFX1_HVT \ram_reg[1][221]  ( .D(n538), .CLK(clk), .Q(\ram[1][221] ) );
  DFFX1_HVT \ram_reg[1][220]  ( .D(n537), .CLK(clk), .Q(\ram[1][220] ) );
  DFFX1_HVT \ram_reg[1][219]  ( .D(n536), .CLK(clk), .Q(\ram[1][219] ) );
  DFFX1_HVT \ram_reg[1][218]  ( .D(n535), .CLK(clk), .Q(\ram[1][218] ) );
  DFFX1_HVT \ram_reg[1][217]  ( .D(n534), .CLK(clk), .Q(\ram[1][217] ) );
  DFFX1_HVT \ram_reg[1][216]  ( .D(n533), .CLK(clk), .Q(\ram[1][216] ) );
  DFFX1_HVT \ram_reg[1][215]  ( .D(n532), .CLK(clk), .Q(\ram[1][215] ) );
  DFFX1_HVT \ram_reg[1][214]  ( .D(n531), .CLK(clk), .Q(\ram[1][214] ) );
  DFFX1_HVT \ram_reg[1][213]  ( .D(n530), .CLK(clk), .Q(\ram[1][213] ) );
  DFFX1_HVT \ram_reg[1][212]  ( .D(n529), .CLK(clk), .Q(\ram[1][212] ) );
  DFFX1_HVT \ram_reg[1][211]  ( .D(n528), .CLK(clk), .Q(\ram[1][211] ) );
  DFFX1_HVT \ram_reg[1][210]  ( .D(n527), .CLK(clk), .Q(\ram[1][210] ) );
  DFFX1_HVT \ram_reg[1][209]  ( .D(n526), .CLK(clk), .Q(\ram[1][209] ) );
  DFFX1_HVT \ram_reg[1][208]  ( .D(n525), .CLK(clk), .Q(\ram[1][208] ) );
  DFFX1_HVT \ram_reg[1][207]  ( .D(n524), .CLK(clk), .Q(\ram[1][207] ) );
  DFFX1_HVT \ram_reg[1][206]  ( .D(n523), .CLK(clk), .Q(\ram[1][206] ) );
  DFFX1_HVT \ram_reg[1][205]  ( .D(n522), .CLK(clk), .Q(\ram[1][205] ) );
  DFFX1_HVT \ram_reg[1][204]  ( .D(n521), .CLK(clk), .Q(\ram[1][204] ) );
  DFFX1_HVT \ram_reg[1][203]  ( .D(n520), .CLK(clk), .Q(\ram[1][203] ) );
  DFFX1_HVT \ram_reg[1][202]  ( .D(n519), .CLK(clk), .Q(\ram[1][202] ) );
  DFFX1_HVT \ram_reg[1][201]  ( .D(n518), .CLK(clk), .Q(\ram[1][201] ) );
  DFFX1_HVT \ram_reg[1][200]  ( .D(n517), .CLK(clk), .Q(\ram[1][200] ) );
  DFFX1_HVT \ram_reg[1][199]  ( .D(n516), .CLK(clk), .Q(\ram[1][199] ) );
  DFFX1_HVT \ram_reg[1][198]  ( .D(n515), .CLK(clk), .Q(\ram[1][198] ) );
  DFFX1_HVT \ram_reg[1][197]  ( .D(n514), .CLK(clk), .Q(\ram[1][197] ) );
  DFFX1_HVT \ram_reg[1][196]  ( .D(n513), .CLK(clk), .Q(\ram[1][196] ) );
  DFFX1_HVT \ram_reg[1][195]  ( .D(n512), .CLK(clk), .Q(\ram[1][195] ) );
  DFFX1_HVT \ram_reg[1][194]  ( .D(n511), .CLK(clk), .Q(\ram[1][194] ) );
  DFFX1_HVT \ram_reg[1][193]  ( .D(n510), .CLK(clk), .Q(\ram[1][193] ) );
  DFFX1_HVT \ram_reg[1][192]  ( .D(n509), .CLK(clk), .Q(\ram[1][192] ) );
  DFFX1_HVT \ram_reg[1][191]  ( .D(n508), .CLK(clk), .Q(\ram[1][191] ) );
  DFFX1_HVT \ram_reg[1][190]  ( .D(n507), .CLK(clk), .Q(\ram[1][190] ) );
  DFFX1_HVT \ram_reg[1][189]  ( .D(n506), .CLK(clk), .Q(\ram[1][189] ) );
  DFFX1_HVT \ram_reg[1][188]  ( .D(n505), .CLK(clk), .Q(\ram[1][188] ) );
  DFFX1_HVT \ram_reg[1][187]  ( .D(n504), .CLK(clk), .Q(\ram[1][187] ) );
  DFFX1_HVT \ram_reg[1][186]  ( .D(n503), .CLK(clk), .Q(\ram[1][186] ) );
  DFFX1_HVT \ram_reg[1][185]  ( .D(n502), .CLK(clk), .Q(\ram[1][185] ) );
  DFFX1_HVT \ram_reg[1][184]  ( .D(n501), .CLK(clk), .Q(\ram[1][184] ) );
  DFFX1_HVT \ram_reg[1][183]  ( .D(n500), .CLK(clk), .Q(\ram[1][183] ) );
  DFFX1_HVT \ram_reg[1][182]  ( .D(n499), .CLK(clk), .Q(\ram[1][182] ) );
  DFFX1_HVT \ram_reg[1][181]  ( .D(n498), .CLK(clk), .Q(\ram[1][181] ) );
  DFFX1_HVT \ram_reg[1][180]  ( .D(n497), .CLK(clk), .Q(\ram[1][180] ) );
  DFFX1_HVT \ram_reg[1][179]  ( .D(n496), .CLK(clk), .Q(\ram[1][179] ) );
  DFFX1_HVT \ram_reg[1][178]  ( .D(n495), .CLK(clk), .Q(\ram[1][178] ) );
  DFFX1_HVT \ram_reg[1][177]  ( .D(n494), .CLK(clk), .Q(\ram[1][177] ) );
  DFFX1_HVT \ram_reg[1][176]  ( .D(n493), .CLK(clk), .Q(\ram[1][176] ) );
  DFFX1_HVT \ram_reg[1][175]  ( .D(n492), .CLK(clk), .Q(\ram[1][175] ) );
  DFFX1_HVT \ram_reg[1][174]  ( .D(n491), .CLK(clk), .Q(\ram[1][174] ) );
  DFFX1_HVT \ram_reg[1][173]  ( .D(n490), .CLK(clk), .Q(\ram[1][173] ) );
  DFFX1_HVT \ram_reg[1][172]  ( .D(n489), .CLK(clk), .Q(\ram[1][172] ) );
  DFFX1_HVT \ram_reg[1][171]  ( .D(n488), .CLK(clk), .Q(\ram[1][171] ) );
  DFFX1_HVT \ram_reg[1][170]  ( .D(n487), .CLK(clk), .Q(\ram[1][170] ) );
  DFFX1_HVT \ram_reg[1][169]  ( .D(n486), .CLK(clk), .Q(\ram[1][169] ) );
  DFFX1_HVT \ram_reg[1][168]  ( .D(n485), .CLK(clk), .Q(\ram[1][168] ), .QN(
        n4887) );
  DFFX1_HVT \ram_reg[1][167]  ( .D(n484), .CLK(clk), .Q(\ram[1][167] ) );
  DFFX1_HVT \ram_reg[1][166]  ( .D(n483), .CLK(clk), .Q(\ram[1][166] ) );
  DFFX1_HVT \ram_reg[1][165]  ( .D(n482), .CLK(clk), .Q(\ram[1][165] ) );
  DFFX1_HVT \ram_reg[1][164]  ( .D(n481), .CLK(clk), .Q(\ram[1][164] ) );
  DFFX1_HVT \ram_reg[1][163]  ( .D(n480), .CLK(clk), .Q(\ram[1][163] ) );
  DFFX1_HVT \ram_reg[1][162]  ( .D(n479), .CLK(clk), .Q(\ram[1][162] ) );
  DFFX1_HVT \ram_reg[1][161]  ( .D(n478), .CLK(clk), .Q(\ram[1][161] ) );
  DFFX1_HVT \ram_reg[1][160]  ( .D(n477), .CLK(clk), .Q(\ram[1][160] ) );
  DFFX1_HVT \ram_reg[1][159]  ( .D(n476), .CLK(clk), .Q(\ram[1][159] ) );
  DFFX1_HVT \ram_reg[1][158]  ( .D(n475), .CLK(clk), .Q(\ram[1][158] ) );
  DFFX1_HVT \ram_reg[1][157]  ( .D(n474), .CLK(clk), .Q(\ram[1][157] ) );
  DFFX1_HVT \ram_reg[1][156]  ( .D(n473), .CLK(clk), .Q(\ram[1][156] ) );
  DFFX1_HVT \ram_reg[1][155]  ( .D(n472), .CLK(clk), .Q(\ram[1][155] ) );
  DFFX1_HVT \ram_reg[1][154]  ( .D(n471), .CLK(clk), .Q(\ram[1][154] ) );
  DFFX1_HVT \ram_reg[1][153]  ( .D(n470), .CLK(clk), .Q(\ram[1][153] ) );
  DFFX1_HVT \ram_reg[1][152]  ( .D(n469), .CLK(clk), .Q(\ram[1][152] ) );
  DFFX1_HVT \ram_reg[1][151]  ( .D(n468), .CLK(clk), .Q(\ram[1][151] ) );
  DFFX1_HVT \ram_reg[1][150]  ( .D(n467), .CLK(clk), .Q(\ram[1][150] ) );
  DFFX1_HVT \ram_reg[1][149]  ( .D(n466), .CLK(clk), .Q(\ram[1][149] ) );
  DFFX1_HVT \ram_reg[1][148]  ( .D(n465), .CLK(clk), .Q(\ram[1][148] ) );
  DFFX1_HVT \ram_reg[1][147]  ( .D(n464), .CLK(clk), .Q(\ram[1][147] ), .QN(
        n866) );
  DFFX1_HVT \ram_reg[1][146]  ( .D(n463), .CLK(clk), .Q(\ram[1][146] ) );
  DFFX1_HVT \ram_reg[1][145]  ( .D(n462), .CLK(clk), .Q(\ram[1][145] ) );
  DFFX1_HVT \ram_reg[1][144]  ( .D(n461), .CLK(clk), .Q(\ram[1][144] ) );
  DFFX1_HVT \ram_reg[1][143]  ( .D(n460), .CLK(clk), .Q(\ram[1][143] ) );
  DFFX1_HVT \ram_reg[1][142]  ( .D(n459), .CLK(clk), .Q(\ram[1][142] ) );
  DFFX1_HVT \ram_reg[1][141]  ( .D(n458), .CLK(clk), .Q(\ram[1][141] ) );
  DFFX1_HVT \ram_reg[1][140]  ( .D(n457), .CLK(clk), .Q(\ram[1][140] ) );
  DFFX1_HVT \ram_reg[1][139]  ( .D(n456), .CLK(clk), .Q(\ram[1][139] ) );
  DFFX1_HVT \ram_reg[1][138]  ( .D(n455), .CLK(clk), .Q(\ram[1][138] ) );
  DFFX1_HVT \ram_reg[1][137]  ( .D(n454), .CLK(clk), .Q(\ram[1][137] ) );
  DFFX1_HVT \ram_reg[1][136]  ( .D(n453), .CLK(clk), .Q(\ram[1][136] ) );
  DFFX1_HVT \ram_reg[1][135]  ( .D(n452), .CLK(clk), .Q(\ram[1][135] ) );
  DFFX1_HVT \ram_reg[1][134]  ( .D(n451), .CLK(clk), .Q(\ram[1][134] ) );
  DFFX1_HVT \ram_reg[1][133]  ( .D(n450), .CLK(clk), .Q(\ram[1][133] ) );
  DFFX1_HVT \ram_reg[1][132]  ( .D(n449), .CLK(clk), .Q(\ram[1][132] ) );
  DFFX1_HVT \ram_reg[1][131]  ( .D(n448), .CLK(clk), .Q(\ram[1][131] ) );
  DFFX1_HVT \ram_reg[1][130]  ( .D(n447), .CLK(clk), .Q(\ram[1][130] ) );
  DFFX1_HVT \ram_reg[1][129]  ( .D(n446), .CLK(clk), .Q(\ram[1][129] ) );
  DFFX1_HVT \ram_reg[1][128]  ( .D(n445), .CLK(clk), .Q(\ram[1][128] ) );
  DFFX1_HVT \ram_reg[1][127]  ( .D(n444), .CLK(clk), .Q(\ram[1][127] ) );
  DFFX1_HVT \ram_reg[1][126]  ( .D(n443), .CLK(clk), .Q(\ram[1][126] ) );
  DFFX1_HVT \ram_reg[1][125]  ( .D(n442), .CLK(clk), .Q(\ram[1][125] ) );
  DFFX1_HVT \ram_reg[1][124]  ( .D(n441), .CLK(clk), .Q(\ram[1][124] ) );
  DFFX1_HVT \ram_reg[1][123]  ( .D(n440), .CLK(clk), .Q(\ram[1][123] ) );
  DFFX1_HVT \ram_reg[1][122]  ( .D(n439), .CLK(clk), .Q(\ram[1][122] ), .QN(
        n4219) );
  DFFX1_HVT \ram_reg[1][121]  ( .D(n438), .CLK(clk), .Q(\ram[1][121] ) );
  DFFX1_HVT \ram_reg[1][120]  ( .D(n437), .CLK(clk), .Q(\ram[1][120] ), .QN(
        n4890) );
  DFFX1_HVT \ram_reg[1][119]  ( .D(n436), .CLK(clk), .Q(\ram[1][119] ) );
  DFFX1_HVT \ram_reg[1][118]  ( .D(n435), .CLK(clk), .Q(\ram[1][118] ) );
  DFFX1_HVT \ram_reg[1][117]  ( .D(n434), .CLK(clk), .Q(\ram[1][117] ) );
  DFFX1_HVT \ram_reg[1][116]  ( .D(n433), .CLK(clk), .Q(\ram[1][116] ) );
  DFFX1_HVT \ram_reg[1][115]  ( .D(n432), .CLK(clk), .Q(\ram[1][115] ) );
  DFFX1_HVT \ram_reg[1][114]  ( .D(n431), .CLK(clk), .Q(\ram[1][114] ) );
  DFFX1_HVT \ram_reg[1][113]  ( .D(n430), .CLK(clk), .Q(\ram[1][113] ) );
  DFFX1_HVT \ram_reg[1][112]  ( .D(n429), .CLK(clk), .Q(\ram[1][112] ), .QN(
        n5439) );
  DFFX1_HVT \ram_reg[1][111]  ( .D(n428), .CLK(clk), .Q(\ram[1][111] ) );
  DFFX1_HVT \ram_reg[1][110]  ( .D(n427), .CLK(clk), .Q(\ram[1][110] ) );
  DFFX1_HVT \ram_reg[1][109]  ( .D(n426), .CLK(clk), .Q(\ram[1][109] ) );
  DFFX1_HVT \ram_reg[1][108]  ( .D(n425), .CLK(clk), .Q(\ram[1][108] ) );
  DFFX1_HVT \ram_reg[1][107]  ( .D(n424), .CLK(clk), .Q(\ram[1][107] ) );
  DFFX1_HVT \ram_reg[1][106]  ( .D(n423), .CLK(clk), .Q(\ram[1][106] ) );
  DFFX1_HVT \ram_reg[1][105]  ( .D(n422), .CLK(clk), .Q(\ram[1][105] ) );
  DFFX1_HVT \ram_reg[1][104]  ( .D(n421), .CLK(clk), .Q(\ram[1][104] ) );
  DFFX1_HVT \ram_reg[1][103]  ( .D(n420), .CLK(clk), .Q(\ram[1][103] ) );
  DFFX1_HVT \ram_reg[1][102]  ( .D(n419), .CLK(clk), .Q(\ram[1][102] ) );
  DFFX1_HVT \ram_reg[1][101]  ( .D(n418), .CLK(clk), .Q(\ram[1][101] ) );
  DFFX1_HVT \ram_reg[1][100]  ( .D(n417), .CLK(clk), .Q(\ram[1][100] ) );
  DFFX1_HVT \ram_reg[1][99]  ( .D(n416), .CLK(clk), .Q(\ram[1][99] ) );
  DFFX1_HVT \ram_reg[1][98]  ( .D(n415), .CLK(clk), .Q(\ram[1][98] ) );
  DFFX1_HVT \ram_reg[1][97]  ( .D(n414), .CLK(clk), .Q(\ram[1][97] ) );
  DFFX1_HVT \ram_reg[1][96]  ( .D(n413), .CLK(clk), .Q(\ram[1][96] ) );
  DFFX1_HVT \ram_reg[1][95]  ( .D(n412), .CLK(clk), .Q(\ram[1][95] ) );
  DFFX1_HVT \ram_reg[1][94]  ( .D(n411), .CLK(clk), .Q(\ram[1][94] ) );
  DFFX1_HVT \ram_reg[1][93]  ( .D(n410), .CLK(clk), .Q(\ram[1][93] ) );
  DFFX1_HVT \ram_reg[1][92]  ( .D(n409), .CLK(clk), .Q(\ram[1][92] ) );
  DFFX1_HVT \ram_reg[1][91]  ( .D(n408), .CLK(clk), .Q(\ram[1][91] ) );
  DFFX1_HVT \ram_reg[1][90]  ( .D(n407), .CLK(clk), .Q(\ram[1][90] ) );
  DFFX1_HVT \ram_reg[1][89]  ( .D(n406), .CLK(clk), .Q(\ram[1][89] ) );
  DFFX1_HVT \ram_reg[1][88]  ( .D(n405), .CLK(clk), .Q(\ram[1][88] ), .QN(
        n5482) );
  DFFX1_HVT \ram_reg[1][87]  ( .D(n404), .CLK(clk), .Q(\ram[1][87] ) );
  DFFX1_HVT \ram_reg[1][86]  ( .D(n403), .CLK(clk), .Q(\ram[1][86] ), .QN(
        n4671) );
  DFFX1_HVT \ram_reg[1][85]  ( .D(n402), .CLK(clk), .Q(\ram[1][85] ) );
  DFFX1_HVT \ram_reg[1][84]  ( .D(n401), .CLK(clk), .Q(\ram[1][84] ) );
  DFFX1_HVT \ram_reg[1][83]  ( .D(n400), .CLK(clk), .Q(\ram[1][83] ) );
  DFFX1_HVT \ram_reg[1][82]  ( .D(n399), .CLK(clk), .Q(\ram[1][82] ) );
  DFFX1_HVT \ram_reg[1][81]  ( .D(n398), .CLK(clk), .Q(\ram[1][81] ) );
  DFFX1_HVT \ram_reg[1][80]  ( .D(n397), .CLK(clk), .Q(\ram[1][80] ) );
  DFFX1_HVT \ram_reg[1][79]  ( .D(n396), .CLK(clk), .Q(\ram[1][79] ) );
  DFFX1_HVT \ram_reg[1][78]  ( .D(n395), .CLK(clk), .Q(\ram[1][78] ) );
  DFFX1_HVT \ram_reg[1][77]  ( .D(n394), .CLK(clk), .Q(\ram[1][77] ) );
  DFFX1_HVT \ram_reg[1][76]  ( .D(n393), .CLK(clk), .Q(\ram[1][76] ) );
  DFFX1_HVT \ram_reg[1][75]  ( .D(n392), .CLK(clk), .Q(\ram[1][75] ) );
  DFFX1_HVT \ram_reg[1][74]  ( .D(n391), .CLK(clk), .Q(\ram[1][74] ) );
  DFFX1_HVT \ram_reg[1][73]  ( .D(n390), .CLK(clk), .Q(\ram[1][73] ) );
  DFFX1_HVT \ram_reg[1][72]  ( .D(n389), .CLK(clk), .Q(\ram[1][72] ) );
  DFFX1_HVT \ram_reg[1][71]  ( .D(n388), .CLK(clk), .Q(\ram[1][71] ) );
  DFFX1_HVT \ram_reg[1][70]  ( .D(n387), .CLK(clk), .Q(\ram[1][70] ) );
  DFFX1_HVT \ram_reg[1][69]  ( .D(n386), .CLK(clk), .Q(\ram[1][69] ) );
  DFFX1_HVT \ram_reg[1][68]  ( .D(n385), .CLK(clk), .Q(\ram[1][68] ) );
  DFFX1_HVT \ram_reg[1][67]  ( .D(n384), .CLK(clk), .Q(\ram[1][67] ) );
  DFFX1_HVT \ram_reg[1][66]  ( .D(n383), .CLK(clk), .Q(\ram[1][66] ) );
  DFFX1_HVT \ram_reg[1][65]  ( .D(n382), .CLK(clk), .Q(\ram[1][65] ) );
  DFFX1_HVT \ram_reg[1][64]  ( .D(n381), .CLK(clk), .Q(\ram[1][64] ) );
  DFFX1_HVT \ram_reg[1][63]  ( .D(n380), .CLK(clk), .Q(\ram[1][63] ) );
  DFFX1_HVT \ram_reg[1][62]  ( .D(n379), .CLK(clk), .Q(\ram[1][62] ) );
  DFFX1_HVT \ram_reg[1][61]  ( .D(n378), .CLK(clk), .Q(\ram[1][61] ) );
  DFFX1_HVT \ram_reg[1][60]  ( .D(n377), .CLK(clk), .Q(\ram[1][60] ) );
  DFFX1_HVT \ram_reg[1][59]  ( .D(n376), .CLK(clk), .Q(\ram[1][59] ) );
  DFFX1_HVT \ram_reg[1][58]  ( .D(n375), .CLK(clk), .Q(\ram[1][58] ) );
  DFFX1_HVT \ram_reg[1][57]  ( .D(n374), .CLK(clk), .Q(\ram[1][57] ) );
  DFFX1_HVT \ram_reg[1][56]  ( .D(n373), .CLK(clk), .Q(\ram[1][56] ) );
  DFFX1_HVT \ram_reg[1][55]  ( .D(n372), .CLK(clk), .Q(\ram[1][55] ) );
  DFFX1_HVT \ram_reg[1][54]  ( .D(n371), .CLK(clk), .Q(\ram[1][54] ) );
  DFFX1_HVT \ram_reg[1][53]  ( .D(n370), .CLK(clk), .Q(\ram[1][53] ) );
  DFFX1_HVT \ram_reg[1][52]  ( .D(n369), .CLK(clk), .Q(\ram[1][52] ) );
  DFFX1_HVT \ram_reg[1][51]  ( .D(n368), .CLK(clk), .Q(\ram[1][51] ) );
  DFFX1_HVT \ram_reg[1][50]  ( .D(n367), .CLK(clk), .Q(\ram[1][50] ) );
  DFFX1_HVT \ram_reg[1][49]  ( .D(n366), .CLK(clk), .Q(\ram[1][49] ) );
  DFFX1_HVT \ram_reg[1][48]  ( .D(n365), .CLK(clk), .Q(\ram[1][48] ) );
  DFFX1_HVT \ram_reg[1][47]  ( .D(n364), .CLK(clk), .Q(\ram[1][47] ) );
  DFFX1_HVT \ram_reg[1][46]  ( .D(n363), .CLK(clk), .Q(\ram[1][46] ) );
  DFFX1_HVT \ram_reg[1][45]  ( .D(n362), .CLK(clk), .Q(\ram[1][45] ), .QN(
        n4674) );
  DFFX1_HVT \ram_reg[1][44]  ( .D(n361), .CLK(clk), .Q(\ram[1][44] ) );
  DFFX1_HVT \ram_reg[1][43]  ( .D(n360), .CLK(clk), .Q(\ram[1][43] ) );
  DFFX1_HVT \ram_reg[1][42]  ( .D(n359), .CLK(clk), .Q(\ram[1][42] ), .QN(
        n4865) );
  DFFX1_HVT \ram_reg[1][41]  ( .D(n358), .CLK(clk), .Q(\ram[1][41] ) );
  DFFX1_HVT \ram_reg[1][40]  ( .D(n357), .CLK(clk), .Q(\ram[1][40] ), .QN(
        n4866) );
  DFFX1_HVT \ram_reg[1][39]  ( .D(n356), .CLK(clk), .Q(\ram[1][39] ) );
  DFFX1_HVT \ram_reg[1][38]  ( .D(n355), .CLK(clk), .Q(\ram[1][38] ) );
  DFFX1_HVT \ram_reg[1][37]  ( .D(n354), .CLK(clk), .Q(\ram[1][37] ) );
  DFFX1_HVT \ram_reg[1][36]  ( .D(n353), .CLK(clk), .Q(\ram[1][36] ) );
  DFFX1_HVT \ram_reg[1][35]  ( .D(n352), .CLK(clk), .Q(\ram[1][35] ) );
  DFFX1_HVT \ram_reg[1][34]  ( .D(n351), .CLK(clk), .Q(\ram[1][34] ) );
  DFFX1_HVT \ram_reg[1][33]  ( .D(n350), .CLK(clk), .Q(\ram[1][33] ) );
  DFFX1_HVT \ram_reg[1][32]  ( .D(n349), .CLK(clk), .Q(\ram[1][32] ) );
  DFFX1_HVT \ram_reg[1][31]  ( .D(n348), .CLK(clk), .Q(\ram[1][31] ) );
  DFFX1_HVT \ram_reg[1][30]  ( .D(n347), .CLK(clk), .Q(\ram[1][30] ) );
  DFFX1_HVT \ram_reg[1][29]  ( .D(n346), .CLK(clk), .Q(\ram[1][29] ), .QN(
        n4603) );
  DFFX1_HVT \ram_reg[1][28]  ( .D(n345), .CLK(clk), .Q(\ram[1][28] ) );
  DFFX1_HVT \ram_reg[1][27]  ( .D(n344), .CLK(clk), .Q(\ram[1][27] ) );
  DFFX1_HVT \ram_reg[1][26]  ( .D(n343), .CLK(clk), .Q(\ram[1][26] ) );
  DFFX1_HVT \ram_reg[1][25]  ( .D(n342), .CLK(clk), .Q(\ram[1][25] ) );
  DFFX1_HVT \ram_reg[1][24]  ( .D(n341), .CLK(clk), .Q(\ram[1][24] ) );
  DFFX1_HVT \ram_reg[1][23]  ( .D(n340), .CLK(clk), .Q(\ram[1][23] ) );
  DFFX1_HVT \ram_reg[1][22]  ( .D(n339), .CLK(clk), .Q(\ram[1][22] ) );
  DFFX1_HVT \ram_reg[1][21]  ( .D(n338), .CLK(clk), .Q(\ram[1][21] ) );
  DFFX1_HVT \ram_reg[1][20]  ( .D(n337), .CLK(clk), .Q(\ram[1][20] ) );
  DFFX1_HVT \ram_reg[1][19]  ( .D(n336), .CLK(clk), .Q(\ram[1][19] ) );
  DFFX1_HVT \ram_reg[1][18]  ( .D(n335), .CLK(clk), .Q(\ram[1][18] ) );
  DFFX1_HVT \ram_reg[1][17]  ( .D(n334), .CLK(clk), .Q(\ram[1][17] ) );
  DFFX1_HVT \ram_reg[1][16]  ( .D(n333), .CLK(clk), .Q(\ram[1][16] ) );
  DFFX1_HVT \ram_reg[1][15]  ( .D(n332), .CLK(clk), .Q(\ram[1][15] ) );
  DFFX1_HVT \ram_reg[1][14]  ( .D(n331), .CLK(clk), .Q(\ram[1][14] ) );
  DFFX1_HVT \ram_reg[1][13]  ( .D(n330), .CLK(clk), .Q(\ram[1][13] ) );
  DFFX1_HVT \ram_reg[1][12]  ( .D(n329), .CLK(clk), .Q(\ram[1][12] ) );
  DFFX1_HVT \ram_reg[1][11]  ( .D(n328), .CLK(clk), .Q(\ram[1][11] ) );
  DFFX1_HVT \ram_reg[1][10]  ( .D(n327), .CLK(clk), .Q(\ram[1][10] ), .QN(
        n4579) );
  DFFX1_HVT \ram_reg[1][9]  ( .D(n326), .CLK(clk), .Q(\ram[1][9] ) );
  DFFX1_HVT \ram_reg[1][8]  ( .D(n325), .CLK(clk), .Q(\ram[1][8] ) );
  DFFX1_HVT \ram_reg[1][7]  ( .D(n324), .CLK(clk), .Q(\ram[1][7] ), .QN(n5440)
         );
  DFFX1_HVT \ram_reg[1][6]  ( .D(n323), .CLK(clk), .Q(\ram[1][6] ) );
  DFFX1_HVT \ram_reg[1][5]  ( .D(n322), .CLK(clk), .Q(\ram[1][5] ) );
  DFFX1_HVT \ram_reg[1][4]  ( .D(n321), .CLK(clk), .Q(\ram[1][4] ) );
  DFFX1_HVT \ram_reg[1][3]  ( .D(n320), .CLK(clk), .Q(\ram[1][3] ) );
  DFFX1_HVT \ram_reg[1][2]  ( .D(n319), .CLK(clk), .Q(\ram[1][2] ) );
  DFFX1_HVT \ram_reg[1][1]  ( .D(n318), .CLK(clk), .Q(\ram[1][1] ) );
  DFFX1_HVT \ram_reg[1][0]  ( .D(n317), .CLK(clk), .Q(\ram[1][0] ) );
  DFFX1_HVT \ram_reg[0][255]  ( .D(n316), .CLK(clk), .Q(\ram[0][255] ) );
  DFFX1_HVT \ram_reg[0][254]  ( .D(n315), .CLK(clk), .Q(\ram[0][254] ) );
  DFFX1_HVT \ram_reg[0][253]  ( .D(n314), .CLK(clk), .Q(\ram[0][253] ) );
  DFFX1_HVT \ram_reg[0][252]  ( .D(n313), .CLK(clk), .Q(\ram[0][252] ) );
  DFFX1_HVT \ram_reg[0][251]  ( .D(n312), .CLK(clk), .Q(\ram[0][251] ) );
  DFFX1_HVT \ram_reg[0][250]  ( .D(n311), .CLK(clk), .Q(\ram[0][250] ) );
  DFFX1_HVT \ram_reg[0][249]  ( .D(n310), .CLK(clk), .Q(\ram[0][249] ) );
  DFFX1_HVT \ram_reg[0][248]  ( .D(n309), .CLK(clk), .Q(\ram[0][248] ) );
  DFFX1_HVT \ram_reg[0][247]  ( .D(n308), .CLK(clk), .Q(\ram[0][247] ) );
  DFFX1_HVT \ram_reg[0][246]  ( .D(n307), .CLK(clk), .Q(\ram[0][246] ) );
  DFFX1_HVT \ram_reg[0][245]  ( .D(n306), .CLK(clk), .Q(\ram[0][245] ) );
  DFFX1_HVT \ram_reg[0][244]  ( .D(n305), .CLK(clk), .Q(\ram[0][244] ) );
  DFFX1_HVT \ram_reg[0][243]  ( .D(n304), .CLK(clk), .Q(\ram[0][243] ) );
  DFFX1_HVT \ram_reg[0][242]  ( .D(n303), .CLK(clk), .Q(\ram[0][242] ) );
  DFFX1_HVT \ram_reg[0][241]  ( .D(n302), .CLK(clk), .Q(\ram[0][241] ) );
  DFFX1_HVT \ram_reg[0][240]  ( .D(n301), .CLK(clk), .Q(\ram[0][240] ) );
  DFFX1_HVT \ram_reg[0][239]  ( .D(n300), .CLK(clk), .Q(\ram[0][239] ) );
  DFFX1_HVT \ram_reg[0][238]  ( .D(n299), .CLK(clk), .Q(\ram[0][238] ) );
  DFFX1_HVT \ram_reg[0][237]  ( .D(n298), .CLK(clk), .Q(\ram[0][237] ) );
  DFFX1_HVT \ram_reg[0][236]  ( .D(n297), .CLK(clk), .Q(\ram[0][236] ) );
  DFFX1_HVT \ram_reg[0][235]  ( .D(n296), .CLK(clk), .Q(\ram[0][235] ) );
  DFFX1_HVT \ram_reg[0][234]  ( .D(n295), .CLK(clk), .Q(\ram[0][234] ) );
  DFFX1_HVT \ram_reg[0][233]  ( .D(n294), .CLK(clk), .Q(\ram[0][233] ) );
  DFFX1_HVT \ram_reg[0][232]  ( .D(n293), .CLK(clk), .Q(\ram[0][232] ) );
  DFFX1_HVT \ram_reg[0][231]  ( .D(n292), .CLK(clk), .Q(\ram[0][231] ) );
  DFFX1_HVT \ram_reg[0][230]  ( .D(n291), .CLK(clk), .Q(\ram[0][230] ) );
  DFFX1_HVT \ram_reg[0][229]  ( .D(n290), .CLK(clk), .Q(\ram[0][229] ) );
  DFFX1_HVT \ram_reg[0][228]  ( .D(n289), .CLK(clk), .Q(\ram[0][228] ) );
  DFFX1_HVT \ram_reg[0][227]  ( .D(n288), .CLK(clk), .Q(\ram[0][227] ) );
  DFFX1_HVT \ram_reg[0][226]  ( .D(n287), .CLK(clk), .Q(\ram[0][226] ) );
  DFFX1_HVT \ram_reg[0][225]  ( .D(n286), .CLK(clk), .Q(\ram[0][225] ) );
  DFFX1_HVT \ram_reg[0][224]  ( .D(n285), .CLK(clk), .Q(\ram[0][224] ), .QN(
        n5168) );
  DFFX1_HVT \ram_reg[0][223]  ( .D(n284), .CLK(clk), .Q(\ram[0][223] ) );
  DFFX1_HVT \ram_reg[0][222]  ( .D(n283), .CLK(clk), .Q(\ram[0][222] ) );
  DFFX1_HVT \ram_reg[0][221]  ( .D(n282), .CLK(clk), .Q(\ram[0][221] ) );
  DFFX1_HVT \ram_reg[0][220]  ( .D(n281), .CLK(clk), .Q(\ram[0][220] ) );
  DFFX1_HVT \ram_reg[0][219]  ( .D(n280), .CLK(clk), .Q(\ram[0][219] ) );
  DFFX1_HVT \ram_reg[0][218]  ( .D(n279), .CLK(clk), .Q(\ram[0][218] ) );
  DFFX1_HVT \ram_reg[0][217]  ( .D(n278), .CLK(clk), .Q(\ram[0][217] ) );
  DFFX1_HVT \ram_reg[0][216]  ( .D(n277), .CLK(clk), .Q(\ram[0][216] ) );
  DFFX1_HVT \ram_reg[0][215]  ( .D(n276), .CLK(clk), .Q(\ram[0][215] ) );
  DFFX1_HVT \ram_reg[0][214]  ( .D(n275), .CLK(clk), .Q(\ram[0][214] ) );
  DFFX1_HVT \ram_reg[0][213]  ( .D(n274), .CLK(clk), .Q(\ram[0][213] ) );
  DFFX1_HVT \ram_reg[0][212]  ( .D(n273), .CLK(clk), .Q(\ram[0][212] ) );
  DFFX1_HVT \ram_reg[0][211]  ( .D(n272), .CLK(clk), .Q(\ram[0][211] ) );
  DFFX1_HVT \ram_reg[0][210]  ( .D(n271), .CLK(clk), .Q(\ram[0][210] ) );
  DFFX1_HVT \ram_reg[0][209]  ( .D(n270), .CLK(clk), .Q(\ram[0][209] ) );
  DFFX1_HVT \ram_reg[0][208]  ( .D(n269), .CLK(clk), .Q(\ram[0][208] ) );
  DFFX1_HVT \ram_reg[0][207]  ( .D(n268), .CLK(clk), .Q(\ram[0][207] ) );
  DFFX1_HVT \ram_reg[0][206]  ( .D(n267), .CLK(clk), .Q(\ram[0][206] ) );
  DFFX1_HVT \ram_reg[0][205]  ( .D(n266), .CLK(clk), .Q(\ram[0][205] ) );
  DFFX1_HVT \ram_reg[0][204]  ( .D(n265), .CLK(clk), .Q(\ram[0][204] ) );
  DFFX1_HVT \ram_reg[0][203]  ( .D(n264), .CLK(clk), .Q(\ram[0][203] ) );
  DFFX1_HVT \ram_reg[0][202]  ( .D(n263), .CLK(clk), .Q(\ram[0][202] ) );
  DFFX1_HVT \ram_reg[0][201]  ( .D(n262), .CLK(clk), .Q(\ram[0][201] ) );
  DFFX1_HVT \ram_reg[0][200]  ( .D(n261), .CLK(clk), .Q(\ram[0][200] ) );
  DFFX1_HVT \ram_reg[0][199]  ( .D(n260), .CLK(clk), .Q(\ram[0][199] ) );
  DFFX1_HVT \ram_reg[0][198]  ( .D(n259), .CLK(clk), .Q(\ram[0][198] ) );
  DFFX1_HVT \ram_reg[0][197]  ( .D(n258), .CLK(clk), .Q(\ram[0][197] ) );
  DFFX1_HVT \ram_reg[0][196]  ( .D(n257), .CLK(clk), .Q(\ram[0][196] ) );
  DFFX1_HVT \ram_reg[0][195]  ( .D(n256), .CLK(clk), .Q(\ram[0][195] ) );
  DFFX1_HVT \ram_reg[0][194]  ( .D(n255), .CLK(clk), .Q(\ram[0][194] ) );
  DFFX1_HVT \ram_reg[0][193]  ( .D(n254), .CLK(clk), .Q(\ram[0][193] ) );
  DFFX1_HVT \ram_reg[0][192]  ( .D(n253), .CLK(clk), .Q(\ram[0][192] ) );
  DFFX1_HVT \ram_reg[0][191]  ( .D(n252), .CLK(clk), .Q(\ram[0][191] ) );
  DFFX1_HVT \ram_reg[0][190]  ( .D(n251), .CLK(clk), .Q(\ram[0][190] ) );
  DFFX1_HVT \ram_reg[0][189]  ( .D(n250), .CLK(clk), .Q(\ram[0][189] ) );
  DFFX1_HVT \ram_reg[0][188]  ( .D(n249), .CLK(clk), .Q(\ram[0][188] ) );
  DFFX1_HVT \ram_reg[0][187]  ( .D(n248), .CLK(clk), .Q(\ram[0][187] ) );
  DFFX1_HVT \ram_reg[0][186]  ( .D(n247), .CLK(clk), .Q(\ram[0][186] ) );
  DFFX1_HVT \ram_reg[0][185]  ( .D(n246), .CLK(clk), .Q(\ram[0][185] ) );
  DFFX1_HVT \ram_reg[0][184]  ( .D(n245), .CLK(clk), .Q(\ram[0][184] ) );
  DFFX1_HVT \ram_reg[0][183]  ( .D(n244), .CLK(clk), .Q(\ram[0][183] ) );
  DFFX1_HVT \ram_reg[0][182]  ( .D(n243), .CLK(clk), .Q(\ram[0][182] ) );
  DFFX1_HVT \ram_reg[0][181]  ( .D(n242), .CLK(clk), .Q(\ram[0][181] ) );
  DFFX1_HVT \ram_reg[0][180]  ( .D(n241), .CLK(clk), .Q(\ram[0][180] ) );
  DFFX1_HVT \ram_reg[0][179]  ( .D(n240), .CLK(clk), .Q(\ram[0][179] ) );
  DFFX1_HVT \ram_reg[0][178]  ( .D(n239), .CLK(clk), .Q(\ram[0][178] ) );
  DFFX1_HVT \ram_reg[0][177]  ( .D(n238), .CLK(clk), .Q(\ram[0][177] ) );
  DFFX1_HVT \ram_reg[0][176]  ( .D(n237), .CLK(clk), .Q(\ram[0][176] ) );
  DFFX1_HVT \ram_reg[0][175]  ( .D(n236), .CLK(clk), .Q(\ram[0][175] ) );
  DFFX1_HVT \ram_reg[0][174]  ( .D(n235), .CLK(clk), .Q(\ram[0][174] ) );
  DFFX1_HVT \ram_reg[0][173]  ( .D(n234), .CLK(clk), .Q(\ram[0][173] ) );
  DFFX1_HVT \ram_reg[0][172]  ( .D(n233), .CLK(clk), .Q(\ram[0][172] ) );
  DFFX1_HVT \ram_reg[0][171]  ( .D(n232), .CLK(clk), .Q(\ram[0][171] ) );
  DFFX1_HVT \ram_reg[0][170]  ( .D(n231), .CLK(clk), .Q(\ram[0][170] ) );
  DFFX1_HVT \ram_reg[0][169]  ( .D(n230), .CLK(clk), .Q(\ram[0][169] ) );
  DFFX1_HVT \ram_reg[0][168]  ( .D(n229), .CLK(clk), .Q(\ram[0][168] ) );
  DFFX1_HVT \ram_reg[0][167]  ( .D(n228), .CLK(clk), .Q(\ram[0][167] ) );
  DFFX1_HVT \ram_reg[0][166]  ( .D(n227), .CLK(clk), .Q(\ram[0][166] ) );
  DFFX1_HVT \ram_reg[0][165]  ( .D(n226), .CLK(clk), .Q(\ram[0][165] ) );
  DFFX1_HVT \ram_reg[0][164]  ( .D(n225), .CLK(clk), .Q(\ram[0][164] ) );
  DFFX1_HVT \ram_reg[0][163]  ( .D(n224), .CLK(clk), .Q(\ram[0][163] ) );
  DFFX1_HVT \ram_reg[0][162]  ( .D(n223), .CLK(clk), .Q(\ram[0][162] ) );
  DFFX1_HVT \ram_reg[0][161]  ( .D(n222), .CLK(clk), .Q(\ram[0][161] ) );
  DFFX1_HVT \ram_reg[0][160]  ( .D(n221), .CLK(clk), .Q(\ram[0][160] ) );
  DFFX1_HVT \ram_reg[0][159]  ( .D(n220), .CLK(clk), .Q(\ram[0][159] ) );
  DFFX1_HVT \ram_reg[0][158]  ( .D(n219), .CLK(clk), .Q(\ram[0][158] ) );
  DFFX1_HVT \ram_reg[0][157]  ( .D(n218), .CLK(clk), .Q(\ram[0][157] ) );
  DFFX1_HVT \ram_reg[0][156]  ( .D(n217), .CLK(clk), .Q(\ram[0][156] ) );
  DFFX1_HVT \ram_reg[0][155]  ( .D(n216), .CLK(clk), .Q(\ram[0][155] ) );
  DFFX1_HVT \ram_reg[0][154]  ( .D(n215), .CLK(clk), .Q(\ram[0][154] ) );
  DFFX1_HVT \ram_reg[0][153]  ( .D(n214), .CLK(clk), .Q(\ram[0][153] ) );
  DFFX1_HVT \ram_reg[0][152]  ( .D(n213), .CLK(clk), .Q(\ram[0][152] ) );
  DFFX1_HVT \ram_reg[0][151]  ( .D(n212), .CLK(clk), .Q(\ram[0][151] ) );
  DFFX1_HVT \ram_reg[0][150]  ( .D(n211), .CLK(clk), .Q(\ram[0][150] ) );
  DFFX1_HVT \ram_reg[0][149]  ( .D(n210), .CLK(clk), .Q(\ram[0][149] ) );
  DFFX1_HVT \ram_reg[0][148]  ( .D(n209), .CLK(clk), .Q(\ram[0][148] ) );
  DFFX1_HVT \ram_reg[0][147]  ( .D(n208), .CLK(clk), .Q(\ram[0][147] ), .QN(
        n877) );
  DFFX1_HVT \ram_reg[0][146]  ( .D(n207), .CLK(clk), .Q(\ram[0][146] ) );
  DFFX1_HVT \ram_reg[0][145]  ( .D(n206), .CLK(clk), .Q(\ram[0][145] ) );
  DFFX1_HVT \ram_reg[0][144]  ( .D(n205), .CLK(clk), .Q(n4877), .QN(n5477) );
  DFFX1_HVT \ram_reg[0][143]  ( .D(n204), .CLK(clk), .Q(\ram[0][143] ) );
  DFFX1_HVT \ram_reg[0][142]  ( .D(n203), .CLK(clk), .Q(\ram[0][142] ) );
  DFFX1_HVT \ram_reg[0][141]  ( .D(n202), .CLK(clk), .Q(\ram[0][141] ) );
  DFFX1_HVT \ram_reg[0][140]  ( .D(n201), .CLK(clk), .Q(\ram[0][140] ) );
  DFFX1_HVT \ram_reg[0][139]  ( .D(n200), .CLK(clk), .Q(\ram[0][139] ) );
  DFFX1_HVT \ram_reg[0][138]  ( .D(n199), .CLK(clk), .Q(\ram[0][138] ) );
  DFFX1_HVT \ram_reg[0][137]  ( .D(n198), .CLK(clk), .Q(\ram[0][137] ) );
  DFFX1_HVT \ram_reg[0][136]  ( .D(n197), .CLK(clk), .Q(\ram[0][136] ) );
  DFFX1_HVT \ram_reg[0][135]  ( .D(n196), .CLK(clk), .Q(\ram[0][135] ) );
  DFFX1_HVT \ram_reg[0][134]  ( .D(n195), .CLK(clk), .Q(\ram[0][134] ) );
  DFFX1_HVT \ram_reg[0][133]  ( .D(n194), .CLK(clk), .Q(\ram[0][133] ) );
  DFFX1_HVT \ram_reg[0][132]  ( .D(n193), .CLK(clk), .Q(\ram[0][132] ) );
  DFFX1_HVT \ram_reg[0][131]  ( .D(n192), .CLK(clk), .Q(\ram[0][131] ) );
  DFFX1_HVT \ram_reg[0][130]  ( .D(n191), .CLK(clk), .Q(\ram[0][130] ) );
  DFFX1_HVT \ram_reg[0][129]  ( .D(n190), .CLK(clk), .Q(\ram[0][129] ) );
  DFFX1_HVT \ram_reg[0][128]  ( .D(n189), .CLK(clk), .Q(\ram[0][128] ) );
  DFFX1_HVT \ram_reg[0][127]  ( .D(n188), .CLK(clk), .Q(\ram[0][127] ) );
  DFFX1_HVT \ram_reg[0][126]  ( .D(n187), .CLK(clk), .Q(\ram[0][126] ) );
  DFFX1_HVT \ram_reg[0][125]  ( .D(n186), .CLK(clk), .Q(\ram[0][125] ) );
  DFFX1_HVT \ram_reg[0][124]  ( .D(n185), .CLK(clk), .Q(\ram[0][124] ), .QN(
        n4561) );
  DFFX1_HVT \ram_reg[0][123]  ( .D(n184), .CLK(clk), .Q(\ram[0][123] ) );
  DFFX1_HVT \ram_reg[0][122]  ( .D(n183), .CLK(clk), .Q(\ram[0][122] ) );
  DFFX1_HVT \ram_reg[0][121]  ( .D(n182), .CLK(clk), .Q(\ram[0][121] ) );
  DFFX1_HVT \ram_reg[0][120]  ( .D(n181), .CLK(clk), .Q(\ram[0][120] ) );
  DFFX1_HVT \ram_reg[0][119]  ( .D(n180), .CLK(clk), .Q(\ram[0][119] ) );
  DFFX1_HVT \ram_reg[0][118]  ( .D(n179), .CLK(clk), .Q(\ram[0][118] ) );
  DFFX1_HVT \ram_reg[0][117]  ( .D(n178), .CLK(clk), .Q(\ram[0][117] ) );
  DFFX1_HVT \ram_reg[0][116]  ( .D(n177), .CLK(clk), .Q(\ram[0][116] ) );
  DFFX1_HVT \ram_reg[0][115]  ( .D(n176), .CLK(clk), .Q(\ram[0][115] ) );
  DFFX1_HVT \ram_reg[0][114]  ( .D(n175), .CLK(clk), .Q(\ram[0][114] ) );
  DFFX1_HVT \ram_reg[0][113]  ( .D(n174), .CLK(clk), .Q(\ram[0][113] ) );
  DFFX1_HVT \ram_reg[0][112]  ( .D(n173), .CLK(clk), .Q(\ram[0][112] ), .QN(
        n5840) );
  DFFX1_HVT \ram_reg[0][111]  ( .D(n172), .CLK(clk), .Q(\ram[0][111] ) );
  DFFX1_HVT \ram_reg[0][110]  ( .D(n171), .CLK(clk), .Q(\ram[0][110] ) );
  DFFX1_HVT \ram_reg[0][109]  ( .D(n170), .CLK(clk), .Q(\ram[0][109] ) );
  DFFX1_HVT \ram_reg[0][108]  ( .D(n169), .CLK(clk), .Q(\ram[0][108] ) );
  DFFX1_HVT \ram_reg[0][107]  ( .D(n168), .CLK(clk), .Q(\ram[0][107] ) );
  DFFX1_HVT \ram_reg[0][106]  ( .D(n167), .CLK(clk), .Q(\ram[0][106] ) );
  DFFX1_HVT \ram_reg[0][105]  ( .D(n166), .CLK(clk), .Q(\ram[0][105] ) );
  DFFX1_HVT \ram_reg[0][104]  ( .D(n165), .CLK(clk), .Q(\ram[0][104] ) );
  DFFX1_HVT \ram_reg[0][103]  ( .D(n164), .CLK(clk), .Q(\ram[0][103] ), .QN(
        n4341) );
  DFFX1_HVT \ram_reg[0][102]  ( .D(n163), .CLK(clk), .Q(\ram[0][102] ) );
  DFFX1_HVT \ram_reg[0][101]  ( .D(n162), .CLK(clk), .Q(\ram[0][101] ) );
  DFFX1_HVT \ram_reg[0][100]  ( .D(n161), .CLK(clk), .Q(\ram[0][100] ) );
  DFFX1_HVT \ram_reg[0][99]  ( .D(n160), .CLK(clk), .Q(\ram[0][99] ) );
  DFFX1_HVT \ram_reg[0][98]  ( .D(n159), .CLK(clk), .Q(\ram[0][98] ) );
  DFFX1_HVT \ram_reg[0][97]  ( .D(n158), .CLK(clk), .Q(\ram[0][97] ) );
  DFFX1_HVT \ram_reg[0][96]  ( .D(n157), .CLK(clk), .Q(\ram[0][96] ) );
  DFFX1_HVT \ram_reg[0][95]  ( .D(n156), .CLK(clk), .Q(\ram[0][95] ) );
  DFFX1_HVT \ram_reg[0][94]  ( .D(n155), .CLK(clk), .Q(\ram[0][94] ) );
  DFFX1_HVT \ram_reg[0][93]  ( .D(n154), .CLK(clk), .Q(\ram[0][93] ) );
  DFFX1_HVT \ram_reg[0][92]  ( .D(n153), .CLK(clk), .Q(\ram[0][92] ) );
  DFFX1_HVT \ram_reg[0][91]  ( .D(n152), .CLK(clk), .Q(\ram[0][91] ) );
  DFFX1_HVT \ram_reg[0][90]  ( .D(n151), .CLK(clk), .Q(\ram[0][90] ) );
  DFFX1_HVT \ram_reg[0][89]  ( .D(n150), .CLK(clk), .Q(\ram[0][89] ) );
  DFFX1_HVT \ram_reg[0][88]  ( .D(n149), .CLK(clk), .Q(\ram[0][88] ) );
  DFFX1_HVT \ram_reg[0][87]  ( .D(n148), .CLK(clk), .Q(\ram[0][87] ) );
  DFFX1_HVT \ram_reg[0][86]  ( .D(n147), .CLK(clk), .Q(\ram[0][86] ) );
  DFFX1_HVT \ram_reg[0][85]  ( .D(n146), .CLK(clk), .Q(\ram[0][85] ) );
  DFFX1_HVT \ram_reg[0][84]  ( .D(n145), .CLK(clk), .Q(\ram[0][84] ) );
  DFFX1_HVT \ram_reg[0][83]  ( .D(n144), .CLK(clk), .Q(\ram[0][83] ) );
  DFFX1_HVT \ram_reg[0][82]  ( .D(n143), .CLK(clk), .Q(\ram[0][82] ) );
  DFFX1_HVT \ram_reg[0][81]  ( .D(n142), .CLK(clk), .Q(\ram[0][81] ) );
  DFFX1_HVT \ram_reg[0][80]  ( .D(n141), .CLK(clk), .Q(\ram[0][80] ) );
  DFFX1_HVT \ram_reg[0][79]  ( .D(n140), .CLK(clk), .Q(\ram[0][79] ) );
  DFFX1_HVT \ram_reg[0][78]  ( .D(n139), .CLK(clk), .Q(\ram[0][78] ) );
  DFFX1_HVT \ram_reg[0][77]  ( .D(n138), .CLK(clk), .Q(\ram[0][77] ) );
  DFFX1_HVT \ram_reg[0][76]  ( .D(n137), .CLK(clk), .Q(\ram[0][76] ) );
  DFFX1_HVT \ram_reg[0][75]  ( .D(n136), .CLK(clk), .Q(\ram[0][75] ) );
  DFFX1_HVT \ram_reg[0][74]  ( .D(n135), .CLK(clk), .Q(\ram[0][74] ) );
  DFFX1_HVT \ram_reg[0][73]  ( .D(n134), .CLK(clk), .Q(\ram[0][73] ) );
  DFFX1_HVT \ram_reg[0][72]  ( .D(n133), .CLK(clk), .Q(\ram[0][72] ) );
  DFFX1_HVT \ram_reg[0][71]  ( .D(n132), .CLK(clk), .Q(\ram[0][71] ) );
  DFFX1_HVT \ram_reg[0][70]  ( .D(n131), .CLK(clk), .Q(\ram[0][70] ) );
  DFFX1_HVT \ram_reg[0][69]  ( .D(n130), .CLK(clk), .Q(\ram[0][69] ) );
  DFFX1_HVT \ram_reg[0][68]  ( .D(n129), .CLK(clk), .Q(\ram[0][68] ) );
  DFFX1_HVT \ram_reg[0][67]  ( .D(n128), .CLK(clk), .Q(\ram[0][67] ) );
  DFFX1_HVT \ram_reg[0][66]  ( .D(n127), .CLK(clk), .Q(\ram[0][66] ) );
  DFFX1_HVT \ram_reg[0][65]  ( .D(n126), .CLK(clk), .Q(\ram[0][65] ) );
  DFFX1_HVT \ram_reg[0][64]  ( .D(n125), .CLK(clk), .Q(\ram[0][64] ) );
  DFFX1_HVT \ram_reg[0][63]  ( .D(n124), .CLK(clk), .Q(\ram[0][63] ) );
  DFFX1_HVT \ram_reg[0][62]  ( .D(n123), .CLK(clk), .Q(\ram[0][62] ) );
  DFFX1_HVT \ram_reg[0][61]  ( .D(n122), .CLK(clk), .Q(\ram[0][61] ) );
  DFFX1_HVT \ram_reg[0][60]  ( .D(n121), .CLK(clk), .Q(\ram[0][60] ) );
  DFFX1_HVT \ram_reg[0][59]  ( .D(n120), .CLK(clk), .Q(\ram[0][59] ) );
  DFFX1_HVT \ram_reg[0][58]  ( .D(n119), .CLK(clk), .Q(\ram[0][58] ) );
  DFFX1_HVT \ram_reg[0][57]  ( .D(n118), .CLK(clk), .Q(\ram[0][57] ) );
  DFFX1_HVT \ram_reg[0][56]  ( .D(n117), .CLK(clk), .Q(\ram[0][56] ) );
  DFFX1_HVT \ram_reg[0][55]  ( .D(n116), .CLK(clk), .Q(\ram[0][55] ) );
  DFFX1_HVT \ram_reg[0][54]  ( .D(n115), .CLK(clk), .Q(\ram[0][54] ) );
  DFFX1_HVT \ram_reg[0][53]  ( .D(n114), .CLK(clk), .Q(\ram[0][53] ) );
  DFFX1_HVT \ram_reg[0][52]  ( .D(n113), .CLK(clk), .Q(\ram[0][52] ) );
  DFFX1_HVT \ram_reg[0][51]  ( .D(n112), .CLK(clk), .Q(\ram[0][51] ) );
  DFFX1_HVT \ram_reg[0][50]  ( .D(n111), .CLK(clk), .Q(\ram[0][50] ), .QN(
        n4443) );
  DFFX1_HVT \ram_reg[0][49]  ( .D(n110), .CLK(clk), .Q(\ram[0][49] ) );
  DFFX1_HVT \ram_reg[0][48]  ( .D(n109), .CLK(clk), .Q(\ram[0][48] ) );
  DFFX1_HVT \ram_reg[0][47]  ( .D(n108), .CLK(clk), .Q(\ram[0][47] ) );
  DFFX1_HVT \ram_reg[0][46]  ( .D(n107), .CLK(clk), .Q(\ram[0][46] ) );
  DFFX1_HVT \ram_reg[0][45]  ( .D(n106), .CLK(clk), .Q(\ram[0][45] ) );
  DFFX1_HVT \ram_reg[0][44]  ( .D(n105), .CLK(clk), .Q(\ram[0][44] ) );
  DFFX1_HVT \ram_reg[0][43]  ( .D(n104), .CLK(clk), .Q(\ram[0][43] ) );
  DFFX1_HVT \ram_reg[0][42]  ( .D(n103), .CLK(clk), .Q(\ram[0][42] ) );
  DFFX1_HVT \ram_reg[0][41]  ( .D(n102), .CLK(clk), .Q(\ram[0][41] ) );
  DFFX1_HVT \ram_reg[0][40]  ( .D(n101), .CLK(clk), .Q(\ram[0][40] ) );
  DFFX1_HVT \ram_reg[0][39]  ( .D(n100), .CLK(clk), .Q(\ram[0][39] ) );
  DFFX1_HVT \ram_reg[0][38]  ( .D(n99), .CLK(clk), .Q(\ram[0][38] ) );
  DFFX1_HVT \ram_reg[0][37]  ( .D(n98), .CLK(clk), .Q(\ram[0][37] ) );
  DFFX1_HVT \ram_reg[0][36]  ( .D(n97), .CLK(clk), .Q(\ram[0][36] ) );
  DFFX1_HVT \ram_reg[0][35]  ( .D(n96), .CLK(clk), .Q(\ram[0][35] ) );
  DFFX1_HVT \ram_reg[0][34]  ( .D(n95), .CLK(clk), .Q(\ram[0][34] ) );
  DFFX1_HVT \ram_reg[0][33]  ( .D(n94), .CLK(clk), .Q(\ram[0][33] ) );
  DFFX1_HVT \ram_reg[0][32]  ( .D(n93), .CLK(clk), .Q(\ram[0][32] ) );
  DFFX1_HVT \ram_reg[0][31]  ( .D(n92), .CLK(clk), .Q(\ram[0][31] ) );
  DFFX1_HVT \ram_reg[0][30]  ( .D(n91), .CLK(clk), .Q(\ram[0][30] ) );
  DFFX1_HVT \ram_reg[0][29]  ( .D(n90), .CLK(clk), .Q(\ram[0][29] ) );
  DFFX1_HVT \ram_reg[0][28]  ( .D(n89), .CLK(clk), .Q(\ram[0][28] ) );
  DFFX1_HVT \ram_reg[0][27]  ( .D(n88), .CLK(clk), .Q(\ram[0][27] ) );
  DFFX1_HVT \ram_reg[0][26]  ( .D(n87), .CLK(clk), .Q(\ram[0][26] ) );
  DFFX1_HVT \ram_reg[0][25]  ( .D(n86), .CLK(clk), .Q(\ram[0][25] ) );
  DFFX1_HVT \ram_reg[0][24]  ( .D(n85), .CLK(clk), .Q(\ram[0][24] ) );
  DFFX1_HVT \ram_reg[0][23]  ( .D(n84), .CLK(clk), .Q(\ram[0][23] ) );
  DFFX1_HVT \ram_reg[0][22]  ( .D(n83), .CLK(clk), .Q(\ram[0][22] ) );
  DFFX1_HVT \ram_reg[0][21]  ( .D(n82), .CLK(clk), .Q(\ram[0][21] ) );
  DFFX1_HVT \ram_reg[0][20]  ( .D(n81), .CLK(clk), .Q(\ram[0][20] ), .QN(n4483) );
  DFFX1_HVT \ram_reg[0][19]  ( .D(n80), .CLK(clk), .Q(\ram[0][19] ) );
  DFFX1_HVT \ram_reg[0][18]  ( .D(n79), .CLK(clk), .Q(\ram[0][18] ) );
  DFFX1_HVT \ram_reg[0][17]  ( .D(n78), .CLK(clk), .Q(\ram[0][17] ) );
  DFFX1_HVT \ram_reg[0][16]  ( .D(n77), .CLK(clk), .Q(\ram[0][16] ) );
  DFFX1_HVT \ram_reg[0][15]  ( .D(n76), .CLK(clk), .Q(\ram[0][15] ) );
  DFFX1_HVT \ram_reg[0][14]  ( .D(n75), .CLK(clk), .Q(\ram[0][14] ) );
  DFFX1_HVT \ram_reg[0][13]  ( .D(n74), .CLK(clk), .Q(\ram[0][13] ) );
  DFFX1_HVT \ram_reg[0][12]  ( .D(n73), .CLK(clk), .Q(\ram[0][12] ) );
  DFFX1_HVT \ram_reg[0][11]  ( .D(n72), .CLK(clk), .Q(\ram[0][11] ) );
  DFFX1_HVT \ram_reg[0][10]  ( .D(n71), .CLK(clk), .Q(\ram[0][10] ) );
  DFFX1_HVT \ram_reg[0][9]  ( .D(n70), .CLK(clk), .Q(\ram[0][9] ) );
  DFFX1_HVT \ram_reg[0][8]  ( .D(n69), .CLK(clk), .Q(\ram[0][8] ) );
  DFFX1_HVT \ram_reg[0][7]  ( .D(n68), .CLK(clk), .Q(\ram[0][7] ), .QN(n6404)
         );
  DFFX1_HVT \ram_reg[0][6]  ( .D(n67), .CLK(clk), .Q(\ram[0][6] ) );
  DFFX1_HVT \ram_reg[0][5]  ( .D(n66), .CLK(clk), .Q(\ram[0][5] ) );
  DFFX1_HVT \ram_reg[0][4]  ( .D(n65), .CLK(clk), .Q(\ram[0][4] ) );
  DFFX1_HVT \ram_reg[0][3]  ( .D(n64), .CLK(clk), .Q(\ram[0][3] ) );
  DFFX1_HVT \ram_reg[0][2]  ( .D(n63), .CLK(clk), .Q(\ram[0][2] ), .QN(n4484)
         );
  DFFX1_HVT \ram_reg[0][1]  ( .D(n62), .CLK(clk), .Q(\ram[0][1] ) );
  DFFX1_HVT \ram_reg[0][0]  ( .D(n61), .CLK(clk), .Q(\ram[0][0] ) );
  AO22X1_HVT U7 ( .A1(\ram[0][0] ), .A2(n6670), .A3(n9307), .A4(n6497), .Y(n61) );
  AO22X1_HVT U8 ( .A1(\ram[0][1] ), .A2(n6707), .A3(n9310), .A4(n6539), .Y(n62) );
  AO22X1_HVT U10 ( .A1(\ram[0][3] ), .A2(n6705), .A3(n9316), .A4(n6536), .Y(
        n64) );
  AO22X1_HVT U11 ( .A1(\ram[0][4] ), .A2(n6704), .A3(n9320), .A4(n6535), .Y(
        n65) );
  AO22X1_HVT U12 ( .A1(\ram[0][5] ), .A2(n6702), .A3(n9323), .A4(n6533), .Y(
        n66) );
  AO22X1_HVT U13 ( .A1(\ram[0][6] ), .A2(n6701), .A3(n9326), .A4(n6532), .Y(
        n67) );
  AO22X1_HVT U14 ( .A1(\ram[0][7] ), .A2(n6672), .A3(n9329), .A4(n6529), .Y(
        n68) );
  AO22X1_HVT U15 ( .A1(\ram[0][8] ), .A2(n6698), .A3(n9332), .A4(n6528), .Y(
        n69) );
  AO22X1_HVT U16 ( .A1(\ram[0][9] ), .A2(n6696), .A3(n9335), .A4(n6526), .Y(
        n70) );
  AO22X1_HVT U17 ( .A1(\ram[0][10] ), .A2(n4385), .A3(n9338), .A4(n6525), .Y(
        n71) );
  AO22X1_HVT U18 ( .A1(\ram[0][11] ), .A2(n6695), .A3(n9341), .A4(n6524), .Y(
        n72) );
  AO22X1_HVT U19 ( .A1(\ram[0][12] ), .A2(n6694), .A3(n9345), .A4(n6523), .Y(
        n73) );
  AO22X1_HVT U20 ( .A1(\ram[0][13] ), .A2(n4385), .A3(n9348), .A4(n6521), .Y(
        n74) );
  AO22X1_HVT U21 ( .A1(\ram[0][14] ), .A2(n6692), .A3(n9351), .A4(n6520), .Y(
        n75) );
  AO22X1_HVT U22 ( .A1(\ram[0][15] ), .A2(n6690), .A3(n9354), .A4(n6518), .Y(
        n76) );
  AO22X1_HVT U23 ( .A1(\ram[0][16] ), .A2(n10368), .A3(n9357), .A4(n6517), .Y(
        n77) );
  AO22X1_HVT U24 ( .A1(\ram[0][17] ), .A2(n6689), .A3(n9360), .A4(n4272), .Y(
        n78) );
  AO22X1_HVT U25 ( .A1(\ram[0][18] ), .A2(n6667), .A3(n9363), .A4(n6513), .Y(
        n79) );
  AO22X1_HVT U26 ( .A1(\ram[0][19] ), .A2(n6685), .A3(n9366), .A4(n6523), .Y(
        n80) );
  AO22X1_HVT U28 ( .A1(\ram[0][21] ), .A2(n6682), .A3(n9371), .A4(n10354), .Y(
        n82) );
  AO22X1_HVT U29 ( .A1(\ram[0][22] ), .A2(n6681), .A3(n9374), .A4(n6509), .Y(
        n83) );
  AO22X1_HVT U30 ( .A1(\ram[0][23] ), .A2(n6677), .A3(n9377), .A4(n6544), .Y(
        n84) );
  AO22X1_HVT U31 ( .A1(\ram[0][24] ), .A2(n6676), .A3(n9380), .A4(n6502), .Y(
        n85) );
  AO22X1_HVT U32 ( .A1(\ram[0][25] ), .A2(n6673), .A3(n9383), .A4(n6501), .Y(
        n86) );
  AO22X1_HVT U33 ( .A1(\ram[0][26] ), .A2(n6699), .A3(n9386), .A4(n6500), .Y(
        n87) );
  AO22X1_HVT U34 ( .A1(\ram[0][27] ), .A2(n6670), .A3(n9389), .A4(n6497), .Y(
        n88) );
  AO22X1_HVT U35 ( .A1(\ram[0][28] ), .A2(n6669), .A3(n9392), .A4(n6496), .Y(
        n89) );
  AO22X1_HVT U36 ( .A1(\ram[0][29] ), .A2(n4398), .A3(n9395), .A4(n6495), .Y(
        n90) );
  AO22X1_HVT U37 ( .A1(\ram[0][30] ), .A2(n6688), .A3(n9398), .A4(n6494), .Y(
        n91) );
  AO22X1_HVT U38 ( .A1(\ram[0][31] ), .A2(n6731), .A3(n9401), .A4(n6490), .Y(
        n92) );
  AO22X1_HVT U39 ( .A1(\ram[0][32] ), .A2(n6730), .A3(n9404), .A4(n6489), .Y(
        n93) );
  AO22X1_HVT U40 ( .A1(\ram[0][33] ), .A2(n6729), .A3(n9407), .A4(n6487), .Y(
        n94) );
  AO22X1_HVT U41 ( .A1(\ram[0][34] ), .A2(n6729), .A3(n9410), .A4(n6487), .Y(
        n95) );
  AO22X1_HVT U42 ( .A1(\ram[0][35] ), .A2(n10368), .A3(n9413), .A4(n6525), .Y(
        n96) );
  AO22X1_HVT U43 ( .A1(\ram[0][36] ), .A2(n6695), .A3(n9416), .A4(n6524), .Y(
        n97) );
  AO22X1_HVT U44 ( .A1(\ram[0][37] ), .A2(n6694), .A3(n9419), .A4(n6523), .Y(
        n98) );
  AO22X1_HVT U45 ( .A1(\ram[0][38] ), .A2(n4385), .A3(n9422), .A4(n6521), .Y(
        n99) );
  AO22X1_HVT U46 ( .A1(\ram[0][39] ), .A2(n6692), .A3(data[39]), .A4(n6520), 
        .Y(n100) );
  AO22X1_HVT U47 ( .A1(\ram[0][40] ), .A2(n6690), .A3(n9428), .A4(n6518), .Y(
        n101) );
  AO22X1_HVT U48 ( .A1(\ram[0][41] ), .A2(n10368), .A3(n9431), .A4(n6517), .Y(
        n102) );
  AO22X1_HVT U49 ( .A1(\ram[0][42] ), .A2(n6689), .A3(n9434), .A4(n6547), .Y(
        n103) );
  AO22X1_HVT U50 ( .A1(\ram[0][43] ), .A2(n6725), .A3(n9437), .A4(n6548), .Y(
        n104) );
  AO22X1_HVT U51 ( .A1(\ram[0][44] ), .A2(n6723), .A3(n9440), .A4(n10357), .Y(
        n105) );
  AO22X1_HVT U52 ( .A1(\ram[0][45] ), .A2(n6722), .A3(n9443), .A4(n4272), .Y(
        n106) );
  AO22X1_HVT U53 ( .A1(\ram[0][46] ), .A2(n6721), .A3(n9446), .A4(n6546), .Y(
        n107) );
  AO22X1_HVT U54 ( .A1(\ram[0][47] ), .A2(n4198), .A3(n9449), .A4(n6507), .Y(
        n108) );
  AO22X1_HVT U55 ( .A1(\ram[0][48] ), .A2(n6720), .A3(n9452), .A4(n6487), .Y(
        n109) );
  AO22X1_HVT U56 ( .A1(\ram[0][49] ), .A2(n6717), .A3(n9455), .A4(n6507), .Y(
        n110) );
  AO22X1_HVT U58 ( .A1(\ram[0][51] ), .A2(n6715), .A3(n9461), .A4(n6495), .Y(
        n112) );
  AO22X1_HVT U59 ( .A1(\ram[0][52] ), .A2(n4198), .A3(n9464), .A4(n6506), .Y(
        n113) );
  AO22X1_HVT U60 ( .A1(\ram[0][53] ), .A2(n6711), .A3(n9467), .A4(n6493), .Y(
        n114) );
  AO22X1_HVT U61 ( .A1(\ram[0][54] ), .A2(n6710), .A3(n9470), .A4(n4397), .Y(
        n115) );
  AO22X1_HVT U62 ( .A1(\ram[0][55] ), .A2(n6707), .A3(n9473), .A4(n6549), .Y(
        n116) );
  AO22X1_HVT U63 ( .A1(\ram[0][56] ), .A2(n6706), .A3(n9476), .A4(n6548), .Y(
        n117) );
  AO22X1_HVT U64 ( .A1(\ram[0][57] ), .A2(n6705), .A3(n9479), .A4(n4396), .Y(
        n118) );
  AO22X1_HVT U65 ( .A1(\ram[0][58] ), .A2(n6704), .A3(n9482), .A4(n6514), .Y(
        n119) );
  AO22X1_HVT U66 ( .A1(\ram[0][59] ), .A2(n6702), .A3(n9485), .A4(n6546), .Y(
        n120) );
  AO22X1_HVT U67 ( .A1(\ram[0][60] ), .A2(n6728), .A3(n9488), .A4(n6545), .Y(
        n121) );
  AO22X1_HVT U68 ( .A1(\ram[0][61] ), .A2(n6714), .A3(n9491), .A4(n6544), .Y(
        n122) );
  AO22X1_HVT U69 ( .A1(\ram[0][62] ), .A2(n6669), .A3(n9494), .A4(n10356), .Y(
        n123) );
  AO22X1_HVT U70 ( .A1(\ram[0][63] ), .A2(n6672), .A3(n9497), .A4(n6543), .Y(
        n124) );
  AO22X1_HVT U71 ( .A1(\ram[0][64] ), .A2(n6684), .A3(n9500), .A4(n6542), .Y(
        n125) );
  AO22X1_HVT U72 ( .A1(\ram[0][65] ), .A2(n6666), .A3(n9503), .A4(n6541), .Y(
        n126) );
  AO22X1_HVT U73 ( .A1(\ram[0][66] ), .A2(n6679), .A3(n9506), .A4(n6540), .Y(
        n127) );
  AO22X1_HVT U74 ( .A1(\ram[0][67] ), .A2(n6726), .A3(n9509), .A4(n6539), .Y(
        n128) );
  AO22X1_HVT U75 ( .A1(\ram[0][68] ), .A2(n6725), .A3(n9512), .A4(n6538), .Y(
        n129) );
  AO22X1_HVT U76 ( .A1(\ram[0][69] ), .A2(n6723), .A3(n9515), .A4(n6536), .Y(
        n130) );
  AO22X1_HVT U77 ( .A1(\ram[0][70] ), .A2(n6722), .A3(n9518), .A4(n6535), .Y(
        n131) );
  AO22X1_HVT U78 ( .A1(\ram[0][71] ), .A2(n6721), .A3(n9521), .A4(n6533), .Y(
        n132) );
  AO22X1_HVT U79 ( .A1(\ram[0][72] ), .A2(n6701), .A3(n9524), .A4(n6532), .Y(
        n133) );
  AO22X1_HVT U80 ( .A1(\ram[0][73] ), .A2(n4398), .A3(n9527), .A4(n6529), .Y(
        n134) );
  AO22X1_HVT U81 ( .A1(\ram[0][74] ), .A2(n6698), .A3(n9530), .A4(n6528), .Y(
        n135) );
  AO22X1_HVT U82 ( .A1(\ram[0][75] ), .A2(n6696), .A3(n9533), .A4(n6526), .Y(
        n136) );
  AO22X1_HVT U83 ( .A1(\ram[0][76] ), .A2(n4343), .A3(n9536), .A4(n6525), .Y(
        n137) );
  AO22X1_HVT U84 ( .A1(\ram[0][77] ), .A2(n6695), .A3(n9539), .A4(n6524), .Y(
        n138) );
  AO22X1_HVT U85 ( .A1(\ram[0][78] ), .A2(n6694), .A3(n9542), .A4(n6523), .Y(
        n139) );
  AO22X1_HVT U86 ( .A1(\ram[0][79] ), .A2(n4385), .A3(n9545), .A4(n6521), .Y(
        n140) );
  AO22X1_HVT U87 ( .A1(\ram[0][80] ), .A2(n6692), .A3(n9548), .A4(n6520), .Y(
        n141) );
  AO22X1_HVT U88 ( .A1(\ram[0][81] ), .A2(n6690), .A3(n9551), .A4(n6518), .Y(
        n142) );
  AO22X1_HVT U89 ( .A1(\ram[0][82] ), .A2(n10370), .A3(n9554), .A4(n6517), .Y(
        n143) );
  AO22X1_HVT U90 ( .A1(\ram[0][83] ), .A2(n6689), .A3(n9557), .A4(n6514), .Y(
        n144) );
  AO22X1_HVT U91 ( .A1(\ram[0][84] ), .A2(n6688), .A3(n9560), .A4(n6513), .Y(
        n145) );
  AO22X1_HVT U92 ( .A1(\ram[0][85] ), .A2(n6685), .A3(n9563), .A4(n6526), .Y(
        n146) );
  AO22X1_HVT U93 ( .A1(\ram[0][86] ), .A2(n6667), .A3(n9566), .A4(n6513), .Y(
        n147) );
  AO22X1_HVT U94 ( .A1(\ram[0][87] ), .A2(n6685), .A3(n9569), .A4(n6525), .Y(
        n148) );
  AO22X1_HVT U95 ( .A1(\ram[0][88] ), .A2(n6678), .A3(n9572), .A4(n6510), .Y(
        n149) );
  AO22X1_HVT U96 ( .A1(\ram[0][89] ), .A2(n6682), .A3(n9575), .A4(n10356), .Y(
        n150) );
  AO22X1_HVT U97 ( .A1(\ram[0][90] ), .A2(n6681), .A3(n9578), .A4(n6509), .Y(
        n151) );
  AO22X1_HVT U98 ( .A1(\ram[0][91] ), .A2(n6677), .A3(n9581), .A4(n6503), .Y(
        n152) );
  AO22X1_HVT U99 ( .A1(\ram[0][92] ), .A2(n6676), .A3(n9584), .A4(n6502), .Y(
        n153) );
  AO22X1_HVT U100 ( .A1(\ram[0][93] ), .A2(n6673), .A3(n9587), .A4(n6501), .Y(
        n154) );
  AO22X1_HVT U101 ( .A1(\ram[0][94] ), .A2(n6720), .A3(n9590), .A4(n6545), .Y(
        n155) );
  AO22X1_HVT U102 ( .A1(\ram[0][95] ), .A2(n6717), .A3(n9593), .A4(n6503), .Y(
        n156) );
  AO22X1_HVT U103 ( .A1(\ram[0][96] ), .A2(n6716), .A3(n9596), .A4(n10356), 
        .Y(n157) );
  AO22X1_HVT U104 ( .A1(\ram[0][97] ), .A2(n6715), .A3(n9599), .A4(n6543), .Y(
        n158) );
  AO22X1_HVT U105 ( .A1(\ram[0][98] ), .A2(n4344), .A3(n9602), .A4(n6506), .Y(
        n159) );
  AO22X1_HVT U106 ( .A1(\ram[0][99] ), .A2(n4344), .A3(n9605), .A4(n6510), .Y(
        n160) );
  AO22X1_HVT U107 ( .A1(\ram[0][100] ), .A2(n6682), .A3(n9608), .A4(n10358), 
        .Y(n161) );
  AO22X1_HVT U108 ( .A1(\ram[0][101] ), .A2(n6667), .A3(n9611), .A4(n6494), 
        .Y(n162) );
  AO22X1_HVT U109 ( .A1(\ram[0][102] ), .A2(n6731), .A3(n9614), .A4(n6490), 
        .Y(n163) );
  AO22X1_HVT U111 ( .A1(\ram[0][104] ), .A2(n6677), .A3(n9620), .A4(n6503), 
        .Y(n165) );
  AO22X1_HVT U112 ( .A1(\ram[0][105] ), .A2(n6676), .A3(n9623), .A4(n6502), 
        .Y(n166) );
  AO22X1_HVT U113 ( .A1(\ram[0][106] ), .A2(n6673), .A3(n9626), .A4(n6501), 
        .Y(n167) );
  AO22X1_HVT U114 ( .A1(\ram[0][107] ), .A2(n6672), .A3(n9629), .A4(n6500), 
        .Y(n168) );
  AO22X1_HVT U115 ( .A1(\ram[0][108] ), .A2(n6670), .A3(n9632), .A4(n6497), 
        .Y(n169) );
  AO22X1_HVT U116 ( .A1(\ram[0][109] ), .A2(n6669), .A3(n9635), .A4(n6496), 
        .Y(n170) );
  AO22X1_HVT U117 ( .A1(\ram[0][110] ), .A2(n6699), .A3(n9638), .A4(n6495), 
        .Y(n171) );
  AO22X1_HVT U118 ( .A1(\ram[0][111] ), .A2(n6688), .A3(n9641), .A4(n6494), 
        .Y(n172) );
  AO22X1_HVT U119 ( .A1(\ram[0][112] ), .A2(n6731), .A3(n9644), .A4(n6490), 
        .Y(n173) );
  AO22X1_HVT U120 ( .A1(\ram[0][113] ), .A2(n6730), .A3(n9647), .A4(n6489), 
        .Y(n174) );
  AO22X1_HVT U121 ( .A1(\ram[0][114] ), .A2(n6729), .A3(n9650), .A4(n6486), 
        .Y(n175) );
  AO22X1_HVT U122 ( .A1(\ram[0][115] ), .A2(n6726), .A3(n9653), .A4(n6486), 
        .Y(n176) );
  AO22X1_HVT U123 ( .A1(\ram[0][116] ), .A2(n6728), .A3(n9656), .A4(n6486), 
        .Y(n177) );
  AO22X1_HVT U124 ( .A1(\ram[0][117] ), .A2(n4342), .A3(n9659), .A4(n6507), 
        .Y(n178) );
  AO22X1_HVT U125 ( .A1(\ram[0][118] ), .A2(n6678), .A3(n9662), .A4(n6506), 
        .Y(n179) );
  AO22X1_HVT U126 ( .A1(\ram[0][119] ), .A2(n6666), .A3(n9665), .A4(n6493), 
        .Y(n180) );
  AO22X1_HVT U127 ( .A1(\ram[0][120] ), .A2(n4342), .A3(n9668), .A4(n6488), 
        .Y(n181) );
  AO22X1_HVT U128 ( .A1(\ram[0][121] ), .A2(n6726), .A3(n9671), .A4(n6488), 
        .Y(n182) );
  AO22X1_HVT U129 ( .A1(\ram[0][122] ), .A2(n6725), .A3(n9674), .A4(n4330), 
        .Y(n183) );
  AO22X1_HVT U130 ( .A1(\ram[0][123] ), .A2(n6723), .A3(n9677), .A4(n6507), 
        .Y(n184) );
  AO22X1_HVT U132 ( .A1(\ram[0][125] ), .A2(n6721), .A3(n9683), .A4(n6493), 
        .Y(n186) );
  AO22X1_HVT U133 ( .A1(\ram[0][126] ), .A2(n6720), .A3(n9686), .A4(n4397), 
        .Y(n187) );
  AO22X1_HVT U134 ( .A1(\ram[0][127] ), .A2(n6717), .A3(n9689), .A4(n6549), 
        .Y(n188) );
  AO22X1_HVT U135 ( .A1(\ram[0][128] ), .A2(n6716), .A3(n9692), .A4(n6486), 
        .Y(n189) );
  AO22X1_HVT U136 ( .A1(\ram[0][129] ), .A2(n6715), .A3(n9695), .A4(n6488), 
        .Y(n190) );
  AO22X1_HVT U137 ( .A1(\ram[0][130] ), .A2(n6679), .A3(n9698), .A4(n6507), 
        .Y(n191) );
  AO22X1_HVT U138 ( .A1(\ram[0][131] ), .A2(n6711), .A3(n9701), .A4(n6506), 
        .Y(n192) );
  AO22X1_HVT U139 ( .A1(\ram[0][132] ), .A2(n6710), .A3(n9704), .A4(n6493), 
        .Y(n193) );
  AO22X1_HVT U140 ( .A1(\ram[0][133] ), .A2(n6707), .A3(n9707), .A4(n4396), 
        .Y(n194) );
  AO22X1_HVT U141 ( .A1(\ram[0][134] ), .A2(n6706), .A3(n9710), .A4(n6549), 
        .Y(n195) );
  AO22X1_HVT U142 ( .A1(\ram[0][135] ), .A2(n6705), .A3(n9713), .A4(n6548), 
        .Y(n196) );
  AO22X1_HVT U143 ( .A1(\ram[0][136] ), .A2(n6704), .A3(n9716), .A4(n6538), 
        .Y(n197) );
  AO22X1_HVT U144 ( .A1(\ram[0][137] ), .A2(n6668), .A3(n9719), .A4(n6536), 
        .Y(n198) );
  AO22X1_HVT U145 ( .A1(\ram[0][138] ), .A2(n6670), .A3(n9722), .A4(n6535), 
        .Y(n199) );
  AO22X1_HVT U146 ( .A1(\ram[0][139] ), .A2(n6669), .A3(n9725), .A4(n6533), 
        .Y(n200) );
  AO22X1_HVT U147 ( .A1(\ram[0][140] ), .A2(n6668), .A3(n9729), .A4(n4397), 
        .Y(n201) );
  AO22X1_HVT U148 ( .A1(\ram[0][141] ), .A2(n6667), .A3(n9732), .A4(n6548), 
        .Y(n202) );
  AO22X1_HVT U149 ( .A1(\ram[0][142] ), .A2(n6731), .A3(data[142]), .A4(n4397), 
        .Y(n203) );
  AO22X1_HVT U150 ( .A1(\ram[0][143] ), .A2(n6730), .A3(n9738), .A4(n4330), 
        .Y(n204) );
  AO22X1_HVT U152 ( .A1(\ram[0][145] ), .A2(n6714), .A3(n9745), .A4(n4272), 
        .Y(n206) );
  AO22X1_HVT U153 ( .A1(\ram[0][146] ), .A2(n6711), .A3(n9748), .A4(n6546), 
        .Y(n207) );
  AO22X1_HVT U154 ( .A1(\ram[0][147] ), .A2(n6710), .A3(n9751), .A4(n6545), 
        .Y(n208) );
  AO22X1_HVT U155 ( .A1(\ram[0][148] ), .A2(n6707), .A3(n9755), .A4(n4273), 
        .Y(n209) );
  AO22X1_HVT U156 ( .A1(\ram[0][149] ), .A2(n6666), .A3(n9758), .A4(n6506), 
        .Y(n210) );
  AO22X1_HVT U157 ( .A1(\ram[0][150] ), .A2(n6702), .A3(n9761), .A4(n6543), 
        .Y(n211) );
  AO22X1_HVT U158 ( .A1(\ram[0][151] ), .A2(n6701), .A3(n9764), .A4(n6542), 
        .Y(n212) );
  AO22X1_HVT U159 ( .A1(\ram[0][152] ), .A2(n6730), .A3(n9767), .A4(n6541), 
        .Y(n213) );
  AO22X1_HVT U160 ( .A1(\ram[0][153] ), .A2(n6729), .A3(n9770), .A4(n6540), 
        .Y(n214) );
  AO22X1_HVT U161 ( .A1(\ram[0][154] ), .A2(n6672), .A3(n9773), .A4(n6539), 
        .Y(n215) );
  AO22X1_HVT U162 ( .A1(\ram[0][155] ), .A2(n6698), .A3(n9776), .A4(n6538), 
        .Y(n216) );
  AO22X1_HVT U163 ( .A1(\ram[0][156] ), .A2(n6696), .A3(n9780), .A4(n6536), 
        .Y(n217) );
  AO22X1_HVT U164 ( .A1(\ram[0][157] ), .A2(n10368), .A3(n9783), .A4(n6535), 
        .Y(n218) );
  AO22X1_HVT U165 ( .A1(\ram[0][158] ), .A2(n6695), .A3(n9786), .A4(n6533), 
        .Y(n219) );
  AO22X1_HVT U166 ( .A1(\ram[0][159] ), .A2(n6694), .A3(n9789), .A4(n6532), 
        .Y(n220) );
  AO22X1_HVT U167 ( .A1(\ram[0][160] ), .A2(n4385), .A3(n9793), .A4(n6529), 
        .Y(n221) );
  AO22X1_HVT U168 ( .A1(\ram[0][161] ), .A2(n6692), .A3(n9796), .A4(n6528), 
        .Y(n222) );
  AO22X1_HVT U169 ( .A1(\ram[0][162] ), .A2(n6690), .A3(n9799), .A4(n6526), 
        .Y(n223) );
  AO22X1_HVT U170 ( .A1(\ram[0][163] ), .A2(n10368), .A3(n9802), .A4(n6525), 
        .Y(n224) );
  AO22X1_HVT U171 ( .A1(\ram[0][164] ), .A2(n6689), .A3(n9805), .A4(n6524), 
        .Y(n225) );
  AO22X1_HVT U172 ( .A1(\ram[0][165] ), .A2(n6688), .A3(n9808), .A4(n6523), 
        .Y(n226) );
  AO22X1_HVT U173 ( .A1(\ram[0][166] ), .A2(n6685), .A3(n9811), .A4(n6521), 
        .Y(n227) );
  AO22X1_HVT U174 ( .A1(\ram[0][167] ), .A2(n6684), .A3(n9814), .A4(n6520), 
        .Y(n228) );
  AO22X1_HVT U175 ( .A1(\ram[0][168] ), .A2(n6682), .A3(n9817), .A4(n6547), 
        .Y(n229) );
  AO22X1_HVT U176 ( .A1(\ram[0][169] ), .A2(n6681), .A3(n9820), .A4(n6546), 
        .Y(n230) );
  AO22X1_HVT U177 ( .A1(\ram[0][170] ), .A2(n6677), .A3(n9823), .A4(n6545), 
        .Y(n231) );
  AO22X1_HVT U178 ( .A1(\ram[0][171] ), .A2(n6676), .A3(n9826), .A4(n4273), 
        .Y(n232) );
  AO22X1_HVT U179 ( .A1(\ram[0][172] ), .A2(n6673), .A3(n9830), .A4(n10356), 
        .Y(n233) );
  AO22X1_HVT U180 ( .A1(\ram[0][173] ), .A2(n6699), .A3(n9833), .A4(n6543), 
        .Y(n234) );
  AO22X1_HVT U181 ( .A1(\ram[0][174] ), .A2(n6670), .A3(n9836), .A4(n6542), 
        .Y(n235) );
  AO22X1_HVT U182 ( .A1(\ram[0][175] ), .A2(n6669), .A3(n9839), .A4(n6532), 
        .Y(n236) );
  AO22X1_HVT U183 ( .A1(\ram[0][176] ), .A2(n4398), .A3(n9843), .A4(n6529), 
        .Y(n237) );
  AO22X1_HVT U184 ( .A1(\ram[0][177] ), .A2(n6667), .A3(n9846), .A4(n6528), 
        .Y(n238) );
  AO22X1_HVT U185 ( .A1(\ram[0][178] ), .A2(n6731), .A3(n9849), .A4(n6526), 
        .Y(n239) );
  AO22X1_HVT U186 ( .A1(\ram[0][179] ), .A2(n6730), .A3(n9852), .A4(n6549), 
        .Y(n240) );
  AO22X1_HVT U187 ( .A1(\ram[0][180] ), .A2(n6729), .A3(n9856), .A4(n6518), 
        .Y(n241) );
  AO22X1_HVT U188 ( .A1(\ram[0][181] ), .A2(n6731), .A3(n9859), .A4(n6517), 
        .Y(n242) );
  AO22X1_HVT U189 ( .A1(\ram[0][182] ), .A2(n6728), .A3(n9862), .A4(n6547), 
        .Y(n243) );
  AO22X1_HVT U190 ( .A1(\ram[0][183] ), .A2(n4198), .A3(n9865), .A4(n6544), 
        .Y(n244) );
  AO22X1_HVT U191 ( .A1(\ram[0][184] ), .A2(n4344), .A3(n9869), .A4(n6521), 
        .Y(n245) );
  AO22X1_HVT U192 ( .A1(\ram[0][185] ), .A2(n6666), .A3(n9872), .A4(n6510), 
        .Y(n246) );
  AO22X1_HVT U193 ( .A1(\ram[0][186] ), .A2(n6679), .A3(n9875), .A4(n10357), 
        .Y(n247) );
  AO22X1_HVT U194 ( .A1(\ram[0][187] ), .A2(n6726), .A3(n9878), .A4(n6509), 
        .Y(n248) );
  AO22X1_HVT U195 ( .A1(\ram[0][188] ), .A2(n6730), .A3(n9881), .A4(n6544), 
        .Y(n249) );
  AO22X1_HVT U196 ( .A1(\ram[0][189] ), .A2(n6728), .A3(n9884), .A4(n6502), 
        .Y(n250) );
  AO22X1_HVT U197 ( .A1(\ram[0][190] ), .A2(n6714), .A3(n9887), .A4(n6501), 
        .Y(n251) );
  AO22X1_HVT U198 ( .A1(\ram[0][191] ), .A2(n6684), .A3(n9890), .A4(n4396), 
        .Y(n252) );
  AO22X1_HVT U199 ( .A1(\ram[0][192] ), .A2(n6666), .A3(n9894), .A4(n4396), 
        .Y(n253) );
  AO22X1_HVT U200 ( .A1(\ram[0][193] ), .A2(n6714), .A3(n9897), .A4(n6549), 
        .Y(n254) );
  AO22X1_HVT U201 ( .A1(\ram[0][194] ), .A2(n6726), .A3(n9900), .A4(n6548), 
        .Y(n255) );
  AO22X1_HVT U202 ( .A1(\ram[0][195] ), .A2(n6725), .A3(n9903), .A4(n10357), 
        .Y(n256) );
  AO22X1_HVT U203 ( .A1(\ram[0][196] ), .A2(n6706), .A3(n9907), .A4(n6547), 
        .Y(n257) );
  AO22X1_HVT U204 ( .A1(\ram[0][197] ), .A2(n6705), .A3(n9910), .A4(n6546), 
        .Y(n258) );
  AO22X1_HVT U205 ( .A1(\ram[0][198] ), .A2(n6704), .A3(n9913), .A4(n6545), 
        .Y(n259) );
  AO22X1_HVT U206 ( .A1(\ram[0][199] ), .A2(n6702), .A3(n9916), .A4(n6503), 
        .Y(n260) );
  AO22X1_HVT U207 ( .A1(\ram[0][200] ), .A2(n4198), .A3(n9920), .A4(n10356), 
        .Y(n261) );
  AO22X1_HVT U208 ( .A1(\ram[0][201] ), .A2(n6725), .A3(n9923), .A4(n6543), 
        .Y(n262) );
  AO22X1_HVT U209 ( .A1(\ram[0][202] ), .A2(n6723), .A3(n9926), .A4(n6542), 
        .Y(n263) );
  AO22X1_HVT U210 ( .A1(\ram[0][203] ), .A2(n6729), .A3(n9929), .A4(n6541), 
        .Y(n264) );
  AO22X1_HVT U211 ( .A1(\ram[0][204] ), .A2(n6728), .A3(n9932), .A4(n6540), 
        .Y(n265) );
  AO22X1_HVT U212 ( .A1(\ram[0][205] ), .A2(n6722), .A3(n9935), .A4(n6539), 
        .Y(n266) );
  AO22X1_HVT U213 ( .A1(\ram[0][206] ), .A2(n6721), .A3(n9938), .A4(n6538), 
        .Y(n267) );
  AO22X1_HVT U214 ( .A1(\ram[0][207] ), .A2(n6720), .A3(n9941), .A4(n6536), 
        .Y(n268) );
  AO22X1_HVT U215 ( .A1(\ram[0][208] ), .A2(n6717), .A3(n9945), .A4(n6535), 
        .Y(n269) );
  AO22X1_HVT U216 ( .A1(\ram[0][209] ), .A2(n6716), .A3(n9948), .A4(n6500), 
        .Y(n270) );
  AO22X1_HVT U217 ( .A1(\ram[0][210] ), .A2(n6715), .A3(n9951), .A4(n6497), 
        .Y(n271) );
  AO22X1_HVT U218 ( .A1(\ram[0][211] ), .A2(n6679), .A3(n9954), .A4(n6496), 
        .Y(n272) );
  AO22X1_HVT U219 ( .A1(\ram[0][212] ), .A2(n6711), .A3(n9957), .A4(n6495), 
        .Y(n273) );
  AO22X1_HVT U220 ( .A1(\ram[0][213] ), .A2(n6710), .A3(n9960), .A4(n6494), 
        .Y(n274) );
  AO22X1_HVT U221 ( .A1(\ram[0][214] ), .A2(n6707), .A3(n9963), .A4(n6490), 
        .Y(n275) );
  AO22X1_HVT U222 ( .A1(\ram[0][215] ), .A2(n6706), .A3(n9966), .A4(n6489), 
        .Y(n276) );
  AO22X1_HVT U223 ( .A1(\ram[0][216] ), .A2(n6705), .A3(n9969), .A4(n4330), 
        .Y(n277) );
  AO22X1_HVT U224 ( .A1(\ram[0][217] ), .A2(n6704), .A3(n9972), .A4(n6542), 
        .Y(n278) );
  AO22X1_HVT U225 ( .A1(\ram[0][218] ), .A2(n6702), .A3(n9975), .A4(n6541), 
        .Y(n279) );
  AO22X1_HVT U226 ( .A1(\ram[0][219] ), .A2(n6701), .A3(n9978), .A4(n6540), 
        .Y(n280) );
  AO22X1_HVT U227 ( .A1(\ram[0][220] ), .A2(n6668), .A3(n9982), .A4(n6539), 
        .Y(n281) );
  AO22X1_HVT U228 ( .A1(\ram[0][221] ), .A2(n6698), .A3(n9985), .A4(n6514), 
        .Y(n282) );
  AO22X1_HVT U229 ( .A1(\ram[0][222] ), .A2(n6696), .A3(n9988), .A4(n6533), 
        .Y(n283) );
  AO22X1_HVT U230 ( .A1(\ram[0][223] ), .A2(n4343), .A3(n9991), .A4(n6532), 
        .Y(n284) );
  AO22X1_HVT U231 ( .A1(\ram[0][224] ), .A2(n6695), .A3(n9994), .A4(n6489), 
        .Y(n285) );
  AO22X1_HVT U232 ( .A1(\ram[0][225] ), .A2(n6694), .A3(n9997), .A4(n6488), 
        .Y(n286) );
  AO22X1_HVT U233 ( .A1(\ram[0][226] ), .A2(n4385), .A3(n10000), .A4(n6529), 
        .Y(n287) );
  AO22X1_HVT U234 ( .A1(\ram[0][227] ), .A2(n6678), .A3(n10003), .A4(n6528), 
        .Y(n288) );
  AO22X1_HVT U235 ( .A1(\ram[0][228] ), .A2(n6690), .A3(n10006), .A4(n6526), 
        .Y(n289) );
  AO22X1_HVT U236 ( .A1(\ram[0][229] ), .A2(n10371), .A3(n10009), .A4(n6525), 
        .Y(n290) );
  AO22X1_HVT U237 ( .A1(\ram[0][230] ), .A2(n6689), .A3(n10012), .A4(n6524), 
        .Y(n291) );
  AO22X1_HVT U238 ( .A1(\ram[0][231] ), .A2(n6688), .A3(n10015), .A4(n6523), 
        .Y(n292) );
  AO22X1_HVT U239 ( .A1(\ram[0][232] ), .A2(n6685), .A3(n10019), .A4(n6521), 
        .Y(n293) );
  AO22X1_HVT U240 ( .A1(\ram[0][233] ), .A2(n6678), .A3(n10022), .A4(n6520), 
        .Y(n294) );
  AO22X1_HVT U241 ( .A1(\ram[0][234] ), .A2(n6682), .A3(n10025), .A4(n6518), 
        .Y(n295) );
  AO22X1_HVT U242 ( .A1(\ram[0][235] ), .A2(n6681), .A3(n10028), .A4(n6517), 
        .Y(n296) );
  AO22X1_HVT U243 ( .A1(\ram[0][236] ), .A2(n6677), .A3(n10031), .A4(n6514), 
        .Y(n297) );
  AO22X1_HVT U244 ( .A1(\ram[0][237] ), .A2(n6676), .A3(n10034), .A4(n6513), 
        .Y(n298) );
  AO22X1_HVT U245 ( .A1(\ram[0][238] ), .A2(n6673), .A3(n10037), .A4(n6524), 
        .Y(n299) );
  AO22X1_HVT U246 ( .A1(\ram[0][239] ), .A2(n6723), .A3(n10040), .A4(n6510), 
        .Y(n300) );
  AO22X1_HVT U247 ( .A1(\ram[0][240] ), .A2(n6722), .A3(n10044), .A4(n10359), 
        .Y(n301) );
  AO22X1_HVT U248 ( .A1(\ram[0][241] ), .A2(n6721), .A3(n10047), .A4(n6509), 
        .Y(n302) );
  AO22X1_HVT U249 ( .A1(\ram[0][242] ), .A2(n6720), .A3(n10050), .A4(n4273), 
        .Y(n303) );
  AO22X1_HVT U250 ( .A1(\ram[0][243] ), .A2(n6717), .A3(n10053), .A4(n6502), 
        .Y(n304) );
  AO22X1_HVT U251 ( .A1(\ram[0][244] ), .A2(n6716), .A3(n10056), .A4(n6501), 
        .Y(n305) );
  AO22X1_HVT U252 ( .A1(\ram[0][245] ), .A2(n6715), .A3(n10059), .A4(n6500), 
        .Y(n306) );
  AO22X1_HVT U253 ( .A1(\ram[0][246] ), .A2(n4342), .A3(n10062), .A4(n6497), 
        .Y(n307) );
  AO22X1_HVT U254 ( .A1(\ram[0][247] ), .A2(n6701), .A3(n10065), .A4(n6496), 
        .Y(n308) );
  AO22X1_HVT U255 ( .A1(\ram[0][248] ), .A2(n6699), .A3(n10069), .A4(n6495), 
        .Y(n309) );
  AO22X1_HVT U256 ( .A1(\ram[0][249] ), .A2(n6698), .A3(n10072), .A4(n6494), 
        .Y(n310) );
  AO22X1_HVT U257 ( .A1(\ram[0][250] ), .A2(n6696), .A3(n10075), .A4(n6490), 
        .Y(n311) );
  AO22X1_HVT U258 ( .A1(\ram[0][251] ), .A2(n6726), .A3(n10078), .A4(n6489), 
        .Y(n312) );
  AO22X1_HVT U259 ( .A1(\ram[0][252] ), .A2(n6728), .A3(n10082), .A4(n6487), 
        .Y(n313) );
  AO22X1_HVT U260 ( .A1(\ram[0][253] ), .A2(n6711), .A3(n10085), .A4(n6541), 
        .Y(n314) );
  AO22X1_HVT U261 ( .A1(\ram[0][254] ), .A2(n6710), .A3(n10088), .A4(n6540), 
        .Y(n315) );
  AO22X1_HVT U262 ( .A1(\ram[0][255] ), .A2(n6668), .A3(n10091), .A4(n6500), 
        .Y(n316) );
  AND2X1_HVT U265 ( .A1(n5822), .A2(n5130), .Y(n7) );
  AO22X1_HVT U266 ( .A1(\ram[1][0] ), .A2(n4615), .A3(n6831), .A4(n9306), .Y(
        n317) );
  AO22X1_HVT U267 ( .A1(\ram[1][1] ), .A2(n7047), .A3(n6830), .A4(n9309), .Y(
        n318) );
  AO22X1_HVT U268 ( .A1(\ram[1][2] ), .A2(n7048), .A3(n6829), .A4(data[2]), 
        .Y(n319) );
  AO22X1_HVT U269 ( .A1(\ram[1][3] ), .A2(n7050), .A3(n6890), .A4(n9315), .Y(
        n320) );
  AO22X1_HVT U270 ( .A1(\ram[1][4] ), .A2(n7042), .A3(n6889), .A4(n9319), .Y(
        n321) );
  AO22X1_HVT U271 ( .A1(\ram[1][5] ), .A2(n4869), .A3(n6888), .A4(n9322), .Y(
        n322) );
  AO22X1_HVT U272 ( .A1(\ram[1][6] ), .A2(n4593), .A3(n6887), .A4(n9325), .Y(
        n323) );
  AO22X1_HVT U273 ( .A1(\ram[1][7] ), .A2(n4419), .A3(n6886), .A4(n9328), .Y(
        n324) );
  AO22X1_HVT U274 ( .A1(\ram[1][8] ), .A2(n7032), .A3(n6828), .A4(n9331), .Y(
        n325) );
  AO22X1_HVT U275 ( .A1(\ram[1][9] ), .A2(n7031), .A3(n6827), .A4(n9334), .Y(
        n326) );
  AO22X1_HVT U277 ( .A1(\ram[1][11] ), .A2(n7029), .A3(n6885), .A4(n9340), .Y(
        n328) );
  AO22X1_HVT U278 ( .A1(\ram[1][12] ), .A2(n7032), .A3(n10342), .A4(n9344), 
        .Y(n329) );
  AO22X1_HVT U279 ( .A1(\ram[1][13] ), .A2(n7031), .A3(n6884), .A4(n9347), .Y(
        n330) );
  AO22X1_HVT U280 ( .A1(\ram[1][14] ), .A2(n7030), .A3(n6883), .A4(n9350), .Y(
        n331) );
  AO22X1_HVT U281 ( .A1(\ram[1][15] ), .A2(n4574), .A3(n6858), .A4(n9353), .Y(
        n332) );
  AO22X1_HVT U282 ( .A1(\ram[1][16] ), .A2(n7069), .A3(n6880), .A4(n9356), .Y(
        n333) );
  AO22X1_HVT U283 ( .A1(\ram[1][17] ), .A2(n4444), .A3(n6878), .A4(n9359), .Y(
        n334) );
  AO22X1_HVT U285 ( .A1(\ram[1][19] ), .A2(n7069), .A3(n6874), .A4(n9365), .Y(
        n336) );
  AO22X1_HVT U286 ( .A1(\ram[1][20] ), .A2(n4723), .A3(n6873), .A4(n9368), .Y(
        n337) );
  AO22X1_HVT U287 ( .A1(\ram[1][21] ), .A2(n4785), .A3(n6872), .A4(n9370), .Y(
        n338) );
  AO22X1_HVT U288 ( .A1(\ram[1][22] ), .A2(n7062), .A3(n4323), .A4(n9373), .Y(
        n339) );
  AO22X1_HVT U289 ( .A1(\ram[1][23] ), .A2(n4722), .A3(n6869), .A4(n9376), .Y(
        n340) );
  AO22X1_HVT U290 ( .A1(\ram[1][24] ), .A2(n7078), .A3(n6868), .A4(n9379), .Y(
        n341) );
  AO22X1_HVT U291 ( .A1(\ram[1][25] ), .A2(n7078), .A3(n6841), .A4(n9382), .Y(
        n342) );
  AO22X1_HVT U292 ( .A1(\ram[1][26] ), .A2(n7075), .A3(n6866), .A4(n9385), .Y(
        n343) );
  AO22X1_HVT U293 ( .A1(\ram[1][27] ), .A2(n7077), .A3(n6865), .A4(n9388), .Y(
        n344) );
  AO22X1_HVT U294 ( .A1(\ram[1][28] ), .A2(n7069), .A3(n6864), .A4(n9391), .Y(
        n345) );
  AO22X1_HVT U296 ( .A1(\ram[1][30] ), .A2(n7069), .A3(n6860), .A4(n9397), .Y(
        n347) );
  AO22X1_HVT U297 ( .A1(\ram[1][31] ), .A2(n7069), .A3(n6859), .A4(n9400), .Y(
        n348) );
  AO22X1_HVT U298 ( .A1(\ram[1][32] ), .A2(n7041), .A3(n6858), .A4(n9403), .Y(
        n349) );
  AO22X1_HVT U299 ( .A1(\ram[1][33] ), .A2(n7033), .A3(n4440), .A4(n9406), .Y(
        n350) );
  AO22X1_HVT U300 ( .A1(\ram[1][34] ), .A2(n4593), .A3(n6856), .A4(n9409), .Y(
        n351) );
  AO22X1_HVT U301 ( .A1(\ram[1][35] ), .A2(n7040), .A3(n6841), .A4(n9412), .Y(
        n352) );
  AO22X1_HVT U302 ( .A1(\ram[1][36] ), .A2(n4869), .A3(n6869), .A4(n9415), .Y(
        n353) );
  AO22X1_HVT U303 ( .A1(\ram[1][37] ), .A2(n7041), .A3(n6868), .A4(n9418), .Y(
        n354) );
  AO22X1_HVT U304 ( .A1(\ram[1][38] ), .A2(n4868), .A3(n6867), .A4(n9421), .Y(
        n355) );
  AO22X1_HVT U305 ( .A1(\ram[1][39] ), .A2(n7040), .A3(n6866), .A4(n9424), .Y(
        n356) );
  AO22X1_HVT U307 ( .A1(\ram[1][41] ), .A2(n4871), .A3(n6864), .A4(n9430), .Y(
        n358) );
  AO22X1_HVT U309 ( .A1(\ram[1][43] ), .A2(n7033), .A3(n6853), .A4(n9436), .Y(
        n360) );
  AO22X1_HVT U310 ( .A1(\ram[1][44] ), .A2(n4444), .A3(n6850), .A4(n9439), .Y(
        n361) );
  AO22X1_HVT U312 ( .A1(\ram[1][46] ), .A2(n7046), .A3(n6847), .A4(n9445), .Y(
        n363) );
  AO22X1_HVT U313 ( .A1(\ram[1][47] ), .A2(n7036), .A3(n6828), .A4(n9448), .Y(
        n364) );
  AO22X1_HVT U315 ( .A1(\ram[1][49] ), .A2(n7051), .A3(n6874), .A4(n9454), .Y(
        n366) );
  AO22X1_HVT U316 ( .A1(\ram[1][50] ), .A2(n7048), .A3(n6873), .A4(n9457), .Y(
        n367) );
  AO22X1_HVT U317 ( .A1(\ram[1][51] ), .A2(n7045), .A3(n6872), .A4(n9460), .Y(
        n368) );
  AO22X1_HVT U318 ( .A1(\ram[1][52] ), .A2(n7046), .A3(n6867), .A4(n9463), .Y(
        n369) );
  AO22X1_HVT U319 ( .A1(\ram[1][53] ), .A2(n7062), .A3(n6869), .A4(n9466), .Y(
        n370) );
  AO22X1_HVT U320 ( .A1(\ram[1][54] ), .A2(n7059), .A3(n6845), .A4(n9469), .Y(
        n371) );
  AO22X1_HVT U321 ( .A1(\ram[1][55] ), .A2(n7060), .A3(n6829), .A4(n9472), .Y(
        n372) );
  AO22X1_HVT U322 ( .A1(\ram[1][56] ), .A2(n4785), .A3(n6844), .A4(n9475), .Y(
        n373) );
  AO22X1_HVT U323 ( .A1(\ram[1][57] ), .A2(n7057), .A3(n6885), .A4(n9478), .Y(
        n374) );
  AO22X1_HVT U324 ( .A1(\ram[1][58] ), .A2(n7057), .A3(n10342), .A4(n9481), 
        .Y(n375) );
  AO22X1_HVT U325 ( .A1(\ram[1][59] ), .A2(n7057), .A3(n6884), .A4(n9484), .Y(
        n376) );
  AO22X1_HVT U326 ( .A1(\ram[1][60] ), .A2(n7035), .A3(n6859), .A4(n9487), .Y(
        n377) );
  AO22X1_HVT U327 ( .A1(\ram[1][61] ), .A2(n4870), .A3(n6858), .A4(n9490), .Y(
        n378) );
  AO22X1_HVT U328 ( .A1(\ram[1][62] ), .A2(n4863), .A3(n6841), .A4(n9493), .Y(
        n379) );
  AO22X1_HVT U329 ( .A1(\ram[1][63] ), .A2(n7045), .A3(n6854), .A4(n9496), .Y(
        n380) );
  AO22X1_HVT U330 ( .A1(\ram[1][64] ), .A2(n7061), .A3(n6853), .A4(n9499), .Y(
        n381) );
  AO22X1_HVT U331 ( .A1(\ram[1][65] ), .A2(n7059), .A3(n6850), .A4(n9502), .Y(
        n382) );
  AO22X1_HVT U332 ( .A1(\ram[1][66] ), .A2(n7059), .A3(n6849), .A4(n9505), .Y(
        n383) );
  AO22X1_HVT U333 ( .A1(\ram[1][67] ), .A2(n7061), .A3(n6847), .A4(n9508), .Y(
        n384) );
  AO22X1_HVT U334 ( .A1(\ram[1][68] ), .A2(n7061), .A3(n6857), .A4(n9511), .Y(
        n385) );
  AO22X1_HVT U335 ( .A1(\ram[1][69] ), .A2(n7062), .A3(n6846), .A4(n9514), .Y(
        n386) );
  AO22X1_HVT U336 ( .A1(\ram[1][70] ), .A2(n4723), .A3(n6845), .A4(n9517), .Y(
        n387) );
  AO22X1_HVT U337 ( .A1(\ram[1][71] ), .A2(n7060), .A3(n6828), .A4(n9520), .Y(
        n388) );
  AO22X1_HVT U338 ( .A1(\ram[1][72] ), .A2(n4722), .A3(n6844), .A4(n9523), .Y(
        n389) );
  AO22X1_HVT U339 ( .A1(\ram[1][73] ), .A2(n4785), .A3(n6885), .A4(n9526), .Y(
        n390) );
  AO22X1_HVT U340 ( .A1(\ram[1][74] ), .A2(n4722), .A3(n6840), .A4(n9529), .Y(
        n391) );
  AO22X1_HVT U341 ( .A1(\ram[1][75] ), .A2(n7061), .A3(n6839), .A4(n9532), .Y(
        n392) );
  AO22X1_HVT U342 ( .A1(\ram[1][76] ), .A2(n4871), .A3(n6836), .A4(n9535), .Y(
        n393) );
  AO22X1_HVT U343 ( .A1(\ram[1][77] ), .A2(n7047), .A3(n6835), .A4(n9538), .Y(
        n394) );
  AO22X1_HVT U344 ( .A1(\ram[1][78] ), .A2(n7048), .A3(n6832), .A4(n9541), .Y(
        n395) );
  AO22X1_HVT U345 ( .A1(\ram[1][79] ), .A2(n7050), .A3(n6835), .A4(n9544), .Y(
        n396) );
  AO22X1_HVT U346 ( .A1(\ram[1][80] ), .A2(n7033), .A3(n6830), .A4(n9547), .Y(
        n397) );
  AO22X1_HVT U347 ( .A1(\ram[1][81] ), .A2(n7041), .A3(n6829), .A4(n9550), .Y(
        n398) );
  AO22X1_HVT U348 ( .A1(\ram[1][82] ), .A2(n4593), .A3(n6890), .A4(n9553), .Y(
        n399) );
  AO22X1_HVT U349 ( .A1(\ram[1][83] ), .A2(n4419), .A3(n6889), .A4(n9556), .Y(
        n400) );
  AO22X1_HVT U350 ( .A1(\ram[1][84] ), .A2(n7045), .A3(n6888), .A4(n9559), .Y(
        n401) );
  AO22X1_HVT U351 ( .A1(\ram[1][85] ), .A2(n7047), .A3(n6887), .A4(n9562), .Y(
        n402) );
  AO22X1_HVT U353 ( .A1(\ram[1][87] ), .A2(n7042), .A3(n6828), .A4(n9568), .Y(
        n404) );
  AO22X1_HVT U355 ( .A1(\ram[1][89] ), .A2(n7065), .A3(n6842), .A4(n9574), .Y(
        n406) );
  AO22X1_HVT U356 ( .A1(\ram[1][90] ), .A2(n7066), .A3(n6871), .A4(n9577), .Y(
        n407) );
  AO22X1_HVT U357 ( .A1(\ram[1][91] ), .A2(n7066), .A3(n6854), .A4(n9580), .Y(
        n408) );
  AO22X1_HVT U358 ( .A1(\ram[1][92] ), .A2(n7067), .A3(n6853), .A4(n9583), .Y(
        n409) );
  AO22X1_HVT U359 ( .A1(\ram[1][93] ), .A2(n7067), .A3(n6850), .A4(n9586), .Y(
        n410) );
  AO22X1_HVT U360 ( .A1(\ram[1][94] ), .A2(n7067), .A3(n6849), .A4(n9589), .Y(
        n411) );
  AO22X1_HVT U361 ( .A1(\ram[1][95] ), .A2(n7065), .A3(n6847), .A4(n9592), .Y(
        n412) );
  AO22X1_HVT U362 ( .A1(\ram[1][96] ), .A2(n7046), .A3(n6827), .A4(n9595), .Y(
        n413) );
  AO22X1_HVT U363 ( .A1(\ram[1][97] ), .A2(n4673), .A3(n6846), .A4(n9598), .Y(
        n414) );
  AO22X1_HVT U364 ( .A1(\ram[1][98] ), .A2(n7034), .A3(n6860), .A4(n9601), .Y(
        n415) );
  AO22X1_HVT U365 ( .A1(\ram[1][99] ), .A2(n4869), .A3(n6859), .A4(n9604), .Y(
        n416) );
  AO22X1_HVT U366 ( .A1(\ram[1][100] ), .A2(n7077), .A3(n6858), .A4(n9607), 
        .Y(n417) );
  AO22X1_HVT U367 ( .A1(\ram[1][101] ), .A2(n5483), .A3(n6857), .A4(n9610), 
        .Y(n418) );
  AO22X1_HVT U368 ( .A1(\ram[1][102] ), .A2(n7077), .A3(n6856), .A4(n9613), 
        .Y(n419) );
  AO22X1_HVT U369 ( .A1(\ram[1][103] ), .A2(n7075), .A3(n6840), .A4(n9616), 
        .Y(n420) );
  AO22X1_HVT U370 ( .A1(\ram[1][104] ), .A2(n7056), .A3(n6839), .A4(n9619), 
        .Y(n421) );
  AO22X1_HVT U371 ( .A1(\ram[1][105] ), .A2(n7055), .A3(n6836), .A4(n9622), 
        .Y(n422) );
  AO22X1_HVT U372 ( .A1(\ram[1][106] ), .A2(n4332), .A3(n10342), .A4(n9625), 
        .Y(n423) );
  AO22X1_HVT U373 ( .A1(\ram[1][107] ), .A2(n7056), .A3(n6846), .A4(n9628), 
        .Y(n424) );
  AO22X1_HVT U374 ( .A1(\ram[1][108] ), .A2(n7032), .A3(n6845), .A4(n9631), 
        .Y(n425) );
  AO22X1_HVT U375 ( .A1(\ram[1][109] ), .A2(n7031), .A3(n6827), .A4(n9634), 
        .Y(n426) );
  AO22X1_HVT U376 ( .A1(\ram[1][110] ), .A2(n7030), .A3(n6827), .A4(n9637), 
        .Y(n427) );
  AO22X1_HVT U377 ( .A1(\ram[1][111] ), .A2(n7029), .A3(n6856), .A4(n9640), 
        .Y(n428) );
  AO22X1_HVT U378 ( .A1(\ram[1][112] ), .A2(n7057), .A3(n6856), .A4(n9643), 
        .Y(n429) );
  AO22X1_HVT U379 ( .A1(\ram[1][113] ), .A2(n4332), .A3(n10342), .A4(n9646), 
        .Y(n430) );
  AO22X1_HVT U380 ( .A1(\ram[1][114] ), .A2(n7055), .A3(n6884), .A4(n9649), 
        .Y(n431) );
  AO22X1_HVT U381 ( .A1(\ram[1][115] ), .A2(n7056), .A3(n6883), .A4(n9652), 
        .Y(n432) );
  AO22X1_HVT U382 ( .A1(\ram[1][116] ), .A2(n4612), .A3(n6881), .A4(n9655), 
        .Y(n433) );
  AO22X1_HVT U383 ( .A1(\ram[1][117] ), .A2(n7058), .A3(n6880), .A4(n9658), 
        .Y(n434) );
  AO22X1_HVT U384 ( .A1(\ram[1][118] ), .A2(n7055), .A3(n6878), .A4(n9661), 
        .Y(n435) );
  AO22X1_HVT U385 ( .A1(\ram[1][119] ), .A2(n7058), .A3(n6877), .A4(n9664), 
        .Y(n436) );
  AO22X1_HVT U387 ( .A1(\ram[1][121] ), .A2(n7071), .A3(n6827), .A4(n9670), 
        .Y(n438) );
  AO22X1_HVT U389 ( .A1(\ram[1][123] ), .A2(n7072), .A3(n6867), .A4(n9676), 
        .Y(n440) );
  AO22X1_HVT U390 ( .A1(\ram[1][124] ), .A2(n4261), .A3(n6854), .A4(n9679), 
        .Y(n441) );
  AO22X1_HVT U391 ( .A1(\ram[1][125] ), .A2(n7081), .A3(n6853), .A4(n9682), 
        .Y(n442) );
  AO22X1_HVT U392 ( .A1(\ram[1][126] ), .A2(n7080), .A3(n6850), .A4(n9685), 
        .Y(n443) );
  AO22X1_HVT U393 ( .A1(\ram[1][127] ), .A2(n4259), .A3(n6849), .A4(n9688), 
        .Y(n444) );
  AO22X1_HVT U394 ( .A1(\ram[1][128] ), .A2(n4747), .A3(n6887), .A4(n9691), 
        .Y(n445) );
  AO22X1_HVT U395 ( .A1(\ram[1][129] ), .A2(n7075), .A3(n6886), .A4(n9694), 
        .Y(n446) );
  AO22X1_HVT U396 ( .A1(\ram[1][130] ), .A2(n5483), .A3(n6828), .A4(n9697), 
        .Y(n447) );
  AO22X1_HVT U397 ( .A1(\ram[1][131] ), .A2(n7076), .A3(n6827), .A4(n9700), 
        .Y(n448) );
  AO22X1_HVT U398 ( .A1(\ram[1][132] ), .A2(n7076), .A3(n6881), .A4(n9703), 
        .Y(n449) );
  AO22X1_HVT U399 ( .A1(\ram[1][133] ), .A2(n7078), .A3(n6880), .A4(n9706), 
        .Y(n450) );
  AO22X1_HVT U400 ( .A1(\ram[1][134] ), .A2(n7077), .A3(n6878), .A4(n9709), 
        .Y(n451) );
  AO22X1_HVT U401 ( .A1(\ram[1][135] ), .A2(n7078), .A3(n6877), .A4(n9712), 
        .Y(n452) );
  AO22X1_HVT U402 ( .A1(\ram[1][136] ), .A2(n7075), .A3(n6874), .A4(n9715), 
        .Y(n453) );
  AO22X1_HVT U403 ( .A1(\ram[1][137] ), .A2(n5483), .A3(n6873), .A4(n9718), 
        .Y(n454) );
  AO22X1_HVT U404 ( .A1(\ram[1][138] ), .A2(n7076), .A3(n6872), .A4(n9721), 
        .Y(n455) );
  AO22X1_HVT U405 ( .A1(\ram[1][139] ), .A2(n7075), .A3(n6871), .A4(n9724), 
        .Y(n456) );
  AO22X1_HVT U406 ( .A1(\ram[1][140] ), .A2(n7052), .A3(n6869), .A4(n9728), 
        .Y(n457) );
  AO22X1_HVT U407 ( .A1(\ram[1][141] ), .A2(n4871), .A3(n6868), .A4(n9731), 
        .Y(n458) );
  AO22X1_HVT U408 ( .A1(\ram[1][142] ), .A2(n4870), .A3(n4323), .A4(n9734), 
        .Y(n459) );
  AO22X1_HVT U409 ( .A1(\ram[1][143] ), .A2(n7050), .A3(n6866), .A4(n9737), 
        .Y(n460) );
  AO22X1_HVT U410 ( .A1(\ram[1][144] ), .A2(n7032), .A3(n6865), .A4(n9741), 
        .Y(n461) );
  AO22X1_HVT U411 ( .A1(\ram[1][145] ), .A2(n7031), .A3(n6864), .A4(n9744), 
        .Y(n462) );
  AO22X1_HVT U412 ( .A1(\ram[1][146] ), .A2(n7030), .A3(n6861), .A4(n9747), 
        .Y(n463) );
  AO22X1_HVT U413 ( .A1(\ram[1][147] ), .A2(n4574), .A3(n6860), .A4(n9750), 
        .Y(n464) );
  AO22X1_HVT U414 ( .A1(\ram[1][148] ), .A2(n4869), .A3(n6859), .A4(n9754), 
        .Y(n465) );
  AO22X1_HVT U415 ( .A1(\ram[1][149] ), .A2(n7042), .A3(n6831), .A4(n9757), 
        .Y(n466) );
  AO22X1_HVT U416 ( .A1(\ram[1][150] ), .A2(n4416), .A3(n6832), .A4(n9760), 
        .Y(n467) );
  AO22X1_HVT U417 ( .A1(\ram[1][151] ), .A2(n7040), .A3(n6835), .A4(n9763), 
        .Y(n468) );
  AO22X1_HVT U418 ( .A1(\ram[1][152] ), .A2(n4863), .A3(n6830), .A4(n9766), 
        .Y(n469) );
  AO22X1_HVT U419 ( .A1(\ram[1][153] ), .A2(n4615), .A3(n6829), .A4(n9769), 
        .Y(n470) );
  AO22X1_HVT U420 ( .A1(\ram[1][154] ), .A2(n7034), .A3(n6890), .A4(n9772), 
        .Y(n471) );
  AO22X1_HVT U421 ( .A1(\ram[1][155] ), .A2(n7033), .A3(n6889), .A4(n9775), 
        .Y(n472) );
  AO22X1_HVT U422 ( .A1(\ram[1][156] ), .A2(n7047), .A3(n6888), .A4(n9779), 
        .Y(n473) );
  AO22X1_HVT U423 ( .A1(\ram[1][157] ), .A2(n4870), .A3(n6844), .A4(n9782), 
        .Y(n474) );
  AO22X1_HVT U424 ( .A1(\ram[1][158] ), .A2(n7036), .A3(n6885), .A4(n9785), 
        .Y(n475) );
  AO22X1_HVT U425 ( .A1(\ram[1][159] ), .A2(n4863), .A3(n10342), .A4(n9788), 
        .Y(n476) );
  AO22X1_HVT U426 ( .A1(\ram[1][160] ), .A2(n4675), .A3(n6884), .A4(n9792), 
        .Y(n477) );
  AO22X1_HVT U427 ( .A1(\ram[1][161] ), .A2(n7051), .A3(n6842), .A4(n9795), 
        .Y(n478) );
  AO22X1_HVT U428 ( .A1(\ram[1][162] ), .A2(n7036), .A3(n6840), .A4(n9798), 
        .Y(n479) );
  AO22X1_HVT U429 ( .A1(\ram[1][163] ), .A2(n4863), .A3(n6839), .A4(n9801), 
        .Y(n480) );
  AO22X1_HVT U430 ( .A1(\ram[1][164] ), .A2(n5483), .A3(n6868), .A4(n9804), 
        .Y(n481) );
  AO22X1_HVT U431 ( .A1(\ram[1][165] ), .A2(n7077), .A3(n6867), .A4(n9807), 
        .Y(n482) );
  AO22X1_HVT U432 ( .A1(\ram[1][166] ), .A2(n7076), .A3(n6866), .A4(n9810), 
        .Y(n483) );
  AO22X1_HVT U433 ( .A1(\ram[1][167] ), .A2(n7076), .A3(n6865), .A4(n9813), 
        .Y(n484) );
  AO22X1_HVT U435 ( .A1(\ram[1][169] ), .A2(n7071), .A3(n6861), .A4(n9819), 
        .Y(n486) );
  AO22X1_HVT U436 ( .A1(\ram[1][170] ), .A2(n7070), .A3(n6860), .A4(n9822), 
        .Y(n487) );
  AO22X1_HVT U437 ( .A1(\ram[1][171] ), .A2(n7070), .A3(n6859), .A4(n9825), 
        .Y(n488) );
  AO22X1_HVT U438 ( .A1(\ram[1][172] ), .A2(n7068), .A3(n6881), .A4(n9829), 
        .Y(n489) );
  AO22X1_HVT U439 ( .A1(\ram[1][173] ), .A2(n5480), .A3(n4440), .A4(n9832), 
        .Y(n490) );
  AO22X1_HVT U440 ( .A1(\ram[1][174] ), .A2(n5480), .A3(n4440), .A4(n9835), 
        .Y(n491) );
  AO22X1_HVT U441 ( .A1(\ram[1][175] ), .A2(n7067), .A3(n6840), .A4(n9838), 
        .Y(n492) );
  AO22X1_HVT U442 ( .A1(\ram[1][176] ), .A2(n7072), .A3(n6881), .A4(n9842), 
        .Y(n493) );
  AO22X1_HVT U443 ( .A1(\ram[1][177] ), .A2(n7071), .A3(n6857), .A4(n9845), 
        .Y(n494) );
  AO22X1_HVT U444 ( .A1(\ram[1][178] ), .A2(n7072), .A3(n4440), .A4(n9848), 
        .Y(n495) );
  AO22X1_HVT U445 ( .A1(\ram[1][179] ), .A2(n7072), .A3(n6840), .A4(n9851), 
        .Y(n496) );
  AO22X1_HVT U446 ( .A1(\ram[1][180] ), .A2(n7070), .A3(n6839), .A4(n9855), 
        .Y(n497) );
  AO22X1_HVT U447 ( .A1(\ram[1][181] ), .A2(n7071), .A3(n6836), .A4(n9858), 
        .Y(n498) );
  AO22X1_HVT U448 ( .A1(\ram[1][182] ), .A2(n7070), .A3(n6831), .A4(n9861), 
        .Y(n499) );
  AO22X1_HVT U449 ( .A1(\ram[1][183] ), .A2(n7070), .A3(n6832), .A4(n9864), 
        .Y(n500) );
  AO22X1_HVT U450 ( .A1(\ram[1][184] ), .A2(n7041), .A3(n6835), .A4(n9868), 
        .Y(n501) );
  AO22X1_HVT U451 ( .A1(\ram[1][185] ), .A2(n7033), .A3(n6830), .A4(n9871), 
        .Y(n502) );
  AO22X1_HVT U452 ( .A1(\ram[1][186] ), .A2(n4416), .A3(n6829), .A4(n9874), 
        .Y(n503) );
  AO22X1_HVT U453 ( .A1(\ram[1][187] ), .A2(n4419), .A3(n6890), .A4(n9877), 
        .Y(n504) );
  AO22X1_HVT U454 ( .A1(\ram[1][188] ), .A2(n4261), .A3(n6889), .A4(n9880), 
        .Y(n505) );
  AO22X1_HVT U455 ( .A1(\ram[1][189] ), .A2(n7081), .A3(n6888), .A4(n9883), 
        .Y(n506) );
  AO22X1_HVT U456 ( .A1(\ram[1][190] ), .A2(n7080), .A3(n6887), .A4(n9886), 
        .Y(n507) );
  AO22X1_HVT U457 ( .A1(\ram[1][191] ), .A2(n7079), .A3(n6886), .A4(n9889), 
        .Y(n508) );
  AO22X1_HVT U458 ( .A1(\ram[1][192] ), .A2(n4673), .A3(n6842), .A4(n9893), 
        .Y(n509) );
  AO22X1_HVT U459 ( .A1(\ram[1][193] ), .A2(n4677), .A3(n4323), .A4(n9896), 
        .Y(n510) );
  AO22X1_HVT U460 ( .A1(\ram[1][194] ), .A2(n7035), .A3(n6854), .A4(n9899), 
        .Y(n511) );
  AO22X1_HVT U461 ( .A1(\ram[1][195] ), .A2(n7050), .A3(n6853), .A4(n9902), 
        .Y(n512) );
  AO22X1_HVT U462 ( .A1(\ram[1][196] ), .A2(n4871), .A3(n6883), .A4(n9906), 
        .Y(n513) );
  AO22X1_HVT U463 ( .A1(\ram[1][197] ), .A2(n7052), .A3(n6858), .A4(n9909), 
        .Y(n514) );
  AO22X1_HVT U464 ( .A1(\ram[1][198] ), .A2(n7051), .A3(n6880), .A4(n9912), 
        .Y(n515) );
  AO22X1_HVT U465 ( .A1(\ram[1][199] ), .A2(n7050), .A3(n6878), .A4(n9915), 
        .Y(n516) );
  AO22X1_HVT U466 ( .A1(\ram[1][200] ), .A2(n7051), .A3(n6871), .A4(n9919), 
        .Y(n517) );
  AO22X1_HVT U467 ( .A1(\ram[1][201] ), .A2(n4675), .A3(n6836), .A4(n9922), 
        .Y(n518) );
  AO22X1_HVT U468 ( .A1(\ram[1][202] ), .A2(n7045), .A3(n6835), .A4(n9925), 
        .Y(n519) );
  AO22X1_HVT U469 ( .A1(\ram[1][203] ), .A2(n7046), .A3(n6839), .A4(n9928), 
        .Y(n520) );
  AO22X1_HVT U470 ( .A1(\ram[1][204] ), .A2(n7062), .A3(n6836), .A4(n9931), 
        .Y(n521) );
  AO22X1_HVT U471 ( .A1(\ram[1][205] ), .A2(n4785), .A3(n6831), .A4(n9934), 
        .Y(n522) );
  AO22X1_HVT U472 ( .A1(\ram[1][206] ), .A2(n7060), .A3(n6832), .A4(n9937), 
        .Y(n523) );
  AO22X1_HVT U473 ( .A1(\ram[1][207] ), .A2(n4723), .A3(n6831), .A4(n9940), 
        .Y(n524) );
  AO22X1_HVT U474 ( .A1(\ram[1][208] ), .A2(n7082), .A3(n6830), .A4(n9944), 
        .Y(n525) );
  AO22X1_HVT U475 ( .A1(\ram[1][209] ), .A2(n7081), .A3(n6829), .A4(n9947), 
        .Y(n526) );
  AO22X1_HVT U476 ( .A1(\ram[1][210] ), .A2(n7080), .A3(n6890), .A4(n9950), 
        .Y(n527) );
  AO22X1_HVT U477 ( .A1(\ram[1][211] ), .A2(n4259), .A3(n6889), .A4(n9953), 
        .Y(n528) );
  AO22X1_HVT U478 ( .A1(\ram[1][212] ), .A2(n7082), .A3(n6888), .A4(n9956), 
        .Y(n529) );
  AO22X1_HVT U479 ( .A1(\ram[1][213] ), .A2(n7081), .A3(n6887), .A4(n9959), 
        .Y(n530) );
  AO22X1_HVT U480 ( .A1(\ram[1][214] ), .A2(n7080), .A3(n6886), .A4(n9962), 
        .Y(n531) );
  AO22X1_HVT U481 ( .A1(\ram[1][215] ), .A2(n7079), .A3(n6847), .A4(n9965), 
        .Y(n532) );
  AO22X1_HVT U482 ( .A1(\ram[1][216] ), .A2(n7068), .A3(n6857), .A4(n9968), 
        .Y(n533) );
  AO22X1_HVT U483 ( .A1(\ram[1][217] ), .A2(n7067), .A3(n6846), .A4(n9971), 
        .Y(n534) );
  AO22X1_HVT U484 ( .A1(\ram[1][218] ), .A2(n7065), .A3(n6845), .A4(n9974), 
        .Y(n535) );
  AO22X1_HVT U485 ( .A1(\ram[1][219] ), .A2(n7066), .A3(n6873), .A4(n9977), 
        .Y(n536) );
  AO22X1_HVT U486 ( .A1(\ram[1][220] ), .A2(n7055), .A3(n6844), .A4(n9981), 
        .Y(n537) );
  AO22X1_HVT U487 ( .A1(\ram[1][221] ), .A2(n4612), .A3(n6885), .A4(n9984), 
        .Y(n538) );
  AO22X1_HVT U488 ( .A1(\ram[1][222] ), .A2(n4332), .A3(n10337), .A4(n9987), 
        .Y(n539) );
  AO22X1_HVT U489 ( .A1(\ram[1][223] ), .A2(n7058), .A3(n6884), .A4(n9990), 
        .Y(n540) );
  AO22X1_HVT U490 ( .A1(\ram[1][224] ), .A2(n5480), .A3(n6883), .A4(n9993), 
        .Y(n541) );
  AO22X1_HVT U491 ( .A1(\ram[1][225] ), .A2(n7066), .A3(n6881), .A4(n9996), 
        .Y(n542) );
  AO22X1_HVT U492 ( .A1(\ram[1][226] ), .A2(n7065), .A3(n6880), .A4(n9999), 
        .Y(n543) );
  AO22X1_HVT U493 ( .A1(\ram[1][227] ), .A2(n5480), .A3(n6878), .A4(n10002), 
        .Y(n544) );
  AO22X1_HVT U494 ( .A1(\ram[1][228] ), .A2(n4673), .A3(n6877), .A4(n10005), 
        .Y(n545) );
  AO22X1_HVT U495 ( .A1(\ram[1][229] ), .A2(n4677), .A3(n6874), .A4(n10008), 
        .Y(n546) );
  AO22X1_HVT U496 ( .A1(\ram[1][230] ), .A2(n7052), .A3(n6873), .A4(n10011), 
        .Y(n547) );
  AO22X1_HVT U497 ( .A1(\ram[1][231] ), .A2(n7050), .A3(n6872), .A4(n10014), 
        .Y(n548) );
  AO22X1_HVT U498 ( .A1(\ram[1][232] ), .A2(n7036), .A3(n6841), .A4(n10018), 
        .Y(n549) );
  AO22X1_HVT U499 ( .A1(\ram[1][233] ), .A2(n4677), .A3(n6869), .A4(n10021), 
        .Y(n550) );
  AO22X1_HVT U500 ( .A1(\ram[1][234] ), .A2(n7034), .A3(n6868), .A4(n10024), 
        .Y(n551) );
  AO22X1_HVT U501 ( .A1(\ram[1][235] ), .A2(n7041), .A3(n6871), .A4(n10027), 
        .Y(n552) );
  AO22X1_HVT U502 ( .A1(\ram[1][236] ), .A2(n7045), .A3(n6866), .A4(n10030), 
        .Y(n553) );
  AO22X1_HVT U503 ( .A1(\ram[1][237] ), .A2(n7052), .A3(n6865), .A4(n10033), 
        .Y(n554) );
  AO22X1_HVT U504 ( .A1(\ram[1][238] ), .A2(n7034), .A3(n6864), .A4(n10036), 
        .Y(n555) );
  AO22X1_HVT U505 ( .A1(\ram[1][239] ), .A2(n7042), .A3(n6850), .A4(n10039), 
        .Y(n556) );
  AO22X1_HVT U506 ( .A1(\ram[1][240] ), .A2(n7058), .A3(n6849), .A4(n10043), 
        .Y(n557) );
  AO22X1_HVT U507 ( .A1(\ram[1][241] ), .A2(n7056), .A3(n6847), .A4(n10046), 
        .Y(n558) );
  AO22X1_HVT U508 ( .A1(\ram[1][242] ), .A2(n7058), .A3(n10342), .A4(n10049), 
        .Y(n559) );
  AO22X1_HVT U509 ( .A1(\ram[1][243] ), .A2(n7057), .A3(n6846), .A4(n10052), 
        .Y(n560) );
  AO22X1_HVT U511 ( .A1(\ram[1][245] ), .A2(n7031), .A3(n10336), .A4(n10058), 
        .Y(n562) );
  AO22X1_HVT U512 ( .A1(\ram[1][246] ), .A2(n7030), .A3(n6844), .A4(n10061), 
        .Y(n563) );
  AO22X1_HVT U513 ( .A1(\ram[1][247] ), .A2(n4574), .A3(n6877), .A4(n10064), 
        .Y(n564) );
  AO22X1_HVT U514 ( .A1(\ram[1][248] ), .A2(n4261), .A3(n6874), .A4(n10068), 
        .Y(n565) );
  AO22X1_HVT U515 ( .A1(\ram[1][249] ), .A2(n7081), .A3(n6873), .A4(n10071), 
        .Y(n566) );
  AO22X1_HVT U516 ( .A1(\ram[1][250] ), .A2(n7080), .A3(n6872), .A4(n10074), 
        .Y(n567) );
  AO22X1_HVT U517 ( .A1(\ram[1][251] ), .A2(n4259), .A3(n6854), .A4(n10077), 
        .Y(n568) );
  AO22X1_HVT U519 ( .A1(\ram[1][253] ), .A2(n7065), .A3(n6861), .A4(n10084), 
        .Y(n570) );
  AO22X1_HVT U520 ( .A1(\ram[1][254] ), .A2(n7066), .A3(n6860), .A4(n10087), 
        .Y(n571) );
  AO22X1_HVT U521 ( .A1(\ram[1][255] ), .A2(n5480), .A3(n6832), .A4(n10090), 
        .Y(n572) );
  AND2X1_HVT U524 ( .A1(n5822), .A2(n5042), .Y(n12) );
  AO22X1_HVT U525 ( .A1(\ram[2][0] ), .A2(n7178), .A3(n6274), .A4(n9306), .Y(
        n573) );
  AO22X1_HVT U526 ( .A1(\ram[2][1] ), .A2(n7179), .A3(n6286), .A4(n9309), .Y(
        n574) );
  AO22X1_HVT U527 ( .A1(\ram[2][2] ), .A2(n7177), .A3(n6313), .A4(n9313), .Y(
        n575) );
  AO22X1_HVT U528 ( .A1(\ram[2][3] ), .A2(n7176), .A3(n10320), .A4(n9315), .Y(
        n576) );
  AO22X1_HVT U529 ( .A1(\ram[2][4] ), .A2(n4709), .A3(n10321), .A4(n9319), .Y(
        n577) );
  AO22X1_HVT U530 ( .A1(\ram[2][5] ), .A2(n4709), .A3(n6311), .A4(n9322), .Y(
        n578) );
  AO22X1_HVT U531 ( .A1(\ram[2][6] ), .A2(n4709), .A3(n6296), .A4(n9325), .Y(
        n579) );
  AO22X1_HVT U533 ( .A1(\ram[2][8] ), .A2(n7173), .A3(n6305), .A4(n9331), .Y(
        n581) );
  AO22X1_HVT U534 ( .A1(\ram[2][9] ), .A2(n7172), .A3(n6304), .A4(n9334), .Y(
        n582) );
  AO22X1_HVT U535 ( .A1(\ram[2][10] ), .A2(n7171), .A3(n6295), .A4(n9337), .Y(
        n583) );
  AO22X1_HVT U536 ( .A1(\ram[2][11] ), .A2(n7170), .A3(n6326), .A4(n9340), .Y(
        n584) );
  AO22X1_HVT U537 ( .A1(\ram[2][12] ), .A2(n7158), .A3(n6325), .A4(n9344), .Y(
        n585) );
  AO22X1_HVT U538 ( .A1(\ram[2][13] ), .A2(n7157), .A3(n6322), .A4(n9347), .Y(
        n586) );
  AO22X1_HVT U539 ( .A1(\ram[2][14] ), .A2(n7156), .A3(n6321), .A4(n9350), .Y(
        n587) );
  AO22X1_HVT U540 ( .A1(\ram[2][15] ), .A2(n7155), .A3(n6319), .A4(n9353), .Y(
        n588) );
  AO22X1_HVT U541 ( .A1(\ram[2][16] ), .A2(n7186), .A3(n6318), .A4(n9356), .Y(
        n589) );
  AO22X1_HVT U542 ( .A1(\ram[2][17] ), .A2(n4316), .A3(n6316), .A4(n9359), .Y(
        n590) );
  AO22X1_HVT U543 ( .A1(\ram[2][18] ), .A2(n7184), .A3(n6315), .A4(n9362), .Y(
        n591) );
  AO22X1_HVT U544 ( .A1(\ram[2][19] ), .A2(n7182), .A3(n6314), .A4(n9365), .Y(
        n592) );
  AO22X1_HVT U545 ( .A1(\ram[2][20] ), .A2(n7193), .A3(n6313), .A4(n9368), .Y(
        n593) );
  AO22X1_HVT U546 ( .A1(\ram[2][21] ), .A2(n4650), .A3(n10320), .A4(n9370), 
        .Y(n594) );
  AO22X1_HVT U547 ( .A1(\ram[2][22] ), .A2(n4303), .A3(n10322), .A4(n9373), 
        .Y(n595) );
  AO22X1_HVT U548 ( .A1(\ram[2][23] ), .A2(n7193), .A3(n6311), .A4(n9376), .Y(
        n596) );
  AO22X1_HVT U549 ( .A1(\ram[2][24] ), .A2(n5160), .A3(n6310), .A4(n9379), .Y(
        n597) );
  AO22X1_HVT U550 ( .A1(\ram[2][25] ), .A2(n7199), .A3(n6309), .A4(n9382), .Y(
        n598) );
  AO22X1_HVT U551 ( .A1(\ram[2][26] ), .A2(n7202), .A3(n6308), .A4(n9385), .Y(
        n599) );
  AO22X1_HVT U552 ( .A1(\ram[2][27] ), .A2(n7202), .A3(n6305), .A4(n9388), .Y(
        n600) );
  AO22X1_HVT U553 ( .A1(\ram[2][28] ), .A2(n7194), .A3(n6304), .A4(n9391), .Y(
        n601) );
  AO22X1_HVT U554 ( .A1(\ram[2][29] ), .A2(n7196), .A3(n6302), .A4(n9394), .Y(
        n602) );
  AO22X1_HVT U555 ( .A1(\ram[2][30] ), .A2(n7195), .A3(n6301), .A4(n9397), .Y(
        n603) );
  AO22X1_HVT U556 ( .A1(\ram[2][31] ), .A2(n7194), .A3(n6298), .A4(n9400), .Y(
        n604) );
  AO22X1_HVT U557 ( .A1(\ram[2][32] ), .A2(n7164), .A3(n6285), .A4(n9403), .Y(
        n605) );
  AO22X1_HVT U558 ( .A1(\ram[2][33] ), .A2(n7166), .A3(n6281), .A4(n9406), .Y(
        n606) );
  AO22X1_HVT U559 ( .A1(\ram[2][34] ), .A2(n7165), .A3(n6326), .A4(n9409), .Y(
        n607) );
  AO22X1_HVT U560 ( .A1(\ram[2][35] ), .A2(n7164), .A3(n6325), .A4(n9412), .Y(
        n608) );
  AO22X1_HVT U561 ( .A1(\ram[2][36] ), .A2(n7165), .A3(n6322), .A4(n9415), .Y(
        n609) );
  AO22X1_HVT U562 ( .A1(\ram[2][37] ), .A2(n7165), .A3(n6321), .A4(n9418), .Y(
        n610) );
  AO22X1_HVT U563 ( .A1(\ram[2][38] ), .A2(n4564), .A3(n6319), .A4(n9421), .Y(
        n611) );
  AO22X1_HVT U564 ( .A1(\ram[2][39] ), .A2(n7165), .A3(n6318), .A4(n9424), .Y(
        n612) );
  AO22X1_HVT U565 ( .A1(\ram[2][40] ), .A2(n7173), .A3(n6316), .A4(n9427), .Y(
        n613) );
  AO22X1_HVT U566 ( .A1(\ram[2][41] ), .A2(n7172), .A3(n6315), .A4(n9430), .Y(
        n614) );
  AO22X1_HVT U567 ( .A1(\ram[2][42] ), .A2(n7171), .A3(n6314), .A4(n9433), .Y(
        n615) );
  AO22X1_HVT U568 ( .A1(\ram[2][43] ), .A2(n7170), .A3(n6313), .A4(n9436), .Y(
        n616) );
  AO22X1_HVT U569 ( .A1(\ram[2][44] ), .A2(n7162), .A3(n10321), .A4(n9439), 
        .Y(n617) );
  AO22X1_HVT U570 ( .A1(\ram[2][45] ), .A2(n7161), .A3(n6308), .A4(n9442), .Y(
        n618) );
  AO22X1_HVT U571 ( .A1(\ram[2][46] ), .A2(n7160), .A3(n6271), .A4(n9445), .Y(
        n619) );
  AO22X1_HVT U572 ( .A1(\ram[2][47] ), .A2(n7159), .A3(n6270), .A4(n9448), .Y(
        n620) );
  AO22X1_HVT U574 ( .A1(\ram[2][49] ), .A2(n7162), .A3(n6311), .A4(n9454), .Y(
        n622) );
  AO22X1_HVT U575 ( .A1(\ram[2][50] ), .A2(n7161), .A3(n6310), .A4(n9457), .Y(
        n623) );
  AO22X1_HVT U576 ( .A1(\ram[2][51] ), .A2(n7160), .A3(n6309), .A4(n9460), .Y(
        n624) );
  AO22X1_HVT U577 ( .A1(\ram[2][52] ), .A2(n7159), .A3(n6308), .A4(n9463), .Y(
        n625) );
  AO22X1_HVT U578 ( .A1(\ram[2][53] ), .A2(n7206), .A3(n6305), .A4(n9466), .Y(
        n626) );
  AO22X1_HVT U580 ( .A1(\ram[2][55] ), .A2(n7204), .A3(n6266), .A4(n9472), .Y(
        n628) );
  AO22X1_HVT U581 ( .A1(\ram[2][56] ), .A2(n7203), .A3(n6265), .A4(n9475), .Y(
        n629) );
  AO22X1_HVT U582 ( .A1(\ram[2][57] ), .A2(n7201), .A3(n6264), .A4(n9478), .Y(
        n630) );
  AO22X1_HVT U583 ( .A1(\ram[2][58] ), .A2(n7201), .A3(n10324), .A4(n9481), 
        .Y(n631) );
  AO22X1_HVT U584 ( .A1(\ram[2][59] ), .A2(n5160), .A3(n6263), .A4(n9484), .Y(
        n632) );
  AO22X1_HVT U585 ( .A1(\ram[2][60] ), .A2(n7173), .A3(n6284), .A4(n9487), .Y(
        n633) );
  AO22X1_HVT U586 ( .A1(\ram[2][61] ), .A2(n7172), .A3(n6263), .A4(n9490), .Y(
        n634) );
  AO22X1_HVT U587 ( .A1(\ram[2][62] ), .A2(n7171), .A3(n6268), .A4(n9493), .Y(
        n635) );
  AO22X1_HVT U588 ( .A1(\ram[2][63] ), .A2(n7170), .A3(n6267), .A4(n9496), .Y(
        n636) );
  AO22X1_HVT U589 ( .A1(\ram[2][64] ), .A2(n7192), .A3(n6296), .A4(n9499), .Y(
        n637) );
  AO22X1_HVT U590 ( .A1(\ram[2][65] ), .A2(n7192), .A3(n6264), .A4(n9502), .Y(
        n638) );
  AO22X1_HVT U591 ( .A1(\ram[2][66] ), .A2(n4408), .A3(n6262), .A4(n9505), .Y(
        n639) );
  AO22X1_HVT U593 ( .A1(\ram[2][68] ), .A2(n7192), .A3(n6268), .A4(n9511), .Y(
        n641) );
  AO22X1_HVT U594 ( .A1(\ram[2][69] ), .A2(n7192), .A3(n6267), .A4(n9514), .Y(
        n642) );
  AO22X1_HVT U595 ( .A1(\ram[2][70] ), .A2(n7190), .A3(n6296), .A4(n9517), .Y(
        n643) );
  AO22X1_HVT U596 ( .A1(\ram[2][71] ), .A2(n7189), .A3(n6295), .A4(n9520), .Y(
        n644) );
  AO22X1_HVT U598 ( .A1(\ram[2][73] ), .A2(n7202), .A3(n6279), .A4(n9526), .Y(
        n646) );
  AO22X1_HVT U599 ( .A1(\ram[2][74] ), .A2(n7199), .A3(n6278), .A4(n9529), .Y(
        n647) );
  AO22X1_HVT U600 ( .A1(\ram[2][75] ), .A2(n7199), .A3(n6275), .A4(n9532), .Y(
        n648) );
  AO22X1_HVT U601 ( .A1(\ram[2][76] ), .A2(n7173), .A3(n6274), .A4(n9535), .Y(
        n649) );
  AO22X1_HVT U602 ( .A1(\ram[2][77] ), .A2(n7172), .A3(n6288), .A4(n9538), .Y(
        n650) );
  AO22X1_HVT U603 ( .A1(\ram[2][78] ), .A2(n7171), .A3(n6272), .A4(n9541), .Y(
        n651) );
  AO22X1_HVT U604 ( .A1(\ram[2][79] ), .A2(n7170), .A3(n6271), .A4(n9544), .Y(
        n652) );
  AO22X1_HVT U605 ( .A1(\ram[2][80] ), .A2(n7182), .A3(n6270), .A4(n9547), .Y(
        n653) );
  AO22X1_HVT U606 ( .A1(\ram[2][81] ), .A2(n7181), .A3(n6266), .A4(n9550), .Y(
        n654) );
  AO22X1_HVT U607 ( .A1(\ram[2][82] ), .A2(n7180), .A3(n6265), .A4(n9553), .Y(
        n655) );
  AO22X1_HVT U608 ( .A1(\ram[2][83] ), .A2(n7179), .A3(n6264), .A4(n9556), .Y(
        n656) );
  AO22X1_HVT U609 ( .A1(\ram[2][84] ), .A2(n7158), .A3(n6315), .A4(n9559), .Y(
        n657) );
  AO22X1_HVT U610 ( .A1(\ram[2][85] ), .A2(n7157), .A3(n6314), .A4(n9562), .Y(
        n658) );
  AO22X1_HVT U611 ( .A1(\ram[2][86] ), .A2(n7156), .A3(n6267), .A4(n9565), .Y(
        n659) );
  AO22X1_HVT U612 ( .A1(\ram[2][87] ), .A2(n7155), .A3(n6309), .A4(n9568), .Y(
        n660) );
  AO22X1_HVT U613 ( .A1(\ram[2][88] ), .A2(n7181), .A3(n6308), .A4(n9571), .Y(
        n661) );
  AO22X1_HVT U614 ( .A1(\ram[2][89] ), .A2(n7181), .A3(n6291), .A4(n9574), .Y(
        n662) );
  AO22X1_HVT U615 ( .A1(\ram[2][90] ), .A2(n7180), .A3(n6290), .A4(n9577), .Y(
        n663) );
  AO22X1_HVT U616 ( .A1(\ram[2][91] ), .A2(n7178), .A3(n6289), .A4(n9580), .Y(
        n664) );
  AO22X1_HVT U617 ( .A1(\ram[2][92] ), .A2(n7196), .A3(n6288), .A4(n9583), .Y(
        n665) );
  AO22X1_HVT U618 ( .A1(\ram[2][93] ), .A2(n7194), .A3(n6287), .A4(n9586), .Y(
        n666) );
  AO22X1_HVT U619 ( .A1(\ram[2][94] ), .A2(n4303), .A3(n6286), .A4(n9589), .Y(
        n667) );
  AO22X1_HVT U620 ( .A1(\ram[2][95] ), .A2(n7194), .A3(n6285), .A4(n9592), .Y(
        n668) );
  AO22X1_HVT U621 ( .A1(\ram[2][96] ), .A2(n7162), .A3(n6266), .A4(n9595), .Y(
        n669) );
  AO22X1_HVT U622 ( .A1(\ram[2][97] ), .A2(n7161), .A3(n6265), .A4(n9598), .Y(
        n670) );
  AO22X1_HVT U623 ( .A1(\ram[2][98] ), .A2(n7160), .A3(n6288), .A4(n9601), .Y(
        n671) );
  AO22X1_HVT U624 ( .A1(\ram[2][99] ), .A2(n7159), .A3(n6287), .A4(n9604), .Y(
        n672) );
  AO22X1_HVT U625 ( .A1(\ram[2][100] ), .A2(n4317), .A3(n6286), .A4(n9607), 
        .Y(n673) );
  AO22X1_HVT U626 ( .A1(\ram[2][101] ), .A2(n7186), .A3(n6285), .A4(n9610), 
        .Y(n674) );
  AO22X1_HVT U627 ( .A1(\ram[2][102] ), .A2(n7184), .A3(n6284), .A4(n9613), 
        .Y(n675) );
  AO22X1_HVT U628 ( .A1(\ram[2][103] ), .A2(n7183), .A3(n6279), .A4(n9616), 
        .Y(n676) );
  AO22X1_HVT U629 ( .A1(\ram[2][104] ), .A2(n7183), .A3(n6278), .A4(n9619), 
        .Y(n677) );
  AO22X1_HVT U630 ( .A1(\ram[2][105] ), .A2(n7182), .A3(n6275), .A4(n9622), 
        .Y(n678) );
  AO22X1_HVT U631 ( .A1(\ram[2][106] ), .A2(n7180), .A3(n6318), .A4(n9625), 
        .Y(n679) );
  AO22X1_HVT U632 ( .A1(\ram[2][107] ), .A2(n7175), .A3(n6316), .A4(n9628), 
        .Y(n680) );
  AO22X1_HVT U633 ( .A1(\ram[2][108] ), .A2(n5209), .A3(n6294), .A4(n9631), 
        .Y(n681) );
  AO22X1_HVT U634 ( .A1(\ram[2][109] ), .A2(n7179), .A3(n6291), .A4(n9634), 
        .Y(n682) );
  AO22X1_HVT U635 ( .A1(\ram[2][110] ), .A2(n7177), .A3(n6285), .A4(n9637), 
        .Y(n683) );
  AO22X1_HVT U636 ( .A1(\ram[2][111] ), .A2(n7176), .A3(n6284), .A4(n9640), 
        .Y(n684) );
  AO22X1_HVT U637 ( .A1(\ram[2][112] ), .A2(n7178), .A3(n6279), .A4(n9643), 
        .Y(n685) );
  AO22X1_HVT U638 ( .A1(\ram[2][113] ), .A2(n7179), .A3(n6278), .A4(n9646), 
        .Y(n686) );
  AO22X1_HVT U639 ( .A1(\ram[2][114] ), .A2(n7177), .A3(n6275), .A4(n9649), 
        .Y(n687) );
  AO22X1_HVT U640 ( .A1(\ram[2][115] ), .A2(n7176), .A3(n6274), .A4(n9652), 
        .Y(n688) );
  AO22X1_HVT U641 ( .A1(\ram[2][116] ), .A2(n4650), .A3(n6284), .A4(n9655), 
        .Y(n689) );
  AO22X1_HVT U642 ( .A1(\ram[2][117] ), .A2(n7194), .A3(n6272), .A4(n9658), 
        .Y(n690) );
  AO22X1_HVT U643 ( .A1(\ram[2][118] ), .A2(n7196), .A3(n6271), .A4(n9661), 
        .Y(n691) );
  AO22X1_HVT U644 ( .A1(\ram[2][119] ), .A2(n7195), .A3(n6270), .A4(n9664), 
        .Y(n692) );
  AO22X1_HVT U645 ( .A1(\ram[2][120] ), .A2(n7202), .A3(n6311), .A4(n9667), 
        .Y(n693) );
  AO22X1_HVT U646 ( .A1(\ram[2][121] ), .A2(n7200), .A3(n6310), .A4(n9670), 
        .Y(n694) );
  AO22X1_HVT U647 ( .A1(\ram[2][122] ), .A2(n7199), .A3(n6309), .A4(n9673), 
        .Y(n695) );
  AO22X1_HVT U648 ( .A1(\ram[2][123] ), .A2(n5160), .A3(n6308), .A4(n9676), 
        .Y(n696) );
  AO22X1_HVT U649 ( .A1(\ram[2][124] ), .A2(n7179), .A3(n6305), .A4(n9679), 
        .Y(n697) );
  AO22X1_HVT U650 ( .A1(\ram[2][125] ), .A2(n5209), .A3(n6304), .A4(n9682), 
        .Y(n698) );
  AO22X1_HVT U651 ( .A1(\ram[2][126] ), .A2(n7177), .A3(n6302), .A4(n9685), 
        .Y(n699) );
  AO22X1_HVT U652 ( .A1(\ram[2][127] ), .A2(n7176), .A3(n6301), .A4(n9688), 
        .Y(n700) );
  AO22X1_HVT U655 ( .A1(\ram[2][130] ), .A2(n7166), .A3(n6281), .A4(n9697), 
        .Y(n703) );
  AO22X1_HVT U656 ( .A1(\ram[2][131] ), .A2(n4709), .A3(n6280), .A4(n9700), 
        .Y(n704) );
  AO22X1_HVT U657 ( .A1(\ram[2][132] ), .A2(n7178), .A3(n6311), .A4(n9703), 
        .Y(n705) );
  AO22X1_HVT U658 ( .A1(\ram[2][133] ), .A2(n7178), .A3(n6310), .A4(n9706), 
        .Y(n706) );
  AO22X1_HVT U659 ( .A1(\ram[2][134] ), .A2(n7177), .A3(n6322), .A4(n9709), 
        .Y(n707) );
  AO22X1_HVT U660 ( .A1(\ram[2][135] ), .A2(n7176), .A3(n6321), .A4(n9712), 
        .Y(n708) );
  AO22X1_HVT U661 ( .A1(\ram[2][136] ), .A2(n7167), .A3(n6319), .A4(n9715), 
        .Y(n709) );
  AO22X1_HVT U662 ( .A1(\ram[2][137] ), .A2(n7164), .A3(n6318), .A4(n9718), 
        .Y(n710) );
  AO22X1_HVT U663 ( .A1(\ram[2][138] ), .A2(n7164), .A3(n6316), .A4(n9721), 
        .Y(n711) );
  AO22X1_HVT U664 ( .A1(\ram[2][139] ), .A2(n7167), .A3(n6315), .A4(n9724), 
        .Y(n712) );
  AO22X1_HVT U665 ( .A1(\ram[2][140] ), .A2(n7173), .A3(n6314), .A4(n9728), 
        .Y(n713) );
  AO22X1_HVT U666 ( .A1(\ram[2][141] ), .A2(n7172), .A3(n6313), .A4(n9731), 
        .Y(n714) );
  AO22X1_HVT U667 ( .A1(\ram[2][142] ), .A2(n7171), .A3(n10323), .A4(n9734), 
        .Y(n715) );
  AO22X1_HVT U668 ( .A1(\ram[2][143] ), .A2(n7170), .A3(n10323), .A4(n9737), 
        .Y(n716) );
  AO22X1_HVT U669 ( .A1(\ram[2][144] ), .A2(n7162), .A3(n6281), .A4(n9741), 
        .Y(n717) );
  AO22X1_HVT U670 ( .A1(\ram[2][145] ), .A2(n7161), .A3(n6280), .A4(n9744), 
        .Y(n718) );
  AO22X1_HVT U671 ( .A1(\ram[2][146] ), .A2(n7160), .A3(n6294), .A4(n9747), 
        .Y(n719) );
  AO22X1_HVT U672 ( .A1(\ram[2][147] ), .A2(n7159), .A3(n6281), .A4(n9750), 
        .Y(n720) );
  AO22X1_HVT U673 ( .A1(\ram[2][148] ), .A2(n4317), .A3(n6291), .A4(n9754), 
        .Y(n721) );
  AO22X1_HVT U674 ( .A1(\ram[2][149] ), .A2(n4315), .A3(n6290), .A4(n9757), 
        .Y(n722) );
  AO22X1_HVT U675 ( .A1(\ram[2][150] ), .A2(n7184), .A3(n6289), .A4(n9760), 
        .Y(n723) );
  AO22X1_HVT U676 ( .A1(\ram[2][151] ), .A2(n7183), .A3(n6325), .A4(n9763), 
        .Y(n724) );
  AO22X1_HVT U677 ( .A1(\ram[2][152] ), .A2(n5160), .A3(n6322), .A4(n9766), 
        .Y(n725) );
  AO22X1_HVT U678 ( .A1(\ram[2][153] ), .A2(n7201), .A3(n6321), .A4(n9769), 
        .Y(n726) );
  AO22X1_HVT U679 ( .A1(\ram[2][154] ), .A2(n7199), .A3(n6319), .A4(n9772), 
        .Y(n727) );
  AO22X1_HVT U680 ( .A1(\ram[2][155] ), .A2(n7201), .A3(n6268), .A4(n9775), 
        .Y(n728) );
  AO22X1_HVT U681 ( .A1(\ram[2][156] ), .A2(n4303), .A3(n6275), .A4(n9779), 
        .Y(n729) );
  AO22X1_HVT U682 ( .A1(\ram[2][157] ), .A2(n7193), .A3(n6281), .A4(n9782), 
        .Y(n730) );
  AO22X1_HVT U683 ( .A1(\ram[2][158] ), .A2(n7196), .A3(n6280), .A4(n9785), 
        .Y(n731) );
  AO22X1_HVT U684 ( .A1(\ram[2][159] ), .A2(n7193), .A3(n6294), .A4(n9788), 
        .Y(n732) );
  AO22X1_HVT U685 ( .A1(\ram[2][160] ), .A2(n7191), .A3(n6294), .A4(n9792), 
        .Y(n733) );
  AO22X1_HVT U686 ( .A1(\ram[2][161] ), .A2(n7191), .A3(n6291), .A4(n9795), 
        .Y(n734) );
  AO22X1_HVT U687 ( .A1(\ram[2][162] ), .A2(n7190), .A3(n6290), .A4(n9798), 
        .Y(n735) );
  AO22X1_HVT U688 ( .A1(\ram[2][163] ), .A2(n7192), .A3(n6289), .A4(n9801), 
        .Y(n736) );
  AO22X1_HVT U689 ( .A1(\ram[2][164] ), .A2(n7206), .A3(n6288), .A4(n9804), 
        .Y(n737) );
  AO22X1_HVT U690 ( .A1(\ram[2][165] ), .A2(n7205), .A3(n6287), .A4(n9807), 
        .Y(n738) );
  AO22X1_HVT U691 ( .A1(\ram[2][166] ), .A2(n7204), .A3(n6286), .A4(n9810), 
        .Y(n739) );
  AO22X1_HVT U692 ( .A1(\ram[2][167] ), .A2(n7203), .A3(n6287), .A4(n9813), 
        .Y(n740) );
  AO22X1_HVT U693 ( .A1(\ram[2][168] ), .A2(n7196), .A3(n6266), .A4(n9816), 
        .Y(n741) );
  AO22X1_HVT U694 ( .A1(\ram[2][169] ), .A2(n7195), .A3(n6265), .A4(n9819), 
        .Y(n742) );
  AO22X1_HVT U695 ( .A1(\ram[2][170] ), .A2(n7195), .A3(n6264), .A4(n9822), 
        .Y(n743) );
  AO22X1_HVT U696 ( .A1(\ram[2][171] ), .A2(n4650), .A3(n10323), .A4(n9825), 
        .Y(n744) );
  AO22X1_HVT U697 ( .A1(\ram[2][172] ), .A2(n7206), .A3(n6263), .A4(n9829), 
        .Y(n745) );
  AO22X1_HVT U698 ( .A1(\ram[2][173] ), .A2(n7205), .A3(n6268), .A4(n9832), 
        .Y(n746) );
  AO22X1_HVT U699 ( .A1(\ram[2][174] ), .A2(n7204), .A3(n6267), .A4(n9835), 
        .Y(n747) );
  AO22X1_HVT U700 ( .A1(\ram[2][175] ), .A2(n7203), .A3(n6296), .A4(n9838), 
        .Y(n748) );
  AO22X1_HVT U701 ( .A1(\ram[2][176] ), .A2(n7166), .A3(n6295), .A4(n9842), 
        .Y(n749) );
  AO22X1_HVT U702 ( .A1(\ram[2][177] ), .A2(n7167), .A3(n6326), .A4(n9845), 
        .Y(n750) );
  AO22X1_HVT U703 ( .A1(\ram[2][178] ), .A2(n7167), .A3(n6325), .A4(n9848), 
        .Y(n751) );
  AO22X1_HVT U704 ( .A1(\ram[2][179] ), .A2(n7166), .A3(n6298), .A4(n9851), 
        .Y(n752) );
  AO22X1_HVT U705 ( .A1(\ram[2][180] ), .A2(n7162), .A3(n6287), .A4(n9855), 
        .Y(n753) );
  AO22X1_HVT U706 ( .A1(\ram[2][181] ), .A2(n7161), .A3(n6286), .A4(n9858), 
        .Y(n754) );
  AO22X1_HVT U707 ( .A1(\ram[2][182] ), .A2(n7160), .A3(n6285), .A4(n9861), 
        .Y(n755) );
  AO22X1_HVT U708 ( .A1(\ram[2][183] ), .A2(n7159), .A3(n6284), .A4(n9864), 
        .Y(n756) );
  AO22X1_HVT U709 ( .A1(\ram[2][184] ), .A2(n4317), .A3(n6279), .A4(n9868), 
        .Y(n757) );
  AO22X1_HVT U710 ( .A1(\ram[2][185] ), .A2(n7183), .A3(n6278), .A4(n9871), 
        .Y(n758) );
  AO22X1_HVT U711 ( .A1(\ram[2][186] ), .A2(n7184), .A3(n6275), .A4(n9874), 
        .Y(n759) );
  AO22X1_HVT U712 ( .A1(\ram[2][187] ), .A2(n4316), .A3(n6274), .A4(n9877), 
        .Y(n760) );
  AO22X1_HVT U713 ( .A1(\ram[2][188] ), .A2(n7185), .A3(n6268), .A4(n9880), 
        .Y(n761) );
  AO22X1_HVT U714 ( .A1(\ram[2][189] ), .A2(n4315), .A3(n6272), .A4(n9883), 
        .Y(n762) );
  AO22X1_HVT U715 ( .A1(\ram[2][190] ), .A2(n7184), .A3(n6271), .A4(n9886), 
        .Y(n763) );
  AO22X1_HVT U716 ( .A1(\ram[2][191] ), .A2(n7181), .A3(n6270), .A4(n9889), 
        .Y(n764) );
  AO22X1_HVT U717 ( .A1(\ram[2][192] ), .A2(n7186), .A3(n6267), .A4(n9893), 
        .Y(n765) );
  AO22X1_HVT U718 ( .A1(\ram[2][193] ), .A2(n7182), .A3(n6296), .A4(n9896), 
        .Y(n766) );
  AO22X1_HVT U719 ( .A1(\ram[2][194] ), .A2(n7184), .A3(n6295), .A4(n9899), 
        .Y(n767) );
  AO22X1_HVT U720 ( .A1(\ram[2][195] ), .A2(n7186), .A3(n6326), .A4(n9902), 
        .Y(n768) );
  AO22X1_HVT U721 ( .A1(\ram[2][196] ), .A2(n7186), .A3(n6325), .A4(n9906), 
        .Y(n769) );
  AO22X1_HVT U722 ( .A1(\ram[2][197] ), .A2(n4316), .A3(n6310), .A4(n9909), 
        .Y(n770) );
  AO22X1_HVT U723 ( .A1(\ram[2][198] ), .A2(n7180), .A3(n6309), .A4(n9912), 
        .Y(n771) );
  AO22X1_HVT U724 ( .A1(\ram[2][199] ), .A2(n7174), .A3(n6308), .A4(n9915), 
        .Y(n772) );
  AO22X1_HVT U725 ( .A1(\ram[2][200] ), .A2(n7206), .A3(n6305), .A4(n9919), 
        .Y(n773) );
  AO22X1_HVT U726 ( .A1(\ram[2][201] ), .A2(n7205), .A3(n6295), .A4(n9922), 
        .Y(n774) );
  AO22X1_HVT U727 ( .A1(\ram[2][202] ), .A2(n7204), .A3(n6302), .A4(n9925), 
        .Y(n775) );
  AO22X1_HVT U728 ( .A1(\ram[2][203] ), .A2(n7203), .A3(n6301), .A4(n9928), 
        .Y(n776) );
  AO22X1_HVT U729 ( .A1(\ram[2][204] ), .A2(n4315), .A3(n6280), .A4(n9931), 
        .Y(n777) );
  AO22X1_HVT U730 ( .A1(\ram[2][205] ), .A2(n7182), .A3(n6294), .A4(n9934), 
        .Y(n778) );
  AO22X1_HVT U731 ( .A1(\ram[2][206] ), .A2(n7180), .A3(n6267), .A4(n9937), 
        .Y(n779) );
  AO22X1_HVT U732 ( .A1(\ram[2][207] ), .A2(n5209), .A3(n6291), .A4(n9940), 
        .Y(n780) );
  AO22X1_HVT U733 ( .A1(\ram[2][208] ), .A2(n7189), .A3(n6290), .A4(n9944), 
        .Y(n781) );
  AO22X1_HVT U734 ( .A1(\ram[2][209] ), .A2(n7189), .A3(n6289), .A4(n9947), 
        .Y(n782) );
  AO22X1_HVT U735 ( .A1(\ram[2][210] ), .A2(n7190), .A3(n6288), .A4(n9950), 
        .Y(n783) );
  AO22X1_HVT U736 ( .A1(\ram[2][211] ), .A2(n7191), .A3(n6287), .A4(n9953), 
        .Y(n784) );
  AO22X1_HVT U737 ( .A1(\ram[2][212] ), .A2(n7191), .A3(n6286), .A4(n9956), 
        .Y(n785) );
  AO22X1_HVT U738 ( .A1(\ram[2][213] ), .A2(n7191), .A3(n6285), .A4(n9959), 
        .Y(n786) );
  AO22X1_HVT U739 ( .A1(\ram[2][214] ), .A2(n7190), .A3(n6284), .A4(n9962), 
        .Y(n787) );
  AO22X1_HVT U740 ( .A1(\ram[2][215] ), .A2(n7192), .A3(n6279), .A4(n9965), 
        .Y(n788) );
  AO22X1_HVT U741 ( .A1(\ram[2][216] ), .A2(n5209), .A3(n6278), .A4(n9968), 
        .Y(n789) );
  AO22X1_HVT U742 ( .A1(\ram[2][217] ), .A2(n5209), .A3(n6275), .A4(n9971), 
        .Y(n790) );
  AO22X1_HVT U743 ( .A1(\ram[2][218] ), .A2(n7177), .A3(n6274), .A4(n9974), 
        .Y(n791) );
  AO22X1_HVT U744 ( .A1(\ram[2][219] ), .A2(n7176), .A3(n6279), .A4(n9977), 
        .Y(n792) );
  AO22X1_HVT U745 ( .A1(\ram[2][220] ), .A2(n7173), .A3(n6272), .A4(n9981), 
        .Y(n793) );
  AO22X1_HVT U746 ( .A1(\ram[2][221] ), .A2(n7172), .A3(n6271), .A4(n9984), 
        .Y(n794) );
  AO22X1_HVT U747 ( .A1(\ram[2][222] ), .A2(n7171), .A3(n6270), .A4(n9987), 
        .Y(n795) );
  AO22X1_HVT U748 ( .A1(\ram[2][223] ), .A2(n7170), .A3(n6266), .A4(n9990), 
        .Y(n796) );
  AO22X1_HVT U749 ( .A1(\ram[2][224] ), .A2(n7162), .A3(n6265), .A4(n9993), 
        .Y(n797) );
  AO22X1_HVT U750 ( .A1(\ram[2][225] ), .A2(n7161), .A3(n6264), .A4(n9996), 
        .Y(n798) );
  AO22X1_HVT U751 ( .A1(\ram[2][226] ), .A2(n7160), .A3(n10324), .A4(n9999), 
        .Y(n799) );
  AO22X1_HVT U752 ( .A1(\ram[2][227] ), .A2(n7159), .A3(n6263), .A4(n10002), 
        .Y(n800) );
  AO22X1_HVT U753 ( .A1(\ram[2][228] ), .A2(n7181), .A3(n6304), .A4(n10005), 
        .Y(n801) );
  AO22X1_HVT U754 ( .A1(\ram[2][229] ), .A2(n7183), .A3(n6302), .A4(n10008), 
        .Y(n802) );
  AO22X1_HVT U755 ( .A1(\ram[2][230] ), .A2(n7180), .A3(n6301), .A4(n10011), 
        .Y(n803) );
  AO22X1_HVT U756 ( .A1(\ram[2][231] ), .A2(n5160), .A3(n6298), .A4(n10014), 
        .Y(n804) );
  AO22X1_HVT U757 ( .A1(\ram[2][232] ), .A2(n7158), .A3(n6290), .A4(n10018), 
        .Y(n805) );
  AO22X1_HVT U758 ( .A1(\ram[2][233] ), .A2(n7157), .A3(n6281), .A4(n10021), 
        .Y(n806) );
  AO22X1_HVT U759 ( .A1(\ram[2][234] ), .A2(n7156), .A3(n6280), .A4(n10024), 
        .Y(n807) );
  AO22X1_HVT U760 ( .A1(\ram[2][235] ), .A2(n7155), .A3(n6294), .A4(n10027), 
        .Y(n808) );
  AO22X1_HVT U761 ( .A1(\ram[2][236] ), .A2(n7206), .A3(n6319), .A4(n10030), 
        .Y(n809) );
  AO22X1_HVT U762 ( .A1(\ram[2][237] ), .A2(n7205), .A3(n6291), .A4(n10033), 
        .Y(n810) );
  AO22X1_HVT U763 ( .A1(\ram[2][238] ), .A2(n7204), .A3(n6290), .A4(n10036), 
        .Y(n811) );
  AO22X1_HVT U764 ( .A1(\ram[2][239] ), .A2(n7203), .A3(n6289), .A4(n10039), 
        .Y(n812) );
  AO22X1_HVT U765 ( .A1(\ram[2][240] ), .A2(n7158), .A3(n6322), .A4(n10043), 
        .Y(n813) );
  AO22X1_HVT U766 ( .A1(\ram[2][241] ), .A2(n7157), .A3(n6321), .A4(n10046), 
        .Y(n814) );
  AO22X1_HVT U767 ( .A1(\ram[2][242] ), .A2(n7156), .A3(n6319), .A4(n10049), 
        .Y(n815) );
  AO22X1_HVT U768 ( .A1(\ram[2][243] ), .A2(n7155), .A3(n6318), .A4(n10052), 
        .Y(n816) );
  AO22X1_HVT U769 ( .A1(\ram[2][244] ), .A2(n7202), .A3(n6316), .A4(n10055), 
        .Y(n817) );
  AO22X1_HVT U770 ( .A1(\ram[2][245] ), .A2(n7200), .A3(n6315), .A4(n10058), 
        .Y(n818) );
  AO22X1_HVT U771 ( .A1(\ram[2][246] ), .A2(n7200), .A3(n6314), .A4(n10061), 
        .Y(n819) );
  AO22X1_HVT U772 ( .A1(\ram[2][247] ), .A2(n4564), .A3(n6313), .A4(n10064), 
        .Y(n820) );
  AO22X1_HVT U773 ( .A1(\ram[2][248] ), .A2(n7158), .A3(n6304), .A4(n10068), 
        .Y(n821) );
  AO22X1_HVT U774 ( .A1(\ram[2][249] ), .A2(n7157), .A3(n6302), .A4(n10071), 
        .Y(n822) );
  AO22X1_HVT U775 ( .A1(\ram[2][250] ), .A2(n7156), .A3(n6301), .A4(n10074), 
        .Y(n823) );
  AO22X1_HVT U776 ( .A1(\ram[2][251] ), .A2(n7155), .A3(n6298), .A4(n10077), 
        .Y(n824) );
  AO22X1_HVT U778 ( .A1(\ram[2][253] ), .A2(n7189), .A3(n10322), .A4(n10084), 
        .Y(n826) );
  AO22X1_HVT U779 ( .A1(\ram[2][254] ), .A2(n7190), .A3(n10323), .A4(n10087), 
        .Y(n827) );
  AO22X1_HVT U780 ( .A1(\ram[2][255] ), .A2(n7191), .A3(n6288), .A4(n10090), 
        .Y(n828) );
  AND2X1_HVT U783 ( .A1(n6644), .A2(n5822), .Y(n16) );
  AO22X1_HVT U790 ( .A1(\ram[3][6] ), .A2(n7123), .A3(n4294), .A4(n9325), .Y(
        n835) );
  AO22X1_HVT U791 ( .A1(\ram[3][7] ), .A2(n7122), .A3(n6767), .A4(n9328), .Y(
        n836) );
  AO22X1_HVT U793 ( .A1(\ram[3][9] ), .A2(n7110), .A3(n5243), .A4(n9334), .Y(
        n838) );
  AO22X1_HVT U794 ( .A1(\ram[3][10] ), .A2(n7109), .A3(n5250), .A4(n9337), .Y(
        n839) );
  AO22X1_HVT U795 ( .A1(\ram[3][11] ), .A2(n7108), .A3(n5267), .A4(n9340), .Y(
        n840) );
  AO22X1_HVT U796 ( .A1(\ram[3][12] ), .A2(n7100), .A3(n5243), .A4(n9344), .Y(
        n841) );
  AO22X1_HVT U797 ( .A1(\ram[3][13] ), .A2(n7099), .A3(n5266), .A4(n9347), .Y(
        n842) );
  AO22X1_HVT U798 ( .A1(\ram[3][14] ), .A2(n7098), .A3(n6768), .A4(n9350), .Y(
        n843) );
  AO22X1_HVT U799 ( .A1(\ram[3][15] ), .A2(n7134), .A3(n5252), .A4(n9353), .Y(
        n844) );
  AO22X1_HVT U803 ( .A1(\ram[3][19] ), .A2(n7103), .A3(n5276), .A4(n9365), .Y(
        n848) );
  AO22X1_HVT U804 ( .A1(\ram[3][20] ), .A2(n7106), .A3(n10308), .A4(n9368), 
        .Y(n849) );
  AO22X1_HVT U805 ( .A1(\ram[3][21] ), .A2(n7105), .A3(n5260), .A4(n9370), .Y(
        n850) );
  AO22X1_HVT U806 ( .A1(\ram[3][22] ), .A2(n7104), .A3(n5270), .A4(n9373), .Y(
        n851) );
  AO22X1_HVT U807 ( .A1(\ram[3][23] ), .A2(n7103), .A3(n5254), .A4(n9376), .Y(
        n852) );
  AO22X1_HVT U808 ( .A1(\ram[3][24] ), .A2(n7125), .A3(n5283), .A4(n9379), .Y(
        n853) );
  AO22X1_HVT U809 ( .A1(\ram[3][25] ), .A2(n7124), .A3(n5240), .A4(n9382), .Y(
        n854) );
  AO22X1_HVT U811 ( .A1(\ram[3][27] ), .A2(n7122), .A3(n5258), .A4(n9388), .Y(
        n856) );
  AO22X1_HVT U812 ( .A1(\ram[3][28] ), .A2(n7111), .A3(n10310), .A4(n9391), 
        .Y(n857) );
  AO22X1_HVT U813 ( .A1(\ram[3][29] ), .A2(n7110), .A3(n5281), .A4(n9394), .Y(
        n858) );
  AO22X1_HVT U814 ( .A1(\ram[3][30] ), .A2(n7109), .A3(n5280), .A4(n9397), .Y(
        n859) );
  AO22X1_HVT U815 ( .A1(\ram[3][31] ), .A2(n7108), .A3(n5260), .A4(n9400), .Y(
        n860) );
  AO22X1_HVT U816 ( .A1(\ram[3][32] ), .A2(n4307), .A3(n4543), .A4(n9403), .Y(
        n861) );
  AO22X1_HVT U817 ( .A1(\ram[3][33] ), .A2(n7099), .A3(n6254), .A4(n9406), .Y(
        n862) );
  AO22X1_HVT U818 ( .A1(\ram[3][34] ), .A2(n7098), .A3(n5251), .A4(n9409), .Y(
        n863) );
  AO22X1_HVT U819 ( .A1(\ram[3][35] ), .A2(n7097), .A3(n5256), .A4(n9412), .Y(
        n864) );
  AO22X1_HVT U820 ( .A1(\ram[3][36] ), .A2(n7135), .A3(n5279), .A4(n9415), .Y(
        n865) );
  AO22X1_HVT U822 ( .A1(\ram[3][38] ), .A2(n7133), .A3(n5272), .A4(n9421), .Y(
        n867) );
  AO22X1_HVT U823 ( .A1(\ram[3][39] ), .A2(n7132), .A3(n4516), .A4(n9424), .Y(
        n868) );
  AO22X1_HVT U824 ( .A1(\ram[3][40] ), .A2(n7135), .A3(n5283), .A4(n9427), .Y(
        n869) );
  AO22X1_HVT U825 ( .A1(\ram[3][41] ), .A2(n7134), .A3(n5247), .A4(n9430), .Y(
        n870) );
  AO22X1_HVT U826 ( .A1(\ram[3][42] ), .A2(n7133), .A3(n5272), .A4(n9433), .Y(
        n871) );
  AO22X1_HVT U827 ( .A1(\ram[3][43] ), .A2(n7132), .A3(n5270), .A4(n9436), .Y(
        n872) );
  AO22X1_HVT U828 ( .A1(\ram[3][44] ), .A2(n7106), .A3(n4516), .A4(n9439), .Y(
        n873) );
  AO22X1_HVT U829 ( .A1(\ram[3][45] ), .A2(n7105), .A3(n5261), .A4(n9442), .Y(
        n874) );
  AO22X1_HVT U830 ( .A1(\ram[3][46] ), .A2(n7104), .A3(n5256), .A4(n9445), .Y(
        n875) );
  AO22X1_HVT U831 ( .A1(\ram[3][47] ), .A2(n7103), .A3(n5281), .A4(n9448), .Y(
        n876) );
  AO22X1_HVT U833 ( .A1(\ram[3][49] ), .A2(n7094), .A3(n5277), .A4(n9454), .Y(
        n878) );
  AO22X1_HVT U834 ( .A1(\ram[3][50] ), .A2(n7093), .A3(n5262), .A4(n9457), .Y(
        n879) );
  AO22X1_HVT U835 ( .A1(\ram[3][51] ), .A2(n7093), .A3(n5266), .A4(n9460), .Y(
        n880) );
  AO22X1_HVT U836 ( .A1(\ram[3][52] ), .A2(n7092), .A3(n5264), .A4(n9463), .Y(
        n881) );
  AO22X1_HVT U837 ( .A1(\ram[3][53] ), .A2(n7139), .A3(n10311), .A4(n9466), 
        .Y(n882) );
  AO22X1_HVT U838 ( .A1(\ram[3][54] ), .A2(n7138), .A3(n5240), .A4(n9469), .Y(
        n883) );
  AO22X1_HVT U839 ( .A1(\ram[3][55] ), .A2(n7137), .A3(n5279), .A4(n9472), .Y(
        n884) );
  AO22X1_HVT U840 ( .A1(\ram[3][56] ), .A2(n7136), .A3(n10311), .A4(n9475), 
        .Y(n885) );
  AO22X1_HVT U842 ( .A1(\ram[3][58] ), .A2(n7134), .A3(n5247), .A4(n9481), .Y(
        n887) );
  AO22X1_HVT U843 ( .A1(\ram[3][59] ), .A2(n7133), .A3(n10313), .A4(n9484), 
        .Y(n888) );
  AO22X1_HVT U844 ( .A1(\ram[3][60] ), .A2(n7115), .A3(n5277), .A4(n9487), .Y(
        n889) );
  AO22X1_HVT U845 ( .A1(\ram[3][61] ), .A2(n4583), .A3(n5270), .A4(n9490), .Y(
        n890) );
  AO22X1_HVT U846 ( .A1(\ram[3][62] ), .A2(n7114), .A3(n5250), .A4(n9493), .Y(
        n891) );
  AO22X1_HVT U847 ( .A1(\ram[3][63] ), .A2(n7113), .A3(n5261), .A4(n9496), .Y(
        n892) );
  AO22X1_HVT U848 ( .A1(\ram[3][64] ), .A2(n7090), .A3(n10307), .A4(n9499), 
        .Y(n893) );
  AO22X1_HVT U849 ( .A1(\ram[3][65] ), .A2(n7093), .A3(n5269), .A4(n9502), .Y(
        n894) );
  AO22X1_HVT U850 ( .A1(\ram[3][66] ), .A2(n7088), .A3(n5245), .A4(n9505), .Y(
        n895) );
  AO22X1_HVT U851 ( .A1(\ram[3][67] ), .A2(n7087), .A3(n4294), .A4(n9508), .Y(
        n896) );
  AO22X1_HVT U852 ( .A1(\ram[3][68] ), .A2(n7090), .A3(n4544), .A4(n9511), .Y(
        n897) );
  AO22X1_HVT U853 ( .A1(\ram[3][69] ), .A2(n7095), .A3(n5250), .A4(n9514), .Y(
        n898) );
  AO22X1_HVT U854 ( .A1(\ram[3][70] ), .A2(n7088), .A3(n5243), .A4(n9517), .Y(
        n899) );
  AO22X1_HVT U855 ( .A1(\ram[3][71] ), .A2(n7087), .A3(n4293), .A4(n9520), .Y(
        n900) );
  AO22X1_HVT U856 ( .A1(\ram[3][72] ), .A2(n7090), .A3(n5255), .A4(n9523), .Y(
        n901) );
  AO22X1_HVT U857 ( .A1(\ram[3][73] ), .A2(n7094), .A3(n5277), .A4(n9526), .Y(
        n902) );
  AO22X1_HVT U858 ( .A1(\ram[3][74] ), .A2(n7088), .A3(n5275), .A4(n9529), .Y(
        n903) );
  AO22X1_HVT U859 ( .A1(\ram[3][75] ), .A2(n7087), .A3(n5245), .A4(n9532), .Y(
        n904) );
  AO22X1_HVT U860 ( .A1(\ram[3][76] ), .A2(n7111), .A3(n5273), .A4(n9535), .Y(
        n905) );
  AO22X1_HVT U861 ( .A1(\ram[3][77] ), .A2(n7110), .A3(n10307), .A4(n9538), 
        .Y(n906) );
  AO22X1_HVT U862 ( .A1(\ram[3][78] ), .A2(n7109), .A3(n4543), .A4(n9541), .Y(
        n907) );
  AO22X1_HVT U863 ( .A1(\ram[3][79] ), .A2(n7108), .A3(n5272), .A4(n9544), .Y(
        n908) );
  AO22X1_HVT U864 ( .A1(\ram[3][80] ), .A2(n7127), .A3(n5281), .A4(n9547), .Y(
        n909) );
  AO22X1_HVT U865 ( .A1(\ram[3][81] ), .A2(n7127), .A3(n5264), .A4(n9550), .Y(
        n910) );
  AO22X1_HVT U866 ( .A1(\ram[3][82] ), .A2(n4737), .A3(n5243), .A4(n9553), .Y(
        n911) );
  AO22X1_HVT U867 ( .A1(\ram[3][83] ), .A2(n4737), .A3(n5273), .A4(n9556), .Y(
        n912) );
  AO22X1_HVT U869 ( .A1(\ram[3][85] ), .A2(n7132), .A3(n10314), .A4(n9562), 
        .Y(n914) );
  AO22X1_HVT U870 ( .A1(\ram[3][86] ), .A2(n7126), .A3(n5247), .A4(n9565), .Y(
        n915) );
  AO22X1_HVT U873 ( .A1(\ram[3][89] ), .A2(n7126), .A3(n4254), .A4(n9574), .Y(
        n918) );
  AO22X1_HVT U874 ( .A1(\ram[3][90] ), .A2(n7125), .A3(n5270), .A4(n9577), .Y(
        n919) );
  AO22X1_HVT U875 ( .A1(\ram[3][91] ), .A2(n7135), .A3(n5279), .A4(n9580), .Y(
        n920) );
  AO22X1_HVT U876 ( .A1(\ram[3][92] ), .A2(n4307), .A3(n5264), .A4(n9583), .Y(
        n921) );
  AO22X1_HVT U877 ( .A1(\ram[3][93] ), .A2(n7099), .A3(n6766), .A4(n9586), .Y(
        n922) );
  AO22X1_HVT U878 ( .A1(\ram[3][94] ), .A2(n7098), .A3(n5260), .A4(n9589), .Y(
        n923) );
  AO22X1_HVT U879 ( .A1(\ram[3][95] ), .A2(n7097), .A3(n5266), .A4(n9592), .Y(
        n924) );
  AO22X1_HVT U880 ( .A1(\ram[3][96] ), .A2(n4307), .A3(n6254), .A4(n9595), .Y(
        n925) );
  AO22X1_HVT U882 ( .A1(\ram[3][98] ), .A2(n7098), .A3(n10313), .A4(n9601), 
        .Y(n927) );
  AO22X1_HVT U883 ( .A1(\ram[3][99] ), .A2(n7097), .A3(n5264), .A4(n9604), .Y(
        n928) );
  AO22X1_HVT U884 ( .A1(\ram[3][100] ), .A2(n7139), .A3(n10310), .A4(n9607), 
        .Y(n929) );
  AO22X1_HVT U885 ( .A1(\ram[3][101] ), .A2(n7138), .A3(n4516), .A4(n9610), 
        .Y(n930) );
  AO22X1_HVT U886 ( .A1(\ram[3][102] ), .A2(n7137), .A3(n5262), .A4(n9613), 
        .Y(n931) );
  AO22X1_HVT U887 ( .A1(\ram[3][103] ), .A2(n7136), .A3(n4517), .A4(n9616), 
        .Y(n932) );
  AO22X1_HVT U888 ( .A1(\ram[3][104] ), .A2(n7135), .A3(n5254), .A4(n9619), 
        .Y(n933) );
  AO22X1_HVT U890 ( .A1(\ram[3][106] ), .A2(n7133), .A3(n5275), .A4(n9625), 
        .Y(n935) );
  AO22X1_HVT U891 ( .A1(\ram[3][107] ), .A2(n7132), .A3(n10313), .A4(n9628), 
        .Y(n936) );
  AO22X1_HVT U892 ( .A1(\ram[3][108] ), .A2(n7129), .A3(n5264), .A4(n9631), 
        .Y(n937) );
  AO22X1_HVT U893 ( .A1(\ram[3][109] ), .A2(n4737), .A3(n6768), .A4(n9634), 
        .Y(n938) );
  AO22X1_HVT U894 ( .A1(\ram[3][110] ), .A2(n7129), .A3(n6766), .A4(n9637), 
        .Y(n939) );
  AO22X1_HVT U895 ( .A1(\ram[3][111] ), .A2(n7129), .A3(n5272), .A4(n9640), 
        .Y(n940) );
  AO22X1_HVT U896 ( .A1(\ram[3][112] ), .A2(n7139), .A3(n5251), .A4(n9643), 
        .Y(n941) );
  AO22X1_HVT U897 ( .A1(\ram[3][113] ), .A2(n7138), .A3(n4544), .A4(n9646), 
        .Y(n942) );
  AO22X1_HVT U899 ( .A1(\ram[3][115] ), .A2(n7136), .A3(n5245), .A4(n9652), 
        .Y(n944) );
  AO22X1_HVT U900 ( .A1(\ram[3][116] ), .A2(n7139), .A3(n5250), .A4(n9655), 
        .Y(n945) );
  AO22X1_HVT U901 ( .A1(\ram[3][117] ), .A2(n7138), .A3(n5269), .A4(n9658), 
        .Y(n946) );
  AO22X1_HVT U903 ( .A1(\ram[3][119] ), .A2(n7136), .A3(n4293), .A4(n9664), 
        .Y(n948) );
  AO22X1_HVT U904 ( .A1(\ram[3][120] ), .A2(n7111), .A3(n5275), .A4(n9667), 
        .Y(n949) );
  AO22X1_HVT U905 ( .A1(\ram[3][121] ), .A2(n7110), .A3(n5252), .A4(n9670), 
        .Y(n950) );
  AO22X1_HVT U906 ( .A1(\ram[3][122] ), .A2(n7109), .A3(n5261), .A4(n9673), 
        .Y(n951) );
  AO22X1_HVT U907 ( .A1(\ram[3][123] ), .A2(n7108), .A3(n10309), .A4(n9676), 
        .Y(n952) );
  AO22X1_HVT U908 ( .A1(\ram[3][124] ), .A2(n7111), .A3(n10313), .A4(n9679), 
        .Y(n953) );
  AO22X1_HVT U909 ( .A1(\ram[3][125] ), .A2(n7110), .A3(n10311), .A4(n9682), 
        .Y(n954) );
  AO22X1_HVT U910 ( .A1(\ram[3][126] ), .A2(n7109), .A3(n10313), .A4(n9685), 
        .Y(n955) );
  AO22X1_HVT U911 ( .A1(\ram[3][127] ), .A2(n7108), .A3(n5251), .A4(n9688), 
        .Y(n956) );
  AO22X1_HVT U912 ( .A1(\ram[3][128] ), .A2(n7115), .A3(n4254), .A4(n9691), 
        .Y(n957) );
  AO22X1_HVT U913 ( .A1(\ram[3][129] ), .A2(n4583), .A3(n5249), .A4(n9694), 
        .Y(n958) );
  AO22X1_HVT U914 ( .A1(\ram[3][130] ), .A2(n7114), .A3(n10314), .A4(n9697), 
        .Y(n959) );
  AO22X1_HVT U915 ( .A1(\ram[3][131] ), .A2(n7113), .A3(n5283), .A4(n9700), 
        .Y(n960) );
  AO22X1_HVT U916 ( .A1(\ram[3][132] ), .A2(n4339), .A3(n5273), .A4(n9703), 
        .Y(n961) );
  AO22X1_HVT U917 ( .A1(\ram[3][133] ), .A2(n7092), .A3(n10311), .A4(n9706), 
        .Y(n962) );
  AO22X1_HVT U918 ( .A1(\ram[3][134] ), .A2(n7119), .A3(n4296), .A4(n9709), 
        .Y(n963) );
  AO22X1_HVT U919 ( .A1(\ram[3][135] ), .A2(n7118), .A3(n5250), .A4(n9712), 
        .Y(n964) );
  AO22X1_HVT U920 ( .A1(\ram[3][136] ), .A2(n7117), .A3(n5254), .A4(n9715), 
        .Y(n965) );
  AO22X1_HVT U921 ( .A1(\ram[3][137] ), .A2(n7116), .A3(n5269), .A4(n9718), 
        .Y(n966) );
  AO22X1_HVT U922 ( .A1(\ram[3][138] ), .A2(n7115), .A3(n5275), .A4(n9721), 
        .Y(n967) );
  AO22X1_HVT U923 ( .A1(\ram[3][139] ), .A2(n7123), .A3(n5256), .A4(n9724), 
        .Y(n968) );
  AO22X1_HVT U924 ( .A1(\ram[3][140] ), .A2(n7119), .A3(n10309), .A4(n9728), 
        .Y(n969) );
  AO22X1_HVT U925 ( .A1(\ram[3][141] ), .A2(n7118), .A3(n4517), .A4(n9731), 
        .Y(n970) );
  AO22X1_HVT U926 ( .A1(\ram[3][142] ), .A2(n7117), .A3(n5250), .A4(n9734), 
        .Y(n971) );
  AO22X1_HVT U927 ( .A1(\ram[3][143] ), .A2(n7116), .A3(n5264), .A4(n9737), 
        .Y(n972) );
  AO22X1_HVT U928 ( .A1(\ram[3][144] ), .A2(n7119), .A3(n5256), .A4(n9741), 
        .Y(n973) );
  AO22X1_HVT U929 ( .A1(\ram[3][145] ), .A2(n7118), .A3(n5255), .A4(n9744), 
        .Y(n974) );
  AO22X1_HVT U930 ( .A1(\ram[3][146] ), .A2(n7117), .A3(n5266), .A4(n9747), 
        .Y(n975) );
  AO22X1_HVT U931 ( .A1(\ram[3][147] ), .A2(n7116), .A3(n5254), .A4(n9750), 
        .Y(n976) );
  AO22X1_HVT U932 ( .A1(\ram[3][148] ), .A2(n7115), .A3(n5250), .A4(n9754), 
        .Y(n977) );
  AO22X1_HVT U933 ( .A1(\ram[3][149] ), .A2(n4583), .A3(n5260), .A4(n9757), 
        .Y(n978) );
  AO22X1_HVT U934 ( .A1(\ram[3][150] ), .A2(n7114), .A3(n5270), .A4(n9760), 
        .Y(n979) );
  AO22X1_HVT U935 ( .A1(\ram[3][151] ), .A2(n7113), .A3(n10313), .A4(n9763), 
        .Y(n980) );
  AO22X1_HVT U936 ( .A1(\ram[3][152] ), .A2(n7090), .A3(n5252), .A4(n9766), 
        .Y(n981) );
  AO22X1_HVT U937 ( .A1(\ram[3][153] ), .A2(n7089), .A3(n10309), .A4(n9769), 
        .Y(n982) );
  AO22X1_HVT U938 ( .A1(\ram[3][154] ), .A2(n7088), .A3(n5281), .A4(n9772), 
        .Y(n983) );
  AO22X1_HVT U939 ( .A1(\ram[3][155] ), .A2(n7087), .A3(n4295), .A4(n9775), 
        .Y(n984) );
  AO22X1_HVT U940 ( .A1(\ram[3][156] ), .A2(n7139), .A3(n5266), .A4(n9779), 
        .Y(n985) );
  AO22X1_HVT U941 ( .A1(\ram[3][157] ), .A2(n7138), .A3(n5240), .A4(n9782), 
        .Y(n986) );
  AO22X1_HVT U942 ( .A1(\ram[3][158] ), .A2(n7137), .A3(n4254), .A4(n9785), 
        .Y(n987) );
  AO22X1_HVT U943 ( .A1(\ram[3][159] ), .A2(n7136), .A3(n5252), .A4(n9788), 
        .Y(n988) );
  AO22X1_HVT U944 ( .A1(\ram[3][160] ), .A2(n7125), .A3(n5275), .A4(n9792), 
        .Y(n989) );
  AO22X1_HVT U945 ( .A1(\ram[3][161] ), .A2(n7124), .A3(n5267), .A4(n9795), 
        .Y(n990) );
  AO22X1_HVT U946 ( .A1(\ram[3][162] ), .A2(n7123), .A3(n4254), .A4(n9798), 
        .Y(n991) );
  AO22X1_HVT U947 ( .A1(\ram[3][163] ), .A2(n7122), .A3(n5240), .A4(n9801), 
        .Y(n992) );
  AO22X1_HVT U949 ( .A1(\ram[3][165] ), .A2(n7124), .A3(n4294), .A4(n9807), 
        .Y(n994) );
  AO22X1_HVT U950 ( .A1(\ram[3][166] ), .A2(n7123), .A3(n5267), .A4(n9810), 
        .Y(n995) );
  AO22X1_HVT U951 ( .A1(\ram[3][167] ), .A2(n7122), .A3(n4517), .A4(n9813), 
        .Y(n996) );
  AO22X1_HVT U952 ( .A1(\ram[3][168] ), .A2(n7119), .A3(n10311), .A4(n9816), 
        .Y(n997) );
  AO22X1_HVT U953 ( .A1(\ram[3][169] ), .A2(n7118), .A3(n5240), .A4(n9819), 
        .Y(n998) );
  AO22X1_HVT U954 ( .A1(\ram[3][170] ), .A2(n7117), .A3(n5283), .A4(n9822), 
        .Y(n999) );
  AO22X1_HVT U955 ( .A1(\ram[3][171] ), .A2(n7116), .A3(n4295), .A4(n9825), 
        .Y(n1000) );
  AO22X1_HVT U956 ( .A1(\ram[3][172] ), .A2(n7106), .A3(n5249), .A4(n9829), 
        .Y(n1001) );
  AO22X1_HVT U957 ( .A1(\ram[3][173] ), .A2(n7105), .A3(n5280), .A4(n9832), 
        .Y(n1002) );
  AO22X1_HVT U958 ( .A1(\ram[3][174] ), .A2(n7104), .A3(n5258), .A4(n9835), 
        .Y(n1003) );
  AO22X1_HVT U960 ( .A1(\ram[3][176] ), .A2(n4583), .A3(n5243), .A4(n9842), 
        .Y(n1005) );
  AO22X1_HVT U961 ( .A1(\ram[3][177] ), .A2(n7114), .A3(n5258), .A4(n9845), 
        .Y(n1006) );
  AO22X1_HVT U962 ( .A1(\ram[3][178] ), .A2(n7113), .A3(n5262), .A4(n9848), 
        .Y(n1007) );
  AO22X1_HVT U963 ( .A1(\ram[3][179] ), .A2(n7090), .A3(n10313), .A4(n9851), 
        .Y(n1008) );
  AO22X1_HVT U964 ( .A1(\ram[3][180] ), .A2(n7095), .A3(n4543), .A4(n9855), 
        .Y(n1009) );
  AO22X1_HVT U965 ( .A1(\ram[3][181] ), .A2(n7088), .A3(n5272), .A4(n9858), 
        .Y(n1010) );
  AO22X1_HVT U967 ( .A1(\ram[3][183] ), .A2(n7122), .A3(n5254), .A4(n9864), 
        .Y(n1012) );
  AO22X1_HVT U968 ( .A1(\ram[3][184] ), .A2(n7115), .A3(n5262), .A4(n9868), 
        .Y(n1013) );
  AO22X1_HVT U969 ( .A1(\ram[3][185] ), .A2(n4583), .A3(n5252), .A4(n9871), 
        .Y(n1014) );
  AO22X1_HVT U970 ( .A1(\ram[3][186] ), .A2(n7114), .A3(n5245), .A4(n9874), 
        .Y(n1015) );
  AO22X1_HVT U971 ( .A1(\ram[3][187] ), .A2(n7113), .A3(n5280), .A4(n9877), 
        .Y(n1016) );
  AO22X1_HVT U972 ( .A1(\ram[3][188] ), .A2(n7115), .A3(n5267), .A4(n9880), 
        .Y(n1017) );
  AO22X1_HVT U973 ( .A1(\ram[3][189] ), .A2(n4583), .A3(n5273), .A4(n9883), 
        .Y(n1018) );
  AO22X1_HVT U974 ( .A1(\ram[3][190] ), .A2(n7114), .A3(n10309), .A4(n9886), 
        .Y(n1019) );
  AO22X1_HVT U975 ( .A1(\ram[3][191] ), .A2(n7113), .A3(n4254), .A4(n9889), 
        .Y(n1020) );
  AO22X1_HVT U976 ( .A1(\ram[3][192] ), .A2(n7135), .A3(n10308), .A4(n9893), 
        .Y(n1021) );
  AO22X1_HVT U977 ( .A1(\ram[3][193] ), .A2(n7134), .A3(n4293), .A4(n9896), 
        .Y(n1022) );
  AO22X1_HVT U979 ( .A1(\ram[3][195] ), .A2(n7132), .A3(n10309), .A4(n9902), 
        .Y(n1024) );
  AO22X1_HVT U980 ( .A1(\ram[3][196] ), .A2(n7128), .A3(n10309), .A4(n9906), 
        .Y(n1025) );
  AO22X1_HVT U981 ( .A1(\ram[3][197] ), .A2(n7129), .A3(n5269), .A4(n9909), 
        .Y(n1026) );
  AO22X1_HVT U982 ( .A1(\ram[3][198] ), .A2(n7127), .A3(n5280), .A4(n9912), 
        .Y(n1027) );
  AO22X1_HVT U983 ( .A1(\ram[3][199] ), .A2(n7127), .A3(n5804), .A4(n9915), 
        .Y(n1028) );
  AO22X1_HVT U984 ( .A1(\ram[3][200] ), .A2(n7125), .A3(n6768), .A4(n9919), 
        .Y(n1029) );
  AO22X1_HVT U985 ( .A1(\ram[3][201] ), .A2(n7124), .A3(n5240), .A4(n9922), 
        .Y(n1030) );
  AO22X1_HVT U986 ( .A1(\ram[3][202] ), .A2(n7123), .A3(n5264), .A4(n9925), 
        .Y(n1031) );
  AO22X1_HVT U988 ( .A1(\ram[3][204] ), .A2(n7111), .A3(n5247), .A4(n9931), 
        .Y(n1033) );
  AO22X1_HVT U989 ( .A1(\ram[3][205] ), .A2(n7110), .A3(n5275), .A4(n9934), 
        .Y(n1034) );
  AO22X1_HVT U990 ( .A1(\ram[3][206] ), .A2(n7109), .A3(n5283), .A4(n9937), 
        .Y(n1035) );
  AO22X1_HVT U991 ( .A1(\ram[3][207] ), .A2(n7108), .A3(n5272), .A4(n9940), 
        .Y(n1036) );
  AO22X1_HVT U992 ( .A1(\ram[3][208] ), .A2(n7097), .A3(n5277), .A4(n9944), 
        .Y(n1037) );
  AO22X1_HVT U993 ( .A1(\ram[3][209] ), .A2(n7106), .A3(n4293), .A4(n9947), 
        .Y(n1038) );
  AO22X1_HVT U994 ( .A1(\ram[3][210] ), .A2(n7105), .A3(n5281), .A4(n9950), 
        .Y(n1039) );
  AO22X1_HVT U995 ( .A1(\ram[3][211] ), .A2(n7104), .A3(n4295), .A4(n9953), 
        .Y(n1040) );
  AO22X1_HVT U996 ( .A1(\ram[3][212] ), .A2(n7103), .A3(n5255), .A4(n9956), 
        .Y(n1041) );
  AO22X1_HVT U997 ( .A1(\ram[3][213] ), .A2(n4338), .A3(n10311), .A4(n9959), 
        .Y(n1042) );
  AO22X1_HVT U998 ( .A1(\ram[3][214] ), .A2(n7093), .A3(n5255), .A4(n9962), 
        .Y(n1043) );
  AO22X1_HVT U999 ( .A1(\ram[3][215] ), .A2(n7124), .A3(n4296), .A4(n9965), 
        .Y(n1044) );
  AO22X1_HVT U1000 ( .A1(\ram[3][216] ), .A2(n7094), .A3(n5266), .A4(n9968), 
        .Y(n1045) );
  AO22X1_HVT U1001 ( .A1(\ram[3][217] ), .A2(n7089), .A3(n4296), .A4(n9971), 
        .Y(n1046) );
  AO22X1_HVT U1002 ( .A1(\ram[3][218] ), .A2(n7095), .A3(n6767), .A4(n9974), 
        .Y(n1047) );
  AO22X1_HVT U1003 ( .A1(\ram[3][219] ), .A2(n7092), .A3(n4295), .A4(n9977), 
        .Y(n1048) );
  AO22X1_HVT U1004 ( .A1(\ram[3][220] ), .A2(n7089), .A3(n5240), .A4(n9981), 
        .Y(n1049) );
  AO22X1_HVT U1005 ( .A1(\ram[3][221] ), .A2(n7094), .A3(n5281), .A4(n9984), 
        .Y(n1050) );
  AO22X1_HVT U1006 ( .A1(\ram[3][222] ), .A2(n7089), .A3(n5245), .A4(n9987), 
        .Y(n1051) );
  AO22X1_HVT U1008 ( .A1(\ram[3][224] ), .A2(n7106), .A3(n5251), .A4(n9993), 
        .Y(n1053) );
  AO22X1_HVT U1009 ( .A1(\ram[3][225] ), .A2(n7105), .A3(n4296), .A4(n9996), 
        .Y(n1054) );
  AO22X1_HVT U1010 ( .A1(\ram[3][226] ), .A2(n7104), .A3(n5249), .A4(n9999), 
        .Y(n1055) );
  AO22X1_HVT U1011 ( .A1(\ram[3][227] ), .A2(n7103), .A3(n6766), .A4(n10002), 
        .Y(n1056) );
  AO22X1_HVT U1012 ( .A1(\ram[3][228] ), .A2(n7093), .A3(n5256), .A4(n10005), 
        .Y(n1057) );
  AO22X1_HVT U1013 ( .A1(\ram[3][229] ), .A2(n4338), .A3(n5260), .A4(n10008), 
        .Y(n1058) );
  AO22X1_HVT U1014 ( .A1(\ram[3][230] ), .A2(n4339), .A3(n5280), .A4(n10011), 
        .Y(n1059) );
  AO22X1_HVT U1015 ( .A1(\ram[3][231] ), .A2(n7092), .A3(n5252), .A4(n10014), 
        .Y(n1060) );
  AO22X1_HVT U1016 ( .A1(\ram[3][232] ), .A2(n7119), .A3(n5240), .A4(n10018), 
        .Y(n1061) );
  AO22X1_HVT U1017 ( .A1(\ram[3][233] ), .A2(n7118), .A3(n10309), .A4(n10021), 
        .Y(n1062) );
  AO22X1_HVT U1018 ( .A1(\ram[3][234] ), .A2(n7117), .A3(n5261), .A4(n10024), 
        .Y(n1063) );
  AO22X1_HVT U1019 ( .A1(\ram[3][235] ), .A2(n7116), .A3(n4517), .A4(n10027), 
        .Y(n1064) );
  AO22X1_HVT U1020 ( .A1(\ram[3][236] ), .A2(n4737), .A3(n5245), .A4(n10030), 
        .Y(n1065) );
  AO22X1_HVT U1021 ( .A1(\ram[3][237] ), .A2(n7126), .A3(n5281), .A4(n10033), 
        .Y(n1066) );
  AO22X1_HVT U1022 ( .A1(\ram[3][238] ), .A2(n7126), .A3(n5256), .A4(n10036), 
        .Y(n1067) );
  AO22X1_HVT U1023 ( .A1(\ram[3][239] ), .A2(n7126), .A3(n5280), .A4(n10039), 
        .Y(n1068) );
  AO22X1_HVT U1024 ( .A1(\ram[3][240] ), .A2(n7128), .A3(n5275), .A4(n10043), 
        .Y(n1069) );
  AO22X1_HVT U1025 ( .A1(\ram[3][241] ), .A2(n7129), .A3(n5279), .A4(n10046), 
        .Y(n1070) );
  AO22X1_HVT U1026 ( .A1(\ram[3][242] ), .A2(n7128), .A3(n5267), .A4(n10049), 
        .Y(n1071) );
  AO22X1_HVT U1027 ( .A1(\ram[3][243] ), .A2(n7128), .A3(n5283), .A4(n10052), 
        .Y(n1072) );
  AO22X1_HVT U1028 ( .A1(\ram[3][244] ), .A2(n7089), .A3(n5272), .A4(n10055), 
        .Y(n1073) );
  AO22X1_HVT U1029 ( .A1(\ram[3][245] ), .A2(n4338), .A3(n5255), .A4(n10058), 
        .Y(n1074) );
  AO22X1_HVT U1030 ( .A1(\ram[3][246] ), .A2(n7094), .A3(n5243), .A4(n10061), 
        .Y(n1075) );
  AO22X1_HVT U1031 ( .A1(\ram[3][247] ), .A2(n7092), .A3(n5250), .A4(n10064), 
        .Y(n1076) );
  AO22X1_HVT U1032 ( .A1(\ram[3][248] ), .A2(n4307), .A3(n4516), .A4(n10068), 
        .Y(n1077) );
  AO22X1_HVT U1034 ( .A1(\ram[3][250] ), .A2(n7098), .A3(n5255), .A4(n10074), 
        .Y(n1079) );
  AO22X1_HVT U1035 ( .A1(\ram[3][251] ), .A2(n7097), .A3(n5273), .A4(n10077), 
        .Y(n1080) );
  AO22X1_HVT U1036 ( .A1(\ram[3][252] ), .A2(n7119), .A3(n4294), .A4(n10081), 
        .Y(n1081) );
  AO22X1_HVT U1037 ( .A1(\ram[3][253] ), .A2(n7118), .A3(n5273), .A4(n10084), 
        .Y(n1082) );
  AO22X1_HVT U1038 ( .A1(\ram[3][254] ), .A2(n7117), .A3(n6768), .A4(n10087), 
        .Y(n1083) );
  AO22X1_HVT U1039 ( .A1(\ram[3][255] ), .A2(n7116), .A3(n5267), .A4(n10090), 
        .Y(n1084) );
  AO22X1_HVT U1045 ( .A1(\ram[4][1] ), .A2(n6176), .A3(n6217), .A4(n9309), .Y(
        n1086) );
  AO22X1_HVT U1046 ( .A1(\ram[4][2] ), .A2(n4970), .A3(n6216), .A4(data[2]), 
        .Y(n1087) );
  AO22X1_HVT U1047 ( .A1(\ram[4][3] ), .A2(n6171), .A3(n6201), .A4(n9315), .Y(
        n1088) );
  AO22X1_HVT U1048 ( .A1(\ram[4][4] ), .A2(n6169), .A3(n6220), .A4(n9319), .Y(
        n1089) );
  AO22X1_HVT U1055 ( .A1(\ram[4][11] ), .A2(n6178), .A3(n6197), .A4(n9340), 
        .Y(n1096) );
  AO22X1_HVT U1057 ( .A1(\ram[4][13] ), .A2(n4395), .A3(n6201), .A4(n9347), 
        .Y(n1098) );
  AO22X1_HVT U1058 ( .A1(\ram[4][14] ), .A2(n6177), .A3(n6249), .A4(n9350), 
        .Y(n1099) );
  AO22X1_HVT U1059 ( .A1(\ram[4][15] ), .A2(n6177), .A3(n6195), .A4(n9353), 
        .Y(n1100) );
  AO22X1_HVT U1060 ( .A1(\ram[4][16] ), .A2(n6177), .A3(n6194), .A4(n9356), 
        .Y(n1101) );
  AO22X1_HVT U1061 ( .A1(\ram[4][17] ), .A2(n4968), .A3(n6191), .A4(n9359), 
        .Y(n1102) );
  AO22X1_HVT U1062 ( .A1(\ram[4][18] ), .A2(n6173), .A3(n6190), .A4(n9362), 
        .Y(n1103) );
  AO22X1_HVT U1063 ( .A1(\ram[4][19] ), .A2(n6171), .A3(n6189), .A4(n9365), 
        .Y(n1104) );
  AO22X1_HVT U1067 ( .A1(\ram[4][23] ), .A2(n4835), .A3(n6205), .A4(n9376), 
        .Y(n1108) );
  AO22X1_HVT U1068 ( .A1(\ram[4][24] ), .A2(n6181), .A3(n6203), .A4(n9379), 
        .Y(n1109) );
  AO22X1_HVT U1072 ( .A1(\ram[4][28] ), .A2(n6154), .A3(n6194), .A4(n9391), 
        .Y(n1113) );
  AO22X1_HVT U1074 ( .A1(\ram[4][30] ), .A2(n6181), .A3(n6211), .A4(n9397), 
        .Y(n1115) );
  AO22X1_HVT U1075 ( .A1(\ram[4][31] ), .A2(n6160), .A3(n6209), .A4(n9400), 
        .Y(n1116) );
  AO22X1_HVT U1076 ( .A1(\ram[4][32] ), .A2(n4706), .A3(n6208), .A4(n9403), 
        .Y(n1117) );
  AO22X1_HVT U1078 ( .A1(\ram[4][34] ), .A2(n6143), .A3(n6205), .A4(n9409), 
        .Y(n1119) );
  AO22X1_HVT U1079 ( .A1(\ram[4][35] ), .A2(n4961), .A3(n6203), .A4(n9412), 
        .Y(n1120) );
  AO22X1_HVT U1081 ( .A1(\ram[4][37] ), .A2(n6172), .A3(n10297), .A4(n9418), 
        .Y(n1122) );
  AO22X1_HVT U1082 ( .A1(\ram[4][38] ), .A2(n6146), .A3(n6217), .A4(n9421), 
        .Y(n1123) );
  AO22X1_HVT U1084 ( .A1(\ram[4][40] ), .A2(n5484), .A3(n6192), .A4(n9427), 
        .Y(n1125) );
  AO22X1_HVT U1085 ( .A1(\ram[4][41] ), .A2(n4965), .A3(n6246), .A4(n9430), 
        .Y(n1126) );
  AO22X1_HVT U1087 ( .A1(\ram[4][43] ), .A2(n4706), .A3(n6227), .A4(n9436), 
        .Y(n1128) );
  AO22X1_HVT U1088 ( .A1(\ram[4][44] ), .A2(n6170), .A3(n6189), .A4(n9439), 
        .Y(n1129) );
  AO22X1_HVT U1089 ( .A1(\ram[4][45] ), .A2(n6150), .A3(n6188), .A4(n9442), 
        .Y(n1130) );
  AO22X1_HVT U1090 ( .A1(\ram[4][46] ), .A2(n6178), .A3(n6187), .A4(n9445), 
        .Y(n1131) );
  AO22X1_HVT U1091 ( .A1(\ram[4][47] ), .A2(n6173), .A3(n6250), .A4(n9448), 
        .Y(n1132) );
  AO22X1_HVT U1093 ( .A1(\ram[4][49] ), .A2(n4439), .A3(n6245), .A4(n9454), 
        .Y(n1134) );
  AO22X1_HVT U1095 ( .A1(\ram[4][51] ), .A2(n6149), .A3(n6242), .A4(n9460), 
        .Y(n1136) );
  AO22X1_HVT U1099 ( .A1(\ram[4][55] ), .A2(n6182), .A3(n6236), .A4(n9472), 
        .Y(n1140) );
  AO22X1_HVT U1100 ( .A1(\ram[4][56] ), .A2(n4836), .A3(n6240), .A4(n9475), 
        .Y(n1141) );
  AO22X1_HVT U1101 ( .A1(\ram[4][57] ), .A2(n4370), .A3(n6237), .A4(n9478), 
        .Y(n1142) );
  AO22X1_HVT U1102 ( .A1(\ram[4][58] ), .A2(n4395), .A3(n6236), .A4(n9481), 
        .Y(n1143) );
  AO22X1_HVT U1104 ( .A1(\ram[4][60] ), .A2(n6154), .A3(n6211), .A4(n9487), 
        .Y(n1145) );
  AO22X1_HVT U1105 ( .A1(\ram[4][61] ), .A2(n6160), .A3(n6209), .A4(n9490), 
        .Y(n1146) );
  AO22X1_HVT U1107 ( .A1(\ram[4][63] ), .A2(n5484), .A3(n6206), .A4(n9496), 
        .Y(n1148) );
  AO22X1_HVT U1108 ( .A1(\ram[4][64] ), .A2(n6160), .A3(n6205), .A4(n9499), 
        .Y(n1149) );
  AO22X1_HVT U1109 ( .A1(\ram[4][65] ), .A2(n6171), .A3(n6203), .A4(n9502), 
        .Y(n1150) );
  AO22X1_HVT U1110 ( .A1(\ram[4][66] ), .A2(n5445), .A3(n6202), .A4(n9505), 
        .Y(n1151) );
  AO22X1_HVT U1112 ( .A1(\ram[4][68] ), .A2(n4823), .A3(n6206), .A4(n9511), 
        .Y(n1153) );
  AO22X1_HVT U1113 ( .A1(\ram[4][69] ), .A2(n6164), .A3(n6205), .A4(n9514), 
        .Y(n1154) );
  AO22X1_HVT U1114 ( .A1(\ram[4][70] ), .A2(n4370), .A3(n6203), .A4(n9517), 
        .Y(n1155) );
  AO22X1_HVT U1115 ( .A1(\ram[4][71] ), .A2(n6161), .A3(n6202), .A4(n9520), 
        .Y(n1156) );
  AO22X1_HVT U1116 ( .A1(\ram[4][72] ), .A2(n4928), .A3(n10296), .A4(n9523), 
        .Y(n1157) );
  AO22X1_HVT U1117 ( .A1(\ram[4][73] ), .A2(n4928), .A3(n6220), .A4(n9526), 
        .Y(n1158) );
  AO22X1_HVT U1118 ( .A1(\ram[4][74] ), .A2(n6151), .A3(n6193), .A4(n9529), 
        .Y(n1159) );
  AO22X1_HVT U1119 ( .A1(\ram[4][75] ), .A2(n6178), .A3(n6192), .A4(n9532), 
        .Y(n1160) );
  AO22X1_HVT U1120 ( .A1(\ram[4][76] ), .A2(n6174), .A3(n6245), .A4(n9535), 
        .Y(n1161) );
  AO22X1_HVT U1121 ( .A1(\ram[4][77] ), .A2(n5460), .A3(n6243), .A4(n9538), 
        .Y(n1162) );
  AO22X1_HVT U1122 ( .A1(\ram[4][78] ), .A2(n6149), .A3(n6242), .A4(n9541), 
        .Y(n1163) );
  AO22X1_HVT U1123 ( .A1(\ram[4][79] ), .A2(n6143), .A3(n6241), .A4(n9544), 
        .Y(n1164) );
  AO22X1_HVT U1124 ( .A1(\ram[4][80] ), .A2(n4823), .A3(n6214), .A4(n9547), 
        .Y(n1165) );
  AO22X1_HVT U1125 ( .A1(\ram[4][81] ), .A2(n6177), .A3(n6188), .A4(n9550), 
        .Y(n1166) );
  AO22X1_HVT U1126 ( .A1(\ram[4][82] ), .A2(n6179), .A3(n6187), .A4(n9553), 
        .Y(n1167) );
  AO22X1_HVT U1127 ( .A1(\ram[4][83] ), .A2(n6161), .A3(n6228), .A4(n9556), 
        .Y(n1168) );
  AO22X1_HVT U1128 ( .A1(\ram[4][84] ), .A2(n4370), .A3(n6227), .A4(n9559), 
        .Y(n1169) );
  AO22X1_HVT U1129 ( .A1(\ram[4][85] ), .A2(n5460), .A3(n6226), .A4(n9562), 
        .Y(n1170) );
  AO22X1_HVT U1130 ( .A1(\ram[4][86] ), .A2(n6168), .A3(n6223), .A4(n9565), 
        .Y(n1171) );
  AO22X1_HVT U1131 ( .A1(\ram[4][87] ), .A2(n5484), .A3(n6222), .A4(n9568), 
        .Y(n1172) );
  AO22X1_HVT U1132 ( .A1(\ram[4][88] ), .A2(n6179), .A3(n6220), .A4(n9571), 
        .Y(n1173) );
  AO22X1_HVT U1134 ( .A1(\ram[4][90] ), .A2(n6163), .A3(n6217), .A4(n9577), 
        .Y(n1175) );
  AO22X1_HVT U1135 ( .A1(\ram[4][91] ), .A2(n5460), .A3(n6216), .A4(n9580), 
        .Y(n1176) );
  AO22X1_HVT U1136 ( .A1(\ram[4][92] ), .A2(n5489), .A3(n6201), .A4(n9583), 
        .Y(n1177) );
  AO22X1_HVT U1137 ( .A1(\ram[4][93] ), .A2(n6174), .A3(n6200), .A4(n9586), 
        .Y(n1178) );
  AO22X1_HVT U1138 ( .A1(\ram[4][94] ), .A2(n6173), .A3(n6198), .A4(n9589), 
        .Y(n1179) );
  AO22X1_HVT U1139 ( .A1(\ram[4][95] ), .A2(n5060), .A3(n6222), .A4(n9592), 
        .Y(n1180) );
  AO22X1_HVT U1140 ( .A1(\ram[4][96] ), .A2(n6154), .A3(n6220), .A4(n9595), 
        .Y(n1181) );
  AO22X1_HVT U1141 ( .A1(\ram[4][97] ), .A2(n4836), .A3(n6241), .A4(n9598), 
        .Y(n1182) );
  AO22X1_HVT U1142 ( .A1(\ram[4][98] ), .A2(n6153), .A3(n6240), .A4(n9601), 
        .Y(n1183) );
  AO22X1_HVT U1143 ( .A1(\ram[4][99] ), .A2(n6181), .A3(n6237), .A4(n9604), 
        .Y(n1184) );
  AO22X1_HVT U1144 ( .A1(\ram[4][100] ), .A2(n6179), .A3(n6236), .A4(n9607), 
        .Y(n1185) );
  AO22X1_HVT U1145 ( .A1(\ram[4][101] ), .A2(n4835), .A3(n6234), .A4(n9610), 
        .Y(n1186) );
  AO22X1_HVT U1146 ( .A1(\ram[4][102] ), .A2(n6144), .A3(n6233), .A4(n9613), 
        .Y(n1187) );
  AO22X1_HVT U1147 ( .A1(\ram[4][103] ), .A2(n4970), .A3(n6231), .A4(n9616), 
        .Y(n1188) );
  AO22X1_HVT U1148 ( .A1(\ram[4][104] ), .A2(n6168), .A3(n6230), .A4(n9619), 
        .Y(n1189) );
  AO22X1_HVT U1149 ( .A1(\ram[4][105] ), .A2(n6153), .A3(n6188), .A4(n9622), 
        .Y(n1190) );
  AO22X1_HVT U1150 ( .A1(\ram[4][106] ), .A2(n6180), .A3(n6228), .A4(n9625), 
        .Y(n1191) );
  AO22X1_HVT U1151 ( .A1(\ram[4][107] ), .A2(n4835), .A3(n6227), .A4(n9628), 
        .Y(n1192) );
  AO22X1_HVT U1152 ( .A1(\ram[4][108] ), .A2(n6143), .A3(n6226), .A4(n9631), 
        .Y(n1193) );
  AO22X1_HVT U1153 ( .A1(\ram[4][109] ), .A2(n6179), .A3(n10294), .A4(n9634), 
        .Y(n1194) );
  AO22X1_HVT U1154 ( .A1(\ram[4][110] ), .A2(n4395), .A3(n6193), .A4(n9637), 
        .Y(n1195) );
  AO22X1_HVT U1155 ( .A1(\ram[4][111] ), .A2(n6180), .A3(n6192), .A4(n9640), 
        .Y(n1196) );
  AO22X1_HVT U1156 ( .A1(\ram[4][112] ), .A2(n6179), .A3(n6246), .A4(n9643), 
        .Y(n1197) );
  AO22X1_HVT U1157 ( .A1(\ram[4][113] ), .A2(n4706), .A3(n6245), .A4(n9646), 
        .Y(n1198) );
  AO22X1_HVT U1158 ( .A1(\ram[4][114] ), .A2(n5490), .A3(n6243), .A4(n9649), 
        .Y(n1199) );
  AO22X1_HVT U1159 ( .A1(\ram[4][115] ), .A2(n6176), .A3(n6242), .A4(n9652), 
        .Y(n1200) );
  AO22X1_HVT U1160 ( .A1(\ram[4][116] ), .A2(n5490), .A3(n6241), .A4(n9655), 
        .Y(n1201) );
  AO22X1_HVT U1161 ( .A1(\ram[4][117] ), .A2(n6173), .A3(n6240), .A4(n9658), 
        .Y(n1202) );
  AO22X1_HVT U1162 ( .A1(\ram[4][118] ), .A2(n6174), .A3(n6237), .A4(n9661), 
        .Y(n1203) );
  AO22X1_HVT U1163 ( .A1(\ram[4][119] ), .A2(n6172), .A3(n6246), .A4(n9664), 
        .Y(n1204) );
  AO22X1_HVT U1164 ( .A1(\ram[4][120] ), .A2(n6150), .A3(n6222), .A4(n9667), 
        .Y(n1205) );
  AO22X1_HVT U1166 ( .A1(\ram[4][122] ), .A2(n6153), .A3(n6219), .A4(n9673), 
        .Y(n1207) );
  AO22X1_HVT U1167 ( .A1(\ram[4][123] ), .A2(n6169), .A3(n6217), .A4(n9676), 
        .Y(n1208) );
  AO22X1_HVT U1168 ( .A1(\ram[4][124] ), .A2(n4961), .A3(n6216), .A4(n9679), 
        .Y(n1209) );
  AO22X1_HVT U1169 ( .A1(\ram[4][125] ), .A2(n5060), .A3(n6201), .A4(n9682), 
        .Y(n1210) );
  AO22X1_HVT U1170 ( .A1(\ram[4][126] ), .A2(n6153), .A3(n6200), .A4(n9685), 
        .Y(n1211) );
  AO22X1_HVT U1171 ( .A1(\ram[4][127] ), .A2(n4836), .A3(n6198), .A4(n9688), 
        .Y(n1212) );
  AO22X1_HVT U1172 ( .A1(\ram[4][128] ), .A2(n6151), .A3(n6197), .A4(n9691), 
        .Y(n1213) );
  AO22X1_HVT U1173 ( .A1(\ram[4][129] ), .A2(n5502), .A3(n6195), .A4(n9694), 
        .Y(n1214) );
  AO22X1_HVT U1174 ( .A1(\ram[4][130] ), .A2(n6168), .A3(n6192), .A4(n9697), 
        .Y(n1215) );
  AO22X1_HVT U1176 ( .A1(\ram[4][132] ), .A2(n6163), .A3(n6214), .A4(n9703), 
        .Y(n1217) );
  AO22X1_HVT U1177 ( .A1(\ram[4][133] ), .A2(n6176), .A3(n6212), .A4(n9706), 
        .Y(n1218) );
  AO22X1_HVT U1178 ( .A1(\ram[4][134] ), .A2(n6177), .A3(n6230), .A4(n9709), 
        .Y(n1219) );
  AO22X1_HVT U1179 ( .A1(\ram[4][135] ), .A2(n6148), .A3(n6190), .A4(n9712), 
        .Y(n1220) );
  AO22X1_HVT U1180 ( .A1(\ram[4][136] ), .A2(n6144), .A3(n6200), .A4(n9715), 
        .Y(n1221) );
  AO22X1_HVT U1181 ( .A1(\ram[4][137] ), .A2(n6167), .A3(n6198), .A4(n9718), 
        .Y(n1222) );
  AO22X1_HVT U1182 ( .A1(\ram[4][138] ), .A2(n6170), .A3(n6197), .A4(n9721), 
        .Y(n1223) );
  AO22X1_HVT U1184 ( .A1(\ram[4][140] ), .A2(n4395), .A3(n6228), .A4(n9728), 
        .Y(n1225) );
  AO22X1_HVT U1186 ( .A1(\ram[4][142] ), .A2(n6150), .A3(n6194), .A4(n9734), 
        .Y(n1227) );
  AO22X1_HVT U1187 ( .A1(\ram[4][143] ), .A2(n4928), .A3(n6191), .A4(n9737), 
        .Y(n1228) );
  AO22X1_HVT U1188 ( .A1(\ram[4][144] ), .A2(n4823), .A3(n6216), .A4(n9741), 
        .Y(n1229) );
  AO22X1_HVT U1190 ( .A1(\ram[4][146] ), .A2(n4706), .A3(n10291), .A4(n9747), 
        .Y(n1231) );
  AO22X1_HVT U1191 ( .A1(\ram[4][147] ), .A2(n5489), .A3(n6194), .A4(n9750), 
        .Y(n1232) );
  AO22X1_HVT U1192 ( .A1(\ram[4][148] ), .A2(n6168), .A3(n6191), .A4(n9754), 
        .Y(n1233) );
  AO22X1_HVT U1193 ( .A1(\ram[4][149] ), .A2(n6146), .A3(n6190), .A4(n9757), 
        .Y(n1234) );
  AO22X1_HVT U1194 ( .A1(\ram[4][150] ), .A2(n4927), .A3(n6189), .A4(n9760), 
        .Y(n1235) );
  AO22X1_HVT U1195 ( .A1(\ram[4][151] ), .A2(n6148), .A3(n6188), .A4(n9763), 
        .Y(n1236) );
  AO22X1_HVT U1196 ( .A1(\ram[4][152] ), .A2(n5502), .A3(n6187), .A4(n9766), 
        .Y(n1237) );
  AO22X1_HVT U1197 ( .A1(\ram[4][153] ), .A2(n5460), .A3(n6250), .A4(n9769), 
        .Y(n1238) );
  AO22X1_HVT U1198 ( .A1(\ram[4][154] ), .A2(n6167), .A3(n6249), .A4(n9772), 
        .Y(n1239) );
  AO22X1_HVT U1199 ( .A1(\ram[4][155] ), .A2(n6170), .A3(n6215), .A4(n9775), 
        .Y(n1240) );
  AO22X1_HVT U1200 ( .A1(\ram[4][156] ), .A2(n6160), .A3(n6217), .A4(n9779), 
        .Y(n1241) );
  AO22X1_HVT U1201 ( .A1(\ram[4][157] ), .A2(n4968), .A3(n6216), .A4(n9782), 
        .Y(n1242) );
  AO22X1_HVT U1202 ( .A1(\ram[4][158] ), .A2(n6155), .A3(n6201), .A4(n9785), 
        .Y(n1243) );
  AO22X1_HVT U1203 ( .A1(\ram[4][159] ), .A2(n5484), .A3(n6200), .A4(n9788), 
        .Y(n1244) );
  AO22X1_HVT U1204 ( .A1(\ram[4][160] ), .A2(n6178), .A3(n6198), .A4(n9792), 
        .Y(n1245) );
  AO22X1_HVT U1205 ( .A1(\ram[4][161] ), .A2(n6154), .A3(n6197), .A4(n9795), 
        .Y(n1246) );
  AO22X1_HVT U1206 ( .A1(\ram[4][162] ), .A2(n4968), .A3(n6195), .A4(n9798), 
        .Y(n1247) );
  AO22X1_HVT U1207 ( .A1(\ram[4][163] ), .A2(n6180), .A3(n6211), .A4(n9801), 
        .Y(n1248) );
  AO22X1_HVT U1208 ( .A1(\ram[4][164] ), .A2(n6161), .A3(n6209), .A4(n9804), 
        .Y(n1249) );
  AO22X1_HVT U1209 ( .A1(\ram[4][165] ), .A2(n6151), .A3(n6208), .A4(n9807), 
        .Y(n1250) );
  AO22X1_HVT U1210 ( .A1(\ram[4][166] ), .A2(n6151), .A3(n6206), .A4(n9810), 
        .Y(n1251) );
  AO22X1_HVT U1211 ( .A1(\ram[4][167] ), .A2(n6164), .A3(n6250), .A4(n9813), 
        .Y(n1252) );
  AO22X1_HVT U1212 ( .A1(\ram[4][168] ), .A2(n6144), .A3(n6220), .A4(n9816), 
        .Y(n1253) );
  AO22X1_HVT U1213 ( .A1(\ram[4][169] ), .A2(n6149), .A3(n6234), .A4(n9819), 
        .Y(n1254) );
  AO22X1_HVT U1214 ( .A1(\ram[4][170] ), .A2(n4965), .A3(n6233), .A4(n9822), 
        .Y(n1255) );
  AO22X1_HVT U1215 ( .A1(\ram[4][171] ), .A2(n6146), .A3(n6231), .A4(n9825), 
        .Y(n1256) );
  AO22X1_HVT U1216 ( .A1(\ram[4][172] ), .A2(n6149), .A3(n6230), .A4(n9829), 
        .Y(n1257) );
  AO22X1_HVT U1217 ( .A1(\ram[4][173] ), .A2(n6143), .A3(n6188), .A4(n9832), 
        .Y(n1258) );
  AO22X1_HVT U1218 ( .A1(\ram[4][174] ), .A2(n6181), .A3(n6228), .A4(n9835), 
        .Y(n1259) );
  AO22X1_HVT U1219 ( .A1(\ram[4][175] ), .A2(n6180), .A3(n6227), .A4(n9838), 
        .Y(n1260) );
  AO22X1_HVT U1221 ( .A1(\ram[4][177] ), .A2(n4823), .A3(n6223), .A4(n9845), 
        .Y(n1262) );
  AO22X1_HVT U1222 ( .A1(\ram[4][178] ), .A2(n6148), .A3(n6222), .A4(n9848), 
        .Y(n1263) );
  AO22X1_HVT U1223 ( .A1(\ram[4][179] ), .A2(n4836), .A3(n6219), .A4(n9851), 
        .Y(n1264) );
  AO22X1_HVT U1224 ( .A1(\ram[4][180] ), .A2(n6174), .A3(n6231), .A4(n9855), 
        .Y(n1265) );
  AO22X1_HVT U1225 ( .A1(\ram[4][181] ), .A2(n6169), .A3(n6236), .A4(n9858), 
        .Y(n1266) );
  AO22X1_HVT U1226 ( .A1(\ram[4][182] ), .A2(n6170), .A3(n6234), .A4(n9861), 
        .Y(n1267) );
  AO22X1_HVT U1227 ( .A1(\ram[4][183] ), .A2(n6170), .A3(n6233), .A4(n9864), 
        .Y(n1268) );
  AO22X1_HVT U1228 ( .A1(\ram[4][184] ), .A2(n4970), .A3(n6231), .A4(n9868), 
        .Y(n1269) );
  AO22X1_HVT U1229 ( .A1(\ram[4][185] ), .A2(n6144), .A3(n6230), .A4(n9871), 
        .Y(n1270) );
  AO22X1_HVT U1230 ( .A1(\ram[4][186] ), .A2(n6146), .A3(n6190), .A4(n9874), 
        .Y(n1271) );
  AO22X1_HVT U1231 ( .A1(\ram[4][187] ), .A2(n4370), .A3(n6228), .A4(n9877), 
        .Y(n1272) );
  AO22X1_HVT U1232 ( .A1(\ram[4][188] ), .A2(n6162), .A3(n6227), .A4(n9880), 
        .Y(n1273) );
  AO22X1_HVT U1233 ( .A1(\ram[4][189] ), .A2(n6163), .A3(n6226), .A4(n9883), 
        .Y(n1274) );
  AO22X1_HVT U1234 ( .A1(\ram[4][190] ), .A2(n5502), .A3(n6223), .A4(n9886), 
        .Y(n1275) );
  AO22X1_HVT U1235 ( .A1(\ram[4][191] ), .A2(n6161), .A3(n6222), .A4(n9889), 
        .Y(n1276) );
  AO22X1_HVT U1236 ( .A1(\ram[4][192] ), .A2(n6177), .A3(n6249), .A4(n9893), 
        .Y(n1277) );
  AO22X1_HVT U1237 ( .A1(\ram[4][193] ), .A2(n6157), .A3(n6215), .A4(n9896), 
        .Y(n1278) );
  AO22X1_HVT U1238 ( .A1(\ram[4][194] ), .A2(n4910), .A3(n6214), .A4(n9899), 
        .Y(n1279) );
  AO22X1_HVT U1240 ( .A1(\ram[4][196] ), .A2(n5060), .A3(n6211), .A4(n9906), 
        .Y(n1281) );
  AO22X1_HVT U1241 ( .A1(\ram[4][197] ), .A2(n5502), .A3(n6209), .A4(n9909), 
        .Y(n1282) );
  AO22X1_HVT U1242 ( .A1(\ram[4][198] ), .A2(n6178), .A3(n6208), .A4(n9912), 
        .Y(n1283) );
  AO22X1_HVT U1244 ( .A1(\ram[4][200] ), .A2(n6157), .A3(n6194), .A4(n9919), 
        .Y(n1285) );
  AO22X1_HVT U1245 ( .A1(\ram[4][201] ), .A2(n4910), .A3(n6191), .A4(n9922), 
        .Y(n1286) );
  AO22X1_HVT U1246 ( .A1(\ram[4][202] ), .A2(n6161), .A3(n6190), .A4(n9925), 
        .Y(n1287) );
  AO22X1_HVT U1247 ( .A1(\ram[4][203] ), .A2(n6144), .A3(n6189), .A4(n9928), 
        .Y(n1288) );
  AO22X1_HVT U1248 ( .A1(\ram[4][204] ), .A2(n6169), .A3(n6188), .A4(n9931), 
        .Y(n1289) );
  AO22X1_HVT U1249 ( .A1(\ram[4][205] ), .A2(n6172), .A3(n6187), .A4(n9934), 
        .Y(n1290) );
  AO22X1_HVT U1250 ( .A1(\ram[4][206] ), .A2(n6162), .A3(n6250), .A4(n9937), 
        .Y(n1291) );
  AO22X1_HVT U1251 ( .A1(\ram[4][207] ), .A2(n6168), .A3(n6249), .A4(n9940), 
        .Y(n1292) );
  AO22X1_HVT U1252 ( .A1(\ram[4][208] ), .A2(n4835), .A3(n6215), .A4(n9944), 
        .Y(n1293) );
  AO22X1_HVT U1254 ( .A1(\ram[4][210] ), .A2(n5460), .A3(n6249), .A4(n9950), 
        .Y(n1295) );
  AO22X1_HVT U1255 ( .A1(\ram[4][211] ), .A2(n6162), .A3(n6215), .A4(n9953), 
        .Y(n1296) );
  AO22X1_HVT U1256 ( .A1(\ram[4][212] ), .A2(n5060), .A3(n6214), .A4(n9956), 
        .Y(n1297) );
  AO22X1_HVT U1258 ( .A1(\ram[4][214] ), .A2(n6176), .A3(n6211), .A4(n9962), 
        .Y(n1299) );
  AO22X1_HVT U1260 ( .A1(\ram[4][216] ), .A2(n6161), .A3(n6208), .A4(n9968), 
        .Y(n1301) );
  AO22X1_HVT U1261 ( .A1(\ram[4][217] ), .A2(n6160), .A3(n6243), .A4(n9971), 
        .Y(n1302) );
  AO22X1_HVT U1262 ( .A1(\ram[4][218] ), .A2(n6172), .A3(n6193), .A4(n9974), 
        .Y(n1303) );
  AO22X1_HVT U1263 ( .A1(\ram[4][219] ), .A2(n5484), .A3(n6192), .A4(n9977), 
        .Y(n1304) );
  AO22X1_HVT U1264 ( .A1(\ram[4][220] ), .A2(n6157), .A3(n6246), .A4(n9981), 
        .Y(n1305) );
  AO22X1_HVT U1265 ( .A1(\ram[4][221] ), .A2(n6156), .A3(n6215), .A4(n9984), 
        .Y(n1306) );
  AO22X1_HVT U1266 ( .A1(\ram[4][222] ), .A2(n4965), .A3(n6190), .A4(n9987), 
        .Y(n1307) );
  AO22X1_HVT U1267 ( .A1(\ram[4][223] ), .A2(n6146), .A3(n6189), .A4(n9990), 
        .Y(n1308) );
  AO22X1_HVT U1268 ( .A1(\ram[4][224] ), .A2(n4439), .A3(n6245), .A4(n9993), 
        .Y(n1309) );
  AO22X1_HVT U1269 ( .A1(\ram[4][225] ), .A2(n6182), .A3(n6243), .A4(n9996), 
        .Y(n1310) );
  AO22X1_HVT U1270 ( .A1(\ram[4][226] ), .A2(n6157), .A3(n6242), .A4(n9999), 
        .Y(n1311) );
  AO22X1_HVT U1271 ( .A1(\ram[4][227] ), .A2(n6156), .A3(n6241), .A4(n10002), 
        .Y(n1312) );
  AO22X1_HVT U1272 ( .A1(\ram[4][228] ), .A2(n5060), .A3(n6240), .A4(n10005), 
        .Y(n1313) );
  AO22X1_HVT U1273 ( .A1(\ram[4][229] ), .A2(n6164), .A3(n6237), .A4(n10008), 
        .Y(n1314) );
  AO22X1_HVT U1274 ( .A1(\ram[4][230] ), .A2(n6163), .A3(n6236), .A4(n10011), 
        .Y(n1315) );
  AO22X1_HVT U1275 ( .A1(\ram[4][231] ), .A2(n6182), .A3(n6234), .A4(n10014), 
        .Y(n1316) );
  AO22X1_HVT U1276 ( .A1(\ram[4][232] ), .A2(n6180), .A3(n6233), .A4(n10018), 
        .Y(n1317) );
  AO22X1_HVT U1277 ( .A1(\ram[4][233] ), .A2(n6178), .A3(n6231), .A4(n10021), 
        .Y(n1318) );
  AO22X1_HVT U1278 ( .A1(\ram[4][234] ), .A2(n5490), .A3(n6230), .A4(n10024), 
        .Y(n1319) );
  AO22X1_HVT U1279 ( .A1(\ram[4][235] ), .A2(n4910), .A3(n6189), .A4(n10027), 
        .Y(n1320) );
  AO22X1_HVT U1280 ( .A1(\ram[4][236] ), .A2(n6182), .A3(n6226), .A4(n10030), 
        .Y(n1321) );
  AO22X1_HVT U1281 ( .A1(\ram[4][237] ), .A2(n6181), .A3(n6223), .A4(n10033), 
        .Y(n1322) );
  AO22X1_HVT U1282 ( .A1(\ram[4][238] ), .A2(n4439), .A3(n6206), .A4(n10036), 
        .Y(n1323) );
  AO22X1_HVT U1283 ( .A1(\ram[4][239] ), .A2(n4961), .A3(n6205), .A4(n10039), 
        .Y(n1324) );
  AO22X1_HVT U1284 ( .A1(\ram[4][240] ), .A2(n5445), .A3(n6203), .A4(n10043), 
        .Y(n1325) );
  AO22X1_HVT U1285 ( .A1(\ram[4][241] ), .A2(n6151), .A3(n6202), .A4(n10046), 
        .Y(n1326) );
  AO22X1_HVT U1286 ( .A1(\ram[4][242] ), .A2(n6167), .A3(n10297), .A4(n10049), 
        .Y(n1327) );
  AO22X1_HVT U1287 ( .A1(\ram[4][243] ), .A2(n6146), .A3(n6212), .A4(n10052), 
        .Y(n1328) );
  AO22X1_HVT U1288 ( .A1(\ram[4][244] ), .A2(n4927), .A3(n6193), .A4(n10055), 
        .Y(n1329) );
  AO22X1_HVT U1289 ( .A1(\ram[4][245] ), .A2(n6162), .A3(n6192), .A4(n10058), 
        .Y(n1330) );
  AO22X1_HVT U1290 ( .A1(\ram[4][246] ), .A2(n6174), .A3(n6246), .A4(n10061), 
        .Y(n1331) );
  AO22X1_HVT U1291 ( .A1(\ram[4][247] ), .A2(n6156), .A3(n6245), .A4(n10064), 
        .Y(n1332) );
  AO22X1_HVT U1292 ( .A1(\ram[4][248] ), .A2(n6148), .A3(n6243), .A4(n10068), 
        .Y(n1333) );
  AO22X1_HVT U1293 ( .A1(\ram[4][249] ), .A2(n5490), .A3(n6242), .A4(n10071), 
        .Y(n1334) );
  AO22X1_HVT U1294 ( .A1(\ram[4][250] ), .A2(n4927), .A3(n6214), .A4(n10074), 
        .Y(n1335) );
  AO22X1_HVT U1295 ( .A1(\ram[4][251] ), .A2(n6167), .A3(n6212), .A4(n10077), 
        .Y(n1336) );
  AO22X1_HVT U1296 ( .A1(\ram[4][252] ), .A2(n6167), .A3(n6187), .A4(n10081), 
        .Y(n1337) );
  AO22X1_HVT U1297 ( .A1(\ram[4][253] ), .A2(n4965), .A3(n6197), .A4(n10084), 
        .Y(n1338) );
  AO22X1_HVT U1298 ( .A1(\ram[4][254] ), .A2(n6146), .A3(n6195), .A4(n10087), 
        .Y(n1339) );
  AO22X1_HVT U1299 ( .A1(\ram[4][255] ), .A2(n4970), .A3(n6223), .A4(n10090), 
        .Y(n1340) );
  AND2X1_HVT U1302 ( .A1(n9), .A2(n5880), .Y(n24) );
  AO22X1_HVT U1303 ( .A1(\ram[5][0] ), .A2(n4938), .A3(n9286), .A4(n9306), .Y(
        n1341) );
  AO22X1_HVT U1304 ( .A1(\ram[5][1] ), .A2(n4897), .A3(n9262), .A4(n9309), .Y(
        n1342) );
  AO22X1_HVT U1308 ( .A1(\ram[5][5] ), .A2(n4954), .A3(n9283), .A4(n9322), .Y(
        n1346) );
  AO22X1_HVT U1310 ( .A1(\ram[5][7] ), .A2(n5710), .A3(n9281), .A4(n9328), .Y(
        n1348) );
  AO22X1_HVT U1312 ( .A1(\ram[5][9] ), .A2(n4795), .A3(n9272), .A4(n9334), .Y(
        n1350) );
  AO22X1_HVT U1314 ( .A1(\ram[5][11] ), .A2(n4838), .A3(n4692), .A4(n9340), 
        .Y(n1352) );
  AO22X1_HVT U1322 ( .A1(\ram[5][19] ), .A2(n4952), .A3(n4646), .A4(n9365), 
        .Y(n1360) );
  AO22X1_HVT U1324 ( .A1(\ram[5][21] ), .A2(n5695), .A3(n4271), .A4(n9370), 
        .Y(n1362) );
  AO22X1_HVT U1325 ( .A1(\ram[5][22] ), .A2(n4529), .A3(n9286), .A4(n9373), 
        .Y(n1363) );
  AO22X1_HVT U1326 ( .A1(\ram[5][23] ), .A2(n5693), .A3(n4646), .A4(n9376), 
        .Y(n1364) );
  AO22X1_HVT U1327 ( .A1(\ram[5][24] ), .A2(n4256), .A3(n9295), .A4(n9379), 
        .Y(n1365) );
  AO22X1_HVT U1328 ( .A1(\ram[5][25] ), .A2(n5701), .A3(n9294), .A4(n9382), 
        .Y(n1366) );
  AO22X1_HVT U1329 ( .A1(\ram[5][26] ), .A2(n4765), .A3(n9293), .A4(n9385), 
        .Y(n1367) );
  AO22X1_HVT U1330 ( .A1(\ram[5][27] ), .A2(n4231), .A3(n9292), .A4(n9388), 
        .Y(n1368) );
  AO22X1_HVT U1334 ( .A1(\ram[5][31] ), .A2(n4915), .A3(n9292), .A4(n9400), 
        .Y(n1372) );
  AO22X1_HVT U1335 ( .A1(\ram[5][32] ), .A2(n4850), .A3(n9290), .A4(n9403), 
        .Y(n1373) );
  AO22X1_HVT U1336 ( .A1(\ram[5][33] ), .A2(n5701), .A3(n9289), .A4(n9406), 
        .Y(n1374) );
  AO22X1_HVT U1338 ( .A1(\ram[5][35] ), .A2(n4896), .A3(n9290), .A4(n9412), 
        .Y(n1376) );
  AO22X1_HVT U1340 ( .A1(\ram[5][37] ), .A2(n5677), .A3(n4691), .A4(n9418), 
        .Y(n1378) );
  AO22X1_HVT U1342 ( .A1(\ram[5][39] ), .A2(n5693), .A3(n9276), .A4(n9424), 
        .Y(n1380) );
  AO22X1_HVT U1343 ( .A1(\ram[5][40] ), .A2(n5686), .A3(n9265), .A4(n9427), 
        .Y(n1381) );
  AO22X1_HVT U1344 ( .A1(\ram[5][41] ), .A2(n4937), .A3(n4695), .A4(n9430), 
        .Y(n1382) );
  AO22X1_HVT U1345 ( .A1(\ram[5][42] ), .A2(n5678), .A3(n9265), .A4(n9433), 
        .Y(n1383) );
  AO22X1_HVT U1346 ( .A1(\ram[5][43] ), .A2(n5696), .A3(n9267), .A4(n9436), 
        .Y(n1384) );
  AO22X1_HVT U1347 ( .A1(\ram[5][44] ), .A2(n4954), .A3(n9256), .A4(n9439), 
        .Y(n1385) );
  AO22X1_HVT U1348 ( .A1(\ram[5][45] ), .A2(n5690), .A3(n9302), .A4(n9442), 
        .Y(n1386) );
  AO22X1_HVT U1349 ( .A1(\ram[5][46] ), .A2(n5686), .A3(n9262), .A4(n9445), 
        .Y(n1387) );
  AO22X1_HVT U1355 ( .A1(\ram[5][52] ), .A2(n5683), .A3(n9273), .A4(n9463), 
        .Y(n1393) );
  AO22X1_HVT U1356 ( .A1(\ram[5][53] ), .A2(n4850), .A3(n9266), .A4(n9466), 
        .Y(n1394) );
  AO22X1_HVT U1357 ( .A1(\ram[5][54] ), .A2(n4938), .A3(n9271), .A4(n9469), 
        .Y(n1395) );
  AO22X1_HVT U1358 ( .A1(\ram[5][55] ), .A2(n5709), .A3(n4691), .A4(n9472), 
        .Y(n1396) );
  AO22X1_HVT U1359 ( .A1(\ram[5][56] ), .A2(n5684), .A3(n4702), .A4(n9475), 
        .Y(n1397) );
  AO22X1_HVT U1360 ( .A1(\ram[5][57] ), .A2(n4728), .A3(n9302), .A4(n9478), 
        .Y(n1398) );
  AO22X1_HVT U1361 ( .A1(\ram[5][58] ), .A2(n4795), .A3(n9303), .A4(n9481), 
        .Y(n1399) );
  AO22X1_HVT U1362 ( .A1(\ram[5][59] ), .A2(n4210), .A3(n9302), .A4(n9484), 
        .Y(n1400) );
  AO22X1_HVT U1363 ( .A1(\ram[5][60] ), .A2(n4210), .A3(n4695), .A4(n9487), 
        .Y(n1401) );
  AO22X1_HVT U1364 ( .A1(\ram[5][61] ), .A2(n4331), .A3(n9272), .A4(n9490), 
        .Y(n1402) );
  AO22X1_HVT U1366 ( .A1(\ram[5][63] ), .A2(n4732), .A3(n9277), .A4(n9496), 
        .Y(n1404) );
  AO22X1_HVT U1367 ( .A1(\ram[5][64] ), .A2(n5678), .A3(n9256), .A4(n9499), 
        .Y(n1405) );
  AO22X1_HVT U1369 ( .A1(\ram[5][66] ), .A2(n5712), .A3(n4689), .A4(n9505), 
        .Y(n1407) );
  AO22X1_HVT U1370 ( .A1(\ram[5][67] ), .A2(n5672), .A3(n9259), .A4(n9508), 
        .Y(n1408) );
  AO22X1_HVT U1372 ( .A1(\ram[5][69] ), .A2(n4773), .A3(n9283), .A4(n9514), 
        .Y(n1410) );
  AO22X1_HVT U1373 ( .A1(\ram[5][70] ), .A2(n5694), .A3(n9282), .A4(n9517), 
        .Y(n1411) );
  AO22X1_HVT U1374 ( .A1(\ram[5][71] ), .A2(n5669), .A3(n9281), .A4(n9520), 
        .Y(n1412) );
  AO22X1_HVT U1375 ( .A1(\ram[5][72] ), .A2(n5672), .A3(n9255), .A4(n9523), 
        .Y(n1413) );
  AO22X1_HVT U1376 ( .A1(\ram[5][73] ), .A2(n5687), .A3(n4422), .A4(n9526), 
        .Y(n1414) );
  AO22X1_HVT U1377 ( .A1(\ram[5][74] ), .A2(n4938), .A3(n9255), .A4(n9529), 
        .Y(n1415) );
  AO22X1_HVT U1378 ( .A1(\ram[5][75] ), .A2(n5686), .A3(n4271), .A4(n9532), 
        .Y(n1416) );
  AO22X1_HVT U1379 ( .A1(\ram[5][76] ), .A2(n4764), .A3(n9284), .A4(n9535), 
        .Y(n1417) );
  AO22X1_HVT U1380 ( .A1(\ram[5][77] ), .A2(n5685), .A3(n9283), .A4(n9538), 
        .Y(n1418) );
  AO22X1_HVT U1381 ( .A1(\ram[5][78] ), .A2(n5695), .A3(n9282), .A4(n9541), 
        .Y(n1419) );
  AO22X1_HVT U1382 ( .A1(\ram[5][79] ), .A2(n5671), .A3(n9281), .A4(n9544), 
        .Y(n1420) );
  AO22X1_HVT U1383 ( .A1(\ram[5][80] ), .A2(n5690), .A3(n4410), .A4(n9547), 
        .Y(n1421) );
  AO22X1_HVT U1384 ( .A1(\ram[5][81] ), .A2(n5677), .A3(n9290), .A4(n9550), 
        .Y(n1422) );
  AO22X1_HVT U1385 ( .A1(\ram[5][82] ), .A2(n5710), .A3(n5011), .A4(n9553), 
        .Y(n1423) );
  AO22X1_HVT U1386 ( .A1(\ram[5][83] ), .A2(n5684), .A3(n9290), .A4(n9556), 
        .Y(n1424) );
  AO22X1_HVT U1387 ( .A1(\ram[5][84] ), .A2(n4628), .A3(n9262), .A4(n9559), 
        .Y(n1425) );
  AO22X1_HVT U1388 ( .A1(\ram[5][85] ), .A2(n5678), .A3(n9261), .A4(n9562), 
        .Y(n1426) );
  AO22X1_HVT U1389 ( .A1(\ram[5][86] ), .A2(n5703), .A3(n4689), .A4(n9565), 
        .Y(n1427) );
  AO22X1_HVT U1390 ( .A1(\ram[5][87] ), .A2(n5672), .A3(n9259), .A4(n9568), 
        .Y(n1428) );
  AO22X1_HVT U1391 ( .A1(\ram[5][88] ), .A2(n5685), .A3(n9285), .A4(n9571), 
        .Y(n1429) );
  AO22X1_HVT U1392 ( .A1(\ram[5][89] ), .A2(n5713), .A3(n9291), .A4(n9574), 
        .Y(n1430) );
  AO22X1_HVT U1393 ( .A1(\ram[5][90] ), .A2(n4917), .A3(n9286), .A4(n9577), 
        .Y(n1431) );
  AO22X1_HVT U1395 ( .A1(\ram[5][92] ), .A2(n5670), .A3(n9284), .A4(n9583), 
        .Y(n1433) );
  AO22X1_HVT U1396 ( .A1(\ram[5][93] ), .A2(n5690), .A3(n9283), .A4(n9586), 
        .Y(n1434) );
  AO22X1_HVT U1397 ( .A1(\ram[5][94] ), .A2(n5691), .A3(n9282), .A4(n9589), 
        .Y(n1435) );
  AO22X1_HVT U1398 ( .A1(\ram[5][95] ), .A2(n4813), .A3(n9281), .A4(n9592), 
        .Y(n1436) );
  AO22X1_HVT U1399 ( .A1(\ram[5][96] ), .A2(n5713), .A3(n9256), .A4(n9595), 
        .Y(n1437) );
  AO22X1_HVT U1401 ( .A1(\ram[5][98] ), .A2(n5675), .A3(n9256), .A4(n9601), 
        .Y(n1439) );
  AO22X1_HVT U1402 ( .A1(\ram[5][99] ), .A2(n4742), .A3(n4271), .A4(n9604), 
        .Y(n1440) );
  AO22X1_HVT U1403 ( .A1(\ram[5][100] ), .A2(n4626), .A3(n4702), .A4(n9607), 
        .Y(n1441) );
  AO22X1_HVT U1404 ( .A1(\ram[5][101] ), .A2(n5671), .A3(n9302), .A4(n9610), 
        .Y(n1442) );
  AO22X1_HVT U1405 ( .A1(\ram[5][102] ), .A2(n5703), .A3(n9304), .A4(n9613), 
        .Y(n1443) );
  AO22X1_HVT U1406 ( .A1(\ram[5][103] ), .A2(n4742), .A3(n9303), .A4(n9616), 
        .Y(n1444) );
  AO22X1_HVT U1407 ( .A1(\ram[5][104] ), .A2(n4838), .A3(n4701), .A4(n9619), 
        .Y(n1445) );
  AO22X1_HVT U1408 ( .A1(\ram[5][105] ), .A2(n4917), .A3(n9301), .A4(n9622), 
        .Y(n1446) );
  AO22X1_HVT U1409 ( .A1(\ram[5][106] ), .A2(n5676), .A3(n9300), .A4(n9625), 
        .Y(n1447) );
  AO22X1_HVT U1410 ( .A1(\ram[5][107] ), .A2(n4938), .A3(n9301), .A4(n9628), 
        .Y(n1448) );
  AO22X1_HVT U1411 ( .A1(\ram[5][108] ), .A2(n5685), .A3(n4646), .A4(n9631), 
        .Y(n1449) );
  AO22X1_HVT U1413 ( .A1(\ram[5][110] ), .A2(n5687), .A3(n9286), .A4(n9637), 
        .Y(n1451) );
  AO22X1_HVT U1414 ( .A1(\ram[5][111] ), .A2(n4749), .A3(n4646), .A4(n9640), 
        .Y(n1452) );
  AO22X1_HVT U1415 ( .A1(\ram[5][112] ), .A2(n5683), .A3(n9266), .A4(n9643), 
        .Y(n1453) );
  AO22X1_HVT U1416 ( .A1(\ram[5][113] ), .A2(n5669), .A3(n4695), .A4(n9646), 
        .Y(n1454) );
  AO22X1_HVT U1417 ( .A1(\ram[5][114] ), .A2(n5687), .A3(n9270), .A4(n9649), 
        .Y(n1455) );
  AO22X1_HVT U1418 ( .A1(\ram[5][115] ), .A2(n5707), .A3(n9270), .A4(n9652), 
        .Y(n1456) );
  AO22X1_HVT U1419 ( .A1(\ram[5][116] ), .A2(n5713), .A3(n4702), .A4(n9655), 
        .Y(n1457) );
  AO22X1_HVT U1420 ( .A1(\ram[5][117] ), .A2(n4626), .A3(n9303), .A4(n9658), 
        .Y(n1458) );
  AO22X1_HVT U1421 ( .A1(\ram[5][118] ), .A2(n4626), .A3(n9304), .A4(n9661), 
        .Y(n1459) );
  AO22X1_HVT U1422 ( .A1(\ram[5][119] ), .A2(n4813), .A3(n9304), .A4(n9664), 
        .Y(n1460) );
  AO22X1_HVT U1424 ( .A1(\ram[5][121] ), .A2(n5675), .A3(n9290), .A4(n9670), 
        .Y(n1462) );
  AO22X1_HVT U1426 ( .A1(\ram[5][123] ), .A2(n4896), .A3(n9291), .A4(n9676), 
        .Y(n1464) );
  AO22X1_HVT U1427 ( .A1(\ram[5][124] ), .A2(n5694), .A3(n9265), .A4(n9679), 
        .Y(n1465) );
  AO22X1_HVT U1428 ( .A1(\ram[5][125] ), .A2(n5703), .A3(n9266), .A4(n9682), 
        .Y(n1466) );
  AO22X1_HVT U1429 ( .A1(\ram[5][126] ), .A2(n4728), .A3(n4692), .A4(n9685), 
        .Y(n1467) );
  AO22X1_HVT U1430 ( .A1(\ram[5][127] ), .A2(n5710), .A3(n9267), .A4(n9688), 
        .Y(n1468) );
  AO22X1_HVT U1431 ( .A1(\ram[5][128] ), .A2(n5697), .A3(n4702), .A4(n9691), 
        .Y(n1469) );
  AO22X1_HVT U1432 ( .A1(\ram[5][129] ), .A2(n5677), .A3(n9302), .A4(n9694), 
        .Y(n1470) );
  AO22X1_HVT U1433 ( .A1(\ram[5][130] ), .A2(n4321), .A3(n9304), .A4(n9697), 
        .Y(n1471) );
  AO22X1_HVT U1434 ( .A1(\ram[5][131] ), .A2(n5662), .A3(n4422), .A4(n9700), 
        .Y(n1472) );
  AO22X1_HVT U1435 ( .A1(\ram[5][132] ), .A2(n5672), .A3(n9264), .A4(n9703), 
        .Y(n1473) );
  AO22X1_HVT U1436 ( .A1(\ram[5][133] ), .A2(n4917), .A3(n9273), .A4(n9706), 
        .Y(n1474) );
  AO22X1_HVT U1437 ( .A1(\ram[5][134] ), .A2(n5675), .A3(n9267), .A4(n9709), 
        .Y(n1475) );
  AO22X1_HVT U1438 ( .A1(\ram[5][135] ), .A2(n4838), .A3(n9264), .A4(n9712), 
        .Y(n1476) );
  AO22X1_HVT U1439 ( .A1(\ram[5][136] ), .A2(n4915), .A3(n9262), .A4(n9715), 
        .Y(n1477) );
  AO22X1_HVT U1440 ( .A1(\ram[5][137] ), .A2(n5675), .A3(n9261), .A4(n9718), 
        .Y(n1478) );
  AO22X1_HVT U1441 ( .A1(\ram[5][138] ), .A2(n4321), .A3(n9260), .A4(n9721), 
        .Y(n1479) );
  AO22X1_HVT U1442 ( .A1(\ram[5][139] ), .A2(n5696), .A3(n9259), .A4(n9724), 
        .Y(n1480) );
  AO22X1_HVT U1443 ( .A1(\ram[5][140] ), .A2(n5671), .A3(n9286), .A4(n9728), 
        .Y(n1481) );
  AO22X1_HVT U1444 ( .A1(\ram[5][141] ), .A2(n5670), .A3(n4830), .A4(n9731), 
        .Y(n1482) );
  AO22X1_HVT U1445 ( .A1(\ram[5][142] ), .A2(n4628), .A3(n9286), .A4(n9734), 
        .Y(n1483) );
  AO22X1_HVT U1446 ( .A1(\ram[5][143] ), .A2(n5689), .A3(n9285), .A4(n9737), 
        .Y(n1484) );
  AO22X1_HVT U1447 ( .A1(\ram[5][144] ), .A2(n5711), .A3(n9284), .A4(n9741), 
        .Y(n1485) );
  AO22X1_HVT U1448 ( .A1(\ram[5][145] ), .A2(n5692), .A3(n9283), .A4(n9744), 
        .Y(n1486) );
  AO22X1_HVT U1449 ( .A1(\ram[5][146] ), .A2(n4208), .A3(n9282), .A4(n9747), 
        .Y(n1487) );
  AO22X1_HVT U1450 ( .A1(\ram[5][147] ), .A2(n4937), .A3(n9281), .A4(n9750), 
        .Y(n1488) );
  AO22X1_HVT U1451 ( .A1(\ram[5][148] ), .A2(n4813), .A3(n4692), .A4(n9754), 
        .Y(n1489) );
  AO22X1_HVT U1452 ( .A1(\ram[5][149] ), .A2(n4795), .A3(n9273), .A4(n9757), 
        .Y(n1490) );
  AO22X1_HVT U1453 ( .A1(\ram[5][150] ), .A2(n5707), .A3(n9264), .A4(n9760), 
        .Y(n1491) );
  AO22X1_HVT U1454 ( .A1(\ram[5][151] ), .A2(n4230), .A3(n9265), .A4(n9763), 
        .Y(n1492) );
  AO22X1_HVT U1455 ( .A1(\ram[5][152] ), .A2(n4529), .A3(n9256), .A4(n9766), 
        .Y(n1493) );
  AO22X1_HVT U1456 ( .A1(\ram[5][153] ), .A2(n4732), .A3(n9261), .A4(n9769), 
        .Y(n1494) );
  AO22X1_HVT U1457 ( .A1(\ram[5][154] ), .A2(n5702), .A3(n4689), .A4(n9772), 
        .Y(n1495) );
  AO22X1_HVT U1458 ( .A1(\ram[5][155] ), .A2(n5710), .A3(n9259), .A4(n9775), 
        .Y(n1496) );
  AO22X1_HVT U1459 ( .A1(\ram[5][156] ), .A2(n4331), .A3(n9276), .A4(n9779), 
        .Y(n1497) );
  AO22X1_HVT U1460 ( .A1(\ram[5][157] ), .A2(n5712), .A3(n9270), .A4(n9782), 
        .Y(n1498) );
  AO22X1_HVT U1461 ( .A1(\ram[5][158] ), .A2(n5687), .A3(n4690), .A4(n9785), 
        .Y(n1499) );
  AO22X1_HVT U1462 ( .A1(\ram[5][159] ), .A2(n4915), .A3(n9278), .A4(n9788), 
        .Y(n1500) );
  AO22X1_HVT U1463 ( .A1(\ram[5][160] ), .A2(n5678), .A3(n4690), .A4(n9792), 
        .Y(n1501) );
  AO22X1_HVT U1464 ( .A1(\ram[5][161] ), .A2(n5671), .A3(n9277), .A4(n9795), 
        .Y(n1502) );
  AO22X1_HVT U1465 ( .A1(\ram[5][162] ), .A2(n5696), .A3(n9275), .A4(n9798), 
        .Y(n1503) );
  AO22X1_HVT U1466 ( .A1(\ram[5][163] ), .A2(n5692), .A3(n4690), .A4(n9801), 
        .Y(n1504) );
  AO22X1_HVT U1467 ( .A1(\ram[5][164] ), .A2(n5684), .A3(n4692), .A4(n9804), 
        .Y(n1505) );
  AO22X1_HVT U1468 ( .A1(\ram[5][165] ), .A2(n5713), .A3(n9266), .A4(n9807), 
        .Y(n1506) );
  AO22X1_HVT U1469 ( .A1(\ram[5][166] ), .A2(n5687), .A3(n9267), .A4(n9810), 
        .Y(n1507) );
  AO22X1_HVT U1470 ( .A1(\ram[5][167] ), .A2(n4915), .A3(n9264), .A4(n9813), 
        .Y(n1508) );
  AO22X1_HVT U1471 ( .A1(\ram[5][168] ), .A2(n5693), .A3(n9255), .A4(n9816), 
        .Y(n1509) );
  AO22X1_HVT U1472 ( .A1(\ram[5][169] ), .A2(n5709), .A3(n9261), .A4(n9819), 
        .Y(n1510) );
  AO22X1_HVT U1474 ( .A1(\ram[5][171] ), .A2(n5705), .A3(n9259), .A4(n9825), 
        .Y(n1512) );
  AO22X1_HVT U1475 ( .A1(\ram[5][172] ), .A2(n5707), .A3(n9299), .A4(n9829), 
        .Y(n1513) );
  AO22X1_HVT U1476 ( .A1(\ram[5][173] ), .A2(n5685), .A3(n9301), .A4(n9832), 
        .Y(n1514) );
  AO22X1_HVT U1477 ( .A1(\ram[5][174] ), .A2(n5701), .A3(n9299), .A4(n9835), 
        .Y(n1515) );
  AO22X1_HVT U1478 ( .A1(\ram[5][175] ), .A2(n5694), .A3(n9298), .A4(n9838), 
        .Y(n1516) );
  AO22X1_HVT U1479 ( .A1(\ram[5][176] ), .A2(n5677), .A3(n9262), .A4(n9842), 
        .Y(n1517) );
  AO22X1_HVT U1480 ( .A1(\ram[5][177] ), .A2(n5707), .A3(n9282), .A4(n9845), 
        .Y(n1518) );
  AO22X1_HVT U1481 ( .A1(\ram[5][178] ), .A2(n4773), .A3(n9255), .A4(n9848), 
        .Y(n1519) );
  AO22X1_HVT U1482 ( .A1(\ram[5][179] ), .A2(n5696), .A3(n4271), .A4(n9851), 
        .Y(n1520) );
  AO22X1_HVT U1483 ( .A1(\ram[5][180] ), .A2(n5697), .A3(n9272), .A4(n9855), 
        .Y(n1521) );
  AO22X1_HVT U1484 ( .A1(\ram[5][181] ), .A2(n4728), .A3(n9273), .A4(n9858), 
        .Y(n1522) );
  AO22X1_HVT U1485 ( .A1(\ram[5][182] ), .A2(n5676), .A3(n9277), .A4(n9861), 
        .Y(n1523) );
  AO22X1_HVT U1486 ( .A1(\ram[5][183] ), .A2(n5694), .A3(n4691), .A4(n9864), 
        .Y(n1524) );
  AO22X1_HVT U1487 ( .A1(\ram[5][184] ), .A2(n5693), .A3(n4702), .A4(n9868), 
        .Y(n1525) );
  AO22X1_HVT U1488 ( .A1(\ram[5][185] ), .A2(n5676), .A3(n4422), .A4(n9871), 
        .Y(n1526) );
  AO22X1_HVT U1489 ( .A1(\ram[5][186] ), .A2(n5712), .A3(n9304), .A4(n9874), 
        .Y(n1527) );
  AO22X1_HVT U1490 ( .A1(\ram[5][187] ), .A2(n4206), .A3(n9303), .A4(n9877), 
        .Y(n1528) );
  AO22X1_HVT U1491 ( .A1(\ram[5][188] ), .A2(n4206), .A3(n9298), .A4(n9880), 
        .Y(n1529) );
  AO22X1_HVT U1492 ( .A1(\ram[5][189] ), .A2(n5695), .A3(n9299), .A4(n9883), 
        .Y(n1530) );
  AO22X1_HVT U1493 ( .A1(\ram[5][190] ), .A2(n4203), .A3(n9298), .A4(n9886), 
        .Y(n1531) );
  AO22X1_HVT U1494 ( .A1(\ram[5][191] ), .A2(n5683), .A3(n4701), .A4(n9889), 
        .Y(n1532) );
  AO22X1_HVT U1495 ( .A1(\ram[5][192] ), .A2(n5697), .A3(n9299), .A4(n9893), 
        .Y(n1533) );
  AO22X1_HVT U1496 ( .A1(\ram[5][193] ), .A2(n4447), .A3(n9298), .A4(n9896), 
        .Y(n1534) );
  AO22X1_HVT U1497 ( .A1(\ram[5][194] ), .A2(n4897), .A3(n4701), .A4(n9899), 
        .Y(n1535) );
  AO22X1_HVT U1498 ( .A1(\ram[5][195] ), .A2(n5697), .A3(n9300), .A4(n9902), 
        .Y(n1536) );
  AO22X1_HVT U1499 ( .A1(\ram[5][196] ), .A2(n4230), .A3(n9295), .A4(n9906), 
        .Y(n1537) );
  AO22X1_HVT U1500 ( .A1(\ram[5][197] ), .A2(n5709), .A3(n9294), .A4(n9909), 
        .Y(n1538) );
  AO22X1_HVT U1501 ( .A1(\ram[5][198] ), .A2(n4749), .A3(n9293), .A4(n9912), 
        .Y(n1539) );
  AO22X1_HVT U1502 ( .A1(\ram[5][199] ), .A2(n5685), .A3(n9292), .A4(n9915), 
        .Y(n1540) );
  AO22X1_HVT U1503 ( .A1(\ram[5][200] ), .A2(n5678), .A3(n9295), .A4(n9919), 
        .Y(n1541) );
  AO22X1_HVT U1504 ( .A1(\ram[5][201] ), .A2(n4795), .A3(n9294), .A4(n9922), 
        .Y(n1542) );
  AO22X1_HVT U1505 ( .A1(\ram[5][202] ), .A2(n5695), .A3(n9293), .A4(n9925), 
        .Y(n1543) );
  AO22X1_HVT U1506 ( .A1(\ram[5][203] ), .A2(n5702), .A3(n9292), .A4(n9928), 
        .Y(n1544) );
  AO22X1_HVT U1507 ( .A1(\ram[5][204] ), .A2(n4203), .A3(n4702), .A4(n9931), 
        .Y(n1545) );
  AO22X1_HVT U1508 ( .A1(\ram[5][205] ), .A2(n4937), .A3(n9303), .A4(n9934), 
        .Y(n1546) );
  AO22X1_HVT U1509 ( .A1(\ram[5][206] ), .A2(n5705), .A3(n4422), .A4(n9937), 
        .Y(n1547) );
  AO22X1_HVT U1510 ( .A1(\ram[5][207] ), .A2(n5702), .A3(n4422), .A4(n9940), 
        .Y(n1548) );
  AO22X1_HVT U1511 ( .A1(\ram[5][208] ), .A2(n5706), .A3(n9298), .A4(n9944), 
        .Y(n1549) );
  AO22X1_HVT U1512 ( .A1(\ram[5][209] ), .A2(n4321), .A3(n9300), .A4(n9947), 
        .Y(n1550) );
  AO22X1_HVT U1513 ( .A1(\ram[5][210] ), .A2(n5693), .A3(n4701), .A4(n9950), 
        .Y(n1551) );
  AO22X1_HVT U1514 ( .A1(\ram[5][211] ), .A2(n5712), .A3(n9301), .A4(n9953), 
        .Y(n1552) );
  AO22X1_HVT U1516 ( .A1(\ram[5][213] ), .A2(n4915), .A3(n9270), .A4(n9959), 
        .Y(n1554) );
  AO22X1_HVT U1517 ( .A1(\ram[5][214] ), .A2(n4203), .A3(n9278), .A4(n9962), 
        .Y(n1555) );
  AO22X1_HVT U1518 ( .A1(\ram[5][215] ), .A2(n5703), .A3(n9275), .A4(n9965), 
        .Y(n1556) );
  AO22X1_HVT U1519 ( .A1(\ram[5][216] ), .A2(n5692), .A3(n4695), .A4(n9968), 
        .Y(n1557) );
  AO22X1_HVT U1520 ( .A1(\ram[5][217] ), .A2(n4742), .A3(n9272), .A4(n9971), 
        .Y(n1558) );
  AO22X1_HVT U1521 ( .A1(\ram[5][218] ), .A2(n5671), .A3(n4691), .A4(n9974), 
        .Y(n1559) );
  AO22X1_HVT U1522 ( .A1(\ram[5][219] ), .A2(n5709), .A3(n9271), .A4(n9977), 
        .Y(n1560) );
  AO22X1_HVT U1525 ( .A1(\ram[5][222] ), .A2(n5687), .A3(n9301), .A4(n9987), 
        .Y(n1563) );
  AO22X1_HVT U1526 ( .A1(\ram[5][223] ), .A2(n5705), .A3(n9300), .A4(n9990), 
        .Y(n1564) );
  AO22X1_HVT U1527 ( .A1(\ram[5][224] ), .A2(n5690), .A3(n9295), .A4(n9993), 
        .Y(n1565) );
  AO22X1_HVT U1528 ( .A1(\ram[5][225] ), .A2(n5686), .A3(n9294), .A4(n9996), 
        .Y(n1566) );
  AO22X1_HVT U1529 ( .A1(\ram[5][226] ), .A2(n5672), .A3(n9293), .A4(n9999), 
        .Y(n1567) );
  AO22X1_HVT U1530 ( .A1(\ram[5][227] ), .A2(n5697), .A3(n9292), .A4(n10002), 
        .Y(n1568) );
  AO22X1_HVT U1531 ( .A1(\ram[5][228] ), .A2(n4850), .A3(n9291), .A4(n10005), 
        .Y(n1569) );
  AO22X1_HVT U1532 ( .A1(\ram[5][229] ), .A2(n4952), .A3(n9289), .A4(n10008), 
        .Y(n1570) );
  AO22X1_HVT U1534 ( .A1(\ram[5][231] ), .A2(n5662), .A3(n9291), .A4(n10014), 
        .Y(n1572) );
  AO22X1_HVT U1535 ( .A1(\ram[5][232] ), .A2(n4838), .A3(n9275), .A4(n10018), 
        .Y(n1573) );
  AO22X1_HVT U1536 ( .A1(\ram[5][233] ), .A2(n4628), .A3(n9277), .A4(n10021), 
        .Y(n1574) );
  AO22X1_HVT U1538 ( .A1(\ram[5][235] ), .A2(n5684), .A3(n4690), .A4(n10027), 
        .Y(n1576) );
  AO22X1_HVT U1539 ( .A1(\ram[5][236] ), .A2(n5705), .A3(n9289), .A4(n10030), 
        .Y(n1577) );
  AO22X1_HVT U1541 ( .A1(\ram[5][238] ), .A2(n4749), .A3(n5011), .A4(n10036), 
        .Y(n1579) );
  AO22X1_HVT U1542 ( .A1(\ram[5][239] ), .A2(n4765), .A3(n9289), .A4(n10039), 
        .Y(n1580) );
  AO22X1_HVT U1543 ( .A1(\ram[5][240] ), .A2(n4208), .A3(n9278), .A4(n10043), 
        .Y(n1581) );
  AO22X1_HVT U1544 ( .A1(\ram[5][241] ), .A2(n4954), .A3(n9271), .A4(n10046), 
        .Y(n1582) );
  AO22X1_HVT U1545 ( .A1(\ram[5][242] ), .A2(n5662), .A3(n9276), .A4(n10049), 
        .Y(n1583) );
  AO22X1_HVT U1546 ( .A1(\ram[5][243] ), .A2(n5706), .A3(n9278), .A4(n10052), 
        .Y(n1584) );
  AO22X1_HVT U1547 ( .A1(\ram[5][244] ), .A2(n5701), .A3(n4830), .A4(n10055), 
        .Y(n1585) );
  AO22X1_HVT U1548 ( .A1(\ram[5][245] ), .A2(n5702), .A3(n9291), .A4(n10058), 
        .Y(n1586) );
  AO22X1_HVT U1549 ( .A1(\ram[5][246] ), .A2(n5703), .A3(n5011), .A4(n10061), 
        .Y(n1587) );
  AO22X1_HVT U1550 ( .A1(\ram[5][247] ), .A2(n4917), .A3(n9289), .A4(n10064), 
        .Y(n1588) );
  AO22X1_HVT U1551 ( .A1(\ram[5][248] ), .A2(n4206), .A3(n9295), .A4(n10068), 
        .Y(n1589) );
  AO22X1_HVT U1552 ( .A1(\ram[5][249] ), .A2(n5684), .A3(n9294), .A4(n10071), 
        .Y(n1590) );
  AO22X1_HVT U1553 ( .A1(\ram[5][250] ), .A2(n5692), .A3(n9293), .A4(n10074), 
        .Y(n1591) );
  AO22X1_HVT U1554 ( .A1(\ram[5][251] ), .A2(n5707), .A3(n9292), .A4(n10077), 
        .Y(n1592) );
  AO22X1_HVT U1555 ( .A1(\ram[5][252] ), .A2(n5692), .A3(n9284), .A4(n10081), 
        .Y(n1593) );
  AO22X1_HVT U1556 ( .A1(\ram[5][253] ), .A2(n5683), .A3(n9283), .A4(n10084), 
        .Y(n1594) );
  AO22X1_HVT U1557 ( .A1(\ram[5][254] ), .A2(n4773), .A3(n9282), .A4(n10087), 
        .Y(n1595) );
  AO22X1_HVT U1558 ( .A1(\ram[5][255] ), .A2(n5691), .A3(n9281), .A4(n10090), 
        .Y(n1596) );
  AND2X1_HVT U1561 ( .A1(n5880), .A2(n5042), .Y(n28) );
  AO22X1_HVT U1563 ( .A1(\ram[6][1] ), .A2(n5944), .A3(n9231), .A4(n9309), .Y(
        n1598) );
  AO22X1_HVT U1565 ( .A1(\ram[6][3] ), .A2(n5944), .A3(n9229), .A4(n9315), .Y(
        n1600) );
  AO22X1_HVT U1566 ( .A1(\ram[6][4] ), .A2(n5587), .A3(n9228), .A4(n9319), .Y(
        n1601) );
  AO22X1_HVT U1568 ( .A1(\ram[6][6] ), .A2(n5517), .A3(n9226), .A4(n9325), .Y(
        n1603) );
  AO22X1_HVT U1569 ( .A1(\ram[6][7] ), .A2(n5944), .A3(n9225), .A4(n9328), .Y(
        n1604) );
  AO22X1_HVT U1570 ( .A1(\ram[6][8] ), .A2(n5949), .A3(n9210), .A4(n9331), .Y(
        n1605) );
  AO22X1_HVT U1571 ( .A1(\ram[6][9] ), .A2(n10274), .A3(n9209), .A4(n9334), 
        .Y(n1606) );
  AO22X1_HVT U1572 ( .A1(\ram[6][10] ), .A2(n10274), .A3(n9208), .A4(n9337), 
        .Y(n1607) );
  AO22X1_HVT U1573 ( .A1(\ram[6][11] ), .A2(n4704), .A3(n9207), .A4(n9340), 
        .Y(n1608) );
  AO22X1_HVT U1574 ( .A1(\ram[6][12] ), .A2(n10274), .A3(n9204), .A4(n9344), 
        .Y(n1609) );
  AO22X1_HVT U1575 ( .A1(\ram[6][13] ), .A2(n10281), .A3(n9203), .A4(n9347), 
        .Y(n1610) );
  AO22X1_HVT U1576 ( .A1(\ram[6][14] ), .A2(n5949), .A3(n9202), .A4(n9350), 
        .Y(n1611) );
  AO22X1_HVT U1577 ( .A1(\ram[6][15] ), .A2(n5514), .A3(n9201), .A4(n9353), 
        .Y(n1612) );
  AO22X1_HVT U1579 ( .A1(\ram[6][17] ), .A2(n4700), .A3(n9231), .A4(n9359), 
        .Y(n1614) );
  AO22X1_HVT U1580 ( .A1(\ram[6][18] ), .A2(n5944), .A3(n9230), .A4(n9362), 
        .Y(n1615) );
  AO22X1_HVT U1581 ( .A1(\ram[6][19] ), .A2(n5944), .A3(n9229), .A4(n9365), 
        .Y(n1616) );
  AO22X1_HVT U1583 ( .A1(\ram[6][21] ), .A2(n5545), .A3(n9231), .A4(n9370), 
        .Y(n1618) );
  AO22X1_HVT U1584 ( .A1(\ram[6][22] ), .A2(n10274), .A3(n9230), .A4(n9373), 
        .Y(n1619) );
  AO22X1_HVT U1585 ( .A1(\ram[6][23] ), .A2(n5949), .A3(n9229), .A4(n9376), 
        .Y(n1620) );
  AO22X1_HVT U1586 ( .A1(\ram[6][24] ), .A2(n5513), .A3(n9241), .A4(n9379), 
        .Y(n1621) );
  AO22X1_HVT U1587 ( .A1(\ram[6][25] ), .A2(n4920), .A3(n9240), .A4(n9382), 
        .Y(n1622) );
  AO22X1_HVT U1588 ( .A1(\ram[6][26] ), .A2(n5949), .A3(n9239), .A4(n9385), 
        .Y(n1623) );
  AO22X1_HVT U1589 ( .A1(\ram[6][27] ), .A2(n5944), .A3(n9238), .A4(n9388), 
        .Y(n1624) );
  AO22X1_HVT U1590 ( .A1(\ram[6][28] ), .A2(n6628), .A3(n9241), .A4(n9391), 
        .Y(n1625) );
  AO22X1_HVT U1591 ( .A1(\ram[6][29] ), .A2(n10274), .A3(n9240), .A4(n9394), 
        .Y(n1626) );
  AO22X1_HVT U1595 ( .A1(\ram[6][33] ), .A2(n5184), .A3(n9236), .A4(n9406), 
        .Y(n1630) );
  AO22X1_HVT U1596 ( .A1(\ram[6][34] ), .A2(n5190), .A3(n9235), .A4(n9409), 
        .Y(n1631) );
  AO22X1_HVT U1597 ( .A1(\ram[6][35] ), .A2(n5194), .A3(n9234), .A4(n9412), 
        .Y(n1632) );
  AO22X1_HVT U1599 ( .A1(\ram[6][37] ), .A2(n5192), .A3(n9221), .A4(n9418), 
        .Y(n1634) );
  AO22X1_HVT U1600 ( .A1(\ram[6][38] ), .A2(n5191), .A3(n9220), .A4(n9421), 
        .Y(n1635) );
  AO22X1_HVT U1603 ( .A1(\ram[6][41] ), .A2(n5185), .A3(n9209), .A4(n9430), 
        .Y(n1638) );
  AO22X1_HVT U1604 ( .A1(\ram[6][42] ), .A2(n5176), .A3(n9208), .A4(n9433), 
        .Y(n1639) );
  AO22X1_HVT U1605 ( .A1(\ram[6][43] ), .A2(n5191), .A3(n9207), .A4(n9436), 
        .Y(n1640) );
  AO22X1_HVT U1606 ( .A1(\ram[6][44] ), .A2(n5186), .A3(n9200), .A4(n9439), 
        .Y(n1641) );
  AO22X1_HVT U1607 ( .A1(\ram[6][45] ), .A2(n5181), .A3(n9199), .A4(n9442), 
        .Y(n1642) );
  AO22X1_HVT U1608 ( .A1(\ram[6][46] ), .A2(n5179), .A3(n9198), .A4(n9445), 
        .Y(n1643) );
  AO22X1_HVT U1614 ( .A1(\ram[6][52] ), .A2(n4858), .A3(n9216), .A4(n9463), 
        .Y(n1649) );
  AO22X1_HVT U1617 ( .A1(\ram[6][55] ), .A2(n10280), .A3(n9213), .A4(n9472), 
        .Y(n1652) );
  AO22X1_HVT U1618 ( .A1(\ram[6][56] ), .A2(n5514), .A3(n9251), .A4(n9475), 
        .Y(n1653) );
  AO22X1_HVT U1619 ( .A1(\ram[6][57] ), .A2(n4704), .A3(n9250), .A4(n9478), 
        .Y(n1654) );
  AO22X1_HVT U1620 ( .A1(\ram[6][58] ), .A2(n10277), .A3(n9249), .A4(n9481), 
        .Y(n1655) );
  AO22X1_HVT U1621 ( .A1(\ram[6][59] ), .A2(n4700), .A3(n9248), .A4(n9484), 
        .Y(n1656) );
  AO22X1_HVT U1622 ( .A1(\ram[6][60] ), .A2(n5514), .A3(n9216), .A4(n9487), 
        .Y(n1657) );
  AO22X1_HVT U1623 ( .A1(\ram[6][61] ), .A2(n10279), .A3(n9215), .A4(n9490), 
        .Y(n1658) );
  AO22X1_HVT U1624 ( .A1(\ram[6][62] ), .A2(n10279), .A3(n9214), .A4(n9493), 
        .Y(n1659) );
  AO22X1_HVT U1625 ( .A1(\ram[6][63] ), .A2(n5545), .A3(n9213), .A4(n9496), 
        .Y(n1660) );
  AO22X1_HVT U1626 ( .A1(\ram[6][64] ), .A2(n10277), .A3(n9204), .A4(n9499), 
        .Y(n1661) );
  AO22X1_HVT U1627 ( .A1(\ram[6][65] ), .A2(n5517), .A3(n9203), .A4(n9502), 
        .Y(n1662) );
  AO22X1_HVT U1628 ( .A1(\ram[6][66] ), .A2(n10279), .A3(n9202), .A4(n9505), 
        .Y(n1663) );
  AO22X1_HVT U1629 ( .A1(\ram[6][67] ), .A2(n6630), .A3(n9201), .A4(n9508), 
        .Y(n1664) );
  AO22X1_HVT U1631 ( .A1(\ram[6][69] ), .A2(n10277), .A3(n9227), .A4(n9514), 
        .Y(n1666) );
  AO22X1_HVT U1632 ( .A1(\ram[6][70] ), .A2(n5513), .A3(n9226), .A4(n9517), 
        .Y(n1667) );
  AO22X1_HVT U1633 ( .A1(\ram[6][71] ), .A2(n4704), .A3(n9225), .A4(n9520), 
        .Y(n1668) );
  AO22X1_HVT U1634 ( .A1(\ram[6][72] ), .A2(n10276), .A3(n9200), .A4(n9523), 
        .Y(n1669) );
  AO22X1_HVT U1635 ( .A1(\ram[6][73] ), .A2(n10280), .A3(n9199), .A4(n9526), 
        .Y(n1670) );
  AO22X1_HVT U1636 ( .A1(\ram[6][74] ), .A2(n5513), .A3(n9198), .A4(n9529), 
        .Y(n1671) );
  AO22X1_HVT U1637 ( .A1(\ram[6][75] ), .A2(n10276), .A3(n9197), .A4(n9532), 
        .Y(n1672) );
  AO22X1_HVT U1638 ( .A1(\ram[6][76] ), .A2(n4720), .A3(n9228), .A4(n9535), 
        .Y(n1673) );
  AO22X1_HVT U1639 ( .A1(\ram[6][77] ), .A2(n4859), .A3(n9227), .A4(n9538), 
        .Y(n1674) );
  AO22X1_HVT U1640 ( .A1(\ram[6][78] ), .A2(n10275), .A3(n9226), .A4(n9541), 
        .Y(n1675) );
  AO22X1_HVT U1641 ( .A1(\ram[6][79] ), .A2(n10275), .A3(n9225), .A4(n9544), 
        .Y(n1676) );
  AO22X1_HVT U1642 ( .A1(\ram[6][80] ), .A2(n10279), .A3(n9237), .A4(n9547), 
        .Y(n1677) );
  AO22X1_HVT U1643 ( .A1(\ram[6][81] ), .A2(n4859), .A3(n9236), .A4(n9550), 
        .Y(n1678) );
  AO22X1_HVT U1644 ( .A1(\ram[6][82] ), .A2(n4858), .A3(n9235), .A4(n9553), 
        .Y(n1679) );
  AO22X1_HVT U1645 ( .A1(\ram[6][83] ), .A2(n4704), .A3(n9234), .A4(n9556), 
        .Y(n1680) );
  AO22X1_HVT U1646 ( .A1(\ram[6][84] ), .A2(n10282), .A3(n9204), .A4(n9559), 
        .Y(n1681) );
  AO22X1_HVT U1647 ( .A1(\ram[6][85] ), .A2(n5516), .A3(n9203), .A4(n9562), 
        .Y(n1682) );
  AO22X1_HVT U1648 ( .A1(\ram[6][86] ), .A2(n10279), .A3(n9202), .A4(n9565), 
        .Y(n1683) );
  AO22X1_HVT U1649 ( .A1(\ram[6][87] ), .A2(n4859), .A3(n9201), .A4(n9568), 
        .Y(n1684) );
  AO22X1_HVT U1650 ( .A1(\ram[6][88] ), .A2(n10280), .A3(n9240), .A4(n9571), 
        .Y(n1685) );
  AO22X1_HVT U1651 ( .A1(\ram[6][89] ), .A2(n6630), .A3(n9231), .A4(n9574), 
        .Y(n1686) );
  AO22X1_HVT U1652 ( .A1(\ram[6][90] ), .A2(n6628), .A3(n9230), .A4(n9577), 
        .Y(n1687) );
  AO22X1_HVT U1653 ( .A1(\ram[6][91] ), .A2(n10277), .A3(n9229), .A4(n9580), 
        .Y(n1688) );
  AO22X1_HVT U1654 ( .A1(\ram[6][92] ), .A2(n10275), .A3(n9228), .A4(n9583), 
        .Y(n1689) );
  AO22X1_HVT U1655 ( .A1(\ram[6][93] ), .A2(n5516), .A3(n9227), .A4(n9586), 
        .Y(n1690) );
  AO22X1_HVT U1656 ( .A1(\ram[6][94] ), .A2(n4859), .A3(n9226), .A4(n9589), 
        .Y(n1691) );
  AO22X1_HVT U1657 ( .A1(\ram[6][95] ), .A2(n10278), .A3(n9225), .A4(n9592), 
        .Y(n1692) );
  AO22X1_HVT U1658 ( .A1(\ram[6][96] ), .A2(n10280), .A3(n9200), .A4(n9595), 
        .Y(n1693) );
  AO22X1_HVT U1659 ( .A1(\ram[6][97] ), .A2(n5517), .A3(n9199), .A4(n9598), 
        .Y(n1694) );
  AO22X1_HVT U1660 ( .A1(\ram[6][98] ), .A2(n10276), .A3(n9198), .A4(n9601), 
        .Y(n1695) );
  AO22X1_HVT U1661 ( .A1(\ram[6][99] ), .A2(n6628), .A3(n9197), .A4(n9604), 
        .Y(n1696) );
  AO22X1_HVT U1662 ( .A1(\ram[6][100] ), .A2(n5587), .A3(n9251), .A4(n9607), 
        .Y(n1697) );
  AO22X1_HVT U1663 ( .A1(\ram[6][101] ), .A2(n4858), .A3(n9250), .A4(n9610), 
        .Y(n1698) );
  AO22X1_HVT U1664 ( .A1(\ram[6][102] ), .A2(n10278), .A3(n9249), .A4(n9613), 
        .Y(n1699) );
  AO22X1_HVT U1665 ( .A1(\ram[6][103] ), .A2(n10275), .A3(n9248), .A4(n9616), 
        .Y(n1700) );
  AO22X1_HVT U1666 ( .A1(\ram[6][104] ), .A2(n5516), .A3(n9246), .A4(n9619), 
        .Y(n1701) );
  AO22X1_HVT U1667 ( .A1(\ram[6][105] ), .A2(n10277), .A3(n9245), .A4(n9622), 
        .Y(n1702) );
  AO22X1_HVT U1668 ( .A1(\ram[6][106] ), .A2(n5516), .A3(n9245), .A4(n9625), 
        .Y(n1703) );
  AO22X1_HVT U1669 ( .A1(\ram[6][107] ), .A2(n10276), .A3(n4350), .A4(n9628), 
        .Y(n1704) );
  AO22X1_HVT U1670 ( .A1(\ram[6][108] ), .A2(n5517), .A3(n9231), .A4(n9631), 
        .Y(n1705) );
  AO22X1_HVT U1671 ( .A1(\ram[6][109] ), .A2(n4858), .A3(n9231), .A4(n9634), 
        .Y(n1706) );
  AO22X1_HVT U1672 ( .A1(\ram[6][110] ), .A2(n10276), .A3(n9230), .A4(n9637), 
        .Y(n1707) );
  AO22X1_HVT U1673 ( .A1(\ram[6][111] ), .A2(n5587), .A3(n9229), .A4(n9640), 
        .Y(n1708) );
  AO22X1_HVT U1674 ( .A1(\ram[6][112] ), .A2(n10275), .A3(n9216), .A4(n9643), 
        .Y(n1709) );
  AO22X1_HVT U1675 ( .A1(\ram[6][113] ), .A2(n10278), .A3(n9215), .A4(n9646), 
        .Y(n1710) );
  AO22X1_HVT U1676 ( .A1(\ram[6][114] ), .A2(n6630), .A3(n9214), .A4(n9649), 
        .Y(n1711) );
  AO22X1_HVT U1677 ( .A1(\ram[6][115] ), .A2(n6629), .A3(n9213), .A4(n9652), 
        .Y(n1712) );
  AO22X1_HVT U1678 ( .A1(\ram[6][116] ), .A2(n10281), .A3(n9251), .A4(n9655), 
        .Y(n1713) );
  AO22X1_HVT U1679 ( .A1(\ram[6][117] ), .A2(n6630), .A3(n9250), .A4(n9658), 
        .Y(n1714) );
  AO22X1_HVT U1681 ( .A1(\ram[6][119] ), .A2(n4859), .A3(n9248), .A4(n9664), 
        .Y(n1716) );
  AO22X1_HVT U1682 ( .A1(\ram[6][120] ), .A2(n10284), .A3(n9237), .A4(n9667), 
        .Y(n1717) );
  AO22X1_HVT U1683 ( .A1(\ram[6][121] ), .A2(n10283), .A3(n9236), .A4(n9670), 
        .Y(n1718) );
  AO22X1_HVT U1684 ( .A1(\ram[6][122] ), .A2(n4415), .A3(n9235), .A4(n9673), 
        .Y(n1719) );
  AO22X1_HVT U1685 ( .A1(\ram[6][123] ), .A2(n6629), .A3(n9234), .A4(n9676), 
        .Y(n1720) );
  AO22X1_HVT U1686 ( .A1(\ram[6][124] ), .A2(n6628), .A3(n9210), .A4(n9679), 
        .Y(n1721) );
  AO22X1_HVT U1687 ( .A1(\ram[6][125] ), .A2(n6627), .A3(n9209), .A4(n9682), 
        .Y(n1722) );
  AO22X1_HVT U1688 ( .A1(\ram[6][126] ), .A2(n5517), .A3(n9208), .A4(n9685), 
        .Y(n1723) );
  AO22X1_HVT U1689 ( .A1(\ram[6][127] ), .A2(n4704), .A3(n9207), .A4(n9688), 
        .Y(n1724) );
  AO22X1_HVT U1690 ( .A1(\ram[6][128] ), .A2(n5545), .A3(n9251), .A4(n9691), 
        .Y(n1725) );
  AO22X1_HVT U1691 ( .A1(\ram[6][129] ), .A2(n10284), .A3(n9250), .A4(n9694), 
        .Y(n1726) );
  AO22X1_HVT U1692 ( .A1(\ram[6][130] ), .A2(n6627), .A3(n9249), .A4(n9697), 
        .Y(n1727) );
  AO22X1_HVT U1693 ( .A1(\ram[6][131] ), .A2(n10285), .A3(n9248), .A4(n9700), 
        .Y(n1728) );
  AO22X1_HVT U1694 ( .A1(\ram[6][132] ), .A2(n5514), .A3(n9210), .A4(n9703), 
        .Y(n1729) );
  AO22X1_HVT U1695 ( .A1(\ram[6][133] ), .A2(n10282), .A3(n9209), .A4(n9706), 
        .Y(n1730) );
  AO22X1_HVT U1696 ( .A1(\ram[6][134] ), .A2(n5516), .A3(n9208), .A4(n9709), 
        .Y(n1731) );
  AO22X1_HVT U1697 ( .A1(\ram[6][135] ), .A2(n4704), .A3(n9207), .A4(n9712), 
        .Y(n1732) );
  AO22X1_HVT U1698 ( .A1(\ram[6][136] ), .A2(n10284), .A3(n9204), .A4(n9715), 
        .Y(n1733) );
  AO22X1_HVT U1699 ( .A1(\ram[6][137] ), .A2(n5546), .A3(n9203), .A4(n9718), 
        .Y(n1734) );
  AO22X1_HVT U1700 ( .A1(\ram[6][138] ), .A2(n10283), .A3(n9202), .A4(n9721), 
        .Y(n1735) );
  AO22X1_HVT U1701 ( .A1(\ram[6][139] ), .A2(n10285), .A3(n9201), .A4(n9724), 
        .Y(n1736) );
  AO22X1_HVT U1702 ( .A1(\ram[6][140] ), .A2(n5513), .A3(n9216), .A4(n9728), 
        .Y(n1737) );
  AO22X1_HVT U1703 ( .A1(\ram[6][141] ), .A2(n5546), .A3(n9231), .A4(n9731), 
        .Y(n1738) );
  AO22X1_HVT U1704 ( .A1(\ram[6][142] ), .A2(n10280), .A3(n9230), .A4(n9734), 
        .Y(n1739) );
  AO22X1_HVT U1705 ( .A1(\ram[6][143] ), .A2(n10278), .A3(n9229), .A4(n9737), 
        .Y(n1740) );
  AO22X1_HVT U1706 ( .A1(\ram[6][144] ), .A2(n10284), .A3(n9228), .A4(n9741), 
        .Y(n1741) );
  AO22X1_HVT U1707 ( .A1(\ram[6][145] ), .A2(n10282), .A3(n9227), .A4(n9744), 
        .Y(n1742) );
  AO22X1_HVT U1708 ( .A1(\ram[6][146] ), .A2(n6627), .A3(n9226), .A4(n9747), 
        .Y(n1743) );
  AO22X1_HVT U1709 ( .A1(\ram[6][147] ), .A2(n10283), .A3(n9225), .A4(n9750), 
        .Y(n1744) );
  AO22X1_HVT U1710 ( .A1(\ram[6][148] ), .A2(n4720), .A3(n9210), .A4(n9754), 
        .Y(n1745) );
  AO22X1_HVT U1711 ( .A1(\ram[6][149] ), .A2(n6627), .A3(n9209), .A4(n9757), 
        .Y(n1746) );
  AO22X1_HVT U1712 ( .A1(\ram[6][150] ), .A2(n6629), .A3(n9208), .A4(n9760), 
        .Y(n1747) );
  AO22X1_HVT U1713 ( .A1(\ram[6][151] ), .A2(n5587), .A3(n9207), .A4(n9763), 
        .Y(n1748) );
  AO22X1_HVT U1714 ( .A1(\ram[6][152] ), .A2(n5513), .A3(n9204), .A4(n9766), 
        .Y(n1749) );
  AO22X1_HVT U1715 ( .A1(\ram[6][153] ), .A2(n10285), .A3(n9203), .A4(n9769), 
        .Y(n1750) );
  AO22X1_HVT U1716 ( .A1(\ram[6][154] ), .A2(n5546), .A3(n9202), .A4(n9772), 
        .Y(n1751) );
  AO22X1_HVT U1717 ( .A1(\ram[6][155] ), .A2(n6627), .A3(n9201), .A4(n9775), 
        .Y(n1752) );
  AO22X1_HVT U1718 ( .A1(\ram[6][156] ), .A2(n6628), .A3(n9222), .A4(n9779), 
        .Y(n1753) );
  AO22X1_HVT U1719 ( .A1(\ram[6][157] ), .A2(n4700), .A3(n9221), .A4(n9782), 
        .Y(n1754) );
  AO22X1_HVT U1720 ( .A1(\ram[6][158] ), .A2(n10279), .A3(n9220), .A4(n9785), 
        .Y(n1755) );
  AO22X1_HVT U1721 ( .A1(\ram[6][159] ), .A2(n10278), .A3(n9219), .A4(n9788), 
        .Y(n1756) );
  AO22X1_HVT U1722 ( .A1(\ram[6][160] ), .A2(n10284), .A3(n9222), .A4(n9792), 
        .Y(n1757) );
  AO22X1_HVT U1723 ( .A1(\ram[6][161] ), .A2(n10282), .A3(n9221), .A4(n9795), 
        .Y(n1758) );
  AO22X1_HVT U1724 ( .A1(\ram[6][162] ), .A2(n6629), .A3(n9220), .A4(n9798), 
        .Y(n1759) );
  AO22X1_HVT U1725 ( .A1(\ram[6][163] ), .A2(n5546), .A3(n9219), .A4(n9801), 
        .Y(n1760) );
  AO22X1_HVT U1726 ( .A1(\ram[6][164] ), .A2(n4415), .A3(n9210), .A4(n9804), 
        .Y(n1761) );
  AO22X1_HVT U1727 ( .A1(\ram[6][165] ), .A2(n6629), .A3(n9209), .A4(n9807), 
        .Y(n1762) );
  AO22X1_HVT U1728 ( .A1(\ram[6][166] ), .A2(n5517), .A3(n9208), .A4(n9810), 
        .Y(n1763) );
  AO22X1_HVT U1729 ( .A1(\ram[6][167] ), .A2(n10281), .A3(n9207), .A4(n9813), 
        .Y(n1764) );
  AO22X1_HVT U1730 ( .A1(\ram[6][168] ), .A2(n10284), .A3(n9204), .A4(n9816), 
        .Y(n1765) );
  AO22X1_HVT U1731 ( .A1(\ram[6][169] ), .A2(n10283), .A3(n9203), .A4(n9819), 
        .Y(n1766) );
  AO22X1_HVT U1732 ( .A1(\ram[6][170] ), .A2(n10283), .A3(n9202), .A4(n9822), 
        .Y(n1767) );
  AO22X1_HVT U1733 ( .A1(\ram[6][171] ), .A2(n4858), .A3(n9201), .A4(n9825), 
        .Y(n1768) );
  AO22X1_HVT U1734 ( .A1(\ram[6][172] ), .A2(n6628), .A3(n9244), .A4(n9829), 
        .Y(n1769) );
  AO22X1_HVT U1735 ( .A1(\ram[6][173] ), .A2(n10285), .A3(n9244), .A4(n9832), 
        .Y(n1770) );
  AO22X1_HVT U1736 ( .A1(\ram[6][174] ), .A2(n4415), .A3(n9247), .A4(n9835), 
        .Y(n1771) );
  AO22X1_HVT U1737 ( .A1(\ram[6][175] ), .A2(n10281), .A3(n9247), .A4(n9838), 
        .Y(n1772) );
  AO22X1_HVT U1738 ( .A1(\ram[6][176] ), .A2(n5514), .A3(n9200), .A4(n9842), 
        .Y(n1773) );
  AO22X1_HVT U1739 ( .A1(\ram[6][177] ), .A2(n6627), .A3(n9199), .A4(n9845), 
        .Y(n1774) );
  AO22X1_HVT U1740 ( .A1(\ram[6][178] ), .A2(n5545), .A3(n9198), .A4(n9848), 
        .Y(n1775) );
  AO22X1_HVT U1741 ( .A1(\ram[6][179] ), .A2(n10285), .A3(n9197), .A4(n9851), 
        .Y(n1776) );
  AO22X1_HVT U1742 ( .A1(\ram[6][180] ), .A2(n5514), .A3(n9216), .A4(n9855), 
        .Y(n1777) );
  AO22X1_HVT U1743 ( .A1(\ram[6][181] ), .A2(n5546), .A3(n9215), .A4(n9858), 
        .Y(n1778) );
  AO22X1_HVT U1744 ( .A1(\ram[6][182] ), .A2(n10280), .A3(n9214), .A4(n9861), 
        .Y(n1779) );
  AO22X1_HVT U1745 ( .A1(\ram[6][183] ), .A2(n10281), .A3(n9213), .A4(n9864), 
        .Y(n1780) );
  AO22X1_HVT U1746 ( .A1(\ram[6][184] ), .A2(n4720), .A3(n9251), .A4(n9868), 
        .Y(n1781) );
  AO22X1_HVT U1747 ( .A1(\ram[6][185] ), .A2(n5546), .A3(n9250), .A4(n9871), 
        .Y(n1782) );
  AO22X1_HVT U1748 ( .A1(\ram[6][186] ), .A2(n10285), .A3(n9249), .A4(n9874), 
        .Y(n1783) );
  AO22X1_HVT U1749 ( .A1(\ram[6][187] ), .A2(n4415), .A3(n9248), .A4(n9877), 
        .Y(n1784) );
  AO22X1_HVT U1750 ( .A1(\ram[6][188] ), .A2(n5513), .A3(n9246), .A4(n9880), 
        .Y(n1785) );
  AO22X1_HVT U1751 ( .A1(\ram[6][189] ), .A2(n10283), .A3(n9246), .A4(n9883), 
        .Y(n1786) );
  AO22X1_HVT U1752 ( .A1(\ram[6][190] ), .A2(n10276), .A3(n9247), .A4(n9886), 
        .Y(n1787) );
  AO22X1_HVT U1753 ( .A1(\ram[6][191] ), .A2(n5587), .A3(n9247), .A4(n9889), 
        .Y(n1788) );
  AO22X1_HVT U1755 ( .A1(\ram[6][193] ), .A2(n5180), .A3(n9246), .A4(n9896), 
        .Y(n1790) );
  AO22X1_HVT U1756 ( .A1(\ram[6][194] ), .A2(n5193), .A3(n9245), .A4(n9899), 
        .Y(n1791) );
  AO22X1_HVT U1758 ( .A1(\ram[6][196] ), .A2(n5185), .A3(n9241), .A4(n9906), 
        .Y(n1793) );
  AO22X1_HVT U1759 ( .A1(\ram[6][197] ), .A2(n5187), .A3(n9240), .A4(n9909), 
        .Y(n1794) );
  AO22X1_HVT U1760 ( .A1(\ram[6][198] ), .A2(n5187), .A3(n9239), .A4(n9912), 
        .Y(n1795) );
  AO22X1_HVT U1761 ( .A1(\ram[6][199] ), .A2(n5182), .A3(n9238), .A4(n9915), 
        .Y(n1796) );
  AO22X1_HVT U1762 ( .A1(\ram[6][200] ), .A2(n5180), .A3(n9241), .A4(n9919), 
        .Y(n1797) );
  AO22X1_HVT U1764 ( .A1(\ram[6][202] ), .A2(n5181), .A3(n9239), .A4(n9925), 
        .Y(n1799) );
  AO22X1_HVT U1765 ( .A1(\ram[6][203] ), .A2(n5175), .A3(n9238), .A4(n9928), 
        .Y(n1800) );
  AO22X1_HVT U1767 ( .A1(\ram[6][205] ), .A2(n5194), .A3(n9250), .A4(n9934), 
        .Y(n1802) );
  AO22X1_HVT U1768 ( .A1(\ram[6][206] ), .A2(n5182), .A3(n9249), .A4(n9937), 
        .Y(n1803) );
  AO22X1_HVT U1769 ( .A1(\ram[6][207] ), .A2(n5179), .A3(n9248), .A4(n9940), 
        .Y(n1804) );
  AO22X1_HVT U1770 ( .A1(\ram[6][208] ), .A2(n5193), .A3(n9244), .A4(n9944), 
        .Y(n1805) );
  AO22X1_HVT U1771 ( .A1(\ram[6][209] ), .A2(n5176), .A3(n9245), .A4(n9947), 
        .Y(n1806) );
  AO22X1_HVT U1772 ( .A1(\ram[6][210] ), .A2(n5194), .A3(n9244), .A4(n9950), 
        .Y(n1807) );
  AO22X1_HVT U1773 ( .A1(\ram[6][211] ), .A2(n5174), .A3(n4227), .A4(n9953), 
        .Y(n1808) );
  AO22X1_HVT U1774 ( .A1(\ram[6][212] ), .A2(n5176), .A3(n9222), .A4(n9956), 
        .Y(n1809) );
  AO22X1_HVT U1775 ( .A1(\ram[6][213] ), .A2(n5191), .A3(n9221), .A4(n9959), 
        .Y(n1810) );
  AO22X1_HVT U1776 ( .A1(\ram[6][214] ), .A2(n5190), .A3(n9220), .A4(n9962), 
        .Y(n1811) );
  AO22X1_HVT U1777 ( .A1(\ram[6][215] ), .A2(n5194), .A3(n9219), .A4(n9965), 
        .Y(n1812) );
  AO22X1_HVT U1778 ( .A1(\ram[6][216] ), .A2(n5179), .A3(n9216), .A4(n9968), 
        .Y(n1813) );
  AO22X1_HVT U1780 ( .A1(\ram[6][218] ), .A2(n5180), .A3(n9214), .A4(n9974), 
        .Y(n1815) );
  AO22X1_HVT U1781 ( .A1(\ram[6][219] ), .A2(n5174), .A3(n9213), .A4(n9977), 
        .Y(n1816) );
  AO22X1_HVT U1782 ( .A1(\ram[6][220] ), .A2(n5188), .A3(n4350), .A4(n9981), 
        .Y(n1817) );
  AO22X1_HVT U1783 ( .A1(\ram[6][221] ), .A2(n5188), .A3(n4350), .A4(n9984), 
        .Y(n1818) );
  AO22X1_HVT U1784 ( .A1(\ram[6][222] ), .A2(n5179), .A3(n4350), .A4(n9987), 
        .Y(n1819) );
  AO22X1_HVT U1785 ( .A1(\ram[6][223] ), .A2(n5193), .A3(n4227), .A4(n9990), 
        .Y(n1820) );
  AO22X1_HVT U1786 ( .A1(\ram[6][224] ), .A2(n5190), .A3(n9241), .A4(n9993), 
        .Y(n1821) );
  AO22X1_HVT U1787 ( .A1(\ram[6][225] ), .A2(n5176), .A3(n9240), .A4(n9996), 
        .Y(n1822) );
  AO22X1_HVT U1788 ( .A1(\ram[6][226] ), .A2(n5180), .A3(n9239), .A4(n9999), 
        .Y(n1823) );
  AO22X1_HVT U1789 ( .A1(\ram[6][227] ), .A2(n5188), .A3(n9238), .A4(n10002), 
        .Y(n1824) );
  AO22X1_HVT U1790 ( .A1(\ram[6][228] ), .A2(n5181), .A3(n9237), .A4(n10005), 
        .Y(n1825) );
  AO22X1_HVT U1791 ( .A1(\ram[6][229] ), .A2(n5192), .A3(n9236), .A4(n10008), 
        .Y(n1826) );
  AO22X1_HVT U1792 ( .A1(\ram[6][230] ), .A2(n5185), .A3(n9235), .A4(n10011), 
        .Y(n1827) );
  AO22X1_HVT U1793 ( .A1(\ram[6][231] ), .A2(n5192), .A3(n9234), .A4(n10014), 
        .Y(n1828) );
  AO22X1_HVT U1794 ( .A1(\ram[6][232] ), .A2(n5174), .A3(n9222), .A4(n10018), 
        .Y(n1829) );
  AO22X1_HVT U1795 ( .A1(\ram[6][233] ), .A2(n5187), .A3(n9221), .A4(n10021), 
        .Y(n1830) );
  AO22X1_HVT U1796 ( .A1(\ram[6][234] ), .A2(n5182), .A3(n9220), .A4(n10024), 
        .Y(n1831) );
  AO22X1_HVT U1798 ( .A1(\ram[6][236] ), .A2(n5175), .A3(n9237), .A4(n10030), 
        .Y(n1833) );
  AO22X1_HVT U1799 ( .A1(\ram[6][237] ), .A2(n5181), .A3(n9236), .A4(n10033), 
        .Y(n1834) );
  AO22X1_HVT U1800 ( .A1(\ram[6][238] ), .A2(n5190), .A3(n9235), .A4(n10036), 
        .Y(n1835) );
  AO22X1_HVT U1801 ( .A1(\ram[6][239] ), .A2(n5187), .A3(n9234), .A4(n10039), 
        .Y(n1836) );
  AO22X1_HVT U1802 ( .A1(\ram[6][240] ), .A2(n5186), .A3(n9222), .A4(n10043), 
        .Y(n1837) );
  AO22X1_HVT U1803 ( .A1(\ram[6][241] ), .A2(n5191), .A3(n9221), .A4(n10046), 
        .Y(n1838) );
  AO22X1_HVT U1804 ( .A1(\ram[6][242] ), .A2(n5179), .A3(n9220), .A4(n10049), 
        .Y(n1839) );
  AO22X1_HVT U1805 ( .A1(\ram[6][243] ), .A2(n5184), .A3(n9219), .A4(n10052), 
        .Y(n1840) );
  AO22X1_HVT U1806 ( .A1(\ram[6][244] ), .A2(n5182), .A3(n9237), .A4(n10055), 
        .Y(n1841) );
  AO22X1_HVT U1807 ( .A1(\ram[6][245] ), .A2(n5186), .A3(n9236), .A4(n10058), 
        .Y(n1842) );
  AO22X1_HVT U1808 ( .A1(\ram[6][246] ), .A2(n5184), .A3(n9235), .A4(n10061), 
        .Y(n1843) );
  AO22X1_HVT U1809 ( .A1(\ram[6][247] ), .A2(n5175), .A3(n9234), .A4(n10064), 
        .Y(n1844) );
  AO22X1_HVT U1810 ( .A1(\ram[6][248] ), .A2(n5192), .A3(n9241), .A4(n10068), 
        .Y(n1845) );
  AO22X1_HVT U1811 ( .A1(\ram[6][249] ), .A2(n5193), .A3(n9240), .A4(n10071), 
        .Y(n1846) );
  AO22X1_HVT U1812 ( .A1(\ram[6][250] ), .A2(n5184), .A3(n9239), .A4(n10074), 
        .Y(n1847) );
  AO22X1_HVT U1813 ( .A1(\ram[6][251] ), .A2(n5180), .A3(n9238), .A4(n10077), 
        .Y(n1848) );
  AO22X1_HVT U1814 ( .A1(\ram[6][252] ), .A2(n5181), .A3(n9228), .A4(n10081), 
        .Y(n1849) );
  AO22X1_HVT U1815 ( .A1(\ram[6][253] ), .A2(n5188), .A3(n9227), .A4(n10084), 
        .Y(n1850) );
  AO22X1_HVT U1816 ( .A1(\ram[6][254] ), .A2(n5186), .A3(n9226), .A4(n10087), 
        .Y(n1851) );
  AO22X1_HVT U1817 ( .A1(\ram[6][255] ), .A2(n5187), .A3(n9225), .A4(n10090), 
        .Y(n1852) );
  AND2X1_HVT U1818 ( .A1(n5626), .A2(n10375), .Y(n30) );
  AO22X1_HVT U1821 ( .A1(\ram[7][0] ), .A2(n6918), .A3(n9174), .A4(n9306), .Y(
        n1853) );
  AO22X1_HVT U1822 ( .A1(\ram[7][1] ), .A2(n6964), .A3(n9173), .A4(data[1]), 
        .Y(n1854) );
  AO22X1_HVT U1823 ( .A1(\ram[7][2] ), .A2(n6953), .A3(n9172), .A4(n9313), .Y(
        n1855) );
  AO22X1_HVT U1824 ( .A1(\ram[7][3] ), .A2(n6952), .A3(n9171), .A4(n9317), .Y(
        n1856) );
  AO22X1_HVT U1825 ( .A1(\ram[7][4] ), .A2(n6952), .A3(n9170), .A4(data[4]), 
        .Y(n1857) );
  AO22X1_HVT U1826 ( .A1(\ram[7][5] ), .A2(n6951), .A3(n9169), .A4(n9322), .Y(
        n1858) );
  AO22X1_HVT U1827 ( .A1(\ram[7][6] ), .A2(n6950), .A3(n9168), .A4(data[6]), 
        .Y(n1859) );
  AO22X1_HVT U1828 ( .A1(\ram[7][7] ), .A2(n6913), .A3(n9167), .A4(data[7]), 
        .Y(n1860) );
  AO22X1_HVT U1829 ( .A1(\ram[7][8] ), .A2(n6912), .A3(n9152), .A4(data[8]), 
        .Y(n1861) );
  AO22X1_HVT U1830 ( .A1(\ram[7][9] ), .A2(n6910), .A3(n9151), .A4(n9335), .Y(
        n1862) );
  AO22X1_HVT U1831 ( .A1(\ram[7][10] ), .A2(n6910), .A3(n9150), .A4(data[10]), 
        .Y(n1863) );
  AO22X1_HVT U1832 ( .A1(\ram[7][11] ), .A2(n6908), .A3(n9149), .A4(n9342), 
        .Y(n1864) );
  AO22X1_HVT U1833 ( .A1(\ram[7][12] ), .A2(n6907), .A3(n9146), .A4(data[12]), 
        .Y(n1865) );
  AO22X1_HVT U1834 ( .A1(\ram[7][13] ), .A2(n6905), .A3(n9145), .A4(data[13]), 
        .Y(n1866) );
  AO22X1_HVT U1835 ( .A1(\ram[7][14] ), .A2(n6904), .A3(n9144), .A4(data[14]), 
        .Y(n1867) );
  AO22X1_HVT U1836 ( .A1(\ram[7][15] ), .A2(n6899), .A3(n9143), .A4(data[15]), 
        .Y(n1868) );
  AO22X1_HVT U1837 ( .A1(\ram[7][16] ), .A2(n6937), .A3(n9174), .A4(data[16]), 
        .Y(n1869) );
  AO22X1_HVT U1838 ( .A1(\ram[7][17] ), .A2(n6936), .A3(n9173), .A4(data[17]), 
        .Y(n1870) );
  AO22X1_HVT U1839 ( .A1(\ram[7][18] ), .A2(n6934), .A3(n9172), .A4(n9363), 
        .Y(n1871) );
  AO22X1_HVT U1840 ( .A1(\ram[7][19] ), .A2(n6933), .A3(n9171), .A4(data[19]), 
        .Y(n1872) );
  AO22X1_HVT U1841 ( .A1(\ram[7][20] ), .A2(n6960), .A3(n9174), .A4(n9368), 
        .Y(n1873) );
  AO22X1_HVT U1842 ( .A1(\ram[7][21] ), .A2(n6959), .A3(n9173), .A4(n9371), 
        .Y(n1874) );
  AO22X1_HVT U1843 ( .A1(\ram[7][22] ), .A2(n6957), .A3(n9172), .A4(data[22]), 
        .Y(n1875) );
  AO22X1_HVT U1844 ( .A1(\ram[7][23] ), .A2(n6956), .A3(n9171), .A4(data[23]), 
        .Y(n1876) );
  AO22X1_HVT U1845 ( .A1(\ram[7][24] ), .A2(n6955), .A3(n9184), .A4(data[24]), 
        .Y(n1877) );
  AO22X1_HVT U1846 ( .A1(\ram[7][25] ), .A2(n6954), .A3(n9183), .A4(data[25]), 
        .Y(n1878) );
  AO22X1_HVT U1847 ( .A1(\ram[7][26] ), .A2(n6954), .A3(n9182), .A4(data[26]), 
        .Y(n1879) );
  AO22X1_HVT U1848 ( .A1(\ram[7][27] ), .A2(n6953), .A3(n9181), .A4(data[27]), 
        .Y(n1880) );
  AO22X1_HVT U1849 ( .A1(\ram[7][28] ), .A2(n6952), .A3(n9184), .A4(data[28]), 
        .Y(n1881) );
  AO22X1_HVT U1850 ( .A1(\ram[7][29] ), .A2(n6951), .A3(n9183), .A4(n9395), 
        .Y(n1882) );
  AO22X1_HVT U1851 ( .A1(\ram[7][30] ), .A2(n6950), .A3(n9182), .A4(n9398), 
        .Y(n1883) );
  AO22X1_HVT U1852 ( .A1(\ram[7][31] ), .A2(n6913), .A3(n9181), .A4(data[31]), 
        .Y(n1884) );
  AO22X1_HVT U1853 ( .A1(\ram[7][32] ), .A2(n6912), .A3(n9180), .A4(data[32]), 
        .Y(n1885) );
  AO22X1_HVT U1854 ( .A1(\ram[7][33] ), .A2(n6910), .A3(n9179), .A4(data[33]), 
        .Y(n1886) );
  AO22X1_HVT U1855 ( .A1(\ram[7][34] ), .A2(n6924), .A3(n9178), .A4(data[34]), 
        .Y(n1887) );
  AO22X1_HVT U1856 ( .A1(\ram[7][35] ), .A2(n6921), .A3(n9177), .A4(data[35]), 
        .Y(n1888) );
  AO22X1_HVT U1857 ( .A1(\ram[7][36] ), .A2(n6920), .A3(n9164), .A4(data[36]), 
        .Y(n1889) );
  AO22X1_HVT U1858 ( .A1(\ram[7][37] ), .A2(n6919), .A3(n9163), .A4(data[37]), 
        .Y(n1890) );
  AO22X1_HVT U1859 ( .A1(\ram[7][38] ), .A2(n6916), .A3(n9162), .A4(data[38]), 
        .Y(n1891) );
  AO22X1_HVT U1860 ( .A1(\ram[7][39] ), .A2(n6963), .A3(n9161), .A4(n9425), 
        .Y(n1892) );
  AO22X1_HVT U1861 ( .A1(\ram[7][40] ), .A2(n6947), .A3(n9152), .A4(data[40]), 
        .Y(n1893) );
  AO22X1_HVT U1862 ( .A1(\ram[7][41] ), .A2(n6946), .A3(n9151), .A4(n9431), 
        .Y(n1894) );
  AO22X1_HVT U1863 ( .A1(\ram[7][42] ), .A2(n6902), .A3(n9150), .A4(n9434), 
        .Y(n1895) );
  AO22X1_HVT U1864 ( .A1(\ram[7][43] ), .A2(n6946), .A3(n9149), .A4(data[43]), 
        .Y(n1896) );
  AO22X1_HVT U1865 ( .A1(\ram[7][44] ), .A2(n10268), .A3(n9142), .A4(data[44]), 
        .Y(n1897) );
  AO22X1_HVT U1866 ( .A1(\ram[7][45] ), .A2(n6944), .A3(n9141), .A4(data[45]), 
        .Y(n1898) );
  AO22X1_HVT U1867 ( .A1(\ram[7][46] ), .A2(n6943), .A3(n9140), .A4(data[46]), 
        .Y(n1899) );
  AO22X1_HVT U1868 ( .A1(\ram[7][47] ), .A2(n6942), .A3(n9139), .A4(data[47]), 
        .Y(n1900) );
  AO22X1_HVT U1869 ( .A1(\ram[7][48] ), .A2(n6921), .A3(n9142), .A4(n9452), 
        .Y(n1901) );
  AO22X1_HVT U1870 ( .A1(\ram[7][49] ), .A2(n6920), .A3(n9141), .A4(data[49]), 
        .Y(n1902) );
  AO22X1_HVT U1871 ( .A1(\ram[7][50] ), .A2(n6919), .A3(n9140), .A4(data[50]), 
        .Y(n1903) );
  AO22X1_HVT U1872 ( .A1(\ram[7][51] ), .A2(n6918), .A3(n9139), .A4(n9461), 
        .Y(n1904) );
  AO22X1_HVT U1873 ( .A1(\ram[7][52] ), .A2(n6964), .A3(n9158), .A4(data[52]), 
        .Y(n1905) );
  AO22X1_HVT U1874 ( .A1(\ram[7][53] ), .A2(n6963), .A3(n9157), .A4(n9467), 
        .Y(n1906) );
  AO22X1_HVT U1875 ( .A1(\ram[7][54] ), .A2(n6947), .A3(n9156), .A4(data[54]), 
        .Y(n1907) );
  AO22X1_HVT U1876 ( .A1(\ram[7][55] ), .A2(n6946), .A3(n9155), .A4(data[55]), 
        .Y(n1908) );
  AO22X1_HVT U1877 ( .A1(\ram[7][56] ), .A2(n10265), .A3(n9194), .A4(data[56]), 
        .Y(n1909) );
  AO22X1_HVT U1878 ( .A1(\ram[7][57] ), .A2(n6944), .A3(n9193), .A4(n9479), 
        .Y(n1910) );
  AO22X1_HVT U1879 ( .A1(\ram[7][58] ), .A2(n6905), .A3(n9192), .A4(n9482), 
        .Y(n1911) );
  AO22X1_HVT U1880 ( .A1(\ram[7][59] ), .A2(n6904), .A3(n9191), .A4(n9485), 
        .Y(n1912) );
  AO22X1_HVT U1881 ( .A1(\ram[7][60] ), .A2(n6899), .A3(n9158), .A4(data[60]), 
        .Y(n1913) );
  AO22X1_HVT U1882 ( .A1(\ram[7][61] ), .A2(n6898), .A3(n9157), .A4(data[61]), 
        .Y(n1914) );
  AO22X1_HVT U1883 ( .A1(\ram[7][62] ), .A2(n6897), .A3(n9156), .A4(data[62]), 
        .Y(n1915) );
  AO22X1_HVT U1884 ( .A1(\ram[7][63] ), .A2(n6896), .A3(n9155), .A4(data[63]), 
        .Y(n1916) );
  AO22X1_HVT U1885 ( .A1(\ram[7][64] ), .A2(n6895), .A3(n9146), .A4(data[64]), 
        .Y(n1917) );
  AO22X1_HVT U1886 ( .A1(\ram[7][65] ), .A2(n6917), .A3(n9145), .A4(data[65]), 
        .Y(n1918) );
  AO22X1_HVT U1887 ( .A1(\ram[7][66] ), .A2(n6916), .A3(n9144), .A4(data[66]), 
        .Y(n1919) );
  AO22X1_HVT U1888 ( .A1(\ram[7][67] ), .A2(n6902), .A3(n9143), .A4(data[67]), 
        .Y(n1920) );
  AO22X1_HVT U1889 ( .A1(\ram[7][68] ), .A2(n6896), .A3(n9170), .A4(data[68]), 
        .Y(n1921) );
  AO22X1_HVT U1890 ( .A1(\ram[7][69] ), .A2(n6895), .A3(n9169), .A4(data[69]), 
        .Y(n1922) );
  AO22X1_HVT U1891 ( .A1(\ram[7][70] ), .A2(n6917), .A3(n9168), .A4(data[70]), 
        .Y(n1923) );
  AO22X1_HVT U1892 ( .A1(\ram[7][71] ), .A2(n6916), .A3(n9167), .A4(n9521), 
        .Y(n1924) );
  AO22X1_HVT U1893 ( .A1(\ram[7][72] ), .A2(n6902), .A3(n9142), .A4(data[72]), 
        .Y(n1925) );
  AO22X1_HVT U1894 ( .A1(\ram[7][73] ), .A2(n6924), .A3(n9141), .A4(data[73]), 
        .Y(n1926) );
  AO22X1_HVT U1895 ( .A1(\ram[7][74] ), .A2(n6931), .A3(n9140), .A4(data[74]), 
        .Y(n1927) );
  AO22X1_HVT U1896 ( .A1(\ram[7][75] ), .A2(n6930), .A3(n9139), .A4(n9533), 
        .Y(n1928) );
  AO22X1_HVT U1897 ( .A1(\ram[7][76] ), .A2(n6946), .A3(n9170), .A4(data[76]), 
        .Y(n1929) );
  AO22X1_HVT U1898 ( .A1(\ram[7][77] ), .A2(n10263), .A3(n9169), .A4(data[77]), 
        .Y(n1930) );
  AO22X1_HVT U1899 ( .A1(\ram[7][78] ), .A2(n6944), .A3(n9168), .A4(data[78]), 
        .Y(n1931) );
  AO22X1_HVT U1900 ( .A1(\ram[7][79] ), .A2(n6943), .A3(n9167), .A4(data[79]), 
        .Y(n1932) );
  AO22X1_HVT U1901 ( .A1(\ram[7][80] ), .A2(n6936), .A3(n9180), .A4(data[80]), 
        .Y(n1933) );
  AO22X1_HVT U1902 ( .A1(\ram[7][81] ), .A2(n6912), .A3(n9179), .A4(data[81]), 
        .Y(n1934) );
  AO22X1_HVT U1903 ( .A1(\ram[7][82] ), .A2(n6910), .A3(n9178), .A4(data[82]), 
        .Y(n1935) );
  AO22X1_HVT U1904 ( .A1(\ram[7][83] ), .A2(n6942), .A3(n9177), .A4(data[83]), 
        .Y(n1936) );
  AO22X1_HVT U1905 ( .A1(\ram[7][84] ), .A2(n6939), .A3(n9146), .A4(data[84]), 
        .Y(n1937) );
  AO22X1_HVT U1906 ( .A1(\ram[7][85] ), .A2(n6952), .A3(n9145), .A4(data[85]), 
        .Y(n1938) );
  AO22X1_HVT U1907 ( .A1(\ram[7][86] ), .A2(n6908), .A3(n9144), .A4(data[86]), 
        .Y(n1939) );
  AO22X1_HVT U1908 ( .A1(\ram[7][87] ), .A2(n6907), .A3(n9143), .A4(n9569), 
        .Y(n1940) );
  AO22X1_HVT U1909 ( .A1(\ram[7][88] ), .A2(n6905), .A3(n9174), .A4(data[88]), 
        .Y(n1941) );
  AO22X1_HVT U1910 ( .A1(\ram[7][89] ), .A2(n6904), .A3(n9173), .A4(data[89]), 
        .Y(n1942) );
  AO22X1_HVT U1911 ( .A1(\ram[7][90] ), .A2(n6899), .A3(n9172), .A4(data[90]), 
        .Y(n1943) );
  AO22X1_HVT U1912 ( .A1(\ram[7][91] ), .A2(n6898), .A3(n9171), .A4(data[91]), 
        .Y(n1944) );
  AO22X1_HVT U1913 ( .A1(\ram[7][92] ), .A2(n6897), .A3(n9170), .A4(data[92]), 
        .Y(n1945) );
  AO22X1_HVT U1914 ( .A1(\ram[7][93] ), .A2(n6896), .A3(n9169), .A4(data[93]), 
        .Y(n1946) );
  AO22X1_HVT U1915 ( .A1(\ram[7][94] ), .A2(n6895), .A3(n9168), .A4(data[94]), 
        .Y(n1947) );
  AO22X1_HVT U1916 ( .A1(\ram[7][95] ), .A2(n6910), .A3(n9167), .A4(data[95]), 
        .Y(n1948) );
  AO22X1_HVT U1917 ( .A1(\ram[7][96] ), .A2(n6937), .A3(n9142), .A4(data[96]), 
        .Y(n1949) );
  AO22X1_HVT U1918 ( .A1(\ram[7][97] ), .A2(n6943), .A3(n9141), .A4(data[97]), 
        .Y(n1950) );
  AO22X1_HVT U1919 ( .A1(\ram[7][98] ), .A2(n6942), .A3(n9140), .A4(data[98]), 
        .Y(n1951) );
  AO22X1_HVT U1920 ( .A1(\ram[7][99] ), .A2(n6939), .A3(n9139), .A4(data[99]), 
        .Y(n1952) );
  AO22X1_HVT U1921 ( .A1(\ram[7][100] ), .A2(n6938), .A3(n9194), .A4(data[100]), .Y(n1953) );
  AO22X1_HVT U1922 ( .A1(\ram[7][101] ), .A2(n6937), .A3(n9193), .A4(data[101]), .Y(n1954) );
  AO22X1_HVT U1923 ( .A1(\ram[7][102] ), .A2(n6936), .A3(n9192), .A4(data[102]), .Y(n1955) );
  AO22X1_HVT U1924 ( .A1(\ram[7][103] ), .A2(n6934), .A3(n9191), .A4(data[103]), .Y(n1956) );
  AO22X1_HVT U1925 ( .A1(\ram[7][104] ), .A2(n6933), .A3(n9190), .A4(data[104]), .Y(n1957) );
  AO22X1_HVT U1926 ( .A1(\ram[7][105] ), .A2(n6960), .A3(n9189), .A4(data[105]), .Y(n1958) );
  AO22X1_HVT U1927 ( .A1(\ram[7][106] ), .A2(n6959), .A3(n9188), .A4(data[106]), .Y(n1959) );
  AO22X1_HVT U1928 ( .A1(\ram[7][107] ), .A2(n6957), .A3(n9187), .A4(data[107]), .Y(n1960) );
  AO22X1_HVT U1929 ( .A1(\ram[7][108] ), .A2(n6956), .A3(n9174), .A4(n9632), 
        .Y(n1961) );
  AO22X1_HVT U1930 ( .A1(\ram[7][109] ), .A2(n6953), .A3(n9173), .A4(data[109]), .Y(n1962) );
  AO22X1_HVT U1931 ( .A1(\ram[7][110] ), .A2(n6931), .A3(n9172), .A4(data[110]), .Y(n1963) );
  AO22X1_HVT U1932 ( .A1(\ram[7][111] ), .A2(n6930), .A3(n9171), .A4(data[111]), .Y(n1964) );
  AO22X1_HVT U1933 ( .A1(\ram[7][112] ), .A2(n6927), .A3(n9158), .A4(data[112]), .Y(n1965) );
  AO22X1_HVT U1934 ( .A1(\ram[7][113] ), .A2(n6926), .A3(n9157), .A4(data[113]), .Y(n1966) );
  AO22X1_HVT U1935 ( .A1(\ram[7][114] ), .A2(n6925), .A3(n9156), .A4(data[114]), .Y(n1967) );
  AO22X1_HVT U1936 ( .A1(\ram[7][115] ), .A2(n6924), .A3(n9155), .A4(data[115]), .Y(n1968) );
  AO22X1_HVT U1937 ( .A1(\ram[7][116] ), .A2(n6921), .A3(n9194), .A4(data[116]), .Y(n1969) );
  AO22X1_HVT U1938 ( .A1(\ram[7][117] ), .A2(n6920), .A3(n9193), .A4(data[117]), .Y(n1970) );
  AO22X1_HVT U1939 ( .A1(\ram[7][118] ), .A2(n6919), .A3(n9192), .A4(data[118]), .Y(n1971) );
  AO22X1_HVT U1940 ( .A1(\ram[7][119] ), .A2(n6927), .A3(n9191), .A4(data[119]), .Y(n1972) );
  AO22X1_HVT U1941 ( .A1(\ram[7][120] ), .A2(n6926), .A3(n9180), .A4(data[120]), .Y(n1973) );
  AO22X1_HVT U1942 ( .A1(\ram[7][121] ), .A2(n6925), .A3(n9179), .A4(data[121]), .Y(n1974) );
  AO22X1_HVT U1943 ( .A1(\ram[7][122] ), .A2(n6924), .A3(n9178), .A4(data[122]), .Y(n1975) );
  AO22X1_HVT U1944 ( .A1(\ram[7][123] ), .A2(n6921), .A3(n9177), .A4(data[123]), .Y(n1976) );
  AO22X1_HVT U1945 ( .A1(\ram[7][124] ), .A2(n6920), .A3(n9152), .A4(data[124]), .Y(n1977) );
  AO22X1_HVT U1946 ( .A1(\ram[7][125] ), .A2(n6919), .A3(n9151), .A4(data[125]), .Y(n1978) );
  AO22X1_HVT U1947 ( .A1(\ram[7][126] ), .A2(n6918), .A3(n9150), .A4(data[126]), .Y(n1979) );
  AO22X1_HVT U1948 ( .A1(\ram[7][127] ), .A2(n6942), .A3(n9149), .A4(data[127]), .Y(n1980) );
  AO22X1_HVT U1949 ( .A1(\ram[7][128] ), .A2(n6939), .A3(n9194), .A4(data[128]), .Y(n1981) );
  AO22X1_HVT U1950 ( .A1(\ram[7][129] ), .A2(n6938), .A3(n9193), .A4(data[129]), .Y(n1982) );
  AO22X1_HVT U1951 ( .A1(\ram[7][130] ), .A2(n6937), .A3(n9192), .A4(data[130]), .Y(n1983) );
  AO22X1_HVT U1952 ( .A1(\ram[7][131] ), .A2(n6931), .A3(n9191), .A4(data[131]), .Y(n1984) );
  AO22X1_HVT U1953 ( .A1(\ram[7][132] ), .A2(n6939), .A3(n9152), .A4(data[132]), .Y(n1985) );
  AO22X1_HVT U1954 ( .A1(\ram[7][133] ), .A2(n6938), .A3(n9151), .A4(data[133]), .Y(n1986) );
  AO22X1_HVT U1955 ( .A1(\ram[7][134] ), .A2(n6937), .A3(n9150), .A4(data[134]), .Y(n1987) );
  AO22X1_HVT U1956 ( .A1(\ram[7][135] ), .A2(n6936), .A3(n9149), .A4(data[135]), .Y(n1988) );
  AO22X1_HVT U1957 ( .A1(\ram[7][136] ), .A2(n6934), .A3(n9146), .A4(n9716), 
        .Y(n1989) );
  AO22X1_HVT U1958 ( .A1(\ram[7][137] ), .A2(n6951), .A3(n9145), .A4(data[137]), .Y(n1990) );
  AO22X1_HVT U1959 ( .A1(\ram[7][138] ), .A2(n6950), .A3(n9144), .A4(n9722), 
        .Y(n1991) );
  AO22X1_HVT U1960 ( .A1(\ram[7][139] ), .A2(n6898), .A3(n9143), .A4(n9726), 
        .Y(n1992) );
  AO22X1_HVT U1961 ( .A1(\ram[7][140] ), .A2(n6897), .A3(n9174), .A4(data[140]), .Y(n1993) );
  AO22X1_HVT U1962 ( .A1(\ram[7][141] ), .A2(n6896), .A3(n9173), .A4(data[141]), .Y(n1994) );
  AO22X1_HVT U1963 ( .A1(\ram[7][142] ), .A2(n6895), .A3(n9172), .A4(n9735), 
        .Y(n1995) );
  AO22X1_HVT U1964 ( .A1(\ram[7][143] ), .A2(n6917), .A3(n9171), .A4(n9739), 
        .Y(n1996) );
  AO22X1_HVT U1965 ( .A1(\ram[7][144] ), .A2(n6916), .A3(n9170), .A4(data[144]), .Y(n1997) );
  AO22X1_HVT U1966 ( .A1(\ram[7][145] ), .A2(n6902), .A3(n9169), .A4(n9745), 
        .Y(n1998) );
  AO22X1_HVT U1967 ( .A1(\ram[7][146] ), .A2(n6938), .A3(n9168), .A4(data[146]), .Y(n1999) );
  AO22X1_HVT U1968 ( .A1(\ram[7][147] ), .A2(n6931), .A3(n9167), .A4(n9752), 
        .Y(n2000) );
  AO22X1_HVT U1969 ( .A1(\ram[7][148] ), .A2(n6930), .A3(n9152), .A4(data[148]), .Y(n2001) );
  AO22X1_HVT U1970 ( .A1(\ram[7][149] ), .A2(n6927), .A3(n9151), .A4(data[149]), .Y(n2002) );
  AO22X1_HVT U1971 ( .A1(\ram[7][150] ), .A2(n6926), .A3(n9150), .A4(data[150]), .Y(n2003) );
  AO22X1_HVT U1972 ( .A1(\ram[7][151] ), .A2(n6953), .A3(n9149), .A4(data[151]), .Y(n2004) );
  AO22X1_HVT U1973 ( .A1(\ram[7][152] ), .A2(n6952), .A3(n9146), .A4(n9767), 
        .Y(n2005) );
  AO22X1_HVT U1974 ( .A1(\ram[7][153] ), .A2(n6951), .A3(n9145), .A4(n9770), 
        .Y(n2006) );
  AO22X1_HVT U1975 ( .A1(\ram[7][154] ), .A2(n6950), .A3(n9144), .A4(data[154]), .Y(n2007) );
  AO22X1_HVT U1976 ( .A1(\ram[7][155] ), .A2(n6913), .A3(n9143), .A4(n9777), 
        .Y(n2008) );
  AO22X1_HVT U1977 ( .A1(\ram[7][156] ), .A2(n6912), .A3(n9164), .A4(data[156]), .Y(n2009) );
  AO22X1_HVT U1978 ( .A1(\ram[7][157] ), .A2(n6910), .A3(n9163), .A4(data[157]), .Y(n2010) );
  AO22X1_HVT U1979 ( .A1(\ram[7][158] ), .A2(n6939), .A3(n9162), .A4(data[158]), .Y(n2011) );
  AO22X1_HVT U1980 ( .A1(\ram[7][159] ), .A2(n6908), .A3(n9161), .A4(n9790), 
        .Y(n2012) );
  AO22X1_HVT U1981 ( .A1(\ram[7][160] ), .A2(n6907), .A3(n9164), .A4(n9793), 
        .Y(n2013) );
  AO22X1_HVT U1982 ( .A1(\ram[7][161] ), .A2(n6907), .A3(n9163), .A4(data[161]), .Y(n2014) );
  AO22X1_HVT U1983 ( .A1(\ram[7][162] ), .A2(n6908), .A3(n9162), .A4(data[162]), .Y(n2015) );
  AO22X1_HVT U1984 ( .A1(\ram[7][163] ), .A2(n6907), .A3(n9161), .A4(data[163]), .Y(n2016) );
  AO22X1_HVT U1985 ( .A1(\ram[7][164] ), .A2(n6905), .A3(n9152), .A4(data[164]), .Y(n2017) );
  AO22X1_HVT U1986 ( .A1(\ram[7][165] ), .A2(n6904), .A3(n9151), .A4(n9808), 
        .Y(n2018) );
  AO22X1_HVT U1987 ( .A1(\ram[7][166] ), .A2(n6899), .A3(n9150), .A4(data[166]), .Y(n2019) );
  AO22X1_HVT U1988 ( .A1(\ram[7][167] ), .A2(n6898), .A3(n9149), .A4(n9814), 
        .Y(n2020) );
  AO22X1_HVT U1989 ( .A1(\ram[7][168] ), .A2(n6897), .A3(n9146), .A4(data[168]), .Y(n2021) );
  AO22X1_HVT U1990 ( .A1(\ram[7][169] ), .A2(n6918), .A3(n9145), .A4(data[169]), .Y(n2022) );
  AO22X1_HVT U1991 ( .A1(\ram[7][170] ), .A2(n6964), .A3(n9144), .A4(data[170]), .Y(n2023) );
  AO22X1_HVT U1992 ( .A1(\ram[7][171] ), .A2(n6963), .A3(n9143), .A4(n9827), 
        .Y(n2024) );
  AO22X1_HVT U1993 ( .A1(\ram[7][172] ), .A2(n6947), .A3(n9190), .A4(data[172]), .Y(n2025) );
  AO22X1_HVT U1994 ( .A1(\ram[7][173] ), .A2(n6902), .A3(n9189), .A4(n9833), 
        .Y(n2026) );
  AO22X1_HVT U1995 ( .A1(\ram[7][174] ), .A2(n6933), .A3(n9188), .A4(data[174]), .Y(n2027) );
  AO22X1_HVT U1996 ( .A1(\ram[7][175] ), .A2(n6960), .A3(n9187), .A4(n9840), 
        .Y(n2028) );
  AO22X1_HVT U1997 ( .A1(\ram[7][176] ), .A2(n6944), .A3(n9142), .A4(data[176]), .Y(n2029) );
  AO22X1_HVT U1998 ( .A1(\ram[7][177] ), .A2(n6943), .A3(n9141), .A4(data[177]), .Y(n2030) );
  AO22X1_HVT U1999 ( .A1(\ram[7][178] ), .A2(n6959), .A3(n9140), .A4(data[178]), .Y(n2031) );
  AO22X1_HVT U2000 ( .A1(\ram[7][179] ), .A2(n6957), .A3(n9139), .A4(n9853), 
        .Y(n2032) );
  AO22X1_HVT U2001 ( .A1(\ram[7][180] ), .A2(n6956), .A3(n9158), .A4(data[180]), .Y(n2033) );
  AO22X1_HVT U2002 ( .A1(\ram[7][181] ), .A2(n6955), .A3(n9157), .A4(data[181]), .Y(n2034) );
  AO22X1_HVT U2003 ( .A1(\ram[7][182] ), .A2(n6954), .A3(n9156), .A4(data[182]), .Y(n2035) );
  AO22X1_HVT U2004 ( .A1(\ram[7][183] ), .A2(n6953), .A3(n9155), .A4(n9866), 
        .Y(n2036) );
  AO22X1_HVT U2005 ( .A1(\ram[7][184] ), .A2(n6952), .A3(n9194), .A4(n9869), 
        .Y(n2037) );
  AO22X1_HVT U2006 ( .A1(\ram[7][185] ), .A2(n6951), .A3(n9193), .A4(data[185]), .Y(n2038) );
  AO22X1_HVT U2007 ( .A1(\ram[7][186] ), .A2(n6950), .A3(n9192), .A4(n9875), 
        .Y(n2039) );
  AO22X1_HVT U2008 ( .A1(\ram[7][187] ), .A2(n6913), .A3(n9191), .A4(data[187]), .Y(n2040) );
  AO22X1_HVT U2009 ( .A1(\ram[7][188] ), .A2(n6913), .A3(n9190), .A4(n9881), 
        .Y(n2041) );
  AO22X1_HVT U2010 ( .A1(\ram[7][189] ), .A2(n6912), .A3(n9189), .A4(data[189]), .Y(n2042) );
  AO22X1_HVT U2011 ( .A1(\ram[7][190] ), .A2(n6925), .A3(n9188), .A4(n9887), 
        .Y(n2043) );
  AO22X1_HVT U2012 ( .A1(\ram[7][191] ), .A2(n6924), .A3(n9187), .A4(n9891), 
        .Y(n2044) );
  AO22X1_HVT U2013 ( .A1(\ram[7][192] ), .A2(n6925), .A3(n9190), .A4(data[192]), .Y(n2045) );
  AO22X1_HVT U2014 ( .A1(\ram[7][193] ), .A2(n6931), .A3(n9189), .A4(data[193]), .Y(n2046) );
  AO22X1_HVT U2015 ( .A1(\ram[7][194] ), .A2(n6963), .A3(n9188), .A4(data[194]), .Y(n2047) );
  AO22X1_HVT U2016 ( .A1(\ram[7][195] ), .A2(n6947), .A3(n9187), .A4(n9904), 
        .Y(n2048) );
  AO22X1_HVT U2017 ( .A1(\ram[7][196] ), .A2(n6930), .A3(n9184), .A4(data[196]), .Y(n2049) );
  AO22X1_HVT U2018 ( .A1(\ram[7][197] ), .A2(n6927), .A3(n9183), .A4(data[197]), .Y(n2050) );
  AO22X1_HVT U2019 ( .A1(\ram[7][198] ), .A2(n6926), .A3(n9182), .A4(data[198]), .Y(n2051) );
  AO22X1_HVT U2020 ( .A1(\ram[7][199] ), .A2(n6925), .A3(n9181), .A4(n9917), 
        .Y(n2052) );
  AO22X1_HVT U2021 ( .A1(\ram[7][200] ), .A2(n6924), .A3(n9184), .A4(data[200]), .Y(n2053) );
  AO22X1_HVT U2022 ( .A1(\ram[7][201] ), .A2(n6921), .A3(n9183), .A4(data[201]), .Y(n2054) );
  AO22X1_HVT U2023 ( .A1(\ram[7][202] ), .A2(n6920), .A3(n9182), .A4(data[202]), .Y(n2055) );
  AO22X1_HVT U2024 ( .A1(\ram[7][203] ), .A2(n6919), .A3(n9181), .A4(n9929), 
        .Y(n2056) );
  AO22X1_HVT U2025 ( .A1(\ram[7][204] ), .A2(n6964), .A3(n9194), .A4(n9932), 
        .Y(n2057) );
  AO22X1_HVT U2026 ( .A1(\ram[7][205] ), .A2(n6905), .A3(n9193), .A4(data[205]), .Y(n2058) );
  AO22X1_HVT U2027 ( .A1(\ram[7][206] ), .A2(n6904), .A3(n9192), .A4(data[206]), .Y(n2059) );
  AO22X1_HVT U2028 ( .A1(\ram[7][207] ), .A2(n6899), .A3(n9191), .A4(n9942), 
        .Y(n2060) );
  AO22X1_HVT U2029 ( .A1(\ram[7][208] ), .A2(n6898), .A3(n9190), .A4(data[208]), .Y(n2061) );
  AO22X1_HVT U2030 ( .A1(\ram[7][209] ), .A2(n6897), .A3(n9189), .A4(n9948), 
        .Y(n2062) );
  AO22X1_HVT U2031 ( .A1(\ram[7][210] ), .A2(n6896), .A3(n9188), .A4(data[210]), .Y(n2063) );
  AO22X1_HVT U2032 ( .A1(\ram[7][211] ), .A2(n6895), .A3(n9187), .A4(data[211]), .Y(n2064) );
  AO22X1_HVT U2033 ( .A1(\ram[7][212] ), .A2(n6917), .A3(n9164), .A4(data[212]), .Y(n2065) );
  AO22X1_HVT U2034 ( .A1(\ram[7][213] ), .A2(n6916), .A3(n9163), .A4(data[213]), .Y(n2066) );
  AO22X1_HVT U2035 ( .A1(\ram[7][214] ), .A2(n6902), .A3(n9162), .A4(data[214]), .Y(n2067) );
  AO22X1_HVT U2036 ( .A1(\ram[7][215] ), .A2(n6955), .A3(n9161), .A4(data[215]), .Y(n2068) );
  AO22X1_HVT U2037 ( .A1(\ram[7][216] ), .A2(n6954), .A3(n9158), .A4(data[216]), .Y(n2069) );
  AO22X1_HVT U2038 ( .A1(\ram[7][217] ), .A2(n6938), .A3(n9157), .A4(data[217]), .Y(n2070) );
  AO22X1_HVT U2039 ( .A1(\ram[7][218] ), .A2(n6937), .A3(n9156), .A4(data[218]), .Y(n2071) );
  AO22X1_HVT U2040 ( .A1(\ram[7][219] ), .A2(n6936), .A3(n9155), .A4(n9979), 
        .Y(n2072) );
  AO22X1_HVT U2041 ( .A1(\ram[7][220] ), .A2(n6934), .A3(n9190), .A4(data[220]), .Y(n2073) );
  AO22X1_HVT U2042 ( .A1(\ram[7][221] ), .A2(n6933), .A3(n9189), .A4(data[221]), .Y(n2074) );
  AO22X1_HVT U2043 ( .A1(\ram[7][222] ), .A2(n6960), .A3(n9188), .A4(n9988), 
        .Y(n2075) );
  AO22X1_HVT U2044 ( .A1(\ram[7][223] ), .A2(n6959), .A3(n9187), .A4(n9991), 
        .Y(n2076) );
  AO22X1_HVT U2045 ( .A1(\ram[7][224] ), .A2(n6957), .A3(n9184), .A4(data[224]), .Y(n2077) );
  AO22X1_HVT U2046 ( .A1(\ram[7][225] ), .A2(n6956), .A3(n9183), .A4(data[225]), .Y(n2078) );
  AO22X1_HVT U2047 ( .A1(\ram[7][226] ), .A2(n6955), .A3(n9182), .A4(data[226]), .Y(n2079) );
  AO22X1_HVT U2048 ( .A1(\ram[7][227] ), .A2(n6954), .A3(n9181), .A4(data[227]), .Y(n2080) );
  AO22X1_HVT U2049 ( .A1(\ram[7][228] ), .A2(n6953), .A3(n9180), .A4(data[228]), .Y(n2081) );
  AO22X1_HVT U2050 ( .A1(\ram[7][229] ), .A2(n6964), .A3(n9179), .A4(data[229]), .Y(n2082) );
  AO22X1_HVT U2051 ( .A1(\ram[7][230] ), .A2(n6963), .A3(n9178), .A4(data[230]), .Y(n2083) );
  AO22X1_HVT U2052 ( .A1(\ram[7][231] ), .A2(n6947), .A3(n9177), .A4(n10016), 
        .Y(n2084) );
  AO22X1_HVT U2053 ( .A1(\ram[7][232] ), .A2(n6946), .A3(n9164), .A4(data[232]), .Y(n2085) );
  AO22X1_HVT U2054 ( .A1(\ram[7][233] ), .A2(n10265), .A3(n9163), .A4(n10022), 
        .Y(n2086) );
  AO22X1_HVT U2055 ( .A1(\ram[7][234] ), .A2(n6944), .A3(n9162), .A4(n10025), 
        .Y(n2087) );
  AO22X1_HVT U2056 ( .A1(\ram[7][235] ), .A2(n6943), .A3(n9161), .A4(data[235]), .Y(n2088) );
  AO22X1_HVT U2057 ( .A1(\ram[7][236] ), .A2(n6942), .A3(n9180), .A4(data[236]), .Y(n2089) );
  AO22X1_HVT U2058 ( .A1(\ram[7][237] ), .A2(n6939), .A3(n9179), .A4(n10034), 
        .Y(n2090) );
  AO22X1_HVT U2059 ( .A1(\ram[7][238] ), .A2(n6938), .A3(n9178), .A4(data[238]), .Y(n2091) );
  AO22X1_HVT U2060 ( .A1(\ram[7][239] ), .A2(n6936), .A3(n9177), .A4(n10041), 
        .Y(n2092) );
  AO22X1_HVT U2061 ( .A1(\ram[7][240] ), .A2(n6934), .A3(n9164), .A4(n10044), 
        .Y(n2093) );
  AO22X1_HVT U2062 ( .A1(\ram[7][241] ), .A2(n6933), .A3(n9163), .A4(data[241]), .Y(n2094) );
  AO22X1_HVT U2063 ( .A1(\ram[7][242] ), .A2(n6960), .A3(n9162), .A4(data[242]), .Y(n2095) );
  AO22X1_HVT U2064 ( .A1(\ram[7][243] ), .A2(n6959), .A3(n9161), .A4(data[243]), .Y(n2096) );
  AO22X1_HVT U2065 ( .A1(\ram[7][244] ), .A2(n6957), .A3(n9180), .A4(data[244]), .Y(n2097) );
  AO22X1_HVT U2066 ( .A1(\ram[7][245] ), .A2(n6956), .A3(n9179), .A4(n10059), 
        .Y(n2098) );
  AO22X1_HVT U2067 ( .A1(\ram[7][246] ), .A2(n6955), .A3(n9178), .A4(data[246]), .Y(n2099) );
  AO22X1_HVT U2068 ( .A1(\ram[7][247] ), .A2(n6930), .A3(n9177), .A4(n10066), 
        .Y(n2100) );
  AO22X1_HVT U2069 ( .A1(\ram[7][248] ), .A2(n6927), .A3(n9184), .A4(data[248]), .Y(n2101) );
  AO22X1_HVT U2070 ( .A1(\ram[7][249] ), .A2(n6926), .A3(n9183), .A4(data[249]), .Y(n2102) );
  AO22X1_HVT U2071 ( .A1(\ram[7][250] ), .A2(n6925), .A3(n9182), .A4(data[250]), .Y(n2103) );
  AO22X1_HVT U2072 ( .A1(\ram[7][251] ), .A2(n6917), .A3(n9181), .A4(n10079), 
        .Y(n2104) );
  AO22X1_HVT U2073 ( .A1(\ram[7][252] ), .A2(n6895), .A3(n9170), .A4(n10082), 
        .Y(n2105) );
  AO22X1_HVT U2074 ( .A1(\ram[7][253] ), .A2(n6908), .A3(n9169), .A4(data[253]), .Y(n2106) );
  AO22X1_HVT U2075 ( .A1(\ram[7][254] ), .A2(n6907), .A3(n9168), .A4(data[254]), .Y(n2107) );
  AO22X1_HVT U2076 ( .A1(\ram[7][255] ), .A2(n6918), .A3(n9167), .A4(n10092), 
        .Y(n2108) );
  AND2X1_HVT U2077 ( .A1(n34), .A2(n5645), .Y(n33) );
  AND2X1_HVT U2079 ( .A1(n5511), .A2(n5620), .Y(n34) );
  AND2X1_HVT U2080 ( .A1(n7714), .A2(n7544), .Y(n25) );
  AO22X1_HVT U2081 ( .A1(\ram[8][0] ), .A2(n4238), .A3(n6040), .A4(n9307), .Y(
        n2109) );
  AO22X1_HVT U2082 ( .A1(\ram[8][1] ), .A2(n7414), .A3(n6070), .A4(n9310), .Y(
        n2110) );
  AO22X1_HVT U2083 ( .A1(\ram[8][2] ), .A2(n4647), .A3(n6039), .A4(n9312), .Y(
        n2111) );
  AO22X1_HVT U2084 ( .A1(\ram[8][3] ), .A2(n7384), .A3(n6075), .A4(n9316), .Y(
        n2112) );
  AO22X1_HVT U2085 ( .A1(\ram[8][4] ), .A2(n7383), .A3(n6074), .A4(n9320), .Y(
        n2113) );
  AO22X1_HVT U2086 ( .A1(\ram[8][5] ), .A2(n4349), .A3(n6073), .A4(n9323), .Y(
        n2114) );
  AO22X1_HVT U2087 ( .A1(\ram[8][6] ), .A2(n4377), .A3(n6072), .A4(n9326), .Y(
        n2115) );
  AO22X1_HVT U2088 ( .A1(\ram[8][7] ), .A2(n7354), .A3(n6071), .A4(n9329), .Y(
        n2116) );
  AO22X1_HVT U2089 ( .A1(\ram[8][8] ), .A2(n7380), .A3(n6070), .A4(n9332), .Y(
        n2117) );
  AO22X1_HVT U2090 ( .A1(\ram[8][9] ), .A2(n10248), .A3(n6068), .A4(n9335), 
        .Y(n2118) );
  AO22X1_HVT U2091 ( .A1(\ram[8][10] ), .A2(n7377), .A3(n6067), .A4(n9338), 
        .Y(n2119) );
  AO22X1_HVT U2093 ( .A1(\ram[8][12] ), .A2(n7361), .A3(n6065), .A4(n9345), 
        .Y(n2121) );
  AO22X1_HVT U2094 ( .A1(\ram[8][13] ), .A2(n7374), .A3(n6062), .A4(n9348), 
        .Y(n2122) );
  AO22X1_HVT U2095 ( .A1(\ram[8][14] ), .A2(n4581), .A3(n6061), .A4(n9351), 
        .Y(n2123) );
  AO22X1_HVT U2097 ( .A1(\ram[8][16] ), .A2(n7390), .A3(n6045), .A4(n9357), 
        .Y(n2125) );
  AO22X1_HVT U2100 ( .A1(\ram[8][19] ), .A2(n7367), .A3(n6049), .A4(n9366), 
        .Y(n2128) );
  AO22X1_HVT U2101 ( .A1(\ram[8][20] ), .A2(n7366), .A3(n6085), .A4(n9368), 
        .Y(n2129) );
  AO22X1_HVT U2102 ( .A1(\ram[8][21] ), .A2(n7365), .A3(n6048), .A4(n9371), 
        .Y(n2130) );
  AO22X1_HVT U2103 ( .A1(\ram[8][22] ), .A2(n7379), .A3(n6042), .A4(n9374), 
        .Y(n2131) );
  AO22X1_HVT U2104 ( .A1(\ram[8][23] ), .A2(n7374), .A3(n6041), .A4(n9377), 
        .Y(n2132) );
  AO22X1_HVT U2105 ( .A1(\ram[8][24] ), .A2(n7395), .A3(n6040), .A4(n9380), 
        .Y(n2133) );
  AO22X1_HVT U2108 ( .A1(\ram[8][27] ), .A2(n7373), .A3(n6065), .A4(n9389), 
        .Y(n2136) );
  AO22X1_HVT U2109 ( .A1(\ram[8][28] ), .A2(n7396), .A3(n6062), .A4(n9392), 
        .Y(n2137) );
  AO22X1_HVT U2110 ( .A1(\ram[8][29] ), .A2(n7388), .A3(n6061), .A4(n9395), 
        .Y(n2138) );
  AO22X1_HVT U2111 ( .A1(\ram[8][30] ), .A2(n7387), .A3(n6042), .A4(data[30]), 
        .Y(n2139) );
  AO22X1_HVT U2112 ( .A1(\ram[8][31] ), .A2(n7369), .A3(n6074), .A4(n9401), 
        .Y(n2140) );
  AO22X1_HVT U2114 ( .A1(\ram[8][33] ), .A2(n7378), .A3(n6108), .A4(n9407), 
        .Y(n2142) );
  AO22X1_HVT U2115 ( .A1(\ram[8][34] ), .A2(n7411), .A3(n6107), .A4(n9410), 
        .Y(n2143) );
  AO22X1_HVT U2116 ( .A1(\ram[8][35] ), .A2(n4345), .A3(n6105), .A4(n9413), 
        .Y(n2144) );
  AO22X1_HVT U2117 ( .A1(\ram[8][36] ), .A2(n7411), .A3(n6104), .A4(n9416), 
        .Y(n2145) );
  AO22X1_HVT U2118 ( .A1(\ram[8][37] ), .A2(n7408), .A3(n6102), .A4(n9419), 
        .Y(n2146) );
  AO22X1_HVT U2119 ( .A1(\ram[8][38] ), .A2(n7406), .A3(n6061), .A4(n9422), 
        .Y(n2147) );
  AO22X1_HVT U2121 ( .A1(\ram[8][40] ), .A2(n7402), .A3(n6099), .A4(n9428), 
        .Y(n2149) );
  AO22X1_HVT U2122 ( .A1(\ram[8][41] ), .A2(n7401), .A3(n6096), .A4(n9431), 
        .Y(n2150) );
  AO22X1_HVT U2123 ( .A1(\ram[8][42] ), .A2(n7400), .A3(n6095), .A4(n9434), 
        .Y(n2151) );
  AO22X1_HVT U2124 ( .A1(\ram[8][43] ), .A2(n7371), .A3(n6093), .A4(n9437), 
        .Y(n2152) );
  AO22X1_HVT U2125 ( .A1(\ram[8][44] ), .A2(n7370), .A3(n6089), .A4(n9440), 
        .Y(n2153) );
  AO22X1_HVT U2126 ( .A1(\ram[8][45] ), .A2(n7369), .A3(n6088), .A4(n9443), 
        .Y(n2154) );
  AO22X1_HVT U2127 ( .A1(\ram[8][46] ), .A2(n4353), .A3(n6100), .A4(n9446), 
        .Y(n2155) );
  AO22X1_HVT U2129 ( .A1(\ram[8][48] ), .A2(n7396), .A3(n6048), .A4(n9452), 
        .Y(n2157) );
  AO22X1_HVT U2130 ( .A1(\ram[8][49] ), .A2(n7361), .A3(n6100), .A4(n9455), 
        .Y(n2158) );
  AO22X1_HVT U2131 ( .A1(\ram[8][50] ), .A2(n7361), .A3(n6087), .A4(n9458), 
        .Y(n2159) );
  AO22X1_HVT U2132 ( .A1(\ram[8][51] ), .A2(n7357), .A3(n6045), .A4(n9461), 
        .Y(n2160) );
  AO22X1_HVT U2133 ( .A1(\ram[8][52] ), .A2(n7356), .A3(n6111), .A4(n9464), 
        .Y(n2161) );
  AO22X1_HVT U2134 ( .A1(\ram[8][53] ), .A2(n7417), .A3(n6104), .A4(n9467), 
        .Y(n2162) );
  AO22X1_HVT U2135 ( .A1(\ram[8][54] ), .A2(n4214), .A3(n6102), .A4(n9470), 
        .Y(n2163) );
  AO22X1_HVT U2136 ( .A1(\ram[8][55] ), .A2(n4238), .A3(n6049), .A4(n9473), 
        .Y(n2164) );
  AO22X1_HVT U2137 ( .A1(\ram[8][56] ), .A2(n7414), .A3(n6101), .A4(n9476), 
        .Y(n2165) );
  AO22X1_HVT U2138 ( .A1(\ram[8][57] ), .A2(n7360), .A3(n6061), .A4(n9479), 
        .Y(n2166) );
  AO22X1_HVT U2140 ( .A1(\ram[8][59] ), .A2(n7383), .A3(n6112), .A4(n9485), 
        .Y(n2168) );
  AO22X1_HVT U2141 ( .A1(\ram[8][60] ), .A2(n4580), .A3(n6041), .A4(n9488), 
        .Y(n2169) );
  AO22X1_HVT U2142 ( .A1(\ram[8][61] ), .A2(n7394), .A3(n6104), .A4(n9491), 
        .Y(n2170) );
  AO22X1_HVT U2143 ( .A1(\ram[8][62] ), .A2(n7371), .A3(n4356), .A4(n9494), 
        .Y(n2171) );
  AO22X1_HVT U2144 ( .A1(\ram[8][63] ), .A2(n7370), .A3(n6111), .A4(n9497), 
        .Y(n2172) );
  AO22X1_HVT U2145 ( .A1(\ram[8][64] ), .A2(n7365), .A3(n6105), .A4(n9500), 
        .Y(n2173) );
  AO22X1_HVT U2146 ( .A1(\ram[8][65] ), .A2(n7364), .A3(n6100), .A4(n9503), 
        .Y(n2174) );
  AO22X1_HVT U2147 ( .A1(\ram[8][66] ), .A2(n7360), .A3(n6042), .A4(n9506), 
        .Y(n2175) );
  AO22X1_HVT U2148 ( .A1(\ram[8][67] ), .A2(n4349), .A3(n6102), .A4(n9509), 
        .Y(n2176) );
  AO22X1_HVT U2149 ( .A1(\ram[8][68] ), .A2(n7357), .A3(n6084), .A4(n9512), 
        .Y(n2177) );
  AO22X1_HVT U2150 ( .A1(\ram[8][69] ), .A2(n7356), .A3(n6112), .A4(n9515), 
        .Y(n2178) );
  AO22X1_HVT U2151 ( .A1(\ram[8][70] ), .A2(n7417), .A3(n6107), .A4(n9518), 
        .Y(n2179) );
  AO22X1_HVT U2152 ( .A1(\ram[8][71] ), .A2(n4606), .A3(n6085), .A4(n9521), 
        .Y(n2180) );
  AO22X1_HVT U2153 ( .A1(\ram[8][72] ), .A2(n7367), .A3(n6051), .A4(n9524), 
        .Y(n2181) );
  AO22X1_HVT U2154 ( .A1(\ram[8][73] ), .A2(n7366), .A3(n6096), .A4(n9527), 
        .Y(n2182) );
  AO22X1_HVT U2155 ( .A1(\ram[8][74] ), .A2(n7391), .A3(n6079), .A4(n9530), 
        .Y(n2183) );
  AO22X1_HVT U2156 ( .A1(\ram[8][75] ), .A2(n7390), .A3(n6107), .A4(n9533), 
        .Y(n2184) );
  AO22X1_HVT U2157 ( .A1(\ram[8][76] ), .A2(n7354), .A3(n6102), .A4(n9536), 
        .Y(n2185) );
  AO22X1_HVT U2158 ( .A1(\ram[8][77] ), .A2(n7354), .A3(n6101), .A4(n9539), 
        .Y(n2186) );
  AO22X1_HVT U2159 ( .A1(\ram[8][78] ), .A2(n7379), .A3(n6050), .A4(n9542), 
        .Y(n2187) );
  AO22X1_HVT U2160 ( .A1(\ram[8][79] ), .A2(n7413), .A3(n6099), .A4(n9545), 
        .Y(n2188) );
  AO22X1_HVT U2161 ( .A1(\ram[8][80] ), .A2(n7377), .A3(n6082), .A4(n9548), 
        .Y(n2189) );
  AO22X1_HVT U2162 ( .A1(\ram[8][81] ), .A2(n7375), .A3(n6108), .A4(n9551), 
        .Y(n2190) );
  AO22X1_HVT U2163 ( .A1(\ram[8][82] ), .A2(n10240), .A3(n6104), .A4(n9554), 
        .Y(n2191) );
  AO22X1_HVT U2164 ( .A1(\ram[8][83] ), .A2(n7374), .A3(n6099), .A4(n9557), 
        .Y(n2192) );
  AO22X1_HVT U2165 ( .A1(\ram[8][84] ), .A2(n7400), .A3(n6105), .A4(n9560), 
        .Y(n2193) );
  AO22X1_HVT U2166 ( .A1(\ram[8][85] ), .A2(n7399), .A3(n6088), .A4(n9563), 
        .Y(n2194) );
  AO22X1_HVT U2167 ( .A1(\ram[8][86] ), .A2(n7398), .A3(n6108), .A4(n9566), 
        .Y(n2195) );
  AO22X1_HVT U2168 ( .A1(\ram[8][87] ), .A2(n10246), .A3(n6085), .A4(n9569), 
        .Y(n2196) );
  AO22X1_HVT U2169 ( .A1(\ram[8][88] ), .A2(n7397), .A3(n6083), .A4(n9572), 
        .Y(n2197) );
  AO22X1_HVT U2170 ( .A1(\ram[8][89] ), .A2(n7372), .A3(n6071), .A4(n9575), 
        .Y(n2198) );
  AO22X1_HVT U2171 ( .A1(\ram[8][90] ), .A2(n7397), .A3(n6083), .A4(n9578), 
        .Y(n2199) );
  AO22X1_HVT U2172 ( .A1(\ram[8][91] ), .A2(n7379), .A3(n6089), .A4(n9581), 
        .Y(n2200) );
  AO22X1_HVT U2173 ( .A1(\ram[8][92] ), .A2(n10248), .A3(n6054), .A4(n9584), 
        .Y(n2201) );
  AO22X1_HVT U2174 ( .A1(\ram[8][93] ), .A2(n7377), .A3(n6062), .A4(n9587), 
        .Y(n2202) );
  AO22X1_HVT U2175 ( .A1(\ram[8][94] ), .A2(n7375), .A3(n6045), .A4(n9590), 
        .Y(n2203) );
  AO22X1_HVT U2176 ( .A1(\ram[8][95] ), .A2(n7384), .A3(n6096), .A4(n9593), 
        .Y(n2204) );
  AO22X1_HVT U2177 ( .A1(\ram[8][96] ), .A2(n7399), .A3(n6084), .A4(n9596), 
        .Y(n2205) );
  AO22X1_HVT U2178 ( .A1(\ram[8][97] ), .A2(n7398), .A3(n6090), .A4(n9599), 
        .Y(n2206) );
  AO22X1_HVT U2179 ( .A1(\ram[8][98] ), .A2(n10246), .A3(n6055), .A4(n9602), 
        .Y(n2207) );
  AO22X1_HVT U2180 ( .A1(\ram[8][99] ), .A2(n7397), .A3(n6062), .A4(n9605), 
        .Y(n2208) );
  AO22X1_HVT U2181 ( .A1(\ram[8][100] ), .A2(n7394), .A3(n6054), .A4(n9608), 
        .Y(n2209) );
  AO22X1_HVT U2182 ( .A1(\ram[8][101] ), .A2(n4580), .A3(n6099), .A4(n9611), 
        .Y(n2210) );
  AO22X1_HVT U2183 ( .A1(\ram[8][102] ), .A2(n7396), .A3(n6039), .A4(n9614), 
        .Y(n2211) );
  AO22X1_HVT U2184 ( .A1(\ram[8][103] ), .A2(n7391), .A3(n6092), .A4(n9617), 
        .Y(n2212) );
  AO22X1_HVT U2185 ( .A1(\ram[8][104] ), .A2(n7390), .A3(n6058), .A4(n9620), 
        .Y(n2213) );
  AO22X1_HVT U2186 ( .A1(\ram[8][105] ), .A2(n7388), .A3(n6085), .A4(n9623), 
        .Y(n2214) );
  AO22X1_HVT U2187 ( .A1(\ram[8][106] ), .A2(n7387), .A3(n6055), .A4(n9626), 
        .Y(n2215) );
  AO22X1_HVT U2188 ( .A1(\ram[8][107] ), .A2(n7401), .A3(n6100), .A4(n9629), 
        .Y(n2216) );
  AO22X1_HVT U2189 ( .A1(\ram[8][108] ), .A2(n7372), .A3(n6042), .A4(n9632), 
        .Y(n2217) );
  AO22X1_HVT U2190 ( .A1(\ram[8][109] ), .A2(n4353), .A3(n6093), .A4(n9635), 
        .Y(n2218) );
  AO22X1_HVT U2191 ( .A1(\ram[8][110] ), .A2(n4353), .A3(n6059), .A4(n9638), 
        .Y(n2219) );
  AO22X1_HVT U2192 ( .A1(\ram[8][111] ), .A2(n7409), .A3(n6065), .A4(n9641), 
        .Y(n2220) );
  AO22X1_HVT U2193 ( .A1(\ram[8][112] ), .A2(n7412), .A3(n6058), .A4(n9644), 
        .Y(n2221) );
  AO22X1_HVT U2194 ( .A1(\ram[8][113] ), .A2(n7409), .A3(n6107), .A4(n9647), 
        .Y(n2222) );
  AO22X1_HVT U2195 ( .A1(\ram[8][114] ), .A2(n7408), .A3(n6040), .A4(n9650), 
        .Y(n2223) );
  AO22X1_HVT U2196 ( .A1(\ram[8][115] ), .A2(n7406), .A3(n6095), .A4(n9653), 
        .Y(n2224) );
  AO22X1_HVT U2197 ( .A1(\ram[8][116] ), .A2(n7405), .A3(n6078), .A4(n9656), 
        .Y(n2225) );
  AO22X1_HVT U2198 ( .A1(\ram[8][117] ), .A2(n7402), .A3(n6066), .A4(n9659), 
        .Y(n2226) );
  AO22X1_HVT U2199 ( .A1(\ram[8][118] ), .A2(n7401), .A3(n6072), .A4(n9662), 
        .Y(n2227) );
  AO22X1_HVT U2200 ( .A1(\ram[8][119] ), .A2(n7400), .A3(n6105), .A4(n9665), 
        .Y(n2228) );
  AO22X1_HVT U2201 ( .A1(\ram[8][120] ), .A2(n4345), .A3(n6039), .A4(n9668), 
        .Y(n2229) );
  AO22X1_HVT U2202 ( .A1(\ram[8][121] ), .A2(n4345), .A3(n6051), .A4(n9671), 
        .Y(n2230) );
  AO22X1_HVT U2203 ( .A1(\ram[8][122] ), .A2(n7412), .A3(n6050), .A4(n9674), 
        .Y(n2231) );
  AO22X1_HVT U2204 ( .A1(\ram[8][123] ), .A2(n7408), .A3(n6049), .A4(n9677), 
        .Y(n2232) );
  AO22X1_HVT U2205 ( .A1(\ram[8][124] ), .A2(n7406), .A3(n6048), .A4(n9680), 
        .Y(n2233) );
  AO22X1_HVT U2206 ( .A1(\ram[8][125] ), .A2(n4647), .A3(n6042), .A4(n9683), 
        .Y(n2234) );
  AO22X1_HVT U2207 ( .A1(\ram[8][126] ), .A2(n7402), .A3(n6041), .A4(n9686), 
        .Y(n2235) );
  AO22X1_HVT U2208 ( .A1(\ram[8][127] ), .A2(n7401), .A3(n6040), .A4(n9689), 
        .Y(n2236) );
  AO22X1_HVT U2209 ( .A1(\ram[8][128] ), .A2(n7400), .A3(n6041), .A4(n9692), 
        .Y(n2237) );
  AO22X1_HVT U2210 ( .A1(\ram[8][129] ), .A2(n7399), .A3(n6039), .A4(n9695), 
        .Y(n2238) );
  AO22X1_HVT U2211 ( .A1(\ram[8][130] ), .A2(n7398), .A3(n6075), .A4(n9698), 
        .Y(n2239) );
  AO22X1_HVT U2212 ( .A1(\ram[8][131] ), .A2(n4647), .A3(n6074), .A4(n9701), 
        .Y(n2240) );
  AO22X1_HVT U2213 ( .A1(\ram[8][132] ), .A2(n7395), .A3(n6101), .A4(n9704), 
        .Y(n2241) );
  AO22X1_HVT U2214 ( .A1(\ram[8][133] ), .A2(n7396), .A3(n6087), .A4(n9707), 
        .Y(n2242) );
  AO22X1_HVT U2215 ( .A1(\ram[8][134] ), .A2(n7395), .A3(n6045), .A4(n9710), 
        .Y(n2243) );
  AO22X1_HVT U2216 ( .A1(\ram[8][135] ), .A2(n7394), .A3(n6112), .A4(n9713), 
        .Y(n2244) );
  AO22X1_HVT U2217 ( .A1(\ram[8][136] ), .A2(n7391), .A3(n6092), .A4(n9716), 
        .Y(n2245) );
  AO22X1_HVT U2218 ( .A1(\ram[8][137] ), .A2(n7364), .A3(n6090), .A4(n9719), 
        .Y(n2246) );
  AO22X1_HVT U2219 ( .A1(\ram[8][138] ), .A2(n4349), .A3(n6111), .A4(n9722), 
        .Y(n2247) );
  AO22X1_HVT U2220 ( .A1(\ram[8][139] ), .A2(n7360), .A3(n6108), .A4(n9725), 
        .Y(n2248) );
  AO22X1_HVT U2221 ( .A1(\ram[8][140] ), .A2(n7357), .A3(n6107), .A4(n9729), 
        .Y(n2249) );
  AO22X1_HVT U2222 ( .A1(\ram[8][141] ), .A2(n7356), .A3(n6105), .A4(n9732), 
        .Y(n2250) );
  AO22X1_HVT U2223 ( .A1(\ram[8][142] ), .A2(n7417), .A3(n6104), .A4(data[142]), .Y(n2251) );
  AO22X1_HVT U2224 ( .A1(\ram[8][143] ), .A2(n4606), .A3(n6102), .A4(n9738), 
        .Y(n2252) );
  AO22X1_HVT U2225 ( .A1(\ram[8][144] ), .A2(n4238), .A3(n6068), .A4(n9742), 
        .Y(n2253) );
  AO22X1_HVT U2226 ( .A1(\ram[8][145] ), .A2(n7371), .A3(n6067), .A4(n9745), 
        .Y(n2254) );
  AO22X1_HVT U2227 ( .A1(\ram[8][146] ), .A2(n7370), .A3(n6066), .A4(n9748), 
        .Y(n2255) );
  AO22X1_HVT U2228 ( .A1(\ram[8][147] ), .A2(n7369), .A3(n6075), .A4(n9751), 
        .Y(n2256) );
  AO22X1_HVT U2229 ( .A1(\ram[8][148] ), .A2(n7378), .A3(n6072), .A4(n9755), 
        .Y(n2257) );
  AO22X1_HVT U2230 ( .A1(\ram[8][149] ), .A2(n10242), .A3(n6071), .A4(n9758), 
        .Y(n2258) );
  AO22X1_HVT U2231 ( .A1(\ram[8][150] ), .A2(n7390), .A3(n6070), .A4(n9761), 
        .Y(n2259) );
  AO22X1_HVT U2232 ( .A1(\ram[8][151] ), .A2(n7388), .A3(n6068), .A4(n9764), 
        .Y(n2260) );
  AO22X1_HVT U2233 ( .A1(\ram[8][152] ), .A2(n7367), .A3(n6067), .A4(n9767), 
        .Y(n2261) );
  AO22X1_HVT U2234 ( .A1(\ram[8][153] ), .A2(n7366), .A3(n6066), .A4(n9770), 
        .Y(n2262) );
  AO22X1_HVT U2235 ( .A1(\ram[8][154] ), .A2(n7399), .A3(n6065), .A4(n9773), 
        .Y(n2263) );
  AO22X1_HVT U2236 ( .A1(\ram[8][155] ), .A2(n7398), .A3(n6062), .A4(n9776), 
        .Y(n2264) );
  AO22X1_HVT U2237 ( .A1(\ram[8][156] ), .A2(n7416), .A3(n6048), .A4(n9780), 
        .Y(n2265) );
  AO22X1_HVT U2238 ( .A1(\ram[8][157] ), .A2(n7373), .A3(n6042), .A4(n9783), 
        .Y(n2266) );
  AO22X1_HVT U2239 ( .A1(\ram[8][158] ), .A2(n7394), .A3(n6041), .A4(n9786), 
        .Y(n2267) );
  AO22X1_HVT U2240 ( .A1(\ram[8][159] ), .A2(n7373), .A3(n6082), .A4(n9789), 
        .Y(n2268) );
  AO22X1_HVT U2241 ( .A1(\ram[8][160] ), .A2(n7372), .A3(n6079), .A4(n9793), 
        .Y(n2269) );
  AO22X1_HVT U2242 ( .A1(\ram[8][161] ), .A2(n7391), .A3(n6078), .A4(n9796), 
        .Y(n2270) );
  AO22X1_HVT U2243 ( .A1(\ram[8][162] ), .A2(n7390), .A3(n6059), .A4(n9799), 
        .Y(n2271) );
  AO22X1_HVT U2244 ( .A1(\ram[8][163] ), .A2(n7388), .A3(n6058), .A4(n9802), 
        .Y(n2272) );
  AO22X1_HVT U2245 ( .A1(\ram[8][164] ), .A2(n7387), .A3(n6055), .A4(n9805), 
        .Y(n2273) );
  AO22X1_HVT U2246 ( .A1(\ram[8][165] ), .A2(n7367), .A3(n6054), .A4(n9808), 
        .Y(n2274) );
  AO22X1_HVT U2247 ( .A1(\ram[8][166] ), .A2(n7387), .A3(n6051), .A4(n9811), 
        .Y(n2275) );
  AO22X1_HVT U2248 ( .A1(\ram[8][167] ), .A2(n7367), .A3(n6070), .A4(n9814), 
        .Y(n2276) );
  AO22X1_HVT U2249 ( .A1(\ram[8][168] ), .A2(n7366), .A3(n6084), .A4(n9817), 
        .Y(n2277) );
  AO22X1_HVT U2250 ( .A1(\ram[8][169] ), .A2(n7365), .A3(n4356), .A4(n9820), 
        .Y(n2278) );
  AO22X1_HVT U2251 ( .A1(\ram[8][170] ), .A2(n7364), .A3(n6082), .A4(n9823), 
        .Y(n2279) );
  AO22X1_HVT U2252 ( .A1(\ram[8][171] ), .A2(n4349), .A3(n6079), .A4(n9826), 
        .Y(n2280) );
  AO22X1_HVT U2253 ( .A1(\ram[8][172] ), .A2(n10242), .A3(n6078), .A4(n9830), 
        .Y(n2281) );
  AO22X1_HVT U2254 ( .A1(\ram[8][173] ), .A2(n7357), .A3(n6059), .A4(n9833), 
        .Y(n2282) );
  AO22X1_HVT U2255 ( .A1(\ram[8][174] ), .A2(n7356), .A3(n6058), .A4(n9836), 
        .Y(n2283) );
  AO22X1_HVT U2256 ( .A1(\ram[8][175] ), .A2(n7417), .A3(n6055), .A4(n9839), 
        .Y(n2284) );
  AO22X1_HVT U2257 ( .A1(\ram[8][176] ), .A2(n4214), .A3(n6054), .A4(n9843), 
        .Y(n2285) );
  AO22X1_HVT U2258 ( .A1(\ram[8][177] ), .A2(n7415), .A3(n6051), .A4(n9846), 
        .Y(n2286) );
  AO22X1_HVT U2259 ( .A1(\ram[8][178] ), .A2(n7414), .A3(n6050), .A4(n9849), 
        .Y(n2287) );
  AO22X1_HVT U2260 ( .A1(\ram[8][179] ), .A2(n7361), .A3(n6049), .A4(n9852), 
        .Y(n2288) );
  AO22X1_HVT U2261 ( .A1(\ram[8][180] ), .A2(n7384), .A3(n6073), .A4(n9856), 
        .Y(n2289) );
  AO22X1_HVT U2262 ( .A1(\ram[8][181] ), .A2(n7383), .A3(n6095), .A4(n9859), 
        .Y(n2290) );
  AO22X1_HVT U2263 ( .A1(\ram[8][182] ), .A2(n4581), .A3(n6093), .A4(n9862), 
        .Y(n2291) );
  AO22X1_HVT U2264 ( .A1(\ram[8][183] ), .A2(n4377), .A3(n6096), .A4(n9865), 
        .Y(n2292) );
  AO22X1_HVT U2265 ( .A1(\ram[8][184] ), .A2(n4377), .A3(n6095), .A4(n9869), 
        .Y(n2293) );
  AO22X1_HVT U2266 ( .A1(\ram[8][185] ), .A2(n7379), .A3(n6093), .A4(n9872), 
        .Y(n2294) );
  AO22X1_HVT U2267 ( .A1(\ram[8][186] ), .A2(n7413), .A3(n6092), .A4(n9875), 
        .Y(n2295) );
  AO22X1_HVT U2268 ( .A1(\ram[8][187] ), .A2(n7377), .A3(n6090), .A4(n9878), 
        .Y(n2296) );
  AO22X1_HVT U2269 ( .A1(\ram[8][188] ), .A2(n7414), .A3(n6089), .A4(n9881), 
        .Y(n2297) );
  AO22X1_HVT U2270 ( .A1(\ram[8][189] ), .A2(n4349), .A3(n6088), .A4(n9884), 
        .Y(n2298) );
  AO22X1_HVT U2271 ( .A1(\ram[8][190] ), .A2(n7384), .A3(n6087), .A4(n9887), 
        .Y(n2299) );
  AO22X1_HVT U2272 ( .A1(\ram[8][191] ), .A2(n7383), .A3(n6085), .A4(n9890), 
        .Y(n2300) );
  AO22X1_HVT U2273 ( .A1(\ram[8][192] ), .A2(n7361), .A3(n6039), .A4(n9894), 
        .Y(n2301) );
  AO22X1_HVT U2274 ( .A1(\ram[8][193] ), .A2(n7380), .A3(n6111), .A4(n9897), 
        .Y(n2302) );
  AO22X1_HVT U2275 ( .A1(\ram[8][194] ), .A2(n7380), .A3(n6067), .A4(n9900), 
        .Y(n2303) );
  AO22X1_HVT U2276 ( .A1(\ram[8][195] ), .A2(n4377), .A3(n6068), .A4(n9903), 
        .Y(n2304) );
  AO22X1_HVT U2277 ( .A1(\ram[8][196] ), .A2(n10248), .A3(n6065), .A4(n9907), 
        .Y(n2305) );
  AO22X1_HVT U2278 ( .A1(\ram[8][197] ), .A2(n7412), .A3(n6070), .A4(n9910), 
        .Y(n2306) );
  AO22X1_HVT U2279 ( .A1(\ram[8][198] ), .A2(n7409), .A3(n6071), .A4(n9913), 
        .Y(n2307) );
  AO22X1_HVT U2280 ( .A1(\ram[8][199] ), .A2(n7409), .A3(n6072), .A4(n9916), 
        .Y(n2308) );
  AO22X1_HVT U2281 ( .A1(\ram[8][200] ), .A2(n7354), .A3(n6073), .A4(n9920), 
        .Y(n2309) );
  AO22X1_HVT U2282 ( .A1(\ram[8][201] ), .A2(n7375), .A3(n6074), .A4(n9923), 
        .Y(n2310) );
  AO22X1_HVT U2283 ( .A1(\ram[8][202] ), .A2(n10247), .A3(n6066), .A4(n9926), 
        .Y(n2311) );
  AO22X1_HVT U2284 ( .A1(\ram[8][203] ), .A2(n7365), .A3(n6075), .A4(n9929), 
        .Y(n2312) );
  AO22X1_HVT U2285 ( .A1(\ram[8][204] ), .A2(n7364), .A3(n6074), .A4(n9932), 
        .Y(n2313) );
  AO22X1_HVT U2286 ( .A1(\ram[8][205] ), .A2(n7366), .A3(n6059), .A4(n9935), 
        .Y(n2314) );
  AO22X1_HVT U2287 ( .A1(\ram[8][206] ), .A2(n7365), .A3(n6073), .A4(n9938), 
        .Y(n2315) );
  AO22X1_HVT U2288 ( .A1(\ram[8][207] ), .A2(n7364), .A3(n6092), .A4(n9941), 
        .Y(n2316) );
  AO22X1_HVT U2289 ( .A1(\ram[8][208] ), .A2(n10242), .A3(n6078), .A4(n9945), 
        .Y(n2317) );
  AO22X1_HVT U2290 ( .A1(\ram[8][209] ), .A2(n10242), .A3(n6112), .A4(n9948), 
        .Y(n2318) );
  AO22X1_HVT U2291 ( .A1(\ram[8][210] ), .A2(n7357), .A3(n6078), .A4(n9951), 
        .Y(n2319) );
  AO22X1_HVT U2292 ( .A1(\ram[8][211] ), .A2(n7356), .A3(n6108), .A4(n9954), 
        .Y(n2320) );
  AO22X1_HVT U2293 ( .A1(\ram[8][212] ), .A2(n7417), .A3(n6093), .A4(n9957), 
        .Y(n2321) );
  AO22X1_HVT U2294 ( .A1(\ram[8][213] ), .A2(n4606), .A3(n6079), .A4(n9960), 
        .Y(n2322) );
  AO22X1_HVT U2295 ( .A1(\ram[8][214] ), .A2(n7415), .A3(n6075), .A4(n9963), 
        .Y(n2323) );
  AO22X1_HVT U2296 ( .A1(\ram[8][215] ), .A2(n7414), .A3(n6040), .A4(n9966), 
        .Y(n2324) );
  AO22X1_HVT U2297 ( .A1(\ram[8][216] ), .A2(n10237), .A3(n6089), .A4(n9969), 
        .Y(n2325) );
  AO22X1_HVT U2298 ( .A1(\ram[8][217] ), .A2(n7374), .A3(n6055), .A4(n9972), 
        .Y(n2326) );
  AO22X1_HVT U2299 ( .A1(\ram[8][218] ), .A2(n4311), .A3(n6072), .A4(n9975), 
        .Y(n2327) );
  AO22X1_HVT U2300 ( .A1(\ram[8][219] ), .A2(n4581), .A3(n6082), .A4(n9978), 
        .Y(n2328) );
  AO22X1_HVT U2301 ( .A1(\ram[8][220] ), .A2(n7371), .A3(n6101), .A4(n9982), 
        .Y(n2329) );
  AO22X1_HVT U2302 ( .A1(\ram[8][221] ), .A2(n7370), .A3(n6090), .A4(n9985), 
        .Y(n2330) );
  AO22X1_HVT U2303 ( .A1(\ram[8][222] ), .A2(n7369), .A3(n6058), .A4(n9988), 
        .Y(n2331) );
  AO22X1_HVT U2304 ( .A1(\ram[8][223] ), .A2(n10248), .A3(n6073), .A4(n9991), 
        .Y(n2332) );
  AO22X1_HVT U2305 ( .A1(\ram[8][224] ), .A2(n7378), .A3(n6079), .A4(n9994), 
        .Y(n2333) );
  AO22X1_HVT U2306 ( .A1(\ram[8][225] ), .A2(n7411), .A3(n6092), .A4(n9997), 
        .Y(n2334) );
  AO22X1_HVT U2307 ( .A1(\ram[8][226] ), .A2(n7411), .A3(n6061), .A4(n10000), 
        .Y(n2335) );
  AO22X1_HVT U2308 ( .A1(\ram[8][227] ), .A2(n7412), .A3(n6059), .A4(n10003), 
        .Y(n2336) );
  AO22X1_HVT U2309 ( .A1(\ram[8][228] ), .A2(n7408), .A3(n6048), .A4(n10006), 
        .Y(n2337) );
  AO22X1_HVT U2310 ( .A1(\ram[8][229] ), .A2(n7406), .A3(n6084), .A4(n10009), 
        .Y(n2338) );
  AO22X1_HVT U2311 ( .A1(\ram[8][230] ), .A2(n4647), .A3(n6088), .A4(n10012), 
        .Y(n2339) );
  AO22X1_HVT U2312 ( .A1(\ram[8][231] ), .A2(n7402), .A3(n4356), .A4(n10015), 
        .Y(n2340) );
  AO22X1_HVT U2313 ( .A1(\ram[8][232] ), .A2(n7401), .A3(n6070), .A4(n10019), 
        .Y(n2341) );
  AO22X1_HVT U2314 ( .A1(\ram[8][233] ), .A2(n7400), .A3(n6101), .A4(n10022), 
        .Y(n2342) );
  AO22X1_HVT U2315 ( .A1(\ram[8][234] ), .A2(n7399), .A3(n6089), .A4(n10025), 
        .Y(n2343) );
  AO22X1_HVT U2316 ( .A1(\ram[8][235] ), .A2(n7398), .A3(n6084), .A4(n10028), 
        .Y(n2344) );
  AO22X1_HVT U2317 ( .A1(\ram[8][236] ), .A2(n4361), .A3(n6082), .A4(n10031), 
        .Y(n2345) );
  AO22X1_HVT U2318 ( .A1(\ram[8][237] ), .A2(n7397), .A3(n6071), .A4(n10034), 
        .Y(n2346) );
  AO22X1_HVT U2319 ( .A1(\ram[8][238] ), .A2(n4581), .A3(n6087), .A4(n10037), 
        .Y(n2347) );
  AO22X1_HVT U2320 ( .A1(\ram[8][239] ), .A2(n7378), .A3(n6090), .A4(n10040), 
        .Y(n2348) );
  AO22X1_HVT U2321 ( .A1(\ram[8][240] ), .A2(n7377), .A3(n6050), .A4(n10044), 
        .Y(n2349) );
  AO22X1_HVT U2322 ( .A1(\ram[8][241] ), .A2(n7375), .A3(n6045), .A4(n10047), 
        .Y(n2350) );
  AO22X1_HVT U2323 ( .A1(\ram[8][242] ), .A2(n7360), .A3(n6040), .A4(n10050), 
        .Y(n2351) );
  AO22X1_HVT U2324 ( .A1(\ram[8][243] ), .A2(n7374), .A3(n6088), .A4(n10053), 
        .Y(n2352) );
  AO22X1_HVT U2325 ( .A1(\ram[8][244] ), .A2(n7373), .A3(n6096), .A4(n10056), 
        .Y(n2353) );
  AO22X1_HVT U2326 ( .A1(\ram[8][245] ), .A2(n7372), .A3(n6051), .A4(n10059), 
        .Y(n2354) );
  AO22X1_HVT U2327 ( .A1(\ram[8][246] ), .A2(n7371), .A3(n6067), .A4(n10062), 
        .Y(n2355) );
  AO22X1_HVT U2328 ( .A1(\ram[8][247] ), .A2(n7408), .A3(n6042), .A4(n10065), 
        .Y(n2356) );
  AO22X1_HVT U2329 ( .A1(\ram[8][248] ), .A2(n7406), .A3(n6083), .A4(n10069), 
        .Y(n2357) );
  AO22X1_HVT U2330 ( .A1(\ram[8][249] ), .A2(n7405), .A3(n6095), .A4(n10072), 
        .Y(n2358) );
  AO22X1_HVT U2331 ( .A1(\ram[8][250] ), .A2(n7402), .A3(n6054), .A4(n10075), 
        .Y(n2359) );
  AO22X1_HVT U2332 ( .A1(\ram[8][251] ), .A2(n7380), .A3(n6068), .A4(n10078), 
        .Y(n2360) );
  AO22X1_HVT U2333 ( .A1(\ram[8][252] ), .A2(n10242), .A3(n6049), .A4(n10082), 
        .Y(n2361) );
  AO22X1_HVT U2334 ( .A1(\ram[8][253] ), .A2(n7370), .A3(n6041), .A4(n10085), 
        .Y(n2362) );
  AO22X1_HVT U2335 ( .A1(\ram[8][254] ), .A2(n7369), .A3(n6087), .A4(n10088), 
        .Y(n2363) );
  AO22X1_HVT U2336 ( .A1(\ram[8][255] ), .A2(n4580), .A3(n6087), .A4(n10091), 
        .Y(n2364) );
  AND2X1_HVT U2339 ( .A1(n38), .A2(n5130), .Y(n37) );
  AO22X1_HVT U2340 ( .A1(\ram[9][0] ), .A2(n10217), .A3(n9124), .A4(data[0]), 
        .Y(n2365) );
  AO22X1_HVT U2341 ( .A1(\ram[9][1] ), .A2(n7641), .A3(n9118), .A4(n9310), .Y(
        n2366) );
  AO22X1_HVT U2342 ( .A1(\ram[9][2] ), .A2(n4682), .A3(n9117), .A4(n9313), .Y(
        n2367) );
  AO22X1_HVT U2343 ( .A1(\ram[9][3] ), .A2(n7588), .A3(n9116), .A4(n9317), .Y(
        n2368) );
  AO22X1_HVT U2344 ( .A1(\ram[9][4] ), .A2(n7611), .A3(n9115), .A4(data[4]), 
        .Y(n2369) );
  AO22X1_HVT U2345 ( .A1(\ram[9][5] ), .A2(n7634), .A3(n9114), .A4(data[5]), 
        .Y(n2370) );
  AO22X1_HVT U2346 ( .A1(\ram[9][6] ), .A2(n7643), .A3(n9113), .A4(data[6]), 
        .Y(n2371) );
  AO22X1_HVT U2347 ( .A1(\ram[9][7] ), .A2(n7642), .A3(n9112), .A4(data[7]), 
        .Y(n2372) );
  AO22X1_HVT U2348 ( .A1(\ram[9][8] ), .A2(n7604), .A3(n9102), .A4(n9332), .Y(
        n2373) );
  AO22X1_HVT U2349 ( .A1(\ram[9][9] ), .A2(n7619), .A3(n9096), .A4(data[9]), 
        .Y(n2374) );
  AO22X1_HVT U2351 ( .A1(\ram[9][11] ), .A2(n4474), .A3(n9094), .A4(n9342), 
        .Y(n2376) );
  AO22X1_HVT U2352 ( .A1(\ram[9][12] ), .A2(n7618), .A3(n4800), .A4(data[12]), 
        .Y(n2377) );
  AO22X1_HVT U2353 ( .A1(\ram[9][13] ), .A2(n7643), .A3(n4801), .A4(data[13]), 
        .Y(n2378) );
  AO22X1_HVT U2354 ( .A1(\ram[9][14] ), .A2(n7617), .A3(n9089), .A4(n9351), 
        .Y(n2379) );
  AO22X1_HVT U2355 ( .A1(\ram[9][15] ), .A2(n7615), .A3(n4736), .A4(data[15]), 
        .Y(n2380) );
  AO22X1_HVT U2356 ( .A1(\ram[9][16] ), .A2(n7614), .A3(n9132), .A4(n9356), 
        .Y(n2381) );
  AO22X1_HVT U2357 ( .A1(\ram[9][17] ), .A2(n7609), .A3(n9118), .A4(n9360), 
        .Y(n2382) );
  AO22X1_HVT U2358 ( .A1(\ram[9][18] ), .A2(n7606), .A3(n9117), .A4(data[18]), 
        .Y(n2383) );
  AO22X1_HVT U2359 ( .A1(\ram[9][19] ), .A2(n4585), .A3(n9116), .A4(n9366), 
        .Y(n2384) );
  AO22X1_HVT U2360 ( .A1(\ram[9][20] ), .A2(n7604), .A3(n4724), .A4(n9368), 
        .Y(n2385) );
  AO22X1_HVT U2361 ( .A1(\ram[9][21] ), .A2(n7662), .A3(n9118), .A4(data[21]), 
        .Y(n2386) );
  AO22X1_HVT U2362 ( .A1(\ram[9][22] ), .A2(n7661), .A3(n9117), .A4(n9374), 
        .Y(n2387) );
  AO22X1_HVT U2363 ( .A1(\ram[9][23] ), .A2(n7660), .A3(n9116), .A4(n9377), 
        .Y(n2388) );
  AO22X1_HVT U2365 ( .A1(\ram[9][25] ), .A2(n7657), .A3(n9125), .A4(n9383), 
        .Y(n2390) );
  AO22X1_HVT U2367 ( .A1(\ram[9][27] ), .A2(n7654), .A3(n4724), .A4(n9389), 
        .Y(n2392) );
  AO22X1_HVT U2368 ( .A1(\ram[9][28] ), .A2(n7653), .A3(n9124), .A4(n9392), 
        .Y(n2393) );
  AO22X1_HVT U2371 ( .A1(\ram[9][31] ), .A2(n7642), .A3(n4658), .A4(data[31]), 
        .Y(n2396) );
  AO22X1_HVT U2372 ( .A1(\ram[9][32] ), .A2(n7638), .A3(n9122), .A4(data[32]), 
        .Y(n2397) );
  AO22X1_HVT U2373 ( .A1(\ram[9][33] ), .A2(n7637), .A3(n4656), .A4(data[33]), 
        .Y(n2398) );
  AO22X1_HVT U2374 ( .A1(\ram[9][34] ), .A2(n7590), .A3(n4656), .A4(n9410), 
        .Y(n2399) );
  AO22X1_HVT U2375 ( .A1(\ram[9][35] ), .A2(n7606), .A3(n4445), .A4(data[35]), 
        .Y(n2400) );
  AO22X1_HVT U2378 ( .A1(\ram[9][38] ), .A2(n7639), .A3(n9107), .A4(n9422), 
        .Y(n2403) );
  AO22X1_HVT U2380 ( .A1(\ram[9][40] ), .A2(n7599), .A3(n4335), .A4(data[40]), 
        .Y(n2405) );
  AO22X1_HVT U2381 ( .A1(\ram[9][41] ), .A2(n10211), .A3(n9105), .A4(data[41]), 
        .Y(n2406) );
  AO22X1_HVT U2382 ( .A1(\ram[9][42] ), .A2(n4585), .A3(n9095), .A4(data[42]), 
        .Y(n2407) );
  AO22X1_HVT U2383 ( .A1(\ram[9][43] ), .A2(n7597), .A3(n4380), .A4(n9437), 
        .Y(n2408) );
  AO22X1_HVT U2384 ( .A1(\ram[9][44] ), .A2(n7596), .A3(n9087), .A4(n9440), 
        .Y(n2409) );
  AO22X1_HVT U2389 ( .A1(\ram[9][49] ), .A2(n7605), .A3(n9086), .A4(n9454), 
        .Y(n2414) );
  AO22X1_HVT U2390 ( .A1(\ram[9][50] ), .A2(n7643), .A3(n9085), .A4(n9457), 
        .Y(n2415) );
  AO22X1_HVT U2391 ( .A1(\ram[9][51] ), .A2(n7642), .A3(n9084), .A4(data[51]), 
        .Y(n2416) );
  AO22X1_HVT U2392 ( .A1(\ram[9][52] ), .A2(n7634), .A3(n9103), .A4(n9464), 
        .Y(n2417) );
  AO22X1_HVT U2393 ( .A1(\ram[9][53] ), .A2(n7604), .A3(n4432), .A4(data[53]), 
        .Y(n2418) );
  AO22X1_HVT U2394 ( .A1(\ram[9][54] ), .A2(n7662), .A3(n9101), .A4(data[54]), 
        .Y(n2419) );
  AO22X1_HVT U2396 ( .A1(\ram[9][56] ), .A2(n7660), .A3(n4665), .A4(n9476), 
        .Y(n2421) );
  AO22X1_HVT U2397 ( .A1(\ram[9][57] ), .A2(n7658), .A3(n4726), .A4(data[57]), 
        .Y(n2422) );
  AO22X1_HVT U2398 ( .A1(\ram[9][58] ), .A2(n7657), .A3(n9134), .A4(data[58]), 
        .Y(n2423) );
  AO22X1_HVT U2399 ( .A1(\ram[9][59] ), .A2(n7656), .A3(n4445), .A4(data[59]), 
        .Y(n2424) );
  AO22X1_HVT U2400 ( .A1(\ram[9][60] ), .A2(n7654), .A3(n9103), .A4(n9488), 
        .Y(n2425) );
  AO22X1_HVT U2401 ( .A1(\ram[9][61] ), .A2(n7653), .A3(n4432), .A4(n9491), 
        .Y(n2426) );
  AO22X1_HVT U2403 ( .A1(\ram[9][63] ), .A2(n7650), .A3(n9100), .A4(data[63]), 
        .Y(n2428) );
  AO22X1_HVT U2404 ( .A1(\ram[9][64] ), .A2(n7649), .A3(n4308), .A4(n9500), 
        .Y(n2429) );
  AO22X1_HVT U2405 ( .A1(\ram[9][65] ), .A2(n7648), .A3(n9090), .A4(n9503), 
        .Y(n2430) );
  AO22X1_HVT U2406 ( .A1(\ram[9][66] ), .A2(n7646), .A3(n9089), .A4(n9506), 
        .Y(n2431) );
  AO22X1_HVT U2407 ( .A1(\ram[9][67] ), .A2(n7645), .A3(n9095), .A4(n9509), 
        .Y(n2432) );
  AO22X1_HVT U2408 ( .A1(\ram[9][68] ), .A2(n7588), .A3(n9115), .A4(n9512), 
        .Y(n2433) );
  AO22X1_HVT U2409 ( .A1(\ram[9][69] ), .A2(n7641), .A3(n9114), .A4(data[69]), 
        .Y(n2434) );
  AO22X1_HVT U2410 ( .A1(\ram[9][70] ), .A2(n7615), .A3(n9113), .A4(data[70]), 
        .Y(n2435) );
  AO22X1_HVT U2411 ( .A1(\ram[9][71] ), .A2(n7619), .A3(n9112), .A4(data[71]), 
        .Y(n2436) );
  AO22X1_HVT U2412 ( .A1(\ram[9][72] ), .A2(n7619), .A3(n9087), .A4(data[72]), 
        .Y(n2437) );
  AO22X1_HVT U2413 ( .A1(\ram[9][73] ), .A2(n7661), .A3(n9086), .A4(n9527), 
        .Y(n2438) );
  AO22X1_HVT U2414 ( .A1(\ram[9][74] ), .A2(n7618), .A3(n9085), .A4(n9530), 
        .Y(n2439) );
  AO22X1_HVT U2415 ( .A1(\ram[9][75] ), .A2(n7617), .A3(n9084), .A4(n9533), 
        .Y(n2440) );
  AO22X1_HVT U2416 ( .A1(\ram[9][76] ), .A2(n7617), .A3(n9115), .A4(data[76]), 
        .Y(n2441) );
  AO22X1_HVT U2417 ( .A1(\ram[9][77] ), .A2(n7615), .A3(n9114), .A4(n9539), 
        .Y(n2442) );
  AO22X1_HVT U2418 ( .A1(\ram[9][78] ), .A2(n7654), .A3(n9113), .A4(n9542), 
        .Y(n2443) );
  AO22X1_HVT U2419 ( .A1(\ram[9][79] ), .A2(n10212), .A3(n9112), .A4(n9545), 
        .Y(n2444) );
  AO22X1_HVT U2420 ( .A1(\ram[9][80] ), .A2(n7614), .A3(n9123), .A4(n9548), 
        .Y(n2445) );
  AO22X1_HVT U2421 ( .A1(\ram[9][81] ), .A2(n7613), .A3(n4503), .A4(n9551), 
        .Y(n2446) );
  AO22X1_HVT U2423 ( .A1(\ram[9][83] ), .A2(n7611), .A3(n4308), .A4(data[83]), 
        .Y(n2448) );
  AO22X1_HVT U2424 ( .A1(\ram[9][84] ), .A2(n7610), .A3(n9091), .A4(n9560), 
        .Y(n2449) );
  AO22X1_HVT U2425 ( .A1(\ram[9][85] ), .A2(n7656), .A3(n4335), .A4(n9563), 
        .Y(n2450) );
  AO22X1_HVT U2426 ( .A1(\ram[9][86] ), .A2(n7632), .A3(n4799), .A4(n9566), 
        .Y(n2451) );
  AO22X1_HVT U2427 ( .A1(\ram[9][87] ), .A2(n7631), .A3(n9094), .A4(data[87]), 
        .Y(n2452) );
  AO22X1_HVT U2428 ( .A1(\ram[9][88] ), .A2(n7630), .A3(n4652), .A4(n9571), 
        .Y(n2453) );
  AO22X1_HVT U2429 ( .A1(\ram[9][89] ), .A2(n7627), .A3(n9118), .A4(n9575), 
        .Y(n2454) );
  AO22X1_HVT U2430 ( .A1(\ram[9][90] ), .A2(n7626), .A3(n9117), .A4(data[90]), 
        .Y(n2455) );
  AO22X1_HVT U2431 ( .A1(\ram[9][91] ), .A2(n7625), .A3(n9116), .A4(data[91]), 
        .Y(n2456) );
  AO22X1_HVT U2432 ( .A1(\ram[9][92] ), .A2(n7624), .A3(n9115), .A4(n9584), 
        .Y(n2457) );
  AO22X1_HVT U2433 ( .A1(\ram[9][93] ), .A2(n7623), .A3(n9114), .A4(n9587), 
        .Y(n2458) );
  AO22X1_HVT U2434 ( .A1(\ram[9][94] ), .A2(n7622), .A3(n9113), .A4(n9590), 
        .Y(n2459) );
  AO22X1_HVT U2435 ( .A1(\ram[9][95] ), .A2(n7618), .A3(n9112), .A4(n9593), 
        .Y(n2460) );
  AO22X1_HVT U2436 ( .A1(\ram[9][96] ), .A2(n7601), .A3(n9087), .A4(n9596), 
        .Y(n2461) );
  AO22X1_HVT U2437 ( .A1(\ram[9][97] ), .A2(n7600), .A3(n9086), .A4(n9599), 
        .Y(n2462) );
  AO22X1_HVT U2438 ( .A1(\ram[9][98] ), .A2(n7599), .A3(n9085), .A4(n9602), 
        .Y(n2463) );
  AO22X1_HVT U2439 ( .A1(\ram[9][99] ), .A2(n4682), .A3(n9084), .A4(n9605), 
        .Y(n2464) );
  AO22X1_HVT U2440 ( .A1(\ram[9][100] ), .A2(n7588), .A3(n4726), .A4(n9608), 
        .Y(n2465) );
  AO22X1_HVT U2441 ( .A1(\ram[9][101] ), .A2(n7597), .A3(n9135), .A4(n9611), 
        .Y(n2466) );
  AO22X1_HVT U2442 ( .A1(\ram[9][102] ), .A2(n7596), .A3(n9135), .A4(n9614), 
        .Y(n2467) );
  AO22X1_HVT U2443 ( .A1(\ram[9][103] ), .A2(n7622), .A3(n9134), .A4(data[103]), .Y(n2468) );
  AO22X1_HVT U2444 ( .A1(\ram[9][104] ), .A2(n7652), .A3(n4663), .A4(n9620), 
        .Y(n2469) );
  AO22X1_HVT U2445 ( .A1(\ram[9][105] ), .A2(n7601), .A3(n4509), .A4(data[105]), .Y(n2470) );
  AO22X1_HVT U2446 ( .A1(\ram[9][106] ), .A2(n7600), .A3(n9133), .A4(n9626), 
        .Y(n2471) );
  AO22X1_HVT U2448 ( .A1(\ram[9][108] ), .A2(n4585), .A3(n9136), .A4(data[108]), .Y(n2473) );
  AO22X1_HVT U2449 ( .A1(\ram[9][109] ), .A2(n10216), .A3(n9118), .A4(n9635), 
        .Y(n2474) );
  AO22X1_HVT U2450 ( .A1(\ram[9][110] ), .A2(n7597), .A3(n9117), .A4(n9638), 
        .Y(n2475) );
  AO22X1_HVT U2451 ( .A1(\ram[9][111] ), .A2(n7596), .A3(n9116), .A4(n9641), 
        .Y(n2476) );
  AO22X1_HVT U2452 ( .A1(\ram[9][112] ), .A2(n7595), .A3(n4308), .A4(n9644), 
        .Y(n2477) );
  AO22X1_HVT U2453 ( .A1(\ram[9][113] ), .A2(n7592), .A3(n4801), .A4(n9647), 
        .Y(n2478) );
  AO22X1_HVT U2454 ( .A1(\ram[9][114] ), .A2(n7591), .A3(n9101), .A4(n9650), 
        .Y(n2479) );
  AO22X1_HVT U2455 ( .A1(\ram[9][115] ), .A2(n7623), .A3(n9100), .A4(data[115]), .Y(n2480) );
  AO22X1_HVT U2456 ( .A1(\ram[9][116] ), .A2(n7622), .A3(n4665), .A4(n9656), 
        .Y(n2481) );
  AO22X1_HVT U2457 ( .A1(\ram[9][117] ), .A2(n10214), .A3(n9129), .A4(
        data[117]), .Y(n2482) );
  AO22X1_HVT U2458 ( .A1(\ram[9][118] ), .A2(n7601), .A3(n9133), .A4(data[118]), .Y(n2483) );
  AO22X1_HVT U2459 ( .A1(\ram[9][119] ), .A2(n7600), .A3(n4726), .A4(n9665), 
        .Y(n2484) );
  AO22X1_HVT U2460 ( .A1(\ram[9][120] ), .A2(n7590), .A3(n9123), .A4(data[120]), .Y(n2485) );
  AO22X1_HVT U2461 ( .A1(\ram[9][121] ), .A2(n10209), .A3(n9121), .A4(
        data[121]), .Y(n2486) );
  AO22X1_HVT U2462 ( .A1(\ram[9][122] ), .A2(n7657), .A3(n9122), .A4(data[122]), .Y(n2487) );
  AO22X1_HVT U2463 ( .A1(\ram[9][123] ), .A2(n10217), .A3(n9123), .A4(n9677), 
        .Y(n2488) );
  AO22X1_HVT U2464 ( .A1(\ram[9][124] ), .A2(n10209), .A3(n4684), .A4(n9680), 
        .Y(n2489) );
  AO22X1_HVT U2465 ( .A1(\ram[9][125] ), .A2(n7587), .A3(n9096), .A4(n9683), 
        .Y(n2490) );
  AO22X1_HVT U2467 ( .A1(\ram[9][127] ), .A2(n7606), .A3(n4736), .A4(n9689), 
        .Y(n2492) );
  AO22X1_HVT U2468 ( .A1(\ram[9][128] ), .A2(n7605), .A3(n4464), .A4(data[128]), .Y(n2493) );
  AO22X1_HVT U2469 ( .A1(\ram[9][129] ), .A2(n7643), .A3(n9133), .A4(n9695), 
        .Y(n2494) );
  AO22X1_HVT U2470 ( .A1(\ram[9][130] ), .A2(n7638), .A3(n9130), .A4(n9698), 
        .Y(n2495) );
  AO22X1_HVT U2471 ( .A1(\ram[9][131] ), .A2(n7637), .A3(n4464), .A4(data[131]), .Y(n2496) );
  AO22X1_HVT U2472 ( .A1(\ram[9][132] ), .A2(n7636), .A3(n4684), .A4(n9704), 
        .Y(n2497) );
  AO22X1_HVT U2473 ( .A1(\ram[9][133] ), .A2(n7635), .A3(n9096), .A4(n9707), 
        .Y(n2498) );
  AO22X1_HVT U2474 ( .A1(\ram[9][134] ), .A2(n7634), .A3(n9088), .A4(n9710), 
        .Y(n2499) );
  AO22X1_HVT U2475 ( .A1(\ram[9][135] ), .A2(n7632), .A3(n9088), .A4(data[135]), .Y(n2500) );
  AO22X1_HVT U2476 ( .A1(\ram[9][136] ), .A2(n7631), .A3(n9103), .A4(data[136]), .Y(n2501) );
  AO22X1_HVT U2477 ( .A1(\ram[9][137] ), .A2(n7630), .A3(n4801), .A4(n9719), 
        .Y(n2502) );
  AO22X1_HVT U2478 ( .A1(\ram[9][138] ), .A2(n7627), .A3(n4799), .A4(data[138]), .Y(n2503) );
  AO22X1_HVT U2479 ( .A1(\ram[9][139] ), .A2(n7626), .A3(n4380), .A4(n9726), 
        .Y(n2504) );
  AO22X1_HVT U2480 ( .A1(\ram[9][140] ), .A2(n7625), .A3(n9134), .A4(n9729), 
        .Y(n2505) );
  AO22X1_HVT U2481 ( .A1(\ram[9][141] ), .A2(n7624), .A3(n9118), .A4(n9732), 
        .Y(n2506) );
  AO22X1_HVT U2482 ( .A1(\ram[9][142] ), .A2(n7623), .A3(n9117), .A4(n9735), 
        .Y(n2507) );
  AO22X1_HVT U2483 ( .A1(\ram[9][143] ), .A2(n7622), .A3(n9116), .A4(n9739), 
        .Y(n2508) );
  AO22X1_HVT U2484 ( .A1(\ram[9][144] ), .A2(n7610), .A3(n9115), .A4(n9742), 
        .Y(n2509) );
  AO22X1_HVT U2485 ( .A1(\ram[9][145] ), .A2(n7590), .A3(n9114), .A4(data[145]), .Y(n2510) );
  AO22X1_HVT U2486 ( .A1(\ram[9][146] ), .A2(n10212), .A3(n9113), .A4(n9748), 
        .Y(n2511) );
  AO22X1_HVT U2487 ( .A1(\ram[9][147] ), .A2(n7614), .A3(n9112), .A4(n9752), 
        .Y(n2512) );
  AO22X1_HVT U2488 ( .A1(\ram[9][148] ), .A2(n7613), .A3(n9090), .A4(n9755), 
        .Y(n2513) );
  AO22X1_HVT U2489 ( .A1(\ram[9][149] ), .A2(n7645), .A3(n9091), .A4(n9758), 
        .Y(n2514) );
  AO22X1_HVT U2490 ( .A1(\ram[9][150] ), .A2(n7611), .A3(n4736), .A4(data[150]), .Y(n2515) );
  AO22X1_HVT U2491 ( .A1(\ram[9][151] ), .A2(n7610), .A3(n9094), .A4(n9764), 
        .Y(n2516) );
  AO22X1_HVT U2492 ( .A1(\ram[9][152] ), .A2(n7609), .A3(n9103), .A4(n9767), 
        .Y(n2517) );
  AO22X1_HVT U2493 ( .A1(\ram[9][153] ), .A2(n7606), .A3(n9102), .A4(data[153]), .Y(n2518) );
  AO22X1_HVT U2494 ( .A1(\ram[9][154] ), .A2(n7605), .A3(n9089), .A4(n9773), 
        .Y(n2519) );
  AO22X1_HVT U2495 ( .A1(\ram[9][155] ), .A2(n7604), .A3(n4857), .A4(n9777), 
        .Y(n2520) );
  AO22X1_HVT U2496 ( .A1(\ram[9][156] ), .A2(n7662), .A3(n4358), .A4(data[156]), .Y(n2521) );
  AO22X1_HVT U2498 ( .A1(\ram[9][158] ), .A2(n7660), .A3(n4797), .A4(data[158]), .Y(n2523) );
  AO22X1_HVT U2499 ( .A1(\ram[9][159] ), .A2(n7658), .A3(n9106), .A4(n9790), 
        .Y(n2524) );
  AO22X1_HVT U2500 ( .A1(\ram[9][160] ), .A2(n7657), .A3(n4503), .A4(data[160]), .Y(n2525) );
  AO22X1_HVT U2501 ( .A1(\ram[9][161] ), .A2(n7656), .A3(n9108), .A4(data[161]), .Y(n2526) );
  AO22X1_HVT U2502 ( .A1(\ram[9][162] ), .A2(n7654), .A3(n4797), .A4(n9799), 
        .Y(n2527) );
  AO22X1_HVT U2503 ( .A1(\ram[9][163] ), .A2(n7652), .A3(n9106), .A4(n9802), 
        .Y(n2528) );
  AO22X1_HVT U2504 ( .A1(\ram[9][164] ), .A2(n7650), .A3(n4801), .A4(data[164]), .Y(n2529) );
  AO22X1_HVT U2505 ( .A1(\ram[9][165] ), .A2(n7649), .A3(n4800), .A4(data[165]), .Y(n2530) );
  AO22X1_HVT U2506 ( .A1(\ram[9][166] ), .A2(n7648), .A3(n4857), .A4(data[166]), .Y(n2531) );
  AO22X1_HVT U2507 ( .A1(\ram[9][167] ), .A2(n7646), .A3(n4857), .A4(data[167]), .Y(n2532) );
  AO22X1_HVT U2508 ( .A1(\ram[9][168] ), .A2(n7645), .A3(n4800), .A4(n9817), 
        .Y(n2533) );
  AO22X1_HVT U2509 ( .A1(\ram[9][169] ), .A2(n7613), .A3(n4684), .A4(n9820), 
        .Y(n2534) );
  AO22X1_HVT U2510 ( .A1(\ram[9][170] ), .A2(n7641), .A3(n4799), .A4(data[170]), .Y(n2535) );
  AO22X1_HVT U2512 ( .A1(\ram[9][172] ), .A2(n7639), .A3(n9129), .A4(data[172]), .Y(n2537) );
  AO22X1_HVT U2513 ( .A1(\ram[9][173] ), .A2(n7650), .A3(n9129), .A4(data[173]), .Y(n2538) );
  AO22X1_HVT U2514 ( .A1(\ram[9][174] ), .A2(n7638), .A3(n9131), .A4(data[174]), .Y(n2539) );
  AO22X1_HVT U2515 ( .A1(\ram[9][175] ), .A2(n7636), .A3(n9131), .A4(n9840), 
        .Y(n2540) );
  AO22X1_HVT U2516 ( .A1(\ram[9][176] ), .A2(n7635), .A3(n9087), .A4(data[176]), .Y(n2541) );
  AO22X1_HVT U2517 ( .A1(\ram[9][177] ), .A2(n7587), .A3(n9086), .A4(data[177]), .Y(n2542) );
  AO22X1_HVT U2518 ( .A1(\ram[9][178] ), .A2(n7632), .A3(n9085), .A4(data[178]), .Y(n2543) );
  AO22X1_HVT U2519 ( .A1(\ram[9][179] ), .A2(n7631), .A3(n9084), .A4(n9853), 
        .Y(n2544) );
  AO22X1_HVT U2520 ( .A1(\ram[9][180] ), .A2(n7595), .A3(n9091), .A4(n9856), 
        .Y(n2545) );
  AO22X1_HVT U2521 ( .A1(\ram[9][181] ), .A2(n7592), .A3(n9097), .A4(data[181]), .Y(n2546) );
  AO22X1_HVT U2522 ( .A1(\ram[9][182] ), .A2(n7591), .A3(n9101), .A4(n9862), 
        .Y(n2547) );
  AO22X1_HVT U2523 ( .A1(\ram[9][183] ), .A2(n7601), .A3(n9100), .A4(n9866), 
        .Y(n2548) );
  AO22X1_HVT U2524 ( .A1(\ram[9][184] ), .A2(n7600), .A3(n4656), .A4(data[184]), .Y(n2549) );
  AO22X1_HVT U2525 ( .A1(\ram[9][185] ), .A2(n7599), .A3(n9135), .A4(n9872), 
        .Y(n2550) );
  AO22X1_HVT U2526 ( .A1(\ram[9][186] ), .A2(n7642), .A3(n9129), .A4(data[186]), .Y(n2551) );
  AO22X1_HVT U2527 ( .A1(\ram[9][187] ), .A2(n7587), .A3(n4466), .A4(data[187]), .Y(n2552) );
  AO22X1_HVT U2528 ( .A1(\ram[9][188] ), .A2(n7619), .A3(n4663), .A4(data[188]), .Y(n2553) );
  AO22X1_HVT U2529 ( .A1(\ram[9][189] ), .A2(n7609), .A3(n9130), .A4(n9884), 
        .Y(n2554) );
  AO22X1_HVT U2530 ( .A1(\ram[9][190] ), .A2(n7661), .A3(n9131), .A4(data[190]), .Y(n2555) );
  AO22X1_HVT U2531 ( .A1(\ram[9][191] ), .A2(n7618), .A3(n9131), .A4(n9891), 
        .Y(n2556) );
  AO22X1_HVT U2532 ( .A1(\ram[9][192] ), .A2(n10212), .A3(n4663), .A4(n9894), 
        .Y(n2557) );
  AO22X1_HVT U2533 ( .A1(\ram[9][193] ), .A2(n7614), .A3(n4725), .A4(n9897), 
        .Y(n2558) );
  AO22X1_HVT U2534 ( .A1(\ram[9][194] ), .A2(n7613), .A3(n4725), .A4(data[194]), .Y(n2559) );
  AO22X1_HVT U2535 ( .A1(\ram[9][195] ), .A2(n10216), .A3(n4358), .A4(n9904), 
        .Y(n2560) );
  AO22X1_HVT U2536 ( .A1(\ram[9][196] ), .A2(n7611), .A3(n4658), .A4(data[196]), .Y(n2561) );
  AO22X1_HVT U2537 ( .A1(\ram[9][197] ), .A2(n7610), .A3(n4658), .A4(data[197]), .Y(n2562) );
  AO22X1_HVT U2538 ( .A1(\ram[9][198] ), .A2(n7609), .A3(n9125), .A4(data[198]), .Y(n2563) );
  AO22X1_HVT U2539 ( .A1(\ram[9][199] ), .A2(n7606), .A3(n4725), .A4(n9917), 
        .Y(n2564) );
  AO22X1_HVT U2540 ( .A1(\ram[9][200] ), .A2(n10216), .A3(n9135), .A4(n9920), 
        .Y(n2565) );
  AO22X1_HVT U2541 ( .A1(\ram[9][201] ), .A2(n10211), .A3(n9135), .A4(
        data[201]), .Y(n2566) );
  AO22X1_HVT U2542 ( .A1(\ram[9][202] ), .A2(n7597), .A3(n4724), .A4(n9926), 
        .Y(n2567) );
  AO22X1_HVT U2543 ( .A1(\ram[9][203] ), .A2(n7596), .A3(n4726), .A4(data[203]), .Y(n2568) );
  AO22X1_HVT U2544 ( .A1(\ram[9][204] ), .A2(n7595), .A3(n4466), .A4(data[204]), .Y(n2569) );
  AO22X1_HVT U2545 ( .A1(\ram[9][205] ), .A2(n7592), .A3(n4665), .A4(data[205]), .Y(n2570) );
  AO22X1_HVT U2546 ( .A1(\ram[9][206] ), .A2(n7591), .A3(n4726), .A4(n9938), 
        .Y(n2571) );
  AO22X1_HVT U2547 ( .A1(\ram[9][207] ), .A2(n7590), .A3(n9130), .A4(n9942), 
        .Y(n2572) );
  AO22X1_HVT U2548 ( .A1(\ram[9][208] ), .A2(n7587), .A3(n9132), .A4(n9945), 
        .Y(n2573) );
  AO22X1_HVT U2549 ( .A1(\ram[9][209] ), .A2(n10212), .A3(n4509), .A4(
        data[209]), .Y(n2574) );
  AO22X1_HVT U2550 ( .A1(\ram[9][210] ), .A2(n10209), .A3(n4725), .A4(n9951), 
        .Y(n2575) );
  AO22X1_HVT U2551 ( .A1(\ram[9][211] ), .A2(n10209), .A3(n9130), .A4(n9954), 
        .Y(n2576) );
  AO22X1_HVT U2552 ( .A1(\ram[9][212] ), .A2(n4682), .A3(n9109), .A4(n9957), 
        .Y(n2577) );
  AO22X1_HVT U2553 ( .A1(\ram[9][213] ), .A2(n7588), .A3(n9108), .A4(data[213]), .Y(n2578) );
  AO22X1_HVT U2554 ( .A1(\ram[9][214] ), .A2(n7658), .A3(n4797), .A4(n9963), 
        .Y(n2579) );
  AO22X1_HVT U2555 ( .A1(\ram[9][215] ), .A2(n7660), .A3(n9106), .A4(data[215]), .Y(n2580) );
  AO22X1_HVT U2556 ( .A1(\ram[9][216] ), .A2(n7653), .A3(n4800), .A4(n9969), 
        .Y(n2581) );
  AO22X1_HVT U2557 ( .A1(\ram[9][217] ), .A2(n7652), .A3(n9097), .A4(n9972), 
        .Y(n2582) );
  AO22X1_HVT U2558 ( .A1(\ram[9][218] ), .A2(n7650), .A3(n9101), .A4(n9975), 
        .Y(n2583) );
  AO22X1_HVT U2559 ( .A1(\ram[9][219] ), .A2(n7649), .A3(n9100), .A4(n9979), 
        .Y(n2584) );
  AO22X1_HVT U2560 ( .A1(\ram[9][220] ), .A2(n7648), .A3(n9132), .A4(n9982), 
        .Y(n2585) );
  AO22X1_HVT U2561 ( .A1(\ram[9][221] ), .A2(n7646), .A3(n9131), .A4(data[221]), .Y(n2586) );
  AO22X1_HVT U2562 ( .A1(\ram[9][222] ), .A2(n7645), .A3(n9133), .A4(data[222]), .Y(n2587) );
  AO22X1_HVT U2563 ( .A1(\ram[9][223] ), .A2(n7648), .A3(n4725), .A4(data[223]), .Y(n2588) );
  AO22X1_HVT U2564 ( .A1(\ram[9][224] ), .A2(n7641), .A3(n9125), .A4(n9994), 
        .Y(n2589) );
  AO22X1_HVT U2567 ( .A1(\ram[9][227] ), .A2(n7649), .A3(n9125), .A4(n10003), 
        .Y(n2592) );
  AO22X1_HVT U2568 ( .A1(\ram[9][228] ), .A2(n7638), .A3(n4684), .A4(data[228]), .Y(n2593) );
  AO22X1_HVT U2569 ( .A1(\ram[9][229] ), .A2(n7637), .A3(n9121), .A4(n10009), 
        .Y(n2594) );
  AO22X1_HVT U2570 ( .A1(\ram[9][230] ), .A2(n7636), .A3(n9122), .A4(n10012), 
        .Y(n2595) );
  AO22X1_HVT U2571 ( .A1(\ram[9][231] ), .A2(n7635), .A3(n4233), .A4(n10016), 
        .Y(n2596) );
  AO22X1_HVT U2572 ( .A1(\ram[9][232] ), .A2(n4585), .A3(n9109), .A4(n10019), 
        .Y(n2597) );
  AO22X1_HVT U2573 ( .A1(\ram[9][233] ), .A2(n7637), .A3(n9108), .A4(data[233]), .Y(n2598) );
  AO22X1_HVT U2574 ( .A1(\ram[9][234] ), .A2(n7636), .A3(n9107), .A4(data[234]), .Y(n2599) );
  AO22X1_HVT U2575 ( .A1(\ram[9][235] ), .A2(n7635), .A3(n9106), .A4(n10028), 
        .Y(n2600) );
  AO22X1_HVT U2576 ( .A1(\ram[9][236] ), .A2(n7605), .A3(n9121), .A4(data[236]), .Y(n2601) );
  AO22X1_HVT U2577 ( .A1(\ram[9][237] ), .A2(n7632), .A3(n4652), .A4(data[237]), .Y(n2602) );
  AO22X1_HVT U2578 ( .A1(\ram[9][238] ), .A2(n7631), .A3(n9122), .A4(n10037), 
        .Y(n2603) );
  AO22X1_HVT U2579 ( .A1(\ram[9][239] ), .A2(n7630), .A3(n9121), .A4(n10041), 
        .Y(n2604) );
  AO22X1_HVT U2580 ( .A1(\ram[9][240] ), .A2(n7627), .A3(n4503), .A4(n10044), 
        .Y(n2605) );
  AO22X1_HVT U2581 ( .A1(\ram[9][241] ), .A2(n7626), .A3(n9108), .A4(n10047), 
        .Y(n2606) );
  AO22X1_HVT U2582 ( .A1(\ram[9][242] ), .A2(n7625), .A3(n9107), .A4(n10050), 
        .Y(n2607) );
  AO22X1_HVT U2583 ( .A1(\ram[9][243] ), .A2(n7624), .A3(n9106), .A4(n10053), 
        .Y(n2608) );
  AO22X1_HVT U2584 ( .A1(\ram[9][244] ), .A2(n7623), .A3(n9121), .A4(data[244]), .Y(n2609) );
  AO22X1_HVT U2585 ( .A1(\ram[9][245] ), .A2(n7630), .A3(n9122), .A4(data[245]), .Y(n2610) );
  AO22X1_HVT U2586 ( .A1(\ram[9][246] ), .A2(n7627), .A3(n4432), .A4(data[246]), .Y(n2611) );
  AO22X1_HVT U2587 ( .A1(\ram[9][247] ), .A2(n7626), .A3(n4503), .A4(n10066), 
        .Y(n2612) );
  AO22X1_HVT U2588 ( .A1(\ram[9][248] ), .A2(n7625), .A3(n4724), .A4(n10069), 
        .Y(n2613) );
  AO22X1_HVT U2589 ( .A1(\ram[9][249] ), .A2(n7624), .A3(n9124), .A4(data[249]), .Y(n2614) );
  AO22X1_HVT U2590 ( .A1(\ram[9][250] ), .A2(n7588), .A3(n4233), .A4(n10075), 
        .Y(n2615) );
  AO22X1_HVT U2591 ( .A1(\ram[9][251] ), .A2(n10217), .A3(n4233), .A4(n10079), 
        .Y(n2616) );
  AO22X1_HVT U2592 ( .A1(\ram[9][252] ), .A2(n7658), .A3(n9115), .A4(data[252]), .Y(n2617) );
  AO22X1_HVT U2593 ( .A1(\ram[9][253] ), .A2(n7617), .A3(n9114), .A4(data[253]), .Y(n2618) );
  AO22X1_HVT U2594 ( .A1(\ram[9][254] ), .A2(n7615), .A3(n9113), .A4(n10088), 
        .Y(n2619) );
  AO22X1_HVT U2595 ( .A1(\ram[9][255] ), .A2(n7653), .A3(n9112), .A4(n10092), 
        .Y(n2620) );
  AND2X1_HVT U2596 ( .A1(n41), .A2(n10375), .Y(n40) );
  AND2X1_HVT U2598 ( .A1(n5563), .A2(n38), .Y(n41) );
  AO22X1_HVT U2599 ( .A1(\ram[10][0] ), .A2(n7481), .A3(n6476), .A4(n9307), 
        .Y(n2621) );
  AO22X1_HVT U2600 ( .A1(\ram[10][1] ), .A2(n7522), .A3(n6474), .A4(n9310), 
        .Y(n2622) );
  AO22X1_HVT U2601 ( .A1(\ram[10][2] ), .A2(n7521), .A3(n6473), .A4(n9312), 
        .Y(n2623) );
  AO22X1_HVT U2602 ( .A1(\ram[10][3] ), .A2(n7519), .A3(n6449), .A4(n9316), 
        .Y(n2624) );
  AO22X1_HVT U2603 ( .A1(\ram[10][4] ), .A2(n7518), .A3(n6425), .A4(n9320), 
        .Y(n2625) );
  AO22X1_HVT U2604 ( .A1(\ram[10][5] ), .A2(n7515), .A3(n6479), .A4(n9323), 
        .Y(n2626) );
  AO22X1_HVT U2605 ( .A1(\ram[10][6] ), .A2(n7514), .A3(n6478), .A4(n9326), 
        .Y(n2627) );
  AO22X1_HVT U2606 ( .A1(\ram[10][7] ), .A2(n7512), .A3(n6477), .A4(n9329), 
        .Y(n2628) );
  AO22X1_HVT U2607 ( .A1(\ram[10][8] ), .A2(n7511), .A3(n6476), .A4(n9332), 
        .Y(n2629) );
  AO22X1_HVT U2608 ( .A1(\ram[10][9] ), .A2(n7509), .A3(n6474), .A4(n9335), 
        .Y(n2630) );
  AO22X1_HVT U2609 ( .A1(\ram[10][10] ), .A2(n7508), .A3(n6473), .A4(n9338), 
        .Y(n2631) );
  AO22X1_HVT U2610 ( .A1(\ram[10][11] ), .A2(n7506), .A3(n6472), .A4(n9341), 
        .Y(n2632) );
  AO22X1_HVT U2611 ( .A1(\ram[10][12] ), .A2(n7505), .A3(n6471), .A4(n9345), 
        .Y(n2633) );
  AO22X1_HVT U2612 ( .A1(\ram[10][13] ), .A2(n7503), .A3(n6466), .A4(n9348), 
        .Y(n2634) );
  AO22X1_HVT U2613 ( .A1(\ram[10][14] ), .A2(n7502), .A3(n6463), .A4(n9351), 
        .Y(n2635) );
  AO22X1_HVT U2614 ( .A1(\ram[10][15] ), .A2(n7500), .A3(n6462), .A4(n9354), 
        .Y(n2636) );
  AO22X1_HVT U2615 ( .A1(\ram[10][16] ), .A2(n7499), .A3(n6460), .A4(n9357), 
        .Y(n2637) );
  AO22X1_HVT U2616 ( .A1(\ram[10][17] ), .A2(n7498), .A3(n6477), .A4(n9360), 
        .Y(n2638) );
  AO22X1_HVT U2617 ( .A1(\ram[10][18] ), .A2(n7497), .A3(n6421), .A4(n9363), 
        .Y(n2639) );
  AO22X1_HVT U2618 ( .A1(\ram[10][19] ), .A2(n7494), .A3(n6420), .A4(n9366), 
        .Y(n2640) );
  AO22X1_HVT U2619 ( .A1(\ram[10][20] ), .A2(n7493), .A3(n6472), .A4(data[20]), 
        .Y(n2641) );
  AO22X1_HVT U2620 ( .A1(\ram[10][21] ), .A2(n7492), .A3(n6469), .A4(n9371), 
        .Y(n2642) );
  AO22X1_HVT U2621 ( .A1(\ram[10][22] ), .A2(n7491), .A3(n6468), .A4(n9374), 
        .Y(n2643) );
  AO22X1_HVT U2622 ( .A1(\ram[10][23] ), .A2(n7486), .A3(n6425), .A4(n9377), 
        .Y(n2644) );
  AO22X1_HVT U2623 ( .A1(\ram[10][24] ), .A2(n7485), .A3(n6467), .A4(n9380), 
        .Y(n2645) );
  AO22X1_HVT U2624 ( .A1(\ram[10][25] ), .A2(n7484), .A3(n6466), .A4(n9383), 
        .Y(n2646) );
  AO22X1_HVT U2625 ( .A1(\ram[10][26] ), .A2(n7483), .A3(n6463), .A4(n9386), 
        .Y(n2647) );
  AO22X1_HVT U2626 ( .A1(\ram[10][27] ), .A2(n7481), .A3(n6462), .A4(n9389), 
        .Y(n2648) );
  AO22X1_HVT U2627 ( .A1(\ram[10][28] ), .A2(n7480), .A3(n6460), .A4(n9392), 
        .Y(n2649) );
  AO22X1_HVT U2628 ( .A1(\ram[10][29] ), .A2(n7479), .A3(n6459), .A4(n9395), 
        .Y(n2650) );
  AO22X1_HVT U2629 ( .A1(\ram[10][30] ), .A2(n7478), .A3(n10185), .A4(data[30]), .Y(n2651) );
  AO22X1_HVT U2630 ( .A1(\ram[10][31] ), .A2(n7542), .A3(n6460), .A4(n9401), 
        .Y(n2652) );
  AO22X1_HVT U2631 ( .A1(\ram[10][32] ), .A2(n7541), .A3(n6459), .A4(n9404), 
        .Y(n2653) );
  AO22X1_HVT U2632 ( .A1(\ram[10][33] ), .A2(n7540), .A3(n10185), .A4(n9407), 
        .Y(n2654) );
  AO22X1_HVT U2633 ( .A1(\ram[10][34] ), .A2(n7539), .A3(n6457), .A4(n9410), 
        .Y(n2655) );
  AO22X1_HVT U2634 ( .A1(\ram[10][35] ), .A2(n7508), .A3(n6456), .A4(n9413), 
        .Y(n2656) );
  AO22X1_HVT U2635 ( .A1(\ram[10][36] ), .A2(n7506), .A3(n6455), .A4(n9416), 
        .Y(n2657) );
  AO22X1_HVT U2636 ( .A1(\ram[10][37] ), .A2(n7505), .A3(n6454), .A4(n9419), 
        .Y(n2658) );
  AO22X1_HVT U2637 ( .A1(\ram[10][38] ), .A2(n7503), .A3(n6453), .A4(n9422), 
        .Y(n2659) );
  AO22X1_HVT U2638 ( .A1(\ram[10][39] ), .A2(n7502), .A3(n4199), .A4(data[39]), 
        .Y(n2660) );
  AO22X1_HVT U2639 ( .A1(\ram[10][40] ), .A2(n7500), .A3(n6424), .A4(n9428), 
        .Y(n2661) );
  AO22X1_HVT U2640 ( .A1(\ram[10][41] ), .A2(n7499), .A3(n6452), .A4(n9431), 
        .Y(n2662) );
  AO22X1_HVT U2641 ( .A1(\ram[10][42] ), .A2(n7498), .A3(n10181), .A4(n9434), 
        .Y(n2663) );
  AO22X1_HVT U2642 ( .A1(\ram[10][43] ), .A2(n10199), .A3(n6447), .A4(n9437), 
        .Y(n2664) );
  AO22X1_HVT U2643 ( .A1(\ram[10][44] ), .A2(n7537), .A3(n6446), .A4(n9440), 
        .Y(n2665) );
  AO22X1_HVT U2644 ( .A1(\ram[10][45] ), .A2(n7536), .A3(n6471), .A4(n9443), 
        .Y(n2666) );
  AO22X1_HVT U2645 ( .A1(\ram[10][46] ), .A2(n7535), .A3(n6470), .A4(n9446), 
        .Y(n2667) );
  AO22X1_HVT U2646 ( .A1(\ram[10][47] ), .A2(n7490), .A3(n6469), .A4(n9449), 
        .Y(n2668) );
  AO22X1_HVT U2647 ( .A1(\ram[10][48] ), .A2(n7509), .A3(n6449), .A4(n9452), 
        .Y(n2669) );
  AO22X1_HVT U2648 ( .A1(\ram[10][49] ), .A2(n7508), .A3(n6421), .A4(n9455), 
        .Y(n2670) );
  AO22X1_HVT U2649 ( .A1(\ram[10][50] ), .A2(n7506), .A3(n6448), .A4(n9458), 
        .Y(n2671) );
  AO22X1_HVT U2650 ( .A1(\ram[10][51] ), .A2(n7505), .A3(n6422), .A4(n9461), 
        .Y(n2672) );
  AO22X1_HVT U2651 ( .A1(\ram[10][52] ), .A2(n7503), .A3(n6448), .A4(n9464), 
        .Y(n2673) );
  AO22X1_HVT U2652 ( .A1(\ram[10][53] ), .A2(n7502), .A3(n6468), .A4(n9467), 
        .Y(n2674) );
  AO22X1_HVT U2653 ( .A1(\ram[10][54] ), .A2(n7500), .A3(n10179), .A4(n9470), 
        .Y(n2675) );
  AO22X1_HVT U2654 ( .A1(\ram[10][55] ), .A2(n7499), .A3(n6467), .A4(n9473), 
        .Y(n2676) );
  AO22X1_HVT U2655 ( .A1(\ram[10][56] ), .A2(n7498), .A3(n6466), .A4(n9476), 
        .Y(n2677) );
  AO22X1_HVT U2656 ( .A1(\ram[10][57] ), .A2(n7497), .A3(n6463), .A4(n9479), 
        .Y(n2678) );
  AO22X1_HVT U2657 ( .A1(\ram[10][58] ), .A2(n7494), .A3(n6462), .A4(n9482), 
        .Y(n2679) );
  AO22X1_HVT U2658 ( .A1(\ram[10][59] ), .A2(n7493), .A3(n6460), .A4(n9485), 
        .Y(n2680) );
  AO22X1_HVT U2659 ( .A1(\ram[10][60] ), .A2(n7475), .A3(n6452), .A4(n9488), 
        .Y(n2681) );
  AO22X1_HVT U2660 ( .A1(\ram[10][61] ), .A2(n7538), .A3(n6449), .A4(n9491), 
        .Y(n2682) );
  AO22X1_HVT U2661 ( .A1(\ram[10][62] ), .A2(n7534), .A3(n6477), .A4(n9494), 
        .Y(n2683) );
  AO22X1_HVT U2662 ( .A1(\ram[10][63] ), .A2(n7537), .A3(n6448), .A4(n9497), 
        .Y(n2684) );
  AO22X1_HVT U2663 ( .A1(\ram[10][64] ), .A2(n7536), .A3(n6447), .A4(n9500), 
        .Y(n2685) );
  AO22X1_HVT U2664 ( .A1(\ram[10][65] ), .A2(n7535), .A3(n6446), .A4(n9503), 
        .Y(n2686) );
  AO22X1_HVT U2665 ( .A1(\ram[10][66] ), .A2(n7534), .A3(n6446), .A4(n9506), 
        .Y(n2687) );
  AO22X1_HVT U2666 ( .A1(\ram[10][67] ), .A2(n7531), .A3(n6445), .A4(n9509), 
        .Y(n2688) );
  AO22X1_HVT U2667 ( .A1(\ram[10][68] ), .A2(n7530), .A3(n6456), .A4(n9512), 
        .Y(n2689) );
  AO22X1_HVT U2668 ( .A1(\ram[10][69] ), .A2(n7527), .A3(n6455), .A4(n9515), 
        .Y(n2690) );
  AO22X1_HVT U2669 ( .A1(\ram[10][70] ), .A2(n7526), .A3(n6454), .A4(n9518), 
        .Y(n2691) );
  AO22X1_HVT U2670 ( .A1(\ram[10][71] ), .A2(n7524), .A3(n6453), .A4(n9521), 
        .Y(n2692) );
  AO22X1_HVT U2671 ( .A1(\ram[10][72] ), .A2(n7523), .A3(n6472), .A4(n9524), 
        .Y(n2693) );
  AO22X1_HVT U2672 ( .A1(\ram[10][73] ), .A2(n7522), .A3(n6471), .A4(n9527), 
        .Y(n2694) );
  AO22X1_HVT U2673 ( .A1(\ram[10][74] ), .A2(n7521), .A3(n6470), .A4(n9530), 
        .Y(n2695) );
  AO22X1_HVT U2674 ( .A1(\ram[10][75] ), .A2(n7519), .A3(n6472), .A4(n9533), 
        .Y(n2696) );
  AO22X1_HVT U2675 ( .A1(\ram[10][76] ), .A2(n7518), .A3(n6471), .A4(n9536), 
        .Y(n2697) );
  AO22X1_HVT U2676 ( .A1(\ram[10][77] ), .A2(n7483), .A3(n6470), .A4(n9539), 
        .Y(n2698) );
  AO22X1_HVT U2677 ( .A1(\ram[10][78] ), .A2(n7481), .A3(n6469), .A4(n9542), 
        .Y(n2699) );
  AO22X1_HVT U2678 ( .A1(\ram[10][79] ), .A2(n7480), .A3(n6468), .A4(n9545), 
        .Y(n2700) );
  AO22X1_HVT U2679 ( .A1(\ram[10][80] ), .A2(n7479), .A3(n10187), .A4(n9548), 
        .Y(n2701) );
  AO22X1_HVT U2680 ( .A1(\ram[10][81] ), .A2(n7478), .A3(n6467), .A4(n9551), 
        .Y(n2702) );
  AO22X1_HVT U2681 ( .A1(\ram[10][82] ), .A2(n7542), .A3(n6466), .A4(n9554), 
        .Y(n2703) );
  AO22X1_HVT U2682 ( .A1(\ram[10][83] ), .A2(n7541), .A3(n6463), .A4(n9557), 
        .Y(n2704) );
  AO22X1_HVT U2683 ( .A1(\ram[10][84] ), .A2(n7540), .A3(n10187), .A4(n9560), 
        .Y(n2705) );
  AO22X1_HVT U2684 ( .A1(\ram[10][85] ), .A2(n7526), .A3(n6467), .A4(n9563), 
        .Y(n2706) );
  AO22X1_HVT U2685 ( .A1(\ram[10][86] ), .A2(n7524), .A3(n6478), .A4(n9566), 
        .Y(n2707) );
  AO22X1_HVT U2686 ( .A1(\ram[10][87] ), .A2(n7523), .A3(n6427), .A4(n9569), 
        .Y(n2708) );
  AO22X1_HVT U2687 ( .A1(\ram[10][88] ), .A2(n7522), .A3(n6422), .A4(n9572), 
        .Y(n2709) );
  AO22X1_HVT U2688 ( .A1(\ram[10][89] ), .A2(n7476), .A3(n6418), .A4(n9575), 
        .Y(n2710) );
  AO22X1_HVT U2689 ( .A1(\ram[10][90] ), .A2(n7515), .A3(n6479), .A4(n9578), 
        .Y(n2711) );
  AO22X1_HVT U2690 ( .A1(\ram[10][91] ), .A2(n7514), .A3(n6478), .A4(n9581), 
        .Y(n2712) );
  AO22X1_HVT U2691 ( .A1(\ram[10][92] ), .A2(n7541), .A3(n6477), .A4(n9584), 
        .Y(n2713) );
  AO22X1_HVT U2692 ( .A1(\ram[10][93] ), .A2(n7540), .A3(n6476), .A4(n9587), 
        .Y(n2714) );
  AO22X1_HVT U2693 ( .A1(\ram[10][94] ), .A2(n7512), .A3(n6474), .A4(n9590), 
        .Y(n2715) );
  AO22X1_HVT U2694 ( .A1(\ram[10][95] ), .A2(n7511), .A3(n6473), .A4(n9593), 
        .Y(n2716) );
  AO22X1_HVT U2695 ( .A1(\ram[10][96] ), .A2(n7492), .A3(n6452), .A4(n9596), 
        .Y(n2717) );
  AO22X1_HVT U2696 ( .A1(\ram[10][97] ), .A2(n7491), .A3(n10180), .A4(n9599), 
        .Y(n2718) );
  AO22X1_HVT U2697 ( .A1(\ram[10][98] ), .A2(n7486), .A3(n6430), .A4(n9602), 
        .Y(n2719) );
  AO22X1_HVT U2698 ( .A1(\ram[10][99] ), .A2(n7485), .A3(n6428), .A4(n9605), 
        .Y(n2720) );
  AO22X1_HVT U2699 ( .A1(\ram[10][100] ), .A2(n7484), .A3(n6427), .A4(n9608), 
        .Y(n2721) );
  AO22X1_HVT U2700 ( .A1(\ram[10][101] ), .A2(n7483), .A3(n6422), .A4(n9611), 
        .Y(n2722) );
  AO22X1_HVT U2701 ( .A1(\ram[10][102] ), .A2(n7481), .A3(n6421), .A4(n9614), 
        .Y(n2723) );
  AO22X1_HVT U2702 ( .A1(\ram[10][103] ), .A2(n7480), .A3(n6420), .A4(n9617), 
        .Y(n2724) );
  AO22X1_HVT U2703 ( .A1(\ram[10][104] ), .A2(n7479), .A3(n6419), .A4(n9620), 
        .Y(n2725) );
  AO22X1_HVT U2704 ( .A1(\ram[10][105] ), .A2(n7478), .A3(n6418), .A4(n9623), 
        .Y(n2726) );
  AO22X1_HVT U2705 ( .A1(\ram[10][106] ), .A2(n7542), .A3(n6469), .A4(n9626), 
        .Y(n2727) );
  AO22X1_HVT U2706 ( .A1(\ram[10][107] ), .A2(n7541), .A3(n6468), .A4(n9629), 
        .Y(n2728) );
  AO22X1_HVT U2707 ( .A1(\ram[10][108] ), .A2(n7540), .A3(n6471), .A4(n9632), 
        .Y(n2729) );
  AO22X1_HVT U2708 ( .A1(\ram[10][109] ), .A2(n7539), .A3(n6449), .A4(n9635), 
        .Y(n2730) );
  AO22X1_HVT U2709 ( .A1(\ram[10][110] ), .A2(n10195), .A3(n6428), .A4(n9638), 
        .Y(n2731) );
  AO22X1_HVT U2710 ( .A1(\ram[10][111] ), .A2(n7490), .A3(n6427), .A4(n9641), 
        .Y(n2732) );
  AO22X1_HVT U2711 ( .A1(\ram[10][112] ), .A2(n7489), .A3(n6422), .A4(n9644), 
        .Y(n2733) );
  AO22X1_HVT U2712 ( .A1(\ram[10][113] ), .A2(n7476), .A3(n6421), .A4(n9647), 
        .Y(n2734) );
  AO22X1_HVT U2713 ( .A1(\ram[10][114] ), .A2(n7475), .A3(n6420), .A4(n9650), 
        .Y(n2735) );
  AO22X1_HVT U2714 ( .A1(\ram[10][115] ), .A2(n7538), .A3(n6419), .A4(n9653), 
        .Y(n2736) );
  AO22X1_HVT U2715 ( .A1(\ram[10][116] ), .A2(n7539), .A3(n6418), .A4(n9656), 
        .Y(n2737) );
  AO22X1_HVT U2716 ( .A1(\ram[10][117] ), .A2(n7499), .A3(n6479), .A4(n9659), 
        .Y(n2738) );
  AO22X1_HVT U2717 ( .A1(\ram[10][118] ), .A2(n7490), .A3(n6478), .A4(n9662), 
        .Y(n2739) );
  AO22X1_HVT U2718 ( .A1(\ram[10][119] ), .A2(n7489), .A3(n6477), .A4(n9665), 
        .Y(n2740) );
  AO22X1_HVT U2719 ( .A1(\ram[10][120] ), .A2(n7539), .A3(n6427), .A4(n9668), 
        .Y(n2741) );
  AO22X1_HVT U2720 ( .A1(\ram[10][121] ), .A2(n7490), .A3(n6422), .A4(n9671), 
        .Y(n2742) );
  AO22X1_HVT U2721 ( .A1(\ram[10][122] ), .A2(n7480), .A3(n6421), .A4(n9674), 
        .Y(n2743) );
  AO22X1_HVT U2722 ( .A1(\ram[10][123] ), .A2(n7479), .A3(n6420), .A4(n9677), 
        .Y(n2744) );
  AO22X1_HVT U2723 ( .A1(\ram[10][124] ), .A2(n7489), .A3(n6419), .A4(n9680), 
        .Y(n2745) );
  AO22X1_HVT U2724 ( .A1(\ram[10][125] ), .A2(n7476), .A3(n6418), .A4(n9683), 
        .Y(n2746) );
  AO22X1_HVT U2725 ( .A1(\ram[10][126] ), .A2(n7475), .A3(n6479), .A4(n9686), 
        .Y(n2747) );
  AO22X1_HVT U2726 ( .A1(\ram[10][127] ), .A2(n7538), .A3(n6478), .A4(n9689), 
        .Y(n2748) );
  AO22X1_HVT U2727 ( .A1(\ram[10][128] ), .A2(n10192), .A3(n6477), .A4(n9692), 
        .Y(n2749) );
  AO22X1_HVT U2728 ( .A1(\ram[10][129] ), .A2(n7537), .A3(n6476), .A4(n9695), 
        .Y(n2750) );
  AO22X1_HVT U2729 ( .A1(\ram[10][130] ), .A2(n7536), .A3(n6474), .A4(n9698), 
        .Y(n2751) );
  AO22X1_HVT U2730 ( .A1(\ram[10][131] ), .A2(n7535), .A3(n6473), .A4(n9701), 
        .Y(n2752) );
  AO22X1_HVT U2731 ( .A1(\ram[10][132] ), .A2(n7534), .A3(n6443), .A4(n9704), 
        .Y(n2753) );
  AO22X1_HVT U2732 ( .A1(\ram[10][133] ), .A2(n7531), .A3(n6440), .A4(n9707), 
        .Y(n2754) );
  AO22X1_HVT U2733 ( .A1(\ram[10][134] ), .A2(n7530), .A3(n6439), .A4(n9710), 
        .Y(n2755) );
  AO22X1_HVT U2734 ( .A1(\ram[10][135] ), .A2(n7527), .A3(n6438), .A4(n9713), 
        .Y(n2756) );
  AO22X1_HVT U2735 ( .A1(\ram[10][136] ), .A2(n7526), .A3(n6437), .A4(n9716), 
        .Y(n2757) );
  AO22X1_HVT U2736 ( .A1(\ram[10][137] ), .A2(n7524), .A3(n6434), .A4(n9719), 
        .Y(n2758) );
  AO22X1_HVT U2737 ( .A1(\ram[10][138] ), .A2(n7523), .A3(n6433), .A4(n9722), 
        .Y(n2759) );
  AO22X1_HVT U2738 ( .A1(\ram[10][139] ), .A2(n7522), .A3(n6431), .A4(n9725), 
        .Y(n2760) );
  AO22X1_HVT U2739 ( .A1(\ram[10][140] ), .A2(n7521), .A3(n6430), .A4(n9729), 
        .Y(n2761) );
  AO22X1_HVT U2740 ( .A1(\ram[10][141] ), .A2(n7519), .A3(n4199), .A4(n9732), 
        .Y(n2762) );
  AO22X1_HVT U2741 ( .A1(\ram[10][142] ), .A2(n7518), .A3(n6424), .A4(
        data[142]), .Y(n2763) );
  AO22X1_HVT U2742 ( .A1(\ram[10][143] ), .A2(n7515), .A3(n6443), .A4(n9738), 
        .Y(n2764) );
  AO22X1_HVT U2743 ( .A1(\ram[10][144] ), .A2(n7514), .A3(n6440), .A4(n9742), 
        .Y(n2765) );
  AO22X1_HVT U2744 ( .A1(\ram[10][145] ), .A2(n7512), .A3(n6439), .A4(n9745), 
        .Y(n2766) );
  AO22X1_HVT U2745 ( .A1(\ram[10][146] ), .A2(n7511), .A3(n6438), .A4(n9748), 
        .Y(n2767) );
  AO22X1_HVT U2746 ( .A1(\ram[10][147] ), .A2(n7509), .A3(n6437), .A4(n9751), 
        .Y(n2768) );
  AO22X1_HVT U2747 ( .A1(\ram[10][148] ), .A2(n7508), .A3(n6434), .A4(n9755), 
        .Y(n2769) );
  AO22X1_HVT U2748 ( .A1(\ram[10][149] ), .A2(n7506), .A3(n6433), .A4(n9758), 
        .Y(n2770) );
  AO22X1_HVT U2749 ( .A1(\ram[10][150] ), .A2(n7505), .A3(n6431), .A4(n9761), 
        .Y(n2771) );
  AO22X1_HVT U2750 ( .A1(\ram[10][151] ), .A2(n7503), .A3(n6430), .A4(n9764), 
        .Y(n2772) );
  AO22X1_HVT U2751 ( .A1(\ram[10][152] ), .A2(n7502), .A3(n6428), .A4(n9767), 
        .Y(n2773) );
  AO22X1_HVT U2752 ( .A1(\ram[10][153] ), .A2(n7500), .A3(n6424), .A4(n9770), 
        .Y(n2774) );
  AO22X1_HVT U2753 ( .A1(\ram[10][154] ), .A2(n7499), .A3(n6452), .A4(n9773), 
        .Y(n2775) );
  AO22X1_HVT U2754 ( .A1(\ram[10][155] ), .A2(n7498), .A3(n6444), .A4(n9776), 
        .Y(n2776) );
  AO22X1_HVT U2755 ( .A1(\ram[10][156] ), .A2(n7497), .A3(n6430), .A4(n9780), 
        .Y(n2777) );
  AO22X1_HVT U2756 ( .A1(\ram[10][157] ), .A2(n7494), .A3(n6428), .A4(n9783), 
        .Y(n2778) );
  AO22X1_HVT U2757 ( .A1(\ram[10][158] ), .A2(n7497), .A3(n6434), .A4(n9786), 
        .Y(n2779) );
  AO22X1_HVT U2758 ( .A1(\ram[10][159] ), .A2(n7494), .A3(n6433), .A4(n9789), 
        .Y(n2780) );
  AO22X1_HVT U2759 ( .A1(\ram[10][160] ), .A2(n7493), .A3(n6431), .A4(n9793), 
        .Y(n2781) );
  AO22X1_HVT U2760 ( .A1(\ram[10][161] ), .A2(n7492), .A3(n6430), .A4(n9796), 
        .Y(n2782) );
  AO22X1_HVT U2761 ( .A1(\ram[10][162] ), .A2(n7491), .A3(n6428), .A4(n9799), 
        .Y(n2783) );
  AO22X1_HVT U2762 ( .A1(\ram[10][163] ), .A2(n7486), .A3(n6427), .A4(n9802), 
        .Y(n2784) );
  AO22X1_HVT U2763 ( .A1(\ram[10][164] ), .A2(n7485), .A3(n6422), .A4(n9805), 
        .Y(n2785) );
  AO22X1_HVT U2764 ( .A1(\ram[10][165] ), .A2(n7484), .A3(n6421), .A4(n9808), 
        .Y(n2786) );
  AO22X1_HVT U2765 ( .A1(\ram[10][166] ), .A2(n7534), .A3(n6420), .A4(n9811), 
        .Y(n2787) );
  AO22X1_HVT U2766 ( .A1(\ram[10][167] ), .A2(n7531), .A3(n6419), .A4(n9814), 
        .Y(n2788) );
  AO22X1_HVT U2767 ( .A1(\ram[10][168] ), .A2(n7530), .A3(n6440), .A4(n9817), 
        .Y(n2789) );
  AO22X1_HVT U2768 ( .A1(\ram[10][169] ), .A2(n7527), .A3(n6439), .A4(n9820), 
        .Y(n2790) );
  AO22X1_HVT U2769 ( .A1(\ram[10][170] ), .A2(n7489), .A3(n6438), .A4(n9823), 
        .Y(n2791) );
  AO22X1_HVT U2770 ( .A1(\ram[10][171] ), .A2(n7493), .A3(n6437), .A4(n9826), 
        .Y(n2792) );
  AO22X1_HVT U2771 ( .A1(\ram[10][172] ), .A2(n7492), .A3(n6434), .A4(n9830), 
        .Y(n2793) );
  AO22X1_HVT U2772 ( .A1(\ram[10][173] ), .A2(n7478), .A3(n6433), .A4(n9833), 
        .Y(n2794) );
  AO22X1_HVT U2773 ( .A1(\ram[10][174] ), .A2(n7542), .A3(n6431), .A4(n9836), 
        .Y(n2795) );
  AO22X1_HVT U2774 ( .A1(\ram[10][175] ), .A2(n7491), .A3(n6473), .A4(n9839), 
        .Y(n2796) );
  AO22X1_HVT U2775 ( .A1(\ram[10][176] ), .A2(n7486), .A3(n6472), .A4(n9843), 
        .Y(n2797) );
  AO22X1_HVT U2776 ( .A1(\ram[10][177] ), .A2(n7485), .A3(n6471), .A4(n9846), 
        .Y(n2798) );
  AO22X1_HVT U2777 ( .A1(\ram[10][178] ), .A2(n7484), .A3(n6470), .A4(n9849), 
        .Y(n2799) );
  AO22X1_HVT U2778 ( .A1(\ram[10][179] ), .A2(n7483), .A3(n6479), .A4(n9852), 
        .Y(n2800) );
  AO22X1_HVT U2779 ( .A1(\ram[10][180] ), .A2(n7481), .A3(n6447), .A4(n9856), 
        .Y(n2801) );
  AO22X1_HVT U2780 ( .A1(\ram[10][181] ), .A2(n7480), .A3(n6446), .A4(n9859), 
        .Y(n2802) );
  AO22X1_HVT U2781 ( .A1(\ram[10][182] ), .A2(n7479), .A3(n6445), .A4(n9862), 
        .Y(n2803) );
  AO22X1_HVT U2782 ( .A1(\ram[10][183] ), .A2(n7478), .A3(n6444), .A4(n9865), 
        .Y(n2804) );
  AO22X1_HVT U2783 ( .A1(\ram[10][184] ), .A2(n7542), .A3(n6443), .A4(n9869), 
        .Y(n2805) );
  AO22X1_HVT U2784 ( .A1(\ram[10][185] ), .A2(n7541), .A3(n6440), .A4(n9872), 
        .Y(n2806) );
  AO22X1_HVT U2785 ( .A1(\ram[10][186] ), .A2(n7540), .A3(n6439), .A4(n9875), 
        .Y(n2807) );
  AO22X1_HVT U2786 ( .A1(\ram[10][187] ), .A2(n7539), .A3(n6438), .A4(n9878), 
        .Y(n2808) );
  AO22X1_HVT U2787 ( .A1(\ram[10][188] ), .A2(n10191), .A3(n6437), .A4(n9881), 
        .Y(n2809) );
  AO22X1_HVT U2788 ( .A1(\ram[10][189] ), .A2(n7490), .A3(n6445), .A4(n9884), 
        .Y(n2810) );
  AO22X1_HVT U2789 ( .A1(\ram[10][190] ), .A2(n7489), .A3(n6444), .A4(n9887), 
        .Y(n2811) );
  AO22X1_HVT U2790 ( .A1(\ram[10][191] ), .A2(n7476), .A3(n6443), .A4(n9890), 
        .Y(n2812) );
  AO22X1_HVT U2791 ( .A1(\ram[10][192] ), .A2(n7476), .A3(n6466), .A4(n9894), 
        .Y(n2813) );
  AO22X1_HVT U2792 ( .A1(\ram[10][193] ), .A2(n7475), .A3(n6463), .A4(n9897), 
        .Y(n2814) );
  AO22X1_HVT U2793 ( .A1(\ram[10][194] ), .A2(n7538), .A3(n6462), .A4(n9900), 
        .Y(n2815) );
  AO22X1_HVT U2794 ( .A1(\ram[10][195] ), .A2(n7512), .A3(n6460), .A4(n9903), 
        .Y(n2816) );
  AO22X1_HVT U2795 ( .A1(\ram[10][196] ), .A2(n7521), .A3(n6459), .A4(n9907), 
        .Y(n2817) );
  AO22X1_HVT U2796 ( .A1(\ram[10][197] ), .A2(n7519), .A3(n10183), .A4(n9910), 
        .Y(n2818) );
  AO22X1_HVT U2797 ( .A1(\ram[10][198] ), .A2(n7518), .A3(n6457), .A4(n9913), 
        .Y(n2819) );
  AO22X1_HVT U2798 ( .A1(\ram[10][199] ), .A2(n7515), .A3(n6455), .A4(n9916), 
        .Y(n2820) );
  AO22X1_HVT U2799 ( .A1(\ram[10][200] ), .A2(n7475), .A3(n6454), .A4(n9920), 
        .Y(n2821) );
  AO22X1_HVT U2800 ( .A1(\ram[10][201] ), .A2(n7535), .A3(n6453), .A4(n9923), 
        .Y(n2822) );
  AO22X1_HVT U2801 ( .A1(\ram[10][202] ), .A2(n7537), .A3(n6425), .A4(n9926), 
        .Y(n2823) );
  AO22X1_HVT U2802 ( .A1(\ram[10][203] ), .A2(n7539), .A3(n6474), .A4(n9929), 
        .Y(n2824) );
  AO22X1_HVT U2803 ( .A1(\ram[10][204] ), .A2(n7486), .A3(n10184), .A4(n9932), 
        .Y(n2825) );
  AO22X1_HVT U2804 ( .A1(\ram[10][205] ), .A2(n7536), .A3(n6457), .A4(n9935), 
        .Y(n2826) );
  AO22X1_HVT U2805 ( .A1(\ram[10][206] ), .A2(n7535), .A3(n6456), .A4(n9938), 
        .Y(n2827) );
  AO22X1_HVT U2806 ( .A1(\ram[10][207] ), .A2(n7534), .A3(n6455), .A4(n9941), 
        .Y(n2828) );
  AO22X1_HVT U2807 ( .A1(\ram[10][208] ), .A2(n7531), .A3(n6454), .A4(n9945), 
        .Y(n2829) );
  AO22X1_HVT U2808 ( .A1(\ram[10][209] ), .A2(n7530), .A3(n6453), .A4(n9948), 
        .Y(n2830) );
  AO22X1_HVT U2809 ( .A1(\ram[10][210] ), .A2(n7527), .A3(n4199), .A4(n9951), 
        .Y(n2831) );
  AO22X1_HVT U2810 ( .A1(\ram[10][211] ), .A2(n7526), .A3(n6424), .A4(n9954), 
        .Y(n2832) );
  AO22X1_HVT U2811 ( .A1(\ram[10][212] ), .A2(n7524), .A3(n6452), .A4(n9957), 
        .Y(n2833) );
  AO22X1_HVT U2812 ( .A1(\ram[10][213] ), .A2(n7523), .A3(n6448), .A4(n9960), 
        .Y(n2834) );
  AO22X1_HVT U2813 ( .A1(\ram[10][214] ), .A2(n7522), .A3(n6447), .A4(n9963), 
        .Y(n2835) );
  AO22X1_HVT U2814 ( .A1(\ram[10][215] ), .A2(n7521), .A3(n6467), .A4(n9966), 
        .Y(n2836) );
  AO22X1_HVT U2815 ( .A1(\ram[10][216] ), .A2(n7519), .A3(n6454), .A4(n9969), 
        .Y(n2837) );
  AO22X1_HVT U2816 ( .A1(\ram[10][217] ), .A2(n7518), .A3(n6453), .A4(n9972), 
        .Y(n2838) );
  AO22X1_HVT U2817 ( .A1(\ram[10][218] ), .A2(n7515), .A3(n4199), .A4(n9975), 
        .Y(n2839) );
  AO22X1_HVT U2818 ( .A1(\ram[10][219] ), .A2(n7514), .A3(n6424), .A4(n9978), 
        .Y(n2840) );
  AO22X1_HVT U2819 ( .A1(\ram[10][220] ), .A2(n7512), .A3(n6452), .A4(n9982), 
        .Y(n2841) );
  AO22X1_HVT U2820 ( .A1(\ram[10][221] ), .A2(n7511), .A3(n6445), .A4(n9985), 
        .Y(n2842) );
  AO22X1_HVT U2821 ( .A1(\ram[10][222] ), .A2(n7509), .A3(n6449), .A4(n9988), 
        .Y(n2843) );
  AO22X1_HVT U2822 ( .A1(\ram[10][223] ), .A2(n7508), .A3(n6419), .A4(n9991), 
        .Y(n2844) );
  AO22X1_HVT U2823 ( .A1(\ram[10][224] ), .A2(n7506), .A3(n6448), .A4(n9994), 
        .Y(n2845) );
  AO22X1_HVT U2824 ( .A1(\ram[10][225] ), .A2(n7505), .A3(n6445), .A4(n9997), 
        .Y(n2846) );
  AO22X1_HVT U2825 ( .A1(\ram[10][226] ), .A2(n7503), .A3(n6444), .A4(n10000), 
        .Y(n2847) );
  AO22X1_HVT U2826 ( .A1(\ram[10][227] ), .A2(n7502), .A3(n6459), .A4(n10003), 
        .Y(n2848) );
  AO22X1_HVT U2827 ( .A1(\ram[10][228] ), .A2(n7500), .A3(n6446), .A4(n10006), 
        .Y(n2849) );
  AO22X1_HVT U2828 ( .A1(\ram[10][229] ), .A2(n7499), .A3(n6445), .A4(n10009), 
        .Y(n2850) );
  AO22X1_HVT U2829 ( .A1(\ram[10][230] ), .A2(n7498), .A3(n6444), .A4(n10012), 
        .Y(n2851) );
  AO22X1_HVT U2830 ( .A1(\ram[10][231] ), .A2(n7497), .A3(n6443), .A4(n10015), 
        .Y(n2852) );
  AO22X1_HVT U2831 ( .A1(\ram[10][232] ), .A2(n7494), .A3(n6440), .A4(n10019), 
        .Y(n2853) );
  AO22X1_HVT U2832 ( .A1(\ram[10][233] ), .A2(n7493), .A3(n6439), .A4(n10022), 
        .Y(n2854) );
  AO22X1_HVT U2833 ( .A1(\ram[10][234] ), .A2(n7492), .A3(n6438), .A4(n10025), 
        .Y(n2855) );
  AO22X1_HVT U2834 ( .A1(\ram[10][235] ), .A2(n7491), .A3(n6437), .A4(n10028), 
        .Y(n2856) );
  AO22X1_HVT U2835 ( .A1(\ram[10][236] ), .A2(n7486), .A3(n6434), .A4(n10031), 
        .Y(n2857) );
  AO22X1_HVT U2836 ( .A1(\ram[10][237] ), .A2(n7485), .A3(n6457), .A4(n10034), 
        .Y(n2858) );
  AO22X1_HVT U2837 ( .A1(\ram[10][238] ), .A2(n7484), .A3(n6456), .A4(n10037), 
        .Y(n2859) );
  AO22X1_HVT U2838 ( .A1(\ram[10][239] ), .A2(n7537), .A3(n6455), .A4(n10040), 
        .Y(n2860) );
  AO22X1_HVT U2839 ( .A1(\ram[10][240] ), .A2(n7536), .A3(n6470), .A4(n10044), 
        .Y(n2861) );
  AO22X1_HVT U2840 ( .A1(\ram[10][241] ), .A2(n7535), .A3(n6469), .A4(n10047), 
        .Y(n2862) );
  AO22X1_HVT U2841 ( .A1(\ram[10][242] ), .A2(n7534), .A3(n6468), .A4(n10050), 
        .Y(n2863) );
  AO22X1_HVT U2842 ( .A1(\ram[10][243] ), .A2(n7531), .A3(n10187), .A4(n10053), 
        .Y(n2864) );
  AO22X1_HVT U2843 ( .A1(\ram[10][244] ), .A2(n7530), .A3(n6459), .A4(n10056), 
        .Y(n2865) );
  AO22X1_HVT U2844 ( .A1(\ram[10][245] ), .A2(n7527), .A3(n10184), .A4(n10059), 
        .Y(n2866) );
  AO22X1_HVT U2845 ( .A1(\ram[10][246] ), .A2(n7526), .A3(n6457), .A4(n10062), 
        .Y(n2867) );
  AO22X1_HVT U2846 ( .A1(\ram[10][247] ), .A2(n7514), .A3(n6456), .A4(n10065), 
        .Y(n2868) );
  AO22X1_HVT U2847 ( .A1(\ram[10][248] ), .A2(n7512), .A3(n6476), .A4(n10069), 
        .Y(n2869) );
  AO22X1_HVT U2848 ( .A1(\ram[10][249] ), .A2(n7511), .A3(n6419), .A4(n10072), 
        .Y(n2870) );
  AO22X1_HVT U2849 ( .A1(\ram[10][250] ), .A2(n7509), .A3(n6418), .A4(n10075), 
        .Y(n2871) );
  AO22X1_HVT U2850 ( .A1(\ram[10][251] ), .A2(n7538), .A3(n6447), .A4(n10078), 
        .Y(n2872) );
  AO22X1_HVT U2851 ( .A1(\ram[10][252] ), .A2(n7540), .A3(n6418), .A4(n10082), 
        .Y(n2873) );
  AO22X1_HVT U2852 ( .A1(\ram[10][253] ), .A2(n7524), .A3(n6433), .A4(n10085), 
        .Y(n2874) );
  AO22X1_HVT U2853 ( .A1(\ram[10][254] ), .A2(n7523), .A3(n6431), .A4(n10088), 
        .Y(n2875) );
  AO22X1_HVT U2854 ( .A1(\ram[10][255] ), .A2(n7483), .A3(n6462), .A4(n10091), 
        .Y(n2876) );
  AND2X1_HVT U2857 ( .A1(n38), .A2(n6644), .Y(n44) );
  AO22X1_HVT U2858 ( .A1(\ram[11][0] ), .A2(n7423), .A3(n6787), .A4(data[0]), 
        .Y(n2877) );
  AO22X1_HVT U2859 ( .A1(\ram[11][1] ), .A2(n7452), .A3(n6771), .A4(data[1]), 
        .Y(n2878) );
  AO22X1_HVT U2860 ( .A1(\ram[11][2] ), .A2(n10169), .A3(n6802), .A4(n9313), 
        .Y(n2879) );
  AO22X1_HVT U2861 ( .A1(\ram[11][3] ), .A2(n7451), .A3(n6825), .A4(n9317), 
        .Y(n2880) );
  AO22X1_HVT U2862 ( .A1(\ram[11][4] ), .A2(n7450), .A3(n6824), .A4(data[4]), 
        .Y(n2881) );
  AO22X1_HVT U2863 ( .A1(\ram[11][5] ), .A2(n7438), .A3(n6823), .A4(data[5]), 
        .Y(n2882) );
  AO22X1_HVT U2864 ( .A1(\ram[11][6] ), .A2(n7467), .A3(n6822), .A4(data[6]), 
        .Y(n2883) );
  AO22X1_HVT U2866 ( .A1(\ram[11][8] ), .A2(n7444), .A3(n10153), .A4(data[8]), 
        .Y(n2885) );
  AO22X1_HVT U2867 ( .A1(\ram[11][9] ), .A2(n7443), .A3(n6820), .A4(data[9]), 
        .Y(n2886) );
  AO22X1_HVT U2868 ( .A1(\ram[11][10] ), .A2(n7442), .A3(n6786), .A4(data[10]), 
        .Y(n2887) );
  AO22X1_HVT U2869 ( .A1(\ram[11][11] ), .A2(n10171), .A3(n6785), .A4(n9342), 
        .Y(n2888) );
  AO22X1_HVT U2870 ( .A1(\ram[11][12] ), .A2(n10168), .A3(n6783), .A4(data[12]), .Y(n2889) );
  AO22X1_HVT U2871 ( .A1(\ram[11][13] ), .A2(n10170), .A3(n6782), .A4(data[13]), .Y(n2890) );
  AO22X1_HVT U2872 ( .A1(\ram[11][14] ), .A2(n7441), .A3(n6779), .A4(data[14]), 
        .Y(n2891) );
  AO22X1_HVT U2873 ( .A1(\ram[11][15] ), .A2(n7440), .A3(n6777), .A4(data[15]), 
        .Y(n2892) );
  AO22X1_HVT U2874 ( .A1(\ram[11][16] ), .A2(n7439), .A3(n6776), .A4(data[16]), 
        .Y(n2893) );
  AO22X1_HVT U2875 ( .A1(\ram[11][17] ), .A2(n7438), .A3(n6774), .A4(data[17]), 
        .Y(n2894) );
  AO22X1_HVT U2876 ( .A1(\ram[11][18] ), .A2(n10168), .A3(n6773), .A4(data[18]), .Y(n2895) );
  AO22X1_HVT U2877 ( .A1(\ram[11][19] ), .A2(n7436), .A3(n6772), .A4(data[19]), 
        .Y(n2896) );
  AO22X1_HVT U2878 ( .A1(\ram[11][20] ), .A2(n7435), .A3(n6771), .A4(data[20]), 
        .Y(n2897) );
  AO22X1_HVT U2879 ( .A1(\ram[11][21] ), .A2(n7434), .A3(n6770), .A4(data[21]), 
        .Y(n2898) );
  AO22X1_HVT U2880 ( .A1(\ram[11][22] ), .A2(n7433), .A3(n6791), .A4(data[22]), 
        .Y(n2899) );
  AO22X1_HVT U2881 ( .A1(\ram[11][23] ), .A2(n7427), .A3(n6789), .A4(data[23]), 
        .Y(n2900) );
  AO22X1_HVT U2882 ( .A1(\ram[11][24] ), .A2(n7435), .A3(n10160), .A4(data[24]), .Y(n2901) );
  AO22X1_HVT U2883 ( .A1(\ram[11][25] ), .A2(n7426), .A3(n6788), .A4(data[25]), 
        .Y(n2902) );
  AO22X1_HVT U2884 ( .A1(\ram[11][26] ), .A2(n7425), .A3(n6801), .A4(data[26]), 
        .Y(n2903) );
  AO22X1_HVT U2885 ( .A1(\ram[11][27] ), .A2(n7422), .A3(n6809), .A4(data[27]), 
        .Y(n2904) );
  AO22X1_HVT U2886 ( .A1(\ram[11][28] ), .A2(n7423), .A3(n10159), .A4(data[28]), .Y(n2905) );
  AO22X1_HVT U2888 ( .A1(\ram[11][30] ), .A2(n7419), .A3(n6825), .A4(n9398), 
        .Y(n2907) );
  AO22X1_HVT U2892 ( .A1(\ram[11][34] ), .A2(n7471), .A3(n6821), .A4(data[34]), 
        .Y(n2911) );
  AO22X1_HVT U2893 ( .A1(\ram[11][35] ), .A2(n7442), .A3(n10152), .A4(data[35]), .Y(n2912) );
  AO22X1_HVT U2894 ( .A1(\ram[11][36] ), .A2(n10166), .A3(n6820), .A4(data[36]), .Y(n2913) );
  AO22X1_HVT U2895 ( .A1(\ram[11][37] ), .A2(n10168), .A3(n6819), .A4(data[37]), .Y(n2914) );
  AO22X1_HVT U2896 ( .A1(\ram[11][38] ), .A2(n10170), .A3(n6814), .A4(data[38]), .Y(n2915) );
  AO22X1_HVT U2897 ( .A1(\ram[11][39] ), .A2(n7441), .A3(n6813), .A4(n9425), 
        .Y(n2916) );
  AO22X1_HVT U2898 ( .A1(\ram[11][40] ), .A2(n7440), .A3(n6811), .A4(data[40]), 
        .Y(n2917) );
  AO22X1_HVT U2899 ( .A1(\ram[11][41] ), .A2(n7439), .A3(n10159), .A4(data[41]), .Y(n2918) );
  AO22X1_HVT U2900 ( .A1(\ram[11][42] ), .A2(n7448), .A3(n6808), .A4(data[42]), 
        .Y(n2919) );
  AO22X1_HVT U2901 ( .A1(\ram[11][43] ), .A2(n7447), .A3(n6823), .A4(data[43]), 
        .Y(n2920) );
  AO22X1_HVT U2902 ( .A1(\ram[11][44] ), .A2(n7431), .A3(n6822), .A4(data[44]), 
        .Y(n2921) );
  AO22X1_HVT U2903 ( .A1(\ram[11][45] ), .A2(n7430), .A3(n6821), .A4(data[45]), 
        .Y(n2922) );
  AO22X1_HVT U2904 ( .A1(\ram[11][46] ), .A2(n7464), .A3(n10160), .A4(data[46]), .Y(n2923) );
  AO22X1_HVT U2905 ( .A1(\ram[11][47] ), .A2(n7431), .A3(n6820), .A4(data[47]), 
        .Y(n2924) );
  AO22X1_HVT U2906 ( .A1(\ram[11][48] ), .A2(n7470), .A3(n6821), .A4(data[48]), 
        .Y(n2925) );
  AO22X1_HVT U2907 ( .A1(\ram[11][49] ), .A2(n4431), .A3(n6774), .A4(data[49]), 
        .Y(n2926) );
  AO22X1_HVT U2908 ( .A1(\ram[11][50] ), .A2(n7422), .A3(n6779), .A4(data[50]), 
        .Y(n2927) );
  AO22X1_HVT U2909 ( .A1(\ram[11][51] ), .A2(n7420), .A3(n6805), .A4(data[51]), 
        .Y(n2928) );
  AO22X1_HVT U2910 ( .A1(\ram[11][52] ), .A2(n4314), .A3(n6777), .A4(data[52]), 
        .Y(n2929) );
  AO22X1_HVT U2911 ( .A1(\ram[11][53] ), .A2(n10168), .A3(n6819), .A4(data[53]), .Y(n2930) );
  AO22X1_HVT U2912 ( .A1(\ram[11][54] ), .A2(n10173), .A3(n6822), .A4(n9469), 
        .Y(n2931) );
  AO22X1_HVT U2913 ( .A1(\ram[11][55] ), .A2(n7468), .A3(n6773), .A4(data[55]), 
        .Y(n2932) );
  AO22X1_HVT U2914 ( .A1(\ram[11][56] ), .A2(n7467), .A3(n6780), .A4(data[56]), 
        .Y(n2933) );
  AO22X1_HVT U2915 ( .A1(\ram[11][57] ), .A2(n4426), .A3(n6817), .A4(data[57]), 
        .Y(n2934) );
  AO22X1_HVT U2916 ( .A1(\ram[11][58] ), .A2(n7430), .A3(n6779), .A4(data[58]), 
        .Y(n2935) );
  AO22X1_HVT U2917 ( .A1(\ram[11][59] ), .A2(n7464), .A3(n6813), .A4(data[59]), 
        .Y(n2936) );
  AO22X1_HVT U2918 ( .A1(\ram[11][60] ), .A2(n7463), .A3(n6824), .A4(data[60]), 
        .Y(n2937) );
  AO22X1_HVT U2919 ( .A1(\ram[11][61] ), .A2(n7461), .A3(n6771), .A4(data[61]), 
        .Y(n2938) );
  AO22X1_HVT U2920 ( .A1(\ram[11][62] ), .A2(n7460), .A3(n6776), .A4(data[62]), 
        .Y(n2939) );
  AO22X1_HVT U2921 ( .A1(\ram[11][63] ), .A2(n7458), .A3(n6786), .A4(data[63]), 
        .Y(n2940) );
  AO22X1_HVT U2922 ( .A1(\ram[11][64] ), .A2(n7457), .A3(n6802), .A4(data[64]), 
        .Y(n2941) );
  AO22X1_HVT U2923 ( .A1(\ram[11][65] ), .A2(n7455), .A3(n6813), .A4(data[65]), 
        .Y(n2942) );
  AO22X1_HVT U2924 ( .A1(\ram[11][66] ), .A2(n7454), .A3(n6823), .A4(data[66]), 
        .Y(n2943) );
  AO22X1_HVT U2925 ( .A1(\ram[11][67] ), .A2(n7452), .A3(n6772), .A4(data[67]), 
        .Y(n2944) );
  AO22X1_HVT U2926 ( .A1(\ram[11][68] ), .A2(n10172), .A3(n6777), .A4(data[68]), .Y(n2945) );
  AO22X1_HVT U2927 ( .A1(\ram[11][69] ), .A2(n7451), .A3(n10152), .A4(data[69]), .Y(n2946) );
  AO22X1_HVT U2928 ( .A1(\ram[11][70] ), .A2(n7450), .A3(n6776), .A4(data[70]), 
        .Y(n2947) );
  AO22X1_HVT U2929 ( .A1(\ram[11][71] ), .A2(n7448), .A3(n6814), .A4(data[71]), 
        .Y(n2948) );
  AO22X1_HVT U2930 ( .A1(\ram[11][72] ), .A2(n7447), .A3(n6797), .A4(n9524), 
        .Y(n2949) );
  AO22X1_HVT U2931 ( .A1(\ram[11][73] ), .A2(n7445), .A3(n6825), .A4(data[73]), 
        .Y(n2950) );
  AO22X1_HVT U2932 ( .A1(\ram[11][74] ), .A2(n7444), .A3(n6805), .A4(data[74]), 
        .Y(n2951) );
  AO22X1_HVT U2933 ( .A1(\ram[11][75] ), .A2(n7443), .A3(n10155), .A4(data[75]), .Y(n2952) );
  AO22X1_HVT U2934 ( .A1(\ram[11][76] ), .A2(n7442), .A3(n6794), .A4(data[76]), 
        .Y(n2953) );
  AO22X1_HVT U2935 ( .A1(\ram[11][77] ), .A2(n10174), .A3(n10158), .A4(
        data[77]), .Y(n2954) );
  AO22X1_HVT U2936 ( .A1(\ram[11][78] ), .A2(n10169), .A3(n6814), .A4(data[78]), .Y(n2955) );
  AO22X1_HVT U2937 ( .A1(\ram[11][79] ), .A2(n10169), .A3(n6799), .A4(data[79]), .Y(n2956) );
  AO22X1_HVT U2938 ( .A1(\ram[11][80] ), .A2(n7441), .A3(n6770), .A4(data[80]), 
        .Y(n2957) );
  AO22X1_HVT U2939 ( .A1(\ram[11][81] ), .A2(n7440), .A3(n10153), .A4(data[81]), .Y(n2958) );
  AO22X1_HVT U2940 ( .A1(\ram[11][82] ), .A2(n7439), .A3(n6796), .A4(data[82]), 
        .Y(n2959) );
  AO22X1_HVT U2941 ( .A1(\ram[11][83] ), .A2(n7448), .A3(n6808), .A4(data[83]), 
        .Y(n2960) );
  AO22X1_HVT U2942 ( .A1(\ram[11][84] ), .A2(n10169), .A3(n6819), .A4(data[84]), .Y(n2961) );
  AO22X1_HVT U2943 ( .A1(\ram[11][85] ), .A2(n7436), .A3(n4211), .A4(data[85]), 
        .Y(n2962) );
  AO22X1_HVT U2944 ( .A1(\ram[11][86] ), .A2(n10166), .A3(n6783), .A4(data[86]), .Y(n2963) );
  AO22X1_HVT U2945 ( .A1(\ram[11][87] ), .A2(n7436), .A3(n6776), .A4(data[87]), 
        .Y(n2964) );
  AO22X1_HVT U2946 ( .A1(\ram[11][88] ), .A2(n7465), .A3(n6797), .A4(data[88]), 
        .Y(n2965) );
  AO22X1_HVT U2947 ( .A1(\ram[11][89] ), .A2(n7434), .A3(n10158), .A4(data[89]), .Y(n2966) );
  AO22X1_HVT U2948 ( .A1(\ram[11][90] ), .A2(n7433), .A3(n6820), .A4(data[90]), 
        .Y(n2967) );
  AO22X1_HVT U2949 ( .A1(\ram[11][91] ), .A2(n7427), .A3(n6801), .A4(data[91]), 
        .Y(n2968) );
  AO22X1_HVT U2950 ( .A1(\ram[11][92] ), .A2(n7445), .A3(n6782), .A4(data[92]), 
        .Y(n2969) );
  AO22X1_HVT U2951 ( .A1(\ram[11][93] ), .A2(n7426), .A3(n6777), .A4(data[93]), 
        .Y(n2970) );
  AO22X1_HVT U2952 ( .A1(\ram[11][94] ), .A2(n7463), .A3(n6798), .A4(data[94]), 
        .Y(n2971) );
  AO22X1_HVT U2953 ( .A1(\ram[11][95] ), .A2(n7461), .A3(n6809), .A4(data[95]), 
        .Y(n2972) );
  AO22X1_HVT U2954 ( .A1(\ram[11][96] ), .A2(n7460), .A3(n10155), .A4(data[96]), .Y(n2973) );
  AO22X1_HVT U2955 ( .A1(\ram[11][97] ), .A2(n7458), .A3(n6770), .A4(data[97]), 
        .Y(n2974) );
  AO22X1_HVT U2956 ( .A1(\ram[11][98] ), .A2(n4314), .A3(n6771), .A4(data[98]), 
        .Y(n2975) );
  AO22X1_HVT U2957 ( .A1(\ram[11][99] ), .A2(n4314), .A3(n6779), .A4(data[99]), 
        .Y(n2976) );
  AO22X1_HVT U2958 ( .A1(\ram[11][100] ), .A2(n7434), .A3(n6799), .A4(
        data[100]), .Y(n2977) );
  AO22X1_HVT U2959 ( .A1(\ram[11][101] ), .A2(n7419), .A3(n6819), .A4(
        data[101]), .Y(n2978) );
  AO22X1_HVT U2960 ( .A1(\ram[11][102] ), .A2(n7474), .A3(n6819), .A4(
        data[102]), .Y(n2979) );
  AO22X1_HVT U2961 ( .A1(\ram[11][103] ), .A2(n7433), .A3(n4211), .A4(
        data[103]), .Y(n2980) );
  AO22X1_HVT U2962 ( .A1(\ram[11][104] ), .A2(n7427), .A3(n6772), .A4(
        data[104]), .Y(n2981) );
  AO22X1_HVT U2963 ( .A1(\ram[11][105] ), .A2(n7465), .A3(n6782), .A4(n9623), 
        .Y(n2982) );
  AO22X1_HVT U2964 ( .A1(\ram[11][106] ), .A2(n7426), .A3(n10157), .A4(
        data[106]), .Y(n2983) );
  AO22X1_HVT U2965 ( .A1(\ram[11][107] ), .A2(n7425), .A3(n6814), .A4(
        data[107]), .Y(n2984) );
  AO22X1_HVT U2966 ( .A1(\ram[11][108] ), .A2(n7423), .A3(n6820), .A4(
        data[108]), .Y(n2985) );
  AO22X1_HVT U2967 ( .A1(\ram[11][109] ), .A2(n7422), .A3(n6802), .A4(
        data[109]), .Y(n2986) );
  AO22X1_HVT U2968 ( .A1(\ram[11][110] ), .A2(n7420), .A3(n6773), .A4(
        data[110]), .Y(n2987) );
  AO22X1_HVT U2969 ( .A1(\ram[11][111] ), .A2(n7419), .A3(n6783), .A4(
        data[111]), .Y(n2988) );
  AO22X1_HVT U2970 ( .A1(\ram[11][112] ), .A2(n7474), .A3(n6806), .A4(
        data[112]), .Y(n2989) );
  AO22X1_HVT U2971 ( .A1(\ram[11][113] ), .A2(n7473), .A3(n6810), .A4(
        data[113]), .Y(n2990) );
  AO22X1_HVT U2972 ( .A1(\ram[11][114] ), .A2(n7472), .A3(n6820), .A4(
        data[114]), .Y(n2991) );
  AO22X1_HVT U2973 ( .A1(\ram[11][115] ), .A2(n7471), .A3(n6770), .A4(
        data[115]), .Y(n2992) );
  AO22X1_HVT U2974 ( .A1(\ram[11][116] ), .A2(n7470), .A3(n6774), .A4(
        data[116]), .Y(n2993) );
  AO22X1_HVT U2975 ( .A1(\ram[11][117] ), .A2(n7445), .A3(n6785), .A4(n9659), 
        .Y(n2994) );
  AO22X1_HVT U2976 ( .A1(\ram[11][118] ), .A2(n7465), .A3(n6780), .A4(n9662), 
        .Y(n2995) );
  AO22X1_HVT U2977 ( .A1(\ram[11][119] ), .A2(n7474), .A3(n6811), .A4(
        data[119]), .Y(n2996) );
  AO22X1_HVT U2978 ( .A1(\ram[11][120] ), .A2(n10166), .A3(n6787), .A4(n9668), 
        .Y(n2997) );
  AO22X1_HVT U2979 ( .A1(\ram[11][121] ), .A2(n7468), .A3(n10151), .A4(n9671), 
        .Y(n2998) );
  AO22X1_HVT U2980 ( .A1(\ram[11][122] ), .A2(n7447), .A3(n6810), .A4(n9674), 
        .Y(n2999) );
  AO22X1_HVT U2981 ( .A1(\ram[11][123] ), .A2(n4426), .A3(n6809), .A4(
        data[123]), .Y(n3000) );
  AO22X1_HVT U2982 ( .A1(\ram[11][124] ), .A2(n4314), .A3(n6789), .A4(
        data[124]), .Y(n3001) );
  AO22X1_HVT U2983 ( .A1(\ram[11][125] ), .A2(n7464), .A3(n10155), .A4(
        data[125]), .Y(n3002) );
  AO22X1_HVT U2984 ( .A1(\ram[11][126] ), .A2(n7463), .A3(n6788), .A4(
        data[126]), .Y(n3003) );
  AO22X1_HVT U2985 ( .A1(\ram[11][127] ), .A2(n7461), .A3(n6787), .A4(
        data[127]), .Y(n3004) );
  AO22X1_HVT U2986 ( .A1(\ram[11][128] ), .A2(n7460), .A3(n6773), .A4(
        data[128]), .Y(n3005) );
  AO22X1_HVT U2987 ( .A1(\ram[11][129] ), .A2(n7458), .A3(n10151), .A4(
        data[129]), .Y(n3006) );
  AO22X1_HVT U2988 ( .A1(\ram[11][130] ), .A2(n7457), .A3(n6825), .A4(
        data[130]), .Y(n3007) );
  AO22X1_HVT U2989 ( .A1(\ram[11][131] ), .A2(n7455), .A3(n6824), .A4(
        data[131]), .Y(n3008) );
  AO22X1_HVT U2990 ( .A1(\ram[11][132] ), .A2(n7454), .A3(n6811), .A4(
        data[132]), .Y(n3009) );
  AO22X1_HVT U2991 ( .A1(\ram[11][133] ), .A2(n7452), .A3(n6810), .A4(
        data[133]), .Y(n3010) );
  AO22X1_HVT U2992 ( .A1(\ram[11][134] ), .A2(n10166), .A3(n6798), .A4(
        data[134]), .Y(n3011) );
  AO22X1_HVT U2993 ( .A1(\ram[11][135] ), .A2(n7451), .A3(n6797), .A4(
        data[135]), .Y(n3012) );
  AO22X1_HVT U2994 ( .A1(\ram[11][136] ), .A2(n7450), .A3(n6796), .A4(
        data[136]), .Y(n3013) );
  AO22X1_HVT U2995 ( .A1(\ram[11][137] ), .A2(n7425), .A3(n6794), .A4(
        data[137]), .Y(n3014) );
  AO22X1_HVT U2996 ( .A1(\ram[11][138] ), .A2(n7422), .A3(n6793), .A4(
        data[138]), .Y(n3015) );
  AO22X1_HVT U2997 ( .A1(\ram[11][139] ), .A2(n7423), .A3(n6792), .A4(n9726), 
        .Y(n3016) );
  AO22X1_HVT U2998 ( .A1(\ram[11][140] ), .A2(n7420), .A3(n6791), .A4(
        data[140]), .Y(n3017) );
  AO22X1_HVT U2999 ( .A1(\ram[11][141] ), .A2(n7419), .A3(n6789), .A4(
        data[141]), .Y(n3018) );
  AO22X1_HVT U3000 ( .A1(\ram[11][142] ), .A2(n7474), .A3(n4211), .A4(n9735), 
        .Y(n3019) );
  AO22X1_HVT U3001 ( .A1(\ram[11][143] ), .A2(n7473), .A3(n6788), .A4(n9739), 
        .Y(n3020) );
  AO22X1_HVT U3002 ( .A1(\ram[11][144] ), .A2(n7472), .A3(n10153), .A4(
        data[144]), .Y(n3021) );
  AO22X1_HVT U3003 ( .A1(\ram[11][145] ), .A2(n7457), .A3(n10152), .A4(
        data[145]), .Y(n3022) );
  AO22X1_HVT U3004 ( .A1(\ram[11][146] ), .A2(n7455), .A3(n6786), .A4(
        data[146]), .Y(n3023) );
  AO22X1_HVT U3005 ( .A1(\ram[11][147] ), .A2(n7454), .A3(n6785), .A4(n9752), 
        .Y(n3024) );
  AO22X1_HVT U3006 ( .A1(\ram[11][148] ), .A2(n7452), .A3(n6783), .A4(
        data[148]), .Y(n3025) );
  AO22X1_HVT U3007 ( .A1(\ram[11][149] ), .A2(n7471), .A3(n6782), .A4(
        data[149]), .Y(n3026) );
  AO22X1_HVT U3008 ( .A1(\ram[11][150] ), .A2(n7438), .A3(n6780), .A4(
        data[150]), .Y(n3027) );
  AO22X1_HVT U3009 ( .A1(\ram[11][151] ), .A2(n7467), .A3(n6796), .A4(
        data[151]), .Y(n3028) );
  AO22X1_HVT U3010 ( .A1(\ram[11][152] ), .A2(n7473), .A3(n6794), .A4(
        data[152]), .Y(n3029) );
  AO22X1_HVT U3011 ( .A1(\ram[11][153] ), .A2(n7472), .A3(n6793), .A4(
        data[153]), .Y(n3030) );
  AO22X1_HVT U3012 ( .A1(\ram[11][154] ), .A2(n7431), .A3(n6792), .A4(
        data[154]), .Y(n3031) );
  AO22X1_HVT U3013 ( .A1(\ram[11][155] ), .A2(n7444), .A3(n6801), .A4(n9777), 
        .Y(n3032) );
  AO22X1_HVT U3014 ( .A1(\ram[11][156] ), .A2(n7443), .A3(n6794), .A4(
        data[156]), .Y(n3033) );
  AO22X1_HVT U3015 ( .A1(\ram[11][157] ), .A2(n7442), .A3(n6793), .A4(
        data[157]), .Y(n3034) );
  AO22X1_HVT U3016 ( .A1(\ram[11][158] ), .A2(n10174), .A3(n6792), .A4(
        data[158]), .Y(n3035) );
  AO22X1_HVT U3017 ( .A1(\ram[11][159] ), .A2(n10169), .A3(n6791), .A4(n9790), 
        .Y(n3036) );
  AO22X1_HVT U3018 ( .A1(\ram[11][160] ), .A2(n10174), .A3(n6789), .A4(
        data[160]), .Y(n3037) );
  AO22X1_HVT U3019 ( .A1(\ram[11][161] ), .A2(n7441), .A3(n10157), .A4(
        data[161]), .Y(n3038) );
  AO22X1_HVT U3020 ( .A1(\ram[11][162] ), .A2(n7440), .A3(n6788), .A4(
        data[162]), .Y(n3039) );
  AO22X1_HVT U3021 ( .A1(\ram[11][163] ), .A2(n7439), .A3(n10155), .A4(
        data[163]), .Y(n3040) );
  AO22X1_HVT U3022 ( .A1(\ram[11][164] ), .A2(n7438), .A3(n6817), .A4(
        data[164]), .Y(n3041) );
  AO22X1_HVT U3023 ( .A1(\ram[11][165] ), .A2(n10166), .A3(n10156), .A4(
        data[165]), .Y(n3042) );
  AO22X1_HVT U3024 ( .A1(\ram[11][166] ), .A2(n7436), .A3(n10152), .A4(
        data[166]), .Y(n3043) );
  AO22X1_HVT U3025 ( .A1(\ram[11][167] ), .A2(n7465), .A3(n6817), .A4(
        data[167]), .Y(n3044) );
  AO22X1_HVT U3026 ( .A1(\ram[11][168] ), .A2(n7434), .A3(n6811), .A4(
        data[168]), .Y(n3045) );
  AO22X1_HVT U3027 ( .A1(\ram[11][169] ), .A2(n7433), .A3(n6799), .A4(
        data[169]), .Y(n3046) );
  AO22X1_HVT U3028 ( .A1(\ram[11][170] ), .A2(n7427), .A3(n6798), .A4(
        data[170]), .Y(n3047) );
  AO22X1_HVT U3029 ( .A1(\ram[11][171] ), .A2(n7431), .A3(n6797), .A4(n9827), 
        .Y(n3048) );
  AO22X1_HVT U3030 ( .A1(\ram[11][172] ), .A2(n7426), .A3(n6796), .A4(n9830), 
        .Y(n3049) );
  AO22X1_HVT U3031 ( .A1(\ram[11][173] ), .A2(n7425), .A3(n6794), .A4(
        data[173]), .Y(n3050) );
  AO22X1_HVT U3032 ( .A1(\ram[11][174] ), .A2(n7423), .A3(n6793), .A4(
        data[174]), .Y(n3051) );
  AO22X1_HVT U3033 ( .A1(\ram[11][175] ), .A2(n7422), .A3(n6792), .A4(n9840), 
        .Y(n3052) );
  AO22X1_HVT U3034 ( .A1(\ram[11][176] ), .A2(n7420), .A3(n6791), .A4(n9843), 
        .Y(n3053) );
  AO22X1_HVT U3035 ( .A1(\ram[11][177] ), .A2(n7419), .A3(n6798), .A4(
        data[177]), .Y(n3054) );
  AO22X1_HVT U3036 ( .A1(\ram[11][178] ), .A2(n7474), .A3(n6797), .A4(
        data[178]), .Y(n3055) );
  AO22X1_HVT U3037 ( .A1(\ram[11][179] ), .A2(n7473), .A3(n6796), .A4(n9853), 
        .Y(n3056) );
  AO22X1_HVT U3038 ( .A1(\ram[11][180] ), .A2(n7472), .A3(n6779), .A4(
        data[180]), .Y(n3057) );
  AO22X1_HVT U3039 ( .A1(\ram[11][181] ), .A2(n7471), .A3(n6777), .A4(n9859), 
        .Y(n3058) );
  AO22X1_HVT U3040 ( .A1(\ram[11][182] ), .A2(n7470), .A3(n6776), .A4(
        data[182]), .Y(n3059) );
  AO22X1_HVT U3041 ( .A1(\ram[11][183] ), .A2(n4431), .A3(n6774), .A4(n9866), 
        .Y(n3060) );
  AO22X1_HVT U3042 ( .A1(\ram[11][184] ), .A2(n7435), .A3(n6773), .A4(
        data[184]), .Y(n3061) );
  AO22X1_HVT U3043 ( .A1(\ram[11][185] ), .A2(n7473), .A3(n6772), .A4(
        data[185]), .Y(n3062) );
  AO22X1_HVT U3044 ( .A1(\ram[11][186] ), .A2(n10165), .A3(n6771), .A4(
        data[186]), .Y(n3063) );
  AO22X1_HVT U3045 ( .A1(\ram[11][187] ), .A2(n7468), .A3(n6770), .A4(
        data[187]), .Y(n3064) );
  AO22X1_HVT U3046 ( .A1(\ram[11][188] ), .A2(n7471), .A3(n10157), .A4(
        data[188]), .Y(n3065) );
  AO22X1_HVT U3047 ( .A1(\ram[11][189] ), .A2(n7470), .A3(n6802), .A4(
        data[189]), .Y(n3066) );
  AO22X1_HVT U3048 ( .A1(\ram[11][190] ), .A2(n4431), .A3(n6799), .A4(
        data[190]), .Y(n3067) );
  AO22X1_HVT U3049 ( .A1(\ram[11][191] ), .A2(n7430), .A3(n6813), .A4(n9891), 
        .Y(n3068) );
  AO22X1_HVT U3050 ( .A1(\ram[11][192] ), .A2(n7472), .A3(n6788), .A4(
        data[192]), .Y(n3069) );
  AO22X1_HVT U3051 ( .A1(\ram[11][193] ), .A2(n10169), .A3(n6787), .A4(
        data[193]), .Y(n3070) );
  AO22X1_HVT U3052 ( .A1(\ram[11][194] ), .A2(n7468), .A3(n6772), .A4(
        data[194]), .Y(n3071) );
  AO22X1_HVT U3053 ( .A1(\ram[11][195] ), .A2(n7467), .A3(n10157), .A4(n9904), 
        .Y(n3072) );
  AO22X1_HVT U3054 ( .A1(\ram[11][196] ), .A2(n10168), .A3(n6824), .A4(
        data[196]), .Y(n3073) );
  AO22X1_HVT U3055 ( .A1(\ram[11][197] ), .A2(n7451), .A3(n6823), .A4(
        data[197]), .Y(n3074) );
  AO22X1_HVT U3056 ( .A1(\ram[11][198] ), .A2(n7450), .A3(n6822), .A4(
        data[198]), .Y(n3075) );
  AO22X1_HVT U3057 ( .A1(\ram[11][199] ), .A2(n7448), .A3(n6821), .A4(n9917), 
        .Y(n3076) );
  AO22X1_HVT U3058 ( .A1(\ram[11][200] ), .A2(n7435), .A3(n6798), .A4(
        data[200]), .Y(n3077) );
  AO22X1_HVT U3059 ( .A1(\ram[11][201] ), .A2(n7467), .A3(n6806), .A4(n9923), 
        .Y(n3078) );
  AO22X1_HVT U3060 ( .A1(\ram[11][202] ), .A2(n4426), .A3(n6805), .A4(
        data[202]), .Y(n3079) );
  AO22X1_HVT U3061 ( .A1(\ram[11][203] ), .A2(n7471), .A3(n6785), .A4(
        data[203]), .Y(n3080) );
  AO22X1_HVT U3062 ( .A1(\ram[11][204] ), .A2(n7470), .A3(n6785), .A4(
        data[204]), .Y(n3081) );
  AO22X1_HVT U3063 ( .A1(\ram[11][205] ), .A2(n7430), .A3(n6783), .A4(
        data[205]), .Y(n3082) );
  AO22X1_HVT U3064 ( .A1(\ram[11][206] ), .A2(n7464), .A3(n6782), .A4(
        data[206]), .Y(n3083) );
  AO22X1_HVT U3065 ( .A1(\ram[11][207] ), .A2(n7463), .A3(n6780), .A4(n9942), 
        .Y(n3084) );
  AO22X1_HVT U3066 ( .A1(\ram[11][208] ), .A2(n7461), .A3(n6774), .A4(
        data[208]), .Y(n3085) );
  AO22X1_HVT U3067 ( .A1(\ram[11][209] ), .A2(n7460), .A3(n6773), .A4(
        data[209]), .Y(n3086) );
  AO22X1_HVT U3068 ( .A1(\ram[11][210] ), .A2(n7458), .A3(n6772), .A4(
        data[210]), .Y(n3087) );
  AO22X1_HVT U3069 ( .A1(\ram[11][211] ), .A2(n7457), .A3(n6771), .A4(
        data[211]), .Y(n3088) );
  AO22X1_HVT U3070 ( .A1(\ram[11][212] ), .A2(n7455), .A3(n6792), .A4(
        data[212]), .Y(n3089) );
  AO22X1_HVT U3071 ( .A1(\ram[11][213] ), .A2(n7454), .A3(n6791), .A4(n9960), 
        .Y(n3090) );
  AO22X1_HVT U3072 ( .A1(\ram[11][214] ), .A2(n7452), .A3(n6789), .A4(
        data[214]), .Y(n3091) );
  AO22X1_HVT U3073 ( .A1(\ram[11][215] ), .A2(n7420), .A3(n10156), .A4(
        data[215]), .Y(n3092) );
  AO22X1_HVT U3074 ( .A1(\ram[11][216] ), .A2(n7451), .A3(n6809), .A4(
        data[216]), .Y(n3093) );
  AO22X1_HVT U3075 ( .A1(\ram[11][217] ), .A2(n7450), .A3(n10160), .A4(
        data[217]), .Y(n3094) );
  AO22X1_HVT U3076 ( .A1(\ram[11][218] ), .A2(n7448), .A3(n6808), .A4(
        data[218]), .Y(n3095) );
  AO22X1_HVT U3077 ( .A1(\ram[11][219] ), .A2(n7447), .A3(n10154), .A4(n9979), 
        .Y(n3096) );
  AO22X1_HVT U3078 ( .A1(\ram[11][220] ), .A2(n7466), .A3(n6806), .A4(
        data[220]), .Y(n3097) );
  AO22X1_HVT U3079 ( .A1(\ram[11][221] ), .A2(n7444), .A3(n6805), .A4(
        data[221]), .Y(n3098) );
  AO22X1_HVT U3080 ( .A1(\ram[11][222] ), .A2(n7443), .A3(n6805), .A4(
        data[222]), .Y(n3099) );
  AO22X1_HVT U3081 ( .A1(\ram[11][223] ), .A2(n7442), .A3(n10155), .A4(
        data[223]), .Y(n3100) );
  AO22X1_HVT U3082 ( .A1(\ram[11][224] ), .A2(n10173), .A3(n6817), .A4(
        data[224]), .Y(n3101) );
  AO22X1_HVT U3083 ( .A1(\ram[11][225] ), .A2(n10168), .A3(n6811), .A4(
        data[225]), .Y(n3102) );
  AO22X1_HVT U3084 ( .A1(\ram[11][226] ), .A2(n10165), .A3(n10152), .A4(
        data[226]), .Y(n3103) );
  AO22X1_HVT U3085 ( .A1(\ram[11][227] ), .A2(n7441), .A3(n6786), .A4(
        data[227]), .Y(n3104) );
  AO22X1_HVT U3086 ( .A1(\ram[11][228] ), .A2(n7440), .A3(n10152), .A4(n10006), 
        .Y(n3105) );
  AO22X1_HVT U3087 ( .A1(\ram[11][229] ), .A2(n7439), .A3(n6806), .A4(
        data[229]), .Y(n3106) );
  AO22X1_HVT U3088 ( .A1(\ram[11][230] ), .A2(n7438), .A3(n6805), .A4(
        data[230]), .Y(n3107) );
  AO22X1_HVT U3089 ( .A1(\ram[11][231] ), .A2(n10166), .A3(n10154), .A4(n10016), .Y(n3108) );
  AO22X1_HVT U3090 ( .A1(\ram[11][232] ), .A2(n7436), .A3(n6817), .A4(
        data[232]), .Y(n3109) );
  AO22X1_HVT U3091 ( .A1(\ram[11][233] ), .A2(n7430), .A3(n6787), .A4(
        data[233]), .Y(n3110) );
  AO22X1_HVT U3092 ( .A1(\ram[11][234] ), .A2(n7434), .A3(n10150), .A4(
        data[234]), .Y(n3111) );
  AO22X1_HVT U3093 ( .A1(\ram[11][235] ), .A2(n7433), .A3(n6786), .A4(
        data[235]), .Y(n3112) );
  AO22X1_HVT U3094 ( .A1(\ram[11][236] ), .A2(n7427), .A3(n10152), .A4(n10031), 
        .Y(n3113) );
  AO22X1_HVT U3095 ( .A1(\ram[11][237] ), .A2(n7445), .A3(n6806), .A4(
        data[237]), .Y(n3114) );
  AO22X1_HVT U3096 ( .A1(\ram[11][238] ), .A2(n7426), .A3(n6811), .A4(
        data[238]), .Y(n3115) );
  AO22X1_HVT U3097 ( .A1(\ram[11][239] ), .A2(n7445), .A3(n6810), .A4(n10041), 
        .Y(n3116) );
  AO22X1_HVT U3098 ( .A1(\ram[11][240] ), .A2(n7435), .A3(n6793), .A4(
        data[240]), .Y(n3117) );
  AO22X1_HVT U3099 ( .A1(\ram[11][241] ), .A2(n7464), .A3(n6787), .A4(
        data[241]), .Y(n3118) );
  AO22X1_HVT U3100 ( .A1(\ram[11][242] ), .A2(n7463), .A3(n6774), .A4(
        data[242]), .Y(n3119) );
  AO22X1_HVT U3101 ( .A1(\ram[11][243] ), .A2(n7461), .A3(n6801), .A4(
        data[243]), .Y(n3120) );
  AO22X1_HVT U3102 ( .A1(\ram[11][244] ), .A2(n7460), .A3(n6825), .A4(n10056), 
        .Y(n3121) );
  AO22X1_HVT U3103 ( .A1(\ram[11][245] ), .A2(n7458), .A3(n6799), .A4(
        data[245]), .Y(n3122) );
  AO22X1_HVT U3104 ( .A1(\ram[11][246] ), .A2(n7457), .A3(n6808), .A4(
        data[246]), .Y(n3123) );
  AO22X1_HVT U3105 ( .A1(\ram[11][247] ), .A2(n7447), .A3(n10153), .A4(n10066), 
        .Y(n3124) );
  AO22X1_HVT U3106 ( .A1(\ram[11][248] ), .A2(n7431), .A3(n6810), .A4(
        data[248]), .Y(n3125) );
  AO22X1_HVT U3107 ( .A1(\ram[11][249] ), .A2(n7444), .A3(n6809), .A4(
        data[249]), .Y(n3126) );
  AO22X1_HVT U3108 ( .A1(\ram[11][250] ), .A2(n7443), .A3(n10160), .A4(
        data[250]), .Y(n3127) );
  AO22X1_HVT U3109 ( .A1(\ram[11][251] ), .A2(n7468), .A3(n6808), .A4(n10079), 
        .Y(n3128) );
  AO22X1_HVT U3110 ( .A1(\ram[11][252] ), .A2(n7470), .A3(n6770), .A4(
        data[252]), .Y(n3129) );
  AO22X1_HVT U3111 ( .A1(\ram[11][253] ), .A2(n7455), .A3(n6814), .A4(n10085), 
        .Y(n3130) );
  AO22X1_HVT U3112 ( .A1(\ram[11][254] ), .A2(n7454), .A3(n6813), .A4(
        data[254]), .Y(n3131) );
  AO22X1_HVT U3113 ( .A1(\ram[11][255] ), .A2(n7425), .A3(n6780), .A4(n10092), 
        .Y(n3132) );
  AND2X1_HVT U3116 ( .A1(n38), .A2(n6013), .Y(n47) );
  AO22X1_HVT U3118 ( .A1(\ram[12][0] ), .A2(n6588), .A3(n6378), .A4(n9307), 
        .Y(n3133) );
  AO22X1_HVT U3119 ( .A1(\ram[12][1] ), .A2(n6592), .A3(n4552), .A4(data[1]), 
        .Y(n3134) );
  AO22X1_HVT U3120 ( .A1(\ram[12][2] ), .A2(n6591), .A3(n4550), .A4(n9313), 
        .Y(n3135) );
  AO22X1_HVT U3121 ( .A1(\ram[12][3] ), .A2(n6590), .A3(n4550), .A4(n9317), 
        .Y(n3136) );
  AO22X1_HVT U3122 ( .A1(\ram[12][4] ), .A2(n10135), .A3(n6377), .A4(n9320), 
        .Y(n3137) );
  AO22X1_HVT U3123 ( .A1(\ram[12][5] ), .A2(n6588), .A3(n4409), .A4(n9323), 
        .Y(n3138) );
  AO22X1_HVT U3124 ( .A1(\ram[12][6] ), .A2(n6587), .A3(n4409), .A4(n9326), 
        .Y(n3139) );
  AO22X1_HVT U3125 ( .A1(\ram[12][7] ), .A2(n6584), .A3(n4409), .A4(n9329), 
        .Y(n3140) );
  AO22X1_HVT U3126 ( .A1(\ram[12][8] ), .A2(n6583), .A3(n4411), .A4(n9331), 
        .Y(n3141) );
  AO22X1_HVT U3127 ( .A1(\ram[12][9] ), .A2(n6580), .A3(n6370), .A4(data[9]), 
        .Y(n3142) );
  AO22X1_HVT U3128 ( .A1(\ram[12][10] ), .A2(n6579), .A3(n6372), .A4(n9338), 
        .Y(n3143) );
  AO22X1_HVT U3129 ( .A1(\ram[12][11] ), .A2(n6610), .A3(n4552), .A4(n9342), 
        .Y(n3144) );
  AO22X1_HVT U3130 ( .A1(\ram[12][12] ), .A2(n6621), .A3(n4557), .A4(n9345), 
        .Y(n3145) );
  AO22X1_HVT U3131 ( .A1(\ram[12][13] ), .A2(n6620), .A3(n4552), .A4(n9348), 
        .Y(n3146) );
  AO22X1_HVT U3133 ( .A1(\ram[12][15] ), .A2(n6618), .A3(n6371), .A4(n9354), 
        .Y(n3148) );
  AO22X1_HVT U3134 ( .A1(\ram[12][16] ), .A2(n6616), .A3(n6371), .A4(data[16]), 
        .Y(n3149) );
  AO22X1_HVT U3135 ( .A1(\ram[12][17] ), .A2(n6615), .A3(n6375), .A4(n9360), 
        .Y(n3150) );
  AO22X1_HVT U3136 ( .A1(\ram[12][18] ), .A2(n6613), .A3(n6372), .A4(n9362), 
        .Y(n3151) );
  AO22X1_HVT U3137 ( .A1(\ram[12][19] ), .A2(n6613), .A3(n4552), .A4(n9366), 
        .Y(n3152) );
  AO22X1_HVT U3138 ( .A1(\ram[12][20] ), .A2(n6612), .A3(n6370), .A4(data[20]), 
        .Y(n3153) );
  AO22X1_HVT U3139 ( .A1(\ram[12][21] ), .A2(n6610), .A3(n4411), .A4(data[21]), 
        .Y(n3154) );
  AO22X1_HVT U3140 ( .A1(\ram[12][22] ), .A2(n6609), .A3(n6366), .A4(data[22]), 
        .Y(n3155) );
  AO22X1_HVT U3141 ( .A1(\ram[12][23] ), .A2(n6606), .A3(n6367), .A4(n9377), 
        .Y(n3156) );
  AO22X1_HVT U3142 ( .A1(\ram[12][24] ), .A2(n6557), .A3(n6367), .A4(n9380), 
        .Y(n3157) );
  AO22X1_HVT U3143 ( .A1(\ram[12][25] ), .A2(n6556), .A3(n6367), .A4(n9382), 
        .Y(n3158) );
  AO22X1_HVT U3144 ( .A1(\ram[12][26] ), .A2(n6587), .A3(n4551), .A4(data[26]), 
        .Y(n3159) );
  AO22X1_HVT U3145 ( .A1(\ram[12][27] ), .A2(n6584), .A3(n6366), .A4(data[27]), 
        .Y(n3160) );
  AO22X1_HVT U3147 ( .A1(\ram[12][29] ), .A2(n6602), .A3(n6334), .A4(n9394), 
        .Y(n3162) );
  AO22X1_HVT U3148 ( .A1(\ram[12][30] ), .A2(n6612), .A3(n6342), .A4(n9398), 
        .Y(n3163) );
  AO22X1_HVT U3149 ( .A1(\ram[12][31] ), .A2(n6601), .A3(n6333), .A4(n9401), 
        .Y(n3164) );
  AO22X1_HVT U3151 ( .A1(\ram[12][33] ), .A2(n6591), .A3(n4744), .A4(n9407), 
        .Y(n3166) );
  AO22X1_HVT U3154 ( .A1(\ram[12][36] ), .A2(n6605), .A3(n4549), .A4(data[36]), 
        .Y(n3169) );
  AO22X1_HVT U3155 ( .A1(\ram[12][37] ), .A2(n6602), .A3(n6377), .A4(n9419), 
        .Y(n3170) );
  AO22X1_HVT U3156 ( .A1(\ram[12][38] ), .A2(n6601), .A3(n6376), .A4(data[38]), 
        .Y(n3171) );
  AO22X1_HVT U3157 ( .A1(\ram[12][39] ), .A2(n6559), .A3(n4707), .A4(n9425), 
        .Y(n3172) );
  AO22X1_HVT U3158 ( .A1(\ram[12][40] ), .A2(n6558), .A3(n6344), .A4(n9428), 
        .Y(n3173) );
  AO22X1_HVT U3159 ( .A1(\ram[12][41] ), .A2(n6572), .A3(n6343), .A4(data[41]), 
        .Y(n3174) );
  AO22X1_HVT U3160 ( .A1(\ram[12][42] ), .A2(n6571), .A3(n4707), .A4(n9433), 
        .Y(n3175) );
  AO22X1_HVT U3161 ( .A1(\ram[12][43] ), .A2(n6624), .A3(n4557), .A4(n9437), 
        .Y(n3176) );
  AO22X1_HVT U3162 ( .A1(\ram[12][44] ), .A2(n6622), .A3(n6378), .A4(n9440), 
        .Y(n3177) );
  AO22X1_HVT U3163 ( .A1(\ram[12][45] ), .A2(n4268), .A3(n4549), .A4(n9443), 
        .Y(n3178) );
  AO22X1_HVT U3164 ( .A1(\ram[12][46] ), .A2(n6621), .A3(n6380), .A4(data[46]), 
        .Y(n3179) );
  AO22X1_HVT U3165 ( .A1(\ram[12][47] ), .A2(n6598), .A3(n6379), .A4(n9449), 
        .Y(n3180) );
  AO22X1_HVT U3166 ( .A1(\ram[12][48] ), .A2(n6577), .A3(n6332), .A4(data[48]), 
        .Y(n3181) );
  AO22X1_HVT U3168 ( .A1(\ram[12][50] ), .A2(n4357), .A3(n4559), .A4(data[50]), 
        .Y(n3183) );
  AO22X1_HVT U3169 ( .A1(\ram[12][51] ), .A2(n6577), .A3(n6351), .A4(n9460), 
        .Y(n3184) );
  AO22X1_HVT U3170 ( .A1(\ram[12][52] ), .A2(n6576), .A3(n6376), .A4(n9464), 
        .Y(n3185) );
  AO22X1_HVT U3171 ( .A1(\ram[12][53] ), .A2(n6606), .A3(n4354), .A4(n9466), 
        .Y(n3186) );
  AO22X1_HVT U3172 ( .A1(\ram[12][54] ), .A2(n6572), .A3(n6338), .A4(data[54]), 
        .Y(n3187) );
  AO22X1_HVT U3173 ( .A1(\ram[12][55] ), .A2(n6571), .A3(n6335), .A4(data[55]), 
        .Y(n3188) );
  AO22X1_HVT U3174 ( .A1(\ram[12][56] ), .A2(n6570), .A3(n4406), .A4(data[56]), 
        .Y(n3189) );
  AO22X1_HVT U3175 ( .A1(\ram[12][57] ), .A2(n6568), .A3(n6337), .A4(data[57]), 
        .Y(n3190) );
  AO22X1_HVT U3176 ( .A1(\ram[12][58] ), .A2(n4360), .A3(n4406), .A4(data[58]), 
        .Y(n3191) );
  AO22X1_HVT U3177 ( .A1(\ram[12][59] ), .A2(n6617), .A3(n6343), .A4(n9485), 
        .Y(n3192) );
  AO22X1_HVT U3178 ( .A1(\ram[12][60] ), .A2(n6618), .A3(n6375), .A4(n9488), 
        .Y(n3193) );
  AO22X1_HVT U3179 ( .A1(\ram[12][61] ), .A2(n6616), .A3(n6370), .A4(n9491), 
        .Y(n3194) );
  AO22X1_HVT U3180 ( .A1(\ram[12][62] ), .A2(n6597), .A3(n6372), .A4(n9494), 
        .Y(n3195) );
  AO22X1_HVT U3181 ( .A1(\ram[12][63] ), .A2(n6562), .A3(n4549), .A4(n9497), 
        .Y(n3196) );
  AO22X1_HVT U3182 ( .A1(\ram[12][64] ), .A2(n6561), .A3(n4409), .A4(data[64]), 
        .Y(n3197) );
  AO22X1_HVT U3183 ( .A1(\ram[12][65] ), .A2(n6583), .A3(n6368), .A4(data[65]), 
        .Y(n3198) );
  AO22X1_HVT U3184 ( .A1(\ram[12][66] ), .A2(n6580), .A3(n6366), .A4(n9506), 
        .Y(n3199) );
  AO22X1_HVT U3185 ( .A1(\ram[12][67] ), .A2(n6587), .A3(n4462), .A4(data[67]), 
        .Y(n3200) );
  AO22X1_HVT U3186 ( .A1(\ram[12][68] ), .A2(n6584), .A3(n4551), .A4(n9512), 
        .Y(n3201) );
  AO22X1_HVT U3188 ( .A1(\ram[12][70] ), .A2(n6580), .A3(n4708), .A4(n9518), 
        .Y(n3203) );
  AO22X1_HVT U3189 ( .A1(\ram[12][71] ), .A2(n6579), .A3(n4707), .A4(data[71]), 
        .Y(n3204) );
  AO22X1_HVT U3190 ( .A1(\ram[12][72] ), .A2(n6565), .A3(n6366), .A4(n9523), 
        .Y(n3205) );
  AO22X1_HVT U3191 ( .A1(\ram[12][73] ), .A2(n6587), .A3(n4411), .A4(n9527), 
        .Y(n3206) );
  AO22X1_HVT U3192 ( .A1(\ram[12][74] ), .A2(n6584), .A3(n6370), .A4(n9530), 
        .Y(n3207) );
  AO22X1_HVT U3193 ( .A1(\ram[12][75] ), .A2(n6583), .A3(n4409), .A4(data[75]), 
        .Y(n3208) );
  AO22X1_HVT U3194 ( .A1(\ram[12][76] ), .A2(n6580), .A3(n6348), .A4(n9536), 
        .Y(n3209) );
  AO22X1_HVT U3195 ( .A1(\ram[12][77] ), .A2(n6579), .A3(n6338), .A4(data[77]), 
        .Y(n3210) );
  AO22X1_HVT U3196 ( .A1(\ram[12][78] ), .A2(n6577), .A3(n6353), .A4(n9542), 
        .Y(n3211) );
  AO22X1_HVT U3197 ( .A1(\ram[12][79] ), .A2(n6576), .A3(n6335), .A4(data[79]), 
        .Y(n3212) );
  AO22X1_HVT U3198 ( .A1(\ram[12][80] ), .A2(n6619), .A3(n6369), .A4(data[80]), 
        .Y(n3213) );
  AO22X1_HVT U3199 ( .A1(\ram[12][81] ), .A2(n6572), .A3(n6346), .A4(data[81]), 
        .Y(n3214) );
  AO22X1_HVT U3200 ( .A1(\ram[12][82] ), .A2(n6571), .A3(n6348), .A4(data[82]), 
        .Y(n3215) );
  AO22X1_HVT U3202 ( .A1(\ram[12][84] ), .A2(n6609), .A3(n6367), .A4(n9560), 
        .Y(n3217) );
  AO22X1_HVT U3204 ( .A1(\ram[12][86] ), .A2(n6605), .A3(n6379), .A4(n9566), 
        .Y(n3219) );
  AO22X1_HVT U3205 ( .A1(\ram[12][87] ), .A2(n6602), .A3(n6346), .A4(data[87]), 
        .Y(n3220) );
  AO22X1_HVT U3206 ( .A1(\ram[12][88] ), .A2(n6601), .A3(n6377), .A4(data[88]), 
        .Y(n3221) );
  AO22X1_HVT U3207 ( .A1(\ram[12][89] ), .A2(n6592), .A3(n6369), .A4(n9575), 
        .Y(n3222) );
  AO22X1_HVT U3208 ( .A1(\ram[12][90] ), .A2(n6591), .A3(n6361), .A4(n9578), 
        .Y(n3223) );
  AO22X1_HVT U3209 ( .A1(\ram[12][91] ), .A2(n6590), .A3(n6359), .A4(n9581), 
        .Y(n3224) );
  AO22X1_HVT U3210 ( .A1(\ram[12][92] ), .A2(n6613), .A3(n4686), .A4(data[92]), 
        .Y(n3225) );
  AO22X1_HVT U3211 ( .A1(\ram[12][93] ), .A2(n6588), .A3(n6380), .A4(n9587), 
        .Y(n3226) );
  AO22X1_HVT U3212 ( .A1(\ram[12][94] ), .A2(n6592), .A3(n6347), .A4(data[94]), 
        .Y(n3227) );
  AO22X1_HVT U3213 ( .A1(\ram[12][95] ), .A2(n6591), .A3(n4744), .A4(data[95]), 
        .Y(n3228) );
  AO22X1_HVT U3214 ( .A1(\ram[12][96] ), .A2(n6590), .A3(n6339), .A4(data[96]), 
        .Y(n3229) );
  AO22X1_HVT U3215 ( .A1(\ram[12][97] ), .A2(n6580), .A3(n6341), .A4(n9599), 
        .Y(n3230) );
  AO22X1_HVT U3217 ( .A1(\ram[12][99] ), .A2(n6587), .A3(n6380), .A4(data[99]), 
        .Y(n3232) );
  AO22X1_HVT U3218 ( .A1(\ram[12][100] ), .A2(n6584), .A3(n6341), .A4(n9608), 
        .Y(n3233) );
  AO22X1_HVT U3219 ( .A1(\ram[12][101] ), .A2(n6583), .A3(n6368), .A4(n9611), 
        .Y(n3234) );
  AO22X1_HVT U3220 ( .A1(\ram[12][102] ), .A2(n6598), .A3(n6339), .A4(
        data[102]), .Y(n3235) );
  AO22X1_HVT U3221 ( .A1(\ram[12][103] ), .A2(n6597), .A3(n6334), .A4(n9617), 
        .Y(n3236) );
  AO22X1_HVT U3222 ( .A1(\ram[12][104] ), .A2(n6570), .A3(n6378), .A4(n9620), 
        .Y(n3237) );
  AO22X1_HVT U3223 ( .A1(\ram[12][105] ), .A2(n6568), .A3(n4462), .A4(
        data[105]), .Y(n3238) );
  AO22X1_HVT U3224 ( .A1(\ram[12][106] ), .A2(n6620), .A3(n6346), .A4(n9626), 
        .Y(n3239) );
  AO22X1_HVT U3225 ( .A1(\ram[12][107] ), .A2(n4357), .A3(n6376), .A4(n9629), 
        .Y(n3240) );
  AO22X1_HVT U3226 ( .A1(\ram[12][108] ), .A2(n6568), .A3(n6369), .A4(
        data[108]), .Y(n3241) );
  AO22X1_HVT U3227 ( .A1(\ram[12][109] ), .A2(n6580), .A3(n6357), .A4(n9635), 
        .Y(n3242) );
  AO22X1_HVT U3228 ( .A1(\ram[12][110] ), .A2(n6579), .A3(n6346), .A4(n9638), 
        .Y(n3243) );
  AO22X1_HVT U3229 ( .A1(\ram[12][111] ), .A2(n6577), .A3(n6363), .A4(n9641), 
        .Y(n3244) );
  AO22X1_HVT U3230 ( .A1(\ram[12][112] ), .A2(n6576), .A3(n4549), .A4(n9644), 
        .Y(n3245) );
  AO22X1_HVT U3231 ( .A1(\ram[12][113] ), .A2(n6573), .A3(n4309), .A4(n9647), 
        .Y(n3246) );
  AO22X1_HVT U3232 ( .A1(\ram[12][114] ), .A2(n6572), .A3(n6352), .A4(n9650), 
        .Y(n3247) );
  AO22X1_HVT U3233 ( .A1(\ram[12][115] ), .A2(n6571), .A3(n6355), .A4(n9653), 
        .Y(n3248) );
  AO22X1_HVT U3234 ( .A1(\ram[12][116] ), .A2(n6570), .A3(n6332), .A4(
        data[116]), .Y(n3249) );
  AO22X1_HVT U3235 ( .A1(\ram[12][117] ), .A2(n6625), .A3(n6379), .A4(n9659), 
        .Y(n3250) );
  AO22X1_HVT U3236 ( .A1(\ram[12][118] ), .A2(n6624), .A3(n6334), .A4(
        data[118]), .Y(n3251) );
  AO22X1_HVT U3237 ( .A1(\ram[12][119] ), .A2(n6567), .A3(n6337), .A4(n9665), 
        .Y(n3252) );
  AO22X1_HVT U3238 ( .A1(\ram[12][120] ), .A2(n6566), .A3(n6357), .A4(n9667), 
        .Y(n3253) );
  AO22X1_HVT U3239 ( .A1(\ram[12][121] ), .A2(n6615), .A3(n4557), .A4(n9670), 
        .Y(n3254) );
  AO22X1_HVT U3240 ( .A1(\ram[12][122] ), .A2(n6613), .A3(n6343), .A4(n9673), 
        .Y(n3255) );
  AO22X1_HVT U3241 ( .A1(\ram[12][123] ), .A2(n6612), .A3(n6357), .A4(
        data[123]), .Y(n3256) );
  AO22X1_HVT U3242 ( .A1(\ram[12][124] ), .A2(n6610), .A3(n4551), .A4(
        data[124]), .Y(n3257) );
  AO22X1_HVT U3243 ( .A1(\ram[12][125] ), .A2(n6562), .A3(n4619), .A4(
        data[125]), .Y(n3258) );
  AO22X1_HVT U3244 ( .A1(\ram[12][126] ), .A2(n6622), .A3(n6335), .A4(n9686), 
        .Y(n3259) );
  AO22X1_HVT U3245 ( .A1(\ram[12][127] ), .A2(n10142), .A3(n4406), .A4(
        data[127]), .Y(n3260) );
  AO22X1_HVT U3246 ( .A1(\ram[12][128] ), .A2(n6579), .A3(n4551), .A4(n9692), 
        .Y(n3261) );
  AO22X1_HVT U3247 ( .A1(\ram[12][129] ), .A2(n6577), .A3(n6366), .A4(n9695), 
        .Y(n3262) );
  AO22X1_HVT U3248 ( .A1(\ram[12][130] ), .A2(n6572), .A3(n4309), .A4(
        data[130]), .Y(n3263) );
  AO22X1_HVT U3249 ( .A1(\ram[12][131] ), .A2(n6571), .A3(n6350), .A4(n9701), 
        .Y(n3264) );
  AO22X1_HVT U3250 ( .A1(\ram[12][132] ), .A2(n6570), .A3(n6348), .A4(
        data[132]), .Y(n3265) );
  AO22X1_HVT U3251 ( .A1(\ram[12][133] ), .A2(n6568), .A3(n4862), .A4(
        data[133]), .Y(n3266) );
  AO22X1_HVT U3252 ( .A1(\ram[12][134] ), .A2(n4360), .A3(n4413), .A4(
        data[134]), .Y(n3267) );
  AO22X1_HVT U3253 ( .A1(\ram[12][135] ), .A2(n6566), .A3(n6359), .A4(n9713), 
        .Y(n3268) );
  AO22X1_HVT U3254 ( .A1(\ram[12][136] ), .A2(n6565), .A3(n6372), .A4(
        data[136]), .Y(n3269) );
  AO22X1_HVT U3255 ( .A1(\ram[12][137] ), .A2(n10146), .A3(n4411), .A4(
        data[137]), .Y(n3270) );
  AO22X1_HVT U3256 ( .A1(\ram[12][138] ), .A2(n10146), .A3(n6334), .A4(
        data[138]), .Y(n3271) );
  AO22X1_HVT U3257 ( .A1(\ram[12][139] ), .A2(n6617), .A3(n4310), .A4(n9726), 
        .Y(n3272) );
  AO22X1_HVT U3259 ( .A1(\ram[12][141] ), .A2(n6595), .A3(n6362), .A4(n9732), 
        .Y(n3274) );
  AO22X1_HVT U3262 ( .A1(\ram[12][144] ), .A2(n6558), .A3(n6337), .A4(
        data[144]), .Y(n3277) );
  AO22X1_HVT U3263 ( .A1(\ram[12][145] ), .A2(n6557), .A3(n6369), .A4(
        data[145]), .Y(n3278) );
  AO22X1_HVT U3264 ( .A1(\ram[12][146] ), .A2(n6556), .A3(n4744), .A4(n9748), 
        .Y(n3279) );
  AO22X1_HVT U3265 ( .A1(\ram[12][147] ), .A2(n6598), .A3(n6363), .A4(n9752), 
        .Y(n3280) );
  AO22X1_HVT U3266 ( .A1(\ram[12][148] ), .A2(n6596), .A3(n6341), .A4(
        data[148]), .Y(n3281) );
  AO22X1_HVT U3267 ( .A1(\ram[12][149] ), .A2(n4346), .A3(n6334), .A4(n9758), 
        .Y(n3282) );
  AO22X1_HVT U3268 ( .A1(\ram[12][150] ), .A2(n6565), .A3(n4552), .A4(n9761), 
        .Y(n3283) );
  AO22X1_HVT U3269 ( .A1(\ram[12][151] ), .A2(n10146), .A3(n6359), .A4(
        data[151]), .Y(n3284) );
  AO22X1_HVT U3270 ( .A1(\ram[12][152] ), .A2(n6566), .A3(n4685), .A4(
        data[152]), .Y(n3285) );
  AO22X1_HVT U3271 ( .A1(\ram[12][153] ), .A2(n6596), .A3(n4310), .A4(
        data[153]), .Y(n3286) );
  AO22X1_HVT U3272 ( .A1(\ram[12][154] ), .A2(n6595), .A3(n6355), .A4(n9773), 
        .Y(n3287) );
  AO22X1_HVT U3273 ( .A1(\ram[12][155] ), .A2(n6560), .A3(n6354), .A4(n9777), 
        .Y(n3288) );
  AO22X1_HVT U3274 ( .A1(\ram[12][156] ), .A2(n6559), .A3(n4622), .A4(n9780), 
        .Y(n3289) );
  AO22X1_HVT U3275 ( .A1(\ram[12][157] ), .A2(n6558), .A3(n4862), .A4(n9783), 
        .Y(n3290) );
  AO22X1_HVT U3276 ( .A1(\ram[12][158] ), .A2(n6557), .A3(n6367), .A4(n9786), 
        .Y(n3291) );
  AO22X1_HVT U3277 ( .A1(\ram[12][159] ), .A2(n6556), .A3(n6353), .A4(n9790), 
        .Y(n3292) );
  AO22X1_HVT U3278 ( .A1(\ram[12][160] ), .A2(n6568), .A3(n6339), .A4(
        data[160]), .Y(n3293) );
  AO22X1_HVT U3279 ( .A1(\ram[12][161] ), .A2(n6567), .A3(n6362), .A4(n9796), 
        .Y(n3294) );
  AO22X1_HVT U3280 ( .A1(\ram[12][162] ), .A2(n4346), .A3(n6338), .A4(
        data[162]), .Y(n3295) );
  AO22X1_HVT U3281 ( .A1(\ram[12][163] ), .A2(n6565), .A3(n6370), .A4(n9802), 
        .Y(n3296) );
  AO22X1_HVT U3282 ( .A1(\ram[12][164] ), .A2(n10146), .A3(n4862), .A4(n9805), 
        .Y(n3297) );
  AO22X1_HVT U3283 ( .A1(\ram[12][165] ), .A2(n6617), .A3(n6332), .A4(
        data[165]), .Y(n3298) );
  AO22X1_HVT U3284 ( .A1(\ram[12][166] ), .A2(n6596), .A3(n6362), .A4(n9811), 
        .Y(n3299) );
  AO22X1_HVT U3285 ( .A1(\ram[12][167] ), .A2(n6595), .A3(n4309), .A4(
        data[167]), .Y(n3300) );
  AO22X1_HVT U3286 ( .A1(\ram[12][168] ), .A2(n6621), .A3(n6358), .A4(n9817), 
        .Y(n3301) );
  AO22X1_HVT U3287 ( .A1(\ram[12][169] ), .A2(n6620), .A3(n6379), .A4(
        data[169]), .Y(n3302) );
  AO22X1_HVT U3288 ( .A1(\ram[12][170] ), .A2(n6565), .A3(n6357), .A4(n9823), 
        .Y(n3303) );
  AO22X1_HVT U3290 ( .A1(\ram[12][172] ), .A2(n6609), .A3(n4310), .A4(n9830), 
        .Y(n3305) );
  AO22X1_HVT U3291 ( .A1(\ram[12][173] ), .A2(n4357), .A3(n4708), .A4(
        data[173]), .Y(n3306) );
  AO22X1_HVT U3292 ( .A1(\ram[12][174] ), .A2(n6605), .A3(n6333), .A4(n9836), 
        .Y(n3307) );
  AO22X1_HVT U3293 ( .A1(\ram[12][175] ), .A2(n6602), .A3(n6352), .A4(n9840), 
        .Y(n3308) );
  AO22X1_HVT U3294 ( .A1(\ram[12][176] ), .A2(n6561), .A3(n6369), .A4(n9843), 
        .Y(n3309) );
  AO22X1_HVT U3295 ( .A1(\ram[12][177] ), .A2(n4275), .A3(n6337), .A4(n9846), 
        .Y(n3310) );
  AO22X1_HVT U3296 ( .A1(\ram[12][178] ), .A2(n6618), .A3(n4708), .A4(n9849), 
        .Y(n3311) );
  AO22X1_HVT U3297 ( .A1(\ram[12][179] ), .A2(n6576), .A3(n6332), .A4(n9853), 
        .Y(n3312) );
  AO22X1_HVT U3298 ( .A1(\ram[12][180] ), .A2(n6588), .A3(n6358), .A4(n9856), 
        .Y(n3313) );
  AO22X1_HVT U3299 ( .A1(\ram[12][181] ), .A2(n6618), .A3(n6359), .A4(n9859), 
        .Y(n3314) );
  AO22X1_HVT U3300 ( .A1(\ram[12][182] ), .A2(n6616), .A3(n4413), .A4(
        data[182]), .Y(n3315) );
  AO22X1_HVT U3301 ( .A1(\ram[12][183] ), .A2(n6615), .A3(n6352), .A4(n9866), 
        .Y(n3316) );
  AO22X1_HVT U3302 ( .A1(\ram[12][184] ), .A2(n6613), .A3(n6335), .A4(
        data[184]), .Y(n3317) );
  AO22X1_HVT U3303 ( .A1(\ram[12][185] ), .A2(n6612), .A3(n6357), .A4(
        data[185]), .Y(n3318) );
  AO22X1_HVT U3304 ( .A1(\ram[12][186] ), .A2(n6610), .A3(n6349), .A4(
        data[186]), .Y(n3319) );
  AO22X1_HVT U3305 ( .A1(\ram[12][187] ), .A2(n6609), .A3(n6362), .A4(n9878), 
        .Y(n3320) );
  AO22X1_HVT U3306 ( .A1(\ram[12][188] ), .A2(n6573), .A3(n6361), .A4(n9881), 
        .Y(n3321) );
  AO22X1_HVT U3307 ( .A1(\ram[12][189] ), .A2(n6616), .A3(n6358), .A4(n9884), 
        .Y(n3322) );
  AO22X1_HVT U3308 ( .A1(\ram[12][190] ), .A2(n6615), .A3(n6339), .A4(n9887), 
        .Y(n3323) );
  AO22X1_HVT U3309 ( .A1(\ram[12][191] ), .A2(n6613), .A3(n6355), .A4(n9891), 
        .Y(n3324) );
  AO22X1_HVT U3310 ( .A1(\ram[12][192] ), .A2(n6598), .A3(n6335), .A4(
        data[192]), .Y(n3325) );
  AO22X1_HVT U3311 ( .A1(\ram[12][193] ), .A2(n6597), .A3(n6375), .A4(
        data[193]), .Y(n3326) );
  AO22X1_HVT U3312 ( .A1(\ram[12][194] ), .A2(n6562), .A3(n6344), .A4(n9900), 
        .Y(n3327) );
  AO22X1_HVT U3313 ( .A1(\ram[12][195] ), .A2(n6616), .A3(n6375), .A4(n9904), 
        .Y(n3328) );
  AO22X1_HVT U3314 ( .A1(\ram[12][196] ), .A2(n6615), .A3(n6376), .A4(n9907), 
        .Y(n3329) );
  AO22X1_HVT U3315 ( .A1(\ram[12][197] ), .A2(n6566), .A3(n6377), .A4(n9910), 
        .Y(n3330) );
  AO22X1_HVT U3316 ( .A1(\ram[12][198] ), .A2(n6596), .A3(n6371), .A4(n9913), 
        .Y(n3331) );
  AO22X1_HVT U3317 ( .A1(\ram[12][199] ), .A2(n6601), .A3(n6372), .A4(n9917), 
        .Y(n3332) );
  AO22X1_HVT U3318 ( .A1(\ram[12][200] ), .A2(n6592), .A3(n4411), .A4(
        data[200]), .Y(n3333) );
  AO22X1_HVT U3319 ( .A1(\ram[12][201] ), .A2(n6591), .A3(n6371), .A4(
        data[201]), .Y(n3334) );
  AO22X1_HVT U3320 ( .A1(\ram[12][202] ), .A2(n6590), .A3(n4708), .A4(
        data[202]), .Y(n3335) );
  AO22X1_HVT U3321 ( .A1(\ram[12][203] ), .A2(n6625), .A3(n6341), .A4(
        data[203]), .Y(n3336) );
  AO22X1_HVT U3322 ( .A1(\ram[12][204] ), .A2(n6624), .A3(n6362), .A4(
        data[204]), .Y(n3337) );
  AO22X1_HVT U3323 ( .A1(\ram[12][205] ), .A2(n6622), .A3(n6354), .A4(
        data[205]), .Y(n3338) );
  AO22X1_HVT U3325 ( .A1(\ram[12][207] ), .A2(n6621), .A3(n4622), .A4(n9942), 
        .Y(n3340) );
  AO22X1_HVT U3326 ( .A1(\ram[12][208] ), .A2(n6620), .A3(n6355), .A4(n9945), 
        .Y(n3341) );
  AO22X1_HVT U3327 ( .A1(\ram[12][209] ), .A2(n6606), .A3(n6358), .A4(
        data[209]), .Y(n3342) );
  AO22X1_HVT U3328 ( .A1(\ram[12][210] ), .A2(n6618), .A3(n6353), .A4(n9951), 
        .Y(n3343) );
  AO22X1_HVT U3329 ( .A1(\ram[12][211] ), .A2(n6560), .A3(n4622), .A4(n9954), 
        .Y(n3344) );
  AO22X1_HVT U3330 ( .A1(\ram[12][212] ), .A2(n6559), .A3(n6338), .A4(n9957), 
        .Y(n3345) );
  AO22X1_HVT U3331 ( .A1(\ram[12][213] ), .A2(n6558), .A3(n4559), .A4(
        data[213]), .Y(n3346) );
  AO22X1_HVT U3332 ( .A1(\ram[12][214] ), .A2(n6557), .A3(n6354), .A4(
        data[214]), .Y(n3347) );
  AO22X1_HVT U3333 ( .A1(\ram[12][215] ), .A2(n6556), .A3(n4619), .A4(n9966), 
        .Y(n3348) );
  AO22X1_HVT U3334 ( .A1(\ram[12][216] ), .A2(n6625), .A3(n6377), .A4(n9969), 
        .Y(n3349) );
  AO22X1_HVT U3335 ( .A1(\ram[12][217] ), .A2(n6624), .A3(n6378), .A4(n9971), 
        .Y(n3350) );
  AO22X1_HVT U3336 ( .A1(\ram[12][218] ), .A2(n6622), .A3(n6334), .A4(n9975), 
        .Y(n3351) );
  AO22X1_HVT U3337 ( .A1(\ram[12][219] ), .A2(n10138), .A3(n6353), .A4(n9979), 
        .Y(n3352) );
  AO22X1_HVT U3338 ( .A1(\ram[12][220] ), .A2(n6621), .A3(n4685), .A4(n9982), 
        .Y(n3353) );
  AO22X1_HVT U3339 ( .A1(\ram[12][221] ), .A2(n6620), .A3(n4549), .A4(n9985), 
        .Y(n3354) );
  AO22X1_HVT U3340 ( .A1(\ram[12][222] ), .A2(n6619), .A3(n6339), .A4(
        data[222]), .Y(n3355) );
  AO22X1_HVT U3341 ( .A1(\ram[12][223] ), .A2(n6598), .A3(n6363), .A4(
        data[223]), .Y(n3356) );
  AO22X1_HVT U3342 ( .A1(\ram[12][224] ), .A2(n6597), .A3(n6352), .A4(n9994), 
        .Y(n3357) );
  AO22X1_HVT U3343 ( .A1(\ram[12][225] ), .A2(n6562), .A3(n4310), .A4(n9997), 
        .Y(n3358) );
  AO22X1_HVT U3344 ( .A1(\ram[12][226] ), .A2(n6561), .A3(n6376), .A4(n10000), 
        .Y(n3359) );
  AO22X1_HVT U3345 ( .A1(\ram[12][227] ), .A2(n6625), .A3(n6361), .A4(
        data[227]), .Y(n3360) );
  AO22X1_HVT U3346 ( .A1(\ram[12][228] ), .A2(n6612), .A3(n4686), .A4(
        data[228]), .Y(n3361) );
  AO22X1_HVT U3347 ( .A1(\ram[12][229] ), .A2(n6610), .A3(n6339), .A4(
        data[229]), .Y(n3362) );
  AO22X1_HVT U3348 ( .A1(\ram[12][230] ), .A2(n6609), .A3(n4707), .A4(
        data[230]), .Y(n3363) );
  AO22X1_HVT U3349 ( .A1(\ram[12][231] ), .A2(n6573), .A3(n6355), .A4(n10016), 
        .Y(n3364) );
  AO22X1_HVT U3350 ( .A1(\ram[12][232] ), .A2(n6605), .A3(n6379), .A4(
        data[232]), .Y(n3365) );
  AO22X1_HVT U3351 ( .A1(\ram[12][233] ), .A2(n6602), .A3(n4550), .A4(
        data[233]), .Y(n3366) );
  AO22X1_HVT U3352 ( .A1(\ram[12][234] ), .A2(n6601), .A3(n6332), .A4(
        data[234]), .Y(n3367) );
  AO22X1_HVT U3353 ( .A1(\ram[12][235] ), .A2(n6561), .A3(n6347), .A4(n10028), 
        .Y(n3368) );
  AO22X1_HVT U3354 ( .A1(\ram[12][236] ), .A2(n6625), .A3(n6358), .A4(n10031), 
        .Y(n3369) );
  AO22X1_HVT U3355 ( .A1(\ram[12][237] ), .A2(n6624), .A3(n6354), .A4(
        data[237]), .Y(n3370) );
  AO22X1_HVT U3356 ( .A1(\ram[12][238] ), .A2(n6622), .A3(n6359), .A4(n10037), 
        .Y(n3371) );
  AO22X1_HVT U3357 ( .A1(\ram[12][239] ), .A2(n6612), .A3(n6333), .A4(n10041), 
        .Y(n3372) );
  AO22X1_HVT U3358 ( .A1(\ram[12][240] ), .A2(n6619), .A3(n6342), .A4(
        data[240]), .Y(n3373) );
  AO22X1_HVT U3359 ( .A1(\ram[12][241] ), .A2(n4346), .A3(n4685), .A4(
        data[241]), .Y(n3374) );
  AO22X1_HVT U3360 ( .A1(\ram[12][242] ), .A2(n4360), .A3(n4550), .A4(
        data[242]), .Y(n3375) );
  AO22X1_HVT U3361 ( .A1(\ram[12][243] ), .A2(n6595), .A3(n4619), .A4(
        data[243]), .Y(n3376) );
  AO22X1_HVT U3362 ( .A1(\ram[12][244] ), .A2(n6560), .A3(n6349), .A4(n10056), 
        .Y(n3377) );
  AO22X1_HVT U3363 ( .A1(\ram[12][245] ), .A2(n6559), .A3(n6348), .A4(
        data[245]), .Y(n3378) );
  AO22X1_HVT U3364 ( .A1(\ram[12][246] ), .A2(n6558), .A3(n4309), .A4(n10062), 
        .Y(n3379) );
  AO22X1_HVT U3365 ( .A1(\ram[12][247] ), .A2(n6557), .A3(n6375), .A4(n10066), 
        .Y(n3380) );
  AO22X1_HVT U3366 ( .A1(\ram[12][248] ), .A2(n6556), .A3(n6380), .A4(
        data[248]), .Y(n3381) );
  AO22X1_HVT U3367 ( .A1(\ram[12][249] ), .A2(n6597), .A3(n6347), .A4(n10072), 
        .Y(n3382) );
  AO22X1_HVT U3368 ( .A1(\ram[12][250] ), .A2(n6562), .A3(n6343), .A4(n10075), 
        .Y(n3383) );
  AO22X1_HVT U3369 ( .A1(\ram[12][251] ), .A2(n6561), .A3(n4686), .A4(n10079), 
        .Y(n3384) );
  AO22X1_HVT U3370 ( .A1(\ram[12][252] ), .A2(n6556), .A3(n6378), .A4(
        data[252]), .Y(n3385) );
  AO22X1_HVT U3371 ( .A1(\ram[12][253] ), .A2(n6595), .A3(n6380), .A4(n10085), 
        .Y(n3386) );
  AO22X1_HVT U3372 ( .A1(\ram[12][254] ), .A2(n6560), .A3(n6337), .A4(
        data[254]), .Y(n3387) );
  AO22X1_HVT U3373 ( .A1(\ram[12][255] ), .A2(n10144), .A3(n6347), .A4(n10092), 
        .Y(n3388) );
  AND2X1_HVT U3374 ( .A1(n50), .A2(n6258), .Y(n49) );
  AND2X1_HVT U3376 ( .A1(n5935), .A2(n5130), .Y(n50) );
  AO22X1_HVT U3378 ( .A1(\ram[13][0] ), .A2(n6982), .A3(n4599), .A4(data[0]), 
        .Y(n3389) );
  AO22X1_HVT U3379 ( .A1(\ram[13][1] ), .A2(n6982), .A3(n8931), .A4(n9309), 
        .Y(n3390) );
  AO22X1_HVT U3380 ( .A1(\ram[13][2] ), .A2(n6976), .A3(n4599), .A4(n9313), 
        .Y(n3391) );
  AO22X1_HVT U3382 ( .A1(\ram[13][4] ), .A2(n6978), .A3(n8943), .A4(n9319), 
        .Y(n3393) );
  AO22X1_HVT U3383 ( .A1(\ram[13][5] ), .A2(n6977), .A3(n8928), .A4(data[5]), 
        .Y(n3394) );
  AO22X1_HVT U3384 ( .A1(\ram[13][6] ), .A2(n4705), .A3(n4299), .A4(n9325), 
        .Y(n3395) );
  AO22X1_HVT U3385 ( .A1(\ram[13][7] ), .A2(n4715), .A3(n8929), .A4(n9328), 
        .Y(n3396) );
  AO22X1_HVT U3386 ( .A1(\ram[13][8] ), .A2(n6978), .A3(n8936), .A4(data[8]), 
        .Y(n3397) );
  AO22X1_HVT U3387 ( .A1(\ram[13][9] ), .A2(n6977), .A3(n4584), .A4(n9334), 
        .Y(n3398) );
  AO22X1_HVT U3388 ( .A1(\ram[13][10] ), .A2(n4542), .A3(n4589), .A4(n9337), 
        .Y(n3399) );
  AO22X1_HVT U3390 ( .A1(\ram[13][12] ), .A2(n7001), .A3(n8942), .A4(n9345), 
        .Y(n3401) );
  AO22X1_HVT U3391 ( .A1(\ram[13][13] ), .A2(n7000), .A3(n8941), .A4(n9348), 
        .Y(n3402) );
  AO22X1_HVT U3392 ( .A1(\ram[13][14] ), .A2(n6999), .A3(n8940), .A4(data[14]), 
        .Y(n3403) );
  AO22X1_HVT U3393 ( .A1(\ram[13][15] ), .A2(n4763), .A3(n8931), .A4(n9354), 
        .Y(n3404) );
  AO22X1_HVT U3394 ( .A1(\ram[13][16] ), .A2(n6996), .A3(n8943), .A4(n9357), 
        .Y(n3405) );
  AO22X1_HVT U3395 ( .A1(\ram[13][17] ), .A2(n6995), .A3(n8942), .A4(data[17]), 
        .Y(n3406) );
  AO22X1_HVT U3396 ( .A1(\ram[13][18] ), .A2(n6994), .A3(n8941), .A4(data[18]), 
        .Y(n3407) );
  AO22X1_HVT U3397 ( .A1(\ram[13][19] ), .A2(n6993), .A3(n8940), .A4(data[19]), 
        .Y(n3408) );
  AO22X1_HVT U3398 ( .A1(\ram[13][20] ), .A2(n7025), .A3(n5455), .A4(data[20]), 
        .Y(n3409) );
  AO22X1_HVT U3399 ( .A1(\ram[13][21] ), .A2(n7024), .A3(n5455), .A4(n9370), 
        .Y(n3410) );
  AO22X1_HVT U3400 ( .A1(\ram[13][22] ), .A2(n7023), .A3(n8944), .A4(n9374), 
        .Y(n3411) );
  AO22X1_HVT U3401 ( .A1(\ram[13][23] ), .A2(n7022), .A3(n4786), .A4(data[23]), 
        .Y(n3412) );
  AO22X1_HVT U3402 ( .A1(\ram[13][24] ), .A2(n7013), .A3(n4698), .A4(data[24]), 
        .Y(n3413) );
  AO22X1_HVT U3403 ( .A1(\ram[13][25] ), .A2(n7010), .A3(n8925), .A4(data[25]), 
        .Y(n3414) );
  AO22X1_HVT U3404 ( .A1(\ram[13][26] ), .A2(n7011), .A3(n4781), .A4(n9386), 
        .Y(n3415) );
  AO22X1_HVT U3407 ( .A1(\ram[13][29] ), .A2(n7000), .A3(n8914), .A4(data[29]), 
        .Y(n3418) );
  AO22X1_HVT U3409 ( .A1(\ram[13][31] ), .A2(n4763), .A3(n8912), .A4(n9401), 
        .Y(n3420) );
  AO22X1_HVT U3410 ( .A1(\ram[13][32] ), .A2(n7012), .A3(n8949), .A4(n9404), 
        .Y(n3421) );
  AO22X1_HVT U3411 ( .A1(\ram[13][33] ), .A2(n7011), .A3(n4852), .A4(n9407), 
        .Y(n3422) );
  AO22X1_HVT U3412 ( .A1(\ram[13][34] ), .A2(n6984), .A3(n4934), .A4(n9410), 
        .Y(n3423) );
  AO22X1_HVT U3413 ( .A1(\ram[13][35] ), .A2(n4715), .A3(n4699), .A4(n9413), 
        .Y(n3424) );
  AO22X1_HVT U3414 ( .A1(\ram[13][36] ), .A2(n7021), .A3(n4853), .A4(n9416), 
        .Y(n3425) );
  AO22X1_HVT U3415 ( .A1(\ram[13][37] ), .A2(n4834), .A3(n8919), .A4(n9418), 
        .Y(n3426) );
  AO22X1_HVT U3416 ( .A1(\ram[13][38] ), .A2(n7020), .A3(n4852), .A4(n9422), 
        .Y(n3427) );
  AO22X1_HVT U3417 ( .A1(\ram[13][39] ), .A2(n7020), .A3(n8917), .A4(n9425), 
        .Y(n3428) );
  AO22X1_HVT U3418 ( .A1(\ram[13][40] ), .A2(n7021), .A3(n4786), .A4(n9428), 
        .Y(n3429) );
  AO22X1_HVT U3419 ( .A1(\ram[13][41] ), .A2(n4448), .A3(n8945), .A4(n9431), 
        .Y(n3430) );
  AO22X1_HVT U3420 ( .A1(\ram[13][42] ), .A2(n7020), .A3(n5455), .A4(data[42]), 
        .Y(n3431) );
  AO22X1_HVT U3421 ( .A1(\ram[13][43] ), .A2(n7019), .A3(n8946), .A4(data[43]), 
        .Y(n3432) );
  AO22X1_HVT U3422 ( .A1(\ram[13][44] ), .A2(n4542), .A3(n8943), .A4(data[44]), 
        .Y(n3433) );
  AO22X1_HVT U3423 ( .A1(\ram[13][45] ), .A2(n6984), .A3(n8942), .A4(data[45]), 
        .Y(n3434) );
  AO22X1_HVT U3424 ( .A1(\ram[13][46] ), .A2(n6981), .A3(n8941), .A4(n9446), 
        .Y(n3435) );
  AO22X1_HVT U3425 ( .A1(\ram[13][47] ), .A2(n6981), .A3(n8940), .A4(data[47]), 
        .Y(n3436) );
  AO22X1_HVT U3426 ( .A1(\ram[13][48] ), .A2(n6978), .A3(n4932), .A4(n9451), 
        .Y(n3437) );
  AO22X1_HVT U3427 ( .A1(\ram[13][49] ), .A2(n6977), .A3(n4936), .A4(data[49]), 
        .Y(n3438) );
  AO22X1_HVT U3428 ( .A1(\ram[13][50] ), .A2(n6990), .A3(n4934), .A4(n9458), 
        .Y(n3439) );
  AO22X1_HVT U3429 ( .A1(\ram[13][51] ), .A2(n4901), .A3(n8950), .A4(data[51]), 
        .Y(n3440) );
  AO22X1_HVT U3430 ( .A1(\ram[13][52] ), .A2(n7021), .A3(n8959), .A4(data[52]), 
        .Y(n3441) );
  AO22X1_HVT U3431 ( .A1(\ram[13][53] ), .A2(n5083), .A3(n8958), .A4(data[53]), 
        .Y(n3442) );
  AO22X1_HVT U3432 ( .A1(\ram[13][54] ), .A2(n4832), .A3(n4788), .A4(n9470), 
        .Y(n3443) );
  AO22X1_HVT U3433 ( .A1(\ram[13][55] ), .A2(n4761), .A3(n8960), .A4(n9473), 
        .Y(n3444) );
  AO22X1_HVT U3434 ( .A1(\ram[13][56] ), .A2(n7000), .A3(n8925), .A4(n9476), 
        .Y(n3445) );
  AO22X1_HVT U3435 ( .A1(\ram[13][57] ), .A2(n6999), .A3(n8925), .A4(n9479), 
        .Y(n3446) );
  AO22X1_HVT U3436 ( .A1(\ram[13][58] ), .A2(n4763), .A3(n8917), .A4(n9482), 
        .Y(n3447) );
  AO22X1_HVT U3440 ( .A1(\ram[13][62] ), .A2(n6993), .A3(n4781), .A4(data[62]), 
        .Y(n3451) );
  AO22X1_HVT U3441 ( .A1(\ram[13][63] ), .A2(n7001), .A3(n8917), .A4(n9497), 
        .Y(n3452) );
  AO22X1_HVT U3442 ( .A1(\ram[13][64] ), .A2(n7001), .A3(n8915), .A4(n9500), 
        .Y(n3453) );
  AO22X1_HVT U3443 ( .A1(\ram[13][65] ), .A2(n7000), .A3(n8914), .A4(n9503), 
        .Y(n3454) );
  AO22X1_HVT U3444 ( .A1(\ram[13][66] ), .A2(n6999), .A3(n8913), .A4(data[66]), 
        .Y(n3455) );
  AO22X1_HVT U3445 ( .A1(\ram[13][67] ), .A2(n4763), .A3(n4698), .A4(n9509), 
        .Y(n3456) );
  AO22X1_HVT U3447 ( .A1(\ram[13][69] ), .A2(n7000), .A3(n8963), .A4(n9515), 
        .Y(n3458) );
  AO22X1_HVT U3448 ( .A1(\ram[13][70] ), .A2(n6999), .A3(n8949), .A4(n9518), 
        .Y(n3459) );
  AO22X1_HVT U3451 ( .A1(\ram[13][73] ), .A2(n6974), .A3(n4698), .A4(data[73]), 
        .Y(n3462) );
  AO22X1_HVT U3452 ( .A1(\ram[13][74] ), .A2(n4828), .A3(n4526), .A4(data[74]), 
        .Y(n3463) );
  AO22X1_HVT U3454 ( .A1(\ram[13][76] ), .A2(n6971), .A3(n8945), .A4(n9536), 
        .Y(n3465) );
  AO22X1_HVT U3456 ( .A1(\ram[13][78] ), .A2(n7004), .A3(n8946), .A4(data[78]), 
        .Y(n3467) );
  AO22X1_HVT U3457 ( .A1(\ram[13][79] ), .A2(n4832), .A3(n8943), .A4(n9545), 
        .Y(n3468) );
  AO22X1_HVT U3458 ( .A1(\ram[13][80] ), .A2(n4831), .A3(n8942), .A4(n9548), 
        .Y(n3469) );
  AO22X1_HVT U3459 ( .A1(\ram[13][81] ), .A2(n7001), .A3(n8941), .A4(n9551), 
        .Y(n3470) );
  AO22X1_HVT U3460 ( .A1(\ram[13][82] ), .A2(n7000), .A3(n8940), .A4(n9554), 
        .Y(n3471) );
  AO22X1_HVT U3462 ( .A1(\ram[13][84] ), .A2(n7005), .A3(n8937), .A4(data[84]), 
        .Y(n3473) );
  AO22X1_HVT U3463 ( .A1(\ram[13][85] ), .A2(n7004), .A3(n8937), .A4(data[85]), 
        .Y(n3474) );
  AO22X1_HVT U3464 ( .A1(\ram[13][86] ), .A2(n7003), .A3(n8935), .A4(data[86]), 
        .Y(n3475) );
  AO22X1_HVT U3465 ( .A1(\ram[13][87] ), .A2(n7002), .A3(n8934), .A4(n9569), 
        .Y(n3476) );
  AO22X1_HVT U3466 ( .A1(\ram[13][88] ), .A2(n4714), .A3(n4932), .A4(n9572), 
        .Y(n3477) );
  AO22X1_HVT U3467 ( .A1(\ram[13][89] ), .A2(n4901), .A3(n4788), .A4(data[89]), 
        .Y(n3478) );
  AO22X1_HVT U3468 ( .A1(\ram[13][90] ), .A2(n4900), .A3(n8952), .A4(n9578), 
        .Y(n3479) );
  AO22X1_HVT U3469 ( .A1(\ram[13][91] ), .A2(n4900), .A3(n8949), .A4(n9581), 
        .Y(n3480) );
  AO22X1_HVT U3470 ( .A1(\ram[13][92] ), .A2(n4541), .A3(n8960), .A4(n9584), 
        .Y(n3481) );
  AO22X1_HVT U3471 ( .A1(\ram[13][93] ), .A2(n6976), .A3(n8959), .A4(data[93]), 
        .Y(n3482) );
  AO22X1_HVT U3472 ( .A1(\ram[13][94] ), .A2(n6988), .A3(n8960), .A4(n9590), 
        .Y(n3483) );
  AO22X1_HVT U3473 ( .A1(\ram[13][95] ), .A2(n6988), .A3(n8960), .A4(n9593), 
        .Y(n3484) );
  AO22X1_HVT U3474 ( .A1(\ram[13][96] ), .A2(n6996), .A3(n8926), .A4(n9596), 
        .Y(n3485) );
  AO22X1_HVT U3475 ( .A1(\ram[13][97] ), .A2(n6995), .A3(n8923), .A4(data[97]), 
        .Y(n3486) );
  AO22X1_HVT U3476 ( .A1(\ram[13][98] ), .A2(n6994), .A3(n8924), .A4(data[98]), 
        .Y(n3487) );
  AO22X1_HVT U3477 ( .A1(\ram[13][99] ), .A2(n4485), .A3(n8915), .A4(n9605), 
        .Y(n3488) );
  AO22X1_HVT U3478 ( .A1(\ram[13][100] ), .A2(n6990), .A3(n8914), .A4(
        data[100]), .Y(n3489) );
  AO22X1_HVT U3480 ( .A1(\ram[13][102] ), .A2(n4824), .A3(n4698), .A4(n9614), 
        .Y(n3491) );
  AO22X1_HVT U3481 ( .A1(\ram[13][103] ), .A2(n6978), .A3(n8965), .A4(n9617), 
        .Y(n3492) );
  AO22X1_HVT U3482 ( .A1(\ram[13][104] ), .A2(n6977), .A3(n8915), .A4(
        data[104]), .Y(n3493) );
  AO22X1_HVT U3483 ( .A1(\ram[13][105] ), .A2(n4705), .A3(n8914), .A4(n9623), 
        .Y(n3494) );
  AO22X1_HVT U3484 ( .A1(\ram[13][106] ), .A2(n6984), .A3(n8913), .A4(
        data[106]), .Y(n3495) );
  AO22X1_HVT U3485 ( .A1(\ram[13][107] ), .A2(n4760), .A3(n8926), .A4(
        data[107]), .Y(n3496) );
  AO22X1_HVT U3486 ( .A1(\ram[13][108] ), .A2(n6978), .A3(n8954), .A4(n9632), 
        .Y(n3497) );
  AO22X1_HVT U3487 ( .A1(\ram[13][109] ), .A2(n6977), .A3(n4932), .A4(
        data[109]), .Y(n3498) );
  AO22X1_HVT U3488 ( .A1(\ram[13][110] ), .A2(n6989), .A3(n8953), .A4(
        data[110]), .Y(n3499) );
  AO22X1_HVT U3489 ( .A1(\ram[13][111] ), .A2(n4901), .A3(n5454), .A4(
        data[111]), .Y(n3500) );
  AO22X1_HVT U3490 ( .A1(\ram[13][112] ), .A2(n7011), .A3(n4932), .A4(
        data[112]), .Y(n3501) );
  AO22X1_HVT U3491 ( .A1(\ram[13][113] ), .A2(n7014), .A3(n8952), .A4(
        data[113]), .Y(n3502) );
  AO22X1_HVT U3492 ( .A1(\ram[13][114] ), .A2(n7014), .A3(n8950), .A4(
        data[114]), .Y(n3503) );
  AO22X1_HVT U3493 ( .A1(\ram[13][115] ), .A2(n7010), .A3(n4936), .A4(n9653), 
        .Y(n3504) );
  AO22X1_HVT U3494 ( .A1(\ram[13][116] ), .A2(n7011), .A3(n8961), .A4(n9656), 
        .Y(n3505) );
  AO22X1_HVT U3495 ( .A1(\ram[13][117] ), .A2(n4669), .A3(n8958), .A4(
        data[117]), .Y(n3506) );
  AO22X1_HVT U3496 ( .A1(\ram[13][118] ), .A2(n4669), .A3(n8959), .A4(n9661), 
        .Y(n3507) );
  AO22X1_HVT U3497 ( .A1(\ram[13][119] ), .A2(n4668), .A3(n8958), .A4(
        data[119]), .Y(n3508) );
  AO22X1_HVT U3498 ( .A1(\ram[13][120] ), .A2(n4714), .A3(n8959), .A4(
        data[120]), .Y(n3509) );
  AO22X1_HVT U3500 ( .A1(\ram[13][122] ), .A2(n6981), .A3(n8912), .A4(
        data[122]), .Y(n3511) );
  AO22X1_HVT U3501 ( .A1(\ram[13][123] ), .A2(n6981), .A3(n8933), .A4(n9677), 
        .Y(n3512) );
  AO22X1_HVT U3502 ( .A1(\ram[13][124] ), .A2(n6976), .A3(n8955), .A4(n9680), 
        .Y(n3513) );
  AO22X1_HVT U3503 ( .A1(\ram[13][125] ), .A2(n4705), .A3(n8962), .A4(n9683), 
        .Y(n3514) );
  AO22X1_HVT U3504 ( .A1(\ram[13][126] ), .A2(n4824), .A3(n8954), .A4(
        data[126]), .Y(n3515) );
  AO22X1_HVT U3505 ( .A1(\ram[13][127] ), .A2(n6987), .A3(n4934), .A4(n9689), 
        .Y(n3516) );
  AO22X1_HVT U3506 ( .A1(\ram[13][128] ), .A2(n6996), .A3(n4526), .A4(n9692), 
        .Y(n3517) );
  AO22X1_HVT U3507 ( .A1(\ram[13][129] ), .A2(n6995), .A3(n8913), .A4(
        data[129]), .Y(n3518) );
  AO22X1_HVT U3508 ( .A1(\ram[13][130] ), .A2(n6994), .A3(n8934), .A4(n9698), 
        .Y(n3519) );
  AO22X1_HVT U3509 ( .A1(\ram[13][131] ), .A2(n6993), .A3(n8930), .A4(n9701), 
        .Y(n3520) );
  AO22X1_HVT U3510 ( .A1(\ram[13][132] ), .A2(n5083), .A3(n8918), .A4(n9704), 
        .Y(n3521) );
  AO22X1_HVT U3511 ( .A1(\ram[13][133] ), .A2(n7014), .A3(n8919), .A4(n9707), 
        .Y(n3522) );
  AO22X1_HVT U3512 ( .A1(\ram[13][134] ), .A2(n7015), .A3(n8961), .A4(n9710), 
        .Y(n3523) );
  AO22X1_HVT U3513 ( .A1(\ram[13][135] ), .A2(n7012), .A3(n4936), .A4(n9713), 
        .Y(n3524) );
  AO22X1_HVT U3515 ( .A1(\ram[13][137] ), .A2(n7011), .A3(n8952), .A4(n9719), 
        .Y(n3526) );
  AO22X1_HVT U3516 ( .A1(\ram[13][138] ), .A2(n7008), .A3(n8926), .A4(n9722), 
        .Y(n3527) );
  AO22X1_HVT U3517 ( .A1(\ram[13][139] ), .A2(n7021), .A3(n8930), .A4(n9726), 
        .Y(n3528) );
  AO22X1_HVT U3518 ( .A1(\ram[13][140] ), .A2(n6990), .A3(n8923), .A4(
        data[140]), .Y(n3529) );
  AO22X1_HVT U3519 ( .A1(\ram[13][141] ), .A2(n6989), .A3(n8920), .A4(
        data[141]), .Y(n3530) );
  AO22X1_HVT U3521 ( .A1(\ram[13][143] ), .A2(n6987), .A3(n5454), .A4(n9739), 
        .Y(n3532) );
  AO22X1_HVT U3523 ( .A1(\ram[13][145] ), .A2(n4714), .A3(n4758), .A4(n9745), 
        .Y(n3534) );
  AO22X1_HVT U3524 ( .A1(\ram[13][146] ), .A2(n6975), .A3(n4781), .A4(
        data[146]), .Y(n3535) );
  AO22X1_HVT U3525 ( .A1(\ram[13][147] ), .A2(n4900), .A3(n8934), .A4(n9752), 
        .Y(n3536) );
  AO22X1_HVT U3526 ( .A1(\ram[13][148] ), .A2(n6982), .A3(n4477), .A4(n9755), 
        .Y(n3537) );
  AO22X1_HVT U3527 ( .A1(\ram[13][149] ), .A2(n6975), .A3(n8936), .A4(
        data[149]), .Y(n3538) );
  AO22X1_HVT U3528 ( .A1(\ram[13][150] ), .A2(n4901), .A3(n8958), .A4(n9761), 
        .Y(n3539) );
  AO22X1_HVT U3529 ( .A1(\ram[13][151] ), .A2(n6982), .A3(n4788), .A4(n9764), 
        .Y(n3540) );
  AO22X1_HVT U3530 ( .A1(\ram[13][152] ), .A2(n4900), .A3(n4788), .A4(
        data[152]), .Y(n3541) );
  AO22X1_HVT U3531 ( .A1(\ram[13][153] ), .A2(n6974), .A3(n8950), .A4(n9770), 
        .Y(n3542) );
  AO22X1_HVT U3532 ( .A1(\ram[13][154] ), .A2(n4828), .A3(n8924), .A4(
        data[154]), .Y(n3543) );
  AO22X1_HVT U3533 ( .A1(\ram[13][155] ), .A2(n4825), .A3(n8935), .A4(n9777), 
        .Y(n3544) );
  AO22X1_HVT U3534 ( .A1(\ram[13][156] ), .A2(n6996), .A3(n8925), .A4(n9780), 
        .Y(n3545) );
  AO22X1_HVT U3535 ( .A1(\ram[13][157] ), .A2(n6995), .A3(n8952), .A4(
        data[157]), .Y(n3546) );
  AO22X1_HVT U3536 ( .A1(\ram[13][158] ), .A2(n6994), .A3(n8965), .A4(n9786), 
        .Y(n3547) );
  AO22X1_HVT U3537 ( .A1(\ram[13][159] ), .A2(n6993), .A3(n8928), .A4(n9790), 
        .Y(n3548) );
  AO22X1_HVT U3538 ( .A1(\ram[13][160] ), .A2(n7015), .A3(n4853), .A4(n9793), 
        .Y(n3549) );
  AO22X1_HVT U3540 ( .A1(\ram[13][162] ), .A2(n7012), .A3(n4758), .A4(n9799), 
        .Y(n3551) );
  AO22X1_HVT U3541 ( .A1(\ram[13][163] ), .A2(n7013), .A3(n8965), .A4(
        data[163]), .Y(n3552) );
  AO22X1_HVT U3542 ( .A1(\ram[13][164] ), .A2(n7005), .A3(n8930), .A4(n9805), 
        .Y(n3553) );
  AO22X1_HVT U3543 ( .A1(\ram[13][165] ), .A2(n4833), .A3(n4526), .A4(n9808), 
        .Y(n3554) );
  AO22X1_HVT U3544 ( .A1(\ram[13][166] ), .A2(n7003), .A3(n8964), .A4(n9811), 
        .Y(n3555) );
  AO22X1_HVT U3545 ( .A1(\ram[13][167] ), .A2(n4831), .A3(n8954), .A4(n9814), 
        .Y(n3556) );
  AO22X1_HVT U3546 ( .A1(\ram[13][168] ), .A2(n4705), .A3(n8960), .A4(
        data[168]), .Y(n3557) );
  AO22X1_HVT U3547 ( .A1(\ram[13][169] ), .A2(n6976), .A3(n8931), .A4(n9820), 
        .Y(n3558) );
  AO22X1_HVT U3548 ( .A1(\ram[13][170] ), .A2(n6987), .A3(n8955), .A4(n9823), 
        .Y(n3559) );
  AO22X1_HVT U3549 ( .A1(\ram[13][171] ), .A2(n6988), .A3(n8964), .A4(n9827), 
        .Y(n3560) );
  AO22X1_HVT U3550 ( .A1(\ram[13][172] ), .A2(n6978), .A3(n8961), .A4(
        data[172]), .Y(n3561) );
  AO22X1_HVT U3551 ( .A1(\ram[13][173] ), .A2(n6977), .A3(n8962), .A4(n9833), 
        .Y(n3562) );
  AO22X1_HVT U3552 ( .A1(\ram[13][174] ), .A2(n6990), .A3(n8929), .A4(n9836), 
        .Y(n3563) );
  AO22X1_HVT U3553 ( .A1(\ram[13][175] ), .A2(n6975), .A3(n8914), .A4(n9840), 
        .Y(n3564) );
  AO22X1_HVT U3554 ( .A1(\ram[13][176] ), .A2(n4828), .A3(n8935), .A4(
        data[176]), .Y(n3565) );
  AO22X1_HVT U3555 ( .A1(\ram[13][177] ), .A2(n6973), .A3(n8929), .A4(n9846), 
        .Y(n3566) );
  AO22X1_HVT U3556 ( .A1(\ram[13][178] ), .A2(n4825), .A3(n8915), .A4(n9849), 
        .Y(n3567) );
  AO22X1_HVT U3557 ( .A1(\ram[13][179] ), .A2(n6971), .A3(n4584), .A4(n9853), 
        .Y(n3568) );
  AO22X1_HVT U3558 ( .A1(\ram[13][180] ), .A2(n4834), .A3(n8945), .A4(
        data[180]), .Y(n3569) );
  AO22X1_HVT U3559 ( .A1(\ram[13][181] ), .A2(n7004), .A3(n8953), .A4(
        data[181]), .Y(n3570) );
  AO22X1_HVT U3560 ( .A1(\ram[13][182] ), .A2(n7003), .A3(n4477), .A4(n9862), 
        .Y(n3571) );
  AO22X1_HVT U3561 ( .A1(\ram[13][183] ), .A2(n7002), .A3(n4786), .A4(n9866), 
        .Y(n3572) );
  AO22X1_HVT U3562 ( .A1(\ram[13][184] ), .A2(n4481), .A3(n5454), .A4(n9869), 
        .Y(n3573) );
  AO22X1_HVT U3563 ( .A1(\ram[13][185] ), .A2(n7024), .A3(n8928), .A4(n9872), 
        .Y(n3574) );
  AO22X1_HVT U3564 ( .A1(\ram[13][186] ), .A2(n7023), .A3(n8945), .A4(n9875), 
        .Y(n3575) );
  AO22X1_HVT U3565 ( .A1(\ram[13][187] ), .A2(n7022), .A3(n8944), .A4(n9878), 
        .Y(n3576) );
  AO22X1_HVT U3566 ( .A1(\ram[13][188] ), .A2(n7025), .A3(n8949), .A4(
        data[188]), .Y(n3577) );
  AO22X1_HVT U3568 ( .A1(\ram[13][190] ), .A2(n7023), .A3(n8930), .A4(
        data[190]), .Y(n3579) );
  AO22X1_HVT U3569 ( .A1(\ram[13][191] ), .A2(n7022), .A3(n4299), .A4(n9891), 
        .Y(n3580) );
  AO22X1_HVT U3570 ( .A1(\ram[13][192] ), .A2(n6972), .A3(n4786), .A4(n9894), 
        .Y(n3581) );
  AO22X1_HVT U3571 ( .A1(\ram[13][193] ), .A2(n7008), .A3(n8944), .A4(n9897), 
        .Y(n3582) );
  AO22X1_HVT U3572 ( .A1(\ram[13][194] ), .A2(n7015), .A3(n8944), .A4(n9899), 
        .Y(n3583) );
  AO22X1_HVT U3573 ( .A1(\ram[13][195] ), .A2(n7015), .A3(n8943), .A4(n9904), 
        .Y(n3584) );
  AO22X1_HVT U3574 ( .A1(\ram[13][196] ), .A2(n7009), .A3(n8942), .A4(n9907), 
        .Y(n3585) );
  AO22X1_HVT U3575 ( .A1(\ram[13][197] ), .A2(n4228), .A3(n8941), .A4(n9910), 
        .Y(n3586) );
  AO22X1_HVT U3576 ( .A1(\ram[13][198] ), .A2(n7024), .A3(n8940), .A4(n9913), 
        .Y(n3587) );
  AO22X1_HVT U3577 ( .A1(\ram[13][199] ), .A2(n7023), .A3(n8931), .A4(n9917), 
        .Y(n3588) );
  AO22X1_HVT U3578 ( .A1(\ram[13][200] ), .A2(n7022), .A3(n8913), .A4(n9920), 
        .Y(n3589) );
  AO22X1_HVT U3579 ( .A1(\ram[13][201] ), .A2(n5083), .A3(n8924), .A4(n9922), 
        .Y(n3590) );
  AO22X1_HVT U3580 ( .A1(\ram[13][202] ), .A2(n6991), .A3(n8915), .A4(n9926), 
        .Y(n3591) );
  AO22X1_HVT U3581 ( .A1(\ram[13][203] ), .A2(n7020), .A3(n8914), .A4(n9928), 
        .Y(n3592) );
  AO22X1_HVT U3582 ( .A1(\ram[13][204] ), .A2(n6973), .A3(n8920), .A4(n9932), 
        .Y(n3593) );
  AO22X1_HVT U3583 ( .A1(\ram[13][205] ), .A2(n6974), .A3(n8919), .A4(n9935), 
        .Y(n3594) );
  AO22X1_HVT U3584 ( .A1(\ram[13][206] ), .A2(n6972), .A3(n8918), .A4(
        data[206]), .Y(n3595) );
  AO22X1_HVT U3585 ( .A1(\ram[13][207] ), .A2(n6971), .A3(n8917), .A4(n9942), 
        .Y(n3596) );
  AO22X1_HVT U3586 ( .A1(\ram[13][208] ), .A2(n6973), .A3(n4925), .A4(
        data[208]), .Y(n3597) );
  AO22X1_HVT U3587 ( .A1(\ram[13][209] ), .A2(n4828), .A3(n4925), .A4(n9948), 
        .Y(n3598) );
  AO22X1_HVT U3588 ( .A1(\ram[13][210] ), .A2(n6972), .A3(n8955), .A4(
        data[210]), .Y(n3599) );
  AO22X1_HVT U3589 ( .A1(\ram[13][211] ), .A2(n6971), .A3(n8955), .A4(
        data[211]), .Y(n3600) );
  AO22X1_HVT U3590 ( .A1(\ram[13][212] ), .A2(n7019), .A3(n4584), .A4(
        data[212]), .Y(n3601) );
  AO22X1_HVT U3591 ( .A1(\ram[13][213] ), .A2(n4761), .A3(n8937), .A4(n9959), 
        .Y(n3602) );
  AO22X1_HVT U3592 ( .A1(\ram[13][214] ), .A2(n5083), .A3(n4589), .A4(n9963), 
        .Y(n3603) );
  AO22X1_HVT U3593 ( .A1(\ram[13][215] ), .A2(n4760), .A3(n8934), .A4(n9966), 
        .Y(n3604) );
  AO22X1_HVT U3594 ( .A1(\ram[13][216] ), .A2(n7015), .A3(n8920), .A4(
        data[216]), .Y(n3605) );
  AO22X1_HVT U3595 ( .A1(\ram[13][217] ), .A2(n7009), .A3(n8919), .A4(
        data[217]), .Y(n3606) );
  AO22X1_HVT U3597 ( .A1(\ram[13][219] ), .A2(n4668), .A3(n8923), .A4(n9979), 
        .Y(n3608) );
  AO22X1_HVT U3598 ( .A1(\ram[13][220] ), .A2(n7009), .A3(n4699), .A4(
        data[220]), .Y(n3609) );
  AO22X1_HVT U3599 ( .A1(\ram[13][221] ), .A2(n7008), .A3(n8952), .A4(n9985), 
        .Y(n3610) );
  AO22X1_HVT U3600 ( .A1(\ram[13][222] ), .A2(n4448), .A3(n4934), .A4(n9988), 
        .Y(n3611) );
  AO22X1_HVT U3601 ( .A1(\ram[13][223] ), .A2(n7014), .A3(n4853), .A4(n9991), 
        .Y(n3612) );
  AO22X1_HVT U3602 ( .A1(\ram[13][224] ), .A2(n7015), .A3(n8919), .A4(
        data[224]), .Y(n3613) );
  AO22X1_HVT U3603 ( .A1(\ram[13][225] ), .A2(n7008), .A3(n8918), .A4(n9997), 
        .Y(n3614) );
  AO22X1_HVT U3604 ( .A1(\ram[13][226] ), .A2(n7010), .A3(n8924), .A4(n10000), 
        .Y(n3615) );
  AO22X1_HVT U3605 ( .A1(\ram[13][227] ), .A2(n7013), .A3(n5455), .A4(n10003), 
        .Y(n3616) );
  AO22X1_HVT U3606 ( .A1(\ram[13][228] ), .A2(n6974), .A3(n4853), .A4(n10006), 
        .Y(n3617) );
  AO22X1_HVT U3607 ( .A1(\ram[13][229] ), .A2(n6972), .A3(n8919), .A4(n10009), 
        .Y(n3618) );
  AO22X1_HVT U3608 ( .A1(\ram[13][230] ), .A2(n4825), .A3(n4852), .A4(n10012), 
        .Y(n3619) );
  AO22X1_HVT U3609 ( .A1(\ram[13][231] ), .A2(n7005), .A3(n4781), .A4(n10016), 
        .Y(n3620) );
  AO22X1_HVT U3610 ( .A1(\ram[13][232] ), .A2(n4833), .A3(n8945), .A4(n10019), 
        .Y(n3621) );
  AO22X1_HVT U3611 ( .A1(\ram[13][233] ), .A2(n7003), .A3(n8944), .A4(n10022), 
        .Y(n3622) );
  AO22X1_HVT U3612 ( .A1(\ram[13][234] ), .A2(n7002), .A3(n5455), .A4(n10025), 
        .Y(n3623) );
  AO22X1_HVT U3613 ( .A1(\ram[13][235] ), .A2(n6973), .A3(n8946), .A4(
        data[235]), .Y(n3624) );
  AO22X1_HVT U3614 ( .A1(\ram[13][236] ), .A2(n7005), .A3(n8943), .A4(
        data[236]), .Y(n3625) );
  AO22X1_HVT U3615 ( .A1(\ram[13][237] ), .A2(n4833), .A3(n8942), .A4(n10034), 
        .Y(n3626) );
  AO22X1_HVT U3616 ( .A1(\ram[13][238] ), .A2(n7003), .A3(n8941), .A4(
        data[238]), .Y(n3627) );
  AO22X1_HVT U3617 ( .A1(\ram[13][239] ), .A2(n4831), .A3(n8940), .A4(n10041), 
        .Y(n3628) );
  AO22X1_HVT U3618 ( .A1(\ram[13][240] ), .A2(n4446), .A3(n8963), .A4(
        data[240]), .Y(n3629) );
  AO22X1_HVT U3619 ( .A1(\ram[13][241] ), .A2(n4669), .A3(n8963), .A4(n10047), 
        .Y(n3630) );
  AO22X1_HVT U3620 ( .A1(\ram[13][242] ), .A2(n4669), .A3(n8964), .A4(n10050), 
        .Y(n3631) );
  AO22X1_HVT U3621 ( .A1(\ram[13][243] ), .A2(n7012), .A3(n8963), .A4(n10053), 
        .Y(n3632) );
  AO22X1_HVT U3622 ( .A1(\ram[13][244] ), .A2(n6989), .A3(n4925), .A4(
        data[244]), .Y(n3633) );
  AO22X1_HVT U3623 ( .A1(\ram[13][245] ), .A2(n4541), .A3(n8963), .A4(n10059), 
        .Y(n3634) );
  AO22X1_HVT U3624 ( .A1(\ram[13][246] ), .A2(n6988), .A3(n4925), .A4(n10062), 
        .Y(n3635) );
  AO22X1_HVT U3625 ( .A1(\ram[13][247] ), .A2(n4824), .A3(n8962), .A4(n10066), 
        .Y(n3636) );
  AO22X1_HVT U3626 ( .A1(\ram[13][248] ), .A2(n4228), .A3(n8958), .A4(n10069), 
        .Y(n3637) );
  AO22X1_HVT U3627 ( .A1(\ram[13][249] ), .A2(n7024), .A3(n8961), .A4(n10071), 
        .Y(n3638) );
  AO22X1_HVT U3628 ( .A1(\ram[13][250] ), .A2(n4480), .A3(n8961), .A4(
        data[250]), .Y(n3639) );
  AO22X1_HVT U3629 ( .A1(\ram[13][251] ), .A2(n4485), .A3(n8959), .A4(n10079), 
        .Y(n3640) );
  AO22X1_HVT U3631 ( .A1(\ram[13][253] ), .A2(n6992), .A3(n4786), .A4(
        data[253]), .Y(n3642) );
  AO22X1_HVT U3632 ( .A1(\ram[13][254] ), .A2(n7013), .A3(n8955), .A4(n10088), 
        .Y(n3643) );
  AO22X1_HVT U3633 ( .A1(\ram[13][255] ), .A2(n4668), .A3(n4758), .A4(n10092), 
        .Y(n3644) );
  AND2X1_HVT U3634 ( .A1(n5645), .A2(n54), .Y(n53) );
  AND2X1_HVT U3636 ( .A1(n5563), .A2(n5935), .Y(n54) );
  AND2X1_HVT U3637 ( .A1(n5659), .A2(n5114), .Y(n13) );
  AO22X1_HVT U3638 ( .A1(\ram[14][0] ), .A2(n7210), .A3(n9069), .A4(n9307), 
        .Y(n3645) );
  AO22X1_HVT U3639 ( .A1(\ram[14][1] ), .A2(n7235), .A3(n9068), .A4(n9310), 
        .Y(n3646) );
  AO22X1_HVT U3640 ( .A1(\ram[14][2] ), .A2(n7232), .A3(n9067), .A4(n9312), 
        .Y(n3647) );
  AO22X1_HVT U3641 ( .A1(\ram[14][3] ), .A2(n4534), .A3(n9068), .A4(n9316), 
        .Y(n3648) );
  AO22X1_HVT U3642 ( .A1(\ram[14][4] ), .A2(n4637), .A3(n9063), .A4(n9320), 
        .Y(n3649) );
  AO22X1_HVT U3643 ( .A1(\ram[14][5] ), .A2(n7223), .A3(n9066), .A4(n9323), 
        .Y(n3650) );
  AO22X1_HVT U3644 ( .A1(\ram[14][6] ), .A2(n7212), .A3(n9066), .A4(n9326), 
        .Y(n3651) );
  AO22X1_HVT U3645 ( .A1(\ram[14][7] ), .A2(n7221), .A3(n9065), .A4(n9329), 
        .Y(n3652) );
  AO22X1_HVT U3646 ( .A1(\ram[14][8] ), .A2(n4638), .A3(n9029), .A4(n9332), 
        .Y(n3653) );
  AO22X1_HVT U3648 ( .A1(\ram[14][10] ), .A2(n4540), .A3(n9048), .A4(n9338), 
        .Y(n3655) );
  AO22X1_HVT U3649 ( .A1(\ram[14][11] ), .A2(n4637), .A3(n9026), .A4(n9341), 
        .Y(n3656) );
  AO22X1_HVT U3650 ( .A1(\ram[14][12] ), .A2(n7221), .A3(n9074), .A4(n9345), 
        .Y(n3657) );
  AO22X1_HVT U3651 ( .A1(\ram[14][13] ), .A2(n7211), .A3(n4278), .A4(n9348), 
        .Y(n3658) );
  AO22X1_HVT U3652 ( .A1(\ram[14][14] ), .A2(n7210), .A3(n9067), .A4(n9351), 
        .Y(n3659) );
  AO22X1_HVT U3653 ( .A1(\ram[14][15] ), .A2(n7222), .A3(n9078), .A4(n9354), 
        .Y(n3660) );
  AO22X1_HVT U3654 ( .A1(\ram[14][16] ), .A2(n7224), .A3(n9060), .A4(n9357), 
        .Y(n3661) );
  AO22X1_HVT U3655 ( .A1(\ram[14][17] ), .A2(n7240), .A3(n9059), .A4(n9360), 
        .Y(n3662) );
  AO22X1_HVT U3656 ( .A1(\ram[14][18] ), .A2(n7242), .A3(n9058), .A4(n9363), 
        .Y(n3663) );
  AO22X1_HVT U3657 ( .A1(\ram[14][19] ), .A2(n7241), .A3(n9057), .A4(n9366), 
        .Y(n3664) );
  AO22X1_HVT U3658 ( .A1(\ram[14][20] ), .A2(n4417), .A3(n9039), .A4(data[20]), 
        .Y(n3665) );
  AO22X1_HVT U3659 ( .A1(\ram[14][21] ), .A2(n7252), .A3(n9032), .A4(n9371), 
        .Y(n3666) );
  AO22X1_HVT U3660 ( .A1(\ram[14][22] ), .A2(n4417), .A3(n9033), .A4(n9374), 
        .Y(n3667) );
  AO22X1_HVT U3661 ( .A1(\ram[14][23] ), .A2(n7251), .A3(n9037), .A4(n9377), 
        .Y(n3668) );
  AO22X1_HVT U3662 ( .A1(\ram[14][24] ), .A2(n4568), .A3(n9080), .A4(n9380), 
        .Y(n3669) );
  AO22X1_HVT U3663 ( .A1(\ram[14][25] ), .A2(n4568), .A3(n4270), .A4(n9383), 
        .Y(n3670) );
  AO22X1_HVT U3664 ( .A1(\ram[14][26] ), .A2(n7257), .A3(n9077), .A4(n9386), 
        .Y(n3671) );
  AO22X1_HVT U3665 ( .A1(\ram[14][27] ), .A2(n7255), .A3(n9077), .A4(n9389), 
        .Y(n3672) );
  AO22X1_HVT U3666 ( .A1(\ram[14][28] ), .A2(n7252), .A3(n9056), .A4(n9392), 
        .Y(n3673) );
  AO22X1_HVT U3667 ( .A1(\ram[14][29] ), .A2(n4197), .A3(n9055), .A4(n9395), 
        .Y(n3674) );
  AO22X1_HVT U3668 ( .A1(\ram[14][30] ), .A2(n7229), .A3(n9054), .A4(data[30]), 
        .Y(n3675) );
  AO22X1_HVT U3669 ( .A1(\ram[14][31] ), .A2(n4417), .A3(n9053), .A4(n9401), 
        .Y(n3676) );
  AO22X1_HVT U3670 ( .A1(\ram[14][32] ), .A2(n4569), .A3(n9029), .A4(n9404), 
        .Y(n3677) );
  AO22X1_HVT U3671 ( .A1(\ram[14][33] ), .A2(n4637), .A3(n9028), .A4(n9407), 
        .Y(n3678) );
  AO22X1_HVT U3672 ( .A1(\ram[14][34] ), .A2(n7209), .A3(n9027), .A4(n9410), 
        .Y(n3679) );
  AO22X1_HVT U3673 ( .A1(\ram[14][35] ), .A2(n7212), .A3(n9026), .A4(n9413), 
        .Y(n3680) );
  AO22X1_HVT U3674 ( .A1(\ram[14][36] ), .A2(n4638), .A3(n4533), .A4(n9416), 
        .Y(n3681) );
  AO22X1_HVT U3675 ( .A1(\ram[14][37] ), .A2(n7222), .A3(n9038), .A4(n9419), 
        .Y(n3682) );
  AO22X1_HVT U3676 ( .A1(\ram[14][38] ), .A2(n7209), .A3(n4531), .A4(n9422), 
        .Y(n3683) );
  AO22X1_HVT U3677 ( .A1(\ram[14][39] ), .A2(n7220), .A3(n9045), .A4(data[39]), 
        .Y(n3684) );
  AO22X1_HVT U3678 ( .A1(\ram[14][40] ), .A2(n7220), .A3(n4533), .A4(n9428), 
        .Y(n3685) );
  AO22X1_HVT U3679 ( .A1(\ram[14][41] ), .A2(n4535), .A3(n9038), .A4(n9431), 
        .Y(n3686) );
  AO22X1_HVT U3680 ( .A1(\ram[14][42] ), .A2(n7227), .A3(n9031), .A4(n9434), 
        .Y(n3687) );
  AO22X1_HVT U3681 ( .A1(\ram[14][43] ), .A2(n7226), .A3(n4610), .A4(n9437), 
        .Y(n3688) );
  AO22X1_HVT U3682 ( .A1(\ram[14][44] ), .A2(n7217), .A3(n9060), .A4(n9440), 
        .Y(n3689) );
  AO22X1_HVT U3683 ( .A1(\ram[14][45] ), .A2(n7216), .A3(n9059), .A4(n9443), 
        .Y(n3690) );
  AO22X1_HVT U3684 ( .A1(\ram[14][46] ), .A2(n7215), .A3(n9058), .A4(n9446), 
        .Y(n3691) );
  AO22X1_HVT U3685 ( .A1(\ram[14][47] ), .A2(n7214), .A3(n9057), .A4(n9449), 
        .Y(n3692) );
  AO22X1_HVT U3687 ( .A1(\ram[14][49] ), .A2(n4540), .A3(n9054), .A4(n9455), 
        .Y(n3694) );
  AO22X1_HVT U3688 ( .A1(\ram[14][50] ), .A2(n4534), .A3(n9053), .A4(n9458), 
        .Y(n3695) );
  AO22X1_HVT U3689 ( .A1(\ram[14][51] ), .A2(n4534), .A3(n9030), .A4(n9461), 
        .Y(n3696) );
  AO22X1_HVT U3690 ( .A1(\ram[14][52] ), .A2(n7234), .A3(n9059), .A4(n9464), 
        .Y(n3697) );
  AO22X1_HVT U3691 ( .A1(\ram[14][53] ), .A2(n7235), .A3(n9038), .A4(n9467), 
        .Y(n3698) );
  AO22X1_HVT U3692 ( .A1(\ram[14][54] ), .A2(n7232), .A3(n9039), .A4(n9470), 
        .Y(n3699) );
  AO22X1_HVT U3694 ( .A1(\ram[14][56] ), .A2(n4195), .A3(n4533), .A4(n9476), 
        .Y(n3701) );
  AO22X1_HVT U3695 ( .A1(\ram[14][57] ), .A2(n4417), .A3(n9070), .A4(n9479), 
        .Y(n3702) );
  AO22X1_HVT U3696 ( .A1(\ram[14][58] ), .A2(n4569), .A3(n9070), .A4(n9482), 
        .Y(n3703) );
  AO22X1_HVT U3697 ( .A1(\ram[14][59] ), .A2(n7250), .A3(n9069), .A4(n9485), 
        .Y(n3704) );
  AO22X1_HVT U3698 ( .A1(\ram[14][60] ), .A2(n7255), .A3(n9068), .A4(n9488), 
        .Y(n3705) );
  AO22X1_HVT U3699 ( .A1(\ram[14][61] ), .A2(n7257), .A3(n4257), .A4(n9491), 
        .Y(n3706) );
  AO22X1_HVT U3700 ( .A1(\ram[14][62] ), .A2(n7258), .A3(n9065), .A4(n9494), 
        .Y(n3707) );
  AO22X1_HVT U3701 ( .A1(\ram[14][63] ), .A2(n7256), .A3(n9063), .A4(n9497), 
        .Y(n3708) );
  AO22X1_HVT U3702 ( .A1(\ram[14][64] ), .A2(n7257), .A3(n9065), .A4(n9500), 
        .Y(n3709) );
  AO22X1_HVT U3703 ( .A1(\ram[14][65] ), .A2(n7256), .A3(n9073), .A4(n9503), 
        .Y(n3710) );
  AO22X1_HVT U3704 ( .A1(\ram[14][66] ), .A2(n4568), .A3(n4278), .A4(n9506), 
        .Y(n3711) );
  AO22X1_HVT U3706 ( .A1(\ram[14][68] ), .A2(n7220), .A3(n9075), .A4(n9512), 
        .Y(n3713) );
  AO22X1_HVT U3707 ( .A1(\ram[14][69] ), .A2(n7211), .A3(n9039), .A4(n9515), 
        .Y(n3714) );
  AO22X1_HVT U3708 ( .A1(\ram[14][70] ), .A2(n7234), .A3(n9032), .A4(n9518), 
        .Y(n3715) );
  AO22X1_HVT U3709 ( .A1(\ram[14][71] ), .A2(n7223), .A3(n9033), .A4(n9521), 
        .Y(n3716) );
  AO22X1_HVT U3710 ( .A1(\ram[14][72] ), .A2(n7211), .A3(n9053), .A4(n9524), 
        .Y(n3717) );
  AO22X1_HVT U3711 ( .A1(\ram[14][73] ), .A2(n7243), .A3(n9044), .A4(n9527), 
        .Y(n3718) );
  AO22X1_HVT U3712 ( .A1(\ram[14][74] ), .A2(n7242), .A3(n9044), .A4(n9530), 
        .Y(n3719) );
  AO22X1_HVT U3713 ( .A1(\ram[14][75] ), .A2(n7241), .A3(n9043), .A4(n9533), 
        .Y(n3720) );
  AO22X1_HVT U3714 ( .A1(\ram[14][76] ), .A2(n7262), .A3(n9042), .A4(n9536), 
        .Y(n3721) );
  AO22X1_HVT U3715 ( .A1(\ram[14][77] ), .A2(n7261), .A3(n9050), .A4(n9539), 
        .Y(n3722) );
  AO22X1_HVT U3716 ( .A1(\ram[14][78] ), .A2(n7260), .A3(n9050), .A4(n9542), 
        .Y(n3723) );
  AO22X1_HVT U3717 ( .A1(\ram[14][79] ), .A2(n7259), .A3(n9048), .A4(n9545), 
        .Y(n3724) );
  AO22X1_HVT U3718 ( .A1(\ram[14][80] ), .A2(n7262), .A3(n9048), .A4(n9548), 
        .Y(n3725) );
  AO22X1_HVT U3719 ( .A1(\ram[14][81] ), .A2(n7261), .A3(n9032), .A4(n9551), 
        .Y(n3726) );
  AO22X1_HVT U3720 ( .A1(\ram[14][82] ), .A2(n7260), .A3(n4611), .A4(n9554), 
        .Y(n3727) );
  AO22X1_HVT U3721 ( .A1(\ram[14][83] ), .A2(n7259), .A3(n9033), .A4(n9557), 
        .Y(n3728) );
  AO22X1_HVT U3722 ( .A1(\ram[14][84] ), .A2(n4497), .A3(n9080), .A4(n9560), 
        .Y(n3729) );
  AO22X1_HVT U3723 ( .A1(\ram[14][85] ), .A2(n7243), .A3(n9080), .A4(n9563), 
        .Y(n3730) );
  AO22X1_HVT U3724 ( .A1(\ram[14][86] ), .A2(n7243), .A3(n9078), .A4(n9566), 
        .Y(n3731) );
  AO22X1_HVT U3725 ( .A1(\ram[14][87] ), .A2(n7237), .A3(n9077), .A4(n9569), 
        .Y(n3732) );
  AO22X1_HVT U3726 ( .A1(\ram[14][88] ), .A2(n7248), .A3(n9077), .A4(n9572), 
        .Y(n3733) );
  AO22X1_HVT U3727 ( .A1(\ram[14][89] ), .A2(n7248), .A3(n9075), .A4(n9575), 
        .Y(n3734) );
  AO22X1_HVT U3728 ( .A1(\ram[14][90] ), .A2(n7246), .A3(n4278), .A4(n9578), 
        .Y(n3735) );
  AO22X1_HVT U3729 ( .A1(\ram[14][91] ), .A2(n4418), .A3(n9079), .A4(n9581), 
        .Y(n3736) );
  AO22X1_HVT U3730 ( .A1(\ram[14][92] ), .A2(n7247), .A3(n9036), .A4(n9584), 
        .Y(n3737) );
  AO22X1_HVT U3731 ( .A1(\ram[14][93] ), .A2(n7247), .A3(n4611), .A4(n9587), 
        .Y(n3738) );
  AO22X1_HVT U3732 ( .A1(\ram[14][94] ), .A2(n4570), .A3(n9050), .A4(n9590), 
        .Y(n3739) );
  AO22X1_HVT U3733 ( .A1(\ram[14][95] ), .A2(n7246), .A3(n9045), .A4(n9593), 
        .Y(n3740) );
  AO22X1_HVT U3734 ( .A1(\ram[14][96] ), .A2(n7210), .A3(n4610), .A4(n9596), 
        .Y(n3741) );
  AO22X1_HVT U3735 ( .A1(\ram[14][97] ), .A2(n7235), .A3(n9045), .A4(n9599), 
        .Y(n3742) );
  AO22X1_HVT U3736 ( .A1(\ram[14][98] ), .A2(n7233), .A3(n9043), .A4(n9602), 
        .Y(n3743) );
  AO22X1_HVT U3737 ( .A1(\ram[14][99] ), .A2(n7232), .A3(n9042), .A4(n9605), 
        .Y(n3744) );
  AO22X1_HVT U3738 ( .A1(\ram[14][100] ), .A2(n7228), .A3(n4531), .A4(n9608), 
        .Y(n3745) );
  AO22X1_HVT U3739 ( .A1(\ram[14][101] ), .A2(n7229), .A3(n9050), .A4(n9611), 
        .Y(n3746) );
  AO22X1_HVT U3741 ( .A1(\ram[14][103] ), .A2(n7226), .A3(n9049), .A4(n9617), 
        .Y(n3748) );
  AO22X1_HVT U3742 ( .A1(\ram[14][104] ), .A2(n4535), .A3(n9060), .A4(n9620), 
        .Y(n3749) );
  AO22X1_HVT U3743 ( .A1(\ram[14][105] ), .A2(n7228), .A3(n9059), .A4(n9623), 
        .Y(n3750) );
  AO22X1_HVT U3744 ( .A1(\ram[14][106] ), .A2(n7227), .A3(n9058), .A4(n9626), 
        .Y(n3751) );
  AO22X1_HVT U3745 ( .A1(\ram[14][107] ), .A2(n7226), .A3(n9057), .A4(n9629), 
        .Y(n3752) );
  AO22X1_HVT U3746 ( .A1(\ram[14][108] ), .A2(n7237), .A3(n9065), .A4(n9632), 
        .Y(n3753) );
  AO22X1_HVT U3747 ( .A1(\ram[14][109] ), .A2(n7240), .A3(n4257), .A4(n9635), 
        .Y(n3754) );
  AO22X1_HVT U3748 ( .A1(\ram[14][110] ), .A2(n7240), .A3(n4257), .A4(n9638), 
        .Y(n3755) );
  AO22X1_HVT U3749 ( .A1(\ram[14][111] ), .A2(n4495), .A3(n9064), .A4(n9641), 
        .Y(n3756) );
  AO22X1_HVT U3750 ( .A1(\ram[14][112] ), .A2(n7221), .A3(n9029), .A4(n9644), 
        .Y(n3757) );
  AO22X1_HVT U3751 ( .A1(\ram[14][113] ), .A2(n7211), .A3(n9028), .A4(n9647), 
        .Y(n3758) );
  AO22X1_HVT U3752 ( .A1(\ram[14][114] ), .A2(n7210), .A3(n9027), .A4(n9650), 
        .Y(n3759) );
  AO22X1_HVT U3753 ( .A1(\ram[14][115] ), .A2(n7223), .A3(n9026), .A4(n9653), 
        .Y(n3760) );
  AO22X1_HVT U3754 ( .A1(\ram[14][116] ), .A2(n7262), .A3(n9074), .A4(n9656), 
        .Y(n3761) );
  AO22X1_HVT U3755 ( .A1(\ram[14][117] ), .A2(n7261), .A3(n9076), .A4(n9659), 
        .Y(n3762) );
  AO22X1_HVT U3756 ( .A1(\ram[14][118] ), .A2(n7260), .A3(n4278), .A4(n9662), 
        .Y(n3763) );
  AO22X1_HVT U3757 ( .A1(\ram[14][119] ), .A2(n7259), .A3(n9074), .A4(n9665), 
        .Y(n3764) );
  AO22X1_HVT U3758 ( .A1(\ram[14][120] ), .A2(n4638), .A3(n4270), .A4(n9668), 
        .Y(n3765) );
  AO22X1_HVT U3759 ( .A1(\ram[14][121] ), .A2(n4499), .A3(n9051), .A4(n9671), 
        .Y(n3766) );
  AO22X1_HVT U3760 ( .A1(\ram[14][122] ), .A2(n7242), .A3(n9051), .A4(n9674), 
        .Y(n3767) );
  AO22X1_HVT U3761 ( .A1(\ram[14][123] ), .A2(n7241), .A3(n9027), .A4(n9677), 
        .Y(n3768) );
  AO22X1_HVT U3762 ( .A1(\ram[14][124] ), .A2(n4540), .A3(n9027), .A4(n9680), 
        .Y(n3769) );
  AO22X1_HVT U3763 ( .A1(\ram[14][125] ), .A2(n7235), .A3(n9029), .A4(n9683), 
        .Y(n3770) );
  AO22X1_HVT U3764 ( .A1(\ram[14][126] ), .A2(n7233), .A3(n9028), .A4(n9686), 
        .Y(n3771) );
  AO22X1_HVT U3765 ( .A1(\ram[14][127] ), .A2(n7233), .A3(n9048), .A4(n9689), 
        .Y(n3772) );
  AO22X1_HVT U3766 ( .A1(\ram[14][128] ), .A2(n4637), .A3(n9026), .A4(n9692), 
        .Y(n3773) );
  AO22X1_HVT U3767 ( .A1(\ram[14][129] ), .A2(n7209), .A3(n9056), .A4(n9695), 
        .Y(n3774) );
  AO22X1_HVT U3768 ( .A1(\ram[14][130] ), .A2(n7212), .A3(n9055), .A4(n9698), 
        .Y(n3775) );
  AO22X1_HVT U3769 ( .A1(\ram[14][131] ), .A2(n7221), .A3(n9054), .A4(n9701), 
        .Y(n3776) );
  AO22X1_HVT U3770 ( .A1(\ram[14][132] ), .A2(n4535), .A3(n4532), .A4(n9704), 
        .Y(n3777) );
  AO22X1_HVT U3771 ( .A1(\ram[14][133] ), .A2(n7228), .A3(n4270), .A4(n9707), 
        .Y(n3778) );
  AO22X1_HVT U3772 ( .A1(\ram[14][134] ), .A2(n4630), .A3(n9079), .A4(n9710), 
        .Y(n3779) );
  AO22X1_HVT U3773 ( .A1(\ram[14][135] ), .A2(n7226), .A3(n9080), .A4(n9713), 
        .Y(n3780) );
  AO22X1_HVT U3774 ( .A1(\ram[14][136] ), .A2(n7246), .A3(n9080), .A4(n9716), 
        .Y(n3781) );
  AO22X1_HVT U3775 ( .A1(\ram[14][137] ), .A2(n7246), .A3(n9074), .A4(n9719), 
        .Y(n3782) );
  AO22X1_HVT U3776 ( .A1(\ram[14][138] ), .A2(n7249), .A3(n9076), .A4(n9722), 
        .Y(n3783) );
  AO22X1_HVT U3777 ( .A1(\ram[14][139] ), .A2(n7248), .A3(n9073), .A4(n9725), 
        .Y(n3784) );
  AO22X1_HVT U3778 ( .A1(\ram[14][140] ), .A2(n7247), .A3(n9076), .A4(n9729), 
        .Y(n3785) );
  AO22X1_HVT U3779 ( .A1(\ram[14][141] ), .A2(n4418), .A3(n9078), .A4(n9732), 
        .Y(n3786) );
  AO22X1_HVT U3780 ( .A1(\ram[14][142] ), .A2(n7246), .A3(n9078), .A4(n9735), 
        .Y(n3787) );
  AO22X1_HVT U3781 ( .A1(\ram[14][143] ), .A2(n7248), .A3(n4270), .A4(n9738), 
        .Y(n3788) );
  AO22X1_HVT U3783 ( .A1(\ram[14][145] ), .A2(n7217), .A3(n9060), .A4(n9745), 
        .Y(n3790) );
  AO22X1_HVT U3784 ( .A1(\ram[14][146] ), .A2(n7216), .A3(n9059), .A4(n9748), 
        .Y(n3791) );
  AO22X1_HVT U3785 ( .A1(\ram[14][147] ), .A2(n7215), .A3(n9058), .A4(n9751), 
        .Y(n3792) );
  AO22X1_HVT U3786 ( .A1(\ram[14][148] ), .A2(n7214), .A3(n9057), .A4(n9755), 
        .Y(n3793) );
  AO22X1_HVT U3787 ( .A1(\ram[14][149] ), .A2(n7262), .A3(n9057), .A4(n9758), 
        .Y(n3794) );
  AO22X1_HVT U3788 ( .A1(\ram[14][150] ), .A2(n7261), .A3(n9056), .A4(n9761), 
        .Y(n3795) );
  AO22X1_HVT U3789 ( .A1(\ram[14][151] ), .A2(n7260), .A3(n9055), .A4(n9764), 
        .Y(n3796) );
  AO22X1_HVT U3790 ( .A1(\ram[14][152] ), .A2(n7259), .A3(n9060), .A4(n9767), 
        .Y(n3797) );
  AO22X1_HVT U3791 ( .A1(\ram[14][153] ), .A2(n7256), .A3(n9031), .A4(n9770), 
        .Y(n3798) );
  AO22X1_HVT U3792 ( .A1(\ram[14][154] ), .A2(n7255), .A3(n9031), .A4(n9773), 
        .Y(n3799) );
  AO22X1_HVT U3793 ( .A1(\ram[14][155] ), .A2(n7256), .A3(n4532), .A4(n9776), 
        .Y(n3800) );
  AO22X1_HVT U3794 ( .A1(\ram[14][156] ), .A2(n7258), .A3(n9029), .A4(n9780), 
        .Y(n3801) );
  AO22X1_HVT U3795 ( .A1(\ram[14][157] ), .A2(n7256), .A3(n9028), .A4(n9783), 
        .Y(n3802) );
  AO22X1_HVT U3796 ( .A1(\ram[14][158] ), .A2(n7257), .A3(n4532), .A4(n9786), 
        .Y(n3803) );
  AO22X1_HVT U3797 ( .A1(\ram[14][159] ), .A2(n4568), .A3(n9026), .A4(n9789), 
        .Y(n3804) );
  AO22X1_HVT U3798 ( .A1(\ram[14][160] ), .A2(n7228), .A3(n9060), .A4(n9793), 
        .Y(n3805) );
  AO22X1_HVT U3799 ( .A1(\ram[14][161] ), .A2(n4535), .A3(n9059), .A4(n9796), 
        .Y(n3806) );
  AO22X1_HVT U3800 ( .A1(\ram[14][162] ), .A2(n4630), .A3(n9058), .A4(n9799), 
        .Y(n3807) );
  AO22X1_HVT U3801 ( .A1(\ram[14][163] ), .A2(n7226), .A3(n9057), .A4(n9802), 
        .Y(n3808) );
  AO22X1_HVT U3802 ( .A1(\ram[14][164] ), .A2(n4495), .A3(n9056), .A4(n9805), 
        .Y(n3809) );
  AO22X1_HVT U3803 ( .A1(\ram[14][165] ), .A2(n7239), .A3(n9055), .A4(n9808), 
        .Y(n3810) );
  AO22X1_HVT U3804 ( .A1(\ram[14][166] ), .A2(n7240), .A3(n9054), .A4(n9811), 
        .Y(n3811) );
  AO22X1_HVT U3805 ( .A1(\ram[14][167] ), .A2(n7238), .A3(n9053), .A4(n9814), 
        .Y(n3812) );
  AO22X1_HVT U3806 ( .A1(\ram[14][168] ), .A2(n7220), .A3(n9037), .A4(n9817), 
        .Y(n3813) );
  AO22X1_HVT U3807 ( .A1(\ram[14][169] ), .A2(n7211), .A3(n4352), .A4(n9820), 
        .Y(n3814) );
  AO22X1_HVT U3808 ( .A1(\ram[14][170] ), .A2(n7234), .A3(n9051), .A4(n9823), 
        .Y(n3815) );
  AO22X1_HVT U3809 ( .A1(\ram[14][171] ), .A2(n7223), .A3(n9030), .A4(n9826), 
        .Y(n3816) );
  AO22X1_HVT U3810 ( .A1(\ram[14][172] ), .A2(n4497), .A3(n9067), .A4(n9830), 
        .Y(n3817) );
  AO22X1_HVT U3811 ( .A1(\ram[14][173] ), .A2(n7239), .A3(n9067), .A4(n9833), 
        .Y(n3818) );
  AO22X1_HVT U3812 ( .A1(\ram[14][174] ), .A2(n7237), .A3(n9069), .A4(n9836), 
        .Y(n3819) );
  AO22X1_HVT U3813 ( .A1(\ram[14][175] ), .A2(n7243), .A3(n9069), .A4(n9839), 
        .Y(n3820) );
  AO22X1_HVT U3814 ( .A1(\ram[14][176] ), .A2(n4497), .A3(n9064), .A4(n9843), 
        .Y(n3821) );
  AO22X1_HVT U3815 ( .A1(\ram[14][177] ), .A2(n7237), .A3(n9064), .A4(n9846), 
        .Y(n3822) );
  AO22X1_HVT U3816 ( .A1(\ram[14][178] ), .A2(n7237), .A3(n9064), .A4(n9849), 
        .Y(n3823) );
  AO22X1_HVT U3817 ( .A1(\ram[14][179] ), .A2(n7243), .A3(n9064), .A4(n9852), 
        .Y(n3824) );
  AO22X1_HVT U3818 ( .A1(\ram[14][180] ), .A2(n7217), .A3(n9045), .A4(n9856), 
        .Y(n3825) );
  AO22X1_HVT U3819 ( .A1(\ram[14][181] ), .A2(n7216), .A3(n9030), .A4(n9859), 
        .Y(n3826) );
  AO22X1_HVT U3820 ( .A1(\ram[14][182] ), .A2(n7215), .A3(n9043), .A4(n9862), 
        .Y(n3827) );
  AO22X1_HVT U3821 ( .A1(\ram[14][183] ), .A2(n7214), .A3(n9042), .A4(n9865), 
        .Y(n3828) );
  AO22X1_HVT U3822 ( .A1(\ram[14][184] ), .A2(n7230), .A3(n4531), .A4(n9869), 
        .Y(n3829) );
  AO22X1_HVT U3823 ( .A1(\ram[14][185] ), .A2(n4499), .A3(n4531), .A4(n9872), 
        .Y(n3830) );
  AO22X1_HVT U3824 ( .A1(\ram[14][186] ), .A2(n7242), .A3(n9049), .A4(n9875), 
        .Y(n3831) );
  AO22X1_HVT U3825 ( .A1(\ram[14][187] ), .A2(n7241), .A3(n9049), .A4(n9878), 
        .Y(n3832) );
  AO22X1_HVT U3826 ( .A1(\ram[14][188] ), .A2(n4497), .A3(n9032), .A4(n9881), 
        .Y(n3833) );
  AO22X1_HVT U3827 ( .A1(\ram[14][189] ), .A2(n4495), .A3(n9039), .A4(n9884), 
        .Y(n3834) );
  AO22X1_HVT U3828 ( .A1(\ram[14][190] ), .A2(n7238), .A3(n9033), .A4(n9887), 
        .Y(n3835) );
  AO22X1_HVT U3829 ( .A1(\ram[14][191] ), .A2(n7240), .A3(n4533), .A4(n9890), 
        .Y(n3836) );
  AO22X1_HVT U3830 ( .A1(\ram[14][192] ), .A2(n7217), .A3(n4257), .A4(n9894), 
        .Y(n3837) );
  AO22X1_HVT U3831 ( .A1(\ram[14][193] ), .A2(n7216), .A3(n9063), .A4(n9897), 
        .Y(n3838) );
  AO22X1_HVT U3832 ( .A1(\ram[14][194] ), .A2(n7215), .A3(n9063), .A4(n9900), 
        .Y(n3839) );
  AO22X1_HVT U3833 ( .A1(\ram[14][195] ), .A2(n7214), .A3(n9066), .A4(n9903), 
        .Y(n3840) );
  AO22X1_HVT U3834 ( .A1(\ram[14][196] ), .A2(n7222), .A3(n9029), .A4(n9907), 
        .Y(n3841) );
  AO22X1_HVT U3835 ( .A1(\ram[14][197] ), .A2(n4499), .A3(n9028), .A4(n9910), 
        .Y(n3842) );
  AO22X1_HVT U3836 ( .A1(\ram[14][198] ), .A2(n7242), .A3(n9049), .A4(n9913), 
        .Y(n3843) );
  AO22X1_HVT U3837 ( .A1(\ram[14][199] ), .A2(n7241), .A3(n9026), .A4(n9916), 
        .Y(n3844) );
  AO22X1_HVT U3838 ( .A1(\ram[14][200] ), .A2(n7225), .A3(n9036), .A4(n9920), 
        .Y(n3845) );
  AO22X1_HVT U3839 ( .A1(\ram[14][201] ), .A2(n7238), .A3(n4611), .A4(n9923), 
        .Y(n3846) );
  AO22X1_HVT U3840 ( .A1(\ram[14][202] ), .A2(n7242), .A3(n9051), .A4(n9926), 
        .Y(n3847) );
  AO22X1_HVT U3841 ( .A1(\ram[14][203] ), .A2(n7241), .A3(n9030), .A4(n9929), 
        .Y(n3848) );
  AO22X1_HVT U3842 ( .A1(\ram[14][204] ), .A2(n7234), .A3(n9073), .A4(n9932), 
        .Y(n3849) );
  AO22X1_HVT U3843 ( .A1(\ram[14][205] ), .A2(n7235), .A3(n9070), .A4(n9935), 
        .Y(n3850) );
  AO22X1_HVT U3844 ( .A1(\ram[14][206] ), .A2(n4534), .A3(n4300), .A4(n9938), 
        .Y(n3851) );
  AO22X1_HVT U3845 ( .A1(\ram[14][207] ), .A2(n7232), .A3(n4300), .A4(n9941), 
        .Y(n3852) );
  AO22X1_HVT U3846 ( .A1(\ram[14][208] ), .A2(n7222), .A3(n4300), .A4(n9945), 
        .Y(n3853) );
  AO22X1_HVT U3847 ( .A1(\ram[14][209] ), .A2(n7209), .A3(n9066), .A4(n9948), 
        .Y(n3854) );
  AO22X1_HVT U3848 ( .A1(\ram[14][210] ), .A2(n7212), .A3(n9066), .A4(n9951), 
        .Y(n3855) );
  AO22X1_HVT U3849 ( .A1(\ram[14][211] ), .A2(n7220), .A3(n9063), .A4(n9954), 
        .Y(n3856) );
  AO22X1_HVT U3850 ( .A1(\ram[14][212] ), .A2(n7229), .A3(n9065), .A4(n9957), 
        .Y(n3857) );
  AO22X1_HVT U3851 ( .A1(\ram[14][213] ), .A2(n7229), .A3(n9044), .A4(n9960), 
        .Y(n3858) );
  AO22X1_HVT U3852 ( .A1(\ram[14][214] ), .A2(n7227), .A3(n9043), .A4(n9963), 
        .Y(n3859) );
  AO22X1_HVT U3853 ( .A1(\ram[14][215] ), .A2(n7226), .A3(n9042), .A4(n9966), 
        .Y(n3860) );
  AO22X1_HVT U3854 ( .A1(\ram[14][216] ), .A2(n7217), .A3(n9037), .A4(n9969), 
        .Y(n3861) );
  AO22X1_HVT U3855 ( .A1(\ram[14][217] ), .A2(n7216), .A3(n9036), .A4(n9972), 
        .Y(n3862) );
  AO22X1_HVT U3856 ( .A1(\ram[14][218] ), .A2(n7215), .A3(n9038), .A4(n9975), 
        .Y(n3863) );
  AO22X1_HVT U3857 ( .A1(\ram[14][219] ), .A2(n7214), .A3(n9031), .A4(n9978), 
        .Y(n3864) );
  AO22X1_HVT U3858 ( .A1(\ram[14][220] ), .A2(n7217), .A3(n9044), .A4(n9982), 
        .Y(n3865) );
  AO22X1_HVT U3859 ( .A1(\ram[14][221] ), .A2(n7216), .A3(n9079), .A4(n9985), 
        .Y(n3866) );
  AO22X1_HVT U3860 ( .A1(\ram[14][222] ), .A2(n7215), .A3(n9079), .A4(n9988), 
        .Y(n3867) );
  AO22X1_HVT U3861 ( .A1(\ram[14][223] ), .A2(n7214), .A3(n9077), .A4(n9991), 
        .Y(n3868) );
  AO22X1_HVT U3862 ( .A1(\ram[14][224] ), .A2(n7255), .A3(n9078), .A4(n9994), 
        .Y(n3869) );
  AO22X1_HVT U3863 ( .A1(\ram[14][225] ), .A2(n7258), .A3(n9076), .A4(n9997), 
        .Y(n3870) );
  AO22X1_HVT U3864 ( .A1(\ram[14][226] ), .A2(n7257), .A3(n9075), .A4(n10000), 
        .Y(n3871) );
  AO22X1_HVT U3865 ( .A1(\ram[14][227] ), .A2(n7258), .A3(n9076), .A4(n10003), 
        .Y(n3872) );
  AO22X1_HVT U3866 ( .A1(\ram[14][228] ), .A2(n7251), .A3(n9056), .A4(n10006), 
        .Y(n3873) );
  AO22X1_HVT U3867 ( .A1(\ram[14][229] ), .A2(n4569), .A3(n9055), .A4(n10009), 
        .Y(n3874) );
  AO22X1_HVT U3868 ( .A1(\ram[14][230] ), .A2(n4195), .A3(n9054), .A4(n10012), 
        .Y(n3875) );
  AO22X1_HVT U3869 ( .A1(\ram[14][231] ), .A2(n7252), .A3(n9053), .A4(n10015), 
        .Y(n3876) );
  AO22X1_HVT U3870 ( .A1(\ram[14][232] ), .A2(n7248), .A3(n9073), .A4(n10019), 
        .Y(n3877) );
  AO22X1_HVT U3871 ( .A1(\ram[14][233] ), .A2(n4570), .A3(n9075), .A4(n10022), 
        .Y(n3878) );
  AO22X1_HVT U3872 ( .A1(\ram[14][234] ), .A2(n7247), .A3(n9075), .A4(n10025), 
        .Y(n3879) );
  AO22X1_HVT U3873 ( .A1(\ram[14][235] ), .A2(n4418), .A3(n9073), .A4(n10028), 
        .Y(n3880) );
  AO22X1_HVT U3874 ( .A1(\ram[14][236] ), .A2(n4569), .A3(n9070), .A4(n10031), 
        .Y(n3881) );
  AO22X1_HVT U3875 ( .A1(\ram[14][237] ), .A2(n7252), .A3(n9068), .A4(n10034), 
        .Y(n3882) );
  AO22X1_HVT U3876 ( .A1(\ram[14][238] ), .A2(n4197), .A3(n9070), .A4(n10037), 
        .Y(n3883) );
  AO22X1_HVT U3877 ( .A1(\ram[14][239] ), .A2(n4195), .A3(n4300), .A4(n10040), 
        .Y(n3884) );
  AO22X1_HVT U3878 ( .A1(\ram[14][240] ), .A2(n7251), .A3(n9056), .A4(n10044), 
        .Y(n3885) );
  AO22X1_HVT U3879 ( .A1(\ram[14][241] ), .A2(n4417), .A3(n9055), .A4(n10047), 
        .Y(n3886) );
  AO22X1_HVT U3880 ( .A1(\ram[14][242] ), .A2(n7250), .A3(n9054), .A4(n10050), 
        .Y(n3887) );
  AO22X1_HVT U3881 ( .A1(\ram[14][243] ), .A2(n7251), .A3(n9053), .A4(n10053), 
        .Y(n3888) );
  AO22X1_HVT U3882 ( .A1(\ram[14][244] ), .A2(n7262), .A3(n4610), .A4(n10056), 
        .Y(n3889) );
  AO22X1_HVT U3883 ( .A1(\ram[14][245] ), .A2(n7261), .A3(n4610), .A4(n10059), 
        .Y(n3890) );
  AO22X1_HVT U3884 ( .A1(\ram[14][246] ), .A2(n7260), .A3(n9043), .A4(n10062), 
        .Y(n3891) );
  AO22X1_HVT U3885 ( .A1(\ram[14][247] ), .A2(n7259), .A3(n9042), .A4(n10065), 
        .Y(n3892) );
  AO22X1_HVT U3886 ( .A1(\ram[14][248] ), .A2(n7223), .A3(n9069), .A4(n10069), 
        .Y(n3893) );
  AO22X1_HVT U3887 ( .A1(\ram[14][249] ), .A2(n7209), .A3(n9068), .A4(n10072), 
        .Y(n3894) );
  AO22X1_HVT U3888 ( .A1(\ram[14][250] ), .A2(n7212), .A3(n9067), .A4(n10075), 
        .Y(n3895) );
  AO22X1_HVT U3889 ( .A1(\ram[14][251] ), .A2(n4638), .A3(n9079), .A4(n10078), 
        .Y(n3896) );
  AO22X1_HVT U3890 ( .A1(\ram[14][252] ), .A2(n4570), .A3(n4352), .A4(n10082), 
        .Y(n3897) );
  AO22X1_HVT U3891 ( .A1(\ram[14][253] ), .A2(n7249), .A3(n4611), .A4(n10085), 
        .Y(n3898) );
  AO22X1_HVT U3892 ( .A1(\ram[14][254] ), .A2(n4570), .A3(n9037), .A4(n10088), 
        .Y(n3899) );
  AO22X1_HVT U3893 ( .A1(\ram[14][255] ), .A2(n7247), .A3(n9036), .A4(n10091), 
        .Y(n3900) );
  AND2X1_HVT U3894 ( .A1(n57), .A2(n5645), .Y(n56) );
  AND2X1_HVT U3896 ( .A1(n5935), .A2(n6644), .Y(n57) );
  AND2X1_HVT U3897 ( .A1(n8801), .A2(n5236), .Y(n17) );
  AO22X1_HVT U3898 ( .A1(\ram[15][0] ), .A2(n5385), .A3(n9013), .A4(n9307), 
        .Y(n3901) );
  AO22X1_HVT U3899 ( .A1(\ram[15][1] ), .A2(n5390), .A3(n9012), .A4(n9310), 
        .Y(n3902) );
  AO22X1_HVT U3900 ( .A1(\ram[15][2] ), .A2(n5413), .A3(n9011), .A4(n9312), 
        .Y(n3903) );
  AO22X1_HVT U3901 ( .A1(\ram[15][3] ), .A2(n5417), .A3(n9010), .A4(n9316), 
        .Y(n3904) );
  AO22X1_HVT U3902 ( .A1(\ram[15][4] ), .A2(n5404), .A3(n9009), .A4(n9320), 
        .Y(n3905) );
  AO22X1_HVT U3903 ( .A1(\ram[15][5] ), .A2(n5392), .A3(n9008), .A4(n9323), 
        .Y(n3906) );
  AO22X1_HVT U3904 ( .A1(\ram[15][6] ), .A2(n5386), .A3(n9007), .A4(n9326), 
        .Y(n3907) );
  AO22X1_HVT U3905 ( .A1(\ram[15][7] ), .A2(n5396), .A3(n9006), .A4(n9329), 
        .Y(n3908) );
  AO22X1_HVT U3906 ( .A1(\ram[15][8] ), .A2(n5416), .A3(n8971), .A4(n9332), 
        .Y(n3909) );
  AO22X1_HVT U3907 ( .A1(\ram[15][9] ), .A2(n5418), .A3(n8970), .A4(n9335), 
        .Y(n3910) );
  AO22X1_HVT U3908 ( .A1(\ram[15][10] ), .A2(n5388), .A3(n8969), .A4(n9338), 
        .Y(n3911) );
  AO22X1_HVT U3909 ( .A1(\ram[15][11] ), .A2(n5391), .A3(n8968), .A4(n9341), 
        .Y(n3912) );
  AO22X1_HVT U3911 ( .A1(\ram[15][13] ), .A2(n5383), .A3(n9012), .A4(n9348), 
        .Y(n3914) );
  AO22X1_HVT U3912 ( .A1(\ram[15][14] ), .A2(n5387), .A3(n9011), .A4(n9351), 
        .Y(n3915) );
  AO22X1_HVT U3913 ( .A1(\ram[15][15] ), .A2(n5421), .A3(n9010), .A4(n9354), 
        .Y(n3916) );
  AO22X1_HVT U3914 ( .A1(\ram[15][16] ), .A2(n5391), .A3(n9003), .A4(n9357), 
        .Y(n3917) );
  AO22X1_HVT U3915 ( .A1(\ram[15][17] ), .A2(n5422), .A3(n9002), .A4(n9360), 
        .Y(n3918) );
  AO22X1_HVT U3916 ( .A1(\ram[15][18] ), .A2(n5400), .A3(n9001), .A4(n9363), 
        .Y(n3919) );
  AO22X1_HVT U3917 ( .A1(\ram[15][19] ), .A2(n5399), .A3(n9000), .A4(n9366), 
        .Y(n3920) );
  AO22X1_HVT U3918 ( .A1(\ram[15][20] ), .A2(n5413), .A3(n9023), .A4(data[20]), 
        .Y(n3921) );
  AO22X1_HVT U3919 ( .A1(\ram[15][21] ), .A2(n5422), .A3(n9022), .A4(n9371), 
        .Y(n3922) );
  AO22X1_HVT U3920 ( .A1(\ram[15][22] ), .A2(n5416), .A3(n9021), .A4(n9374), 
        .Y(n3923) );
  AO22X1_HVT U3921 ( .A1(\ram[15][23] ), .A2(n5389), .A3(n9020), .A4(n9377), 
        .Y(n3924) );
  AO22X1_HVT U3922 ( .A1(\ram[15][24] ), .A2(n5424), .A3(n9019), .A4(n9380), 
        .Y(n3925) );
  AO22X1_HVT U3923 ( .A1(\ram[15][25] ), .A2(n5390), .A3(n9018), .A4(n9383), 
        .Y(n3926) );
  AO22X1_HVT U3927 ( .A1(\ram[15][29] ), .A2(n5410), .A3(n8998), .A4(n9395), 
        .Y(n3930) );
  AO22X1_HVT U3929 ( .A1(\ram[15][31] ), .A2(n6893), .A3(n8996), .A4(n9401), 
        .Y(n3932) );
  AO22X1_HVT U3930 ( .A1(\ram[15][32] ), .A2(n10107), .A3(n8976), .A4(n9404), 
        .Y(n3933) );
  AO22X1_HVT U3931 ( .A1(\ram[15][33] ), .A2(n5394), .A3(n8975), .A4(n9407), 
        .Y(n3934) );
  AO22X1_HVT U3932 ( .A1(\ram[15][34] ), .A2(n5383), .A3(n8974), .A4(n9410), 
        .Y(n3935) );
  AO22X1_HVT U3933 ( .A1(\ram[15][35] ), .A2(n5399), .A3(n8973), .A4(n9413), 
        .Y(n3936) );
  AO22X1_HVT U3934 ( .A1(\ram[15][36] ), .A2(n5392), .A3(n8968), .A4(n9416), 
        .Y(n3937) );
  AO22X1_HVT U3935 ( .A1(\ram[15][37] ), .A2(n5385), .A3(n8976), .A4(n9419), 
        .Y(n3938) );
  AO22X1_HVT U3936 ( .A1(\ram[15][38] ), .A2(n5383), .A3(n8975), .A4(n9422), 
        .Y(n3939) );
  AO22X1_HVT U3937 ( .A1(\ram[15][39] ), .A2(n5424), .A3(n8973), .A4(data[39]), 
        .Y(n3940) );
  AO22X1_HVT U3938 ( .A1(\ram[15][40] ), .A2(n5407), .A3(n8976), .A4(n9428), 
        .Y(n3941) );
  AO22X1_HVT U3939 ( .A1(\ram[15][41] ), .A2(n5418), .A3(n8975), .A4(n9431), 
        .Y(n3942) );
  AO22X1_HVT U3940 ( .A1(\ram[15][42] ), .A2(n5422), .A3(n8974), .A4(n9434), 
        .Y(n3943) );
  AO22X1_HVT U3941 ( .A1(\ram[15][43] ), .A2(n5423), .A3(n8973), .A4(n9437), 
        .Y(n3944) );
  AO22X1_HVT U3942 ( .A1(\ram[15][44] ), .A2(n5419), .A3(n9003), .A4(n9440), 
        .Y(n3945) );
  AO22X1_HVT U3943 ( .A1(\ram[15][45] ), .A2(n5405), .A3(n9002), .A4(n9443), 
        .Y(n3946) );
  AO22X1_HVT U3944 ( .A1(\ram[15][46] ), .A2(n5404), .A3(n9001), .A4(n9446), 
        .Y(n3947) );
  AO22X1_HVT U3945 ( .A1(\ram[15][47] ), .A2(n5409), .A3(n9000), .A4(n9449), 
        .Y(n3948) );
  AO22X1_HVT U3947 ( .A1(\ram[15][49] ), .A2(n5912), .A3(n9009), .A4(n9455), 
        .Y(n3950) );
  AO22X1_HVT U3948 ( .A1(\ram[15][50] ), .A2(n5910), .A3(n9008), .A4(n9458), 
        .Y(n3951) );
  AO22X1_HVT U3949 ( .A1(\ram[15][51] ), .A2(n5918), .A3(n9007), .A4(n9461), 
        .Y(n3952) );
  AO22X1_HVT U3950 ( .A1(\ram[15][52] ), .A2(n5917), .A3(n9006), .A4(n9464), 
        .Y(n3953) );
  AO22X1_HVT U3951 ( .A1(\ram[15][53] ), .A2(n5915), .A3(n9019), .A4(n9467), 
        .Y(n3954) );
  AO22X1_HVT U3952 ( .A1(\ram[15][54] ), .A2(n5917), .A3(n9018), .A4(n9470), 
        .Y(n3955) );
  AO22X1_HVT U3953 ( .A1(\ram[15][55] ), .A2(n5915), .A3(n9017), .A4(n9473), 
        .Y(n3956) );
  AO22X1_HVT U3954 ( .A1(\ram[15][56] ), .A2(n5914), .A3(n9016), .A4(n9476), 
        .Y(n3957) );
  AO22X1_HVT U3955 ( .A1(\ram[15][57] ), .A2(n5911), .A3(n8996), .A4(n9479), 
        .Y(n3958) );
  AO22X1_HVT U3956 ( .A1(\ram[15][58] ), .A2(n5917), .A3(n8981), .A4(n9482), 
        .Y(n3959) );
  AO22X1_HVT U3957 ( .A1(\ram[15][59] ), .A2(n5915), .A3(n8980), .A4(n9485), 
        .Y(n3960) );
  AO22X1_HVT U3958 ( .A1(\ram[15][60] ), .A2(n5390), .A3(n8978), .A4(n9488), 
        .Y(n3961) );
  AO22X1_HVT U3959 ( .A1(\ram[15][61] ), .A2(n5403), .A3(n9023), .A4(n9491), 
        .Y(n3962) );
  AO22X1_HVT U3960 ( .A1(\ram[15][62] ), .A2(n5403), .A3(n9022), .A4(n9494), 
        .Y(n3963) );
  AO22X1_HVT U3961 ( .A1(\ram[15][63] ), .A2(n5398), .A3(n9021), .A4(n9497), 
        .Y(n3964) );
  AO22X1_HVT U3962 ( .A1(\ram[15][64] ), .A2(n10109), .A3(n9020), .A4(n9500), 
        .Y(n3965) );
  AO22X1_HVT U3963 ( .A1(\ram[15][65] ), .A2(n5407), .A3(n8976), .A4(n9503), 
        .Y(n3966) );
  AO22X1_HVT U3964 ( .A1(\ram[15][66] ), .A2(n5408), .A3(n8975), .A4(n9506), 
        .Y(n3967) );
  AO22X1_HVT U3965 ( .A1(\ram[15][67] ), .A2(n5418), .A3(n8974), .A4(n9509), 
        .Y(n3968) );
  AO22X1_HVT U3966 ( .A1(\ram[15][68] ), .A2(n5386), .A3(n8973), .A4(n9512), 
        .Y(n3969) );
  AO22X1_HVT U3967 ( .A1(\ram[15][69] ), .A2(n5414), .A3(n9003), .A4(n9515), 
        .Y(n3970) );
  AO22X1_HVT U3968 ( .A1(\ram[15][70] ), .A2(n5425), .A3(n9002), .A4(n9518), 
        .Y(n3971) );
  AO22X1_HVT U3969 ( .A1(\ram[15][71] ), .A2(n5397), .A3(n9001), .A4(n9521), 
        .Y(n3972) );
  AO22X1_HVT U3970 ( .A1(\ram[15][72] ), .A2(n5407), .A3(n9010), .A4(n9524), 
        .Y(n3973) );
  AO22X1_HVT U3971 ( .A1(\ram[15][73] ), .A2(n5401), .A3(n9009), .A4(n9527), 
        .Y(n3974) );
  AO22X1_HVT U3972 ( .A1(\ram[15][74] ), .A2(n5402), .A3(n9008), .A4(n9530), 
        .Y(n3975) );
  AO22X1_HVT U3974 ( .A1(\ram[15][76] ), .A2(n5400), .A3(n9006), .A4(n9536), 
        .Y(n3977) );
  AO22X1_HVT U3975 ( .A1(\ram[15][77] ), .A2(n5402), .A3(n8971), .A4(n9539), 
        .Y(n3978) );
  AO22X1_HVT U3976 ( .A1(\ram[15][78] ), .A2(n5391), .A3(n8970), .A4(n9542), 
        .Y(n3979) );
  AO22X1_HVT U3977 ( .A1(\ram[15][79] ), .A2(n5403), .A3(n8969), .A4(n9545), 
        .Y(n3980) );
  AO22X1_HVT U3978 ( .A1(\ram[15][80] ), .A2(n5423), .A3(n8968), .A4(n9548), 
        .Y(n3981) );
  AO22X1_HVT U3979 ( .A1(\ram[15][81] ), .A2(n6893), .A3(n8981), .A4(n9551), 
        .Y(n3982) );
  AO22X1_HVT U3980 ( .A1(\ram[15][82] ), .A2(n5397), .A3(n8980), .A4(n9554), 
        .Y(n3983) );
  AO22X1_HVT U3982 ( .A1(\ram[15][84] ), .A2(n5420), .A3(n8999), .A4(n9560), 
        .Y(n3985) );
  AO22X1_HVT U3983 ( .A1(\ram[15][85] ), .A2(n10107), .A3(n8998), .A4(n9563), 
        .Y(n3986) );
  AO22X1_HVT U3984 ( .A1(\ram[15][86] ), .A2(n5412), .A3(n8997), .A4(n9566), 
        .Y(n3987) );
  AO22X1_HVT U3985 ( .A1(\ram[15][87] ), .A2(n5400), .A3(n8996), .A4(n9569), 
        .Y(n3988) );
  AO22X1_HVT U3986 ( .A1(\ram[15][88] ), .A2(n5423), .A3(n9003), .A4(n9572), 
        .Y(n3989) );
  AO22X1_HVT U3987 ( .A1(\ram[15][89] ), .A2(n5405), .A3(n9002), .A4(n9575), 
        .Y(n3990) );
  AO22X1_HVT U3988 ( .A1(\ram[15][90] ), .A2(n6893), .A3(n9001), .A4(n9578), 
        .Y(n3991) );
  AO22X1_HVT U3989 ( .A1(\ram[15][91] ), .A2(n5420), .A3(n9000), .A4(n9581), 
        .Y(n3992) );
  AO22X1_HVT U3990 ( .A1(\ram[15][92] ), .A2(n5391), .A3(n8993), .A4(n9584), 
        .Y(n3993) );
  AO22X1_HVT U3991 ( .A1(\ram[15][93] ), .A2(n5396), .A3(n8992), .A4(n9587), 
        .Y(n3994) );
  AO22X1_HVT U3992 ( .A1(\ram[15][94] ), .A2(n5384), .A3(n8991), .A4(n9590), 
        .Y(n3995) );
  AO22X1_HVT U3993 ( .A1(\ram[15][95] ), .A2(n5393), .A3(n8990), .A4(n9593), 
        .Y(n3996) );
  AO22X1_HVT U3994 ( .A1(\ram[15][96] ), .A2(n5398), .A3(n8999), .A4(n9596), 
        .Y(n3997) );
  AO22X1_HVT U3995 ( .A1(\ram[15][97] ), .A2(n5407), .A3(n8998), .A4(n9599), 
        .Y(n3998) );
  AO22X1_HVT U3996 ( .A1(\ram[15][98] ), .A2(n5423), .A3(n8997), .A4(n9602), 
        .Y(n3999) );
  AO22X1_HVT U3997 ( .A1(\ram[15][99] ), .A2(n5403), .A3(n8996), .A4(n9605), 
        .Y(n4000) );
  AO22X1_HVT U3998 ( .A1(\ram[15][100] ), .A2(n5404), .A3(n9013), .A4(n9608), 
        .Y(n4001) );
  AO22X1_HVT U3999 ( .A1(\ram[15][101] ), .A2(n5421), .A3(n9012), .A4(n9611), 
        .Y(n4002) );
  AO22X1_HVT U4000 ( .A1(\ram[15][102] ), .A2(n5401), .A3(n9011), .A4(n9614), 
        .Y(n4003) );
  AO22X1_HVT U4002 ( .A1(\ram[15][104] ), .A2(n10100), .A3(n9009), .A4(n9620), 
        .Y(n4005) );
  AO22X1_HVT U4003 ( .A1(\ram[15][105] ), .A2(n5385), .A3(n9008), .A4(n9623), 
        .Y(n4006) );
  AO22X1_HVT U4004 ( .A1(\ram[15][106] ), .A2(n5406), .A3(n9007), .A4(n9626), 
        .Y(n4007) );
  AO22X1_HVT U4005 ( .A1(\ram[15][107] ), .A2(n5414), .A3(n9006), .A4(n9629), 
        .Y(n4008) );
  AO22X1_HVT U4006 ( .A1(\ram[15][108] ), .A2(n5422), .A3(n8999), .A4(n9632), 
        .Y(n4009) );
  AO22X1_HVT U4007 ( .A1(\ram[15][109] ), .A2(n10106), .A3(n8998), .A4(n9635), 
        .Y(n4010) );
  AO22X1_HVT U4008 ( .A1(\ram[15][110] ), .A2(n5392), .A3(n8997), .A4(n9638), 
        .Y(n4011) );
  AO22X1_HVT U4009 ( .A1(\ram[15][111] ), .A2(n5405), .A3(n8996), .A4(n9641), 
        .Y(n4012) );
  AO22X1_HVT U4010 ( .A1(\ram[15][112] ), .A2(n5390), .A3(n8981), .A4(n9644), 
        .Y(n4013) );
  AO22X1_HVT U4011 ( .A1(\ram[15][113] ), .A2(n5394), .A3(n8980), .A4(n9647), 
        .Y(n4014) );
  AO22X1_HVT U4012 ( .A1(\ram[15][114] ), .A2(n5422), .A3(n8979), .A4(n9650), 
        .Y(n4015) );
  AO22X1_HVT U4013 ( .A1(\ram[15][115] ), .A2(n5415), .A3(n8978), .A4(n9653), 
        .Y(n4016) );
  AO22X1_HVT U4014 ( .A1(\ram[15][116] ), .A2(n5399), .A3(n9009), .A4(n9656), 
        .Y(n4017) );
  AO22X1_HVT U4015 ( .A1(\ram[15][117] ), .A2(n10103), .A3(n9008), .A4(n9659), 
        .Y(n4018) );
  AO22X1_HVT U4016 ( .A1(\ram[15][118] ), .A2(n5414), .A3(n9007), .A4(n9662), 
        .Y(n4019) );
  AO22X1_HVT U4017 ( .A1(\ram[15][119] ), .A2(n5385), .A3(n9006), .A4(n9665), 
        .Y(n4020) );
  AO22X1_HVT U4018 ( .A1(\ram[15][120] ), .A2(n5917), .A3(n8993), .A4(n9668), 
        .Y(n4021) );
  AO22X1_HVT U4019 ( .A1(\ram[15][121] ), .A2(n5918), .A3(n8992), .A4(n9671), 
        .Y(n4022) );
  AO22X1_HVT U4020 ( .A1(\ram[15][122] ), .A2(n5912), .A3(n8991), .A4(n9674), 
        .Y(n4023) );
  AO22X1_HVT U4021 ( .A1(\ram[15][123] ), .A2(n5911), .A3(n8990), .A4(n9677), 
        .Y(n4024) );
  AO22X1_HVT U4022 ( .A1(\ram[15][124] ), .A2(n5910), .A3(n8987), .A4(n9680), 
        .Y(n4025) );
  AO22X1_HVT U4023 ( .A1(\ram[15][125] ), .A2(n5918), .A3(n8986), .A4(n9683), 
        .Y(n4026) );
  AO22X1_HVT U4024 ( .A1(\ram[15][126] ), .A2(n5915), .A3(n8985), .A4(n9686), 
        .Y(n4027) );
  AO22X1_HVT U4025 ( .A1(\ram[15][127] ), .A2(n5914), .A3(n8984), .A4(n9689), 
        .Y(n4028) );
  AO22X1_HVT U4026 ( .A1(\ram[15][128] ), .A2(n5911), .A3(n9023), .A4(n9692), 
        .Y(n4029) );
  AO22X1_HVT U4027 ( .A1(\ram[15][129] ), .A2(n5917), .A3(n9022), .A4(n9695), 
        .Y(n4030) );
  AO22X1_HVT U4028 ( .A1(\ram[15][130] ), .A2(n5910), .A3(n9021), .A4(n9698), 
        .Y(n4031) );
  AO22X1_HVT U4029 ( .A1(\ram[15][131] ), .A2(n5918), .A3(n9020), .A4(n9701), 
        .Y(n4032) );
  AO22X1_HVT U4030 ( .A1(\ram[15][132] ), .A2(n5398), .A3(n8987), .A4(n9704), 
        .Y(n4033) );
  AO22X1_HVT U4031 ( .A1(\ram[15][133] ), .A2(n5425), .A3(n8986), .A4(n9707), 
        .Y(n4034) );
  AO22X1_HVT U4032 ( .A1(\ram[15][134] ), .A2(n5395), .A3(n8985), .A4(n9710), 
        .Y(n4035) );
  AO22X1_HVT U4033 ( .A1(\ram[15][135] ), .A2(n5401), .A3(n8984), .A4(n9713), 
        .Y(n4036) );
  AO22X1_HVT U4034 ( .A1(\ram[15][136] ), .A2(n5421), .A3(n9023), .A4(n9716), 
        .Y(n4037) );
  AO22X1_HVT U4035 ( .A1(\ram[15][137] ), .A2(n5409), .A3(n9022), .A4(n9719), 
        .Y(n4038) );
  AO22X1_HVT U4036 ( .A1(\ram[15][138] ), .A2(n5408), .A3(n9021), .A4(n9722), 
        .Y(n4039) );
  AO22X1_HVT U4037 ( .A1(\ram[15][139] ), .A2(n10105), .A3(n9020), .A4(n9725), 
        .Y(n4040) );
  AO22X1_HVT U4038 ( .A1(\ram[15][140] ), .A2(n5415), .A3(n8987), .A4(n9729), 
        .Y(n4041) );
  AO22X1_HVT U4039 ( .A1(\ram[15][141] ), .A2(n5420), .A3(n8986), .A4(n9732), 
        .Y(n4042) );
  AO22X1_HVT U4040 ( .A1(\ram[15][142] ), .A2(n5399), .A3(n8985), .A4(
        data[142]), .Y(n4043) );
  AO22X1_HVT U4041 ( .A1(\ram[15][143] ), .A2(n5395), .A3(n8984), .A4(n9738), 
        .Y(n4044) );
  AO22X1_HVT U4042 ( .A1(\ram[15][144] ), .A2(n5411), .A3(n8993), .A4(n9742), 
        .Y(n4045) );
  AO22X1_HVT U4043 ( .A1(\ram[15][145] ), .A2(n5419), .A3(n8992), .A4(n9745), 
        .Y(n4046) );
  AO22X1_HVT U4044 ( .A1(\ram[15][146] ), .A2(n5403), .A3(n8991), .A4(n9748), 
        .Y(n4047) );
  AO22X1_HVT U4045 ( .A1(\ram[15][147] ), .A2(n10100), .A3(n8990), .A4(n9751), 
        .Y(n4048) );
  AO22X1_HVT U4047 ( .A1(\ram[15][149] ), .A2(n6760), .A3(n9012), .A4(n9758), 
        .Y(n4050) );
  AO22X1_HVT U4048 ( .A1(\ram[15][150] ), .A2(n5387), .A3(n9011), .A4(n9761), 
        .Y(n4051) );
  AO22X1_HVT U4049 ( .A1(\ram[15][151] ), .A2(n5388), .A3(n9010), .A4(n9764), 
        .Y(n4052) );
  AO22X1_HVT U4051 ( .A1(\ram[15][153] ), .A2(n5386), .A3(n8980), .A4(n9770), 
        .Y(n4054) );
  AO22X1_HVT U4052 ( .A1(\ram[15][154] ), .A2(n5389), .A3(n8979), .A4(n9773), 
        .Y(n4055) );
  AO22X1_HVT U4053 ( .A1(\ram[15][155] ), .A2(n5384), .A3(n8978), .A4(n9776), 
        .Y(n4056) );
  AO22X1_HVT U4054 ( .A1(\ram[15][156] ), .A2(n5420), .A3(n9023), .A4(n9780), 
        .Y(n4057) );
  AO22X1_HVT U4055 ( .A1(\ram[15][157] ), .A2(n5393), .A3(n9022), .A4(n9783), 
        .Y(n4058) );
  AO22X1_HVT U4056 ( .A1(\ram[15][158] ), .A2(n5417), .A3(n9021), .A4(n9786), 
        .Y(n4059) );
  AO22X1_HVT U4057 ( .A1(\ram[15][159] ), .A2(n5416), .A3(n9020), .A4(n9789), 
        .Y(n4060) );
  AO22X1_HVT U4058 ( .A1(\ram[15][160] ), .A2(n5387), .A3(n9019), .A4(n9793), 
        .Y(n4061) );
  AO22X1_HVT U4059 ( .A1(\ram[15][161] ), .A2(n5402), .A3(n9018), .A4(n9796), 
        .Y(n4062) );
  AO22X1_HVT U4060 ( .A1(\ram[15][162] ), .A2(n5401), .A3(n9017), .A4(n9799), 
        .Y(n4063) );
  AO22X1_HVT U4061 ( .A1(\ram[15][163] ), .A2(n5396), .A3(n9016), .A4(n9802), 
        .Y(n4064) );
  AO22X1_HVT U4062 ( .A1(\ram[15][164] ), .A2(n10110), .A3(n8976), .A4(n9805), 
        .Y(n4065) );
  AO22X1_HVT U4063 ( .A1(\ram[15][165] ), .A2(n5398), .A3(n8975), .A4(n9808), 
        .Y(n4066) );
  AO22X1_HVT U4064 ( .A1(\ram[15][166] ), .A2(n5388), .A3(n8974), .A4(n9811), 
        .Y(n4067) );
  AO22X1_HVT U4065 ( .A1(\ram[15][167] ), .A2(n5392), .A3(n8973), .A4(n9814), 
        .Y(n4068) );
  AO22X1_HVT U4066 ( .A1(\ram[15][168] ), .A2(n5411), .A3(n8993), .A4(n9817), 
        .Y(n4069) );
  AO22X1_HVT U4067 ( .A1(\ram[15][169] ), .A2(n5408), .A3(n8992), .A4(n9820), 
        .Y(n4070) );
  AO22X1_HVT U4068 ( .A1(\ram[15][170] ), .A2(n5389), .A3(n8991), .A4(n9823), 
        .Y(n4071) );
  AO22X1_HVT U4069 ( .A1(\ram[15][171] ), .A2(n5405), .A3(n8990), .A4(n9826), 
        .Y(n4072) );
  AO22X1_HVT U4070 ( .A1(\ram[15][172] ), .A2(n5397), .A3(n8987), .A4(n9830), 
        .Y(n4073) );
  AO22X1_HVT U4071 ( .A1(\ram[15][173] ), .A2(n5419), .A3(n8986), .A4(n9833), 
        .Y(n4074) );
  AO22X1_HVT U4072 ( .A1(\ram[15][174] ), .A2(n5409), .A3(n8985), .A4(n9836), 
        .Y(n4075) );
  AO22X1_HVT U4073 ( .A1(\ram[15][175] ), .A2(n5412), .A3(n8984), .A4(n9839), 
        .Y(n4076) );
  AO22X1_HVT U4074 ( .A1(\ram[15][176] ), .A2(n6764), .A3(n9003), .A4(n9843), 
        .Y(n4077) );
  AO22X1_HVT U4075 ( .A1(\ram[15][177] ), .A2(n5416), .A3(n9002), .A4(n9846), 
        .Y(n4078) );
  AO22X1_HVT U4076 ( .A1(\ram[15][178] ), .A2(n5399), .A3(n9001), .A4(n9849), 
        .Y(n4079) );
  AO22X1_HVT U4077 ( .A1(\ram[15][179] ), .A2(n5749), .A3(n9000), .A4(n9852), 
        .Y(n4080) );
  AO22X1_HVT U4078 ( .A1(\ram[15][180] ), .A2(n5406), .A3(n8971), .A4(n9856), 
        .Y(n4081) );
  AO22X1_HVT U4079 ( .A1(\ram[15][181] ), .A2(n5407), .A3(n8970), .A4(n9859), 
        .Y(n4082) );
  AO22X1_HVT U4080 ( .A1(\ram[15][182] ), .A2(n5390), .A3(n8969), .A4(n9862), 
        .Y(n4083) );
  AO22X1_HVT U4081 ( .A1(\ram[15][183] ), .A2(n5384), .A3(n8968), .A4(n9865), 
        .Y(n4084) );
  AO22X1_HVT U4082 ( .A1(\ram[15][184] ), .A2(n5413), .A3(n8971), .A4(n9869), 
        .Y(n4085) );
  AO22X1_HVT U4083 ( .A1(\ram[15][185] ), .A2(n5410), .A3(n8970), .A4(n9872), 
        .Y(n4086) );
  AO22X1_HVT U4084 ( .A1(\ram[15][186] ), .A2(n5419), .A3(n8969), .A4(n9875), 
        .Y(n4087) );
  AO22X1_HVT U4085 ( .A1(\ram[15][187] ), .A2(n5409), .A3(n8974), .A4(n9878), 
        .Y(n4088) );
  AO22X1_HVT U4086 ( .A1(\ram[15][188] ), .A2(n10098), .A3(n9019), .A4(n9881), 
        .Y(n4089) );
  AO22X1_HVT U4087 ( .A1(\ram[15][189] ), .A2(n6764), .A3(n9018), .A4(n9884), 
        .Y(n4090) );
  AO22X1_HVT U4088 ( .A1(\ram[15][190] ), .A2(n5424), .A3(n9017), .A4(n9887), 
        .Y(n4091) );
  AO22X1_HVT U4089 ( .A1(\ram[15][191] ), .A2(n5401), .A3(n9016), .A4(n9890), 
        .Y(n4092) );
  AO22X1_HVT U4090 ( .A1(\ram[15][192] ), .A2(n5393), .A3(n9020), .A4(n9894), 
        .Y(n4093) );
  AO22X1_HVT U4091 ( .A1(\ram[15][193] ), .A2(n5394), .A3(n8999), .A4(n9897), 
        .Y(n4094) );
  AO22X1_HVT U4092 ( .A1(\ram[15][194] ), .A2(n5408), .A3(n8998), .A4(n9900), 
        .Y(n4095) );
  AO22X1_HVT U4093 ( .A1(\ram[15][195] ), .A2(n5417), .A3(n8997), .A4(n9903), 
        .Y(n4096) );
  AO22X1_HVT U4094 ( .A1(\ram[15][196] ), .A2(n10104), .A3(n8979), .A4(n9907), 
        .Y(n4097) );
  AO22X1_HVT U4095 ( .A1(\ram[15][197] ), .A2(n5397), .A3(n9019), .A4(n9910), 
        .Y(n4098) );
  AO22X1_HVT U4096 ( .A1(\ram[15][198] ), .A2(n6893), .A3(n9018), .A4(n9913), 
        .Y(n4099) );
  AO22X1_HVT U4097 ( .A1(\ram[15][199] ), .A2(n5423), .A3(n9017), .A4(n9916), 
        .Y(n4100) );
  AO22X1_HVT U4098 ( .A1(\ram[15][200] ), .A2(n10102), .A3(n9016), .A4(n9920), 
        .Y(n4101) );
  AO22X1_HVT U4099 ( .A1(\ram[15][201] ), .A2(n5412), .A3(n9013), .A4(n9923), 
        .Y(n4102) );
  AO22X1_HVT U4100 ( .A1(\ram[15][202] ), .A2(n5410), .A3(n9012), .A4(n9926), 
        .Y(n4103) );
  AO22X1_HVT U4101 ( .A1(\ram[15][203] ), .A2(n5404), .A3(n9011), .A4(n9929), 
        .Y(n4104) );
  AO22X1_HVT U4104 ( .A1(\ram[15][206] ), .A2(n5389), .A3(n8970), .A4(n9938), 
        .Y(n4107) );
  AO22X1_HVT U4105 ( .A1(\ram[15][207] ), .A2(n5386), .A3(n8969), .A4(n9941), 
        .Y(n4108) );
  AO22X1_HVT U4106 ( .A1(\ram[15][208] ), .A2(n5395), .A3(n8968), .A4(n9945), 
        .Y(n4109) );
  AO22X1_HVT U4107 ( .A1(\ram[15][209] ), .A2(n10104), .A3(n9013), .A4(n9948), 
        .Y(n4110) );
  AO22X1_HVT U4108 ( .A1(\ram[15][210] ), .A2(n5417), .A3(n9012), .A4(n9951), 
        .Y(n4111) );
  AO22X1_HVT U4109 ( .A1(\ram[15][211] ), .A2(n5387), .A3(n9011), .A4(n9954), 
        .Y(n4112) );
  AO22X1_HVT U4110 ( .A1(\ram[15][212] ), .A2(n10098), .A3(n9010), .A4(n9957), 
        .Y(n4113) );
  AO22X1_HVT U4111 ( .A1(\ram[15][213] ), .A2(n5415), .A3(n9023), .A4(n9960), 
        .Y(n4114) );
  AO22X1_HVT U4112 ( .A1(\ram[15][214] ), .A2(n5396), .A3(n9022), .A4(n9963), 
        .Y(n4115) );
  AO22X1_HVT U4113 ( .A1(\ram[15][215] ), .A2(n10103), .A3(n9021), .A4(n9966), 
        .Y(n4116) );
  AO22X1_HVT U4115 ( .A1(\ram[15][217] ), .A2(n5914), .A3(n8999), .A4(n9972), 
        .Y(n4118) );
  AO22X1_HVT U4116 ( .A1(\ram[15][218] ), .A2(n5912), .A3(n8998), .A4(n9975), 
        .Y(n4119) );
  AO22X1_HVT U4117 ( .A1(\ram[15][219] ), .A2(n10099), .A3(n8997), .A4(n9978), 
        .Y(n4120) );
  AO22X1_HVT U4118 ( .A1(\ram[15][220] ), .A2(n5912), .A3(n8996), .A4(n9982), 
        .Y(n4121) );
  AO22X1_HVT U4119 ( .A1(\ram[15][221] ), .A2(n5911), .A3(n8987), .A4(n9985), 
        .Y(n4122) );
  AO22X1_HVT U4120 ( .A1(\ram[15][222] ), .A2(n5910), .A3(n8986), .A4(n9988), 
        .Y(n4123) );
  AO22X1_HVT U4121 ( .A1(\ram[15][223] ), .A2(n5914), .A3(n8985), .A4(n9991), 
        .Y(n4124) );
  AO22X1_HVT U4122 ( .A1(\ram[15][224] ), .A2(n5915), .A3(n8984), .A4(n9994), 
        .Y(n4125) );
  AO22X1_HVT U4123 ( .A1(\ram[15][225] ), .A2(n5912), .A3(n9009), .A4(n9997), 
        .Y(n4126) );
  AO22X1_HVT U4124 ( .A1(\ram[15][226] ), .A2(n5911), .A3(n9008), .A4(n10000), 
        .Y(n4127) );
  AO22X1_HVT U4125 ( .A1(\ram[15][227] ), .A2(n5910), .A3(n9007), .A4(n10003), 
        .Y(n4128) );
  AO22X1_HVT U4126 ( .A1(\ram[15][228] ), .A2(n5411), .A3(n8971), .A4(n10006), 
        .Y(n4129) );
  AO22X1_HVT U4127 ( .A1(\ram[15][229] ), .A2(n5408), .A3(n8970), .A4(n10009), 
        .Y(n4130) );
  AO22X1_HVT U4128 ( .A1(\ram[15][230] ), .A2(n5411), .A3(n8969), .A4(n10012), 
        .Y(n4131) );
  AO22X1_HVT U4129 ( .A1(\ram[15][231] ), .A2(n5391), .A3(n8968), .A4(n10015), 
        .Y(n4132) );
  AO22X1_HVT U4130 ( .A1(\ram[15][232] ), .A2(n5388), .A3(n8976), .A4(n10019), 
        .Y(n4133) );
  AO22X1_HVT U4131 ( .A1(\ram[15][233] ), .A2(n5415), .A3(n8975), .A4(n10022), 
        .Y(n4134) );
  AO22X1_HVT U4132 ( .A1(\ram[15][234] ), .A2(n5420), .A3(n8974), .A4(n10025), 
        .Y(n4135) );
  AO22X1_HVT U4133 ( .A1(\ram[15][235] ), .A2(n5400), .A3(n8973), .A4(n10028), 
        .Y(n4136) );
  AO22X1_HVT U4134 ( .A1(\ram[15][236] ), .A2(n5410), .A3(n9003), .A4(n10031), 
        .Y(n4137) );
  AO22X1_HVT U4135 ( .A1(\ram[15][237] ), .A2(n5397), .A3(n9002), .A4(n10034), 
        .Y(n4138) );
  AO22X1_HVT U4136 ( .A1(\ram[15][238] ), .A2(n5424), .A3(n9001), .A4(n10037), 
        .Y(n4139) );
  AO22X1_HVT U4137 ( .A1(\ram[15][239] ), .A2(n5414), .A3(n9000), .A4(n10040), 
        .Y(n4140) );
  AO22X1_HVT U4139 ( .A1(\ram[15][241] ), .A2(n5389), .A3(n8980), .A4(n10047), 
        .Y(n4142) );
  AO22X1_HVT U4140 ( .A1(\ram[15][242] ), .A2(n5412), .A3(n8979), .A4(n10050), 
        .Y(n4143) );
  AO22X1_HVT U4141 ( .A1(\ram[15][243] ), .A2(n5398), .A3(n8978), .A4(n10053), 
        .Y(n4144) );
  AO22X1_HVT U4142 ( .A1(\ram[15][244] ), .A2(n5400), .A3(n8993), .A4(n10056), 
        .Y(n4145) );
  AO22X1_HVT U4143 ( .A1(\ram[15][245] ), .A2(n5424), .A3(n8992), .A4(n10059), 
        .Y(n4146) );
  AO22X1_HVT U4144 ( .A1(\ram[15][246] ), .A2(n5384), .A3(n8991), .A4(n10062), 
        .Y(n4147) );
  AO22X1_HVT U4146 ( .A1(\ram[15][248] ), .A2(n5425), .A3(n8987), .A4(n10069), 
        .Y(n4149) );
  AO22X1_HVT U4147 ( .A1(\ram[15][249] ), .A2(n5402), .A3(n8986), .A4(n10072), 
        .Y(n4150) );
  AO22X1_HVT U4148 ( .A1(\ram[15][250] ), .A2(n5385), .A3(n8985), .A4(n10075), 
        .Y(n4151) );
  AO22X1_HVT U4149 ( .A1(\ram[15][251] ), .A2(n5421), .A3(n8984), .A4(n10078), 
        .Y(n4152) );
  AO22X1_HVT U4150 ( .A1(\ram[15][252] ), .A2(n10102), .A3(n9019), .A4(n10082), 
        .Y(n4153) );
  AO22X1_HVT U4151 ( .A1(\ram[15][253] ), .A2(n5409), .A3(n9018), .A4(n10085), 
        .Y(n4154) );
  AO22X1_HVT U4152 ( .A1(\ram[15][254] ), .A2(n5387), .A3(n9017), .A4(n10088), 
        .Y(n4155) );
  AO22X1_HVT U4153 ( .A1(\ram[15][255] ), .A2(n5418), .A3(n9016), .A4(n10091), 
        .Y(n4156) );
  AND2X1_HVT U4154 ( .A1(n60), .A2(n10377), .Y(n59) );
  INVX0_HVT U3 ( .A(n5608), .Y(n4918) );
  INVX1_HVT U4 ( .A(n5336), .Y(n5512) );
  MUX41X1_HVT U5 ( .A1(n8283), .A3(n8285), .A2(n8282), .A4(n8284), .S0(n7567), 
        .S1(n1), .Y(q[138]) );
  IBUFFX16_HVT U6 ( .A(n5631), .Y(n1) );
  MUX41X1_HVT U9 ( .A1(\ram[10][185] ), .A3(\ram[8][185] ), .A2(\ram[11][185] ), .A4(\ram[9][185] ), .S0(n3), .S1(n6738), .Y(n8470) );
  IBUFFX2_HVT U27 ( .A(n8788), .Y(n8810) );
  INVX1_HVT U57 ( .A(n2), .Y(n3) );
  IBUFFX2_HVT U110 ( .A(n5345), .Y(n5346) );
  INVX0_HVT U131 ( .A(n5346), .Y(n5447) );
  INVX0_HVT U151 ( .A(n5346), .Y(n6411) );
  INVX0_HVT U263 ( .A(n5346), .Y(n4982) );
  INVX0_HVT U264 ( .A(n5314), .Y(n5457) );
  INVX0_HVT U276 ( .A(n5314), .Y(n43) );
  INVX0_HVT U284 ( .A(n6003), .Y(n2) );
  IBUFFX2_HVT U295 ( .A(n7343), .Y(n6003) );
  MUX41X1_HVT U306 ( .A1(n8551), .A3(n8552), .A2(n8549), .A4(n8550), .S0(n5737), .S1(n5654), .Y(q[205]) );
  MUX41X2_HVT U308 ( .A1(\ram[11][205] ), .A3(\ram[9][205] ), .A2(
        \ram[10][205] ), .A4(\ram[8][205] ), .S0(n5976), .S1(n7294), .Y(n8550)
         );
  IBUFFX2_HVT U311 ( .A(n6131), .Y(n6006) );
  MUX41X1_HVT U314 ( .A1(\ram[11][236] ), .A3(\ram[9][236] ), .A2(
        \ram[10][236] ), .A4(\ram[8][236] ), .S0(n5968), .S1(n4165), .Y(n8672)
         );
  IBUFFX2_HVT U352 ( .A(n6663), .Y(n7700) );
  IBUFFX2_HVT U354 ( .A(n5987), .Y(n5972) );
  INVX0_HVT U386 ( .A(n6765), .Y(n5796) );
  MUX41X1_HVT U388 ( .A1(n8715), .A3(n8717), .A2(n8716), .A4(n8718), .S0(n4), 
        .S1(n5), .Y(q[247]) );
  IBUFFX16_HVT U434 ( .A(n5323), .Y(n4) );
  IBUFFX16_HVT U510 ( .A(n8767), .Y(n5) );
  INVX0_HVT U518 ( .A(n8833), .Y(n7277) );
  IBUFFX2_HVT U522 ( .A(n8833), .Y(n5741) );
  MUX41X1_HVT U523 ( .A1(\ram[11][189] ), .A3(\ram[9][189] ), .A2(
        \ram[10][189] ), .A4(\ram[8][189] ), .S0(n6), .S1(n4888), .Y(n8486) );
  IBUFFX16_HVT U532 ( .A(n6018), .Y(n6) );
  INVX0_HVT U573 ( .A(n6126), .Y(n6965) );
  MUX41X1_HVT U579 ( .A1(n8257), .A3(n8255), .A2(n8256), .A4(n8254), .S0(n11), 
        .S1(n14), .Y(q[131]) );
  IBUFFX16_HVT U592 ( .A(n5831), .Y(n11) );
  IBUFFX16_HVT U597 ( .A(n6643), .Y(n14) );
  MUX41X1_HVT U653 ( .A1(\ram[11][72] ), .A3(\ram[9][72] ), .A2(\ram[10][72] ), 
        .A4(\ram[8][72] ), .S0(n5125), .S1(n15), .Y(n8019) );
  IBUFFX16_HVT U654 ( .A(n5964), .Y(n15) );
  IBUFFX2_HVT U777 ( .A(n8781), .Y(n8821) );
  INVX0_HVT U781 ( .A(n6823), .Y(n4389) );
  INVX0_HVT U782 ( .A(n6815), .Y(n6823) );
  INVX1_HVT U784 ( .A(n7577), .Y(n5628) );
  MUX41X1_HVT U785 ( .A1(\ram[15][216] ), .A3(\ram[13][216] ), .A2(
        \ram[14][216] ), .A4(\ram[12][216] ), .S0(n4161), .S1(n19), .Y(n8593)
         );
  IBUFFX16_HVT U786 ( .A(n5147), .Y(n19) );
  IBUFFX4_HVT U787 ( .A(n8826), .Y(n4161) );
  INVX1_HVT U788 ( .A(n5632), .Y(n5090) );
  INVX1_HVT U789 ( .A(n5646), .Y(n7303) );
  INVX0_HVT U792 ( .A(n9028), .Y(n4596) );
  MUX41X1_HVT U800 ( .A1(\ram[0][241] ), .A3(\ram[2][241] ), .A2(\ram[1][241] ), .A4(\ram[3][241] ), .S0(n5946), .S1(n23), .Y(n8694) );
  IBUFFX16_HVT U801 ( .A(n4987), .Y(n23) );
  INVX1_HVT U802 ( .A(n6392), .Y(n8794) );
  MUX41X1_HVT U810 ( .A1(\ram[12][171] ), .A3(\ram[14][171] ), .A2(
        \ram[13][171] ), .A4(\ram[15][171] ), .S0(n26), .S1(n7696), .Y(n8413)
         );
  IBUFFX16_HVT U821 ( .A(n6645), .Y(n26) );
  IBUFFX2_HVT U832 ( .A(n7565), .Y(n5836) );
  INVX1_HVT U841 ( .A(n7311), .Y(n5294) );
  IBUFFX2_HVT U868 ( .A(n6406), .Y(n5970) );
  IBUFFX2_HVT U871 ( .A(n8874), .Y(n5127) );
  INVX1_HVT U872 ( .A(n8834), .Y(n6392) );
  INVX0_HVT U881 ( .A(n8778), .Y(n7271) );
  INVX0_HVT U889 ( .A(n7271), .Y(n5635) );
  MUX41X1_HVT U898 ( .A1(\ram[3][154] ), .A3(\ram[1][154] ), .A2(\ram[2][154] ), .A4(\ram[0][154] ), .S0(n5985), .S1(n27), .Y(n8348) );
  IBUFFX16_HVT U902 ( .A(n8860), .Y(n27) );
  IBUFFX2_HVT U948 ( .A(n7565), .Y(n7576) );
  INVX0_HVT U959 ( .A(n7551), .Y(n6742) );
  INVX0_HVT U966 ( .A(n5984), .Y(n6410) );
  MUX41X1_HVT U978 ( .A1(n8508), .A3(n8507), .A2(n8506), .A4(n8505), .S0(n6388), .S1(n6259), .Y(q[194]) );
  MUX41X2_HVT U987 ( .A1(\ram[15][194] ), .A3(\ram[13][194] ), .A2(
        \ram[14][194] ), .A4(\ram[12][194] ), .S0(n5941), .S1(n5567), .Y(n8505) );
  INVX0_HVT U1007 ( .A(n5660), .Y(n6388) );
  MUX41X1_HVT U1033 ( .A1(\ram[14][177] ), .A3(\ram[12][177] ), .A2(
        \ram[15][177] ), .A4(\ram[13][177] ), .S0(n5738), .S1(n8877), .Y(n8437) );
  IBUFFX2_HVT U1040 ( .A(n5610), .Y(n5638) );
  IBUFFX2_HVT U1041 ( .A(n5610), .Y(n7572) );
  IBUFFX2_HVT U1042 ( .A(n5610), .Y(n7281) );
  IBUFFX2_HVT U1043 ( .A(n8787), .Y(n8804) );
  IBUFFX2_HVT U1044 ( .A(n8787), .Y(n8816) );
  MUX41X1_HVT U1049 ( .A1(\ram[2][235] ), .A3(\ram[0][235] ), .A2(
        \ram[3][235] ), .A4(\ram[1][235] ), .S0(n6405), .S1(n6010), .Y(n8670)
         );
  INVX0_HVT U1050 ( .A(n7292), .Y(n7141) );
  INVX1_HVT U1051 ( .A(n5898), .Y(n5087) );
  MUX41X1_HVT U1052 ( .A1(n8428), .A3(n8426), .A2(n8427), .A4(n8425), .S0(n29), 
        .S1(n31), .Y(q[174]) );
  IBUFFX16_HVT U1053 ( .A(n5151), .Y(n29) );
  IBUFFX16_HVT U1054 ( .A(n5637), .Y(n31) );
  INVX0_HVT U1056 ( .A(n7705), .Y(n7668) );
  MUX41X1_HVT U1064 ( .A1(\ram[13][229] ), .A3(\ram[15][229] ), .A2(
        \ram[12][229] ), .A4(\ram[14][229] ), .S0(n5733), .S1(n5556), .Y(n8645) );
  MUX41X1_HVT U1065 ( .A1(n36), .A3(n35), .A2(n39), .A4(n42), .S0(n6645), .S1(
        n5616), .Y(n32) );
  IBUFFX16_HVT U1066 ( .A(n32), .Y(n8555) );
  IBUFFX16_HVT U1069 ( .A(\ram[4][206] ), .Y(n35) );
  IBUFFX2_HVT U1070 ( .A(n3), .Y(n8830) );
  MUX41X1_HVT U1071 ( .A1(\ram[7][162] ), .A3(\ram[5][162] ), .A2(
        \ram[6][162] ), .A4(\ram[4][162] ), .S0(n4989), .S1(n5457), .Y(n8379)
         );
  MUX41X1_HVT U1073 ( .A1(\ram[2][251] ), .A3(\ram[0][251] ), .A2(
        \ram[3][251] ), .A4(\ram[1][251] ), .S0(n4993), .S1(n5138), .Y(n8734)
         );
  INVX0_HVT U1077 ( .A(n5987), .Y(n6113) );
  MUX41X1_HVT U1080 ( .A1(n8384), .A3(n8383), .A2(n8382), .A4(n8381), .S0(
        n5092), .S1(n45), .Y(q[163]) );
  IBUFFX16_HVT U1083 ( .A(n5131), .Y(n45) );
  INVX1_HVT U1086 ( .A(n7310), .Y(n7584) );
  IBUFFX2_HVT U1092 ( .A(n8813), .Y(n6133) );
  IBUFFX2_HVT U1094 ( .A(n8813), .Y(n5794) );
  MUX41X1_HVT U1096 ( .A1(\ram[5][209] ), .A3(\ram[7][209] ), .A2(
        \ram[4][209] ), .A4(\ram[6][209] ), .S0(n6021), .S1(n5118), .Y(n8567)
         );
  IBUFFX2_HVT U1097 ( .A(n3), .Y(n8829) );
  INVX0_HVT U1098 ( .A(n7672), .Y(n1023) );
  MUX41X1_HVT U1103 ( .A1(n8525), .A3(n8527), .A2(n8526), .A4(n8528), .S0(n46), 
        .S1(n48), .Y(q[199]) );
  IBUFFX16_HVT U1106 ( .A(n5289), .Y(n46) );
  IBUFFX16_HVT U1111 ( .A(n5800), .Y(n48) );
  MUX41X1_HVT U1133 ( .A1(n8442), .A3(n8444), .A2(n8441), .A4(n8443), .S0(n58), 
        .S1(n7666), .Y(q[178]) );
  IBUFFX16_HVT U1165 ( .A(n6658), .Y(n58) );
  MUX41X1_HVT U1175 ( .A1(\ram[6][134] ), .A3(\ram[4][134] ), .A2(
        \ram[7][134] ), .A4(\ram[5][134] ), .S0(n6389), .S1(n8903), .Y(n8268)
         );
  INVX0_HVT U1183 ( .A(n7344), .Y(n6389) );
  IBUFFX2_HVT U1185 ( .A(n8812), .Y(n5984) );
  IBUFFX2_HVT U1189 ( .A(n8812), .Y(n6414) );
  INVX1_HVT U1220 ( .A(n8812), .Y(n7571) );
  IBUFFX2_HVT U1239 ( .A(n7668), .Y(n6038) );
  NBUFFX2_HVT U1243 ( .A(n5008), .Y(n5807) );
  IBUFFX2_HVT U1253 ( .A(n7550), .Y(n5602) );
  MUX41X1_HVT U1257 ( .A1(n866), .A3(n833), .A2(n877), .A4(n917), .S0(n5014), 
        .S1(n7331), .Y(n829) );
  IBUFFX16_HVT U1259 ( .A(n829), .Y(n8320) );
  IBUFFX16_HVT U1300 ( .A(\ram[3][147] ), .Y(n833) );
  INVX0_HVT U1301 ( .A(n6645), .Y(n8791) );
  INVX1_HVT U1305 ( .A(n6131), .Y(n6966) );
  INVX1_HVT U1306 ( .A(n7546), .Y(n7550) );
  IBUFFX2_HVT U1307 ( .A(n6641), .Y(n4177) );
  INVX1_HVT U1309 ( .A(n6733), .Y(n6136) );
  MUX41X1_HVT U1311 ( .A1(\ram[0][142] ), .A3(\ram[2][142] ), .A2(
        \ram[1][142] ), .A4(\ram[3][142] ), .S0(n8805), .S1(n1023), .Y(n8301)
         );
  IBUFFX2_HVT U1313 ( .A(n7551), .Y(n5594) );
  MUX41X1_HVT U1315 ( .A1(n8703), .A3(n8705), .A2(n8704), .A4(n8706), .S0(
        n5352), .S1(n5020), .Y(q[244]) );
  IBUFFX4_HVT U1316 ( .A(n5800), .Y(n5020) );
  NBUFFX2_HVT U1317 ( .A(n5661), .Y(n7344) );
  IBUFFX2_HVT U1318 ( .A(n7319), .Y(n7321) );
  IBUFFX2_HVT U1319 ( .A(n7319), .Y(n7325) );
  INVX1_HVT U1320 ( .A(n5785), .Y(n7546) );
  NBUFFX2_HVT U1321 ( .A(n7344), .Y(n1078) );
  MUX41X1_HVT U1323 ( .A1(n8586), .A3(n8588), .A2(n8585), .A4(n8587), .S0(
        n1137), .S1(n5239), .Y(q[214]) );
  IBUFFX16_HVT U1331 ( .A(n5156), .Y(n1137) );
  IBUFFX2_HVT U1332 ( .A(n8786), .Y(n8807) );
  INVX1_HVT U1333 ( .A(n8834), .Y(n5651) );
  INVX1_HVT U1337 ( .A(n5651), .Y(n8840) );
  INVX0_HVT U1339 ( .A(n5091), .Y(n4162) );
  IBUFFX2_HVT U1341 ( .A(n7347), .Y(n8784) );
  MUX41X1_HVT U1350 ( .A1(\ram[1][166] ), .A3(\ram[3][166] ), .A2(
        \ram[0][166] ), .A4(\ram[2][166] ), .S0(n4162), .S1(n5607), .Y(n8396)
         );
  IBUFFX2_HVT U1351 ( .A(n6023), .Y(n5738) );
  INVX0_HVT U1352 ( .A(n6003), .Y(n5957) );
  NBUFFX2_HVT U1353 ( .A(n5659), .Y(n8859) );
  IBUFFX2_HVT U1354 ( .A(n7546), .Y(n6005) );
  INVX0_HVT U1365 ( .A(n5895), .Y(n7292) );
  IBUFFX2_HVT U1368 ( .A(n5895), .Y(n5091) );
  IBUFFX2_HVT U1371 ( .A(n8786), .Y(n6183) );
  IBUFFX2_HVT U1394 ( .A(n5346), .Y(n7691) );
  IBUFFX2_HVT U1400 ( .A(n8833), .Y(n5640) );
  IBUFFX2_HVT U1412 ( .A(n8833), .Y(n5743) );
  IBUFFX2_HVT U1423 ( .A(n7284), .Y(n6021) );
  INVX0_HVT U1425 ( .A(N26), .Y(n7144) );
  MUX41X1_HVT U1473 ( .A1(n8658), .A3(n8660), .A2(n8657), .A4(n8659), .S0(
        n5575), .S1(n5087), .Y(q[232]) );
  MUX41X1_HVT U1515 ( .A1(n1357), .A3(n1344), .A2(n1359), .A4(n1361), .S0(
        n7313), .S1(n7580), .Y(n1144) );
  IBUFFX16_HVT U1523 ( .A(n1144), .Y(n7884) );
  IBUFFX16_HVT U1524 ( .A(\ram[8][38] ), .Y(n1344) );
  IBUFFX2_HVT U1533 ( .A(n8781), .Y(n5993) );
  IBUFFX2_HVT U1537 ( .A(n7319), .Y(n5866) );
  INVX0_HVT U1540 ( .A(n4165), .Y(n1389) );
  INVX0_HVT U1559 ( .A(n8860), .Y(n4165) );
  INVX0_HVT U1560 ( .A(n6736), .Y(n5819) );
  NBUFFX4_HVT U1562 ( .A(n4930), .Y(n7696) );
  INVX1_HVT U1564 ( .A(n8874), .Y(n5230) );
  INVX0_HVT U1567 ( .A(n8790), .Y(n1391) );
  INVX0_HVT U1578 ( .A(n1391), .Y(n1461) );
  INVX1_HVT U1582 ( .A(n4703), .Y(n6034) );
  MUX41X1_HVT U1592 ( .A1(\ram[15][185] ), .A3(\ram[13][185] ), .A2(
        \ram[14][185] ), .A4(\ram[12][185] ), .S0(n7561), .S1(n6732), .Y(n8469) );
  INVX0_HVT U1593 ( .A(n5155), .Y(n7338) );
  MUX41X1_HVT U1594 ( .A1(n8683), .A3(n8685), .A2(n8684), .A4(n8686), .S0(
        n1463), .S1(n5995), .Y(q[239]) );
  IBUFFX16_HVT U1598 ( .A(n6383), .Y(n1463) );
  INVX0_HVT U1601 ( .A(n5885), .Y(n4183) );
  MUX41X1_HVT U1602 ( .A1(\ram[9][216] ), .A3(\ram[11][216] ), .A2(
        \ram[8][216] ), .A4(\ram[10][216] ), .S0(n5657), .S1(n1633), .Y(n8594)
         );
  INVX0_HVT U1609 ( .A(n5566), .Y(n5956) );
  INVX1_HVT U1610 ( .A(n8885), .Y(n5730) );
  IBUFFX2_HVT U1611 ( .A(n7316), .Y(n7330) );
  IBUFFX2_HVT U1612 ( .A(n7316), .Y(n6024) );
  MUX41X1_HVT U1613 ( .A1(n8522), .A3(n8524), .A2(n8521), .A4(n8523), .S0(
        n1597), .S1(n4177), .Y(q[198]) );
  IBUFFX16_HVT U1615 ( .A(n5654), .Y(n1597) );
  IBUFFX2_HVT U1616 ( .A(n6001), .Y(n7266) );
  INVX0_HVT U1630 ( .A(n7334), .Y(n5231) );
  IBUFFX2_HVT U1680 ( .A(n5235), .Y(n4888) );
  IBUFFX2_HVT U1754 ( .A(n5235), .Y(n5377) );
  INVX0_HVT U1757 ( .A(n6646), .Y(n6408) );
  INVX0_HVT U1763 ( .A(n6646), .Y(n7678) );
  INVX0_HVT U1766 ( .A(n5260), .Y(n4518) );
  IBUFFX2_HVT U1779 ( .A(n7708), .Y(n1633) );
  INVX0_HVT U1797 ( .A(n5972), .Y(n1651) );
  INVX0_HVT U1819 ( .A(n6408), .Y(n7708) );
  MUX41X1_HVT U1820 ( .A1(n8337), .A3(n8339), .A2(n8338), .A4(n8340), .S0(
        n1798), .S1(n7702), .Y(q[152]) );
  IBUFFX16_HVT U2078 ( .A(n6415), .Y(n1798) );
  MUX41X1_HVT U2092 ( .A1(n3949), .A3(n3929), .A2(n4105), .A4(n4157), .S0(
        n7303), .S1(n5138), .Y(n1801) );
  IBUFFX16_HVT U2096 ( .A(n1801), .Y(n8378) );
  IBUFFX16_HVT U2098 ( .A(\ram[8][162] ), .Y(n3929) );
  INVX1_HVT U2099 ( .A(n5565), .Y(n5566) );
  INVX1_HVT U2106 ( .A(n5583), .Y(n5000) );
  IBUFFX2_HVT U2107 ( .A(n5905), .Y(n6022) );
  MUX41X1_HVT U2113 ( .A1(\ram[7][163] ), .A3(\ram[5][163] ), .A2(
        \ram[6][163] ), .A4(\ram[4][163] ), .S0(n4158), .S1(n5084), .Y(n8383)
         );
  IBUFFX16_HVT U2120 ( .A(n7145), .Y(n4158) );
  INVX0_HVT U2128 ( .A(n5127), .Y(n5108) );
  INVX1_HVT U2139 ( .A(n4772), .Y(n5084) );
  MUX21X2_HVT U2337 ( .A1(n5320), .A2(n5319), .S0(n5562), .Y(n8703) );
  INVX0_HVT U2338 ( .A(n7283), .Y(n5134) );
  INVX1_HVT U2350 ( .A(n8882), .Y(n7283) );
  MUX41X1_HVT U2364 ( .A1(\ram[8][190] ), .A3(\ram[10][190] ), .A2(
        \ram[9][190] ), .A4(\ram[11][190] ), .S0(n4159), .S1(n8881), .Y(n8490)
         );
  IBUFFX16_HVT U2366 ( .A(n7682), .Y(n4159) );
  INVX0_HVT U2369 ( .A(n7564), .Y(n5488) );
  MUX41X1_HVT U2370 ( .A1(\ram[4][128] ), .A3(\ram[6][128] ), .A2(
        \ram[5][128] ), .A4(\ram[7][128] ), .S0(n4160), .S1(n5147), .Y(n8244)
         );
  IBUFFX16_HVT U2376 ( .A(n7147), .Y(n4160) );
  IBUFFX2_HVT U2377 ( .A(n5996), .Y(n6384) );
  MUX41X1_HVT U2379 ( .A1(\ram[2][245] ), .A3(\ram[0][245] ), .A2(
        \ram[3][245] ), .A4(\ram[1][245] ), .S0(n5738), .S1(n5147), .Y(n8710)
         );
  IBUFFX2_HVT U2385 ( .A(n8888), .Y(n5229) );
  INVX0_HVT U2386 ( .A(n7315), .Y(n5147) );
  MUX41X1_HVT U2387 ( .A1(\ram[7][183] ), .A3(\ram[5][183] ), .A2(
        \ram[6][183] ), .A4(\ram[4][183] ), .S0(n4161), .S1(n5141), .Y(n8463)
         );
  DELLN1X2_HVT U2388 ( .A(n5819), .Y(n8870) );
  IBUFFX2_HVT U2395 ( .A(n5565), .Y(n5141) );
  IBUFFX2_HVT U2402 ( .A(n5984), .Y(n8793) );
  IBUFFX2_HVT U2422 ( .A(n5984), .Y(n5132) );
  INVX0_HVT U2447 ( .A(n7549), .Y(n4178) );
  INVX1_HVT U2466 ( .A(n7283), .Y(n5562) );
  IBUFFX2_HVT U2497 ( .A(n5583), .Y(n7264) );
  IBUFFX2_HVT U2511 ( .A(n5583), .Y(n8818) );
  MUX41X1_HVT U2565 ( .A1(n8656), .A3(n8654), .A2(n8655), .A4(n8653), .S0(
        n5752), .S1(n5980), .Y(q[231]) );
  IBUFFX2_HVT U2566 ( .A(n5980), .Y(n5868) );
  MUX41X1_HVT U2597 ( .A1(\ram[1][156] ), .A3(\ram[3][156] ), .A2(
        \ram[0][156] ), .A4(\ram[2][156] ), .S0(n5310), .S1(n7315), .Y(n8356)
         );
  INVX1_HVT U2855 ( .A(n8900), .Y(n5715) );
  NOR2X4_HVT U2856 ( .A1(n6114), .A2(n1461), .Y(n9) );
  MUX41X1_HVT U2865 ( .A1(n7914), .A3(n7912), .A2(n7913), .A4(n7911), .S0(
        n4163), .S1(n4164), .Y(q[45]) );
  IBUFFX16_HVT U2887 ( .A(n5015), .Y(n4163) );
  IBUFFX16_HVT U2889 ( .A(n4999), .Y(n4164) );
  INVX1_HVT U2890 ( .A(n5715), .Y(n5656) );
  MUX41X1_HVT U2891 ( .A1(\ram[7][146] ), .A3(\ram[5][146] ), .A2(
        \ram[6][146] ), .A4(\ram[4][146] ), .S0(n5824), .S1(n4165), .Y(n8315)
         );
  INVX0_HVT U3114 ( .A(n5311), .Y(n8790) );
  IBUFFX2_HVT U3115 ( .A(n8780), .Y(n7291) );
  INVX0_HVT U3117 ( .A(n5342), .Y(n4166) );
  INVX0_HVT U3132 ( .A(n6395), .Y(n4167) );
  NBUFFX2_HVT U3146 ( .A(n7692), .Y(n5342) );
  NBUFFX2_HVT U3150 ( .A(n5797), .Y(n6395) );
  MUX41X1_HVT U3152 ( .A1(n4170), .A3(n4169), .A2(n4171), .A4(n4172), .S0(
        n6018), .S1(n5084), .Y(n4168) );
  IBUFFX16_HVT U3153 ( .A(n4168), .Y(n8275) );
  IBUFFX16_HVT U3167 ( .A(\ram[11][136] ), .Y(n4169) );
  MUX41X1_HVT U3187 ( .A1(\ram[6][151] ), .A3(\ram[4][151] ), .A2(
        \ram[7][151] ), .A4(\ram[5][151] ), .S0(n5884), .S1(n6747), .Y(n8335)
         );
  INVX0_HVT U3201 ( .A(n8945), .Y(n4678) );
  MUX41X1_HVT U3203 ( .A1(\ram[0][188] ), .A3(\ram[2][188] ), .A2(
        \ram[1][188] ), .A4(\ram[3][188] ), .S0(n4173), .S1(n6132), .Y(n8484)
         );
  IBUFFX16_HVT U3216 ( .A(n7314), .Y(n4173) );
  INVX0_HVT U3258 ( .A(n7671), .Y(n6251) );
  IBUFFX2_HVT U3260 ( .A(n6126), .Y(n6132) );
  INVX0_HVT U3261 ( .A(N26), .Y(n7295) );
  INVX0_HVT U3289 ( .A(n7692), .Y(n5641) );
  INVX0_HVT U3324 ( .A(n6113), .Y(n4174) );
  INVX0_HVT U3375 ( .A(n5298), .Y(n5016) );
  INVX0_HVT U3377 ( .A(n10379), .Y(n6123) );
  INVX0_HVT U3381 ( .A(n7547), .Y(n5012) );
  INVX1_HVT U3389 ( .A(n7664), .Y(n4175) );
  IBUFFX2_HVT U3405 ( .A(n8813), .Y(n5357) );
  NBUFFX2_HVT U3406 ( .A(n6737), .Y(n8855) );
  NBUFFX2_HVT U3408 ( .A(n6394), .Y(n4176) );
  INVX1_HVT U3437 ( .A(n5129), .Y(n6735) );
  IBUFFX2_HVT U3438 ( .A(n5906), .Y(n6126) );
  IBUFFX2_HVT U3439 ( .A(n5087), .Y(n5369) );
  IBUFFX2_HVT U3446 ( .A(n7664), .Y(n7688) );
  INVX1_HVT U3449 ( .A(n5617), .Y(n5608) );
  MUX41X1_HVT U3450 ( .A1(\ram[14][137] ), .A3(\ram[12][137] ), .A2(
        \ram[15][137] ), .A4(\ram[13][137] ), .S0(n4178), .S1(n4189), .Y(n8278) );
  INVX0_HVT U3453 ( .A(n5729), .Y(n5724) );
  NBUFFX4_HVT U3455 ( .A(n4848), .Y(n7681) );
  INVX0_HVT U3461 ( .A(n7333), .Y(n5007) );
  IBUFFX2_HVT U3479 ( .A(n7710), .Y(n6655) );
  IBUFFX2_HVT U3499 ( .A(n7710), .Y(n5818) );
  MUX41X1_HVT U3514 ( .A1(n8650), .A3(n8652), .A2(n8649), .A4(n8651), .S0(
        n4179), .S1(n4180), .Y(q[230]) );
  IBUFFX16_HVT U3520 ( .A(n4998), .Y(n4179) );
  IBUFFX16_HVT U3522 ( .A(n5039), .Y(n4180) );
  INVX1_HVT U3539 ( .A(n8883), .Y(n6551) );
  INVX0_HVT U3567 ( .A(n6551), .Y(n5621) );
  DELLN2X2_HVT U3596 ( .A(n8882), .Y(n8909) );
  IBUFFX2_HVT U3630 ( .A(n5729), .Y(n6734) );
  INVX0_HVT U3635 ( .A(n8790), .Y(n8782) );
  NBUFFX4_HVT U3647 ( .A(n7710), .Y(n6382) );
  INVX1_HVT U3686 ( .A(n5094), .Y(n8783) );
  MUX41X1_HVT U3693 ( .A1(\ram[14][128] ), .A3(\ram[12][128] ), .A2(
        \ram[15][128] ), .A4(\ram[13][128] ), .S0(n4193), .S1(n4181), .Y(n8242) );
  IBUFFX16_HVT U3705 ( .A(n6393), .Y(n4181) );
  IBUFFX2_HVT U3740 ( .A(n8786), .Y(n8809) );
  INVX1_HVT U3782 ( .A(n7664), .Y(n4847) );
  NBUFFX4_HVT U3895 ( .A(n7318), .Y(n8863) );
  INVX0_HVT U3910 ( .A(n8883), .Y(n5825) );
  INVX0_HVT U3924 ( .A(n8883), .Y(n7331) );
  NBUFFX2_HVT U3925 ( .A(n6395), .Y(n4182) );
  MUX41X1_HVT U3926 ( .A1(n8354), .A3(n8356), .A2(n8353), .A4(n8355), .S0(
        n5623), .S1(n4183), .Y(q[156]) );
  INVX1_HVT U3928 ( .A(n8783), .Y(n7551) );
  INVX1_HVT U3946 ( .A(n5653), .Y(n5572) );
  INVX1_HVT U3973 ( .A(n5486), .Y(n5479) );
  INVX0_HVT U3981 ( .A(n5796), .Y(n5797) );
  IBUFFX2_HVT U4001 ( .A(n6663), .Y(n6640) );
  INVX0_HVT U4046 ( .A(n5103), .Y(n5071) );
  INVX0_HVT U4050 ( .A(n4193), .Y(n4184) );
  INVX0_HVT U4102 ( .A(n7325), .Y(n4193) );
  MUX41X1_HVT U4103 ( .A1(n8460), .A3(n8458), .A2(n8459), .A4(n8457), .S0(
        n4185), .S1(n5239), .Y(q[182]) );
  IBUFFX4_HVT U4114 ( .A(n5623), .Y(n4185) );
  MUX41X1_HVT U4138 ( .A1(n8674), .A3(n8672), .A2(n8673), .A4(n8671), .S0(
        n4185), .S1(n4186), .Y(q[236]) );
  IBUFFX16_HVT U4145 ( .A(n5338), .Y(n4186) );
  MUX41X1_HVT U4155 ( .A1(n8489), .A3(n8491), .A2(n8490), .A4(n8492), .S0(
        n4187), .S1(n4190), .Y(q[190]) );
  IBUFFX16_HVT U4156 ( .A(n5925), .Y(n4187) );
  IBUFFX2_HVT U4157 ( .A(n1461), .Y(n5961) );
  INVX1_HVT U4158 ( .A(n7292), .Y(n5751) );
  INVX1_HVT U4159 ( .A(n4192), .Y(n7582) );
  INVX1_HVT U4160 ( .A(n5377), .Y(n7671) );
  IBUFFX2_HVT U4161 ( .A(n6126), .Y(n4188) );
  INVX1_HVT U4162 ( .A(n5106), .Y(n6754) );
  INVX0_HVT U4163 ( .A(n7280), .Y(n4190) );
  INVX0_HVT U4164 ( .A(n7299), .Y(n7280) );
  DELLN2X2_HVT U4165 ( .A(n8882), .Y(n7704) );
  IBUFFX2_HVT U4166 ( .A(n5426), .Y(n5967) );
  IBUFFX2_HVT U4167 ( .A(n8782), .Y(n5859) );
  IBUFFX2_HVT U4168 ( .A(n5091), .Y(n6652) );
  IBUFFX2_HVT U4169 ( .A(n7347), .Y(n5518) );
  IBUFFX2_HVT U4170 ( .A(n4703), .Y(n4189) );
  IBUFFX2_HVT U4171 ( .A(n5583), .Y(n8824) );
  IBUFFX2_HVT U4172 ( .A(n5583), .Y(n6007) );
  IBUFFX2_HVT U4173 ( .A(n7263), .Y(n7313) );
  INVX1_HVT U4174 ( .A(n6138), .Y(n5875) );
  INVX0_HVT U4175 ( .A(n7705), .Y(n4191) );
  INVX0_HVT U4176 ( .A(n4191), .Y(n4192) );
  IBUFFX2_HVT U4177 ( .A(n5651), .Y(n7324) );
  MUX41X1_HVT U4178 ( .A1(\ram[15][250] ), .A3(\ram[13][250] ), .A2(
        \ram[14][250] ), .A4(\ram[12][250] ), .S0(n4193), .S1(n7688), .Y(n8727) );
  NBUFFX4_HVT U4179 ( .A(n6737), .Y(n7676) );
  INVX1_HVT U4180 ( .A(n8871), .Y(n6138) );
  INVX1_HVT U4181 ( .A(n7676), .Y(n5077) );
  INVX0_HVT U4182 ( .A(n6052), .Y(n6054) );
  INVX0_HVT U4183 ( .A(n7250), .Y(n4194) );
  INVX0_HVT U4184 ( .A(n4194), .Y(n4195) );
  INVX0_HVT U4185 ( .A(n9015), .Y(n9021) );
  OAI22X1_HVT U4186 ( .A1(n4196), .A2(n5378), .A3(n5603), .A4(n4594), .Y(n3927) );
  INVX0_HVT U4187 ( .A(n9014), .Y(n9017) );
  IBUFFX4_HVT U4188 ( .A(n9386), .Y(n4594) );
  INVX0_HVT U4189 ( .A(n4496), .Y(n4197) );
  NBUFFX2_HVT U4190 ( .A(n10370), .Y(n4198) );
  INVX0_HVT U4191 ( .A(n10370), .Y(n6712) );
  INVX0_HVT U4192 ( .A(n6876), .Y(n6885) );
  INVX0_HVT U4193 ( .A(n6876), .Y(n6847) );
  INVX0_HVT U4194 ( .A(n6876), .Y(n6878) );
  NBUFFX2_HVT U4195 ( .A(n6425), .Y(n4199) );
  INVX0_HVT U4196 ( .A(n4262), .Y(n4200) );
  INVX0_HVT U4197 ( .A(n5680), .Y(n5689) );
  OAI22X1_HVT U4198 ( .A1(n4201), .A2(n4202), .A3(n4645), .A4(n9579), .Y(n1432) );
  INVX0_HVT U4199 ( .A(n4773), .Y(n4202) );
  INVX0_HVT U4200 ( .A(n4202), .Y(n4203) );
  OAI22X1_HVT U4201 ( .A1(n4204), .A2(n4205), .A3(n5951), .A4(n4768), .Y(n1409) );
  IBUFFX4_HVT U4202 ( .A(data[68]), .Y(n4768) );
  INVX0_HVT U4203 ( .A(n4331), .Y(n4205) );
  INVX0_HVT U4204 ( .A(n4205), .Y(n4206) );
  INVX0_HVT U4205 ( .A(n7446), .Y(n7438) );
  INVX0_HVT U4206 ( .A(n7446), .Y(n7448) );
  INVX0_HVT U4207 ( .A(n7449), .Y(n7447) );
  INVX0_HVT U4208 ( .A(n7449), .Y(n7467) );
  INVX0_HVT U4209 ( .A(n7421), .Y(n7423) );
  INVX0_HVT U4210 ( .A(n7421), .Y(n7422) );
  INVX0_HVT U4211 ( .A(n5669), .Y(n4207) );
  INVX0_HVT U4212 ( .A(n4207), .Y(n4208) );
  INVX0_HVT U4213 ( .A(n5670), .Y(n4209) );
  INVX0_HVT U4214 ( .A(n4209), .Y(n4210) );
  INVX0_HVT U4215 ( .A(n6716), .Y(n4441) );
  INVX0_HVT U4216 ( .A(n6718), .Y(n6716) );
  INVX0_HVT U4217 ( .A(n6800), .Y(n4211) );
  OAI22X1_HVT U4218 ( .A1(n4213), .A2(n4605), .A3(n6109), .A4(n4212), .Y(n2120) );
  IBUFFX16_HVT U4219 ( .A(n9341), .Y(n4212) );
  INVX0_HVT U4220 ( .A(n7389), .Y(n7375) );
  INVX0_HVT U4221 ( .A(n6064), .Y(n6066) );
  INVX0_HVT U4222 ( .A(n4222), .Y(n4214) );
  INVX0_HVT U4223 ( .A(n7405), .Y(n4222) );
  INVX0_HVT U4224 ( .A(n7449), .Y(n7450) );
  INVX0_HVT U4225 ( .A(n7421), .Y(n7452) );
  INVX0_HVT U4226 ( .A(n7446), .Y(n7439) );
  INVX0_HVT U4227 ( .A(n30), .Y(n4215) );
  INVX0_HVT U4228 ( .A(n4215), .Y(n4216) );
  INVX0_HVT U4229 ( .A(n6530), .Y(n6546) );
  INVX0_HVT U4230 ( .A(n6530), .Y(n6549) );
  INVX0_HVT U4231 ( .A(n6530), .Y(n6532) );
  INVX0_HVT U4232 ( .A(n6534), .Y(n6541) );
  INVX0_HVT U4233 ( .A(n6534), .Y(n6540) );
  INVX0_HVT U4234 ( .A(n6534), .Y(n6536) );
  INVX0_HVT U4235 ( .A(n6527), .Y(n6535) );
  INVX0_HVT U4236 ( .A(n6527), .Y(n6529) );
  INVX0_HVT U4237 ( .A(n6527), .Y(n6528) );
  OAI22X1_HVT U4238 ( .A1(n4219), .A2(n4260), .A3(n4217), .A4(n4218), .Y(n439)
         );
  IBUFFX16_HVT U4239 ( .A(n6842), .Y(n4217) );
  IBUFFX16_HVT U4240 ( .A(n9673), .Y(n4218) );
  INVX0_HVT U4241 ( .A(n5271), .Y(n5281) );
  INVX0_HVT U4242 ( .A(n7121), .Y(n7127) );
  INVX0_HVT U4243 ( .A(n6060), .Y(n6061) );
  INVX0_HVT U4244 ( .A(n6060), .Y(n6101) );
  INVX0_HVT U4245 ( .A(n6060), .Y(n6085) );
  OAI22X1_HVT U4246 ( .A1(n4221), .A2(n4281), .A3(n4280), .A4(n4220), .Y(n2156) );
  IBUFFX16_HVT U4247 ( .A(n9449), .Y(n4220) );
  INVX0_HVT U4248 ( .A(n6097), .Y(n6099) );
  OAI22X1_HVT U4249 ( .A1(n4224), .A2(n4222), .A3(n4280), .A4(n4223), .Y(n2148) );
  IBUFFX16_HVT U4250 ( .A(n9425), .Y(n4223) );
  INVX0_HVT U4251 ( .A(n6098), .Y(n6100) );
  OAI22X1_HVT U4252 ( .A1(n4226), .A2(n4225), .A3(n4232), .A4(n9995), .Y(n2590) );
  IBUFFX16_HVT U4253 ( .A(n7640), .Y(n4225) );
  INVX0_HVT U4254 ( .A(n4874), .Y(n4227) );
  INVX0_HVT U4255 ( .A(n9228), .Y(n4874) );
  NBUFFX2_HVT U4256 ( .A(n4481), .Y(n4228) );
  INVX0_HVT U4257 ( .A(n6060), .Y(n6068) );
  INVX0_HVT U4258 ( .A(n5674), .Y(n4229) );
  INVX0_HVT U4259 ( .A(n4229), .Y(n4230) );
  INVX0_HVT U4260 ( .A(n4566), .Y(n4231) );
  INVX0_HVT U4261 ( .A(n4937), .Y(n4566) );
  INVX0_HVT U4262 ( .A(n9126), .Y(n4232) );
  INVX0_HVT U4263 ( .A(n4232), .Y(n4233) );
  OAI22X1_HVT U4264 ( .A1(n4235), .A2(n4234), .A3(n4502), .A4(n9998), .Y(n2591) );
  IBUFFX16_HVT U4265 ( .A(n7639), .Y(n4234) );
  OAI22X1_HVT U4266 ( .A1(n4237), .A2(n4258), .A3(n4236), .A4(n4576), .Y(n569)
         );
  IBUFFX16_HVT U4267 ( .A(n6886), .Y(n4236) );
  IBUFFX4_HVT U4268 ( .A(n10081), .Y(n4576) );
  NBUFFX2_HVT U4269 ( .A(n7415), .Y(n4238) );
  INVX0_HVT U4270 ( .A(n10362), .Y(n4239) );
  OAI22X1_HVT U4271 ( .A1(n4241), .A2(n4849), .A3(n4729), .A4(n4240), .Y(n1438) );
  IBUFFX16_HVT U4272 ( .A(n9598), .Y(n4240) );
  OAI22X1_HVT U4273 ( .A1(n4244), .A2(n4306), .A3(n4242), .A4(n4243), .Y(n847)
         );
  IBUFFX16_HVT U4274 ( .A(n6768), .Y(n4242) );
  IBUFFX16_HVT U4275 ( .A(n9362), .Y(n4243) );
  OAI22X1_HVT U4276 ( .A1(n4247), .A2(n5374), .A3(n4245), .A4(n4246), .Y(n846)
         );
  IBUFFX16_HVT U4277 ( .A(n5249), .Y(n4245) );
  IBUFFX16_HVT U4278 ( .A(n9359), .Y(n4246) );
  OA22X1_HVT U4279 ( .A1(n4250), .A2(n4306), .A3(n4249), .A4(n4711), .Y(n4248)
         );
  IBUFFX16_HVT U4280 ( .A(n4248), .Y(n837) );
  IBUFFX16_HVT U4281 ( .A(n4544), .Y(n4249) );
  IBUFFX4_HVT U4282 ( .A(n9331), .Y(n4711) );
  OAI22X1_HVT U4283 ( .A1(n4252), .A2(n5374), .A3(n5253), .A4(n4251), .Y(n832)
         );
  IBUFFX16_HVT U4284 ( .A(n9315), .Y(n4251) );
  INVX0_HVT U4285 ( .A(n5257), .Y(n5258) );
  OAI22X1_HVT U4286 ( .A1(n4253), .A2(n5374), .A3(n5265), .A4(n9837), .Y(n1004) );
  INVX1_HVT U4287 ( .A(data[175]), .Y(n9837) );
  INVX0_HVT U4288 ( .A(n5242), .Y(n4254) );
  INVX0_HVT U4289 ( .A(n5674), .Y(n4255) );
  INVX0_HVT U4290 ( .A(n4255), .Y(n4256) );
  INVX0_HVT U4291 ( .A(n9061), .Y(n4257) );
  INVX0_HVT U4292 ( .A(n7079), .Y(n4258) );
  INVX0_HVT U4293 ( .A(n4258), .Y(n4259) );
  INVX0_HVT U4294 ( .A(n7082), .Y(n4260) );
  INVX0_HVT U4295 ( .A(n4260), .Y(n4261) );
  INVX0_HVT U4296 ( .A(n10305), .Y(n6159) );
  INVX0_HVT U4297 ( .A(n7027), .Y(n7074) );
  INVX0_HVT U4298 ( .A(n10349), .Y(n4262) );
  INVX0_HVT U4299 ( .A(n4262), .Y(n4263) );
  INVX0_HVT U4300 ( .A(n7413), .Y(n4281) );
  INVX1_HVT U4301 ( .A(n10108), .Y(n5748) );
  INVX0_HVT U4302 ( .A(n5920), .Y(n5383) );
  INVX0_HVT U4303 ( .A(n4265), .Y(n4264) );
  INVX0_HVT U4304 ( .A(n7038), .Y(n4265) );
  INVX0_HVT U4305 ( .A(n4265), .Y(n4266) );
  OAI22X1_HVT U4306 ( .A1(n4267), .A2(n4670), .A3(n7269), .A4(n9821), .Y(n1511) );
  INVX0_HVT U4307 ( .A(n4402), .Y(n4268) );
  INVX0_HVT U4308 ( .A(n6605), .Y(n4402) );
  INVX0_HVT U4309 ( .A(n6103), .Y(n6104) );
  INVX1_HVT U4310 ( .A(n10227), .Y(n6103) );
  NBUFFX2_HVT U4311 ( .A(n4683), .Y(n4269) );
  INVX0_HVT U4312 ( .A(n9072), .Y(n4270) );
  NBUFFX2_HVT U4313 ( .A(n9257), .Y(n4271) );
  NOR2X1_HVT U4314 ( .A1(n7292), .A2(n5543), .Y(n21) );
  INVX0_HVT U4315 ( .A(n9015), .Y(n9023) );
  INVX0_HVT U4316 ( .A(n6512), .Y(n4272) );
  INVX0_HVT U4317 ( .A(n6511), .Y(n4273) );
  INVX0_HVT U4318 ( .A(n9081), .Y(n9119) );
  INVX0_HVT U4319 ( .A(n10133), .Y(n6356) );
  INVX0_HVT U4320 ( .A(n4354), .Y(n4274) );
  INVX0_HVT U4321 ( .A(n4400), .Y(n4275) );
  INVX0_HVT U4322 ( .A(n6592), .Y(n4400) );
  OAI22X1_HVT U4323 ( .A1(n4276), .A2(n4283), .A3(n4368), .A4(n9561), .Y(n3218) );
  OAI22X1_HVT U4324 ( .A1(n4277), .A2(n4283), .A3(n4368), .A4(n9349), .Y(n3147) );
  INVX0_HVT U4325 ( .A(n6567), .Y(n4283) );
  INVX0_HVT U4326 ( .A(n6559), .Y(n4546) );
  INVX0_HVT U4327 ( .A(n9071), .Y(n4278) );
  INVX0_HVT U4328 ( .A(n5190), .Y(n4279) );
  INVX0_HVT U4329 ( .A(n5189), .Y(n5190) );
  INVX0_HVT U4330 ( .A(n10229), .Y(n4280) );
  INVX0_HVT U4331 ( .A(n4631), .Y(n1216) );
  OAI22X1_HVT U4332 ( .A1(n4282), .A2(n4281), .A3(n4436), .A4(n4390), .Y(n2141) );
  INVX0_HVT U4333 ( .A(n6109), .Y(n6111) );
  IBUFFX4_HVT U4334 ( .A(data[32]), .Y(n4390) );
  INVX0_HVT U4335 ( .A(n6312), .Y(n6314) );
  INVX0_HVT U4336 ( .A(n7197), .Y(n7200) );
  OAI22X1_HVT U4337 ( .A1(n4284), .A2(n4283), .A3(n4304), .A4(n9727), .Y(n3273) );
  OA22X1_HVT U4338 ( .A1(n4287), .A2(n4320), .A3(n4688), .A4(n4286), .Y(n4285)
         );
  IBUFFX16_HVT U4339 ( .A(n4285), .Y(n1353) );
  IBUFFX16_HVT U4340 ( .A(n9344), .Y(n4286) );
  OAI22X1_HVT U4341 ( .A1(n4288), .A2(n4494), .A3(n4478), .A4(n4449), .Y(n3693) );
  IBUFFX4_HVT U4342 ( .A(data[48]), .Y(n4449) );
  INVX0_HVT U4343 ( .A(n8948), .Y(n5454) );
  OAI22X1_HVT U4344 ( .A1(n4290), .A2(n4498), .A3(n4301), .A4(n4289), .Y(n3700) );
  IBUFFX16_HVT U4345 ( .A(n9473), .Y(n4289) );
  OA22X1_HVT U4346 ( .A1(n4292), .A2(n4964), .A3(n6229), .A4(n9730), .Y(n4291)
         );
  IBUFFX16_HVT U4347 ( .A(n4291), .Y(n1226) );
  INVX0_HVT U4348 ( .A(n6069), .Y(n6070) );
  INVX1_HVT U4349 ( .A(n10235), .Y(n6069) );
  INVX0_HVT U4350 ( .A(n5278), .Y(n4293) );
  INVX0_HVT U4351 ( .A(n5278), .Y(n4294) );
  INVX0_HVT U4352 ( .A(n5248), .Y(n4295) );
  INVX0_HVT U4353 ( .A(n5248), .Y(n4296) );
  INVX0_HVT U4354 ( .A(n10119), .Y(n4297) );
  INVX0_HVT U4355 ( .A(n4297), .Y(n4298) );
  NBUFFX2_HVT U4356 ( .A(n4513), .Y(n4299) );
  INVX0_HVT U4357 ( .A(n9062), .Y(n4300) );
  INVX0_HVT U4358 ( .A(n9046), .Y(n4301) );
  INVX0_HVT U4359 ( .A(n4301), .Y(n4302) );
  INVX0_HVT U4360 ( .A(n4582), .Y(n4303) );
  INVX0_HVT U4361 ( .A(n6800), .Y(n6801) );
  INVX0_HVT U4362 ( .A(n6800), .Y(n6802) );
  INVX0_HVT U4363 ( .A(n6331), .Y(n4304) );
  INVX0_HVT U4364 ( .A(n4304), .Y(n4305) );
  INVX0_HVT U4365 ( .A(n7100), .Y(n4306) );
  INVX0_HVT U4366 ( .A(n4306), .Y(n4307) );
  NBUFFX2_HVT U4367 ( .A(n4334), .Y(n4308) );
  NBUFFX2_HVT U4368 ( .A(n6361), .Y(n4309) );
  NBUFFX2_HVT U4369 ( .A(n6363), .Y(n4310) );
  INVX0_HVT U4370 ( .A(n4365), .Y(n4311) );
  INVX0_HVT U4371 ( .A(n7388), .Y(n4365) );
  INVX0_HVT U4372 ( .A(n6077), .Y(n6079) );
  INVX0_HVT U4373 ( .A(n4861), .Y(n4312) );
  INVX0_HVT U4374 ( .A(n4312), .Y(n4313) );
  INVX0_HVT U4375 ( .A(n7428), .Y(n4314) );
  NBUFFX2_HVT U4376 ( .A(n7185), .Y(n4315) );
  NBUFFX2_HVT U4377 ( .A(n7185), .Y(n4316) );
  NBUFFX2_HVT U4378 ( .A(n7185), .Y(n4317) );
  INVX0_HVT U4379 ( .A(n6511), .Y(n6544) );
  INVX0_HVT U4380 ( .A(n6511), .Y(n6503) );
  INVX0_HVT U4381 ( .A(n6511), .Y(n6513) );
  INVX0_HVT U4382 ( .A(n6512), .Y(n6547) );
  INVX0_HVT U4383 ( .A(n6512), .Y(n6493) );
  INVX0_HVT U4384 ( .A(n6512), .Y(n6514) );
  OAI22X1_HVT U4385 ( .A1(n4319), .A2(n4964), .A3(n4318), .A4(n9901), .Y(n1280) );
  IBUFFX16_HVT U4386 ( .A(n6212), .Y(n4318) );
  INVX1_HVT U4387 ( .A(data[195]), .Y(n9901) );
  INVX0_HVT U4388 ( .A(n4607), .Y(n3304) );
  INVX0_HVT U4389 ( .A(n5691), .Y(n4320) );
  INVX0_HVT U4390 ( .A(n4320), .Y(n4321) );
  INVX0_HVT U4391 ( .A(n4447), .Y(n4322) );
  INVX0_HVT U4392 ( .A(n6870), .Y(n4323) );
  INVX0_HVT U4393 ( .A(n4649), .Y(n4324) );
  INVX0_HVT U4394 ( .A(n4324), .Y(n4325) );
  INVX0_HVT U4395 ( .A(n10347), .Y(n4326) );
  INVX0_HVT U4396 ( .A(n4326), .Y(n4327) );
  OA22X1_HVT U4397 ( .A1(n4329), .A2(n5679), .A3(n5010), .A4(n10032), .Y(n4328) );
  IBUFFX16_HVT U4398 ( .A(n4328), .Y(n1578) );
  NBUFFX2_HVT U4399 ( .A(n4507), .Y(n4330) );
  INVX0_HVT U4400 ( .A(n5700), .Y(n4331) );
  INVX0_HVT U4401 ( .A(n7359), .Y(n7361) );
  INVX0_HVT U4402 ( .A(n4200), .Y(n4332) );
  INVX0_HVT U4403 ( .A(n7453), .Y(n7468) );
  INVX0_HVT U4404 ( .A(n7453), .Y(n7451) );
  INVX0_HVT U4405 ( .A(n7453), .Y(n7455) );
  INVX0_HVT U4406 ( .A(n7453), .Y(n7454) );
  INVX0_HVT U4407 ( .A(n6833), .Y(n6831) );
  INVX0_HVT U4408 ( .A(n6833), .Y(n6835) );
  INVX0_HVT U4409 ( .A(n6834), .Y(n6881) );
  INVX0_HVT U4410 ( .A(n6834), .Y(n6858) );
  INVX0_HVT U4411 ( .A(n6870), .Y(n6867) );
  INVX0_HVT U4412 ( .A(n6882), .Y(n6841) );
  INVX0_HVT U4413 ( .A(n9093), .Y(n4333) );
  INVX0_HVT U4414 ( .A(n4333), .Y(n4334) );
  INVX0_HVT U4415 ( .A(n4683), .Y(n4335) );
  OAI22X1_HVT U4416 ( .A1(n4336), .A2(n4337), .A3(n5253), .A4(n9989), .Y(n1052) );
  INVX0_HVT U4417 ( .A(n7095), .Y(n4337) );
  INVX0_HVT U4418 ( .A(n4337), .Y(n4338) );
  INVX0_HVT U4419 ( .A(n5349), .Y(n4339) );
  OAI22X1_HVT U4420 ( .A1(n4341), .A2(n6674), .A3(n4340), .A4(n6508), .Y(n164)
         );
  IBUFFX16_HVT U4421 ( .A(n9617), .Y(n4340) );
  INVX0_HVT U4422 ( .A(n6680), .Y(n6681) );
  INVX0_HVT U4423 ( .A(n6508), .Y(n6509) );
  INVX0_HVT U4424 ( .A(n6712), .Y(n4342) );
  INVX0_HVT U4425 ( .A(n7428), .Y(n7465) );
  INVX0_HVT U4426 ( .A(n5278), .Y(n5277) );
  INVX0_HVT U4427 ( .A(n5278), .Y(n5279) );
  INVX0_HVT U4428 ( .A(n5248), .Y(n5270) );
  INVX0_HVT U4429 ( .A(n5248), .Y(n5249) );
  INVX0_HVT U4430 ( .A(n6834), .Y(n6836) );
  INVX0_HVT U4431 ( .A(n6833), .Y(n6868) );
  INVX0_HVT U4432 ( .A(n6870), .Y(n6871) );
  INVX0_HVT U4433 ( .A(n4560), .Y(n4343) );
  INVX0_HVT U4434 ( .A(n6722), .Y(n4560) );
  INVX0_HVT U4435 ( .A(n6683), .Y(n4344) );
  INVX0_HVT U4436 ( .A(n7591), .Y(n4451) );
  INVX0_HVT U4437 ( .A(n7589), .Y(n7591) );
  INVX1_HVT U4438 ( .A(n4667), .Y(n7091) );
  INVX0_HVT U4439 ( .A(n4281), .Y(n4345) );
  INVX0_HVT U4440 ( .A(n6564), .Y(n4346) );
  OAI22X1_HVT U4441 ( .A1(n4348), .A2(n4614), .A3(n4347), .A4(n10054), .Y(n561) );
  IBUFFX16_HVT U4442 ( .A(n6845), .Y(n4347) );
  INVX0_HVT U4443 ( .A(n7359), .Y(n4349) );
  INVX0_HVT U4444 ( .A(n9242), .Y(n4350) );
  OAI22X1_HVT U4445 ( .A1(n4351), .A2(n4489), .A3(n4502), .A4(n4608), .Y(n2536) );
  INVX0_HVT U4446 ( .A(n7628), .Y(n7640) );
  INVX0_HVT U4447 ( .A(n9824), .Y(n9827) );
  IBUFFX4_HVT U4448 ( .A(n9827), .Y(n4608) );
  INVX0_HVT U4449 ( .A(n4478), .Y(n4352) );
  INVX0_HVT U4450 ( .A(n4532), .Y(n4478) );
  INVX0_HVT U4451 ( .A(n7376), .Y(n4353) );
  INVX0_HVT U4452 ( .A(n4368), .Y(n4354) );
  INVX0_HVT U4453 ( .A(n4305), .Y(n4368) );
  AOI21X1_HVT U4454 ( .A1(n20), .A2(n10377), .A3(n10381), .Y(n4355) );
  NBUFFX2_HVT U4455 ( .A(n6083), .Y(n4356) );
  INVX0_HVT U4456 ( .A(n6604), .Y(n4357) );
  INVX0_HVT U4457 ( .A(n9061), .Y(n9066) );
  INVX0_HVT U4458 ( .A(n9061), .Y(n9064) );
  INVX0_HVT U4459 ( .A(n9061), .Y(n9063) );
  INVX0_HVT U4460 ( .A(n4379), .Y(n4358) );
  OAI22X1_HVT U4461 ( .A1(n4359), .A2(n6255), .A3(n5265), .A4(n9803), .Y(n993)
         );
  INVX0_HVT U4462 ( .A(n7120), .Y(n7125) );
  INVX0_HVT U4463 ( .A(n5265), .Y(n5267) );
  INVX0_HVT U4464 ( .A(n6594), .Y(n4360) );
  INVX0_HVT U4465 ( .A(n4362), .Y(n4361) );
  INVX0_HVT U4466 ( .A(n7387), .Y(n4362) );
  OAI22X1_HVT U4467 ( .A1(n4364), .A2(n4362), .A3(n4436), .A4(n4363), .Y(n2127) );
  IBUFFX16_HVT U4468 ( .A(n9363), .Y(n4363) );
  INVX0_HVT U4469 ( .A(n6076), .Y(n6050) );
  IBUFFX4_HVT U4470 ( .A(n10226), .Y(n4436) );
  OAI22X1_HVT U4471 ( .A1(n4366), .A2(n4365), .A3(n6110), .A4(n9358), .Y(n2126) );
  INVX0_HVT U4472 ( .A(n6110), .Y(n6112) );
  OAI22X1_HVT U4473 ( .A1(n4367), .A2(n5349), .A3(n5282), .A4(n9621), .Y(n934)
         );
  INVX0_HVT U4474 ( .A(n7130), .Y(n7134) );
  INVX0_HVT U4475 ( .A(n5282), .Y(n5283) );
  INVX0_HVT U4476 ( .A(n10314), .Y(n5282) );
  OAI22X1_HVT U4477 ( .A1(n4369), .A2(n6593), .A3(n4368), .A4(n9600), .Y(n3231) );
  INVX0_HVT U4478 ( .A(n6586), .Y(n6588) );
  INVX0_HVT U4479 ( .A(n6159), .Y(n4370) );
  INVX0_HVT U4480 ( .A(n4908), .Y(n4371) );
  INVX0_HVT U4481 ( .A(n4908), .Y(n4909) );
  INVX0_HVT U4482 ( .A(n6671), .Y(n6692) );
  INVX0_HVT U4483 ( .A(n4239), .Y(n6678) );
  INVX0_HVT U4484 ( .A(n6193), .Y(n4966) );
  INVX0_HVT U4485 ( .A(n6232), .Y(n6193) );
  INVX0_HVT U4486 ( .A(n9072), .Y(n9080) );
  INVX0_HVT U4487 ( .A(n9072), .Y(n9079) );
  INVX0_HVT U4488 ( .A(n9072), .Y(n9077) );
  INVX0_HVT U4489 ( .A(n7592), .Y(n4453) );
  INVX0_HVT U4490 ( .A(n9025), .Y(n9072) );
  INVX0_HVT U4491 ( .A(n9025), .Y(n9071) );
  OAI22X1_HVT U4492 ( .A1(n4373), .A2(n6255), .A3(n5274), .A4(n4372), .Y(n845)
         );
  IBUFFX16_HVT U4493 ( .A(n9356), .Y(n4372) );
  INVX0_HVT U4494 ( .A(n4371), .Y(n4374) );
  INVX0_HVT U4495 ( .A(n4909), .Y(n4375) );
  OAI22X1_HVT U4496 ( .A1(n4376), .A2(n4562), .A3(n4520), .A4(n9567), .Y(n916)
         );
  INVX0_HVT U4497 ( .A(n7121), .Y(n7128) );
  INVX0_HVT U4498 ( .A(n5265), .Y(n5266) );
  INVX0_HVT U4499 ( .A(n4545), .Y(n4377) );
  INVX0_HVT U4500 ( .A(n4956), .Y(n4378) );
  INVX0_HVT U4501 ( .A(n10204), .Y(n9098) );
  INVX0_HVT U4502 ( .A(n9095), .Y(n4379) );
  INVX0_HVT U4503 ( .A(n4379), .Y(n4380) );
  OAI22X1_HVT U4504 ( .A1(n4381), .A2(n4504), .A3(n4662), .A4(n9684), .Y(n2491) );
  OAI22X1_HVT U4505 ( .A1(n4383), .A2(n4489), .A3(n4657), .A4(n4382), .Y(n2375) );
  IBUFFX16_HVT U4506 ( .A(data[10]), .Y(n4382) );
  INVX0_HVT U4507 ( .A(n7661), .Y(n4489) );
  OAI22X1_HVT U4508 ( .A1(n4384), .A2(n5860), .A3(n5244), .A4(n9860), .Y(n1011) );
  INVX0_HVT U4509 ( .A(n5253), .Y(n5254) );
  OAI21X2_HVT U4510 ( .A1(n6118), .A2(n5802), .A3(n5835), .Y(n5754) );
  INVX0_HVT U4511 ( .A(n5189), .Y(n5192) );
  INVX0_HVT U4512 ( .A(n6564), .Y(n6566) );
  INVX0_HVT U4513 ( .A(n6564), .Y(n6617) );
  INVX0_HVT U4514 ( .A(n9061), .Y(n9065) );
  NBUFFX2_HVT U4515 ( .A(n4399), .Y(n4385) );
  OAI22X1_HVT U4516 ( .A1(n4388), .A2(n4430), .A3(n4386), .A4(n4387), .Y(n2910) );
  IBUFFX16_HVT U4517 ( .A(n6822), .Y(n4386) );
  IBUFFX16_HVT U4518 ( .A(data[33]), .Y(n4387) );
  OAI22X1_HVT U4519 ( .A1(n4391), .A2(n4425), .A3(n4389), .A4(n4390), .Y(n2909) );
  OAI22X1_HVT U4520 ( .A1(n4394), .A2(n4425), .A3(n4392), .A4(n4393), .Y(n2908) );
  IBUFFX16_HVT U4521 ( .A(n6824), .Y(n4392) );
  IBUFFX16_HVT U4522 ( .A(data[31]), .Y(n4393) );
  NBUFFX2_HVT U4523 ( .A(n6142), .Y(n4395) );
  INVX0_HVT U4524 ( .A(n6142), .Y(n6175) );
  NBUFFX2_HVT U4525 ( .A(n6492), .Y(n4396) );
  NBUFFX2_HVT U4526 ( .A(n6485), .Y(n4397) );
  INVX0_HVT U4527 ( .A(n4239), .Y(n4398) );
  INVX0_HVT U4528 ( .A(n4528), .Y(n4399) );
  OAI22X1_HVT U4529 ( .A1(n4401), .A2(n4400), .A3(n4405), .A4(n9402), .Y(n3165) );
  OAI22X1_HVT U4530 ( .A1(n4404), .A2(n4402), .A3(n4405), .A4(n4403), .Y(n3161) );
  IBUFFX16_HVT U4531 ( .A(data[28]), .Y(n4403) );
  INVX0_HVT U4532 ( .A(n6333), .Y(n4405) );
  INVX0_HVT U4533 ( .A(n4405), .Y(n4406) );
  INVX0_HVT U4534 ( .A(n7154), .Y(n4407) );
  INVX0_HVT U4535 ( .A(n4407), .Y(n4408) );
  NBUFFX2_HVT U4536 ( .A(n6330), .Y(n4409) );
  INVX0_HVT U4537 ( .A(n6330), .Y(n6373) );
  NBUFFX2_HVT U4538 ( .A(n9252), .Y(n4410) );
  INVX0_HVT U4539 ( .A(n9252), .Y(n9287) );
  NBUFFX2_HVT U4540 ( .A(n6329), .Y(n4411) );
  INVX0_HVT U4541 ( .A(n6329), .Y(n6365) );
  INVX0_HVT U4542 ( .A(n6368), .Y(n4412) );
  INVX0_HVT U4543 ( .A(n4412), .Y(n4413) );
  INVX0_HVT U4544 ( .A(n6594), .Y(n6567) );
  INVX0_HVT U4545 ( .A(n6594), .Y(n6596) );
  INVX1_HVT U4546 ( .A(n5544), .Y(n10286) );
  INVX0_HVT U4547 ( .A(n5545), .Y(n4414) );
  INVX0_HVT U4548 ( .A(n4414), .Y(n4415) );
  INVX0_HVT U4549 ( .A(n9071), .Y(n9073) );
  INVX0_HVT U4550 ( .A(n9071), .Y(n9075) );
  INVX0_HVT U4551 ( .A(n9071), .Y(n9076) );
  INVX0_HVT U4552 ( .A(n7410), .Y(n7411) );
  INVX0_HVT U4553 ( .A(n7410), .Y(n7409) );
  INVX0_HVT U4554 ( .A(n9062), .Y(n9070) );
  INVX0_HVT U4555 ( .A(n9062), .Y(n9067) );
  INVX0_HVT U4556 ( .A(n9062), .Y(n9068) );
  INVX0_HVT U4557 ( .A(n9062), .Y(n9069) );
  INVX0_HVT U4558 ( .A(n9024), .Y(n9062) );
  INVX1_HVT U4559 ( .A(\ram[14][65] ), .Y(n4879) );
  INVX0_HVT U4560 ( .A(n4573), .Y(n4416) );
  NBUFFX2_HVT U4561 ( .A(n7207), .Y(n4417) );
  INVX0_HVT U4562 ( .A(n7207), .Y(n7245) );
  NBUFFX2_HVT U4563 ( .A(n7249), .Y(n4418) );
  INVX0_HVT U4564 ( .A(n6686), .Y(n6667) );
  INVX0_HVT U4565 ( .A(n6686), .Y(n6688) );
  NBUFFX2_HVT U4566 ( .A(n7037), .Y(n4419) );
  OAI22X1_HVT U4567 ( .A1(n4421), .A2(n4455), .A3(n4420), .A4(n9669), .Y(n3510) );
  IBUFFX16_HVT U4568 ( .A(n8950), .Y(n4420) );
  INVX0_HVT U4569 ( .A(n9297), .Y(n4422) );
  INVX0_HVT U4570 ( .A(n4639), .Y(n4423) );
  INVX0_HVT U4571 ( .A(n4423), .Y(n4424) );
  INVX0_HVT U4572 ( .A(n7466), .Y(n4425) );
  INVX0_HVT U4573 ( .A(n4425), .Y(n4426) );
  OAI22X1_HVT U4574 ( .A1(n4429), .A2(n4430), .A3(n4427), .A4(n4428), .Y(n2884) );
  IBUFFX16_HVT U4575 ( .A(n6821), .Y(n4427) );
  IBUFFX16_HVT U4576 ( .A(data[7]), .Y(n4428) );
  INVX0_HVT U4577 ( .A(n7466), .Y(n4430) );
  INVX0_HVT U4578 ( .A(n4430), .Y(n4431) );
  INVX0_HVT U4579 ( .A(n7410), .Y(n7412) );
  NBUFFX2_HVT U4580 ( .A(n4537), .Y(n4432) );
  INVX0_HVT U4581 ( .A(n6712), .Y(n6714) );
  INVX0_HVT U4582 ( .A(n6671), .Y(n6668) );
  INVX0_HVT U4583 ( .A(n6683), .Y(n6672) );
  INVX0_HVT U4584 ( .A(n4433), .Y(n7413) );
  INVX0_HVT U4585 ( .A(n7376), .Y(n7378) );
  INVX0_HVT U4586 ( .A(n10244), .Y(n4433) );
  INVX0_HVT U4587 ( .A(n4433), .Y(n4434) );
  OA22X1_HVT U4588 ( .A1(n4437), .A2(n4472), .A3(n4436), .A4(n9352), .Y(n4435)
         );
  IBUFFX16_HVT U4589 ( .A(n4435), .Y(n2124) );
  INVX0_HVT U4590 ( .A(n10352), .Y(n4438) );
  INVX0_HVT U4591 ( .A(n6175), .Y(n4439) );
  INVX0_HVT U4592 ( .A(n4461), .Y(n4440) );
  OAI22X1_HVT U4593 ( .A1(n4443), .A2(n4441), .A3(n4442), .A4(n6508), .Y(n111)
         );
  IBUFFX16_HVT U4594 ( .A(n9458), .Y(n4442) );
  INVX0_HVT U4595 ( .A(n6516), .Y(n6496) );
  INVX0_HVT U4596 ( .A(n4592), .Y(n4444) );
  INVX0_HVT U4597 ( .A(n4655), .Y(n4445) );
  INVX0_HVT U4598 ( .A(n4455), .Y(n4446) );
  INVX0_HVT U4599 ( .A(n7009), .Y(n4455) );
  INVX0_HVT U4600 ( .A(n4738), .Y(n4447) );
  INVX0_HVT U4601 ( .A(n4896), .Y(n4738) );
  INVX0_HVT U4602 ( .A(n4457), .Y(n4448) );
  INVX0_HVT U4603 ( .A(n6987), .Y(n4457) );
  OAI22X1_HVT U4604 ( .A1(n4450), .A2(n7651), .A3(n4508), .A4(n4449), .Y(n2413) );
  INVX0_HVT U4605 ( .A(n10220), .Y(n10217) );
  OAI22X1_HVT U4606 ( .A1(n4452), .A2(n4451), .A3(n4508), .A4(n9447), .Y(n2412) );
  OAI22X1_HVT U4607 ( .A1(n4454), .A2(n4453), .A3(n4508), .A4(n9444), .Y(n2411) );
  INVX0_HVT U4608 ( .A(n7599), .Y(n4467) );
  OAI22X1_HVT U4609 ( .A1(n4456), .A2(n4455), .A3(n4525), .A4(n9794), .Y(n3550) );
  OAI22X1_HVT U4610 ( .A1(n4458), .A2(n4457), .A3(n4476), .A4(n9733), .Y(n3531) );
  INVX1_HVT U4611 ( .A(n7652), .Y(n4487) );
  OA22X1_HVT U4612 ( .A1(n4460), .A2(n4601), .A3(n4512), .A4(n9519), .Y(n4459)
         );
  IBUFFX16_HVT U4613 ( .A(n4459), .Y(n3460) );
  INVX1_HVT U4614 ( .A(n4600), .Y(n4601) );
  INVX0_HVT U4615 ( .A(n10344), .Y(n4461) );
  INVX0_HVT U4616 ( .A(n4556), .Y(n4462) );
  INVX0_HVT U4617 ( .A(n10207), .Y(n4463) );
  INVX0_HVT U4618 ( .A(n4508), .Y(n4464) );
  INVX0_HVT U4619 ( .A(n9136), .Y(n4465) );
  INVX0_HVT U4620 ( .A(n4465), .Y(n4466) );
  OAI22X1_HVT U4621 ( .A1(n4468), .A2(n4467), .A3(n4664), .A4(n9627), .Y(n2472) );
  NOR2X1_HVT U4622 ( .A1(n5246), .A2(n9477), .Y(n4469) );
  IBUFFX16_HVT U4623 ( .A(n4469), .Y(n6000) );
  INVX0_HVT U4624 ( .A(n5244), .Y(n5245) );
  OAI22X1_HVT U4625 ( .A1(n4471), .A2(n4472), .A3(n6052), .A4(n4470), .Y(n2134) );
  IBUFFX16_HVT U4626 ( .A(n9383), .Y(n4470) );
  INVX0_HVT U4627 ( .A(n4280), .Y(n6045) );
  INVX0_HVT U4628 ( .A(n4434), .Y(n4472) );
  OAI22X1_HVT U4629 ( .A1(n4473), .A2(n5329), .A3(n4520), .A4(n4891), .Y(n831)
         );
  INVX0_HVT U4630 ( .A(n5246), .Y(n5247) );
  INVX0_HVT U4631 ( .A(n4467), .Y(n4474) );
  INVX0_HVT U4632 ( .A(n4955), .Y(n4475) );
  INVX0_HVT U4633 ( .A(n8936), .Y(n4476) );
  INVX0_HVT U4634 ( .A(n4476), .Y(n4477) );
  OAI22X1_HVT U4635 ( .A1(n4479), .A2(n4494), .A3(n4478), .A4(n9612), .Y(n3747) );
  INVX0_HVT U4636 ( .A(n4538), .Y(n4480) );
  INVX0_HVT U4637 ( .A(n4668), .Y(n4538) );
  NBUFFX2_HVT U4638 ( .A(n7025), .Y(n4481) );
  INVX0_HVT U4639 ( .A(n6522), .Y(n6523) );
  OA22X1_HVT U4640 ( .A1(n4483), .A2(n6693), .A3(n9367), .A4(n6537), .Y(n4482)
         );
  IBUFFX16_HVT U4641 ( .A(n4482), .Y(n81) );
  INVX0_HVT U4642 ( .A(n6671), .Y(n6684) );
  OAI22X1_HVT U4643 ( .A1(n4484), .A2(n6719), .A3(n4891), .A4(n4506), .Y(n63)
         );
  INVX0_HVT U4644 ( .A(n6708), .Y(n6706) );
  INVX0_HVT U4645 ( .A(n6515), .Y(n6538) );
  INVX0_HVT U4646 ( .A(n4527), .Y(n4485) );
  INVX0_HVT U4647 ( .A(n4824), .Y(n4527) );
  OAI22X1_HVT U4648 ( .A1(n4486), .A2(n4538), .A3(n4525), .A4(n9489), .Y(n3450) );
  OAI22X1_HVT U4649 ( .A1(n4488), .A2(n4487), .A3(n4269), .A4(n9492), .Y(n2427) );
  OAI22X1_HVT U4650 ( .A1(n4490), .A2(n4489), .A3(n4502), .A4(n9471), .Y(n2420) );
  OAI22X1_HVT U4651 ( .A1(n4491), .A2(n4453), .A3(n4657), .A4(n9441), .Y(n2410) );
  INVX0_HVT U4652 ( .A(n7053), .Y(n4492) );
  INVX0_HVT U4653 ( .A(n4492), .Y(n4493) );
  INVX0_HVT U4654 ( .A(n7238), .Y(n4494) );
  INVX0_HVT U4655 ( .A(n4494), .Y(n4495) );
  INVX0_HVT U4656 ( .A(n7239), .Y(n4496) );
  INVX0_HVT U4657 ( .A(n4496), .Y(n4497) );
  INVX0_HVT U4658 ( .A(n7239), .Y(n4498) );
  INVX0_HVT U4659 ( .A(n4498), .Y(n4499) );
  OAI22X1_HVT U4660 ( .A1(n4500), .A2(n5329), .A3(n4520), .A4(n9597), .Y(n926)
         );
  INVX0_HVT U4661 ( .A(n5259), .Y(n5255) );
  IBUFFX4_HVT U4662 ( .A(n5276), .Y(n4520) );
  INVX0_HVT U4663 ( .A(n7661), .Y(n4504) );
  OAI22X1_HVT U4664 ( .A1(n4501), .A2(n6574), .A3(n4621), .A4(n4770), .Y(n3216) );
  INVX0_HVT U4665 ( .A(n6569), .Y(n6570) );
  IBUFFX4_HVT U4666 ( .A(n9557), .Y(n4770) );
  INVX0_HVT U4667 ( .A(n9109), .Y(n4502) );
  INVX0_HVT U4668 ( .A(n4333), .Y(n4503) );
  OAI22X1_HVT U4669 ( .A1(n4505), .A2(n4504), .A3(n4269), .A4(n9781), .Y(n2522) );
  INVX0_HVT U4670 ( .A(n10353), .Y(n4506) );
  INVX0_HVT U4671 ( .A(n4506), .Y(n4507) );
  INVX0_HVT U4672 ( .A(n9082), .Y(n9128) );
  INVX0_HVT U4673 ( .A(n9083), .Y(n4508) );
  INVX0_HVT U4674 ( .A(n4465), .Y(n4509) );
  INVX0_HVT U4675 ( .A(n6611), .Y(n4510) );
  INVX0_HVT U4676 ( .A(n4510), .Y(n4511) );
  INVX0_HVT U4677 ( .A(n8927), .Y(n4512) );
  INVX0_HVT U4678 ( .A(n4512), .Y(n4513) );
  INVX0_HVT U4679 ( .A(n10380), .Y(n4514) );
  IBUFFX2_HVT U4680 ( .A(n8760), .Y(n5015) );
  INVX0_HVT U4681 ( .A(n9074), .Y(n4616) );
  INVX0_HVT U4682 ( .A(n9071), .Y(n9074) );
  OAI22X1_HVT U4683 ( .A1(n4515), .A2(n4670), .A3(n5010), .A4(n4903), .Y(n1370) );
  INVX0_HVT U4684 ( .A(n9288), .Y(n9294) );
  INVX0_HVT U4685 ( .A(n5268), .Y(n4516) );
  INVX0_HVT U4686 ( .A(n5268), .Y(n4517) );
  INVX0_HVT U4687 ( .A(n5268), .Y(n5276) );
  OAI22X1_HVT U4688 ( .A1(n4519), .A2(n5860), .A3(n4518), .A4(n9558), .Y(n913)
         );
  INVX0_HVT U4689 ( .A(n7130), .Y(n7133) );
  OAI22X1_HVT U4690 ( .A1(n4522), .A2(n4562), .A3(n4520), .A4(n4521), .Y(n855)
         );
  IBUFFX16_HVT U4691 ( .A(n9385), .Y(n4521) );
  INVX0_HVT U4692 ( .A(n7120), .Y(n7123) );
  OAI22X1_HVT U4693 ( .A1(n4524), .A2(n4562), .A3(n5257), .A4(n4523), .Y(n947)
         );
  IBUFFX16_HVT U4694 ( .A(n9661), .Y(n4523) );
  INVX0_HVT U4695 ( .A(n7131), .Y(n7137) );
  IBUFFX4_HVT U4696 ( .A(n7137), .Y(n4562) );
  INVX0_HVT U4697 ( .A(n5246), .Y(n5256) );
  AO22X1_HVT U4698 ( .A1(\ram[4][89] ), .A2(n6164), .A3(n6219), .A4(n9574), 
        .Y(n1174) );
  INVX0_HVT U4699 ( .A(n7662), .Y(n4752) );
  INVX0_HVT U4700 ( .A(n8912), .Y(n4525) );
  INVX0_HVT U4701 ( .A(n4525), .Y(n4526) );
  OAI22X1_HVT U4702 ( .A1(n4810), .A2(n4527), .A3(n4931), .A4(n9609), .Y(n3490) );
  INVX0_HVT U4703 ( .A(n10367), .Y(n4528) );
  INVX0_HVT U4704 ( .A(n4625), .Y(n4529) );
  INVX0_HVT U4705 ( .A(n7350), .Y(n8827) );
  INVX0_HVT U4706 ( .A(n7350), .Y(n6029) );
  INVX0_HVT U4707 ( .A(n7350), .Y(n8836) );
  NBUFFX2_HVT U4708 ( .A(n9052), .Y(n4530) );
  NBUFFX2_HVT U4709 ( .A(n9047), .Y(n4531) );
  NBUFFX2_HVT U4710 ( .A(n9046), .Y(n4532) );
  NBUFFX2_HVT U4711 ( .A(n9034), .Y(n4533) );
  INVX0_HVT U4712 ( .A(n6159), .Y(n6163) );
  NBUFFX2_HVT U4713 ( .A(n7230), .Y(n4534) );
  NBUFFX2_HVT U4714 ( .A(n7225), .Y(n4535) );
  INVX0_HVT U4715 ( .A(n9099), .Y(n4536) );
  INVX0_HVT U4716 ( .A(n4536), .Y(n4537) );
  OAI22X1_HVT U4717 ( .A1(n4539), .A2(n4538), .A3(n4643), .A4(n9973), .Y(n3607) );
  NBUFFX2_HVT U4718 ( .A(n7231), .Y(n4540) );
  INVX0_HVT U4719 ( .A(n7646), .Y(n4653) );
  NBUFFX2_HVT U4720 ( .A(n6989), .Y(n4541) );
  INVX0_HVT U4721 ( .A(n4575), .Y(n4542) );
  INVX0_HVT U4722 ( .A(n7010), .Y(n4575) );
  INVX0_HVT U4723 ( .A(n5257), .Y(n4543) );
  INVX0_HVT U4724 ( .A(n5257), .Y(n4544) );
  INVX0_HVT U4725 ( .A(n5257), .Y(n5251) );
  INVX0_HVT U4726 ( .A(n10238), .Y(n4545) );
  INVX0_HVT U4727 ( .A(n10238), .Y(n7358) );
  OAI22X1_HVT U4728 ( .A1(n4548), .A2(n4546), .A3(n4558), .A4(n4547), .Y(n3276) );
  IBUFFX16_HVT U4729 ( .A(n9739), .Y(n4547) );
  INVX0_HVT U4730 ( .A(n6373), .Y(n4549) );
  INVX0_HVT U4731 ( .A(n6374), .Y(n4550) );
  INVX0_HVT U4732 ( .A(n6364), .Y(n4551) );
  INVX0_HVT U4733 ( .A(n6365), .Y(n4552) );
  INVX0_HVT U4734 ( .A(n5200), .Y(n10331) );
  INVX0_HVT U4735 ( .A(n10315), .Y(n6767) );
  OAI22X1_HVT U4736 ( .A1(n4554), .A2(n6574), .A3(n4743), .A4(n4553), .Y(n3182) );
  IBUFFX16_HVT U4737 ( .A(n9455), .Y(n4553) );
  INVX0_HVT U4738 ( .A(n6574), .Y(n6576) );
  OAI22X1_HVT U4739 ( .A1(n4555), .A2(n6589), .A3(n4274), .A4(n9411), .Y(n3168) );
  INVX0_HVT U4740 ( .A(n6342), .Y(n4556) );
  INVX0_HVT U4741 ( .A(n4743), .Y(n4557) );
  INVX0_HVT U4742 ( .A(n6349), .Y(n4558) );
  INVX0_HVT U4743 ( .A(n4558), .Y(n4559) );
  OAI22X1_HVT U4744 ( .A1(n4561), .A2(n4560), .A3(n9678), .A4(n6504), .Y(n185)
         );
  OAI22X1_HVT U4745 ( .A1(n4563), .A2(n4562), .A3(n5263), .A4(n9648), .Y(n943)
         );
  INVX0_HVT U4746 ( .A(n4463), .Y(n7627) );
  INVX0_HVT U4747 ( .A(n7602), .Y(n7590) );
  INVX0_HVT U4748 ( .A(n7153), .Y(n7198) );
  INVX0_HVT U4749 ( .A(n5467), .Y(n4564) );
  INVX0_HVT U4750 ( .A(n6767), .Y(n5274) );
  OAI22X1_HVT U4751 ( .A1(n4565), .A2(n4755), .A3(n4588), .A4(n9882), .Y(n3578) );
  OAI22X1_HVT U4752 ( .A1(n4567), .A2(n4566), .A3(n4645), .A4(n9633), .Y(n1450) );
  INVX0_HVT U4753 ( .A(n7253), .Y(n4568) );
  INVX0_HVT U4754 ( .A(n7245), .Y(n4569) );
  INVX0_HVT U4755 ( .A(n7244), .Y(n4570) );
  INVX0_HVT U4756 ( .A(n6152), .Y(n4571) );
  INVX0_HVT U4757 ( .A(n4571), .Y(n4572) );
  INVX0_HVT U4758 ( .A(n7029), .Y(n4573) );
  INVX0_HVT U4759 ( .A(n4573), .Y(n4574) );
  OAI22X1_HVT U4760 ( .A1(n4577), .A2(n4575), .A3(n4588), .A4(n4576), .Y(n3641) );
  OAI22X1_HVT U4761 ( .A1(n4579), .A2(n4672), .A3(n4578), .A4(n4693), .Y(n327)
         );
  IBUFFX16_HVT U4762 ( .A(n6842), .Y(n4578) );
  IBUFFX4_HVT U4763 ( .A(n9337), .Y(n4693) );
  INVX0_HVT U4764 ( .A(n7253), .Y(n7257) );
  INVX0_HVT U4765 ( .A(n4472), .Y(n4580) );
  INVX0_HVT U4766 ( .A(n7392), .Y(n4581) );
  NBUFFX2_HVT U4767 ( .A(n7188), .Y(n4582) );
  NBUFFX2_HVT U4768 ( .A(n18), .Y(n4583) );
  INVX0_HVT U4769 ( .A(n18), .Y(n7112) );
  IBUFFX2_HVT U4770 ( .A(n4759), .Y(n8) );
  INVX0_HVT U4771 ( .A(n7074), .Y(n7082) );
  INVX0_HVT U4772 ( .A(n7074), .Y(n7081) );
  INVX0_HVT U4773 ( .A(n7074), .Y(n7080) );
  INVX0_HVT U4774 ( .A(n7074), .Y(n7079) );
  INVX0_HVT U4775 ( .A(n10171), .Y(n7429) );
  NBUFFX2_HVT U4776 ( .A(n8933), .Y(n4584) );
  INVX0_HVT U4777 ( .A(n7359), .Y(n7360) );
  INVX0_HVT U4778 ( .A(n7603), .Y(n4585) );
  OAI22X1_HVT U4779 ( .A1(n4587), .A2(n4627), .A3(n4586), .A4(n9983), .Y(n1562) );
  IBUFFX16_HVT U4780 ( .A(n9299), .Y(n4586) );
  INVX0_HVT U4781 ( .A(n8935), .Y(n4588) );
  INVX0_HVT U4782 ( .A(n4588), .Y(n4589) );
  OAI22X1_HVT U4783 ( .A1(n4591), .A2(n4762), .A3(n4590), .A4(n9723), .Y(n1224) );
  IBUFFX16_HVT U4784 ( .A(n6195), .Y(n4590) );
  INVX1_HVT U4785 ( .A(data[139]), .Y(n9723) );
  INVX0_HVT U4786 ( .A(n7040), .Y(n4592) );
  INVX0_HVT U4787 ( .A(n4592), .Y(n4593) );
  OAI22X1_HVT U4788 ( .A1(n4595), .A2(n7363), .A3(n6053), .A4(n4594), .Y(n2135) );
  INVX0_HVT U4789 ( .A(n7381), .Y(n7383) );
  MUX41X1_HVT U4790 ( .A1(n7836), .A3(n7838), .A2(n7837), .A4(n7839), .S0(
        n6399), .S1(n5637), .Y(q[26]) );
  INVX0_HVT U4791 ( .A(n6233), .Y(n4632) );
  INVX0_HVT U4792 ( .A(n6232), .Y(n6233) );
  OAI22X1_HVT U4793 ( .A1(n4818), .A2(n4605), .A3(n6052), .A4(n9480), .Y(n2167) );
  INVX0_HVT U4794 ( .A(n7382), .Y(n7384) );
  INVX0_HVT U4795 ( .A(n7603), .Y(n7605) );
  INVX0_HVT U4796 ( .A(n7602), .Y(n7634) );
  OAI22X1_HVT U4797 ( .A1(n4598), .A2(n4629), .A3(n4596), .A4(n4597), .Y(n3654) );
  IBUFFX16_HVT U4798 ( .A(n9335), .Y(n4597) );
  NBUFFX2_HVT U4799 ( .A(n4513), .Y(n4599) );
  INVX0_HVT U4800 ( .A(n7633), .Y(n7635) );
  INVX0_HVT U4801 ( .A(n4463), .Y(n7637) );
  INVX0_HVT U4802 ( .A(n7602), .Y(n7636) );
  INVX0_HVT U4803 ( .A(n7603), .Y(n7639) );
  INVX0_HVT U4804 ( .A(n6998), .Y(n4600) );
  OAI22X1_HVT U4805 ( .A1(n4603), .A2(n4614), .A3(n4602), .A4(n4903), .Y(n346)
         );
  IBUFFX16_HVT U4806 ( .A(n6861), .Y(n4602) );
  IBUFFX4_HVT U4807 ( .A(data[29]), .Y(n4903) );
  INVX0_HVT U4808 ( .A(n7017), .Y(n7025) );
  INVX0_HVT U4809 ( .A(n7017), .Y(n7024) );
  INVX0_HVT U4810 ( .A(n7017), .Y(n7023) );
  INVX0_HVT U4811 ( .A(n7017), .Y(n7022) );
  INVX0_HVT U4812 ( .A(n6968), .Y(n7017) );
  INVX0_HVT U4813 ( .A(n7727), .Y(n4604) );
  INVX0_HVT U4814 ( .A(n6012), .Y(n6013) );
  INVX0_HVT U4815 ( .A(n7253), .Y(n7258) );
  INVX0_HVT U4816 ( .A(n7416), .Y(n4605) );
  INVX0_HVT U4817 ( .A(n4605), .Y(n4606) );
  OA22X1_HVT U4818 ( .A1(n4609), .A2(n6564), .A3(n4743), .A4(n4608), .Y(n4607)
         );
  NBUFFX2_HVT U4819 ( .A(n9041), .Y(n4610) );
  NBUFFX2_HVT U4820 ( .A(n9035), .Y(n4611) );
  INVX0_HVT U4821 ( .A(n4200), .Y(n4612) );
  INVX0_HVT U4822 ( .A(n7585), .Y(n4613) );
  INVX0_HVT U4823 ( .A(n7016), .Y(n7021) );
  INVX0_HVT U4824 ( .A(n7355), .Y(n7390) );
  INVX0_HVT U4825 ( .A(n7355), .Y(n7370) );
  INVX0_HVT U4826 ( .A(n7355), .Y(n7357) );
  INVX0_HVT U4827 ( .A(n7355), .Y(n7356) );
  INVX1_HVT U4828 ( .A(n10237), .Y(n7355) );
  INVX0_HVT U4829 ( .A(n7044), .Y(n4614) );
  INVX0_HVT U4830 ( .A(n4614), .Y(n4615) );
  INVX0_HVT U4831 ( .A(n4896), .Y(n4680) );
  INVX0_HVT U4832 ( .A(n10113), .Y(n9034) );
  INVX0_HVT U4833 ( .A(n10113), .Y(n9046) );
  INVX1_HVT U4834 ( .A(n10115), .Y(n10113) );
  OAI22X1_HVT U4835 ( .A1(n4618), .A2(n4629), .A3(n4616), .A4(n4617), .Y(n3712) );
  IBUFFX16_HVT U4836 ( .A(n9509), .Y(n4617) );
  NBUFFX2_HVT U4837 ( .A(n6338), .Y(n4619) );
  OAI22X1_HVT U4838 ( .A1(n4620), .A2(n4546), .A3(n4621), .A4(n9936), .Y(n3339) );
  INVX0_HVT U4839 ( .A(n6344), .Y(n4621) );
  INVX0_HVT U4840 ( .A(n4621), .Y(n4622) );
  INVX0_HVT U4841 ( .A(n7393), .Y(n7394) );
  INVX0_HVT U4842 ( .A(n7393), .Y(n7372) );
  INVX0_HVT U4843 ( .A(n7392), .Y(n7396) );
  INVX0_HVT U4844 ( .A(n4472), .Y(n7395) );
  INVX0_HVT U4845 ( .A(n7392), .Y(n7397) );
  INVX0_HVT U4846 ( .A(n7393), .Y(n7373) );
  OAI22X1_HVT U4847 ( .A1(n4624), .A2(n4627), .A3(n4623), .A4(n9980), .Y(n1561) );
  IBUFFX16_HVT U4848 ( .A(n9300), .Y(n4623) );
  INVX0_HVT U4849 ( .A(n5706), .Y(n4625) );
  INVX0_HVT U4850 ( .A(n4625), .Y(n4626) );
  INVX0_HVT U4851 ( .A(n5704), .Y(n4627) );
  INVX0_HVT U4852 ( .A(n4627), .Y(n4628) );
  INVX0_HVT U4853 ( .A(n6604), .Y(n6606) );
  INVX0_HVT U4854 ( .A(n6604), .Y(n6573) );
  INVX0_HVT U4855 ( .A(n6604), .Y(n6619) );
  INVX0_HVT U4856 ( .A(n7227), .Y(n4629) );
  INVX0_HVT U4857 ( .A(n4629), .Y(n4630) );
  INVX0_HVT U4858 ( .A(n10149), .Y(n10147) );
  INVX0_HVT U4859 ( .A(n7253), .Y(n7255) );
  OA22X1_HVT U4860 ( .A1(n4633), .A2(n5501), .A3(n4632), .A4(n9699), .Y(n4631)
         );
  OAI22X1_HVT U4861 ( .A1(n4636), .A2(n5442), .A3(n4634), .A4(n4635), .Y(n640)
         );
  IBUFFX16_HVT U4862 ( .A(n6263), .Y(n4634) );
  IBUFFX16_HVT U4863 ( .A(n9508), .Y(n4635) );
  NBUFFX2_HVT U4864 ( .A(n7219), .Y(n4637) );
  NBUFFX2_HVT U4865 ( .A(n7218), .Y(n4638) );
  NAND2X0_HVT U4866 ( .A1(n28), .A2(n10377), .Y(n4639) );
  INVX0_HVT U4867 ( .A(n4648), .Y(n4640) );
  OAI22X1_HVT U4868 ( .A1(n4641), .A2(n4914), .A3(n4645), .A4(n10010), .Y(
        n1571) );
  OAI22X1_HVT U4869 ( .A1(n4642), .A2(n4755), .A3(n4643), .A4(n9486), .Y(n3449) );
  IBUFFX4_HVT U4870 ( .A(n8923), .Y(n4643) );
  OAI22X1_HVT U4871 ( .A1(n4644), .A2(n4755), .A3(n4643), .A4(n9483), .Y(n3448) );
  INVX0_HVT U4872 ( .A(n5200), .Y(n10334) );
  MUX41X1_HVT U4873 ( .A1(n7905), .A3(n7903), .A2(n7906), .A4(n7904), .S0(
        n8761), .S1(n5828), .Y(q[43]) );
  INVX0_HVT U4874 ( .A(n9285), .Y(n4645) );
  INVX0_HVT U4875 ( .A(n4645), .Y(n4646) );
  INVX0_HVT U4876 ( .A(n7362), .Y(n4647) );
  INVX0_HVT U4877 ( .A(n5681), .Y(n4648) );
  INVX0_HVT U4878 ( .A(n4648), .Y(n4649) );
  MUX41X1_HVT U4879 ( .A1(\ram[2][116] ), .A3(\ram[0][116] ), .A2(
        \ram[3][116] ), .A4(\ram[1][116] ), .S0(n5863), .S1(n5134), .Y(n8197)
         );
  INVX0_HVT U4880 ( .A(n4582), .Y(n4650) );
  INVX0_HVT U4881 ( .A(n7152), .Y(n7188) );
  MUX41X1_HVT U4882 ( .A1(\ram[4][0] ), .A3(\ram[6][0] ), .A2(\ram[5][0] ), 
        .A4(\ram[7][0] ), .S0(n4883), .S1(n5165), .Y(n7736) );
  MUX41X1_HVT U4883 ( .A1(\ram[7][13] ), .A3(\ram[5][13] ), .A2(\ram[6][13] ), 
        .A4(\ram[4][13] ), .S0(n5125), .S1(n4666), .Y(n7788) );
  INVX0_HVT U4884 ( .A(n5576), .Y(n5580) );
  IBUFFX4_HVT U4885 ( .A(n7695), .Y(n4666) );
  INVX0_HVT U4886 ( .A(n9257), .Y(n4729) );
  INVX0_HVT U4887 ( .A(n9082), .Y(n4651) );
  INVX0_HVT U4888 ( .A(n9082), .Y(n9127) );
  INVX0_HVT U4889 ( .A(n4655), .Y(n4652) );
  OAI22X1_HVT U4890 ( .A1(n4654), .A2(n4653), .A3(n4657), .A4(n9552), .Y(n2447) );
  INVX0_HVT U4891 ( .A(n9123), .Y(n4655) );
  INVX0_HVT U4892 ( .A(n4655), .Y(n4656) );
  INVX0_HVT U4893 ( .A(n9124), .Y(n4657) );
  INVX0_HVT U4894 ( .A(n4465), .Y(n4658) );
  OAI22X1_HVT U4895 ( .A1(n4660), .A2(n4659), .A3(n4664), .A4(n9384), .Y(n2391) );
  IBUFFX16_HVT U4896 ( .A(n7656), .Y(n4659) );
  OAI22X1_HVT U4897 ( .A1(n4661), .A2(n7598), .A3(n4662), .A4(n9378), .Y(n2389) );
  INVX0_HVT U4898 ( .A(n9132), .Y(n4662) );
  INVX0_HVT U4899 ( .A(n4662), .Y(n4663) );
  INVX0_HVT U4900 ( .A(n9134), .Y(n4664) );
  INVX0_HVT U4901 ( .A(n4664), .Y(n4665) );
  MUX41X1_HVT U4902 ( .A1(\ram[13][99] ), .A3(\ram[15][99] ), .A2(
        \ram[12][99] ), .A4(\ram[14][99] ), .S0(n8826), .S1(n5337), .Y(n8126)
         );
  MUX41X1_HVT U4903 ( .A1(\ram[11][61] ), .A3(\ram[9][61] ), .A2(\ram[10][61] ), .A4(\ram[8][61] ), .S0(n4898), .S1(n4666), .Y(n7975) );
  INVX0_HVT U4904 ( .A(n18), .Y(n4667) );
  INVX0_HVT U4905 ( .A(n5934), .Y(n5935) );
  INVX0_HVT U4906 ( .A(n51), .Y(n5934) );
  INVX0_HVT U4907 ( .A(n7007), .Y(n4668) );
  INVX0_HVT U4908 ( .A(n7006), .Y(n4669) );
  INVX0_HVT U4909 ( .A(n4952), .Y(n4670) );
  OAI22X1_HVT U4910 ( .A1(n4671), .A2(n4672), .A3(n6838), .A4(n9564), .Y(n403)
         );
  INVX0_HVT U4911 ( .A(n7035), .Y(n4672) );
  INVX0_HVT U4912 ( .A(n4672), .Y(n4673) );
  OAI22X1_HVT U4913 ( .A1(n4674), .A2(n4676), .A3(n6852), .A4(n9441), .Y(n362)
         );
  INVX0_HVT U4914 ( .A(n6848), .Y(n6849) );
  INVX0_HVT U4915 ( .A(n4676), .Y(n4675) );
  INVX0_HVT U4916 ( .A(n7044), .Y(n4676) );
  INVX0_HVT U4917 ( .A(n4676), .Y(n4677) );
  INVX0_HVT U4918 ( .A(n5631), .Y(n5622) );
  NBUFFX2_HVT U4919 ( .A(n6019), .Y(n7352) );
  OAI22X1_HVT U4920 ( .A1(n4679), .A2(n4854), .A3(n4678), .A4(n9537), .Y(n3466) );
  OAI22X1_HVT U4921 ( .A1(n4681), .A2(n4680), .A3(n4839), .A4(n9352), .Y(n1356) );
  INVX0_HVT U4922 ( .A(n4750), .Y(n4682) );
  INVX0_HVT U4923 ( .A(n7640), .Y(n4750) );
  INVX0_HVT U4924 ( .A(n9090), .Y(n4683) );
  INVX0_HVT U4925 ( .A(n4536), .Y(n4684) );
  INVX0_HVT U4926 ( .A(n10204), .Y(n9105) );
  NBUFFX2_HVT U4927 ( .A(n6360), .Y(n4685) );
  NBUFFX2_HVT U4928 ( .A(n6360), .Y(n4686) );
  OAI22X1_HVT U4929 ( .A1(n4687), .A2(n6586), .A3(n4313), .A4(n9513), .Y(n3202) );
  INVX0_HVT U4930 ( .A(n6581), .Y(n6583) );
  INVX0_HVT U4931 ( .A(n9260), .Y(n4688) );
  INVX0_HVT U4932 ( .A(n4688), .Y(n4689) );
  NBUFFX2_HVT U4933 ( .A(n9274), .Y(n4690) );
  NBUFFX2_HVT U4934 ( .A(n9268), .Y(n4691) );
  NBUFFX2_HVT U4935 ( .A(n9263), .Y(n4692) );
  OAI22X1_HVT U4936 ( .A1(n4694), .A2(n4727), .A3(n4780), .A4(n4693), .Y(n1351) );
  NBUFFX2_HVT U4937 ( .A(n9269), .Y(n4695) );
  INVX0_HVT U4938 ( .A(n6147), .Y(n4696) );
  INVX0_HVT U4939 ( .A(n4696), .Y(n4697) );
  NBUFFX2_HVT U4940 ( .A(n8922), .Y(n4698) );
  INVX0_HVT U4941 ( .A(n4933), .Y(n4699) );
  INVX0_HVT U4942 ( .A(n4719), .Y(n4700) );
  INVX0_HVT U4943 ( .A(n9296), .Y(n4701) );
  NBUFFX2_HVT U4944 ( .A(n9253), .Y(n4702) );
  INVX0_HVT U4945 ( .A(n5052), .Y(n9253) );
  INVX0_HVT U4946 ( .A(n9253), .Y(n9297) );
  INVX0_HVT U4947 ( .A(n8895), .Y(n4703) );
  NBUFFX2_HVT U4948 ( .A(n7268), .Y(n4704) );
  INVX0_HVT U4949 ( .A(n7268), .Y(n5762) );
  IBUFFX2_HVT U4950 ( .A(n9275), .Y(n4893) );
  INVX0_HVT U4951 ( .A(n9276), .Y(n4780) );
  NBUFFX2_HVT U4952 ( .A(n4776), .Y(n4705) );
  INVX0_HVT U4953 ( .A(n4778), .Y(n6161) );
  INVX0_HVT U4954 ( .A(n5501), .Y(n4706) );
  NBUFFX2_HVT U4955 ( .A(n6340), .Y(n4707) );
  NBUFFX2_HVT U4956 ( .A(n6345), .Y(n4708) );
  NBUFFX2_HVT U4957 ( .A(n7163), .Y(n4709) );
  INVX0_HVT U4958 ( .A(n5777), .Y(n4734) );
  INVX0_HVT U4959 ( .A(n5663), .Y(n4710) );
  OAI22X1_HVT U4960 ( .A1(n4712), .A2(n4741), .A3(n4943), .A4(n4711), .Y(n1349) );
  OAI22X1_HVT U4961 ( .A1(n4713), .A2(n4741), .A3(n4729), .A4(n4891), .Y(n1343) );
  IBUFFX4_HVT U4962 ( .A(data[2]), .Y(n4891) );
  NBUFFX2_HVT U4963 ( .A(n6983), .Y(n4714) );
  NBUFFX2_HVT U4964 ( .A(n6983), .Y(n4715) );
  INVX0_HVT U4965 ( .A(n4957), .Y(n4716) );
  MUX41X1_HVT U4966 ( .A1(\ram[14][113] ), .A3(\ram[12][113] ), .A2(
        \ram[15][113] ), .A4(\ram[13][113] ), .S0(n5821), .S1(n7691), .Y(n8182) );
  OAI22X1_HVT U4967 ( .A1(n4717), .A2(n4741), .A3(n4729), .A4(n9501), .Y(n1406) );
  INVX0_HVT U4968 ( .A(n6036), .Y(n4718) );
  INVX0_HVT U4969 ( .A(n10282), .Y(n4719) );
  INVX0_HVT U4970 ( .A(n4719), .Y(n4720) );
  OR2X1_HVT U4971 ( .A1(n4721), .A2(n4755), .Y(n5081) );
  NBUFFX2_HVT U4972 ( .A(n7059), .Y(n4722) );
  NBUFFX2_HVT U4973 ( .A(n7060), .Y(n4723) );
  INVX0_HVT U4974 ( .A(n9120), .Y(n4724) );
  INVX0_HVT U4975 ( .A(n9128), .Y(n4725) );
  INVX0_HVT U4976 ( .A(n4651), .Y(n4726) );
  INVX0_HVT U4977 ( .A(n5688), .Y(n4727) );
  INVX0_HVT U4978 ( .A(n4727), .Y(n4728) );
  OAI22X1_HVT U4979 ( .A1(n4730), .A2(n4731), .A3(n4729), .A4(n9447), .Y(n1388) );
  INVX0_HVT U4980 ( .A(n5711), .Y(n4731) );
  INVX0_HVT U4981 ( .A(n4953), .Y(n4732) );
  OAI22X1_HVT U4982 ( .A1(n4733), .A2(n4914), .A3(n4943), .A4(n9358), .Y(n1358) );
  MUX41X1_HVT U4983 ( .A1(\ram[7][52] ), .A3(\ram[5][52] ), .A2(\ram[6][52] ), 
        .A4(\ram[4][52] ), .S0(n5894), .S1(n4734), .Y(n7941) );
  INVX0_HVT U4984 ( .A(n9088), .Y(n4735) );
  INVX0_HVT U4985 ( .A(n4735), .Y(n4736) );
  INVX1_HVT U4986 ( .A(n7121), .Y(n4737) );
  OAI22X1_HVT U4987 ( .A1(n4739), .A2(n4738), .A3(n4893), .A4(n9955), .Y(n1553) );
  OAI22X1_HVT U4988 ( .A1(n4740), .A2(n4741), .A3(n4780), .A4(n9420), .Y(n1379) );
  INVX0_HVT U4989 ( .A(n5689), .Y(n4741) );
  INVX0_HVT U4990 ( .A(n4727), .Y(n4742) );
  INVX0_HVT U4991 ( .A(n6344), .Y(n4743) );
  INVX0_HVT U4992 ( .A(n4743), .Y(n4744) );
  OAI22X1_HVT U4993 ( .A1(n4746), .A2(n6574), .A3(n4313), .A4(n4745), .Y(n3167) );
  IBUFFX16_HVT U4994 ( .A(data[34]), .Y(n4745) );
  INVX0_HVT U4995 ( .A(n6589), .Y(n6590) );
  INVX0_HVT U4996 ( .A(n10350), .Y(n4747) );
  INVX0_HVT U4997 ( .A(n10351), .Y(n10350) );
  INVX0_HVT U4998 ( .A(n4947), .Y(n4748) );
  INVX0_HVT U4999 ( .A(n4748), .Y(n4749) );
  INVX0_HVT U5000 ( .A(n4774), .Y(n4755) );
  OAI22X1_HVT U5001 ( .A1(n4751), .A2(n4750), .A3(n4798), .A4(n9417), .Y(n2402) );
  OAI22X1_HVT U5002 ( .A1(n4753), .A2(n4752), .A3(n4796), .A4(n4894), .Y(n2401) );
  IBUFFX4_HVT U5003 ( .A(n9415), .Y(n4894) );
  OAI22X1_HVT U5004 ( .A1(n5842), .A2(n4851), .A3(n5841), .A4(n9468), .Y(n4754) );
  OAI22X1_HVT U5005 ( .A1(n4757), .A2(n4755), .A3(n4931), .A4(n4756), .Y(n3400) );
  IBUFFX16_HVT U5006 ( .A(n9342), .Y(n4756) );
  INVX0_HVT U5007 ( .A(n9296), .Y(n9298) );
  INVX0_HVT U5008 ( .A(n9296), .Y(n9299) );
  INVX0_HVT U5009 ( .A(n9296), .Y(n9300) );
  INVX0_HVT U5010 ( .A(n9297), .Y(n9304) );
  INVX0_HVT U5011 ( .A(n9297), .Y(n9302) );
  INVX0_HVT U5012 ( .A(n9297), .Y(n9303) );
  INVX0_HVT U5013 ( .A(n4933), .Y(n4758) );
  INVX0_HVT U5014 ( .A(n8785), .Y(n5888) );
  NAND2X0_HVT U5015 ( .A1(n5106), .A2(n7544), .Y(n4759) );
  NBUFFX2_HVT U5016 ( .A(n7019), .Y(n4760) );
  NBUFFX2_HVT U5017 ( .A(n7018), .Y(n4761) );
  INVX0_HVT U5018 ( .A(n6142), .Y(n4762) );
  NBUFFX2_HVT U5019 ( .A(n52), .Y(n4763) );
  INVX0_HVT U5020 ( .A(n52), .Y(n6998) );
  INVX0_HVT U5021 ( .A(n9296), .Y(n9301) );
  INVX0_HVT U5022 ( .A(n4948), .Y(n4764) );
  INVX0_HVT U5023 ( .A(n4948), .Y(n4765) );
  OAI22X1_HVT U5024 ( .A1(n4767), .A2(n4849), .A3(n4766), .A4(n9346), .Y(n1354) );
  IBUFFX16_HVT U5025 ( .A(n9261), .Y(n4766) );
  OAI22X1_HVT U5026 ( .A1(n4769), .A2(n4844), .A3(n4935), .A4(n4768), .Y(n3457) );
  OAI22X1_HVT U5027 ( .A1(n4771), .A2(n4854), .A3(n4931), .A4(n4770), .Y(n3472) );
  INVX0_HVT U5028 ( .A(n4847), .Y(n4772) );
  INVX0_HVT U5029 ( .A(n9120), .Y(n9124) );
  INVX0_HVT U5030 ( .A(n9120), .Y(n9126) );
  INVX0_HVT U5031 ( .A(n5698), .Y(n4773) );
  INVX0_HVT U5032 ( .A(n4775), .Y(n4774) );
  INVX0_HVT U5033 ( .A(n6986), .Y(n4775) );
  INVX0_HVT U5034 ( .A(n4775), .Y(n4776) );
  INVX0_HVT U5035 ( .A(n7011), .Y(n4782) );
  INVX0_HVT U5036 ( .A(n10123), .Y(n8922) );
  INVX0_HVT U5037 ( .A(n10125), .Y(n10123) );
  MUX41X1_HVT U5038 ( .A1(n7876), .A3(n7878), .A2(n7875), .A4(n7877), .S0(
        n5101), .S1(n5622), .Y(q[36]) );
  INVX0_HVT U5039 ( .A(n6158), .Y(n4777) );
  INVX0_HVT U5040 ( .A(n4777), .Y(n4778) );
  OAI22X1_HVT U5041 ( .A1(n4779), .A2(n4680), .A3(n4780), .A4(n10023), .Y(
        n1575) );
  IBUFFX16_HVT U5042 ( .A(\ram[5][234] ), .Y(n4779) );
  MUX41X1_HVT U5043 ( .A1(\ram[13][78] ), .A3(\ram[15][78] ), .A2(
        \ram[12][78] ), .A4(\ram[14][78] ), .S0(n4939), .S1(n5658), .Y(n8042)
         );
  NBUFFX2_HVT U5044 ( .A(n8921), .Y(n4781) );
  OAI22X1_HVT U5045 ( .A1(n4784), .A2(n4782), .A3(n4935), .A4(n4783), .Y(n3416) );
  IBUFFX16_HVT U5046 ( .A(n9389), .Y(n4783) );
  INVX0_HVT U5047 ( .A(n9119), .Y(n9122) );
  INVX0_HVT U5048 ( .A(n9119), .Y(n9121) );
  INVX0_HVT U5049 ( .A(n9119), .Y(n9123) );
  INVX0_HVT U5050 ( .A(n4651), .Y(n9131) );
  INVX0_HVT U5051 ( .A(n9127), .Y(n9130) );
  INVX0_HVT U5052 ( .A(n9127), .Y(n9129) );
  INVX0_HVT U5053 ( .A(n9127), .Y(n9133) );
  INVX0_HVT U5054 ( .A(n9127), .Y(n9136) );
  INVX0_HVT U5055 ( .A(n9128), .Y(n9135) );
  INVX0_HVT U5056 ( .A(n7297), .Y(n8828) );
  INVX0_HVT U5057 ( .A(n7054), .Y(n4785) );
  MUX41X1_HVT U5058 ( .A1(\ram[0][40] ), .A3(\ram[2][40] ), .A2(\ram[1][40] ), 
        .A4(\ram[3][40] ), .S0(n8817), .S1(n4793), .Y(n7894) );
  NBUFFX2_HVT U5059 ( .A(n4924), .Y(n4786) );
  INVX0_HVT U5060 ( .A(n8946), .Y(n4787) );
  INVX0_HVT U5061 ( .A(n4787), .Y(n4788) );
  INVX0_HVT U5062 ( .A(n4808), .Y(n4789) );
  INVX0_HVT U5063 ( .A(n8855), .Y(n4808) );
  INVX0_HVT U5064 ( .A(n10133), .Y(n4790) );
  INVX0_HVT U5065 ( .A(n4790), .Y(n4791) );
  INVX0_HVT U5066 ( .A(n9128), .Y(n9132) );
  INVX0_HVT U5067 ( .A(n4651), .Y(n9134) );
  AOI21X1_HVT U5068 ( .A1(n57), .A2(n4792), .A3(n10381), .Y(n55) );
  IBUFFX16_HVT U5069 ( .A(n5802), .Y(n4792) );
  INVX0_HVT U5070 ( .A(n4803), .Y(n4793) );
  INVX0_HVT U5071 ( .A(n7578), .Y(n4803) );
  MUX41X1_HVT U5072 ( .A1(\ram[13][18] ), .A3(\ram[15][18] ), .A2(
        \ram[12][18] ), .A4(\ram[14][18] ), .S0(n5523), .S1(n5300), .Y(n7806)
         );
  MUX41X1_HVT U5073 ( .A1(\ram[2][192] ), .A3(\ram[0][192] ), .A2(
        \ram[3][192] ), .A4(\ram[1][192] ), .S0(n5113), .S1(n5593), .Y(n8500)
         );
  INVX0_HVT U5074 ( .A(n7324), .Y(n5125) );
  INVX0_HVT U5075 ( .A(n5487), .Y(n5593) );
  INVX0_HVT U5076 ( .A(n8787), .Y(n4794) );
  INVX0_HVT U5077 ( .A(n4371), .Y(n10128) );
  NBUFFX2_HVT U5078 ( .A(n4942), .Y(n4795) );
  INVX0_HVT U5079 ( .A(n9107), .Y(n4796) );
  INVX0_HVT U5080 ( .A(n4796), .Y(n4797) );
  INVX0_HVT U5081 ( .A(n9089), .Y(n4798) );
  INVX0_HVT U5082 ( .A(n4798), .Y(n4799) );
  NBUFFX2_HVT U5083 ( .A(n9093), .Y(n4800) );
  NBUFFX2_HVT U5084 ( .A(n9099), .Y(n4801) );
  MUX41X1_HVT U5085 ( .A1(n4804), .A3(n4805), .A2(n5842), .A4(n4806), .S0(
        n5803), .S1(n4803), .Y(n4802) );
  IBUFFX16_HVT U5086 ( .A(n4802), .Y(n7949) );
  INVX0_HVT U5087 ( .A(n8781), .Y(n5994) );
  INVX0_HVT U5088 ( .A(n8781), .Y(n6741) );
  MUX41X1_HVT U5089 ( .A1(n4809), .A3(n4810), .A2(n4811), .A4(n4812), .S0(
        n5085), .S1(n4808), .Y(n4807) );
  IBUFFX16_HVT U5090 ( .A(n4807), .Y(n8134) );
  MUX41X1_HVT U5091 ( .A1(n7754), .A3(n7756), .A2(n7755), .A4(n7757), .S0(
        n5723), .S1(n5809), .Y(q[5]) );
  INVX0_HVT U5092 ( .A(n4748), .Y(n4813) );
  INVX0_HVT U5093 ( .A(n5459), .Y(n6181) );
  INVX1_HVT U5094 ( .A(n6145), .Y(n5459) );
  MUX41X1_HVT U5095 ( .A1(n4815), .A3(n4816), .A2(n4817), .A4(n4818), .S0(
        n5574), .S1(n5874), .Y(n4814) );
  NBUFFX2_HVT U5096 ( .A(n8896), .Y(n4819) );
  NBUFFX2_HVT U5097 ( .A(n5107), .Y(n4820) );
  OAI22X1_HVT U5098 ( .A1(n4821), .A2(n4822), .A3(n6207), .A4(n9507), .Y(n1152) );
  INVX0_HVT U5099 ( .A(n6150), .Y(n4822) );
  INVX0_HVT U5100 ( .A(n4822), .Y(n4823) );
  NBUFFX2_HVT U5101 ( .A(n4909), .Y(n4824) );
  NBUFFX2_HVT U5102 ( .A(n6969), .Y(n4825) );
  OAI22X1_HVT U5103 ( .A1(n4827), .A2(n4782), .A3(n4935), .A4(n4826), .Y(n3464) );
  IBUFFX16_HVT U5104 ( .A(data[75]), .Y(n4826) );
  NBUFFX2_HVT U5105 ( .A(n6970), .Y(n4828) );
  INVX0_HVT U5106 ( .A(n4774), .Y(n4829) );
  INVX0_HVT U5107 ( .A(n6864), .Y(n4886) );
  INVX0_HVT U5108 ( .A(n6862), .Y(n6864) );
  INVX0_HVT U5109 ( .A(n5155), .Y(n8825) );
  INVX0_HVT U5110 ( .A(n4839), .Y(n4830) );
  INVX0_HVT U5111 ( .A(n9260), .Y(n4839) );
  INVX0_HVT U5112 ( .A(n5145), .Y(n5054) );
  INVX0_HVT U5113 ( .A(n10203), .Y(n9099) );
  NBUFFX2_HVT U5114 ( .A(n7002), .Y(n4831) );
  INVX0_HVT U5115 ( .A(n4854), .Y(n4832) );
  INVX0_HVT U5116 ( .A(n6999), .Y(n4854) );
  NBUFFX2_HVT U5117 ( .A(n7004), .Y(n4833) );
  INVX0_HVT U5118 ( .A(n7308), .Y(n5826) );
  INVX0_HVT U5119 ( .A(n4844), .Y(n4834) );
  INVX0_HVT U5120 ( .A(n7001), .Y(n4844) );
  NBUFFX2_HVT U5121 ( .A(n4572), .Y(n4835) );
  NBUFFX2_HVT U5122 ( .A(n6152), .Y(n4836) );
  NBUFFX2_HVT U5123 ( .A(n5094), .Y(n4837) );
  MUX41X1_HVT U5124 ( .A1(\ram[6][153] ), .A3(\ram[4][153] ), .A2(
        \ram[7][153] ), .A4(\ram[5][153] ), .S0(n5124), .S1(n7555), .Y(n8343)
         );
  INVX0_HVT U5125 ( .A(n6967), .Y(n7006) );
  INVX0_HVT U5126 ( .A(n6967), .Y(n7007) );
  INVX1_HVT U5127 ( .A(n4924), .Y(n8938) );
  INVX0_HVT U5128 ( .A(n4924), .Y(n8939) );
  INVX0_HVT U5129 ( .A(n8780), .Y(n8785) );
  NBUFFX2_HVT U5130 ( .A(n5688), .Y(n4838) );
  OAI22X1_HVT U5131 ( .A1(n4840), .A2(n4670), .A3(n4839), .A4(n9349), .Y(n1355) );
  OAI22X1_HVT U5132 ( .A1(n4842), .A2(n4916), .A3(n5951), .A4(n4841), .Y(n1392) );
  IBUFFX16_HVT U5133 ( .A(n9460), .Y(n4841) );
  OAI22X1_HVT U5134 ( .A1(n4843), .A2(n4670), .A3(n5010), .A4(n9408), .Y(n1375) );
  OAI22X1_HVT U5135 ( .A1(n4846), .A2(n4844), .A3(n4931), .A4(n4845), .Y(n3417) );
  IBUFFX16_HVT U5136 ( .A(n9392), .Y(n4845) );
  INVX0_HVT U5137 ( .A(n5072), .Y(n6986) );
  INVX0_HVT U5138 ( .A(n9287), .Y(n9289) );
  INVX0_HVT U5139 ( .A(n9287), .Y(n9291) );
  INVX0_HVT U5140 ( .A(n4847), .Y(n4848) );
  INVX0_HVT U5141 ( .A(n6166), .Y(n5484) );
  MUX41X1_HVT U5142 ( .A1(n8111), .A3(n8113), .A2(n8110), .A4(n8112), .S0(
        n5343), .S1(n5339), .Y(q[95]) );
  INVX0_HVT U5143 ( .A(n5676), .Y(n4849) );
  INVX0_HVT U5144 ( .A(n4849), .Y(n4850) );
  INVX0_HVT U5145 ( .A(n4920), .Y(n4851) );
  NBUFFX2_HVT U5146 ( .A(n8918), .Y(n4852) );
  NBUFFX2_HVT U5147 ( .A(n8920), .Y(n4853) );
  OAI22X1_HVT U5148 ( .A1(n4856), .A2(n4854), .A3(n4935), .A4(n4855), .Y(n3419) );
  IBUFFX16_HVT U5149 ( .A(n9398), .Y(n4855) );
  INVX0_HVT U5150 ( .A(n4325), .Y(n5702) );
  NBUFFX2_HVT U5151 ( .A(n9092), .Y(n4857) );
  INVX0_HVT U5152 ( .A(n5525), .Y(n4858) );
  INVX0_HVT U5153 ( .A(n5525), .Y(n4859) );
  MUX41X1_HVT U5154 ( .A1(n8192), .A3(n8190), .A2(n8193), .A4(n8191), .S0(
        n5289), .S1(n6396), .Y(q[115]) );
  INVX0_HVT U5155 ( .A(n5760), .Y(n6393) );
  MUX41X1_HVT U5156 ( .A1(n8202), .A3(n8204), .A2(n8203), .A4(n8205), .S0(
        n5015), .S1(n5868), .Y(q[118]) );
  INVX0_HVT U5157 ( .A(n5347), .Y(n4860) );
  INVX0_HVT U5158 ( .A(n4640), .Y(n5694) );
  INVX0_HVT U5159 ( .A(n5618), .Y(n8841) );
  INVX0_HVT U5160 ( .A(n6360), .Y(n4861) );
  INVX0_HVT U5161 ( .A(n4861), .Y(n4862) );
  INVX0_HVT U5162 ( .A(n5618), .Y(n8835) );
  NBUFFX2_HVT U5163 ( .A(n7043), .Y(n4863) );
  OAI22X1_HVT U5164 ( .A1(n4865), .A2(n4867), .A3(n6851), .A4(n4864), .Y(n359)
         );
  IBUFFX16_HVT U5165 ( .A(n9433), .Y(n4864) );
  INVX0_HVT U5166 ( .A(n6851), .Y(n6861) );
  INVX1_HVT U5167 ( .A(n10344), .Y(n6851) );
  OAI22X1_HVT U5168 ( .A1(n4866), .A2(n4867), .A3(n6870), .A4(n9426), .Y(n357)
         );
  INVX0_HVT U5169 ( .A(n6863), .Y(n6865) );
  INVX0_HVT U5170 ( .A(n7039), .Y(n4867) );
  INVX0_HVT U5171 ( .A(n4867), .Y(n4868) );
  NBUFFX2_HVT U5172 ( .A(n4266), .Y(n4869) );
  NBUFFX2_HVT U5173 ( .A(n4264), .Y(n4870) );
  NBUFFX2_HVT U5174 ( .A(n7049), .Y(n4871) );
  MUX41X1_HVT U5175 ( .A1(\ram[15][126] ), .A3(\ram[13][126] ), .A2(
        \ram[14][126] ), .A4(\ram[12][126] ), .S0(n7305), .S1(n4872), .Y(n8234) );
  INVX0_HVT U5176 ( .A(n5939), .Y(n4872) );
  INVX1_HVT U5177 ( .A(n4872), .Y(n4873) );
  INVX0_HVT U5178 ( .A(n5983), .Y(n5939) );
  OAI22X1_HVT U5179 ( .A1(n4875), .A2(n4919), .A3(n4874), .A4(n9510), .Y(n1665) );
  MUX41X1_HVT U5180 ( .A1(n8012), .A3(n8010), .A2(n8013), .A4(n8011), .S0(
        n5172), .S1(n5776), .Y(q[70]) );
  INVX0_HVT U5181 ( .A(n6381), .Y(n7332) );
  NBUFFX2_HVT U5182 ( .A(n6019), .Y(n8767) );
  MUX41X1_HVT U5183 ( .A1(\ram[15][14] ), .A3(\ram[13][14] ), .A2(
        \ram[14][14] ), .A4(\ram[12][14] ), .S0(n5814), .S1(n4888), .Y(n7790)
         );
  MUX41X1_HVT U5184 ( .A1(\ram[3][144] ), .A3(\ram[1][144] ), .A2(
        \ram[2][144] ), .A4(n4877), .S0(n5816), .S1(n6390), .Y(n4876) );
  INVX0_HVT U5185 ( .A(n5164), .Y(n7699) );
  INVX0_HVT U5186 ( .A(n10), .Y(n7053) );
  INVX0_HVT U5187 ( .A(n5013), .Y(n10) );
  MUX41X1_HVT U5188 ( .A1(n4880), .A3(n4879), .A2(n4881), .A4(n4882), .S0(
        n8800), .S1(n4921), .Y(n4878) );
  IBUFFX16_HVT U5189 ( .A(n4878), .Y(n7990) );
  MUX41X1_HVT U5190 ( .A1(n7760), .A3(n7758), .A2(n7761), .A4(n7759), .S0(
        n4998), .S1(n6400), .Y(q[6]) );
  INVX0_HVT U5191 ( .A(n4898), .Y(n4883) );
  INVX0_HVT U5192 ( .A(n7324), .Y(n4898) );
  NBUFFX2_HVT U5193 ( .A(n7320), .Y(n4884) );
  INVX0_HVT U5194 ( .A(n4375), .Y(n6970) );
  INVX0_HVT U5195 ( .A(n4899), .Y(n4885) );
  INVX0_HVT U5196 ( .A(n6657), .Y(n4899) );
  OAI22X1_HVT U5197 ( .A1(n4887), .A2(n5481), .A3(n4886), .A4(n9815), .Y(n485)
         );
  INVX0_HVT U5198 ( .A(n5235), .Y(n5236) );
  INVX0_HVT U5199 ( .A(n7026), .Y(n7064) );
  OAI22X1_HVT U5200 ( .A1(n4890), .A2(n5481), .A3(n6837), .A4(n4889), .Y(n437)
         );
  IBUFFX16_HVT U5201 ( .A(n9667), .Y(n4889) );
  OAI22X1_HVT U5202 ( .A1(n4892), .A2(n4851), .A3(n5841), .A4(n4891), .Y(n1599) );
  OAI22X1_HVT U5203 ( .A1(n4895), .A2(n4322), .A3(n4893), .A4(n4894), .Y(n1377) );
  INVX0_HVT U5204 ( .A(n4325), .Y(n4896) );
  INVX0_HVT U5205 ( .A(n4914), .Y(n4897) );
  INVX0_HVT U5206 ( .A(n5972), .Y(n6417) );
  INVX0_HVT U5207 ( .A(n1633), .Y(n5515) );
  INVX0_HVT U5208 ( .A(n6113), .Y(n6748) );
  INVX0_HVT U5209 ( .A(n10378), .Y(n10375) );
  INVX0_HVT U5210 ( .A(n9242), .Y(n9246) );
  INVX0_HVT U5211 ( .A(n9242), .Y(n9245) );
  INVX0_HVT U5212 ( .A(n6392), .Y(n8798) );
  INVX0_HVT U5213 ( .A(n6392), .Y(n7298) );
  MUX41X1_HVT U5214 ( .A1(\ram[14][124] ), .A3(\ram[12][124] ), .A2(
        \ram[15][124] ), .A4(\ram[13][124] ), .S0(n4898), .S1(n4899), .Y(n8226) );
  IBUFFX2_HVT U5215 ( .A(n9271), .Y(n4943) );
  NBUFFX2_HVT U5216 ( .A(n6979), .Y(n4900) );
  NBUFFX2_HVT U5217 ( .A(n6980), .Y(n4901) );
  OA22X1_HVT U5218 ( .A1(n4904), .A2(n7418), .A3(n6781), .A4(n4903), .Y(n4902)
         );
  IBUFFX16_HVT U5219 ( .A(n4902), .Y(n2906) );
  INVX0_HVT U5220 ( .A(n4906), .Y(n4905) );
  INVX0_HVT U5221 ( .A(n8837), .Y(n4906) );
  INVX0_HVT U5222 ( .A(n6656), .Y(n5609) );
  MUX41X1_HVT U5223 ( .A1(\ram[11][94] ), .A3(\ram[9][94] ), .A2(\ram[10][94] ), .A4(\ram[8][94] ), .S0(n4906), .S1(n4911), .Y(n8107) );
  INVX1_HVT U5224 ( .A(n5636), .Y(n4911) );
  INVX1_HVT U5225 ( .A(n5426), .Y(n4907) );
  INVX0_HVT U5226 ( .A(n10129), .Y(n4908) );
  NBUFFX2_HVT U5227 ( .A(n6155), .Y(n4910) );
  INVX0_HVT U5228 ( .A(n4922), .Y(n5636) );
  INVX0_HVT U5229 ( .A(n4988), .Y(n5953) );
  INVX0_HVT U5230 ( .A(n6002), .Y(n4912) );
  INVX0_HVT U5231 ( .A(n4912), .Y(n4913) );
  MUX41X1_HVT U5232 ( .A1(\ram[15][165] ), .A3(\ram[13][165] ), .A2(
        \ram[14][165] ), .A4(\ram[12][165] ), .S0(n5234), .S1(n6732), .Y(n8389) );
  INVX0_HVT U5233 ( .A(n5689), .Y(n4914) );
  INVX0_HVT U5234 ( .A(n4941), .Y(n4915) );
  INVX0_HVT U5235 ( .A(n5688), .Y(n4916) );
  INVX0_HVT U5236 ( .A(n4916), .Y(n4917) );
  MUX41X1_HVT U5237 ( .A1(n8391), .A3(n8389), .A2(n8392), .A4(n8390), .S0(
        n4998), .S1(n4997), .Y(q[165]) );
  IBUFFX4_HVT U5238 ( .A(n5372), .Y(n4998) );
  IBUFFX4_HVT U5239 ( .A(n5980), .Y(n4997) );
  MUX41X1_HVT U5240 ( .A1(\ram[7][171] ), .A3(\ram[5][171] ), .A2(
        \ram[6][171] ), .A4(\ram[4][171] ), .S0(n7305), .S1(n5882), .Y(n8415)
         );
  MUX41X1_HVT U5241 ( .A1(n7820), .A3(n7822), .A2(n7821), .A4(n7823), .S0(
        n5207), .S1(n5832), .Y(q[22]) );
  INVX0_HVT U5242 ( .A(n7545), .Y(n5646) );
  INVX0_HVT U5243 ( .A(n7545), .Y(n8826) );
  INVX0_HVT U5244 ( .A(n5949), .Y(n4919) );
  INVX0_HVT U5245 ( .A(n4919), .Y(n4920) );
  MUX41X1_HVT U5246 ( .A1(\ram[15][187] ), .A3(\ram[13][187] ), .A2(
        \ram[14][187] ), .A4(\ram[12][187] ), .S0(n7583), .S1(n4922), .Y(n8477) );
  INVX0_HVT U5247 ( .A(n4922), .Y(n4921) );
  INVX0_HVT U5248 ( .A(n8895), .Y(n6656) );
  INVX0_HVT U5249 ( .A(n8895), .Y(n7290) );
  INVX0_HVT U5250 ( .A(n4926), .Y(n4922) );
  INVX0_HVT U5251 ( .A(n7263), .Y(n5817) );
  INVX0_HVT U5252 ( .A(n7582), .Y(n7151) );
  INVX0_HVT U5253 ( .A(n53), .Y(n4923) );
  INVX0_HVT U5254 ( .A(n4923), .Y(n4924) );
  NBUFFX2_HVT U5255 ( .A(n8953), .Y(n4925) );
  INVX0_HVT U5256 ( .A(n4929), .Y(n4926) );
  NBUFFX2_HVT U5257 ( .A(n4697), .Y(n4927) );
  NBUFFX2_HVT U5258 ( .A(n4697), .Y(n4928) );
  INVX1_HVT U5259 ( .A(n8876), .Y(n5719) );
  INVX0_HVT U5260 ( .A(n8849), .Y(n5979) );
  INVX0_HVT U5261 ( .A(n8849), .Y(n5742) );
  INVX0_HVT U5262 ( .A(n5525), .Y(n10275) );
  INVX0_HVT U5263 ( .A(n5525), .Y(n10277) );
  INVX1_HVT U5264 ( .A(n7268), .Y(n5525) );
  INVX0_HVT U5265 ( .A(n5573), .Y(n5767) );
  NBUFFX2_HVT U5266 ( .A(n6662), .Y(n8889) );
  MUX41X1_HVT U5267 ( .A1(\ram[2][102] ), .A3(\ram[0][102] ), .A2(
        \ram[3][102] ), .A4(\ram[1][102] ), .S0(n5821), .S1(n8889), .Y(n8141)
         );
  INVX0_HVT U5268 ( .A(n7291), .Y(n8832) );
  IBUFFX2_HVT U5269 ( .A(n5626), .Y(n6118) );
  MUX41X1_HVT U5270 ( .A1(\ram[5][235] ), .A3(\ram[7][235] ), .A2(
        \ram[4][235] ), .A4(\ram[6][235] ), .S0(n8808), .S1(n5882), .Y(n8669)
         );
  INVX0_HVT U5271 ( .A(n6408), .Y(n7664) );
  INVX0_HVT U5272 ( .A(n6001), .Y(n4929) );
  INVX0_HVT U5273 ( .A(n4929), .Y(n4930) );
  MUX41X1_HVT U5274 ( .A1(\ram[2][69] ), .A3(\ram[0][69] ), .A2(\ram[3][69] ), 
        .A4(\ram[1][69] ), .S0(n5824), .S1(n5589), .Y(n8009) );
  MUX41X1_HVT U5275 ( .A1(\ram[6][3] ), .A3(\ram[4][3] ), .A2(\ram[7][3] ), 
        .A4(\ram[5][3] ), .S0(n5942), .S1(n5444), .Y(n7748) );
  INVX0_HVT U5276 ( .A(n7545), .Y(n6008) );
  INVX0_HVT U5277 ( .A(n8951), .Y(n4931) );
  INVX0_HVT U5278 ( .A(n4787), .Y(n4932) );
  INVX0_HVT U5279 ( .A(n8951), .Y(n4933) );
  INVX0_HVT U5280 ( .A(n4787), .Y(n4934) );
  INVX0_HVT U5281 ( .A(n8951), .Y(n4935) );
  INVX0_HVT U5282 ( .A(n4933), .Y(n4936) );
  MUX41X1_HVT U5283 ( .A1(\ram[2][11] ), .A3(\ram[0][11] ), .A2(\ram[3][11] ), 
        .A4(\ram[1][11] ), .S0(n5201), .S1(n5287), .Y(n7781) );
  INVX0_HVT U5284 ( .A(n5114), .Y(n5945) );
  NBUFFX2_HVT U5285 ( .A(n5662), .Y(n4937) );
  NBUFFX2_HVT U5286 ( .A(n5708), .Y(n4938) );
  INVX0_HVT U5287 ( .A(n5663), .Y(n5699) );
  INVX0_HVT U5288 ( .A(n4958), .Y(n4939) );
  INVX0_HVT U5289 ( .A(n6410), .Y(n4958) );
  NBUFFX2_HVT U5290 ( .A(n5621), .Y(n4940) );
  INVX1_HVT U5291 ( .A(n22), .Y(n10306) );
  INVX0_HVT U5292 ( .A(n5668), .Y(n4941) );
  INVX0_HVT U5293 ( .A(n4941), .Y(n4942) );
  INVX0_HVT U5294 ( .A(n6656), .Y(n5614) );
  INVX0_HVT U5295 ( .A(n5699), .Y(n5690) );
  INVX0_HVT U5296 ( .A(n4948), .Y(n5708) );
  INVX1_HVT U5297 ( .A(n4947), .Y(n4948) );
  INVX0_HVT U5298 ( .A(n4649), .Y(n5691) );
  INVX0_HVT U5299 ( .A(n4640), .Y(n5695) );
  OAI22X1_HVT U5300 ( .A1(n4944), .A2(n5665), .A3(n4943), .A4(n9492), .Y(n1403) );
  OAI22X1_HVT U5301 ( .A1(n4946), .A2(n4731), .A3(n5782), .A4(n4945), .Y(n1369) );
  IBUFFX16_HVT U5302 ( .A(n9391), .Y(n4945) );
  INVX0_HVT U5303 ( .A(n9288), .Y(n9295) );
  OR2X1_HVT U5304 ( .A1(n10381), .A2(n5051), .Y(n5771) );
  INVX0_HVT U5305 ( .A(n5771), .Y(n4947) );
  NBUFFX2_HVT U5306 ( .A(n7287), .Y(n4949) );
  INVX0_HVT U5307 ( .A(n7287), .Y(n7297) );
  OAI22X1_HVT U5308 ( .A1(n4951), .A2(n4953), .A3(n5951), .A4(n4950), .Y(n1347) );
  IBUFFX16_HVT U5309 ( .A(n9325), .Y(n4950) );
  INVX0_HVT U5310 ( .A(n4941), .Y(n4952) );
  INVX0_HVT U5311 ( .A(n5711), .Y(n4953) );
  INVX0_HVT U5312 ( .A(n4916), .Y(n4954) );
  INVX0_HVT U5313 ( .A(n7350), .Y(n6028) );
  INVX0_HVT U5314 ( .A(n55), .Y(n4955) );
  INVX0_HVT U5315 ( .A(n4955), .Y(n4956) );
  INVX0_HVT U5316 ( .A(n7245), .Y(n7252) );
  INVX0_HVT U5317 ( .A(n7245), .Y(n7250) );
  INVX0_HVT U5318 ( .A(n7244), .Y(n7249) );
  INVX0_HVT U5319 ( .A(n7244), .Y(n7247) );
  INVX0_HVT U5320 ( .A(n7244), .Y(n7246) );
  MUX41X1_HVT U5321 ( .A1(n7853), .A3(n5977), .A2(n7854), .A4(n7852), .S0(
        n7543), .S1(n4999), .Y(q[30]) );
  IBUFFX4_HVT U5322 ( .A(n7352), .Y(n4999) );
  AND2X1_HVT U5323 ( .A1(n5217), .A2(n5218), .Y(n4957) );
  MUX41X1_HVT U5324 ( .A1(\ram[3][194] ), .A3(\ram[1][194] ), .A2(
        \ram[2][194] ), .A4(\ram[0][194] ), .S0(n4958), .S1(n5002), .Y(n8508)
         );
  INVX1_HVT U5325 ( .A(n7695), .Y(n5002) );
  NBUFFX2_HVT U5326 ( .A(n6032), .Y(n8873) );
  OAI22X1_HVT U5327 ( .A1(n4960), .A2(n4964), .A3(n6210), .A4(n4959), .Y(n1133) );
  IBUFFX16_HVT U5328 ( .A(n9451), .Y(n4959) );
  INVX0_HVT U5329 ( .A(n6210), .Y(n6212) );
  INVX0_HVT U5330 ( .A(n4964), .Y(n4961) );
  MUX41X1_HVT U5331 ( .A1(n8273), .A3(n8272), .A2(n8271), .A4(n8270), .S0(
        n5295), .S1(n5003), .Y(q[135]) );
  INVX2_HVT U5332 ( .A(n5898), .Y(n5295) );
  MUX41X1_HVT U5333 ( .A1(\ram[3][196] ), .A3(\ram[1][196] ), .A2(
        \ram[2][196] ), .A4(\ram[0][196] ), .S0(n5942), .S1(n5145), .Y(n8516)
         );
  INVX0_HVT U5334 ( .A(n5953), .Y(n5145) );
  OAI22X1_HVT U5335 ( .A1(n4963), .A2(n5664), .A3(n5951), .A4(n4962), .Y(n1371) );
  IBUFFX16_HVT U5336 ( .A(n9397), .Y(n4962) );
  INVX0_HVT U5337 ( .A(n9288), .Y(n9293) );
  INVX0_HVT U5338 ( .A(n4777), .Y(n4964) );
  INVX0_HVT U5339 ( .A(n4964), .Y(n4965) );
  OAI22X1_HVT U5340 ( .A1(n4967), .A2(n4969), .A3(n4966), .A4(n9423), .Y(n1124) );
  INVX0_HVT U5341 ( .A(n4969), .Y(n4968) );
  INVX0_HVT U5342 ( .A(n5489), .Y(n4969) );
  INVX0_HVT U5343 ( .A(n4969), .Y(n4970) );
  NBUFFX2_HVT U5344 ( .A(n6036), .Y(n4971) );
  INVX0_HVT U5345 ( .A(n5544), .Y(n4972) );
  INVX0_HVT U5346 ( .A(n7673), .Y(n4973) );
  INVX0_HVT U5347 ( .A(n4977), .Y(n4974) );
  INVX0_HVT U5348 ( .A(n7583), .Y(n4975) );
  INVX0_HVT U5349 ( .A(n7670), .Y(n5576) );
  INVX0_HVT U5350 ( .A(n7670), .Y(n5883) );
  INVX0_HVT U5351 ( .A(n6663), .Y(n5053) );
  INVX0_HVT U5352 ( .A(n7678), .Y(n6662) );
  MUX41X1_HVT U5353 ( .A1(\ram[10][153] ), .A3(\ram[8][153] ), .A2(
        \ram[11][153] ), .A4(\ram[9][153] ), .S0(n5527), .S1(n4994), .Y(n8342)
         );
  INVX0_HVT U5354 ( .A(n5608), .Y(n8843) );
  INVX0_HVT U5355 ( .A(n5608), .Y(n8820) );
  INVX0_HVT U5356 ( .A(n6119), .Y(n5949) );
  INVX0_HVT U5357 ( .A(n4978), .Y(n4976) );
  INVX0_HVT U5358 ( .A(n7328), .Y(n4977) );
  NBUFFX2_HVT U5359 ( .A(n8882), .Y(n7328) );
  INVX0_HVT U5360 ( .A(n7663), .Y(n4978) );
  INVX0_HVT U5361 ( .A(n4978), .Y(n4979) );
  INVX0_HVT U5362 ( .A(n5552), .Y(n5650) );
  INVX0_HVT U5363 ( .A(n5961), .Y(n4980) );
  INVX0_HVT U5364 ( .A(n5356), .Y(n4981) );
  INVX0_HVT U5365 ( .A(n5961), .Y(n7336) );
  INVX0_HVT U5366 ( .A(n7582), .Y(n5008) );
  INVX0_HVT U5367 ( .A(n5961), .Y(n5360) );
  INVX0_HVT U5368 ( .A(n8782), .Y(n5322) );
  MUX41X1_HVT U5369 ( .A1(\ram[6][252] ), .A3(\ram[4][252] ), .A2(
        \ram[7][252] ), .A4(\ram[5][252] ), .S0(n6746), .S1(n5656), .Y(n8737)
         );
  MUX41X1_HVT U5370 ( .A1(\ram[12][91] ), .A3(\ram[14][91] ), .A2(
        \ram[13][91] ), .A4(\ram[15][91] ), .S0(n8799), .S1(n5506), .Y(n8094)
         );
  MUX41X1_HVT U5371 ( .A1(\ram[11][171] ), .A3(\ram[9][171] ), .A2(
        \ram[10][171] ), .A4(\ram[8][171] ), .S0(n4986), .S1(n7698), .Y(n8414)
         );
  INVX0_HVT U5372 ( .A(n4948), .Y(n5662) );
  INVX0_HVT U5373 ( .A(n5059), .Y(n8795) );
  INVX0_HVT U5374 ( .A(n5059), .Y(n7549) );
  INVX0_HVT U5375 ( .A(n5059), .Y(n6757) );
  NBUFFX2_HVT U5376 ( .A(n8871), .Y(n8866) );
  INVX0_HVT U5377 ( .A(n7308), .Y(n6732) );
  INVX0_HVT U5378 ( .A(n4913), .Y(n5996) );
  NBUFFX2_HVT U5379 ( .A(n6038), .Y(n8868) );
  INVX0_HVT U5380 ( .A(n5345), .Y(n5331) );
  INVX0_HVT U5381 ( .A(n7684), .Y(n5958) );
  INVX0_HVT U5382 ( .A(n7684), .Y(n7716) );
  INVX0_HVT U5383 ( .A(n7684), .Y(n7709) );
  NBUFFX2_HVT U5384 ( .A(n5615), .Y(n4983) );
  MUX41X1_HVT U5385 ( .A1(n8461), .A3(n8463), .A2(n8462), .A4(n8464), .S0(
        n5015), .S1(n5039), .Y(q[183]) );
  INVX0_HVT U5386 ( .A(n5617), .Y(n8781) );
  INVX0_HVT U5387 ( .A(n5617), .Y(n5618) );
  INVX0_HVT U5388 ( .A(n6038), .Y(n7315) );
  INVX0_HVT U5389 ( .A(n6184), .Y(n6185) );
  INVX0_HVT U5390 ( .A(n8809), .Y(n6645) );
  INVX0_HVT U5391 ( .A(n8809), .Y(n5829) );
  MUX41X1_HVT U5392 ( .A1(\ram[3][185] ), .A3(\ram[1][185] ), .A2(
        \ram[2][185] ), .A4(\ram[0][185] ), .S0(n4986), .S1(n5836), .Y(n8472)
         );
  NBUFFX2_HVT U5393 ( .A(n6115), .Y(n4984) );
  INVX0_HVT U5394 ( .A(n6138), .Y(n6115) );
  INVX0_HVT U5395 ( .A(n7263), .Y(n6626) );
  INVX0_HVT U5396 ( .A(n4986), .Y(n4985) );
  INVX0_HVT U5397 ( .A(n8807), .Y(n4986) );
  MUX41X1_HVT U5398 ( .A1(\ram[6][227] ), .A3(\ram[4][227] ), .A2(
        \ram[7][227] ), .A4(\ram[5][227] ), .S0(n5942), .S1(n6411), .Y(n8639)
         );
  INVX0_HVT U5399 ( .A(n7703), .Y(n4987) );
  INVX0_HVT U5400 ( .A(n7703), .Y(n7698) );
  INVX0_HVT U5401 ( .A(n5632), .Y(n5895) );
  INVX1_HVT U5402 ( .A(n7703), .Y(n6745) );
  INVX0_HVT U5403 ( .A(n5984), .Y(n8805) );
  INVX0_HVT U5404 ( .A(n4192), .Y(n4988) );
  INVX0_HVT U5405 ( .A(n5346), .Y(n5314) );
  INVX0_HVT U5406 ( .A(n7263), .Y(n7265) );
  NBUFFX2_HVT U5407 ( .A(n6626), .Y(n4989) );
  NBUFFX2_HVT U5408 ( .A(n6653), .Y(n4990) );
  INVX0_HVT U5409 ( .A(n5651), .Y(n6653) );
  INVX0_HVT U5410 ( .A(n5798), .Y(n4991) );
  NBUFFX2_HVT U5411 ( .A(n7559), .Y(n4992) );
  MUX41X1_HVT U5412 ( .A1(\ram[14][129] ), .A3(\ram[12][129] ), .A2(
        \ram[15][129] ), .A4(\ram[13][129] ), .S0(n7314), .S1(n5907), .Y(n8246) );
  NBUFFX2_HVT U5413 ( .A(n6626), .Y(n4993) );
  INVX0_HVT U5414 ( .A(n7295), .Y(n6646) );
  MUX41X1_HVT U5415 ( .A1(\ram[7][212] ), .A3(\ram[5][212] ), .A2(
        \ram[6][212] ), .A4(\ram[4][212] ), .S0(n5555), .S1(n5002), .Y(n8579)
         );
  NBUFFX2_HVT U5416 ( .A(n4188), .Y(n8861) );
  MUX41X1_HVT U5417 ( .A1(n7857), .A3(n7855), .A2(n7858), .A4(n7856), .S0(
        n5003), .S1(n5887), .Y(q[31]) );
  IBUFFX4_HVT U5418 ( .A(n5326), .Y(n5003) );
  INVX0_HVT U5419 ( .A(n7144), .Y(n7712) );
  NBUFFX2_HVT U5420 ( .A(n5943), .Y(n4994) );
  INVX0_HVT U5421 ( .A(n5988), .Y(n5943) );
  INVX0_HVT U5422 ( .A(n7343), .Y(n7319) );
  NBUFFX2_HVT U5423 ( .A(n6743), .Y(n4995) );
  MUX41X1_HVT U5424 ( .A1(n8641), .A3(n8643), .A2(n8642), .A4(n8644), .S0(
        n4996), .S1(n4997), .Y(q[228]) );
  IBUFFX16_HVT U5425 ( .A(n5867), .Y(n4996) );
  INVX1_HVT U5426 ( .A(n7311), .Y(n6413) );
  INVX0_HVT U5427 ( .A(n5366), .Y(n5001) );
  NBUFFX2_HVT U5428 ( .A(n6114), .Y(n5366) );
  NBUFFX2_HVT U5429 ( .A(n6185), .Y(n7695) );
  MUX41X1_HVT U5430 ( .A1(n8416), .A3(n8414), .A2(n8415), .A4(n8413), .S0(
        n5003), .S1(n5746), .Y(q[171]) );
  INVX0_HVT U5431 ( .A(n4926), .Y(n5568) );
  NBUFFX2_HVT U5432 ( .A(n8807), .Y(n5004) );
  INVX1_HVT U5433 ( .A(n6126), .Y(n5729) );
  IBUFFX2_HVT U5434 ( .A(n7301), .Y(n5018) );
  INVX0_HVT U5435 ( .A(n5370), .Y(n5005) );
  INVX0_HVT U5436 ( .A(n5005), .Y(n5006) );
  INVX0_HVT U5437 ( .A(n5153), .Y(n5370) );
  MUX41X1_HVT U5438 ( .A1(n8646), .A3(n8648), .A2(n8645), .A4(n8647), .S0(
        n7548), .S1(n5007), .Y(q[229]) );
  INVX0_HVT U5439 ( .A(n4639), .Y(n5009) );
  INVX0_HVT U5440 ( .A(n4410), .Y(n5010) );
  INVX0_HVT U5441 ( .A(n5010), .Y(n5011) );
  INVX0_HVT U5442 ( .A(n7582), .Y(n7565) );
  INVX0_HVT U5443 ( .A(n7147), .Y(n5014) );
  IBUFFX2_HVT U5444 ( .A(n6032), .Y(n5919) );
  MUX41X1_HVT U5445 ( .A1(n8387), .A3(n8385), .A2(n8388), .A4(n8386), .S0(
        n5172), .S1(n5012), .Y(q[164]) );
  IBUFFX2_HVT U5446 ( .A(n7297), .Y(n8844) );
  AO21X1_HVT U5447 ( .A1(n12), .A2(we), .A3(rst), .Y(n5013) );
  INVX0_HVT U5448 ( .A(n9287), .Y(n9290) );
  MUX41X1_HVT U5449 ( .A1(\ram[8][249] ), .A3(\ram[10][249] ), .A2(
        \ram[9][249] ), .A4(\ram[11][249] ), .S0(n5014), .S1(n5143), .Y(n8724)
         );
  MUX41X1_HVT U5450 ( .A1(n8082), .A3(n8084), .A2(n8083), .A4(n8085), .S0(
        n5015), .S1(n5016), .Y(q[88]) );
  MUX41X1_HVT U5451 ( .A1(n7928), .A3(n7930), .A2(n7927), .A4(n7929), .S0(
        n5017), .S1(n5018), .Y(q[49]) );
  IBUFFX16_HVT U5452 ( .A(n5171), .Y(n5017) );
  MUX41X1_HVT U5453 ( .A1(n8529), .A3(n8531), .A2(n8530), .A4(n8532), .S0(
        n5019), .S1(n5020), .Y(q[200]) );
  IBUFFX16_HVT U5454 ( .A(n5799), .Y(n5019) );
  NAND2X0_HVT U5455 ( .A1(\ram[1][18] ), .A2(n7069), .Y(n5021) );
  NAND2X0_HVT U5456 ( .A1(n6877), .A2(n9362), .Y(n5022) );
  NAND2X0_HVT U5457 ( .A1(n5021), .A2(n5022), .Y(n335) );
  INVX0_HVT U5458 ( .A(n6875), .Y(n6877) );
  INVX0_HVT U5459 ( .A(n5084), .Y(n5055) );
  NBUFFX2_HVT U5460 ( .A(n6117), .Y(n8895) );
  NBUFFX2_HVT U5461 ( .A(n6022), .Y(n8878) );
  NAND2X0_HVT U5462 ( .A1(n5769), .A2(n5055), .Y(n5056) );
  INVX0_HVT U5463 ( .A(n10315), .Y(n10314) );
  INVX1_HVT U5464 ( .A(n10381), .Y(n5218) );
  INVX1_HVT U5465 ( .A(n5835), .Y(n10381) );
  NBUFFX2_HVT U5466 ( .A(n6022), .Y(n7580) );
  INVX0_HVT U5467 ( .A(n6656), .Y(n5758) );
  NBUFFX2_HVT U5468 ( .A(n7718), .Y(n7577) );
  INVX0_HVT U5469 ( .A(n8833), .Y(n7311) );
  INVX1_HVT U5470 ( .A(n6759), .Y(n7294) );
  IBUFFX2_HVT U5471 ( .A(n6135), .Y(n5080) );
  INVX1_HVT U5472 ( .A(n6022), .Y(n5732) );
  NBUFFX2_HVT U5473 ( .A(n6662), .Y(n8857) );
  IBUFFX2_HVT U5474 ( .A(n5983), .Y(n5143) );
  INVX0_HVT U5475 ( .A(n6252), .Y(n5974) );
  INVX0_HVT U5476 ( .A(n6750), .Y(n8756) );
  INVX0_HVT U5477 ( .A(n4327), .Y(n10345) );
  INVX0_HVT U5478 ( .A(n4778), .Y(n6152) );
  INVX0_HVT U5479 ( .A(n7725), .Y(n6186) );
  INVX0_HVT U5480 ( .A(n5170), .Y(n5668) );
  INVX0_HVT U5481 ( .A(n10221), .Y(n10218) );
  INVX0_HVT U5482 ( .A(n52), .Y(n6997) );
  INVX1_HVT U5483 ( .A(n8769), .Y(n5902) );
  NBUFFX2_HVT U5484 ( .A(n5853), .Y(n8902) );
  INVX0_HVT U5485 ( .A(n8763), .Y(n8753) );
  INVX0_HVT U5486 ( .A(n5734), .Y(n5335) );
  INVX0_HVT U5487 ( .A(n8800), .Y(n5426) );
  INVX0_HVT U5488 ( .A(n5972), .Y(n6747) );
  NBUFFX2_HVT U5489 ( .A(n5447), .Y(n8854) );
  INVX0_HVT U5490 ( .A(n8775), .Y(n5102) );
  INVX0_HVT U5491 ( .A(n8754), .Y(n8759) );
  INVX0_HVT U5492 ( .A(n6894), .Y(n5770) );
  NBUFFX2_HVT U5493 ( .A(n5641), .Y(n7701) );
  INVX0_HVT U5494 ( .A(n8754), .Y(n8760) );
  NBUFFX2_HVT U5495 ( .A(n6022), .Y(n8886) );
  NBUFFX2_HVT U5496 ( .A(n6892), .Y(n8908) );
  INVX1_HVT U5497 ( .A(n5721), .Y(n5926) );
  INVX0_HVT U5498 ( .A(n6113), .Y(n6035) );
  NBUFFX2_HVT U5499 ( .A(n5947), .Y(n8769) );
  INVX0_HVT U5500 ( .A(n5923), .Y(n5234) );
  INVX0_HVT U5501 ( .A(n6406), .Y(n5356) );
  INVX1_HVT U5502 ( .A(n8867), .Y(n7345) );
  MUX41X1_HVT U5503 ( .A1(\ram[15][190] ), .A3(\ram[13][190] ), .A2(
        \ram[14][190] ), .A4(\ram[12][190] ), .S0(n5903), .S1(n7149), .Y(n8489) );
  IBUFFX2_HVT U5504 ( .A(n5312), .Y(n5355) );
  INVX0_HVT U5505 ( .A(n7697), .Y(n5122) );
  INVX0_HVT U5506 ( .A(n6397), .Y(n5340) );
  IBUFFX2_HVT U5507 ( .A(n8756), .Y(n5372) );
  INVX0_HVT U5508 ( .A(n8787), .Y(n6018) );
  NBUFFX2_HVT U5509 ( .A(n5553), .Y(n6385) );
  INVX0_HVT U5510 ( .A(n5543), .Y(n5505) );
  INVX0_HVT U5511 ( .A(n7197), .Y(n5160) );
  INVX0_HVT U5512 ( .A(n6166), .Y(n6171) );
  INVX0_HVT U5513 ( .A(n6159), .Y(n6162) );
  INVX0_HVT U5514 ( .A(n6159), .Y(n6164) );
  NBUFFX2_HVT U5515 ( .A(n10101), .Y(n5384) );
  INVX0_HVT U5516 ( .A(n5904), .Y(n5109) );
  INVX0_HVT U5517 ( .A(n6397), .Y(n5171) );
  OR2X1_HVT U5518 ( .A1(n6273), .A2(n9522), .Y(n5159) );
  INVX0_HVT U5519 ( .A(n7100), .Y(n5374) );
  NAND2X0_HVT U5520 ( .A1(\ram[3][1] ), .A2(n7099), .Y(n5327) );
  INVX0_HVT U5521 ( .A(n7134), .Y(n5349) );
  INVX0_HVT U5522 ( .A(n7127), .Y(n5285) );
  NAND2X0_HVT U5523 ( .A1(\ram[3][203] ), .A2(n7122), .Y(n5643) );
  INVX0_HVT U5524 ( .A(n7099), .Y(n5329) );
  AO22X1_HVT U5525 ( .A1(\ram[4][215] ), .A2(n4836), .A3(n6209), .A4(n9965), 
        .Y(n1300) );
  INVX1_HVT U5526 ( .A(n5116), .Y(n1617) );
  INVX0_HVT U5527 ( .A(n9444), .Y(n9446) );
  INVX0_HVT U5528 ( .A(n9675), .Y(n9677) );
  INVX0_HVT U5529 ( .A(n9318), .Y(n9320) );
  INVX0_HVT U5530 ( .A(data[54]), .Y(n9468) );
  INVX0_HVT U5531 ( .A(n9468), .Y(n9470) );
  INVX0_HVT U5532 ( .A(n9955), .Y(n9957) );
  INVX0_HVT U5533 ( .A(n5183), .Y(n5184) );
  INVX0_HVT U5534 ( .A(n9797), .Y(n9799) );
  INVX0_HVT U5535 ( .A(n7729), .Y(n10140) );
  INVX0_HVT U5536 ( .A(n10140), .Y(n6578) );
  INVX0_HVT U5537 ( .A(n4978), .Y(n7555) );
  INVX0_HVT U5538 ( .A(n9645), .Y(n9647) );
  INVX0_HVT U5539 ( .A(n9672), .Y(n9674) );
  INVX0_HVT U5540 ( .A(n9627), .Y(n9629) );
  INVX0_HVT U5541 ( .A(n9522), .Y(n9524) );
  INVX0_HVT U5542 ( .A(n9525), .Y(n9527) );
  INVX0_HVT U5543 ( .A(n9519), .Y(n9521) );
  INVX0_HVT U5544 ( .A(n9375), .Y(n9377) );
  INVX0_HVT U5545 ( .A(n10073), .Y(n10075) );
  INVX0_HVT U5546 ( .A(n9417), .Y(n9419) );
  INVX0_HVT U5547 ( .A(n9492), .Y(n9494) );
  INVX0_HVT U5548 ( .A(n9474), .Y(n9476) );
  INVX0_HVT U5549 ( .A(n9480), .Y(n9482) );
  INVX0_HVT U5550 ( .A(n9516), .Y(n9518) );
  INVX0_HVT U5551 ( .A(n9794), .Y(n9796) );
  INVX0_HVT U5552 ( .A(n9870), .Y(n9872) );
  INVX0_HVT U5553 ( .A(n10083), .Y(n10085) );
  INVX0_HVT U5554 ( .A(n10045), .Y(n10047) );
  INVX0_HVT U5555 ( .A(data[217]), .Y(n9970) );
  INVX0_HVT U5556 ( .A(n9970), .Y(n9972) );
  INVX0_HVT U5557 ( .A(n9324), .Y(n9326) );
  INVX0_HVT U5558 ( .A(n9534), .Y(n9536) );
  INVX0_HVT U5559 ( .A(n9311), .Y(n9312) );
  INVX0_HVT U5560 ( .A(n9311), .Y(n9313) );
  INVX0_HVT U5561 ( .A(n9399), .Y(n9401) );
  INVX0_HVT U5562 ( .A(n9678), .Y(n9680) );
  INVX0_HVT U5563 ( .A(n9579), .Y(n9581) );
  INVX0_HVT U5564 ( .A(n9471), .Y(n9473) );
  INVX0_HVT U5565 ( .A(n9564), .Y(n9566) );
  INVX0_HVT U5566 ( .A(n9414), .Y(n9416) );
  INVX0_HVT U5567 ( .A(n9720), .Y(n9722) );
  INVX0_HVT U5568 ( .A(n5062), .Y(n6142) );
  INVX0_HVT U5569 ( .A(n6803), .Y(n6805) );
  INVX0_HVT U5570 ( .A(n7719), .Y(n10164) );
  INVX0_HVT U5571 ( .A(n6816), .Y(n6787) );
  INVX0_HVT U5572 ( .A(n6816), .Y(n6811) );
  INVX0_HVT U5573 ( .A(n6292), .Y(n10324) );
  INVX0_HVT U5574 ( .A(n10315), .Y(n10309) );
  INVX0_HVT U5575 ( .A(n5244), .Y(n5252) );
  INVX0_HVT U5576 ( .A(n5301), .Y(n10307) );
  INVX0_HVT U5577 ( .A(n10238), .Y(n7359) );
  INVX0_HVT U5578 ( .A(n6749), .Y(n8757) );
  INVX0_HVT U5579 ( .A(n5321), .Y(n5297) );
  INVX0_HVT U5580 ( .A(n5321), .Y(n5305) );
  INVX0_HVT U5581 ( .A(n5305), .Y(n6259) );
  INVX0_HVT U5582 ( .A(n5625), .Y(n5131) );
  INVX0_HVT U5583 ( .A(n6658), .Y(n6651) );
  NBUFFX2_HVT U5584 ( .A(n5819), .Y(n5795) );
  INVX0_HVT U5585 ( .A(n7323), .Y(n5309) );
  INVX1_HVT U5586 ( .A(n5795), .Y(n5161) );
  INVX0_HVT U5587 ( .A(n5987), .Y(n5988) );
  INVX0_HVT U5588 ( .A(n8876), .Y(n6252) );
  INVX0_HVT U5589 ( .A(n8906), .Y(n7289) );
  NBUFFX2_HVT U5590 ( .A(n5862), .Y(n7578) );
  INVX0_HVT U5591 ( .A(n5853), .Y(n5588) );
  INVX0_HVT U5592 ( .A(n6891), .Y(n6135) );
  INVX0_HVT U5593 ( .A(n5827), .Y(n5039) );
  INVX1_HVT U5594 ( .A(n7573), .Y(n5581) );
  INVX0_HVT U5595 ( .A(n5877), .Y(n5873) );
  INVX0_HVT U5596 ( .A(n5199), .Y(n5092) );
  INVX1_HVT U5597 ( .A(n5995), .Y(n5339) );
  INVX1_HVT U5598 ( .A(n8778), .Y(n5871) );
  INVX0_HVT U5599 ( .A(n5093), .Y(n5308) );
  INVX1_HVT U5600 ( .A(n5873), .Y(n5157) );
  INVX0_HVT U5601 ( .A(n5827), .Y(n5199) );
  INVX0_HVT U5602 ( .A(n9952), .Y(n9954) );
  INVX0_HVT U5603 ( .A(n10051), .Y(n10053) );
  INVX0_HVT U5604 ( .A(n9876), .Y(n9878) );
  INVX0_HVT U5605 ( .A(n9711), .Y(n9713) );
  INVX0_HVT U5606 ( .A(n9815), .Y(n9817) );
  INVX0_HVT U5607 ( .A(n9943), .Y(n9945) );
  INVX0_HVT U5608 ( .A(n9690), .Y(n9692) );
  INVX0_HVT U5609 ( .A(n9828), .Y(n9830) );
  INVX0_HVT U5610 ( .A(n9992), .Y(n9994) );
  INVX0_HVT U5611 ( .A(n9964), .Y(n9966) );
  INVX0_HVT U5612 ( .A(n9702), .Y(n9704) );
  INVX0_HVT U5613 ( .A(n10029), .Y(n10031) );
  INVX0_HVT U5614 ( .A(n9727), .Y(n9729) );
  INVX0_HVT U5615 ( .A(n9841), .Y(n9843) );
  INVX0_HVT U5616 ( .A(n9791), .Y(n9793) );
  INVX0_HVT U5617 ( .A(n9905), .Y(n9907) );
  INVX0_HVT U5618 ( .A(n9918), .Y(n9920) );
  INVX0_HVT U5619 ( .A(n9867), .Y(n9869) );
  INVX0_HVT U5620 ( .A(n9967), .Y(n9969) );
  INVX0_HVT U5621 ( .A(n9980), .Y(n9982) );
  INVX0_HVT U5622 ( .A(n10017), .Y(n10019) );
  INVX0_HVT U5623 ( .A(n9762), .Y(n9764) );
  INVX0_HVT U5624 ( .A(n10004), .Y(n10006) );
  INVX0_HVT U5625 ( .A(n9778), .Y(n9780) );
  INVX0_HVT U5626 ( .A(n10067), .Y(n10069) );
  INVX0_HVT U5627 ( .A(n9892), .Y(n9894) );
  INVX0_HVT U5628 ( .A(n9803), .Y(n9805) );
  INVX0_HVT U5629 ( .A(n10054), .Y(n10056) );
  INVX0_HVT U5630 ( .A(n9879), .Y(n9881) );
  INVX0_HVT U5631 ( .A(data[252]), .Y(n10080) );
  INVX0_HVT U5632 ( .A(n10080), .Y(n10082) );
  INVX0_HVT U5633 ( .A(n9714), .Y(n9716) );
  INVX0_HVT U5634 ( .A(n9753), .Y(n9755) );
  INVX0_HVT U5635 ( .A(n9740), .Y(n9742) );
  INVX0_HVT U5636 ( .A(n10042), .Y(n10044) );
  INVX0_HVT U5637 ( .A(n9812), .Y(n9814) );
  INVX0_HVT U5638 ( .A(n9927), .Y(n9929) );
  INVX0_HVT U5639 ( .A(n9927), .Y(n9928) );
  INVX0_HVT U5640 ( .A(n9765), .Y(n9767) );
  INVX0_HVT U5641 ( .A(n9930), .Y(n9932) );
  INVX0_HVT U5642 ( .A(data[204]), .Y(n9930) );
  INVX0_HVT U5643 ( .A(n9699), .Y(n9701) );
  INVX0_HVT U5644 ( .A(n10001), .Y(n10003) );
  INVX0_HVT U5645 ( .A(n9989), .Y(n9991) );
  INVX0_HVT U5646 ( .A(n10026), .Y(n10028) );
  INVX0_HVT U5647 ( .A(n9800), .Y(n9802) );
  INVX0_HVT U5648 ( .A(n9280), .Y(n9258) );
  INVX0_HVT U5649 ( .A(n9995), .Y(n9997) );
  OAI22X1_HVT U5650 ( .A1(n5526), .A2(n4279), .A3(n5117), .A4(n9921), .Y(n5023) );
  INVX0_HVT U5651 ( .A(n9873), .Y(n9875) );
  INVX0_HVT U5652 ( .A(n10048), .Y(n10050) );
  OAI22X1_HVT U5653 ( .A1(n5897), .A2(n5380), .A3(n6015), .A4(n9930), .Y(n5024) );
  OAI22X1_HVT U5654 ( .A1(n6011), .A2(n5173), .A3(n5117), .A4(n9414), .Y(n5025) );
  OAI22X1_HVT U5655 ( .A1(n5532), .A2(n4971), .A3(n5846), .A4(n9305), .Y(n5026) );
  AO22X1_HVT U5656 ( .A1(\ram[4][59] ), .A2(n6162), .A3(n6234), .A4(n9484), 
        .Y(n5027) );
  AO22X1_HVT U5657 ( .A1(\ram[4][52] ), .A2(n6163), .A3(n6241), .A4(n9463), 
        .Y(n5028) );
  OAI22X1_HVT U5658 ( .A1(n5330), .A2(n5329), .A3(n5284), .A4(n10070), .Y(
        n5029) );
  OAI22X1_HVT U5659 ( .A1(n5350), .A2(n5349), .A3(n5253), .A4(n9417), .Y(n5030) );
  OAI22X1_HVT U5660 ( .A1(n6256), .A2(n6255), .A3(n5284), .A4(n9318), .Y(n5031) );
  OAI22X1_HVT U5661 ( .A1(n5375), .A2(n5374), .A3(n5284), .A4(n9305), .Y(n5032) );
  OAI22X1_HVT U5662 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n9570), .Y(n5034) );
  INVX0_HVT U5663 ( .A(n9687), .Y(n9689) );
  INVX0_HVT U5664 ( .A(n9633), .Y(n9635) );
  INVX0_HVT U5665 ( .A(n9946), .Y(n9948) );
  INVX0_HVT U5666 ( .A(n10057), .Y(n10059) );
  INVX0_HVT U5667 ( .A(n9447), .Y(n9449) );
  INVX0_HVT U5668 ( .A(n9594), .Y(n9596) );
  INVX0_HVT U5669 ( .A(n9540), .Y(n9542) );
  INVX0_HVT U5670 ( .A(n9537), .Y(n9539) );
  INVX0_HVT U5671 ( .A(n9908), .Y(n9910) );
  INVX0_HVT U5672 ( .A(n9857), .Y(n9859) );
  INVX0_HVT U5673 ( .A(n9717), .Y(n9719) );
  INVX0_HVT U5674 ( .A(n9669), .Y(n9671) );
  INVX0_HVT U5675 ( .A(n9549), .Y(n9551) );
  INVX0_HVT U5676 ( .A(n9844), .Y(n9846) );
  INVX0_HVT U5677 ( .A(n9743), .Y(n9745) );
  INVX0_HVT U5678 ( .A(n10007), .Y(n10009) );
  INVX0_HVT U5679 ( .A(n9818), .Y(n9820) );
  INVX0_HVT U5680 ( .A(n9983), .Y(n9985) );
  INVX0_HVT U5681 ( .A(n9895), .Y(n9897) );
  INVX0_HVT U5682 ( .A(n9756), .Y(n9758) );
  INVX0_HVT U5683 ( .A(n9882), .Y(n9884) );
  INVX0_HVT U5684 ( .A(n9507), .Y(n9509) );
  INVX0_HVT U5685 ( .A(n9831), .Y(n9833) );
  INVX0_HVT U5686 ( .A(n10020), .Y(n10022) );
  INVX0_HVT U5687 ( .A(n9693), .Y(n9695) );
  INVX0_HVT U5688 ( .A(n9730), .Y(n9732) );
  INVX0_HVT U5689 ( .A(n9781), .Y(n9783) );
  INVX0_HVT U5690 ( .A(n9806), .Y(n9808) );
  INVX0_HVT U5691 ( .A(n9933), .Y(n9935) );
  INVX0_HVT U5692 ( .A(data[201]), .Y(n9921) );
  INVX0_HVT U5693 ( .A(n9921), .Y(n9923) );
  INVX0_HVT U5694 ( .A(n9681), .Y(n9683) );
  INVX0_HVT U5695 ( .A(n9630), .Y(n9632) );
  INVX0_HVT U5696 ( .A(n9573), .Y(n9575) );
  INVX0_HVT U5697 ( .A(n9498), .Y(n9500) );
  INVX0_HVT U5698 ( .A(n9501), .Y(n9503) );
  INVX0_HVT U5699 ( .A(n9513), .Y(n9515) );
  INVX0_HVT U5700 ( .A(data[213]), .Y(n9958) );
  INVX0_HVT U5701 ( .A(n9958), .Y(n9960) );
  INVX0_HVT U5702 ( .A(n9705), .Y(n9707) );
  OAI22X1_HVT U5703 ( .A1(n6016), .A2(n5380), .A3(n6015), .A4(n9450), .Y(n5035) );
  INVX0_HVT U5704 ( .A(n10032), .Y(n10034) );
  INVX0_HVT U5705 ( .A(n9768), .Y(n9770) );
  INVX0_HVT U5706 ( .A(n9642), .Y(n9644) );
  INVX0_HVT U5707 ( .A(n9308), .Y(n9310) );
  INVX0_HVT U5708 ( .A(n9308), .Y(n9309) );
  INVX0_HVT U5709 ( .A(n9854), .Y(n9856) );
  INVX0_HVT U5710 ( .A(n9588), .Y(n9590) );
  INVX0_HVT U5711 ( .A(n9597), .Y(n9599) );
  INVX0_HVT U5712 ( .A(n9663), .Y(n9665) );
  INVX0_HVT U5713 ( .A(n10070), .Y(n10072) );
  INVX0_HVT U5714 ( .A(n9657), .Y(n9659) );
  INVX0_HVT U5715 ( .A(n9358), .Y(n9360) );
  INVX0_HVT U5716 ( .A(n9528), .Y(n9530) );
  INVX0_HVT U5717 ( .A(n9591), .Y(n9593) );
  INVX0_HVT U5718 ( .A(n9621), .Y(n9623) );
  INVX0_HVT U5719 ( .A(n9651), .Y(n9653) );
  INVX0_HVT U5720 ( .A(data[42]), .Y(n9432) );
  INVX0_HVT U5721 ( .A(n9432), .Y(n9434) );
  INVX0_HVT U5722 ( .A(n9477), .Y(n9479) );
  INVX0_HVT U5723 ( .A(n9495), .Y(n9497) );
  INVX0_HVT U5724 ( .A(n9372), .Y(n9374) );
  INVX0_HVT U5725 ( .A(n9384), .Y(n9386) );
  INVX0_HVT U5726 ( .A(n9336), .Y(n9338) );
  INVX0_HVT U5727 ( .A(n9346), .Y(n9348) );
  INVX0_HVT U5728 ( .A(n9327), .Y(n9329) );
  INVX0_HVT U5729 ( .A(data[5]), .Y(n9321) );
  INVX0_HVT U5730 ( .A(n9321), .Y(n9323) );
  INVX0_HVT U5731 ( .A(n9429), .Y(n9431) );
  INVX0_HVT U5732 ( .A(n9618), .Y(n9620) );
  INVX0_HVT U5733 ( .A(n9504), .Y(n9506) );
  INVX0_HVT U5734 ( .A(n9609), .Y(n9611) );
  INVX0_HVT U5735 ( .A(n9510), .Y(n9512) );
  INVX0_HVT U5736 ( .A(n9585), .Y(n9587) );
  INVX0_HVT U5737 ( .A(n9402), .Y(n9404) );
  INVX0_HVT U5738 ( .A(n9352), .Y(n9354) );
  INVX0_HVT U5739 ( .A(data[9]), .Y(n9333) );
  INVX0_HVT U5740 ( .A(n9333), .Y(n9335) );
  INVX0_HVT U5741 ( .A(data[21]), .Y(n9369) );
  INVX0_HVT U5742 ( .A(n9369), .Y(n9371) );
  INVX0_HVT U5743 ( .A(data[8]), .Y(n9330) );
  INVX0_HVT U5744 ( .A(n9330), .Y(n9332) );
  INVX0_HVT U5745 ( .A(n9364), .Y(n9366) );
  INVX0_HVT U5746 ( .A(n9408), .Y(n9410) );
  INVX0_HVT U5747 ( .A(n9423), .Y(n9425) );
  INVX0_HVT U5748 ( .A(n9654), .Y(n9656) );
  INVX0_HVT U5749 ( .A(n9684), .Y(n9686) );
  INVX0_HVT U5750 ( .A(n9600), .Y(n9602) );
  INVX0_HVT U5751 ( .A(n9636), .Y(n9638) );
  INVX0_HVT U5752 ( .A(n9486), .Y(n9488) );
  INVX0_HVT U5753 ( .A(n9603), .Y(n9605) );
  INVX0_HVT U5754 ( .A(n9561), .Y(n9563) );
  INVX0_HVT U5755 ( .A(n9483), .Y(n9485) );
  INVX0_HVT U5756 ( .A(n9552), .Y(n9554) );
  INVX0_HVT U5757 ( .A(n9405), .Y(n9407) );
  INVX0_HVT U5758 ( .A(n9576), .Y(n9578) );
  INVX0_HVT U5759 ( .A(n9639), .Y(n9641) );
  INVX0_HVT U5760 ( .A(n9624), .Y(n9626) );
  INVX0_HVT U5761 ( .A(n9612), .Y(n9614) );
  INVX0_HVT U5762 ( .A(n9606), .Y(n9608) );
  INVX0_HVT U5763 ( .A(n9582), .Y(n9584) );
  INVX0_HVT U5764 ( .A(n9546), .Y(n9548) );
  INVX0_HVT U5765 ( .A(n9543), .Y(n9545) );
  INVX0_HVT U5766 ( .A(n9462), .Y(n9464) );
  INVX0_HVT U5767 ( .A(n9489), .Y(n9491) );
  INVX0_HVT U5768 ( .A(data[53]), .Y(n9465) );
  INVX0_HVT U5769 ( .A(n9465), .Y(n9467) );
  INVX0_HVT U5770 ( .A(data[51]), .Y(n9459) );
  INVX0_HVT U5771 ( .A(n9459), .Y(n9461) );
  INVX0_HVT U5772 ( .A(n9567), .Y(n9569) );
  INVX0_HVT U5773 ( .A(data[18]), .Y(n9361) );
  INVX0_HVT U5774 ( .A(n9361), .Y(n9363) );
  INVX0_HVT U5775 ( .A(n9558), .Y(n9560) );
  INVX0_HVT U5776 ( .A(n9378), .Y(n9380) );
  INVX0_HVT U5777 ( .A(data[25]), .Y(n9381) );
  INVX0_HVT U5778 ( .A(n9381), .Y(n9383) );
  INVX0_HVT U5779 ( .A(n9435), .Y(n9437) );
  INVX0_HVT U5780 ( .A(n9420), .Y(n9422) );
  INVX0_HVT U5781 ( .A(n9441), .Y(n9443) );
  INVX0_HVT U5782 ( .A(data[29]), .Y(n9393) );
  INVX0_HVT U5783 ( .A(n9393), .Y(n9395) );
  INVX0_HVT U5784 ( .A(n9349), .Y(n9351) );
  INVX0_HVT U5785 ( .A(data[118]), .Y(n9660) );
  INVX0_HVT U5786 ( .A(n9660), .Y(n9662) );
  INVX0_HVT U5787 ( .A(n9648), .Y(n9650) );
  INVX0_HVT U5788 ( .A(n9666), .Y(n9668) );
  INVX0_HVT U5789 ( .A(n9438), .Y(n9440) );
  INVX0_HVT U5790 ( .A(n9426), .Y(n9428) );
  INVX0_HVT U5791 ( .A(n9411), .Y(n9413) );
  INVX0_HVT U5792 ( .A(n9456), .Y(n9458) );
  INVX0_HVT U5793 ( .A(n5183), .Y(n5185) );
  INVX0_HVT U5794 ( .A(n9615), .Y(n9617) );
  INVX0_HVT U5795 ( .A(data[88]), .Y(n9570) );
  INVX0_HVT U5796 ( .A(n9570), .Y(n9572) );
  INVX0_HVT U5797 ( .A(n9555), .Y(n9557) );
  INVX0_HVT U5798 ( .A(n9531), .Y(n9533) );
  INVX0_HVT U5799 ( .A(n9390), .Y(n9392) );
  INVX0_HVT U5800 ( .A(n9450), .Y(n9452) );
  INVX0_HVT U5801 ( .A(data[48]), .Y(n9450) );
  INVX0_HVT U5802 ( .A(n5175), .Y(n5173) );
  INVX0_HVT U5803 ( .A(n5183), .Y(n5187) );
  INVX0_HVT U5804 ( .A(n5183), .Y(n5186) );
  INVX0_HVT U5805 ( .A(n5183), .Y(n5188) );
  INVX0_HVT U5806 ( .A(n9343), .Y(n9345) );
  INVX0_HVT U5807 ( .A(data[16]), .Y(n9355) );
  INVX0_HVT U5808 ( .A(n9355), .Y(n9357) );
  INVX0_HVT U5809 ( .A(data[49]), .Y(n9453) );
  INVX0_HVT U5810 ( .A(n9453), .Y(n9455) );
  INVX0_HVT U5811 ( .A(n9387), .Y(n9389) );
  INVX0_HVT U5812 ( .A(data[27]), .Y(n9387) );
  INVX0_HVT U5813 ( .A(data[0]), .Y(n9305) );
  INVX0_HVT U5814 ( .A(n9305), .Y(n9307) );
  INVX0_HVT U5815 ( .A(n9885), .Y(n9887) );
  INVX0_HVT U5816 ( .A(n9949), .Y(n9951) );
  INVX0_HVT U5817 ( .A(n10023), .Y(n10025) );
  INVX0_HVT U5818 ( .A(n9784), .Y(n9786) );
  INVX0_HVT U5819 ( .A(n9759), .Y(n9761) );
  INVX0_HVT U5820 ( .A(n9733), .Y(n9735) );
  INVX0_HVT U5821 ( .A(n9973), .Y(n9975) );
  INVX0_HVT U5822 ( .A(n9986), .Y(n9988) );
  INVX0_HVT U5823 ( .A(n9834), .Y(n9836) );
  INVX0_HVT U5824 ( .A(n9898), .Y(n9900) );
  INVX0_HVT U5825 ( .A(n9936), .Y(n9938) );
  INVX0_HVT U5826 ( .A(n9847), .Y(n9849) );
  INVX0_HVT U5827 ( .A(n10060), .Y(n10062) );
  INVX0_HVT U5828 ( .A(n9821), .Y(n9823) );
  INVX0_HVT U5829 ( .A(n9924), .Y(n9926) );
  INVX0_HVT U5830 ( .A(n9771), .Y(n9773) );
  INVX0_HVT U5831 ( .A(n10086), .Y(n10088) );
  INVX0_HVT U5832 ( .A(n9696), .Y(n9698) );
  INVX0_HVT U5833 ( .A(n9860), .Y(n9862) );
  INVX0_HVT U5834 ( .A(n9911), .Y(n9913) );
  INVX0_HVT U5835 ( .A(n9961), .Y(n9963) );
  INVX0_HVT U5836 ( .A(n9708), .Y(n9710) );
  INVX0_HVT U5837 ( .A(n10010), .Y(n10012) );
  INVX0_HVT U5838 ( .A(n9746), .Y(n9748) );
  INVX0_HVT U5839 ( .A(n9809), .Y(n9811) );
  INVX0_HVT U5840 ( .A(n9998), .Y(n10000) );
  INVX0_HVT U5841 ( .A(n10035), .Y(n10037) );
  INVX0_HVT U5842 ( .A(n10334), .Y(n7175) );
  INVX0_HVT U5843 ( .A(n9233), .Y(n9239) );
  INVX0_HVT U5844 ( .A(n9205), .Y(n5117) );
  INVX0_HVT U5845 ( .A(n9233), .Y(n9240) );
  INVX0_HVT U5846 ( .A(n4778), .Y(n6160) );
  OAI22X1_HVT U5847 ( .A1(n5604), .A2(n5382), .A3(n5603), .A4(n9390), .Y(n5036) );
  INVX0_HVT U5848 ( .A(n10163), .Y(n10156) );
  INVX0_HVT U5849 ( .A(n6800), .Y(n10157) );
  INVX0_HVT U5850 ( .A(n6812), .Y(n10155) );
  INVX0_HVT U5851 ( .A(n7428), .Y(n7430) );
  INVX0_HVT U5852 ( .A(n7429), .Y(n7431) );
  INVX0_HVT U5853 ( .A(n7429), .Y(n7466) );
  INVX0_HVT U5854 ( .A(n7429), .Y(n7445) );
  INVX0_HVT U5855 ( .A(n7428), .Y(n7435) );
  INVX0_HVT U5856 ( .A(n7418), .Y(n7420) );
  INVX1_HVT U5857 ( .A(n10187), .Y(n6442) );
  INVX0_HVT U5858 ( .A(n6423), .Y(n6425) );
  INVX0_HVT U5859 ( .A(n6475), .Y(n6477) );
  INVX0_HVT U5860 ( .A(n10251), .Y(n10241) );
  INVX0_HVT U5861 ( .A(n7358), .Y(n10240) );
  INVX1_HVT U5862 ( .A(n10301), .Y(n10295) );
  INVX0_HVT U5863 ( .A(n6248), .Y(n6220) );
  INVX0_HVT U5864 ( .A(n6221), .Y(n6217) );
  INVX0_HVT U5865 ( .A(n10301), .Y(n10297) );
  INVX0_HVT U5866 ( .A(n10301), .Y(n10296) );
  INVX0_HVT U5867 ( .A(n6244), .Y(n6195) );
  INVX0_HVT U5868 ( .A(n6225), .Y(n6216) );
  INVX0_HVT U5869 ( .A(n6247), .Y(n6228) );
  INVX0_HVT U5870 ( .A(n6247), .Y(n6249) );
  INVX0_HVT U5871 ( .A(n6221), .Y(n6201) );
  INVX1_HVT U5872 ( .A(n10360), .Y(n10359) );
  INVX0_HVT U5873 ( .A(n6504), .Y(n6506) );
  INVX0_HVT U5874 ( .A(n6491), .Y(n6492) );
  INVX0_HVT U5875 ( .A(n6519), .Y(n6526) );
  INVX0_HVT U5876 ( .A(n6522), .Y(n6521) );
  INVX0_HVT U5877 ( .A(n4438), .Y(n6525) );
  INVX0_HVT U5878 ( .A(n6519), .Y(n6524) );
  INVX0_HVT U5879 ( .A(n6306), .Y(n6319) );
  INVX0_HVT U5880 ( .A(n6293), .Y(n6267) );
  INVX0_HVT U5881 ( .A(n6293), .Y(n6291) );
  INVX0_HVT U5882 ( .A(n6293), .Y(n6294) );
  INVX0_HVT U5883 ( .A(n10329), .Y(n10320) );
  INVX0_HVT U5884 ( .A(n10329), .Y(n10321) );
  INVX0_HVT U5885 ( .A(n10329), .Y(n10323) );
  INVX0_HVT U5886 ( .A(n10329), .Y(n10322) );
  INVX0_HVT U5887 ( .A(n6277), .Y(n6268) );
  INVX0_HVT U5888 ( .A(n6277), .Y(n6279) );
  INVX0_HVT U5889 ( .A(n6282), .Y(n6290) );
  INVX0_HVT U5890 ( .A(n6283), .Y(n6287) );
  INVX0_HVT U5891 ( .A(n6283), .Y(n6285) );
  INVX0_HVT U5892 ( .A(n6282), .Y(n6275) );
  INVX0_HVT U5893 ( .A(n6283), .Y(n10325) );
  INVX0_HVT U5894 ( .A(n4461), .Y(n6857) );
  INVX0_HVT U5895 ( .A(n4461), .Y(n6856) );
  INVX1_HVT U5896 ( .A(n10343), .Y(n6848) );
  INVX0_HVT U5897 ( .A(n10345), .Y(n6828) );
  INVX0_HVT U5898 ( .A(n6843), .Y(n6829) );
  INVX0_HVT U5899 ( .A(n10340), .Y(n6855) );
  INVX0_HVT U5900 ( .A(n6901), .Y(n10268) );
  INVX0_HVT U5901 ( .A(n6900), .Y(n6902) );
  INVX0_HVT U5902 ( .A(n10269), .Y(n6900) );
  INVX0_HVT U5903 ( .A(n10269), .Y(n6901) );
  INVX0_HVT U5904 ( .A(n6900), .Y(n10265) );
  INVX0_HVT U5905 ( .A(n6923), .Y(n6953) );
  INVX0_HVT U5906 ( .A(n6923), .Y(n6925) );
  INVX0_HVT U5907 ( .A(n6922), .Y(n6938) );
  INVX0_HVT U5908 ( .A(n6922), .Y(n6924) );
  INVX1_HVT U5909 ( .A(n10262), .Y(n6948) );
  INVX1_HVT U5910 ( .A(n10267), .Y(n6949) );
  INVX0_HVT U5911 ( .A(n6935), .Y(n6937) );
  INVX0_HVT U5912 ( .A(n6909), .Y(n6952) );
  INVX0_HVT U5913 ( .A(n6906), .Y(n6939) );
  INVX0_HVT U5914 ( .A(n6906), .Y(n6907) );
  INVX0_HVT U5915 ( .A(n10111), .Y(n10110) );
  INVX0_HVT U5916 ( .A(n10111), .Y(n6893) );
  INVX0_HVT U5917 ( .A(n5749), .Y(n10111) );
  INVX0_HVT U5918 ( .A(n10111), .Y(n10102) );
  INVX0_HVT U5919 ( .A(n6081), .Y(n6083) );
  INVX1_HVT U5920 ( .A(n10230), .Y(n6060) );
  INVX1_HVT U5921 ( .A(n10372), .Y(n6724) );
  INVX0_HVT U5922 ( .A(n10372), .Y(n10374) );
  INVX0_HVT U5923 ( .A(n4511), .Y(n6612) );
  INVX0_HVT U5924 ( .A(n10140), .Y(n6611) );
  INVX0_HVT U5925 ( .A(n4511), .Y(n6613) );
  INVX0_HVT U5926 ( .A(n4511), .Y(n6580) );
  INVX1_HVT U5927 ( .A(n10194), .Y(n7517) );
  INVX1_HVT U5928 ( .A(n10195), .Y(n7516) );
  INVX0_HVT U5929 ( .A(n10193), .Y(n7510) );
  INVX0_HVT U5930 ( .A(n10193), .Y(n7532) );
  INVX0_HVT U5931 ( .A(n7533), .Y(n7535) );
  INVX0_HVT U5932 ( .A(n7510), .Y(n7512) );
  INVX0_HVT U5933 ( .A(n5248), .Y(n5262) );
  INVX0_HVT U5934 ( .A(n5278), .Y(n5261) );
  INVX0_HVT U5935 ( .A(n10307), .Y(n5278) );
  INVX0_HVT U5936 ( .A(n5241), .Y(n5240) );
  INVX0_HVT U5937 ( .A(n5274), .Y(n10311) );
  INVX0_HVT U5938 ( .A(n5348), .Y(n5271) );
  INVX0_HVT U5939 ( .A(n6004), .Y(n5284) );
  INVX0_HVT U5940 ( .A(n10312), .Y(n5241) );
  INVX0_HVT U5941 ( .A(n7589), .Y(n7642) );
  INVX0_HVT U5942 ( .A(n7647), .Y(n7649) );
  INVX0_HVT U5943 ( .A(n7731), .Y(n10221) );
  INVX0_HVT U5944 ( .A(n7647), .Y(n7648) );
  INVX0_HVT U5945 ( .A(n7644), .Y(n7646) );
  INVX0_HVT U5946 ( .A(n7644), .Y(n7645) );
  INVX0_HVT U5947 ( .A(n7620), .Y(n7617) );
  INVX0_HVT U5948 ( .A(n7616), .Y(n7658) );
  INVX0_HVT U5949 ( .A(n7616), .Y(n7643) );
  INVX0_HVT U5950 ( .A(n7633), .Y(n7587) );
  INVX0_HVT U5951 ( .A(n7659), .Y(n7660) );
  INVX0_HVT U5952 ( .A(n7651), .Y(n7654) );
  INVX0_HVT U5953 ( .A(n7651), .Y(n7653) );
  INVX0_HVT U5954 ( .A(n7612), .Y(n7614) );
  INVX0_HVT U5955 ( .A(n7607), .Y(n7618) );
  INVX0_HVT U5956 ( .A(n7607), .Y(n7652) );
  INVX0_HVT U5957 ( .A(n10219), .Y(n10213) );
  INVX0_HVT U5958 ( .A(n7659), .Y(n7662) );
  INVX0_HVT U5959 ( .A(n10220), .Y(n7661) );
  INVX0_HVT U5960 ( .A(n7608), .Y(n7619) );
  INVX0_HVT U5961 ( .A(n7608), .Y(n7609) );
  INVX0_HVT U5962 ( .A(n7608), .Y(n7611) );
  INVX0_HVT U5963 ( .A(n10221), .Y(n10219) );
  INVX0_HVT U5964 ( .A(n10219), .Y(n7588) );
  INVX0_HVT U5965 ( .A(n7731), .Y(n7585) );
  INVX0_HVT U5966 ( .A(n7655), .Y(n7656) );
  INVX0_HVT U5967 ( .A(n7655), .Y(n7657) );
  INVX0_HVT U5968 ( .A(n4463), .Y(n7606) );
  INVX0_HVT U5969 ( .A(n7633), .Y(n7604) );
  INVX0_HVT U5970 ( .A(n7585), .Y(n10220) );
  INVX0_HVT U5971 ( .A(n7593), .Y(n7615) );
  INVX1_HVT U5972 ( .A(n8755), .Y(n6658) );
  INVX0_HVT U5973 ( .A(n5870), .Y(n5318) );
  INVX0_HVT U5974 ( .A(n5805), .Y(n5289) );
  INVX0_HVT U5975 ( .A(n7339), .Y(n5110) );
  INVX0_HVT U5976 ( .A(n5323), .Y(n5101) );
  INVX0_HVT U5977 ( .A(n5306), .Y(n6750) );
  INVX0_HVT U5978 ( .A(n7570), .Y(n5156) );
  INVX0_HVT U5979 ( .A(n5297), .Y(n5867) );
  INVX0_HVT U5980 ( .A(n5901), .Y(n6415) );
  INVX0_HVT U5981 ( .A(n6750), .Y(n6383) );
  INVX0_HVT U5982 ( .A(n6383), .Y(n5207) );
  INVX0_HVT U5983 ( .A(n6383), .Y(n5151) );
  INVX0_HVT U5984 ( .A(n7567), .Y(n7300) );
  INVX0_HVT U5985 ( .A(n7567), .Y(n6756) );
  INVX0_HVT U5986 ( .A(n5623), .Y(n5225) );
  INVX0_HVT U5987 ( .A(n8751), .Y(n8752) );
  INVX0_HVT U5988 ( .A(n6659), .Y(n7685) );
  INVX0_HVT U5989 ( .A(n6749), .Y(n6416) );
  INVX0_HVT U5990 ( .A(n6661), .Y(n5111) );
  INVX0_HVT U5991 ( .A(n6661), .Y(n5354) );
  INVX0_HVT U5992 ( .A(n6383), .Y(n5364) );
  INVX1_HVT U5993 ( .A(n5306), .Y(n6749) );
  INVX0_HVT U5994 ( .A(n8755), .Y(n5321) );
  INVX0_HVT U5995 ( .A(n7339), .Y(n5323) );
  INVX0_HVT U5996 ( .A(n5326), .Y(n5097) );
  INVX0_HVT U5997 ( .A(n5297), .Y(n5172) );
  INVX0_HVT U5998 ( .A(n8760), .Y(n5343) );
  INVX0_HVT U5999 ( .A(n5990), .Y(n5752) );
  INVX0_HVT U6000 ( .A(n7570), .Y(n5078) );
  INVX0_HVT U6001 ( .A(n5634), .Y(n5363) );
  INVX0_HVT U6002 ( .A(n5870), .Y(n5317) );
  INVX0_HVT U6003 ( .A(n8758), .Y(n5352) );
  INVX0_HVT U6004 ( .A(n8760), .Y(n5326) );
  INVX0_HVT U6005 ( .A(n5752), .Y(n7349) );
  INVX1_HVT U6006 ( .A(n5078), .Y(n5634) );
  INVX0_HVT U6007 ( .A(n8782), .Y(n8850) );
  INVX0_HVT U6008 ( .A(n8845), .Y(n6746) );
  INVX0_HVT U6009 ( .A(n8845), .Y(n5201) );
  INVX0_HVT U6010 ( .A(n5448), .Y(n5238) );
  INVX0_HVT U6011 ( .A(n5751), .Y(n5299) );
  INVX0_HVT U6012 ( .A(n8840), .Y(n5113) );
  INVX0_HVT U6013 ( .A(n4837), .Y(n5124) );
  INVX0_HVT U6014 ( .A(n5794), .Y(n5126) );
  INVX0_HVT U6015 ( .A(n5356), .Y(n8823) );
  INVX0_HVT U6016 ( .A(n8813), .Y(n7334) );
  INVX0_HVT U6017 ( .A(n5076), .Y(n5333) );
  INVX0_HVT U6018 ( .A(n8789), .Y(n5982) );
  INVX0_HVT U6019 ( .A(n8823), .Y(n5085) );
  INVX0_HVT U6020 ( .A(n7553), .Y(n5942) );
  INVX0_HVT U6021 ( .A(n8789), .Y(n7557) );
  INVX0_HVT U6022 ( .A(n6136), .Y(n5076) );
  INVX0_HVT U6023 ( .A(n8788), .Y(n8797) );
  INVX0_HVT U6024 ( .A(n5966), .Y(n5633) );
  INVX0_HVT U6025 ( .A(n8788), .Y(n8838) );
  INVX0_HVT U6026 ( .A(n7291), .Y(n7553) );
  INVX0_HVT U6027 ( .A(n2), .Y(n5142) );
  INVX0_HVT U6028 ( .A(n5537), .Y(n5574) );
  INVX0_HVT U6029 ( .A(n5966), .Y(n6031) );
  INVX0_HVT U6030 ( .A(n5571), .Y(n5050) );
  INVX0_HVT U6031 ( .A(n8789), .Y(n5975) );
  INVX0_HVT U6032 ( .A(n8789), .Y(n5966) );
  INVX0_HVT U6033 ( .A(n8789), .Y(n5976) );
  INVX0_HVT U6034 ( .A(n6023), .Y(n5152) );
  NBUFFX2_HVT U6035 ( .A(n5659), .Y(n7706) );
  INVX0_HVT U6036 ( .A(n8905), .Y(n5508) );
  INVX0_HVT U6037 ( .A(n6252), .Y(n5560) );
  INVX0_HVT U6038 ( .A(n5552), .Y(n5950) );
  INVX0_HVT U6039 ( .A(n6663), .Y(n5290) );
  INVX0_HVT U6040 ( .A(n6252), .Y(n5971) );
  INVX0_HVT U6041 ( .A(n7674), .Y(n5336) );
  INVX0_HVT U6042 ( .A(n7148), .Y(n5924) );
  INVX0_HVT U6043 ( .A(n6184), .Y(n7674) );
  INVX0_HVT U6044 ( .A(n5588), .Y(n5584) );
  INVX0_HVT U6045 ( .A(n5986), .Y(n6738) );
  INVX0_HVT U6046 ( .A(n7675), .Y(n5337) );
  INVX0_HVT U6047 ( .A(n6409), .Y(n7340) );
  INVX1_HVT U6048 ( .A(n4926), .Y(n5882) );
  INVX0_HVT U6049 ( .A(n7717), .Y(n5898) );
  INVX0_HVT U6050 ( .A(n7573), .Y(n5093) );
  INVX1_HVT U6051 ( .A(n7677), .Y(n5079) );
  INVX0_HVT U6052 ( .A(n8765), .Y(n7574) );
  INVX0_HVT U6053 ( .A(n7333), .Y(n5298) );
  INVX0_HVT U6054 ( .A(n5312), .Y(n5237) );
  INVX1_HVT U6055 ( .A(n7299), .Y(n5112) );
  INVX0_HVT U6056 ( .A(n7558), .Y(n7272) );
  INVX0_HVT U6057 ( .A(n8770), .Y(n5312) );
  INVX0_HVT U6058 ( .A(n5355), .Y(n5359) );
  INVX0_HVT U6059 ( .A(n5315), .Y(n5307) );
  INVX0_HVT U6060 ( .A(n6033), .Y(n5344) );
  INVX0_HVT U6061 ( .A(n5239), .Y(n5887) );
  INVX0_HVT U6062 ( .A(n5770), .Y(n5291) );
  INVX0_HVT U6063 ( .A(n8770), .Y(n5631) );
  INVX0_HVT U6064 ( .A(n5315), .Y(n5896) );
  INVX0_HVT U6065 ( .A(n8770), .Y(n5721) );
  INVX0_HVT U6066 ( .A(n5770), .Y(n5362) );
  INVX0_HVT U6067 ( .A(n6894), .Y(n7307) );
  INVX1_HVT U6068 ( .A(n7307), .Y(n5536) );
  INVX0_HVT U6069 ( .A(n6033), .Y(n5315) );
  INVX0_HVT U6070 ( .A(n5291), .Y(n5233) );
  INVX0_HVT U6071 ( .A(n5376), .Y(n5136) );
  INVX0_HVT U6072 ( .A(n5827), .Y(n5773) );
  INVX0_HVT U6073 ( .A(n7717), .Y(n5991) );
  INVX0_HVT U6074 ( .A(n8774), .Y(n5373) );
  INVX0_HVT U6075 ( .A(n8770), .Y(n5624) );
  INVX0_HVT U6076 ( .A(n6033), .Y(n5376) );
  INVX0_HVT U6077 ( .A(n5660), .Y(n5162) );
  INVX0_HVT U6078 ( .A(n5877), .Y(n5040) );
  INVX1_HVT U6079 ( .A(n5041), .Y(n5042) );
  MUX41X1_HVT U6080 ( .A1(\ram[5][187] ), .A3(\ram[7][187] ), .A2(
        \ram[4][187] ), .A4(\ram[6][187] ), .S0(n5537), .S1(n5739), .Y(n8479)
         );
  INVX1_HVT U6081 ( .A(n5943), .Y(n5922) );
  INVX0_HVT U6082 ( .A(n5062), .Y(n6147) );
  NAND2X0_HVT U6083 ( .A1(\ram[4][26] ), .A2(n6149), .Y(n5037) );
  NAND2X0_HVT U6084 ( .A1(n10295), .A2(n9385), .Y(n5038) );
  NAND2X0_HVT U6085 ( .A1(n5037), .A2(n5038), .Y(n1111) );
  INVX0_HVT U6086 ( .A(n6758), .Y(n5986) );
  MUX41X1_HVT U6087 ( .A1(n8690), .A3(n8688), .A2(n8689), .A4(n8687), .S0(
        n5156), .S1(n5040), .Y(q[240]) );
  INVX0_HVT U6088 ( .A(n13), .Y(n5041) );
  NAND2X0_HVT U6089 ( .A1(\ram[9][39] ), .A2(n7634), .Y(n5043) );
  NAND2X0_HVT U6090 ( .A1(n9106), .A2(n9425), .Y(n5044) );
  NAND2X0_HVT U6091 ( .A1(n5043), .A2(n5044), .Y(n2404) );
  NAND2X0_HVT U6092 ( .A1(\ram[9][30] ), .A2(n7639), .Y(n5045) );
  NAND2X0_HVT U6093 ( .A1(n9126), .A2(n9398), .Y(n5046) );
  NAND2X0_HVT U6094 ( .A1(n5045), .A2(n5046), .Y(n2395) );
  INVX0_HVT U6095 ( .A(n9396), .Y(n9398) );
  NAND2X0_HVT U6096 ( .A1(\ram[9][29] ), .A2(n7640), .Y(n5047) );
  NAND2X0_HVT U6097 ( .A1(n9126), .A2(data[29]), .Y(n5048) );
  NAND2X0_HVT U6098 ( .A1(n5047), .A2(n5048), .Y(n2394) );
  INVX0_HVT U6099 ( .A(n9120), .Y(n9125) );
  INVX0_HVT U6100 ( .A(n7275), .Y(n8834) );
  INVX0_HVT U6101 ( .A(n7727), .Y(n10178) );
  INVX0_HVT U6102 ( .A(n7263), .Y(n7314) );
  NBUFFX2_HVT U6103 ( .A(n6892), .Y(n5528) );
  INVX0_HVT U6104 ( .A(n5073), .Y(n5049) );
  INVX1_HVT U6105 ( .A(n5732), .Y(n5073) );
  MUX41X1_HVT U6106 ( .A1(\ram[8][242] ), .A3(\ram[10][242] ), .A2(
        \ram[9][242] ), .A4(\ram[11][242] ), .S0(n5537), .S1(n5053), .Y(n8696)
         );
  INVX0_HVT U6107 ( .A(n7319), .Y(n8833) );
  IBUFFX2_HVT U6108 ( .A(n7316), .Y(n8819) );
  MUX41X1_HVT U6109 ( .A1(\ram[10][172] ), .A3(\ram[8][172] ), .A2(
        \ram[11][172] ), .A4(\ram[9][172] ), .S0(n5982), .S1(n6035), .Y(n8418)
         );
  INVX0_HVT U6110 ( .A(n5834), .Y(n5051) );
  INVX0_HVT U6111 ( .A(n5051), .Y(n5052) );
  INVX1_HVT U6112 ( .A(n5049), .Y(n5589) );
  MUX41X1_HVT U6113 ( .A1(\ram[8][155] ), .A3(\ram[10][155] ), .A2(
        \ram[9][155] ), .A4(\ram[11][155] ), .S0(n5058), .S1(n5053), .Y(n8350)
         );
  MUX21X2_HVT U6114 ( .A1(n5744), .A2(n5745), .S0(n5228), .Y(n8062) );
  IBUFFX2_HVT U6115 ( .A(n7286), .Y(n8815) );
  NAND2X0_HVT U6116 ( .A1(n5768), .A2(n5084), .Y(n5057) );
  NAND2X0_HVT U6117 ( .A1(n5056), .A2(n5057), .Y(n7926) );
  INVX0_HVT U6118 ( .A(n8785), .Y(n5058) );
  INVX0_HVT U6119 ( .A(n5058), .Y(n5059) );
  INVX1_HVT U6120 ( .A(n8788), .Y(n5948) );
  IBUFFX2_HVT U6121 ( .A(n7732), .Y(n5663) );
  INVX0_HVT U6122 ( .A(n8839), .Y(n7561) );
  INVX0_HVT U6123 ( .A(n7546), .Y(n8839) );
  MUX41X1_HVT U6124 ( .A1(n8181), .A3(n8179), .A2(n8180), .A4(n8178), .S0(
        n5289), .S1(n8766), .Y(q[112]) );
  INVX0_HVT U6125 ( .A(n10304), .Y(n5060) );
  INVX0_HVT U6126 ( .A(n5060), .Y(n5061) );
  INVX0_HVT U6127 ( .A(n6145), .Y(n10304) );
  MUX41X1_HVT U6128 ( .A1(n8560), .A3(n8558), .A2(n8559), .A4(n8557), .S0(
        n5752), .S1(n5087), .Y(q[207]) );
  INVX0_HVT U6129 ( .A(n7315), .Y(n5107) );
  AO22X1_HVT U6130 ( .A1(\ram[4][209] ), .A2(n4370), .A3(n6250), .A4(n9947), 
        .Y(n1294) );
  AO22X1_HVT U6131 ( .A1(\ram[4][53] ), .A2(n6164), .A3(n6240), .A4(n9466), 
        .Y(n1138) );
  MUX41X1_HVT U6132 ( .A1(n8730), .A3(n8729), .A2(n8728), .A4(n8727), .S0(
        n5162), .S1(n5318), .Y(q[250]) );
  INVX0_HVT U6133 ( .A(n5890), .Y(n5104) );
  IBUFFX2_HVT U6134 ( .A(n5960), .Y(n5759) );
  INVX0_HVT U6135 ( .A(n10305), .Y(n5062) );
  NAND2X0_HVT U6136 ( .A1(\ram[4][62] ), .A2(n4927), .Y(n5063) );
  NAND2X0_HVT U6137 ( .A1(n6208), .A2(n9493), .Y(n5064) );
  NAND2X0_HVT U6138 ( .A1(n5063), .A2(n5064), .Y(n1147) );
  OAI22X1_HVT U6139 ( .A1(n5065), .A2(n5501), .A3(n6247), .A4(n9456), .Y(n1135) );
  INVX0_HVT U6140 ( .A(n6238), .Y(n6243) );
  NAND2X0_HVT U6141 ( .A1(\ram[4][22] ), .A2(n6143), .Y(n5066) );
  NAND2X0_HVT U6142 ( .A1(n6187), .A2(n9373), .Y(n5067) );
  NAND2X0_HVT U6143 ( .A1(n5066), .A2(n5067), .Y(n1107) );
  OAI22X1_HVT U6144 ( .A1(n5068), .A2(n5501), .A3(n6196), .A4(n9336), .Y(n1095) );
  INVX0_HVT U6145 ( .A(n6196), .Y(n6198) );
  NAND2X0_HVT U6146 ( .A1(\ram[4][199] ), .A2(n4928), .Y(n5069) );
  NAND2X0_HVT U6147 ( .A1(n10293), .A2(n9915), .Y(n5070) );
  NAND2X0_HVT U6148 ( .A1(n5069), .A2(n5070), .Y(n1284) );
  INVX0_HVT U6149 ( .A(n7291), .Y(n5793) );
  INVX1_HVT U6150 ( .A(n8893), .Y(n5103) );
  MUX41X1_HVT U6151 ( .A1(\ram[2][9] ), .A3(\ram[0][9] ), .A2(\ram[3][9] ), 
        .A4(\ram[1][9] ), .S0(n5333), .S1(n5316), .Y(n7773) );
  IBUFFX2_HVT U6152 ( .A(n5091), .Y(n8822) );
  MUX41X1_HVT U6153 ( .A1(n8472), .A3(n8470), .A2(n8471), .A4(n8469), .S0(
        n5172), .S1(n5093), .Y(q[185]) );
  INVX0_HVT U6154 ( .A(n5542), .Y(n5487) );
  INVX0_HVT U6155 ( .A(n5487), .Y(n7689) );
  INVX0_HVT U6156 ( .A(n5919), .Y(n5889) );
  AO21X1_HVT U6157 ( .A1(n54), .A2(n10375), .A3(rst), .Y(n5072) );
  MUX41X1_HVT U6158 ( .A1(\ram[4][207] ), .A3(\ram[6][207] ), .A2(
        \ram[5][207] ), .A4(\ram[7][207] ), .S0(n5657), .S1(n5073), .Y(n8559)
         );
  MUX41X1_HVT U6159 ( .A1(\ram[14][203] ), .A3(\ram[12][203] ), .A2(
        \ram[15][203] ), .A4(\ram[13][203] ), .S0(n6660), .S1(n8857), .Y(n8541) );
  MUX21X1_HVT U6160 ( .A1(\ram[12][244] ), .A2(\ram[14][244] ), .S0(n5895), 
        .Y(n5320) );
  INVX1_HVT U6161 ( .A(n5553), .Y(n7146) );
  INVX0_HVT U6162 ( .A(n5166), .Y(n8628) );
  NAND2X0_HVT U6163 ( .A1(\ram[4][54] ), .A2(n5445), .Y(n5074) );
  NAND2X0_HVT U6164 ( .A1(n6237), .A2(n9469), .Y(n5075) );
  NAND2X0_HVT U6165 ( .A1(n5074), .A2(n5075), .Y(n1139) );
  NBUFFX2_HVT U6166 ( .A(n5008), .Y(n7564) );
  MUX41X1_HVT U6167 ( .A1(\ram[0][152] ), .A3(\ram[2][152] ), .A2(
        \ram[1][152] ), .A4(\ram[3][152] ), .S0(n5076), .S1(n5080), .Y(n8340)
         );
  NBUFFX2_HVT U6168 ( .A(n5129), .Y(n6146) );
  INVX0_HVT U6169 ( .A(n7267), .Y(n6407) );
  MUX41X1_HVT U6170 ( .A1(\ram[11][174] ), .A3(\ram[9][174] ), .A2(
        \ram[10][174] ), .A4(\ram[8][174] ), .S0(n5357), .S1(n5077), .Y(n8426)
         );
  MUX41X1_HVT U6171 ( .A1(n8484), .A3(n8482), .A2(n8483), .A4(n8481), .S0(
        n5078), .S1(n5079), .Y(q[188]) );
  MUX41X1_HVT U6172 ( .A1(\ram[12][211] ), .A3(\ram[14][211] ), .A2(
        \ram[13][211] ), .A4(\ram[15][211] ), .S0(n5509), .S1(n5080), .Y(n8573) );
  INVX1_HVT U6173 ( .A(n8898), .Y(n5606) );
  MUX41X1_HVT U6174 ( .A1(\ram[11][253] ), .A3(\ram[9][253] ), .A2(
        \ram[10][253] ), .A4(\ram[8][253] ), .S0(n5299), .S1(n5883), .Y(n8740)
         );
  INVX0_HVT U6175 ( .A(n5740), .Y(n5731) );
  MUX41X1_HVT U6176 ( .A1(\ram[14][200] ), .A3(\ram[12][200] ), .A2(
        \ram[15][200] ), .A4(\ram[13][200] ), .S0(n5124), .S1(n5642), .Y(n8529) );
  IBUFFX2_HVT U6177 ( .A(n5753), .Y(n7317) );
  MUX41X1_HVT U6178 ( .A1(\ram[2][12] ), .A3(\ram[0][12] ), .A2(\ram[3][12] ), 
        .A4(\ram[1][12] ), .S0(n5142), .S1(n5788), .Y(n7785) );
  INVX0_HVT U6179 ( .A(n8790), .Y(n5583) );
  INVX0_HVT U6180 ( .A(n6166), .Y(n6173) );
  NAND2X0_HVT U6181 ( .A1(n8928), .A2(n9317), .Y(n5082) );
  NAND2X0_HVT U6182 ( .A1(n5081), .A2(n5082), .Y(n3392) );
  INVX0_HVT U6183 ( .A(n7016), .Y(n5083) );
  INVX0_HVT U6184 ( .A(n9314), .Y(n9317) );
  MUX21X1_HVT U6185 ( .A1(\ram[0][48] ), .A2(\ram[2][48] ), .S0(n5132), .Y(
        n5768) );
  MUX41X1_HVT U6186 ( .A1(\ram[3][225] ), .A3(\ram[1][225] ), .A2(
        \ram[2][225] ), .A4(\ram[0][225] ), .S0(n5085), .S1(n5230), .Y(n8632)
         );
  INVX0_HVT U6187 ( .A(n5986), .Y(n5964) );
  INVX0_HVT U6188 ( .A(n6166), .Y(n6174) );
  OAI22X1_HVT U6189 ( .A1(n5086), .A2(n5461), .A3(n6225), .A4(n9327), .Y(n1092) );
  INVX0_HVT U6190 ( .A(n5960), .Y(n5155) );
  INVX0_HVT U6191 ( .A(n5960), .Y(n7545) );
  INVX1_HVT U6192 ( .A(n8877), .Y(n5740) );
  INVX0_HVT U6193 ( .A(n5741), .Y(n5353) );
  NAND2X0_HVT U6194 ( .A1(\ram[4][176] ), .A2(n4910), .Y(n5088) );
  NAND2X0_HVT U6195 ( .A1(n6226), .A2(n9842), .Y(n5089) );
  NAND2X0_HVT U6196 ( .A1(n5088), .A2(n5089), .Y(n1261) );
  INVX0_HVT U6197 ( .A(n6224), .Y(n6226) );
  NBUFFX2_HVT U6198 ( .A(n5853), .Y(n8896) );
  MUX41X1_HVT U6199 ( .A1(n8606), .A3(n8605), .A2(n8608), .A4(n8607), .S0(
        n7309), .S1(n6120), .Y(q[219]) );
  INVX0_HVT U6200 ( .A(n5356), .Y(n5310) );
  MUX41X1_HVT U6201 ( .A1(\ram[3][134] ), .A3(\ram[1][134] ), .A2(
        \ram[2][134] ), .A4(\ram[0][134] ), .S0(n5966), .S1(n5118), .Y(n8269)
         );
  INVX0_HVT U6202 ( .A(n6113), .Y(n6755) );
  INVX1_HVT U6203 ( .A(n5128), .Y(n5118) );
  MUX41X1_HVT U6204 ( .A1(n8572), .A3(n8570), .A2(n8571), .A4(n8569), .S0(
        n5799), .S1(n5295), .Y(q[210]) );
  INVX0_HVT U6205 ( .A(n7291), .Y(n5940) );
  MUX41X1_HVT U6206 ( .A1(\ram[5][166] ), .A3(\ram[7][166] ), .A2(
        \ram[4][166] ), .A4(\ram[6][166] ), .S0(n5294), .S1(n5792), .Y(n8395)
         );
  INVX0_HVT U6207 ( .A(n7286), .Y(n5094) );
  INVX0_HVT U6208 ( .A(n7286), .Y(n7287) );
  NBUFFX2_HVT U6209 ( .A(n7708), .Y(n6763) );
  NAND2X0_HVT U6210 ( .A1(\ram[4][5] ), .A2(n6173), .Y(n5095) );
  NAND2X0_HVT U6211 ( .A1(n6219), .A2(n9322), .Y(n5096) );
  NAND2X0_HVT U6212 ( .A1(n5095), .A2(n5096), .Y(n1090) );
  MUX41X1_HVT U6213 ( .A1(n8140), .A3(n8138), .A2(n8141), .A4(n8139), .S0(
        n5097), .S1(n5039), .Y(q[102]) );
  NAND2X0_HVT U6214 ( .A1(\ram[4][145] ), .A2(n6156), .Y(n5098) );
  NAND2X0_HVT U6215 ( .A1(n10294), .A2(n9744), .Y(n5099) );
  NAND2X0_HVT U6216 ( .A1(n5098), .A2(n5099), .Y(n1230) );
  OAI22X1_HVT U6217 ( .A1(n5100), .A2(n4762), .A3(n6248), .A4(n9669), .Y(n1206) );
  INVX0_HVT U6218 ( .A(n8780), .Y(n8786) );
  INVX0_HVT U6219 ( .A(n6733), .Y(n6412) );
  INVX0_HVT U6220 ( .A(n7316), .Y(n6023) );
  INVX0_HVT U6221 ( .A(n4191), .Y(n6765) );
  INVX0_HVT U6222 ( .A(n8852), .Y(n6002) );
  INVX0_HVT U6223 ( .A(n7553), .Y(n5903) );
  IBUFFX2_HVT U6224 ( .A(n5906), .Y(n6131) );
  MUX41X1_HVT U6225 ( .A1(n7931), .A3(n7933), .A2(n7932), .A4(n7934), .S0(
        n5101), .S1(n5102), .Y(q[50]) );
  NBUFFX2_HVT U6226 ( .A(n6386), .Y(n8887) );
  MUX41X1_HVT U6227 ( .A1(\ram[7][251] ), .A3(\ram[5][251] ), .A2(
        \ram[6][251] ), .A4(\ram[4][251] ), .S0(n7314), .S1(n5103), .Y(n8733)
         );
  INVX0_HVT U6228 ( .A(n5961), .Y(n5892) );
  MUX41X1_HVT U6229 ( .A1(\ram[1][148] ), .A3(\ram[3][148] ), .A2(
        \ram[0][148] ), .A4(\ram[2][148] ), .S0(n5750), .S1(n5336), .Y(n8324)
         );
  INVX0_HVT U6230 ( .A(n8862), .Y(n5347) );
  INVX0_HVT U6231 ( .A(n7558), .Y(n5105) );
  INVX0_HVT U6232 ( .A(n5105), .Y(n5106) );
  IBUFFX2_HVT U6233 ( .A(n7319), .Y(n5504) );
  MUX41X1_HVT U6234 ( .A1(\ram[10][228] ), .A3(\ram[8][228] ), .A2(
        \ram[11][228] ), .A4(\ram[9][228] ), .S0(n6660), .S1(n4995), .Y(n8642)
         );
  INVX0_HVT U6235 ( .A(n8780), .Y(n8788) );
  MUX41X1_HVT U6236 ( .A1(\ram[12][225] ), .A3(\ram[14][225] ), .A2(
        \ram[13][225] ), .A4(\ram[15][225] ), .S0(n5294), .S1(n5107), .Y(n8629) );
  NBUFFX2_HVT U6237 ( .A(n7712), .Y(n8882) );
  INVX0_HVT U6238 ( .A(n8327), .Y(n6635) );
  MUX41X1_HVT U6239 ( .A1(n7926), .A3(n7925), .A2(n7924), .A4(n7923), .S0(
        n5109), .S1(n5110), .Y(q[48]) );
  INVX0_HVT U6240 ( .A(n8851), .Y(n6116) );
  MUX41X1_HVT U6241 ( .A1(n7767), .A3(n7769), .A2(n7766), .A4(n7768), .S0(
        n5111), .S1(n5112), .Y(q[8]) );
  MUX41X1_HVT U6242 ( .A1(\ram[1][233] ), .A3(\ram[3][233] ), .A2(
        \ram[0][233] ), .A4(\ram[2][233] ), .S0(n5569), .S1(n7290), .Y(n5115)
         );
  NBUFFX2_HVT U6243 ( .A(n5518), .Y(n5114) );
  MUX41X1_HVT U6244 ( .A1(\ram[15][204] ), .A3(\ram[13][204] ), .A2(
        \ram[14][204] ), .A4(\ram[12][204] ), .S0(n5741), .S1(n7699), .Y(n8545) );
  IBUFFX2_HVT U6245 ( .A(n7267), .Y(n5728) );
  IBUFFX2_HVT U6246 ( .A(n6391), .Y(n5733) );
  NBUFFX2_HVT U6247 ( .A(n6114), .Y(n8874) );
  INVX0_HVT U6248 ( .A(n5651), .Y(n7326) );
  NBUFFX2_HVT U6249 ( .A(n6038), .Y(n7683) );
  MUX41X1_HVT U6250 ( .A1(\ram[15][95] ), .A3(\ram[13][95] ), .A2(
        \ram[14][95] ), .A4(\ram[12][95] ), .S0(n5574), .S1(n5137), .Y(n8110)
         );
  INVX1_HVT U6251 ( .A(n5358), .Y(n5137) );
  MUX41X1_HVT U6252 ( .A1(\ram[2][150] ), .A3(\ram[0][150] ), .A2(
        \ram[3][150] ), .A4(\ram[1][150] ), .S0(n5766), .S1(n5777), .Y(n8332)
         );
  NBUFFX2_HVT U6253 ( .A(n4976), .Y(n7568) );
  NBUFFX2_HVT U6254 ( .A(n5996), .Y(n8905) );
  OA22X2_HVT U6255 ( .A1(n6554), .A2(n6119), .A3(n5117), .A4(n9367), .Y(n5116)
         );
  MUX41X1_HVT U6256 ( .A1(\ram[7][193] ), .A3(\ram[5][193] ), .A2(
        \ram[6][193] ), .A4(\ram[4][193] ), .S0(n5955), .S1(n5137), .Y(n8503)
         );
  INVX0_HVT U6257 ( .A(n6391), .Y(n8849) );
  INVX0_HVT U6258 ( .A(n5747), .Y(n5128) );
  INVX0_HVT U6259 ( .A(n6652), .Y(n5140) );
  NAND2X0_HVT U6260 ( .A1(\ram[5][4] ), .A2(n5677), .Y(n5119) );
  NAND2X0_HVT U6261 ( .A1(n9284), .A2(n9319), .Y(n5120) );
  NAND2X0_HVT U6262 ( .A1(n5119), .A2(n5120), .Y(n1345) );
  INVX0_HVT U6263 ( .A(n5771), .Y(n5121) );
  INVX1_HVT U6264 ( .A(n7703), .Y(n5653) );
  INVX1_HVT U6265 ( .A(n6551), .Y(n5591) );
  MUX41X1_HVT U6266 ( .A1(\ram[12][226] ), .A3(\ram[14][226] ), .A2(
        \ram[13][226] ), .A4(\ram[15][226] ), .S0(n5122), .S1(n8891), .Y(n8633) );
  INVX0_HVT U6267 ( .A(n5907), .Y(n5899) );
  INVX1_HVT U6268 ( .A(n5336), .Y(n5123) );
  MUX41X1_HVT U6269 ( .A1(\ram[2][97] ), .A3(\ram[0][97] ), .A2(\ram[3][97] ), 
        .A4(\ram[1][97] ), .S0(n5787), .S1(n5788), .Y(n8121) );
  INVX0_HVT U6270 ( .A(N29), .Y(n8751) );
  INVX0_HVT U6271 ( .A(n5775), .Y(n5154) );
  MUX41X1_HVT U6272 ( .A1(\ram[7][130] ), .A3(\ram[5][130] ), .A2(
        \ram[6][130] ), .A4(\ram[4][130] ), .S0(n5124), .S1(n7672), .Y(n8252)
         );
  MUX41X1_HVT U6273 ( .A1(\ram[10][176] ), .A3(\ram[8][176] ), .A2(
        \ram[11][176] ), .A4(\ram[9][176] ), .S0(n7306), .S1(n7278), .Y(n8434)
         );
  NBUFFX2_HVT U6274 ( .A(n6030), .Y(n7327) );
  MUX41X1_HVT U6275 ( .A1(\ram[10][117] ), .A3(\ram[8][117] ), .A2(
        \ram[11][117] ), .A4(\ram[9][117] ), .S0(n5125), .S1(n7327), .Y(n8199)
         );
  NBUFFX2_HVT U6276 ( .A(n5008), .Y(n8875) );
  IBUFFX2_HVT U6277 ( .A(n5052), .Y(n10290) );
  IBUFFX2_HVT U6278 ( .A(n8906), .Y(n5874) );
  MUX41X1_HVT U6279 ( .A1(\ram[11][150] ), .A3(\ram[9][150] ), .A2(
        \ram[10][150] ), .A4(\ram[8][150] ), .S0(n5142), .S1(n5127), .Y(n8330)
         );
  IBUFFX2_HVT U6280 ( .A(n7297), .Y(n8831) );
  MUX41X1_HVT U6281 ( .A1(\ram[8][226] ), .A3(\ram[9][226] ), .A2(
        \ram[10][226] ), .A4(\ram[11][226] ), .S0(n5128), .S1(n7554), .Y(n8634) );
  MUX41X1_HVT U6282 ( .A1(n8678), .A3(n8677), .A2(n8676), .A4(n8675), .S0(
        n5136), .S1(n5163), .Y(q[237]) );
  IBUFFX2_HVT U6283 ( .A(n5990), .Y(n5163) );
  INVX0_HVT U6284 ( .A(n10306), .Y(n5129) );
  NBUFFX2_HVT U6285 ( .A(n9), .Y(n5130) );
  MUX41X1_HVT U6286 ( .A1(\ram[7][250] ), .A3(\ram[6][250] ), .A2(
        \ram[5][250] ), .A4(\ram[4][250] ), .S0(n5456), .S1(n5794), .Y(n8729)
         );
  MUX41X1_HVT U6287 ( .A1(n8393), .A3(n8395), .A2(n8394), .A4(n8396), .S0(
        n5326), .S1(n5157), .Y(q[166]) );
  MUX41X1_HVT U6288 ( .A1(\ram[0][133] ), .A3(\ram[2][133] ), .A2(
        \ram[1][133] ), .A4(\ram[3][133] ), .S0(n5132), .S1(n5227), .Y(n8265)
         );
  INVX0_HVT U6289 ( .A(n6127), .Y(n6753) );
  INVX0_HVT U6290 ( .A(n5227), .Y(n5133) );
  INVX0_HVT U6291 ( .A(n7148), .Y(n5227) );
  MUX41X1_HVT U6292 ( .A1(\ram[0][203] ), .A3(\ram[2][203] ), .A2(
        \ram[1][203] ), .A4(\ram[3][203] ), .S0(n5334), .S1(n5134), .Y(n8544)
         );
  NBUFFX2_HVT U6293 ( .A(n5953), .Y(n5135) );
  INVX1_HVT U6294 ( .A(n5137), .Y(n5138) );
  INVX0_HVT U6295 ( .A(n6252), .Y(n5139) );
  INVX0_HVT U6296 ( .A(n5296), .Y(n5358) );
  INVX0_HVT U6297 ( .A(n5651), .Y(n8803) );
  MUX41X1_HVT U6298 ( .A1(\ram[10][181] ), .A3(\ram[8][181] ), .A2(
        \ram[11][181] ), .A4(\ram[9][181] ), .S0(n5142), .S1(n5165), .Y(n8454)
         );
  MUX41X1_HVT U6299 ( .A1(\ram[15][34] ), .A3(\ram[13][34] ), .A2(
        \ram[14][34] ), .A4(\ram[12][34] ), .S0(n6742), .S1(n5735), .Y(n7867)
         );
  INVX1_HVT U6300 ( .A(n7278), .Y(n5735) );
  MUX41X1_HVT U6301 ( .A1(\ram[3][222] ), .A3(\ram[1][222] ), .A2(
        \ram[2][222] ), .A4(\ram[0][222] ), .S0(n5140), .S1(n5351), .Y(n8620)
         );
  IBUFFX2_HVT U6302 ( .A(n5469), .Y(n5611) );
  MUX41X1_HVT U6303 ( .A1(\ram[7][154] ), .A3(\ram[5][154] ), .A2(
        \ram[6][154] ), .A4(\ram[4][154] ), .S0(n7334), .S1(n5141), .Y(n8347)
         );
  INVX0_HVT U6304 ( .A(n5236), .Y(n7710) );
  MUX41X1_HVT U6305 ( .A1(n8122), .A3(n8123), .A2(n8124), .A4(n8125), .S0(
        n6643), .S1(n5575), .Y(q[98]) );
  INVX1_HVT U6306 ( .A(n7566), .Y(n6643) );
  INVX0_HVT U6307 ( .A(n7550), .Y(n5371) );
  INVX0_HVT U6308 ( .A(n8820), .Y(n5955) );
  MUX41X1_HVT U6309 ( .A1(\ram[14][241] ), .A3(\ram[12][241] ), .A2(
        \ram[15][241] ), .A4(\ram[13][241] ), .S0(n5142), .S1(n5143), .Y(n8691) );
  MUX41X1_HVT U6310 ( .A1(\ram[12][231] ), .A3(\ram[14][231] ), .A2(
        \ram[13][231] ), .A4(\ram[15][231] ), .S0(n6021), .S1(n5143), .Y(n8653) );
  INVX1_HVT U6311 ( .A(n5351), .Y(n5144) );
  INVX1_HVT U6312 ( .A(n7568), .Y(n5351) );
  MUX41X1_HVT U6313 ( .A1(\ram[15][116] ), .A3(\ram[13][116] ), .A2(
        \ram[14][116] ), .A4(\ram[12][116] ), .S0(n5152), .S1(n5145), .Y(n8194) );
  IBUFFX2_HVT U6314 ( .A(n6391), .Y(n7084) );
  OAI22X1_HVT U6315 ( .A1(n5146), .A2(n4762), .A3(n6221), .A4(n9324), .Y(n1091) );
  INVX0_HVT U6316 ( .A(n8783), .Y(n8813) );
  INVX1_HVT U6317 ( .A(n5588), .Y(n5148) );
  INVX1_HVT U6318 ( .A(n6135), .Y(n5907) );
  INVX0_HVT U6319 ( .A(n5153), .Y(n5149) );
  INVX0_HVT U6320 ( .A(n5943), .Y(n5153) );
  INVX0_HVT U6321 ( .A(n5208), .Y(n5150) );
  IBUFFX2_HVT U6322 ( .A(n7318), .Y(n5208) );
  MUX41X1_HVT U6323 ( .A1(\ram[12][238] ), .A3(\ram[14][238] ), .A2(
        \ram[13][238] ), .A4(\ram[15][238] ), .S0(n5126), .S1(n5615), .Y(n8679) );
  MUX41X1_HVT U6324 ( .A1(n8513), .A3(n8515), .A2(n8514), .A4(n8516), .S0(
        n5151), .S1(n5199), .Y(q[196]) );
  INVX0_HVT U6325 ( .A(n5785), .Y(n8787) );
  MUX41X1_HVT U6326 ( .A1(\ram[11][35] ), .A3(\ram[9][35] ), .A2(\ram[10][35] ), .A4(\ram[8][35] ), .S0(n5152), .S1(n5747), .Y(n7872) );
  INVX0_HVT U6327 ( .A(n8880), .Y(n5747) );
  MUX41X1_HVT U6328 ( .A1(n8330), .A3(n8332), .A2(n8329), .A4(n8331), .S0(
        n5634), .S1(n5079), .Y(q[150]) );
  MUX41X1_HVT U6329 ( .A1(n8732), .A3(n8731), .A2(n8734), .A4(n8733), .S0(
        n5362), .S1(n5575), .Y(q[251]) );
  MUX41X1_HVT U6330 ( .A1(\ram[13][252] ), .A3(\ram[15][252] ), .A2(
        \ram[12][252] ), .A4(\ram[14][252] ), .S0(n5793), .S1(n5568), .Y(n8735) );
  INVX0_HVT U6331 ( .A(n10304), .Y(n6155) );
  MUX41X1_HVT U6332 ( .A1(\ram[8][191] ), .A3(\ram[10][191] ), .A2(
        \ram[9][191] ), .A4(\ram[11][191] ), .S0(n5360), .S1(n5154), .Y(n8494)
         );
  INVX0_HVT U6333 ( .A(n7674), .Y(n5983) );
  IBUFFX2_HVT U6334 ( .A(n4930), .Y(n5933) );
  MUX41X1_HVT U6335 ( .A1(n8701), .A3(n8699), .A2(n8702), .A4(n8700), .S0(
        n5156), .S1(n5157), .Y(q[243]) );
  OR2X1_HVT U6336 ( .A1(n5468), .A2(n5467), .Y(n5158) );
  NAND2X0_HVT U6337 ( .A1(n5158), .A2(n5159), .Y(n645) );
  INVX0_HVT U6338 ( .A(data[72]), .Y(n9522) );
  NBUFFX2_HVT U6339 ( .A(n17), .Y(n6644) );
  INVX0_HVT U6340 ( .A(n7153), .Y(n7197) );
  MUX41X1_HVT U6341 ( .A1(n8486), .A3(n8488), .A2(n8485), .A4(n8487), .S0(
        n5372), .S1(n5112), .Y(q[189]) );
  MUX41X1_HVT U6342 ( .A1(\ram[7][131] ), .A3(\ram[5][131] ), .A2(
        \ram[6][131] ), .A4(\ram[4][131] ), .S0(n5426), .S1(n5161), .Y(n8256)
         );
  MUX41X1_HVT U6343 ( .A1(n8500), .A3(n8498), .A2(n8499), .A4(n8497), .S0(
        n5225), .S1(n5162), .Y(q[192]) );
  IBUFFX2_HVT U6344 ( .A(n7678), .Y(n5164) );
  INVX0_HVT U6345 ( .A(n6175), .Y(n6182) );
  INVX0_HVT U6346 ( .A(n6252), .Y(n5642) );
  INVX1_HVT U6347 ( .A(n5230), .Y(n5165) );
  MUX41X1_HVT U6348 ( .A1(n5167), .A3(n5033), .A2(n5168), .A4(n5169), .S0(
        n7264), .S1(n7146), .Y(n5166) );
  INVX1_HVT U6349 ( .A(n5753), .Y(n5469) );
  NBUFFX2_HVT U6350 ( .A(n7732), .Y(n5170) );
  INVX0_HVT U6351 ( .A(n5459), .Y(n6180) );
  MUX41X1_HVT U6352 ( .A1(n8300), .A3(n8298), .A2(n8301), .A4(n8299), .S0(
        n6756), .S1(n7301), .Y(q[142]) );
  MUX41X1_HVT U6353 ( .A1(n5115), .A3(n8661), .A2(n8662), .A4(n5965), .S0(
        n5172), .S1(n5808), .Y(q[233]) );
  NBUFFX2_HVT U6354 ( .A(n5178), .Y(n5174) );
  NBUFFX2_HVT U6355 ( .A(n5195), .Y(n5175) );
  NBUFFX2_HVT U6356 ( .A(n5178), .Y(n5176) );
  INVX0_HVT U6357 ( .A(n5754), .Y(n5177) );
  INVX0_HVT U6358 ( .A(n5754), .Y(n5178) );
  NBUFFX2_HVT U6359 ( .A(n5177), .Y(n5179) );
  NBUFFX2_HVT U6360 ( .A(n5177), .Y(n5180) );
  NBUFFX2_HVT U6361 ( .A(n5178), .Y(n5181) );
  NBUFFX2_HVT U6362 ( .A(n5178), .Y(n5182) );
  INVX1_HVT U6363 ( .A(n5195), .Y(n5183) );
  INVX1_HVT U6364 ( .A(n5177), .Y(n5189) );
  INVX1_HVT U6365 ( .A(n5189), .Y(n5191) );
  INVX1_HVT U6366 ( .A(n5189), .Y(n5193) );
  INVX1_HVT U6367 ( .A(n5189), .Y(n5194) );
  OA21X1_HVT U6368 ( .A1(n6118), .A2(n5802), .A3(n5835), .Y(n5195) );
  INVX0_HVT U6369 ( .A(n7715), .Y(n5332) );
  INVX0_HVT U6370 ( .A(n5311), .Y(n5960) );
  IBUFFX2_HVT U6371 ( .A(n5091), .Y(n8796) );
  INVX0_HVT U6372 ( .A(n5947), .Y(n5338) );
  INVX1_HVT U6373 ( .A(n5338), .Y(n5239) );
  NAND2X0_HVT U6374 ( .A1(\ram[4][33] ), .A2(n4395), .Y(n5196) );
  NAND2X0_HVT U6375 ( .A1(n6206), .A2(n9406), .Y(n5197) );
  NAND2X0_HVT U6376 ( .A1(n5196), .A2(n5197), .Y(n1118) );
  OAI22X1_HVT U6377 ( .A1(n5198), .A2(n4762), .A3(n6248), .A4(n9343), .Y(n1097) );
  INVX1_HVT U6378 ( .A(n7279), .Y(n5739) );
  INVX0_HVT U6379 ( .A(n7345), .Y(n5210) );
  INVX0_HVT U6380 ( .A(n5373), .Y(n5324) );
  NBUFFX2_HVT U6381 ( .A(n6739), .Y(n8885) );
  INVX0_HVT U6382 ( .A(n5170), .Y(n5673) );
  AND2X1_HVT U6383 ( .A1(n5217), .A2(n5218), .Y(n5200) );
  MUX41X1_HVT U6384 ( .A1(\ram[7][157] ), .A3(\ram[5][157] ), .A2(
        \ram[6][157] ), .A4(\ram[4][157] ), .S0(n5201), .S1(n5208), .Y(n8359)
         );
  NAND2X0_HVT U6385 ( .A1(\ram[6][47] ), .A2(n5175), .Y(n5202) );
  NAND2X0_HVT U6386 ( .A1(n9197), .A2(n9448), .Y(n5203) );
  NAND2X0_HVT U6387 ( .A1(n5202), .A2(n5203), .Y(n1644) );
  NAND2X0_HVT U6388 ( .A1(\ram[6][39] ), .A2(n5176), .Y(n5204) );
  NAND2X0_HVT U6389 ( .A1(n9219), .A2(n9424), .Y(n5205) );
  NAND2X0_HVT U6390 ( .A1(n5204), .A2(n5205), .Y(n1636) );
  OAI22X1_HVT U6391 ( .A1(n5206), .A2(n5173), .A3(n5117), .A4(n9396), .Y(n1627) );
  MUX41X1_HVT U6392 ( .A1(n8692), .A3(n8694), .A2(n8691), .A4(n8693), .S0(
        n5207), .S1(n5808), .Y(q[241]) );
  MUX41X1_HVT U6393 ( .A1(\ram[7][37] ), .A3(\ram[5][37] ), .A2(\ram[6][37] ), 
        .A4(\ram[4][37] ), .S0(n7572), .S1(n5208), .Y(n7881) );
  NBUFFX2_HVT U6394 ( .A(n7175), .Y(n5209) );
  MUX41X1_HVT U6395 ( .A1(\ram[14][209] ), .A3(\ram[12][209] ), .A2(
        \ram[15][209] ), .A4(\ram[13][209] ), .S0(n7682), .S1(n5210), .Y(n8565) );
  NAND2X0_HVT U6396 ( .A1(\ram[2][129] ), .A2(n7164), .Y(n5211) );
  NAND2X0_HVT U6397 ( .A1(n10324), .A2(n9694), .Y(n5212) );
  NAND2X0_HVT U6398 ( .A1(n5211), .A2(n5212), .Y(n702) );
  NAND2X0_HVT U6399 ( .A1(\ram[2][128] ), .A2(n7167), .Y(n5213) );
  NAND2X0_HVT U6400 ( .A1(n6298), .A2(n9691), .Y(n5214) );
  NAND2X0_HVT U6401 ( .A1(n5213), .A2(n5214), .Y(n701) );
  NAND2X0_HVT U6402 ( .A1(\ram[2][7] ), .A2(n7166), .Y(n5215) );
  NAND2X0_HVT U6403 ( .A1(n6272), .A2(n9328), .Y(n5216) );
  NAND2X0_HVT U6404 ( .A1(n5215), .A2(n5216), .Y(n580) );
  NAND2X0_HVT U6405 ( .A1(n16), .A2(n5645), .Y(n5217) );
  INVX0_HVT U6406 ( .A(n6269), .Y(n6272) );
  INVX0_HVT U6407 ( .A(n10378), .Y(n5645) );
  MUX41X1_HVT U6408 ( .A1(\ram[6][191] ), .A3(\ram[4][191] ), .A2(
        \ram[7][191] ), .A4(\ram[5][191] ), .S0(n5982), .S1(n5290), .Y(n8495)
         );
  IBUFFX2_HVT U6409 ( .A(n5988), .Y(n7329) );
  NAND2X0_HVT U6410 ( .A1(\ram[6][32] ), .A2(n5188), .Y(n5219) );
  NAND2X0_HVT U6411 ( .A1(n9237), .A2(n9403), .Y(n5220) );
  NAND2X0_HVT U6412 ( .A1(n5219), .A2(n5220), .Y(n1629) );
  INVX0_HVT U6413 ( .A(n9232), .Y(n9237) );
  NAND2X0_HVT U6414 ( .A1(\ram[6][31] ), .A2(n5185), .Y(n5221) );
  NAND2X0_HVT U6415 ( .A1(n9238), .A2(n9400), .Y(n5222) );
  NAND2X0_HVT U6416 ( .A1(n5221), .A2(n5222), .Y(n1628) );
  INVX0_HVT U6417 ( .A(n9233), .Y(n9238) );
  NAND2X0_HVT U6418 ( .A1(\ram[6][235] ), .A2(n5186), .Y(n5223) );
  NAND2X0_HVT U6419 ( .A1(n9219), .A2(n10027), .Y(n5224) );
  NAND2X0_HVT U6420 ( .A1(n5223), .A2(n5224), .Y(n1832) );
  INVX0_HVT U6421 ( .A(n7326), .Y(n5878) );
  MUX41X1_HVT U6422 ( .A1(\ram[15][127] ), .A3(\ram[13][127] ), .A2(
        \ram[14][127] ), .A4(\ram[12][127] ), .S0(n5113), .S1(n5228), .Y(n8238) );
  MUX41X1_HVT U6423 ( .A1(n7897), .A3(n7895), .A2(n7898), .A4(n7896), .S0(
        n5225), .S1(n5757), .Y(q[41]) );
  MUX41X1_HVT U6424 ( .A1(\ram[6][41] ), .A3(\ram[4][41] ), .A2(\ram[7][41] ), 
        .A4(\ram[5][41] ), .S0(n6742), .S1(n7579), .Y(n7897) );
  INVX0_HVT U6425 ( .A(n5972), .Y(n5226) );
  MUX41X1_HVT U6426 ( .A1(\ram[0][151] ), .A3(\ram[1][151] ), .A2(
        \ram[2][151] ), .A4(\ram[3][151] ), .S0(n5227), .S1(n7264), .Y(n8336)
         );
  NBUFFX2_HVT U6427 ( .A(n6135), .Y(n5228) );
  INVX0_HVT U6428 ( .A(n5588), .Y(n5869) );
  INVX1_HVT U6429 ( .A(n6637), .Y(n6736) );
  INVX0_HVT U6430 ( .A(n7693), .Y(n5293) );
  NBUFFX2_HVT U6431 ( .A(n6032), .Y(n8888) );
  INVX1_HVT U6432 ( .A(n6747), .Y(n5485) );
  INVX0_HVT U6433 ( .A(n6116), .Y(n6117) );
  INVX0_HVT U6434 ( .A(n5739), .Y(n5578) );
  MUX41X1_HVT U6435 ( .A1(\ram[12][45] ), .A3(\ram[14][45] ), .A2(
        \ram[13][45] ), .A4(\ram[15][45] ), .S0(n5231), .S1(n5505), .Y(n7911)
         );
  INVX1_HVT U6436 ( .A(n7279), .Y(n5607) );
  INVX0_HVT U6437 ( .A(n5505), .Y(n5232) );
  INVX0_HVT U6438 ( .A(n6637), .Y(n7150) );
  MUX41X1_HVT U6439 ( .A1(\ram[11][22] ), .A3(\ram[10][22] ), .A2(\ram[9][22] ), .A4(\ram[8][22] ), .S0(n5336), .S1(n5335), .Y(n7821) );
  MUX41X1_HVT U6440 ( .A1(n8747), .A3(n8749), .A2(n8748), .A4(n8750), .S0(
        n6120), .S1(n5233), .Y(q[255]) );
  INVX1_HVT U6441 ( .A(n10380), .Y(n8763) );
  INVX0_HVT U6442 ( .A(n4514), .Y(n8754) );
  MUX41X1_HVT U6443 ( .A1(\ram[14][254] ), .A3(\ram[12][254] ), .A2(
        \ram[15][254] ), .A4(\ram[13][254] ), .S0(n5955), .S1(n5505), .Y(n8743) );
  INVX0_HVT U6444 ( .A(n5921), .Y(n6638) );
  MUX41X1_HVT U6445 ( .A1(\ram[4][150] ), .A3(\ram[6][150] ), .A2(
        \ram[5][150] ), .A4(\ram[7][150] ), .S0(n8841), .S1(n6417), .Y(n8331)
         );
  MUX41X1_HVT U6446 ( .A1(\ram[3][174] ), .A3(\ram[1][174] ), .A2(
        \ram[2][174] ), .A4(\ram[0][174] ), .S0(n5234), .S1(n43), .Y(n8428) );
  INVX0_HVT U6447 ( .A(n7678), .Y(n5235) );
  MUX41X1_HVT U6448 ( .A1(\ram[11][251] ), .A3(\ram[10][251] ), .A2(
        \ram[9][251] ), .A4(\ram[8][251] ), .S0(n5351), .S1(n7303), .Y(n8732)
         );
  MUX41X1_HVT U6449 ( .A1(n8071), .A3(n8073), .A2(n8070), .A4(n8072), .S0(
        n5736), .S1(n5237), .Y(q[85]) );
  MUX41X1_HVT U6450 ( .A1(\ram[8][254] ), .A3(\ram[10][254] ), .A2(
        \ram[9][254] ), .A4(\ram[11][254] ), .S0(n5238), .S1(n4995), .Y(n8744)
         );
  INVX0_HVT U6451 ( .A(n8787), .Y(n6017) );
  INVX1_HVT U6452 ( .A(n5296), .Y(n7318) );
  INVX0_HVT U6453 ( .A(n8863), .Y(n5486) );
  MUX41X1_HVT U6454 ( .A1(\ram[0][231] ), .A3(\ram[2][231] ), .A2(
        \ram[1][231] ), .A4(\ram[3][231] ), .S0(n5360), .S1(n5572), .Y(n8656)
         );
  IBUFFX2_HVT U6455 ( .A(n5785), .Y(n6405) );
  NBUFFX2_HVT U6456 ( .A(n8871), .Y(n6137) );
  IBUFFX2_HVT U6457 ( .A(n6391), .Y(n8847) );
  MUX41X1_HVT U6458 ( .A1(\ram[7][164] ), .A3(\ram[5][164] ), .A2(
        \ram[6][164] ), .A4(\ram[4][164] ), .S0(n6742), .S1(n5658), .Y(n8387)
         );
  INVX0_HVT U6459 ( .A(n5367), .Y(n5242) );
  INVX1_HVT U6460 ( .A(n5242), .Y(n5243) );
  INVX0_HVT U6461 ( .A(n10310), .Y(n5244) );
  INVX0_HVT U6462 ( .A(n10308), .Y(n5246) );
  INVX0_HVT U6463 ( .A(n10307), .Y(n5248) );
  INVX1_HVT U6464 ( .A(n5241), .Y(n5250) );
  INVX0_HVT U6465 ( .A(n6004), .Y(n5253) );
  INVX0_HVT U6466 ( .A(n6766), .Y(n5257) );
  INVX0_HVT U6467 ( .A(n10310), .Y(n5259) );
  INVX1_HVT U6468 ( .A(n5259), .Y(n5260) );
  INVX0_HVT U6469 ( .A(n6254), .Y(n5263) );
  INVX1_HVT U6470 ( .A(n5263), .Y(n5264) );
  INVX0_HVT U6471 ( .A(n5804), .Y(n5265) );
  INVX0_HVT U6472 ( .A(n10308), .Y(n5268) );
  INVX1_HVT U6473 ( .A(n5268), .Y(n5269) );
  INVX1_HVT U6474 ( .A(n5271), .Y(n5272) );
  INVX1_HVT U6475 ( .A(n5271), .Y(n5273) );
  INVX1_HVT U6476 ( .A(n5274), .Y(n5275) );
  INVX1_HVT U6477 ( .A(n5282), .Y(n5280) );
  INVX0_HVT U6478 ( .A(n5367), .Y(n5368) );
  INVX0_HVT U6479 ( .A(n5271), .Y(n10313) );
  INVX0_HVT U6480 ( .A(n5242), .Y(n6768) );
  INVX0_HVT U6481 ( .A(n5241), .Y(n6766) );
  INVX0_HVT U6482 ( .A(n5242), .Y(n6004) );
  INVX0_HVT U6483 ( .A(n5368), .Y(n6254) );
  INVX0_HVT U6484 ( .A(n5368), .Y(n5804) );
  NBUFFX2_HVT U6485 ( .A(n5819), .Y(n7569) );
  INVX1_HVT U6486 ( .A(n5303), .Y(n5302) );
  INVX0_HVT U6487 ( .A(n5309), .Y(n5287) );
  INVX0_HVT U6488 ( .A(n5791), .Y(n5341) );
  MUX41X1_HVT U6489 ( .A1(\ram[3][207] ), .A3(\ram[1][207] ), .A2(
        \ram[2][207] ), .A4(\ram[0][207] ), .S0(n5817), .S1(n5161), .Y(n8560)
         );
  INVX0_HVT U6490 ( .A(n6626), .Y(n8802) );
  INVX0_HVT U6491 ( .A(n5608), .Y(n5865) );
  INVX0_HVT U6492 ( .A(n8884), .Y(n5288) );
  NBUFFX2_HVT U6493 ( .A(n4976), .Y(n8884) );
  IBUFFX2_HVT U6494 ( .A(n6381), .Y(n5800) );
  NBUFFX2_HVT U6495 ( .A(n5331), .Y(n6663) );
  MUX41X1_HVT U6496 ( .A1(\ram[15][186] ), .A3(\ram[13][186] ), .A2(
        \ram[14][186] ), .A4(\ram[12][186] ), .S0(n7557), .S1(n5300), .Y(n8473) );
  INVX1_HVT U6497 ( .A(n8904), .Y(n5792) );
  NBUFFX2_HVT U6498 ( .A(n8885), .Y(n5292) );
  MUX41X1_HVT U6499 ( .A1(n8713), .A3(n8714), .A2(n8711), .A4(n8712), .S0(
        n5308), .S1(n5318), .Y(q[246]) );
  MUX41X1_HVT U6500 ( .A1(\ram[10][90] ), .A3(\ram[11][90] ), .A2(\ram[8][90] ), .A4(\ram[9][90] ), .S0(n5506), .S1(n7304), .Y(n8091) );
  INVX0_HVT U6501 ( .A(n5510), .Y(n5506) );
  MUX41X1_HVT U6502 ( .A1(\ram[9][184] ), .A3(\ram[11][184] ), .A2(
        \ram[8][184] ), .A4(\ram[10][184] ), .S0(n5322), .S1(n5293), .Y(n8466)
         );
  MUX41X1_HVT U6503 ( .A1(\ram[12][148] ), .A3(\ram[14][148] ), .A2(
        \ram[13][148] ), .A4(\ram[15][148] ), .S0(n5294), .S1(n5138), .Y(n8321) );
  MUX41X1_HVT U6504 ( .A1(\ram[12][251] ), .A3(\ram[14][251] ), .A2(
        \ram[13][251] ), .A4(\ram[15][251] ), .S0(n8796), .S1(n5924), .Y(n8731) );
  MUX41X1_HVT U6505 ( .A1(n8094), .A3(n8096), .A2(n8095), .A4(n8097), .S0(
        n5305), .S1(n6396), .Y(q[91]) );
  MUX41X1_HVT U6506 ( .A1(n8091), .A3(n8093), .A2(n8090), .A4(n8092), .S0(
        n5723), .S1(n5295), .Y(q[90]) );
  INVX0_HVT U6507 ( .A(n7711), .Y(n5570) );
  INVX0_HVT U6508 ( .A(n6117), .Y(n5296) );
  MUX41X1_HVT U6509 ( .A1(n8107), .A3(n8109), .A2(n8106), .A4(n8108), .S0(
        n5297), .S1(n5298), .Y(q[94]) );
  INVX0_HVT U6510 ( .A(n10112), .Y(n5749) );
  IBUFFX2_HVT U6511 ( .A(n7711), .Y(n5629) );
  IBUFFX2_HVT U6512 ( .A(n7711), .Y(n5470) );
  MUX41X1_HVT U6513 ( .A1(\ram[11][91] ), .A3(\ram[9][91] ), .A2(\ram[10][91] ), .A4(\ram[8][91] ), .S0(n5357), .S1(n5541), .Y(n8095) );
  INVX1_HVT U6514 ( .A(n8904), .Y(n5541) );
  MUX41X1_HVT U6515 ( .A1(\ram[15][191] ), .A3(\ram[13][191] ), .A2(
        \ram[14][191] ), .A4(\ram[12][191] ), .S0(n5299), .S1(n5325), .Y(n8493) );
  INVX0_HVT U6516 ( .A(n6763), .Y(n5325) );
  MUX41X1_HVT U6517 ( .A1(\ram[9][204] ), .A3(\ram[11][204] ), .A2(
        \ram[8][204] ), .A4(\ram[10][204] ), .S0(n5238), .S1(n5457), .Y(n8546)
         );
  INVX0_HVT U6518 ( .A(n7279), .Y(n5300) );
  NBUFFX2_HVT U6519 ( .A(n7151), .Y(n8892) );
  NAND2X0_HVT U6520 ( .A1(n8), .A2(n5619), .Y(n5301) );
  NBUFFX2_HVT U6521 ( .A(n7151), .Y(n6743) );
  INVX1_HVT U6522 ( .A(n5309), .Y(n5303) );
  INVX0_HVT U6523 ( .A(n5573), .Y(n5304) );
  NBUFFX2_HVT U6524 ( .A(n6038), .Y(n5573) );
  INVX1_HVT U6525 ( .A(n8867), .Y(n7711) );
  INVX0_HVT U6526 ( .A(n7346), .Y(n7347) );
  MUX41X1_HVT U6527 ( .A1(n8276), .A3(n8274), .A2(n8277), .A4(n8275), .S0(
        n5317), .S1(n5871), .Y(q[136]) );
  INVX0_HVT U6528 ( .A(n7284), .Y(n5334) );
  INVX0_HVT U6529 ( .A(n8751), .Y(n5306) );
  MUX41X1_HVT U6530 ( .A1(n8432), .A3(n8430), .A2(n8431), .A4(n8429), .S0(
        n5867), .S1(n5307), .Y(q[175]) );
  MUX41X1_HVT U6531 ( .A1(\ram[2][175] ), .A3(\ram[0][175] ), .A2(
        \ram[3][175] ), .A4(\ram[1][175] ), .S0(n5104), .S1(n8885), .Y(n8432)
         );
  INVX0_HVT U6532 ( .A(n5356), .Y(n8817) );
  MUX41X1_HVT U6533 ( .A1(\ram[15][202] ), .A3(\ram[13][202] ), .A2(
        \ram[14][202] ), .A4(\ram[12][202] ), .S0(n5942), .S1(n7340), .Y(n8537) );
  INVX0_HVT U6534 ( .A(n8752), .Y(n7544) );
  MUX41X1_HVT U6535 ( .A1(\ram[3][232] ), .A3(\ram[1][232] ), .A2(
        \ram[2][232] ), .A4(\ram[0][232] ), .S0(n5371), .S1(n5309), .Y(n8660)
         );
  INVX1_HVT U6536 ( .A(n5325), .Y(n5316) );
  INVX0_HVT U6537 ( .A(n5501), .Y(n5502) );
  INVX0_HVT U6538 ( .A(n4777), .Y(n5501) );
  NBUFFX2_HVT U6539 ( .A(n8779), .Y(n5311) );
  INVX0_HVT U6540 ( .A(n8779), .Y(n8780) );
  MUX41X1_HVT U6541 ( .A1(n8306), .A3(n8308), .A2(n8307), .A4(n4876), .S0(
        n5372), .S1(n5312), .Y(q[144]) );
  MUX41X1_HVT U6542 ( .A1(n8473), .A3(n8475), .A2(n8474), .A4(n8476), .S0(
        n7567), .S1(n5871), .Y(q[186]) );
  MUX41X1_HVT U6543 ( .A1(n8024), .A3(n8022), .A2(n8025), .A4(n8023), .S0(
        n8760), .S1(n5376), .Y(q[73]) );
  IBUFFX2_HVT U6544 ( .A(n5610), .Y(n7682) );
  NBUFFX2_HVT U6545 ( .A(n6035), .Y(n5313) );
  INVX0_HVT U6546 ( .A(n7712), .Y(n6184) );
  INVX1_HVT U6547 ( .A(n5983), .Y(n5921) );
  MUX41X1_HVT U6548 ( .A1(n8477), .A3(n8479), .A2(n8478), .A4(n8480), .S0(
        n5891), .S1(n5315), .Y(q[187]) );
  MUX21X1_HVT U6549 ( .A1(\ram[15][244] ), .A2(\ram[13][244] ), .S0(n5371), 
        .Y(n5319) );
  MUX41X1_HVT U6550 ( .A1(\ram[4][91] ), .A3(\ram[6][91] ), .A2(\ram[5][91] ), 
        .A4(\ram[7][91] ), .S0(n5000), .S1(n6411), .Y(n8096) );
  MUX41X1_HVT U6551 ( .A1(n7910), .A3(n7908), .A2(n7909), .A4(n7907), .S0(
        n5323), .S1(n5324), .Y(q[44]) );
  MUX41X1_HVT U6552 ( .A1(\ram[11][215] ), .A3(\ram[9][215] ), .A2(
        \ram[10][215] ), .A4(\ram[8][215] ), .S0(n5970), .S1(n5325), .Y(n8590)
         );
  NAND2X0_HVT U6553 ( .A1(n5280), .A2(n9309), .Y(n5328) );
  NAND2X0_HVT U6554 ( .A1(n5327), .A2(n5328), .Y(n830) );
  MUX41X1_HVT U6555 ( .A1(n8020), .A3(n8018), .A2(n8021), .A4(n8019), .S0(
        n5110), .S1(n5332), .Y(q[72]) );
  INVX0_HVT U6556 ( .A(n5331), .Y(n7663) );
  NBUFFX2_HVT U6557 ( .A(n5358), .Y(n7323) );
  MUX41X1_HVT U6558 ( .A1(\ram[3][71] ), .A3(\ram[1][71] ), .A2(\ram[2][71] ), 
        .A4(\ram[0][71] ), .S0(n5333), .S1(n1633), .Y(n8017) );
  INVX0_HVT U6559 ( .A(n5293), .Y(n5788) );
  NBUFFX2_HVT U6560 ( .A(n6891), .Y(n7686) );
  INVX0_HVT U6561 ( .A(N27), .Y(n7346) );
  MUX41X1_HVT U6562 ( .A1(\ram[8][214] ), .A3(\ram[10][214] ), .A2(
        \ram[9][214] ), .A4(\ram[11][214] ), .S0(n5334), .S1(n5950), .Y(n8586)
         );
  INVX0_HVT U6563 ( .A(n6116), .Y(n8852) );
  NBUFFX2_HVT U6564 ( .A(n7151), .Y(n7575) );
  INVX0_HVT U6565 ( .A(n7663), .Y(n5552) );
  MUX41X1_HVT U6566 ( .A1(n8669), .A3(n8667), .A2(n8670), .A4(n8668), .S0(
        n5163), .S1(n5820), .Y(q[235]) );
  NBUFFX2_HVT U6567 ( .A(n6737), .Y(n7675) );
  INVX1_HVT U6568 ( .A(n5653), .Y(n5365) );
  MUX41X1_HVT U6569 ( .A1(\ram[7][10] ), .A3(\ram[5][10] ), .A2(\ram[6][10] ), 
        .A4(\ram[4][10] ), .S0(n5824), .S1(n7331), .Y(n7776) );
  MUX41X1_HVT U6570 ( .A1(\ram[11][115] ), .A3(\ram[9][115] ), .A2(
        \ram[10][115] ), .A4(\ram[8][115] ), .S0(n5970), .S1(n5229), .Y(n8191)
         );
  MUX41X1_HVT U6571 ( .A1(n8002), .A3(n8004), .A2(n8003), .A4(n8005), .S0(
        n5343), .S1(n5373), .Y(q[68]) );
  MUX41X1_HVT U6572 ( .A1(n8548), .A3(n8546), .A2(n8547), .A4(n8545), .S0(
        n5110), .S1(n5339), .Y(q[204]) );
  MUX41X1_HVT U6573 ( .A1(n8635), .A3(n8633), .A2(n8636), .A4(n8634), .S0(
        n5340), .S1(n5341), .Y(q[226]) );
  MUX41X1_HVT U6574 ( .A1(\ram[3][217] ), .A3(\ram[1][217] ), .A2(
        \ram[2][217] ), .A4(\ram[0][217] ), .S0(n5605), .S1(n7331), .Y(n8600)
         );
  MUX41X1_HVT U6575 ( .A1(n8154), .A3(n8156), .A2(n8155), .A4(n8157), .S0(
        n5343), .S1(n5344), .Y(q[106]) );
  INVX0_HVT U6576 ( .A(n7668), .Y(n5345) );
  NBUFFX2_HVT U6577 ( .A(n6765), .Y(n8883) );
  INVX0_HVT U6578 ( .A(n5906), .Y(n7692) );
  NBUFFX2_HVT U6579 ( .A(n8871), .Y(n8862) );
  INVX0_HVT U6580 ( .A(n5301), .Y(n5348) );
  INVX0_HVT U6581 ( .A(n7701), .Y(n5658) );
  MUX41X1_HVT U6582 ( .A1(\ram[11][12] ), .A3(\ram[9][12] ), .A2(\ram[10][12] ), .A4(\ram[8][12] ), .S0(n5201), .S1(n6655), .Y(n7783) );
  INVX0_HVT U6583 ( .A(n7150), .Y(n6891) );
  MUX41X1_HVT U6584 ( .A1(\ram[11][247] ), .A3(\ram[9][247] ), .A2(
        \ram[10][247] ), .A4(\ram[8][247] ), .S0(n5085), .S1(n5496), .Y(n8716)
         );
  MUX41X1_HVT U6585 ( .A1(n8666), .A3(n8664), .A2(n8665), .A4(n8663), .S0(
        n5156), .S1(n5093), .Y(q[234]) );
  INVX0_HVT U6586 ( .A(N27), .Y(n8779) );
  MUX41X1_HVT U6587 ( .A1(n8617), .A3(n8619), .A2(n8618), .A4(n8620), .S0(
        n5352), .S1(n5308), .Y(q[222]) );
  INVX1_HVT U6588 ( .A(n5796), .Y(n5760) );
  MUX41X1_HVT U6589 ( .A1(n8566), .A3(n8568), .A2(n8565), .A4(n8567), .S0(
        n5354), .S1(n5355), .Y(q[209]) );
  MUX41X1_HVT U6590 ( .A1(\ram[7][158] ), .A3(\ram[5][158] ), .A2(
        \ram[6][158] ), .A4(\ram[4][158] ), .S0(n5299), .S1(n5722), .Y(n8363)
         );
  MUX41X1_HVT U6591 ( .A1(\ram[7][152] ), .A3(\ram[5][152] ), .A2(
        \ram[6][152] ), .A4(\ram[4][152] ), .S0(n5357), .S1(n5722), .Y(n8339)
         );
  MUX41X1_HVT U6592 ( .A1(n8294), .A3(n8295), .A2(n8296), .A4(n8297), .S0(
        n5359), .S1(n5131), .Y(q[141]) );
  INVX0_HVT U6593 ( .A(n5496), .Y(n5361) );
  NBUFFX2_HVT U6594 ( .A(n6030), .Y(n8891) );
  INVX0_HVT U6595 ( .A(n7144), .Y(n6637) );
  MUX41X1_HVT U6596 ( .A1(\ram[11][244] ), .A3(\ram[9][244] ), .A2(
        \ram[10][244] ), .A4(\ram[8][244] ), .S0(n5969), .S1(n5377), .Y(n8704)
         );
  MUX41X1_HVT U6597 ( .A1(n8269), .A3(n8267), .A2(n8268), .A4(n8266), .S0(
        n5363), .S1(n5635), .Y(q[134]) );
  MUX41X1_HVT U6598 ( .A1(n8263), .A3(n8265), .A2(n8262), .A4(n8264), .S0(
        n5364), .S1(n6388), .Y(q[133]) );
  MUX41X1_HVT U6599 ( .A1(\ram[0][198] ), .A3(\ram[2][198] ), .A2(
        \ram[1][198] ), .A4(\ram[3][198] ), .S0(n5750), .S1(n5365), .Y(n8524)
         );
  INVX0_HVT U6600 ( .A(n5936), .Y(n5367) );
  MUX41X1_HVT U6601 ( .A1(\ram[14][153] ), .A3(\ram[12][153] ), .A2(
        \ram[15][153] ), .A4(\ram[13][153] ), .S0(n5970), .S1(n5370), .Y(n8341) );
  INVX0_HVT U6602 ( .A(n5981), .Y(n10312) );
  INVX0_HVT U6603 ( .A(N29), .Y(n10380) );
  MUX41X1_HVT U6604 ( .A1(n8453), .A3(n8455), .A2(n8454), .A4(n8456), .S0(
        n5297), .S1(n5376), .Y(q[181]) );
  INVX1_HVT U6605 ( .A(n5358), .Y(n5722) );
  MUX41X1_HVT U6606 ( .A1(\ram[15][176] ), .A3(\ram[14][176] ), .A2(
        \ram[13][176] ), .A4(\ram[12][176] ), .S0(n5377), .S1(n7284), .Y(n8433) );
  INVX0_HVT U6607 ( .A(n5406), .Y(n5378) );
  INVX0_HVT U6608 ( .A(n5425), .Y(n5379) );
  INVX0_HVT U6609 ( .A(n5406), .Y(n5380) );
  INVX0_HVT U6610 ( .A(n5421), .Y(n5381) );
  INVX0_HVT U6611 ( .A(n5413), .Y(n5382) );
  NBUFFX2_HVT U6612 ( .A(n6761), .Y(n5385) );
  NBUFFX2_HVT U6613 ( .A(n10098), .Y(n5386) );
  NBUFFX2_HVT U6614 ( .A(n5600), .Y(n5387) );
  NBUFFX2_HVT U6615 ( .A(n6760), .Y(n5388) );
  NBUFFX2_HVT U6616 ( .A(n10104), .Y(n5389) );
  NBUFFX2_HVT U6617 ( .A(n10101), .Y(n5390) );
  NBUFFX2_HVT U6618 ( .A(n10101), .Y(n5391) );
  NBUFFX2_HVT U6619 ( .A(n10100), .Y(n5392) );
  NBUFFX2_HVT U6620 ( .A(n10100), .Y(n5393) );
  NBUFFX2_HVT U6621 ( .A(n10107), .Y(n5394) );
  NBUFFX2_HVT U6622 ( .A(n10107), .Y(n5395) );
  NBUFFX2_HVT U6623 ( .A(n10098), .Y(n5396) );
  NBUFFX2_HVT U6624 ( .A(n10101), .Y(n5397) );
  NBUFFX2_HVT U6625 ( .A(n10101), .Y(n5398) );
  NBUFFX2_HVT U6626 ( .A(n10104), .Y(n5399) );
  NBUFFX2_HVT U6627 ( .A(n10104), .Y(n5400) );
  NBUFFX2_HVT U6628 ( .A(n10105), .Y(n5401) );
  NBUFFX2_HVT U6629 ( .A(n6760), .Y(n5402) );
  NBUFFX2_HVT U6630 ( .A(n6761), .Y(n5403) );
  NBUFFX2_HVT U6631 ( .A(n6760), .Y(n5404) );
  NBUFFX2_HVT U6632 ( .A(n6760), .Y(n5405) );
  NBUFFX2_HVT U6633 ( .A(n6761), .Y(n5406) );
  NBUFFX2_HVT U6634 ( .A(n6761), .Y(n5407) );
  NBUFFX2_HVT U6635 ( .A(n10105), .Y(n5408) );
  NBUFFX2_HVT U6636 ( .A(n10105), .Y(n5409) );
  NBUFFX2_HVT U6637 ( .A(n6764), .Y(n5410) );
  NBUFFX2_HVT U6638 ( .A(n6764), .Y(n5411) );
  NBUFFX2_HVT U6639 ( .A(n10109), .Y(n5412) );
  NBUFFX2_HVT U6640 ( .A(n10109), .Y(n5413) );
  NBUFFX2_HVT U6641 ( .A(n10103), .Y(n5414) );
  NBUFFX2_HVT U6642 ( .A(n10103), .Y(n5415) );
  NBUFFX2_HVT U6643 ( .A(n10106), .Y(n5416) );
  NBUFFX2_HVT U6644 ( .A(n10106), .Y(n5417) );
  NBUFFX2_HVT U6645 ( .A(n10106), .Y(n5418) );
  NBUFFX2_HVT U6646 ( .A(n10109), .Y(n5419) );
  NBUFFX2_HVT U6647 ( .A(n10110), .Y(n5420) );
  NBUFFX2_HVT U6648 ( .A(n10110), .Y(n5421) );
  NBUFFX2_HVT U6649 ( .A(n10102), .Y(n5422) );
  NBUFFX2_HVT U6650 ( .A(n10102), .Y(n5423) );
  NBUFFX2_HVT U6651 ( .A(n10110), .Y(n5424) );
  NBUFFX2_HVT U6652 ( .A(n6893), .Y(n5425) );
  IBUFFX2_HVT U6653 ( .A(n10112), .Y(n10101) );
  INVX0_HVT U6654 ( .A(n5748), .Y(n6760) );
  INVX0_HVT U6655 ( .A(n5748), .Y(n6761) );
  INVX0_HVT U6656 ( .A(n7140), .Y(n6764) );
  INVX0_HVT U6657 ( .A(n7140), .Y(n10109) );
  INVX0_HVT U6658 ( .A(n7140), .Y(n10103) );
  INVX0_HVT U6659 ( .A(n7140), .Y(n10106) );
  IBUFFX2_HVT U6660 ( .A(n5749), .Y(n7140) );
  MUX41X1_HVT U6661 ( .A1(\ram[3][23] ), .A3(\ram[1][23] ), .A2(\ram[2][23] ), 
        .A4(\ram[0][23] ), .S0(n5426), .S1(n5883), .Y(n7827) );
  INVX0_HVT U6662 ( .A(n7267), .Y(n7713) );
  INVX0_HVT U6663 ( .A(n6160), .Y(n5461) );
  INVX0_HVT U6664 ( .A(n6165), .Y(n5489) );
  NBUFFX2_HVT U6665 ( .A(n7584), .Y(n8778) );
  INVX0_HVT U6666 ( .A(n7545), .Y(n7554) );
  INVX0_HVT U6667 ( .A(n6023), .Y(n7305) );
  INVX1_HVT U6668 ( .A(n6749), .Y(n6659) );
  INVX0_HVT U6669 ( .A(n7571), .Y(n5630) );
  INVX0_HVT U6670 ( .A(n7326), .Y(n5863) );
  INVX0_HVT U6671 ( .A(n6125), .Y(n5780) );
  INVX0_HVT U6672 ( .A(n6124), .Y(n5779) );
  INVX0_HVT U6673 ( .A(n4528), .Y(n6727) );
  INVX0_HVT U6674 ( .A(n22), .Y(n6158) );
  INVX0_HVT U6675 ( .A(n7965), .Y(n5472) );
  INVX0_HVT U6676 ( .A(n7964), .Y(n5473) );
  NBUFFX2_HVT U6677 ( .A(n5947), .Y(n6894) );
  INVX0_HVT U6678 ( .A(n5155), .Y(n7320) );
  INVX0_HVT U6679 ( .A(n5855), .Y(n8142) );
  INVX0_HVT U6680 ( .A(n8845), .Y(n5969) );
  INVX0_HVT U6681 ( .A(n7685), .Y(n7562) );
  INVX0_HVT U6682 ( .A(n5383), .Y(n5531) );
  INVX0_HVT U6683 ( .A(n10096), .Y(n10095) );
  INVX0_HVT U6684 ( .A(n8999), .Y(n5603) );
  INVX0_HVT U6685 ( .A(n21), .Y(n6012) );
  INVX0_HVT U6686 ( .A(n10205), .Y(n10204) );
  INVX0_HVT U6687 ( .A(n7150), .Y(n5853) );
  INVX0_HVT U6688 ( .A(n5625), .Y(n5655) );
  INVX0_HVT U6689 ( .A(n8825), .Y(n5527) );
  INVX0_HVT U6690 ( .A(n6491), .Y(n6485) );
  INVX0_HVT U6691 ( .A(n10328), .Y(n6262) );
  INVX0_HVT U6692 ( .A(n4718), .Y(n10287) );
  INVX0_HVT U6693 ( .A(n10128), .Y(n6969) );
  INVX0_HVT U6694 ( .A(n5896), .Y(n5809) );
  INVX0_HVT U6695 ( .A(n7581), .Y(n5496) );
  INVX0_HVT U6696 ( .A(n8764), .Y(n6399) );
  NBUFFX2_HVT U6697 ( .A(n5519), .Y(n6650) );
  INVX0_HVT U6698 ( .A(n7334), .Y(n5978) );
  IBUFFX2_HVT U6699 ( .A(n8771), .Y(n5757) );
  INVX0_HVT U6700 ( .A(n8820), .Y(n5772) );
  INVX1_HVT U6701 ( .A(n7693), .Y(n5864) );
  INVX0_HVT U6702 ( .A(n7352), .Y(n5776) );
  NBUFFX2_HVT U6703 ( .A(n5938), .Y(n8777) );
  INVX0_HVT U6704 ( .A(n7690), .Y(n7335) );
  INVX0_HVT U6705 ( .A(n5317), .Y(n5736) );
  NBUFFX2_HVT U6706 ( .A(n5938), .Y(n8770) );
  INVX0_HVT U6707 ( .A(n6133), .Y(n5750) );
  INVX0_HVT U6708 ( .A(n8753), .Y(n8762) );
  INVX0_HVT U6709 ( .A(n6416), .Y(n5623) );
  INVX0_HVT U6710 ( .A(n8773), .Y(n5959) );
  INVX0_HVT U6711 ( .A(n5364), .Y(n5756) );
  INVX0_HVT U6712 ( .A(n7352), .Y(n5637) );
  INVX0_HVT U6713 ( .A(n8850), .Y(n5821) );
  INVX0_HVT U6714 ( .A(n6658), .Y(n7570) );
  INVX0_HVT U6715 ( .A(n5877), .Y(n5827) );
  INVX0_HVT U6716 ( .A(n7562), .Y(n5891) );
  INVX0_HVT U6717 ( .A(n5990), .Y(n5799) );
  INVX0_HVT U6718 ( .A(n5969), .Y(n5657) );
  NBUFFX2_HVT U6719 ( .A(n5581), .Y(n8768) );
  INVX0_HVT U6720 ( .A(n6659), .Y(n5901) );
  NBUFFX2_HVT U6721 ( .A(n5581), .Y(n8772) );
  INVX1_HVT U6722 ( .A(n6661), .Y(n6397) );
  NBUFFX2_HVT U6723 ( .A(n7272), .Y(n8774) );
  INVX0_HVT U6724 ( .A(n5714), .Y(n8665) );
  INVX0_HVT U6725 ( .A(n5805), .Y(n5654) );
  INVX0_HVT U6726 ( .A(n5854), .Y(n5449) );
  INVX0_HVT U6727 ( .A(n8756), .Y(n5990) );
  INVX0_HVT U6728 ( .A(n5778), .Y(n8739) );
  INVX0_HVT U6729 ( .A(n8758), .Y(n6120) );
  INVX0_HVT U6730 ( .A(n5936), .Y(n10310) );
  INVX0_HVT U6731 ( .A(n7359), .Y(n10242) );
  INVX0_HVT U6732 ( .A(n8947), .Y(n8952) );
  INVX0_HVT U6733 ( .A(n8956), .Y(n8960) );
  INVX0_HVT U6734 ( .A(n5471), .Y(q[58]) );
  INVX0_HVT U6735 ( .A(n7963), .Y(n5474) );
  INVX0_HVT U6736 ( .A(n6415), .Y(n5575) );
  INVX0_HVT U6737 ( .A(n7068), .Y(n5481) );
  INVX0_HVT U6738 ( .A(n7200), .Y(n5467) );
  INVX0_HVT U6739 ( .A(n7189), .Y(n5442) );
  INVX0_HVT U6740 ( .A(n5848), .Y(n1646) );
  INVX0_HVT U6741 ( .A(n9199), .Y(n5849) );
  INVX0_HVT U6742 ( .A(n5845), .Y(n1648) );
  INVX0_HVT U6743 ( .A(n9197), .Y(n5846) );
  INVX0_HVT U6744 ( .A(n5843), .Y(n1650) );
  INVX0_HVT U6745 ( .A(n9214), .Y(n5841) );
  INVX0_HVT U6746 ( .A(n5494), .Y(n3525) );
  INVX1_HVT U6747 ( .A(n10065), .Y(n5596) );
  INVX0_HVT U6748 ( .A(n7673), .Y(n5592) );
  INVX0_HVT U6749 ( .A(n7293), .Y(n5805) );
  INVX0_HVT U6750 ( .A(n10252), .Y(n10250) );
  INVX0_HVT U6751 ( .A(n5613), .Y(n7293) );
  INVX0_HVT U6752 ( .A(n5613), .Y(n5625) );
  INVX0_HVT U6753 ( .A(n7570), .Y(n5925) );
  INVX0_HVT U6754 ( .A(n4545), .Y(n7379) );
  INVX0_HVT U6755 ( .A(n6751), .Y(n5774) );
  INVX0_HVT U6756 ( .A(n5881), .Y(n5538) );
  INVX1_HVT U6757 ( .A(n7288), .Y(n5808) );
  INVX0_HVT U6758 ( .A(n6641), .Y(n5791) );
  INVX0_HVT U6759 ( .A(n6416), .Y(n5831) );
  INVX0_HVT U6760 ( .A(n5953), .Y(n7348) );
  INVX0_HVT U6761 ( .A(n5931), .Y(n5806) );
  INVX0_HVT U6762 ( .A(n4912), .Y(n7672) );
  INVX0_HVT U6763 ( .A(n9014), .Y(n9016) );
  INVX1_HVT U6764 ( .A(n5898), .Y(n5755) );
  INVX0_HVT U6765 ( .A(n9258), .Y(n5782) );
  INVX0_HVT U6766 ( .A(n8759), .Y(n5886) );
  INVX0_HVT U6767 ( .A(n7723), .Y(n10347) );
  INVX0_HVT U6768 ( .A(n9227), .Y(n5533) );
  INVX0_HVT U6769 ( .A(n6069), .Y(n10230) );
  INVX0_HVT U6770 ( .A(n6069), .Y(n10231) );
  INVX0_HVT U6771 ( .A(n10116), .Y(n10115) );
  INVX1_HVT U6772 ( .A(n56), .Y(n10116) );
  INVX0_HVT U6773 ( .A(n9000), .Y(n6015) );
  INVX0_HVT U6774 ( .A(n5681), .Y(n5688) );
  INVX0_HVT U6775 ( .A(n8911), .Y(n8957) );
  INVX0_HVT U6776 ( .A(n8957), .Y(n8965) );
  INVX0_HVT U6777 ( .A(n8947), .Y(n8949) );
  INVX0_HVT U6778 ( .A(n7566), .Y(n7301) );
  INVX1_HVT U6779 ( .A(n7309), .Y(n5503) );
  INVX0_HVT U6780 ( .A(n7733), .Y(n10269) );
  INVX0_HVT U6781 ( .A(n10256), .Y(n10255) );
  INVX0_HVT U6782 ( .A(n6659), .Y(n7548) );
  INVX0_HVT U6783 ( .A(n5954), .Y(n5916) );
  INVX0_HVT U6784 ( .A(n5913), .Y(n5915) );
  INVX0_HVT U6785 ( .A(n4956), .Y(n7236) );
  INVX0_HVT U6786 ( .A(n7724), .Y(n10330) );
  INVX0_HVT U6787 ( .A(n7720), .Y(n10361) );
  INVX0_HVT U6788 ( .A(n10116), .Y(n9025) );
  INVX0_HVT U6789 ( .A(n10116), .Y(n9024) );
  INVX0_HVT U6790 ( .A(n8997), .Y(n5520) );
  INVX0_HVT U6791 ( .A(n10206), .Y(n10205) );
  INVX0_HVT U6792 ( .A(n6003), .Y(n6733) );
  INVX0_HVT U6793 ( .A(n7665), .Y(n5450) );
  INVX0_HVT U6794 ( .A(n9166), .Y(n9154) );
  INVX0_HVT U6795 ( .A(n9165), .Y(n9153) );
  INVX0_HVT U6796 ( .A(n9257), .Y(n7269) );
  INVX0_HVT U6797 ( .A(n10096), .Y(n10094) );
  INVX0_HVT U6798 ( .A(n10099), .Y(n5913) );
  INVX0_HVT U6799 ( .A(n7583), .Y(n6642) );
  INVX1_HVT U6800 ( .A(n10205), .Y(n10203) );
  INVX0_HVT U6801 ( .A(n5291), .Y(n5737) );
  INVX0_HVT U6802 ( .A(n4424), .Y(n9254) );
  INVX0_HVT U6803 ( .A(n10273), .Y(n10272) );
  INVX0_HVT U6804 ( .A(n9111), .Y(n9083) );
  INVX0_HVT U6805 ( .A(n6651), .Y(n6130) );
  INVX1_HVT U6806 ( .A(n5873), .Y(n5904) );
  INVX0_HVT U6807 ( .A(n10289), .Y(n9274) );
  INVX0_HVT U6808 ( .A(n10289), .Y(n9268) );
  INVX0_HVT U6809 ( .A(n6423), .Y(n10182) );
  INVX0_HVT U6810 ( .A(n10254), .Y(n9159) );
  INVX0_HVT U6811 ( .A(n10253), .Y(n9148) );
  INVX0_HVT U6812 ( .A(n10253), .Y(n9147) );
  INVX0_HVT U6813 ( .A(n10114), .Y(n9041) );
  INVX0_HVT U6814 ( .A(n10113), .Y(n9047) );
  INVX0_HVT U6815 ( .A(n10114), .Y(n9035) );
  INVX0_HVT U6816 ( .A(n5954), .Y(n10099) );
  INVX0_HVT U6817 ( .A(n5909), .Y(n5911) );
  INVX0_HVT U6818 ( .A(n5909), .Y(n5912) );
  INVX0_HVT U6819 ( .A(n6036), .Y(n5544) );
  INVX0_HVT U6820 ( .A(n6735), .Y(n5490) );
  INVX0_HVT U6821 ( .A(n10304), .Y(n6178) );
  INVX0_HVT U6822 ( .A(n10204), .Y(n9092) );
  INVX0_HVT U6823 ( .A(n10203), .Y(n9104) );
  INVX0_HVT U6824 ( .A(n10203), .Y(n9093) );
  INVX0_HVT U6825 ( .A(n10123), .Y(n8921) );
  INVX0_HVT U6826 ( .A(n6651), .Y(n5815) );
  INVX0_HVT U6827 ( .A(n10288), .Y(n9263) );
  INVX0_HVT U6828 ( .A(n10288), .Y(n9269) );
  INVX0_HVT U6829 ( .A(n8773), .Y(n7299) );
  INVX0_HVT U6830 ( .A(n5487), .Y(n5478) );
  INVX0_HVT U6831 ( .A(n4791), .Y(n10131) );
  INVX0_HVT U6832 ( .A(n4791), .Y(n10132) );
  INVX0_HVT U6833 ( .A(n4956), .Y(n10118) );
  INVX0_HVT U6834 ( .A(n10120), .Y(n10119) );
  INVX0_HVT U6835 ( .A(n10190), .Y(n6423) );
  INVX0_HVT U6836 ( .A(n10271), .Y(n9206) );
  INVX0_HVT U6837 ( .A(n10270), .Y(n9217) );
  INVX0_HVT U6838 ( .A(n9224), .Y(n9205) );
  INVX0_HVT U6839 ( .A(n4355), .Y(n10316) );
  INVX0_HVT U6840 ( .A(n4355), .Y(n10318) );
  INVX0_HVT U6841 ( .A(n6037), .Y(n5802) );
  OAI22X1_HVT U6842 ( .A1(n7270), .A2(n5667), .A3(n7269), .A4(n9450), .Y(n5427) );
  OAI22X1_HVT U6843 ( .A1(n5876), .A2(n5665), .A3(n7269), .A4(n9456), .Y(n5428) );
  OAI22X1_HVT U6844 ( .A1(n6631), .A2(n5173), .A3(n5533), .A4(n9930), .Y(n5429) );
  OAI22X1_HVT U6845 ( .A1(n5963), .A2(n5664), .A3(n9287), .A4(n9666), .Y(n5430) );
  OAI22X1_HVT U6846 ( .A1(n6553), .A2(n5666), .A3(n5782), .A4(n9367), .Y(n5431) );
  OAI22X1_HVT U6847 ( .A1(n5872), .A2(n5667), .A3(n5782), .A4(n9314), .Y(n5432) );
  OAI22X1_HVT U6848 ( .A1(n5783), .A2(n5665), .A3(n5782), .A4(n9355), .Y(n5433) );
  OAI22X1_HVT U6849 ( .A1(n5781), .A2(n5666), .A3(n5782), .A4(n9361), .Y(n5434) );
  OAI22X1_HVT U6850 ( .A1(n5952), .A2(n5664), .A3(n5951), .A4(n9672), .Y(n5435) );
  INVX0_HVT U6851 ( .A(n7729), .Y(n10149) );
  INVX0_HVT U6852 ( .A(n7726), .Y(n10252) );
  INVX0_HVT U6853 ( .A(n7728), .Y(n10202) );
  INVX0_HVT U6854 ( .A(n7721), .Y(n10236) );
  INVX0_HVT U6855 ( .A(n7725), .Y(n10303) );
  INVX0_HVT U6856 ( .A(n6191), .Y(n5451) );
  INVX0_HVT U6857 ( .A(n10134), .Y(n6336) );
  INVX0_HVT U6858 ( .A(n55), .Y(n10121) );
  INVX0_HVT U6859 ( .A(n10121), .Y(n7213) );
  INVX0_HVT U6860 ( .A(n7574), .Y(n7310) );
  INVX0_HVT U6861 ( .A(n5991), .Y(n5801) );
  INVX0_HVT U6862 ( .A(n10290), .Y(n10288) );
  INVX0_HVT U6863 ( .A(n10290), .Y(n10289) );
  INVX0_HVT U6864 ( .A(n10115), .Y(n10114) );
  INVX0_HVT U6865 ( .A(n5531), .Y(n10100) );
  INVX0_HVT U6866 ( .A(n10097), .Y(n8972) );
  NBUFFX2_HVT U6867 ( .A(n6763), .Y(n5441) );
  INVX0_HVT U6868 ( .A(n6025), .Y(n20) );
  OAI22X1_HVT U6869 ( .A1(n5443), .A2(n5442), .A3(n6276), .A4(n10080), .Y(n825) );
  INVX0_HVT U6870 ( .A(n6373), .Y(n6376) );
  INVX0_HVT U6871 ( .A(n6373), .Y(n6375) );
  INVX0_HVT U6872 ( .A(n6364), .Y(n6369) );
  INVX0_HVT U6873 ( .A(n6364), .Y(n6368) );
  INVX0_HVT U6874 ( .A(n6364), .Y(n6366) );
  INVX0_HVT U6875 ( .A(n6365), .Y(n6372) );
  INVX0_HVT U6876 ( .A(n6365), .Y(n6370) );
  INVX0_HVT U6877 ( .A(n5608), .Y(n8837) );
  INVX0_HVT U6878 ( .A(n5456), .Y(n5444) );
  INVX0_HVT U6879 ( .A(n7559), .Y(n5456) );
  NBUFFX2_HVT U6880 ( .A(n6171), .Y(n5445) );
  IBUFFX2_HVT U6881 ( .A(n6166), .Y(n6172) );
  OAI22X1_HVT U6882 ( .A1(n5477), .A2(n6713), .A3(n9740), .A4(n6498), .Y(n205)
         );
  INVX0_HVT U6883 ( .A(n6374), .Y(n6380) );
  INVX0_HVT U6884 ( .A(n6374), .Y(n6379) );
  INVX0_HVT U6885 ( .A(n5450), .Y(n5446) );
  INVX0_HVT U6886 ( .A(n6373), .Y(n6377) );
  INVX0_HVT U6887 ( .A(n6364), .Y(n6367) );
  INVX0_HVT U6888 ( .A(n6365), .Y(n6371) );
  INVX0_HVT U6889 ( .A(n6374), .Y(n6378) );
  NBUFFX2_HVT U6890 ( .A(n7690), .Y(n5448) );
  IBUFFX2_HVT U6891 ( .A(n7685), .Y(n6661) );
  INVX0_HVT U6892 ( .A(n8910), .Y(n8947) );
  INVX0_HVT U6893 ( .A(n6165), .Y(n6169) );
  MUX41X1_HVT U6894 ( .A1(\ram[3][243] ), .A3(\ram[1][243] ), .A2(
        \ram[2][243] ), .A4(\ram[0][243] ), .S0(n5449), .S1(n5450), .Y(n8702)
         );
  INVX0_HVT U6895 ( .A(n5062), .Y(n6177) );
  INVX0_HVT U6896 ( .A(n6165), .Y(n6170) );
  OAI22X1_HVT U6897 ( .A1(n5452), .A2(n4762), .A3(n5451), .A4(n9393), .Y(n1114) );
  OAI22X1_HVT U6898 ( .A1(n5453), .A2(n6175), .A3(n6235), .A4(n9958), .Y(n1298) );
  INVX0_HVT U6899 ( .A(n6735), .Y(n6176) );
  INVX0_HVT U6900 ( .A(n5879), .Y(n5880) );
  INVX0_HVT U6901 ( .A(n8910), .Y(n8948) );
  INVX0_HVT U6902 ( .A(n8939), .Y(n5455) );
  INVX0_HVT U6903 ( .A(n5837), .Y(n8181) );
  MUX41X1_HVT U6904 ( .A1(\ram[7][19] ), .A3(\ram[5][19] ), .A2(\ram[6][19] ), 
        .A4(\ram[4][19] ), .S0(n5738), .S1(n5628), .Y(n7812) );
  IBUFFX2_HVT U6905 ( .A(n6391), .Y(n5734) );
  INVX0_HVT U6906 ( .A(n10361), .Y(n6491) );
  MUX41X1_HVT U6907 ( .A1(\ram[7][192] ), .A3(\ram[5][192] ), .A2(
        \ram[6][192] ), .A4(\ram[4][192] ), .S0(n5201), .S1(n43), .Y(n8499) );
  INVX0_HVT U6908 ( .A(n4327), .Y(n6826) );
  INVX0_HVT U6909 ( .A(n5465), .Y(n5458) );
  INVX0_HVT U6910 ( .A(n8881), .Y(n5465) );
  INVX0_HVT U6911 ( .A(n5459), .Y(n5460) );
  INVX0_HVT U6912 ( .A(n6401), .Y(n7765) );
  INVX0_HVT U6913 ( .A(n5704), .Y(n5664) );
  OAI22X1_HVT U6914 ( .A1(n5861), .A2(n5860), .A3(n5284), .A4(n9898), .Y(n5462) );
  INVX0_HVT U6915 ( .A(n5704), .Y(n5667) );
  MUX41X1_HVT U6916 ( .A1(\ram[3][43] ), .A3(\ram[1][43] ), .A2(\ram[2][43] ), 
        .A4(\ram[0][43] ), .S0(n5878), .S1(n5813), .Y(n7906) );
  INVX0_HVT U6917 ( .A(n5469), .Y(n5463) );
  INVX0_HVT U6918 ( .A(n5762), .Y(n10278) );
  OAI22X1_HVT U6919 ( .A1(n5464), .A2(n5762), .A3(n5533), .A4(n9660), .Y(n1715) );
  IBUFFX2_HVT U6920 ( .A(n9243), .Y(n9249) );
  IBUFFX2_HVT U6921 ( .A(n10126), .Y(n8916) );
  MUX41X1_HVT U6922 ( .A1(\ram[15][67] ), .A3(\ram[13][67] ), .A2(
        \ram[14][67] ), .A4(\ram[12][67] ), .S0(n7556), .S1(n5465), .Y(n7998)
         );
  AO22X1_HVT U6923 ( .A1(\ram[3][48] ), .A2(n7132), .A3(n5273), .A4(n9451), 
        .Y(n5466) );
  INVX0_HVT U6924 ( .A(n6282), .Y(n6284) );
  MUX41X1_HVT U6925 ( .A1(\ram[3][135] ), .A3(\ram[1][135] ), .A2(
        \ram[2][135] ), .A4(\ram[0][135] ), .S0(n6654), .S1(n5469), .Y(n8273)
         );
  IBUFFX2_HVT U6926 ( .A(n8867), .Y(n7143) );
  IBUFFX2_HVT U6927 ( .A(n8948), .Y(n8954) );
  IBUFFX2_HVT U6928 ( .A(n7187), .Y(n7190) );
  MUX41X1_HVT U6929 ( .A1(n5474), .A3(n5473), .A2(n4814), .A4(n5472), .S0(
        n5736), .S1(n5904), .Y(n5471) );
  MUX41X1_HVT U6930 ( .A1(\ram[11][57] ), .A3(\ram[9][57] ), .A2(\ram[10][57] ), .A4(\ram[8][57] ), .S0(n7281), .S1(n5133), .Y(n7960) );
  INVX0_HVT U6931 ( .A(n10236), .Y(n6043) );
  INVX0_HVT U6932 ( .A(n10236), .Y(n6044) );
  INVX1_HVT U6933 ( .A(n6654), .Y(n5475) );
  INVX0_HVT U6934 ( .A(n5825), .Y(n6387) );
  INVX0_HVT U6935 ( .A(n7142), .Y(n5476) );
  INVX0_HVT U6936 ( .A(n7133), .Y(n5860) );
  INVX0_HVT U6937 ( .A(n7322), .Y(n7142) );
  MUX41X1_HVT U6938 ( .A1(\ram[10][105] ), .A3(\ram[8][105] ), .A2(
        \ram[11][105] ), .A4(\ram[9][105] ), .S0(n4986), .S1(n5812), .Y(n8151)
         );
  INVX0_HVT U6939 ( .A(n8956), .Y(n8961) );
  INVX0_HVT U6940 ( .A(n8956), .Y(n8959) );
  INVX0_HVT U6941 ( .A(n7063), .Y(n5480) );
  OAI22X1_HVT U6942 ( .A1(n5482), .A2(n5481), .A3(n6826), .A4(n9570), .Y(n405)
         );
  INVX0_HVT U6943 ( .A(n10346), .Y(n6827) );
  INVX0_HVT U6944 ( .A(n7073), .Y(n5483) );
  MUX41X1_HVT U6945 ( .A1(\ram[15][118] ), .A3(\ram[13][118] ), .A2(
        \ram[14][118] ), .A4(\ram[12][118] ), .S0(n5640), .S1(n5485), .Y(n8202) );
  MUX41X1_HVT U6946 ( .A1(\ram[15][88] ), .A3(\ram[13][88] ), .A2(
        \ram[14][88] ), .A4(\ram[12][88] ), .S0(n5803), .S1(n5485), .Y(n8082)
         );
  INVX0_HVT U6947 ( .A(n8956), .Y(n8958) );
  MUX41X1_HVT U6948 ( .A1(\ram[11][225] ), .A3(\ram[9][225] ), .A2(
        \ram[10][225] ), .A4(\ram[8][225] ), .S0(n5787), .S1(n5337), .Y(n8630)
         );
  INVX0_HVT U6949 ( .A(n7325), .Y(n5787) );
  MUX41X1_HVT U6950 ( .A1(\ram[11][245] ), .A3(\ram[9][245] ), .A2(
        \ram[10][245] ), .A4(\ram[8][245] ), .S0(n5884), .S1(n5893), .Y(n8708)
         );
  INVX0_HVT U6951 ( .A(n10221), .Y(n7586) );
  INVX0_HVT U6952 ( .A(n5689), .Y(n5666) );
  INVX0_HVT U6953 ( .A(n8957), .Y(n8964) );
  INVX0_HVT U6954 ( .A(n8957), .Y(n8962) );
  INVX0_HVT U6955 ( .A(n8957), .Y(n8963) );
  INVX0_HVT U6956 ( .A(n8947), .Y(n8951) );
  INVX0_HVT U6957 ( .A(n8947), .Y(n8950) );
  INVX0_HVT U6958 ( .A(n8948), .Y(n8955) );
  INVX0_HVT U6959 ( .A(n8948), .Y(n8953) );
  MUX41X1_HVT U6960 ( .A1(\ram[7][216] ), .A3(\ram[5][216] ), .A2(
        \ram[6][216] ), .A4(\ram[4][216] ), .S0(n5234), .S1(n5486), .Y(n8595)
         );
  MUX41X1_HVT U6961 ( .A1(\ram[11][8] ), .A3(\ram[9][8] ), .A2(\ram[10][8] ), 
        .A4(\ram[8][8] ), .S0(n5814), .S1(n5488), .Y(n7767) );
  INVX0_HVT U6962 ( .A(n6023), .Y(n5814) );
  IBUFFX2_HVT U6963 ( .A(n7064), .Y(n7071) );
  INVX0_HVT U6964 ( .A(n5646), .Y(n6654) );
  MUX41X1_HVT U6965 ( .A1(\ram[7][85] ), .A3(\ram[5][85] ), .A2(\ram[6][85] ), 
        .A4(\ram[4][85] ), .S0(n6136), .S1(n5775), .Y(n8072) );
  INVX0_HVT U6966 ( .A(n7188), .Y(n7196) );
  INVX0_HVT U6967 ( .A(n7188), .Y(n7194) );
  INVX0_HVT U6968 ( .A(n4582), .Y(n7193) );
  INVX0_HVT U6969 ( .A(n7187), .Y(n7192) );
  INVX0_HVT U6970 ( .A(n7187), .Y(n7191) );
  INVX0_HVT U6971 ( .A(n7187), .Y(n7189) );
  MUX41X1_HVT U6972 ( .A1(\ram[14][82] ), .A3(\ram[12][82] ), .A2(
        \ram[15][82] ), .A4(\ram[13][82] ), .S0(n5638), .S1(n5512), .Y(n8058)
         );
  MUX41X1_HVT U6973 ( .A1(n8054), .A3(n8055), .A2(n8056), .A4(n8057), .S0(
        n5648), .S1(n5655), .Y(q[81]) );
  INVX0_HVT U6974 ( .A(n7282), .Y(n5491) );
  INVX0_HVT U6975 ( .A(n5493), .Y(n5492) );
  INVX0_HVT U6976 ( .A(n8881), .Y(n5493) );
  MUX41X1_HVT U6977 ( .A1(\ram[1][3] ), .A3(\ram[3][3] ), .A2(\ram[0][3] ), 
        .A4(\ram[2][3] ), .S0(n5122), .S1(n7148), .Y(n7749) );
  MUX41X1_HVT U6978 ( .A1(\ram[3][52] ), .A3(\ram[1][52] ), .A2(\ram[2][52] ), 
        .A4(\ram[0][52] ), .S0(n5602), .S1(n5493), .Y(n7942) );
  AOI21X1_HVT U6979 ( .A1(n54), .A2(n10375), .A3(rst), .Y(n52) );
  INVX0_HVT U6980 ( .A(n5833), .Y(n5723) );
  INVX0_HVT U6981 ( .A(n8754), .Y(n5833) );
  OA22X1_HVT U6982 ( .A1(n5495), .A2(n4601), .A3(n8938), .A4(n9714), .Y(n5494)
         );
  IBUFFX2_HVT U6983 ( .A(n7007), .Y(n7012) );
  MUX41X1_HVT U6984 ( .A1(\ram[3][8] ), .A3(\ram[1][8] ), .A2(\ram[2][8] ), 
        .A4(\ram[0][8] ), .S0(n7281), .S1(n5496), .Y(n7769) );
  OAI22X1_HVT U6985 ( .A1(n5497), .A2(n5173), .A3(n5533), .A4(n9970), .Y(n1814) );
  OAI22X1_HVT U6986 ( .A1(n5498), .A2(n5378), .A3(n5520), .A4(n9531), .Y(n3976) );
  IBUFFX2_HVT U6987 ( .A(n9004), .Y(n9007) );
  INVX0_HVT U6988 ( .A(n5696), .Y(n5665) );
  NBUFFX2_HVT U6989 ( .A(n5661), .Y(n5499) );
  NBUFFX2_HVT U6990 ( .A(n7564), .Y(n5500) );
  INVX0_HVT U6991 ( .A(n4972), .Y(n5514) );
  MUX41X1_HVT U6992 ( .A1(n7982), .A3(n7984), .A2(n7983), .A4(n7985), .S0(
        n7349), .S1(n5503), .Y(q[63]) );
  INVX0_HVT U6993 ( .A(n7063), .Y(n7067) );
  INVX0_HVT U6994 ( .A(n7063), .Y(n7066) );
  INVX0_HVT U6995 ( .A(n7063), .Y(n7065) );
  INVX0_HVT U6996 ( .A(n7073), .Y(n7077) );
  INVX0_HVT U6997 ( .A(n7073), .Y(n7076) );
  INVX0_HVT U6998 ( .A(n7073), .Y(n7075) );
  INVX0_HVT U6999 ( .A(n7064), .Y(n7072) );
  INVX0_HVT U7000 ( .A(n7064), .Y(n7070) );
  INVX0_HVT U7001 ( .A(n7064), .Y(n7069) );
  NBUFFX2_HVT U7002 ( .A(n6892), .Y(n8898) );
  INVX0_HVT U7003 ( .A(n7569), .Y(n5510) );
  INVX0_HVT U7004 ( .A(n5525), .Y(n6630) );
  MUX41X1_HVT U7005 ( .A1(n8171), .A3(n8173), .A2(n8170), .A4(n8172), .S0(
        n5830), .S1(n5926), .Y(q[110]) );
  IBUFFX2_HVT U7006 ( .A(n7006), .Y(n7010) );
  INVX0_HVT U7007 ( .A(n7553), .Y(n5507) );
  MUX41X1_HVT U7008 ( .A1(\ram[13][166] ), .A3(\ram[15][166] ), .A2(
        \ram[12][166] ), .A4(\ram[14][166] ), .S0(n4985), .S1(n5049), .Y(n8393) );
  INVX0_HVT U7009 ( .A(n7690), .Y(n8799) );
  MUX41X1_HVT U7010 ( .A1(\ram[15][56] ), .A3(\ram[13][56] ), .A2(
        \ram[14][56] ), .A4(\ram[12][56] ), .S0(n5507), .S1(n5508), .Y(n7955)
         );
  INVX0_HVT U7011 ( .A(n5555), .Y(n5509) );
  INVX0_HVT U7012 ( .A(n7264), .Y(n5555) );
  IBUFFX2_HVT U7013 ( .A(n10125), .Y(n10122) );
  MUX41X1_HVT U7014 ( .A1(\ram[7][103] ), .A3(\ram[5][103] ), .A2(
        \ram[6][103] ), .A4(\ram[4][103] ), .S0(n5647), .S1(n5510), .Y(n8144)
         );
  INVX1_HVT U7015 ( .A(n5879), .Y(n5511) );
  MUX41X1_HVT U7016 ( .A1(\ram[3][74] ), .A3(\ram[1][74] ), .A2(\ram[2][74] ), 
        .A4(\ram[0][74] ), .S0(n5937), .S1(n5232), .Y(n8029) );
  INVX0_HVT U7017 ( .A(n5762), .Y(n10281) );
  IBUFFX2_HVT U7018 ( .A(n5761), .Y(n5513) );
  MUX41X1_HVT U7019 ( .A1(\ram[3][70] ), .A3(\ram[1][70] ), .A2(\ram[2][70] ), 
        .A4(\ram[0][70] ), .S0(n5998), .S1(n5826), .Y(n8013) );
  INVX0_HVT U7020 ( .A(n10287), .Y(n5516) );
  INVX0_HVT U7021 ( .A(n5761), .Y(n5517) );
  INVX0_HVT U7022 ( .A(n5518), .Y(n5519) );
  MUX41X1_HVT U7023 ( .A1(n7899), .A3(n7901), .A2(n7900), .A4(n7902), .S0(
        n5305), .S1(n6398), .Y(q[42]) );
  OAI22X1_HVT U7024 ( .A1(n5521), .A2(n5531), .A3(n5520), .A4(n9396), .Y(n3931) );
  OAI22X1_HVT U7025 ( .A1(n5522), .A2(n5540), .A3(n6015), .A4(n9555), .Y(n3984) );
  INVX0_HVT U7026 ( .A(n10252), .Y(n7353) );
  INVX0_HVT U7027 ( .A(n5627), .Y(n5523) );
  INVX0_HVT U7028 ( .A(n6008), .Y(n5627) );
  AO21X1_HVT U7029 ( .A1(n7), .A2(n6258), .A3(n10381), .Y(n7730) );
  IBUFFX2_HVT U7030 ( .A(n7291), .Y(n6009) );
  INVX0_HVT U7031 ( .A(n8806), .Y(n5941) );
  INVX0_HVT U7032 ( .A(n8806), .Y(n6128) );
  MUX41X1_HVT U7033 ( .A1(\ram[2][249] ), .A3(\ram[0][249] ), .A2(
        \ram[3][249] ), .A4(\ram[1][249] ), .S0(n5507), .S1(n5573), .Y(n8726)
         );
  MUX41X1_HVT U7034 ( .A1(\ram[11][54] ), .A3(\ram[9][54] ), .A2(\ram[10][54] ), .A4(\ram[8][54] ), .S0(n5772), .S1(n5456), .Y(n7948) );
  INVX0_HVT U7035 ( .A(n8845), .Y(n5605) );
  MUX41X1_HVT U7036 ( .A1(n7738), .A3(n7740), .A2(n7739), .A4(n7741), .S0(
        n7276), .S1(n5904), .Y(q[1]) );
  OAI22X1_HVT U7037 ( .A1(n5524), .A2(n5379), .A3(n6015), .A4(n9387), .Y(n3928) );
  MUX41X1_HVT U7038 ( .A1(n8174), .A3(n8176), .A2(n8175), .A4(n8177), .S0(
        n5886), .S1(n5332), .Y(q[111]) );
  MUX41X1_HVT U7039 ( .A1(n8234), .A3(n8236), .A2(n8235), .A4(n8237), .S0(
        n7570), .S1(n5959), .Y(q[126]) );
  INVX0_HVT U7040 ( .A(n8839), .Y(n7673) );
  MUX41X1_HVT U7041 ( .A1(\ram[14][92] ), .A3(\ram[12][92] ), .A2(
        \ram[15][92] ), .A4(\ram[13][92] ), .S0(n5574), .S1(n7667), .Y(n8098)
         );
  MUX41X1_HVT U7042 ( .A1(\ram[3][248] ), .A3(\ram[1][248] ), .A2(
        \ram[2][248] ), .A4(\ram[0][248] ), .S0(n5527), .S1(n5300), .Y(n8722)
         );
  INVX0_HVT U7043 ( .A(n7150), .Y(n6892) );
  OAI22X1_HVT U7044 ( .A1(n5529), .A2(n5381), .A3(n5520), .A4(n9343), .Y(n3913) );
  IBUFFX2_HVT U7045 ( .A(n9005), .Y(n9013) );
  OAI22X1_HVT U7046 ( .A1(n5530), .A2(n5378), .A3(n5520), .A4(n9765), .Y(n4053) );
  OAI22X1_HVT U7047 ( .A1(n5856), .A2(n5380), .A3(n5603), .A4(n9615), .Y(n4004) );
  IBUFFX2_HVT U7048 ( .A(n9005), .Y(n9010) );
  INVX0_HVT U7049 ( .A(n6626), .Y(n5558) );
  MUX41X1_HVT U7050 ( .A1(\ram[3][132] ), .A3(\ram[1][132] ), .A2(
        \ram[2][132] ), .A4(\ram[0][132] ), .S0(n5571), .S1(n5818), .Y(n8261)
         );
  MUX41X1_HVT U7051 ( .A1(n7747), .A3(n7749), .A2(n7746), .A4(n7748), .S0(
        n6399), .S1(n5536), .Y(q[3]) );
  INVX0_HVT U7052 ( .A(n5566), .Y(n5659) );
  MUX41X1_HVT U7053 ( .A1(n7862), .A3(n7860), .A2(n7861), .A4(n7859), .S0(
        n5756), .S1(n5136), .Y(q[32]) );
  MUX41X1_HVT U7054 ( .A1(\ram[11][59] ), .A3(\ram[9][59] ), .A2(\ram[10][59] ), .A4(\ram[8][59] ), .S0(n5140), .S1(n5607), .Y(n7967) );
  MUX41X1_HVT U7055 ( .A1(n7770), .A3(n7772), .A2(n7771), .A4(n7773), .S0(
        n6399), .S1(n5809), .Y(q[9]) );
  MUX41X1_HVT U7056 ( .A1(\ram[11][173] ), .A3(\ram[9][173] ), .A2(
        \ram[10][173] ), .A4(\ram[8][173] ), .S0(n5571), .S1(n5628), .Y(n8422)
         );
  OAI22X1_HVT U7057 ( .A1(n5534), .A2(n5762), .A3(n5533), .A4(n9321), .Y(n1602) );
  NBUFFX2_HVT U7058 ( .A(n7674), .Y(n5535) );
  INVX0_HVT U7059 ( .A(n4829), .Y(n7015) );
  INVX0_HVT U7060 ( .A(n7006), .Y(n7014) );
  INVX0_HVT U7061 ( .A(n7007), .Y(n7013) );
  INVX0_HVT U7062 ( .A(n7016), .Y(n7020) );
  INVX0_HVT U7063 ( .A(n7016), .Y(n7019) );
  INVX0_HVT U7064 ( .A(n5009), .Y(n9279) );
  INVX0_HVT U7065 ( .A(n5009), .Y(n9280) );
  INVX0_HVT U7066 ( .A(n5571), .Y(n5537) );
  INVX0_HVT U7067 ( .A(n2), .Y(n5571) );
  MUX41X1_HVT U7068 ( .A1(\ram[15][173] ), .A3(\ram[13][173] ), .A2(
        \ram[14][173] ), .A4(\ram[12][173] ), .S0(n5894), .S1(n5739), .Y(n8421) );
  INVX0_HVT U7069 ( .A(n5348), .Y(n10315) );
  MUX41X1_HVT U7070 ( .A1(\ram[11][240] ), .A3(\ram[9][240] ), .A2(
        \ram[10][240] ), .A4(\ram[8][240] ), .S0(n7277), .S1(n7149), .Y(n8688)
         );
  AOI21X1_HVT U7071 ( .A1(n24), .A2(n10376), .A3(n10381), .Y(n22) );
  INVX0_HVT U7072 ( .A(n5541), .Y(n5539) );
  MUX41X1_HVT U7073 ( .A1(\ram[11][158] ), .A3(\ram[9][158] ), .A2(
        \ram[10][158] ), .A4(\ram[8][158] ), .S0(n5743), .S1(n7143), .Y(n8362)
         );
  IBUFFX2_HVT U7074 ( .A(n5236), .Y(n7679) );
  INVX0_HVT U7075 ( .A(n5600), .Y(n5540) );
  NBUFFX2_HVT U7076 ( .A(n5797), .Y(n8893) );
  MUX41X1_HVT U7077 ( .A1(\ram[15][183] ), .A3(\ram[13][183] ), .A2(
        \ram[14][183] ), .A4(\ram[12][183] ), .S0(n5527), .S1(n5541), .Y(n8461) );
  INVX0_HVT U7078 ( .A(n6408), .Y(n5542) );
  INVX0_HVT U7079 ( .A(n5542), .Y(n5543) );
  IBUFFX2_HVT U7080 ( .A(n5566), .Y(n7667) );
  INVX0_HVT U7081 ( .A(n7683), .Y(n5556) );
  MUX41X1_HVT U7082 ( .A1(\ram[7][194] ), .A3(\ram[5][194] ), .A2(
        \ram[6][194] ), .A4(\ram[4][194] ), .S0(n7265), .S1(n5715), .Y(n8507)
         );
  MUX41X1_HVT U7083 ( .A1(\ram[7][87] ), .A3(\ram[5][87] ), .A2(\ram[6][87] ), 
        .A4(\ram[4][87] ), .S0(n7313), .S1(n5986), .Y(n8080) );
  INVX0_HVT U7084 ( .A(n10286), .Y(n5545) );
  INVX0_HVT U7085 ( .A(n10287), .Y(n5546) );
  INVX0_HVT U7086 ( .A(n5761), .Y(n10285) );
  INVX0_HVT U7087 ( .A(n10306), .Y(n6145) );
  OAI22X1_HVT U7088 ( .A1(n5547), .A2(n5061), .A3(n6232), .A4(n9432), .Y(n1127) );
  OAI22X1_HVT U7089 ( .A1(n5548), .A2(n6175), .A3(n6199), .A4(n9414), .Y(n1121) );
  INVX0_HVT U7090 ( .A(n5451), .Y(n6202) );
  OAI22X1_HVT U7091 ( .A1(n5549), .A2(n5061), .A3(n6247), .A4(n9387), .Y(n1112) );
  OAI22X1_HVT U7092 ( .A1(n5550), .A2(n6735), .A3(n6199), .A4(n9381), .Y(n1110) );
  NBUFFX2_HVT U7093 ( .A(n8884), .Y(n5551) );
  INVX0_HVT U7094 ( .A(n5552), .Y(n5553) );
  NBUFFX2_HVT U7095 ( .A(n8893), .Y(n5554) );
  MUX41X1_HVT U7096 ( .A1(n8099), .A3(n8101), .A2(n8098), .A4(n8100), .S0(
        n5720), .S1(n7280), .Y(q[92]) );
  MUX41X1_HVT U7097 ( .A1(\ram[7][84] ), .A3(\ram[5][84] ), .A2(\ram[6][84] ), 
        .A4(\ram[4][84] ), .S0(n6128), .S1(n7348), .Y(n8068) );
  IBUFFX2_HVT U7098 ( .A(n7297), .Y(n8842) );
  INVX1_HVT U7099 ( .A(n8328), .Y(n6633) );
  MUX41X1_HVT U7100 ( .A1(\ram[15][64] ), .A3(\ram[13][64] ), .A2(
        \ram[14][64] ), .A4(\ram[12][64] ), .S0(n5555), .S1(n5556), .Y(n7986)
         );
  INVX0_HVT U7101 ( .A(n5576), .Y(n5557) );
  MUX41X1_HVT U7102 ( .A1(\ram[15][151] ), .A3(\ram[13][151] ), .A2(
        \ram[14][151] ), .A4(\ram[12][151] ), .S0(n5884), .S1(n7294), .Y(n8333) );
  MUX41X1_HVT U7103 ( .A1(\ram[7][118] ), .A3(\ram[5][118] ), .A2(
        \ram[6][118] ), .A4(\ram[4][118] ), .S0(n5941), .S1(n4888), .Y(n8204)
         );
  MUX41X1_HVT U7104 ( .A1(n8119), .A3(n8121), .A2(n8118), .A4(n8120), .S0(
        n5352), .S1(n5873), .Y(q[97]) );
  MUX41X1_HVT U7105 ( .A1(n8210), .A3(n8212), .A2(n8211), .A4(n8213), .S0(
        n7276), .S1(n7299), .Y(q[120]) );
  MUX41X1_HVT U7106 ( .A1(\ram[14][10] ), .A3(\ram[12][10] ), .A2(
        \ram[15][10] ), .A4(\ram[13][10] ), .S0(n6128), .S1(n5851), .Y(n7774)
         );
  IBUFFX2_HVT U7107 ( .A(n8769), .Y(n5820) );
  MUX41X1_HVT U7108 ( .A1(\ram[12][158] ), .A3(\ram[14][158] ), .A2(
        \ram[13][158] ), .A4(\ram[15][158] ), .S0(n5558), .S1(n5642), .Y(n8361) );
  NOR2X4_HVT U7109 ( .A1(n6129), .A2(n7272), .Y(n38) );
  MUX41X1_HVT U7110 ( .A1(\ram[8][218] ), .A3(\ram[10][218] ), .A2(
        \ram[9][218] ), .A4(\ram[11][218] ), .S0(n5558), .S1(n8901), .Y(n8602)
         );
  INVX0_HVT U7111 ( .A(n5816), .Y(n5559) );
  INVX0_HVT U7112 ( .A(n8849), .Y(n5816) );
  OAI22X1_HVT U7113 ( .A1(n5561), .A2(n10286), .A3(n5849), .A4(n9355), .Y(
        n1613) );
  IBUFFX2_HVT U7114 ( .A(n4971), .Y(n5944) );
  INVX0_HVT U7115 ( .A(n25), .Y(n5879) );
  INVX0_HVT U7116 ( .A(n5590), .Y(n7268) );
  INVX0_HVT U7117 ( .A(n4972), .Y(n10276) );
  INVX0_HVT U7118 ( .A(n10287), .Y(n10280) );
  INVX0_HVT U7119 ( .A(n10286), .Y(n10282) );
  INVX0_HVT U7120 ( .A(n4972), .Y(n10279) );
  INVX0_HVT U7121 ( .A(n7583), .Y(n5564) );
  NBUFFX2_HVT U7122 ( .A(n13), .Y(n5563) );
  INVX0_HVT U7123 ( .A(n8806), .Y(n7583) );
  MUX41X1_HVT U7124 ( .A1(\ram[14][102] ), .A3(\ram[12][102] ), .A2(
        \ram[15][102] ), .A4(\ram[13][102] ), .S0(n7690), .S1(n5950), .Y(n8138) );
  NBUFFX2_HVT U7125 ( .A(n6127), .Y(n8890) );
  INVX0_HVT U7126 ( .A(n7692), .Y(n5565) );
  NBUFFX2_HVT U7127 ( .A(n8801), .Y(n5854) );
  NBUFFX2_HVT U7128 ( .A(n5986), .Y(n5567) );
  INVX0_HVT U7129 ( .A(n6018), .Y(n5973) );
  MUX41X1_HVT U7130 ( .A1(n8134), .A3(n8136), .A2(n8135), .A4(n8137), .S0(
        n5720), .S1(n5820), .Y(q[101]) );
  INVX0_HVT U7131 ( .A(n5618), .Y(n5569) );
  MUX41X1_HVT U7132 ( .A1(n8014), .A3(n8016), .A2(n8015), .A4(n8017), .S0(
        n5720), .S1(n5648), .Y(q[71]) );
  INVX0_HVT U7133 ( .A(n6659), .Y(n5720) );
  INVX0_HVT U7134 ( .A(n5040), .Y(n5648) );
  MUX41X1_HVT U7135 ( .A1(n7784), .A3(n7782), .A2(n7785), .A4(n7783), .S0(
        n5815), .S1(n5332), .Y(q[12]) );
  INVX0_HVT U7136 ( .A(n6119), .Y(n10274) );
  INVX0_HVT U7137 ( .A(n7326), .Y(n5998) );
  MUX41X1_HVT U7138 ( .A1(n8222), .A3(n8224), .A2(n8223), .A4(n8225), .S0(
        n5886), .S1(n7288), .Y(q[123]) );
  NBUFFX2_HVT U7139 ( .A(n7584), .Y(n7715) );
  INVX0_HVT U7140 ( .A(n8806), .Y(n7697) );
  MUX41X1_HVT U7141 ( .A1(n7880), .A3(n7882), .A2(n7879), .A4(n7881), .S0(
        n5886), .S1(n5622), .Y(q[37]) );
  INVX0_HVT U7142 ( .A(n5618), .Y(n8806) );
  INVX0_HVT U7143 ( .A(n5784), .Y(n5785) );
  NBUFFX2_HVT U7144 ( .A(n7565), .Y(n7670) );
  NBUFFX2_HVT U7145 ( .A(n5853), .Y(n8858) );
  NBUFFX2_HVT U7146 ( .A(n6891), .Y(n7707) );
  INVX0_HVT U7147 ( .A(n5487), .Y(n6253) );
  MUX41X1_HVT U7148 ( .A1(n8009), .A3(n8007), .A2(n8008), .A4(n8006), .S0(
        n5815), .S1(n5801), .Y(q[69]) );
  INVX0_HVT U7149 ( .A(n6392), .Y(n5577) );
  INVX0_HVT U7150 ( .A(n5813), .Y(n5579) );
  INVX0_HVT U7151 ( .A(n5478), .Y(n5813) );
  NBUFFX2_HVT U7152 ( .A(n6758), .Y(n7342) );
  NBUFFX2_HVT U7153 ( .A(n6030), .Y(n6744) );
  INVX1_HVT U7154 ( .A(n5881), .Y(n5582) );
  MUX41X1_HVT U7155 ( .A1(n8150), .A3(n8152), .A2(n8151), .A4(n8153), .S0(
        n5111), .S1(n5637), .Y(q[105]) );
  INVX0_HVT U7156 ( .A(n7323), .Y(n5881) );
  NBUFFX2_HVT U7157 ( .A(n6010), .Y(n5585) );
  IBUFFX2_HVT U7158 ( .A(n7267), .Y(n6010) );
  NBUFFX2_HVT U7159 ( .A(n7581), .Y(n5586) );
  INVX0_HVT U7160 ( .A(n5762), .Y(n5587) );
  NAND2X0_HVT U7161 ( .A1(n5765), .A2(n5835), .Y(n5590) );
  MUX41X1_HVT U7162 ( .A1(\ram[3][15] ), .A3(\ram[1][15] ), .A2(\ram[2][15] ), 
        .A4(\ram[0][15] ), .S0(n5903), .S1(n5724), .Y(n7797) );
  INVX0_HVT U7163 ( .A(n5927), .Y(n8610) );
  NBUFFX2_HVT U7164 ( .A(n8882), .Y(n7279) );
  INVX0_HVT U7165 ( .A(n6007), .Y(n5803) );
  INVX0_HVT U7166 ( .A(n5905), .Y(n6030) );
  NBUFFX2_HVT U7167 ( .A(n6739), .Y(n8876) );
  MUX41X1_HVT U7168 ( .A1(\ram[4][136] ), .A3(\ram[6][136] ), .A2(
        \ram[5][136] ), .A4(\ram[7][136] ), .S0(n5997), .S1(n5539), .Y(n8276)
         );
  INVX0_HVT U7169 ( .A(n5154), .Y(n5595) );
  MUX41X1_HVT U7170 ( .A1(\ram[11][198] ), .A3(\ram[9][198] ), .A2(
        \ram[10][198] ), .A4(\ram[8][198] ), .S0(n5594), .S1(n4977), .Y(n8522)
         );
  IBUFFX2_HVT U7171 ( .A(n7566), .Y(n7288) );
  MUX41X1_HVT U7172 ( .A1(\ram[4][138] ), .A3(\ram[6][138] ), .A2(
        \ram[5][138] ), .A4(\ram[7][138] ), .S0(n5932), .S1(n8880), .Y(n8284)
         );
  MUX41X1_HVT U7173 ( .A1(\ram[15][87] ), .A3(\ram[13][87] ), .A2(
        \ram[14][87] ), .A4(\ram[12][87] ), .S0(n5772), .S1(n7672), .Y(n8078)
         );
  OAI22X1_HVT U7174 ( .A1(n5597), .A2(n5379), .A3(n5603), .A4(n5596), .Y(n4148) );
  OAI22X1_HVT U7175 ( .A1(n5598), .A2(n5381), .A3(n10093), .A4(n10042), .Y(
        n4141) );
  IBUFFX2_HVT U7176 ( .A(n10096), .Y(n10093) );
  OAI22X1_HVT U7177 ( .A1(n5599), .A2(n5378), .A3(n10095), .A4(n9753), .Y(
        n4049) );
  INVX0_HVT U7178 ( .A(n5531), .Y(n5600) );
  INVX0_HVT U7179 ( .A(n5784), .Y(n5661) );
  NBUFFX2_HVT U7180 ( .A(n6253), .Y(n5601) );
  INVX0_HVT U7181 ( .A(n8775), .Y(n5828) );
  MUX41X1_HVT U7182 ( .A1(\ram[11][48] ), .A3(\ram[9][48] ), .A2(\ram[10][48] ), .A4(\ram[8][48] ), .S0(n5602), .S1(n5493), .Y(n7924) );
  NBUFFX2_HVT U7183 ( .A(n6185), .Y(n7665) );
  MUX41X1_HVT U7184 ( .A1(\ram[3][41] ), .A3(\ram[1][41] ), .A2(\ram[2][41] ), 
        .A4(\ram[0][41] ), .S0(n5605), .S1(n5606), .Y(n7898) );
  NBUFFX2_HVT U7185 ( .A(n5641), .Y(n8853) );
  IBUFFX2_HVT U7186 ( .A(n8774), .Y(n5877) );
  NBUFFX2_HVT U7187 ( .A(n5164), .Y(n8907) );
  INVX0_HVT U7188 ( .A(n8763), .Y(n6129) );
  MUX41X1_HVT U7189 ( .A1(n7812), .A3(n7810), .A2(n7813), .A4(n7811), .S0(
        n5156), .S1(n5828), .Y(q[19]) );
  NBUFFX2_HVT U7190 ( .A(n6759), .Y(n5989) );
  NBUFFX2_HVT U7191 ( .A(n5661), .Y(n5610) );
  NBUFFX2_HVT U7192 ( .A(n5862), .Y(n8899) );
  NBUFFX2_HVT U7193 ( .A(n5661), .Y(n5612) );
  INVX0_HVT U7194 ( .A(n8757), .Y(n5613) );
  NBUFFX2_HVT U7195 ( .A(n7670), .Y(n5615) );
  INVX0_HVT U7196 ( .A(n5902), .Y(n5746) );
  INVX1_HVT U7197 ( .A(n5747), .Y(n5616) );
  INVX0_HVT U7198 ( .A(n8784), .Y(n5617) );
  NBUFFX2_HVT U7199 ( .A(n7287), .Y(n6406) );
  MUX41X1_HVT U7200 ( .A1(\ram[11][40] ), .A3(\ram[9][40] ), .A2(\ram[10][40] ), .A4(\ram[8][40] ), .S0(n5998), .S1(n5005), .Y(n7892) );
  INVX0_HVT U7201 ( .A(n10378), .Y(n10377) );
  INVX0_HVT U7202 ( .A(n5682), .Y(n5697) );
  INVX0_HVT U7203 ( .A(n5682), .Y(n5696) );
  INVX0_HVT U7204 ( .A(n5673), .Y(n5682) );
  NBUFFX2_HVT U7205 ( .A(n4979), .Y(n7684) );
  NBUFFX2_HVT U7206 ( .A(n6030), .Y(n7581) );
  MUX41X1_HVT U7207 ( .A1(n8632), .A3(n8630), .A2(n8631), .A4(n8629), .S0(
        n5317), .S1(n8772), .Y(q[225]) );
  NAND2X0_HVT U7208 ( .A1(n8), .A2(n5619), .Y(n5981) );
  AND2X1_HVT U7209 ( .A1(n10377), .A2(n6013), .Y(n5619) );
  INVX0_HVT U7210 ( .A(n6012), .Y(n5620) );
  MUX41X1_HVT U7211 ( .A1(\ram[3][252] ), .A3(\ram[1][252] ), .A2(
        \ram[2][252] ), .A4(\ram[0][252] ), .S0(n5863), .S1(n7142), .Y(n8738)
         );
  MUX41X1_HVT U7212 ( .A1(n8542), .A3(n8541), .A2(n8544), .A4(n8543), .S0(
        n7352), .S1(n7548), .Y(q[203]) );
  INVX0_HVT U7213 ( .A(n4162), .Y(n5884) );
  MUX41X1_HVT U7214 ( .A1(n7959), .A3(n7961), .A2(n7960), .A4(n7962), .S0(
        n5723), .S1(n5809), .Y(q[57]) );
  AOI21X1_HVT U7215 ( .A1(n20), .A2(n10377), .A3(n10381), .Y(n18) );
  MUX41X1_HVT U7216 ( .A1(\ram[12][195] ), .A3(\ram[14][195] ), .A2(
        \ram[13][195] ), .A4(\ram[15][195] ), .S0(n5733), .S1(n4921), .Y(n8509) );
  MUX41X1_HVT U7217 ( .A1(\ram[3][250] ), .A3(\ram[1][250] ), .A2(
        \ram[2][250] ), .A4(\ram[0][250] ), .S0(n5975), .S1(n5141), .Y(n8730)
         );
  MUX41X1_HVT U7218 ( .A1(\ram[11][237] ), .A3(\ram[9][237] ), .A2(
        \ram[10][237] ), .A4(\ram[8][237] ), .S0(n5937), .S1(n5288), .Y(n8676)
         );
  MUX41X1_HVT U7219 ( .A1(n8333), .A3(n8334), .A2(n8335), .A4(n8336), .S0(
        n5624), .S1(n5634), .Y(q[151]) );
  INVX0_HVT U7220 ( .A(n5518), .Y(n7263) );
  MUX41X1_HVT U7221 ( .A1(n8576), .A3(n8574), .A2(n8575), .A4(n8573), .S0(
        n5625), .S1(n5307), .Y(q[211]) );
  AND2X1_HVT U7222 ( .A1(n25), .A2(n17), .Y(n5626) );
  MUX41X1_HVT U7223 ( .A1(\ram[11][4] ), .A3(\ram[9][4] ), .A2(\ram[10][4] ), 
        .A4(\ram[8][4] ), .S0(n5627), .S1(n7146), .Y(n7751) );
  NBUFFX2_HVT U7224 ( .A(n7674), .Y(n8901) );
  MUX41X1_HVT U7225 ( .A1(\ram[7][145] ), .A3(\ram[5][145] ), .A2(
        \ram[6][145] ), .A4(\ram[4][145] ), .S0(n5937), .S1(n5568), .Y(n8311)
         );
  MUX41X1_HVT U7226 ( .A1(\ram[8][230] ), .A3(\ram[10][230] ), .A2(
        \ram[9][230] ), .A4(\ram[11][230] ), .S0(n5630), .S1(n5629), .Y(n8650)
         );
  NBUFFX2_HVT U7227 ( .A(n6132), .Y(n8894) );
  MUX41X1_HVT U7228 ( .A1(\ram[12][163] ), .A3(\ram[14][163] ), .A2(
        \ram[13][163] ), .A4(\ram[15][163] ), .S0(n5294), .S1(n8861), .Y(n8381) );
  INVX0_HVT U7229 ( .A(n9243), .Y(n9251) );
  NBUFFX2_HVT U7230 ( .A(n7346), .Y(n5632) );
  MUX41X1_HVT U7231 ( .A1(\ram[15][192] ), .A3(\ram[13][192] ), .A2(
        \ram[14][192] ), .A4(\ram[12][192] ), .S0(n5638), .S1(n7709), .Y(n8497) );
  MUX41X1_HVT U7232 ( .A1(\ram[15][43] ), .A3(\ram[14][43] ), .A2(
        \ram[13][43] ), .A4(\ram[12][43] ), .S0(n5001), .S1(n7277), .Y(n7903)
         );
  NBUFFX2_HVT U7233 ( .A(n8888), .Y(n5639) );
  INVX0_HVT U7234 ( .A(n6131), .Y(n7693) );
  MUX41X1_HVT U7235 ( .A1(\ram[7][236] ), .A3(\ram[6][236] ), .A2(
        \ram[5][236] ), .A4(\ram[4][236] ), .S0(n6740), .S1(n5742), .Y(n8673)
         );
  MUX41X1_HVT U7236 ( .A1(\ram[15][245] ), .A3(\ram[13][245] ), .A2(
        \ram[14][245] ), .A4(\ram[12][245] ), .S0(n5743), .S1(n5077), .Y(n8707) );
  INVX0_HVT U7237 ( .A(n5537), .Y(n5647) );
  NAND2X0_HVT U7238 ( .A1(n5247), .A2(n9928), .Y(n5644) );
  NAND2X0_HVT U7239 ( .A1(n5644), .A2(n5643), .Y(n1032) );
  INVX0_HVT U7240 ( .A(n7120), .Y(n7122) );
  INVX0_HVT U7241 ( .A(n8789), .Y(n5824) );
  INVX0_HVT U7242 ( .A(n7322), .Y(n6390) );
  INVX0_HVT U7243 ( .A(n8782), .Y(n8808) );
  INVX0_HVT U7244 ( .A(n7308), .Y(n7267) );
  MUX41X1_HVT U7245 ( .A1(\ram[7][90] ), .A3(\ram[5][90] ), .A2(\ram[6][90] ), 
        .A4(\ram[4][90] ), .S0(n5647), .S1(n5719), .Y(n8092) );
  MUX41X1_HVT U7246 ( .A1(\ram[11][31] ), .A3(\ram[9][31] ), .A2(\ram[10][31] ), .A4(\ram[8][31] ), .S0(n5333), .S1(n5730), .Y(n7856) );
  INVX0_HVT U7247 ( .A(n5866), .Y(n6660) );
  MUX41X1_HVT U7248 ( .A1(n8102), .A3(n8104), .A2(n8103), .A4(n8105), .S0(
        n5830), .S1(n5648), .Y(q[93]) );
  NBUFFX2_HVT U7249 ( .A(n7279), .Y(n5649) );
  INVX0_HVT U7250 ( .A(n5988), .Y(n6114) );
  INVX0_HVT U7251 ( .A(n8765), .Y(n10379) );
  MUX41X1_HVT U7252 ( .A1(\ram[8][148] ), .A3(\ram[10][148] ), .A2(
        \ram[9][148] ), .A4(\ram[11][148] ), .S0(n5000), .S1(n5652), .Y(n8322)
         );
  NBUFFX2_HVT U7253 ( .A(n5947), .Y(n7547) );
  INVX0_HVT U7254 ( .A(n5719), .Y(n5652) );
  INVX0_HVT U7255 ( .A(n7125), .Y(n6255) );
  INVX0_HVT U7256 ( .A(n7130), .Y(n7132) );
  MUX41X1_HVT U7257 ( .A1(n8553), .A3(n8555), .A2(n8554), .A4(n8556), .S0(
        n5655), .S1(n5737), .Y(q[206]) );
  NBUFFX2_HVT U7258 ( .A(n7708), .Y(n8867) );
  MUX41X1_HVT U7259 ( .A1(\ram[15][135] ), .A3(\ram[14][135] ), .A2(
        \ram[13][135] ), .A4(\ram[12][135] ), .S0(n5813), .S1(n5605), .Y(n8270) );
  INVX0_HVT U7260 ( .A(n7717), .Y(n5660) );
  MUX41X1_HVT U7261 ( .A1(\ram[11][76] ), .A3(\ram[9][76] ), .A2(\ram[10][76] ), .A4(\ram[8][76] ), .S0(n5878), .S1(n6753), .Y(n8035) );
  IBUFFX2_HVT U7262 ( .A(n7297), .Y(n8814) );
  MUX41X1_HVT U7263 ( .A1(n8419), .A3(n8417), .A2(n8420), .A4(n8418), .S0(
        n5867), .S1(n5660), .Y(q[172]) );
  NBUFFX2_HVT U7264 ( .A(n4942), .Y(n5669) );
  NBUFFX2_HVT U7265 ( .A(n4942), .Y(n5670) );
  NBUFFX2_HVT U7266 ( .A(n5668), .Y(n5671) );
  NBUFFX2_HVT U7267 ( .A(n5668), .Y(n5672) );
  NBUFFX2_HVT U7268 ( .A(n4765), .Y(n5674) );
  NBUFFX2_HVT U7269 ( .A(n4764), .Y(n5675) );
  NBUFFX2_HVT U7270 ( .A(n5121), .Y(n5676) );
  NBUFFX2_HVT U7271 ( .A(n5708), .Y(n5677) );
  NBUFFX2_HVT U7272 ( .A(n5121), .Y(n5678) );
  INVX0_HVT U7273 ( .A(n5121), .Y(n5679) );
  INVX0_HVT U7274 ( .A(n5673), .Y(n5680) );
  INVX0_HVT U7275 ( .A(n5673), .Y(n5681) );
  INVX0_HVT U7276 ( .A(n4748), .Y(n5683) );
  INVX0_HVT U7277 ( .A(n5679), .Y(n5684) );
  INVX0_HVT U7278 ( .A(n5679), .Y(n5685) );
  INVX0_HVT U7279 ( .A(n4748), .Y(n5686) );
  INVX0_HVT U7280 ( .A(n5680), .Y(n5687) );
  INVX0_HVT U7281 ( .A(n5680), .Y(n5692) );
  INVX0_HVT U7282 ( .A(n5682), .Y(n5693) );
  INVX0_HVT U7283 ( .A(n5663), .Y(n5698) );
  INVX0_HVT U7284 ( .A(n5663), .Y(n5700) );
  INVX0_HVT U7285 ( .A(n5698), .Y(n5701) );
  INVX0_HVT U7286 ( .A(n4710), .Y(n5703) );
  INVX0_HVT U7287 ( .A(n5699), .Y(n5704) );
  INVX0_HVT U7288 ( .A(n5700), .Y(n5705) );
  INVX0_HVT U7289 ( .A(n4710), .Y(n5706) );
  INVX0_HVT U7290 ( .A(n4640), .Y(n5707) );
  INVX0_HVT U7291 ( .A(n5699), .Y(n5709) );
  INVX0_HVT U7292 ( .A(n5698), .Y(n5710) );
  INVX0_HVT U7293 ( .A(n4710), .Y(n5711) );
  INVX0_HVT U7294 ( .A(n5700), .Y(n5712) );
  INVX0_HVT U7295 ( .A(n4710), .Y(n5713) );
  MUX41X1_HVT U7296 ( .A1(n5716), .A3(n5436), .A2(n5717), .A4(n5718), .S0(
        n6389), .S1(n5715), .Y(n5714) );
  INVX0_HVT U7297 ( .A(n9004), .Y(n9006) );
  MUX41X1_HVT U7298 ( .A1(\ram[3][128] ), .A3(\ram[1][128] ), .A2(
        \ram[2][128] ), .A4(\ram[0][128] ), .S0(n5742), .S1(n5719), .Y(n8245)
         );
  NBUFFX2_HVT U7299 ( .A(n6662), .Y(n8900) );
  MUX41X1_HVT U7300 ( .A1(\ram[6][108] ), .A3(\ram[4][108] ), .A2(
        \ram[7][108] ), .A4(\ram[5][108] ), .S0(n5969), .S1(n5292), .Y(n8164)
         );
  INVX0_HVT U7301 ( .A(n6733), .Y(n7690) );
  MUX41X1_HVT U7302 ( .A1(n6555), .A3(n6554), .A2(n6553), .A4(n6552), .S0(
        n5978), .S1(n7700), .Y(n6550) );
  MUX41X1_HVT U7303 ( .A1(n8062), .A3(n8064), .A2(n8063), .A4(n8065), .S0(
        n5151), .S1(n5776), .Y(q[83]) );
  MUX41X1_HVT U7304 ( .A1(n8114), .A3(n8116), .A2(n8115), .A4(n8117), .S0(
        n5720), .S1(n5721), .Y(q[96]) );
  INVX0_HVT U7305 ( .A(n8782), .Y(n8792) );
  INVX0_HVT U7306 ( .A(n5338), .Y(n5931) );
  MUX41X1_HVT U7307 ( .A1(\ram[3][229] ), .A3(\ram[1][229] ), .A2(
        \ram[2][229] ), .A4(\ram[0][229] ), .S0(n7334), .S1(n5722), .Y(n8648)
         );
  NBUFFX2_HVT U7308 ( .A(n7693), .Y(n7669) );
  MUX41X1_HVT U7309 ( .A1(n8357), .A3(n8359), .A2(n8358), .A4(n8360), .S0(
        n5343), .S1(n5721), .Y(q[157]) );
  INVX0_HVT U7310 ( .A(n5078), .Y(n5830) );
  NBUFFX2_HVT U7311 ( .A(n5314), .Y(n7560) );
  IBUFFX2_HVT U7312 ( .A(n7318), .Y(n6657) );
  INVX0_HVT U7313 ( .A(n4829), .Y(n7011) );
  INVX0_HVT U7314 ( .A(n7007), .Y(n7009) );
  INVX0_HVT U7315 ( .A(n7006), .Y(n7008) );
  INVX0_HVT U7316 ( .A(n7197), .Y(n7202) );
  INVX0_HVT U7317 ( .A(n7197), .Y(n7201) );
  INVX0_HVT U7318 ( .A(n9072), .Y(n9078) );
  INVX0_HVT U7319 ( .A(n7253), .Y(n7256) );
  INVX0_HVT U7320 ( .A(n7245), .Y(n7251) );
  INVX0_HVT U7321 ( .A(n4582), .Y(n7195) );
  INVX0_HVT U7322 ( .A(n7063), .Y(n7068) );
  INVX0_HVT U7323 ( .A(n7073), .Y(n7078) );
  INVX0_HVT U7324 ( .A(n7244), .Y(n7248) );
  INVX0_HVT U7325 ( .A(n7197), .Y(n7199) );
  INVX0_HVT U7326 ( .A(n5748), .Y(n10104) );
  INVX0_HVT U7327 ( .A(n5531), .Y(n10098) );
  MUX41X1_HVT U7328 ( .A1(n7943), .A3(n7945), .A2(n7944), .A4(n7946), .S0(
        n5720), .S1(n5344), .Y(q[53]) );
  NBUFFX2_HVT U7329 ( .A(n7565), .Y(n8872) );
  MUX41X1_HVT U7330 ( .A1(\ram[3][190] ), .A3(\ram[2][190] ), .A2(
        \ram[1][190] ), .A4(\ram[0][190] ), .S0(n5304), .S1(n5829), .Y(n8492)
         );
  INVX0_HVT U7331 ( .A(n5852), .Y(n5832) );
  AO22X1_HVT U7332 ( .A1(\ram[13][144] ), .A2(n7018), .A3(n8916), .A4(n9742), 
        .Y(n3533) );
  INVX0_HVT U7333 ( .A(n7016), .Y(n7018) );
  OAI22X1_HVT U7334 ( .A1(n5725), .A2(n6735), .A3(n6229), .A4(n9369), .Y(n1106) );
  OAI22X1_HVT U7335 ( .A1(n5726), .A2(n5061), .A3(n5451), .A4(n9333), .Y(n1094) );
  OAI22X1_HVT U7336 ( .A1(n5727), .A2(n6735), .A3(n6238), .A4(n9330), .Y(n1093) );
  OAI22X1_HVT U7337 ( .A1(n6555), .A2(n5061), .A3(n6196), .A4(n9367), .Y(n1105) );
  INVX0_HVT U7338 ( .A(n6736), .Y(n6737) );
  INVX0_HVT U7339 ( .A(n8779), .Y(n7343) );
  MUX41X1_HVT U7340 ( .A1(\ram[11][196] ), .A3(\ram[9][196] ), .A2(
        \ram[10][196] ), .A4(\ram[8][196] ), .S0(n7305), .S1(n5730), .Y(n8514)
         );
  MUX41X1_HVT U7341 ( .A1(n8258), .A3(n8260), .A2(n8259), .A4(n8261), .S0(
        n5736), .S1(n5373), .Y(q[132]) );
  MUX41X1_HVT U7342 ( .A1(n8207), .A3(n8209), .A2(n8206), .A4(n8208), .S0(
        n6120), .S1(n5755), .Y(q[119]) );
  MUX41X1_HVT U7343 ( .A1(\ram[3][93] ), .A3(\ram[1][93] ), .A2(\ram[2][93] ), 
        .A4(\ram[0][93] ), .S0(n5979), .S1(n5304), .Y(n8105) );
  INVX0_HVT U7344 ( .A(n6391), .Y(n7312) );
  MUX41X1_HVT U7345 ( .A1(n8682), .A3(n8680), .A2(n8681), .A4(n8679), .S0(
        n5833), .S1(n8768), .Y(q[238]) );
  NBUFFX2_HVT U7346 ( .A(n4848), .Y(n7278) );
  MUX41X1_HVT U7347 ( .A1(n8279), .A3(n8281), .A2(n8278), .A4(n8280), .S0(
        n5655), .S1(n5852), .Y(q[137]) );
  INVX0_HVT U7348 ( .A(n5646), .Y(n5894) );
  MUX41X1_HVT U7349 ( .A1(\ram[7][82] ), .A3(\ram[5][82] ), .A2(\ram[6][82] ), 
        .A4(\ram[4][82] ), .S0(n4958), .S1(n5864), .Y(n8060) );
  INVX0_HVT U7350 ( .A(n5652), .Y(n7282) );
  NBUFFX2_HVT U7351 ( .A(n5641), .Y(n7563) );
  NBUFFX2_HVT U7352 ( .A(n5996), .Y(n8877) );
  NBUFFX2_HVT U7353 ( .A(n5553), .Y(n6386) );
  MUX41X1_HVT U7354 ( .A1(n8725), .A3(n8723), .A2(n8726), .A4(n8724), .S0(
        n5625), .S1(n5773), .Y(q[249]) );
  INVX0_HVT U7355 ( .A(n5540), .Y(n10107) );
  INVX0_HVT U7356 ( .A(n10108), .Y(n10112) );
  MUX41X1_HVT U7357 ( .A1(\ram[11][177] ), .A3(\ram[9][177] ), .A2(
        \ram[10][177] ), .A4(\ram[8][177] ), .S0(n5507), .S1(n7283), .Y(n8438)
         );
  NBUFFX2_HVT U7358 ( .A(n7718), .Y(n7559) );
  INVX0_HVT U7359 ( .A(n8759), .Y(n7276) );
  INVX0_HVT U7360 ( .A(n5905), .Y(n6001) );
  MUX21X1_HVT U7361 ( .A1(\ram[15][83] ), .A2(\ram[13][83] ), .S0(n5941), .Y(
        n5744) );
  MUX21X1_HVT U7362 ( .A1(\ram[14][83] ), .A2(\ram[12][83] ), .S0(n6128), .Y(
        n5745) );
  NBUFFX2_HVT U7363 ( .A(n8801), .Y(n5900) );
  MUX41X1_HVT U7364 ( .A1(n8496), .A3(n8494), .A2(n8495), .A4(n8493), .S0(
        n5654), .S1(n5746), .Y(q[191]) );
  INVX0_HVT U7365 ( .A(N28), .Y(n8765) );
  INVX0_HVT U7366 ( .A(n8900), .Y(n7285) );
  MUX41X1_HVT U7367 ( .A1(\ram[8][234] ), .A3(\ram[10][234] ), .A2(
        \ram[9][234] ), .A4(\ram[11][234] ), .S0(n8832), .S1(n6763), .Y(n8664)
         );
  MUX41X1_HVT U7368 ( .A1(\ram[7][5] ), .A3(\ram[5][5] ), .A2(\ram[6][5] ), 
        .A4(\ram[4][5] ), .S0(n5759), .S1(n6393), .Y(n7756) );
  MUX41X1_HVT U7369 ( .A1(\ram[10][187] ), .A3(\ram[11][187] ), .A2(
        \ram[8][187] ), .A4(\ram[9][187] ), .S0(n5760), .S1(n5863), .Y(n8478)
         );
  NBUFFX2_HVT U7370 ( .A(n7584), .Y(n8771) );
  INVX0_HVT U7371 ( .A(n5543), .Y(n5753) );
  MUX41X1_HVT U7372 ( .A1(n8408), .A3(n8406), .A2(n8407), .A4(n8405), .S0(
        n5756), .S1(n5755), .Y(q[169]) );
  INVX0_HVT U7373 ( .A(n4913), .Y(n7718) );
  MUX41X1_HVT U7374 ( .A1(n8372), .A3(n8370), .A2(n8371), .A4(n8369), .S0(
        n5756), .S1(n5808), .Y(q[160]) );
  MUX41X1_HVT U7375 ( .A1(n8286), .A3(n8288), .A2(n8287), .A4(n8289), .S0(
        n5151), .S1(n5757), .Y(q[139]) );
  NBUFFX2_HVT U7376 ( .A(n5590), .Y(n6119) );
  INVX0_HVT U7377 ( .A(n4718), .Y(n5761) );
  NAND2X0_HVT U7378 ( .A1(\ram[6][50] ), .A2(n5516), .Y(n5763) );
  NAND2X0_HVT U7379 ( .A1(n9198), .A2(n9457), .Y(n5764) );
  NAND2X0_HVT U7380 ( .A1(n5763), .A2(n5764), .Y(n1647) );
  NAND2X0_HVT U7381 ( .A1(n6037), .A2(n5626), .Y(n5765) );
  NAND2X0_HVT U7382 ( .A1(n5765), .A2(n5835), .Y(n6036) );
  INVX0_HVT U7383 ( .A(n8820), .Y(n5766) );
  NBUFFX2_HVT U7384 ( .A(n6754), .Y(n7309) );
  MUX41X1_HVT U7385 ( .A1(n8599), .A3(n8600), .A2(n8597), .A4(n8598), .S0(
        n5773), .S1(n7300), .Y(q[217]) );
  INVX1_HVT U7386 ( .A(n6381), .Y(n5980) );
  MUX21X1_HVT U7387 ( .A1(\ram[1][48] ), .A2(\ram[3][48] ), .S0(n5888), .Y(
        n5769) );
  NBUFFX2_HVT U7388 ( .A(n6891), .Y(n8881) );
  INVX0_HVT U7389 ( .A(n8757), .Y(n7339) );
  MUX41X1_HVT U7390 ( .A1(n7998), .A3(n8000), .A2(n7999), .A4(n8001), .S0(
        n5830), .S1(n5770), .Y(q[67]) );
  INVX1_HVT U7391 ( .A(rst), .Y(n5835) );
  NBUFFX2_HVT U7392 ( .A(n6185), .Y(n8903) );
  MUX41X1_HVT U7393 ( .A1(\ram[7][66] ), .A3(\ram[5][66] ), .A2(\ram[6][66] ), 
        .A4(\ram[4][66] ), .S0(n5772), .S1(n7716), .Y(n7996) );
  NBUFFX2_HVT U7394 ( .A(n6662), .Y(n7694) );
  INVX0_HVT U7395 ( .A(we), .Y(n10378) );
  INVX0_HVT U7396 ( .A(we), .Y(n6639) );
  MUX41X1_HVT U7397 ( .A1(n8735), .A3(n8737), .A2(n8736), .A4(n8738), .S0(
        n5364), .S1(n5773), .Y(q[252]) );
  MUX41X1_HVT U7398 ( .A1(n8409), .A3(n8411), .A2(n8410), .A4(n8412), .S0(
        n5830), .S1(n5774), .Y(q[170]) );
  INVX0_HVT U7399 ( .A(n8900), .Y(n5775) );
  MUX41X1_HVT U7400 ( .A1(n7885), .A3(n7883), .A2(n7886), .A4(n7884), .S0(
        n5363), .S1(n5776), .Y(q[38]) );
  NBUFFX2_HVT U7401 ( .A(n6001), .Y(n5777) );
  INVX0_HVT U7402 ( .A(n5759), .Y(n5890) );
  MUX41X1_HVT U7403 ( .A1(\ram[15][50] ), .A3(\ram[13][50] ), .A2(
        \ram[14][50] ), .A4(\ram[12][50] ), .S0(n5602), .S1(n5826), .Y(n7931)
         );
  INVX0_HVT U7404 ( .A(n7668), .Y(n5906) );
  MUX21X1_HVT U7405 ( .A1(\ram[12][253] ), .A2(\ram[14][253] ), .S0(n7553), 
        .Y(n6125) );
  MUX21X1_HVT U7406 ( .A1(n5780), .A2(n5779), .S0(n5573), .Y(n5778) );
  MUX41X1_HVT U7407 ( .A1(n8740), .A3(n8742), .A2(n8739), .A4(n8741), .S0(
        n5352), .S1(n7280), .Y(q[253]) );
  MUX41X1_HVT U7408 ( .A1(n8242), .A3(n8244), .A2(n8243), .A4(n8245), .S0(
        n5372), .S1(n5199), .Y(q[128]) );
  INVX0_HVT U7409 ( .A(n7347), .Y(n5784) );
  MUX41X1_HVT U7410 ( .A1(\ram[15][221] ), .A3(\ram[14][221] ), .A2(
        \ram[13][221] ), .A4(\ram[12][221] ), .S0(n6393), .S1(n5759), .Y(n8613) );
  OAI22X1_HVT U7411 ( .A1(n5786), .A2(n5667), .A3(n7269), .A4(n9453), .Y(n1390) );
  MUX41X1_HVT U7412 ( .A1(\ram[13][174] ), .A3(\ram[15][174] ), .A2(
        \ram[12][174] ), .A4(\ram[14][174] ), .S0(n5793), .S1(n5893), .Y(n8425) );
  MUX41X1_HVT U7413 ( .A1(\ram[15][1] ), .A3(\ram[13][1] ), .A2(\ram[14][1] ), 
        .A4(\ram[12][1] ), .S0(n5787), .S1(n6657), .Y(n7738) );
  NAND2X0_HVT U7414 ( .A1(\ram[6][195] ), .A2(n5182), .Y(n5789) );
  NAND2X0_HVT U7415 ( .A1(n9244), .A2(n9902), .Y(n5790) );
  NAND2X0_HVT U7416 ( .A1(n5789), .A2(n5790), .Y(n1792) );
  INVX0_HVT U7417 ( .A(n9242), .Y(n9244) );
  MUX41X1_HVT U7418 ( .A1(n8710), .A3(n8709), .A2(n8708), .A4(n8707), .S0(
        n5801), .S1(n5815), .Y(q[245]) );
  MUX41X1_HVT U7419 ( .A1(n8398), .A3(n8400), .A2(n8397), .A4(n8399), .S0(
        n5901), .S1(n5791), .Y(q[167]) );
  NBUFFX2_HVT U7420 ( .A(n5862), .Y(n8904) );
  MUX41X1_HVT U7421 ( .A1(\ram[7][231] ), .A3(\ram[6][231] ), .A2(
        \ram[5][231] ), .A4(\ram[4][231] ), .S0(n5881), .S1(n5817), .Y(n8655)
         );
  MUX41X1_HVT U7422 ( .A1(\ram[12][172] ), .A3(\ram[14][172] ), .A2(
        \ram[13][172] ), .A4(\ram[15][172] ), .S0(n5940), .S1(n7342), .Y(n8417) );
  MUX41X1_HVT U7423 ( .A1(\ram[6][249] ), .A3(\ram[4][249] ), .A2(
        \ram[7][249] ), .A4(\ram[5][249] ), .S0(n5894), .S1(n5108), .Y(n8725)
         );
  MUX41X1_HVT U7424 ( .A1(n8079), .A3(n8081), .A2(n8078), .A4(n8080), .S0(
        n5831), .S1(n5896), .Y(q[87]) );
  MUX41X1_HVT U7425 ( .A1(\ram[7][59] ), .A3(\ram[5][59] ), .A2(\ram[6][59] ), 
        .A4(\ram[4][59] ), .S0(n5969), .S1(n6138), .Y(n7968) );
  INVX0_HVT U7426 ( .A(n5519), .Y(n5798) );
  INVX0_HVT U7427 ( .A(n4410), .Y(n5951) );
  MUX41X1_HVT U7428 ( .A1(\ram[7][142] ), .A3(\ram[5][142] ), .A2(
        \ram[6][142] ), .A4(\ram[4][142] ), .S0(n5803), .S1(n5874), .Y(n8300)
         );
  MUX41X1_HVT U7429 ( .A1(n8345), .A3(n8347), .A2(n8346), .A4(n8348), .S0(
        n5805), .S1(n5806), .Y(q[154]) );
  MUX41X1_HVT U7430 ( .A1(n8465), .A3(n8467), .A2(n8466), .A4(n8468), .S0(
        n5364), .S1(n7702), .Y(q[184]) );
  NAND2X0_HVT U7431 ( .A1(\ram[15][205] ), .A2(n5600), .Y(n5810) );
  NAND2X0_HVT U7432 ( .A1(n8971), .A2(n9935), .Y(n5811) );
  NAND2X0_HVT U7433 ( .A1(n5810), .A2(n5811), .Y(n4106) );
  INVX0_HVT U7434 ( .A(n5239), .Y(n6398) );
  NBUFFX2_HVT U7435 ( .A(n7559), .Y(n5812) );
  NBUFFX2_HVT U7436 ( .A(n6185), .Y(n8906) );
  MUX41X1_HVT U7437 ( .A1(\ram[11][166] ), .A3(\ram[9][166] ), .A2(
        \ram[10][166] ), .A4(\ram[8][166] ), .S0(n5814), .S1(n5836), .Y(n8394)
         );
  MUX41X1_HVT U7438 ( .A1(n8402), .A3(n8404), .A2(n8401), .A4(n8403), .S0(
        n5151), .S1(n5755), .Y(q[168]) );
  MUX41X1_HVT U7439 ( .A1(\ram[14][4] ), .A3(\ram[12][4] ), .A2(\ram[15][4] ), 
        .A4(\ram[13][4] ), .S0(n5152), .S1(n8906), .Y(n7750) );
  MUX41X1_HVT U7440 ( .A1(\ram[15][234] ), .A3(\ram[13][234] ), .A2(
        \ram[14][234] ), .A4(\ram[12][234] ), .S0(n5816), .S1(n5230), .Y(n8663) );
  INVX0_HVT U7441 ( .A(n6751), .Y(n5885) );
  MUX41X1_HVT U7442 ( .A1(\ram[15][249] ), .A3(\ram[13][249] ), .A2(
        \ram[14][249] ), .A4(\ram[12][249] ), .S0(n7313), .S1(n5740), .Y(n8723) );
  MUX41X1_HVT U7443 ( .A1(\ram[3][246] ), .A3(\ram[1][246] ), .A2(
        \ram[2][246] ), .A4(\ram[0][246] ), .S0(n5829), .S1(n4888), .Y(n8714)
         );
  MUX41X1_HVT U7444 ( .A1(n8561), .A3(n8563), .A2(n8562), .A4(n8564), .S0(
        n7276), .S1(n5157), .Y(q[208]) );
  NBUFFX2_HVT U7445 ( .A(n4188), .Y(n8864) );
  INVX0_HVT U7446 ( .A(n6023), .Y(n7304) );
  MUX41X1_HVT U7447 ( .A1(\ram[3][182] ), .A3(\ram[1][182] ), .A2(
        \ram[2][182] ), .A4(\ram[0][182] ), .S0(n5821), .S1(n4911), .Y(n8460)
         );
  INVX0_HVT U7448 ( .A(n4759), .Y(n5822) );
  MUX41X1_HVT U7449 ( .A1(n8509), .A3(n8510), .A2(n8511), .A4(n8512), .S0(
        n5904), .S1(n5870), .Y(q[195]) );
  INVX0_HVT U7450 ( .A(n8756), .Y(n5870) );
  NBUFFX2_HVT U7451 ( .A(n7584), .Y(n7666) );
  MUX41X1_HVT U7452 ( .A1(\ram[11][222] ), .A3(\ram[9][222] ), .A2(
        \ram[10][222] ), .A4(\ram[8][222] ), .S0(n7304), .S1(n5347), .Y(n8618)
         );
  NBUFFX2_HVT U7453 ( .A(n6765), .Y(n8871) );
  MUX41X1_HVT U7454 ( .A1(\ram[3][173] ), .A3(\ram[1][173] ), .A2(
        \ram[2][173] ), .A4(\ram[0][173] ), .S0(n5968), .S1(n6384), .Y(n8424)
         );
  MUX41X1_HVT U7455 ( .A1(\ram[3][16] ), .A3(\ram[1][16] ), .A2(\ram[2][16] ), 
        .A4(\ram[0][16] ), .S0(n6742), .S1(n5826), .Y(n7801) );
  MUX41X1_HVT U7456 ( .A1(n7800), .A3(n7798), .A2(n7801), .A4(n7799), .S0(
        n8764), .S1(n5902), .Y(q[16]) );
  INVX1_HVT U7457 ( .A(n5293), .Y(n5823) );
  MUX41X1_HVT U7458 ( .A1(\ram[3][211] ), .A3(\ram[1][211] ), .A2(
        \ram[2][211] ), .A4(\ram[0][211] ), .S0(n5824), .S1(n5595), .Y(n8576)
         );
  MUX41X1_HVT U7459 ( .A1(\ram[11][209] ), .A3(\ram[9][209] ), .A2(
        \ram[10][209] ), .A4(\ram[8][209] ), .S0(n7313), .S1(n5825), .Y(n8566)
         );
  NBUFFX2_HVT U7460 ( .A(n5938), .Y(n8766) );
  INVX0_HVT U7461 ( .A(n8766), .Y(n6257) );
  INVX0_HVT U7462 ( .A(n5114), .Y(n8800) );
  INVX0_HVT U7463 ( .A(n5798), .Y(n8845) );
  INVX0_HVT U7464 ( .A(n6002), .Y(n7308) );
  NBUFFX2_HVT U7465 ( .A(n6759), .Y(n8897) );
  MUX41X1_HVT U7466 ( .A1(\ram[15][22] ), .A3(\ram[13][22] ), .A2(
        \ram[14][22] ), .A4(\ram[12][22] ), .S0(n5448), .S1(n5836), .Y(n7820)
         );
  MUX41X1_HVT U7467 ( .A1(n8422), .A3(n8424), .A2(n8421), .A4(n8423), .S0(
        n7339), .S1(n5079), .Y(q[173]) );
  MUX41X1_HVT U7468 ( .A1(n8146), .A3(n8148), .A2(n8147), .A4(n8149), .S0(
        n5723), .S1(n7333), .Y(q[104]) );
  DELLN2X2_HVT U7469 ( .A(n6019), .Y(n8775) );
  MUX41X1_HVT U7470 ( .A1(n8058), .A3(n8060), .A2(n8059), .A4(n8061), .S0(
        n5831), .S1(n5832), .Y(q[82]) );
  MUX41X1_HVT U7471 ( .A1(n7968), .A3(n7966), .A2(n7969), .A4(n7967), .S0(
        n5833), .S1(n5991), .Y(q[59]) );
  NAND2X0_HVT U7472 ( .A1(n28), .A2(n6258), .Y(n5834) );
  NAND2X0_HVT U7473 ( .A1(n5834), .A2(n5835), .Y(n7732) );
  MUX41X1_HVT U7474 ( .A1(n5838), .A3(n5439), .A2(n5839), .A4(n5840), .S0(
        n6136), .S1(n5893), .Y(n5837) );
  OA22X1_HVT U7475 ( .A1(n6119), .A2(n5844), .A3(n5117), .A4(n9465), .Y(n5843)
         );
  OA22X1_HVT U7476 ( .A1(n5847), .A2(n6119), .A3(n5846), .A4(n9459), .Y(n5845)
         );
  OA22X1_HVT U7477 ( .A1(n5850), .A2(n6119), .A3(n5849), .A4(n9453), .Y(n5848)
         );
  NBUFFX2_HVT U7478 ( .A(n7278), .Y(n5851) );
  INVX0_HVT U7479 ( .A(n5959), .Y(n5852) );
  MUX41X1_HVT U7480 ( .A1(n8182), .A3(n8184), .A2(n8183), .A4(n8185), .S0(
        n5305), .S1(n6641), .Y(q[113]) );
  INVX0_HVT U7481 ( .A(n7275), .Y(n8801) );
  MUX41X1_HVT U7482 ( .A1(\ram[6][253] ), .A3(\ram[4][253] ), .A2(
        \ram[7][253] ), .A4(\ram[5][253] ), .S0(n7306), .S1(n4984), .Y(n8741)
         );
  MUX41X1_HVT U7483 ( .A1(n8613), .A3(n8615), .A2(n8614), .A4(n8616), .S0(
        n5354), .S1(n6643), .Y(q[221]) );
  MUX41X1_HVT U7484 ( .A1(n5856), .A3(n5437), .A2(n5857), .A4(n5858), .S0(
        n5766), .S1(n5302), .Y(n5855) );
  INVX0_HVT U7485 ( .A(n5796), .Y(n5862) );
  MUX41X1_HVT U7486 ( .A1(\ram[6][147] ), .A3(\ram[4][147] ), .A2(
        \ram[7][147] ), .A4(\ram[5][147] ), .S0(n5448), .S1(n5921), .Y(n8319)
         );
  MUX41X1_HVT U7487 ( .A1(\ram[13][228] ), .A3(\ram[15][228] ), .A2(
        \ram[12][228] ), .A4(\ram[14][228] ), .S0(n6652), .S1(n5864), .Y(n8641) );
  INVX0_HVT U7488 ( .A(n4988), .Y(n5987) );
  NBUFFX2_HVT U7489 ( .A(n6117), .Y(n6759) );
  MUX41X1_HVT U7490 ( .A1(\ram[11][160] ), .A3(\ram[9][160] ), .A2(
        \ram[10][160] ), .A4(\ram[8][160] ), .S0(n5903), .S1(n5229), .Y(n8370)
         );
  MUX41X1_HVT U7491 ( .A1(\ram[10][195] ), .A3(\ram[8][195] ), .A2(
        \ram[11][195] ), .A4(\ram[9][195] ), .S0(n7561), .S1(n6137), .Y(n8510)
         );
  INVX0_HVT U7492 ( .A(n5610), .Y(n7284) );
  NBUFFX2_HVT U7493 ( .A(n5164), .Y(n8880) );
  INVX0_HVT U7494 ( .A(n6123), .Y(n5947) );
  INVX0_HVT U7495 ( .A(n6416), .Y(n7567) );
  MUX41X1_HVT U7496 ( .A1(\ram[6][165] ), .A3(\ram[4][165] ), .A2(
        \ram[7][165] ), .A4(\ram[5][165] ), .S0(n7305), .S1(n8862), .Y(n8391)
         );
  IBUFFX2_HVT U7497 ( .A(n7665), .Y(n5893) );
  MUX41X1_HVT U7498 ( .A1(\ram[11][87] ), .A3(\ram[9][87] ), .A2(\ram[10][87] ), .A4(\ram[8][87] ), .S0(n5979), .S1(n5288), .Y(n8079) );
  INVX0_HVT U7499 ( .A(n7295), .Y(n7705) );
  MUX41X1_HVT U7500 ( .A1(\ram[7][241] ), .A3(\ram[5][241] ), .A2(
        \ram[6][241] ), .A4(\ram[4][241] ), .S0(n5878), .S1(n5792), .Y(n8693)
         );
  NBUFFX2_HVT U7501 ( .A(n4848), .Y(n7341) );
  MUX41X1_HVT U7502 ( .A1(\ram[3][237] ), .A3(\ram[1][237] ), .A2(
        \ram[2][237] ), .A4(\ram[0][237] ), .S0(n5638), .S1(n5882), .Y(n8678)
         );
  MUX41X1_HVT U7503 ( .A1(\ram[7][229] ), .A3(\ram[5][229] ), .A2(
        \ram[6][229] ), .A4(\ram[4][229] ), .S0(n5973), .S1(n5576), .Y(n8647)
         );
  MUX41X1_HVT U7504 ( .A1(\ram[7][217] ), .A3(\ram[5][217] ), .A2(
        \ram[6][217] ), .A4(\ram[4][217] ), .S0(n5884), .S1(n5228), .Y(n8599)
         );
  MUX41X1_HVT U7505 ( .A1(n7990), .A3(n7992), .A2(n7991), .A4(n7993), .S0(
        n5886), .S1(n5887), .Y(q[65]) );
  INVX0_HVT U7506 ( .A(n8785), .Y(n8789) );
  MUX41X1_HVT U7507 ( .A1(n8625), .A3(n8627), .A2(n8626), .A4(n8628), .S0(
        n5901), .S1(n5631), .Y(q[224]) );
  MUX41X1_HVT U7508 ( .A1(\ram[0][213] ), .A3(\ram[2][213] ), .A2(
        \ram[1][213] ), .A4(\ram[3][213] ), .S0(n5890), .S1(n5446), .Y(n8584)
         );
  MUX41X1_HVT U7509 ( .A1(n8517), .A3(n8519), .A2(n8518), .A4(n8520), .S0(
        n5891), .S1(n5369), .Y(q[197]) );
  MUX41X1_HVT U7510 ( .A1(\ram[0][155] ), .A3(\ram[2][155] ), .A2(
        \ram[1][155] ), .A4(\ram[3][155] ), .S0(n8820), .S1(n5512), .Y(n8352)
         );
  NBUFFX2_HVT U7511 ( .A(n4979), .Y(n8865) );
  MUX41X1_HVT U7512 ( .A1(\ram[11][183] ), .A3(\ram[9][183] ), .A2(
        \ram[10][183] ), .A4(\ram[8][183] ), .S0(n8788), .S1(n6384), .Y(n8462)
         );
  MUX41X1_HVT U7513 ( .A1(\ram[3][90] ), .A3(\ram[1][90] ), .A2(\ram[2][90] ), 
        .A4(\ram[0][90] ), .S0(n5985), .S1(n6638), .Y(n8093) );
  INVX0_HVT U7514 ( .A(n5920), .Y(n10108) );
  NBUFFX2_HVT U7515 ( .A(n7712), .Y(n6758) );
  MUX41X1_HVT U7516 ( .A1(\ram[3][201] ), .A3(\ram[1][201] ), .A2(
        \ram[2][201] ), .A4(\ram[0][201] ), .S0(n5640), .S1(n5767), .Y(n8536)
         );
  INVX0_HVT U7517 ( .A(n8851), .Y(n5905) );
  NBUFFX2_HVT U7518 ( .A(n7272), .Y(n7717) );
  MUX41X1_HVT U7519 ( .A1(\ram[12][215] ), .A3(\ram[14][215] ), .A2(
        \ram[13][215] ), .A4(\ram[15][215] ), .S0(n6020), .S1(n5907), .Y(n8589) );
  IBUFFX2_HVT U7520 ( .A(n5798), .Y(n8846) );
  INVX0_HVT U7521 ( .A(n6736), .Y(n6739) );
  INVX0_HVT U7522 ( .A(n5748), .Y(n10105) );
  MUX41X1_HVT U7523 ( .A1(\ram[3][158] ), .A3(\ram[1][158] ), .A2(
        \ram[2][158] ), .A4(\ram[0][158] ), .S0(n5829), .S1(n7711), .Y(n8364)
         );
  INVX1_HVT U7524 ( .A(n5916), .Y(n5908) );
  INVX1_HVT U7525 ( .A(n10099), .Y(n5909) );
  INVX1_HVT U7526 ( .A(n5908), .Y(n5910) );
  INVX1_HVT U7527 ( .A(n5913), .Y(n5914) );
  NBUFFX2_HVT U7528 ( .A(n5916), .Y(n5917) );
  NBUFFX2_HVT U7529 ( .A(n5916), .Y(n5918) );
  OAI21X1_HVT U7530 ( .A1(n5992), .A2(n5802), .A3(n5835), .Y(n5954) );
  AO21X1_HVT U7531 ( .A1(n60), .A2(n6037), .A3(n10381), .Y(n5920) );
  MUX41X1_HVT U7532 ( .A1(n8312), .A3(n8310), .A2(n8311), .A4(n8309), .S0(
        n5163), .S1(n8768), .Y(q[145]) );
  MUX41X1_HVT U7533 ( .A1(n8533), .A3(n8535), .A2(n8534), .A4(n8536), .S0(
        n5354), .S1(n5233), .Y(q[201]) );
  MUX41X1_HVT U7534 ( .A1(\ram[7][248] ), .A3(\ram[5][248] ), .A2(
        \ram[6][248] ), .A4(\ram[4][248] ), .S0(n5829), .S1(n5922), .Y(n8721)
         );
  NBUFFX2_HVT U7535 ( .A(n8809), .Y(n5923) );
  MUX41X1_HVT U7536 ( .A1(n8743), .A3(n8745), .A2(n8744), .A4(n8746), .S0(
        n5831), .S1(n7307), .Y(q[254]) );
  MUX41X1_HVT U7537 ( .A1(\ram[6][188] ), .A3(\ram[4][188] ), .A2(
        \ram[7][188] ), .A4(\ram[5][188] ), .S0(n7306), .S1(n6387), .Y(n8483)
         );
  MUX41X1_HVT U7538 ( .A1(\ram[11][6] ), .A3(\ram[9][6] ), .A2(\ram[10][6] ), 
        .A4(\ram[8][6] ), .S0(n7265), .S1(n4734), .Y(n7759) );
  MUX41X1_HVT U7539 ( .A1(\ram[11][165] ), .A3(\ram[9][165] ), .A2(
        \ram[10][165] ), .A4(\ram[8][165] ), .S0(n6414), .S1(n5826), .Y(n8390)
         );
  IBUFFX2_HVT U7540 ( .A(n7316), .Y(n8811) );
  INVX0_HVT U7541 ( .A(n5953), .Y(n7148) );
  IBUFFX2_HVT U7542 ( .A(n7326), .Y(n5937) );
  MUX41X1_HVT U7543 ( .A1(\ram[11][131] ), .A3(\ram[9][131] ), .A2(
        \ram[10][131] ), .A4(\ram[8][131] ), .S0(n6414), .S1(n7317), .Y(n8255)
         );
  MUX41X1_HVT U7544 ( .A1(\ram[3][131] ), .A3(\ram[1][131] ), .A2(
        \ram[2][131] ), .A4(\ram[0][131] ), .S0(n7277), .S1(n7266), .Y(n8257)
         );
  INVX0_HVT U7545 ( .A(n8776), .Y(n6400) );
  MUX41X1_HVT U7546 ( .A1(\ram[11][164] ), .A3(\ram[9][164] ), .A2(
        \ram[10][164] ), .A4(\ram[8][164] ), .S0(n7313), .S1(n4167), .Y(n8386)
         );
  IBUFFX2_HVT U7547 ( .A(n8773), .Y(n6641) );
  MUX41X1_HVT U7548 ( .A1(n5928), .A3(n5438), .A2(n5929), .A4(n5930), .S0(
        n8835), .S1(n5365), .Y(n5927) );
  NBUFFX2_HVT U7549 ( .A(n5314), .Y(n7579) );
  MUX41X1_HVT U7550 ( .A1(n8637), .A3(n8639), .A2(n8638), .A4(n8640), .S0(
        n5354), .S1(n5806), .Y(q[227]) );
  NBUFFX2_HVT U7551 ( .A(n6385), .Y(n8869) );
  INVX0_HVT U7552 ( .A(n7311), .Y(n5932) );
  INVX0_HVT U7553 ( .A(n10312), .Y(n5936) );
  MUX41X1_HVT U7554 ( .A1(\ram[11][223] ), .A3(\ram[9][223] ), .A2(
        \ram[10][223] ), .A4(\ram[8][223] ), .S0(n5937), .S1(n5813), .Y(n8622)
         );
  MUX41X1_HVT U7555 ( .A1(n8380), .A3(n8378), .A2(n8379), .A4(n8377), .S0(
        n7562), .S1(n5980), .Y(q[162]) );
  INVX0_HVT U7556 ( .A(n6123), .Y(n5938) );
  MUX41X1_HVT U7557 ( .A1(\ram[11][138] ), .A3(\ram[9][138] ), .A2(
        \ram[10][138] ), .A4(\ram[8][138] ), .S0(n5941), .S1(n5469), .Y(n8283)
         );
  INVX0_HVT U7558 ( .A(n8844), .Y(n5968) );
  INVX0_HVT U7559 ( .A(n8786), .Y(n8812) );
  INVX0_HVT U7560 ( .A(n6131), .Y(n6127) );
  INVX0_HVT U7561 ( .A(n5798), .Y(n5946) );
  MUX41X1_HVT U7562 ( .A1(n7950), .A3(n7948), .A2(n7949), .A4(n7947), .S0(
        n6416), .S1(n5801), .Y(q[54]) );
  INVX0_HVT U7563 ( .A(n5992), .Y(n60) );
  IBUFFX2_HVT U7564 ( .A(n5613), .Y(n8761) );
  MUX41X1_HVT U7565 ( .A1(n8449), .A3(n8451), .A2(n8450), .A4(n8452), .S0(
        n6397), .S1(n5868), .Y(q[180]) );
  MUX41X1_HVT U7566 ( .A1(n8361), .A3(n8363), .A2(n8362), .A4(n8364), .S0(
        n5111), .S1(n5959), .Y(q[158]) );
  NBUFFX2_HVT U7567 ( .A(n6411), .Y(n5962) );
  NOR2X0_HVT U7568 ( .A1(n6129), .A2(n7310), .Y(n51) );
  MUX41X1_HVT U7569 ( .A1(\ram[15][233] ), .A3(\ram[13][233] ), .A2(
        \ram[14][233] ), .A4(\ram[12][233] ), .S0(n5982), .S1(n5775), .Y(n5965) );
  INVX0_HVT U7570 ( .A(n8325), .Y(n6636) );
  MUX41X1_HVT U7571 ( .A1(\ram[15][6] ), .A3(\ram[13][6] ), .A2(\ram[14][6] ), 
        .A4(\ram[12][6] ), .S0(n6392), .S1(n5724), .Y(n7758) );
  MUX41X1_HVT U7572 ( .A1(\ram[11][201] ), .A3(\ram[10][201] ), .A2(
        \ram[9][201] ), .A4(\ram[8][201] ), .S0(n6638), .S1(n7561), .Y(n8534)
         );
  MUX41X1_HVT U7573 ( .A1(\ram[11][203] ), .A3(\ram[9][203] ), .A2(
        \ram[10][203] ), .A4(\ram[8][203] ), .S0(n5973), .S1(n6390), .Y(n8542)
         );
  MUX41X1_HVT U7574 ( .A1(\ram[11][231] ), .A3(\ram[9][231] ), .A2(
        \ram[10][231] ), .A4(\ram[8][231] ), .S0(n7557), .S1(n5302), .Y(n8654)
         );
  MUX41X1_HVT U7575 ( .A1(n8695), .A3(n8697), .A2(n8696), .A4(n8698), .S0(
        n5891), .S1(n7301), .Y(q[242]) );
  INVX1_HVT U7576 ( .A(n7714), .Y(n6752) );
  INVX0_HVT U7577 ( .A(n8771), .Y(n5995) );
  INVX0_HVT U7578 ( .A(n5504), .Y(n5985) );
  MUX41X1_HVT U7579 ( .A1(\ram[12][30] ), .A3(\ram[14][30] ), .A2(
        \ram[13][30] ), .A4(\ram[15][30] ), .S0(n5978), .S1(n5313), .Y(n5977)
         );
  MUX41X1_HVT U7580 ( .A1(\ram[14][232] ), .A3(\ram[12][232] ), .A2(
        \ram[15][232] ), .A4(\ram[13][232] ), .S0(n5975), .S1(n5950), .Y(n8657) );
  MUX41X1_HVT U7581 ( .A1(\ram[7][218] ), .A3(\ram[5][218] ), .A2(
        \ram[6][218] ), .A4(\ram[4][218] ), .S0(n5979), .S1(n5606), .Y(n8603)
         );
  NBUFFX2_HVT U7582 ( .A(n5478), .Y(n8860) );
  MUX41X1_HVT U7583 ( .A1(\ram[5][199] ), .A3(\ram[7][199] ), .A2(
        \ram[4][199] ), .A4(\ram[6][199] ), .S0(n7552), .S1(n6134), .Y(n8527)
         );
  INVX1_HVT U7584 ( .A(n7694), .Y(n6134) );
  MUX41X1_HVT U7585 ( .A1(\ram[3][161] ), .A3(\ram[1][161] ), .A2(
        \ram[2][161] ), .A4(\ram[0][161] ), .S0(n7571), .S1(n6251), .Y(n8376)
         );
  MUX41X1_HVT U7586 ( .A1(n8341), .A3(n8343), .A2(n8342), .A4(n8344), .S0(
        n5990), .S1(n5991), .Y(q[153]) );
  MUX41X1_HVT U7587 ( .A1(\ram[7][247] ), .A3(\ram[5][247] ), .A2(
        \ram[6][247] ), .A4(\ram[4][247] ), .S0(n7314), .S1(n6134), .Y(n8717)
         );
  NAND2X0_HVT U7588 ( .A1(n21), .A2(n51), .Y(n5992) );
  INVX0_HVT U7589 ( .A(n5090), .Y(n6391) );
  INVX0_HVT U7590 ( .A(n7673), .Y(n5997) );
  INVX0_HVT U7591 ( .A(n8839), .Y(n7147) );
  MUX41X1_HVT U7592 ( .A1(\ram[15][243] ), .A3(\ram[13][243] ), .A2(
        \ram[14][243] ), .A4(\ram[12][243] ), .S0(n5998), .S1(n5825), .Y(n8699) );
  MUX41X1_HVT U7593 ( .A1(\ram[15][132] ), .A3(\ram[13][132] ), .A2(
        \ram[14][132] ), .A4(\ram[12][132] ), .S0(n7265), .S1(n5730), .Y(n8258) );
  MUX41X1_HVT U7594 ( .A1(\ram[11][156] ), .A3(\ram[9][156] ), .A2(
        \ram[10][156] ), .A4(\ram[8][156] ), .S0(n7697), .S1(n5818), .Y(n8354)
         );
  MUX41X1_HVT U7595 ( .A1(n8304), .A3(n8302), .A2(n8305), .A4(n8303), .S0(
        n7562), .S1(n5344), .Y(q[143]) );
  MUX41X1_HVT U7596 ( .A1(\ram[2][205] ), .A3(\ram[0][205] ), .A2(
        \ram[3][205] ), .A4(\ram[1][205] ), .S0(n6136), .S1(n7686), .Y(n8552)
         );
  INVX0_HVT U7597 ( .A(n7343), .Y(n7286) );
  NAND2X0_HVT U7598 ( .A1(\ram[3][57] ), .A2(n7135), .Y(n5999) );
  NAND2X0_HVT U7599 ( .A1(n5999), .A2(n6000), .Y(n886) );
  INVX0_HVT U7600 ( .A(n7130), .Y(n7135) );
  MUX41X1_HVT U7601 ( .A1(\ram[3][247] ), .A3(\ram[1][247] ), .A2(
        \ram[2][247] ), .A4(\ram[0][247] ), .S0(n5976), .S1(n7709), .Y(n8718)
         );
  MUX41X1_HVT U7602 ( .A1(\ram[3][160] ), .A3(\ram[1][160] ), .A2(
        \ram[2][160] ), .A4(\ram[0][160] ), .S0(n6133), .S1(n7285), .Y(n8372)
         );
  MUX41X1_HVT U7603 ( .A1(\ram[11][13] ), .A3(\ram[9][13] ), .A2(\ram[10][13] ), .A4(\ram[8][13] ), .S0(n6133), .S1(n7285), .Y(n7787) );
  INVX0_HVT U7604 ( .A(n6639), .Y(n6037) );
  INVX0_HVT U7605 ( .A(n5087), .Y(n7333) );
  NBUFFX2_HVT U7606 ( .A(n8857), .Y(n6014) );
  INVX0_HVT U7607 ( .A(n6632), .Y(q[149]) );
  INVX1_HVT U7608 ( .A(n8326), .Y(n6634) );
  NBUFFX2_HVT U7609 ( .A(n7574), .Y(n6019) );
  INVX0_HVT U7610 ( .A(n5798), .Y(n6020) );
  MUX41X1_HVT U7611 ( .A1(\ram[11][63] ), .A3(\ram[9][63] ), .A2(\ram[10][63] ), .A4(\ram[8][63] ), .S0(n5608), .S1(n5508), .Y(n7983) );
  MUX41X1_HVT U7612 ( .A1(\ram[8][179] ), .A3(\ram[10][179] ), .A2(
        \ram[9][179] ), .A4(\ram[11][179] ), .S0(n8848), .S1(n6034), .Y(n8446)
         );
  MUX41X1_HVT U7613 ( .A1(\ram[1][54] ), .A3(\ram[3][54] ), .A2(\ram[0][54] ), 
        .A4(\ram[2][54] ), .S0(n5577), .S1(n7290), .Y(n7950) );
  NAND2X0_HVT U7614 ( .A1(n5620), .A2(n8), .Y(n6025) );
  NAND2X0_HVT U7615 ( .A1(\ram[3][5] ), .A2(n7124), .Y(n6026) );
  NAND2X0_HVT U7616 ( .A1(n5279), .A2(n9322), .Y(n6027) );
  NAND2X0_HVT U7617 ( .A1(n6026), .A2(n6027), .Y(n834) );
  INVX0_HVT U7618 ( .A(n7120), .Y(n7124) );
  MUX41X1_HVT U7619 ( .A1(n8349), .A3(n8350), .A2(n8351), .A4(n8352), .S0(
        n5344), .S1(n7302), .Y(q[155]) );
  INVX0_HVT U7620 ( .A(n8762), .Y(n7302) );
  MUX41X1_HVT U7621 ( .A1(\ram[11][33] ), .A3(\ram[9][33] ), .A2(\ram[10][33] ), .A4(\ram[8][33] ), .S0(n6746), .S1(n5792), .Y(n7864) );
  INVX0_HVT U7622 ( .A(N28), .Y(n7558) );
  INVX0_HVT U7623 ( .A(n7144), .Y(n8851) );
  NBUFFX2_HVT U7624 ( .A(n8852), .Y(n6032) );
  INVX0_HVT U7625 ( .A(n6123), .Y(n6033) );
  MUX41X1_HVT U7626 ( .A1(\ram[7][203] ), .A3(\ram[5][203] ), .A2(
        \ram[6][203] ), .A4(\ram[4][203] ), .S0(n5638), .S1(n5002), .Y(n8543)
         );
  IBUFFX2_HVT U7627 ( .A(n10286), .Y(n6629) );
  IBUFFX2_HVT U7628 ( .A(n4971), .Y(n10284) );
  IBUFFX2_HVT U7629 ( .A(n4971), .Y(n10283) );
  IBUFFX2_HVT U7630 ( .A(n5761), .Y(n6627) );
  IBUFFX2_HVT U7631 ( .A(n4972), .Y(n6628) );
  INVX0_HVT U7632 ( .A(n8767), .Y(n6396) );
  NBUFFX2_HVT U7633 ( .A(n10233), .Y(n6039) );
  NBUFFX2_HVT U7634 ( .A(n10227), .Y(n6040) );
  NBUFFX2_HVT U7635 ( .A(n10234), .Y(n6041) );
  NBUFFX2_HVT U7636 ( .A(n10235), .Y(n6042) );
  INVX0_HVT U7637 ( .A(n10222), .Y(n6046) );
  INVX0_HVT U7638 ( .A(n10222), .Y(n6047) );
  INVX1_HVT U7639 ( .A(n6046), .Y(n6048) );
  INVX1_HVT U7640 ( .A(n6047), .Y(n6049) );
  INVX1_HVT U7641 ( .A(n6076), .Y(n6051) );
  INVX0_HVT U7642 ( .A(n10223), .Y(n6052) );
  INVX0_HVT U7643 ( .A(n10223), .Y(n6053) );
  INVX1_HVT U7644 ( .A(n6053), .Y(n6055) );
  INVX0_HVT U7645 ( .A(n10224), .Y(n6056) );
  INVX0_HVT U7646 ( .A(n10224), .Y(n6057) );
  INVX1_HVT U7647 ( .A(n6056), .Y(n6058) );
  INVX1_HVT U7648 ( .A(n6057), .Y(n6059) );
  INVX1_HVT U7649 ( .A(n6094), .Y(n6062) );
  INVX0_HVT U7650 ( .A(n10231), .Y(n6063) );
  INVX0_HVT U7651 ( .A(n10231), .Y(n6064) );
  INVX1_HVT U7652 ( .A(n6063), .Y(n6065) );
  INVX1_HVT U7653 ( .A(n6094), .Y(n6067) );
  INVX1_HVT U7654 ( .A(n6063), .Y(n6071) );
  INVX1_HVT U7655 ( .A(n6052), .Y(n6072) );
  INVX1_HVT U7656 ( .A(n6094), .Y(n6073) );
  INVX1_HVT U7657 ( .A(n6063), .Y(n6074) );
  INVX1_HVT U7658 ( .A(n6053), .Y(n6075) );
  INVX0_HVT U7659 ( .A(n10234), .Y(n6076) );
  INVX0_HVT U7660 ( .A(n10234), .Y(n6077) );
  INVX1_HVT U7661 ( .A(n6076), .Y(n6078) );
  INVX0_HVT U7662 ( .A(n10233), .Y(n6080) );
  INVX0_HVT U7663 ( .A(n10233), .Y(n6081) );
  INVX1_HVT U7664 ( .A(n6080), .Y(n6082) );
  INVX1_HVT U7665 ( .A(n6064), .Y(n6084) );
  INVX0_HVT U7666 ( .A(n10230), .Y(n6086) );
  INVX1_HVT U7667 ( .A(n6086), .Y(n6087) );
  INVX1_HVT U7668 ( .A(n6091), .Y(n6088) );
  INVX1_HVT U7669 ( .A(n6097), .Y(n6089) );
  INVX1_HVT U7670 ( .A(n6098), .Y(n6090) );
  INVX0_HVT U7671 ( .A(n10232), .Y(n6091) );
  INVX1_HVT U7672 ( .A(n6057), .Y(n6092) );
  INVX1_HVT U7673 ( .A(n6091), .Y(n6093) );
  INVX0_HVT U7674 ( .A(n10229), .Y(n6094) );
  INVX1_HVT U7675 ( .A(n6094), .Y(n6095) );
  INVX1_HVT U7676 ( .A(n6086), .Y(n6096) );
  INVX0_HVT U7677 ( .A(n10228), .Y(n6097) );
  INVX0_HVT U7678 ( .A(n10228), .Y(n6098) );
  INVX1_HVT U7679 ( .A(n6064), .Y(n6102) );
  INVX1_HVT U7680 ( .A(n6056), .Y(n6105) );
  INVX0_HVT U7681 ( .A(n10226), .Y(n6106) );
  INVX1_HVT U7682 ( .A(n6106), .Y(n6107) );
  INVX1_HVT U7683 ( .A(n6106), .Y(n6108) );
  INVX0_HVT U7684 ( .A(n10225), .Y(n6109) );
  INVX0_HVT U7685 ( .A(n10225), .Y(n6110) );
  INVX0_HVT U7686 ( .A(n6077), .Y(n10222) );
  INVX0_HVT U7687 ( .A(n6043), .Y(n10223) );
  INVX0_HVT U7688 ( .A(n6103), .Y(n10224) );
  MUX41X1_HVT U7689 ( .A1(n8540), .A3(n8538), .A2(n8539), .A4(n8537), .S0(
        n6259), .S1(n5237), .Y(q[202]) );
  MUX41X1_HVT U7690 ( .A1(\ram[7][221] ), .A3(\ram[5][221] ), .A2(
        \ram[6][221] ), .A4(\ram[4][221] ), .S0(n4993), .S1(n5767), .Y(n8615)
         );
  INVX0_HVT U7691 ( .A(n10379), .Y(n7573) );
  NAND2X0_HVT U7692 ( .A1(\ram[6][40] ), .A2(n5174), .Y(n6121) );
  NAND2X0_HVT U7693 ( .A1(n9210), .A2(n9427), .Y(n6122) );
  NAND2X0_HVT U7694 ( .A1(n6121), .A2(n6122), .Y(n1637) );
  MUX21X1_HVT U7695 ( .A1(\ram[15][253] ), .A2(\ram[13][253] ), .S0(n7673), 
        .Y(n6124) );
  MUX41X1_HVT U7696 ( .A1(\ram[15][242] ), .A3(\ram[13][242] ), .A2(
        \ram[14][242] ), .A4(\ram[12][242] ), .S0(n6128), .S1(n7709), .Y(n8695) );
  INVX0_HVT U7697 ( .A(n8774), .Y(n6381) );
  MUX41X1_HVT U7698 ( .A1(n8440), .A3(n8438), .A2(n8439), .A4(n8437), .S0(
        n6130), .S1(n5896), .Y(q[177]) );
  MUX41X1_HVT U7699 ( .A1(\ram[11][32] ), .A3(\ram[9][32] ), .A2(\ram[10][32] ), .A4(\ram[8][32] ), .S0(n6133), .S1(n6134), .Y(n7860) );
  INVX0_HVT U7700 ( .A(n7721), .Y(n10235) );
  MUX41X1_HVT U7701 ( .A1(\ram[15][214] ), .A3(\ram[13][214] ), .A2(
        \ram[14][214] ), .A4(\ram[12][214] ), .S0(n7265), .S1(n5153), .Y(n8585) );
  MUX41X1_HVT U7702 ( .A1(\ram[7][181] ), .A3(\ram[5][181] ), .A2(
        \ram[6][181] ), .A4(\ram[4][181] ), .S0(n5817), .S1(n6138), .Y(n8455)
         );
  NAND2X0_HVT U7703 ( .A1(\ram[4][0] ), .A2(n4961), .Y(n6139) );
  NAND2X0_HVT U7704 ( .A1(n6219), .A2(n9306), .Y(n6140) );
  NAND2X0_HVT U7705 ( .A1(n6139), .A2(n6140), .Y(n1085) );
  INVX0_HVT U7706 ( .A(n6158), .Y(n6141) );
  NBUFFX2_HVT U7707 ( .A(n6152), .Y(n6143) );
  NBUFFX2_HVT U7708 ( .A(n6147), .Y(n6144) );
  NBUFFX2_HVT U7709 ( .A(n4697), .Y(n6148) );
  NBUFFX2_HVT U7710 ( .A(n6147), .Y(n6149) );
  NBUFFX2_HVT U7711 ( .A(n5129), .Y(n6150) );
  NBUFFX2_HVT U7712 ( .A(n5129), .Y(n6151) );
  NBUFFX2_HVT U7713 ( .A(n4572), .Y(n6153) );
  NBUFFX2_HVT U7714 ( .A(n4572), .Y(n6154) );
  NBUFFX2_HVT U7715 ( .A(n6155), .Y(n6156) );
  NBUFFX2_HVT U7716 ( .A(n6155), .Y(n6157) );
  INVX1_HVT U7717 ( .A(n6141), .Y(n6165) );
  INVX1_HVT U7718 ( .A(n6141), .Y(n6166) );
  IBUFFX2_HVT U7719 ( .A(n6165), .Y(n6167) );
  IBUFFX2_HVT U7720 ( .A(n6165), .Y(n6168) );
  IBUFFX2_HVT U7721 ( .A(n5459), .Y(n6179) );
  INVX0_HVT U7722 ( .A(n6218), .Y(n6219) );
  INVX0_HVT U7723 ( .A(n10306), .Y(n10305) );
  NBUFFX2_HVT U7724 ( .A(n6186), .Y(n6187) );
  NBUFFX2_HVT U7725 ( .A(n6186), .Y(n6188) );
  NBUFFX2_HVT U7726 ( .A(n6186), .Y(n6189) );
  NBUFFX2_HVT U7727 ( .A(n6186), .Y(n6190) );
  NBUFFX2_HVT U7728 ( .A(n6186), .Y(n6191) );
  INVX1_HVT U7729 ( .A(n6224), .Y(n6192) );
  INVX1_HVT U7730 ( .A(n6229), .Y(n6194) );
  INVX0_HVT U7731 ( .A(n10291), .Y(n6196) );
  INVX1_HVT U7732 ( .A(n6218), .Y(n6197) );
  INVX0_HVT U7733 ( .A(n10291), .Y(n6199) );
  INVX1_HVT U7734 ( .A(n6199), .Y(n6200) );
  INVX1_HVT U7735 ( .A(n6213), .Y(n6203) );
  INVX0_HVT U7736 ( .A(n10296), .Y(n6204) );
  INVX1_HVT U7737 ( .A(n6204), .Y(n6205) );
  INVX1_HVT U7738 ( .A(n6204), .Y(n6206) );
  INVX0_HVT U7739 ( .A(n10297), .Y(n6207) );
  INVX1_HVT U7740 ( .A(n6207), .Y(n6208) );
  INVX1_HVT U7741 ( .A(n6239), .Y(n6209) );
  INVX0_HVT U7742 ( .A(n10296), .Y(n6210) );
  INVX1_HVT U7743 ( .A(n6204), .Y(n6211) );
  INVX0_HVT U7744 ( .A(n10295), .Y(n6213) );
  INVX1_HVT U7745 ( .A(n6213), .Y(n6214) );
  INVX1_HVT U7746 ( .A(n6213), .Y(n6215) );
  INVX0_HVT U7747 ( .A(n10298), .Y(n6218) );
  INVX0_HVT U7748 ( .A(n10299), .Y(n6221) );
  INVX1_HVT U7749 ( .A(n6221), .Y(n6222) );
  INVX1_HVT U7750 ( .A(n6224), .Y(n6223) );
  INVX0_HVT U7751 ( .A(n10298), .Y(n6224) );
  INVX0_HVT U7752 ( .A(n10295), .Y(n6225) );
  INVX1_HVT U7753 ( .A(n6225), .Y(n6227) );
  INVX0_HVT U7754 ( .A(n10292), .Y(n6229) );
  INVX1_HVT U7755 ( .A(n6229), .Y(n6230) );
  INVX1_HVT U7756 ( .A(n6207), .Y(n6231) );
  INVX0_HVT U7757 ( .A(n10294), .Y(n6232) );
  INVX1_HVT U7758 ( .A(n6239), .Y(n6234) );
  INVX0_HVT U7759 ( .A(n10292), .Y(n6235) );
  INVX1_HVT U7760 ( .A(n6235), .Y(n6236) );
  INVX1_HVT U7761 ( .A(n6235), .Y(n6237) );
  INVX0_HVT U7762 ( .A(n10293), .Y(n6238) );
  INVX0_HVT U7763 ( .A(n10293), .Y(n6239) );
  INVX1_HVT U7764 ( .A(n6238), .Y(n6240) );
  INVX1_HVT U7765 ( .A(n6239), .Y(n6241) );
  INVX1_HVT U7766 ( .A(n6210), .Y(n6242) );
  INVX0_HVT U7767 ( .A(n10299), .Y(n6244) );
  INVX1_HVT U7768 ( .A(n6244), .Y(n6245) );
  INVX1_HVT U7769 ( .A(n6244), .Y(n6246) );
  INVX0_HVT U7770 ( .A(n10299), .Y(n6247) );
  INVX0_HVT U7771 ( .A(n10298), .Y(n6248) );
  INVX1_HVT U7772 ( .A(n6248), .Y(n6250) );
  INVX0_HVT U7773 ( .A(n6218), .Y(n10291) );
  MUX41X1_HVT U7774 ( .A1(\ram[15][77] ), .A3(\ram[13][77] ), .A2(
        \ram[14][77] ), .A4(\ram[12][77] ), .S0(n5817), .S1(n6251), .Y(n8038)
         );
  MUX41X1_HVT U7775 ( .A1(\ram[11][135] ), .A3(\ram[9][135] ), .A2(
        \ram[10][135] ), .A4(\ram[8][135] ), .S0(n7546), .S1(n5722), .Y(n8271)
         );
  MUX41X1_HVT U7776 ( .A1(\ram[14][133] ), .A3(\ram[12][133] ), .A2(
        \ram[15][133] ), .A4(\ram[13][133] ), .S0(n5961), .S1(n6253), .Y(n8262) );
  MUX41X1_HVT U7777 ( .A1(n8323), .A3(n8321), .A2(n8324), .A4(n8322), .S0(
        n5925), .S1(n6643), .Y(q[148]) );
  MUX41X1_HVT U7778 ( .A1(\ram[11][15] ), .A3(\ram[9][15] ), .A2(\ram[10][15] ), .A4(\ram[8][15] ), .S0(n5985), .S1(n5899), .Y(n7795) );
  MUX41X1_HVT U7779 ( .A1(\ram[11][232] ), .A3(\ram[10][232] ), .A2(
        \ram[9][232] ), .A4(\ram[8][232] ), .S0(n6390), .S1(n6389), .Y(n8658)
         );
  INVX0_HVT U7780 ( .A(n5936), .Y(n10308) );
  MUX41X1_HVT U7781 ( .A1(n8050), .A3(n8052), .A2(n8051), .A4(n8053), .S0(
        n7276), .S1(n6257), .Y(q[80]) );
  NBUFFX2_HVT U7782 ( .A(n10376), .Y(n6258) );
  INVX0_HVT U7783 ( .A(n6639), .Y(n10376) );
  AO21X1_HVT U7784 ( .A1(n50), .A2(n6258), .A3(n10381), .Y(n7729) );
  MUX41X1_HVT U7785 ( .A1(\ram[3][226] ), .A3(\ram[1][226] ), .A2(
        \ram[2][226] ), .A4(\ram[0][226] ), .S0(n6412), .S1(n7716), .Y(n8636)
         );
  NAND2X0_HVT U7786 ( .A1(\ram[2][54] ), .A2(n7205), .Y(n6260) );
  NAND2X0_HVT U7787 ( .A1(n6326), .A2(n9469), .Y(n6261) );
  NAND2X0_HVT U7788 ( .A1(n6260), .A2(n6261), .Y(n627) );
  NBUFFX2_HVT U7789 ( .A(n6262), .Y(n6263) );
  NBUFFX2_HVT U7790 ( .A(n6262), .Y(n6264) );
  NBUFFX2_HVT U7791 ( .A(n6262), .Y(n6265) );
  NBUFFX2_HVT U7792 ( .A(n6262), .Y(n6266) );
  INVX0_HVT U7793 ( .A(n10319), .Y(n6269) );
  INVX1_HVT U7794 ( .A(n6269), .Y(n6270) );
  INVX1_HVT U7795 ( .A(n6276), .Y(n6271) );
  INVX0_HVT U7796 ( .A(n10319), .Y(n6273) );
  INVX1_HVT U7797 ( .A(n6273), .Y(n6274) );
  INVX0_HVT U7798 ( .A(n10322), .Y(n6276) );
  INVX0_HVT U7799 ( .A(n10326), .Y(n6277) );
  INVX1_HVT U7800 ( .A(n6276), .Y(n6278) );
  INVX1_HVT U7801 ( .A(n6299), .Y(n6280) );
  INVX1_HVT U7802 ( .A(n6292), .Y(n6281) );
  INVX0_HVT U7803 ( .A(n10326), .Y(n6282) );
  INVX0_HVT U7804 ( .A(n10326), .Y(n6283) );
  INVX1_HVT U7805 ( .A(n6277), .Y(n6286) );
  INVX1_HVT U7806 ( .A(n6306), .Y(n6288) );
  INVX1_HVT U7807 ( .A(n6300), .Y(n6289) );
  INVX0_HVT U7808 ( .A(n10327), .Y(n6292) );
  INVX0_HVT U7809 ( .A(n10327), .Y(n6293) );
  INVX1_HVT U7810 ( .A(n6323), .Y(n6295) );
  INVX1_HVT U7811 ( .A(n6317), .Y(n6296) );
  INVX0_HVT U7812 ( .A(n10325), .Y(n6297) );
  INVX1_HVT U7813 ( .A(n6297), .Y(n6298) );
  INVX0_HVT U7814 ( .A(n10325), .Y(n6299) );
  INVX0_HVT U7815 ( .A(n10325), .Y(n6300) );
  INVX1_HVT U7816 ( .A(n6299), .Y(n6301) );
  INVX1_HVT U7817 ( .A(n6300), .Y(n6302) );
  INVX0_HVT U7818 ( .A(n10319), .Y(n6303) );
  INVX1_HVT U7819 ( .A(n6303), .Y(n6304) );
  INVX1_HVT U7820 ( .A(n6303), .Y(n6305) );
  INVX0_HVT U7821 ( .A(n10327), .Y(n6306) );
  INVX0_HVT U7822 ( .A(n10322), .Y(n6307) );
  INVX1_HVT U7823 ( .A(n6306), .Y(n6308) );
  INVX1_HVT U7824 ( .A(n6307), .Y(n6309) );
  INVX1_HVT U7825 ( .A(n6297), .Y(n6310) );
  INVX1_HVT U7826 ( .A(n6324), .Y(n6311) );
  INVX0_HVT U7827 ( .A(n10323), .Y(n6312) );
  INVX1_HVT U7828 ( .A(n6312), .Y(n6313) );
  INVX1_HVT U7829 ( .A(n6307), .Y(n6315) );
  INVX1_HVT U7830 ( .A(n6307), .Y(n6316) );
  INVX0_HVT U7831 ( .A(n10321), .Y(n6317) );
  INVX1_HVT U7832 ( .A(n6317), .Y(n6318) );
  INVX0_HVT U7833 ( .A(n10321), .Y(n6320) );
  INVX1_HVT U7834 ( .A(n6320), .Y(n6321) );
  INVX1_HVT U7835 ( .A(n6320), .Y(n6322) );
  INVX0_HVT U7836 ( .A(n10320), .Y(n6323) );
  INVX0_HVT U7837 ( .A(n10320), .Y(n6324) );
  INVX1_HVT U7838 ( .A(n6323), .Y(n6325) );
  INVX1_HVT U7839 ( .A(n6324), .Y(n6326) );
  INVX0_HVT U7840 ( .A(n7198), .Y(n7205) );
  INVX0_HVT U7841 ( .A(n6292), .Y(n10319) );
  INVX0_HVT U7842 ( .A(n10330), .Y(n10329) );
  NAND2X0_HVT U7843 ( .A1(\ram[12][142] ), .A2(n6560), .Y(n6327) );
  NAND2X0_HVT U7844 ( .A1(n4550), .A2(n9735), .Y(n6328) );
  NAND2X0_HVT U7845 ( .A1(n6327), .A2(n6328), .Y(n3275) );
  INVX0_HVT U7846 ( .A(n10130), .Y(n6329) );
  INVX0_HVT U7847 ( .A(n10130), .Y(n6330) );
  INVX0_HVT U7848 ( .A(n10130), .Y(n6331) );
  NBUFFX2_HVT U7849 ( .A(n4305), .Y(n6332) );
  NBUFFX2_HVT U7850 ( .A(n6331), .Y(n6333) );
  NBUFFX2_HVT U7851 ( .A(n6336), .Y(n6334) );
  NBUFFX2_HVT U7852 ( .A(n4305), .Y(n6335) );
  NBUFFX2_HVT U7853 ( .A(n6336), .Y(n6337) );
  NBUFFX2_HVT U7854 ( .A(n6336), .Y(n6338) );
  NBUFFX2_HVT U7855 ( .A(n6336), .Y(n6339) );
  INVX0_HVT U7856 ( .A(n10131), .Y(n6340) );
  NBUFFX2_HVT U7857 ( .A(n6340), .Y(n6341) );
  NBUFFX2_HVT U7858 ( .A(n6340), .Y(n6342) );
  NBUFFX2_HVT U7859 ( .A(n6350), .Y(n6343) );
  NBUFFX2_HVT U7860 ( .A(n6331), .Y(n6344) );
  INVX0_HVT U7861 ( .A(n10131), .Y(n6345) );
  NBUFFX2_HVT U7862 ( .A(n6345), .Y(n6346) );
  NBUFFX2_HVT U7863 ( .A(n6345), .Y(n6347) );
  NBUFFX2_HVT U7864 ( .A(n6340), .Y(n6348) );
  NBUFFX2_HVT U7865 ( .A(n6345), .Y(n6349) );
  INVX0_HVT U7866 ( .A(n10132), .Y(n6350) );
  INVX0_HVT U7867 ( .A(n10132), .Y(n6351) );
  NBUFFX2_HVT U7868 ( .A(n6350), .Y(n6352) );
  NBUFFX2_HVT U7869 ( .A(n6350), .Y(n6353) );
  NBUFFX2_HVT U7870 ( .A(n6351), .Y(n6354) );
  NBUFFX2_HVT U7871 ( .A(n6351), .Y(n6355) );
  INVX0_HVT U7872 ( .A(n6356), .Y(n6357) );
  INVX0_HVT U7873 ( .A(n6356), .Y(n6358) );
  INVX0_HVT U7874 ( .A(n6356), .Y(n6359) );
  INVX0_HVT U7875 ( .A(n6356), .Y(n6360) );
  INVX0_HVT U7876 ( .A(n10131), .Y(n6361) );
  INVX0_HVT U7877 ( .A(n6356), .Y(n6362) );
  INVX0_HVT U7878 ( .A(n10132), .Y(n6363) );
  INVX1_HVT U7879 ( .A(n6329), .Y(n6364) );
  INVX1_HVT U7880 ( .A(n6330), .Y(n6374) );
  INVX0_HVT U7881 ( .A(n10134), .Y(n10133) );
  INVX0_HVT U7882 ( .A(n6044), .Y(n10229) );
  INVX0_HVT U7883 ( .A(n6080), .Y(n10228) );
  IBUFFX2_HVT U7884 ( .A(n8753), .Y(n8764) );
  MUX41X1_HVT U7885 ( .A1(\ram[11][25] ), .A3(\ram[9][25] ), .A2(\ram[10][25] ), .A4(\ram[8][25] ), .S0(n6412), .S1(n7348), .Y(n7833) );
  NBUFFX2_HVT U7886 ( .A(n6754), .Y(n8773) );
  MUX41X1_HVT U7887 ( .A1(\ram[15][125] ), .A3(\ram[13][125] ), .A2(
        \ram[14][125] ), .A4(\ram[12][125] ), .S0(n6405), .S1(n6384), .Y(n8230) );
  IBUFFX2_HVT U7888 ( .A(n8769), .Y(n7702) );
  INVX0_HVT U7889 ( .A(n49), .Y(n10130) );
  MUX41X1_HVT U7890 ( .A1(\ram[14][79] ), .A3(\ram[12][79] ), .A2(
        \ram[15][79] ), .A4(\ram[13][79] ), .S0(n7281), .S1(n6748), .Y(n8046)
         );
  MUX41X1_HVT U7891 ( .A1(n8580), .A3(n8578), .A2(n8579), .A4(n8577), .S0(
        n6130), .S1(n6388), .Y(q[212]) );
  INVX0_HVT U7892 ( .A(n10302), .Y(n10294) );
  INVX0_HVT U7893 ( .A(n10302), .Y(n10293) );
  INVX0_HVT U7894 ( .A(n10302), .Y(n10292) );
  MUX41X1_HVT U7895 ( .A1(\ram[3][10] ), .A3(\ram[1][10] ), .A2(\ram[2][10] ), 
        .A4(\ram[0][10] ), .S0(n6405), .S1(n7576), .Y(n7777) );
  NBUFFX2_HVT U7896 ( .A(n5797), .Y(n6394) );
  MUX41X1_HVT U7897 ( .A1(n8188), .A3(n8186), .A2(n8189), .A4(n8187), .S0(
        n5097), .S1(n5308), .Y(q[114]) );
  MUX41X1_HVT U7898 ( .A1(n7824), .A3(n7826), .A2(n7825), .A4(n7827), .S0(
        n6397), .S1(n5624), .Y(q[23]) );
  MUX41X1_HVT U7899 ( .A1(n7796), .A3(n7794), .A2(n7797), .A4(n7795), .S0(
        n8762), .S1(n5624), .Y(q[15]) );
  MUX41X1_HVT U7900 ( .A1(n7790), .A3(n7792), .A2(n7791), .A4(n7793), .S0(
        n6651), .S1(n5359), .Y(q[14]) );
  MUX41X1_HVT U7901 ( .A1(n7778), .A3(n7780), .A2(n7779), .A4(n7781), .S0(
        n6399), .S1(n6400), .Y(q[11]) );
  MUX41X1_HVT U7902 ( .A1(n7775), .A3(n7777), .A2(n7774), .A4(n7776), .S0(
        n7349), .S1(n5162), .Y(q[10]) );
  MUX41X1_HVT U7903 ( .A1(n6402), .A3(n5440), .A2(n6403), .A4(n6404), .S0(
        n6405), .S1(n6740), .Y(n6401) );
  NBUFFX2_HVT U7904 ( .A(n6892), .Y(n6409) );
  MUX41X1_HVT U7905 ( .A1(\ram[15][201] ), .A3(\ram[13][201] ), .A2(
        \ram[14][201] ), .A4(\ram[12][201] ), .S0(n6412), .S1(n5653), .Y(n8533) );
  MUX41X1_HVT U7906 ( .A1(\ram[15][159] ), .A3(\ram[13][159] ), .A2(
        \ram[14][159] ), .A4(\ram[12][159] ), .S0(n7571), .S1(n7289), .Y(n8365) );
  INVX0_HVT U7907 ( .A(n7814), .Y(n6649) );
  NBUFFX2_HVT U7908 ( .A(n10182), .Y(n6418) );
  NBUFFX2_HVT U7909 ( .A(n10182), .Y(n6419) );
  NBUFFX2_HVT U7910 ( .A(n10180), .Y(n6420) );
  NBUFFX2_HVT U7911 ( .A(n10179), .Y(n6421) );
  NBUFFX2_HVT U7912 ( .A(n10179), .Y(n6422) );
  INVX1_HVT U7913 ( .A(n6426), .Y(n6424) );
  INVX0_HVT U7914 ( .A(n10181), .Y(n6426) );
  INVX1_HVT U7915 ( .A(n6429), .Y(n6427) );
  INVX1_HVT U7916 ( .A(n6426), .Y(n6428) );
  INVX0_HVT U7917 ( .A(n10179), .Y(n6429) );
  INVX1_HVT U7918 ( .A(n6464), .Y(n6430) );
  INVX1_HVT U7919 ( .A(n6429), .Y(n6431) );
  INVX0_HVT U7920 ( .A(n10180), .Y(n6432) );
  INVX1_HVT U7921 ( .A(n6432), .Y(n6433) );
  INVX1_HVT U7922 ( .A(n6432), .Y(n6434) );
  INVX0_HVT U7923 ( .A(n10181), .Y(n6435) );
  INVX0_HVT U7924 ( .A(n10181), .Y(n6436) );
  INVX1_HVT U7925 ( .A(n6435), .Y(n6437) );
  INVX1_HVT U7926 ( .A(n6436), .Y(n6438) );
  INVX1_HVT U7927 ( .A(n6436), .Y(n6439) );
  INVX1_HVT U7928 ( .A(n6426), .Y(n6440) );
  INVX0_HVT U7929 ( .A(n10186), .Y(n6441) );
  INVX1_HVT U7930 ( .A(n6441), .Y(n6443) );
  INVX1_HVT U7931 ( .A(n6442), .Y(n6444) );
  INVX1_HVT U7932 ( .A(n6450), .Y(n6445) );
  INVX1_HVT U7933 ( .A(n6441), .Y(n6446) );
  INVX1_HVT U7934 ( .A(n6441), .Y(n6447) );
  INVX1_HVT U7935 ( .A(n6451), .Y(n6448) );
  INVX1_HVT U7936 ( .A(n6465), .Y(n6449) );
  INVX0_HVT U7937 ( .A(n10186), .Y(n6450) );
  INVX0_HVT U7938 ( .A(n10186), .Y(n6451) );
  INVX1_HVT U7939 ( .A(n6451), .Y(n6452) );
  INVX1_HVT U7940 ( .A(n6451), .Y(n6453) );
  INVX1_HVT U7941 ( .A(n6441), .Y(n6454) );
  INVX1_HVT U7942 ( .A(n6464), .Y(n6455) );
  INVX1_HVT U7943 ( .A(n6461), .Y(n6456) );
  INVX1_HVT U7944 ( .A(n6458), .Y(n6457) );
  INVX0_HVT U7945 ( .A(n10185), .Y(n6458) );
  INVX1_HVT U7946 ( .A(n6458), .Y(n6459) );
  INVX1_HVT U7947 ( .A(n6465), .Y(n6460) );
  INVX0_HVT U7948 ( .A(n10184), .Y(n6461) );
  INVX1_HVT U7949 ( .A(n6458), .Y(n6462) );
  INVX1_HVT U7950 ( .A(n6461), .Y(n6463) );
  INVX0_HVT U7951 ( .A(n10183), .Y(n6464) );
  INVX0_HVT U7952 ( .A(n10183), .Y(n6465) );
  INVX1_HVT U7953 ( .A(n6464), .Y(n6466) );
  INVX1_HVT U7954 ( .A(n6465), .Y(n6467) );
  INVX1_HVT U7955 ( .A(n6442), .Y(n6468) );
  INVX1_HVT U7956 ( .A(n6450), .Y(n6469) );
  INVX1_HVT U7957 ( .A(n6429), .Y(n6470) );
  INVX1_HVT U7958 ( .A(n6450), .Y(n6471) );
  INVX1_HVT U7959 ( .A(n6435), .Y(n6472) );
  INVX1_HVT U7960 ( .A(n6429), .Y(n6473) );
  INVX1_HVT U7961 ( .A(n6461), .Y(n6474) );
  INVX0_HVT U7962 ( .A(n10182), .Y(n6475) );
  INVX1_HVT U7963 ( .A(n6436), .Y(n6476) );
  INVX1_HVT U7964 ( .A(n6442), .Y(n6478) );
  INVX1_HVT U7965 ( .A(n6435), .Y(n6479) );
  INVX0_HVT U7966 ( .A(n7722), .Y(n10179) );
  INVX0_HVT U7967 ( .A(n6475), .Y(n10180) );
  INVX0_HVT U7968 ( .A(n6423), .Y(n10181) );
  MUX41X1_HVT U7969 ( .A1(n6481), .A3(n6482), .A2(n6483), .A4(n6484), .S0(
        n5975), .S1(n6551), .Y(n6480) );
  NBUFFX2_HVT U7970 ( .A(n4507), .Y(n6486) );
  NBUFFX2_HVT U7971 ( .A(n4507), .Y(n6487) );
  NBUFFX2_HVT U7972 ( .A(n6485), .Y(n6488) );
  NBUFFX2_HVT U7973 ( .A(n6485), .Y(n6489) );
  NBUFFX2_HVT U7974 ( .A(n6492), .Y(n6490) );
  INVX1_HVT U7975 ( .A(n6498), .Y(n6494) );
  INVX1_HVT U7976 ( .A(n6515), .Y(n6495) );
  INVX1_HVT U7977 ( .A(n6499), .Y(n6497) );
  INVX0_HVT U7978 ( .A(n10353), .Y(n6498) );
  INVX0_HVT U7979 ( .A(n10353), .Y(n6499) );
  INVX1_HVT U7980 ( .A(n6498), .Y(n6500) );
  INVX1_HVT U7981 ( .A(n6499), .Y(n6501) );
  INVX1_HVT U7982 ( .A(n6499), .Y(n6502) );
  INVX0_HVT U7983 ( .A(n10359), .Y(n6504) );
  INVX0_HVT U7984 ( .A(n10359), .Y(n6505) );
  INVX1_HVT U7985 ( .A(n6505), .Y(n6507) );
  INVX0_HVT U7986 ( .A(n10357), .Y(n6508) );
  INVX1_HVT U7987 ( .A(n6516), .Y(n6510) );
  INVX0_HVT U7988 ( .A(n10354), .Y(n6511) );
  INVX0_HVT U7989 ( .A(n10354), .Y(n6512) );
  INVX0_HVT U7990 ( .A(n10355), .Y(n6515) );
  INVX0_HVT U7991 ( .A(n10355), .Y(n6516) );
  INVX1_HVT U7992 ( .A(n6515), .Y(n6517) );
  INVX1_HVT U7993 ( .A(n6516), .Y(n6518) );
  INVX0_HVT U7994 ( .A(n10352), .Y(n6519) );
  INVX1_HVT U7995 ( .A(n6537), .Y(n6520) );
  INVX0_HVT U7996 ( .A(n10352), .Y(n6522) );
  INVX0_HVT U7997 ( .A(n10358), .Y(n6527) );
  INVX0_HVT U7998 ( .A(n10358), .Y(n6530) );
  INVX0_HVT U7999 ( .A(n10359), .Y(n6531) );
  INVX1_HVT U8000 ( .A(n6531), .Y(n6533) );
  INVX0_HVT U8001 ( .A(n10358), .Y(n6534) );
  INVX0_HVT U8002 ( .A(n10355), .Y(n6537) );
  INVX1_HVT U8003 ( .A(n6537), .Y(n6539) );
  INVX1_HVT U8004 ( .A(n6505), .Y(n6542) );
  INVX1_HVT U8005 ( .A(n6505), .Y(n6543) );
  INVX1_HVT U8006 ( .A(n6531), .Y(n6545) );
  INVX1_HVT U8007 ( .A(n6531), .Y(n6548) );
  INVX0_HVT U8008 ( .A(n7720), .Y(n10352) );
  INVX0_HVT U8009 ( .A(n6491), .Y(n10353) );
  INVX0_HVT U8010 ( .A(n6522), .Y(n10357) );
  INVX0_HVT U8011 ( .A(n6519), .Y(n10354) );
  INVX0_HVT U8012 ( .A(n4438), .Y(n10355) );
  INVX0_HVT U8013 ( .A(n10360), .Y(n10358) );
  INVX0_HVT U8014 ( .A(n6504), .Y(n10356) );
  INVX0_HVT U8015 ( .A(n7722), .Y(n10190) );
  NBUFFX2_HVT U8016 ( .A(n10136), .Y(n6556) );
  NBUFFX2_HVT U8017 ( .A(n10138), .Y(n6557) );
  NBUFFX2_HVT U8018 ( .A(n10141), .Y(n6558) );
  NBUFFX2_HVT U8019 ( .A(n10145), .Y(n6559) );
  NBUFFX2_HVT U8020 ( .A(n10136), .Y(n6560) );
  INVX1_HVT U8021 ( .A(n6585), .Y(n6561) );
  INVX1_HVT U8022 ( .A(n6607), .Y(n6562) );
  INVX0_HVT U8023 ( .A(n10135), .Y(n6563) );
  INVX0_HVT U8024 ( .A(n10135), .Y(n6564) );
  INVX1_HVT U8025 ( .A(n6563), .Y(n6565) );
  INVX1_HVT U8026 ( .A(n6623), .Y(n6568) );
  INVX0_HVT U8027 ( .A(n10144), .Y(n6569) );
  INVX1_HVT U8028 ( .A(n6569), .Y(n6571) );
  INVX1_HVT U8029 ( .A(n6563), .Y(n6572) );
  INVX0_HVT U8030 ( .A(n10139), .Y(n6574) );
  INVX0_HVT U8031 ( .A(n10139), .Y(n6575) );
  INVX1_HVT U8032 ( .A(n6575), .Y(n6577) );
  INVX1_HVT U8033 ( .A(n6608), .Y(n6579) );
  INVX0_HVT U8034 ( .A(n10145), .Y(n6581) );
  INVX0_HVT U8035 ( .A(n10137), .Y(n6582) );
  INVX1_HVT U8036 ( .A(n6582), .Y(n6584) );
  INVX0_HVT U8037 ( .A(n10137), .Y(n6585) );
  INVX0_HVT U8038 ( .A(n10137), .Y(n6586) );
  INVX1_HVT U8039 ( .A(n6585), .Y(n6587) );
  INVX0_HVT U8040 ( .A(n10143), .Y(n6589) );
  INVX1_HVT U8041 ( .A(n6589), .Y(n6591) );
  INVX1_HVT U8042 ( .A(n6575), .Y(n6592) );
  INVX0_HVT U8043 ( .A(n4510), .Y(n6593) );
  INVX0_HVT U8044 ( .A(n10136), .Y(n6594) );
  INVX1_HVT U8045 ( .A(n6593), .Y(n6595) );
  INVX1_HVT U8046 ( .A(n6600), .Y(n6597) );
  INVX1_HVT U8047 ( .A(n6599), .Y(n6598) );
  INVX0_HVT U8048 ( .A(n10141), .Y(n6599) );
  INVX0_HVT U8049 ( .A(n10141), .Y(n6600) );
  INVX1_HVT U8050 ( .A(n6599), .Y(n6601) );
  INVX1_HVT U8051 ( .A(n6600), .Y(n6602) );
  INVX0_HVT U8052 ( .A(n10142), .Y(n6603) );
  INVX0_HVT U8053 ( .A(n10142), .Y(n6604) );
  INVX1_HVT U8054 ( .A(n6603), .Y(n6605) );
  INVX0_HVT U8055 ( .A(n10138), .Y(n6607) );
  INVX0_HVT U8056 ( .A(n10143), .Y(n6608) );
  INVX1_HVT U8057 ( .A(n6607), .Y(n6609) );
  INVX1_HVT U8058 ( .A(n6608), .Y(n6610) );
  INVX0_HVT U8059 ( .A(n10143), .Y(n6614) );
  INVX1_HVT U8060 ( .A(n6614), .Y(n6615) );
  INVX1_HVT U8061 ( .A(n6614), .Y(n6616) );
  INVX1_HVT U8062 ( .A(n6581), .Y(n6618) );
  INVX1_HVT U8063 ( .A(n6603), .Y(n6620) );
  INVX1_HVT U8064 ( .A(n6582), .Y(n6621) );
  INVX1_HVT U8065 ( .A(n6581), .Y(n6622) );
  INVX0_HVT U8066 ( .A(n10144), .Y(n6623) );
  INVX1_HVT U8067 ( .A(n6593), .Y(n6624) );
  INVX1_HVT U8068 ( .A(n6623), .Y(n6625) );
  INVX0_HVT U8069 ( .A(n6586), .Y(n10146) );
  MUX41X1_HVT U8070 ( .A1(\ram[7][40] ), .A3(\ram[5][40] ), .A2(\ram[6][40] ), 
        .A4(\ram[4][40] ), .S0(n5794), .S1(n6740), .Y(n7893) );
  INVX0_HVT U8071 ( .A(n10190), .Y(n10188) );
  MUX41X1_HVT U8072 ( .A1(\ram[15][59] ), .A3(\ram[13][59] ), .A2(
        \ram[14][59] ), .A4(\ram[12][59] ), .S0(n4993), .S1(n5933), .Y(n7966)
         );
  INVX0_HVT U8073 ( .A(n6647), .Y(q[20]) );
  INVX0_HVT U8074 ( .A(n7815), .Y(n6648) );
  MUX41X1_HVT U8075 ( .A1(\ram[11][139] ), .A3(\ram[9][139] ), .A2(
        \ram[10][139] ), .A4(\ram[8][139] ), .S0(n7572), .S1(n4885), .Y(n8287)
         );
  MUX41X1_HVT U8076 ( .A1(\ram[11][194] ), .A3(\ram[9][194] ), .A2(
        \ram[10][194] ), .A4(\ram[8][194] ), .S0(n5966), .S1(n7146), .Y(n8506)
         );
  MUX41X1_HVT U8077 ( .A1(n6635), .A3(n6636), .A2(n6633), .A4(n6634), .S0(
        n6756), .S1(n6752), .Y(n6632) );
  MUX41X1_HVT U8078 ( .A1(\ram[12][212] ), .A3(\ram[14][212] ), .A2(
        \ram[13][212] ), .A4(\ram[15][212] ), .S0(n6642), .S1(n6387), .Y(n8577) );
  MUX41X1_HVT U8079 ( .A1(\ram[15][184] ), .A3(\ram[13][184] ), .A2(
        \ram[14][184] ), .A4(\ram[12][184] ), .S0(n6645), .S1(n6655), .Y(n8465) );
  MUX41X1_HVT U8080 ( .A1(n6649), .A3(n6550), .A2(n6480), .A4(n6648), .S0(
        n8753), .S1(n6752), .Y(n6647) );
  MUX41X1_HVT U8081 ( .A1(n7806), .A3(n7808), .A2(n7807), .A4(n7809), .S0(
        n6651), .S1(n7271), .Y(q[18]) );
  INVX0_HVT U8082 ( .A(n5646), .Y(n7556) );
  MUX41X1_HVT U8083 ( .A1(n7762), .A3(n7764), .A2(n7763), .A4(n7765), .S0(
        n7349), .S1(n7271), .Y(q[7]) );
  DELLN2X2_HVT U8084 ( .A(n5581), .Y(n7351) );
  INVX0_HVT U8085 ( .A(n5090), .Y(n7275) );
  MUX41X1_HVT U8086 ( .A1(\ram[3][105] ), .A3(\ram[1][105] ), .A2(
        \ram[2][105] ), .A4(\ram[0][105] ), .S0(n6654), .S1(n5133), .Y(n8153)
         );
  MUX41X1_HVT U8087 ( .A1(\ram[15][80] ), .A3(\ram[13][80] ), .A2(
        \ram[14][80] ), .A4(\ram[12][80] ), .S0(n5449), .S1(n5001), .Y(n8050)
         );
  IBUFFX2_HVT U8088 ( .A(n5114), .Y(n7083) );
  NBUFFX2_HVT U8089 ( .A(n5311), .Y(n7350) );
  INVX0_HVT U8090 ( .A(n6752), .Y(n6751) );
  NAND2X0_HVT U8091 ( .A1(\ram[6][192] ), .A2(n5174), .Y(n6664) );
  NAND2X0_HVT U8092 ( .A1(n9247), .A2(n9893), .Y(n6665) );
  NAND2X0_HVT U8093 ( .A1(n6664), .A2(n6665), .Y(n1789) );
  INVX0_HVT U8094 ( .A(n9242), .Y(n9247) );
  MUX41X1_HVT U8095 ( .A1(\ram[15][26] ), .A3(\ram[13][26] ), .A2(
        \ram[14][26] ), .A4(\ram[12][26] ), .S0(n8781), .S1(n7289), .Y(n7836)
         );
  INVX0_HVT U8096 ( .A(n5478), .Y(n6740) );
  INVX1_HVT U8097 ( .A(n6713), .Y(n6666) );
  INVX1_HVT U8098 ( .A(n6708), .Y(n6669) );
  INVX1_HVT U8099 ( .A(n6709), .Y(n6670) );
  INVX0_HVT U8100 ( .A(n10362), .Y(n6671) );
  INVX1_HVT U8101 ( .A(n6687), .Y(n6673) );
  INVX0_HVT U8102 ( .A(n10363), .Y(n6674) );
  INVX0_HVT U8103 ( .A(n10363), .Y(n6675) );
  INVX1_HVT U8104 ( .A(n6674), .Y(n6676) );
  INVX1_HVT U8105 ( .A(n6675), .Y(n6677) );
  INVX0_HVT U8106 ( .A(n6712), .Y(n6679) );
  INVX0_HVT U8107 ( .A(n10364), .Y(n6680) );
  INVX0_HVT U8108 ( .A(n6680), .Y(n6682) );
  INVX0_HVT U8109 ( .A(n10362), .Y(n6683) );
  INVX0_HVT U8110 ( .A(n6687), .Y(n6685) );
  INVX0_HVT U8111 ( .A(n10365), .Y(n6686) );
  INVX0_HVT U8112 ( .A(n10365), .Y(n6687) );
  INVX0_HVT U8113 ( .A(n6687), .Y(n6689) );
  INVX0_HVT U8114 ( .A(n6709), .Y(n6690) );
  INVX0_HVT U8115 ( .A(n4399), .Y(n6691) );
  INVX0_HVT U8116 ( .A(n10366), .Y(n6693) );
  INVX1_HVT U8117 ( .A(n6693), .Y(n6694) );
  INVX0_HVT U8118 ( .A(n6693), .Y(n6695) );
  INVX0_HVT U8119 ( .A(n6674), .Y(n6696) );
  INVX0_HVT U8120 ( .A(n10371), .Y(n6697) );
  INVX1_HVT U8121 ( .A(n6697), .Y(n6698) );
  INVX0_HVT U8122 ( .A(n6683), .Y(n6699) );
  INVX0_HVT U8123 ( .A(n10366), .Y(n6700) );
  INVX1_HVT U8124 ( .A(n6700), .Y(n6701) );
  INVX0_HVT U8125 ( .A(n6700), .Y(n6702) );
  INVX0_HVT U8126 ( .A(n10365), .Y(n6703) );
  INVX1_HVT U8127 ( .A(n6703), .Y(n6704) );
  INVX0_HVT U8128 ( .A(n6703), .Y(n6705) );
  INVX0_HVT U8129 ( .A(n6686), .Y(n6707) );
  INVX0_HVT U8130 ( .A(n10369), .Y(n6708) );
  INVX0_HVT U8131 ( .A(n10369), .Y(n6709) );
  INVX1_HVT U8132 ( .A(n6708), .Y(n6710) );
  INVX0_HVT U8133 ( .A(n6709), .Y(n6711) );
  INVX0_HVT U8134 ( .A(n10366), .Y(n6713) );
  INVX0_HVT U8135 ( .A(n6713), .Y(n6715) );
  INVX0_HVT U8136 ( .A(n6680), .Y(n6717) );
  INVX0_HVT U8137 ( .A(n10371), .Y(n6718) );
  INVX0_HVT U8138 ( .A(n10364), .Y(n6719) );
  INVX1_HVT U8139 ( .A(n6718), .Y(n6720) );
  INVX0_HVT U8140 ( .A(n6719), .Y(n6721) );
  INVX1_HVT U8141 ( .A(n6675), .Y(n6722) );
  INVX0_HVT U8142 ( .A(n6697), .Y(n6723) );
  INVX1_HVT U8143 ( .A(n6719), .Y(n6725) );
  INVX0_HVT U8144 ( .A(n6724), .Y(n6726) );
  NBUFFX2_HVT U8145 ( .A(n6727), .Y(n6728) );
  NBUFFX2_HVT U8146 ( .A(n6727), .Y(n6729) );
  NBUFFX2_HVT U8147 ( .A(n6727), .Y(n6730) );
  NBUFFX2_HVT U8148 ( .A(n6727), .Y(n6731) );
  INVX0_HVT U8149 ( .A(n6691), .Y(n10362) );
  INVX0_HVT U8150 ( .A(n10374), .Y(n10363) );
  INVX0_HVT U8151 ( .A(n6724), .Y(n10364) );
  INVX0_HVT U8152 ( .A(n10373), .Y(n10365) );
  INVX0_HVT U8153 ( .A(n10374), .Y(n10366) );
  INVX0_HVT U8154 ( .A(n7730), .Y(n10367) );
  INVX0_HVT U8155 ( .A(n6700), .Y(n10368) );
  INVX0_HVT U8156 ( .A(n10373), .Y(n10369) );
  INVX0_HVT U8157 ( .A(n6691), .Y(n10370) );
  INVX0_HVT U8158 ( .A(n6724), .Y(n10371) );
  INVX0_HVT U8159 ( .A(n7730), .Y(n10372) );
  MUX41X1_HVT U8160 ( .A1(\ram[11][221] ), .A3(\ram[9][221] ), .A2(
        \ram[10][221] ), .A4(\ram[8][221] ), .S0(n8782), .S1(n6745), .Y(n8614)
         );
  MUX41X1_HVT U8161 ( .A1(\ram[11][71] ), .A3(\ram[9][71] ), .A2(\ram[10][71] ), .A4(\ram[8][71] ), .S0(n5738), .S1(n5127), .Y(n8015) );
  MUX41X1_HVT U8162 ( .A1(\ram[15][219] ), .A3(\ram[13][219] ), .A2(
        \ram[14][219] ), .A4(\ram[12][219] ), .S0(n5155), .S1(n6740), .Y(n8605) );
  MUX41X1_HVT U8163 ( .A1(\ram[14][75] ), .A3(\ram[12][75] ), .A2(
        \ram[15][75] ), .A4(\ram[13][75] ), .S0(n5448), .S1(n7555), .Y(n8030)
         );
  MUX41X1_HVT U8164 ( .A1(\ram[15][227] ), .A3(\ram[13][227] ), .A2(
        \ram[14][227] ), .A4(\ram[12][227] ), .S0(n5743), .S1(n6734), .Y(n8637) );
  MUX41X1_HVT U8165 ( .A1(\ram[15][248] ), .A3(\ram[13][248] ), .A2(
        \ram[14][248] ), .A4(\ram[12][248] ), .S0(n7561), .S1(n6745), .Y(n8719) );
  MUX41X1_HVT U8166 ( .A1(\ram[3][236] ), .A3(\ram[1][236] ), .A2(
        \ram[2][236] ), .A4(\ram[0][236] ), .S0(n6746), .S1(n5488), .Y(n8674)
         );
  MUX41X1_HVT U8167 ( .A1(\ram[15][94] ), .A3(\ram[13][94] ), .A2(
        \ram[14][94] ), .A4(\ram[12][94] ), .S0(n7277), .S1(n6732), .Y(n8106)
         );
  INVX0_HVT U8168 ( .A(n8752), .Y(n8755) );
  MUX41X1_HVT U8169 ( .A1(\ram[0][77] ), .A3(\ram[2][77] ), .A2(\ram[1][77] ), 
        .A4(\ram[3][77] ), .S0(n5630), .S1(n5656), .Y(n8041) );
  MUX41X1_HVT U8170 ( .A1(\ram[0][127] ), .A3(\ram[2][127] ), .A2(
        \ram[1][127] ), .A4(\ram[3][127] ), .S0(n8804), .S1(n6748), .Y(n8241)
         );
  MUX41X1_HVT U8171 ( .A1(\ram[15][41] ), .A3(\ram[13][41] ), .A2(
        \ram[14][41] ), .A4(\ram[12][41] ), .S0(n7572), .S1(n7142), .Y(n7895)
         );
  IBUFFX2_HVT U8172 ( .A(n8753), .Y(n7543) );
  MUX41X1_HVT U8173 ( .A1(\ram[14][152] ), .A3(\ram[12][152] ), .A2(
        \ram[15][152] ), .A4(\ram[13][152] ), .S0(n7556), .S1(n6137), .Y(n8337) );
  NBUFFX2_HVT U8174 ( .A(n5797), .Y(n7687) );
  MUX41X1_HVT U8175 ( .A1(\ram[3][180] ), .A3(\ram[1][180] ), .A2(
        \ram[2][180] ), .A4(\ram[0][180] ), .S0(n5903), .S1(n6656), .Y(n8452)
         );
  MUX41X1_HVT U8176 ( .A1(\ram[3][163] ), .A3(\ram[1][163] ), .A2(
        \ram[2][163] ), .A4(\ram[0][163] ), .S0(n7557), .S1(n7576), .Y(n8384)
         );
  MUX41X1_HVT U8177 ( .A1(\ram[12][220] ), .A3(\ram[14][220] ), .A2(
        \ram[13][220] ), .A4(\ram[15][220] ), .S0(n7321), .S1(n8907), .Y(n8609) );
  MUX41X1_HVT U8178 ( .A1(\ram[1][220] ), .A3(\ram[3][220] ), .A2(
        \ram[0][220] ), .A4(\ram[2][220] ), .S0(n7141), .S1(n5567), .Y(n8612)
         );
  NBUFFX2_HVT U8179 ( .A(n4930), .Y(n6762) );
  IBUFFX2_HVT U8180 ( .A(n7664), .Y(n7149) );
  IBUFFX2_HVT U8181 ( .A(n7719), .Y(n6769) );
  NBUFFX2_HVT U8182 ( .A(n6769), .Y(n6770) );
  NBUFFX2_HVT U8183 ( .A(n6769), .Y(n6771) );
  NBUFFX2_HVT U8184 ( .A(n6769), .Y(n6772) );
  NBUFFX2_HVT U8185 ( .A(n6769), .Y(n6773) );
  NBUFFX2_HVT U8186 ( .A(n6769), .Y(n6774) );
  INVX0_HVT U8187 ( .A(n10150), .Y(n6775) );
  INVX1_HVT U8188 ( .A(n6775), .Y(n6776) );
  INVX1_HVT U8189 ( .A(n6775), .Y(n6777) );
  INVX0_HVT U8190 ( .A(n10151), .Y(n6778) );
  INVX1_HVT U8191 ( .A(n6778), .Y(n6779) );
  INVX1_HVT U8192 ( .A(n6778), .Y(n6780) );
  INVX0_HVT U8193 ( .A(n10150), .Y(n6781) );
  INVX1_HVT U8194 ( .A(n6781), .Y(n6782) );
  INVX1_HVT U8195 ( .A(n6781), .Y(n6783) );
  INVX0_HVT U8196 ( .A(n10151), .Y(n6784) );
  INVX1_HVT U8197 ( .A(n6784), .Y(n6785) );
  INVX1_HVT U8198 ( .A(n6778), .Y(n6786) );
  INVX1_HVT U8199 ( .A(n6818), .Y(n6788) );
  INVX1_HVT U8200 ( .A(n6784), .Y(n6789) );
  INVX0_HVT U8201 ( .A(n10156), .Y(n6790) );
  INVX1_HVT U8202 ( .A(n6795), .Y(n6791) );
  INVX1_HVT U8203 ( .A(n6790), .Y(n6792) );
  INVX1_HVT U8204 ( .A(n6790), .Y(n6793) );
  INVX1_HVT U8205 ( .A(n6790), .Y(n6794) );
  INVX0_HVT U8206 ( .A(n10156), .Y(n6795) );
  INVX1_HVT U8207 ( .A(n6795), .Y(n6796) );
  INVX1_HVT U8208 ( .A(n6795), .Y(n6797) );
  INVX1_HVT U8209 ( .A(n6807), .Y(n6798) );
  INVX1_HVT U8210 ( .A(n6804), .Y(n6799) );
  INVX0_HVT U8211 ( .A(n10160), .Y(n6800) );
  INVX0_HVT U8212 ( .A(n10159), .Y(n6803) );
  INVX0_HVT U8213 ( .A(n10159), .Y(n6804) );
  INVX1_HVT U8214 ( .A(n6804), .Y(n6806) );
  INVX0_HVT U8215 ( .A(n10158), .Y(n6807) );
  INVX1_HVT U8216 ( .A(n6807), .Y(n6808) );
  INVX1_HVT U8217 ( .A(n6815), .Y(n6809) );
  INVX1_HVT U8218 ( .A(n6807), .Y(n6810) );
  INVX0_HVT U8219 ( .A(n10158), .Y(n6812) );
  INVX1_HVT U8220 ( .A(n6812), .Y(n6813) );
  INVX1_HVT U8221 ( .A(n6812), .Y(n6814) );
  INVX0_HVT U8222 ( .A(n10153), .Y(n6815) );
  INVX0_HVT U8223 ( .A(n10154), .Y(n6816) );
  INVX1_HVT U8224 ( .A(n6818), .Y(n6817) );
  INVX0_HVT U8225 ( .A(n10154), .Y(n6818) );
  INVX1_HVT U8226 ( .A(n6818), .Y(n6819) );
  INVX1_HVT U8227 ( .A(n6803), .Y(n6820) );
  INVX1_HVT U8228 ( .A(n6804), .Y(n6821) );
  INVX1_HVT U8229 ( .A(n6781), .Y(n6822) );
  INVX1_HVT U8230 ( .A(n6784), .Y(n6824) );
  INVX1_HVT U8231 ( .A(n6775), .Y(n6825) );
  INVX0_HVT U8232 ( .A(n10163), .Y(n10150) );
  INVX0_HVT U8233 ( .A(n10163), .Y(n10151) );
  INVX0_HVT U8234 ( .A(n10161), .Y(n10160) );
  INVX0_HVT U8235 ( .A(n10162), .Y(n10153) );
  INVX0_HVT U8236 ( .A(n10162), .Y(n10154) );
  INVX1_HVT U8237 ( .A(n6882), .Y(n6830) );
  INVX1_HVT U8238 ( .A(n6875), .Y(n6832) );
  INVX0_HVT U8239 ( .A(n10335), .Y(n6833) );
  INVX0_HVT U8240 ( .A(n10335), .Y(n6834) );
  INVX0_HVT U8241 ( .A(n10337), .Y(n6837) );
  INVX0_HVT U8242 ( .A(n10343), .Y(n6838) );
  INVX1_HVT U8243 ( .A(n6837), .Y(n6839) );
  INVX1_HVT U8244 ( .A(n6838), .Y(n6840) );
  INVX1_HVT U8245 ( .A(n6863), .Y(n6842) );
  INVX0_HVT U8246 ( .A(n10340), .Y(n6843) );
  INVX1_HVT U8247 ( .A(n6862), .Y(n6844) );
  INVX1_HVT U8248 ( .A(n6879), .Y(n6845) );
  INVX1_HVT U8249 ( .A(n6879), .Y(n6846) );
  INVX1_HVT U8250 ( .A(n6862), .Y(n6850) );
  INVX0_HVT U8251 ( .A(n10344), .Y(n6852) );
  INVX1_HVT U8252 ( .A(n6851), .Y(n6853) );
  INVX1_HVT U8253 ( .A(n6852), .Y(n6854) );
  INVX1_HVT U8254 ( .A(n6875), .Y(n6859) );
  INVX1_HVT U8255 ( .A(n6837), .Y(n6860) );
  INVX0_HVT U8256 ( .A(n10336), .Y(n6862) );
  INVX0_HVT U8257 ( .A(n10336), .Y(n6863) );
  INVX1_HVT U8258 ( .A(n6848), .Y(n6866) );
  INVX1_HVT U8259 ( .A(n6852), .Y(n6869) );
  INVX0_HVT U8260 ( .A(n10338), .Y(n6870) );
  INVX1_HVT U8261 ( .A(n6848), .Y(n6872) );
  INVX1_HVT U8262 ( .A(n6843), .Y(n6873) );
  INVX1_HVT U8263 ( .A(n6863), .Y(n6874) );
  INVX0_HVT U8264 ( .A(n10339), .Y(n6875) );
  INVX0_HVT U8265 ( .A(n10339), .Y(n6876) );
  INVX0_HVT U8266 ( .A(n10341), .Y(n6879) );
  INVX1_HVT U8267 ( .A(n6879), .Y(n6880) );
  INVX0_HVT U8268 ( .A(n10338), .Y(n6882) );
  INVX1_HVT U8269 ( .A(n6838), .Y(n6883) );
  INVX1_HVT U8270 ( .A(n6882), .Y(n6884) );
  NBUFFX2_HVT U8271 ( .A(n10343), .Y(n6886) );
  NBUFFX2_HVT U8272 ( .A(n10341), .Y(n6887) );
  NBUFFX2_HVT U8273 ( .A(n10335), .Y(n6888) );
  NBUFFX2_HVT U8274 ( .A(n10338), .Y(n6889) );
  NBUFFX2_HVT U8275 ( .A(n10337), .Y(n6890) );
  INVX0_HVT U8276 ( .A(n10346), .Y(n10335) );
  INVX0_HVT U8277 ( .A(n6843), .Y(n10336) );
  INVX0_HVT U8278 ( .A(n10345), .Y(n10338) );
  INVX0_HVT U8279 ( .A(n6826), .Y(n10339) );
  INVX0_HVT U8280 ( .A(n10345), .Y(n10337) );
  MUX41X1_HVT U8281 ( .A1(n8164), .A3(n8162), .A2(n8165), .A4(n8163), .S0(
        n5097), .S1(n5369), .Y(q[108]) );
  MUX41X1_HVT U8282 ( .A1(\ram[7][175] ), .A3(\ram[5][175] ), .A2(
        \ram[6][175] ), .A4(\ram[4][175] ), .S0(n5741), .S1(n7285), .Y(n8431)
         );
  MUX41X1_HVT U8283 ( .A1(\ram[11][246] ), .A3(\ram[9][246] ), .A2(
        \ram[10][246] ), .A4(\ram[8][246] ), .S0(n5878), .S1(n5465), .Y(n8712)
         );
  MUX41X1_HVT U8284 ( .A1(\ram[15][46] ), .A3(\ram[13][46] ), .A2(
        \ram[14][46] ), .A4(\ram[12][46] ), .S0(n5741), .S1(n7317), .Y(n7915)
         );
  MUX41X1_HVT U8285 ( .A1(\ram[12][49] ), .A3(\ram[14][49] ), .A2(
        \ram[13][49] ), .A4(\ram[15][49] ), .S0(n8838), .S1(n5807), .Y(n7927)
         );
  NBUFFX2_HVT U8286 ( .A(n10258), .Y(n6895) );
  NBUFFX2_HVT U8287 ( .A(n10264), .Y(n6896) );
  NBUFFX2_HVT U8288 ( .A(n10259), .Y(n6897) );
  NBUFFX2_HVT U8289 ( .A(n10257), .Y(n6898) );
  NBUFFX2_HVT U8290 ( .A(n10265), .Y(n6899) );
  INVX0_HVT U8291 ( .A(n10257), .Y(n6903) );
  INVX1_HVT U8292 ( .A(n6903), .Y(n6904) );
  INVX1_HVT U8293 ( .A(n6903), .Y(n6905) );
  INVX0_HVT U8294 ( .A(n10258), .Y(n6906) );
  INVX1_HVT U8295 ( .A(n6940), .Y(n6908) );
  INVX0_HVT U8296 ( .A(n10258), .Y(n6909) );
  INVX1_HVT U8297 ( .A(n6909), .Y(n6910) );
  INVX0_HVT U8298 ( .A(n10259), .Y(n6911) );
  INVX1_HVT U8299 ( .A(n6911), .Y(n6912) );
  INVX1_HVT U8300 ( .A(n6911), .Y(n6913) );
  INVX0_HVT U8301 ( .A(n10268), .Y(n6914) );
  INVX0_HVT U8302 ( .A(n10268), .Y(n6915) );
  INVX1_HVT U8303 ( .A(n6914), .Y(n6916) );
  INVX1_HVT U8304 ( .A(n6915), .Y(n6917) );
  INVX1_HVT U8305 ( .A(n6915), .Y(n6918) );
  INVX1_HVT U8306 ( .A(n6914), .Y(n6919) );
  INVX1_HVT U8307 ( .A(n6962), .Y(n6920) );
  INVX1_HVT U8308 ( .A(n6961), .Y(n6921) );
  INVX0_HVT U8309 ( .A(n10266), .Y(n6922) );
  INVX0_HVT U8310 ( .A(n10266), .Y(n6923) );
  INVX1_HVT U8311 ( .A(n6949), .Y(n6926) );
  INVX1_HVT U8312 ( .A(n6949), .Y(n6927) );
  INVX0_HVT U8313 ( .A(n10260), .Y(n6928) );
  INVX0_HVT U8314 ( .A(n10263), .Y(n6929) );
  INVX1_HVT U8315 ( .A(n6928), .Y(n6930) );
  INVX1_HVT U8316 ( .A(n6929), .Y(n6931) );
  INVX0_HVT U8317 ( .A(n10260), .Y(n6932) );
  INVX1_HVT U8318 ( .A(n6928), .Y(n6933) );
  INVX1_HVT U8319 ( .A(n6932), .Y(n6934) );
  INVX0_HVT U8320 ( .A(n10266), .Y(n6935) );
  INVX1_HVT U8321 ( .A(n6935), .Y(n6936) );
  INVX0_HVT U8322 ( .A(n10261), .Y(n6940) );
  INVX0_HVT U8323 ( .A(n10261), .Y(n6941) );
  INVX1_HVT U8324 ( .A(n6940), .Y(n6942) );
  INVX1_HVT U8325 ( .A(n6941), .Y(n6943) );
  INVX1_HVT U8326 ( .A(n6941), .Y(n6944) );
  INVX0_HVT U8327 ( .A(n10263), .Y(n6945) );
  INVX1_HVT U8328 ( .A(n6945), .Y(n6946) );
  INVX1_HVT U8329 ( .A(n6945), .Y(n6947) );
  INVX1_HVT U8330 ( .A(n6948), .Y(n6950) );
  INVX1_HVT U8331 ( .A(n6949), .Y(n6951) );
  INVX1_HVT U8332 ( .A(n6948), .Y(n6954) );
  INVX1_HVT U8333 ( .A(n6948), .Y(n6955) );
  INVX1_HVT U8334 ( .A(n6929), .Y(n6956) );
  INVX1_HVT U8335 ( .A(n6932), .Y(n6957) );
  INVX0_HVT U8336 ( .A(n10264), .Y(n6958) );
  INVX1_HVT U8337 ( .A(n6958), .Y(n6959) );
  INVX1_HVT U8338 ( .A(n6958), .Y(n6960) );
  INVX0_HVT U8339 ( .A(n10260), .Y(n6961) );
  INVX0_HVT U8340 ( .A(n10264), .Y(n6962) );
  INVX1_HVT U8341 ( .A(n6961), .Y(n6963) );
  INVX1_HVT U8342 ( .A(n6962), .Y(n6964) );
  INVX0_HVT U8343 ( .A(n6923), .Y(n10257) );
  INVX0_HVT U8344 ( .A(n7733), .Y(n10258) );
  INVX0_HVT U8345 ( .A(n6922), .Y(n10259) );
  INVX0_HVT U8346 ( .A(n7733), .Y(n10266) );
  INVX0_HVT U8347 ( .A(n6906), .Y(n10267) );
  INVX0_HVT U8348 ( .A(n6935), .Y(n10262) );
  INVX0_HVT U8349 ( .A(n6901), .Y(n10263) );
  INVX0_HVT U8350 ( .A(n6900), .Y(n10264) );
  INVX0_HVT U8351 ( .A(n10127), .Y(n6967) );
  INVX0_HVT U8352 ( .A(n10127), .Y(n6968) );
  NBUFFX2_HVT U8353 ( .A(n6969), .Y(n6971) );
  NBUFFX2_HVT U8354 ( .A(n6969), .Y(n6972) );
  NBUFFX2_HVT U8355 ( .A(n6970), .Y(n6973) );
  NBUFFX2_HVT U8356 ( .A(n6970), .Y(n6974) );
  NBUFFX2_HVT U8357 ( .A(n6980), .Y(n6975) );
  NBUFFX2_HVT U8358 ( .A(n4776), .Y(n6976) );
  NBUFFX2_HVT U8359 ( .A(n6986), .Y(n6977) );
  NBUFFX2_HVT U8360 ( .A(n6986), .Y(n6978) );
  INVX0_HVT U8361 ( .A(n6997), .Y(n6979) );
  INVX0_HVT U8362 ( .A(n4374), .Y(n6980) );
  NBUFFX2_HVT U8363 ( .A(n6979), .Y(n6981) );
  NBUFFX2_HVT U8364 ( .A(n6979), .Y(n6982) );
  NBUFFX2_HVT U8365 ( .A(n6980), .Y(n6983) );
  NBUFFX2_HVT U8366 ( .A(n6980), .Y(n6984) );
  INVX0_HVT U8367 ( .A(n4375), .Y(n6985) );
  NBUFFX2_HVT U8368 ( .A(n6985), .Y(n6987) );
  NBUFFX2_HVT U8369 ( .A(n6985), .Y(n6988) );
  NBUFFX2_HVT U8370 ( .A(n4776), .Y(n6989) );
  NBUFFX2_HVT U8371 ( .A(n4776), .Y(n6990) );
  INVX0_HVT U8372 ( .A(n10128), .Y(n6991) );
  INVX0_HVT U8373 ( .A(n4374), .Y(n6992) );
  NBUFFX2_HVT U8374 ( .A(n6991), .Y(n6993) );
  NBUFFX2_HVT U8375 ( .A(n6991), .Y(n6994) );
  NBUFFX2_HVT U8376 ( .A(n6992), .Y(n6995) );
  NBUFFX2_HVT U8377 ( .A(n6992), .Y(n6996) );
  INVX0_HVT U8378 ( .A(n6997), .Y(n6999) );
  INVX0_HVT U8379 ( .A(n6997), .Y(n7000) );
  INVX0_HVT U8380 ( .A(n6997), .Y(n7001) );
  INVX0_HVT U8381 ( .A(n6998), .Y(n7002) );
  INVX0_HVT U8382 ( .A(n4601), .Y(n7003) );
  INVX0_HVT U8383 ( .A(n6998), .Y(n7004) );
  INVX0_HVT U8384 ( .A(n4601), .Y(n7005) );
  INVX1_HVT U8385 ( .A(n6968), .Y(n7016) );
  INVX0_HVT U8386 ( .A(n5072), .Y(n10129) );
  INVX0_HVT U8387 ( .A(n10348), .Y(n7026) );
  INVX0_HVT U8388 ( .A(n10348), .Y(n7027) );
  INVX0_HVT U8389 ( .A(n4263), .Y(n7028) );
  NBUFFX2_HVT U8390 ( .A(n7028), .Y(n7029) );
  NBUFFX2_HVT U8391 ( .A(n7028), .Y(n7030) );
  NBUFFX2_HVT U8392 ( .A(n7039), .Y(n7031) );
  NBUFFX2_HVT U8393 ( .A(n7028), .Y(n7032) );
  NBUFFX2_HVT U8394 ( .A(n7038), .Y(n7033) );
  NBUFFX2_HVT U8395 ( .A(n7044), .Y(n7034) );
  NBUFFX2_HVT U8396 ( .A(n4492), .Y(n7035) );
  NBUFFX2_HVT U8397 ( .A(n7043), .Y(n7036) );
  INVX0_HVT U8398 ( .A(n10350), .Y(n7037) );
  INVX0_HVT U8399 ( .A(n10349), .Y(n7038) );
  NBUFFX2_HVT U8400 ( .A(n7037), .Y(n7039) );
  NBUFFX2_HVT U8401 ( .A(n7037), .Y(n7040) );
  NBUFFX2_HVT U8402 ( .A(n7038), .Y(n7041) );
  NBUFFX2_HVT U8403 ( .A(n4266), .Y(n7042) );
  INVX0_HVT U8404 ( .A(n4263), .Y(n7043) );
  INVX0_HVT U8405 ( .A(n10350), .Y(n7044) );
  NBUFFX2_HVT U8406 ( .A(n7043), .Y(n7045) );
  NBUFFX2_HVT U8407 ( .A(n4264), .Y(n7046) );
  NBUFFX2_HVT U8408 ( .A(n4747), .Y(n7047) );
  NBUFFX2_HVT U8409 ( .A(n7049), .Y(n7048) );
  INVX0_HVT U8410 ( .A(n10350), .Y(n7049) );
  NBUFFX2_HVT U8411 ( .A(n4492), .Y(n7050) );
  NBUFFX2_HVT U8412 ( .A(n7049), .Y(n7051) );
  NBUFFX2_HVT U8413 ( .A(n4747), .Y(n7052) );
  IBUFFX2_HVT U8414 ( .A(n10351), .Y(n7054) );
  INVX0_HVT U8415 ( .A(n4493), .Y(n7055) );
  INVX0_HVT U8416 ( .A(n4493), .Y(n7056) );
  INVX0_HVT U8417 ( .A(n7053), .Y(n7057) );
  INVX0_HVT U8418 ( .A(n7053), .Y(n7058) );
  INVX0_HVT U8419 ( .A(n7054), .Y(n7059) );
  INVX0_HVT U8420 ( .A(n7054), .Y(n7060) );
  INVX0_HVT U8421 ( .A(n7054), .Y(n7061) );
  INVX0_HVT U8422 ( .A(n7054), .Y(n7062) );
  INVX1_HVT U8423 ( .A(n7026), .Y(n7063) );
  INVX1_HVT U8424 ( .A(n7027), .Y(n7073) );
  INVX0_HVT U8425 ( .A(n5013), .Y(n10351) );
  INVX0_HVT U8426 ( .A(n10), .Y(n10348) );
  IBUFFX2_HVT U8427 ( .A(n10351), .Y(n10349) );
  MUX41X1_HVT U8428 ( .A1(\ram[7][161] ), .A3(\ram[5][161] ), .A2(
        \ram[6][161] ), .A4(\ram[4][161] ), .S0(n6645), .S1(n5922), .Y(n8375)
         );
  INVX0_HVT U8429 ( .A(n10129), .Y(n10127) );
  INVX0_HVT U8430 ( .A(n10317), .Y(n7085) );
  INVX0_HVT U8431 ( .A(n10317), .Y(n7086) );
  NBUFFX2_HVT U8432 ( .A(n7101), .Y(n7087) );
  NBUFFX2_HVT U8433 ( .A(n7096), .Y(n7088) );
  NBUFFX2_HVT U8434 ( .A(n7091), .Y(n7089) );
  NBUFFX2_HVT U8435 ( .A(n7102), .Y(n7090) );
  NBUFFX2_HVT U8436 ( .A(n7091), .Y(n7092) );
  NBUFFX2_HVT U8437 ( .A(n7091), .Y(n7093) );
  NBUFFX2_HVT U8438 ( .A(n7091), .Y(n7094) );
  NBUFFX2_HVT U8439 ( .A(n7091), .Y(n7095) );
  INVX0_HVT U8440 ( .A(n10318), .Y(n7096) );
  NBUFFX2_HVT U8441 ( .A(n7096), .Y(n7097) );
  NBUFFX2_HVT U8442 ( .A(n7096), .Y(n7098) );
  NBUFFX2_HVT U8443 ( .A(n7096), .Y(n7099) );
  NBUFFX2_HVT U8444 ( .A(n7102), .Y(n7100) );
  INVX0_HVT U8445 ( .A(n10316), .Y(n7101) );
  INVX0_HVT U8446 ( .A(n10318), .Y(n7102) );
  NBUFFX2_HVT U8447 ( .A(n7101), .Y(n7103) );
  NBUFFX2_HVT U8448 ( .A(n7101), .Y(n7104) );
  NBUFFX2_HVT U8449 ( .A(n7102), .Y(n7105) );
  NBUFFX2_HVT U8450 ( .A(n7102), .Y(n7106) );
  INVX0_HVT U8451 ( .A(n10316), .Y(n7107) );
  NBUFFX2_HVT U8452 ( .A(n7107), .Y(n7108) );
  NBUFFX2_HVT U8453 ( .A(n7107), .Y(n7109) );
  NBUFFX2_HVT U8454 ( .A(n7107), .Y(n7110) );
  NBUFFX2_HVT U8455 ( .A(n7101), .Y(n7111) );
  INVX0_HVT U8456 ( .A(n10318), .Y(n7113) );
  INVX0_HVT U8457 ( .A(n10316), .Y(n7114) );
  INVX0_HVT U8458 ( .A(n7112), .Y(n7115) );
  INVX0_HVT U8459 ( .A(n7112), .Y(n7116) );
  INVX0_HVT U8460 ( .A(n7112), .Y(n7117) );
  INVX0_HVT U8461 ( .A(n7112), .Y(n7118) );
  INVX0_HVT U8462 ( .A(n7112), .Y(n7119) );
  INVX1_HVT U8463 ( .A(n7085), .Y(n7120) );
  INVX1_HVT U8464 ( .A(n7085), .Y(n7121) );
  INVX1_HVT U8465 ( .A(n7121), .Y(n7126) );
  INVX1_HVT U8466 ( .A(n7121), .Y(n7129) );
  INVX1_HVT U8467 ( .A(n7086), .Y(n7130) );
  INVX1_HVT U8468 ( .A(n7086), .Y(n7131) );
  INVX1_HVT U8469 ( .A(n7131), .Y(n7136) );
  INVX1_HVT U8470 ( .A(n7131), .Y(n7138) );
  INVX1_HVT U8471 ( .A(n7131), .Y(n7139) );
  INVX0_HVT U8472 ( .A(n4355), .Y(n10317) );
  MUX41X1_HVT U8473 ( .A1(\ram[15][105] ), .A3(\ram[13][105] ), .A2(
        \ram[14][105] ), .A4(\ram[12][105] ), .S0(n5759), .S1(n5883), .Y(n8150) );
  MUX41X1_HVT U8474 ( .A1(\ram[15][54] ), .A3(\ram[13][54] ), .A2(
        \ram[14][54] ), .A4(\ram[12][54] ), .S0(n5759), .S1(n7345), .Y(n7947)
         );
  MUX41X1_HVT U8475 ( .A1(n7752), .A3(n7750), .A2(n7753), .A4(n7751), .S0(
        n7562), .S1(n6257), .Y(q[4]) );
  AO22X1_HVT U8476 ( .A1(\ram[13][72] ), .A2(n4763), .A3(n4786), .A4(data[72]), 
        .Y(n3461) );
  IBUFFX2_HVT U8477 ( .A(n8783), .Y(n7145) );
  MUX41X1_HVT U8478 ( .A1(\ram[3][81] ), .A3(\ram[1][81] ), .A2(\ram[2][81] ), 
        .A4(\ram[0][81] ), .S0(n5894), .S1(n4175), .Y(n8057) );
  MUX41X1_HVT U8479 ( .A1(\ram[3][218] ), .A3(\ram[1][218] ), .A2(
        \ram[2][218] ), .A4(\ram[0][218] ), .S0(n5640), .S1(n5567), .Y(n8604)
         );
  MUX41X1_HVT U8480 ( .A1(\ram[3][165] ), .A3(\ram[1][165] ), .A2(
        \ram[2][165] ), .A4(\ram[0][165] ), .S0(n7303), .S1(n7294), .Y(n8392)
         );
  INVX0_HVT U8481 ( .A(n10332), .Y(n7152) );
  INVX0_HVT U8482 ( .A(n10332), .Y(n7153) );
  INVX0_HVT U8483 ( .A(n4716), .Y(n7154) );
  NBUFFX2_HVT U8484 ( .A(n4408), .Y(n7155) );
  NBUFFX2_HVT U8485 ( .A(n4408), .Y(n7156) );
  NBUFFX2_HVT U8486 ( .A(n7154), .Y(n7157) );
  NBUFFX2_HVT U8487 ( .A(n7154), .Y(n7158) );
  NBUFFX2_HVT U8488 ( .A(n7153), .Y(n7159) );
  NBUFFX2_HVT U8489 ( .A(n7152), .Y(n7160) );
  NBUFFX2_HVT U8490 ( .A(n7168), .Y(n7161) );
  NBUFFX2_HVT U8491 ( .A(n7169), .Y(n7162) );
  INVX0_HVT U8492 ( .A(n10334), .Y(n7163) );
  NBUFFX2_HVT U8493 ( .A(n7163), .Y(n7164) );
  NBUFFX2_HVT U8494 ( .A(n7163), .Y(n7165) );
  NBUFFX2_HVT U8495 ( .A(n7163), .Y(n7166) );
  NBUFFX2_HVT U8496 ( .A(n7163), .Y(n7167) );
  INVX0_HVT U8497 ( .A(n10333), .Y(n7168) );
  INVX0_HVT U8498 ( .A(n10333), .Y(n7169) );
  NBUFFX2_HVT U8499 ( .A(n7168), .Y(n7170) );
  NBUFFX2_HVT U8500 ( .A(n7168), .Y(n7171) );
  NBUFFX2_HVT U8501 ( .A(n7169), .Y(n7172) );
  NBUFFX2_HVT U8502 ( .A(n7169), .Y(n7173) );
  INVX0_HVT U8503 ( .A(n10334), .Y(n7174) );
  NBUFFX2_HVT U8504 ( .A(n7174), .Y(n7176) );
  NBUFFX2_HVT U8505 ( .A(n7174), .Y(n7177) );
  NBUFFX2_HVT U8506 ( .A(n7175), .Y(n7178) );
  NBUFFX2_HVT U8507 ( .A(n7175), .Y(n7179) );
  INVX0_HVT U8508 ( .A(n4716), .Y(n7180) );
  INVX0_HVT U8509 ( .A(n10331), .Y(n7181) );
  INVX0_HVT U8510 ( .A(n10331), .Y(n7182) );
  INVX0_HVT U8511 ( .A(n10331), .Y(n7183) );
  INVX0_HVT U8512 ( .A(n4716), .Y(n7184) );
  INVX0_HVT U8513 ( .A(n10331), .Y(n7185) );
  INVX0_HVT U8514 ( .A(n10331), .Y(n7186) );
  INVX1_HVT U8515 ( .A(n7152), .Y(n7187) );
  INVX1_HVT U8516 ( .A(n7198), .Y(n7203) );
  INVX1_HVT U8517 ( .A(n7198), .Y(n7204) );
  INVX1_HVT U8518 ( .A(n7198), .Y(n7206) );
  INVX0_HVT U8519 ( .A(n4957), .Y(n10332) );
  IBUFFX2_HVT U8520 ( .A(n4957), .Y(n10333) );
  AO22X1_HVT U8521 ( .A1(\ram[15][216] ), .A2(n5918), .A3(n8978), .A4(n9969), 
        .Y(n4117) );
  INVX0_HVT U8522 ( .A(n10117), .Y(n7207) );
  INVX0_HVT U8523 ( .A(n10117), .Y(n7208) );
  NBUFFX2_HVT U8524 ( .A(n4475), .Y(n7209) );
  NBUFFX2_HVT U8525 ( .A(n7231), .Y(n7210) );
  NBUFFX2_HVT U8526 ( .A(n4475), .Y(n7211) );
  NBUFFX2_HVT U8527 ( .A(n7213), .Y(n7212) );
  NBUFFX2_HVT U8528 ( .A(n4475), .Y(n7214) );
  NBUFFX2_HVT U8529 ( .A(n4475), .Y(n7215) );
  NBUFFX2_HVT U8530 ( .A(n7213), .Y(n7216) );
  NBUFFX2_HVT U8531 ( .A(n7213), .Y(n7217) );
  INVX0_HVT U8532 ( .A(n4298), .Y(n7218) );
  INVX0_HVT U8533 ( .A(n4298), .Y(n7219) );
  NBUFFX2_HVT U8534 ( .A(n7218), .Y(n7220) );
  NBUFFX2_HVT U8535 ( .A(n7218), .Y(n7221) );
  NBUFFX2_HVT U8536 ( .A(n7219), .Y(n7222) );
  NBUFFX2_HVT U8537 ( .A(n7219), .Y(n7223) );
  INVX0_HVT U8538 ( .A(n10119), .Y(n7224) );
  INVX0_HVT U8539 ( .A(n10118), .Y(n7225) );
  NBUFFX2_HVT U8540 ( .A(n7224), .Y(n7226) );
  NBUFFX2_HVT U8541 ( .A(n7224), .Y(n7227) );
  NBUFFX2_HVT U8542 ( .A(n7225), .Y(n7228) );
  NBUFFX2_HVT U8543 ( .A(n7225), .Y(n7229) );
  INVX0_HVT U8544 ( .A(n4378), .Y(n7230) );
  INVX0_HVT U8545 ( .A(n4378), .Y(n7231) );
  NBUFFX2_HVT U8546 ( .A(n7230), .Y(n7232) );
  NBUFFX2_HVT U8547 ( .A(n7230), .Y(n7233) );
  NBUFFX2_HVT U8548 ( .A(n7231), .Y(n7234) );
  NBUFFX2_HVT U8549 ( .A(n7213), .Y(n7235) );
  INVX0_HVT U8550 ( .A(n7236), .Y(n7237) );
  INVX0_HVT U8551 ( .A(n10118), .Y(n7238) );
  INVX0_HVT U8552 ( .A(n7236), .Y(n7239) );
  INVX0_HVT U8553 ( .A(n10118), .Y(n7240) );
  INVX0_HVT U8554 ( .A(n4298), .Y(n7241) );
  INVX0_HVT U8555 ( .A(n7236), .Y(n7242) );
  INVX0_HVT U8556 ( .A(n4378), .Y(n7243) );
  INVX1_HVT U8557 ( .A(n7207), .Y(n7244) );
  INVX1_HVT U8558 ( .A(n7208), .Y(n7253) );
  INVX1_HVT U8559 ( .A(n7208), .Y(n7254) );
  INVX1_HVT U8560 ( .A(n7254), .Y(n7259) );
  INVX1_HVT U8561 ( .A(n7254), .Y(n7260) );
  INVX1_HVT U8562 ( .A(n7254), .Y(n7261) );
  INVX1_HVT U8563 ( .A(n7254), .Y(n7262) );
  INVX0_HVT U8564 ( .A(n10121), .Y(n10120) );
  INVX0_HVT U8565 ( .A(n10120), .Y(n10117) );
  AO22X1_HVT U8566 ( .A1(\ram[14][144] ), .A2(n7258), .A3(n9058), .A4(n9742), 
        .Y(n3789) );
  INVX0_HVT U8567 ( .A(n7326), .Y(n7296) );
  INVX0_HVT U8568 ( .A(n10164), .Y(n10161) );
  INVX0_HVT U8569 ( .A(n10164), .Y(n10162) );
  MUX41X1_HVT U8570 ( .A1(n8581), .A3(n8583), .A2(n8582), .A4(n8584), .S0(
        n7548), .S1(n5774), .Y(q[213]) );
  MUX41X1_HVT U8571 ( .A1(\ram[15][37] ), .A3(\ram[13][37] ), .A2(
        \ram[14][37] ), .A4(\ram[12][37] ), .S0(n7314), .S1(n7266), .Y(n7879)
         );
  MUX41X1_HVT U8572 ( .A1(\ram[3][66] ), .A3(\ram[1][66] ), .A2(\ram[2][66] ), 
        .A4(\ram[0][66] ), .S0(n5982), .S1(n6655), .Y(n7997) );
  MUX41X1_HVT U8573 ( .A1(n7994), .A3(n7996), .A2(n7995), .A4(n7997), .S0(
        n5207), .S1(n5503), .Y(q[66]) );
  NAND2X0_HVT U8574 ( .A1(\ram[6][48] ), .A2(n6630), .Y(n7273) );
  NAND2X0_HVT U8575 ( .A1(n9200), .A2(n9451), .Y(n7274) );
  NAND2X0_HVT U8576 ( .A1(n7273), .A2(n7274), .Y(n1645) );
  MUX41X1_HVT U8577 ( .A1(\ram[3][72] ), .A3(\ram[1][72] ), .A2(\ram[2][72] ), 
        .A4(\ram[0][72] ), .S0(n6412), .S1(n5933), .Y(n8021) );
  MUX41X1_HVT U8578 ( .A1(\ram[11][70] ), .A3(\ram[9][70] ), .A2(\ram[10][70] ), .A4(\ram[8][70] ), .S0(n7281), .S1(n7282), .Y(n8011) );
  MUX41X1_HVT U8579 ( .A1(\ram[11][69] ), .A3(\ram[9][69] ), .A2(\ram[10][69] ), .A4(\ram[8][69] ), .S0(n7682), .S1(n7283), .Y(n8007) );
  MUX41X1_HVT U8580 ( .A1(\ram[15][81] ), .A3(\ram[13][81] ), .A2(
        \ram[14][81] ), .A4(\ram[12][81] ), .S0(n5743), .S1(n6135), .Y(n8054)
         );
  MUX41X1_HVT U8581 ( .A1(\ram[11][145] ), .A3(\ram[9][145] ), .A2(
        \ram[10][145] ), .A4(\ram[8][145] ), .S0(n7296), .S1(n5958), .Y(n8310)
         );
  MUX41X1_HVT U8582 ( .A1(n8313), .A3(n8315), .A2(n8314), .A4(n8316), .S0(
        n7685), .S1(n7288), .Y(q[146]) );
  MUX41X1_HVT U8583 ( .A1(\ram[15][72] ), .A3(\ram[13][72] ), .A2(
        \ram[14][72] ), .A4(\ram[12][72] ), .S0(n7557), .S1(n5933), .Y(n8018)
         );
  MUX41X1_HVT U8584 ( .A1(\ram[15][48] ), .A3(\ram[13][48] ), .A2(
        \ram[14][48] ), .A4(\ram[12][48] ), .S0(n5976), .S1(n7290), .Y(n7923)
         );
  MUX41X1_HVT U8585 ( .A1(\ram[15][213] ), .A3(\ram[13][213] ), .A2(
        \ram[14][213] ), .A4(\ram[12][213] ), .S0(n7296), .S1(n5568), .Y(n8581) );
  INVX0_HVT U8586 ( .A(n8839), .Y(n7306) );
  MUX41X1_HVT U8587 ( .A1(\ram[14][145] ), .A3(\ram[12][145] ), .A2(
        \ram[15][145] ), .A4(\ram[13][145] ), .S0(n7296), .S1(n7329), .Y(n8309) );
  MUX41X1_HVT U8588 ( .A1(n8367), .A3(n8365), .A2(n8368), .A4(n8366), .S0(
        n7300), .S1(n7301), .Y(q[159]) );
  MUX41X1_HVT U8589 ( .A1(\ram[13][134] ), .A3(\ram[15][134] ), .A2(
        \ram[12][134] ), .A4(\ram[14][134] ), .S0(n8803), .S1(n5958), .Y(n8266) );
  MUX41X1_HVT U8590 ( .A1(\ram[11][186] ), .A3(\ram[9][186] ), .A2(
        \ram[10][186] ), .A4(\ram[8][186] ), .S0(n5976), .S1(n6745), .Y(n8474)
         );
  MUX41X1_HVT U8591 ( .A1(\ram[11][170] ), .A3(\ram[9][170] ), .A2(
        \ram[10][170] ), .A4(\ram[8][170] ), .S0(n7303), .S1(n6657), .Y(n8410)
         );
  MUX41X1_HVT U8592 ( .A1(\ram[11][167] ), .A3(\ram[9][167] ), .A2(
        \ram[10][167] ), .A4(\ram[8][167] ), .S0(n7304), .S1(n7699), .Y(n8398)
         );
  MUX41X1_HVT U8593 ( .A1(\ram[3][159] ), .A3(\ram[1][159] ), .A2(
        \ram[2][159] ), .A4(\ram[0][159] ), .S0(n5507), .S1(n4987), .Y(n8368)
         );
  MUX41X1_HVT U8594 ( .A1(\ram[15][57] ), .A3(\ram[13][57] ), .A2(
        \ram[14][57] ), .A4(\ram[12][57] ), .S0(n4993), .S1(n5922), .Y(n7959)
         );
  MUX41X1_HVT U8595 ( .A1(\ram[15][36] ), .A3(\ram[13][36] ), .A2(
        \ram[14][36] ), .A4(\ram[12][36] ), .S0(n4989), .S1(n7317), .Y(n7875)
         );
  NBUFFX2_HVT U8596 ( .A(n8784), .Y(n7316) );
  NBUFFX2_HVT U8597 ( .A(n5164), .Y(n8856) );
  IBUFFX2_HVT U8598 ( .A(n5091), .Y(n8848) );
  NBUFFX2_HVT U8599 ( .A(n6758), .Y(n7322) );
  MUX41X1_HVT U8600 ( .A1(\ram[11][233] ), .A3(\ram[9][233] ), .A2(
        \ram[10][233] ), .A4(\ram[8][233] ), .S0(n7284), .S1(n5732), .Y(n8661)
         );
  MUX41X1_HVT U8601 ( .A1(\ram[15][239] ), .A3(\ram[13][239] ), .A2(
        \ram[14][239] ), .A4(\ram[12][239] ), .S0(n5594), .S1(n7331), .Y(n8683) );
  MUX41X1_HVT U8602 ( .A1(n8318), .A3(n8320), .A2(n8317), .A4(n8319), .S0(
        n5111), .S1(n7332), .Y(q[147]) );
  MUX41X1_HVT U8603 ( .A1(\ram[15][182] ), .A3(\ram[13][182] ), .A2(
        \ram[14][182] ), .A4(\ram[12][182] ), .S0(n5142), .S1(n5342), .Y(n8457) );
  IBUFFX2_HVT U8604 ( .A(n5155), .Y(n7337) );
  MUX41X1_HVT U8605 ( .A1(\ram[15][130] ), .A3(\ram[13][130] ), .A2(
        \ram[14][130] ), .A4(\ram[12][130] ), .S0(n5975), .S1(n7340), .Y(n8250) );
  MUX41X1_HVT U8606 ( .A1(\ram[15][237] ), .A3(\ram[13][237] ), .A2(
        \ram[14][237] ), .A4(\ram[12][237] ), .S0(n6405), .S1(n5304), .Y(n8675) );
  MUX41X1_HVT U8607 ( .A1(\ram[3][129] ), .A3(\ram[1][129] ), .A2(
        \ram[2][129] ), .A4(\ram[0][129] ), .S0(n5640), .S1(n5732), .Y(n8249)
         );
  NBUFFX2_HVT U8608 ( .A(n6132), .Y(n8879) );
  MUX41X1_HVT U8609 ( .A1(\ram[3][209] ), .A3(\ram[1][209] ), .A2(
        \ram[2][209] ), .A4(\ram[0][209] ), .S0(n6414), .S1(n7143), .Y(n8568)
         );
  MUX41X1_HVT U8610 ( .A1(\ram[3][78] ), .A3(\ram[1][78] ), .A2(\ram[2][78] ), 
        .A4(\ram[0][78] ), .S0(n6414), .S1(n7266), .Y(n8045) );
  MUX41X1_HVT U8611 ( .A1(n8042), .A3(n8044), .A2(n8043), .A4(n8045), .S0(
        n7548), .S1(n6398), .Y(q[78]) );
  MUX41X1_HVT U8612 ( .A1(\ram[15][123] ), .A3(\ram[13][123] ), .A2(
        \ram[14][123] ), .A4(\ram[12][123] ), .S0(n4989), .S1(n6734), .Y(n8222) );
  MUX41X1_HVT U8613 ( .A1(\ram[15][27] ), .A3(\ram[13][27] ), .A2(
        \ram[14][27] ), .A4(\ram[12][27] ), .S0(n5998), .S1(n6657), .Y(n7840)
         );
  INVX0_HVT U8614 ( .A(n10162), .Y(n10152) );
  INVX0_HVT U8615 ( .A(n10188), .Y(n10186) );
  INVX0_HVT U8616 ( .A(n10188), .Y(n10187) );
  IBUFFX2_HVT U8617 ( .A(n10189), .Y(n10183) );
  IBUFFX2_HVT U8618 ( .A(n10189), .Y(n10184) );
  IBUFFX2_HVT U8619 ( .A(n10189), .Y(n10185) );
  INVX0_HVT U8620 ( .A(n6103), .Y(n10232) );
  INVX0_HVT U8621 ( .A(n6043), .Y(n10233) );
  INVX0_HVT U8622 ( .A(n6044), .Y(n10234) );
  INVX0_HVT U8623 ( .A(n10161), .Y(n10158) );
  INVX0_HVT U8624 ( .A(n10161), .Y(n10159) );
  INVX0_HVT U8625 ( .A(n6077), .Y(n10225) );
  INVX0_HVT U8626 ( .A(n6081), .Y(n10226) );
  INVX0_HVT U8627 ( .A(n6043), .Y(n10227) );
  MUX41X1_HVT U8628 ( .A1(n8246), .A3(n8248), .A2(n8247), .A4(n8249), .S0(
        n5207), .S1(n5885), .Y(q[129]) );
  INVX1_HVT U8629 ( .A(n4545), .Y(n7354) );
  INVX0_HVT U8630 ( .A(n10239), .Y(n7362) );
  INVX0_HVT U8631 ( .A(n10239), .Y(n7363) );
  INVX1_HVT U8632 ( .A(n7362), .Y(n7364) );
  INVX1_HVT U8633 ( .A(n7363), .Y(n7365) );
  INVX1_HVT U8634 ( .A(n7403), .Y(n7366) );
  INVX1_HVT U8635 ( .A(n7404), .Y(n7367) );
  INVX0_HVT U8636 ( .A(n10240), .Y(n7368) );
  INVX1_HVT U8637 ( .A(n7368), .Y(n7369) );
  INVX1_HVT U8638 ( .A(n7389), .Y(n7371) );
  INVX1_HVT U8639 ( .A(n7368), .Y(n7374) );
  INVX0_HVT U8640 ( .A(n10241), .Y(n7376) );
  INVX1_HVT U8641 ( .A(n7382), .Y(n7377) );
  INVX1_HVT U8642 ( .A(n4545), .Y(n7380) );
  INVX0_HVT U8643 ( .A(n10249), .Y(n7381) );
  INVX0_HVT U8644 ( .A(n10249), .Y(n7382) );
  INVX0_HVT U8645 ( .A(n10243), .Y(n7385) );
  INVX0_HVT U8646 ( .A(n10243), .Y(n7386) );
  INVX1_HVT U8647 ( .A(n7385), .Y(n7387) );
  INVX1_HVT U8648 ( .A(n7386), .Y(n7388) );
  INVX0_HVT U8649 ( .A(n10244), .Y(n7389) );
  INVX1_HVT U8650 ( .A(n7389), .Y(n7391) );
  INVX0_HVT U8651 ( .A(n10245), .Y(n7392) );
  INVX0_HVT U8652 ( .A(n10245), .Y(n7393) );
  INVX1_HVT U8653 ( .A(n7385), .Y(n7398) );
  INVX1_HVT U8654 ( .A(n7362), .Y(n7399) );
  INVX1_HVT U8655 ( .A(n7363), .Y(n7400) );
  INVX1_HVT U8656 ( .A(n7381), .Y(n7401) );
  INVX1_HVT U8657 ( .A(n7386), .Y(n7402) );
  INVX0_HVT U8658 ( .A(n10246), .Y(n7403) );
  INVX0_HVT U8659 ( .A(n10246), .Y(n7404) );
  INVX1_HVT U8660 ( .A(n7403), .Y(n7405) );
  INVX1_HVT U8661 ( .A(n7404), .Y(n7406) );
  INVX0_HVT U8662 ( .A(n10241), .Y(n7407) );
  INVX1_HVT U8663 ( .A(n7407), .Y(n7408) );
  INVX0_HVT U8664 ( .A(n10247), .Y(n7410) );
  NBUFFX2_HVT U8665 ( .A(n10245), .Y(n7414) );
  NBUFFX2_HVT U8666 ( .A(n4434), .Y(n7415) );
  NBUFFX2_HVT U8667 ( .A(n10247), .Y(n7416) );
  NBUFFX2_HVT U8668 ( .A(n10240), .Y(n7417) );
  INVX0_HVT U8669 ( .A(n7353), .Y(n10237) );
  INVX0_HVT U8670 ( .A(n7726), .Y(n10238) );
  INVX0_HVT U8671 ( .A(n10250), .Y(n10239) );
  INVX0_HVT U8672 ( .A(n7407), .Y(n10249) );
  INVX0_HVT U8673 ( .A(n10251), .Y(n10243) );
  INVX0_HVT U8674 ( .A(n7358), .Y(n10244) );
  INVX0_HVT U8675 ( .A(n7353), .Y(n10245) );
  INVX0_HVT U8676 ( .A(n10251), .Y(n10246) );
  INVX0_HVT U8677 ( .A(n10250), .Y(n10247) );
  INVX0_HVT U8678 ( .A(n7376), .Y(n10248) );
  INVX0_HVT U8679 ( .A(n10165), .Y(n7418) );
  INVX1_HVT U8680 ( .A(n7418), .Y(n7419) );
  INVX0_HVT U8681 ( .A(n10165), .Y(n7421) );
  INVX0_HVT U8682 ( .A(n10173), .Y(n7424) );
  INVX1_HVT U8683 ( .A(n7424), .Y(n7425) );
  INVX1_HVT U8684 ( .A(n7424), .Y(n7426) );
  INVX1_HVT U8685 ( .A(n7424), .Y(n7427) );
  INVX0_HVT U8686 ( .A(n10172), .Y(n7428) );
  INVX0_HVT U8687 ( .A(n10167), .Y(n7432) );
  INVX1_HVT U8688 ( .A(n7432), .Y(n7433) );
  INVX1_HVT U8689 ( .A(n7432), .Y(n7434) );
  INVX1_HVT U8690 ( .A(n7456), .Y(n7436) );
  INVX0_HVT U8691 ( .A(n10167), .Y(n7437) );
  INVX1_HVT U8692 ( .A(n7437), .Y(n7440) );
  INVX1_HVT U8693 ( .A(n7437), .Y(n7441) );
  INVX1_HVT U8694 ( .A(n7459), .Y(n7442) );
  INVX1_HVT U8695 ( .A(n7459), .Y(n7443) );
  INVX1_HVT U8696 ( .A(n7456), .Y(n7444) );
  INVX0_HVT U8697 ( .A(n10170), .Y(n7446) );
  INVX0_HVT U8698 ( .A(n10170), .Y(n7449) );
  INVX0_HVT U8699 ( .A(n10171), .Y(n7453) );
  INVX0_HVT U8700 ( .A(n10172), .Y(n7456) );
  INVX1_HVT U8701 ( .A(n7456), .Y(n7457) );
  INVX1_HVT U8702 ( .A(n7456), .Y(n7458) );
  INVX0_HVT U8703 ( .A(n10173), .Y(n7459) );
  INVX1_HVT U8704 ( .A(n7462), .Y(n7460) );
  INVX1_HVT U8705 ( .A(n7459), .Y(n7461) );
  INVX0_HVT U8706 ( .A(n10174), .Y(n7462) );
  INVX1_HVT U8707 ( .A(n7462), .Y(n7463) );
  INVX1_HVT U8708 ( .A(n7462), .Y(n7464) );
  IBUFFX2_HVT U8709 ( .A(n7727), .Y(n7469) );
  NBUFFX2_HVT U8710 ( .A(n7469), .Y(n7470) );
  NBUFFX2_HVT U8711 ( .A(n7469), .Y(n7471) );
  NBUFFX2_HVT U8712 ( .A(n7469), .Y(n7472) );
  NBUFFX2_HVT U8713 ( .A(n7469), .Y(n7473) );
  NBUFFX2_HVT U8714 ( .A(n7469), .Y(n7474) );
  INVX0_HVT U8715 ( .A(n10176), .Y(n10165) );
  INVX0_HVT U8716 ( .A(n10177), .Y(n10166) );
  INVX0_HVT U8717 ( .A(n10177), .Y(n10167) );
  INVX0_HVT U8718 ( .A(n10177), .Y(n10168) );
  INVX0_HVT U8719 ( .A(n10177), .Y(n10169) );
  INVX0_HVT U8720 ( .A(n10176), .Y(n10170) );
  INVX0_HVT U8721 ( .A(n10176), .Y(n10171) );
  INVX0_HVT U8722 ( .A(n10175), .Y(n10172) );
  INVX0_HVT U8723 ( .A(n10175), .Y(n10173) );
  INVX0_HVT U8724 ( .A(n10175), .Y(n10174) );
  INVX1_HVT U8725 ( .A(n7528), .Y(n7475) );
  INVX1_HVT U8726 ( .A(n7513), .Y(n7476) );
  INVX0_HVT U8727 ( .A(n10197), .Y(n7477) );
  INVX1_HVT U8728 ( .A(n7477), .Y(n7478) );
  INVX1_HVT U8729 ( .A(n7477), .Y(n7479) );
  INVX1_HVT U8730 ( .A(n7513), .Y(n7480) );
  INVX1_HVT U8731 ( .A(n7487), .Y(n7481) );
  INVX0_HVT U8732 ( .A(n10192), .Y(n7482) );
  INVX1_HVT U8733 ( .A(n7507), .Y(n7483) );
  INVX1_HVT U8734 ( .A(n7482), .Y(n7484) );
  INVX1_HVT U8735 ( .A(n7488), .Y(n7485) );
  INVX1_HVT U8736 ( .A(n7533), .Y(n7486) );
  INVX0_HVT U8737 ( .A(n10194), .Y(n7487) );
  INVX0_HVT U8738 ( .A(n10191), .Y(n7488) );
  INVX1_HVT U8739 ( .A(n7487), .Y(n7489) );
  INVX1_HVT U8740 ( .A(n7488), .Y(n7490) );
  INVX1_HVT U8741 ( .A(n7504), .Y(n7491) );
  INVX1_HVT U8742 ( .A(n7488), .Y(n7492) );
  INVX1_HVT U8743 ( .A(n7516), .Y(n7493) );
  INVX1_HVT U8744 ( .A(n7517), .Y(n7494) );
  INVX0_HVT U8745 ( .A(n10196), .Y(n7495) );
  INVX0_HVT U8746 ( .A(n10196), .Y(n7496) );
  INVX1_HVT U8747 ( .A(n7495), .Y(n7497) );
  INVX1_HVT U8748 ( .A(n7496), .Y(n7498) );
  INVX1_HVT U8749 ( .A(n7510), .Y(n7499) );
  INVX1_HVT U8750 ( .A(n7496), .Y(n7500) );
  INVX0_HVT U8751 ( .A(n10199), .Y(n7501) );
  INVX1_HVT U8752 ( .A(n7501), .Y(n7502) );
  INVX1_HVT U8753 ( .A(n7501), .Y(n7503) );
  INVX0_HVT U8754 ( .A(n10195), .Y(n7504) );
  INVX1_HVT U8755 ( .A(n7504), .Y(n7505) );
  INVX1_HVT U8756 ( .A(n7504), .Y(n7506) );
  INVX0_HVT U8757 ( .A(n10192), .Y(n7507) );
  INVX1_HVT U8758 ( .A(n7507), .Y(n7508) );
  INVX1_HVT U8759 ( .A(n7482), .Y(n7509) );
  INVX1_HVT U8760 ( .A(n7529), .Y(n7511) );
  INVX0_HVT U8761 ( .A(n10194), .Y(n7513) );
  INVX1_HVT U8762 ( .A(n7513), .Y(n7514) );
  INVX1_HVT U8763 ( .A(n7487), .Y(n7515) );
  INVX1_HVT U8764 ( .A(n7516), .Y(n7518) );
  INVX1_HVT U8765 ( .A(n7517), .Y(n7519) );
  INVX0_HVT U8766 ( .A(n10198), .Y(n7520) );
  INVX1_HVT U8767 ( .A(n7525), .Y(n7521) );
  INVX1_HVT U8768 ( .A(n7520), .Y(n7522) );
  INVX1_HVT U8769 ( .A(n7517), .Y(n7523) );
  INVX1_HVT U8770 ( .A(n7516), .Y(n7524) );
  INVX0_HVT U8771 ( .A(n10198), .Y(n7525) );
  INVX1_HVT U8772 ( .A(n7520), .Y(n7526) );
  INVX1_HVT U8773 ( .A(n7525), .Y(n7527) );
  INVX0_HVT U8774 ( .A(n10197), .Y(n7528) );
  INVX0_HVT U8775 ( .A(n10197), .Y(n7529) );
  INVX1_HVT U8776 ( .A(n7528), .Y(n7530) );
  INVX1_HVT U8777 ( .A(n7529), .Y(n7531) );
  INVX0_HVT U8778 ( .A(n10193), .Y(n7533) );
  INVX1_HVT U8779 ( .A(n7532), .Y(n7534) );
  INVX1_HVT U8780 ( .A(n7520), .Y(n7536) );
  INVX1_HVT U8781 ( .A(n7525), .Y(n7537) );
  INVX1_HVT U8782 ( .A(n7495), .Y(n7538) );
  NBUFFX2_HVT U8783 ( .A(n10191), .Y(n7539) );
  NBUFFX2_HVT U8784 ( .A(n10198), .Y(n7540) );
  NBUFFX2_HVT U8785 ( .A(n10199), .Y(n7541) );
  NBUFFX2_HVT U8786 ( .A(n10196), .Y(n7542) );
  INVX0_HVT U8787 ( .A(n10201), .Y(n10191) );
  INVX0_HVT U8788 ( .A(n10200), .Y(n10194) );
  INVX0_HVT U8789 ( .A(n10200), .Y(n10195) );
  INVX0_HVT U8790 ( .A(n7532), .Y(n10196) );
  INVX0_HVT U8791 ( .A(n7532), .Y(n10192) );
  INVX0_HVT U8792 ( .A(n7728), .Y(n10193) );
  INVX0_HVT U8793 ( .A(n7533), .Y(n10197) );
  INVX0_HVT U8794 ( .A(n10201), .Y(n10198) );
  INVX0_HVT U8795 ( .A(n7510), .Y(n10199) );
  INVX0_HVT U8796 ( .A(n6626), .Y(n7552) );
  MUX41X1_HVT U8797 ( .A1(\ram[11][197] ), .A3(\ram[9][197] ), .A2(
        \ram[10][197] ), .A4(\ram[8][197] ), .S0(n7147), .S1(n5919), .Y(n8518)
         );
  MUX41X1_HVT U8798 ( .A1(\ram[7][178] ), .A3(\ram[5][178] ), .A2(
        \ram[6][178] ), .A4(\ram[4][178] ), .S0(n7556), .S1(n5588), .Y(n8443)
         );
  MUX41X1_HVT U8799 ( .A1(\ram[15][240] ), .A3(\ram[13][240] ), .A2(
        \ram[14][240] ), .A4(\ram[12][240] ), .S0(n7571), .S1(n6753), .Y(n8687) );
  MUX41X1_HVT U8800 ( .A1(\ram[7][195] ), .A3(\ram[5][195] ), .A2(
        \ram[6][195] ), .A4(\ram[4][195] ), .S0(n5059), .S1(n5342), .Y(n8511)
         );
  AO22X1_HVT U8801 ( .A1(\ram[2][48] ), .A2(n7175), .A3(n6268), .A4(n9451), 
        .Y(n621) );
  MUX41X1_HVT U8802 ( .A1(\ram[12][156] ), .A3(\ram[14][156] ), .A2(
        \ram[13][156] ), .A4(\ram[15][156] ), .S0(n6653), .S1(n6382), .Y(n8353) );
  INVX0_HVT U8803 ( .A(n7573), .Y(n7566) );
  MUX41X1_HVT U8804 ( .A1(\ram[8][193] ), .A3(\ram[10][193] ), .A2(
        \ram[9][193] ), .A4(\ram[11][193] ), .S0(n5854), .S1(n6382), .Y(n8502)
         );
  MUX41X1_HVT U8805 ( .A1(n8374), .A3(n8376), .A2(n8373), .A4(n8375), .S0(
        n5655), .S1(n8767), .Y(q[161]) );
  AO22X1_HVT U8806 ( .A1(\ram[1][48] ), .A2(n4612), .A3(n6883), .A4(n9451), 
        .Y(n365) );
  MUX41X1_HVT U8807 ( .A1(\ram[7][133] ), .A3(\ram[5][133] ), .A2(
        \ram[6][133] ), .A4(\ram[4][133] ), .S0(n7571), .S1(n7266), .Y(n8264)
         );
  NBUFFX2_HVT U8808 ( .A(n6739), .Y(n7703) );
  MUX41X1_HVT U8809 ( .A1(\ram[15][160] ), .A3(\ram[13][160] ), .A2(
        \ram[14][160] ), .A4(\ram[12][160] ), .S0(n6414), .S1(n5919), .Y(n8369) );
  MUX41X1_HVT U8810 ( .A1(\ram[15][230] ), .A3(\ram[13][230] ), .A2(
        \ram[14][230] ), .A4(\ram[12][230] ), .S0(n7572), .S1(n5342), .Y(n8649) );
  MUX41X1_HVT U8811 ( .A1(n8601), .A3(n8603), .A2(n8602), .A4(n8604), .S0(
        n5343), .S1(n7677), .Y(q[218]) );
  IBUFFX2_HVT U8812 ( .A(n6750), .Y(n8758) );
  MUX41X1_HVT U8813 ( .A1(\ram[13][255] ), .A3(\ram[15][255] ), .A2(
        \ram[12][255] ), .A4(\ram[14][255] ), .S0(n7298), .S1(n6113), .Y(n8747) );
  MUX41X1_HVT U8814 ( .A1(\ram[15][108] ), .A3(\ram[13][108] ), .A2(
        \ram[14][108] ), .A4(\ram[12][108] ), .S0(n5357), .S1(n5818), .Y(n8162) );
  MUX41X1_HVT U8815 ( .A1(\ram[3][177] ), .A3(\ram[1][177] ), .A2(
        \ram[2][177] ), .A4(\ram[0][177] ), .S0(n7265), .S1(n4167), .Y(n8440)
         );
  MUX41X1_HVT U8816 ( .A1(\ram[15][222] ), .A3(\ram[13][222] ), .A2(
        \ram[14][222] ), .A4(\ram[12][222] ), .S0(n5968), .S1(n5919), .Y(n8617) );
  MUX41X1_HVT U8817 ( .A1(\ram[15][138] ), .A3(\ram[13][138] ), .A2(
        \ram[14][138] ), .A4(\ram[12][138] ), .S0(n6405), .S1(n5607), .Y(n8282) );
  INVX0_HVT U8818 ( .A(n10207), .Y(n7589) );
  INVX1_HVT U8819 ( .A(n7589), .Y(n7592) );
  INVX0_HVT U8820 ( .A(n10208), .Y(n7593) );
  INVX0_HVT U8821 ( .A(n10208), .Y(n7594) );
  INVX1_HVT U8822 ( .A(n7593), .Y(n7595) );
  INVX1_HVT U8823 ( .A(n7594), .Y(n7596) );
  INVX1_HVT U8824 ( .A(n7594), .Y(n7597) );
  INVX0_HVT U8825 ( .A(n10209), .Y(n7598) );
  INVX1_HVT U8826 ( .A(n7598), .Y(n7599) );
  INVX1_HVT U8827 ( .A(n7594), .Y(n7600) );
  INVX1_HVT U8828 ( .A(n7593), .Y(n7601) );
  INVX0_HVT U8829 ( .A(n10210), .Y(n7602) );
  INVX0_HVT U8830 ( .A(n10210), .Y(n7603) );
  INVX0_HVT U8831 ( .A(n10208), .Y(n7607) );
  INVX0_HVT U8832 ( .A(n10213), .Y(n7608) );
  INVX1_HVT U8833 ( .A(n7607), .Y(n7610) );
  INVX0_HVT U8834 ( .A(n10211), .Y(n7612) );
  INVX1_HVT U8835 ( .A(n7612), .Y(n7613) );
  INVX0_HVT U8836 ( .A(n10213), .Y(n7616) );
  INVX0_HVT U8837 ( .A(n10214), .Y(n7620) );
  INVX0_HVT U8838 ( .A(n10214), .Y(n7621) );
  INVX1_HVT U8839 ( .A(n7620), .Y(n7622) );
  INVX1_HVT U8840 ( .A(n7621), .Y(n7623) );
  INVX1_HVT U8841 ( .A(n7620), .Y(n7624) );
  INVX1_HVT U8842 ( .A(n7621), .Y(n7625) );
  INVX1_HVT U8843 ( .A(n7621), .Y(n7626) );
  INVX0_HVT U8844 ( .A(n10215), .Y(n7628) );
  INVX0_HVT U8845 ( .A(n10215), .Y(n7629) );
  INVX1_HVT U8846 ( .A(n7629), .Y(n7630) );
  INVX1_HVT U8847 ( .A(n7628), .Y(n7631) );
  INVX1_HVT U8848 ( .A(n7629), .Y(n7632) );
  INVX0_HVT U8849 ( .A(n10210), .Y(n7633) );
  INVX1_HVT U8850 ( .A(n7628), .Y(n7638) );
  INVX1_HVT U8851 ( .A(n7629), .Y(n7641) );
  INVX0_HVT U8852 ( .A(n10216), .Y(n7644) );
  INVX0_HVT U8853 ( .A(n10207), .Y(n7647) );
  INVX1_HVT U8854 ( .A(n7647), .Y(n7650) );
  INVX0_HVT U8855 ( .A(n10211), .Y(n7651) );
  INVX0_HVT U8856 ( .A(n10217), .Y(n7655) );
  INVX0_HVT U8857 ( .A(n10213), .Y(n7659) );
  INVX0_HVT U8858 ( .A(n4613), .Y(n10207) );
  INVX0_HVT U8859 ( .A(n10219), .Y(n10208) );
  INVX0_HVT U8860 ( .A(n10220), .Y(n10209) );
  INVX0_HVT U8861 ( .A(n7586), .Y(n10214) );
  INVX0_HVT U8862 ( .A(n10218), .Y(n10215) );
  INVX0_HVT U8863 ( .A(n10218), .Y(n10216) );
  IBUFFX2_HVT U8864 ( .A(n5581), .Y(n7677) );
  MUX41X1_HVT U8865 ( .A1(\ram[15][71] ), .A3(\ram[13][71] ), .A2(
        \ram[14][71] ), .A4(\ram[12][71] ), .S0(n7147), .S1(n7149), .Y(n8014)
         );
  MUX41X1_HVT U8866 ( .A1(\ram[15][167] ), .A3(\ram[13][167] ), .A2(
        \ram[14][167] ), .A4(\ram[12][167] ), .S0(n7306), .S1(n7688), .Y(n8397) );
  MUX41X1_HVT U8867 ( .A1(\ram[3][137] ), .A3(\ram[1][137] ), .A2(
        \ram[2][137] ), .A4(\ram[0][137] ), .S0(n4989), .S1(n7290), .Y(n8281)
         );
  MUX41X1_HVT U8868 ( .A1(\ram[11][128] ), .A3(\ram[9][128] ), .A2(
        \ram[10][128] ), .A4(\ram[8][128] ), .S0(n5357), .S1(n4175), .Y(n8243)
         );
  MUX41X1_HVT U8869 ( .A1(n7891), .A3(n7893), .A2(n7892), .A4(n7894), .S0(
        n5101), .S1(n7677), .Y(q[40]) );
  MUX41X1_HVT U8870 ( .A1(\ram[1][169] ), .A3(\ram[3][169] ), .A2(
        \ram[0][169] ), .A4(\ram[2][169] ), .S0(n5940), .S1(n7576), .Y(n8408)
         );
  MUX41X1_HVT U8871 ( .A1(n8501), .A3(n8503), .A2(n8502), .A4(n8504), .S0(
        n7685), .S1(n5503), .Y(q[193]) );
  NBUFFX2_HVT U8872 ( .A(n5943), .Y(n7680) );
  MUX41X1_HVT U8873 ( .A1(\ram[15][58] ), .A3(\ram[13][58] ), .A2(
        \ram[14][58] ), .A4(\ram[12][58] ), .S0(n5152), .S1(n5450), .Y(n7963)
         );
  MUX41X1_HVT U8874 ( .A1(\ram[15][147] ), .A3(\ram[13][147] ), .A2(
        \ram[14][147] ), .A4(\ram[12][147] ), .S0(n7682), .S1(n6732), .Y(n8317) );
  MUX41X1_HVT U8875 ( .A1(\ram[15][96] ), .A3(\ram[13][96] ), .A2(
        \ram[14][96] ), .A4(\ram[12][96] ), .S0(n7697), .S1(n4175), .Y(n8114)
         );
  MUX41X1_HVT U8876 ( .A1(\ram[15][38] ), .A3(\ram[13][38] ), .A2(
        \ram[14][38] ), .A4(\ram[12][38] ), .S0(n5647), .S1(n7688), .Y(n7883)
         );
  MUX41X1_HVT U8877 ( .A1(\ram[15][142] ), .A3(\ram[13][142] ), .A2(
        \ram[14][142] ), .A4(\ram[12][142] ), .S0(n6746), .S1(n7699), .Y(n8298) );
  MUX41X1_HVT U8878 ( .A1(\ram[15][7] ), .A3(\ram[13][7] ), .A2(\ram[14][7] ), 
        .A4(\ram[12][7] ), .S0(n7697), .S1(n5735), .Y(n7762) );
  MUX41X1_HVT U8879 ( .A1(\ram[15][139] ), .A3(\ram[13][139] ), .A2(
        \ram[14][139] ), .A4(\ram[12][139] ), .S0(n5594), .S1(n7576), .Y(n8286) );
  MUX41X1_HVT U8880 ( .A1(\ram[15][16] ), .A3(\ram[13][16] ), .A2(
        \ram[14][16] ), .A4(\ram[12][16] ), .S0(n7296), .S1(n5735), .Y(n7798)
         );
  MUX41X1_HVT U8881 ( .A1(\ram[15][223] ), .A3(\ram[13][223] ), .A2(
        \ram[14][223] ), .A4(\ram[12][223] ), .S0(n8787), .S1(n5232), .Y(n8621) );
  MUX41X1_HVT U8882 ( .A1(\ram[15][247] ), .A3(\ram[13][247] ), .A2(
        \ram[14][247] ), .A4(\ram[12][247] ), .S0(n7350), .S1(n7698), .Y(n8715) );
  MUX41X1_HVT U8883 ( .A1(\ram[15][55] ), .A3(\ram[13][55] ), .A2(
        \ram[14][55] ), .A4(\ram[12][55] ), .S0(n6412), .S1(n7699), .Y(n7951)
         );
  MUX41X1_HVT U8884 ( .A1(\ram[13][21] ), .A3(\ram[15][21] ), .A2(
        \ram[12][21] ), .A4(\ram[14][21] ), .S0(n5945), .S1(n7143), .Y(n7816)
         );
  MUX41X1_HVT U8885 ( .A1(\ram[13][69] ), .A3(\ram[15][69] ), .A2(
        \ram[12][69] ), .A4(\ram[14][69] ), .S0(n8827), .S1(n7348), .Y(n8006)
         );
  MUX41X1_HVT U8886 ( .A1(\ram[13][39] ), .A3(\ram[15][39] ), .A2(
        \ram[12][39] ), .A4(\ram[14][39] ), .S0(n7551), .S1(n7345), .Y(n7887)
         );
  MUX41X1_HVT U8887 ( .A1(\ram[13][9] ), .A3(\ram[15][9] ), .A2(\ram[12][9] ), 
        .A4(\ram[14][9] ), .S0(n6020), .S1(n7143), .Y(n7770) );
  MUX41X1_HVT U8888 ( .A1(\ram[11][159] ), .A3(\ram[9][159] ), .A2(
        \ram[10][159] ), .A4(\ram[8][159] ), .S0(n5794), .S1(n5958), .Y(n8366)
         );
  MUX41X1_HVT U8889 ( .A1(\ram[11][217] ), .A3(\ram[9][217] ), .A2(
        \ram[10][217] ), .A4(\ram[8][217] ), .S0(n7556), .S1(n5825), .Y(n8598)
         );
  MUX41X1_HVT U8890 ( .A1(\ram[11][161] ), .A3(\ram[9][161] ), .A2(
        \ram[10][161] ), .A4(\ram[8][161] ), .S0(n5814), .S1(n5899), .Y(n8374)
         );
  MUX41X1_HVT U8891 ( .A1(\ram[11][178] ), .A3(\ram[9][178] ), .A2(
        \ram[10][178] ), .A4(\ram[8][178] ), .S0(n5970), .S1(n7345), .Y(n8442)
         );
  MUX41X1_HVT U8892 ( .A1(\ram[13][197] ), .A3(\ram[15][197] ), .A2(
        \ram[12][197] ), .A4(\ram[14][197] ), .S0(n8805), .S1(n6753), .Y(n8517) );
  MUX41X1_HVT U8893 ( .A1(\ram[13][193] ), .A3(\ram[15][193] ), .A2(
        \ram[12][193] ), .A4(\ram[14][193] ), .S0(n8804), .S1(n5864), .Y(n8501) );
  MUX41X1_HVT U8894 ( .A1(\ram[13][150] ), .A3(\ram[15][150] ), .A2(
        \ram[12][150] ), .A4(\ram[14][150] ), .S0(n4837), .S1(n7294), .Y(n8329) );
  MUX41X1_HVT U8895 ( .A1(\ram[13][162] ), .A3(\ram[15][162] ), .A2(
        \ram[12][162] ), .A4(\ram[14][162] ), .S0(n8844), .S1(n7698), .Y(n8377) );
  MUX41X1_HVT U8896 ( .A1(\ram[13][169] ), .A3(\ram[15][169] ), .A2(
        \ram[12][169] ), .A4(\ram[14][169] ), .S0(n5322), .S1(n4987), .Y(n8405) );
  NBUFFX2_HVT U8897 ( .A(n5105), .Y(n7714) );
  MUX41X1_HVT U8898 ( .A1(\ram[13][161] ), .A3(\ram[15][161] ), .A2(
        \ram[12][161] ), .A4(\ram[14][161] ), .S0(n8832), .S1(n7716), .Y(n8373) );
  INVX0_HVT U8899 ( .A(n10095), .Y(n8982) );
  INVX0_HVT U8900 ( .A(n10095), .Y(n8977) );
  INVX0_HVT U8901 ( .A(n10094), .Y(n8967) );
  INVX0_HVT U8902 ( .A(n10094), .Y(n8966) );
  INVX0_HVT U8903 ( .A(n10097), .Y(n10096) );
  INVX0_HVT U8904 ( .A(n9450), .Y(n9451) );
  INVX0_HVT U8905 ( .A(n9305), .Y(n9306) );
  INVX0_HVT U8906 ( .A(n9314), .Y(n9315) );
  INVX0_HVT U8907 ( .A(n9318), .Y(n9319) );
  INVX0_HVT U8908 ( .A(n9321), .Y(n9322) );
  INVX0_HVT U8909 ( .A(n9324), .Y(n9325) );
  INVX0_HVT U8910 ( .A(n9327), .Y(n9328) );
  INVX0_HVT U8911 ( .A(n9330), .Y(n9331) );
  INVX0_HVT U8912 ( .A(n9333), .Y(n9334) );
  INVX0_HVT U8913 ( .A(n9336), .Y(n9337) );
  INVX0_HVT U8914 ( .A(n9339), .Y(n9340) );
  INVX0_HVT U8915 ( .A(n9343), .Y(n9344) );
  INVX0_HVT U8916 ( .A(n9346), .Y(n9347) );
  INVX0_HVT U8917 ( .A(n9349), .Y(n9350) );
  INVX0_HVT U8918 ( .A(n9352), .Y(n9353) );
  INVX0_HVT U8919 ( .A(n9355), .Y(n9356) );
  INVX0_HVT U8920 ( .A(n9358), .Y(n9359) );
  INVX0_HVT U8921 ( .A(n9361), .Y(n9362) );
  INVX0_HVT U8922 ( .A(n9364), .Y(n9365) );
  INVX0_HVT U8923 ( .A(n9367), .Y(n9368) );
  INVX0_HVT U8924 ( .A(n9369), .Y(n9370) );
  INVX0_HVT U8925 ( .A(n9372), .Y(n9373) );
  INVX0_HVT U8926 ( .A(n9375), .Y(n9376) );
  INVX0_HVT U8927 ( .A(n9378), .Y(n9379) );
  INVX0_HVT U8928 ( .A(n9381), .Y(n9382) );
  INVX0_HVT U8929 ( .A(n9384), .Y(n9385) );
  INVX0_HVT U8930 ( .A(n9387), .Y(n9388) );
  INVX0_HVT U8931 ( .A(n9390), .Y(n9391) );
  INVX0_HVT U8932 ( .A(n9393), .Y(n9394) );
  INVX0_HVT U8933 ( .A(n9396), .Y(n9397) );
  INVX0_HVT U8934 ( .A(n9399), .Y(n9400) );
  INVX0_HVT U8935 ( .A(n9402), .Y(n9403) );
  INVX0_HVT U8936 ( .A(n9405), .Y(n9406) );
  INVX0_HVT U8937 ( .A(n9408), .Y(n9409) );
  INVX0_HVT U8938 ( .A(n9411), .Y(n9412) );
  INVX0_HVT U8939 ( .A(n9414), .Y(n9415) );
  INVX0_HVT U8940 ( .A(n9417), .Y(n9418) );
  INVX0_HVT U8941 ( .A(n9420), .Y(n9421) );
  INVX0_HVT U8942 ( .A(n9423), .Y(n9424) );
  INVX0_HVT U8943 ( .A(n9426), .Y(n9427) );
  INVX0_HVT U8944 ( .A(n9429), .Y(n9430) );
  INVX0_HVT U8945 ( .A(n9432), .Y(n9433) );
  INVX0_HVT U8946 ( .A(n9435), .Y(n9436) );
  INVX0_HVT U8947 ( .A(n9438), .Y(n9439) );
  INVX0_HVT U8948 ( .A(n9441), .Y(n9442) );
  INVX0_HVT U8949 ( .A(n9444), .Y(n9445) );
  INVX0_HVT U8950 ( .A(n9447), .Y(n9448) );
  INVX0_HVT U8951 ( .A(n9453), .Y(n9454) );
  INVX0_HVT U8952 ( .A(n9456), .Y(n9457) );
  INVX0_HVT U8953 ( .A(n9459), .Y(n9460) );
  INVX0_HVT U8954 ( .A(n9462), .Y(n9463) );
  INVX0_HVT U8955 ( .A(n9465), .Y(n9466) );
  INVX0_HVT U8956 ( .A(n9468), .Y(n9469) );
  INVX0_HVT U8957 ( .A(n9471), .Y(n9472) );
  INVX0_HVT U8958 ( .A(n9474), .Y(n9475) );
  INVX0_HVT U8959 ( .A(n9477), .Y(n9478) );
  INVX0_HVT U8960 ( .A(n9480), .Y(n9481) );
  INVX0_HVT U8961 ( .A(n9483), .Y(n9484) );
  INVX0_HVT U8962 ( .A(n9486), .Y(n9487) );
  INVX0_HVT U8963 ( .A(n9489), .Y(n9490) );
  INVX0_HVT U8964 ( .A(n9492), .Y(n9493) );
  INVX0_HVT U8965 ( .A(n9495), .Y(n9496) );
  INVX0_HVT U8966 ( .A(n9498), .Y(n9499) );
  INVX0_HVT U8967 ( .A(n9501), .Y(n9502) );
  INVX0_HVT U8968 ( .A(n9504), .Y(n9505) );
  INVX0_HVT U8969 ( .A(n9507), .Y(n9508) );
  INVX0_HVT U8970 ( .A(n9510), .Y(n9511) );
  INVX0_HVT U8971 ( .A(n9513), .Y(n9514) );
  INVX0_HVT U8972 ( .A(n9516), .Y(n9517) );
  INVX0_HVT U8973 ( .A(n9519), .Y(n9520) );
  INVX0_HVT U8974 ( .A(n9522), .Y(n9523) );
  INVX0_HVT U8975 ( .A(n9525), .Y(n9526) );
  INVX0_HVT U8976 ( .A(n9528), .Y(n9529) );
  INVX0_HVT U8977 ( .A(n9531), .Y(n9532) );
  INVX0_HVT U8978 ( .A(n9534), .Y(n9535) );
  INVX0_HVT U8979 ( .A(n9537), .Y(n9538) );
  INVX0_HVT U8980 ( .A(n9540), .Y(n9541) );
  INVX0_HVT U8981 ( .A(n9543), .Y(n9544) );
  INVX0_HVT U8982 ( .A(n9546), .Y(n9547) );
  INVX0_HVT U8983 ( .A(n9549), .Y(n9550) );
  INVX0_HVT U8984 ( .A(n9552), .Y(n9553) );
  INVX0_HVT U8985 ( .A(n9555), .Y(n9556) );
  INVX0_HVT U8986 ( .A(n9558), .Y(n9559) );
  INVX0_HVT U8987 ( .A(n9561), .Y(n9562) );
  INVX0_HVT U8988 ( .A(n9564), .Y(n9565) );
  INVX0_HVT U8989 ( .A(n9567), .Y(n9568) );
  INVX0_HVT U8990 ( .A(n9570), .Y(n9571) );
  INVX0_HVT U8991 ( .A(n9573), .Y(n9574) );
  INVX0_HVT U8992 ( .A(n9576), .Y(n9577) );
  INVX0_HVT U8993 ( .A(n9579), .Y(n9580) );
  INVX0_HVT U8994 ( .A(n9582), .Y(n9583) );
  INVX0_HVT U8995 ( .A(n9585), .Y(n9586) );
  INVX0_HVT U8996 ( .A(n9588), .Y(n9589) );
  INVX0_HVT U8997 ( .A(n9591), .Y(n9592) );
  INVX0_HVT U8998 ( .A(n9594), .Y(n9595) );
  INVX0_HVT U8999 ( .A(n9597), .Y(n9598) );
  INVX0_HVT U9000 ( .A(n9600), .Y(n9601) );
  INVX0_HVT U9001 ( .A(n9603), .Y(n9604) );
  INVX0_HVT U9002 ( .A(n9606), .Y(n9607) );
  INVX0_HVT U9003 ( .A(n9609), .Y(n9610) );
  INVX0_HVT U9004 ( .A(n9612), .Y(n9613) );
  INVX0_HVT U9005 ( .A(n9615), .Y(n9616) );
  INVX0_HVT U9006 ( .A(n9618), .Y(n9619) );
  INVX0_HVT U9007 ( .A(n9621), .Y(n9622) );
  INVX0_HVT U9008 ( .A(n9624), .Y(n9625) );
  INVX0_HVT U9009 ( .A(n9627), .Y(n9628) );
  INVX0_HVT U9010 ( .A(n9630), .Y(n9631) );
  INVX0_HVT U9011 ( .A(n9633), .Y(n9634) );
  INVX0_HVT U9012 ( .A(n9636), .Y(n9637) );
  INVX0_HVT U9013 ( .A(n9639), .Y(n9640) );
  INVX0_HVT U9014 ( .A(n9642), .Y(n9643) );
  INVX0_HVT U9015 ( .A(n9645), .Y(n9646) );
  INVX0_HVT U9016 ( .A(n9648), .Y(n9649) );
  INVX0_HVT U9017 ( .A(n9651), .Y(n9652) );
  INVX0_HVT U9018 ( .A(n9654), .Y(n9655) );
  INVX0_HVT U9019 ( .A(n9657), .Y(n9658) );
  INVX0_HVT U9020 ( .A(n9660), .Y(n9661) );
  INVX0_HVT U9021 ( .A(n9663), .Y(n9664) );
  INVX0_HVT U9022 ( .A(n9666), .Y(n9667) );
  INVX0_HVT U9023 ( .A(n9669), .Y(n9670) );
  INVX0_HVT U9024 ( .A(n9672), .Y(n9673) );
  INVX0_HVT U9025 ( .A(n9675), .Y(n9676) );
  INVX0_HVT U9026 ( .A(n9678), .Y(n9679) );
  INVX0_HVT U9027 ( .A(n9681), .Y(n9682) );
  INVX0_HVT U9028 ( .A(n9684), .Y(n9685) );
  INVX0_HVT U9029 ( .A(n9687), .Y(n9688) );
  INVX0_HVT U9030 ( .A(n9690), .Y(n9691) );
  INVX0_HVT U9031 ( .A(n9693), .Y(n9694) );
  INVX0_HVT U9032 ( .A(n9696), .Y(n9697) );
  INVX0_HVT U9033 ( .A(n9699), .Y(n9700) );
  INVX0_HVT U9034 ( .A(n9702), .Y(n9703) );
  INVX0_HVT U9035 ( .A(n9705), .Y(n9706) );
  INVX0_HVT U9036 ( .A(n9708), .Y(n9709) );
  INVX0_HVT U9037 ( .A(n9711), .Y(n9712) );
  INVX0_HVT U9038 ( .A(n9714), .Y(n9715) );
  INVX0_HVT U9039 ( .A(n9717), .Y(n9718) );
  INVX0_HVT U9040 ( .A(n9720), .Y(n9721) );
  INVX0_HVT U9041 ( .A(n9723), .Y(n9724) );
  INVX0_HVT U9042 ( .A(n9727), .Y(n9728) );
  INVX0_HVT U9043 ( .A(n9730), .Y(n9731) );
  INVX0_HVT U9044 ( .A(n9733), .Y(n9734) );
  INVX0_HVT U9045 ( .A(n9736), .Y(n9737) );
  INVX0_HVT U9046 ( .A(n9740), .Y(n9741) );
  INVX0_HVT U9047 ( .A(n9743), .Y(n9744) );
  INVX0_HVT U9048 ( .A(n9746), .Y(n9747) );
  INVX0_HVT U9049 ( .A(n9749), .Y(n9750) );
  INVX0_HVT U9050 ( .A(n9753), .Y(n9754) );
  INVX0_HVT U9051 ( .A(n9756), .Y(n9757) );
  INVX0_HVT U9052 ( .A(n9759), .Y(n9760) );
  INVX0_HVT U9053 ( .A(n9762), .Y(n9763) );
  INVX0_HVT U9054 ( .A(n9765), .Y(n9766) );
  INVX0_HVT U9055 ( .A(n9768), .Y(n9769) );
  INVX0_HVT U9056 ( .A(n9771), .Y(n9772) );
  INVX0_HVT U9057 ( .A(n9774), .Y(n9775) );
  INVX0_HVT U9058 ( .A(n9778), .Y(n9779) );
  INVX0_HVT U9059 ( .A(n9781), .Y(n9782) );
  INVX0_HVT U9060 ( .A(n9784), .Y(n9785) );
  INVX0_HVT U9061 ( .A(n9787), .Y(n9788) );
  INVX0_HVT U9062 ( .A(n9791), .Y(n9792) );
  INVX0_HVT U9063 ( .A(n9794), .Y(n9795) );
  INVX0_HVT U9064 ( .A(n9797), .Y(n9798) );
  INVX0_HVT U9065 ( .A(n9800), .Y(n9801) );
  INVX0_HVT U9066 ( .A(n9803), .Y(n9804) );
  INVX0_HVT U9067 ( .A(n9806), .Y(n9807) );
  INVX0_HVT U9068 ( .A(n9809), .Y(n9810) );
  INVX0_HVT U9069 ( .A(n9812), .Y(n9813) );
  INVX0_HVT U9070 ( .A(n9815), .Y(n9816) );
  INVX0_HVT U9071 ( .A(n9818), .Y(n9819) );
  INVX0_HVT U9072 ( .A(n9821), .Y(n9822) );
  INVX0_HVT U9073 ( .A(n9824), .Y(n9825) );
  INVX0_HVT U9074 ( .A(n9828), .Y(n9829) );
  INVX0_HVT U9075 ( .A(n9831), .Y(n9832) );
  INVX0_HVT U9076 ( .A(n9834), .Y(n9835) );
  INVX0_HVT U9077 ( .A(n9837), .Y(n9838) );
  INVX0_HVT U9078 ( .A(n9841), .Y(n9842) );
  INVX0_HVT U9079 ( .A(n9844), .Y(n9845) );
  INVX0_HVT U9080 ( .A(n9847), .Y(n9848) );
  INVX0_HVT U9081 ( .A(n9850), .Y(n9851) );
  INVX0_HVT U9082 ( .A(n9854), .Y(n9855) );
  INVX0_HVT U9083 ( .A(n9857), .Y(n9858) );
  INVX0_HVT U9084 ( .A(n9860), .Y(n9861) );
  INVX0_HVT U9085 ( .A(n9863), .Y(n9864) );
  INVX0_HVT U9086 ( .A(n9867), .Y(n9868) );
  INVX0_HVT U9087 ( .A(n9870), .Y(n9871) );
  INVX0_HVT U9088 ( .A(n9873), .Y(n9874) );
  INVX0_HVT U9089 ( .A(n9876), .Y(n9877) );
  INVX0_HVT U9090 ( .A(n9879), .Y(n9880) );
  INVX0_HVT U9091 ( .A(n9882), .Y(n9883) );
  INVX0_HVT U9092 ( .A(n9885), .Y(n9886) );
  INVX0_HVT U9093 ( .A(n9888), .Y(n9889) );
  INVX0_HVT U9094 ( .A(n9892), .Y(n9893) );
  INVX0_HVT U9095 ( .A(n9895), .Y(n9896) );
  INVX0_HVT U9096 ( .A(n9898), .Y(n9899) );
  INVX0_HVT U9097 ( .A(n9901), .Y(n9902) );
  INVX0_HVT U9098 ( .A(n9905), .Y(n9906) );
  INVX0_HVT U9099 ( .A(n9908), .Y(n9909) );
  INVX0_HVT U9100 ( .A(n9911), .Y(n9912) );
  INVX0_HVT U9101 ( .A(n9914), .Y(n9915) );
  INVX0_HVT U9102 ( .A(n9918), .Y(n9919) );
  INVX0_HVT U9103 ( .A(n9921), .Y(n9922) );
  INVX0_HVT U9104 ( .A(n9924), .Y(n9925) );
  INVX0_HVT U9105 ( .A(n9930), .Y(n9931) );
  INVX0_HVT U9106 ( .A(n9933), .Y(n9934) );
  INVX0_HVT U9107 ( .A(n9936), .Y(n9937) );
  INVX0_HVT U9108 ( .A(n9939), .Y(n9940) );
  INVX0_HVT U9109 ( .A(n9943), .Y(n9944) );
  INVX0_HVT U9110 ( .A(n9946), .Y(n9947) );
  INVX0_HVT U9111 ( .A(n9949), .Y(n9950) );
  INVX0_HVT U9112 ( .A(n9952), .Y(n9953) );
  INVX0_HVT U9113 ( .A(n9955), .Y(n9956) );
  INVX0_HVT U9114 ( .A(n9958), .Y(n9959) );
  INVX0_HVT U9115 ( .A(n9961), .Y(n9962) );
  INVX0_HVT U9116 ( .A(n9964), .Y(n9965) );
  INVX0_HVT U9117 ( .A(n9967), .Y(n9968) );
  INVX0_HVT U9118 ( .A(n9970), .Y(n9971) );
  INVX0_HVT U9119 ( .A(n9973), .Y(n9974) );
  INVX0_HVT U9120 ( .A(n9976), .Y(n9977) );
  INVX0_HVT U9121 ( .A(n9980), .Y(n9981) );
  INVX0_HVT U9122 ( .A(n9983), .Y(n9984) );
  INVX0_HVT U9123 ( .A(n9986), .Y(n9987) );
  INVX0_HVT U9124 ( .A(n9989), .Y(n9990) );
  INVX0_HVT U9125 ( .A(n9992), .Y(n9993) );
  INVX0_HVT U9126 ( .A(n9995), .Y(n9996) );
  INVX0_HVT U9127 ( .A(n9998), .Y(n9999) );
  INVX0_HVT U9128 ( .A(n10001), .Y(n10002) );
  INVX0_HVT U9129 ( .A(n10004), .Y(n10005) );
  INVX0_HVT U9130 ( .A(n10007), .Y(n10008) );
  INVX0_HVT U9131 ( .A(n10010), .Y(n10011) );
  INVX0_HVT U9132 ( .A(n10013), .Y(n10014) );
  INVX0_HVT U9133 ( .A(n10017), .Y(n10018) );
  INVX0_HVT U9134 ( .A(n10020), .Y(n10021) );
  INVX0_HVT U9135 ( .A(n10023), .Y(n10024) );
  INVX0_HVT U9136 ( .A(n10026), .Y(n10027) );
  INVX0_HVT U9137 ( .A(n10029), .Y(n10030) );
  INVX0_HVT U9138 ( .A(n10032), .Y(n10033) );
  INVX0_HVT U9139 ( .A(n10035), .Y(n10036) );
  INVX0_HVT U9140 ( .A(n10038), .Y(n10039) );
  INVX0_HVT U9141 ( .A(n10042), .Y(n10043) );
  INVX0_HVT U9142 ( .A(n10045), .Y(n10046) );
  INVX0_HVT U9143 ( .A(n10048), .Y(n10049) );
  INVX0_HVT U9144 ( .A(n10051), .Y(n10052) );
  INVX0_HVT U9145 ( .A(n10054), .Y(n10055) );
  INVX0_HVT U9146 ( .A(n10057), .Y(n10058) );
  INVX0_HVT U9147 ( .A(n10060), .Y(n10061) );
  INVX0_HVT U9148 ( .A(n10063), .Y(n10064) );
  INVX0_HVT U9149 ( .A(n10067), .Y(n10068) );
  INVX0_HVT U9150 ( .A(n10070), .Y(n10071) );
  INVX0_HVT U9151 ( .A(n10073), .Y(n10074) );
  INVX0_HVT U9152 ( .A(n10076), .Y(n10077) );
  INVX0_HVT U9153 ( .A(n10080), .Y(n10081) );
  INVX0_HVT U9154 ( .A(n10083), .Y(n10084) );
  INVX0_HVT U9155 ( .A(n10086), .Y(n10087) );
  INVX0_HVT U9156 ( .A(n10089), .Y(n10090) );
  INVX0_HVT U9157 ( .A(data[144]), .Y(n9740) );
  INVX0_HVT U9158 ( .A(data[216]), .Y(n9967) );
  INVX0_HVT U9159 ( .A(data[145]), .Y(n9743) );
  INVX0_HVT U9160 ( .A(data[146]), .Y(n9746) );
  INVX0_HVT U9161 ( .A(data[147]), .Y(n9749) );
  INVX0_HVT U9162 ( .A(data[148]), .Y(n9753) );
  INVX0_HVT U9163 ( .A(data[149]), .Y(n9756) );
  INVX0_HVT U9164 ( .A(data[150]), .Y(n9759) );
  INVX0_HVT U9165 ( .A(data[151]), .Y(n9762) );
  INVX0_HVT U9166 ( .A(data[152]), .Y(n9765) );
  INVX0_HVT U9167 ( .A(data[153]), .Y(n9768) );
  INVX0_HVT U9168 ( .A(data[154]), .Y(n9771) );
  INVX0_HVT U9169 ( .A(data[155]), .Y(n9774) );
  INVX0_HVT U9170 ( .A(data[228]), .Y(n10004) );
  INVX0_HVT U9171 ( .A(data[229]), .Y(n10007) );
  INVX0_HVT U9172 ( .A(data[230]), .Y(n10010) );
  INVX0_HVT U9173 ( .A(data[231]), .Y(n10013) );
  INVX0_HVT U9174 ( .A(data[232]), .Y(n10017) );
  INVX0_HVT U9175 ( .A(data[233]), .Y(n10020) );
  INVX0_HVT U9176 ( .A(data[234]), .Y(n10023) );
  INVX0_HVT U9177 ( .A(data[235]), .Y(n10026) );
  INVX0_HVT U9178 ( .A(data[236]), .Y(n10029) );
  INVX0_HVT U9179 ( .A(data[237]), .Y(n10032) );
  INVX0_HVT U9180 ( .A(data[238]), .Y(n10035) );
  INVX0_HVT U9181 ( .A(data[239]), .Y(n10038) );
  INVX0_HVT U9182 ( .A(data[73]), .Y(n9525) );
  INVX0_HVT U9183 ( .A(data[74]), .Y(n9528) );
  INVX0_HVT U9184 ( .A(data[75]), .Y(n9531) );
  INVX0_HVT U9185 ( .A(data[76]), .Y(n9534) );
  INVX0_HVT U9186 ( .A(data[77]), .Y(n9537) );
  INVX0_HVT U9187 ( .A(data[78]), .Y(n9540) );
  INVX0_HVT U9188 ( .A(data[79]), .Y(n9543) );
  INVX0_HVT U9189 ( .A(data[80]), .Y(n9546) );
  INVX0_HVT U9190 ( .A(data[81]), .Y(n9549) );
  INVX0_HVT U9191 ( .A(data[82]), .Y(n9552) );
  INVX0_HVT U9192 ( .A(data[83]), .Y(n9555) );
  INVX0_HVT U9193 ( .A(data[84]), .Y(n9558) );
  INVX0_HVT U9194 ( .A(data[85]), .Y(n9561) );
  INVX0_HVT U9195 ( .A(data[86]), .Y(n9564) );
  INVX0_HVT U9196 ( .A(data[87]), .Y(n9567) );
  INVX0_HVT U9197 ( .A(data[89]), .Y(n9573) );
  INVX0_HVT U9198 ( .A(data[90]), .Y(n9576) );
  INVX0_HVT U9199 ( .A(data[91]), .Y(n9579) );
  INVX0_HVT U9200 ( .A(data[92]), .Y(n9582) );
  INVX0_HVT U9201 ( .A(data[93]), .Y(n9585) );
  INVX0_HVT U9202 ( .A(data[94]), .Y(n9588) );
  INVX0_HVT U9203 ( .A(data[95]), .Y(n9591) );
  INVX0_HVT U9204 ( .A(data[96]), .Y(n9594) );
  INVX0_HVT U9205 ( .A(data[97]), .Y(n9597) );
  INVX0_HVT U9206 ( .A(data[98]), .Y(n9600) );
  INVX0_HVT U9207 ( .A(data[99]), .Y(n9603) );
  INVX0_HVT U9208 ( .A(data[100]), .Y(n9606) );
  INVX0_HVT U9209 ( .A(data[101]), .Y(n9609) );
  INVX0_HVT U9210 ( .A(data[102]), .Y(n9612) );
  INVX0_HVT U9211 ( .A(data[103]), .Y(n9615) );
  INVX0_HVT U9212 ( .A(data[104]), .Y(n9618) );
  INVX0_HVT U9213 ( .A(data[105]), .Y(n9621) );
  INVX0_HVT U9214 ( .A(data[106]), .Y(n9624) );
  INVX0_HVT U9215 ( .A(data[107]), .Y(n9627) );
  INVX0_HVT U9216 ( .A(data[192]), .Y(n9892) );
  INVX0_HVT U9217 ( .A(data[193]), .Y(n9895) );
  INVX0_HVT U9218 ( .A(data[194]), .Y(n9898) );
  INVX0_HVT U9219 ( .A(data[196]), .Y(n9905) );
  INVX0_HVT U9220 ( .A(data[197]), .Y(n9908) );
  INVX0_HVT U9221 ( .A(data[198]), .Y(n9911) );
  INVX0_HVT U9222 ( .A(data[199]), .Y(n9914) );
  INVX0_HVT U9223 ( .A(data[200]), .Y(n9918) );
  INVX0_HVT U9224 ( .A(data[202]), .Y(n9924) );
  INVX0_HVT U9225 ( .A(data[203]), .Y(n9927) );
  INVX0_HVT U9226 ( .A(data[205]), .Y(n9933) );
  INVX0_HVT U9227 ( .A(data[206]), .Y(n9936) );
  INVX0_HVT U9228 ( .A(data[207]), .Y(n9939) );
  INVX0_HVT U9229 ( .A(data[208]), .Y(n9943) );
  INVX0_HVT U9230 ( .A(data[209]), .Y(n9946) );
  INVX0_HVT U9231 ( .A(data[210]), .Y(n9949) );
  INVX0_HVT U9232 ( .A(data[211]), .Y(n9952) );
  INVX0_HVT U9233 ( .A(data[212]), .Y(n9955) );
  INVX0_HVT U9234 ( .A(data[214]), .Y(n9961) );
  INVX0_HVT U9235 ( .A(data[215]), .Y(n9964) );
  INVX0_HVT U9236 ( .A(data[218]), .Y(n9973) );
  INVX0_HVT U9237 ( .A(data[219]), .Y(n9976) );
  INVX0_HVT U9238 ( .A(data[220]), .Y(n9980) );
  INVX0_HVT U9239 ( .A(data[221]), .Y(n9983) );
  INVX0_HVT U9240 ( .A(data[222]), .Y(n9986) );
  INVX0_HVT U9241 ( .A(data[223]), .Y(n9989) );
  INVX0_HVT U9242 ( .A(data[224]), .Y(n9992) );
  INVX0_HVT U9243 ( .A(data[225]), .Y(n9995) );
  INVX0_HVT U9244 ( .A(data[226]), .Y(n9998) );
  INVX0_HVT U9245 ( .A(data[227]), .Y(n10001) );
  INVX0_HVT U9246 ( .A(data[240]), .Y(n10042) );
  INVX0_HVT U9247 ( .A(data[241]), .Y(n10045) );
  INVX0_HVT U9248 ( .A(data[242]), .Y(n10048) );
  INVX0_HVT U9249 ( .A(data[243]), .Y(n10051) );
  INVX0_HVT U9250 ( .A(data[244]), .Y(n10054) );
  INVX0_HVT U9251 ( .A(data[245]), .Y(n10057) );
  INVX0_HVT U9252 ( .A(data[246]), .Y(n10060) );
  INVX0_HVT U9253 ( .A(data[247]), .Y(n10063) );
  INVX0_HVT U9254 ( .A(data[248]), .Y(n10067) );
  INVX0_HVT U9255 ( .A(data[249]), .Y(n10070) );
  INVX0_HVT U9256 ( .A(data[250]), .Y(n10073) );
  INVX0_HVT U9257 ( .A(data[251]), .Y(n10076) );
  INVX0_HVT U9258 ( .A(data[120]), .Y(n9666) );
  INVX0_HVT U9259 ( .A(data[121]), .Y(n9669) );
  INVX0_HVT U9260 ( .A(data[122]), .Y(n9672) );
  INVX0_HVT U9261 ( .A(data[123]), .Y(n9675) );
  INVX0_HVT U9262 ( .A(data[124]), .Y(n9678) );
  INVX0_HVT U9263 ( .A(data[125]), .Y(n9681) );
  INVX0_HVT U9264 ( .A(data[126]), .Y(n9684) );
  INVX0_HVT U9265 ( .A(data[127]), .Y(n9687) );
  INVX0_HVT U9266 ( .A(data[128]), .Y(n9690) );
  INVX0_HVT U9267 ( .A(data[129]), .Y(n9693) );
  INVX0_HVT U9268 ( .A(data[130]), .Y(n9696) );
  INVX0_HVT U9269 ( .A(data[131]), .Y(n9699) );
  INVX0_HVT U9270 ( .A(data[132]), .Y(n9702) );
  INVX0_HVT U9271 ( .A(data[133]), .Y(n9705) );
  INVX0_HVT U9272 ( .A(data[134]), .Y(n9708) );
  INVX0_HVT U9273 ( .A(data[135]), .Y(n9711) );
  INVX0_HVT U9274 ( .A(data[136]), .Y(n9714) );
  INVX0_HVT U9275 ( .A(data[137]), .Y(n9717) );
  INVX0_HVT U9276 ( .A(data[138]), .Y(n9720) );
  INVX0_HVT U9277 ( .A(data[140]), .Y(n9727) );
  INVX0_HVT U9278 ( .A(data[141]), .Y(n9730) );
  INVX0_HVT U9279 ( .A(data[142]), .Y(n9733) );
  INVX0_HVT U9280 ( .A(data[143]), .Y(n9736) );
  INVX0_HVT U9281 ( .A(data[1]), .Y(n9308) );
  INVX0_HVT U9282 ( .A(data[2]), .Y(n9311) );
  INVX0_HVT U9283 ( .A(data[3]), .Y(n9314) );
  INVX0_HVT U9284 ( .A(data[4]), .Y(n9318) );
  INVX0_HVT U9285 ( .A(data[6]), .Y(n9324) );
  INVX0_HVT U9286 ( .A(data[7]), .Y(n9327) );
  INVX0_HVT U9287 ( .A(data[10]), .Y(n9336) );
  INVX0_HVT U9288 ( .A(data[11]), .Y(n9339) );
  INVX0_HVT U9289 ( .A(data[12]), .Y(n9343) );
  INVX0_HVT U9290 ( .A(data[13]), .Y(n9346) );
  INVX0_HVT U9291 ( .A(data[14]), .Y(n9349) );
  INVX0_HVT U9292 ( .A(data[15]), .Y(n9352) );
  INVX0_HVT U9293 ( .A(data[17]), .Y(n9358) );
  INVX0_HVT U9294 ( .A(data[19]), .Y(n9364) );
  INVX0_HVT U9295 ( .A(data[20]), .Y(n9367) );
  INVX0_HVT U9296 ( .A(data[22]), .Y(n9372) );
  INVX0_HVT U9297 ( .A(data[23]), .Y(n9375) );
  INVX0_HVT U9298 ( .A(data[24]), .Y(n9378) );
  INVX0_HVT U9299 ( .A(data[26]), .Y(n9384) );
  INVX0_HVT U9300 ( .A(data[28]), .Y(n9390) );
  INVX0_HVT U9301 ( .A(data[30]), .Y(n9396) );
  INVX0_HVT U9302 ( .A(data[31]), .Y(n9399) );
  INVX0_HVT U9303 ( .A(data[32]), .Y(n9402) );
  INVX0_HVT U9304 ( .A(data[33]), .Y(n9405) );
  INVX0_HVT U9305 ( .A(data[34]), .Y(n9408) );
  INVX0_HVT U9306 ( .A(data[35]), .Y(n9411) );
  INVX0_HVT U9307 ( .A(data[36]), .Y(n9414) );
  INVX0_HVT U9308 ( .A(data[37]), .Y(n9417) );
  INVX0_HVT U9309 ( .A(data[38]), .Y(n9420) );
  INVX0_HVT U9310 ( .A(data[39]), .Y(n9423) );
  INVX0_HVT U9311 ( .A(data[40]), .Y(n9426) );
  INVX0_HVT U9312 ( .A(data[41]), .Y(n9429) );
  INVX0_HVT U9313 ( .A(data[43]), .Y(n9435) );
  INVX0_HVT U9314 ( .A(data[44]), .Y(n9438) );
  INVX0_HVT U9315 ( .A(data[45]), .Y(n9441) );
  INVX0_HVT U9316 ( .A(data[46]), .Y(n9444) );
  INVX0_HVT U9317 ( .A(data[47]), .Y(n9447) );
  INVX0_HVT U9318 ( .A(data[60]), .Y(n9486) );
  INVX0_HVT U9319 ( .A(data[61]), .Y(n9489) );
  INVX0_HVT U9320 ( .A(data[62]), .Y(n9492) );
  INVX0_HVT U9321 ( .A(data[63]), .Y(n9495) );
  INVX0_HVT U9322 ( .A(data[64]), .Y(n9498) );
  INVX0_HVT U9323 ( .A(data[65]), .Y(n9501) );
  INVX0_HVT U9324 ( .A(data[66]), .Y(n9504) );
  INVX0_HVT U9325 ( .A(data[67]), .Y(n9507) );
  INVX0_HVT U9326 ( .A(data[68]), .Y(n9510) );
  INVX0_HVT U9327 ( .A(data[69]), .Y(n9513) );
  INVX0_HVT U9328 ( .A(data[70]), .Y(n9516) );
  INVX0_HVT U9329 ( .A(data[71]), .Y(n9519) );
  INVX0_HVT U9330 ( .A(data[108]), .Y(n9630) );
  INVX0_HVT U9331 ( .A(data[109]), .Y(n9633) );
  INVX0_HVT U9332 ( .A(data[110]), .Y(n9636) );
  INVX0_HVT U9333 ( .A(data[111]), .Y(n9639) );
  INVX0_HVT U9334 ( .A(data[112]), .Y(n9642) );
  INVX0_HVT U9335 ( .A(data[113]), .Y(n9645) );
  INVX0_HVT U9336 ( .A(data[114]), .Y(n9648) );
  INVX0_HVT U9337 ( .A(data[115]), .Y(n9651) );
  INVX0_HVT U9338 ( .A(data[116]), .Y(n9654) );
  INVX0_HVT U9339 ( .A(data[117]), .Y(n9657) );
  INVX0_HVT U9340 ( .A(data[119]), .Y(n9663) );
  INVX0_HVT U9341 ( .A(data[156]), .Y(n9778) );
  INVX0_HVT U9342 ( .A(data[157]), .Y(n9781) );
  INVX0_HVT U9343 ( .A(data[158]), .Y(n9784) );
  INVX0_HVT U9344 ( .A(data[159]), .Y(n9787) );
  INVX0_HVT U9345 ( .A(data[160]), .Y(n9791) );
  INVX0_HVT U9346 ( .A(data[161]), .Y(n9794) );
  INVX0_HVT U9347 ( .A(data[162]), .Y(n9797) );
  INVX0_HVT U9348 ( .A(data[163]), .Y(n9800) );
  INVX0_HVT U9349 ( .A(data[164]), .Y(n9803) );
  INVX0_HVT U9350 ( .A(data[165]), .Y(n9806) );
  INVX0_HVT U9351 ( .A(data[166]), .Y(n9809) );
  INVX0_HVT U9352 ( .A(data[167]), .Y(n9812) );
  INVX0_HVT U9353 ( .A(data[168]), .Y(n9815) );
  INVX0_HVT U9354 ( .A(data[169]), .Y(n9818) );
  INVX0_HVT U9355 ( .A(data[170]), .Y(n9821) );
  INVX0_HVT U9356 ( .A(data[171]), .Y(n9824) );
  INVX0_HVT U9357 ( .A(data[172]), .Y(n9828) );
  INVX0_HVT U9358 ( .A(data[173]), .Y(n9831) );
  INVX0_HVT U9359 ( .A(data[174]), .Y(n9834) );
  INVX0_HVT U9360 ( .A(data[176]), .Y(n9841) );
  INVX0_HVT U9361 ( .A(data[177]), .Y(n9844) );
  INVX0_HVT U9362 ( .A(data[178]), .Y(n9847) );
  INVX0_HVT U9363 ( .A(data[179]), .Y(n9850) );
  INVX0_HVT U9364 ( .A(data[180]), .Y(n9854) );
  INVX0_HVT U9365 ( .A(data[181]), .Y(n9857) );
  INVX0_HVT U9366 ( .A(data[182]), .Y(n9860) );
  INVX0_HVT U9367 ( .A(data[183]), .Y(n9863) );
  INVX0_HVT U9368 ( .A(data[184]), .Y(n9867) );
  INVX0_HVT U9369 ( .A(data[185]), .Y(n9870) );
  INVX0_HVT U9370 ( .A(data[186]), .Y(n9873) );
  INVX0_HVT U9371 ( .A(data[187]), .Y(n9876) );
  INVX0_HVT U9372 ( .A(data[188]), .Y(n9879) );
  INVX0_HVT U9373 ( .A(data[189]), .Y(n9882) );
  INVX0_HVT U9374 ( .A(data[190]), .Y(n9885) );
  INVX0_HVT U9375 ( .A(data[191]), .Y(n9888) );
  INVX0_HVT U9376 ( .A(data[50]), .Y(n9456) );
  INVX0_HVT U9377 ( .A(data[52]), .Y(n9462) );
  INVX0_HVT U9378 ( .A(data[55]), .Y(n9471) );
  INVX0_HVT U9379 ( .A(data[56]), .Y(n9474) );
  INVX0_HVT U9380 ( .A(data[57]), .Y(n9477) );
  INVX0_HVT U9381 ( .A(data[58]), .Y(n9480) );
  INVX0_HVT U9382 ( .A(data[59]), .Y(n9483) );
  INVX0_HVT U9383 ( .A(data[253]), .Y(n10083) );
  INVX0_HVT U9384 ( .A(data[254]), .Y(n10086) );
  INVX0_HVT U9385 ( .A(data[255]), .Y(n10089) );
  NBUFFX2_HVT U9386 ( .A(n8922), .Y(n8912) );
  NBUFFX2_HVT U9387 ( .A(n8916), .Y(n8913) );
  NBUFFX2_HVT U9388 ( .A(n8921), .Y(n8924) );
  NBUFFX2_HVT U9389 ( .A(n8921), .Y(n8923) );
  NBUFFX2_HVT U9390 ( .A(n8989), .Y(n8993) );
  NBUFFX2_HVT U9391 ( .A(n8989), .Y(n8992) );
  NBUFFX2_HVT U9392 ( .A(n8988), .Y(n8991) );
  NBUFFX2_HVT U9393 ( .A(n8988), .Y(n8990) );
  NBUFFX2_HVT U9394 ( .A(n9047), .Y(n9051) );
  NBUFFX2_HVT U9395 ( .A(n9047), .Y(n9050) );
  NBUFFX2_HVT U9396 ( .A(n4302), .Y(n9049) );
  NBUFFX2_HVT U9397 ( .A(n4302), .Y(n9048) );
  NBUFFX2_HVT U9398 ( .A(n9041), .Y(n9045) );
  NBUFFX2_HVT U9399 ( .A(n9041), .Y(n9044) );
  NBUFFX2_HVT U9400 ( .A(n9040), .Y(n9043) );
  NBUFFX2_HVT U9401 ( .A(n9040), .Y(n9042) );
  NBUFFX2_HVT U9402 ( .A(n9034), .Y(n9037) );
  NBUFFX2_HVT U9403 ( .A(n9034), .Y(n9036) );
  NBUFFX2_HVT U9404 ( .A(n8982), .Y(n8985) );
  NBUFFX2_HVT U9405 ( .A(n8982), .Y(n8984) );
  NBUFFX2_HVT U9406 ( .A(n8977), .Y(n8978) );
  NBUFFX2_HVT U9407 ( .A(n8989), .Y(n8981) );
  NBUFFX2_HVT U9408 ( .A(n8988), .Y(n8980) );
  NBUFFX2_HVT U9409 ( .A(n8977), .Y(n8979) );
  NBUFFX2_HVT U9410 ( .A(n8982), .Y(n8969) );
  NBUFFX2_HVT U9411 ( .A(n8982), .Y(n8968) );
  NBUFFX2_HVT U9412 ( .A(n4302), .Y(n9027) );
  NBUFFX2_HVT U9413 ( .A(n9025), .Y(n9026) );
  INVX1_HVT U9414 ( .A(n10270), .Y(n9218) );
  INVX1_HVT U9415 ( .A(n10254), .Y(n9160) );
  INVX0_HVT U9416 ( .A(n10093), .Y(n8989) );
  INVX0_HVT U9417 ( .A(n10093), .Y(n8988) );
  INVX1_HVT U9418 ( .A(n10114), .Y(n9040) );
  INVX0_HVT U9419 ( .A(n10093), .Y(n8983) );
  INVX1_HVT U9420 ( .A(n10271), .Y(n9212) );
  INVX1_HVT U9421 ( .A(n10271), .Y(n9211) );
  INVX0_HVT U9422 ( .A(n10272), .Y(n10270) );
  INVX0_HVT U9423 ( .A(n10255), .Y(n10253) );
  INVX0_HVT U9424 ( .A(n10255), .Y(n10254) );
  INVX0_HVT U9425 ( .A(n10272), .Y(n10271) );
  INVX0_HVT U9426 ( .A(n7723), .Y(n10340) );
  INVX0_HVT U9427 ( .A(n10346), .Y(n10341) );
  INVX0_HVT U9428 ( .A(n6826), .Y(n10342) );
  INVX0_HVT U9429 ( .A(n6855), .Y(n10343) );
  INVX0_HVT U9430 ( .A(n6855), .Y(n10344) );
  INVX0_HVT U9431 ( .A(n10328), .Y(n10326) );
  INVX0_HVT U9432 ( .A(n10328), .Y(n10327) );
  INVX0_HVT U9433 ( .A(n10300), .Y(n10298) );
  INVX0_HVT U9434 ( .A(n10300), .Y(n10299) );
  INVX0_HVT U9435 ( .A(n10126), .Y(n10125) );
  NBUFFX2_HVT U9436 ( .A(n5938), .Y(n8776) );
  INVX0_HVT U9437 ( .A(n10148), .Y(n10141) );
  INVX0_HVT U9438 ( .A(n10147), .Y(n10142) );
  INVX0_HVT U9439 ( .A(n10361), .Y(n10360) );
  INVX0_HVT U9440 ( .A(n10303), .Y(n10302) );
  INVX0_HVT U9441 ( .A(n10347), .Y(n10346) );
  INVX0_HVT U9442 ( .A(n10303), .Y(n10301) );
  INVX0_HVT U9443 ( .A(n10147), .Y(n10135) );
  INVX0_HVT U9444 ( .A(n10148), .Y(n10136) );
  INVX0_HVT U9445 ( .A(n7586), .Y(n10210) );
  INVX0_HVT U9446 ( .A(n4613), .Y(n10211) );
  INVX0_HVT U9447 ( .A(n7616), .Y(n10212) );
  INVX0_HVT U9448 ( .A(n6901), .Y(n10260) );
  INVX0_HVT U9449 ( .A(n6909), .Y(n10261) );
  INVX0_HVT U9450 ( .A(n6578), .Y(n10143) );
  INVX0_HVT U9451 ( .A(n10190), .Y(n10189) );
  INVX0_HVT U9452 ( .A(n6611), .Y(n10139) );
  INVX0_HVT U9453 ( .A(n10164), .Y(n10163) );
  INVX0_HVT U9454 ( .A(n59), .Y(n10097) );
  INVX0_HVT U9455 ( .A(n59), .Y(n8994) );
  INVX0_HVT U9456 ( .A(n59), .Y(n8995) );
  INVX0_HVT U9457 ( .A(n56), .Y(n9052) );
  INVX0_HVT U9458 ( .A(n4216), .Y(n9224) );
  INVX0_HVT U9459 ( .A(n4216), .Y(n9223) );
  INVX0_HVT U9460 ( .A(n33), .Y(n9166) );
  INVX0_HVT U9461 ( .A(n33), .Y(n9165) );
  INVX0_HVT U9462 ( .A(n40), .Y(n9111) );
  INVX0_HVT U9463 ( .A(n40), .Y(n9110) );
  INVX0_HVT U9464 ( .A(n49), .Y(n10134) );
  INVX0_HVT U9465 ( .A(n10178), .Y(n10177) );
  NAND2X0_HVT U9466 ( .A1(n47), .A2(n5645), .Y(n7719) );
  NAND2X0_HVT U9467 ( .A1(n7), .A2(n6258), .Y(n7720) );
  NAND2X0_HVT U9468 ( .A1(n37), .A2(n10376), .Y(n7721) );
  NAND2X0_HVT U9469 ( .A1(n44), .A2(n6258), .Y(n7722) );
  NAND2X0_HVT U9470 ( .A1(n12), .A2(n10375), .Y(n7723) );
  NAND2X0_HVT U9471 ( .A1(n16), .A2(n6258), .Y(n7724) );
  NAND2X0_HVT U9472 ( .A1(n24), .A2(n10376), .Y(n7725) );
  INVX0_HVT U9473 ( .A(n10178), .Y(n10176) );
  INVX0_HVT U9474 ( .A(n10202), .Y(n10200) );
  INVX0_HVT U9475 ( .A(n4604), .Y(n10175) );
  INVX0_HVT U9476 ( .A(n10252), .Y(n10251) );
  INVX0_HVT U9477 ( .A(n10367), .Y(n10373) );
  INVX0_HVT U9478 ( .A(n10202), .Y(n10201) );
  AO21X1_HVT U9479 ( .A1(n37), .A2(n5645), .A3(n10381), .Y(n7726) );
  AO21X1_HVT U9480 ( .A1(n47), .A2(n10375), .A3(rst), .Y(n7727) );
  AO21X1_HVT U9481 ( .A1(n44), .A2(n5645), .A3(n10381), .Y(n7728) );
  AO21X1_HVT U9482 ( .A1(n41), .A2(n10375), .A3(rst), .Y(n7731) );
  AO21X1_HVT U9483 ( .A1(n34), .A2(n10377), .A3(n10381), .Y(n7733) );
  INVX1_HVT U9484 ( .A(n9314), .Y(n9316) );
  INVX1_HVT U9485 ( .A(n9339), .Y(n9341) );
  INVX1_HVT U9486 ( .A(n9723), .Y(n9725) );
  INVX1_HVT U9487 ( .A(n9736), .Y(n9738) );
  INVX1_HVT U9488 ( .A(n9749), .Y(n9751) );
  INVX1_HVT U9489 ( .A(n9774), .Y(n9776) );
  INVX1_HVT U9490 ( .A(n9787), .Y(n9789) );
  INVX1_HVT U9491 ( .A(n9824), .Y(n9826) );
  INVX1_HVT U9492 ( .A(n9837), .Y(n9839) );
  INVX1_HVT U9493 ( .A(n9850), .Y(n9852) );
  INVX1_HVT U9494 ( .A(n9863), .Y(n9865) );
  INVX1_HVT U9495 ( .A(n9888), .Y(n9890) );
  INVX1_HVT U9496 ( .A(n9901), .Y(n9903) );
  INVX1_HVT U9497 ( .A(n9914), .Y(n9916) );
  INVX1_HVT U9498 ( .A(n9939), .Y(n9941) );
  INVX1_HVT U9499 ( .A(n9976), .Y(n9978) );
  INVX1_HVT U9500 ( .A(n10013), .Y(n10015) );
  INVX1_HVT U9501 ( .A(n10038), .Y(n10040) );
  INVX1_HVT U9502 ( .A(n10063), .Y(n10065) );
  INVX1_HVT U9503 ( .A(n10076), .Y(n10078) );
  INVX1_HVT U9504 ( .A(n10089), .Y(n10091) );
  INVX1_HVT U9505 ( .A(n10013), .Y(n10016) );
  INVX1_HVT U9506 ( .A(n10038), .Y(n10041) );
  INVX1_HVT U9507 ( .A(n9749), .Y(n9752) );
  INVX1_HVT U9508 ( .A(n9774), .Y(n9777) );
  INVX1_HVT U9509 ( .A(n9901), .Y(n9904) );
  INVX1_HVT U9510 ( .A(n9914), .Y(n9917) );
  INVX1_HVT U9511 ( .A(n9939), .Y(n9942) );
  INVX1_HVT U9512 ( .A(n9976), .Y(n9979) );
  INVX1_HVT U9513 ( .A(n10063), .Y(n10066) );
  INVX1_HVT U9514 ( .A(n10076), .Y(n10079) );
  INVX1_HVT U9515 ( .A(n9723), .Y(n9726) );
  INVX1_HVT U9516 ( .A(n9736), .Y(n9739) );
  INVX1_HVT U9517 ( .A(n9339), .Y(n9342) );
  INVX1_HVT U9518 ( .A(n9787), .Y(n9790) );
  INVX1_HVT U9519 ( .A(n9837), .Y(n9840) );
  INVX1_HVT U9520 ( .A(n9850), .Y(n9853) );
  INVX1_HVT U9521 ( .A(n9863), .Y(n9866) );
  INVX1_HVT U9522 ( .A(n9888), .Y(n9891) );
  INVX1_HVT U9523 ( .A(n10089), .Y(n10092) );
  MUX41X1_HVT U9524 ( .A1(\ram[12][0] ), .A3(\ram[14][0] ), .A2(\ram[13][0] ), 
        .A4(\ram[15][0] ), .S0(n5004), .S1(n8896), .Y(n7734) );
  MUX41X1_HVT U9525 ( .A1(\ram[8][0] ), .A3(\ram[10][0] ), .A2(\ram[9][0] ), 
        .A4(\ram[11][0] ), .S0(n4981), .S1(n8872), .Y(n7735) );
  MUX41X1_HVT U9526 ( .A1(\ram[0][0] ), .A3(\ram[2][0] ), .A2(\ram[1][0] ), 
        .A4(\ram[3][0] ), .S0(n8835), .S1(n8863), .Y(n7737) );
  MUX41X1_HVT U9527 ( .A1(n7737), .A3(n7735), .A2(n7736), .A4(n7734), .S0(
        n5799), .S1(n7547), .Y(q[0]) );
  MUX41X1_HVT U9528 ( .A1(\ram[8][1] ), .A3(\ram[10][1] ), .A2(\ram[9][1] ), 
        .A4(\ram[11][1] ), .S0(n5592), .S1(n8863), .Y(n7739) );
  MUX41X1_HVT U9529 ( .A1(\ram[4][1] ), .A3(\ram[6][1] ), .A2(\ram[5][1] ), 
        .A4(\ram[7][1] ), .S0(n5948), .S1(n5054), .Y(n7740) );
  MUX41X1_HVT U9530 ( .A1(\ram[0][1] ), .A3(\ram[2][1] ), .A2(\ram[1][1] ), 
        .A4(\ram[3][1] ), .S0(n6005), .S1(n5149), .Y(n7741) );
  MUX41X1_HVT U9531 ( .A1(\ram[12][2] ), .A3(\ram[14][2] ), .A2(\ram[13][2] ), 
        .A4(\ram[15][2] ), .S0(n5633), .S1(n7577), .Y(n7742) );
  MUX41X1_HVT U9532 ( .A1(\ram[8][2] ), .A3(\ram[10][2] ), .A2(\ram[9][2] ), 
        .A4(\ram[11][2] ), .S0(n5948), .S1(n5611), .Y(n7743) );
  MUX41X1_HVT U9533 ( .A1(\ram[4][2] ), .A3(\ram[6][2] ), .A2(\ram[5][2] ), 
        .A4(\ram[7][2] ), .S0(n5793), .S1(n5562), .Y(n7744) );
  MUX41X1_HVT U9534 ( .A1(\ram[0][2] ), .A3(\ram[2][2] ), .A2(\ram[1][2] ), 
        .A4(\ram[3][2] ), .S0(n8810), .S1(n8899), .Y(n7745) );
  MUX41X1_HVT U9535 ( .A1(n7745), .A3(n7743), .A2(n7744), .A4(n7742), .S0(
        n8764), .S1(n8772), .Y(q[2]) );
  MUX41X1_HVT U9536 ( .A1(\ram[12][3] ), .A3(\ram[14][3] ), .A2(\ram[13][3] ), 
        .A4(\ram[15][3] ), .S0(n7337), .S1(n5812), .Y(n7746) );
  MUX41X1_HVT U9537 ( .A1(\ram[8][3] ), .A3(\ram[10][3] ), .A2(\ram[9][3] ), 
        .A4(\ram[11][3] ), .S0(n7338), .S1(n5139), .Y(n7747) );
  MUX41X1_HVT U9538 ( .A1(\ram[4][4] ), .A3(\ram[6][4] ), .A2(\ram[5][4] ), 
        .A4(\ram[7][4] ), .S0(n6007), .S1(n7689), .Y(n7752) );
  MUX41X1_HVT U9539 ( .A1(\ram[0][4] ), .A3(\ram[2][4] ), .A2(\ram[1][4] ), 
        .A4(\ram[3][4] ), .S0(n8826), .S1(n5586), .Y(n7753) );
  MUX41X1_HVT U9540 ( .A1(\ram[12][5] ), .A3(\ram[14][5] ), .A2(\ram[13][5] ), 
        .A4(\ram[15][5] ), .S0(n6008), .S1(n5585), .Y(n7754) );
  MUX41X1_HVT U9541 ( .A1(\ram[8][5] ), .A3(\ram[10][5] ), .A2(\ram[9][5] ), 
        .A4(\ram[11][5] ), .S0(n5475), .S1(n7680), .Y(n7755) );
  MUX41X1_HVT U9542 ( .A1(\ram[0][5] ), .A3(\ram[2][5] ), .A2(\ram[1][5] ), 
        .A4(\ram[3][5] ), .S0(n7338), .S1(n5823), .Y(n7757) );
  MUX41X1_HVT U9543 ( .A1(\ram[4][6] ), .A3(\ram[6][6] ), .A2(\ram[5][6] ), 
        .A4(\ram[7][6] ), .S0(n6650), .S1(n8897), .Y(n7760) );
  MUX41X1_HVT U9544 ( .A1(\ram[0][6] ), .A3(\ram[2][6] ), .A2(\ram[1][6] ), 
        .A4(\ram[3][6] ), .S0(n5967), .S1(n8866), .Y(n7761) );
  MUX41X1_HVT U9545 ( .A1(\ram[8][7] ), .A3(\ram[10][7] ), .A2(\ram[9][7] ), 
        .A4(\ram[11][7] ), .S0(n8847), .S1(n8908), .Y(n7763) );
  MUX41X1_HVT U9546 ( .A1(\ram[4][7] ), .A3(\ram[6][7] ), .A2(\ram[5][7] ), 
        .A4(\ram[7][7] ), .S0(n8847), .S1(n8891), .Y(n7764) );
  MUX41X1_HVT U9547 ( .A1(\ram[12][8] ), .A3(\ram[14][8] ), .A2(\ram[13][8] ), 
        .A4(\ram[15][8] ), .S0(n8794), .S1(n5589), .Y(n7766) );
  MUX41X1_HVT U9548 ( .A1(\ram[4][8] ), .A3(\ram[6][8] ), .A2(\ram[5][8] ), 
        .A4(\ram[7][8] ), .S0(n6410), .S1(n8908), .Y(n7768) );
  MUX41X1_HVT U9549 ( .A1(\ram[8][9] ), .A3(\ram[10][9] ), .A2(\ram[9][9] ), 
        .A4(\ram[11][9] ), .S0(n4907), .S1(n8886), .Y(n7771) );
  MUX41X1_HVT U9550 ( .A1(\ram[4][9] ), .A3(\ram[6][9] ), .A2(\ram[5][9] ), 
        .A4(\ram[7][9] ), .S0(n5967), .S1(n5616), .Y(n7772) );
  MUX41X1_HVT U9551 ( .A1(\ram[8][10] ), .A3(\ram[10][10] ), .A2(\ram[9][10] ), 
        .A4(\ram[11][10] ), .S0(n7084), .S1(n5492), .Y(n7775) );
  MUX41X1_HVT U9552 ( .A1(\ram[12][11] ), .A3(\ram[14][11] ), .A2(
        \ram[13][11] ), .A4(\ram[15][11] ), .S0(n8798), .S1(n6762), .Y(n7778)
         );
  MUX41X1_HVT U9553 ( .A1(\ram[8][11] ), .A3(\ram[10][11] ), .A2(\ram[9][11] ), 
        .A4(\ram[11][11] ), .S0(n7312), .S1(n5964), .Y(n7779) );
  MUX41X1_HVT U9554 ( .A1(\ram[4][11] ), .A3(\ram[6][11] ), .A2(\ram[5][11] ), 
        .A4(\ram[7][11] ), .S0(n6410), .S1(n8869), .Y(n7780) );
  MUX41X1_HVT U9555 ( .A1(\ram[12][12] ), .A3(\ram[14][12] ), .A2(
        \ram[13][12] ), .A4(\ram[15][12] ), .S0(n4907), .S1(n6762), .Y(n7782)
         );
  MUX41X1_HVT U9556 ( .A1(\ram[4][12] ), .A3(\ram[6][12] ), .A2(\ram[5][12] ), 
        .A4(\ram[7][12] ), .S0(n4991), .S1(n5290), .Y(n7784) );
  MUX41X1_HVT U9557 ( .A1(\ram[12][13] ), .A3(\ram[14][13] ), .A2(
        \ram[13][13] ), .A4(\ram[15][13] ), .S0(n5946), .S1(n8902), .Y(n7786)
         );
  MUX41X1_HVT U9558 ( .A1(\ram[0][13] ), .A3(\ram[2][13] ), .A2(\ram[1][13] ), 
        .A4(\ram[3][13] ), .S0(n7312), .S1(n5758), .Y(n7789) );
  MUX41X1_HVT U9559 ( .A1(n7789), .A3(n7787), .A2(n7788), .A4(n7786), .S0(
        n6415), .S1(n8777), .Y(q[13]) );
  MUX41X1_HVT U9560 ( .A1(\ram[8][14] ), .A3(\ram[10][14] ), .A2(\ram[9][14] ), 
        .A4(\ram[11][14] ), .S0(n8847), .S1(n8896), .Y(n7791) );
  MUX41X1_HVT U9561 ( .A1(\ram[4][14] ), .A3(\ram[6][14] ), .A2(\ram[5][14] ), 
        .A4(\ram[7][14] ), .S0(n7312), .S1(n7707), .Y(n7792) );
  MUX41X1_HVT U9562 ( .A1(\ram[0][14] ), .A3(\ram[2][14] ), .A2(\ram[1][14] ), 
        .A4(\ram[3][14] ), .S0(n5733), .S1(n5851), .Y(n7793) );
  MUX41X1_HVT U9563 ( .A1(\ram[12][15] ), .A3(\ram[14][15] ), .A2(
        \ram[13][15] ), .A4(\ram[15][15] ), .S0(n7084), .S1(n7575), .Y(n7794)
         );
  MUX41X1_HVT U9564 ( .A1(\ram[4][15] ), .A3(\ram[6][15] ), .A2(\ram[5][15] ), 
        .A4(\ram[7][15] ), .S0(n8822), .S1(n5593), .Y(n7796) );
  MUX41X1_HVT U9565 ( .A1(\ram[8][16] ), .A3(\ram[10][16] ), .A2(\ram[9][16] ), 
        .A4(\ram[11][16] ), .S0(n8847), .S1(n7696), .Y(n7799) );
  MUX41X1_HVT U9566 ( .A1(\ram[4][16] ), .A3(\ram[6][16] ), .A2(\ram[5][16] ), 
        .A4(\ram[7][16] ), .S0(n5577), .S1(n8902), .Y(n7800) );
  MUX41X1_HVT U9567 ( .A1(\ram[12][17] ), .A3(\ram[14][17] ), .A2(
        \ram[13][17] ), .A4(\ram[15][17] ), .S0(n7312), .S1(n8862), .Y(n7802)
         );
  MUX41X1_HVT U9568 ( .A1(\ram[8][17] ), .A3(\ram[10][17] ), .A2(\ram[9][17] ), 
        .A4(\ram[11][17] ), .S0(n8848), .S1(n8902), .Y(n7803) );
  MUX41X1_HVT U9569 ( .A1(\ram[4][17] ), .A3(\ram[6][17] ), .A2(\ram[5][17] ), 
        .A4(\ram[7][17] ), .S0(n4991), .S1(n8901), .Y(n7804) );
  MUX41X1_HVT U9570 ( .A1(\ram[0][17] ), .A3(\ram[2][17] ), .A2(\ram[1][17] ), 
        .A4(\ram[3][17] ), .S0(n5945), .S1(n5528), .Y(n7805) );
  MUX41X1_HVT U9571 ( .A1(n7805), .A3(n7803), .A2(n7804), .A4(n7802), .S0(
        n5317), .S1(n7547), .Y(q[17]) );
  MUX41X1_HVT U9572 ( .A1(\ram[8][18] ), .A3(\ram[10][18] ), .A2(\ram[9][18] ), 
        .A4(\ram[11][18] ), .S0(n8822), .S1(n8899), .Y(n7807) );
  MUX41X1_HVT U9573 ( .A1(\ram[4][18] ), .A3(\ram[6][18] ), .A2(\ram[5][18] ), 
        .A4(\ram[7][18] ), .S0(n5945), .S1(n8879), .Y(n7808) );
  MUX41X1_HVT U9574 ( .A1(\ram[0][18] ), .A3(\ram[2][18] ), .A2(\ram[1][18] ), 
        .A4(\ram[3][18] ), .S0(n6650), .S1(n5621), .Y(n7809) );
  MUX41X1_HVT U9575 ( .A1(\ram[12][19] ), .A3(\ram[14][19] ), .A2(
        \ram[13][19] ), .A4(\ram[15][19] ), .S0(n5733), .S1(n4995), .Y(n7810)
         );
  MUX41X1_HVT U9576 ( .A1(\ram[8][19] ), .A3(\ram[10][19] ), .A2(\ram[9][19] ), 
        .A4(\ram[11][19] ), .S0(n7298), .S1(n5492), .Y(n7811) );
  MUX41X1_HVT U9577 ( .A1(\ram[0][19] ), .A3(\ram[2][19] ), .A2(\ram[1][19] ), 
        .A4(\ram[3][19] ), .S0(n7084), .S1(n4982), .Y(n7813) );
  MUX41X1_HVT U9578 ( .A1(\ram[12][20] ), .A3(\ram[14][20] ), .A2(
        \ram[13][20] ), .A4(\ram[15][20] ), .S0(n8848), .S1(n5601), .Y(n7814)
         );
  MUX41X1_HVT U9579 ( .A1(\ram[0][20] ), .A3(\ram[2][20] ), .A2(\ram[1][20] ), 
        .A4(\ram[3][20] ), .S0(n8848), .S1(n8859), .Y(n7815) );
  MUX41X1_HVT U9580 ( .A1(\ram[8][21] ), .A3(\ram[10][21] ), .A2(\ram[9][21] ), 
        .A4(\ram[11][21] ), .S0(n6020), .S1(n5939), .Y(n7817) );
  MUX41X1_HVT U9581 ( .A1(\ram[4][21] ), .A3(\ram[6][21] ), .A2(\ram[5][21] ), 
        .A4(\ram[7][21] ), .S0(n5523), .S1(n7713), .Y(n7818) );
  MUX41X1_HVT U9582 ( .A1(\ram[0][21] ), .A3(\ram[2][21] ), .A2(\ram[1][21] ), 
        .A4(\ram[3][21] ), .S0(n8822), .S1(n7713), .Y(n7819) );
  MUX41X1_HVT U9583 ( .A1(n7819), .A3(n7817), .A2(n7818), .A4(n7816), .S0(
        n8762), .S1(n8778), .Y(q[21]) );
  MUX41X1_HVT U9584 ( .A1(\ram[4][22] ), .A3(\ram[6][22] ), .A2(\ram[5][22] ), 
        .A4(\ram[7][22] ), .S0(n5734), .S1(n7713), .Y(n7822) );
  MUX41X1_HVT U9585 ( .A1(\ram[0][22] ), .A3(\ram[2][22] ), .A2(\ram[1][22] ), 
        .A4(\ram[3][22] ), .S0(n5577), .S1(n7713), .Y(n7823) );
  MUX41X1_HVT U9586 ( .A1(\ram[12][23] ), .A3(\ram[14][23] ), .A2(
        \ram[13][23] ), .A4(\ram[15][23] ), .S0(n8794), .S1(n4873), .Y(n7824)
         );
  MUX41X1_HVT U9587 ( .A1(\ram[8][23] ), .A3(\ram[10][23] ), .A2(\ram[9][23] ), 
        .A4(\ram[11][23] ), .S0(n7084), .S1(n5123), .Y(n7825) );
  MUX41X1_HVT U9588 ( .A1(\ram[4][23] ), .A3(\ram[6][23] ), .A2(\ram[5][23] ), 
        .A4(\ram[7][23] ), .S0(n6410), .S1(n5650), .Y(n7826) );
  MUX41X1_HVT U9589 ( .A1(\ram[12][24] ), .A3(\ram[14][24] ), .A2(
        \ram[13][24] ), .A4(\ram[15][24] ), .S0(n5504), .S1(n5470), .Y(n7828)
         );
  MUX41X1_HVT U9590 ( .A1(\ram[8][24] ), .A3(\ram[10][24] ), .A2(\ram[9][24] ), 
        .A4(\ram[11][24] ), .S0(n6757), .S1(n5586), .Y(n7829) );
  MUX41X1_HVT U9591 ( .A1(\ram[4][24] ), .A3(\ram[6][24] ), .A2(\ram[5][24] ), 
        .A4(\ram[7][24] ), .S0(n4883), .S1(n8872), .Y(n7830) );
  MUX41X1_HVT U9592 ( .A1(\ram[0][24] ), .A3(\ram[2][24] ), .A2(\ram[1][24] ), 
        .A4(\ram[3][24] ), .S0(n8819), .S1(n7706), .Y(n7831) );
  MUX41X1_HVT U9593 ( .A1(n7831), .A3(n7829), .A2(n7830), .A4(n7828), .S0(
        n8762), .S1(n8772), .Y(q[24]) );
  MUX41X1_HVT U9594 ( .A1(\ram[12][25] ), .A3(\ram[14][25] ), .A2(
        \ram[13][25] ), .A4(\ram[15][25] ), .S0(n8814), .S1(n5580), .Y(n7832)
         );
  MUX41X1_HVT U9595 ( .A1(\ram[4][25] ), .A3(\ram[6][25] ), .A2(\ram[5][25] ), 
        .A4(\ram[7][25] ), .S0(n6024), .S1(n7706), .Y(n7834) );
  MUX41X1_HVT U9596 ( .A1(\ram[0][25] ), .A3(\ram[2][25] ), .A2(\ram[1][25] ), 
        .A4(\ram[3][25] ), .S0(n8815), .S1(n8868), .Y(n7835) );
  MUX41X1_HVT U9597 ( .A1(n7835), .A3(n7833), .A2(n7834), .A4(n7832), .S0(
        n7543), .S1(n8771), .Y(q[25]) );
  MUX41X1_HVT U9598 ( .A1(\ram[8][26] ), .A3(\ram[10][26] ), .A2(\ram[9][26] ), 
        .A4(\ram[11][26] ), .S0(n5076), .S1(n7707), .Y(n7837) );
  MUX41X1_HVT U9599 ( .A1(\ram[4][26] ), .A3(\ram[6][26] ), .A2(\ram[5][26] ), 
        .A4(\ram[7][26] ), .S0(n7141), .S1(n8863), .Y(n7838) );
  MUX41X1_HVT U9600 ( .A1(\ram[0][26] ), .A3(\ram[2][26] ), .A2(\ram[1][26] ), 
        .A4(\ram[3][26] ), .S0(n8811), .S1(n4819), .Y(n7839) );
  MUX41X1_HVT U9601 ( .A1(\ram[8][27] ), .A3(\ram[10][27] ), .A2(\ram[9][27] ), 
        .A4(\ram[11][27] ), .S0(n8840), .S1(n8907), .Y(n7841) );
  MUX41X1_HVT U9602 ( .A1(\ram[4][27] ), .A3(\ram[6][27] ), .A2(\ram[5][27] ), 
        .A4(\ram[7][27] ), .S0(n4918), .S1(n4182), .Y(n7842) );
  MUX41X1_HVT U9603 ( .A1(\ram[0][27] ), .A3(\ram[2][27] ), .A2(\ram[1][27] ), 
        .A4(\ram[3][27] ), .S0(n4794), .S1(n5962), .Y(n7843) );
  MUX41X1_HVT U9604 ( .A1(n7843), .A3(n7841), .A2(n7842), .A4(n7840), .S0(
        n5925), .S1(n5536), .Y(q[27]) );
  MUX41X1_HVT U9605 ( .A1(\ram[12][28] ), .A3(\ram[14][28] ), .A2(
        \ram[13][28] ), .A4(\ram[15][28] ), .S0(n4794), .S1(n5290), .Y(n7844)
         );
  MUX41X1_HVT U9606 ( .A1(\ram[8][28] ), .A3(\ram[10][28] ), .A2(\ram[9][28] ), 
        .A4(\ram[11][28] ), .S0(n5859), .S1(n5006), .Y(n7845) );
  MUX41X1_HVT U9607 ( .A1(\ram[4][28] ), .A3(\ram[6][28] ), .A2(\ram[5][28] ), 
        .A4(\ram[7][28] ), .S0(n4939), .S1(n6748), .Y(n7846) );
  MUX41X1_HVT U9608 ( .A1(\ram[0][28] ), .A3(\ram[2][28] ), .A2(\ram[1][28] ), 
        .A4(\ram[3][28] ), .S0(n5854), .S1(n5491), .Y(n7847) );
  MUX41X1_HVT U9609 ( .A1(n7847), .A3(n7845), .A2(n7846), .A4(n7844), .S0(
        n7543), .S1(n5931), .Y(q[28]) );
  MUX41X1_HVT U9610 ( .A1(\ram[12][29] ), .A3(\ram[14][29] ), .A2(
        \ram[13][29] ), .A4(\ram[15][29] ), .S0(n8804), .S1(n7689), .Y(n7848)
         );
  MUX41X1_HVT U9611 ( .A1(\ram[8][29] ), .A3(\ram[10][29] ), .A2(\ram[9][29] ), 
        .A4(\ram[11][29] ), .S0(n5334), .S1(n8858), .Y(n7849) );
  MUX41X1_HVT U9612 ( .A1(\ram[4][29] ), .A3(\ram[6][29] ), .A2(\ram[5][29] ), 
        .A4(\ram[7][29] ), .S0(n8840), .S1(n4873), .Y(n7850) );
  MUX41X1_HVT U9613 ( .A1(\ram[0][29] ), .A3(\ram[2][29] ), .A2(\ram[1][29] ), 
        .A4(\ram[3][29] ), .S0(n7312), .S1(n6014), .Y(n7851) );
  MUX41X1_HVT U9614 ( .A1(n7851), .A3(n7849), .A2(n7850), .A4(n7848), .S0(
        n8762), .S1(n7351), .Y(q[29]) );
  MUX41X1_HVT U9615 ( .A1(\ram[8][30] ), .A3(\ram[10][30] ), .A2(\ram[9][30] ), 
        .A4(\ram[11][30] ), .S0(n8828), .S1(n5444), .Y(n7852) );
  MUX41X1_HVT U9616 ( .A1(\ram[4][30] ), .A3(\ram[6][30] ), .A2(\ram[5][30] ), 
        .A4(\ram[7][30] ), .S0(n4949), .S1(n5585), .Y(n7853) );
  MUX41X1_HVT U9617 ( .A1(\ram[0][30] ), .A3(\ram[2][30] ), .A2(\ram[1][30] ), 
        .A4(\ram[3][30] ), .S0(n7145), .S1(n5621), .Y(n7854) );
  MUX41X1_HVT U9618 ( .A1(\ram[12][31] ), .A3(\ram[14][31] ), .A2(
        \ram[13][31] ), .A4(\ram[15][31] ), .S0(n8814), .S1(n8878), .Y(n7855)
         );
  MUX41X1_HVT U9619 ( .A1(\ram[4][31] ), .A3(\ram[6][31] ), .A2(\ram[5][31] ), 
        .A4(\ram[7][31] ), .S0(n4837), .S1(n8889), .Y(n7857) );
  MUX41X1_HVT U9620 ( .A1(\ram[0][31] ), .A3(\ram[2][31] ), .A2(\ram[1][31] ), 
        .A4(\ram[3][31] ), .S0(n8831), .S1(n4772), .Y(n7858) );
  MUX41X1_HVT U9621 ( .A1(\ram[12][32] ), .A3(\ram[14][32] ), .A2(
        \ram[13][32] ), .A4(\ram[15][32] ), .S0(n7552), .S1(n6006), .Y(n7859)
         );
  MUX41X1_HVT U9622 ( .A1(\ram[4][32] ), .A3(\ram[6][32] ), .A2(\ram[5][32] ), 
        .A4(\ram[7][32] ), .S0(n8846), .S1(n5144), .Y(n7861) );
  MUX41X1_HVT U9623 ( .A1(\ram[0][32] ), .A3(\ram[2][32] ), .A2(\ram[1][32] ), 
        .A4(\ram[3][32] ), .S0(n5310), .S1(n7680), .Y(n7862) );
  MUX41X1_HVT U9624 ( .A1(\ram[12][33] ), .A3(\ram[14][33] ), .A2(
        \ram[13][33] ), .A4(\ram[15][33] ), .S0(n5892), .S1(n8901), .Y(n7863)
         );
  MUX41X1_HVT U9625 ( .A1(\ram[4][33] ), .A3(\ram[6][33] ), .A2(\ram[5][33] ), 
        .A4(\ram[7][33] ), .S0(n6024), .S1(n5642), .Y(n7865) );
  MUX41X1_HVT U9626 ( .A1(\ram[0][33] ), .A3(\ram[2][33] ), .A2(\ram[1][33] ), 
        .A4(\ram[3][33] ), .S0(n6024), .S1(n5609), .Y(n7866) );
  MUX41X1_HVT U9627 ( .A1(n7866), .A3(n7864), .A2(n7865), .A4(n7863), .S0(
        n8762), .S1(n8776), .Y(q[33]) );
  MUX41X1_HVT U9628 ( .A1(\ram[8][34] ), .A3(\ram[10][34] ), .A2(\ram[9][34] ), 
        .A4(\ram[11][34] ), .S0(n5504), .S1(n5560), .Y(n7868) );
  MUX41X1_HVT U9629 ( .A1(\ram[4][34] ), .A3(\ram[6][34] ), .A2(\ram[5][34] ), 
        .A4(\ram[7][34] ), .S0(n5888), .S1(n8878), .Y(n7869) );
  MUX41X1_HVT U9630 ( .A1(\ram[0][34] ), .A3(\ram[2][34] ), .A2(\ram[1][34] ), 
        .A4(\ram[3][34] ), .S0(n5569), .S1(n7327), .Y(n7870) );
  MUX41X1_HVT U9631 ( .A1(n7870), .A3(n7868), .A2(n7869), .A4(n7867), .S0(
        n5925), .S1(n5362), .Y(q[34]) );
  MUX41X1_HVT U9632 ( .A1(\ram[12][35] ), .A3(\ram[14][35] ), .A2(
        \ram[13][35] ), .A4(\ram[15][35] ), .S0(n7321), .S1(n6010), .Y(n7871)
         );
  MUX41X1_HVT U9633 ( .A1(\ram[4][35] ), .A3(\ram[6][35] ), .A2(\ram[5][35] ), 
        .A4(\ram[7][35] ), .S0(n7330), .S1(n7694), .Y(n7873) );
  MUX41X1_HVT U9634 ( .A1(\ram[0][35] ), .A3(\ram[2][35] ), .A2(\ram[1][35] ), 
        .A4(\ram[3][35] ), .S0(n7330), .S1(n5535), .Y(n7874) );
  MUX41X1_HVT U9635 ( .A1(n7874), .A3(n7872), .A2(n7873), .A4(n7871), .S0(
        n7543), .S1(n5112), .Y(q[35]) );
  MUX41X1_HVT U9636 ( .A1(\ram[8][36] ), .A3(\ram[10][36] ), .A2(\ram[9][36] ), 
        .A4(\ram[11][36] ), .S0(n5994), .S1(n7669), .Y(n7876) );
  MUX41X1_HVT U9637 ( .A1(\ram[4][36] ), .A3(\ram[6][36] ), .A2(\ram[5][36] ), 
        .A4(\ram[7][36] ), .S0(n8836), .S1(n8899), .Y(n7877) );
  MUX41X1_HVT U9638 ( .A1(\ram[0][36] ), .A3(\ram[2][36] ), .A2(\ram[1][36] ), 
        .A4(\ram[3][36] ), .S0(n8836), .S1(n8886), .Y(n7878) );
  MUX41X1_HVT U9639 ( .A1(\ram[8][37] ), .A3(\ram[10][37] ), .A2(\ram[9][37] ), 
        .A4(\ram[11][37] ), .S0(n8825), .S1(n7327), .Y(n7880) );
  MUX41X1_HVT U9640 ( .A1(\ram[0][37] ), .A3(\ram[2][37] ), .A2(\ram[1][37] ), 
        .A4(\ram[3][37] ), .S0(n6029), .S1(n6744), .Y(n7882) );
  MUX41X1_HVT U9641 ( .A1(\ram[4][38] ), .A3(\ram[6][38] ), .A2(\ram[5][38] ), 
        .A4(\ram[7][38] ), .S0(n8827), .S1(n5650), .Y(n7885) );
  MUX41X1_HVT U9642 ( .A1(\ram[0][38] ), .A3(\ram[2][38] ), .A2(\ram[1][38] ), 
        .A4(\ram[3][38] ), .S0(n6028), .S1(n8899), .Y(n7886) );
  MUX41X1_HVT U9643 ( .A1(\ram[8][39] ), .A3(\ram[10][39] ), .A2(\ram[9][39] ), 
        .A4(\ram[11][39] ), .S0(n5750), .S1(n5869), .Y(n7888) );
  MUX41X1_HVT U9644 ( .A1(\ram[4][39] ), .A3(\ram[6][39] ), .A2(\ram[5][39] ), 
        .A4(\ram[7][39] ), .S0(n5997), .S1(n8894), .Y(n7889) );
  MUX41X1_HVT U9645 ( .A1(\ram[0][39] ), .A3(\ram[2][39] ), .A2(\ram[1][39] ), 
        .A4(\ram[3][39] ), .S0(n7551), .S1(n7579), .Y(n7890) );
  MUX41X1_HVT U9646 ( .A1(n7890), .A3(n7888), .A2(n7889), .A4(n7887), .S0(
        n7543), .S1(n8777), .Y(q[39]) );
  MUX41X1_HVT U9647 ( .A1(\ram[12][40] ), .A3(\ram[14][40] ), .A2(
        \ram[13][40] ), .A4(\ram[15][40] ), .S0(n6029), .S1(n6747), .Y(n7891)
         );
  MUX41X1_HVT U9648 ( .A1(\ram[8][41] ), .A3(\ram[10][41] ), .A2(\ram[9][41] ), 
        .A4(\ram[11][41] ), .S0(n8827), .S1(n8894), .Y(n7896) );
  MUX41X1_HVT U9649 ( .A1(\ram[12][42] ), .A3(\ram[14][42] ), .A2(
        \ram[13][42] ), .A4(\ram[15][42] ), .S0(n6183), .S1(n8873), .Y(n7899)
         );
  MUX41X1_HVT U9650 ( .A1(\ram[8][42] ), .A3(\ram[10][42] ), .A2(\ram[9][42] ), 
        .A4(\ram[11][42] ), .S0(n5238), .S1(n4176), .Y(n7900) );
  MUX41X1_HVT U9651 ( .A1(\ram[4][42] ), .A3(\ram[6][42] ), .A2(\ram[5][42] ), 
        .A4(\ram[7][42] ), .S0(n8824), .S1(n8897), .Y(n7901) );
  MUX41X1_HVT U9652 ( .A1(\ram[0][42] ), .A3(\ram[2][42] ), .A2(\ram[1][42] ), 
        .A4(\ram[3][42] ), .S0(n8817), .S1(n8866), .Y(n7902) );
  MUX41X1_HVT U9653 ( .A1(\ram[8][43] ), .A3(\ram[10][43] ), .A2(\ram[9][43] ), 
        .A4(\ram[11][43] ), .S0(n7321), .S1(n7679), .Y(n7904) );
  MUX41X1_HVT U9654 ( .A1(\ram[4][43] ), .A3(\ram[6][43] ), .A2(\ram[5][43] ), 
        .A4(\ram[7][43] ), .S0(n7325), .S1(n5989), .Y(n7905) );
  MUX41X1_HVT U9655 ( .A1(\ram[12][44] ), .A3(\ram[14][44] ), .A2(
        \ram[13][44] ), .A4(\ram[15][44] ), .S0(n8797), .S1(n1651), .Y(n7907)
         );
  MUX41X1_HVT U9656 ( .A1(\ram[8][44] ), .A3(\ram[10][44] ), .A2(\ram[9][44] ), 
        .A4(\ram[11][44] ), .S0(n6031), .S1(n5313), .Y(n7908) );
  MUX41X1_HVT U9657 ( .A1(\ram[4][44] ), .A3(\ram[6][44] ), .A2(\ram[5][44] ), 
        .A4(\ram[7][44] ), .S0(n4973), .S1(n6394), .Y(n7909) );
  MUX41X1_HVT U9658 ( .A1(\ram[0][44] ), .A3(\ram[2][44] ), .A2(\ram[1][44] ), 
        .A4(\ram[3][44] ), .S0(n7338), .S1(n5316), .Y(n7910) );
  MUX41X1_HVT U9659 ( .A1(\ram[8][45] ), .A3(\ram[10][45] ), .A2(\ram[9][45] ), 
        .A4(\ram[11][45] ), .S0(n8803), .S1(n5812), .Y(n7912) );
  MUX41X1_HVT U9660 ( .A1(\ram[4][45] ), .A3(\ram[6][45] ), .A2(\ram[5][45] ), 
        .A4(\ram[7][45] ), .S0(n5751), .S1(n5807), .Y(n7913) );
  MUX41X1_HVT U9661 ( .A1(\ram[0][45] ), .A3(\ram[2][45] ), .A2(\ram[1][45] ), 
        .A4(\ram[3][45] ), .S0(n8803), .S1(n5795), .Y(n7914) );
  MUX41X1_HVT U9662 ( .A1(\ram[8][46] ), .A3(\ram[10][46] ), .A2(\ram[9][46] ), 
        .A4(\ram[11][46] ), .S0(n8798), .S1(n5614), .Y(n7916) );
  MUX41X1_HVT U9663 ( .A1(\ram[4][46] ), .A3(\ram[6][46] ), .A2(\ram[5][46] ), 
        .A4(\ram[7][46] ), .S0(n5854), .S1(n7687), .Y(n7917) );
  MUX41X1_HVT U9664 ( .A1(\ram[0][46] ), .A3(\ram[2][46] ), .A2(\ram[1][46] ), 
        .A4(\ram[3][46] ), .S0(n8796), .S1(n5591), .Y(n7918) );
  MUX41X1_HVT U9665 ( .A1(n7918), .A3(n7916), .A2(n7917), .A4(n7915), .S0(
        n5321), .S1(n7309), .Y(q[46]) );
  MUX41X1_HVT U9666 ( .A1(\ram[12][47] ), .A3(\ram[14][47] ), .A2(
        \ram[13][47] ), .A4(\ram[15][47] ), .S0(n6652), .S1(n5226), .Y(n7919)
         );
  MUX41X1_HVT U9667 ( .A1(\ram[8][47] ), .A3(\ram[10][47] ), .A2(\ram[9][47] ), 
        .A4(\ram[11][47] ), .S0(n8796), .S1(n8870), .Y(n7920) );
  MUX41X1_HVT U9668 ( .A1(\ram[4][47] ), .A3(\ram[6][47] ), .A2(\ram[5][47] ), 
        .A4(\ram[7][47] ), .S0(n5900), .S1(n8854), .Y(n7921) );
  MUX41X1_HVT U9669 ( .A1(\ram[0][47] ), .A3(\ram[2][47] ), .A2(\ram[1][47] ), 
        .A4(\ram[3][47] ), .S0(n4990), .S1(n8889), .Y(n7922) );
  MUX41X1_HVT U9670 ( .A1(n7922), .A3(n7920), .A2(n7921), .A4(n7919), .S0(
        n8764), .S1(n7666), .Y(q[47]) );
  MUX41X1_HVT U9671 ( .A1(\ram[4][48] ), .A3(\ram[6][48] ), .A2(\ram[5][48] ), 
        .A4(\ram[7][48] ), .S0(n6018), .S1(n5123), .Y(n7925) );
  MUX41X1_HVT U9672 ( .A1(\ram[8][49] ), .A3(\ram[10][49] ), .A2(\ram[9][49] ), 
        .A4(\ram[11][49] ), .S0(n5946), .S1(n5777), .Y(n7928) );
  MUX41X1_HVT U9673 ( .A1(\ram[4][49] ), .A3(\ram[6][49] ), .A2(\ram[5][49] ), 
        .A4(\ram[7][49] ), .S0(n7084), .S1(n8891), .Y(n7929) );
  MUX41X1_HVT U9674 ( .A1(\ram[0][49] ), .A3(\ram[2][49] ), .A2(\ram[1][49] ), 
        .A4(\ram[3][49] ), .S0(n7550), .S1(n8878), .Y(n7930) );
  MUX41X1_HVT U9675 ( .A1(\ram[8][50] ), .A3(\ram[10][50] ), .A2(\ram[9][50] ), 
        .A4(\ram[11][50] ), .S0(n6031), .S1(n6744), .Y(n7932) );
  MUX41X1_HVT U9676 ( .A1(\ram[4][50] ), .A3(\ram[6][50] ), .A2(\ram[5][50] ), 
        .A4(\ram[7][50] ), .S0(n6642), .S1(n8878), .Y(n7933) );
  MUX41X1_HVT U9677 ( .A1(\ram[0][50] ), .A3(\ram[2][50] ), .A2(\ram[1][50] ), 
        .A4(\ram[3][50] ), .S0(n4907), .S1(n4860), .Y(n7934) );
  MUX41X1_HVT U9678 ( .A1(\ram[12][51] ), .A3(\ram[14][51] ), .A2(
        \ram[13][51] ), .A4(\ram[15][51] ), .S0(n8802), .S1(n5441), .Y(n7935)
         );
  MUX41X1_HVT U9679 ( .A1(\ram[8][51] ), .A3(\ram[10][51] ), .A2(\ram[9][51] ), 
        .A4(\ram[11][51] ), .S0(n7549), .S1(n7560), .Y(n7936) );
  MUX41X1_HVT U9680 ( .A1(\ram[4][51] ), .A3(\ram[6][51] ), .A2(\ram[5][51] ), 
        .A4(\ram[7][51] ), .S0(n8794), .S1(n5470), .Y(n7937) );
  MUX41X1_HVT U9681 ( .A1(\ram[0][51] ), .A3(\ram[2][51] ), .A2(\ram[1][51] ), 
        .A4(\ram[3][51] ), .S0(n7549), .S1(n4983), .Y(n7938) );
  MUX41X1_HVT U9682 ( .A1(n7938), .A3(n7936), .A2(n7937), .A4(n7935), .S0(
        n7293), .S1(n5237), .Y(q[51]) );
  MUX41X1_HVT U9683 ( .A1(\ram[12][52] ), .A3(\ram[14][52] ), .A2(
        \ram[13][52] ), .A4(\ram[15][52] ), .S0(n8842), .S1(n8862), .Y(n7939)
         );
  MUX41X1_HVT U9684 ( .A1(\ram[8][52] ), .A3(\ram[10][52] ), .A2(\ram[9][52] ), 
        .A4(\ram[11][52] ), .S0(n4907), .S1(n5580), .Y(n7940) );
  MUX41X1_HVT U9685 ( .A1(n7942), .A3(n7940), .A2(n7941), .A4(n7939), .S0(
        n8761), .S1(n5926), .Y(q[52]) );
  MUX41X1_HVT U9686 ( .A1(\ram[12][53] ), .A3(\ram[14][53] ), .A2(
        \ram[13][53] ), .A4(\ram[15][53] ), .S0(n7141), .S1(n5593), .Y(n7943)
         );
  MUX41X1_HVT U9687 ( .A1(\ram[8][53] ), .A3(\ram[10][53] ), .A2(\ram[9][53] ), 
        .A4(\ram[11][53] ), .S0(n7549), .S1(n5528), .Y(n7944) );
  MUX41X1_HVT U9688 ( .A1(\ram[4][53] ), .A3(\ram[6][53] ), .A2(\ram[5][53] ), 
        .A4(\ram[7][53] ), .S0(n7141), .S1(n7560), .Y(n7945) );
  MUX41X1_HVT U9689 ( .A1(\ram[0][53] ), .A3(\ram[2][53] ), .A2(\ram[1][53] ), 
        .A4(\ram[3][53] ), .S0(n6757), .S1(n5869), .Y(n7946) );
  MUX41X1_HVT U9690 ( .A1(\ram[8][55] ), .A3(\ram[10][55] ), .A2(\ram[9][55] ), 
        .A4(\ram[11][55] ), .S0(n8793), .S1(n8854), .Y(n7952) );
  MUX41X1_HVT U9691 ( .A1(\ram[4][55] ), .A3(\ram[6][55] ), .A2(\ram[5][55] ), 
        .A4(\ram[7][55] ), .S0(n5940), .S1(n8859), .Y(n7953) );
  MUX41X1_HVT U9692 ( .A1(\ram[0][55] ), .A3(\ram[2][55] ), .A2(\ram[1][55] ), 
        .A4(\ram[3][55] ), .S0(n5050), .S1(n5614), .Y(n7954) );
  MUX41X1_HVT U9693 ( .A1(n7954), .A3(n7952), .A2(n7953), .A4(n7951), .S0(
        n8759), .S1(n5536), .Y(q[55]) );
  MUX41X1_HVT U9694 ( .A1(\ram[8][56] ), .A3(\ram[10][56] ), .A2(\ram[9][56] ), 
        .A4(\ram[11][56] ), .S0(n5793), .S1(n5570), .Y(n7956) );
  MUX41X1_HVT U9695 ( .A1(\ram[4][56] ), .A3(\ram[6][56] ), .A2(\ram[5][56] ), 
        .A4(\ram[7][56] ), .S0(n8810), .S1(n7559), .Y(n7957) );
  MUX41X1_HVT U9696 ( .A1(\ram[0][56] ), .A3(\ram[2][56] ), .A2(\ram[1][56] ), 
        .A4(\ram[3][56] ), .S0(n8838), .S1(n5570), .Y(n7958) );
  MUX41X1_HVT U9697 ( .A1(n7958), .A3(n7956), .A2(n7957), .A4(n7955), .S0(
        n8759), .S1(n8776), .Y(q[56]) );
  MUX41X1_HVT U9698 ( .A1(\ram[4][57] ), .A3(\ram[6][57] ), .A2(\ram[5][57] ), 
        .A4(\ram[7][57] ), .S0(n6029), .S1(n5584), .Y(n7961) );
  MUX41X1_HVT U9699 ( .A1(\ram[0][57] ), .A3(\ram[2][57] ), .A2(\ram[1][57] ), 
        .A4(\ram[3][57] ), .S0(n8836), .S1(n5476), .Y(n7962) );
  MUX41X1_HVT U9700 ( .A1(\ram[4][58] ), .A3(\ram[6][58] ), .A2(\ram[5][58] ), 
        .A4(\ram[7][58] ), .S0(n6028), .S1(n8894), .Y(n7964) );
  MUX41X1_HVT U9701 ( .A1(\ram[0][58] ), .A3(\ram[2][58] ), .A2(\ram[1][58] ), 
        .A4(\ram[3][58] ), .S0(n6031), .S1(n8887), .Y(n7965) );
  MUX41X1_HVT U9702 ( .A1(\ram[0][59] ), .A3(\ram[2][59] ), .A2(\ram[1][59] ), 
        .A4(\ram[3][59] ), .S0(n6029), .S1(n5210), .Y(n7969) );
  MUX41X1_HVT U9703 ( .A1(\ram[12][60] ), .A3(\ram[14][60] ), .A2(
        \ram[13][60] ), .A4(\ram[15][60] ), .S0(n8847), .S1(n5950), .Y(n7970)
         );
  MUX41X1_HVT U9704 ( .A1(\ram[8][60] ), .A3(\ram[10][60] ), .A2(\ram[9][60] ), 
        .A4(\ram[11][60] ), .S0(n5892), .S1(n8873), .Y(n7971) );
  MUX41X1_HVT U9705 ( .A1(\ram[4][60] ), .A3(\ram[6][60] ), .A2(\ram[5][60] ), 
        .A4(\ram[7][60] ), .S0(n5504), .S1(n5889), .Y(n7972) );
  MUX41X1_HVT U9706 ( .A1(\ram[0][60] ), .A3(\ram[2][60] ), .A2(\ram[1][60] ), 
        .A4(\ram[3][60] ), .S0(n5322), .S1(n6762), .Y(n7973) );
  MUX41X1_HVT U9707 ( .A1(n7973), .A3(n7971), .A2(n7972), .A4(n7970), .S0(
        n8761), .S1(n7332), .Y(q[60]) );
  MUX41X1_HVT U9708 ( .A1(\ram[12][61] ), .A3(\ram[14][61] ), .A2(
        \ram[13][61] ), .A4(\ram[15][61] ), .S0(n4884), .S1(n5614), .Y(n7974)
         );
  MUX41X1_HVT U9709 ( .A1(\ram[4][61] ), .A3(\ram[6][61] ), .A2(\ram[5][61] ), 
        .A4(\ram[7][61] ), .S0(n8815), .S1(n6744), .Y(n7976) );
  MUX41X1_HVT U9710 ( .A1(\ram[0][61] ), .A3(\ram[2][61] ), .A2(\ram[1][61] ), 
        .A4(\ram[3][61] ), .S0(n8828), .S1(n6034), .Y(n7977) );
  MUX41X1_HVT U9711 ( .A1(n7977), .A3(n7975), .A2(n7976), .A4(n7974), .S0(
        n8759), .S1(n5136), .Y(q[61]) );
  MUX41X1_HVT U9712 ( .A1(\ram[12][62] ), .A3(\ram[14][62] ), .A2(
        \ram[13][62] ), .A4(\ram[15][62] ), .S0(n5000), .S1(n1389), .Y(n7978)
         );
  MUX41X1_HVT U9713 ( .A1(\ram[8][62] ), .A3(\ram[10][62] ), .A2(\ram[9][62] ), 
        .A4(\ram[11][62] ), .S0(n8815), .S1(n5601), .Y(n7979) );
  MUX41X1_HVT U9714 ( .A1(\ram[4][62] ), .A3(\ram[6][62] ), .A2(\ram[5][62] ), 
        .A4(\ram[7][62] ), .S0(n5000), .S1(n5582), .Y(n7980) );
  MUX41X1_HVT U9715 ( .A1(\ram[0][62] ), .A3(\ram[2][62] ), .A2(\ram[1][62] ), 
        .A4(\ram[3][62] ), .S0(n7324), .S1(n5758), .Y(n7981) );
  MUX41X1_HVT U9716 ( .A1(n7981), .A3(n7979), .A2(n7980), .A4(n7978), .S0(
        n5289), .S1(n8771), .Y(q[62]) );
  MUX41X1_HVT U9717 ( .A1(\ram[12][63] ), .A3(\ram[14][63] ), .A2(
        \ram[13][63] ), .A4(\ram[15][63] ), .S0(n5994), .S1(n8875), .Y(n7982)
         );
  MUX41X1_HVT U9718 ( .A1(\ram[4][63] ), .A3(\ram[6][63] ), .A2(\ram[5][63] ), 
        .A4(\ram[7][63] ), .S0(n5050), .S1(n6394), .Y(n7984) );
  MUX41X1_HVT U9719 ( .A1(\ram[0][63] ), .A3(\ram[2][63] ), .A2(\ram[1][63] ), 
        .A4(\ram[3][63] ), .S0(n6652), .S1(n6407), .Y(n7985) );
  MUX41X1_HVT U9720 ( .A1(\ram[8][64] ), .A3(\ram[10][64] ), .A2(\ram[9][64] ), 
        .A4(\ram[11][64] ), .S0(n8829), .S1(n5458), .Y(n7987) );
  MUX41X1_HVT U9721 ( .A1(\ram[4][64] ), .A3(\ram[6][64] ), .A2(\ram[5][64] ), 
        .A4(\ram[7][64] ), .S0(n7321), .S1(n8875), .Y(n7988) );
  MUX41X1_HVT U9722 ( .A1(\ram[0][64] ), .A3(\ram[2][64] ), .A2(\ram[1][64] ), 
        .A4(\ram[3][64] ), .S0(n8798), .S1(n6407), .Y(n7989) );
  MUX41X1_HVT U9723 ( .A1(n7989), .A3(n7987), .A2(n7988), .A4(n7986), .S0(
        n5110), .S1(n8766), .Y(q[64]) );
  MUX41X1_HVT U9724 ( .A1(\ram[8][65] ), .A3(\ram[10][65] ), .A2(\ram[9][65] ), 
        .A4(\ram[11][65] ), .S0(n5865), .S1(n5591), .Y(n7991) );
  MUX41X1_HVT U9725 ( .A1(\ram[4][65] ), .A3(\ram[6][65] ), .A2(\ram[5][65] ), 
        .A4(\ram[7][65] ), .S0(n5558), .S1(n7683), .Y(n7992) );
  MUX41X1_HVT U9726 ( .A1(\ram[0][65] ), .A3(\ram[2][65] ), .A2(\ram[1][65] ), 
        .A4(\ram[3][65] ), .S0(n5900), .S1(n7687), .Y(n7993) );
  MUX41X1_HVT U9727 ( .A1(\ram[12][66] ), .A3(\ram[14][66] ), .A2(
        \ram[13][66] ), .A4(\ram[15][66] ), .S0(n8821), .S1(n8892), .Y(n7994)
         );
  MUX41X1_HVT U9728 ( .A1(\ram[8][66] ), .A3(\ram[10][66] ), .A2(\ram[9][66] ), 
        .A4(\ram[11][66] ), .S0(n5866), .S1(n7681), .Y(n7995) );
  MUX41X1_HVT U9729 ( .A1(\ram[8][67] ), .A3(\ram[10][67] ), .A2(\ram[9][67] ), 
        .A4(\ram[11][67] ), .S0(n7325), .S1(n5971), .Y(n7999) );
  MUX41X1_HVT U9730 ( .A1(\ram[4][67] ), .A3(\ram[6][67] ), .A2(\ram[5][67] ), 
        .A4(\ram[7][67] ), .S0(n5865), .S1(n5535), .Y(n8000) );
  MUX41X1_HVT U9731 ( .A1(\ram[0][67] ), .A3(\ram[2][67] ), .A2(\ram[1][67] ), 
        .A4(\ram[3][67] ), .S0(n7325), .S1(n5584), .Y(n8001) );
  MUX41X1_HVT U9732 ( .A1(\ram[12][68] ), .A3(\ram[14][68] ), .A2(
        \ram[13][68] ), .A4(\ram[15][68] ), .S0(n8821), .S1(n7681), .Y(n8002)
         );
  MUX41X1_HVT U9733 ( .A1(\ram[8][68] ), .A3(\ram[10][68] ), .A2(\ram[9][68] ), 
        .A4(\ram[11][68] ), .S0(n5993), .S1(n8892), .Y(n8003) );
  MUX41X1_HVT U9734 ( .A1(\ram[4][68] ), .A3(\ram[6][68] ), .A2(\ram[5][68] ), 
        .A4(\ram[7][68] ), .S0(n4990), .S1(n7681), .Y(n8004) );
  MUX41X1_HVT U9735 ( .A1(\ram[0][68] ), .A3(\ram[2][68] ), .A2(\ram[1][68] ), 
        .A4(\ram[3][68] ), .S0(n5866), .S1(n8892), .Y(n8005) );
  MUX41X1_HVT U9736 ( .A1(\ram[4][69] ), .A3(\ram[6][69] ), .A2(\ram[5][69] ), 
        .A4(\ram[7][69] ), .S0(n5360), .S1(n5956), .Y(n8008) );
  MUX41X1_HVT U9737 ( .A1(\ram[12][70] ), .A3(\ram[14][70] ), .A2(
        \ram[13][70] ), .A4(\ram[15][70] ), .S0(n5892), .S1(n5578), .Y(n8010)
         );
  MUX41X1_HVT U9738 ( .A1(\ram[4][70] ), .A3(\ram[6][70] ), .A2(\ram[5][70] ), 
        .A4(\ram[7][70] ), .S0(n8837), .S1(n6966), .Y(n8012) );
  MUX41X1_HVT U9739 ( .A1(\ram[4][71] ), .A3(\ram[6][71] ), .A2(\ram[5][71] ), 
        .A4(\ram[7][71] ), .S0(n5859), .S1(n5971), .Y(n8016) );
  MUX41X1_HVT U9740 ( .A1(\ram[4][72] ), .A3(\ram[6][72] ), .A2(\ram[5][72] ), 
        .A4(\ram[7][72] ), .S0(n5866), .S1(n6640), .Y(n8020) );
  MUX41X1_HVT U9741 ( .A1(\ram[12][73] ), .A3(\ram[14][73] ), .A2(
        \ram[13][73] ), .A4(\ram[15][73] ), .S0(n5957), .S1(n4983), .Y(n8022)
         );
  MUX41X1_HVT U9742 ( .A1(\ram[8][73] ), .A3(\ram[10][73] ), .A2(\ram[9][73] ), 
        .A4(\ram[11][73] ), .S0(n8829), .S1(n5629), .Y(n8023) );
  MUX41X1_HVT U9743 ( .A1(\ram[4][73] ), .A3(\ram[6][73] ), .A2(\ram[5][73] ), 
        .A4(\ram[7][73] ), .S0(n8829), .S1(n5505), .Y(n8024) );
  MUX41X1_HVT U9744 ( .A1(\ram[0][73] ), .A3(\ram[2][73] ), .A2(\ram[1][73] ), 
        .A4(\ram[3][73] ), .S0(n5967), .S1(n6640), .Y(n8025) );
  MUX41X1_HVT U9745 ( .A1(\ram[12][74] ), .A3(\ram[14][74] ), .A2(
        \ram[13][74] ), .A4(\ram[15][74] ), .S0(n5523), .S1(n5851), .Y(n8026)
         );
  MUX41X1_HVT U9746 ( .A1(\ram[8][74] ), .A3(\ram[10][74] ), .A2(\ram[9][74] ), 
        .A4(\ram[11][74] ), .S0(n5993), .S1(n7555), .Y(n8027) );
  MUX41X1_HVT U9747 ( .A1(\ram[4][74] ), .A3(\ram[6][74] ), .A2(\ram[5][74] ), 
        .A4(\ram[7][74] ), .S0(n5633), .S1(n4182), .Y(n8028) );
  MUX41X1_HVT U9748 ( .A1(n8029), .A3(n8027), .A2(n8028), .A4(n8026), .S0(
        n5654), .S1(n5755), .Y(q[74]) );
  MUX41X1_HVT U9749 ( .A1(\ram[8][75] ), .A3(\ram[10][75] ), .A2(\ram[9][75] ), 
        .A4(\ram[11][75] ), .S0(n8831), .S1(n7671), .Y(n8031) );
  MUX41X1_HVT U9750 ( .A1(\ram[4][75] ), .A3(\ram[6][75] ), .A2(\ram[5][75] ), 
        .A4(\ram[7][75] ), .S0(n7298), .S1(n5538), .Y(n8032) );
  MUX41X1_HVT U9751 ( .A1(\ram[0][75] ), .A3(\ram[2][75] ), .A2(\ram[1][75] ), 
        .A4(\ram[3][75] ), .S0(n8828), .S1(n5292), .Y(n8033) );
  MUX41X1_HVT U9752 ( .A1(n8033), .A3(n8031), .A2(n8032), .A4(n8030), .S0(
        n5363), .S1(n5092), .Y(q[75]) );
  MUX41X1_HVT U9753 ( .A1(\ram[12][76] ), .A3(\ram[14][76] ), .A2(
        \ram[13][76] ), .A4(\ram[15][76] ), .S0(n8835), .S1(n7671), .Y(n8034)
         );
  MUX41X1_HVT U9754 ( .A1(\ram[4][76] ), .A3(\ram[6][76] ), .A2(\ram[5][76] ), 
        .A4(\ram[7][76] ), .S0(n8831), .S1(n5055), .Y(n8036) );
  MUX41X1_HVT U9755 ( .A1(\ram[0][76] ), .A3(\ram[2][76] ), .A2(\ram[1][76] ), 
        .A4(\ram[3][76] ), .S0(n4949), .S1(n5538), .Y(n8037) );
  MUX41X1_HVT U9756 ( .A1(n8037), .A3(n8035), .A2(n8036), .A4(n8034), .S0(
        n5833), .S1(n6894), .Y(q[76]) );
  MUX41X1_HVT U9757 ( .A1(\ram[8][77] ), .A3(\ram[10][77] ), .A2(\ram[9][77] ), 
        .A4(\ram[11][77] ), .S0(n8794), .S1(n5476), .Y(n8039) );
  MUX41X1_HVT U9758 ( .A1(\ram[4][77] ), .A3(\ram[6][77] ), .A2(\ram[5][77] ), 
        .A4(\ram[7][77] ), .S0(n8842), .S1(n5962), .Y(n8040) );
  MUX41X1_HVT U9759 ( .A1(n8041), .A3(n8039), .A2(n8040), .A4(n8038), .S0(
        n5318), .S1(n7351), .Y(q[77]) );
  MUX41X1_HVT U9760 ( .A1(\ram[8][78] ), .A3(\ram[10][78] ), .A2(\ram[9][78] ), 
        .A4(\ram[11][78] ), .S0(n4981), .S1(n7578), .Y(n8043) );
  MUX41X1_HVT U9761 ( .A1(\ram[4][78] ), .A3(\ram[6][78] ), .A2(\ram[5][78] ), 
        .A4(\ram[7][78] ), .S0(n6009), .S1(n7578), .Y(n8044) );
  MUX41X1_HVT U9762 ( .A1(\ram[8][79] ), .A3(\ram[10][79] ), .A2(\ram[9][79] ), 
        .A4(\ram[11][79] ), .S0(n8832), .S1(n7569), .Y(n8047) );
  MUX41X1_HVT U9763 ( .A1(\ram[4][79] ), .A3(\ram[6][79] ), .A2(\ram[5][79] ), 
        .A4(\ram[7][79] ), .S0(n5751), .S1(n8890), .Y(n8048) );
  MUX41X1_HVT U9764 ( .A1(\ram[0][79] ), .A3(\ram[2][79] ), .A2(\ram[1][79] ), 
        .A4(\ram[3][79] ), .S0(n8838), .S1(n6407), .Y(n8049) );
  MUX41X1_HVT U9765 ( .A1(n8049), .A3(n8047), .A2(n8048), .A4(n8046), .S0(
        n6130), .S1(n5931), .Y(q[79]) );
  MUX41X1_HVT U9766 ( .A1(\ram[8][80] ), .A3(\ram[10][80] ), .A2(\ram[9][80] ), 
        .A4(\ram[11][80] ), .S0(n5564), .S1(n7701), .Y(n8051) );
  MUX41X1_HVT U9767 ( .A1(\ram[4][80] ), .A3(\ram[6][80] ), .A2(\ram[5][80] ), 
        .A4(\ram[7][80] ), .S0(n4980), .S1(n4940), .Y(n8052) );
  MUX41X1_HVT U9768 ( .A1(\ram[0][80] ), .A3(\ram[2][80] ), .A2(\ram[1][80] ), 
        .A4(\ram[3][80] ), .S0(n5940), .S1(n5150), .Y(n8053) );
  MUX41X1_HVT U9769 ( .A1(\ram[8][81] ), .A3(\ram[10][81] ), .A2(\ram[9][81] ), 
        .A4(\ram[11][81] ), .S0(n4949), .S1(n8866), .Y(n8055) );
  MUX41X1_HVT U9770 ( .A1(\ram[4][81] ), .A3(\ram[6][81] ), .A2(\ram[5][81] ), 
        .A4(\ram[7][81] ), .S0(n8815), .S1(n5639), .Y(n8056) );
  MUX41X1_HVT U9771 ( .A1(\ram[8][82] ), .A3(\ram[10][82] ), .A2(\ram[9][82] ), 
        .A4(\ram[11][82] ), .S0(n8843), .S1(n8897), .Y(n8059) );
  MUX41X1_HVT U9772 ( .A1(\ram[0][82] ), .A3(\ram[2][82] ), .A2(\ram[1][82] ), 
        .A4(\ram[3][82] ), .S0(n5932), .S1(n5458), .Y(n8061) );
  MUX41X1_HVT U9773 ( .A1(\ram[8][83] ), .A3(\ram[10][83] ), .A2(\ram[9][83] ), 
        .A4(\ram[11][83] ), .S0(n4905), .S1(n5551), .Y(n8063) );
  MUX41X1_HVT U9774 ( .A1(\ram[4][83] ), .A3(\ram[6][83] ), .A2(\ram[5][83] ), 
        .A4(\ram[7][83] ), .S0(n8830), .S1(n8890), .Y(n8064) );
  MUX41X1_HVT U9775 ( .A1(\ram[0][83] ), .A3(\ram[2][83] ), .A2(\ram[1][83] ), 
        .A4(\ram[3][83] ), .S0(n5499), .S1(n8888), .Y(n8065) );
  MUX41X1_HVT U9776 ( .A1(\ram[12][84] ), .A3(\ram[14][84] ), .A2(
        \ram[13][84] ), .A4(\ram[15][84] ), .S0(n6650), .S1(n6006), .Y(n8066)
         );
  MUX41X1_HVT U9777 ( .A1(\ram[8][84] ), .A3(\ram[10][84] ), .A2(\ram[9][84] ), 
        .A4(\ram[11][84] ), .S0(n7298), .S1(n5578), .Y(n8067) );
  MUX41X1_HVT U9778 ( .A1(\ram[0][84] ), .A3(\ram[2][84] ), .A2(\ram[1][84] ), 
        .A4(\ram[3][84] ), .S0(n8814), .S1(n6006), .Y(n8069) );
  MUX41X1_HVT U9779 ( .A1(n8069), .A3(n8067), .A2(n8068), .A4(n8066), .S0(
        n5225), .S1(n7666), .Y(q[84]) );
  MUX41X1_HVT U9780 ( .A1(\ram[12][85] ), .A3(\ram[14][85] ), .A2(
        \ram[13][85] ), .A4(\ram[15][85] ), .S0(n6650), .S1(n5585), .Y(n8070)
         );
  MUX41X1_HVT U9781 ( .A1(\ram[8][85] ), .A3(\ram[10][85] ), .A2(\ram[9][85] ), 
        .A4(\ram[11][85] ), .S0(n5577), .S1(n6014), .Y(n8071) );
  MUX41X1_HVT U9782 ( .A1(\ram[0][85] ), .A3(\ram[2][85] ), .A2(\ram[1][85] ), 
        .A4(\ram[3][85] ), .S0(n5004), .S1(n5611), .Y(n8073) );
  MUX41X1_HVT U9783 ( .A1(\ram[12][86] ), .A3(\ram[14][86] ), .A2(
        \ram[13][86] ), .A4(\ram[15][86] ), .S0(n8798), .S1(n8858), .Y(n8074)
         );
  MUX41X1_HVT U9784 ( .A1(\ram[8][86] ), .A3(\ram[10][86] ), .A2(\ram[9][86] ), 
        .A4(\ram[11][86] ), .S0(n8842), .S1(n6385), .Y(n8075) );
  MUX41X1_HVT U9785 ( .A1(\ram[4][86] ), .A3(\ram[6][86] ), .A2(\ram[5][86] ), 
        .A4(\ram[7][86] ), .S0(n8824), .S1(n7580), .Y(n8076) );
  MUX41X1_HVT U9786 ( .A1(\ram[0][86] ), .A3(\ram[2][86] ), .A2(\ram[1][86] ), 
        .A4(\ram[3][86] ), .S0(n4985), .S1(n8865), .Y(n8077) );
  MUX41X1_HVT U9787 ( .A1(n8077), .A3(n8075), .A2(n8076), .A4(n8074), .S0(
        n6130), .S1(n8775), .Y(q[86]) );
  MUX41X1_HVT U9788 ( .A1(\ram[0][87] ), .A3(\ram[2][87] ), .A2(\ram[1][87] ), 
        .A4(\ram[3][87] ), .S0(n8821), .S1(n4940), .Y(n8081) );
  MUX41X1_HVT U9789 ( .A1(\ram[8][88] ), .A3(\ram[10][88] ), .A2(\ram[9][88] ), 
        .A4(\ram[11][88] ), .S0(n5994), .S1(n5807), .Y(n8083) );
  MUX41X1_HVT U9790 ( .A1(\ram[4][88] ), .A3(\ram[6][88] ), .A2(\ram[5][88] ), 
        .A4(\ram[7][88] ), .S0(n5993), .S1(n5562), .Y(n8084) );
  MUX41X1_HVT U9791 ( .A1(\ram[0][88] ), .A3(\ram[2][88] ), .A2(\ram[1][88] ), 
        .A4(\ram[3][88] ), .S0(n8843), .S1(n4984), .Y(n8085) );
  MUX41X1_HVT U9792 ( .A1(\ram[12][89] ), .A3(\ram[14][89] ), .A2(
        \ram[13][89] ), .A4(\ram[15][89] ), .S0(n8829), .S1(n6755), .Y(n8086)
         );
  MUX41X1_HVT U9793 ( .A1(\ram[8][89] ), .A3(\ram[10][89] ), .A2(\ram[9][89] ), 
        .A4(\ram[11][89] ), .S0(n6741), .S1(n5361), .Y(n8087) );
  MUX41X1_HVT U9794 ( .A1(\ram[4][89] ), .A3(\ram[6][89] ), .A2(\ram[5][89] ), 
        .A4(\ram[7][89] ), .S0(n5957), .S1(n8891), .Y(n8088) );
  MUX41X1_HVT U9795 ( .A1(\ram[0][89] ), .A3(\ram[2][89] ), .A2(\ram[1][89] ), 
        .A4(\ram[3][89] ), .S0(n5859), .S1(n8886), .Y(n8089) );
  MUX41X1_HVT U9796 ( .A1(n8089), .A3(n8087), .A2(n8088), .A4(n8086), .S0(
        n5321), .S1(n8777), .Y(q[89]) );
  MUX41X1_HVT U9797 ( .A1(\ram[12][90] ), .A3(\ram[14][90] ), .A2(
        \ram[13][90] ), .A4(\ram[15][90] ), .S0(n8827), .S1(n5551), .Y(n8090)
         );
  MUX41X1_HVT U9798 ( .A1(\ram[0][91] ), .A3(\ram[2][91] ), .A2(\ram[1][91] ), 
        .A4(\ram[3][91] ), .S0(n5569), .S1(n8897), .Y(n8097) );
  MUX41X1_HVT U9799 ( .A1(\ram[8][92] ), .A3(\ram[10][92] ), .A2(\ram[9][92] ), 
        .A4(\ram[11][92] ), .S0(n5994), .S1(n7569), .Y(n8099) );
  MUX41X1_HVT U9800 ( .A1(\ram[4][92] ), .A3(\ram[6][92] ), .A2(\ram[5][92] ), 
        .A4(\ram[7][92] ), .S0(n4975), .S1(n6137), .Y(n8100) );
  MUX41X1_HVT U9801 ( .A1(\ram[0][92] ), .A3(\ram[2][92] ), .A2(\ram[1][92] ), 
        .A4(\ram[3][92] ), .S0(n6413), .S1(n5639), .Y(n8101) );
  MUX41X1_HVT U9802 ( .A1(\ram[12][93] ), .A3(\ram[14][93] ), .A2(
        \ram[13][93] ), .A4(\ram[15][93] ), .S0(n8827), .S1(n5584), .Y(n8102)
         );
  MUX41X1_HVT U9803 ( .A1(\ram[8][93] ), .A3(\ram[10][93] ), .A2(\ram[9][93] ), 
        .A4(\ram[11][93] ), .S0(n5353), .S1(n8898), .Y(n8103) );
  MUX41X1_HVT U9804 ( .A1(\ram[4][93] ), .A3(\ram[6][93] ), .A2(\ram[5][93] ), 
        .A4(\ram[7][93] ), .S0(n7324), .S1(n8898), .Y(n8104) );
  MUX41X1_HVT U9805 ( .A1(\ram[4][94] ), .A3(\ram[6][94] ), .A2(\ram[5][94] ), 
        .A4(\ram[7][94] ), .S0(n5993), .S1(n6417), .Y(n8108) );
  MUX41X1_HVT U9806 ( .A1(\ram[0][94] ), .A3(\ram[2][94] ), .A2(\ram[1][94] ), 
        .A4(\ram[3][94] ), .S0(n4918), .S1(n4974), .Y(n8109) );
  MUX41X1_HVT U9807 ( .A1(\ram[8][95] ), .A3(\ram[10][95] ), .A2(\ram[9][95] ), 
        .A4(\ram[11][95] ), .S0(n8818), .S1(n4789), .Y(n8111) );
  MUX41X1_HVT U9808 ( .A1(\ram[4][95] ), .A3(\ram[6][95] ), .A2(\ram[5][95] ), 
        .A4(\ram[7][95] ), .S0(n8811), .S1(n8898), .Y(n8112) );
  MUX41X1_HVT U9809 ( .A1(\ram[0][95] ), .A3(\ram[2][95] ), .A2(\ram[1][95] ), 
        .A4(\ram[3][95] ), .S0(n8829), .S1(n7579), .Y(n8113) );
  MUX41X1_HVT U9810 ( .A1(\ram[8][96] ), .A3(\ram[10][96] ), .A2(\ram[9][96] ), 
        .A4(\ram[11][96] ), .S0(n6029), .S1(n7327), .Y(n8115) );
  MUX41X1_HVT U9811 ( .A1(\ram[4][96] ), .A3(\ram[6][96] ), .A2(\ram[5][96] ), 
        .A4(\ram[7][96] ), .S0(n5322), .S1(n7580), .Y(n8116) );
  MUX41X1_HVT U9812 ( .A1(\ram[0][96] ), .A3(\ram[2][96] ), .A2(\ram[1][96] ), 
        .A4(\ram[3][96] ), .S0(n8810), .S1(n7581), .Y(n8117) );
  MUX41X1_HVT U9813 ( .A1(\ram[12][97] ), .A3(\ram[14][97] ), .A2(
        \ram[13][97] ), .A4(\ram[15][97] ), .S0(n5994), .S1(n5123), .Y(n8118)
         );
  MUX41X1_HVT U9814 ( .A1(\ram[8][97] ), .A3(\ram[10][97] ), .A2(\ram[9][97] ), 
        .A4(\ram[11][97] ), .S0(n6028), .S1(n7669), .Y(n8119) );
  MUX41X1_HVT U9815 ( .A1(\ram[4][97] ), .A3(\ram[6][97] ), .A2(\ram[5][97] ), 
        .A4(\ram[7][97] ), .S0(n7549), .S1(n7580), .Y(n8120) );
  MUX41X1_HVT U9816 ( .A1(\ram[12][98] ), .A3(\ram[14][98] ), .A2(
        \ram[13][98] ), .A4(\ram[15][98] ), .S0(n8822), .S1(n6744), .Y(n8122)
         );
  MUX41X1_HVT U9817 ( .A1(\ram[8][98] ), .A3(\ram[10][98] ), .A2(\ram[9][98] ), 
        .A4(\ram[11][98] ), .S0(n8836), .S1(n8886), .Y(n8123) );
  MUX41X1_HVT U9818 ( .A1(\ram[4][98] ), .A3(\ram[6][98] ), .A2(\ram[5][98] ), 
        .A4(\ram[7][98] ), .S0(n6028), .S1(n4166), .Y(n8124) );
  MUX41X1_HVT U9819 ( .A1(\ram[0][98] ), .A3(\ram[2][98] ), .A2(\ram[1][98] ), 
        .A4(\ram[3][98] ), .S0(n5360), .S1(n7669), .Y(n8125) );
  MUX41X1_HVT U9820 ( .A1(\ram[8][99] ), .A3(\ram[10][99] ), .A2(\ram[9][99] ), 
        .A4(\ram[11][99] ), .S0(n6008), .S1(n5924), .Y(n8127) );
  MUX41X1_HVT U9821 ( .A1(\ram[4][99] ), .A3(\ram[6][99] ), .A2(\ram[5][99] ), 
        .A4(\ram[7][99] ), .S0(n5475), .S1(n5636), .Y(n8128) );
  MUX41X1_HVT U9822 ( .A1(\ram[0][99] ), .A3(\ram[2][99] ), .A2(\ram[1][99] ), 
        .A4(\ram[3][99] ), .S0(n7336), .S1(n7676), .Y(n8129) );
  MUX41X1_HVT U9823 ( .A1(n8129), .A3(n8127), .A2(n8128), .A4(n8126), .S0(
        n5323), .S1(n8768), .Y(q[99]) );
  MUX41X1_HVT U9824 ( .A1(\ram[12][100] ), .A3(\ram[14][100] ), .A2(
        \ram[13][100] ), .A4(\ram[15][100] ), .S0(n7320), .S1(n7676), .Y(n8130) );
  MUX41X1_HVT U9825 ( .A1(\ram[8][100] ), .A3(\ram[10][100] ), .A2(
        \ram[9][100] ), .A4(\ram[11][100] ), .S0(n6007), .S1(n7676), .Y(n8131)
         );
  MUX41X1_HVT U9826 ( .A1(\ram[4][100] ), .A3(\ram[6][100] ), .A2(
        \ram[5][100] ), .A4(\ram[7][100] ), .S0(n7554), .S1(n7675), .Y(n8132)
         );
  MUX41X1_HVT U9827 ( .A1(\ram[0][100] ), .A3(\ram[2][100] ), .A2(
        \ram[1][100] ), .A4(\ram[3][100] ), .S0(n8792), .S1(n7675), .Y(n8133)
         );
  MUX41X1_HVT U9828 ( .A1(n8133), .A3(n8131), .A2(n8132), .A4(n8130), .S0(
        n5799), .S1(n8776), .Y(q[100]) );
  MUX41X1_HVT U9829 ( .A1(\ram[8][101] ), .A3(\ram[10][101] ), .A2(
        \ram[9][101] ), .A4(\ram[11][101] ), .S0(n4884), .S1(n5292), .Y(n8135)
         );
  MUX41X1_HVT U9830 ( .A1(\ram[4][101] ), .A3(\ram[6][101] ), .A2(
        \ram[5][101] ), .A4(\ram[7][101] ), .S0(n7336), .S1(n7675), .Y(n8136)
         );
  MUX41X1_HVT U9831 ( .A1(\ram[0][101] ), .A3(\ram[2][101] ), .A2(
        \ram[1][101] ), .A4(\ram[3][101] ), .S0(n8826), .S1(n5924), .Y(n8137)
         );
  MUX41X1_HVT U9832 ( .A1(\ram[8][102] ), .A3(\ram[10][102] ), .A2(
        \ram[9][102] ), .A4(\ram[11][102] ), .S0(n8818), .S1(n5144), .Y(n8139)
         );
  MUX41X1_HVT U9833 ( .A1(\ram[4][102] ), .A3(\ram[6][102] ), .A2(
        \ram[5][102] ), .A4(\ram[7][102] ), .S0(n8818), .S1(n6034), .Y(n8140)
         );
  MUX41X1_HVT U9834 ( .A1(\ram[8][103] ), .A3(\ram[10][103] ), .A2(
        \ram[9][103] ), .A4(\ram[11][103] ), .S0(n7335), .S1(n5652), .Y(n8143)
         );
  MUX41X1_HVT U9835 ( .A1(\ram[0][103] ), .A3(\ram[2][103] ), .A2(
        \ram[1][103] ), .A4(\ram[3][103] ), .S0(n4980), .S1(n8908), .Y(n8145)
         );
  MUX41X1_HVT U9836 ( .A1(n8145), .A3(n8143), .A2(n8144), .A4(n8142), .S0(
        n7293), .S1(n7547), .Y(q[103]) );
  MUX41X1_HVT U9837 ( .A1(\ram[12][104] ), .A3(\ram[14][104] ), .A2(
        \ram[13][104] ), .A4(\ram[15][104] ), .S0(n8836), .S1(n8908), .Y(n8146) );
  MUX41X1_HVT U9838 ( .A1(\ram[8][104] ), .A3(\ram[10][104] ), .A2(
        \ram[9][104] ), .A4(\ram[11][104] ), .S0(n8818), .S1(n5639), .Y(n8147)
         );
  MUX41X1_HVT U9839 ( .A1(\ram[4][104] ), .A3(\ram[6][104] ), .A2(
        \ram[5][104] ), .A4(\ram[7][104] ), .S0(n7335), .S1(n8866), .Y(n8148)
         );
  MUX41X1_HVT U9840 ( .A1(\ram[0][104] ), .A3(\ram[2][104] ), .A2(
        \ram[1][104] ), .A4(\ram[3][104] ), .S0(n8818), .S1(n6034), .Y(n8149)
         );
  MUX41X1_HVT U9841 ( .A1(\ram[4][105] ), .A3(\ram[6][105] ), .A2(
        \ram[5][105] ), .A4(\ram[7][105] ), .S0(n5948), .S1(n5570), .Y(n8152)
         );
  MUX41X1_HVT U9842 ( .A1(\ram[12][106] ), .A3(\ram[14][106] ), .A2(
        \ram[13][106] ), .A4(\ram[15][106] ), .S0(n8838), .S1(n5572), .Y(n8154) );
  MUX41X1_HVT U9843 ( .A1(\ram[8][106] ), .A3(\ram[10][106] ), .A2(
        \ram[9][106] ), .A4(\ram[11][106] ), .S0(n8824), .S1(n5582), .Y(n8155)
         );
  MUX41X1_HVT U9844 ( .A1(\ram[4][106] ), .A3(\ram[6][106] ), .A2(
        \ram[5][106] ), .A4(\ram[7][106] ), .S0(n5475), .S1(n5479), .Y(n8156)
         );
  MUX41X1_HVT U9845 ( .A1(\ram[0][106] ), .A3(\ram[2][106] ), .A2(
        \ram[1][106] ), .A4(\ram[3][106] ), .S0(n6183), .S1(n7329), .Y(n8157)
         );
  MUX41X1_HVT U9846 ( .A1(\ram[12][107] ), .A3(\ram[14][107] ), .A2(
        \ram[13][107] ), .A4(\ram[15][107] ), .S0(n5932), .S1(n5447), .Y(n8158) );
  MUX41X1_HVT U9847 ( .A1(\ram[8][107] ), .A3(\ram[10][107] ), .A2(
        \ram[9][107] ), .A4(\ram[11][107] ), .S0(n4884), .S1(n5889), .Y(n8159)
         );
  MUX41X1_HVT U9848 ( .A1(\ram[4][107] ), .A3(\ram[6][107] ), .A2(
        \ram[5][107] ), .A4(\ram[7][107] ), .S0(n6009), .S1(n1389), .Y(n8160)
         );
  MUX41X1_HVT U9849 ( .A1(\ram[0][107] ), .A3(\ram[2][107] ), .A2(
        \ram[1][107] ), .A4(\ram[3][107] ), .S0(n8793), .S1(n8854), .Y(n8161)
         );
  MUX41X1_HVT U9850 ( .A1(n8161), .A3(n8159), .A2(n8160), .A4(n8158), .S0(
        n5097), .S1(n5324), .Y(q[107]) );
  MUX41X1_HVT U9851 ( .A1(\ram[8][108] ), .A3(\ram[10][108] ), .A2(
        \ram[9][108] ), .A4(\ram[11][108] ), .S0(n8816), .S1(n4940), .Y(n8163)
         );
  MUX41X1_HVT U9852 ( .A1(\ram[0][108] ), .A3(\ram[2][108] ), .A2(
        \ram[1][108] ), .A4(\ram[3][108] ), .S0(n5612), .S1(n5500), .Y(n8165)
         );
  MUX41X1_HVT U9853 ( .A1(\ram[12][109] ), .A3(\ram[14][109] ), .A2(
        \ram[13][109] ), .A4(\ram[15][109] ), .S0(n6017), .S1(n6253), .Y(n8166) );
  MUX41X1_HVT U9854 ( .A1(\ram[8][109] ), .A3(\ram[10][109] ), .A2(
        \ram[9][109] ), .A4(\ram[11][109] ), .S0(n5499), .S1(n4921), .Y(n8167)
         );
  MUX41X1_HVT U9855 ( .A1(\ram[4][109] ), .A3(\ram[6][109] ), .A2(
        \ram[5][109] ), .A4(\ram[7][109] ), .S0(n8841), .S1(n5500), .Y(n8168)
         );
  MUX41X1_HVT U9856 ( .A1(\ram[0][109] ), .A3(\ram[2][109] ), .A2(
        \ram[1][109] ), .A4(\ram[3][109] ), .S0(n5499), .S1(n5500), .Y(n8169)
         );
  MUX41X1_HVT U9857 ( .A1(n8169), .A3(n8167), .A2(n8168), .A4(n8166), .S0(
        n5323), .S1(n5092), .Y(q[109]) );
  MUX41X1_HVT U9858 ( .A1(\ram[12][110] ), .A3(\ram[14][110] ), .A2(
        \ram[13][110] ), .A4(\ram[15][110] ), .S0(n6757), .S1(n6966), .Y(n8170) );
  MUX41X1_HVT U9859 ( .A1(\ram[8][110] ), .A3(\ram[10][110] ), .A2(
        \ram[9][110] ), .A4(\ram[11][110] ), .S0(n7550), .S1(n5135), .Y(n8171)
         );
  MUX41X1_HVT U9860 ( .A1(\ram[4][110] ), .A3(\ram[6][110] ), .A2(
        \ram[5][110] ), .A4(\ram[7][110] ), .S0(n5888), .S1(n8904), .Y(n8172)
         );
  MUX41X1_HVT U9861 ( .A1(\ram[0][110] ), .A3(\ram[2][110] ), .A2(
        \ram[1][110] ), .A4(\ram[3][110] ), .S0(n5592), .S1(n7564), .Y(n8173)
         );
  MUX41X1_HVT U9862 ( .A1(\ram[12][111] ), .A3(\ram[14][111] ), .A2(
        \ram[13][111] ), .A4(\ram[15][111] ), .S0(n8791), .S1(n5729), .Y(n8174) );
  MUX41X1_HVT U9863 ( .A1(\ram[8][111] ), .A3(\ram[10][111] ), .A2(
        \ram[9][111] ), .A4(\ram[11][111] ), .S0(n5633), .S1(n7329), .Y(n8175)
         );
  MUX41X1_HVT U9864 ( .A1(\ram[4][111] ), .A3(\ram[6][111] ), .A2(
        \ram[5][111] ), .A4(\ram[7][111] ), .S0(n5050), .S1(n5729), .Y(n8176)
         );
  MUX41X1_HVT U9865 ( .A1(\ram[0][111] ), .A3(\ram[2][111] ), .A2(
        \ram[1][111] ), .A4(\ram[3][111] ), .S0(n7335), .S1(n5139), .Y(n8177)
         );
  MUX41X1_HVT U9866 ( .A1(\ram[12][112] ), .A3(\ram[14][112] ), .A2(
        \ram[13][112] ), .A4(\ram[15][112] ), .S0(n5050), .S1(n5939), .Y(n8178) );
  MUX41X1_HVT U9867 ( .A1(\ram[8][112] ), .A3(\ram[10][112] ), .A2(
        \ram[9][112] ), .A4(\ram[11][112] ), .S0(n8792), .S1(n5728), .Y(n8179)
         );
  MUX41X1_HVT U9868 ( .A1(\ram[4][112] ), .A3(\ram[6][112] ), .A2(
        \ram[5][112] ), .A4(\ram[7][112] ), .S0(n8791), .S1(n5807), .Y(n8180)
         );
  MUX41X1_HVT U9869 ( .A1(\ram[8][113] ), .A3(\ram[10][113] ), .A2(
        \ram[9][113] ), .A4(\ram[11][113] ), .S0(n4980), .S1(n8905), .Y(n8183)
         );
  MUX41X1_HVT U9870 ( .A1(\ram[4][113] ), .A3(\ram[6][113] ), .A2(
        \ram[5][113] ), .A4(\ram[7][113] ), .S0(n8850), .S1(n5728), .Y(n8184)
         );
  MUX41X1_HVT U9871 ( .A1(\ram[0][113] ), .A3(\ram[2][113] ), .A2(
        \ram[1][113] ), .A4(\ram[3][113] ), .S0(n8791), .S1(n6137), .Y(n8185)
         );
  MUX41X1_HVT U9872 ( .A1(\ram[12][114] ), .A3(\ram[14][114] ), .A2(
        \ram[13][114] ), .A4(\ram[15][114] ), .S0(n6020), .S1(n7680), .Y(n8186) );
  MUX41X1_HVT U9873 ( .A1(\ram[8][114] ), .A3(\ram[10][114] ), .A2(
        \ram[9][114] ), .A4(\ram[11][114] ), .S0(n6650), .S1(n5538), .Y(n8187)
         );
  MUX41X1_HVT U9874 ( .A1(\ram[4][114] ), .A3(\ram[6][114] ), .A2(
        \ram[5][114] ), .A4(\ram[7][114] ), .S0(n8822), .S1(n5823), .Y(n8188)
         );
  MUX41X1_HVT U9875 ( .A1(\ram[0][114] ), .A3(\ram[2][114] ), .A2(
        \ram[1][114] ), .A4(\ram[3][114] ), .S0(n5946), .S1(n5609), .Y(n8189)
         );
  MUX41X1_HVT U9876 ( .A1(\ram[12][115] ), .A3(\ram[14][115] ), .A2(
        \ram[13][115] ), .A4(\ram[15][115] ), .S0(n5733), .S1(n4994), .Y(n8190) );
  MUX41X1_HVT U9877 ( .A1(\ram[4][115] ), .A3(\ram[6][115] ), .A2(
        \ram[5][115] ), .A4(\ram[7][115] ), .S0(n7298), .S1(n8892), .Y(n8192)
         );
  MUX41X1_HVT U9878 ( .A1(\ram[0][115] ), .A3(\ram[2][115] ), .A2(
        \ram[1][115] ), .A4(\ram[3][115] ), .S0(n5734), .S1(n7681), .Y(n8193)
         );
  MUX41X1_HVT U9879 ( .A1(\ram[8][116] ), .A3(\ram[10][116] ), .A2(
        \ram[9][116] ), .A4(\ram[11][116] ), .S0(n8848), .S1(n5535), .Y(n8195)
         );
  MUX41X1_HVT U9880 ( .A1(\ram[4][116] ), .A3(\ram[6][116] ), .A2(
        \ram[5][116] ), .A4(\ram[7][116] ), .S0(n8846), .S1(n5055), .Y(n8196)
         );
  MUX41X1_HVT U9881 ( .A1(n8197), .A3(n8195), .A2(n8196), .A4(n8194), .S0(
        n5756), .S1(n6751), .Y(q[116]) );
  MUX41X1_HVT U9882 ( .A1(\ram[12][117] ), .A3(\ram[14][117] ), .A2(
        \ram[13][117] ), .A4(\ram[15][117] ), .S0(n8830), .S1(n6965), .Y(n8198) );
  MUX41X1_HVT U9883 ( .A1(\ram[4][117] ), .A3(\ram[6][117] ), .A2(
        \ram[5][117] ), .A4(\ram[7][117] ), .S0(n6741), .S1(n5515), .Y(n8200)
         );
  MUX41X1_HVT U9884 ( .A1(\ram[0][117] ), .A3(\ram[2][117] ), .A2(
        \ram[1][117] ), .A4(\ram[3][117] ), .S0(n8843), .S1(n8858), .Y(n8201)
         );
  MUX41X1_HVT U9885 ( .A1(n8201), .A3(n8199), .A2(n8200), .A4(n8198), .S0(
        n8761), .S1(n5362), .Y(q[117]) );
  MUX41X1_HVT U9886 ( .A1(\ram[8][118] ), .A3(\ram[10][118] ), .A2(
        \ram[9][118] ), .A4(\ram[11][118] ), .S0(n5076), .S1(n5515), .Y(n8203)
         );
  MUX41X1_HVT U9887 ( .A1(\ram[0][118] ), .A3(\ram[2][118] ), .A2(
        \ram[1][118] ), .A4(\ram[3][118] ), .S0(n8830), .S1(n6965), .Y(n8205)
         );
  MUX41X1_HVT U9888 ( .A1(\ram[12][119] ), .A3(\ram[14][119] ), .A2(
        \ram[13][119] ), .A4(\ram[15][119] ), .S0(n8830), .S1(n5515), .Y(n8206) );
  MUX41X1_HVT U9889 ( .A1(\ram[8][119] ), .A3(\ram[10][119] ), .A2(
        \ram[9][119] ), .A4(\ram[11][119] ), .S0(n5751), .S1(n5962), .Y(n8207)
         );
  MUX41X1_HVT U9890 ( .A1(\ram[4][119] ), .A3(\ram[6][119] ), .A2(
        \ram[5][119] ), .A4(\ram[7][119] ), .S0(n5865), .S1(n6965), .Y(n8208)
         );
  MUX41X1_HVT U9891 ( .A1(\ram[0][119] ), .A3(\ram[2][119] ), .A2(
        \ram[1][119] ), .A4(\ram[3][119] ), .S0(n6741), .S1(n5290), .Y(n8209)
         );
  MUX41X1_HVT U9892 ( .A1(\ram[12][120] ), .A3(\ram[14][120] ), .A2(
        \ram[13][120] ), .A4(\ram[15][120] ), .S0(n6741), .S1(n5144), .Y(n8210) );
  MUX41X1_HVT U9893 ( .A1(\ram[8][120] ), .A3(\ram[10][120] ), .A2(
        \ram[9][120] ), .A4(\ram[11][120] ), .S0(n8830), .S1(n8889), .Y(n8211)
         );
  MUX41X1_HVT U9894 ( .A1(\ram[4][120] ), .A3(\ram[6][120] ), .A2(
        \ram[5][120] ), .A4(\ram[7][120] ), .S0(n5957), .S1(n7564), .Y(n8212)
         );
  MUX41X1_HVT U9895 ( .A1(\ram[0][120] ), .A3(\ram[2][120] ), .A2(
        \ram[1][120] ), .A4(\ram[3][120] ), .S0(n5967), .S1(n7563), .Y(n8213)
         );
  MUX41X1_HVT U9896 ( .A1(\ram[12][121] ), .A3(\ram[14][121] ), .A2(
        \ram[13][121] ), .A4(\ram[15][121] ), .S0(n5957), .S1(n7563), .Y(n8214) );
  MUX41X1_HVT U9897 ( .A1(\ram[8][121] ), .A3(\ram[10][121] ), .A2(
        \ram[9][121] ), .A4(\ram[11][121] ), .S0(n5558), .S1(n7687), .Y(n8215)
         );
  MUX41X1_HVT U9898 ( .A1(\ram[4][121] ), .A3(\ram[6][121] ), .A2(
        \ram[5][121] ), .A4(\ram[7][121] ), .S0(n8837), .S1(n7689), .Y(n8216)
         );
  MUX41X1_HVT U9899 ( .A1(\ram[0][121] ), .A3(\ram[2][121] ), .A2(
        \ram[1][121] ), .A4(\ram[3][121] ), .S0(n6741), .S1(n5579), .Y(n8217)
         );
  MUX41X1_HVT U9900 ( .A1(n8217), .A3(n8215), .A2(n8216), .A4(n8214), .S0(
        n6259), .S1(n7666), .Y(q[121]) );
  MUX41X1_HVT U9901 ( .A1(\ram[12][122] ), .A3(\ram[14][122] ), .A2(
        \ram[13][122] ), .A4(\ram[15][122] ), .S0(n7321), .S1(n6035), .Y(n8218) );
  MUX41X1_HVT U9902 ( .A1(\ram[8][122] ), .A3(\ram[10][122] ), .A2(
        \ram[9][122] ), .A4(\ram[11][122] ), .S0(n5859), .S1(n7694), .Y(n8219)
         );
  MUX41X1_HVT U9903 ( .A1(\ram[4][122] ), .A3(\ram[6][122] ), .A2(
        \ram[5][122] ), .A4(\ram[7][122] ), .S0(n5957), .S1(n5956), .Y(n8220)
         );
  MUX41X1_HVT U9904 ( .A1(\ram[0][122] ), .A3(\ram[2][122] ), .A2(
        \ram[1][122] ), .A4(\ram[3][122] ), .S0(n8821), .S1(n7687), .Y(n8221)
         );
  MUX41X1_HVT U9905 ( .A1(n8221), .A3(n8219), .A2(n8220), .A4(n8218), .S0(
        n6756), .S1(n8778), .Y(q[122]) );
  MUX41X1_HVT U9906 ( .A1(\ram[8][123] ), .A3(\ram[10][123] ), .A2(
        \ram[9][123] ), .A4(\ram[11][123] ), .S0(n8819), .S1(n6762), .Y(n8223)
         );
  MUX41X1_HVT U9907 ( .A1(\ram[4][123] ), .A3(\ram[6][123] ), .A2(
        \ram[5][123] ), .A4(\ram[7][123] ), .S0(n8811), .S1(n8856), .Y(n8224)
         );
  MUX41X1_HVT U9908 ( .A1(\ram[0][123] ), .A3(\ram[2][123] ), .A2(
        \ram[1][123] ), .A4(\ram[3][123] ), .S0(n7330), .S1(n5006), .Y(n8225)
         );
  MUX41X1_HVT U9909 ( .A1(\ram[8][124] ), .A3(\ram[10][124] ), .A2(
        \ram[9][124] ), .A4(\ram[11][124] ), .S0(n8819), .S1(n5758), .Y(n8227)
         );
  MUX41X1_HVT U9910 ( .A1(\ram[4][124] ), .A3(\ram[6][124] ), .A2(
        \ram[5][124] ), .A4(\ram[7][124] ), .S0(n7330), .S1(n5869), .Y(n8228)
         );
  MUX41X1_HVT U9911 ( .A1(\ram[0][124] ), .A3(\ram[2][124] ), .A2(
        \ram[1][124] ), .A4(\ram[3][124] ), .S0(n8819), .S1(n5731), .Y(n8229)
         );
  MUX41X1_HVT U9912 ( .A1(n8229), .A3(n8227), .A2(n8228), .A4(n8226), .S0(
        n8761), .S1(n8769), .Y(q[124]) );
  MUX41X1_HVT U9913 ( .A1(\ram[8][125] ), .A3(\ram[10][125] ), .A2(
        \ram[9][125] ), .A4(\ram[11][125] ), .S0(n6024), .S1(n6395), .Y(n8231)
         );
  MUX41X1_HVT U9914 ( .A1(\ram[4][125] ), .A3(\ram[6][125] ), .A2(
        \ram[5][125] ), .A4(\ram[7][125] ), .S0(n7330), .S1(n5609), .Y(n8232)
         );
  MUX41X1_HVT U9915 ( .A1(\ram[0][125] ), .A3(\ram[2][125] ), .A2(
        \ram[1][125] ), .A4(\ram[3][125] ), .S0(n8811), .S1(n7695), .Y(n8233)
         );
  MUX41X1_HVT U9916 ( .A1(n8233), .A3(n8231), .A2(n8232), .A4(n8230), .S0(
        n5225), .S1(n7351), .Y(q[125]) );
  MUX41X1_HVT U9917 ( .A1(\ram[8][126] ), .A3(\ram[10][126] ), .A2(
        \ram[9][126] ), .A4(\ram[11][126] ), .S0(n6017), .S1(n8888), .Y(n8235)
         );
  MUX41X1_HVT U9918 ( .A1(\ram[4][126] ), .A3(\ram[6][126] ), .A2(
        \ram[5][126] ), .A4(\ram[7][126] ), .S0(n8816), .S1(n6738), .Y(n8236)
         );
  MUX41X1_HVT U9919 ( .A1(\ram[0][126] ), .A3(\ram[2][126] ), .A2(
        \ram[1][126] ), .A4(\ram[3][126] ), .S0(n8808), .S1(n6738), .Y(n8237)
         );
  MUX41X1_HVT U9920 ( .A1(\ram[8][127] ), .A3(\ram[10][127] ), .A2(
        \ram[9][127] ), .A4(\ram[11][127] ), .S0(n6757), .S1(n6755), .Y(n8239)
         );
  MUX41X1_HVT U9921 ( .A1(\ram[4][127] ), .A3(\ram[6][127] ), .A2(
        \ram[5][127] ), .A4(\ram[7][127] ), .S0(n8832), .S1(n4820), .Y(n8240)
         );
  MUX41X1_HVT U9922 ( .A1(n8241), .A3(n8239), .A2(n8240), .A4(n8238), .S0(
        n7543), .S1(n8777), .Y(q[127]) );
  MUX41X1_HVT U9923 ( .A1(\ram[8][129] ), .A3(\ram[10][129] ), .A2(
        \ram[9][129] ), .A4(\ram[11][129] ), .S0(n7551), .S1(n8905), .Y(n8247)
         );
  MUX41X1_HVT U9924 ( .A1(\ram[4][129] ), .A3(\ram[6][129] ), .A2(
        \ram[5][129] ), .A4(\ram[7][129] ), .S0(n8844), .S1(n5226), .Y(n8248)
         );
  MUX41X1_HVT U9925 ( .A1(\ram[8][130] ), .A3(\ram[10][130] ), .A2(
        \ram[9][130] ), .A4(\ram[11][130] ), .S0(n5231), .S1(n4992), .Y(n8251)
         );
  MUX41X1_HVT U9926 ( .A1(\ram[0][130] ), .A3(\ram[2][130] ), .A2(
        \ram[1][130] ), .A4(\ram[3][130] ), .S0(n8823), .S1(n4992), .Y(n8253)
         );
  MUX41X1_HVT U9927 ( .A1(n8253), .A3(n8251), .A2(n8252), .A4(n8250), .S0(
        n5833), .S1(n5307), .Y(q[130]) );
  MUX41X1_HVT U9928 ( .A1(\ram[12][131] ), .A3(\ram[14][131] ), .A2(
        \ram[13][131] ), .A4(\ram[15][131] ), .S0(n8831), .S1(n5054), .Y(n8254) );
  MUX41X1_HVT U9929 ( .A1(\ram[8][132] ), .A3(\ram[10][132] ), .A2(
        \ram[9][132] ), .A4(\ram[11][132] ), .S0(n4981), .S1(n7679), .Y(n8259)
         );
  MUX41X1_HVT U9930 ( .A1(\ram[4][132] ), .A3(\ram[6][132] ), .A2(
        \ram[5][132] ), .A4(\ram[7][132] ), .S0(n7335), .S1(n5921), .Y(n8260)
         );
  MUX41X1_HVT U9931 ( .A1(\ram[8][133] ), .A3(\ram[10][133] ), .A2(
        \ram[9][133] ), .A4(\ram[11][133] ), .S0(n8825), .S1(n6755), .Y(n8263)
         );
  MUX41X1_HVT U9932 ( .A1(\ram[8][134] ), .A3(\ram[10][134] ), .A2(
        \ram[9][134] ), .A4(\ram[11][134] ), .S0(n8817), .S1(n7679), .Y(n8267)
         );
  MUX41X1_HVT U9933 ( .A1(\ram[4][135] ), .A3(\ram[6][135] ), .A2(
        \ram[5][135] ), .A4(\ram[7][135] ), .S0(n5564), .S1(n7667), .Y(n8272)
         );
  MUX41X1_HVT U9934 ( .A1(\ram[12][136] ), .A3(\ram[14][136] ), .A2(
        \ram[13][136] ), .A4(\ram[15][136] ), .S0(n5888), .S1(n5148), .Y(n8274) );
  MUX41X1_HVT U9935 ( .A1(\ram[0][136] ), .A3(\ram[2][136] ), .A2(
        \ram[1][136] ), .A4(\ram[3][136] ), .S0(n6413), .S1(n5135), .Y(n8277)
         );
  MUX41X1_HVT U9936 ( .A1(\ram[8][137] ), .A3(\ram[10][137] ), .A2(
        \ram[9][137] ), .A4(\ram[11][137] ), .S0(n6005), .S1(n8853), .Y(n8279)
         );
  MUX41X1_HVT U9937 ( .A1(\ram[4][137] ), .A3(\ram[6][137] ), .A2(
        \ram[5][137] ), .A4(\ram[7][137] ), .S0(n5888), .S1(n5148), .Y(n8280)
         );
  MUX41X1_HVT U9938 ( .A1(\ram[0][138] ), .A3(\ram[2][138] ), .A2(
        \ram[1][138] ), .A4(\ram[3][138] ), .S0(n4973), .S1(n5512), .Y(n8285)
         );
  MUX41X1_HVT U9939 ( .A1(\ram[4][139] ), .A3(\ram[6][139] ), .A2(
        \ram[5][139] ), .A4(\ram[7][139] ), .S0(n8841), .S1(n8877), .Y(n8288)
         );
  MUX41X1_HVT U9940 ( .A1(\ram[0][139] ), .A3(\ram[2][139] ), .A2(
        \ram[1][139] ), .A4(\ram[3][139] ), .S0(n8817), .S1(n6743), .Y(n8289)
         );
  MUX41X1_HVT U9941 ( .A1(\ram[12][140] ), .A3(\ram[14][140] ), .A2(
        \ram[13][140] ), .A4(\ram[15][140] ), .S0(n8835), .S1(n8861), .Y(n8290) );
  MUX41X1_HVT U9942 ( .A1(\ram[8][140] ), .A3(\ram[10][140] ), .A2(
        \ram[9][140] ), .A4(\ram[11][140] ), .S0(n8797), .S1(n8864), .Y(n8291)
         );
  MUX41X1_HVT U9943 ( .A1(\ram[4][140] ), .A3(\ram[6][140] ), .A2(
        \ram[5][140] ), .A4(\ram[7][140] ), .S0(n8797), .S1(n7575), .Y(n8292)
         );
  MUX41X1_HVT U9944 ( .A1(\ram[0][140] ), .A3(\ram[2][140] ), .A2(
        \ram[1][140] ), .A4(\ram[3][140] ), .S0(n8797), .S1(n7686), .Y(n8293)
         );
  MUX41X1_HVT U9945 ( .A1(n8293), .A3(n8291), .A2(n8292), .A4(n8290), .S0(
        n5752), .S1(n6754), .Y(q[140]) );
  MUX41X1_HVT U9946 ( .A1(\ram[12][141] ), .A3(\ram[14][141] ), .A2(
        \ram[13][141] ), .A4(\ram[15][141] ), .S0(n6008), .S1(n7328), .Y(n8294) );
  MUX41X1_HVT U9947 ( .A1(\ram[8][141] ), .A3(\ram[10][141] ), .A2(
        \ram[9][141] ), .A4(\ram[11][141] ), .S0(n7337), .S1(n5560), .Y(n8295)
         );
  MUX41X1_HVT U9948 ( .A1(\ram[4][141] ), .A3(\ram[6][141] ), .A2(
        \ram[5][141] ), .A4(\ram[7][141] ), .S0(n7338), .S1(n7328), .Y(n8296)
         );
  MUX41X1_HVT U9949 ( .A1(\ram[0][141] ), .A3(\ram[2][141] ), .A2(
        \ram[1][141] ), .A4(\ram[3][141] ), .S0(n5475), .S1(n7328), .Y(n8297)
         );
  MUX41X1_HVT U9950 ( .A1(\ram[8][142] ), .A3(\ram[10][142] ), .A2(
        \ram[9][142] ), .A4(\ram[11][142] ), .S0(n8826), .S1(n8875), .Y(n8299)
         );
  MUX41X1_HVT U9951 ( .A1(\ram[12][143] ), .A3(\ram[14][143] ), .A2(
        \ram[13][143] ), .A4(\ram[15][143] ), .S0(n8808), .S1(n6386), .Y(n8302) );
  MUX41X1_HVT U9952 ( .A1(\ram[8][143] ), .A3(\ram[10][143] ), .A2(
        \ram[9][143] ), .A4(\ram[11][143] ), .S0(n7337), .S1(n5560), .Y(n8303)
         );
  MUX41X1_HVT U9953 ( .A1(\ram[4][143] ), .A3(\ram[6][143] ), .A2(
        \ram[5][143] ), .A4(\ram[7][143] ), .S0(n7320), .S1(n7683), .Y(n8304)
         );
  MUX41X1_HVT U9954 ( .A1(\ram[0][143] ), .A3(\ram[2][143] ), .A2(
        \ram[1][143] ), .A4(\ram[3][143] ), .S0(n4980), .S1(n8875), .Y(n8305)
         );
  MUX41X1_HVT U9955 ( .A1(\ram[12][144] ), .A3(\ram[14][144] ), .A2(
        \ram[13][144] ), .A4(\ram[15][144] ), .S0(n5014), .S1(n6385), .Y(n8306) );
  MUX41X1_HVT U9956 ( .A1(\ram[8][144] ), .A3(\ram[10][144] ), .A2(
        \ram[9][144] ), .A4(\ram[11][144] ), .S0(n5509), .S1(n7577), .Y(n8307)
         );
  MUX41X1_HVT U9957 ( .A1(\ram[4][144] ), .A3(\ram[6][144] ), .A2(
        \ram[5][144] ), .A4(\ram[7][144] ), .S0(n6652), .S1(n6115), .Y(n8308)
         );
  MUX41X1_HVT U9958 ( .A1(\ram[0][145] ), .A3(\ram[2][145] ), .A2(
        \ram[1][145] ), .A4(\ram[3][145] ), .S0(n5865), .S1(n7329), .Y(n8312)
         );
  MUX41X1_HVT U9959 ( .A1(\ram[12][146] ), .A3(\ram[14][146] ), .A2(
        \ram[13][146] ), .A4(\ram[15][146] ), .S0(n8824), .S1(n7683), .Y(n8313) );
  MUX41X1_HVT U9960 ( .A1(\ram[8][146] ), .A3(\ram[10][146] ), .A2(
        \ram[9][146] ), .A4(\ram[11][146] ), .S0(n4973), .S1(n5760), .Y(n8314)
         );
  MUX41X1_HVT U9961 ( .A1(\ram[0][146] ), .A3(\ram[2][146] ), .A2(
        \ram[1][146] ), .A4(\ram[3][146] ), .S0(n8846), .S1(n7342), .Y(n8316)
         );
  MUX41X1_HVT U9962 ( .A1(\ram[8][147] ), .A3(\ram[10][147] ), .A2(
        \ram[9][147] ), .A4(\ram[11][147] ), .S0(n4794), .S1(n6409), .Y(n8318)
         );
  MUX41X1_HVT U9963 ( .A1(\ram[4][148] ), .A3(\ram[6][148] ), .A2(
        \ram[5][148] ), .A4(\ram[7][148] ), .S0(n5948), .S1(n7569), .Y(n8323)
         );
  MUX41X1_HVT U9964 ( .A1(\ram[12][149] ), .A3(\ram[14][149] ), .A2(
        \ram[13][149] ), .A4(\ram[15][149] ), .S0(n8840), .S1(n5366), .Y(n8325) );
  MUX41X1_HVT U9965 ( .A1(\ram[8][149] ), .A3(\ram[10][149] ), .A2(
        \ram[9][149] ), .A4(\ram[11][149] ), .S0(n8796), .S1(n5366), .Y(n8326)
         );
  MUX41X1_HVT U9966 ( .A1(\ram[4][149] ), .A3(\ram[6][149] ), .A2(
        \ram[5][149] ), .A4(\ram[7][149] ), .S0(n6007), .S1(n8887), .Y(n8327)
         );
  MUX41X1_HVT U9967 ( .A1(\ram[0][149] ), .A3(\ram[2][149] ), .A2(
        \ram[1][149] ), .A4(\ram[3][149] ), .S0(n8808), .S1(n8887), .Y(n8328)
         );
  MUX41X1_HVT U9968 ( .A1(\ram[8][151] ), .A3(\ram[10][151] ), .A2(
        \ram[9][151] ), .A4(\ram[11][151] ), .S0(n6406), .S1(n8903), .Y(n8334)
         );
  MUX41X1_HVT U9969 ( .A1(\ram[8][152] ), .A3(\ram[10][152] ), .A2(
        \ram[9][152] ), .A4(\ram[11][152] ), .S0(n5978), .S1(n5974), .Y(n8338)
         );
  MUX41X1_HVT U9970 ( .A1(\ram[0][153] ), .A3(\ram[2][153] ), .A2(
        \ram[1][153] ), .A4(\ram[3][153] ), .S0(n6406), .S1(n1651), .Y(n8344)
         );
  MUX41X1_HVT U9971 ( .A1(\ram[12][154] ), .A3(\ram[14][154] ), .A2(
        \ram[13][154] ), .A4(\ram[15][154] ), .S0(n4991), .S1(n5303), .Y(n8345) );
  MUX41X1_HVT U9972 ( .A1(\ram[8][154] ), .A3(\ram[10][154] ), .A2(
        \ram[9][154] ), .A4(\ram[11][154] ), .S0(n6020), .S1(n7700), .Y(n8346)
         );
  MUX41X1_HVT U9973 ( .A1(\ram[12][155] ), .A3(\ram[14][155] ), .A2(
        \ram[13][155] ), .A4(\ram[15][155] ), .S0(n8814), .S1(n5149), .Y(n8349) );
  MUX41X1_HVT U9974 ( .A1(\ram[4][155] ), .A3(\ram[6][155] ), .A2(
        \ram[5][155] ), .A4(\ram[7][155] ), .S0(n5231), .S1(n7700), .Y(n8351)
         );
  MUX41X1_HVT U9975 ( .A1(\ram[4][156] ), .A3(\ram[6][156] ), .A2(
        \ram[5][156] ), .A4(\ram[7][156] ), .S0(n4837), .S1(n6395), .Y(n8355)
         );
  MUX41X1_HVT U9976 ( .A1(\ram[12][157] ), .A3(\ram[14][157] ), .A2(
        \ram[13][157] ), .A4(\ram[15][157] ), .S0(n7320), .S1(n8873), .Y(n8357) );
  MUX41X1_HVT U9977 ( .A1(\ram[8][157] ), .A3(\ram[10][157] ), .A2(
        \ram[9][157] ), .A4(\ram[11][157] ), .S0(n8828), .S1(n7341), .Y(n8358)
         );
  MUX41X1_HVT U9978 ( .A1(\ram[0][157] ), .A3(\ram[2][157] ), .A2(
        \ram[1][157] ), .A4(\ram[3][157] ), .S0(n4949), .S1(n7577), .Y(n8360)
         );
  MUX41X1_HVT U9979 ( .A1(\ram[4][159] ), .A3(\ram[6][159] ), .A2(
        \ram[5][159] ), .A4(\ram[7][159] ), .S0(n6183), .S1(n5139), .Y(n8367)
         );
  MUX41X1_HVT U9980 ( .A1(\ram[4][160] ), .A3(\ram[6][160] ), .A2(
        \ram[5][160] ), .A4(\ram[7][160] ), .S0(n6183), .S1(n7706), .Y(n8371)
         );
  MUX41X1_HVT U9981 ( .A1(\ram[0][162] ), .A3(\ram[2][162] ), .A2(
        \ram[1][162] ), .A4(\ram[3][162] ), .S0(n8842), .S1(n7689), .Y(n8380)
         );
  MUX41X1_HVT U9982 ( .A1(\ram[8][163] ), .A3(\ram[10][163] ), .A2(
        \ram[9][163] ), .A4(\ram[11][163] ), .S0(n7145), .S1(n5650), .Y(n8382)
         );
  MUX41X1_HVT U9983 ( .A1(\ram[12][164] ), .A3(\ram[14][164] ), .A2(
        \ram[13][164] ), .A4(\ram[15][164] ), .S0(n8844), .S1(n7342), .Y(n8385) );
  MUX41X1_HVT U9984 ( .A1(\ram[0][164] ), .A3(\ram[2][164] ), .A2(
        \ram[1][164] ), .A4(\ram[3][164] ), .S0(n8846), .S1(n8864), .Y(n8388)
         );
  MUX41X1_HVT U9985 ( .A1(\ram[4][167] ), .A3(\ram[6][167] ), .A2(
        \ram[5][167] ), .A4(\ram[7][167] ), .S0(n8819), .S1(n8906), .Y(n8399)
         );
  MUX41X1_HVT U9986 ( .A1(\ram[0][167] ), .A3(\ram[2][167] ), .A2(
        \ram[1][167] ), .A4(\ram[3][167] ), .S0(n8811), .S1(n5150), .Y(n8400)
         );
  MUX41X1_HVT U9987 ( .A1(\ram[12][168] ), .A3(\ram[14][168] ), .A2(
        \ram[13][168] ), .A4(\ram[15][168] ), .S0(n5978), .S1(n5054), .Y(n8401) );
  MUX41X1_HVT U9988 ( .A1(\ram[8][168] ), .A3(\ram[10][168] ), .A2(
        \ram[9][168] ), .A4(\ram[11][168] ), .S0(n8824), .S1(n8907), .Y(n8402)
         );
  MUX41X1_HVT U9989 ( .A1(\ram[4][168] ), .A3(\ram[6][168] ), .A2(
        \ram[5][168] ), .A4(\ram[7][168] ), .S0(n5940), .S1(n8909), .Y(n8403)
         );
  MUX41X1_HVT U9990 ( .A1(\ram[0][168] ), .A3(\ram[2][168] ), .A2(
        \ram[1][168] ), .A4(\ram[3][168] ), .S0(n8838), .S1(n5441), .Y(n8404)
         );
  MUX41X1_HVT U9991 ( .A1(\ram[8][169] ), .A3(\ram[10][169] ), .A2(
        \ram[9][169] ), .A4(\ram[11][169] ), .S0(n8792), .S1(n5649), .Y(n8406)
         );
  MUX41X1_HVT U9992 ( .A1(\ram[4][169] ), .A3(\ram[6][169] ), .A2(
        \ram[5][169] ), .A4(\ram[7][169] ), .S0(n6028), .S1(n7704), .Y(n8407)
         );
  MUX41X1_HVT U9993 ( .A1(\ram[12][170] ), .A3(\ram[14][170] ), .A2(
        \ram[13][170] ), .A4(\ram[15][170] ), .S0(n8793), .S1(n5753), .Y(n8409) );
  MUX41X1_HVT U9994 ( .A1(\ram[4][170] ), .A3(\ram[6][170] ), .A2(
        \ram[5][170] ), .A4(\ram[7][170] ), .S0(n5132), .S1(n5777), .Y(n8411)
         );
  MUX41X1_HVT U9995 ( .A1(\ram[0][170] ), .A3(\ram[2][170] ), .A2(
        \ram[1][170] ), .A4(\ram[3][170] ), .S0(n6008), .S1(n5539), .Y(n8412)
         );
  MUX41X1_HVT U9996 ( .A1(\ram[0][171] ), .A3(\ram[2][171] ), .A2(
        \ram[1][171] ), .A4(\ram[3][171] ), .S0(n6009), .S1(n5447), .Y(n8416)
         );
  MUX41X1_HVT U9997 ( .A1(\ram[4][172] ), .A3(\ram[6][172] ), .A2(
        \ram[5][172] ), .A4(\ram[7][172] ), .S0(n5231), .S1(n5956), .Y(n8419)
         );
  MUX41X1_HVT U9998 ( .A1(\ram[0][172] ), .A3(\ram[2][172] ), .A2(
        \ram[1][172] ), .A4(\ram[3][172] ), .S0(n5923), .S1(n5989), .Y(n8420)
         );
  MUX41X1_HVT U9999 ( .A1(\ram[4][173] ), .A3(\ram[6][173] ), .A2(
        \ram[5][173] ), .A4(\ram[7][173] ), .S0(n4991), .S1(n5989), .Y(n8423)
         );
  MUX41X1_HVT U10000 ( .A1(\ram[4][174] ), .A3(\ram[6][174] ), .A2(
        \ram[5][174] ), .A4(\ram[7][174] ), .S0(n5923), .S1(n8893), .Y(n8427)
         );
  MUX41X1_HVT U10001 ( .A1(\ram[12][175] ), .A3(\ram[14][175] ), .A2(
        \ram[13][175] ), .A4(\ram[15][175] ), .S0(n8807), .S1(n5591), .Y(n8429) );
  MUX41X1_HVT U10002 ( .A1(\ram[8][175] ), .A3(\ram[10][175] ), .A2(
        \ram[9][175] ), .A4(\ram[11][175] ), .S0(n5004), .S1(n8855), .Y(n8430)
         );
  MUX41X1_HVT U10003 ( .A1(\ram[4][176] ), .A3(\ram[6][176] ), .A2(
        \ram[5][176] ), .A4(\ram[7][176] ), .S0(n5004), .S1(n8855), .Y(n8435)
         );
  MUX41X1_HVT U10004 ( .A1(\ram[0][176] ), .A3(\ram[2][176] ), .A2(
        \ram[1][176] ), .A4(\ram[3][176] ), .S0(n6413), .S1(n8855), .Y(n8436)
         );
  MUX41X1_HVT U10005 ( .A1(n8436), .A3(n8434), .A2(n8435), .A4(n8433), .S0(
        n6756), .S1(n7332), .Y(q[176]) );
  MUX41X1_HVT U10006 ( .A1(\ram[4][177] ), .A3(\ram[6][177] ), .A2(
        \ram[5][177] ), .A4(\ram[7][177] ), .S0(n8810), .S1(n8877), .Y(n8439)
         );
  MUX41X1_HVT U10007 ( .A1(\ram[12][178] ), .A3(\ram[14][178] ), .A2(
        \ram[13][178] ), .A4(\ram[15][178] ), .S0(n7336), .S1(n8853), .Y(n8441) );
  MUX41X1_HVT U10008 ( .A1(\ram[0][178] ), .A3(\ram[2][178] ), .A2(
        \ram[1][178] ), .A4(\ram[3][178] ), .S0(n5948), .S1(n8905), .Y(n8444)
         );
  MUX41X1_HVT U10009 ( .A1(\ram[12][179] ), .A3(\ram[14][179] ), .A2(
        \ram[13][179] ), .A4(\ram[15][179] ), .S0(n5890), .S1(n5150), .Y(n8445) );
  MUX41X1_HVT U10010 ( .A1(\ram[4][179] ), .A3(\ram[6][179] ), .A2(
        \ram[5][179] ), .A4(\ram[7][179] ), .S0(n8832), .S1(n5974), .Y(n8447)
         );
  MUX41X1_HVT U10011 ( .A1(\ram[0][179] ), .A3(\ram[2][179] ), .A2(
        \ram[1][179] ), .A4(\ram[3][179] ), .S0(n5793), .S1(n7563), .Y(n8448)
         );
  MUX41X1_HVT U10012 ( .A1(n8448), .A3(n8446), .A2(n8447), .A4(n8445), .S0(
        n7300), .S1(n7715), .Y(q[179]) );
  MUX41X1_HVT U10013 ( .A1(\ram[12][180] ), .A3(\ram[14][180] ), .A2(
        \ram[13][180] ), .A4(\ram[15][180] ), .S0(n8799), .S1(n5135), .Y(n8449) );
  MUX41X1_HVT U10014 ( .A1(\ram[8][180] ), .A3(\ram[10][180] ), .A2(
        \ram[9][180] ), .A4(\ram[11][180] ), .S0(n7336), .S1(n6409), .Y(n8450)
         );
  MUX41X1_HVT U10015 ( .A1(\ram[4][180] ), .A3(\ram[6][180] ), .A2(
        \ram[5][180] ), .A4(\ram[7][180] ), .S0(n8841), .S1(n6409), .Y(n8451)
         );
  MUX41X1_HVT U10016 ( .A1(\ram[12][181] ), .A3(\ram[14][181] ), .A2(
        \ram[13][181] ), .A4(\ram[15][181] ), .S0(n5923), .S1(n5971), .Y(n8453) );
  MUX41X1_HVT U10017 ( .A1(\ram[0][181] ), .A3(\ram[2][181] ), .A2(
        \ram[1][181] ), .A4(\ram[3][181] ), .S0(n5734), .S1(n8903), .Y(n8456)
         );
  MUX41X1_HVT U10018 ( .A1(\ram[8][182] ), .A3(\ram[10][182] ), .A2(
        \ram[9][182] ), .A4(\ram[11][182] ), .S0(n5004), .S1(n5148), .Y(n8458)
         );
  MUX41X1_HVT U10019 ( .A1(\ram[4][182] ), .A3(\ram[6][182] ), .A2(
        \ram[5][182] ), .A4(\ram[7][182] ), .S0(n8792), .S1(n8893), .Y(n8459)
         );
  MUX41X1_HVT U10020 ( .A1(\ram[0][183] ), .A3(\ram[2][183] ), .A2(
        \ram[1][183] ), .A4(\ram[3][183] ), .S0(n7554), .S1(n5557), .Y(n8464)
         );
  MUX41X1_HVT U10021 ( .A1(\ram[4][184] ), .A3(\ram[6][184] ), .A2(
        \ram[5][184] ), .A4(\ram[7][184] ), .S0(n6183), .S1(n8872), .Y(n8467)
         );
  MUX41X1_HVT U10022 ( .A1(\ram[0][184] ), .A3(\ram[2][184] ), .A2(
        \ram[1][184] ), .A4(\ram[3][184] ), .S0(n6009), .S1(n7707), .Y(n8468)
         );
  MUX41X1_HVT U10023 ( .A1(\ram[4][185] ), .A3(\ram[6][185] ), .A2(
        \ram[5][185] ), .A4(\ram[7][185] ), .S0(n6024), .S1(n8907), .Y(n8471)
         );
  MUX41X1_HVT U10024 ( .A1(\ram[4][186] ), .A3(\ram[6][186] ), .A2(
        \ram[5][186] ), .A4(\ram[7][186] ), .S0(n8795), .S1(n8868), .Y(n8475)
         );
  MUX41X1_HVT U10025 ( .A1(\ram[0][186] ), .A3(\ram[2][186] ), .A2(
        \ram[1][186] ), .A4(\ram[3][186] ), .S0(n7550), .S1(n8896), .Y(n8476)
         );
  MUX41X1_HVT U10026 ( .A1(\ram[0][187] ), .A3(\ram[2][187] ), .A2(
        \ram[1][187] ), .A4(\ram[3][187] ), .S0(n8795), .S1(n8868), .Y(n8480)
         );
  MUX41X1_HVT U10027 ( .A1(\ram[12][188] ), .A3(\ram[14][188] ), .A2(
        \ram[13][188] ), .A4(\ram[15][188] ), .S0(n5997), .S1(n4174), .Y(n8481) );
  MUX41X1_HVT U10028 ( .A1(\ram[8][188] ), .A3(\ram[10][188] ), .A2(
        \ram[9][188] ), .A4(\ram[11][188] ), .S0(n4975), .S1(n5535), .Y(n8482)
         );
  MUX41X1_HVT U10029 ( .A1(\ram[12][189] ), .A3(\ram[14][189] ), .A2(
        \ram[13][189] ), .A4(\ram[15][189] ), .S0(n5499), .S1(n4982), .Y(n8485) );
  MUX41X1_HVT U10030 ( .A1(\ram[4][189] ), .A3(\ram[6][189] ), .A2(
        \ram[5][189] ), .A4(\ram[7][189] ), .S0(n6017), .S1(n7581), .Y(n8487)
         );
  MUX41X1_HVT U10031 ( .A1(\ram[0][189] ), .A3(\ram[2][189] ), .A2(
        \ram[1][189] ), .A4(\ram[3][189] ), .S0(n4794), .S1(n7704), .Y(n8488)
         );
  MUX41X1_HVT U10032 ( .A1(\ram[4][190] ), .A3(\ram[6][190] ), .A2(
        \ram[5][190] ), .A4(\ram[7][190] ), .S0(n5751), .S1(n5875), .Y(n8491)
         );
  MUX41X1_HVT U10033 ( .A1(\ram[0][191] ), .A3(\ram[2][191] ), .A2(
        \ram[1][191] ), .A4(\ram[3][191] ), .S0(n6757), .S1(n6006), .Y(n8496)
         );
  MUX41X1_HVT U10034 ( .A1(\ram[8][192] ), .A3(\ram[10][192] ), .A2(
        \ram[9][192] ), .A4(\ram[11][192] ), .S0(n8805), .S1(n7691), .Y(n8498)
         );
  MUX41X1_HVT U10035 ( .A1(\ram[0][193] ), .A3(\ram[2][193] ), .A2(
        \ram[1][193] ), .A4(\ram[3][193] ), .S0(n5612), .S1(n8909), .Y(n8504)
         );
  MUX41X1_HVT U10036 ( .A1(\ram[0][195] ), .A3(\ram[2][195] ), .A2(
        \ram[1][195] ), .A4(\ram[3][195] ), .S0(n8795), .S1(n7341), .Y(n8512)
         );
  MUX41X1_HVT U10037 ( .A1(\ram[12][196] ), .A3(\ram[14][196] ), .A2(
        \ram[13][196] ), .A4(\ram[15][196] ), .S0(n8816), .S1(n7560), .Y(n8513) );
  MUX41X1_HVT U10038 ( .A1(\ram[4][196] ), .A3(\ram[6][196] ), .A2(
        \ram[5][196] ), .A4(\ram[7][196] ), .S0(n5945), .S1(n5557), .Y(n8515)
         );
  MUX41X1_HVT U10039 ( .A1(\ram[4][197] ), .A3(\ram[6][197] ), .A2(
        \ram[5][197] ), .A4(\ram[7][197] ), .S0(n8805), .S1(n7665), .Y(n8519)
         );
  MUX41X1_HVT U10040 ( .A1(\ram[0][197] ), .A3(\ram[2][197] ), .A2(
        \ram[1][197] ), .A4(\ram[3][197] ), .S0(n5592), .S1(n5528), .Y(n8520)
         );
  MUX41X1_HVT U10041 ( .A1(\ram[12][198] ), .A3(\ram[14][198] ), .A2(
        \ram[13][198] ), .A4(\ram[15][198] ), .S0(n4837), .S1(n5528), .Y(n8521) );
  MUX41X1_HVT U10042 ( .A1(\ram[4][198] ), .A3(\ram[6][198] ), .A2(
        \ram[5][198] ), .A4(\ram[7][198] ), .S0(n4162), .S1(n7568), .Y(n8523)
         );
  MUX41X1_HVT U10043 ( .A1(\ram[12][199] ), .A3(\ram[14][199] ), .A2(
        \ram[13][199] ), .A4(\ram[15][199] ), .S0(n7145), .S1(n8853), .Y(n8525) );
  MUX41X1_HVT U10044 ( .A1(\ram[8][199] ), .A3(\ram[10][199] ), .A2(
        \ram[9][199] ), .A4(\ram[11][199] ), .S0(n7145), .S1(n8884), .Y(n8526)
         );
  MUX41X1_HVT U10045 ( .A1(\ram[0][199] ), .A3(\ram[2][199] ), .A2(
        \ram[1][199] ), .A4(\ram[3][199] ), .S0(n7552), .S1(n5463), .Y(n8528)
         );
  MUX41X1_HVT U10046 ( .A1(\ram[8][200] ), .A3(\ram[10][200] ), .A2(
        \ram[9][200] ), .A4(\ram[11][200] ), .S0(n5126), .S1(n5875), .Y(n8530)
         );
  MUX41X1_HVT U10047 ( .A1(\ram[4][200] ), .A3(\ram[6][200] ), .A2(
        \ram[5][200] ), .A4(\ram[7][200] ), .S0(n4162), .S1(n7578), .Y(n8531)
         );
  MUX41X1_HVT U10048 ( .A1(\ram[0][200] ), .A3(\ram[2][200] ), .A2(
        \ram[1][200] ), .A4(\ram[3][200] ), .S0(n7552), .S1(n8890), .Y(n8532)
         );
  MUX41X1_HVT U10049 ( .A1(\ram[4][201] ), .A3(\ram[6][201] ), .A2(
        \ram[5][201] ), .A4(\ram[7][201] ), .S0(n5612), .S1(n8858), .Y(n8535)
         );
  MUX41X1_HVT U10050 ( .A1(\ram[8][202] ), .A3(\ram[10][202] ), .A2(
        \ram[9][202] ), .A4(\ram[11][202] ), .S0(n5559), .S1(n5554), .Y(n8538)
         );
  MUX41X1_HVT U10051 ( .A1(\ram[4][202] ), .A3(\ram[6][202] ), .A2(
        \ram[5][202] ), .A4(\ram[7][202] ), .S0(n5559), .S1(n4982), .Y(n8539)
         );
  MUX41X1_HVT U10052 ( .A1(\ram[0][202] ), .A3(\ram[2][202] ), .A2(
        \ram[1][202] ), .A4(\ram[3][202] ), .S0(n6650), .S1(n7691), .Y(n8540)
         );
  MUX41X1_HVT U10053 ( .A1(\ram[4][204] ), .A3(\ram[6][204] ), .A2(
        \ram[5][204] ), .A4(\ram[7][204] ), .S0(n5132), .S1(n8880), .Y(n8547)
         );
  MUX41X1_HVT U10054 ( .A1(\ram[0][204] ), .A3(\ram[2][204] ), .A2(
        \ram[1][204] ), .A4(\ram[3][204] ), .S0(n5000), .S1(n7686), .Y(n8548)
         );
  MUX41X1_HVT U10055 ( .A1(\ram[12][205] ), .A3(\ram[14][205] ), .A2(
        \ram[13][205] ), .A4(\ram[15][205] ), .S0(n8837), .S1(n6966), .Y(n8549) );
  MUX41X1_HVT U10056 ( .A1(\ram[4][205] ), .A3(\ram[6][205] ), .A2(
        \ram[5][205] ), .A4(\ram[7][205] ), .S0(n5957), .S1(n5728), .Y(n8551)
         );
  MUX41X1_HVT U10057 ( .A1(\ram[12][206] ), .A3(\ram[14][206] ), .A2(
        \ram[13][206] ), .A4(\ram[15][206] ), .S0(n4918), .S1(n6386), .Y(n8553) );
  MUX41X1_HVT U10058 ( .A1(\ram[8][206] ), .A3(\ram[10][206] ), .A2(
        \ram[9][206] ), .A4(\ram[11][206] ), .S0(n4949), .S1(n5441), .Y(n8554)
         );
  MUX41X1_HVT U10059 ( .A1(\ram[0][206] ), .A3(\ram[2][206] ), .A2(
        \ram[1][206] ), .A4(\ram[3][206] ), .S0(n5310), .S1(n5650), .Y(n8556)
         );
  MUX41X1_HVT U10060 ( .A1(\ram[12][207] ), .A3(\ram[14][207] ), .A2(
        \ram[13][207] ), .A4(\ram[15][207] ), .S0(n8794), .S1(n4820), .Y(n8557) );
  MUX41X1_HVT U10061 ( .A1(\ram[8][207] ), .A3(\ram[10][207] ), .A2(
        \ram[9][207] ), .A4(\ram[11][207] ), .S0(n8802), .S1(n7696), .Y(n8558)
         );
  MUX41X1_HVT U10062 ( .A1(\ram[12][208] ), .A3(\ram[14][208] ), .A2(
        \ram[13][208] ), .A4(\ram[15][208] ), .S0(n8835), .S1(n4992), .Y(n8561) );
  MUX41X1_HVT U10063 ( .A1(\ram[8][208] ), .A3(\ram[10][208] ), .A2(
        \ram[9][208] ), .A4(\ram[11][208] ), .S0(n5946), .S1(n8870), .Y(n8562)
         );
  MUX41X1_HVT U10064 ( .A1(\ram[4][208] ), .A3(\ram[6][208] ), .A2(
        \ram[5][208] ), .A4(\ram[7][208] ), .S0(n5504), .S1(n5554), .Y(n8563)
         );
  MUX41X1_HVT U10065 ( .A1(\ram[0][208] ), .A3(\ram[2][208] ), .A2(
        \ram[1][208] ), .A4(\ram[3][208] ), .S0(n8849), .S1(n8884), .Y(n8564)
         );
  MUX41X1_HVT U10066 ( .A1(\ram[12][210] ), .A3(\ram[14][210] ), .A2(
        \ram[13][210] ), .A4(\ram[15][210] ), .S0(n4991), .S1(n6763), .Y(n8569) );
  MUX41X1_HVT U10067 ( .A1(\ram[8][210] ), .A3(\ram[10][210] ), .A2(
        \ram[9][210] ), .A4(\ram[11][210] ), .S0(n8802), .S1(n8870), .Y(n8570)
         );
  MUX41X1_HVT U10068 ( .A1(\ram[4][210] ), .A3(\ram[6][210] ), .A2(
        \ram[5][210] ), .A4(\ram[7][210] ), .S0(n5932), .S1(n8864), .Y(n8571)
         );
  MUX41X1_HVT U10069 ( .A1(\ram[0][210] ), .A3(\ram[2][210] ), .A2(
        \ram[1][210] ), .A4(\ram[3][210] ), .S0(n7083), .S1(n7575), .Y(n8572)
         );
  MUX41X1_HVT U10070 ( .A1(\ram[8][211] ), .A3(\ram[10][211] ), .A2(
        \ram[9][211] ), .A4(\ram[11][211] ), .S0(n7083), .S1(n5446), .Y(n8574)
         );
  MUX41X1_HVT U10071 ( .A1(\ram[4][211] ), .A3(\ram[6][211] ), .A2(
        \ram[5][211] ), .A4(\ram[7][211] ), .S0(n8800), .S1(n4189), .Y(n8575)
         );
  MUX41X1_HVT U10072 ( .A1(\ram[8][212] ), .A3(\ram[10][212] ), .A2(
        \ram[9][212] ), .A4(\ram[11][212] ), .S0(n8815), .S1(n6743), .Y(n8578)
         );
  MUX41X1_HVT U10073 ( .A1(\ram[0][212] ), .A3(\ram[2][212] ), .A2(
        \ram[1][212] ), .A4(\ram[3][212] ), .S0(n7083), .S1(n7341), .Y(n8580)
         );
  MUX41X1_HVT U10074 ( .A1(\ram[8][213] ), .A3(\ram[10][213] ), .A2(
        \ram[9][213] ), .A4(\ram[11][213] ), .S0(n1078), .S1(n7704), .Y(n8582)
         );
  MUX41X1_HVT U10075 ( .A1(\ram[4][213] ), .A3(\ram[6][213] ), .A2(
        \ram[5][213] ), .A4(\ram[7][213] ), .S0(n1078), .S1(n5989), .Y(n8583)
         );
  MUX41X1_HVT U10076 ( .A1(\ram[4][214] ), .A3(\ram[6][214] ), .A2(
        \ram[5][214] ), .A4(\ram[7][214] ), .S0(n7344), .S1(n8856), .Y(n8587)
         );
  MUX41X1_HVT U10077 ( .A1(\ram[0][214] ), .A3(\ram[2][214] ), .A2(
        \ram[1][214] ), .A4(\ram[3][214] ), .S0(n7344), .S1(n7701), .Y(n8588)
         );
  MUX41X1_HVT U10078 ( .A1(\ram[4][215] ), .A3(\ram[6][215] ), .A2(
        \ram[5][215] ), .A4(\ram[7][215] ), .S0(n7344), .S1(n4166), .Y(n8591)
         );
  MUX41X1_HVT U10079 ( .A1(\ram[0][215] ), .A3(\ram[2][215] ), .A2(
        \ram[1][215] ), .A4(\ram[3][215] ), .S0(n1078), .S1(n8879), .Y(n8592)
         );
  MUX41X1_HVT U10080 ( .A1(n8592), .A3(n8590), .A2(n8591), .A4(n8589), .S0(
        n5867), .S1(n8767), .Y(q[215]) );
  MUX41X1_HVT U10081 ( .A1(\ram[0][216] ), .A3(\ram[2][216] ), .A2(
        \ram[1][216] ), .A4(\ram[3][216] ), .S0(n5577), .S1(n5615), .Y(n8596)
         );
  MUX41X1_HVT U10082 ( .A1(n8596), .A3(n8594), .A2(n8595), .A4(n8593), .S0(
        n8758), .S1(n7715), .Y(q[216]) );
  MUX41X1_HVT U10083 ( .A1(\ram[12][217] ), .A3(\ram[14][217] ), .A2(
        \ram[13][217] ), .A4(\ram[15][217] ), .S0(n7083), .S1(n8860), .Y(n8597) );
  MUX41X1_HVT U10084 ( .A1(\ram[12][218] ), .A3(\ram[14][218] ), .A2(
        \ram[13][218] ), .A4(\ram[15][218] ), .S0(n7141), .S1(n8902), .Y(n8601) );
  MUX41X1_HVT U10085 ( .A1(\ram[8][219] ), .A3(\ram[10][219] ), .A2(
        \ram[9][219] ), .A4(\ram[11][219] ), .S0(n4184), .S1(n7693), .Y(n8606)
         );
  MUX41X1_HVT U10086 ( .A1(\ram[4][219] ), .A3(\ram[6][219] ), .A2(
        \ram[5][219] ), .A4(\ram[7][219] ), .S0(n8799), .S1(n8900), .Y(n8607)
         );
  MUX41X1_HVT U10087 ( .A1(\ram[0][219] ), .A3(\ram[2][219] ), .A2(
        \ram[1][219] ), .A4(\ram[3][219] ), .S0(n4184), .S1(n6640), .Y(n8608)
         );
  MUX41X1_HVT U10088 ( .A1(\ram[4][220] ), .A3(\ram[6][220] ), .A2(
        \ram[5][220] ), .A4(\ram[7][220] ), .S0(n4985), .S1(n5470), .Y(n8611)
         );
  MUX41X1_HVT U10089 ( .A1(n8612), .A3(n8610), .A2(n8611), .A4(n8609), .S0(
        n8758), .S1(n8768), .Y(q[220]) );
  MUX41X1_HVT U10090 ( .A1(\ram[0][221] ), .A3(\ram[2][221] ), .A2(
        \ram[1][221] ), .A4(\ram[3][221] ), .S0(n8799), .S1(n8901), .Y(n8616)
         );
  MUX41X1_HVT U10091 ( .A1(\ram[4][222] ), .A3(\ram[6][222] ), .A2(
        \ram[5][222] ), .A4(\ram[7][222] ), .S0(n4990), .S1(n5071), .Y(n8619)
         );
  MUX41X1_HVT U10092 ( .A1(\ram[4][223] ), .A3(\ram[6][223] ), .A2(
        \ram[5][223] ), .A4(\ram[7][223] ), .S0(n8803), .S1(n5649), .Y(n8623)
         );
  MUX41X1_HVT U10093 ( .A1(\ram[0][223] ), .A3(\ram[2][223] ), .A2(
        \ram[1][223] ), .A4(\ram[3][223] ), .S0(n8798), .S1(n5795), .Y(n8624)
         );
  MUX41X1_HVT U10094 ( .A1(n8624), .A3(n8622), .A2(n8623), .A4(n8621), .S0(
        n8758), .S1(n5291), .Y(q[223]) );
  MUX41X1_HVT U10095 ( .A1(\ram[12][224] ), .A3(\ram[14][224] ), .A2(
        \ram[13][224] ), .A4(\ram[15][224] ), .S0(n8796), .S1(n8861), .Y(n8625) );
  MUX41X1_HVT U10096 ( .A1(\ram[8][224] ), .A3(\ram[10][224] ), .A2(
        \ram[9][224] ), .A4(\ram[11][224] ), .S0(n5854), .S1(n7575), .Y(n8626)
         );
  MUX41X1_HVT U10097 ( .A1(\ram[4][224] ), .A3(\ram[6][224] ), .A2(
        \ram[5][224] ), .A4(\ram[7][224] ), .S0(n6413), .S1(n5593), .Y(n8627)
         );
  MUX41X1_HVT U10098 ( .A1(\ram[4][225] ), .A3(\ram[6][225] ), .A2(
        \ram[5][225] ), .A4(\ram[7][225] ), .S0(n5866), .S1(n5921), .Y(n8631)
         );
  MUX41X1_HVT U10099 ( .A1(\ram[4][226] ), .A3(\ram[6][226] ), .A2(
        \ram[5][226] ), .A4(\ram[7][226] ), .S0(n8850), .S1(n7686), .Y(n8635)
         );
  MUX41X1_HVT U10100 ( .A1(\ram[8][227] ), .A3(\ram[10][227] ), .A2(
        \ram[9][227] ), .A4(\ram[11][227] ), .S0(n5353), .S1(n8865), .Y(n8638)
         );
  MUX41X1_HVT U10101 ( .A1(\ram[0][227] ), .A3(\ram[2][227] ), .A2(
        \ram[1][227] ), .A4(\ram[3][227] ), .S0(n5569), .S1(n1023), .Y(n8640)
         );
  MUX41X1_HVT U10102 ( .A1(\ram[4][228] ), .A3(\ram[6][228] ), .A2(
        \ram[5][228] ), .A4(\ram[7][228] ), .S0(n5499), .S1(n8872), .Y(n8643)
         );
  MUX41X1_HVT U10103 ( .A1(\ram[0][228] ), .A3(\ram[2][228] ), .A2(
        \ram[1][228] ), .A4(\ram[3][228] ), .S0(n5854), .S1(n8874), .Y(n8644)
         );
  MUX41X1_HVT U10104 ( .A1(\ram[8][229] ), .A3(\ram[10][229] ), .A2(
        \ram[9][229] ), .A4(\ram[11][229] ), .S0(n5892), .S1(n5629), .Y(n8646)
         );
  MUX41X1_HVT U10105 ( .A1(\ram[4][230] ), .A3(\ram[6][230] ), .A2(
        \ram[5][230] ), .A4(\ram[7][230] ), .S0(n5945), .S1(n7707), .Y(n8651)
         );
  MUX41X1_HVT U10106 ( .A1(\ram[0][230] ), .A3(\ram[2][230] ), .A2(
        \ram[1][230] ), .A4(\ram[3][230] ), .S0(n8841), .S1(n6127), .Y(n8652)
         );
  MUX41X1_HVT U10107 ( .A1(\ram[4][232] ), .A3(\ram[6][232] ), .A2(
        \ram[5][232] ), .A4(\ram[7][232] ), .S0(n8795), .S1(n8859), .Y(n8659)
         );
  MUX41X1_HVT U10108 ( .A1(\ram[4][233] ), .A3(\ram[6][233] ), .A2(
        \ram[5][233] ), .A4(\ram[7][233] ), .S0(n6642), .S1(n4994), .Y(n8662)
         );
  MUX41X1_HVT U10109 ( .A1(\ram[0][234] ), .A3(\ram[2][234] ), .A2(
        \ram[1][234] ), .A4(\ram[3][234] ), .S0(n8849), .S1(n6966), .Y(n8666)
         );
  MUX41X1_HVT U10110 ( .A1(\ram[12][235] ), .A3(\ram[14][235] ), .A2(
        \ram[13][235] ), .A4(\ram[15][235] ), .S0(n7083), .S1(n7667), .Y(n8667) );
  MUX41X1_HVT U10111 ( .A1(\ram[8][235] ), .A3(\ram[10][235] ), .A2(
        \ram[9][235] ), .A4(\ram[11][235] ), .S0(n5564), .S1(n8857), .Y(n8668)
         );
  MUX41X1_HVT U10112 ( .A1(\ram[12][236] ), .A3(\ram[14][236] ), .A2(
        \ram[13][236] ), .A4(\ram[15][236] ), .S0(n5734), .S1(n5366), .Y(n8671) );
  MUX41X1_HVT U10113 ( .A1(\ram[4][237] ), .A3(\ram[6][237] ), .A2(
        \ram[5][237] ), .A4(\ram[7][237] ), .S0(n5569), .S1(n8909), .Y(n8677)
         );
  MUX41X1_HVT U10114 ( .A1(\ram[8][238] ), .A3(\ram[10][238] ), .A2(
        \ram[9][238] ), .A4(\ram[11][238] ), .S0(n8843), .S1(n5649), .Y(n8680)
         );
  MUX41X1_HVT U10115 ( .A1(\ram[4][238] ), .A3(\ram[6][238] ), .A2(
        \ram[5][238] ), .A4(\ram[7][238] ), .S0(n5612), .S1(n8857), .Y(n8681)
         );
  MUX41X1_HVT U10116 ( .A1(\ram[0][238] ), .A3(\ram[2][238] ), .A2(
        \ram[1][238] ), .A4(\ram[3][238] ), .S0(n7337), .S1(n7323), .Y(n8682)
         );
  MUX41X1_HVT U10117 ( .A1(\ram[8][239] ), .A3(\ram[10][239] ), .A2(
        \ram[9][239] ), .A4(\ram[11][239] ), .S0(n6005), .S1(n7679), .Y(n8684)
         );
  MUX41X1_HVT U10118 ( .A1(\ram[4][239] ), .A3(\ram[6][239] ), .A2(
        \ram[5][239] ), .A4(\ram[7][239] ), .S0(n6017), .S1(n6385), .Y(n8685)
         );
  MUX41X1_HVT U10119 ( .A1(\ram[0][239] ), .A3(\ram[2][239] ), .A2(
        \ram[1][239] ), .A4(\ram[3][239] ), .S0(n6653), .S1(n8865), .Y(n8686)
         );
  MUX41X1_HVT U10120 ( .A1(\ram[4][240] ), .A3(\ram[6][240] ), .A2(
        \ram[5][240] ), .A4(\ram[7][240] ), .S0(n8797), .S1(n7322), .Y(n8689)
         );
  MUX41X1_HVT U10121 ( .A1(\ram[0][240] ), .A3(\ram[2][240] ), .A2(
        \ram[1][240] ), .A4(\ram[3][240] ), .S0(n8793), .S1(n8879), .Y(n8690)
         );
  MUX41X1_HVT U10122 ( .A1(\ram[8][241] ), .A3(\ram[10][241] ), .A2(
        \ram[9][241] ), .A4(\ram[11][241] ), .S0(n6005), .S1(n8856), .Y(n8692)
         );
  MUX41X1_HVT U10123 ( .A1(\ram[4][242] ), .A3(\ram[6][242] ), .A2(
        \ram[5][242] ), .A4(\ram[7][242] ), .S0(n4918), .S1(n5582), .Y(n8697)
         );
  MUX41X1_HVT U10124 ( .A1(\ram[0][242] ), .A3(\ram[2][242] ), .A2(
        \ram[1][242] ), .A4(\ram[3][242] ), .S0(n6009), .S1(n7322), .Y(n8698)
         );
  MUX41X1_HVT U10125 ( .A1(\ram[8][243] ), .A3(\ram[10][243] ), .A2(
        \ram[9][243] ), .A4(\ram[11][243] ), .S0(n6653), .S1(n6382), .Y(n8700)
         );
  MUX41X1_HVT U10126 ( .A1(\ram[4][243] ), .A3(\ram[6][243] ), .A2(
        \ram[5][243] ), .A4(\ram[7][243] ), .S0(n7554), .S1(n8903), .Y(n8701)
         );
  MUX41X1_HVT U10127 ( .A1(\ram[4][244] ), .A3(\ram[6][244] ), .A2(
        \ram[5][244] ), .A4(\ram[7][244] ), .S0(n8816), .S1(n5974), .Y(n8705)
         );
  MUX41X1_HVT U10128 ( .A1(\ram[0][244] ), .A3(\ram[2][244] ), .A2(
        \ram[1][244] ), .A4(\ram[3][244] ), .S0(n8804), .S1(n5287), .Y(n8706)
         );
  MUX41X1_HVT U10129 ( .A1(\ram[4][245] ), .A3(\ram[6][245] ), .A2(
        \ram[5][245] ), .A4(\ram[7][245] ), .S0(n7324), .S1(n7342), .Y(n8709)
         );
  MUX41X1_HVT U10130 ( .A1(\ram[12][246] ), .A3(\ram[14][246] ), .A2(
        \ram[13][246] ), .A4(\ram[15][246] ), .S0(n8823), .S1(n6253), .Y(n8711) );
  MUX41X1_HVT U10131 ( .A1(\ram[4][246] ), .A3(\ram[6][246] ), .A2(
        \ram[5][246] ), .A4(\ram[7][246] ), .S0(n8825), .S1(n8885), .Y(n8713)
         );
  MUX41X1_HVT U10132 ( .A1(\ram[8][248] ), .A3(\ram[10][248] ), .A2(
        \ram[9][248] ), .A4(\ram[11][248] ), .S0(n4981), .S1(n5964), .Y(n8720)
         );
  MUX41X1_HVT U10133 ( .A1(n8722), .A3(n8720), .A2(n8721), .A4(n8719), .S0(
        n8756), .S1(n8775), .Y(q[248]) );
  MUX41X1_HVT U10134 ( .A1(\ram[8][250] ), .A3(\ram[10][250] ), .A2(
        \ram[9][250] ), .A4(\ram[11][250] ), .S0(n5612), .S1(n5053), .Y(n8728)
         );
  MUX41X1_HVT U10135 ( .A1(\ram[8][252] ), .A3(\ram[10][252] ), .A2(
        \ram[9][252] ), .A4(\ram[11][252] ), .S0(n6005), .S1(n8856), .Y(n8736)
         );
  MUX41X1_HVT U10136 ( .A1(\ram[0][253] ), .A3(\ram[2][253] ), .A2(
        \ram[1][253] ), .A4(\ram[3][253] ), .S0(n5900), .S1(n5463), .Y(n8742)
         );
  MUX41X1_HVT U10137 ( .A1(\ram[4][254] ), .A3(\ram[6][254] ), .A2(
        \ram[5][254] ), .A4(\ram[7][254] ), .S0(n5900), .S1(n6394), .Y(n8745)
         );
  MUX41X1_HVT U10138 ( .A1(\ram[0][254] ), .A3(\ram[2][254] ), .A2(
        \ram[1][254] ), .A4(\ram[3][254] ), .S0(n4975), .S1(n5557), .Y(n8746)
         );
  MUX41X1_HVT U10139 ( .A1(\ram[8][255] ), .A3(\ram[10][255] ), .A2(
        \ram[9][255] ), .A4(\ram[11][255] ), .S0(n5900), .S1(n4189), .Y(n8748)
         );
  MUX41X1_HVT U10140 ( .A1(\ram[4][255] ), .A3(\ram[6][255] ), .A2(
        \ram[5][255] ), .A4(\ram[7][255] ), .S0(n8803), .S1(n8873), .Y(n8749)
         );
  MUX41X1_HVT U10141 ( .A1(\ram[0][255] ), .A3(\ram[2][255] ), .A2(
        \ram[1][255] ), .A4(\ram[3][255] ), .S0(n8840), .S1(n6382), .Y(n8750)
         );
  INVX0_HVT U10142 ( .A(n10124), .Y(n8910) );
  INVX0_HVT U10143 ( .A(n10124), .Y(n8911) );
  NBUFFX2_HVT U10144 ( .A(n8911), .Y(n8914) );
  NBUFFX2_HVT U10145 ( .A(n8910), .Y(n8915) );
  NBUFFX2_HVT U10146 ( .A(n8921), .Y(n8917) );
  NBUFFX2_HVT U10147 ( .A(n8916), .Y(n8918) );
  NBUFFX2_HVT U10148 ( .A(n8916), .Y(n8919) );
  NBUFFX2_HVT U10149 ( .A(n8916), .Y(n8920) );
  NBUFFX2_HVT U10150 ( .A(n8922), .Y(n8925) );
  NBUFFX2_HVT U10151 ( .A(n8922), .Y(n8926) );
  INVX0_HVT U10152 ( .A(n10122), .Y(n8927) );
  NBUFFX2_HVT U10153 ( .A(n8927), .Y(n8928) );
  NBUFFX2_HVT U10154 ( .A(n4513), .Y(n8929) );
  NBUFFX2_HVT U10155 ( .A(n8927), .Y(n8930) );
  NBUFFX2_HVT U10156 ( .A(n8932), .Y(n8931) );
  INVX0_HVT U10157 ( .A(n10122), .Y(n8932) );
  INVX0_HVT U10158 ( .A(n10122), .Y(n8933) );
  NBUFFX2_HVT U10159 ( .A(n8932), .Y(n8934) );
  NBUFFX2_HVT U10160 ( .A(n8932), .Y(n8935) );
  NBUFFX2_HVT U10161 ( .A(n8933), .Y(n8936) );
  NBUFFX2_HVT U10162 ( .A(n8933), .Y(n8937) );
  INVX0_HVT U10163 ( .A(n8938), .Y(n8940) );
  INVX0_HVT U10164 ( .A(n8938), .Y(n8941) );
  INVX0_HVT U10165 ( .A(n8938), .Y(n8942) );
  INVX0_HVT U10166 ( .A(n8938), .Y(n8943) );
  INVX0_HVT U10167 ( .A(n8939), .Y(n8944) );
  INVX0_HVT U10168 ( .A(n8939), .Y(n8945) );
  INVX0_HVT U10169 ( .A(n8939), .Y(n8946) );
  INVX1_HVT U10170 ( .A(n8911), .Y(n8956) );
  INVX0_HVT U10171 ( .A(n10125), .Y(n10124) );
  INVX0_HVT U10172 ( .A(n53), .Y(n10126) );
  NBUFFX2_HVT U10173 ( .A(n8977), .Y(n8970) );
  NBUFFX2_HVT U10174 ( .A(n8972), .Y(n8971) );
  NBUFFX2_HVT U10175 ( .A(n8972), .Y(n8973) );
  NBUFFX2_HVT U10176 ( .A(n8972), .Y(n8974) );
  NBUFFX2_HVT U10177 ( .A(n8972), .Y(n8975) );
  NBUFFX2_HVT U10178 ( .A(n8972), .Y(n8976) );
  NBUFFX2_HVT U10179 ( .A(n8983), .Y(n8986) );
  NBUFFX2_HVT U10180 ( .A(n8983), .Y(n8987) );
  INVX0_HVT U10181 ( .A(n8994), .Y(n8996) );
  INVX0_HVT U10182 ( .A(n8994), .Y(n8997) );
  INVX0_HVT U10183 ( .A(n8994), .Y(n8998) );
  INVX0_HVT U10184 ( .A(n8994), .Y(n8999) );
  INVX0_HVT U10185 ( .A(n8995), .Y(n9000) );
  INVX0_HVT U10186 ( .A(n8995), .Y(n9001) );
  INVX0_HVT U10187 ( .A(n8995), .Y(n9002) );
  INVX0_HVT U10188 ( .A(n8995), .Y(n9003) );
  INVX1_HVT U10189 ( .A(n8966), .Y(n9004) );
  INVX1_HVT U10190 ( .A(n8966), .Y(n9005) );
  INVX1_HVT U10191 ( .A(n9004), .Y(n9008) );
  INVX1_HVT U10192 ( .A(n9004), .Y(n9009) );
  INVX1_HVT U10193 ( .A(n9005), .Y(n9011) );
  INVX1_HVT U10194 ( .A(n9005), .Y(n9012) );
  INVX1_HVT U10195 ( .A(n8967), .Y(n9014) );
  INVX1_HVT U10196 ( .A(n8967), .Y(n9015) );
  INVX1_HVT U10197 ( .A(n9014), .Y(n9018) );
  INVX1_HVT U10198 ( .A(n9014), .Y(n9019) );
  INVX1_HVT U10199 ( .A(n9015), .Y(n9020) );
  INVX1_HVT U10200 ( .A(n9015), .Y(n9022) );
  NBUFFX2_HVT U10201 ( .A(n9040), .Y(n9028) );
  NBUFFX2_HVT U10202 ( .A(n9024), .Y(n9029) );
  NBUFFX2_HVT U10203 ( .A(n9041), .Y(n9030) );
  NBUFFX2_HVT U10204 ( .A(n9047), .Y(n9031) );
  NBUFFX2_HVT U10205 ( .A(n9035), .Y(n9032) );
  NBUFFX2_HVT U10206 ( .A(n9034), .Y(n9033) );
  NBUFFX2_HVT U10207 ( .A(n9035), .Y(n9038) );
  NBUFFX2_HVT U10208 ( .A(n9035), .Y(n9039) );
  INVX0_HVT U10209 ( .A(n4530), .Y(n9053) );
  INVX0_HVT U10210 ( .A(n4530), .Y(n9054) );
  INVX0_HVT U10211 ( .A(n9052), .Y(n9055) );
  INVX0_HVT U10212 ( .A(n9052), .Y(n9056) );
  INVX0_HVT U10213 ( .A(n10114), .Y(n9057) );
  INVX0_HVT U10214 ( .A(n10113), .Y(n9058) );
  INVX0_HVT U10215 ( .A(n4530), .Y(n9059) );
  INVX0_HVT U10216 ( .A(n4530), .Y(n9060) );
  INVX1_HVT U10217 ( .A(n9024), .Y(n9061) );
  INVX0_HVT U10218 ( .A(n10206), .Y(n9081) );
  INVX0_HVT U10219 ( .A(n10206), .Y(n9082) );
  NBUFFX2_HVT U10220 ( .A(n9083), .Y(n9084) );
  NBUFFX2_HVT U10221 ( .A(n9083), .Y(n9085) );
  NBUFFX2_HVT U10222 ( .A(n9098), .Y(n9086) );
  NBUFFX2_HVT U10223 ( .A(n9083), .Y(n9087) );
  NBUFFX2_HVT U10224 ( .A(n9092), .Y(n9088) );
  NBUFFX2_HVT U10225 ( .A(n9104), .Y(n9089) );
  NBUFFX2_HVT U10226 ( .A(n9099), .Y(n9090) );
  NBUFFX2_HVT U10227 ( .A(n4334), .Y(n9091) );
  NBUFFX2_HVT U10228 ( .A(n9092), .Y(n9094) );
  NBUFFX2_HVT U10229 ( .A(n9092), .Y(n9095) );
  NBUFFX2_HVT U10230 ( .A(n4334), .Y(n9096) );
  NBUFFX2_HVT U10231 ( .A(n4537), .Y(n9097) );
  NBUFFX2_HVT U10232 ( .A(n9098), .Y(n9100) );
  NBUFFX2_HVT U10233 ( .A(n9098), .Y(n9101) );
  NBUFFX2_HVT U10234 ( .A(n4537), .Y(n9102) );
  NBUFFX2_HVT U10235 ( .A(n9093), .Y(n9103) );
  NBUFFX2_HVT U10236 ( .A(n9104), .Y(n9106) );
  NBUFFX2_HVT U10237 ( .A(n9104), .Y(n9107) );
  NBUFFX2_HVT U10238 ( .A(n9105), .Y(n9108) );
  NBUFFX2_HVT U10239 ( .A(n9105), .Y(n9109) );
  INVX0_HVT U10240 ( .A(n9110), .Y(n9112) );
  INVX0_HVT U10241 ( .A(n9110), .Y(n9113) );
  INVX0_HVT U10242 ( .A(n9110), .Y(n9114) );
  INVX0_HVT U10243 ( .A(n9110), .Y(n9115) );
  INVX0_HVT U10244 ( .A(n9111), .Y(n9116) );
  INVX0_HVT U10245 ( .A(n9111), .Y(n9117) );
  INVX0_HVT U10246 ( .A(n9111), .Y(n9118) );
  INVX1_HVT U10247 ( .A(n9081), .Y(n9120) );
  INVX0_HVT U10248 ( .A(n40), .Y(n10206) );
  INVX0_HVT U10249 ( .A(n10256), .Y(n9137) );
  INVX0_HVT U10250 ( .A(n10256), .Y(n9138) );
  NBUFFX2_HVT U10251 ( .A(n9153), .Y(n9139) );
  NBUFFX2_HVT U10252 ( .A(n9154), .Y(n9140) );
  NBUFFX2_HVT U10253 ( .A(n9153), .Y(n9141) );
  NBUFFX2_HVT U10254 ( .A(n9154), .Y(n9142) );
  NBUFFX2_HVT U10255 ( .A(n9160), .Y(n9143) );
  NBUFFX2_HVT U10256 ( .A(n9148), .Y(n9144) );
  NBUFFX2_HVT U10257 ( .A(n9147), .Y(n9145) );
  NBUFFX2_HVT U10258 ( .A(n9159), .Y(n9146) );
  NBUFFX2_HVT U10259 ( .A(n9147), .Y(n9149) );
  NBUFFX2_HVT U10260 ( .A(n9147), .Y(n9150) );
  NBUFFX2_HVT U10261 ( .A(n9148), .Y(n9151) );
  NBUFFX2_HVT U10262 ( .A(n9148), .Y(n9152) );
  NBUFFX2_HVT U10263 ( .A(n9153), .Y(n9155) );
  NBUFFX2_HVT U10264 ( .A(n9153), .Y(n9156) );
  NBUFFX2_HVT U10265 ( .A(n9154), .Y(n9157) );
  NBUFFX2_HVT U10266 ( .A(n9154), .Y(n9158) );
  NBUFFX2_HVT U10267 ( .A(n9159), .Y(n9161) );
  NBUFFX2_HVT U10268 ( .A(n9159), .Y(n9162) );
  NBUFFX2_HVT U10269 ( .A(n9160), .Y(n9163) );
  NBUFFX2_HVT U10270 ( .A(n9160), .Y(n9164) );
  INVX0_HVT U10271 ( .A(n9165), .Y(n9167) );
  INVX0_HVT U10272 ( .A(n9165), .Y(n9168) );
  INVX0_HVT U10273 ( .A(n9165), .Y(n9169) );
  INVX0_HVT U10274 ( .A(n9165), .Y(n9170) );
  INVX0_HVT U10275 ( .A(n9166), .Y(n9171) );
  INVX0_HVT U10276 ( .A(n9166), .Y(n9172) );
  INVX0_HVT U10277 ( .A(n9166), .Y(n9173) );
  INVX0_HVT U10278 ( .A(n9166), .Y(n9174) );
  INVX1_HVT U10279 ( .A(n9137), .Y(n9175) );
  INVX1_HVT U10280 ( .A(n9137), .Y(n9176) );
  INVX1_HVT U10281 ( .A(n9175), .Y(n9177) );
  INVX1_HVT U10282 ( .A(n9175), .Y(n9178) );
  INVX1_HVT U10283 ( .A(n9175), .Y(n9179) );
  INVX1_HVT U10284 ( .A(n9175), .Y(n9180) );
  INVX1_HVT U10285 ( .A(n9176), .Y(n9181) );
  INVX1_HVT U10286 ( .A(n9176), .Y(n9182) );
  INVX1_HVT U10287 ( .A(n9176), .Y(n9183) );
  INVX1_HVT U10288 ( .A(n9176), .Y(n9184) );
  INVX1_HVT U10289 ( .A(n9138), .Y(n9185) );
  INVX1_HVT U10290 ( .A(n9138), .Y(n9186) );
  INVX1_HVT U10291 ( .A(n9185), .Y(n9187) );
  INVX1_HVT U10292 ( .A(n9185), .Y(n9188) );
  INVX1_HVT U10293 ( .A(n9185), .Y(n9189) );
  INVX1_HVT U10294 ( .A(n9185), .Y(n9190) );
  INVX1_HVT U10295 ( .A(n9186), .Y(n9191) );
  INVX1_HVT U10296 ( .A(n9186), .Y(n9192) );
  INVX1_HVT U10297 ( .A(n9186), .Y(n9193) );
  INVX1_HVT U10298 ( .A(n9186), .Y(n9194) );
  INVX0_HVT U10299 ( .A(n33), .Y(n10256) );
  INVX0_HVT U10300 ( .A(n10273), .Y(n9195) );
  INVX0_HVT U10301 ( .A(n10270), .Y(n9196) );
  NBUFFX2_HVT U10302 ( .A(n9211), .Y(n9197) );
  NBUFFX2_HVT U10303 ( .A(n9215), .Y(n9198) );
  NBUFFX2_HVT U10304 ( .A(n9211), .Y(n9199) );
  NBUFFX2_HVT U10305 ( .A(n9217), .Y(n9200) );
  NBUFFX2_HVT U10306 ( .A(n9212), .Y(n9201) );
  NBUFFX2_HVT U10307 ( .A(n9217), .Y(n9202) );
  NBUFFX2_HVT U10308 ( .A(n9205), .Y(n9203) );
  NBUFFX2_HVT U10309 ( .A(n9206), .Y(n9204) );
  NBUFFX2_HVT U10310 ( .A(n9205), .Y(n9207) );
  NBUFFX2_HVT U10311 ( .A(n9205), .Y(n9208) );
  NBUFFX2_HVT U10312 ( .A(n9206), .Y(n9209) );
  NBUFFX2_HVT U10313 ( .A(n9206), .Y(n9210) );
  NBUFFX2_HVT U10314 ( .A(n9211), .Y(n9213) );
  NBUFFX2_HVT U10315 ( .A(n9211), .Y(n9214) );
  NBUFFX2_HVT U10316 ( .A(n9212), .Y(n9215) );
  NBUFFX2_HVT U10317 ( .A(n9212), .Y(n9216) );
  NBUFFX2_HVT U10318 ( .A(n9217), .Y(n9219) );
  NBUFFX2_HVT U10319 ( .A(n9217), .Y(n9220) );
  NBUFFX2_HVT U10320 ( .A(n9218), .Y(n9221) );
  NBUFFX2_HVT U10321 ( .A(n9218), .Y(n9222) );
  INVX0_HVT U10322 ( .A(n9223), .Y(n9225) );
  INVX0_HVT U10323 ( .A(n9223), .Y(n9226) );
  INVX0_HVT U10324 ( .A(n9223), .Y(n9227) );
  INVX0_HVT U10325 ( .A(n9223), .Y(n9228) );
  INVX0_HVT U10326 ( .A(n9224), .Y(n9229) );
  INVX0_HVT U10327 ( .A(n9224), .Y(n9230) );
  INVX0_HVT U10328 ( .A(n9224), .Y(n9231) );
  INVX1_HVT U10329 ( .A(n9195), .Y(n9232) );
  INVX1_HVT U10330 ( .A(n9195), .Y(n9233) );
  INVX1_HVT U10331 ( .A(n9232), .Y(n9234) );
  INVX1_HVT U10332 ( .A(n9232), .Y(n9235) );
  INVX1_HVT U10333 ( .A(n9232), .Y(n9236) );
  INVX1_HVT U10334 ( .A(n9233), .Y(n9241) );
  INVX1_HVT U10335 ( .A(n9196), .Y(n9242) );
  INVX1_HVT U10336 ( .A(n9196), .Y(n9243) );
  INVX1_HVT U10337 ( .A(n9243), .Y(n9248) );
  INVX1_HVT U10338 ( .A(n9243), .Y(n9250) );
  INVX0_HVT U10339 ( .A(n30), .Y(n10273) );
  INVX0_HVT U10340 ( .A(n4424), .Y(n9252) );
  NBUFFX2_HVT U10341 ( .A(n9254), .Y(n9255) );
  NBUFFX2_HVT U10342 ( .A(n9254), .Y(n9256) );
  NBUFFX2_HVT U10343 ( .A(n9254), .Y(n9257) );
  NBUFFX2_HVT U10344 ( .A(n9258), .Y(n9259) );
  NBUFFX2_HVT U10345 ( .A(n9258), .Y(n9260) );
  NBUFFX2_HVT U10346 ( .A(n9258), .Y(n9261) );
  NBUFFX2_HVT U10347 ( .A(n9254), .Y(n9262) );
  NBUFFX2_HVT U10348 ( .A(n9263), .Y(n9264) );
  NBUFFX2_HVT U10349 ( .A(n9263), .Y(n9265) );
  NBUFFX2_HVT U10350 ( .A(n9269), .Y(n9266) );
  NBUFFX2_HVT U10351 ( .A(n9263), .Y(n9267) );
  NBUFFX2_HVT U10352 ( .A(n9268), .Y(n9270) );
  NBUFFX2_HVT U10353 ( .A(n9268), .Y(n9271) );
  NBUFFX2_HVT U10354 ( .A(n9269), .Y(n9272) );
  NBUFFX2_HVT U10355 ( .A(n9269), .Y(n9273) );
  NBUFFX2_HVT U10356 ( .A(n9274), .Y(n9275) );
  NBUFFX2_HVT U10357 ( .A(n9274), .Y(n9276) );
  NBUFFX2_HVT U10358 ( .A(n9268), .Y(n9277) );
  NBUFFX2_HVT U10359 ( .A(n9274), .Y(n9278) );
  INVX0_HVT U10360 ( .A(n9279), .Y(n9281) );
  INVX0_HVT U10361 ( .A(n9279), .Y(n9282) );
  INVX0_HVT U10362 ( .A(n9279), .Y(n9283) );
  INVX0_HVT U10363 ( .A(n9279), .Y(n9284) );
  INVX0_HVT U10364 ( .A(n9280), .Y(n9285) );
  INVX0_HVT U10365 ( .A(n9280), .Y(n9286) );
  INVX1_HVT U10366 ( .A(n9252), .Y(n9288) );
  INVX1_HVT U10367 ( .A(n9288), .Y(n9292) );
  INVX1_HVT U10368 ( .A(n9253), .Y(n9296) );
  INVX0_HVT U10369 ( .A(n10303), .Y(n10300) );
  INVX0_HVT U10370 ( .A(n10330), .Y(n10328) );
  INVX0_HVT U10371 ( .A(n10149), .Y(n10148) );
  INVX0_HVT U10372 ( .A(n6578), .Y(n10138) );
  INVX0_HVT U10373 ( .A(n10147), .Y(n10137) );
  INVX0_HVT U10374 ( .A(n6578), .Y(n10144) );
  INVX0_HVT U10375 ( .A(n10148), .Y(n10145) );
endmodule

