
module sbox_7 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n50, n210, n211, n212, n213, n216, n217, n218, n219, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  NAND2X0_HVT U3 ( .A1(n294), .A2(n289), .Y(n582) );
  NAND2X0_HVT U4 ( .A1(n288), .A2(n582), .Y(n581) );
  NAND2X0_HVT U5 ( .A1(n292), .A2(n275), .Y(n579) );
  NAND2X0_HVT U13 ( .A1(n571), .A2(n291), .Y(n572) );
  NAND2X0_HVT U15 ( .A1(n582), .A2(n277), .Y(n569) );
  NAND2X0_HVT U21 ( .A1(n288), .A2(n298), .Y(n563) );
  NAND2X0_HVT U24 ( .A1(n283), .A2(n50), .Y(n561) );
  NAND2X0_HVT U33 ( .A1(n359), .A2(n23), .Y(n552) );
  NAND2X0_HVT U35 ( .A1(n281), .A2(n50), .Y(n550) );
  NAND2X0_HVT U42 ( .A1(n296), .A2(n283), .Y(n543) );
  MUX41X1_HVT U51 ( .A1(n347), .A3(n305), .A2(n322), .A4(n323), .S0(n303), 
        .S1(n269), .Y(n535) );
  NAND2X0_HVT U53 ( .A1(n532), .A2(n542), .Y(n533) );
  NAND2X0_HVT U56 ( .A1(n288), .A2(n528), .Y(n529) );
  MUX41X1_HVT U57 ( .A1(n348), .A3(n565), .A2(n529), .A4(n574), .S0(n303), 
        .S1(n269), .Y(n527) );
  NAND2X0_HVT U58 ( .A1(n291), .A2(n582), .Y(n526) );
  MUX41X1_HVT U59 ( .A1(n263), .A3(n526), .A2(n261), .A4(n321), .S0(n303), 
        .S1(n269), .Y(n525) );
  MUX41X1_HVT U61 ( .A1(n260), .A3(n320), .A2(n319), .A4(n276), .S0(n303), 
        .S1(n269), .Y(n523) );
  NAND2X0_HVT U62 ( .A1(n23), .A2(n290), .Y(n522) );
  MUX41X1_HVT U63 ( .A1(n522), .A3(n312), .A2(n342), .A4(n318), .S0(n303), 
        .S1(n269), .Y(n521) );
  AO21X1_HVT U66 ( .A1(n316), .A2(n271), .A3(n341), .Y(n518) );
  MUX41X1_HVT U68 ( .A1(n314), .A3(n518), .A2(n517), .A4(n519), .S0(n264), 
        .S1(n240), .Y(n516) );
  MUX41X1_HVT U69 ( .A1(n516), .A3(n524), .A2(n520), .A4(n530), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n285), .A2(n511), .Y(n512) );
  MUX41X1_HVT U74 ( .A1(n513), .A3(n559), .A2(n512), .A4(n561), .S0(n267), 
        .S1(n302), .Y(n510) );
  MUX41X1_HVT U75 ( .A1(n345), .A3(n350), .A2(n363), .A4(n325), .S0(n264), 
        .S1(n239), .Y(n509) );
  MUX41X1_HVT U77 ( .A1(n576), .A3(n352), .A2(n508), .A4(n351), .S0(n272), 
        .S1(n300), .Y(n507) );
  AND3X1_HVT U80 ( .A1(n289), .A2(n528), .A3(n503), .Y(n504) );
  MUX41X1_HVT U82 ( .A1(n540), .A3(n323), .A2(n306), .A4(n570), .S0(n264), 
        .S1(n302), .Y(n501) );
  AND2X1_HVT U83 ( .A1(n296), .A2(n241), .Y(n500) );
  MUX41X1_HVT U84 ( .A1(n324), .A3(n578), .A2(n568), .A4(n500), .S0(n264), 
        .S1(n239), .Y(n499) );
  NAND2X0_HVT U85 ( .A1(n23), .A2(n362), .Y(n498) );
  MUX41X1_HVT U86 ( .A1(n350), .A3(n498), .A2(n258), .A4(n256), .S0(n264), 
        .S1(n239), .Y(n497) );
  MUX41X1_HVT U87 ( .A1(n497), .A3(n501), .A2(n499), .A4(n502), .S0(in[0]), 
        .S1(n247), .Y(n496) );
  MUX41X1_HVT U90 ( .A1(n539), .A3(n543), .A2(n347), .A4(n495), .S0(n265), 
        .S1(n302), .Y(n494) );
  AO21X1_HVT U93 ( .A1(n274), .A2(n490), .A3(n346), .Y(n491) );
  MUX41X1_HVT U96 ( .A1(n306), .A3(n259), .A2(n349), .A4(n488), .S0(n264), 
        .S1(n239), .Y(n487) );
  MUX41X1_HVT U97 ( .A1(n345), .A3(n259), .A2(n218), .A4(n569), .S0(n264), 
        .S1(n240), .Y(n486) );
  MUX41X1_HVT U98 ( .A1(n486), .A3(n489), .A2(n487), .A4(n494), .S0(n282), 
        .S1(n247), .Y(n485) );
  NAND2X0_HVT U101 ( .A1(n481), .A2(n480), .Y(n482) );
  MUX41X1_HVT U103 ( .A1(n582), .A3(n315), .A2(n328), .A4(n550), .S0(n264), 
        .S1(n240), .Y(n478) );
  MUX41X1_HVT U105 ( .A1(n327), .A3(n537), .A2(n477), .A4(n344), .S0(n264), 
        .S1(n272), .Y(n476) );
  NAND2X0_HVT U110 ( .A1(n289), .A2(n471), .Y(n472) );
  AND2X1_HVT U115 ( .A1(n217), .A2(n276), .Y(n466) );
  NAND2X0_HVT U123 ( .A1(n457), .A2(n456), .Y(n458) );
  MUX41X1_HVT U125 ( .A1(n563), .A3(n263), .A2(n314), .A4(n354), .S0(n265), 
        .S1(n303), .Y(n454) );
  AND3X1_HVT U128 ( .A1(n267), .A2(n23), .A3(n241), .Y(n451) );
  MUX41X1_HVT U131 ( .A1(n449), .A3(n451), .A2(n450), .A4(n452), .S0(n271), 
        .S1(n303), .Y(n448) );
  MUX41X1_HVT U136 ( .A1(n256), .A3(n552), .A2(n356), .A4(n549), .S0(n265), 
        .S1(n303), .Y(n444) );
  MUX41X1_HVT U139 ( .A1(n442), .A3(n445), .A2(n444), .A4(n446), .S0(n282), 
        .S1(n270), .Y(n441) );
  AND2X1_HVT U140 ( .A1(n284), .A2(n23), .Y(n440) );
  NAND2X0_HVT U146 ( .A1(n293), .A2(n291), .Y(n511) );
  MUX41X1_HVT U147 ( .A1(n356), .A3(n511), .A2(n345), .A4(n539), .S0(n267), 
        .S1(n303), .Y(n434) );
  MUX41X1_HVT U148 ( .A1(n434), .A3(n438), .A2(n435), .A4(n439), .S0(in[0]), 
        .S1(n247), .Y(n433) );
  OA21X1_HVT U151 ( .A1(n545), .A2(n250), .A3(n430), .Y(n431) );
  MUX41X1_HVT U153 ( .A1(n472), .A3(n260), .A2(n289), .A4(n308), .S0(n265), 
        .S1(n239), .Y(n428) );
  AND2X1_HVT U154 ( .A1(n274), .A2(n283), .Y(n427) );
  NAND2X0_HVT U158 ( .A1(n296), .A2(n362), .Y(n423) );
  MUX41X1_HVT U159 ( .A1(n572), .A3(n276), .A2(n423), .A4(n245), .S0(n300), 
        .S1(n239), .Y(n422) );
  MUX41X1_HVT U160 ( .A1(n422), .A3(n428), .A2(n424), .A4(n429), .S0(n282), 
        .S1(n270), .Y(n421) );
  AND2X1_HVT U162 ( .A1(n578), .A2(n511), .Y(n419) );
  MUX41X1_HVT U163 ( .A1(n320), .A3(n419), .A2(n257), .A4(n420), .S0(n300), 
        .S1(n302), .Y(n418) );
  MUX41X1_HVT U165 ( .A1(n563), .A3(n329), .A2(n539), .A4(n417), .S0(n303), 
        .S1(n299), .Y(n416) );
  NAND2X0_HVT U166 ( .A1(n291), .A2(n528), .Y(n415) );
  NAND2X0_HVT U167 ( .A1(n363), .A2(n50), .Y(n414) );
  MUX41X1_HVT U168 ( .A1(n348), .A3(n284), .A2(n414), .A4(n415), .S0(n300), 
        .S1(n239), .Y(n413) );
  MUX41X1_HVT U172 ( .A1(n410), .A3(n416), .A2(n413), .A4(n418), .S0(n282), 
        .S1(in[5]), .Y(n409) );
  NAND2X0_HVT U174 ( .A1(n218), .A2(n578), .Y(n571) );
  MUX41X1_HVT U176 ( .A1(n279), .A3(n408), .A2(n353), .A4(n571), .S0(n303), 
        .S1(n299), .Y(n407) );
  NAND2X0_HVT U177 ( .A1(n294), .A2(n280), .Y(n406) );
  MUX41X1_HVT U178 ( .A1(n567), .A3(n406), .A2(n357), .A4(n547), .S0(n264), 
        .S1(n302), .Y(n405) );
  MUX41X1_HVT U179 ( .A1(n557), .A3(n358), .A2(n310), .A4(n357), .S0(n299), 
        .S1(n273), .Y(n404) );
  MUX41X1_HVT U180 ( .A1(n313), .A3(n576), .A2(n572), .A4(n255), .S0(n272), 
        .S1(n299), .Y(n403) );
  MUX41X1_HVT U181 ( .A1(n403), .A3(n405), .A2(n404), .A4(n407), .S0(n282), 
        .S1(n270), .Y(n402) );
  MUX41X1_HVT U182 ( .A1(n337), .A3(n287), .A2(n339), .A4(n326), .S0(n303), 
        .S1(n300), .Y(n401) );
  OA21X1_HVT U184 ( .A1(n551), .A2(n250), .A3(n324), .Y(n399) );
  MUX41X1_HVT U186 ( .A1(n259), .A3(n546), .A2(n511), .A4(n539), .S0(n299), 
        .S1(n240), .Y(n397) );
  MUX41X1_HVT U189 ( .A1(n395), .A3(n571), .A2(n396), .A4(n344), .S0(n272), 
        .S1(n300), .Y(n394) );
  MUX41X1_HVT U190 ( .A1(n394), .A3(n397), .A2(n398), .A4(n401), .S0(n270), 
        .S1(in[0]), .Y(n393) );
  MUX41X1_HVT U194 ( .A1(n544), .A3(n558), .A2(n355), .A4(n284), .S0(n272), 
        .S1(n299), .Y(n390) );
  AO21X1_HVT U197 ( .A1(n258), .A2(n273), .A3(n346), .Y(n387) );
  OA21X1_HVT U201 ( .A1(n577), .A2(n250), .A3(n336), .Y(n383) );
  MUX41X1_HVT U205 ( .A1(n241), .A3(n582), .A2(n358), .A4(n331), .S0(n300), 
        .S1(n240), .Y(n379) );
  NAND2X0_HVT U208 ( .A1(n295), .A2(n288), .Y(n471) );
  NAND2X0_HVT U212 ( .A1(n295), .A2(n285), .Y(n528) );
  NAND2X0_HVT U214 ( .A1(n578), .A2(n298), .Y(n377) );
  NAND2X0_HVT U215 ( .A1(n471), .A2(n286), .Y(n376) );
  NAND2X0_HVT U218 ( .A1(n360), .A2(n293), .Y(n430) );
  NAND2X0_HVT U220 ( .A1(n273), .A2(n377), .Y(n503) );
  INVX2_HVT U1 ( .A(n219), .Y(n300) );
  NAND2X2_HVT U2 ( .A1(n237), .A2(n238), .Y(out[4]) );
  INVX2_HVT U6 ( .A(in[7]), .Y(n250) );
  IBUFFX2_HVT U7 ( .A(in[1]), .Y(n23) );
  IBUFFX2_HVT U8 ( .A(in[1]), .Y(n50) );
  INVX0_HVT U9 ( .A(in[1]), .Y(n297) );
  AO21X2_HVT U10 ( .A1(n50), .A2(n360), .A3(n250), .Y(n481) );
  MUX21X1_HVT U11 ( .A1(n255), .A2(n568), .S0(n212), .Y(n384) );
  MUX21X1_HVT U12 ( .A1(n278), .A2(n283), .S0(n296), .Y(n562) );
  OA21X1_HVT U14 ( .A1(n261), .A2(n304), .A3(n554), .Y(n411) );
  XNOR2X2_HVT U16 ( .A1(n279), .A2(in[3]), .Y(n210) );
  INVX8_HVT U17 ( .A(n210), .Y(n578) );
  MUX41X1_HVT U18 ( .A1(n572), .A3(n529), .A2(n562), .A4(n333), .S0(n211), 
        .S1(n240), .Y(n380) );
  IBUFFX16_HVT U19 ( .A(n299), .Y(n211) );
  NBUFFX2_HVT U20 ( .A(n210), .Y(n278) );
  IBUFFX16_HVT U22 ( .A(n272), .Y(n212) );
  MUX21X2_HVT U23 ( .A1(n443), .A2(n581), .S0(n268), .Y(n442) );
  MUX21X2_HVT U25 ( .A1(n496), .A2(n506), .S0(in[6]), .Y(out[1]) );
  INVX1_HVT U26 ( .A(n297), .Y(n217) );
  AO21X2_HVT U27 ( .A1(n268), .A2(n284), .A3(n578), .Y(n463) );
  MUX21X2_HVT U28 ( .A1(n562), .A2(n337), .S0(n273), .Y(n443) );
  INVX2_HVT U29 ( .A(n250), .Y(n303) );
  MUX41X1_HVT U30 ( .A1(n380), .A3(n382), .A2(n379), .A4(n381), .S0(n213), 
        .S1(n216), .Y(n378) );
  IBUFFX16_HVT U31 ( .A(n231), .Y(n213) );
  IBUFFX16_HVT U32 ( .A(n270), .Y(n216) );
  NBUFFX4_HVT U34 ( .A(n364), .Y(n279) );
  MUX21X1_HVT U36 ( .A1(n475), .A2(n485), .S0(in[6]), .Y(out[2]) );
  INVX0_HVT U37 ( .A(in[7]), .Y(n304) );
  MUX21X2_HVT U38 ( .A1(n378), .A2(n385), .S0(in[6]), .Y(out[7]) );
  INVX1_HVT U39 ( .A(n469), .Y(n252) );
  INVX1_HVT U40 ( .A(n235), .Y(n299) );
  MUX21X1_HVT U41 ( .A1(n387), .A2(n388), .S0(n219), .Y(n386) );
  NAND2X0_HVT U43 ( .A1(n340), .A2(n232), .Y(n233) );
  INVX0_HVT U44 ( .A(n543), .Y(n340) );
  INVX0_HVT U45 ( .A(n254), .Y(n236) );
  INVX0_HVT U46 ( .A(n298), .Y(n293) );
  INVX1_HVT U47 ( .A(n273), .Y(n232) );
  NBUFFX2_HVT U48 ( .A(in[7]), .Y(n273) );
  INVX1_HVT U49 ( .A(n301), .Y(n247) );
  INVX1_HVT U50 ( .A(n265), .Y(n235) );
  INVX0_HVT U52 ( .A(n268), .Y(n219) );
  INVX1_HVT U54 ( .A(n282), .Y(n231) );
  MUX21X1_HVT U55 ( .A1(n402), .A2(n393), .S0(n254), .Y(out[6]) );
  MUX21X1_HVT U60 ( .A1(n409), .A2(n421), .S0(in[6]), .Y(out[5]) );
  MUX41X1_HVT U64 ( .A1(n284), .A3(n343), .A2(n276), .A4(n324), .S0(n235), 
        .S1(n232), .Y(n438) );
  INVX1_HVT U65 ( .A(n297), .Y(n218) );
  INVX0_HVT U67 ( .A(n297), .Y(n294) );
  MUX41X1_HVT U70 ( .A1(n550), .A3(n543), .A2(n392), .A4(n536), .S0(n235), 
        .S1(n240), .Y(n391) );
  MUX21X1_HVT U71 ( .A1(n459), .A2(n458), .S0(n274), .Y(n455) );
  MUX21X2_HVT U72 ( .A1(n307), .A2(n460), .S0(n267), .Y(n459) );
  MUX21X2_HVT U76 ( .A1(n570), .A2(n331), .S0(n219), .Y(n484) );
  MUX21X1_HVT U78 ( .A1(n472), .A2(n554), .S0(n235), .Y(n470) );
  OA21X2_HVT U79 ( .A1(n309), .A2(n304), .A3(n554), .Y(n436) );
  MUX21X2_HVT U81 ( .A1(n362), .A2(n349), .S0(n274), .Y(n515) );
  INVX1_HVT U88 ( .A(n553), .Y(n332) );
  MUX41X1_HVT U89 ( .A1(n548), .A3(n584), .A2(n349), .A4(n578), .S0(n235), 
        .S1(n232), .Y(n389) );
  MUX41X1_HVT U91 ( .A1(n514), .A3(n509), .A2(n510), .A4(n507), .S0(n231), 
        .S1(n301), .Y(n506) );
  IBUFFX2_HVT U92 ( .A(n548), .Y(n335) );
  MUX21X2_HVT U94 ( .A1(n462), .A2(n465), .S0(n271), .Y(n461) );
  NAND2X0_HVT U95 ( .A1(n357), .A2(n273), .Y(n234) );
  NAND2X0_HVT U99 ( .A1(n233), .A2(n234), .Y(n388) );
  MUX41X1_HVT U100 ( .A1(n573), .A3(n553), .A2(n549), .A4(n338), .S0(n268), 
        .S1(n304), .Y(n381) );
  IBUFFX2_HVT U102 ( .A(n304), .Y(n302) );
  IBUFFX2_HVT U104 ( .A(n549), .Y(n334) );
  IBUFFX2_HVT U106 ( .A(in[1]), .Y(n298) );
  MUX41X1_HVT U107 ( .A1(n483), .A3(n478), .A2(n479), .A4(n476), .S0(n231), 
        .S1(n301), .Y(n475) );
  MUX21X2_HVT U108 ( .A1(n541), .A2(n515), .S0(n266), .Y(n514) );
  INVX1_HVT U109 ( .A(n373), .Y(n349) );
  INVX1_HVT U111 ( .A(n366), .Y(n357) );
  MUX41X1_HVT U112 ( .A1(n554), .A3(n325), .A2(n466), .A4(n572), .S0(n235), 
        .S1(n232), .Y(n465) );
  NAND2X0_HVT U113 ( .A1(n441), .A2(n236), .Y(n237) );
  NAND2X0_HVT U114 ( .A1(n433), .A2(n254), .Y(n238) );
  INVX1_HVT U116 ( .A(n304), .Y(n239) );
  INVX1_HVT U117 ( .A(n304), .Y(n240) );
  MUX41X1_HVT U118 ( .A1(n391), .A3(n389), .A2(n390), .A4(n386), .S0(n231), 
        .S1(n301), .Y(n385) );
  MUX21X1_HVT U119 ( .A1(n278), .A2(n362), .S0(n294), .Y(n577) );
  OA21X1_HVT U120 ( .A1(n335), .A2(n235), .A3(n321), .Y(n473) );
  INVX1_HVT U121 ( .A(n244), .Y(n445) );
  INVX0_HVT U122 ( .A(n558), .Y(n246) );
  INVX0_HVT U124 ( .A(n579), .Y(n245) );
  NBUFFX2_HVT U126 ( .A(in[5]), .Y(n271) );
  INVX1_HVT U127 ( .A(in[5]), .Y(n301) );
  INVX0_HVT U129 ( .A(in[6]), .Y(n254) );
  INVX1_HVT U130 ( .A(n281), .Y(n241) );
  NAND2X0_HVT U132 ( .A1(n383), .A2(n219), .Y(n242) );
  NAND2X0_HVT U133 ( .A1(n384), .A2(n266), .Y(n243) );
  NAND2X0_HVT U134 ( .A1(n242), .A2(n243), .Y(n382) );
  MUX21X1_HVT U135 ( .A1(n275), .A2(n277), .S0(n298), .Y(n568) );
  NBUFFX2_HVT U137 ( .A(n210), .Y(n277) );
  MUX41X1_HVT U138 ( .A1(n332), .A3(n440), .A2(n336), .A4(n560), .S0(n235), 
        .S1(n232), .Y(n439) );
  INVX0_HVT U141 ( .A(n568), .Y(n319) );
  IBUFFX2_HVT U142 ( .A(n23), .Y(n295) );
  MUX41X1_HVT U143 ( .A1(n246), .A3(n245), .A2(n284), .A4(n368), .S0(n219), 
        .S1(n232), .Y(n244) );
  INVX1_HVT U144 ( .A(n368), .Y(n355) );
  MUX41X1_HVT U145 ( .A1(n461), .A3(n448), .A2(n467), .A4(n453), .S0(n254), 
        .S1(in[0]), .Y(out[3]) );
  NAND2X0_HVT U149 ( .A1(n455), .A2(n247), .Y(n248) );
  NAND2X0_HVT U150 ( .A1(n454), .A2(n301), .Y(n249) );
  NAND2X0_HVT U152 ( .A1(n248), .A2(n249), .Y(n453) );
  MUX21X2_HVT U155 ( .A1(n525), .A2(n527), .S0(n266), .Y(n524) );
  MUX21X2_HVT U156 ( .A1(n531), .A2(n535), .S0(n267), .Y(n530) );
  MUX41X1_HVT U157 ( .A1(n468), .A3(n470), .A2(n474), .A4(n473), .S0(n239), 
        .S1(n271), .Y(n467) );
  INVX0_HVT U161 ( .A(n251), .Y(n468) );
  XOR2X1_HVT U164 ( .A1(n235), .A2(n304), .Y(n538) );
  MUX21X1_HVT U169 ( .A1(n363), .A2(n252), .S0(n253), .Y(n251) );
  XNOR2X1_HVT U170 ( .A1(n217), .A2(n300), .Y(n253) );
  INVX0_HVT U171 ( .A(in[3]), .Y(n361) );
  MUX21X2_HVT U173 ( .A1(n260), .A2(n484), .S0(n538), .Y(n483) );
  INVX1_HVT U175 ( .A(n287), .Y(n359) );
  AND2X1_HVT U183 ( .A1(n278), .A2(n528), .Y(n255) );
  MUX21X1_HVT U185 ( .A1(n257), .A2(n319), .S0(n265), .Y(n450) );
  NBUFFX2_HVT U187 ( .A(n210), .Y(n276) );
  NBUFFX2_HVT U188 ( .A(n580), .Y(n287) );
  INVX1_HVT U191 ( .A(n583), .Y(n363) );
  MUX21X1_HVT U192 ( .A1(n359), .A2(n362), .S0(n271), .Y(n532) );
  NBUFFX2_HVT U193 ( .A(n580), .Y(n288) );
  MUX21X1_HVT U195 ( .A1(n315), .A2(n360), .S0(n271), .Y(n517) );
  AND2X1_HVT U196 ( .A1(n289), .A2(n511), .Y(n256) );
  MUX21X1_HVT U198 ( .A1(n289), .A2(n277), .S0(n217), .Y(n544) );
  MUX21X1_HVT U199 ( .A1(n288), .A2(n578), .S0(n294), .Y(n548) );
  MUX21X1_HVT U200 ( .A1(n276), .A2(n281), .S0(n294), .Y(n480) );
  MUX21X1_HVT U202 ( .A1(n359), .A2(n363), .S0(n295), .Y(n408) );
  MUX21X1_HVT U203 ( .A1(n277), .A2(n359), .S0(n296), .Y(n488) );
  MUX21X1_HVT U204 ( .A1(n363), .A2(n362), .S0(n292), .Y(n558) );
  MUX21X1_HVT U206 ( .A1(n362), .A2(n359), .S0(n296), .Y(n547) );
  MUX21X1_HVT U207 ( .A1(n275), .A2(n363), .S0(n218), .Y(n545) );
  MUX21X1_HVT U209 ( .A1(n578), .A2(n360), .S0(n293), .Y(n368) );
  NAND2X0_HVT U210 ( .A1(n279), .A2(n361), .Y(n580) );
  MUX21X1_HVT U211 ( .A1(n578), .A2(n363), .S0(n296), .Y(n560) );
  MUX21X1_HVT U213 ( .A1(n362), .A2(n277), .S0(n293), .Y(n420) );
  MUX21X1_HVT U216 ( .A1(n288), .A2(n286), .S0(n218), .Y(n495) );
  MUX21X1_HVT U217 ( .A1(n578), .A2(n281), .S0(n292), .Y(n508) );
  XOR2X1_HVT U219 ( .A1(n578), .A2(n295), .Y(n539) );
  INVX1_HVT U221 ( .A(n284), .Y(n360) );
  INVX1_HVT U222 ( .A(n584), .Y(n362) );
  MUX21X1_HVT U223 ( .A1(n362), .A2(n275), .S0(n217), .Y(n551) );
  MUX21X1_HVT U224 ( .A1(n281), .A2(n359), .S0(n293), .Y(n556) );
  MUX21X1_HVT U225 ( .A1(n330), .A2(n447), .S0(n267), .Y(n446) );
  MUX21X1_HVT U226 ( .A1(n354), .A2(n286), .S0(n273), .Y(n447) );
  MUX21X1_HVT U227 ( .A1(n463), .A2(n464), .S0(n273), .Y(n462) );
  MUX21X1_HVT U228 ( .A1(n308), .A2(n333), .S0(n265), .Y(n464) );
  NBUFFX2_HVT U229 ( .A(n583), .Y(n289) );
  MUX21X1_HVT U230 ( .A1(n275), .A2(n281), .S0(n294), .Y(n392) );
  XOR2X1_HVT U231 ( .A1(n289), .A2(n292), .Y(n536) );
  MUX21X1_HVT U232 ( .A1(n359), .A2(n280), .S0(n295), .Y(n369) );
  MUX21X1_HVT U233 ( .A1(n275), .A2(n578), .S0(n295), .Y(n371) );
  MUX21X1_HVT U234 ( .A1(n291), .A2(n285), .S0(n218), .Y(n554) );
  MUX21X1_HVT U235 ( .A1(n288), .A2(n275), .S0(n294), .Y(n573) );
  MUX21X1_HVT U236 ( .A1(n280), .A2(n275), .S0(n293), .Y(n460) );
  XOR2X1_HVT U237 ( .A1(n217), .A2(n360), .Y(n540) );
  MUX21X1_HVT U238 ( .A1(n275), .A2(n291), .S0(n293), .Y(n395) );
  MUX21X1_HVT U239 ( .A1(n584), .A2(n289), .S0(n295), .Y(n396) );
  MUX21X1_HVT U240 ( .A1(n360), .A2(n359), .S0(n295), .Y(n566) );
  MUX21X1_HVT U241 ( .A1(n290), .A2(n285), .S0(n296), .Y(n570) );
  MUX21X1_HVT U242 ( .A1(n287), .A2(n291), .S0(n295), .Y(n490) );
  MUX21X1_HVT U243 ( .A1(n275), .A2(n362), .S0(n292), .Y(n574) );
  NBUFFX2_HVT U244 ( .A(n583), .Y(n290) );
  MUX21X1_HVT U245 ( .A1(n285), .A2(n275), .S0(n296), .Y(n373) );
  MUX21X1_HVT U246 ( .A1(n290), .A2(n280), .S0(n293), .Y(n375) );
  XNOR2X1_HVT U247 ( .A1(n287), .A2(n217), .Y(n257) );
  XNOR2X1_HVT U248 ( .A1(n584), .A2(n296), .Y(n258) );
  AND2X1_HVT U249 ( .A1(n218), .A2(n363), .Y(n259) );
  MUX21X1_HVT U250 ( .A1(n290), .A2(n288), .S0(n218), .Y(n367) );
  AND2X1_HVT U251 ( .A1(n291), .A2(n471), .Y(n260) );
  MUX21X1_HVT U252 ( .A1(n286), .A2(n280), .S0(n293), .Y(n513) );
  MUX21X1_HVT U253 ( .A1(n286), .A2(n291), .S0(n267), .Y(n457) );
  XOR2X1_HVT U254 ( .A1(n279), .A2(n217), .Y(n559) );
  NBUFFX2_HVT U255 ( .A(in[7]), .Y(n272) );
  NBUFFX2_HVT U256 ( .A(n361), .Y(n275) );
  NBUFFX2_HVT U257 ( .A(in[7]), .Y(n274) );
  NBUFFX2_HVT U258 ( .A(in[2]), .Y(n265) );
  NBUFFX2_HVT U259 ( .A(n268), .Y(n266) );
  NBUFFX2_HVT U260 ( .A(in[5]), .Y(n270) );
  NBUFFX2_HVT U261 ( .A(in[2]), .Y(n267) );
  NBUFFX2_HVT U262 ( .A(in[2]), .Y(n268) );
  NBUFFX2_HVT U263 ( .A(n247), .Y(n269) );
  NBUFFX2_HVT U264 ( .A(in[2]), .Y(n264) );
  MUX21X1_HVT U265 ( .A1(n482), .A2(n330), .S0(n267), .Y(n479) );
  MUX21X1_HVT U266 ( .A1(n399), .A2(n400), .S0(n266), .Y(n398) );
  MUX21X1_HVT U267 ( .A1(n498), .A2(n283), .S0(n273), .Y(n400) );
  MUX21X1_HVT U268 ( .A1(n521), .A2(n523), .S0(n266), .Y(n520) );
  XOR2X1_HVT U269 ( .A1(n217), .A2(n283), .Y(n537) );
  MUX21X1_HVT U270 ( .A1(n285), .A2(n278), .S0(n218), .Y(n477) );
  NAND2X0_HVT U271 ( .A1(in[3]), .A2(n281), .Y(n583) );
  NBUFFX2_HVT U272 ( .A(n364), .Y(n281) );
  MUX21X1_HVT U273 ( .A1(n505), .A2(n504), .S0(n268), .Y(n502) );
  MUX21X1_HVT U274 ( .A1(n564), .A2(n286), .S0(n274), .Y(n505) );
  AND2X1_HVT U275 ( .A1(n278), .A2(n23), .Y(n261) );
  NBUFFX2_HVT U276 ( .A(n575), .Y(n284) );
  MUX21X1_HVT U277 ( .A1(n283), .A2(n359), .S0(n294), .Y(n546) );
  MUX21X1_HVT U278 ( .A1(n431), .A2(n432), .S0(n268), .Y(n429) );
  MUX21X1_HVT U279 ( .A1(n351), .A2(n360), .S0(n273), .Y(n432) );
  XOR2X1_HVT U280 ( .A1(n250), .A2(n558), .Y(n541) );
  MUX21X1_HVT U281 ( .A1(n412), .A2(n411), .S0(n267), .Y(n410) );
  MUX21X1_HVT U282 ( .A1(n286), .A2(n349), .S0(n274), .Y(n412) );
  MUX21X1_HVT U283 ( .A1(n437), .A2(n436), .S0(n267), .Y(n435) );
  MUX21X1_HVT U284 ( .A1(n556), .A2(n311), .S0(n274), .Y(n437) );
  MUX21X1_HVT U285 ( .A1(n567), .A2(n332), .S0(n268), .Y(n449) );
  MUX21X1_HVT U286 ( .A1(n360), .A2(n363), .S0(n217), .Y(n417) );
  MUX21X1_HVT U287 ( .A1(n363), .A2(n283), .S0(n218), .Y(n565) );
  MUX21X1_HVT U288 ( .A1(n334), .A2(n582), .S0(n264), .Y(n474) );
  MUX21X1_HVT U289 ( .A1(n533), .A2(n534), .S0(n272), .Y(n531) );
  MUX21X1_HVT U290 ( .A1(n283), .A2(n550), .S0(n271), .Y(n534) );
  XOR2X1_HVT U291 ( .A1(n292), .A2(n270), .Y(n542) );
  MUX21X1_HVT U292 ( .A1(n582), .A2(n50), .S0(n266), .Y(n456) );
  NBUFFX2_HVT U293 ( .A(n575), .Y(n285) );
  MUX21X1_HVT U294 ( .A1(n425), .A2(n426), .S0(n268), .Y(n424) );
  MUX21X1_HVT U295 ( .A1(n427), .A2(n290), .S0(n262), .Y(n426) );
  MUX21X1_HVT U296 ( .A1(n547), .A2(n352), .S0(n272), .Y(n425) );
  MUX21X1_HVT U297 ( .A1(n283), .A2(n360), .S0(n292), .Y(n372) );
  MUX21X1_HVT U298 ( .A1(n555), .A2(n376), .S0(n272), .Y(n370) );
  MUX21X1_HVT U299 ( .A1(n288), .A2(n283), .S0(n294), .Y(n576) );
  MUX21X1_HVT U300 ( .A1(n317), .A2(n50), .S0(n271), .Y(n519) );
  NBUFFX2_HVT U301 ( .A(n584), .Y(n291) );
  MUX21X1_HVT U302 ( .A1(n327), .A2(n555), .S0(n267), .Y(n452) );
  MUX21X1_HVT U303 ( .A1(n290), .A2(n493), .S0(n262), .Y(n492) );
  MUX21X1_HVT U304 ( .A1(n283), .A2(n280), .S0(n274), .Y(n493) );
  NBUFFX2_HVT U305 ( .A(n364), .Y(n280) );
  NBUFFX2_HVT U306 ( .A(n575), .Y(n286) );
  INVX1_HVT U307 ( .A(n298), .Y(n292) );
  XNOR2X1_HVT U308 ( .A1(n304), .A2(n218), .Y(n262) );
  INVX1_HVT U309 ( .A(n297), .Y(n296) );
  AND2X1_HVT U310 ( .A1(n275), .A2(n50), .Y(n263) );
  INVX0_HVT U311 ( .A(in[4]), .Y(n364) );
  MUX21X1_HVT U312 ( .A1(n491), .A2(n492), .S0(n268), .Y(n489) );
  MUX21X1_HVT U313 ( .A1(n359), .A2(n241), .S0(n294), .Y(n553) );
  MUX21X1_HVT U314 ( .A1(n241), .A2(n362), .S0(n292), .Y(n549) );
  NAND2X0_HVT U315 ( .A1(in[4]), .A2(n361), .Y(n575) );
  NAND2X0_HVT U316 ( .A1(in[3]), .A2(in[4]), .Y(n584) );
  MUX21X1_HVT U317 ( .A1(n241), .A2(n578), .S0(n295), .Y(n374) );
  MUX21X1_HVT U318 ( .A1(n241), .A2(n360), .S0(n296), .Y(n567) );
  MUX21X1_HVT U319 ( .A1(n241), .A2(n290), .S0(n217), .Y(n564) );
  MUX21X1_HVT U320 ( .A1(n241), .A2(n285), .S0(n292), .Y(n366) );
  MUX21X1_HVT U321 ( .A1(n241), .A2(n291), .S0(n218), .Y(n365) );
  MUX21X1_HVT U322 ( .A1(n291), .A2(n241), .S0(n293), .Y(n557) );
  MUX21X1_HVT U323 ( .A1(n283), .A2(n241), .S0(n265), .Y(n469) );
  MUX21X1_HVT U324 ( .A1(n275), .A2(n241), .S0(n292), .Y(n555) );
  NBUFFX2_HVT U325 ( .A(in[3]), .Y(n283) );
  NBUFFX2_HVT U326 ( .A(in[0]), .Y(n282) );
  INVX0_HVT U327 ( .A(n563), .Y(n305) );
  INVX0_HVT U328 ( .A(n561), .Y(n306) );
  INVX0_HVT U329 ( .A(n552), .Y(n307) );
  INVX0_HVT U330 ( .A(n550), .Y(n308) );
  INVX0_HVT U331 ( .A(n414), .Y(n309) );
  INVX0_HVT U332 ( .A(n377), .Y(n310) );
  INVX0_HVT U333 ( .A(n582), .Y(n311) );
  INVX0_HVT U334 ( .A(n569), .Y(n312) );
  INVX0_HVT U335 ( .A(n581), .Y(n313) );
  INVX0_HVT U336 ( .A(n577), .Y(n314) );
  INVX0_HVT U337 ( .A(n576), .Y(n315) );
  INVX0_HVT U338 ( .A(n574), .Y(n316) );
  INVX0_HVT U339 ( .A(n573), .Y(n317) );
  INVX0_HVT U340 ( .A(n570), .Y(n318) );
  INVX0_HVT U341 ( .A(n567), .Y(n320) );
  INVX0_HVT U342 ( .A(n566), .Y(n321) );
  INVX0_HVT U343 ( .A(n565), .Y(n322) );
  INVX0_HVT U344 ( .A(n564), .Y(n323) );
  INVX0_HVT U345 ( .A(n562), .Y(n324) );
  INVX0_HVT U346 ( .A(n560), .Y(n325) );
  INVX0_HVT U347 ( .A(n559), .Y(n326) );
  INVX0_HVT U348 ( .A(n557), .Y(n327) );
  INVX0_HVT U349 ( .A(n556), .Y(n328) );
  INVX0_HVT U350 ( .A(n555), .Y(n329) );
  INVX0_HVT U351 ( .A(n370), .Y(n330) );
  INVX0_HVT U352 ( .A(n554), .Y(n331) );
  INVX0_HVT U353 ( .A(n551), .Y(n333) );
  INVX0_HVT U354 ( .A(n547), .Y(n336) );
  INVX0_HVT U355 ( .A(n546), .Y(n337) );
  INVX0_HVT U356 ( .A(n545), .Y(n338) );
  INVX0_HVT U357 ( .A(n544), .Y(n339) );
  INVX0_HVT U358 ( .A(n511), .Y(n341) );
  INVX0_HVT U359 ( .A(n572), .Y(n342) );
  INVX0_HVT U360 ( .A(n471), .Y(n343) );
  INVX0_HVT U361 ( .A(n376), .Y(n344) );
  INVX0_HVT U362 ( .A(n528), .Y(n345) );
  INVX0_HVT U363 ( .A(n430), .Y(n346) );
  INVX0_HVT U364 ( .A(n375), .Y(n347) );
  INVX0_HVT U365 ( .A(n374), .Y(n348) );
  INVX0_HVT U366 ( .A(n372), .Y(n350) );
  INVX0_HVT U367 ( .A(n371), .Y(n351) );
  INVX0_HVT U368 ( .A(n490), .Y(n352) );
  INVX0_HVT U369 ( .A(n480), .Y(n353) );
  INVX0_HVT U370 ( .A(n369), .Y(n354) );
  INVX0_HVT U371 ( .A(n367), .Y(n356) );
  INVX0_HVT U372 ( .A(n365), .Y(n358) );
endmodule

