
module ram_dp_DATA_WIDTH4_ADDR_WIDTH4_0 ( clk, rst, write, a_addr, a_din, 
        b_din, b_dout );
  input [3:0] a_addr;
  input [3:0] a_din;
  input [3:0] b_din;
  output [15:0] b_dout;
  input clk, rst, write;
  wire   N17, N18, N19, N20, \mem[15][15] , \mem[15][14] , \mem[15][13] ,
         \mem[15][12] , \mem[15][11] , \mem[15][10] , \mem[15][9] ,
         \mem[15][8] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][15] ,
         \mem[14][14] , \mem[14][13] , \mem[14][12] , \mem[14][11] ,
         \mem[14][10] , \mem[14][9] , \mem[14][8] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][15] , \mem[13][14] , \mem[13][13] ,
         \mem[13][12] , \mem[13][11] , \mem[13][10] , \mem[13][9] ,
         \mem[13][8] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][15] ,
         \mem[12][14] , \mem[12][13] , \mem[12][12] , \mem[12][11] ,
         \mem[12][10] , \mem[12][9] , \mem[12][8] , \mem[12][7] , \mem[12][6] ,
         \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] , \mem[12][1] ,
         \mem[12][0] , \mem[11][15] , \mem[11][14] , \mem[11][13] ,
         \mem[11][12] , \mem[11][11] , \mem[11][10] , \mem[11][9] ,
         \mem[11][8] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][15] , \mem[9][14] , \mem[9][13] , \mem[9][12] ,
         \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] , \mem[9][7] ,
         \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] ,
         \mem[9][1] , \mem[9][0] , \mem[8][15] , \mem[8][14] , \mem[8][13] ,
         \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] , \mem[8][8] ,
         \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] , \mem[8][3] ,
         \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][15] , \mem[7][14] ,
         \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] ,
         \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][15] ,
         \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] ,
         \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][15] , \mem[3][14] , \mem[3][13] ,
         \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] ,
         \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] ,
         \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][15] ,
         \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N539, N540, N541, N542, N543, N544, N545, N546, N547,
         N548, N549, N550, N551, N552, N553, N554, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n302, n320, n338, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020;
  assign N17 = b_din[0];
  assign N18 = b_din[1];
  assign N19 = b_din[2];
  assign N20 = b_din[3];

  DFFNX1_HVT \b_dout_reg[15]  ( .D(N539), .CLK(clk), .Q(b_dout[15]) );
  DFFNX1_HVT \b_dout_reg[14]  ( .D(N540), .CLK(clk), .Q(b_dout[14]) );
  DFFNX1_HVT \b_dout_reg[13]  ( .D(N541), .CLK(clk), .Q(b_dout[13]) );
  DFFNX1_HVT \b_dout_reg[12]  ( .D(N542), .CLK(clk), .Q(b_dout[12]) );
  DFFNX1_HVT \b_dout_reg[11]  ( .D(N543), .CLK(clk), .Q(b_dout[11]) );
  DFFNX1_HVT \b_dout_reg[10]  ( .D(N544), .CLK(clk), .Q(b_dout[10]) );
  DFFNX1_HVT \b_dout_reg[9]  ( .D(N545), .CLK(clk), .Q(b_dout[9]) );
  DFFNX1_HVT \b_dout_reg[8]  ( .D(N546), .CLK(clk), .Q(b_dout[8]) );
  DFFNX1_HVT \b_dout_reg[7]  ( .D(N547), .CLK(clk), .Q(b_dout[7]) );
  DFFNX1_HVT \b_dout_reg[6]  ( .D(N548), .CLK(clk), .Q(b_dout[6]) );
  DFFNX1_HVT \b_dout_reg[5]  ( .D(N549), .CLK(clk), .Q(b_dout[5]) );
  DFFNX1_HVT \b_dout_reg[4]  ( .D(N550), .CLK(clk), .Q(b_dout[4]) );
  DFFNX1_HVT \b_dout_reg[3]  ( .D(N551), .CLK(clk), .Q(b_dout[3]) );
  DFFNX1_HVT \b_dout_reg[2]  ( .D(N552), .CLK(clk), .Q(b_dout[2]) );
  DFFNX1_HVT \b_dout_reg[1]  ( .D(N553), .CLK(clk), .Q(b_dout[1]) );
  DFFNX1_HVT \b_dout_reg[0]  ( .D(N554), .CLK(clk), .Q(b_dout[0]) );
  DFFNX1_HVT \mem_reg[15][15]  ( .D(n825), .CLK(clk), .Q(\mem[15][15] ) );
  DFFNX1_HVT \mem_reg[15][14]  ( .D(n824), .CLK(clk), .Q(\mem[15][14] ) );
  DFFNX1_HVT \mem_reg[15][13]  ( .D(n823), .CLK(clk), .Q(\mem[15][13] ) );
  DFFNX1_HVT \mem_reg[15][12]  ( .D(n822), .CLK(clk), .Q(\mem[15][12] ) );
  DFFNX1_HVT \mem_reg[15][11]  ( .D(n821), .CLK(clk), .Q(\mem[15][11] ) );
  DFFNX1_HVT \mem_reg[15][10]  ( .D(n820), .CLK(clk), .Q(\mem[15][10] ) );
  DFFNX1_HVT \mem_reg[15][9]  ( .D(n819), .CLK(clk), .Q(\mem[15][9] ) );
  DFFNX1_HVT \mem_reg[15][8]  ( .D(n818), .CLK(clk), .Q(\mem[15][8] ) );
  DFFNX1_HVT \mem_reg[15][7]  ( .D(n817), .CLK(clk), .Q(\mem[15][7] ) );
  DFFNX1_HVT \mem_reg[15][6]  ( .D(n816), .CLK(clk), .Q(\mem[15][6] ) );
  DFFNX1_HVT \mem_reg[15][5]  ( .D(n815), .CLK(clk), .Q(\mem[15][5] ) );
  DFFNX1_HVT \mem_reg[15][4]  ( .D(n814), .CLK(clk), .Q(\mem[15][4] ) );
  DFFNX1_HVT \mem_reg[15][3]  ( .D(n813), .CLK(clk), .Q(\mem[15][3] ) );
  DFFNX1_HVT \mem_reg[15][2]  ( .D(n812), .CLK(clk), .Q(\mem[15][2] ) );
  DFFNX1_HVT \mem_reg[15][1]  ( .D(n811), .CLK(clk), .Q(\mem[15][1] ) );
  DFFNX1_HVT \mem_reg[15][0]  ( .D(n810), .CLK(clk), .Q(\mem[15][0] ) );
  DFFNX1_HVT \mem_reg[14][15]  ( .D(n809), .CLK(clk), .Q(\mem[14][15] ) );
  DFFNX1_HVT \mem_reg[14][14]  ( .D(n808), .CLK(clk), .Q(\mem[14][14] ) );
  DFFNX1_HVT \mem_reg[14][13]  ( .D(n807), .CLK(clk), .Q(\mem[14][13] ) );
  DFFNX1_HVT \mem_reg[14][12]  ( .D(n806), .CLK(clk), .Q(\mem[14][12] ) );
  DFFNX1_HVT \mem_reg[14][11]  ( .D(n805), .CLK(clk), .Q(\mem[14][11] ) );
  DFFNX1_HVT \mem_reg[14][10]  ( .D(n804), .CLK(clk), .Q(\mem[14][10] ) );
  DFFNX1_HVT \mem_reg[14][9]  ( .D(n803), .CLK(clk), .Q(\mem[14][9] ) );
  DFFNX1_HVT \mem_reg[14][8]  ( .D(n802), .CLK(clk), .Q(\mem[14][8] ) );
  DFFNX1_HVT \mem_reg[14][7]  ( .D(n801), .CLK(clk), .Q(\mem[14][7] ) );
  DFFNX1_HVT \mem_reg[14][6]  ( .D(n800), .CLK(clk), .Q(\mem[14][6] ) );
  DFFNX1_HVT \mem_reg[14][5]  ( .D(n799), .CLK(clk), .Q(\mem[14][5] ) );
  DFFNX1_HVT \mem_reg[14][4]  ( .D(n798), .CLK(clk), .Q(\mem[14][4] ) );
  DFFNX1_HVT \mem_reg[14][3]  ( .D(n797), .CLK(clk), .Q(\mem[14][3] ) );
  DFFNX1_HVT \mem_reg[14][2]  ( .D(n796), .CLK(clk), .Q(\mem[14][2] ) );
  DFFNX1_HVT \mem_reg[14][1]  ( .D(n795), .CLK(clk), .Q(\mem[14][1] ) );
  DFFNX1_HVT \mem_reg[14][0]  ( .D(n794), .CLK(clk), .Q(\mem[14][0] ) );
  DFFNX1_HVT \mem_reg[13][15]  ( .D(n793), .CLK(clk), .Q(\mem[13][15] ) );
  DFFNX1_HVT \mem_reg[13][14]  ( .D(n792), .CLK(clk), .Q(\mem[13][14] ) );
  DFFNX1_HVT \mem_reg[13][13]  ( .D(n791), .CLK(clk), .Q(\mem[13][13] ) );
  DFFNX1_HVT \mem_reg[13][12]  ( .D(n790), .CLK(clk), .Q(\mem[13][12] ) );
  DFFNX1_HVT \mem_reg[13][11]  ( .D(n789), .CLK(clk), .Q(\mem[13][11] ) );
  DFFNX1_HVT \mem_reg[13][10]  ( .D(n788), .CLK(clk), .Q(\mem[13][10] ) );
  DFFNX1_HVT \mem_reg[13][9]  ( .D(n787), .CLK(clk), .Q(\mem[13][9] ) );
  DFFNX1_HVT \mem_reg[13][8]  ( .D(n786), .CLK(clk), .Q(\mem[13][8] ) );
  DFFNX1_HVT \mem_reg[13][7]  ( .D(n785), .CLK(clk), .Q(\mem[13][7] ) );
  DFFNX1_HVT \mem_reg[13][6]  ( .D(n784), .CLK(clk), .Q(\mem[13][6] ) );
  DFFNX1_HVT \mem_reg[13][5]  ( .D(n783), .CLK(clk), .Q(\mem[13][5] ) );
  DFFNX1_HVT \mem_reg[13][4]  ( .D(n782), .CLK(clk), .Q(\mem[13][4] ) );
  DFFNX1_HVT \mem_reg[13][3]  ( .D(n781), .CLK(clk), .Q(\mem[13][3] ) );
  DFFNX1_HVT \mem_reg[13][2]  ( .D(n780), .CLK(clk), .Q(\mem[13][2] ) );
  DFFNX1_HVT \mem_reg[13][1]  ( .D(n779), .CLK(clk), .Q(\mem[13][1] ) );
  DFFNX1_HVT \mem_reg[13][0]  ( .D(n778), .CLK(clk), .Q(\mem[13][0] ) );
  DFFNX1_HVT \mem_reg[12][15]  ( .D(n777), .CLK(clk), .Q(\mem[12][15] ) );
  DFFNX1_HVT \mem_reg[12][14]  ( .D(n776), .CLK(clk), .Q(\mem[12][14] ) );
  DFFNX1_HVT \mem_reg[12][13]  ( .D(n775), .CLK(clk), .Q(\mem[12][13] ) );
  DFFNX1_HVT \mem_reg[12][12]  ( .D(n774), .CLK(clk), .Q(\mem[12][12] ) );
  DFFNX1_HVT \mem_reg[12][11]  ( .D(n773), .CLK(clk), .Q(\mem[12][11] ) );
  DFFNX1_HVT \mem_reg[12][10]  ( .D(n772), .CLK(clk), .Q(\mem[12][10] ) );
  DFFNX1_HVT \mem_reg[12][9]  ( .D(n771), .CLK(clk), .Q(\mem[12][9] ) );
  DFFNX1_HVT \mem_reg[12][8]  ( .D(n770), .CLK(clk), .Q(\mem[12][8] ) );
  DFFNX1_HVT \mem_reg[12][7]  ( .D(n769), .CLK(clk), .Q(\mem[12][7] ) );
  DFFNX1_HVT \mem_reg[12][6]  ( .D(n768), .CLK(clk), .Q(\mem[12][6] ) );
  DFFNX1_HVT \mem_reg[12][5]  ( .D(n767), .CLK(clk), .Q(\mem[12][5] ) );
  DFFNX1_HVT \mem_reg[12][4]  ( .D(n766), .CLK(clk), .Q(\mem[12][4] ) );
  DFFNX1_HVT \mem_reg[12][3]  ( .D(n765), .CLK(clk), .Q(\mem[12][3] ) );
  DFFNX1_HVT \mem_reg[12][2]  ( .D(n764), .CLK(clk), .Q(\mem[12][2] ) );
  DFFNX1_HVT \mem_reg[12][1]  ( .D(n763), .CLK(clk), .Q(\mem[12][1] ) );
  DFFNX1_HVT \mem_reg[12][0]  ( .D(n762), .CLK(clk), .Q(\mem[12][0] ) );
  DFFNX1_HVT \mem_reg[11][15]  ( .D(n761), .CLK(clk), .Q(\mem[11][15] ) );
  DFFNX1_HVT \mem_reg[11][14]  ( .D(n760), .CLK(clk), .Q(\mem[11][14] ) );
  DFFNX1_HVT \mem_reg[11][13]  ( .D(n759), .CLK(clk), .Q(\mem[11][13] ) );
  DFFNX1_HVT \mem_reg[11][12]  ( .D(n758), .CLK(clk), .Q(\mem[11][12] ) );
  DFFNX1_HVT \mem_reg[11][11]  ( .D(n757), .CLK(clk), .Q(\mem[11][11] ) );
  DFFNX1_HVT \mem_reg[11][10]  ( .D(n756), .CLK(clk), .Q(\mem[11][10] ) );
  DFFNX1_HVT \mem_reg[11][9]  ( .D(n755), .CLK(clk), .Q(\mem[11][9] ) );
  DFFNX1_HVT \mem_reg[11][8]  ( .D(n754), .CLK(clk), .Q(\mem[11][8] ) );
  DFFNX1_HVT \mem_reg[11][7]  ( .D(n753), .CLK(clk), .Q(\mem[11][7] ) );
  DFFNX1_HVT \mem_reg[11][6]  ( .D(n752), .CLK(clk), .Q(\mem[11][6] ) );
  DFFNX1_HVT \mem_reg[11][5]  ( .D(n751), .CLK(clk), .Q(\mem[11][5] ) );
  DFFNX1_HVT \mem_reg[11][4]  ( .D(n750), .CLK(clk), .Q(\mem[11][4] ) );
  DFFNX1_HVT \mem_reg[11][3]  ( .D(n749), .CLK(clk), .Q(\mem[11][3] ) );
  DFFNX1_HVT \mem_reg[11][2]  ( .D(n748), .CLK(clk), .Q(\mem[11][2] ) );
  DFFNX1_HVT \mem_reg[11][1]  ( .D(n747), .CLK(clk), .Q(\mem[11][1] ) );
  DFFNX1_HVT \mem_reg[11][0]  ( .D(n746), .CLK(clk), .Q(\mem[11][0] ) );
  DFFNX1_HVT \mem_reg[10][15]  ( .D(n745), .CLK(clk), .Q(\mem[10][15] ) );
  DFFNX1_HVT \mem_reg[10][14]  ( .D(n744), .CLK(clk), .Q(\mem[10][14] ) );
  DFFNX1_HVT \mem_reg[10][13]  ( .D(n743), .CLK(clk), .Q(\mem[10][13] ) );
  DFFNX1_HVT \mem_reg[10][12]  ( .D(n742), .CLK(clk), .Q(\mem[10][12] ) );
  DFFNX1_HVT \mem_reg[10][11]  ( .D(n741), .CLK(clk), .Q(\mem[10][11] ) );
  DFFNX1_HVT \mem_reg[10][10]  ( .D(n740), .CLK(clk), .Q(\mem[10][10] ) );
  DFFNX1_HVT \mem_reg[10][9]  ( .D(n739), .CLK(clk), .Q(\mem[10][9] ) );
  DFFNX1_HVT \mem_reg[10][8]  ( .D(n738), .CLK(clk), .Q(\mem[10][8] ) );
  DFFNX1_HVT \mem_reg[10][7]  ( .D(n737), .CLK(clk), .Q(\mem[10][7] ) );
  DFFNX1_HVT \mem_reg[10][6]  ( .D(n736), .CLK(clk), .Q(\mem[10][6] ) );
  DFFNX1_HVT \mem_reg[10][5]  ( .D(n735), .CLK(clk), .Q(\mem[10][5] ) );
  DFFNX1_HVT \mem_reg[10][4]  ( .D(n734), .CLK(clk), .Q(\mem[10][4] ) );
  DFFNX1_HVT \mem_reg[10][3]  ( .D(n733), .CLK(clk), .Q(\mem[10][3] ) );
  DFFNX1_HVT \mem_reg[10][2]  ( .D(n732), .CLK(clk), .Q(\mem[10][2] ) );
  DFFNX1_HVT \mem_reg[10][1]  ( .D(n731), .CLK(clk), .Q(\mem[10][1] ) );
  DFFNX1_HVT \mem_reg[10][0]  ( .D(n730), .CLK(clk), .Q(\mem[10][0] ) );
  DFFNX1_HVT \mem_reg[9][15]  ( .D(n729), .CLK(clk), .Q(\mem[9][15] ) );
  DFFNX1_HVT \mem_reg[9][14]  ( .D(n728), .CLK(clk), .Q(\mem[9][14] ) );
  DFFNX1_HVT \mem_reg[9][13]  ( .D(n727), .CLK(clk), .Q(\mem[9][13] ) );
  DFFNX1_HVT \mem_reg[9][12]  ( .D(n726), .CLK(clk), .Q(\mem[9][12] ) );
  DFFNX1_HVT \mem_reg[9][11]  ( .D(n725), .CLK(clk), .Q(\mem[9][11] ) );
  DFFNX1_HVT \mem_reg[9][10]  ( .D(n724), .CLK(clk), .Q(\mem[9][10] ) );
  DFFNX1_HVT \mem_reg[9][9]  ( .D(n723), .CLK(clk), .Q(\mem[9][9] ) );
  DFFNX1_HVT \mem_reg[9][8]  ( .D(n722), .CLK(clk), .Q(\mem[9][8] ) );
  DFFNX1_HVT \mem_reg[9][7]  ( .D(n721), .CLK(clk), .Q(\mem[9][7] ) );
  DFFNX1_HVT \mem_reg[9][6]  ( .D(n720), .CLK(clk), .Q(\mem[9][6] ) );
  DFFNX1_HVT \mem_reg[9][5]  ( .D(n719), .CLK(clk), .Q(\mem[9][5] ) );
  DFFNX1_HVT \mem_reg[9][4]  ( .D(n718), .CLK(clk), .Q(\mem[9][4] ) );
  DFFNX1_HVT \mem_reg[9][3]  ( .D(n717), .CLK(clk), .Q(\mem[9][3] ) );
  DFFNX1_HVT \mem_reg[9][2]  ( .D(n716), .CLK(clk), .Q(\mem[9][2] ) );
  DFFNX1_HVT \mem_reg[9][1]  ( .D(n715), .CLK(clk), .Q(\mem[9][1] ) );
  DFFNX1_HVT \mem_reg[9][0]  ( .D(n714), .CLK(clk), .Q(\mem[9][0] ) );
  DFFNX1_HVT \mem_reg[8][15]  ( .D(n713), .CLK(clk), .Q(\mem[8][15] ) );
  DFFNX1_HVT \mem_reg[8][14]  ( .D(n712), .CLK(clk), .Q(\mem[8][14] ) );
  DFFNX1_HVT \mem_reg[8][13]  ( .D(n711), .CLK(clk), .Q(\mem[8][13] ) );
  DFFNX1_HVT \mem_reg[8][12]  ( .D(n710), .CLK(clk), .Q(\mem[8][12] ) );
  DFFNX1_HVT \mem_reg[8][11]  ( .D(n709), .CLK(clk), .Q(\mem[8][11] ) );
  DFFNX1_HVT \mem_reg[8][10]  ( .D(n708), .CLK(clk), .Q(\mem[8][10] ) );
  DFFNX1_HVT \mem_reg[8][9]  ( .D(n707), .CLK(clk), .Q(\mem[8][9] ) );
  DFFNX1_HVT \mem_reg[8][8]  ( .D(n706), .CLK(clk), .Q(\mem[8][8] ) );
  DFFNX1_HVT \mem_reg[8][7]  ( .D(n705), .CLK(clk), .Q(\mem[8][7] ) );
  DFFNX1_HVT \mem_reg[8][6]  ( .D(n704), .CLK(clk), .Q(\mem[8][6] ) );
  DFFNX1_HVT \mem_reg[8][5]  ( .D(n703), .CLK(clk), .Q(\mem[8][5] ) );
  DFFNX1_HVT \mem_reg[8][4]  ( .D(n702), .CLK(clk), .Q(\mem[8][4] ) );
  DFFNX1_HVT \mem_reg[8][3]  ( .D(n701), .CLK(clk), .Q(\mem[8][3] ) );
  DFFNX1_HVT \mem_reg[8][2]  ( .D(n700), .CLK(clk), .Q(\mem[8][2] ) );
  DFFNX1_HVT \mem_reg[8][1]  ( .D(n699), .CLK(clk), .Q(\mem[8][1] ) );
  DFFNX1_HVT \mem_reg[8][0]  ( .D(n698), .CLK(clk), .Q(\mem[8][0] ) );
  DFFNX1_HVT \mem_reg[7][15]  ( .D(n697), .CLK(clk), .Q(\mem[7][15] ) );
  DFFNX1_HVT \mem_reg[7][14]  ( .D(n696), .CLK(clk), .Q(\mem[7][14] ) );
  DFFNX1_HVT \mem_reg[7][13]  ( .D(n695), .CLK(clk), .Q(\mem[7][13] ) );
  DFFNX1_HVT \mem_reg[7][12]  ( .D(n694), .CLK(clk), .Q(\mem[7][12] ) );
  DFFNX1_HVT \mem_reg[7][11]  ( .D(n693), .CLK(clk), .Q(\mem[7][11] ) );
  DFFNX1_HVT \mem_reg[7][10]  ( .D(n692), .CLK(clk), .Q(\mem[7][10] ) );
  DFFNX1_HVT \mem_reg[7][9]  ( .D(n691), .CLK(clk), .Q(\mem[7][9] ) );
  DFFNX1_HVT \mem_reg[7][8]  ( .D(n690), .CLK(clk), .Q(\mem[7][8] ) );
  DFFNX1_HVT \mem_reg[7][7]  ( .D(n689), .CLK(clk), .Q(\mem[7][7] ) );
  DFFNX1_HVT \mem_reg[7][6]  ( .D(n688), .CLK(clk), .Q(\mem[7][6] ) );
  DFFNX1_HVT \mem_reg[7][5]  ( .D(n687), .CLK(clk), .Q(\mem[7][5] ) );
  DFFNX1_HVT \mem_reg[7][4]  ( .D(n686), .CLK(clk), .Q(\mem[7][4] ) );
  DFFNX1_HVT \mem_reg[7][3]  ( .D(n685), .CLK(clk), .Q(\mem[7][3] ) );
  DFFNX1_HVT \mem_reg[7][2]  ( .D(n684), .CLK(clk), .Q(\mem[7][2] ) );
  DFFNX1_HVT \mem_reg[7][1]  ( .D(n683), .CLK(clk), .Q(\mem[7][1] ) );
  DFFNX1_HVT \mem_reg[7][0]  ( .D(n682), .CLK(clk), .Q(\mem[7][0] ) );
  DFFNX1_HVT \mem_reg[6][15]  ( .D(n681), .CLK(clk), .Q(\mem[6][15] ) );
  DFFNX1_HVT \mem_reg[6][14]  ( .D(n680), .CLK(clk), .Q(\mem[6][14] ) );
  DFFNX1_HVT \mem_reg[6][13]  ( .D(n679), .CLK(clk), .Q(\mem[6][13] ) );
  DFFNX1_HVT \mem_reg[6][12]  ( .D(n678), .CLK(clk), .Q(\mem[6][12] ) );
  DFFNX1_HVT \mem_reg[6][11]  ( .D(n677), .CLK(clk), .Q(\mem[6][11] ) );
  DFFNX1_HVT \mem_reg[6][10]  ( .D(n676), .CLK(clk), .Q(\mem[6][10] ) );
  DFFNX1_HVT \mem_reg[6][9]  ( .D(n675), .CLK(clk), .Q(\mem[6][9] ) );
  DFFNX1_HVT \mem_reg[6][8]  ( .D(n674), .CLK(clk), .Q(\mem[6][8] ) );
  DFFNX1_HVT \mem_reg[6][7]  ( .D(n673), .CLK(clk), .Q(\mem[6][7] ) );
  DFFNX1_HVT \mem_reg[6][6]  ( .D(n672), .CLK(clk), .Q(\mem[6][6] ) );
  DFFNX1_HVT \mem_reg[6][5]  ( .D(n671), .CLK(clk), .Q(\mem[6][5] ) );
  DFFNX1_HVT \mem_reg[6][4]  ( .D(n670), .CLK(clk), .Q(\mem[6][4] ) );
  DFFNX1_HVT \mem_reg[6][3]  ( .D(n669), .CLK(clk), .Q(\mem[6][3] ) );
  DFFNX1_HVT \mem_reg[6][2]  ( .D(n668), .CLK(clk), .Q(\mem[6][2] ) );
  DFFNX1_HVT \mem_reg[6][1]  ( .D(n667), .CLK(clk), .Q(\mem[6][1] ) );
  DFFNX1_HVT \mem_reg[6][0]  ( .D(n666), .CLK(clk), .Q(\mem[6][0] ) );
  DFFNX1_HVT \mem_reg[5][15]  ( .D(n665), .CLK(clk), .Q(\mem[5][15] ) );
  DFFNX1_HVT \mem_reg[5][14]  ( .D(n664), .CLK(clk), .Q(\mem[5][14] ) );
  DFFNX1_HVT \mem_reg[5][13]  ( .D(n663), .CLK(clk), .Q(\mem[5][13] ) );
  DFFNX1_HVT \mem_reg[5][12]  ( .D(n662), .CLK(clk), .Q(\mem[5][12] ) );
  DFFNX1_HVT \mem_reg[5][11]  ( .D(n661), .CLK(clk), .Q(\mem[5][11] ) );
  DFFNX1_HVT \mem_reg[5][10]  ( .D(n660), .CLK(clk), .Q(\mem[5][10] ) );
  DFFNX1_HVT \mem_reg[5][9]  ( .D(n659), .CLK(clk), .Q(\mem[5][9] ) );
  DFFNX1_HVT \mem_reg[5][8]  ( .D(n658), .CLK(clk), .Q(\mem[5][8] ) );
  DFFNX1_HVT \mem_reg[5][7]  ( .D(n657), .CLK(clk), .Q(\mem[5][7] ) );
  DFFNX1_HVT \mem_reg[5][6]  ( .D(n656), .CLK(clk), .Q(\mem[5][6] ) );
  DFFNX1_HVT \mem_reg[5][5]  ( .D(n655), .CLK(clk), .Q(\mem[5][5] ) );
  DFFNX1_HVT \mem_reg[5][4]  ( .D(n654), .CLK(clk), .Q(\mem[5][4] ) );
  DFFNX1_HVT \mem_reg[5][3]  ( .D(n653), .CLK(clk), .Q(\mem[5][3] ) );
  DFFNX1_HVT \mem_reg[5][2]  ( .D(n652), .CLK(clk), .Q(\mem[5][2] ) );
  DFFNX1_HVT \mem_reg[5][1]  ( .D(n651), .CLK(clk), .Q(\mem[5][1] ) );
  DFFNX1_HVT \mem_reg[5][0]  ( .D(n650), .CLK(clk), .Q(\mem[5][0] ) );
  DFFNX1_HVT \mem_reg[4][15]  ( .D(n649), .CLK(clk), .Q(\mem[4][15] ) );
  DFFNX1_HVT \mem_reg[4][14]  ( .D(n648), .CLK(clk), .Q(\mem[4][14] ) );
  DFFNX1_HVT \mem_reg[4][13]  ( .D(n647), .CLK(clk), .Q(\mem[4][13] ) );
  DFFNX1_HVT \mem_reg[4][12]  ( .D(n646), .CLK(clk), .Q(\mem[4][12] ) );
  DFFNX1_HVT \mem_reg[4][11]  ( .D(n645), .CLK(clk), .Q(\mem[4][11] ) );
  DFFNX1_HVT \mem_reg[4][10]  ( .D(n644), .CLK(clk), .Q(\mem[4][10] ) );
  DFFNX1_HVT \mem_reg[4][9]  ( .D(n643), .CLK(clk), .Q(\mem[4][9] ) );
  DFFNX1_HVT \mem_reg[4][8]  ( .D(n642), .CLK(clk), .Q(\mem[4][8] ) );
  DFFNX1_HVT \mem_reg[4][7]  ( .D(n641), .CLK(clk), .Q(\mem[4][7] ) );
  DFFNX1_HVT \mem_reg[4][6]  ( .D(n640), .CLK(clk), .Q(\mem[4][6] ) );
  DFFNX1_HVT \mem_reg[4][5]  ( .D(n639), .CLK(clk), .Q(\mem[4][5] ) );
  DFFNX1_HVT \mem_reg[4][4]  ( .D(n638), .CLK(clk), .Q(\mem[4][4] ) );
  DFFNX1_HVT \mem_reg[4][3]  ( .D(n637), .CLK(clk), .Q(\mem[4][3] ) );
  DFFNX1_HVT \mem_reg[4][2]  ( .D(n636), .CLK(clk), .Q(\mem[4][2] ) );
  DFFNX1_HVT \mem_reg[4][1]  ( .D(n635), .CLK(clk), .Q(\mem[4][1] ) );
  DFFNX1_HVT \mem_reg[4][0]  ( .D(n634), .CLK(clk), .Q(\mem[4][0] ) );
  DFFNX1_HVT \mem_reg[3][15]  ( .D(n633), .CLK(clk), .Q(\mem[3][15] ) );
  DFFNX1_HVT \mem_reg[3][14]  ( .D(n632), .CLK(clk), .Q(\mem[3][14] ) );
  DFFNX1_HVT \mem_reg[3][13]  ( .D(n631), .CLK(clk), .Q(\mem[3][13] ) );
  DFFNX1_HVT \mem_reg[3][12]  ( .D(n630), .CLK(clk), .Q(\mem[3][12] ) );
  DFFNX1_HVT \mem_reg[3][11]  ( .D(n629), .CLK(clk), .Q(\mem[3][11] ) );
  DFFNX1_HVT \mem_reg[3][10]  ( .D(n628), .CLK(clk), .Q(\mem[3][10] ) );
  DFFNX1_HVT \mem_reg[3][9]  ( .D(n627), .CLK(clk), .Q(\mem[3][9] ) );
  DFFNX1_HVT \mem_reg[3][8]  ( .D(n626), .CLK(clk), .Q(\mem[3][8] ) );
  DFFNX1_HVT \mem_reg[3][7]  ( .D(n625), .CLK(clk), .Q(\mem[3][7] ) );
  DFFNX1_HVT \mem_reg[3][6]  ( .D(n624), .CLK(clk), .Q(\mem[3][6] ) );
  DFFNX1_HVT \mem_reg[3][5]  ( .D(n623), .CLK(clk), .Q(\mem[3][5] ) );
  DFFNX1_HVT \mem_reg[3][4]  ( .D(n622), .CLK(clk), .Q(\mem[3][4] ) );
  DFFNX1_HVT \mem_reg[3][3]  ( .D(n621), .CLK(clk), .Q(\mem[3][3] ) );
  DFFNX1_HVT \mem_reg[3][2]  ( .D(n620), .CLK(clk), .Q(\mem[3][2] ) );
  DFFNX1_HVT \mem_reg[3][1]  ( .D(n619), .CLK(clk), .Q(\mem[3][1] ) );
  DFFNX1_HVT \mem_reg[3][0]  ( .D(n618), .CLK(clk), .Q(\mem[3][0] ) );
  DFFNX1_HVT \mem_reg[2][15]  ( .D(n617), .CLK(clk), .Q(\mem[2][15] ) );
  DFFNX1_HVT \mem_reg[2][14]  ( .D(n616), .CLK(clk), .Q(\mem[2][14] ) );
  DFFNX1_HVT \mem_reg[2][13]  ( .D(n615), .CLK(clk), .Q(\mem[2][13] ) );
  DFFNX1_HVT \mem_reg[2][12]  ( .D(n614), .CLK(clk), .Q(\mem[2][12] ) );
  DFFNX1_HVT \mem_reg[2][11]  ( .D(n613), .CLK(clk), .Q(\mem[2][11] ) );
  DFFNX1_HVT \mem_reg[2][10]  ( .D(n612), .CLK(clk), .Q(\mem[2][10] ) );
  DFFNX1_HVT \mem_reg[2][9]  ( .D(n611), .CLK(clk), .Q(\mem[2][9] ) );
  DFFNX1_HVT \mem_reg[2][8]  ( .D(n610), .CLK(clk), .Q(\mem[2][8] ) );
  DFFNX1_HVT \mem_reg[2][7]  ( .D(n609), .CLK(clk), .Q(\mem[2][7] ) );
  DFFNX1_HVT \mem_reg[2][6]  ( .D(n608), .CLK(clk), .Q(\mem[2][6] ) );
  DFFNX1_HVT \mem_reg[2][5]  ( .D(n607), .CLK(clk), .Q(\mem[2][5] ) );
  DFFNX1_HVT \mem_reg[2][4]  ( .D(n606), .CLK(clk), .Q(\mem[2][4] ) );
  DFFNX1_HVT \mem_reg[2][3]  ( .D(n605), .CLK(clk), .Q(\mem[2][3] ) );
  DFFNX1_HVT \mem_reg[2][2]  ( .D(n604), .CLK(clk), .Q(\mem[2][2] ) );
  DFFNX1_HVT \mem_reg[2][1]  ( .D(n603), .CLK(clk), .Q(\mem[2][1] ) );
  DFFNX1_HVT \mem_reg[2][0]  ( .D(n602), .CLK(clk), .Q(\mem[2][0] ) );
  DFFNX1_HVT \mem_reg[1][15]  ( .D(n601), .CLK(clk), .Q(\mem[1][15] ) );
  DFFNX1_HVT \mem_reg[1][14]  ( .D(n600), .CLK(clk), .Q(\mem[1][14] ) );
  DFFNX1_HVT \mem_reg[1][13]  ( .D(n599), .CLK(clk), .Q(\mem[1][13] ) );
  DFFNX1_HVT \mem_reg[1][12]  ( .D(n598), .CLK(clk), .Q(\mem[1][12] ) );
  DFFNX1_HVT \mem_reg[1][11]  ( .D(n597), .CLK(clk), .Q(\mem[1][11] ) );
  DFFNX1_HVT \mem_reg[1][10]  ( .D(n596), .CLK(clk), .Q(\mem[1][10] ) );
  DFFNX1_HVT \mem_reg[1][9]  ( .D(n595), .CLK(clk), .Q(\mem[1][9] ) );
  DFFNX1_HVT \mem_reg[1][8]  ( .D(n594), .CLK(clk), .Q(\mem[1][8] ) );
  DFFNX1_HVT \mem_reg[1][7]  ( .D(n593), .CLK(clk), .Q(\mem[1][7] ) );
  DFFNX1_HVT \mem_reg[1][6]  ( .D(n592), .CLK(clk), .Q(\mem[1][6] ) );
  DFFNX1_HVT \mem_reg[1][5]  ( .D(n591), .CLK(clk), .Q(\mem[1][5] ) );
  DFFNX1_HVT \mem_reg[1][4]  ( .D(n590), .CLK(clk), .Q(\mem[1][4] ) );
  DFFNX1_HVT \mem_reg[1][3]  ( .D(n589), .CLK(clk), .Q(\mem[1][3] ) );
  DFFNX1_HVT \mem_reg[1][2]  ( .D(n588), .CLK(clk), .Q(\mem[1][2] ) );
  DFFNX1_HVT \mem_reg[1][1]  ( .D(n587), .CLK(clk), .Q(\mem[1][1] ) );
  DFFNX1_HVT \mem_reg[1][0]  ( .D(n586), .CLK(clk), .Q(\mem[1][0] ) );
  DFFNX1_HVT \mem_reg[0][15]  ( .D(n585), .CLK(clk), .Q(\mem[0][15] ) );
  DFFNX1_HVT \mem_reg[0][14]  ( .D(n584), .CLK(clk), .Q(\mem[0][14] ) );
  DFFNX1_HVT \mem_reg[0][13]  ( .D(n583), .CLK(clk), .Q(\mem[0][13] ) );
  DFFNX1_HVT \mem_reg[0][12]  ( .D(n582), .CLK(clk), .Q(\mem[0][12] ) );
  DFFNX1_HVT \mem_reg[0][11]  ( .D(n581), .CLK(clk), .Q(\mem[0][11] ) );
  DFFNX1_HVT \mem_reg[0][10]  ( .D(n580), .CLK(clk), .Q(\mem[0][10] ) );
  DFFNX1_HVT \mem_reg[0][9]  ( .D(n579), .CLK(clk), .Q(\mem[0][9] ) );
  DFFNX1_HVT \mem_reg[0][8]  ( .D(n578), .CLK(clk), .Q(\mem[0][8] ) );
  DFFNX1_HVT \mem_reg[0][7]  ( .D(n577), .CLK(clk), .Q(\mem[0][7] ) );
  DFFNX1_HVT \mem_reg[0][6]  ( .D(n576), .CLK(clk), .Q(\mem[0][6] ) );
  DFFNX1_HVT \mem_reg[0][5]  ( .D(n575), .CLK(clk), .Q(\mem[0][5] ) );
  DFFNX1_HVT \mem_reg[0][4]  ( .D(n574), .CLK(clk), .Q(\mem[0][4] ) );
  DFFNX1_HVT \mem_reg[0][3]  ( .D(n573), .CLK(clk), .Q(\mem[0][3] ) );
  DFFNX1_HVT \mem_reg[0][2]  ( .D(n572), .CLK(clk), .Q(\mem[0][2] ) );
  DFFNX1_HVT \mem_reg[0][1]  ( .D(n571), .CLK(clk), .Q(\mem[0][1] ) );
  DFFNX1_HVT \mem_reg[0][0]  ( .D(n570), .CLK(clk), .Q(\mem[0][0] ) );
  AO22X1_HVT U268 ( .A1(n266), .A2(n186), .A3(\mem[0][0] ), .A4(n890), .Y(n570) );
  AO21X1_HVT U269 ( .A1(n267), .A2(n147), .A3(n162), .Y(n266) );
  AO22X1_HVT U270 ( .A1(n269), .A2(n186), .A3(\mem[0][1] ), .A4(n889), .Y(n571) );
  AO21X1_HVT U271 ( .A1(n270), .A2(n149), .A3(n163), .Y(n269) );
  AO22X1_HVT U272 ( .A1(n271), .A2(n186), .A3(\mem[0][2] ), .A4(n888), .Y(n572) );
  AO21X1_HVT U273 ( .A1(n272), .A2(n148), .A3(n180), .Y(n271) );
  AO22X1_HVT U274 ( .A1(n273), .A2(n186), .A3(\mem[0][3] ), .A4(n887), .Y(n573) );
  AO21X1_HVT U275 ( .A1(n274), .A2(n147), .A3(n163), .Y(n273) );
  AO22X1_HVT U276 ( .A1(n275), .A2(n186), .A3(\mem[0][4] ), .A4(n886), .Y(n574) );
  AO21X1_HVT U277 ( .A1(n276), .A2(n149), .A3(n163), .Y(n275) );
  AO22X1_HVT U278 ( .A1(n277), .A2(n186), .A3(\mem[0][5] ), .A4(n885), .Y(n575) );
  AO21X1_HVT U279 ( .A1(n278), .A2(n148), .A3(n163), .Y(n277) );
  AO22X1_HVT U280 ( .A1(n279), .A2(n186), .A3(\mem[0][6] ), .A4(n884), .Y(n576) );
  AO21X1_HVT U281 ( .A1(n280), .A2(n147), .A3(n163), .Y(n279) );
  AO22X1_HVT U282 ( .A1(n281), .A2(n186), .A3(\mem[0][7] ), .A4(n883), .Y(n577) );
  AO21X1_HVT U283 ( .A1(n282), .A2(n149), .A3(n163), .Y(n281) );
  AO22X1_HVT U284 ( .A1(n283), .A2(n186), .A3(\mem[0][8] ), .A4(n882), .Y(n578) );
  AO21X1_HVT U285 ( .A1(n284), .A2(n148), .A3(n163), .Y(n283) );
  AO22X1_HVT U286 ( .A1(n285), .A2(n186), .A3(\mem[0][9] ), .A4(n881), .Y(n579) );
  AO21X1_HVT U287 ( .A1(n286), .A2(n147), .A3(n164), .Y(n285) );
  AO22X1_HVT U288 ( .A1(n287), .A2(n186), .A3(\mem[0][10] ), .A4(n880), .Y(
        n580) );
  AO21X1_HVT U289 ( .A1(n288), .A2(n149), .A3(n164), .Y(n287) );
  AO22X1_HVT U290 ( .A1(n289), .A2(n186), .A3(\mem[0][11] ), .A4(n879), .Y(
        n581) );
  AO21X1_HVT U291 ( .A1(n290), .A2(n148), .A3(n164), .Y(n289) );
  AO22X1_HVT U292 ( .A1(n291), .A2(n187), .A3(\mem[0][12] ), .A4(n878), .Y(
        n582) );
  AO21X1_HVT U293 ( .A1(n292), .A2(n147), .A3(n164), .Y(n291) );
  AO22X1_HVT U294 ( .A1(n293), .A2(n187), .A3(\mem[0][13] ), .A4(n877), .Y(
        n583) );
  AO21X1_HVT U295 ( .A1(n294), .A2(n149), .A3(n164), .Y(n293) );
  AO22X1_HVT U296 ( .A1(n295), .A2(n187), .A3(\mem[0][14] ), .A4(n876), .Y(
        n584) );
  AO21X1_HVT U297 ( .A1(n296), .A2(n148), .A3(n164), .Y(n295) );
  AO22X1_HVT U298 ( .A1(n297), .A2(n187), .A3(\mem[0][15] ), .A4(n875), .Y(
        n585) );
  AO21X1_HVT U299 ( .A1(n298), .A2(n147), .A3(n164), .Y(n297) );
  AND3X1_HVT U300 ( .A1(n299), .A2(n160), .A3(n300), .Y(n268) );
  AO22X1_HVT U301 ( .A1(n301), .A2(n187), .A3(\mem[1][0] ), .A4(n874), .Y(n586) );
  AO21X1_HVT U302 ( .A1(n146), .A2(n267), .A3(n164), .Y(n301) );
  AO22X1_HVT U303 ( .A1(n303), .A2(n187), .A3(\mem[1][1] ), .A4(n873), .Y(n587) );
  AO21X1_HVT U304 ( .A1(n146), .A2(n270), .A3(n164), .Y(n303) );
  AO22X1_HVT U305 ( .A1(n304), .A2(n187), .A3(\mem[1][2] ), .A4(n872), .Y(n588) );
  AO21X1_HVT U306 ( .A1(n146), .A2(n272), .A3(n164), .Y(n304) );
  AO22X1_HVT U307 ( .A1(n305), .A2(n187), .A3(\mem[1][3] ), .A4(n871), .Y(n589) );
  AO21X1_HVT U308 ( .A1(n146), .A2(n274), .A3(n164), .Y(n305) );
  AO22X1_HVT U309 ( .A1(n306), .A2(n187), .A3(\mem[1][4] ), .A4(n870), .Y(n590) );
  AO21X1_HVT U310 ( .A1(n146), .A2(n276), .A3(n164), .Y(n306) );
  AO22X1_HVT U311 ( .A1(n307), .A2(n187), .A3(\mem[1][5] ), .A4(n869), .Y(n591) );
  AO21X1_HVT U312 ( .A1(n146), .A2(n278), .A3(n164), .Y(n307) );
  AO22X1_HVT U313 ( .A1(n308), .A2(n187), .A3(\mem[1][6] ), .A4(n868), .Y(n592) );
  AO21X1_HVT U314 ( .A1(n146), .A2(n280), .A3(n164), .Y(n308) );
  AO22X1_HVT U315 ( .A1(n309), .A2(n187), .A3(\mem[1][7] ), .A4(n867), .Y(n593) );
  AO21X1_HVT U316 ( .A1(n146), .A2(n282), .A3(n164), .Y(n309) );
  AO22X1_HVT U317 ( .A1(n310), .A2(n188), .A3(\mem[1][8] ), .A4(n866), .Y(n594) );
  AO21X1_HVT U318 ( .A1(n145), .A2(n284), .A3(n165), .Y(n310) );
  AO22X1_HVT U319 ( .A1(n311), .A2(n188), .A3(\mem[1][9] ), .A4(n865), .Y(n595) );
  AO21X1_HVT U320 ( .A1(n145), .A2(n286), .A3(n165), .Y(n311) );
  AO22X1_HVT U321 ( .A1(n312), .A2(n188), .A3(\mem[1][10] ), .A4(n864), .Y(
        n596) );
  AO21X1_HVT U322 ( .A1(n145), .A2(n288), .A3(n165), .Y(n312) );
  AO22X1_HVT U323 ( .A1(n313), .A2(n188), .A3(\mem[1][11] ), .A4(n863), .Y(
        n597) );
  AO21X1_HVT U324 ( .A1(n145), .A2(n290), .A3(n165), .Y(n313) );
  AO22X1_HVT U325 ( .A1(n314), .A2(n188), .A3(\mem[1][12] ), .A4(n862), .Y(
        n598) );
  AO21X1_HVT U326 ( .A1(n145), .A2(n292), .A3(n165), .Y(n314) );
  AO22X1_HVT U327 ( .A1(n315), .A2(n188), .A3(\mem[1][13] ), .A4(n861), .Y(
        n599) );
  AO21X1_HVT U328 ( .A1(n145), .A2(n294), .A3(n165), .Y(n315) );
  AO22X1_HVT U329 ( .A1(n316), .A2(n188), .A3(\mem[1][14] ), .A4(n860), .Y(
        n600) );
  AO21X1_HVT U330 ( .A1(n145), .A2(n296), .A3(n165), .Y(n316) );
  AO22X1_HVT U331 ( .A1(n317), .A2(n188), .A3(\mem[1][15] ), .A4(n859), .Y(
        n601) );
  AO21X1_HVT U332 ( .A1(n145), .A2(n298), .A3(n165), .Y(n317) );
  AO22X1_HVT U334 ( .A1(n319), .A2(n188), .A3(\mem[2][0] ), .A4(n858), .Y(n602) );
  AO21X1_HVT U335 ( .A1(n144), .A2(n267), .A3(n165), .Y(n319) );
  AO22X1_HVT U336 ( .A1(n321), .A2(n188), .A3(\mem[2][1] ), .A4(n857), .Y(n603) );
  AO21X1_HVT U337 ( .A1(n144), .A2(n270), .A3(n165), .Y(n321) );
  AO22X1_HVT U338 ( .A1(n322), .A2(n188), .A3(\mem[2][2] ), .A4(n856), .Y(n604) );
  AO21X1_HVT U339 ( .A1(n144), .A2(n272), .A3(n165), .Y(n322) );
  AO22X1_HVT U340 ( .A1(n323), .A2(n188), .A3(\mem[2][3] ), .A4(n855), .Y(n605) );
  AO21X1_HVT U341 ( .A1(n144), .A2(n274), .A3(n165), .Y(n323) );
  AO22X1_HVT U342 ( .A1(n324), .A2(n189), .A3(\mem[2][4] ), .A4(n854), .Y(n606) );
  AO21X1_HVT U343 ( .A1(n144), .A2(n276), .A3(n165), .Y(n324) );
  AO22X1_HVT U344 ( .A1(n325), .A2(n189), .A3(\mem[2][5] ), .A4(n853), .Y(n607) );
  AO21X1_HVT U345 ( .A1(n144), .A2(n278), .A3(n165), .Y(n325) );
  AO22X1_HVT U346 ( .A1(n326), .A2(n189), .A3(\mem[2][6] ), .A4(n852), .Y(n608) );
  AO21X1_HVT U347 ( .A1(n144), .A2(n280), .A3(n165), .Y(n326) );
  AO22X1_HVT U348 ( .A1(n327), .A2(n189), .A3(\mem[2][7] ), .A4(n851), .Y(n609) );
  AO21X1_HVT U349 ( .A1(n144), .A2(n282), .A3(n166), .Y(n327) );
  AO22X1_HVT U350 ( .A1(n328), .A2(n189), .A3(\mem[2][8] ), .A4(n850), .Y(n610) );
  AO21X1_HVT U351 ( .A1(n143), .A2(n284), .A3(n166), .Y(n328) );
  AO22X1_HVT U352 ( .A1(n329), .A2(n189), .A3(\mem[2][9] ), .A4(n849), .Y(n611) );
  AO21X1_HVT U353 ( .A1(n143), .A2(n286), .A3(n166), .Y(n329) );
  AO22X1_HVT U354 ( .A1(n330), .A2(n189), .A3(\mem[2][10] ), .A4(n848), .Y(
        n612) );
  AO21X1_HVT U355 ( .A1(n143), .A2(n288), .A3(n166), .Y(n330) );
  AO22X1_HVT U356 ( .A1(n331), .A2(n189), .A3(\mem[2][11] ), .A4(n847), .Y(
        n613) );
  AO21X1_HVT U357 ( .A1(n143), .A2(n290), .A3(n166), .Y(n331) );
  AO22X1_HVT U358 ( .A1(n332), .A2(n189), .A3(\mem[2][12] ), .A4(n846), .Y(
        n614) );
  AO21X1_HVT U359 ( .A1(n143), .A2(n292), .A3(n166), .Y(n332) );
  AO22X1_HVT U360 ( .A1(n333), .A2(n189), .A3(\mem[2][13] ), .A4(n845), .Y(
        n615) );
  AO21X1_HVT U361 ( .A1(n143), .A2(n294), .A3(n166), .Y(n333) );
  AO22X1_HVT U362 ( .A1(n334), .A2(n189), .A3(\mem[2][14] ), .A4(n844), .Y(
        n616) );
  AO21X1_HVT U363 ( .A1(n143), .A2(n296), .A3(n166), .Y(n334) );
  AO22X1_HVT U364 ( .A1(n335), .A2(n189), .A3(\mem[2][15] ), .A4(n843), .Y(
        n617) );
  AO21X1_HVT U365 ( .A1(n143), .A2(n298), .A3(n166), .Y(n335) );
  AO22X1_HVT U367 ( .A1(n337), .A2(n185), .A3(\mem[3][0] ), .A4(n842), .Y(n618) );
  AO21X1_HVT U368 ( .A1(n142), .A2(n267), .A3(n166), .Y(n337) );
  AO22X1_HVT U369 ( .A1(n339), .A2(n205), .A3(\mem[3][1] ), .A4(n841), .Y(n619) );
  AO21X1_HVT U370 ( .A1(n142), .A2(n270), .A3(n166), .Y(n339) );
  AO22X1_HVT U371 ( .A1(n340), .A2(n181), .A3(\mem[3][2] ), .A4(n840), .Y(n620) );
  AO21X1_HVT U372 ( .A1(n142), .A2(n272), .A3(n166), .Y(n340) );
  AO22X1_HVT U373 ( .A1(n341), .A2(n182), .A3(\mem[3][3] ), .A4(n839), .Y(n621) );
  AO21X1_HVT U374 ( .A1(n142), .A2(n274), .A3(n166), .Y(n341) );
  AO22X1_HVT U375 ( .A1(n342), .A2(n183), .A3(\mem[3][4] ), .A4(n838), .Y(n622) );
  AO21X1_HVT U376 ( .A1(n142), .A2(n276), .A3(n166), .Y(n342) );
  AO22X1_HVT U377 ( .A1(n343), .A2(n185), .A3(\mem[3][5] ), .A4(n837), .Y(n623) );
  AO21X1_HVT U378 ( .A1(n142), .A2(n278), .A3(n166), .Y(n343) );
  AO22X1_HVT U379 ( .A1(n344), .A2(n205), .A3(\mem[3][6] ), .A4(n836), .Y(n624) );
  AO21X1_HVT U380 ( .A1(n142), .A2(n280), .A3(n167), .Y(n344) );
  AO22X1_HVT U381 ( .A1(n345), .A2(n185), .A3(\mem[3][7] ), .A4(n835), .Y(n625) );
  AO21X1_HVT U382 ( .A1(n142), .A2(n282), .A3(n167), .Y(n345) );
  AO22X1_HVT U383 ( .A1(n346), .A2(n205), .A3(\mem[3][8] ), .A4(n834), .Y(n626) );
  AO21X1_HVT U384 ( .A1(n141), .A2(n284), .A3(n167), .Y(n346) );
  AO22X1_HVT U385 ( .A1(n347), .A2(n185), .A3(\mem[3][9] ), .A4(n833), .Y(n627) );
  AO21X1_HVT U386 ( .A1(n141), .A2(n286), .A3(n167), .Y(n347) );
  AO22X1_HVT U387 ( .A1(n348), .A2(n205), .A3(\mem[3][10] ), .A4(n832), .Y(
        n628) );
  AO21X1_HVT U388 ( .A1(n141), .A2(n288), .A3(n167), .Y(n348) );
  AO22X1_HVT U389 ( .A1(n349), .A2(n205), .A3(\mem[3][11] ), .A4(n831), .Y(
        n629) );
  AO21X1_HVT U390 ( .A1(n141), .A2(n290), .A3(n167), .Y(n349) );
  AO22X1_HVT U391 ( .A1(n350), .A2(n190), .A3(\mem[3][12] ), .A4(n830), .Y(
        n630) );
  AO21X1_HVT U392 ( .A1(n141), .A2(n292), .A3(n167), .Y(n350) );
  AO22X1_HVT U393 ( .A1(n351), .A2(n190), .A3(\mem[3][13] ), .A4(n829), .Y(
        n631) );
  AO21X1_HVT U394 ( .A1(n141), .A2(n294), .A3(n167), .Y(n351) );
  AO22X1_HVT U395 ( .A1(n352), .A2(n190), .A3(\mem[3][14] ), .A4(n828), .Y(
        n632) );
  AO21X1_HVT U396 ( .A1(n141), .A2(n296), .A3(n167), .Y(n352) );
  AO22X1_HVT U397 ( .A1(n353), .A2(n190), .A3(\mem[3][15] ), .A4(n827), .Y(
        n633) );
  AO21X1_HVT U398 ( .A1(n141), .A2(n298), .A3(n167), .Y(n353) );
  AND2X1_HVT U400 ( .A1(n1020), .A2(n891), .Y(n300) );
  AO22X1_HVT U401 ( .A1(n355), .A2(n190), .A3(\mem[4][0] ), .A4(n826), .Y(n634) );
  AO21X1_HVT U402 ( .A1(n138), .A2(n267), .A3(n167), .Y(n355) );
  AO22X1_HVT U403 ( .A1(n357), .A2(n190), .A3(\mem[4][1] ), .A4(n338), .Y(n635) );
  AO21X1_HVT U404 ( .A1(n140), .A2(n270), .A3(n167), .Y(n357) );
  AO22X1_HVT U405 ( .A1(n358), .A2(n190), .A3(\mem[4][2] ), .A4(n320), .Y(n636) );
  AO21X1_HVT U406 ( .A1(n139), .A2(n272), .A3(n167), .Y(n358) );
  AO22X1_HVT U407 ( .A1(n359), .A2(n190), .A3(\mem[4][3] ), .A4(n302), .Y(n637) );
  AO21X1_HVT U408 ( .A1(n138), .A2(n274), .A3(n167), .Y(n359) );
  AO22X1_HVT U409 ( .A1(n360), .A2(n190), .A3(\mem[4][4] ), .A4(n265), .Y(n638) );
  AO21X1_HVT U410 ( .A1(n140), .A2(n276), .A3(n167), .Y(n360) );
  AO22X1_HVT U411 ( .A1(n361), .A2(n190), .A3(\mem[4][5] ), .A4(n264), .Y(n639) );
  AO21X1_HVT U412 ( .A1(n139), .A2(n278), .A3(n168), .Y(n361) );
  AO22X1_HVT U413 ( .A1(n362), .A2(n190), .A3(\mem[4][6] ), .A4(n263), .Y(n640) );
  AO21X1_HVT U414 ( .A1(n138), .A2(n280), .A3(n168), .Y(n362) );
  AO22X1_HVT U415 ( .A1(n363), .A2(n190), .A3(\mem[4][7] ), .A4(n262), .Y(n641) );
  AO21X1_HVT U416 ( .A1(n140), .A2(n282), .A3(n168), .Y(n363) );
  AO22X1_HVT U417 ( .A1(n364), .A2(n191), .A3(\mem[4][8] ), .A4(n261), .Y(n642) );
  AO21X1_HVT U418 ( .A1(n139), .A2(n284), .A3(n168), .Y(n364) );
  AO22X1_HVT U419 ( .A1(n365), .A2(n191), .A3(\mem[4][9] ), .A4(n260), .Y(n643) );
  AO21X1_HVT U420 ( .A1(n138), .A2(n286), .A3(n168), .Y(n365) );
  AO22X1_HVT U421 ( .A1(n366), .A2(n191), .A3(\mem[4][10] ), .A4(n259), .Y(
        n644) );
  AO21X1_HVT U422 ( .A1(n140), .A2(n288), .A3(n168), .Y(n366) );
  AO22X1_HVT U423 ( .A1(n367), .A2(n191), .A3(\mem[4][11] ), .A4(n258), .Y(
        n645) );
  AO21X1_HVT U424 ( .A1(n139), .A2(n290), .A3(n168), .Y(n367) );
  AO22X1_HVT U425 ( .A1(n368), .A2(n191), .A3(\mem[4][12] ), .A4(n257), .Y(
        n646) );
  AO21X1_HVT U426 ( .A1(n138), .A2(n292), .A3(n168), .Y(n368) );
  AO22X1_HVT U427 ( .A1(n369), .A2(n191), .A3(\mem[4][13] ), .A4(n256), .Y(
        n647) );
  AO21X1_HVT U428 ( .A1(n140), .A2(n294), .A3(n168), .Y(n369) );
  AO22X1_HVT U429 ( .A1(n370), .A2(n191), .A3(\mem[4][14] ), .A4(n255), .Y(
        n648) );
  AO21X1_HVT U430 ( .A1(n139), .A2(n296), .A3(n168), .Y(n370) );
  AO22X1_HVT U431 ( .A1(n371), .A2(n191), .A3(\mem[4][15] ), .A4(n254), .Y(
        n649) );
  AO21X1_HVT U432 ( .A1(n138), .A2(n298), .A3(n168), .Y(n371) );
  AND3X1_HVT U433 ( .A1(n299), .A2(n159), .A3(n372), .Y(n356) );
  AO22X1_HVT U434 ( .A1(n373), .A2(n191), .A3(\mem[5][0] ), .A4(n253), .Y(n650) );
  AO21X1_HVT U435 ( .A1(n135), .A2(n267), .A3(n168), .Y(n373) );
  AO22X1_HVT U436 ( .A1(n375), .A2(n191), .A3(\mem[5][1] ), .A4(n252), .Y(n651) );
  AO21X1_HVT U437 ( .A1(n137), .A2(n270), .A3(n168), .Y(n375) );
  AO22X1_HVT U438 ( .A1(n376), .A2(n191), .A3(\mem[5][2] ), .A4(n251), .Y(n652) );
  AO21X1_HVT U439 ( .A1(n136), .A2(n272), .A3(n168), .Y(n376) );
  AO22X1_HVT U440 ( .A1(n377), .A2(n191), .A3(\mem[5][3] ), .A4(n250), .Y(n653) );
  AO21X1_HVT U441 ( .A1(n135), .A2(n274), .A3(n168), .Y(n377) );
  AO22X1_HVT U442 ( .A1(n378), .A2(n192), .A3(\mem[5][4] ), .A4(n249), .Y(n654) );
  AO21X1_HVT U443 ( .A1(n137), .A2(n276), .A3(n169), .Y(n378) );
  AO22X1_HVT U444 ( .A1(n379), .A2(n192), .A3(\mem[5][5] ), .A4(n248), .Y(n655) );
  AO21X1_HVT U445 ( .A1(n136), .A2(n278), .A3(n169), .Y(n379) );
  AO22X1_HVT U446 ( .A1(n380), .A2(n192), .A3(\mem[5][6] ), .A4(n247), .Y(n656) );
  AO21X1_HVT U447 ( .A1(n135), .A2(n280), .A3(n169), .Y(n380) );
  AO22X1_HVT U448 ( .A1(n381), .A2(n192), .A3(\mem[5][7] ), .A4(n246), .Y(n657) );
  AO21X1_HVT U449 ( .A1(n137), .A2(n282), .A3(n169), .Y(n381) );
  AO22X1_HVT U450 ( .A1(n382), .A2(n192), .A3(\mem[5][8] ), .A4(n245), .Y(n658) );
  AO21X1_HVT U451 ( .A1(n136), .A2(n284), .A3(n169), .Y(n382) );
  AO22X1_HVT U452 ( .A1(n383), .A2(n192), .A3(\mem[5][9] ), .A4(n244), .Y(n659) );
  AO21X1_HVT U453 ( .A1(n135), .A2(n286), .A3(n169), .Y(n383) );
  AO22X1_HVT U454 ( .A1(n384), .A2(n192), .A3(\mem[5][10] ), .A4(n243), .Y(
        n660) );
  AO21X1_HVT U455 ( .A1(n137), .A2(n288), .A3(n169), .Y(n384) );
  AO22X1_HVT U456 ( .A1(n385), .A2(n192), .A3(\mem[5][11] ), .A4(n242), .Y(
        n661) );
  AO21X1_HVT U457 ( .A1(n136), .A2(n290), .A3(n169), .Y(n385) );
  AO22X1_HVT U458 ( .A1(n386), .A2(n192), .A3(\mem[5][12] ), .A4(n241), .Y(
        n662) );
  AO21X1_HVT U459 ( .A1(n135), .A2(n292), .A3(n169), .Y(n386) );
  AO22X1_HVT U460 ( .A1(n387), .A2(n192), .A3(\mem[5][13] ), .A4(n240), .Y(
        n663) );
  AO21X1_HVT U461 ( .A1(n137), .A2(n294), .A3(n169), .Y(n387) );
  AO22X1_HVT U462 ( .A1(n388), .A2(n192), .A3(\mem[5][14] ), .A4(n239), .Y(
        n664) );
  AO21X1_HVT U463 ( .A1(n136), .A2(n296), .A3(n169), .Y(n388) );
  AO22X1_HVT U464 ( .A1(n389), .A2(n192), .A3(\mem[5][15] ), .A4(n238), .Y(
        n665) );
  AO21X1_HVT U465 ( .A1(n135), .A2(n298), .A3(n169), .Y(n389) );
  AND3X1_HVT U466 ( .A1(n318), .A2(n159), .A3(n372), .Y(n374) );
  AO22X1_HVT U467 ( .A1(n390), .A2(n205), .A3(\mem[6][0] ), .A4(n237), .Y(n666) );
  AO21X1_HVT U468 ( .A1(n132), .A2(n267), .A3(n169), .Y(n390) );
  AO22X1_HVT U469 ( .A1(n392), .A2(n181), .A3(\mem[6][1] ), .A4(n236), .Y(n667) );
  AO21X1_HVT U470 ( .A1(n134), .A2(n270), .A3(n169), .Y(n392) );
  AO22X1_HVT U471 ( .A1(n393), .A2(n182), .A3(\mem[6][2] ), .A4(n235), .Y(n668) );
  AO21X1_HVT U472 ( .A1(n133), .A2(n272), .A3(n169), .Y(n393) );
  AO22X1_HVT U473 ( .A1(n394), .A2(n183), .A3(\mem[6][3] ), .A4(n234), .Y(n669) );
  AO21X1_HVT U474 ( .A1(n132), .A2(n274), .A3(n170), .Y(n394) );
  AO22X1_HVT U475 ( .A1(n395), .A2(n185), .A3(\mem[6][4] ), .A4(n233), .Y(n670) );
  AO21X1_HVT U476 ( .A1(n134), .A2(n276), .A3(n170), .Y(n395) );
  AO22X1_HVT U477 ( .A1(n396), .A2(n205), .A3(\mem[6][5] ), .A4(n232), .Y(n671) );
  AO21X1_HVT U478 ( .A1(n133), .A2(n278), .A3(n170), .Y(n396) );
  AO22X1_HVT U479 ( .A1(n397), .A2(n181), .A3(\mem[6][6] ), .A4(n231), .Y(n672) );
  AO21X1_HVT U480 ( .A1(n132), .A2(n280), .A3(n170), .Y(n397) );
  AO22X1_HVT U481 ( .A1(n398), .A2(n182), .A3(\mem[6][7] ), .A4(n230), .Y(n673) );
  AO21X1_HVT U482 ( .A1(n134), .A2(n282), .A3(n170), .Y(n398) );
  AO22X1_HVT U483 ( .A1(n399), .A2(n183), .A3(\mem[6][8] ), .A4(n229), .Y(n674) );
  AO21X1_HVT U484 ( .A1(n133), .A2(n284), .A3(n170), .Y(n399) );
  AO22X1_HVT U485 ( .A1(n400), .A2(n185), .A3(\mem[6][9] ), .A4(n228), .Y(n675) );
  AO21X1_HVT U486 ( .A1(n132), .A2(n286), .A3(n170), .Y(n400) );
  AO22X1_HVT U487 ( .A1(n401), .A2(n185), .A3(\mem[6][10] ), .A4(n227), .Y(
        n676) );
  AO21X1_HVT U488 ( .A1(n134), .A2(n288), .A3(n170), .Y(n401) );
  AO22X1_HVT U489 ( .A1(n402), .A2(n185), .A3(\mem[6][11] ), .A4(n226), .Y(
        n677) );
  AO21X1_HVT U490 ( .A1(n133), .A2(n290), .A3(n170), .Y(n402) );
  AO22X1_HVT U491 ( .A1(n403), .A2(n193), .A3(\mem[6][12] ), .A4(n225), .Y(
        n678) );
  AO21X1_HVT U492 ( .A1(n132), .A2(n292), .A3(n170), .Y(n403) );
  AO22X1_HVT U493 ( .A1(n404), .A2(n193), .A3(\mem[6][13] ), .A4(n224), .Y(
        n679) );
  AO21X1_HVT U494 ( .A1(n134), .A2(n294), .A3(n170), .Y(n404) );
  AO22X1_HVT U495 ( .A1(n405), .A2(n193), .A3(\mem[6][14] ), .A4(n223), .Y(
        n680) );
  AO21X1_HVT U496 ( .A1(n133), .A2(n296), .A3(n170), .Y(n405) );
  AO22X1_HVT U497 ( .A1(n406), .A2(n193), .A3(\mem[6][15] ), .A4(n222), .Y(
        n681) );
  AO21X1_HVT U498 ( .A1(n132), .A2(n298), .A3(n170), .Y(n406) );
  AND3X1_HVT U499 ( .A1(n336), .A2(n159), .A3(n372), .Y(n391) );
  AO22X1_HVT U500 ( .A1(n407), .A2(n193), .A3(\mem[7][0] ), .A4(n221), .Y(n682) );
  AO21X1_HVT U501 ( .A1(n129), .A2(n267), .A3(n170), .Y(n407) );
  AO22X1_HVT U502 ( .A1(n409), .A2(n193), .A3(\mem[7][1] ), .A4(n220), .Y(n683) );
  AO21X1_HVT U503 ( .A1(n131), .A2(n270), .A3(n170), .Y(n409) );
  AO22X1_HVT U504 ( .A1(n410), .A2(n193), .A3(\mem[7][2] ), .A4(n219), .Y(n684) );
  AO21X1_HVT U505 ( .A1(n130), .A2(n272), .A3(n171), .Y(n410) );
  AO22X1_HVT U506 ( .A1(n411), .A2(n193), .A3(\mem[7][3] ), .A4(n218), .Y(n685) );
  AO21X1_HVT U507 ( .A1(n129), .A2(n274), .A3(n171), .Y(n411) );
  AO22X1_HVT U508 ( .A1(n412), .A2(n193), .A3(\mem[7][4] ), .A4(n217), .Y(n686) );
  AO21X1_HVT U509 ( .A1(n131), .A2(n276), .A3(n171), .Y(n412) );
  AO22X1_HVT U510 ( .A1(n413), .A2(n193), .A3(\mem[7][5] ), .A4(n216), .Y(n687) );
  AO21X1_HVT U511 ( .A1(n130), .A2(n278), .A3(n171), .Y(n413) );
  AO22X1_HVT U512 ( .A1(n414), .A2(n193), .A3(\mem[7][6] ), .A4(n215), .Y(n688) );
  AO21X1_HVT U513 ( .A1(n129), .A2(n280), .A3(n171), .Y(n414) );
  AO22X1_HVT U514 ( .A1(n415), .A2(n193), .A3(\mem[7][7] ), .A4(n214), .Y(n689) );
  AO21X1_HVT U515 ( .A1(n131), .A2(n282), .A3(n171), .Y(n415) );
  AO22X1_HVT U516 ( .A1(n416), .A2(n194), .A3(\mem[7][8] ), .A4(n213), .Y(n690) );
  AO21X1_HVT U517 ( .A1(n130), .A2(n284), .A3(n171), .Y(n416) );
  AO22X1_HVT U518 ( .A1(n417), .A2(n194), .A3(\mem[7][9] ), .A4(n212), .Y(n691) );
  AO21X1_HVT U519 ( .A1(n129), .A2(n286), .A3(n171), .Y(n417) );
  AO22X1_HVT U520 ( .A1(n418), .A2(n194), .A3(\mem[7][10] ), .A4(n211), .Y(
        n692) );
  AO21X1_HVT U521 ( .A1(n131), .A2(n288), .A3(n171), .Y(n418) );
  AO22X1_HVT U522 ( .A1(n419), .A2(n194), .A3(\mem[7][11] ), .A4(n210), .Y(
        n693) );
  AO21X1_HVT U523 ( .A1(n130), .A2(n290), .A3(n171), .Y(n419) );
  AO22X1_HVT U524 ( .A1(n420), .A2(n194), .A3(\mem[7][12] ), .A4(n209), .Y(
        n694) );
  AO21X1_HVT U525 ( .A1(n129), .A2(n292), .A3(n171), .Y(n420) );
  AO22X1_HVT U526 ( .A1(n421), .A2(n194), .A3(\mem[7][13] ), .A4(n208), .Y(
        n695) );
  AO21X1_HVT U527 ( .A1(n131), .A2(n294), .A3(n171), .Y(n421) );
  AO22X1_HVT U528 ( .A1(n422), .A2(n194), .A3(\mem[7][14] ), .A4(n207), .Y(
        n696) );
  AO21X1_HVT U529 ( .A1(n130), .A2(n296), .A3(n171), .Y(n422) );
  AO22X1_HVT U530 ( .A1(n423), .A2(n194), .A3(\mem[7][15] ), .A4(n206), .Y(
        n697) );
  AO21X1_HVT U531 ( .A1(n129), .A2(n298), .A3(n171), .Y(n423) );
  AND3X1_HVT U532 ( .A1(n354), .A2(n159), .A3(n372), .Y(n408) );
  AND2X1_HVT U533 ( .A1(a_din[2]), .A2(n891), .Y(n372) );
  AO22X1_HVT U534 ( .A1(n424), .A2(n194), .A3(\mem[8][0] ), .A4(n955), .Y(n698) );
  AO21X1_HVT U535 ( .A1(n126), .A2(n267), .A3(n171), .Y(n424) );
  AO22X1_HVT U536 ( .A1(n426), .A2(n194), .A3(\mem[8][1] ), .A4(n954), .Y(n699) );
  AO21X1_HVT U537 ( .A1(n128), .A2(n270), .A3(n172), .Y(n426) );
  AO22X1_HVT U538 ( .A1(n427), .A2(n194), .A3(\mem[8][2] ), .A4(n953), .Y(n700) );
  AO21X1_HVT U539 ( .A1(n127), .A2(n272), .A3(n172), .Y(n427) );
  AO22X1_HVT U540 ( .A1(n428), .A2(n194), .A3(\mem[8][3] ), .A4(n952), .Y(n701) );
  AO21X1_HVT U541 ( .A1(n126), .A2(n274), .A3(n172), .Y(n428) );
  AO22X1_HVT U542 ( .A1(n429), .A2(n195), .A3(\mem[8][4] ), .A4(n951), .Y(n702) );
  AO21X1_HVT U543 ( .A1(n128), .A2(n276), .A3(n172), .Y(n429) );
  AO22X1_HVT U544 ( .A1(n430), .A2(n195), .A3(\mem[8][5] ), .A4(n950), .Y(n703) );
  AO21X1_HVT U545 ( .A1(n127), .A2(n278), .A3(n172), .Y(n430) );
  AO22X1_HVT U546 ( .A1(n431), .A2(n195), .A3(\mem[8][6] ), .A4(n949), .Y(n704) );
  AO21X1_HVT U547 ( .A1(n126), .A2(n280), .A3(n172), .Y(n431) );
  AO22X1_HVT U548 ( .A1(n432), .A2(n195), .A3(\mem[8][7] ), .A4(n948), .Y(n705) );
  AO21X1_HVT U549 ( .A1(n128), .A2(n282), .A3(n172), .Y(n432) );
  AO22X1_HVT U550 ( .A1(n433), .A2(n195), .A3(\mem[8][8] ), .A4(n947), .Y(n706) );
  AO21X1_HVT U551 ( .A1(n127), .A2(n284), .A3(n172), .Y(n433) );
  AO22X1_HVT U552 ( .A1(n434), .A2(n195), .A3(\mem[8][9] ), .A4(n946), .Y(n707) );
  AO21X1_HVT U553 ( .A1(n126), .A2(n286), .A3(n172), .Y(n434) );
  AO22X1_HVT U554 ( .A1(n435), .A2(n195), .A3(\mem[8][10] ), .A4(n945), .Y(
        n708) );
  AO21X1_HVT U555 ( .A1(n128), .A2(n288), .A3(n172), .Y(n435) );
  AO22X1_HVT U556 ( .A1(n436), .A2(n195), .A3(\mem[8][11] ), .A4(n944), .Y(
        n709) );
  AO21X1_HVT U557 ( .A1(n127), .A2(n290), .A3(n172), .Y(n436) );
  AO22X1_HVT U558 ( .A1(n437), .A2(n195), .A3(\mem[8][12] ), .A4(n943), .Y(
        n710) );
  AO21X1_HVT U559 ( .A1(n126), .A2(n292), .A3(n172), .Y(n437) );
  AO22X1_HVT U560 ( .A1(n438), .A2(n195), .A3(\mem[8][13] ), .A4(n942), .Y(
        n711) );
  AO21X1_HVT U561 ( .A1(n128), .A2(n294), .A3(n172), .Y(n438) );
  AO22X1_HVT U562 ( .A1(n439), .A2(n195), .A3(\mem[8][14] ), .A4(n941), .Y(
        n712) );
  AO21X1_HVT U563 ( .A1(n127), .A2(n296), .A3(n172), .Y(n439) );
  AO22X1_HVT U564 ( .A1(n440), .A2(n195), .A3(\mem[8][15] ), .A4(n940), .Y(
        n713) );
  AO21X1_HVT U565 ( .A1(n126), .A2(n298), .A3(n172), .Y(n440) );
  AND3X1_HVT U566 ( .A1(n299), .A2(n4), .A3(n441), .Y(n425) );
  AO22X1_HVT U567 ( .A1(n442), .A2(n196), .A3(\mem[9][0] ), .A4(n939), .Y(n714) );
  AO21X1_HVT U568 ( .A1(n123), .A2(n267), .A3(n173), .Y(n442) );
  AO22X1_HVT U569 ( .A1(n444), .A2(n196), .A3(\mem[9][1] ), .A4(n938), .Y(n715) );
  AO21X1_HVT U570 ( .A1(n125), .A2(n270), .A3(n173), .Y(n444) );
  AO22X1_HVT U571 ( .A1(n445), .A2(n196), .A3(\mem[9][2] ), .A4(n937), .Y(n716) );
  AO21X1_HVT U572 ( .A1(n124), .A2(n272), .A3(n173), .Y(n445) );
  AO22X1_HVT U573 ( .A1(n446), .A2(n196), .A3(\mem[9][3] ), .A4(n936), .Y(n717) );
  AO21X1_HVT U574 ( .A1(n123), .A2(n274), .A3(n173), .Y(n446) );
  AO22X1_HVT U575 ( .A1(n447), .A2(n196), .A3(\mem[9][4] ), .A4(n935), .Y(n718) );
  AO21X1_HVT U576 ( .A1(n125), .A2(n276), .A3(n173), .Y(n447) );
  AO22X1_HVT U577 ( .A1(n448), .A2(n196), .A3(\mem[9][5] ), .A4(n934), .Y(n719) );
  AO21X1_HVT U578 ( .A1(n124), .A2(n278), .A3(n173), .Y(n448) );
  AO22X1_HVT U579 ( .A1(n449), .A2(n196), .A3(\mem[9][6] ), .A4(n933), .Y(n720) );
  AO21X1_HVT U580 ( .A1(n123), .A2(n280), .A3(n173), .Y(n449) );
  AO22X1_HVT U581 ( .A1(n450), .A2(n196), .A3(\mem[9][7] ), .A4(n932), .Y(n721) );
  AO21X1_HVT U582 ( .A1(n125), .A2(n282), .A3(n173), .Y(n450) );
  AO22X1_HVT U583 ( .A1(n451), .A2(n196), .A3(\mem[9][8] ), .A4(n931), .Y(n722) );
  AO21X1_HVT U584 ( .A1(n124), .A2(n284), .A3(n173), .Y(n451) );
  AO22X1_HVT U585 ( .A1(n452), .A2(n196), .A3(\mem[9][9] ), .A4(n930), .Y(n723) );
  AO21X1_HVT U586 ( .A1(n123), .A2(n286), .A3(n173), .Y(n452) );
  AO22X1_HVT U587 ( .A1(n453), .A2(n196), .A3(\mem[9][10] ), .A4(n929), .Y(
        n724) );
  AO21X1_HVT U588 ( .A1(n125), .A2(n288), .A3(n173), .Y(n453) );
  AO22X1_HVT U589 ( .A1(n454), .A2(n196), .A3(\mem[9][11] ), .A4(n928), .Y(
        n725) );
  AO21X1_HVT U590 ( .A1(n124), .A2(n290), .A3(n173), .Y(n454) );
  AO22X1_HVT U591 ( .A1(n455), .A2(n197), .A3(\mem[9][12] ), .A4(n927), .Y(
        n726) );
  AO21X1_HVT U592 ( .A1(n123), .A2(n292), .A3(n173), .Y(n455) );
  AO22X1_HVT U593 ( .A1(n456), .A2(n197), .A3(\mem[9][13] ), .A4(n926), .Y(
        n727) );
  AO21X1_HVT U594 ( .A1(n125), .A2(n294), .A3(n173), .Y(n456) );
  AO22X1_HVT U595 ( .A1(n457), .A2(n197), .A3(\mem[9][14] ), .A4(n925), .Y(
        n728) );
  AO21X1_HVT U596 ( .A1(n124), .A2(n296), .A3(n173), .Y(n457) );
  AO22X1_HVT U597 ( .A1(n458), .A2(n197), .A3(\mem[9][15] ), .A4(n924), .Y(
        n729) );
  AO21X1_HVT U598 ( .A1(n123), .A2(n298), .A3(n174), .Y(n458) );
  AND3X1_HVT U599 ( .A1(n318), .A2(n3), .A3(n441), .Y(n443) );
  AO22X1_HVT U600 ( .A1(n459), .A2(n197), .A3(\mem[10][0] ), .A4(n923), .Y(
        n730) );
  AO21X1_HVT U601 ( .A1(n120), .A2(n267), .A3(n174), .Y(n459) );
  AO22X1_HVT U602 ( .A1(n461), .A2(n197), .A3(\mem[10][1] ), .A4(n922), .Y(
        n731) );
  AO21X1_HVT U603 ( .A1(n122), .A2(n270), .A3(n174), .Y(n461) );
  AO22X1_HVT U604 ( .A1(n462), .A2(n197), .A3(\mem[10][2] ), .A4(n921), .Y(
        n732) );
  AO21X1_HVT U605 ( .A1(n121), .A2(n272), .A3(n174), .Y(n462) );
  AO22X1_HVT U606 ( .A1(n463), .A2(n197), .A3(\mem[10][3] ), .A4(n920), .Y(
        n733) );
  AO21X1_HVT U607 ( .A1(n120), .A2(n274), .A3(n174), .Y(n463) );
  AO22X1_HVT U608 ( .A1(n464), .A2(n197), .A3(\mem[10][4] ), .A4(n919), .Y(
        n734) );
  AO21X1_HVT U609 ( .A1(n122), .A2(n276), .A3(n174), .Y(n464) );
  AO22X1_HVT U610 ( .A1(n465), .A2(n197), .A3(\mem[10][5] ), .A4(n918), .Y(
        n735) );
  AO21X1_HVT U611 ( .A1(n121), .A2(n278), .A3(n174), .Y(n465) );
  AO22X1_HVT U612 ( .A1(n466), .A2(n197), .A3(\mem[10][6] ), .A4(n917), .Y(
        n736) );
  AO21X1_HVT U613 ( .A1(n120), .A2(n280), .A3(n174), .Y(n466) );
  AO22X1_HVT U614 ( .A1(n467), .A2(n197), .A3(\mem[10][7] ), .A4(n916), .Y(
        n737) );
  AO21X1_HVT U615 ( .A1(n122), .A2(n282), .A3(n174), .Y(n467) );
  AO22X1_HVT U616 ( .A1(n468), .A2(n198), .A3(\mem[10][8] ), .A4(n915), .Y(
        n738) );
  AO21X1_HVT U617 ( .A1(n121), .A2(n284), .A3(n174), .Y(n468) );
  AO22X1_HVT U618 ( .A1(n469), .A2(n198), .A3(\mem[10][9] ), .A4(n914), .Y(
        n739) );
  AO21X1_HVT U619 ( .A1(n120), .A2(n286), .A3(n174), .Y(n469) );
  AO22X1_HVT U620 ( .A1(n470), .A2(n198), .A3(\mem[10][10] ), .A4(n913), .Y(
        n740) );
  AO21X1_HVT U621 ( .A1(n122), .A2(n288), .A3(n174), .Y(n470) );
  AO22X1_HVT U622 ( .A1(n471), .A2(n198), .A3(\mem[10][11] ), .A4(n912), .Y(
        n741) );
  AO21X1_HVT U623 ( .A1(n121), .A2(n290), .A3(n174), .Y(n471) );
  AO22X1_HVT U624 ( .A1(n472), .A2(n198), .A3(\mem[10][12] ), .A4(n911), .Y(
        n742) );
  AO21X1_HVT U625 ( .A1(n120), .A2(n292), .A3(n174), .Y(n472) );
  AO22X1_HVT U626 ( .A1(n473), .A2(n198), .A3(\mem[10][13] ), .A4(n910), .Y(
        n743) );
  AO21X1_HVT U627 ( .A1(n122), .A2(n294), .A3(n174), .Y(n473) );
  AO22X1_HVT U628 ( .A1(n474), .A2(n198), .A3(\mem[10][14] ), .A4(n909), .Y(
        n744) );
  AO21X1_HVT U629 ( .A1(n121), .A2(n296), .A3(n175), .Y(n474) );
  AO22X1_HVT U630 ( .A1(n475), .A2(n198), .A3(\mem[10][15] ), .A4(n908), .Y(
        n745) );
  AO21X1_HVT U631 ( .A1(n120), .A2(n298), .A3(n175), .Y(n475) );
  AND3X1_HVT U632 ( .A1(n336), .A2(n160), .A3(n441), .Y(n460) );
  AO22X1_HVT U633 ( .A1(n476), .A2(n198), .A3(\mem[11][0] ), .A4(n907), .Y(
        n746) );
  AO21X1_HVT U634 ( .A1(n117), .A2(n267), .A3(n175), .Y(n476) );
  AO22X1_HVT U635 ( .A1(n478), .A2(n198), .A3(\mem[11][1] ), .A4(n906), .Y(
        n747) );
  AO21X1_HVT U636 ( .A1(n119), .A2(n270), .A3(n175), .Y(n478) );
  AO22X1_HVT U637 ( .A1(n479), .A2(n198), .A3(\mem[11][2] ), .A4(n905), .Y(
        n748) );
  AO21X1_HVT U638 ( .A1(n118), .A2(n272), .A3(n175), .Y(n479) );
  AO22X1_HVT U639 ( .A1(n480), .A2(n198), .A3(\mem[11][3] ), .A4(n904), .Y(
        n749) );
  AO21X1_HVT U640 ( .A1(n117), .A2(n274), .A3(n175), .Y(n480) );
  AO22X1_HVT U641 ( .A1(n481), .A2(n199), .A3(\mem[11][4] ), .A4(n903), .Y(
        n750) );
  AO21X1_HVT U642 ( .A1(n119), .A2(n276), .A3(n175), .Y(n481) );
  AO22X1_HVT U643 ( .A1(n482), .A2(n199), .A3(\mem[11][5] ), .A4(n902), .Y(
        n751) );
  AO21X1_HVT U644 ( .A1(n118), .A2(n278), .A3(n175), .Y(n482) );
  AO22X1_HVT U645 ( .A1(n483), .A2(n199), .A3(\mem[11][6] ), .A4(n901), .Y(
        n752) );
  AO21X1_HVT U646 ( .A1(n117), .A2(n280), .A3(n175), .Y(n483) );
  AO22X1_HVT U647 ( .A1(n484), .A2(n199), .A3(\mem[11][7] ), .A4(n900), .Y(
        n753) );
  AO21X1_HVT U648 ( .A1(n119), .A2(n282), .A3(n175), .Y(n484) );
  AO22X1_HVT U649 ( .A1(n485), .A2(n199), .A3(\mem[11][8] ), .A4(n899), .Y(
        n754) );
  AO21X1_HVT U650 ( .A1(n118), .A2(n284), .A3(n175), .Y(n485) );
  AO22X1_HVT U651 ( .A1(n486), .A2(n199), .A3(\mem[11][9] ), .A4(n898), .Y(
        n755) );
  AO21X1_HVT U652 ( .A1(n117), .A2(n286), .A3(n175), .Y(n486) );
  AO22X1_HVT U653 ( .A1(n487), .A2(n199), .A3(\mem[11][10] ), .A4(n897), .Y(
        n756) );
  AO21X1_HVT U654 ( .A1(n119), .A2(n288), .A3(n175), .Y(n487) );
  AO22X1_HVT U655 ( .A1(n488), .A2(n199), .A3(\mem[11][11] ), .A4(n896), .Y(
        n757) );
  AO21X1_HVT U656 ( .A1(n118), .A2(n290), .A3(n175), .Y(n488) );
  AO22X1_HVT U657 ( .A1(n489), .A2(n199), .A3(\mem[11][12] ), .A4(n895), .Y(
        n758) );
  AO21X1_HVT U658 ( .A1(n117), .A2(n292), .A3(n175), .Y(n489) );
  AO22X1_HVT U659 ( .A1(n490), .A2(n199), .A3(\mem[11][13] ), .A4(n894), .Y(
        n759) );
  AO21X1_HVT U660 ( .A1(n119), .A2(n294), .A3(n176), .Y(n490) );
  AO22X1_HVT U661 ( .A1(n491), .A2(n199), .A3(\mem[11][14] ), .A4(n893), .Y(
        n760) );
  AO21X1_HVT U662 ( .A1(n118), .A2(n296), .A3(n176), .Y(n491) );
  AO22X1_HVT U663 ( .A1(n492), .A2(n199), .A3(\mem[11][15] ), .A4(n892), .Y(
        n761) );
  AO21X1_HVT U664 ( .A1(n117), .A2(n298), .A3(n176), .Y(n492) );
  AND3X1_HVT U665 ( .A1(n354), .A2(n4), .A3(n441), .Y(n477) );
  AND2X1_HVT U666 ( .A1(a_din[3]), .A2(n1020), .Y(n441) );
  AO22X1_HVT U667 ( .A1(n493), .A2(n200), .A3(\mem[12][0] ), .A4(n1019), .Y(
        n762) );
  AO21X1_HVT U668 ( .A1(n114), .A2(n267), .A3(n176), .Y(n493) );
  AO22X1_HVT U669 ( .A1(n495), .A2(n200), .A3(\mem[12][1] ), .A4(n1018), .Y(
        n763) );
  AO21X1_HVT U670 ( .A1(n116), .A2(n270), .A3(n176), .Y(n495) );
  AO22X1_HVT U671 ( .A1(n496), .A2(n200), .A3(\mem[12][2] ), .A4(n1017), .Y(
        n764) );
  AO21X1_HVT U672 ( .A1(n115), .A2(n272), .A3(n176), .Y(n496) );
  AO22X1_HVT U673 ( .A1(n497), .A2(n200), .A3(\mem[12][3] ), .A4(n1016), .Y(
        n765) );
  AO21X1_HVT U674 ( .A1(n114), .A2(n274), .A3(n176), .Y(n497) );
  AO22X1_HVT U675 ( .A1(n498), .A2(n200), .A3(\mem[12][4] ), .A4(n1015), .Y(
        n766) );
  AO21X1_HVT U676 ( .A1(n116), .A2(n276), .A3(n176), .Y(n498) );
  AO22X1_HVT U677 ( .A1(n499), .A2(n200), .A3(\mem[12][5] ), .A4(n1014), .Y(
        n767) );
  AO21X1_HVT U678 ( .A1(n115), .A2(n278), .A3(n176), .Y(n499) );
  AO22X1_HVT U679 ( .A1(n500), .A2(n200), .A3(\mem[12][6] ), .A4(n1013), .Y(
        n768) );
  AO21X1_HVT U680 ( .A1(n114), .A2(n280), .A3(n176), .Y(n500) );
  AO22X1_HVT U681 ( .A1(n501), .A2(n200), .A3(\mem[12][7] ), .A4(n1012), .Y(
        n769) );
  AO21X1_HVT U682 ( .A1(n116), .A2(n282), .A3(n176), .Y(n501) );
  AO22X1_HVT U683 ( .A1(n502), .A2(n200), .A3(\mem[12][8] ), .A4(n1011), .Y(
        n770) );
  AO21X1_HVT U684 ( .A1(n115), .A2(n284), .A3(n176), .Y(n502) );
  AO22X1_HVT U685 ( .A1(n503), .A2(n200), .A3(\mem[12][9] ), .A4(n1010), .Y(
        n771) );
  AO21X1_HVT U686 ( .A1(n114), .A2(n286), .A3(n176), .Y(n503) );
  AO22X1_HVT U687 ( .A1(n504), .A2(n200), .A3(\mem[12][10] ), .A4(n1009), .Y(
        n772) );
  AO21X1_HVT U688 ( .A1(n116), .A2(n288), .A3(n176), .Y(n504) );
  AO22X1_HVT U689 ( .A1(n505), .A2(n200), .A3(\mem[12][11] ), .A4(n1008), .Y(
        n773) );
  AO21X1_HVT U690 ( .A1(n115), .A2(n290), .A3(n176), .Y(n505) );
  AO22X1_HVT U691 ( .A1(n506), .A2(n201), .A3(\mem[12][12] ), .A4(n1007), .Y(
        n774) );
  AO21X1_HVT U692 ( .A1(n114), .A2(n292), .A3(n177), .Y(n506) );
  AO22X1_HVT U693 ( .A1(n507), .A2(n201), .A3(\mem[12][13] ), .A4(n1006), .Y(
        n775) );
  AO21X1_HVT U694 ( .A1(n116), .A2(n294), .A3(n177), .Y(n507) );
  AO22X1_HVT U695 ( .A1(n508), .A2(n201), .A3(\mem[12][14] ), .A4(n1005), .Y(
        n776) );
  AO21X1_HVT U696 ( .A1(n115), .A2(n296), .A3(n177), .Y(n508) );
  AO22X1_HVT U697 ( .A1(n509), .A2(n201), .A3(\mem[12][15] ), .A4(n1004), .Y(
        n777) );
  AO21X1_HVT U698 ( .A1(n114), .A2(n298), .A3(n177), .Y(n509) );
  AND3X1_HVT U699 ( .A1(n299), .A2(n3), .A3(n510), .Y(n494) );
  AND2X1_HVT U700 ( .A1(n150), .A2(n152), .Y(n299) );
  AO22X1_HVT U701 ( .A1(n511), .A2(n201), .A3(\mem[13][0] ), .A4(n1003), .Y(
        n778) );
  AO21X1_HVT U702 ( .A1(n111), .A2(n267), .A3(n177), .Y(n511) );
  AO22X1_HVT U703 ( .A1(n513), .A2(n201), .A3(\mem[13][1] ), .A4(n1002), .Y(
        n779) );
  AO21X1_HVT U704 ( .A1(n113), .A2(n270), .A3(n177), .Y(n513) );
  AO22X1_HVT U705 ( .A1(n514), .A2(n201), .A3(\mem[13][2] ), .A4(n1001), .Y(
        n780) );
  AO21X1_HVT U706 ( .A1(n112), .A2(n272), .A3(n177), .Y(n514) );
  AO22X1_HVT U707 ( .A1(n515), .A2(n201), .A3(\mem[13][3] ), .A4(n1000), .Y(
        n781) );
  AO21X1_HVT U708 ( .A1(n111), .A2(n274), .A3(n177), .Y(n515) );
  AO22X1_HVT U709 ( .A1(n516), .A2(n201), .A3(\mem[13][4] ), .A4(n999), .Y(
        n782) );
  AO21X1_HVT U710 ( .A1(n113), .A2(n276), .A3(n177), .Y(n516) );
  AO22X1_HVT U711 ( .A1(n517), .A2(n201), .A3(\mem[13][5] ), .A4(n998), .Y(
        n783) );
  AO21X1_HVT U712 ( .A1(n112), .A2(n278), .A3(n177), .Y(n517) );
  AO22X1_HVT U713 ( .A1(n518), .A2(n201), .A3(\mem[13][6] ), .A4(n997), .Y(
        n784) );
  AO21X1_HVT U714 ( .A1(n111), .A2(n280), .A3(n177), .Y(n518) );
  AO22X1_HVT U715 ( .A1(n519), .A2(n201), .A3(\mem[13][7] ), .A4(n996), .Y(
        n785) );
  AO21X1_HVT U716 ( .A1(n113), .A2(n282), .A3(n177), .Y(n519) );
  AO22X1_HVT U717 ( .A1(n520), .A2(n202), .A3(\mem[13][8] ), .A4(n995), .Y(
        n786) );
  AO21X1_HVT U718 ( .A1(n112), .A2(n284), .A3(n177), .Y(n520) );
  AO22X1_HVT U719 ( .A1(n521), .A2(n202), .A3(\mem[13][9] ), .A4(n994), .Y(
        n787) );
  AO21X1_HVT U720 ( .A1(n111), .A2(n286), .A3(n177), .Y(n521) );
  AO22X1_HVT U721 ( .A1(n522), .A2(n202), .A3(\mem[13][10] ), .A4(n993), .Y(
        n788) );
  AO21X1_HVT U722 ( .A1(n113), .A2(n288), .A3(n177), .Y(n522) );
  AO22X1_HVT U723 ( .A1(n523), .A2(n202), .A3(\mem[13][11] ), .A4(n992), .Y(
        n789) );
  AO21X1_HVT U724 ( .A1(n112), .A2(n290), .A3(n178), .Y(n523) );
  AO22X1_HVT U725 ( .A1(n524), .A2(n202), .A3(\mem[13][12] ), .A4(n991), .Y(
        n790) );
  AO21X1_HVT U726 ( .A1(n111), .A2(n292), .A3(n178), .Y(n524) );
  AO22X1_HVT U727 ( .A1(n525), .A2(n202), .A3(\mem[13][13] ), .A4(n990), .Y(
        n791) );
  AO21X1_HVT U728 ( .A1(n113), .A2(n294), .A3(n178), .Y(n525) );
  AO22X1_HVT U729 ( .A1(n526), .A2(n202), .A3(\mem[13][14] ), .A4(n989), .Y(
        n792) );
  AO21X1_HVT U730 ( .A1(n112), .A2(n296), .A3(n178), .Y(n526) );
  AO22X1_HVT U731 ( .A1(n527), .A2(n202), .A3(\mem[13][15] ), .A4(n988), .Y(
        n793) );
  AO21X1_HVT U732 ( .A1(n111), .A2(n298), .A3(n178), .Y(n527) );
  AND3X1_HVT U733 ( .A1(n318), .A2(n160), .A3(n510), .Y(n512) );
  AND2X1_HVT U734 ( .A1(a_din[0]), .A2(n152), .Y(n318) );
  AO22X1_HVT U735 ( .A1(n528), .A2(n202), .A3(\mem[14][0] ), .A4(n987), .Y(
        n794) );
  AO21X1_HVT U736 ( .A1(n108), .A2(n267), .A3(n178), .Y(n528) );
  AO22X1_HVT U737 ( .A1(n530), .A2(n202), .A3(\mem[14][1] ), .A4(n986), .Y(
        n795) );
  AO21X1_HVT U738 ( .A1(n110), .A2(n270), .A3(n178), .Y(n530) );
  AO22X1_HVT U739 ( .A1(n531), .A2(n202), .A3(\mem[14][2] ), .A4(n985), .Y(
        n796) );
  AO21X1_HVT U740 ( .A1(n109), .A2(n272), .A3(n178), .Y(n531) );
  AO22X1_HVT U741 ( .A1(n532), .A2(n202), .A3(\mem[14][3] ), .A4(n984), .Y(
        n797) );
  AO21X1_HVT U742 ( .A1(n108), .A2(n274), .A3(n178), .Y(n532) );
  AO22X1_HVT U743 ( .A1(n533), .A2(n203), .A3(\mem[14][4] ), .A4(n983), .Y(
        n798) );
  AO21X1_HVT U744 ( .A1(n110), .A2(n276), .A3(n178), .Y(n533) );
  AO22X1_HVT U745 ( .A1(n534), .A2(n203), .A3(\mem[14][5] ), .A4(n982), .Y(
        n799) );
  AO21X1_HVT U746 ( .A1(n109), .A2(n278), .A3(n178), .Y(n534) );
  AO22X1_HVT U747 ( .A1(n535), .A2(n203), .A3(\mem[14][6] ), .A4(n981), .Y(
        n800) );
  AO21X1_HVT U748 ( .A1(n108), .A2(n280), .A3(n178), .Y(n535) );
  AO22X1_HVT U749 ( .A1(n536), .A2(n203), .A3(\mem[14][7] ), .A4(n980), .Y(
        n801) );
  AO21X1_HVT U750 ( .A1(n110), .A2(n282), .A3(n178), .Y(n536) );
  AO22X1_HVT U751 ( .A1(n537), .A2(n203), .A3(\mem[14][8] ), .A4(n979), .Y(
        n802) );
  AO21X1_HVT U752 ( .A1(n109), .A2(n284), .A3(n178), .Y(n537) );
  AO22X1_HVT U753 ( .A1(n538), .A2(n203), .A3(\mem[14][9] ), .A4(n978), .Y(
        n803) );
  AO21X1_HVT U754 ( .A1(n108), .A2(n286), .A3(n178), .Y(n538) );
  AO22X1_HVT U755 ( .A1(n539), .A2(n203), .A3(\mem[14][10] ), .A4(n977), .Y(
        n804) );
  AO21X1_HVT U756 ( .A1(n110), .A2(n288), .A3(n179), .Y(n539) );
  AO22X1_HVT U757 ( .A1(n540), .A2(n203), .A3(\mem[14][11] ), .A4(n976), .Y(
        n805) );
  AO21X1_HVT U758 ( .A1(n109), .A2(n290), .A3(n179), .Y(n540) );
  AO22X1_HVT U759 ( .A1(n541), .A2(n203), .A3(\mem[14][12] ), .A4(n975), .Y(
        n806) );
  AO21X1_HVT U760 ( .A1(n108), .A2(n292), .A3(n179), .Y(n541) );
  AO22X1_HVT U761 ( .A1(n542), .A2(n203), .A3(\mem[14][13] ), .A4(n974), .Y(
        n807) );
  AO21X1_HVT U762 ( .A1(n110), .A2(n294), .A3(n179), .Y(n542) );
  AO22X1_HVT U763 ( .A1(n543), .A2(n203), .A3(\mem[14][14] ), .A4(n973), .Y(
        n808) );
  AO21X1_HVT U764 ( .A1(n109), .A2(n296), .A3(n179), .Y(n543) );
  AO22X1_HVT U765 ( .A1(n544), .A2(n203), .A3(\mem[14][15] ), .A4(n972), .Y(
        n809) );
  AO21X1_HVT U766 ( .A1(n108), .A2(n298), .A3(n179), .Y(n544) );
  AND3X1_HVT U767 ( .A1(n336), .A2(n4), .A3(n510), .Y(n529) );
  AND2X1_HVT U768 ( .A1(n151), .A2(n150), .Y(n336) );
  AO22X1_HVT U769 ( .A1(n545), .A2(n204), .A3(\mem[15][0] ), .A4(n971), .Y(
        n810) );
  AO21X1_HVT U770 ( .A1(n105), .A2(n267), .A3(n179), .Y(n545) );
  AND2X1_HVT U771 ( .A1(n547), .A2(n548), .Y(n267) );
  AO22X1_HVT U772 ( .A1(n549), .A2(n204), .A3(\mem[15][1] ), .A4(n970), .Y(
        n811) );
  AO21X1_HVT U773 ( .A1(n107), .A2(n270), .A3(n179), .Y(n549) );
  AND2X1_HVT U774 ( .A1(n550), .A2(n547), .Y(n270) );
  AO22X1_HVT U775 ( .A1(n551), .A2(n204), .A3(\mem[15][2] ), .A4(n969), .Y(
        n812) );
  AO21X1_HVT U776 ( .A1(n106), .A2(n272), .A3(n179), .Y(n551) );
  AND2X1_HVT U777 ( .A1(n552), .A2(n547), .Y(n272) );
  AO22X1_HVT U778 ( .A1(n553), .A2(n204), .A3(\mem[15][3] ), .A4(n968), .Y(
        n813) );
  AO21X1_HVT U779 ( .A1(n105), .A2(n274), .A3(n179), .Y(n553) );
  AND2X1_HVT U780 ( .A1(n554), .A2(n547), .Y(n274) );
  AND2X1_HVT U781 ( .A1(n156), .A2(n158), .Y(n547) );
  AO22X1_HVT U782 ( .A1(n555), .A2(n204), .A3(\mem[15][4] ), .A4(n967), .Y(
        n814) );
  AO21X1_HVT U783 ( .A1(n107), .A2(n276), .A3(n179), .Y(n555) );
  AND2X1_HVT U784 ( .A1(n556), .A2(n548), .Y(n276) );
  AO22X1_HVT U785 ( .A1(n557), .A2(n204), .A3(\mem[15][5] ), .A4(n966), .Y(
        n815) );
  AO21X1_HVT U786 ( .A1(n106), .A2(n278), .A3(n179), .Y(n557) );
  AND2X1_HVT U787 ( .A1(n556), .A2(n550), .Y(n278) );
  AO22X1_HVT U788 ( .A1(n558), .A2(n204), .A3(\mem[15][6] ), .A4(n965), .Y(
        n816) );
  AO21X1_HVT U789 ( .A1(n105), .A2(n280), .A3(n179), .Y(n558) );
  AND2X1_HVT U790 ( .A1(n556), .A2(n552), .Y(n280) );
  AO22X1_HVT U791 ( .A1(n559), .A2(n204), .A3(\mem[15][7] ), .A4(n964), .Y(
        n817) );
  AO21X1_HVT U792 ( .A1(n107), .A2(n282), .A3(n179), .Y(n559) );
  AND2X1_HVT U793 ( .A1(n556), .A2(n554), .Y(n282) );
  AND2X1_HVT U794 ( .A1(a_addr[2]), .A2(n158), .Y(n556) );
  AO22X1_HVT U795 ( .A1(n560), .A2(n204), .A3(\mem[15][8] ), .A4(n963), .Y(
        n818) );
  AO21X1_HVT U796 ( .A1(n106), .A2(n284), .A3(n179), .Y(n560) );
  AND2X1_HVT U797 ( .A1(n561), .A2(n548), .Y(n284) );
  AO22X1_HVT U798 ( .A1(n562), .A2(n204), .A3(\mem[15][9] ), .A4(n962), .Y(
        n819) );
  AO21X1_HVT U799 ( .A1(n105), .A2(n286), .A3(n180), .Y(n562) );
  AND2X1_HVT U800 ( .A1(n561), .A2(n550), .Y(n286) );
  AO22X1_HVT U801 ( .A1(n563), .A2(n204), .A3(\mem[15][10] ), .A4(n961), .Y(
        n820) );
  AO21X1_HVT U802 ( .A1(n107), .A2(n288), .A3(n180), .Y(n563) );
  AND2X1_HVT U803 ( .A1(n561), .A2(n552), .Y(n288) );
  AO22X1_HVT U804 ( .A1(n564), .A2(n204), .A3(\mem[15][11] ), .A4(n960), .Y(
        n821) );
  AO21X1_HVT U805 ( .A1(n106), .A2(n290), .A3(n180), .Y(n564) );
  AND2X1_HVT U806 ( .A1(n561), .A2(n554), .Y(n290) );
  AND2X1_HVT U807 ( .A1(n157), .A2(n156), .Y(n561) );
  AO22X1_HVT U808 ( .A1(n565), .A2(n205), .A3(\mem[15][12] ), .A4(n959), .Y(
        n822) );
  AO21X1_HVT U809 ( .A1(n105), .A2(n292), .A3(n180), .Y(n565) );
  AND2X1_HVT U810 ( .A1(n566), .A2(n548), .Y(n292) );
  AND2X1_HVT U811 ( .A1(n153), .A2(n155), .Y(n548) );
  AO22X1_HVT U812 ( .A1(n567), .A2(n205), .A3(\mem[15][13] ), .A4(n958), .Y(
        n823) );
  AO21X1_HVT U813 ( .A1(n107), .A2(n294), .A3(n180), .Y(n567) );
  AND2X1_HVT U814 ( .A1(n566), .A2(n550), .Y(n294) );
  AND2X1_HVT U815 ( .A1(a_addr[0]), .A2(n155), .Y(n550) );
  AO22X1_HVT U816 ( .A1(n568), .A2(n205), .A3(\mem[15][14] ), .A4(n957), .Y(
        n824) );
  AO21X1_HVT U817 ( .A1(n106), .A2(n296), .A3(n180), .Y(n568) );
  AND2X1_HVT U818 ( .A1(n566), .A2(n552), .Y(n296) );
  AND2X1_HVT U819 ( .A1(n154), .A2(n153), .Y(n552) );
  AO22X1_HVT U820 ( .A1(n569), .A2(n205), .A3(\mem[15][15] ), .A4(n956), .Y(
        n825) );
  AO21X1_HVT U821 ( .A1(n105), .A2(n298), .A3(n180), .Y(n569) );
  AND2X1_HVT U822 ( .A1(n566), .A2(n554), .Y(n298) );
  AND2X1_HVT U823 ( .A1(n154), .A2(a_addr[0]), .Y(n554) );
  AND2X1_HVT U824 ( .A1(n157), .A2(a_addr[2]), .Y(n566) );
  AND3X1_HVT U825 ( .A1(n354), .A2(n3), .A3(n510), .Y(n546) );
  AND2X1_HVT U826 ( .A1(a_din[3]), .A2(a_din[2]), .Y(n510) );
  AND2X1_HVT U827 ( .A1(n151), .A2(a_din[0]), .Y(n354) );
  INVX0_HVT U3 ( .A(N17), .Y(n1) );
  INVX1_HVT U4 ( .A(n1), .Y(n2) );
  INVX0_HVT U5 ( .A(n161), .Y(n3) );
  INVX0_HVT U6 ( .A(n161), .Y(n4) );
  INVX0_HVT U7 ( .A(n161), .Y(n159) );
  IBUFFX2_HVT U8 ( .A(write), .Y(n161) );
  INVX1_HVT U9 ( .A(n184), .Y(n190) );
  INVX1_HVT U10 ( .A(n184), .Y(n191) );
  INVX1_HVT U11 ( .A(n184), .Y(n192) );
  INVX1_HVT U12 ( .A(n184), .Y(n193) );
  INVX1_HVT U13 ( .A(n162), .Y(n194) );
  INVX1_HVT U14 ( .A(n184), .Y(n195) );
  INVX1_HVT U15 ( .A(n180), .Y(n196) );
  INVX1_HVT U16 ( .A(n162), .Y(n197) );
  INVX1_HVT U17 ( .A(n184), .Y(n198) );
  INVX1_HVT U18 ( .A(n180), .Y(n199) );
  INVX1_HVT U19 ( .A(n162), .Y(n200) );
  INVX1_HVT U20 ( .A(n162), .Y(n201) );
  INVX1_HVT U21 ( .A(n162), .Y(n202) );
  INVX1_HVT U22 ( .A(n162), .Y(n203) );
  INVX1_HVT U23 ( .A(n162), .Y(n204) );
  INVX1_HVT U24 ( .A(n162), .Y(n205) );
  INVX1_HVT U25 ( .A(n163), .Y(n186) );
  INVX1_HVT U26 ( .A(n163), .Y(n187) );
  INVX1_HVT U27 ( .A(n163), .Y(n188) );
  INVX1_HVT U28 ( .A(n163), .Y(n189) );
  INVX1_HVT U29 ( .A(n161), .Y(n160) );
  INVX1_HVT U30 ( .A(n185), .Y(n162) );
  INVX1_HVT U31 ( .A(n183), .Y(n168) );
  INVX1_HVT U32 ( .A(n182), .Y(n174) );
  INVX1_HVT U33 ( .A(n181), .Y(n179) );
  INVX1_HVT U34 ( .A(n183), .Y(n164) );
  INVX1_HVT U35 ( .A(n183), .Y(n165) );
  INVX1_HVT U36 ( .A(n183), .Y(n166) );
  INVX1_HVT U37 ( .A(n183), .Y(n167) );
  INVX1_HVT U38 ( .A(n182), .Y(n169) );
  INVX1_HVT U39 ( .A(n182), .Y(n170) );
  INVX1_HVT U40 ( .A(n182), .Y(n171) );
  INVX1_HVT U41 ( .A(n182), .Y(n172) );
  INVX1_HVT U42 ( .A(n182), .Y(n173) );
  INVX1_HVT U43 ( .A(n181), .Y(n175) );
  INVX1_HVT U44 ( .A(n181), .Y(n176) );
  INVX1_HVT U45 ( .A(n181), .Y(n177) );
  INVX1_HVT U46 ( .A(n181), .Y(n178) );
  INVX1_HVT U47 ( .A(n183), .Y(n163) );
  INVX1_HVT U48 ( .A(n181), .Y(n180) );
  INVX1_HVT U49 ( .A(n184), .Y(n183) );
  INVX1_HVT U50 ( .A(n184), .Y(n182) );
  INVX1_HVT U51 ( .A(n184), .Y(n181) );
  NBUFFX2_HVT U52 ( .A(n268), .Y(n147) );
  NBUFFX2_HVT U53 ( .A(n268), .Y(n149) );
  NBUFFX2_HVT U54 ( .A(n268), .Y(n148) );
  INVX1_HVT U55 ( .A(n5), .Y(n144) );
  INVX1_HVT U56 ( .A(n5), .Y(n143) );
  INVX1_HVT U57 ( .A(n185), .Y(n184) );
  INVX1_HVT U58 ( .A(rst), .Y(n185) );
  INVX1_HVT U59 ( .A(n158), .Y(n157) );
  INVX1_HVT U60 ( .A(n155), .Y(n154) );
  NBUFFX2_HVT U61 ( .A(n460), .Y(n120) );
  NBUFFX2_HVT U62 ( .A(n529), .Y(n108) );
  NBUFFX2_HVT U63 ( .A(n356), .Y(n138) );
  NBUFFX2_HVT U64 ( .A(n391), .Y(n132) );
  NBUFFX2_HVT U65 ( .A(n425), .Y(n126) );
  NBUFFX2_HVT U66 ( .A(n494), .Y(n114) );
  NBUFFX2_HVT U67 ( .A(n460), .Y(n122) );
  NBUFFX2_HVT U68 ( .A(n460), .Y(n121) );
  NBUFFX2_HVT U69 ( .A(n529), .Y(n110) );
  NBUFFX2_HVT U70 ( .A(n529), .Y(n109) );
  NBUFFX2_HVT U71 ( .A(n356), .Y(n140) );
  NBUFFX2_HVT U72 ( .A(n356), .Y(n139) );
  NBUFFX2_HVT U73 ( .A(n391), .Y(n134) );
  NBUFFX2_HVT U74 ( .A(n391), .Y(n133) );
  NBUFFX2_HVT U75 ( .A(n425), .Y(n128) );
  NBUFFX2_HVT U76 ( .A(n425), .Y(n127) );
  NBUFFX2_HVT U77 ( .A(n494), .Y(n116) );
  NBUFFX2_HVT U78 ( .A(n494), .Y(n115) );
  NBUFFX2_HVT U79 ( .A(n546), .Y(n105) );
  NBUFFX2_HVT U80 ( .A(n374), .Y(n135) );
  NBUFFX2_HVT U81 ( .A(n443), .Y(n123) );
  NBUFFX2_HVT U82 ( .A(n408), .Y(n129) );
  NBUFFX2_HVT U83 ( .A(n477), .Y(n117) );
  NBUFFX2_HVT U84 ( .A(n512), .Y(n111) );
  NBUFFX2_HVT U85 ( .A(n546), .Y(n107) );
  NBUFFX2_HVT U86 ( .A(n546), .Y(n106) );
  NBUFFX2_HVT U87 ( .A(n374), .Y(n137) );
  NBUFFX2_HVT U88 ( .A(n374), .Y(n136) );
  NBUFFX2_HVT U89 ( .A(n408), .Y(n131) );
  NBUFFX2_HVT U90 ( .A(n408), .Y(n130) );
  NBUFFX2_HVT U91 ( .A(n477), .Y(n119) );
  NBUFFX2_HVT U92 ( .A(n477), .Y(n118) );
  NBUFFX2_HVT U93 ( .A(n443), .Y(n125) );
  NBUFFX2_HVT U94 ( .A(n443), .Y(n124) );
  NBUFFX2_HVT U95 ( .A(n512), .Y(n113) );
  NBUFFX2_HVT U96 ( .A(n512), .Y(n112) );
  NAND3X0_HVT U97 ( .A1(n300), .A2(n4), .A3(n336), .Y(n5) );
  INVX1_HVT U98 ( .A(n6), .Y(n142) );
  INVX1_HVT U99 ( .A(n6), .Y(n141) );
  INVX1_HVT U100 ( .A(n7), .Y(n146) );
  INVX1_HVT U101 ( .A(n7), .Y(n145) );
  INVX1_HVT U102 ( .A(a_addr[1]), .Y(n155) );
  INVX1_HVT U103 ( .A(a_addr[3]), .Y(n158) );
  INVX1_HVT U104 ( .A(a_addr[2]), .Y(n156) );
  INVX1_HVT U105 ( .A(a_addr[0]), .Y(n153) );
  NBUFFX2_HVT U106 ( .A(n83), .Y(n103) );
  NBUFFX2_HVT U107 ( .A(n83), .Y(n100) );
  NBUFFX2_HVT U108 ( .A(n82), .Y(n97) );
  NBUFFX2_HVT U109 ( .A(n81), .Y(n94) );
  NBUFFX2_HVT U110 ( .A(n80), .Y(n91) );
  NBUFFX2_HVT U111 ( .A(n82), .Y(n104) );
  NBUFFX2_HVT U112 ( .A(n83), .Y(n101) );
  NBUFFX2_HVT U113 ( .A(n82), .Y(n98) );
  NBUFFX2_HVT U114 ( .A(n81), .Y(n95) );
  NBUFFX2_HVT U115 ( .A(n80), .Y(n92) );
  NBUFFX2_HVT U116 ( .A(n81), .Y(n102) );
  NBUFFX2_HVT U117 ( .A(n83), .Y(n99) );
  NBUFFX2_HVT U118 ( .A(n82), .Y(n96) );
  NBUFFX2_HVT U119 ( .A(n81), .Y(n93) );
  NBUFFX2_HVT U120 ( .A(n80), .Y(n90) );
  NAND3X0_HVT U121 ( .A1(n300), .A2(n3), .A3(n354), .Y(n6) );
  NAND3X0_HVT U122 ( .A1(n300), .A2(n160), .A3(n318), .Y(n7) );
  INVX1_HVT U123 ( .A(n72), .Y(n78) );
  INVX1_HVT U124 ( .A(n72), .Y(n77) );
  INVX1_HVT U125 ( .A(n72), .Y(n76) );
  INVX1_HVT U126 ( .A(n72), .Y(n75) );
  INVX1_HVT U127 ( .A(n72), .Y(n74) );
  INVX1_HVT U128 ( .A(n72), .Y(n73) );
  INVX1_HVT U129 ( .A(n86), .Y(n84) );
  INVX1_HVT U130 ( .A(n86), .Y(n85) );
  INVX1_HVT U131 ( .A(n152), .Y(n151) );
  INVX1_HVT U132 ( .A(n89), .Y(n87) );
  INVX1_HVT U133 ( .A(n89), .Y(n88) );
  INVX0_HVT U134 ( .A(a_din[0]), .Y(n150) );
  NBUFFX2_HVT U135 ( .A(n2), .Y(n83) );
  NBUFFX2_HVT U136 ( .A(n2), .Y(n82) );
  NBUFFX2_HVT U137 ( .A(n2), .Y(n81) );
  NBUFFX2_HVT U138 ( .A(n2), .Y(n80) );
  NBUFFX2_HVT U139 ( .A(n2), .Y(n79) );
  INVX1_HVT U140 ( .A(N18), .Y(n72) );
  INVX0_HVT U141 ( .A(N19), .Y(n86) );
  INVX0_HVT U142 ( .A(a_din[1]), .Y(n152) );
  INVX0_HVT U143 ( .A(N20), .Y(n89) );
  MUX41X1_HVT U144 ( .A1(\mem[12][0] ), .A3(\mem[14][0] ), .A2(\mem[13][0] ), 
        .A4(\mem[15][0] ), .S0(n78), .S1(n103), .Y(n8) );
  MUX41X1_HVT U145 ( .A1(\mem[8][0] ), .A3(\mem[10][0] ), .A2(\mem[9][0] ), 
        .A4(\mem[11][0] ), .S0(n78), .S1(n102), .Y(n9) );
  MUX41X1_HVT U146 ( .A1(\mem[4][0] ), .A3(\mem[6][0] ), .A2(\mem[5][0] ), 
        .A4(\mem[7][0] ), .S0(n78), .S1(n103), .Y(n10) );
  MUX41X1_HVT U147 ( .A1(\mem[0][0] ), .A3(\mem[2][0] ), .A2(\mem[1][0] ), 
        .A4(\mem[3][0] ), .S0(n78), .S1(n102), .Y(n11) );
  MUX41X1_HVT U148 ( .A1(n11), .A3(n9), .A2(n10), .A4(n8), .S0(n87), .S1(n84), 
        .Y(N554) );
  MUX41X1_HVT U149 ( .A1(\mem[12][1] ), .A3(\mem[14][1] ), .A2(\mem[13][1] ), 
        .A4(\mem[15][1] ), .S0(n78), .S1(n103), .Y(n12) );
  MUX41X1_HVT U150 ( .A1(\mem[8][1] ), .A3(\mem[10][1] ), .A2(\mem[9][1] ), 
        .A4(\mem[11][1] ), .S0(n78), .S1(n102), .Y(n13) );
  MUX41X1_HVT U151 ( .A1(\mem[4][1] ), .A3(\mem[6][1] ), .A2(\mem[5][1] ), 
        .A4(\mem[7][1] ), .S0(n78), .S1(n103), .Y(n14) );
  MUX41X1_HVT U152 ( .A1(\mem[0][1] ), .A3(\mem[2][1] ), .A2(\mem[1][1] ), 
        .A4(\mem[3][1] ), .S0(n78), .S1(n102), .Y(n15) );
  MUX41X1_HVT U153 ( .A1(n15), .A3(n13), .A2(n14), .A4(n12), .S0(n87), .S1(n84), .Y(N553) );
  MUX41X1_HVT U154 ( .A1(\mem[12][2] ), .A3(\mem[14][2] ), .A2(\mem[13][2] ), 
        .A4(\mem[15][2] ), .S0(n78), .S1(n104), .Y(n16) );
  MUX41X1_HVT U155 ( .A1(\mem[8][2] ), .A3(\mem[10][2] ), .A2(\mem[9][2] ), 
        .A4(\mem[11][2] ), .S0(n78), .S1(n104), .Y(n17) );
  MUX41X1_HVT U156 ( .A1(\mem[4][2] ), .A3(\mem[6][2] ), .A2(\mem[5][2] ), 
        .A4(\mem[7][2] ), .S0(n78), .S1(n104), .Y(n18) );
  MUX41X1_HVT U157 ( .A1(\mem[0][2] ), .A3(\mem[2][2] ), .A2(\mem[1][2] ), 
        .A4(\mem[3][2] ), .S0(n78), .S1(n104), .Y(n19) );
  MUX41X1_HVT U158 ( .A1(n19), .A3(n17), .A2(n18), .A4(n16), .S0(n87), .S1(n84), .Y(N552) );
  MUX41X1_HVT U159 ( .A1(\mem[12][3] ), .A3(\mem[14][3] ), .A2(\mem[13][3] ), 
        .A4(\mem[15][3] ), .S0(n77), .S1(n100), .Y(n20) );
  MUX41X1_HVT U160 ( .A1(\mem[8][3] ), .A3(\mem[10][3] ), .A2(\mem[9][3] ), 
        .A4(\mem[11][3] ), .S0(n77), .S1(n99), .Y(n21) );
  MUX41X1_HVT U161 ( .A1(\mem[4][3] ), .A3(\mem[6][3] ), .A2(\mem[5][3] ), 
        .A4(\mem[7][3] ), .S0(n77), .S1(n100), .Y(n22) );
  MUX41X1_HVT U162 ( .A1(\mem[0][3] ), .A3(\mem[2][3] ), .A2(\mem[1][3] ), 
        .A4(\mem[3][3] ), .S0(n77), .S1(n99), .Y(n23) );
  MUX41X1_HVT U163 ( .A1(n23), .A3(n21), .A2(n22), .A4(n20), .S0(n87), .S1(n84), .Y(N551) );
  MUX41X1_HVT U164 ( .A1(\mem[12][4] ), .A3(\mem[14][4] ), .A2(\mem[13][4] ), 
        .A4(\mem[15][4] ), .S0(n77), .S1(n100), .Y(n24) );
  MUX41X1_HVT U165 ( .A1(\mem[8][4] ), .A3(\mem[10][4] ), .A2(\mem[9][4] ), 
        .A4(\mem[11][4] ), .S0(n77), .S1(n99), .Y(n25) );
  MUX41X1_HVT U166 ( .A1(\mem[4][4] ), .A3(\mem[6][4] ), .A2(\mem[5][4] ), 
        .A4(\mem[7][4] ), .S0(n77), .S1(n100), .Y(n26) );
  MUX41X1_HVT U167 ( .A1(\mem[0][4] ), .A3(\mem[2][4] ), .A2(\mem[1][4] ), 
        .A4(\mem[3][4] ), .S0(n77), .S1(n99), .Y(n27) );
  MUX41X1_HVT U168 ( .A1(n27), .A3(n25), .A2(n26), .A4(n24), .S0(n87), .S1(n84), .Y(N550) );
  MUX41X1_HVT U169 ( .A1(\mem[12][5] ), .A3(\mem[14][5] ), .A2(\mem[13][5] ), 
        .A4(\mem[15][5] ), .S0(n77), .S1(n101), .Y(n28) );
  MUX41X1_HVT U170 ( .A1(\mem[8][5] ), .A3(\mem[10][5] ), .A2(\mem[9][5] ), 
        .A4(\mem[11][5] ), .S0(n77), .S1(n101), .Y(n29) );
  MUX41X1_HVT U171 ( .A1(\mem[4][5] ), .A3(\mem[6][5] ), .A2(\mem[5][5] ), 
        .A4(\mem[7][5] ), .S0(n77), .S1(n101), .Y(n30) );
  MUX41X1_HVT U172 ( .A1(\mem[0][5] ), .A3(\mem[2][5] ), .A2(\mem[1][5] ), 
        .A4(\mem[3][5] ), .S0(n77), .S1(n101), .Y(n31) );
  MUX41X1_HVT U173 ( .A1(n31), .A3(n29), .A2(n30), .A4(n28), .S0(n87), .S1(n84), .Y(N549) );
  MUX41X1_HVT U174 ( .A1(\mem[12][6] ), .A3(\mem[14][6] ), .A2(\mem[13][6] ), 
        .A4(\mem[15][6] ), .S0(n76), .S1(n97), .Y(n32) );
  MUX41X1_HVT U175 ( .A1(\mem[8][6] ), .A3(\mem[10][6] ), .A2(\mem[9][6] ), 
        .A4(\mem[11][6] ), .S0(n76), .S1(n96), .Y(n33) );
  MUX41X1_HVT U176 ( .A1(\mem[4][6] ), .A3(\mem[6][6] ), .A2(\mem[5][6] ), 
        .A4(\mem[7][6] ), .S0(n76), .S1(n97), .Y(n34) );
  MUX41X1_HVT U177 ( .A1(\mem[0][6] ), .A3(\mem[2][6] ), .A2(\mem[1][6] ), 
        .A4(\mem[3][6] ), .S0(n76), .S1(n96), .Y(n35) );
  MUX41X1_HVT U178 ( .A1(n35), .A3(n33), .A2(n34), .A4(n32), .S0(n87), .S1(n84), .Y(N548) );
  MUX41X1_HVT U179 ( .A1(\mem[12][7] ), .A3(\mem[14][7] ), .A2(\mem[13][7] ), 
        .A4(\mem[15][7] ), .S0(n76), .S1(n97), .Y(n36) );
  MUX41X1_HVT U180 ( .A1(\mem[8][7] ), .A3(\mem[10][7] ), .A2(\mem[9][7] ), 
        .A4(\mem[11][7] ), .S0(n76), .S1(n96), .Y(n37) );
  MUX41X1_HVT U181 ( .A1(\mem[4][7] ), .A3(\mem[6][7] ), .A2(\mem[5][7] ), 
        .A4(\mem[7][7] ), .S0(n76), .S1(n97), .Y(n38) );
  MUX41X1_HVT U182 ( .A1(\mem[0][7] ), .A3(\mem[2][7] ), .A2(\mem[1][7] ), 
        .A4(\mem[3][7] ), .S0(n76), .S1(n96), .Y(n39) );
  MUX41X1_HVT U183 ( .A1(n39), .A3(n37), .A2(n38), .A4(n36), .S0(n87), .S1(n84), .Y(N547) );
  MUX41X1_HVT U184 ( .A1(\mem[12][8] ), .A3(\mem[14][8] ), .A2(\mem[13][8] ), 
        .A4(\mem[15][8] ), .S0(n76), .S1(n98), .Y(n40) );
  MUX41X1_HVT U185 ( .A1(\mem[8][8] ), .A3(\mem[10][8] ), .A2(\mem[9][8] ), 
        .A4(\mem[11][8] ), .S0(n76), .S1(n98), .Y(n41) );
  MUX41X1_HVT U186 ( .A1(\mem[4][8] ), .A3(\mem[6][8] ), .A2(\mem[5][8] ), 
        .A4(\mem[7][8] ), .S0(n76), .S1(n98), .Y(n42) );
  MUX41X1_HVT U187 ( .A1(\mem[0][8] ), .A3(\mem[2][8] ), .A2(\mem[1][8] ), 
        .A4(\mem[3][8] ), .S0(n76), .S1(n98), .Y(n43) );
  MUX41X1_HVT U188 ( .A1(n43), .A3(n41), .A2(n42), .A4(n40), .S0(n88), .S1(n85), .Y(N546) );
  MUX41X1_HVT U189 ( .A1(\mem[12][9] ), .A3(\mem[14][9] ), .A2(\mem[13][9] ), 
        .A4(\mem[15][9] ), .S0(n75), .S1(n94), .Y(n44) );
  MUX41X1_HVT U190 ( .A1(\mem[8][9] ), .A3(\mem[10][9] ), .A2(\mem[9][9] ), 
        .A4(\mem[11][9] ), .S0(n75), .S1(n93), .Y(n45) );
  MUX41X1_HVT U191 ( .A1(\mem[4][9] ), .A3(\mem[6][9] ), .A2(\mem[5][9] ), 
        .A4(\mem[7][9] ), .S0(n75), .S1(n94), .Y(n46) );
  MUX41X1_HVT U192 ( .A1(\mem[0][9] ), .A3(\mem[2][9] ), .A2(\mem[1][9] ), 
        .A4(\mem[3][9] ), .S0(n75), .S1(n93), .Y(n47) );
  MUX41X1_HVT U193 ( .A1(n47), .A3(n45), .A2(n46), .A4(n44), .S0(n88), .S1(n85), .Y(N545) );
  MUX41X1_HVT U194 ( .A1(\mem[12][10] ), .A3(\mem[14][10] ), .A2(\mem[13][10] ), .A4(\mem[15][10] ), .S0(n75), .S1(n94), .Y(n48) );
  MUX41X1_HVT U195 ( .A1(\mem[8][10] ), .A3(\mem[10][10] ), .A2(\mem[9][10] ), 
        .A4(\mem[11][10] ), .S0(n75), .S1(n93), .Y(n49) );
  MUX41X1_HVT U196 ( .A1(\mem[4][10] ), .A3(\mem[6][10] ), .A2(\mem[5][10] ), 
        .A4(\mem[7][10] ), .S0(n75), .S1(n94), .Y(n50) );
  MUX41X1_HVT U197 ( .A1(\mem[0][10] ), .A3(\mem[2][10] ), .A2(\mem[1][10] ), 
        .A4(\mem[3][10] ), .S0(n75), .S1(n93), .Y(n51) );
  MUX41X1_HVT U198 ( .A1(n51), .A3(n49), .A2(n50), .A4(n48), .S0(n88), .S1(n85), .Y(N544) );
  MUX41X1_HVT U199 ( .A1(\mem[12][11] ), .A3(\mem[14][11] ), .A2(\mem[13][11] ), .A4(\mem[15][11] ), .S0(n75), .S1(n95), .Y(n52) );
  MUX41X1_HVT U200 ( .A1(\mem[8][11] ), .A3(\mem[10][11] ), .A2(\mem[9][11] ), 
        .A4(\mem[11][11] ), .S0(n75), .S1(n95), .Y(n53) );
  MUX41X1_HVT U201 ( .A1(\mem[4][11] ), .A3(\mem[6][11] ), .A2(\mem[5][11] ), 
        .A4(\mem[7][11] ), .S0(n75), .S1(n95), .Y(n54) );
  MUX41X1_HVT U202 ( .A1(\mem[0][11] ), .A3(\mem[2][11] ), .A2(\mem[1][11] ), 
        .A4(\mem[3][11] ), .S0(n75), .S1(n95), .Y(n55) );
  MUX41X1_HVT U203 ( .A1(n55), .A3(n53), .A2(n54), .A4(n52), .S0(n88), .S1(n85), .Y(N543) );
  MUX41X1_HVT U204 ( .A1(\mem[12][12] ), .A3(\mem[14][12] ), .A2(\mem[13][12] ), .A4(\mem[15][12] ), .S0(n74), .S1(n91), .Y(n56) );
  MUX41X1_HVT U205 ( .A1(\mem[8][12] ), .A3(\mem[10][12] ), .A2(\mem[9][12] ), 
        .A4(\mem[11][12] ), .S0(n74), .S1(n90), .Y(n57) );
  MUX41X1_HVT U206 ( .A1(\mem[4][12] ), .A3(\mem[6][12] ), .A2(\mem[5][12] ), 
        .A4(\mem[7][12] ), .S0(n74), .S1(n91), .Y(n58) );
  MUX41X1_HVT U207 ( .A1(\mem[0][12] ), .A3(\mem[2][12] ), .A2(\mem[1][12] ), 
        .A4(\mem[3][12] ), .S0(n74), .S1(n90), .Y(n59) );
  MUX41X1_HVT U208 ( .A1(n59), .A3(n57), .A2(n58), .A4(n56), .S0(n88), .S1(n85), .Y(N542) );
  MUX41X1_HVT U209 ( .A1(\mem[12][13] ), .A3(\mem[14][13] ), .A2(\mem[13][13] ), .A4(\mem[15][13] ), .S0(n74), .S1(n91), .Y(n60) );
  MUX41X1_HVT U210 ( .A1(\mem[8][13] ), .A3(\mem[10][13] ), .A2(\mem[9][13] ), 
        .A4(\mem[11][13] ), .S0(n74), .S1(n90), .Y(n61) );
  MUX41X1_HVT U211 ( .A1(\mem[4][13] ), .A3(\mem[6][13] ), .A2(\mem[5][13] ), 
        .A4(\mem[7][13] ), .S0(n74), .S1(n91), .Y(n62) );
  MUX41X1_HVT U212 ( .A1(\mem[0][13] ), .A3(\mem[2][13] ), .A2(\mem[1][13] ), 
        .A4(\mem[3][13] ), .S0(n74), .S1(n90), .Y(n63) );
  MUX41X1_HVT U213 ( .A1(n63), .A3(n61), .A2(n62), .A4(n60), .S0(n88), .S1(n85), .Y(N541) );
  MUX41X1_HVT U214 ( .A1(\mem[12][14] ), .A3(\mem[14][14] ), .A2(\mem[13][14] ), .A4(\mem[15][14] ), .S0(n74), .S1(n92), .Y(n64) );
  MUX41X1_HVT U215 ( .A1(\mem[8][14] ), .A3(\mem[10][14] ), .A2(\mem[9][14] ), 
        .A4(\mem[11][14] ), .S0(n74), .S1(n92), .Y(n65) );
  MUX41X1_HVT U216 ( .A1(\mem[4][14] ), .A3(\mem[6][14] ), .A2(\mem[5][14] ), 
        .A4(\mem[7][14] ), .S0(n74), .S1(n92), .Y(n66) );
  MUX41X1_HVT U217 ( .A1(\mem[0][14] ), .A3(\mem[2][14] ), .A2(\mem[1][14] ), 
        .A4(\mem[3][14] ), .S0(n74), .S1(n92), .Y(n67) );
  MUX41X1_HVT U218 ( .A1(n67), .A3(n65), .A2(n66), .A4(n64), .S0(n88), .S1(n85), .Y(N540) );
  MUX41X1_HVT U219 ( .A1(\mem[12][15] ), .A3(\mem[14][15] ), .A2(\mem[13][15] ), .A4(\mem[15][15] ), .S0(n73), .S1(n79), .Y(n68) );
  MUX41X1_HVT U220 ( .A1(\mem[8][15] ), .A3(\mem[10][15] ), .A2(\mem[9][15] ), 
        .A4(\mem[11][15] ), .S0(n73), .S1(n79), .Y(n69) );
  MUX41X1_HVT U221 ( .A1(\mem[4][15] ), .A3(\mem[6][15] ), .A2(\mem[5][15] ), 
        .A4(\mem[7][15] ), .S0(n73), .S1(n79), .Y(n70) );
  MUX41X1_HVT U222 ( .A1(\mem[0][15] ), .A3(\mem[2][15] ), .A2(\mem[1][15] ), 
        .A4(\mem[3][15] ), .S0(n73), .S1(n79), .Y(n71) );
  MUX41X1_HVT U223 ( .A1(n71), .A3(n69), .A2(n70), .A4(n68), .S0(n88), .S1(n85), .Y(N539) );
  INVX0_HVT U224 ( .A(n423), .Y(n206) );
  INVX0_HVT U225 ( .A(n422), .Y(n207) );
  INVX0_HVT U226 ( .A(n421), .Y(n208) );
  INVX0_HVT U227 ( .A(n420), .Y(n209) );
  INVX0_HVT U228 ( .A(n419), .Y(n210) );
  INVX0_HVT U229 ( .A(n418), .Y(n211) );
  INVX0_HVT U230 ( .A(n417), .Y(n212) );
  INVX0_HVT U231 ( .A(n416), .Y(n213) );
  INVX0_HVT U232 ( .A(n415), .Y(n214) );
  INVX0_HVT U233 ( .A(n414), .Y(n215) );
  INVX0_HVT U234 ( .A(n413), .Y(n216) );
  INVX0_HVT U235 ( .A(n412), .Y(n217) );
  INVX0_HVT U236 ( .A(n411), .Y(n218) );
  INVX0_HVT U237 ( .A(n410), .Y(n219) );
  INVX0_HVT U238 ( .A(n409), .Y(n220) );
  INVX0_HVT U239 ( .A(n407), .Y(n221) );
  INVX0_HVT U240 ( .A(n406), .Y(n222) );
  INVX0_HVT U241 ( .A(n405), .Y(n223) );
  INVX0_HVT U242 ( .A(n404), .Y(n224) );
  INVX0_HVT U243 ( .A(n403), .Y(n225) );
  INVX0_HVT U244 ( .A(n402), .Y(n226) );
  INVX0_HVT U245 ( .A(n401), .Y(n227) );
  INVX0_HVT U246 ( .A(n400), .Y(n228) );
  INVX0_HVT U247 ( .A(n399), .Y(n229) );
  INVX0_HVT U248 ( .A(n398), .Y(n230) );
  INVX0_HVT U249 ( .A(n397), .Y(n231) );
  INVX0_HVT U250 ( .A(n396), .Y(n232) );
  INVX0_HVT U251 ( .A(n395), .Y(n233) );
  INVX0_HVT U252 ( .A(n394), .Y(n234) );
  INVX0_HVT U253 ( .A(n393), .Y(n235) );
  INVX0_HVT U254 ( .A(n392), .Y(n236) );
  INVX0_HVT U255 ( .A(n390), .Y(n237) );
  INVX0_HVT U256 ( .A(n389), .Y(n238) );
  INVX0_HVT U257 ( .A(n388), .Y(n239) );
  INVX0_HVT U258 ( .A(n387), .Y(n240) );
  INVX0_HVT U259 ( .A(n386), .Y(n241) );
  INVX0_HVT U260 ( .A(n385), .Y(n242) );
  INVX0_HVT U261 ( .A(n384), .Y(n243) );
  INVX0_HVT U262 ( .A(n383), .Y(n244) );
  INVX0_HVT U263 ( .A(n382), .Y(n245) );
  INVX0_HVT U264 ( .A(n381), .Y(n246) );
  INVX0_HVT U265 ( .A(n380), .Y(n247) );
  INVX0_HVT U266 ( .A(n379), .Y(n248) );
  INVX0_HVT U267 ( .A(n378), .Y(n249) );
  INVX0_HVT U333 ( .A(n377), .Y(n250) );
  INVX0_HVT U366 ( .A(n376), .Y(n251) );
  INVX0_HVT U399 ( .A(n375), .Y(n252) );
  INVX0_HVT U828 ( .A(n373), .Y(n253) );
  INVX0_HVT U829 ( .A(n371), .Y(n254) );
  INVX0_HVT U830 ( .A(n370), .Y(n255) );
  INVX0_HVT U831 ( .A(n369), .Y(n256) );
  INVX0_HVT U832 ( .A(n368), .Y(n257) );
  INVX0_HVT U833 ( .A(n367), .Y(n258) );
  INVX0_HVT U834 ( .A(n366), .Y(n259) );
  INVX0_HVT U835 ( .A(n365), .Y(n260) );
  INVX0_HVT U836 ( .A(n364), .Y(n261) );
  INVX0_HVT U837 ( .A(n363), .Y(n262) );
  INVX0_HVT U838 ( .A(n362), .Y(n263) );
  INVX0_HVT U839 ( .A(n361), .Y(n264) );
  INVX0_HVT U840 ( .A(n360), .Y(n265) );
  INVX0_HVT U841 ( .A(n359), .Y(n302) );
  INVX0_HVT U842 ( .A(n358), .Y(n320) );
  INVX0_HVT U843 ( .A(n357), .Y(n338) );
  INVX0_HVT U844 ( .A(n355), .Y(n826) );
  INVX0_HVT U845 ( .A(n353), .Y(n827) );
  INVX0_HVT U846 ( .A(n352), .Y(n828) );
  INVX0_HVT U847 ( .A(n351), .Y(n829) );
  INVX0_HVT U848 ( .A(n350), .Y(n830) );
  INVX0_HVT U849 ( .A(n349), .Y(n831) );
  INVX0_HVT U850 ( .A(n348), .Y(n832) );
  INVX0_HVT U851 ( .A(n347), .Y(n833) );
  INVX0_HVT U852 ( .A(n346), .Y(n834) );
  INVX0_HVT U853 ( .A(n345), .Y(n835) );
  INVX0_HVT U854 ( .A(n344), .Y(n836) );
  INVX0_HVT U855 ( .A(n343), .Y(n837) );
  INVX0_HVT U856 ( .A(n342), .Y(n838) );
  INVX0_HVT U857 ( .A(n341), .Y(n839) );
  INVX0_HVT U858 ( .A(n340), .Y(n840) );
  INVX0_HVT U859 ( .A(n339), .Y(n841) );
  INVX0_HVT U860 ( .A(n337), .Y(n842) );
  INVX0_HVT U861 ( .A(n335), .Y(n843) );
  INVX0_HVT U862 ( .A(n334), .Y(n844) );
  INVX0_HVT U863 ( .A(n333), .Y(n845) );
  INVX0_HVT U864 ( .A(n332), .Y(n846) );
  INVX0_HVT U865 ( .A(n331), .Y(n847) );
  INVX0_HVT U866 ( .A(n330), .Y(n848) );
  INVX0_HVT U867 ( .A(n329), .Y(n849) );
  INVX0_HVT U868 ( .A(n328), .Y(n850) );
  INVX0_HVT U869 ( .A(n327), .Y(n851) );
  INVX0_HVT U870 ( .A(n326), .Y(n852) );
  INVX0_HVT U871 ( .A(n325), .Y(n853) );
  INVX0_HVT U872 ( .A(n324), .Y(n854) );
  INVX0_HVT U873 ( .A(n323), .Y(n855) );
  INVX0_HVT U874 ( .A(n322), .Y(n856) );
  INVX0_HVT U875 ( .A(n321), .Y(n857) );
  INVX0_HVT U876 ( .A(n319), .Y(n858) );
  INVX0_HVT U877 ( .A(n317), .Y(n859) );
  INVX0_HVT U878 ( .A(n316), .Y(n860) );
  INVX0_HVT U879 ( .A(n315), .Y(n861) );
  INVX0_HVT U880 ( .A(n314), .Y(n862) );
  INVX0_HVT U881 ( .A(n313), .Y(n863) );
  INVX0_HVT U882 ( .A(n312), .Y(n864) );
  INVX0_HVT U883 ( .A(n311), .Y(n865) );
  INVX0_HVT U884 ( .A(n310), .Y(n866) );
  INVX0_HVT U885 ( .A(n309), .Y(n867) );
  INVX0_HVT U886 ( .A(n308), .Y(n868) );
  INVX0_HVT U887 ( .A(n307), .Y(n869) );
  INVX0_HVT U888 ( .A(n306), .Y(n870) );
  INVX0_HVT U889 ( .A(n305), .Y(n871) );
  INVX0_HVT U890 ( .A(n304), .Y(n872) );
  INVX0_HVT U891 ( .A(n303), .Y(n873) );
  INVX0_HVT U892 ( .A(n301), .Y(n874) );
  INVX0_HVT U893 ( .A(n297), .Y(n875) );
  INVX0_HVT U894 ( .A(n295), .Y(n876) );
  INVX0_HVT U895 ( .A(n293), .Y(n877) );
  INVX0_HVT U896 ( .A(n291), .Y(n878) );
  INVX0_HVT U897 ( .A(n289), .Y(n879) );
  INVX0_HVT U898 ( .A(n287), .Y(n880) );
  INVX0_HVT U899 ( .A(n285), .Y(n881) );
  INVX0_HVT U900 ( .A(n283), .Y(n882) );
  INVX0_HVT U901 ( .A(n281), .Y(n883) );
  INVX0_HVT U902 ( .A(n279), .Y(n884) );
  INVX0_HVT U903 ( .A(n277), .Y(n885) );
  INVX0_HVT U904 ( .A(n275), .Y(n886) );
  INVX0_HVT U905 ( .A(n273), .Y(n887) );
  INVX0_HVT U906 ( .A(n271), .Y(n888) );
  INVX0_HVT U907 ( .A(n269), .Y(n889) );
  INVX0_HVT U908 ( .A(n266), .Y(n890) );
  INVX0_HVT U909 ( .A(a_din[3]), .Y(n891) );
  INVX0_HVT U910 ( .A(n492), .Y(n892) );
  INVX0_HVT U911 ( .A(n491), .Y(n893) );
  INVX0_HVT U912 ( .A(n490), .Y(n894) );
  INVX0_HVT U913 ( .A(n489), .Y(n895) );
  INVX0_HVT U914 ( .A(n488), .Y(n896) );
  INVX0_HVT U915 ( .A(n487), .Y(n897) );
  INVX0_HVT U916 ( .A(n486), .Y(n898) );
  INVX0_HVT U917 ( .A(n485), .Y(n899) );
  INVX0_HVT U918 ( .A(n484), .Y(n900) );
  INVX0_HVT U919 ( .A(n483), .Y(n901) );
  INVX0_HVT U920 ( .A(n482), .Y(n902) );
  INVX0_HVT U921 ( .A(n481), .Y(n903) );
  INVX0_HVT U922 ( .A(n480), .Y(n904) );
  INVX0_HVT U923 ( .A(n479), .Y(n905) );
  INVX0_HVT U924 ( .A(n478), .Y(n906) );
  INVX0_HVT U925 ( .A(n476), .Y(n907) );
  INVX0_HVT U926 ( .A(n475), .Y(n908) );
  INVX0_HVT U927 ( .A(n474), .Y(n909) );
  INVX0_HVT U928 ( .A(n473), .Y(n910) );
  INVX0_HVT U929 ( .A(n472), .Y(n911) );
  INVX0_HVT U930 ( .A(n471), .Y(n912) );
  INVX0_HVT U931 ( .A(n470), .Y(n913) );
  INVX0_HVT U932 ( .A(n469), .Y(n914) );
  INVX0_HVT U933 ( .A(n468), .Y(n915) );
  INVX0_HVT U934 ( .A(n467), .Y(n916) );
  INVX0_HVT U935 ( .A(n466), .Y(n917) );
  INVX0_HVT U936 ( .A(n465), .Y(n918) );
  INVX0_HVT U937 ( .A(n464), .Y(n919) );
  INVX0_HVT U938 ( .A(n463), .Y(n920) );
  INVX0_HVT U939 ( .A(n462), .Y(n921) );
  INVX0_HVT U940 ( .A(n461), .Y(n922) );
  INVX0_HVT U941 ( .A(n459), .Y(n923) );
  INVX0_HVT U942 ( .A(n458), .Y(n924) );
  INVX0_HVT U943 ( .A(n457), .Y(n925) );
  INVX0_HVT U944 ( .A(n456), .Y(n926) );
  INVX0_HVT U945 ( .A(n455), .Y(n927) );
  INVX0_HVT U946 ( .A(n454), .Y(n928) );
  INVX0_HVT U947 ( .A(n453), .Y(n929) );
  INVX0_HVT U948 ( .A(n452), .Y(n930) );
  INVX0_HVT U949 ( .A(n451), .Y(n931) );
  INVX0_HVT U950 ( .A(n450), .Y(n932) );
  INVX0_HVT U951 ( .A(n449), .Y(n933) );
  INVX0_HVT U952 ( .A(n448), .Y(n934) );
  INVX0_HVT U953 ( .A(n447), .Y(n935) );
  INVX0_HVT U954 ( .A(n446), .Y(n936) );
  INVX0_HVT U955 ( .A(n445), .Y(n937) );
  INVX0_HVT U956 ( .A(n444), .Y(n938) );
  INVX0_HVT U957 ( .A(n442), .Y(n939) );
  INVX0_HVT U958 ( .A(n440), .Y(n940) );
  INVX0_HVT U959 ( .A(n439), .Y(n941) );
  INVX0_HVT U960 ( .A(n438), .Y(n942) );
  INVX0_HVT U961 ( .A(n437), .Y(n943) );
  INVX0_HVT U962 ( .A(n436), .Y(n944) );
  INVX0_HVT U963 ( .A(n435), .Y(n945) );
  INVX0_HVT U964 ( .A(n434), .Y(n946) );
  INVX0_HVT U965 ( .A(n433), .Y(n947) );
  INVX0_HVT U966 ( .A(n432), .Y(n948) );
  INVX0_HVT U967 ( .A(n431), .Y(n949) );
  INVX0_HVT U968 ( .A(n430), .Y(n950) );
  INVX0_HVT U969 ( .A(n429), .Y(n951) );
  INVX0_HVT U970 ( .A(n428), .Y(n952) );
  INVX0_HVT U971 ( .A(n427), .Y(n953) );
  INVX0_HVT U972 ( .A(n426), .Y(n954) );
  INVX0_HVT U973 ( .A(n424), .Y(n955) );
  INVX0_HVT U974 ( .A(n569), .Y(n956) );
  INVX0_HVT U975 ( .A(n568), .Y(n957) );
  INVX0_HVT U976 ( .A(n567), .Y(n958) );
  INVX0_HVT U977 ( .A(n565), .Y(n959) );
  INVX0_HVT U978 ( .A(n564), .Y(n960) );
  INVX0_HVT U979 ( .A(n563), .Y(n961) );
  INVX0_HVT U980 ( .A(n562), .Y(n962) );
  INVX0_HVT U981 ( .A(n560), .Y(n963) );
  INVX0_HVT U982 ( .A(n559), .Y(n964) );
  INVX0_HVT U983 ( .A(n558), .Y(n965) );
  INVX0_HVT U984 ( .A(n557), .Y(n966) );
  INVX0_HVT U985 ( .A(n555), .Y(n967) );
  INVX0_HVT U986 ( .A(n553), .Y(n968) );
  INVX0_HVT U987 ( .A(n551), .Y(n969) );
  INVX0_HVT U988 ( .A(n549), .Y(n970) );
  INVX0_HVT U989 ( .A(n545), .Y(n971) );
  INVX0_HVT U990 ( .A(n544), .Y(n972) );
  INVX0_HVT U991 ( .A(n543), .Y(n973) );
  INVX0_HVT U992 ( .A(n542), .Y(n974) );
  INVX0_HVT U993 ( .A(n541), .Y(n975) );
  INVX0_HVT U994 ( .A(n540), .Y(n976) );
  INVX0_HVT U995 ( .A(n539), .Y(n977) );
  INVX0_HVT U996 ( .A(n538), .Y(n978) );
  INVX0_HVT U997 ( .A(n537), .Y(n979) );
  INVX0_HVT U998 ( .A(n536), .Y(n980) );
  INVX0_HVT U999 ( .A(n535), .Y(n981) );
  INVX0_HVT U1000 ( .A(n534), .Y(n982) );
  INVX0_HVT U1001 ( .A(n533), .Y(n983) );
  INVX0_HVT U1002 ( .A(n532), .Y(n984) );
  INVX0_HVT U1003 ( .A(n531), .Y(n985) );
  INVX0_HVT U1004 ( .A(n530), .Y(n986) );
  INVX0_HVT U1005 ( .A(n528), .Y(n987) );
  INVX0_HVT U1006 ( .A(n527), .Y(n988) );
  INVX0_HVT U1007 ( .A(n526), .Y(n989) );
  INVX0_HVT U1008 ( .A(n525), .Y(n990) );
  INVX0_HVT U1009 ( .A(n524), .Y(n991) );
  INVX0_HVT U1010 ( .A(n523), .Y(n992) );
  INVX0_HVT U1011 ( .A(n522), .Y(n993) );
  INVX0_HVT U1012 ( .A(n521), .Y(n994) );
  INVX0_HVT U1013 ( .A(n520), .Y(n995) );
  INVX0_HVT U1014 ( .A(n519), .Y(n996) );
  INVX0_HVT U1015 ( .A(n518), .Y(n997) );
  INVX0_HVT U1016 ( .A(n517), .Y(n998) );
  INVX0_HVT U1017 ( .A(n516), .Y(n999) );
  INVX0_HVT U1018 ( .A(n515), .Y(n1000) );
  INVX0_HVT U1019 ( .A(n514), .Y(n1001) );
  INVX0_HVT U1020 ( .A(n513), .Y(n1002) );
  INVX0_HVT U1021 ( .A(n511), .Y(n1003) );
  INVX0_HVT U1022 ( .A(n509), .Y(n1004) );
  INVX0_HVT U1023 ( .A(n508), .Y(n1005) );
  INVX0_HVT U1024 ( .A(n507), .Y(n1006) );
  INVX0_HVT U1025 ( .A(n506), .Y(n1007) );
  INVX0_HVT U1026 ( .A(n505), .Y(n1008) );
  INVX0_HVT U1027 ( .A(n504), .Y(n1009) );
  INVX0_HVT U1028 ( .A(n503), .Y(n1010) );
  INVX0_HVT U1029 ( .A(n502), .Y(n1011) );
  INVX0_HVT U1030 ( .A(n501), .Y(n1012) );
  INVX0_HVT U1031 ( .A(n500), .Y(n1013) );
  INVX0_HVT U1032 ( .A(n499), .Y(n1014) );
  INVX0_HVT U1033 ( .A(n498), .Y(n1015) );
  INVX0_HVT U1034 ( .A(n497), .Y(n1016) );
  INVX0_HVT U1035 ( .A(n496), .Y(n1017) );
  INVX0_HVT U1036 ( .A(n495), .Y(n1018) );
  INVX0_HVT U1037 ( .A(n493), .Y(n1019) );
  INVX0_HVT U1038 ( .A(a_din[2]), .Y(n1020) );
endmodule

