
module inv_sbox_7 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n1, n6, n196, n197, n198, n199, n200, n201, n202, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584;

  NAND2X0_HVT U5 ( .A1(n582), .A2(n243), .Y(n581) );
  NAND2X0_HVT U6 ( .A1(n235), .A2(n253), .Y(n580) );
  NAND2X0_HVT U7 ( .A1(n304), .A2(n298), .Y(n579) );
  NAND2X0_HVT U8 ( .A1(n234), .A2(n243), .Y(n578) );
  NAND2X0_HVT U9 ( .A1(n268), .A2(n578), .Y(n577) );
  NAND2X0_HVT U10 ( .A1(n268), .A2(n575), .Y(n576) );
  NAND2X0_HVT U11 ( .A1(n223), .A2(n584), .Y(n574) );
  NAND2X0_HVT U12 ( .A1(n234), .A2(n289), .Y(n573) );
  NAND2X0_HVT U13 ( .A1(n298), .A2(n578), .Y(n572) );
  NAND2X0_HVT U15 ( .A1(n265), .A2(n305), .Y(n570) );
  NAND2X0_HVT U19 ( .A1(n234), .A2(n374), .Y(n565) );
  NAND2X0_HVT U32 ( .A1(n292), .A2(n222), .Y(n553) );
  NAND2X0_HVT U35 ( .A1(n578), .A2(n262), .Y(n550) );
  NAND2X0_HVT U38 ( .A1(n289), .A2(n222), .Y(n547) );
  NAND2X0_HVT U42 ( .A1(n262), .A2(n580), .Y(n543) );
  OA21X1_HVT U53 ( .A1(n313), .A2(n535), .A3(n342), .Y(n533) );
  NAND2X0_HVT U55 ( .A1(n298), .A2(n582), .Y(n531) );
  MUX41X1_HVT U56 ( .A1(n355), .A3(n266), .A2(n340), .A4(n531), .S0(n284), 
        .S1(n311), .Y(n530) );
  AO21X1_HVT U60 ( .A1(n525), .A2(n309), .A3(n564), .Y(n526) );
  MUX41X1_HVT U62 ( .A1(n524), .A3(n530), .A2(n528), .A4(n532), .S0(n238), 
        .S1(in[1]), .Y(n523) );
  MUX41X1_HVT U65 ( .A1(n332), .A3(n334), .A2(n333), .A4(n547), .S0(n284), 
        .S1(n309), .Y(n520) );
  NAND2X0_HVT U66 ( .A1(n301), .A2(n247), .Y(n519) );
  MUX41X1_HVT U67 ( .A1(n329), .A3(n356), .A2(n331), .A4(n519), .S0(n288), 
        .S1(n281), .Y(n518) );
  MUX41X1_HVT U68 ( .A1(n329), .A3(n244), .A2(n330), .A4(n253), .S0(n283), 
        .S1(n236), .Y(n517) );
  MUX41X1_HVT U69 ( .A1(n517), .A3(n520), .A2(n518), .A4(n521), .S0(in[5]), 
        .S1(n202), .Y(n516) );
  NAND2X0_HVT U72 ( .A1(n266), .A2(n199), .Y(n514) );
  MUX41X1_HVT U73 ( .A1(n558), .A3(n514), .A2(n357), .A4(n289), .S0(n287), 
        .S1(n280), .Y(n513) );
  NAND2X0_HVT U81 ( .A1(n584), .A2(n579), .Y(n505) );
  AND2X1_HVT U82 ( .A1(n269), .A2(n583), .Y(n504) );
  MUX41X1_HVT U83 ( .A1(n504), .A3(n344), .A2(n360), .A4(n505), .S0(n283), 
        .S1(n309), .Y(n503) );
  MUX41X1_HVT U87 ( .A1(n319), .A3(n276), .A2(n362), .A4(n340), .S0(n282), 
        .S1(n308), .Y(n500) );
  NAND2X0_HVT U89 ( .A1(n223), .A2(n241), .Y(n498) );
  MUX41X1_HVT U90 ( .A1(n373), .A3(n199), .A2(n538), .A4(n498), .S0(n283), 
        .S1(n311), .Y(n497) );
  MUX41X1_HVT U95 ( .A1(n493), .A3(n499), .A2(n497), .A4(n500), .S0(n297), 
        .S1(n202), .Y(n492) );
  MUX41X1_HVT U96 ( .A1(n356), .A3(n572), .A2(n341), .A4(n363), .S0(n284), 
        .S1(n311), .Y(n491) );
  MUX41X1_HVT U98 ( .A1(n490), .A3(n364), .A2(n349), .A4(n557), .S0(n284), 
        .S1(n308), .Y(n489) );
  MUX41X1_HVT U99 ( .A1(n553), .A3(n333), .A2(n537), .A4(n265), .S0(n309), 
        .S1(n281), .Y(n488) );
  NAND2X0_HVT U100 ( .A1(n223), .A2(n248), .Y(n487) );
  MUX41X1_HVT U101 ( .A1(n365), .A3(n573), .A2(n348), .A4(n487), .S0(n309), 
        .S1(n282), .Y(n486) );
  MUX41X1_HVT U102 ( .A1(n486), .A3(n489), .A2(n488), .A4(n491), .S0(n297), 
        .S1(n295), .Y(n485) );
  AND2X1_HVT U104 ( .A1(n199), .A2(n242), .Y(n484) );
  NAND2X0_HVT U114 ( .A1(n268), .A2(n199), .Y(n474) );
  MUX41X1_HVT U115 ( .A1(n474), .A3(n574), .A2(n351), .A4(n583), .S0(n308), 
        .S1(n281), .Y(n473) );
  MUX41X1_HVT U116 ( .A1(n350), .A3(n343), .A2(n316), .A4(n570), .S0(n282), 
        .S1(n311), .Y(n472) );
  NAND2X0_HVT U118 ( .A1(n223), .A2(n244), .Y(n470) );
  MUX41X1_HVT U119 ( .A1(n367), .A3(n471), .A2(n548), .A4(n470), .S0(n282), 
        .S1(n236), .Y(n469) );
  MUX41X1_HVT U120 ( .A1(n469), .A3(n473), .A2(n472), .A4(n475), .S0(n297), 
        .S1(n295), .Y(n468) );
  MUX41X1_HVT U122 ( .A1(n354), .A3(n273), .A2(n539), .A4(n358), .S0(n282), 
        .S1(n311), .Y(n467) );
  MUX41X1_HVT U124 ( .A1(n275), .A3(n466), .A2(n562), .A4(n337), .S0(n237), 
        .S1(n282), .Y(n465) );
  AOI21X1_HVT U127 ( .A1(n286), .A2(n461), .A3(n323), .Y(n462) );
  NAND2X0_HVT U129 ( .A1(in[2]), .A2(n249), .Y(n459) );
  MUX41X1_HVT U130 ( .A1(n459), .A3(n460), .A2(n463), .A4(n462), .S0(n288), 
        .S1(n295), .Y(n458) );
  AND2X1_HVT U131 ( .A1(n247), .A2(n222), .Y(n457) );
  MUX41X1_HVT U132 ( .A1(n320), .A3(n457), .A2(n369), .A4(n329), .S0(n287), 
        .S1(n280), .Y(n456) );
  MUX41X1_HVT U133 ( .A1(n370), .A3(n322), .A2(n531), .A4(n255), .S0(n237), 
        .S1(n285), .Y(n455) );
  MUX41X1_HVT U136 ( .A1(n536), .A3(n487), .A2(n453), .A4(n327), .S0(n285), 
        .S1(n308), .Y(n452) );
  MUX41X1_HVT U137 ( .A1(n578), .A3(n556), .A2(n560), .A4(n363), .S0(n288), 
        .S1(n283), .Y(n451) );
  MUX41X1_HVT U140 ( .A1(n346), .A3(n274), .A2(n339), .A4(n574), .S0(n287), 
        .S1(n281), .Y(n449) );
  NAND2X0_HVT U141 ( .A1(n266), .A2(n222), .Y(n448) );
  MUX41X1_HVT U142 ( .A1(n448), .A3(n546), .A2(n368), .A4(n339), .S0(n286), 
        .S1(n236), .Y(n447) );
  MUX41X1_HVT U145 ( .A1(n554), .A3(n366), .A2(n445), .A4(n505), .S0(n286), 
        .S1(n309), .Y(n444) );
  MUX41X1_HVT U146 ( .A1(n444), .A3(n446), .A2(n447), .A4(n449), .S0(n202), 
        .S1(n238), .Y(n443) );
  AO21X1_HVT U148 ( .A1(n288), .A2(n324), .A3(n248), .Y(n441) );
  MUX41X1_HVT U151 ( .A1(n360), .A3(n349), .A2(n336), .A4(n439), .S0(n309), 
        .S1(n281), .Y(n438) );
  MUX41X1_HVT U155 ( .A1(n339), .A3(n574), .A2(n566), .A4(n341), .S0(n285), 
        .S1(n237), .Y(n434) );
  MUX41X1_HVT U156 ( .A1(n434), .A3(n438), .A2(n435), .A4(n440), .S0(n297), 
        .S1(n295), .Y(n433) );
  NAND2X0_HVT U159 ( .A1(n430), .A2(n429), .Y(n431) );
  MUX41X1_HVT U162 ( .A1(n270), .A3(n334), .A2(n550), .A4(n427), .S0(n285), 
        .S1(n236), .Y(n426) );
  NAND2X0_HVT U163 ( .A1(n234), .A2(n240), .Y(n425) );
  MUX41X1_HVT U164 ( .A1(n577), .A3(n425), .A2(n548), .A4(n335), .S0(n282), 
        .S1(n308), .Y(n424) );
  NAND2X0_HVT U166 ( .A1(n421), .A2(n575), .Y(n422) );
  MUX41X1_HVT U172 ( .A1(n498), .A3(n416), .A2(n272), .A4(n563), .S0(n285), 
        .S1(n311), .Y(n415) );
  MUX41X1_HVT U174 ( .A1(n362), .A3(n531), .A2(n370), .A4(n263), .S0(n285), 
        .S1(n236), .Y(n413) );
  MUX41X1_HVT U175 ( .A1(n413), .A3(n414), .A2(n415), .A4(n417), .S0(n202), 
        .S1(n238), .Y(n412) );
  NAND2X0_HVT U177 ( .A1(n305), .A2(n244), .Y(n411) );
  MUX41X1_HVT U178 ( .A1(n277), .A3(n411), .A2(n252), .A4(n541), .S0(n285), 
        .S1(n308), .Y(n410) );
  MUX41X1_HVT U182 ( .A1(n322), .A3(n582), .A2(n319), .A4(n360), .S0(n282), 
        .S1(n237), .Y(n406) );
  AND2X1_HVT U185 ( .A1(n263), .A2(n223), .Y(n403) );
  MUX41X1_HVT U190 ( .A1(n400), .A3(n401), .A2(n399), .A4(n402), .S0(n202), 
        .S1(n280), .Y(n398) );
  NAND2X0_HVT U191 ( .A1(n313), .A2(n328), .Y(n397) );
  AND2X1_HVT U192 ( .A1(n347), .A2(n395), .Y(n396) );
  NAND2X0_HVT U194 ( .A1(n543), .A2(n395), .Y(n393) );
  MUX41X1_HVT U195 ( .A1(n394), .A3(n393), .A2(n396), .A4(n397), .S0(n283), 
        .S1(n294), .Y(n392) );
  NAND2X0_HVT U198 ( .A1(n301), .A2(n263), .Y(n575) );
  NAND2X0_HVT U200 ( .A1(n243), .A2(n223), .Y(n461) );
  NAND2X0_HVT U207 ( .A1(n222), .A2(n252), .Y(n525) );
  IBUFFX2_HVT U1 ( .A(n306), .Y(n235) );
  INVX0_HVT U2 ( .A(n288), .Y(n198) );
  MUX21X2_HVT U3 ( .A1(n537), .A2(n276), .S0(n198), .Y(n401) );
  INVX2_HVT U4 ( .A(in[0]), .Y(n306) );
  AO21X2_HVT U14 ( .A1(n265), .A2(n582), .A3(n313), .Y(n421) );
  IBUFFX2_HVT U16 ( .A(in[4]), .Y(n313) );
  IBUFFX2_HVT U17 ( .A(n312), .Y(n311) );
  IBUFFX2_HVT U18 ( .A(n312), .Y(n309) );
  NOR2X0_HVT U20 ( .A1(n376), .A2(n6), .Y(n1) );
  IBUFFX16_HVT U21 ( .A(n290), .Y(n6) );
  IBUFFX2_HVT U22 ( .A(n376), .Y(n247) );
  MUX41X1_HVT U23 ( .A1(n484), .A3(n366), .A2(n505), .A4(n571), .S0(n196), 
        .S1(n197), .Y(n483) );
  IBUFFX16_HVT U24 ( .A(n237), .Y(n196) );
  IBUFFX16_HVT U25 ( .A(n284), .Y(n197) );
  AO21X2_HVT U26 ( .A1(n351), .A2(n287), .A3(n561), .Y(n476) );
  MUX21X2_HVT U27 ( .A1(n247), .A2(n374), .S0(n302), .Y(n544) );
  MUX21X2_HVT U28 ( .A1(n323), .A2(n544), .S0(n288), .Y(n477) );
  INVX1_HVT U29 ( .A(n387), .Y(n359) );
  INVX2_HVT U30 ( .A(n221), .Y(n303) );
  XNOR2X1_HVT U31 ( .A1(n1), .A2(n235), .Y(n537) );
  INVX1_HVT U33 ( .A(n1), .Y(n243) );
  INVX1_HVT U34 ( .A(n323), .Y(n199) );
  INVX1_HVT U36 ( .A(n579), .Y(n323) );
  NAND2X2_HVT U37 ( .A1(in[3]), .A2(in[6]), .Y(n583) );
  MUX41X1_HVT U39 ( .A1(n325), .A3(n373), .A2(n574), .A4(n269), .S0(n313), 
        .S1(n233), .Y(n515) );
  IBUFFX32_HVT U40 ( .A(n321), .Y(n269) );
  MUX41X1_HVT U41 ( .A1(n506), .A3(n502), .A2(n507), .A4(n503), .S0(n200), 
        .S1(n201), .Y(n501) );
  IBUFFX16_HVT U43 ( .A(n297), .Y(n200) );
  IBUFFX16_HVT U44 ( .A(n293), .Y(n201) );
  MUX21X2_HVT U45 ( .A1(n410), .A2(n408), .S0(n293), .Y(n407) );
  MUX21X2_HVT U46 ( .A1(n534), .A2(n533), .S0(n281), .Y(n532) );
  MUX21X1_HVT U47 ( .A1(n527), .A2(n526), .S0(n281), .Y(n524) );
  MUX41X1_HVT U48 ( .A1(n454), .A3(n450), .A2(n464), .A4(n458), .S0(n296), 
        .S1(in[7]), .Y(out[4]) );
  NBUFFX2_HVT U49 ( .A(n294), .Y(n202) );
  NAND2X0_HVT U50 ( .A1(n369), .A2(n218), .Y(n219) );
  NAND2X0_HVT U51 ( .A1(n320), .A2(n310), .Y(n220) );
  NAND2X0_HVT U52 ( .A1(n219), .A2(n220), .Y(n442) );
  IBUFFX2_HVT U54 ( .A(n310), .Y(n218) );
  MUX21X1_HVT U57 ( .A1(n441), .A2(n442), .S0(n233), .Y(n440) );
  IBUFFX2_HVT U58 ( .A(n582), .Y(n319) );
  NBUFFX2_HVT U59 ( .A(n306), .Y(n221) );
  NBUFFX2_HVT U61 ( .A(n306), .Y(n222) );
  NBUFFX2_HVT U63 ( .A(n306), .Y(n223) );
  INVX0_HVT U64 ( .A(in[4]), .Y(n312) );
  NAND2X0_HVT U70 ( .A1(n485), .A2(n257), .Y(n231) );
  INVX0_HVT U71 ( .A(n306), .Y(n304) );
  MUX21X1_HVT U74 ( .A1(n254), .A2(n242), .S0(n271), .Y(n270) );
  OA21X1_HVT U75 ( .A1(n317), .A2(n312), .A3(n326), .Y(n436) );
  INVX0_HVT U76 ( .A(n306), .Y(n234) );
  MUX21X1_HVT U77 ( .A1(n583), .A2(n496), .S0(n271), .Y(n495) );
  NAND2X0_HVT U78 ( .A1(n301), .A2(n300), .Y(n582) );
  INVX1_HVT U79 ( .A(n306), .Y(n301) );
  MUX21X1_HVT U80 ( .A1(n359), .A2(n403), .S0(n218), .Y(n402) );
  INVX1_HVT U84 ( .A(n284), .Y(n233) );
  INVX1_HVT U85 ( .A(n284), .Y(n224) );
  INVX1_HVT U86 ( .A(in[1]), .Y(n293) );
  INVX1_HVT U88 ( .A(n293), .Y(n294) );
  INVX1_HVT U91 ( .A(n293), .Y(n295) );
  INVX1_HVT U92 ( .A(in[5]), .Y(n296) );
  INVX0_HVT U93 ( .A(n252), .Y(n253) );
  INVX1_HVT U94 ( .A(n254), .Y(n373) );
  INVX0_HVT U97 ( .A(in[7]), .Y(n257) );
  INVX0_HVT U103 ( .A(n310), .Y(n258) );
  INVX0_HVT U105 ( .A(n312), .Y(n310) );
  INVX1_HVT U106 ( .A(n378), .Y(n369) );
  INVX0_HVT U107 ( .A(n581), .Y(n320) );
  INVX1_HVT U108 ( .A(n306), .Y(n302) );
  MUX21X1_HVT U109 ( .A1(n336), .A2(n582), .S0(n285), .Y(n522) );
  MUX41X1_HVT U110 ( .A1(n562), .A3(n565), .A2(n250), .A4(n240), .S0(n224), 
        .S1(n218), .Y(n446) );
  IBUFFX2_HVT U111 ( .A(n250), .Y(n542) );
  OA21X1_HVT U112 ( .A1(n318), .A2(n312), .A3(n564), .Y(n510) );
  INVX0_HVT U113 ( .A(n564), .Y(n335) );
  MUX41X1_HVT U117 ( .A1(n560), .A3(n361), .A2(n343), .A4(n276), .S0(n224), 
        .S1(n313), .Y(n502) );
  IBUFFX2_HVT U121 ( .A(n312), .Y(n236) );
  NAND2X0_HVT U123 ( .A1(n431), .A2(n224), .Y(n225) );
  NAND2X0_HVT U125 ( .A1(n432), .A2(n286), .Y(n226) );
  NAND2X0_HVT U126 ( .A1(n225), .A2(n226), .Y(n428) );
  NAND2X0_HVT U128 ( .A1(n412), .A2(n257), .Y(n227) );
  NAND2X0_HVT U134 ( .A1(n419), .A2(in[7]), .Y(n228) );
  NAND2X0_HVT U135 ( .A1(n227), .A2(n228), .Y(out[6]) );
  MUX41X1_HVT U138 ( .A1(n407), .A3(n404), .A2(n398), .A4(n392), .S0(n296), 
        .S1(n257), .Y(out[7]) );
  OA21X2_HVT U139 ( .A1(n343), .A2(n313), .A3(n525), .Y(n399) );
  AO21X2_HVT U143 ( .A1(n305), .A2(n248), .A3(n312), .Y(n395) );
  NAND2X0_HVT U144 ( .A1(n494), .A2(n224), .Y(n229) );
  NAND2X0_HVT U147 ( .A1(n495), .A2(n281), .Y(n230) );
  NAND2X0_HVT U149 ( .A1(n229), .A2(n230), .Y(n493) );
  NAND2X0_HVT U150 ( .A1(n492), .A2(in[7]), .Y(n232) );
  NAND2X0_HVT U152 ( .A1(n231), .A2(n232), .Y(out[2]) );
  MUX21X1_HVT U153 ( .A1(n251), .A2(n256), .S0(n287), .Y(n496) );
  MUX41X1_HVT U154 ( .A1(n335), .A3(n346), .A2(n347), .A4(n576), .S0(n233), 
        .S1(n313), .Y(n512) );
  MUX41X1_HVT U157 ( .A1(n512), .A3(n515), .A2(n509), .A4(n513), .S0(n297), 
        .S1(n293), .Y(n508) );
  AO21X2_HVT U158 ( .A1(n223), .A2(n268), .A3(n313), .Y(n429) );
  MUX21X2_HVT U160 ( .A1(n476), .A2(n477), .S0(n286), .Y(n475) );
  MUX41X1_HVT U161 ( .A1(n335), .A3(n340), .A2(n265), .A4(n584), .S0(n309), 
        .S1(n284), .Y(n480) );
  MUX41X1_HVT U165 ( .A1(n479), .A3(n480), .A2(n481), .A4(n483), .S0(in[1]), 
        .S1(n238), .Y(n478) );
  MUX21X2_HVT U167 ( .A1(n465), .A2(n467), .S0(n294), .Y(n464) );
  MUX41X1_HVT U168 ( .A1(n272), .A3(n418), .A2(n277), .A4(n275), .S0(n309), 
        .S1(n224), .Y(n417) );
  IBUFFX2_HVT U169 ( .A(n312), .Y(n308) );
  MUX41X1_HVT U170 ( .A1(n568), .A3(n345), .A2(n567), .A4(n343), .S0(n233), 
        .S1(n313), .Y(n507) );
  MUX21X1_HVT U171 ( .A1(n542), .A2(n358), .S0(n287), .Y(n432) );
  MUX21X1_HVT U173 ( .A1(n371), .A2(n264), .S0(n221), .Y(n563) );
  MUX21X1_HVT U176 ( .A1(n373), .A2(n374), .S0(n301), .Y(n418) );
  MUX21X1_HVT U179 ( .A1(n544), .A2(n357), .S0(n258), .Y(n400) );
  INVX0_HVT U180 ( .A(n270), .Y(n541) );
  INVX0_HVT U181 ( .A(n539), .Y(n353) );
  NBUFFX2_HVT U183 ( .A(n376), .Y(n291) );
  INVX1_HVT U184 ( .A(n291), .Y(n279) );
  INVX1_HVT U186 ( .A(n386), .Y(n360) );
  INVX0_HVT U187 ( .A(n372), .Y(n267) );
  INVX0_HVT U188 ( .A(n305), .Y(n271) );
  INVX1_HVT U189 ( .A(n258), .Y(n237) );
  MUX41X1_HVT U193 ( .A1(n364), .A3(n361), .A2(n316), .A4(n353), .S0(n237), 
        .S1(n283), .Y(n479) );
  MUX21X2_HVT U196 ( .A1(n478), .A2(n468), .S0(n257), .Y(out[3]) );
  MUX41X1_HVT U197 ( .A1(n581), .A3(n577), .A2(n355), .A4(n359), .S0(n224), 
        .S1(n313), .Y(n506) );
  INVX1_HVT U199 ( .A(n296), .Y(n238) );
  MUX41X1_HVT U201 ( .A1(n365), .A3(n482), .A2(n583), .A4(n322), .S0(n236), 
        .S1(n283), .Y(n481) );
  INVX1_HVT U202 ( .A(n381), .Y(n365) );
  INVX0_HVT U203 ( .A(n1), .Y(n239) );
  INVX1_HVT U204 ( .A(n239), .Y(n240) );
  INVX1_HVT U205 ( .A(n239), .Y(n241) );
  INVX1_HVT U206 ( .A(n1), .Y(n242) );
  INVX0_HVT U208 ( .A(n290), .Y(n244) );
  NAND2X0_HVT U209 ( .A1(n406), .A2(n294), .Y(n245) );
  NAND2X0_HVT U210 ( .A1(n405), .A2(n293), .Y(n246) );
  NAND2X0_HVT U211 ( .A1(n245), .A2(n246), .Y(n404) );
  INVX0_HVT U212 ( .A(in[3]), .Y(n372) );
  INVX1_HVT U213 ( .A(n391), .Y(n355) );
  INVX1_HVT U214 ( .A(in[6]), .Y(n376) );
  MUX21X1_HVT U215 ( .A1(n371), .A2(n244), .S0(n304), .Y(n562) );
  IBUFFX2_HVT U216 ( .A(n568), .Y(n331) );
  INVX1_HVT U217 ( .A(n375), .Y(n261) );
  MUX41X1_HVT U218 ( .A1(n335), .A3(n543), .A2(n250), .A4(n355), .S0(n311), 
        .S1(n233), .Y(n405) );
  INVX1_HVT U219 ( .A(n299), .Y(n248) );
  INVX0_HVT U220 ( .A(n563), .Y(n336) );
  MUX41X1_HVT U221 ( .A1(n539), .A3(n555), .A2(n316), .A4(n331), .S0(n224), 
        .S1(n218), .Y(n499) );
  MUX21X1_HVT U222 ( .A1(n256), .A2(n371), .S0(n223), .Y(n389) );
  MUX21X1_HVT U223 ( .A1(n256), .A2(n264), .S0(n302), .Y(n549) );
  INVX0_HVT U224 ( .A(n252), .Y(n249) );
  MUX41X1_HVT U225 ( .A1(n549), .A3(n299), .A2(n252), .A4(n268), .S0(n233), 
        .S1(n258), .Y(n414) );
  INVX1_HVT U226 ( .A(n261), .Y(n262) );
  IBUFFX2_HVT U227 ( .A(n549), .Y(n348) );
  INVX1_HVT U228 ( .A(n254), .Y(n252) );
  MUX21X1_HVT U229 ( .A1(n298), .A2(n267), .S0(n221), .Y(n250) );
  OR2X1_HVT U230 ( .A1(n372), .A2(n279), .Y(n254) );
  XNOR2X1_HVT U231 ( .A1(n279), .A2(n267), .Y(n251) );
  INVX0_HVT U232 ( .A(n264), .Y(n265) );
  INVX0_HVT U233 ( .A(n569), .Y(n264) );
  INVX1_HVT U234 ( .A(n569), .Y(n375) );
  MUX21X1_HVT U235 ( .A1(n289), .A2(n251), .S0(n221), .Y(n564) );
  INVX0_HVT U236 ( .A(n269), .Y(n255) );
  XNOR2X2_HVT U237 ( .A1(n279), .A2(n267), .Y(n569) );
  NOR2X1_HVT U238 ( .A1(n321), .A2(n240), .Y(n409) );
  MUX21X2_HVT U239 ( .A1(n508), .A2(n501), .S0(n257), .Y(out[1]) );
  INVX1_HVT U240 ( .A(n299), .Y(n371) );
  INVX1_HVT U241 ( .A(n545), .Y(n351) );
  NBUFFX2_HVT U242 ( .A(n291), .Y(n256) );
  MUX41X1_HVT U243 ( .A1(n420), .A3(n426), .A2(n424), .A4(n428), .S0(n297), 
        .S1(n295), .Y(n419) );
  MUX21X2_HVT U244 ( .A1(n422), .A2(n423), .S0(n307), .Y(n420) );
  MUX21X2_HVT U245 ( .A1(n335), .A2(n522), .S0(n278), .Y(n521) );
  MUX21X2_HVT U246 ( .A1(n516), .A2(n523), .S0(in[7]), .Y(out[0]) );
  MUX21X2_HVT U247 ( .A1(n443), .A2(n433), .S0(n257), .Y(out[5]) );
  MUX21X1_HVT U248 ( .A1(n569), .A2(n256), .S0(n305), .Y(n560) );
  INVX1_HVT U249 ( .A(n389), .Y(n357) );
  NAND2X0_HVT U250 ( .A1(n559), .A2(n258), .Y(n259) );
  NAND2X0_HVT U251 ( .A1(n562), .A2(n311), .Y(n260) );
  NAND2X0_HVT U252 ( .A1(n260), .A2(n259), .Y(n423) );
  INVX1_HVT U253 ( .A(n251), .Y(n263) );
  INVX0_HVT U254 ( .A(n264), .Y(n266) );
  INVX1_HVT U255 ( .A(n252), .Y(n268) );
  MUX41X1_HVT U256 ( .A1(n409), .A3(n540), .A2(n553), .A4(n314), .S0(n285), 
        .S1(n313), .Y(n408) );
  AND2X1_HVT U257 ( .A1(n269), .A2(n300), .Y(n272) );
  NBUFFX2_HVT U258 ( .A(n584), .Y(n299) );
  NBUFFX2_HVT U259 ( .A(n584), .Y(n300) );
  AND2X1_HVT U260 ( .A1(n300), .A2(n570), .Y(n273) );
  MUX21X1_HVT U261 ( .A1(n352), .A2(n275), .S0(n236), .Y(n394) );
  MUX21X1_HVT U262 ( .A1(n263), .A2(n290), .S0(n235), .Y(n546) );
  MUX21X1_HVT U263 ( .A1(n373), .A2(n241), .S0(n305), .Y(n557) );
  MUX21X1_HVT U264 ( .A1(n248), .A2(n262), .S0(n302), .Y(n552) );
  MUX21X1_HVT U265 ( .A1(n265), .A2(n373), .S0(n235), .Y(n554) );
  MUX21X1_HVT U266 ( .A1(n256), .A2(n371), .S0(n303), .Y(n559) );
  MUX21X1_HVT U267 ( .A1(n337), .A2(n531), .S0(n287), .Y(n527) );
  MUX21X1_HVT U268 ( .A1(n242), .A2(n298), .S0(n234), .Y(n427) );
  MUX21X1_HVT U269 ( .A1(n256), .A2(n241), .S0(n235), .Y(n439) );
  MUX21X1_HVT U270 ( .A1(n373), .A2(n292), .S0(n301), .Y(n416) );
  XOR2X1_HVT U271 ( .A1(n253), .A2(n301), .Y(n548) );
  NAND2X0_HVT U272 ( .A1(n372), .A2(n376), .Y(n584) );
  MUX21X1_HVT U273 ( .A1(n373), .A2(n266), .S0(n301), .Y(n384) );
  MUX21X1_HVT U274 ( .A1(n262), .A2(n292), .S0(n302), .Y(n379) );
  MUX21X1_HVT U275 ( .A1(n290), .A2(n248), .S0(n235), .Y(n555) );
  MUX21X1_HVT U276 ( .A1(n325), .A2(n266), .S0(n288), .Y(n494) );
  MUX21X1_HVT U277 ( .A1(n292), .A2(n584), .S0(n234), .Y(n482) );
  MUX21X1_HVT U278 ( .A1(n242), .A2(n584), .S0(n303), .Y(n378) );
  MUX21X1_HVT U279 ( .A1(n292), .A2(n251), .S0(n301), .Y(n545) );
  XNOR2X1_HVT U280 ( .A1(n299), .A2(n304), .Y(n274) );
  MUX21X1_HVT U281 ( .A1(n298), .A2(n300), .S0(n302), .Y(n567) );
  MUX21X1_HVT U282 ( .A1(n552), .A2(n273), .S0(n286), .Y(n460) );
  MUX21X1_HVT U283 ( .A1(n368), .A2(n274), .S0(n281), .Y(n463) );
  MUX21X1_HVT U284 ( .A1(n261), .A2(n241), .S0(n301), .Y(n551) );
  XOR2X1_HVT U285 ( .A1(n583), .A2(n302), .Y(n538) );
  XOR2X1_HVT U286 ( .A1(n261), .A2(n234), .Y(n539) );
  MUX21X1_HVT U287 ( .A1(n374), .A2(n289), .S0(n305), .Y(n388) );
  MUX21X1_HVT U288 ( .A1(n289), .A2(n300), .S0(n303), .Y(n387) );
  MUX21X1_HVT U289 ( .A1(n249), .A2(n584), .S0(n235), .Y(n571) );
  MUX21X1_HVT U290 ( .A1(n583), .A2(n290), .S0(n304), .Y(n566) );
  MUX21X1_HVT U291 ( .A1(n290), .A2(n292), .S0(n305), .Y(n540) );
  MUX21X1_HVT U292 ( .A1(n289), .A2(n583), .S0(n304), .Y(n381) );
  AND2X1_HVT U293 ( .A1(n303), .A2(n256), .Y(n275) );
  MUX21X1_HVT U294 ( .A1(n298), .A2(n292), .S0(n303), .Y(n466) );
  NBUFFX2_HVT U295 ( .A(n310), .Y(n288) );
  NBUFFX2_HVT U296 ( .A(n310), .Y(n287) );
  NBUFFX2_HVT U297 ( .A(n376), .Y(n292) );
  MUX21X1_HVT U298 ( .A1(n436), .A2(n437), .S0(n286), .Y(n435) );
  MUX21X1_HVT U299 ( .A1(n560), .A2(n276), .S0(n287), .Y(n437) );
  MUX21X1_HVT U300 ( .A1(n584), .A2(n242), .S0(n304), .Y(n445) );
  MUX21X1_HVT U301 ( .A1(n341), .A2(n330), .S0(n288), .Y(n534) );
  MUX21X1_HVT U302 ( .A1(n371), .A2(n374), .S0(n305), .Y(n535) );
  MUX21X1_HVT U303 ( .A1(n338), .A2(n529), .S0(n278), .Y(n528) );
  MUX21X1_HVT U304 ( .A1(n339), .A2(n581), .S0(n286), .Y(n529) );
  MUX21X1_HVT U305 ( .A1(n511), .A2(n510), .S0(n286), .Y(n509) );
  MUX21X1_HVT U306 ( .A1(n358), .A2(n315), .S0(n288), .Y(n511) );
  AND2X1_HVT U307 ( .A1(n298), .A2(n222), .Y(n276) );
  AND2X1_HVT U308 ( .A1(n374), .A2(n222), .Y(n277) );
  NBUFFX2_HVT U309 ( .A(n583), .Y(n298) );
  NBUFFX2_HVT U310 ( .A(n372), .Y(n290) );
  NBUFFX2_HVT U311 ( .A(n372), .Y(n289) );
  NBUFFX2_HVT U312 ( .A(n307), .Y(n285) );
  XNOR2X1_HVT U313 ( .A1(n312), .A2(n282), .Y(n278) );
  NBUFFX2_HVT U314 ( .A(n280), .Y(n286) );
  INVX1_HVT U315 ( .A(n306), .Y(n305) );
  NBUFFX2_HVT U316 ( .A(n307), .Y(n282) );
  NBUFFX2_HVT U317 ( .A(n307), .Y(n284) );
  NBUFFX2_HVT U318 ( .A(n280), .Y(n283) );
  NBUFFX2_HVT U319 ( .A(n307), .Y(n280) );
  NBUFFX2_HVT U320 ( .A(n307), .Y(n281) );
  INVX1_HVT U321 ( .A(n296), .Y(n297) );
  MUX21X1_HVT U322 ( .A1(n247), .A2(n253), .S0(n234), .Y(n568) );
  MUX21X1_HVT U323 ( .A1(n247), .A2(n373), .S0(n304), .Y(n561) );
  MUX21X1_HVT U324 ( .A1(n243), .A2(n244), .S0(n234), .Y(n490) );
  MUX21X1_HVT U325 ( .A1(n373), .A2(n244), .S0(n235), .Y(n377) );
  MUX21X1_HVT U326 ( .A1(n268), .A2(n244), .S0(n303), .Y(n430) );
  MUX21X1_HVT U327 ( .A1(n374), .A2(n240), .S0(n302), .Y(n471) );
  MUX21X1_HVT U328 ( .A1(n451), .A2(n452), .S0(n294), .Y(n450) );
  MUX21X1_HVT U329 ( .A1(n244), .A2(n268), .S0(n305), .Y(n383) );
  MUX21X1_HVT U330 ( .A1(n455), .A2(n456), .S0(n295), .Y(n454) );
  XOR2X1_HVT U331 ( .A1(n302), .A2(n247), .Y(n536) );
  MUX21X1_HVT U332 ( .A1(n248), .A2(n247), .S0(n234), .Y(n453) );
  MUX21X1_HVT U333 ( .A1(n247), .A2(n240), .S0(n235), .Y(n391) );
  MUX21X1_HVT U334 ( .A1(n243), .A2(n247), .S0(n301), .Y(n556) );
  MUX21X1_HVT U335 ( .A1(n292), .A2(n244), .S0(n304), .Y(n558) );
  MUX21X1_HVT U336 ( .A1(n583), .A2(n247), .S0(n302), .Y(n385) );
  MUX21X1_HVT U337 ( .A1(n244), .A2(n242), .S0(n303), .Y(n382) );
  MUX21X1_HVT U338 ( .A1(n247), .A2(n298), .S0(n303), .Y(n390) );
  MUX21X1_HVT U339 ( .A1(n289), .A2(n247), .S0(n303), .Y(n380) );
  NBUFFX2_HVT U340 ( .A(in[2]), .Y(n307) );
  MUX21X1_HVT U341 ( .A1(n289), .A2(n375), .S0(n304), .Y(n386) );
  INVX0_HVT U342 ( .A(n574), .Y(n314) );
  INVX0_HVT U343 ( .A(n553), .Y(n315) );
  INVX0_HVT U344 ( .A(n547), .Y(n316) );
  INVX0_HVT U345 ( .A(n487), .Y(n317) );
  INVX0_HVT U346 ( .A(n448), .Y(n318) );
  INVX0_HVT U347 ( .A(n580), .Y(n321) );
  INVX0_HVT U348 ( .A(n543), .Y(n322) );
  INVX0_HVT U349 ( .A(n578), .Y(n324) );
  INVX0_HVT U350 ( .A(n550), .Y(n325) );
  INVX0_HVT U351 ( .A(n572), .Y(n326) );
  INVX0_HVT U352 ( .A(n577), .Y(n327) );
  INVX0_HVT U353 ( .A(n573), .Y(n328) );
  INVX0_HVT U354 ( .A(n571), .Y(n329) );
  INVX0_HVT U355 ( .A(n570), .Y(n330) );
  INVX0_HVT U356 ( .A(n567), .Y(n332) );
  INVX0_HVT U357 ( .A(n566), .Y(n333) );
  INVX0_HVT U358 ( .A(n565), .Y(n334) );
  INVX0_HVT U359 ( .A(n562), .Y(n337) );
  INVX0_HVT U360 ( .A(n561), .Y(n338) );
  INVX0_HVT U361 ( .A(n560), .Y(n339) );
  INVX0_HVT U362 ( .A(n559), .Y(n340) );
  INVX0_HVT U363 ( .A(n558), .Y(n341) );
  INVX0_HVT U364 ( .A(n557), .Y(n342) );
  INVX0_HVT U365 ( .A(n556), .Y(n343) );
  INVX0_HVT U366 ( .A(n555), .Y(n344) );
  INVX0_HVT U367 ( .A(n554), .Y(n345) );
  INVX0_HVT U368 ( .A(n552), .Y(n346) );
  INVX0_HVT U369 ( .A(n551), .Y(n347) );
  INVX0_HVT U370 ( .A(n548), .Y(n349) );
  INVX0_HVT U371 ( .A(n546), .Y(n350) );
  INVX0_HVT U372 ( .A(n540), .Y(n352) );
  INVX0_HVT U373 ( .A(n576), .Y(n354) );
  INVX0_HVT U374 ( .A(n390), .Y(n356) );
  INVX0_HVT U375 ( .A(n388), .Y(n358) );
  INVX0_HVT U376 ( .A(n385), .Y(n361) );
  INVX0_HVT U377 ( .A(n384), .Y(n362) );
  INVX0_HVT U378 ( .A(n383), .Y(n363) );
  INVX0_HVT U379 ( .A(n382), .Y(n364) );
  INVX0_HVT U380 ( .A(n380), .Y(n366) );
  INVX0_HVT U381 ( .A(n430), .Y(n367) );
  INVX0_HVT U382 ( .A(n379), .Y(n368) );
  INVX0_HVT U383 ( .A(n377), .Y(n370) );
  INVX0_HVT U384 ( .A(n583), .Y(n374) );
endmodule

