
module inv_sbox_12 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n196, n197, n198, n199, n200, n201, n202, n205, n208, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626;

  NAND2X0_HVT U1 ( .A1(in[3]), .A2(n333), .Y(n626) );
  NAND2X0_HVT U3 ( .A1(n304), .A2(n309), .Y(n624) );
  NAND2X0_HVT U5 ( .A1(n623), .A2(n343), .Y(n622) );
  NAND2X0_HVT U8 ( .A1(n245), .A2(n343), .Y(n618) );
  NAND2X0_HVT U9 ( .A1(n350), .A2(n618), .Y(n617) );
  NAND2X0_HVT U10 ( .A1(n350), .A2(n615), .Y(n616) );
  NAND2X0_HVT U11 ( .A1(n235), .A2(n349), .Y(n614) );
  NAND2X0_HVT U12 ( .A1(n275), .A2(n415), .Y(n613) );
  NAND2X0_HVT U13 ( .A1(n346), .A2(n618), .Y(n612) );
  NAND2X0_HVT U15 ( .A1(n339), .A2(n352), .Y(n610) );
  NAND2X0_HVT U19 ( .A1(n237), .A2(n417), .Y(n605) );
  NAND2X0_HVT U25 ( .A1(n309), .A2(n331), .Y(n621) );
  NAND2X0_HVT U32 ( .A1(n333), .A2(n235), .Y(n593) );
  NAND2X0_HVT U35 ( .A1(n618), .A2(n418), .Y(n590) );
  NAND2X0_HVT U38 ( .A1(n330), .A2(n235), .Y(n587) );
  NAND2X0_HVT U42 ( .A1(n620), .A2(n418), .Y(n583) );
  OA21X1_HVT U53 ( .A1(n270), .A2(n575), .A3(n221), .Y(n573) );
  NAND2X0_HVT U55 ( .A1(n345), .A2(n623), .Y(n571) );
  AO21X1_HVT U60 ( .A1(n565), .A2(n327), .A3(n604), .Y(n566) );
  NAND2X0_HVT U66 ( .A1(n237), .A2(n309), .Y(n559) );
  MUX41X1_HVT U67 ( .A1(n377), .A3(n400), .A2(n379), .A4(n559), .S0(n328), 
        .S1(n320), .Y(n558) );
  MUX41X1_HVT U71 ( .A1(n277), .A3(n416), .A2(n614), .A4(n373), .S0(n322), 
        .S1(n360), .Y(n555) );
  NAND2X0_HVT U72 ( .A1(n341), .A2(n619), .Y(n554) );
  MUX41X1_HVT U73 ( .A1(n598), .A3(n554), .A2(n308), .A4(n330), .S0(n328), 
        .S1(n319), .Y(n553) );
  MUX41X1_HVT U74 ( .A1(n616), .A3(n391), .A2(n390), .A4(n383), .S0(n323), 
        .S1(n360), .Y(n552) );
  MUX41X1_HVT U80 ( .A1(n402), .A3(n399), .A2(n617), .A4(n622), .S0(n322), 
        .S1(n360), .Y(n546) );
  NAND2X0_HVT U81 ( .A1(n349), .A2(n619), .Y(n545) );
  AND2X1_HVT U82 ( .A1(n277), .A2(n345), .Y(n544) );
  MUX41X1_HVT U83 ( .A1(n544), .A3(n388), .A2(n305), .A4(n545), .S0(n322), 
        .S1(n360), .Y(n543) );
  MUX41X1_HVT U84 ( .A1(n315), .A3(n387), .A2(n403), .A4(n600), .S0(n323), 
        .S1(n360), .Y(n542) );
  MUX41X1_HVT U85 ( .A1(n542), .A3(n546), .A2(n543), .A4(n547), .S0(n338), 
        .S1(n335), .Y(n541) );
  MUX41X1_HVT U88 ( .A1(n379), .A3(n364), .A2(n595), .A4(n579), .S0(n322), 
        .S1(n359), .Y(n539) );
  NAND2X0_HVT U89 ( .A1(n235), .A2(n414), .Y(n538) );
  MUX41X1_HVT U90 ( .A1(n416), .A3(n619), .A2(n578), .A4(n538), .S0(n322), 
        .S1(n360), .Y(n537) );
  MUX41X1_HVT U95 ( .A1(n533), .A3(n539), .A2(n537), .A4(n540), .S0(n338), 
        .S1(n335), .Y(n532) );
  MUX41X1_HVT U96 ( .A1(n400), .A3(n612), .A2(n386), .A4(n405), .S0(n323), 
        .S1(n359), .Y(n531) );
  MUX41X1_HVT U98 ( .A1(n530), .A3(n406), .A2(n392), .A4(n597), .S0(n323), 
        .S1(n359), .Y(n529) );
  MUX41X1_HVT U99 ( .A1(n593), .A3(n381), .A2(n577), .A4(n341), .S0(n360), 
        .S1(n320), .Y(n528) );
  NAND2X0_HVT U100 ( .A1(n355), .A2(n413), .Y(n527) );
  MUX41X1_HVT U101 ( .A1(n407), .A3(n613), .A2(n246), .A4(n527), .S0(n360), 
        .S1(n318), .Y(n526) );
  AND2X1_HVT U104 ( .A1(n619), .A2(n342), .Y(n524) );
  MUX41X1_HVT U110 ( .A1(n519), .A3(n521), .A2(n520), .A4(n523), .S0(n338), 
        .S1(n300), .Y(n518) );
  AO21X1_HVT U112 ( .A1(n394), .A2(n328), .A3(n601), .Y(n516) );
  NAND2X0_HVT U114 ( .A1(n350), .A2(n619), .Y(n514) );
  MUX41X1_HVT U115 ( .A1(n514), .A3(n614), .A2(n394), .A4(n345), .S0(n360), 
        .S1(n320), .Y(n513) );
  MUX41X1_HVT U116 ( .A1(n393), .A3(n387), .A2(n364), .A4(n610), .S0(n321), 
        .S1(n359), .Y(n512) );
  NAND2X0_HVT U118 ( .A1(n355), .A2(n202), .Y(n510) );
  MUX41X1_HVT U119 ( .A1(n409), .A3(n511), .A2(n588), .A4(n510), .S0(n321), 
        .S1(n359), .Y(n509) );
  MUX41X1_HVT U120 ( .A1(n509), .A3(n513), .A2(n512), .A4(n515), .S0(n338), 
        .S1(n300), .Y(n508) );
  MUX41X1_HVT U122 ( .A1(n398), .A3(n311), .A2(n579), .A4(n401), .S0(n321), 
        .S1(n359), .Y(n507) );
  MUX41X1_HVT U124 ( .A1(n314), .A3(n506), .A2(n602), .A4(n306), .S0(n329), 
        .S1(n321), .Y(n505) );
  AOI21X1_HVT U127 ( .A1(n326), .A2(n501), .A3(n371), .Y(n502) );
  NAND2X0_HVT U129 ( .A1(n325), .A2(n626), .Y(n499) );
  MUX41X1_HVT U130 ( .A1(n499), .A3(n500), .A2(n503), .A4(n502), .S0(n329), 
        .S1(n300), .Y(n498) );
  AND2X1_HVT U131 ( .A1(n309), .A2(n354), .Y(n497) );
  MUX41X1_HVT U132 ( .A1(n368), .A3(n497), .A2(n411), .A4(n377), .S0(n329), 
        .S1(n319), .Y(n496) );
  MUX41X1_HVT U133 ( .A1(n412), .A3(n370), .A2(n262), .A4(n369), .S0(n329), 
        .S1(n318), .Y(n495) );
  MUX41X1_HVT U136 ( .A1(n576), .A3(n527), .A2(n493), .A4(n375), .S0(n325), 
        .S1(n359), .Y(n492) );
  MUX41X1_HVT U137 ( .A1(n618), .A3(n596), .A2(n600), .A4(n405), .S0(n328), 
        .S1(n318), .Y(n491) );
  MUX41X1_HVT U139 ( .A1(n490), .A3(n494), .A2(n498), .A4(n504), .S0(in[5]), 
        .S1(n303), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n390), .A3(n312), .A2(n385), .A4(n614), .S0(n328), 
        .S1(n320), .Y(n489) );
  NAND2X0_HVT U141 ( .A1(n340), .A2(n355), .Y(n488) );
  MUX41X1_HVT U142 ( .A1(n488), .A3(n586), .A2(n410), .A4(n385), .S0(n326), 
        .S1(n359), .Y(n487) );
  MUX41X1_HVT U145 ( .A1(n594), .A3(n408), .A2(n485), .A4(n545), .S0(n326), 
        .S1(n361), .Y(n484) );
  MUX41X1_HVT U151 ( .A1(n305), .A3(n392), .A2(n234), .A4(n479), .S0(n329), 
        .S1(n318), .Y(n478) );
  MUX41X1_HVT U155 ( .A1(n385), .A3(n614), .A2(n606), .A4(n386), .S0(n324), 
        .S1(n361), .Y(n474) );
  NAND2X0_HVT U159 ( .A1(n470), .A2(n469), .Y(n471) );
  MUX41X1_HVT U162 ( .A1(n307), .A3(n382), .A2(n590), .A4(n467), .S0(n324), 
        .S1(n358), .Y(n466) );
  NAND2X0_HVT U163 ( .A1(n351), .A2(n414), .Y(n465) );
  MUX41X1_HVT U164 ( .A1(n617), .A3(n465), .A2(n588), .A4(n383), .S0(n321), 
        .S1(n361), .Y(n464) );
  NAND2X0_HVT U166 ( .A1(n615), .A2(n461), .Y(n462) );
  MUX41X1_HVT U172 ( .A1(n538), .A3(n456), .A2(n313), .A4(n603), .S0(n324), 
        .S1(n361), .Y(n455) );
  MUX41X1_HVT U173 ( .A1(n626), .A3(n416), .A2(n347), .A4(n589), .S0(n324), 
        .S1(n361), .Y(n454) );
  MUX41X1_HVT U175 ( .A1(n453), .A3(n454), .A2(n455), .A4(n457), .S0(n336), 
        .S1(n338), .Y(n452) );
  NAND2X0_HVT U177 ( .A1(n275), .A2(n202), .Y(n451) );
  MUX41X1_HVT U178 ( .A1(n316), .A3(n451), .A2(n416), .A4(n581), .S0(n324), 
        .S1(n361), .Y(n450) );
  AND2X1_HVT U179 ( .A1(n277), .A2(n342), .Y(n449) );
  MUX41X1_HVT U182 ( .A1(n370), .A3(n623), .A2(n367), .A4(n305), .S0(n321), 
        .S1(n358), .Y(n446) );
  AND2X1_HVT U185 ( .A1(n418), .A2(n354), .Y(n443) );
  AND2X1_HVT U192 ( .A1(n391), .A2(n435), .Y(n436) );
  NAND2X0_HVT U194 ( .A1(n435), .A2(n205), .Y(n433) );
  NAND2X0_HVT U198 ( .A1(n351), .A2(n200), .Y(n615) );
  NAND2X0_HVT U200 ( .A1(n343), .A2(n258), .Y(n501) );
  NAND2X0_HVT U207 ( .A1(n258), .A2(n416), .Y(n565) );
  MUX21X2_HVT U2 ( .A1(n396), .A2(n314), .S0(n327), .Y(n434) );
  MUX21X1_HVT U4 ( .A1(n197), .A2(n347), .S0(n218), .Y(n196) );
  IBUFFX16_HVT U6 ( .A(n196), .Y(n599) );
  IBUFFX16_HVT U7 ( .A(n333), .Y(n197) );
  IBUFFX2_HVT U14 ( .A(n300), .Y(n242) );
  IBUFFX2_HVT U16 ( .A(n415), .Y(n304) );
  MUX21X2_HVT U17 ( .A1(n463), .A2(n462), .S0(n230), .Y(n460) );
  XOR2X2_HVT U18 ( .A1(n340), .A2(n276), .Y(n579) );
  INVX2_HVT U20 ( .A(n291), .Y(n362) );
  MUX41X1_HVT U21 ( .A1(n313), .A3(n316), .A2(n458), .A4(n314), .S0(n198), 
        .S1(n361), .Y(n457) );
  IBUFFX16_HVT U22 ( .A(n324), .Y(n198) );
  INVX0_HVT U23 ( .A(n309), .Y(n199) );
  INVX0_HVT U24 ( .A(n340), .Y(n200) );
  INVX0_HVT U26 ( .A(in[6]), .Y(n310) );
  INVX0_HVT U27 ( .A(n339), .Y(n418) );
  INVX1_HVT U28 ( .A(n304), .Y(n201) );
  INVX1_HVT U29 ( .A(n201), .Y(n202) );
  INVX0_HVT U30 ( .A(n370), .Y(n205) );
  MUX21X2_HVT U31 ( .A1(n535), .A2(n534), .S0(n208), .Y(n533) );
  IBUFFX16_HVT U33 ( .A(n325), .Y(n208) );
  MUX41X1_HVT U34 ( .A1(n196), .A3(n404), .A2(n315), .A4(n367), .S0(n236), 
        .S1(n270), .Y(n540) );
  MUX41X1_HVT U36 ( .A1(n434), .A3(n436), .A2(n433), .A4(n437), .S0(n336), 
        .S1(n322), .Y(n432) );
  INVX1_HVT U37 ( .A(n235), .Y(n218) );
  NAND2X1_HVT U39 ( .A1(n299), .A2(n376), .Y(n437) );
  INVX1_HVT U40 ( .A(n278), .Y(n235) );
  IBUFFX2_HVT U41 ( .A(n354), .Y(n352) );
  INVX1_HVT U43 ( .A(n327), .Y(n219) );
  MUX41X1_HVT U44 ( .A1(n442), .A3(n439), .A2(n441), .A4(n440), .S0(n334), 
        .S1(n238), .Y(n438) );
  MUX21X2_HVT U45 ( .A1(n401), .A2(n582), .S0(n219), .Y(n472) );
  INVX0_HVT U46 ( .A(n396), .Y(n220) );
  INVX1_HVT U47 ( .A(n580), .Y(n396) );
  IBUFFX16_HVT U48 ( .A(n362), .Y(n361) );
  XOR2X1_HVT U49 ( .A1(n350), .A2(n237), .Y(n588) );
  MUX21X1_HVT U50 ( .A1(n371), .A2(n584), .S0(n328), .Y(n517) );
  MUX21X1_HVT U51 ( .A1(n373), .A2(n339), .S0(n329), .Y(n534) );
  MUX41X1_HVT U52 ( .A1(n583), .A3(n399), .A2(n383), .A4(n395), .S0(n233), 
        .S1(n232), .Y(n445) );
  IBUFFX2_HVT U54 ( .A(n327), .Y(n232) );
  IBUFFX2_HVT U56 ( .A(n319), .Y(n233) );
  INVX0_HVT U57 ( .A(n582), .Y(n395) );
  MUX21X1_HVT U58 ( .A1(n626), .A2(n222), .S0(n353), .Y(n221) );
  INVX8_HVT U59 ( .A(n221), .Y(n597) );
  IBUFFX16_HVT U61 ( .A(n414), .Y(n222) );
  MUX21X2_HVT U62 ( .A1(n443), .A2(n402), .S0(n327), .Y(n442) );
  NAND2X0_HVT U63 ( .A1(n518), .A2(n223), .Y(n224) );
  NAND2X0_HVT U64 ( .A1(n508), .A2(n253), .Y(n225) );
  NAND2X0_HVT U65 ( .A1(n224), .A2(n225), .Y(out[3]) );
  IBUFFX2_HVT U68 ( .A(n253), .Y(n223) );
  MUX41X1_HVT U69 ( .A1(n363), .A3(n593), .A2(n220), .A4(n449), .S0(n226), 
        .S1(n358), .Y(n448) );
  IBUFFX16_HVT U70 ( .A(n324), .Y(n226) );
  INVX1_HVT U75 ( .A(n327), .Y(n239) );
  NAND2X0_HVT U76 ( .A1(n602), .A2(n227), .Y(n228) );
  NAND2X0_HVT U77 ( .A1(n599), .A2(n239), .Y(n229) );
  NAND2X0_HVT U78 ( .A1(n228), .A2(n229), .Y(n463) );
  INVX0_HVT U79 ( .A(n239), .Y(n227) );
  IBUFFX16_HVT U86 ( .A(n325), .Y(n230) );
  XOR2X2_HVT U87 ( .A1(n231), .A2(n258), .Y(n577) );
  IBUFFX16_HVT U91 ( .A(n342), .Y(n231) );
  INVX0_HVT U92 ( .A(n354), .Y(n353) );
  IBUFFX2_HVT U93 ( .A(n291), .Y(n270) );
  IBUFFX2_HVT U94 ( .A(n290), .Y(n359) );
  MUX21X2_HVT U97 ( .A1(n551), .A2(n550), .S0(n326), .Y(n549) );
  INVX0_HVT U102 ( .A(n285), .Y(n551) );
  IBUFFX2_HVT U103 ( .A(n354), .Y(n237) );
  MUX21X1_HVT U105 ( .A1(n347), .A2(n339), .S0(n258), .Y(n234) );
  INVX8_HVT U106 ( .A(n234), .Y(n603) );
  IBUFFX2_HVT U107 ( .A(n618), .Y(n372) );
  MUX21X2_HVT U108 ( .A1(n247), .A2(n417), .S0(n245), .Y(n584) );
  AO21X2_HVT U109 ( .A1(n328), .A2(n372), .A3(n413), .Y(n481) );
  AO21X1_HVT U111 ( .A1(n351), .A2(n413), .A3(n299), .Y(n435) );
  IBUFFX16_HVT U113 ( .A(n321), .Y(n236) );
  INVX4_HVT U117 ( .A(n362), .Y(n360) );
  XNOR2X2_HVT U121 ( .A1(n332), .A2(n331), .Y(n609) );
  IBUFFX2_HVT U123 ( .A(n332), .Y(n247) );
  MUX21X1_HVT U125 ( .A1(n340), .A2(n332), .S0(n351), .Y(n600) );
  NBUFFX4_HVT U126 ( .A(n310), .Y(n332) );
  MUX41X1_HVT U128 ( .A1(n397), .A3(n403), .A2(n364), .A4(n406), .S0(n271), 
        .S1(n239), .Y(n519) );
  IBUFFX16_HVT U134 ( .A(n319), .Y(n238) );
  MUX21X2_HVT U135 ( .A1(n315), .A2(n600), .S0(n239), .Y(n477) );
  MUX21X1_HVT U138 ( .A1(n346), .A2(n536), .S0(n258), .Y(n535) );
  INVX1_HVT U143 ( .A(n428), .Y(n402) );
  INVX2_HVT U144 ( .A(n362), .Y(n358) );
  MUX41X1_HVT U146 ( .A1(n262), .A3(n404), .A2(n200), .A4(n412), .S0(n240), 
        .S1(n361), .Y(n453) );
  IBUFFX16_HVT U147 ( .A(n324), .Y(n240) );
  AO21X1_HVT U148 ( .A1(n339), .A2(n623), .A3(n299), .Y(n461) );
  MUX21X2_HVT U149 ( .A1(n384), .A2(n569), .S0(n317), .Y(n568) );
  INVX0_HVT U150 ( .A(n600), .Y(n385) );
  MUX21X2_HVT U152 ( .A1(n566), .A2(n567), .S0(n241), .Y(n564) );
  IBUFFX16_HVT U153 ( .A(n325), .Y(n241) );
  MUX41X1_HVT U154 ( .A1(n572), .A3(n568), .A2(n570), .A4(n564), .S0(n337), 
        .S1(n242), .Y(n563) );
  INVX2_HVT U156 ( .A(n337), .Y(n338) );
  INVX1_HVT U157 ( .A(n354), .Y(n275) );
  INVX1_HVT U158 ( .A(n290), .Y(n291) );
  INVX1_HVT U160 ( .A(n278), .Y(n355) );
  NAND2X0_HVT U161 ( .A1(n516), .A2(n271), .Y(n259) );
  INVX0_HVT U165 ( .A(n348), .Y(n296) );
  INVX0_HVT U167 ( .A(n327), .Y(n286) );
  INVX0_HVT U168 ( .A(n429), .Y(n401) );
  INVX1_HVT U169 ( .A(in[5]), .Y(n337) );
  INVX1_HVT U170 ( .A(n335), .Y(n287) );
  INVX0_HVT U171 ( .A(n335), .Y(n269) );
  INVX0_HVT U174 ( .A(in[3]), .Y(n415) );
  INVX0_HVT U176 ( .A(in[7]), .Y(n253) );
  INVX1_HVT U180 ( .A(n355), .Y(n245) );
  INVX0_HVT U181 ( .A(n278), .Y(n258) );
  NBUFFX2_HVT U183 ( .A(in[0]), .Y(n278) );
  INVX1_HVT U184 ( .A(n323), .Y(n271) );
  INVX0_HVT U186 ( .A(n323), .Y(n279) );
  NAND2X0_HVT U187 ( .A1(n483), .A2(in[7]), .Y(n243) );
  NAND2X0_HVT U188 ( .A1(n473), .A2(n253), .Y(n244) );
  NAND2X0_HVT U189 ( .A1(n243), .A2(n244), .Y(out[5]) );
  INVX1_HVT U190 ( .A(n246), .Y(n589) );
  IBUFFX2_HVT U191 ( .A(n619), .Y(n371) );
  NAND2X0_HVT U193 ( .A1(n278), .A2(n344), .Y(n619) );
  MUX41X1_HVT U195 ( .A1(n484), .A3(n486), .A2(n487), .A4(n489), .S0(n336), 
        .S1(n338), .Y(n483) );
  MUX21X1_HVT U196 ( .A1(n247), .A2(n339), .S0(n245), .Y(n246) );
  NAND2X0_HVT U197 ( .A1(n341), .A2(n299), .Y(n248) );
  NAND2X0_HVT U199 ( .A1(n199), .A2(n327), .Y(n249) );
  NAND2X0_HVT U201 ( .A1(n248), .A2(n249), .Y(n536) );
  NBUFFX2_HVT U202 ( .A(n358), .Y(n328) );
  NAND2X0_HVT U203 ( .A1(n383), .A2(n250), .Y(n251) );
  NAND2X0_HVT U204 ( .A1(n562), .A2(n317), .Y(n252) );
  NAND2X0_HVT U205 ( .A1(n251), .A2(n252), .Y(n561) );
  IBUFFX2_HVT U206 ( .A(n317), .Y(n250) );
  NAND2X0_HVT U208 ( .A1(n556), .A2(n253), .Y(n254) );
  NAND2X0_HVT U209 ( .A1(n563), .A2(n303), .Y(n255) );
  NAND2X0_HVT U210 ( .A1(n255), .A2(n254), .Y(out[0]) );
  INVX1_HVT U211 ( .A(n604), .Y(n383) );
  NAND2X0_HVT U212 ( .A1(n541), .A2(n253), .Y(n256) );
  NAND2X0_HVT U213 ( .A1(n548), .A2(n303), .Y(n257) );
  NAND2X0_HVT U214 ( .A1(n256), .A2(n257), .Y(out[1]) );
  MUX21X2_HVT U215 ( .A1(n476), .A2(n477), .S0(n326), .Y(n475) );
  INVX1_HVT U216 ( .A(n596), .Y(n387) );
  NAND2X0_HVT U217 ( .A1(n517), .A2(n326), .Y(n260) );
  NAND2X0_HVT U218 ( .A1(n259), .A2(n260), .Y(n515) );
  INVX1_HVT U219 ( .A(in[0]), .Y(n354) );
  INVX1_HVT U220 ( .A(n344), .Y(n417) );
  MUX21X1_HVT U221 ( .A1(n304), .A2(n341), .S0(n278), .Y(n305) );
  MUX41X1_HVT U222 ( .A1(n438), .A3(n432), .A2(n447), .A4(n444), .S0(n337), 
        .S1(n303), .Y(out[7]) );
  INVX0_HVT U223 ( .A(n571), .Y(n261) );
  INVX1_HVT U224 ( .A(n261), .Y(n262) );
  NBUFFX2_HVT U225 ( .A(n362), .Y(n299) );
  MUX21X2_HVT U226 ( .A1(n482), .A2(n481), .S0(n325), .Y(n480) );
  INVX1_HVT U227 ( .A(n354), .Y(n276) );
  MUX41X1_HVT U228 ( .A1(n347), .A3(n196), .A2(n340), .A4(n383), .S0(n271), 
        .S1(n299), .Y(n520) );
  NBUFFX2_HVT U229 ( .A(n310), .Y(n333) );
  MUX41X1_HVT U230 ( .A1(n350), .A3(n378), .A2(n202), .A4(n377), .S0(n271), 
        .S1(n270), .Y(n557) );
  INVX1_HVT U231 ( .A(in[4]), .Y(n290) );
  NAND2X0_HVT U232 ( .A1(n385), .A2(n279), .Y(n263) );
  NAND2X0_HVT U233 ( .A1(n622), .A2(n326), .Y(n264) );
  NAND2X0_HVT U234 ( .A1(n264), .A2(n263), .Y(n569) );
  NAND2X0_HVT U235 ( .A1(n234), .A2(n279), .Y(n265) );
  NAND2X0_HVT U236 ( .A1(n623), .A2(n325), .Y(n266) );
  NAND2X0_HVT U237 ( .A1(n265), .A2(n266), .Y(n562) );
  NAND2X0_HVT U238 ( .A1(n306), .A2(n299), .Y(n267) );
  NAND2X0_HVT U239 ( .A1(n571), .A2(n328), .Y(n268) );
  NAND2X0_HVT U240 ( .A1(n268), .A2(n267), .Y(n567) );
  OR2X1_HVT U241 ( .A1(n235), .A2(n296), .Y(n623) );
  MUX41X1_HVT U242 ( .A1(n558), .A3(n561), .A2(n557), .A4(n560), .S0(n338), 
        .S1(n269), .Y(n556) );
  NAND2X0_HVT U243 ( .A1(n411), .A2(n272), .Y(n273) );
  NAND2X0_HVT U244 ( .A1(n368), .A2(n328), .Y(n274) );
  NAND2X0_HVT U245 ( .A1(n274), .A2(n273), .Y(n482) );
  IBUFFX2_HVT U246 ( .A(n329), .Y(n272) );
  INVX1_HVT U247 ( .A(n420), .Y(n411) );
  MUX41X1_HVT U248 ( .A1(n480), .A3(n475), .A2(n478), .A4(n474), .S0(n337), 
        .S1(n269), .Y(n473) );
  INVX0_HVT U249 ( .A(n354), .Y(n351) );
  INVX1_HVT U250 ( .A(n369), .Y(n277) );
  INVX1_HVT U251 ( .A(n620), .Y(n369) );
  NAND2X0_HVT U252 ( .A1(n278), .A2(n626), .Y(n620) );
  INVX0_HVT U253 ( .A(n617), .Y(n375) );
  MUX41X1_HVT U254 ( .A1(n608), .A3(n389), .A2(n607), .A4(n387), .S0(n279), 
        .S1(n270), .Y(n547) );
  MUX41X1_HVT U255 ( .A1(n555), .A3(n552), .A2(n553), .A4(n549), .S0(n337), 
        .S1(n287), .Y(n548) );
  MUX21X2_HVT U256 ( .A1(n495), .A2(n496), .S0(n336), .Y(n494) );
  NAND2X0_HVT U257 ( .A1(n573), .A2(n322), .Y(n280) );
  NAND2X0_HVT U258 ( .A1(n574), .A2(n279), .Y(n281) );
  NAND2X0_HVT U259 ( .A1(n280), .A2(n281), .Y(n572) );
  MUX21X1_HVT U260 ( .A1(n386), .A2(n378), .S0(n329), .Y(n574) );
  NAND2X0_HVT U261 ( .A1(n315), .A2(n282), .Y(n283) );
  NAND2X0_HVT U262 ( .A1(n577), .A2(n329), .Y(n284) );
  NAND2X0_HVT U263 ( .A1(n283), .A2(n284), .Y(n441) );
  IBUFFX2_HVT U264 ( .A(n327), .Y(n282) );
  MUX21X1_HVT U265 ( .A1(n593), .A2(n429), .S0(n286), .Y(n285) );
  MUX41X1_HVT U266 ( .A1(n370), .A3(n346), .A2(n522), .A4(n407), .S0(n270), 
        .S1(n279), .Y(n521) );
  NAND2X0_HVT U267 ( .A1(n308), .A2(n299), .Y(n288) );
  NAND2X0_HVT U268 ( .A1(n584), .A2(n328), .Y(n289) );
  NAND2X0_HVT U269 ( .A1(n288), .A2(n289), .Y(n440) );
  OA21X1_HVT U270 ( .A1(n387), .A2(n299), .A3(n565), .Y(n439) );
  NAND2X0_HVT U271 ( .A1(n471), .A2(n271), .Y(n292) );
  NAND2X0_HVT U272 ( .A1(n472), .A2(n326), .Y(n293) );
  NAND2X0_HVT U273 ( .A1(n292), .A2(n293), .Y(n468) );
  NAND2X0_HVT U274 ( .A1(n452), .A2(n253), .Y(n294) );
  NAND2X0_HVT U275 ( .A1(n459), .A2(n303), .Y(n295) );
  NAND2X0_HVT U276 ( .A1(n294), .A2(n295), .Y(out[6]) );
  MUX41X1_HVT U277 ( .A1(n464), .A3(n468), .A2(n460), .A4(n466), .S0(n338), 
        .S1(n269), .Y(n459) );
  NAND2X0_HVT U278 ( .A1(n446), .A2(n300), .Y(n297) );
  NAND2X0_HVT U279 ( .A1(n445), .A2(n287), .Y(n298) );
  NAND2X0_HVT U280 ( .A1(n298), .A2(n297), .Y(n444) );
  INVX1_HVT U281 ( .A(n347), .Y(n413) );
  NBUFFX2_HVT U282 ( .A(n626), .Y(n350) );
  INVX0_HVT U283 ( .A(n333), .Y(n309) );
  INVX1_HVT U284 ( .A(n598), .Y(n386) );
  NAND2X0_HVT U285 ( .A1(n450), .A2(n300), .Y(n301) );
  NAND2X0_HVT U286 ( .A1(n448), .A2(n269), .Y(n302) );
  NAND2X0_HVT U287 ( .A1(n301), .A2(n302), .Y(n447) );
  INVX0_HVT U288 ( .A(n334), .Y(n300) );
  INVX0_HVT U289 ( .A(n307), .Y(n581) );
  MUX41X1_HVT U290 ( .A1(n262), .A3(n196), .A2(n340), .A4(n399), .S0(n271), 
        .S1(n299), .Y(n570) );
  MUX21X1_HVT U291 ( .A1(n415), .A2(n349), .S0(n354), .Y(n306) );
  MUX21X1_HVT U292 ( .A1(n339), .A2(n330), .S0(n218), .Y(n604) );
  MUX41X1_HVT U293 ( .A1(n611), .A3(n545), .A2(n408), .A4(n524), .S0(n359), 
        .S1(n323), .Y(n523) );
  MUX41X1_HVT U294 ( .A1(n531), .A3(n528), .A2(n529), .A4(n526), .S0(n337), 
        .S1(n287), .Y(n525) );
  MUX21X2_HVT U295 ( .A1(n525), .A2(n532), .S0(n303), .Y(out[2]) );
  INVX0_HVT U296 ( .A(n306), .Y(n602) );
  OA21X2_HVT U297 ( .A1(n366), .A2(n270), .A3(n604), .Y(n550) );
  OA21X2_HVT U298 ( .A1(n365), .A2(n270), .A3(n374), .Y(n476) );
  AO21X2_HVT U299 ( .A1(n354), .A2(n350), .A3(n270), .Y(n469) );
  MUX41X1_HVT U300 ( .A1(n587), .A3(n381), .A2(n382), .A4(n380), .S0(n279), 
        .S1(n270), .Y(n560) );
  NBUFFX2_HVT U301 ( .A(in[7]), .Y(n303) );
  INVX1_HVT U302 ( .A(n431), .Y(n399) );
  NBUFFX2_HVT U303 ( .A(n415), .Y(n330) );
  MUX41X1_HVT U304 ( .A1(n602), .A3(n605), .A2(n395), .A4(n414), .S0(n271), 
        .S1(n272), .Y(n486) );
  MUX21X1_HVT U305 ( .A1(n350), .A2(n342), .S0(n355), .Y(n307) );
  INVX1_HVT U306 ( .A(n626), .Y(n416) );
  MUX21X1_HVT U307 ( .A1(n309), .A2(n347), .S0(n354), .Y(n308) );
  NBUFFX2_HVT U308 ( .A(n609), .Y(n341) );
  INVX0_HVT U309 ( .A(in[1]), .Y(n334) );
  NBUFFX2_HVT U310 ( .A(n625), .Y(n347) );
  NBUFFX2_HVT U311 ( .A(n625), .Y(n349) );
  NBUFFX2_HVT U312 ( .A(n625), .Y(n348) );
  AND2X1_HVT U313 ( .A1(n348), .A2(n610), .Y(n311) );
  MUX21X1_HVT U314 ( .A1(n341), .A2(n416), .S0(n275), .Y(n594) );
  MUX21X1_HVT U315 ( .A1(n342), .A2(n345), .S0(n278), .Y(n467) );
  MUX21X1_HVT U316 ( .A1(n418), .A2(n331), .S0(n278), .Y(n586) );
  MUX21X1_HVT U317 ( .A1(n413), .A2(n418), .S0(n353), .Y(n592) );
  MUX21X1_HVT U318 ( .A1(n416), .A2(n417), .S0(n352), .Y(n458) );
  MUX21X1_HVT U319 ( .A1(n332), .A2(n414), .S0(n276), .Y(n479) );
  MUX21X1_HVT U320 ( .A1(n416), .A2(n332), .S0(n276), .Y(n456) );
  NAND2X0_HVT U321 ( .A1(n330), .A2(n332), .Y(n625) );
  MUX21X1_HVT U322 ( .A1(n416), .A2(n341), .S0(n351), .Y(n426) );
  MUX21X1_HVT U323 ( .A1(n331), .A2(n413), .S0(n353), .Y(n595) );
  MUX21X1_HVT U324 ( .A1(n332), .A2(n349), .S0(n352), .Y(n522) );
  MUX21X1_HVT U325 ( .A1(n200), .A2(n199), .S0(n275), .Y(n421) );
  MUX21X1_HVT U326 ( .A1(n332), .A2(n340), .S0(n237), .Y(n585) );
  XNOR2X1_HVT U327 ( .A1(n347), .A2(n276), .Y(n312) );
  MUX21X1_HVT U328 ( .A1(n346), .A2(n348), .S0(n276), .Y(n607) );
  MUX21X1_HVT U329 ( .A1(n592), .A2(n311), .S0(n326), .Y(n500) );
  MUX21X1_HVT U330 ( .A1(n339), .A2(n414), .S0(n275), .Y(n591) );
  MUX21X1_HVT U331 ( .A1(n342), .A2(n349), .S0(n245), .Y(n420) );
  INVX1_HVT U332 ( .A(n342), .Y(n414) );
  MUX21X1_HVT U333 ( .A1(n350), .A2(n349), .S0(n218), .Y(n611) );
  MUX21X1_HVT U334 ( .A1(n330), .A2(n417), .S0(n353), .Y(n582) );
  MUX21X1_HVT U335 ( .A1(n410), .A2(n312), .S0(n325), .Y(n503) );
  MUX21X1_HVT U336 ( .A1(n417), .A2(n330), .S0(n275), .Y(n429) );
  MUX21X1_HVT U337 ( .A1(n330), .A2(n348), .S0(n237), .Y(n428) );
  AND2X1_HVT U338 ( .A1(n277), .A2(n348), .Y(n313) );
  XOR2X1_HVT U339 ( .A1(n346), .A2(n352), .Y(n578) );
  MUX21X1_HVT U340 ( .A1(n345), .A2(n331), .S0(n245), .Y(n606) );
  MUX21X1_HVT U341 ( .A1(n331), .A2(n333), .S0(n275), .Y(n580) );
  AND2X1_HVT U342 ( .A1(n237), .A2(n332), .Y(n314) );
  MUX21X1_HVT U343 ( .A1(n330), .A2(n346), .S0(n275), .Y(n423) );
  MUX21X1_HVT U344 ( .A1(n345), .A2(n333), .S0(n351), .Y(n506) );
  NBUFFX2_HVT U345 ( .A(n358), .Y(n327) );
  NBUFFX2_HVT U346 ( .A(n358), .Y(n329) );
  NBUFFX2_HVT U347 ( .A(n609), .Y(n339) );
  NBUFFX2_HVT U348 ( .A(n609), .Y(n340) );
  MUX21X1_HVT U349 ( .A1(n413), .A2(n417), .S0(n276), .Y(n575) );
  MUX21X1_HVT U350 ( .A1(n347), .A2(n343), .S0(n237), .Y(n485) );
  MUX21X1_HVT U351 ( .A1(n505), .A2(n507), .S0(n336), .Y(n504) );
  NBUFFX2_HVT U352 ( .A(n621), .Y(n342) );
  AND2X1_HVT U353 ( .A1(n345), .A2(n258), .Y(n315) );
  AND2X1_HVT U354 ( .A1(n417), .A2(n355), .Y(n316) );
  NBUFFX2_HVT U355 ( .A(n624), .Y(n344) );
  NBUFFX2_HVT U356 ( .A(n624), .Y(n346) );
  NBUFFX2_HVT U357 ( .A(n624), .Y(n345) );
  NBUFFX2_HVT U358 ( .A(n621), .Y(n343) );
  NBUFFX2_HVT U359 ( .A(n415), .Y(n331) );
  NBUFFX2_HVT U360 ( .A(n356), .Y(n324) );
  NBUFFX2_HVT U361 ( .A(n356), .Y(n326) );
  NBUFFX2_HVT U362 ( .A(n356), .Y(n325) );
  XNOR2X1_HVT U363 ( .A1(n299), .A2(n321), .Y(n317) );
  NBUFFX2_HVT U364 ( .A(n357), .Y(n323) );
  NBUFFX2_HVT U365 ( .A(n357), .Y(n321) );
  NBUFFX2_HVT U366 ( .A(n357), .Y(n322) );
  NBUFFX2_HVT U367 ( .A(n356), .Y(n319) );
  NBUFFX2_HVT U368 ( .A(n356), .Y(n320) );
  NBUFFX2_HVT U369 ( .A(n356), .Y(n318) );
  INVX1_HVT U370 ( .A(n334), .Y(n336) );
  INVX1_HVT U371 ( .A(n334), .Y(n335) );
  MUX21X1_HVT U372 ( .A1(n416), .A2(n202), .S0(n237), .Y(n419) );
  MUX21X1_HVT U373 ( .A1(n350), .A2(n202), .S0(n352), .Y(n470) );
  MUX21X1_HVT U374 ( .A1(n417), .A2(n414), .S0(n218), .Y(n511) );
  MUX21X1_HVT U375 ( .A1(n491), .A2(n492), .S0(n336), .Y(n490) );
  MUX21X1_HVT U376 ( .A1(n343), .A2(n202), .S0(n276), .Y(n530) );
  MUX21X1_HVT U377 ( .A1(n332), .A2(n304), .S0(n351), .Y(n598) );
  MUX21X1_HVT U378 ( .A1(n202), .A2(n350), .S0(n278), .Y(n425) );
  MUX21X1_HVT U379 ( .A1(n202), .A2(n343), .S0(n278), .Y(n424) );
  NBUFFX2_HVT U380 ( .A(in[2]), .Y(n357) );
  NBUFFX2_HVT U381 ( .A(in[2]), .Y(n356) );
  MUX21X1_HVT U382 ( .A1(n413), .A2(n247), .S0(n352), .Y(n493) );
  XOR2X1_HVT U383 ( .A1(n353), .A2(n247), .Y(n576) );
  MUX21X1_HVT U384 ( .A1(n247), .A2(n346), .S0(n353), .Y(n430) );
  MUX21X1_HVT U385 ( .A1(n345), .A2(n247), .S0(n276), .Y(n427) );
  MUX21X1_HVT U386 ( .A1(n247), .A2(n416), .S0(n353), .Y(n601) );
  MUX21X1_HVT U387 ( .A1(n330), .A2(n247), .S0(n351), .Y(n422) );
  MUX21X1_HVT U388 ( .A1(n343), .A2(n247), .S0(n218), .Y(n596) );
  MUX21X1_HVT U389 ( .A1(n247), .A2(n414), .S0(n245), .Y(n431) );
  MUX21X1_HVT U390 ( .A1(n247), .A2(n626), .S0(n352), .Y(n608) );
  INVX0_HVT U391 ( .A(n614), .Y(n363) );
  INVX0_HVT U392 ( .A(n587), .Y(n364) );
  INVX0_HVT U393 ( .A(n527), .Y(n365) );
  INVX0_HVT U394 ( .A(n488), .Y(n366) );
  INVX0_HVT U395 ( .A(n623), .Y(n367) );
  INVX0_HVT U396 ( .A(n622), .Y(n368) );
  INVX0_HVT U397 ( .A(n583), .Y(n370) );
  INVX0_HVT U398 ( .A(n590), .Y(n373) );
  INVX0_HVT U399 ( .A(n612), .Y(n374) );
  INVX0_HVT U400 ( .A(n613), .Y(n376) );
  INVX0_HVT U401 ( .A(n611), .Y(n377) );
  INVX0_HVT U402 ( .A(n610), .Y(n378) );
  INVX0_HVT U403 ( .A(n608), .Y(n379) );
  INVX0_HVT U404 ( .A(n607), .Y(n380) );
  INVX0_HVT U405 ( .A(n606), .Y(n381) );
  INVX0_HVT U406 ( .A(n605), .Y(n382) );
  INVX0_HVT U407 ( .A(n601), .Y(n384) );
  INVX0_HVT U408 ( .A(n595), .Y(n388) );
  INVX0_HVT U409 ( .A(n594), .Y(n389) );
  INVX0_HVT U410 ( .A(n592), .Y(n390) );
  INVX0_HVT U411 ( .A(n591), .Y(n391) );
  INVX0_HVT U412 ( .A(n588), .Y(n392) );
  INVX0_HVT U413 ( .A(n586), .Y(n393) );
  INVX0_HVT U414 ( .A(n585), .Y(n394) );
  INVX0_HVT U415 ( .A(n579), .Y(n397) );
  INVX0_HVT U416 ( .A(n616), .Y(n398) );
  INVX0_HVT U417 ( .A(n430), .Y(n400) );
  INVX0_HVT U418 ( .A(n427), .Y(n403) );
  INVX0_HVT U419 ( .A(n426), .Y(n404) );
  INVX0_HVT U420 ( .A(n425), .Y(n405) );
  INVX0_HVT U421 ( .A(n424), .Y(n406) );
  INVX0_HVT U422 ( .A(n423), .Y(n407) );
  INVX0_HVT U423 ( .A(n422), .Y(n408) );
  INVX0_HVT U424 ( .A(n470), .Y(n409) );
  INVX0_HVT U425 ( .A(n421), .Y(n410) );
  INVX0_HVT U426 ( .A(n419), .Y(n412) );
endmodule

