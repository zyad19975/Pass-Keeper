
module Mix_Column ( in, out );
  input [127:0] in;
  output [127:0] out;
  wire   n15, n16, n17, n19, n21, n22, n23, n24, n26, n27, n28, n29, n30, n31,
         n32, n34, n35, n36, n38, n39, n44, n45, n46, n47, n50, n53, n54, n57,
         n58, n60, n61, n63, n64, n65, n66, n67, n69, n70, n71, n72, n74, n75,
         n76, n77, n78, n80, n81, n83, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n99, n100, n101, n102, n104, n105, n106, n108, n111,
         n115, n116, n117, n118, n119, n121, n122, n123, n124, n129, n130,
         n133, n135, n136, n137, n138, n140, n141, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n153, n154, n155, n157, n158, n159,
         n160, n162, n163, n167, n168, n169, n170, n172, n174, n176, n177,
         n178, n179, n180, n181, n183, n184, n186, n187, n188, n189, n190,
         n193, n195, n196, n197, n199, n200, n201, n202, n204, n207, n208,
         n209, n211, n212, n215, n217, n218, n219, n221, n1, n2, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n18, n20, n25, n33, n37, n40,
         n41, n42, n43, n48, n49, n51, n52, n55, n56, n59, n62, n68, n73, n79,
         n82, n84, n85, n97, n98, n103, n107, n109, n110, n112, n113, n114,
         n120, n125, n126, n127, n128, n131, n132, n134, n139, n142, n152,
         n156, n161, n164, n165, n166, n171, n173, n175, n182, n185, n191,
         n192, n194, n198, n203, n205, n206, n210, n213, n214, n216, n220,
         n222, n223, n224, n225, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2X2_HVT U21 ( .A1(in[78]), .A2(in[70]), .Y(n29) );
  XOR2X2_HVT U24 ( .A1(n67), .A2(n66), .Y(out[76]) );
  XOR2X2_HVT U63 ( .A1(n117), .A2(n116), .Y(out[4]) );
  XOR2X2_HVT U155 ( .A1(n212), .A2(n211), .Y(out[108]) );
  XNOR3X1_HVT U225 ( .A1(n559), .A2(n460), .A3(n457), .Y(n69) );
  INVX1_HVT U1 ( .A(n236), .Y(n1) );
  INVX1_HVT U2 ( .A(in[39]), .Y(n236) );
  XOR3X2_HVT U3 ( .A1(n105), .A2(n2), .A3(n104), .Y(out[56]) );
  IBUFFX16_HVT U4 ( .A(n581), .Y(n2) );
  XOR3X2_HVT U5 ( .A1(n102), .A2(n511), .A3(n130), .Y(out[42]) );
  INVX1_HVT U6 ( .A(in[56]), .Y(n386) );
  XOR2X1_HVT U7 ( .A1(in[118]), .A2(n569), .Y(n197) );
  XOR3X2_HVT U8 ( .A1(n263), .A2(n492), .A3(n143), .Y(n141) );
  INVX1_HVT U9 ( .A(n503), .Y(n4) );
  INVX1_HVT U10 ( .A(in[99]), .Y(n503) );
  INVX1_HVT U11 ( .A(in[89]), .Y(n305) );
  XOR2X2_HVT U12 ( .A1(n269), .A2(n7), .Y(n365) );
  XNOR2X2_HVT U13 ( .A1(n210), .A2(n206), .Y(n489) );
  XOR2X1_HVT U14 ( .A1(n550), .A2(in[24]), .Y(n159) );
  IBUFFX2_HVT U15 ( .A(in[24]), .Y(n576) );
  INVX1_HVT U16 ( .A(in[11]), .Y(n521) );
  IBUFFX2_HVT U17 ( .A(n22), .Y(n48) );
  INVX2_HVT U18 ( .A(n521), .Y(n522) );
  INVX1_HVT U19 ( .A(in[89]), .Y(n165) );
  INVX2_HVT U20 ( .A(in[108]), .Y(n103) );
  INVX0_HVT U22 ( .A(n164), .Y(n5) );
  INVX1_HVT U23 ( .A(in[8]), .Y(n164) );
  NBUFFX2_HVT U25 ( .A(in[53]), .Y(n391) );
  XOR3X1_HVT U26 ( .A1(in[123]), .A2(in[115]), .A3(n215), .Y(n431) );
  XOR3X2_HVT U27 ( .A1(n148), .A2(n163), .A3(n318), .Y(out[17]) );
  INVX1_HVT U28 ( .A(in[35]), .Y(n6) );
  INVX2_HVT U29 ( .A(n6), .Y(n7) );
  XOR3X2_HVT U30 ( .A1(n252), .A2(n56), .A3(n253), .Y(n139) );
  INVX1_HVT U31 ( .A(n133), .Y(n401) );
  INVX0_HVT U32 ( .A(in[83]), .Y(n49) );
  XNOR2X1_HVT U33 ( .A1(in[12]), .A2(n480), .Y(n154) );
  XOR3X2_HVT U34 ( .A1(in[35]), .A2(n8), .A3(n9), .Y(n366) );
  IBUFFX16_HVT U35 ( .A(n353), .Y(n8) );
  IBUFFX16_HVT U36 ( .A(n352), .Y(n9) );
  INVX0_HVT U37 ( .A(in[119]), .Y(n532) );
  XOR3X2_HVT U38 ( .A1(n89), .A2(n391), .A3(n321), .Y(out[61]) );
  XOR2X1_HVT U39 ( .A1(in[8]), .A2(n545), .Y(n15) );
  XOR2X1_HVT U40 ( .A1(in[125]), .A2(in[110]), .Y(n219) );
  INVX1_HVT U41 ( .A(in[125]), .Y(n309) );
  INVX1_HVT U42 ( .A(n346), .Y(n10) );
  INVX1_HVT U43 ( .A(in[22]), .Y(n346) );
  INVX1_HVT U44 ( .A(n199), .Y(n340) );
  NAND2X0_HVT U45 ( .A1(n18), .A2(n12), .Y(n13) );
  NAND2X0_HVT U46 ( .A1(n11), .A2(in[90]), .Y(n14) );
  NAND2X0_HVT U47 ( .A1(n13), .A2(n14), .Y(n71) );
  INVX0_HVT U48 ( .A(in[82]), .Y(n11) );
  IBUFFX2_HVT U49 ( .A(in[90]), .Y(n12) );
  INVX0_HVT U50 ( .A(n11), .Y(n18) );
  INVX1_HVT U51 ( .A(in[34]), .Y(n20) );
  INVX1_HVT U52 ( .A(n20), .Y(n25) );
  XOR2X2_HVT U53 ( .A1(in[126]), .A2(n568), .Y(n218) );
  XOR3X2_HVT U54 ( .A1(n399), .A2(n562), .A3(n423), .Y(n54) );
  XOR3X1_HVT U55 ( .A1(n528), .A2(n323), .A3(n118), .Y(n117) );
  IBUFFX2_HVT U56 ( .A(in[86]), .Y(n471) );
  XNOR2X2_HVT U57 ( .A1(n582), .A2(in[104]), .Y(n26) );
  INVX0_HVT U58 ( .A(in[98]), .Y(n504) );
  XOR2X2_HVT U59 ( .A1(in[98]), .A2(n571), .Y(n308) );
  NBUFFX2_HVT U60 ( .A(n71), .Y(n33) );
  NAND2X0_HVT U61 ( .A1(n478), .A2(n135), .Y(n41) );
  NAND2X0_HVT U62 ( .A1(n37), .A2(n40), .Y(n42) );
  NAND2X0_HVT U64 ( .A1(n41), .A2(n42), .Y(out[3]) );
  INVX0_HVT U65 ( .A(n478), .Y(n37) );
  INVX1_HVT U66 ( .A(n135), .Y(n40) );
  INVX0_HVT U67 ( .A(in[11]), .Y(n412) );
  XOR3X2_HVT U68 ( .A1(n190), .A2(n43), .A3(n48), .Y(out[106]) );
  IBUFFX16_HVT U69 ( .A(n504), .Y(n43) );
  IBUFFX2_HVT U70 ( .A(in[77]), .Y(n459) );
  XNOR2X2_HVT U71 ( .A1(n264), .A2(in[97]), .Y(n190) );
  INVX1_HVT U72 ( .A(n264), .Y(n265) );
  XOR3X2_HVT U73 ( .A1(n103), .A2(n274), .A3(n301), .Y(n201) );
  INVX2_HVT U74 ( .A(in[99]), .Y(n529) );
  XOR2X2_HVT U75 ( .A1(in[44]), .A2(in[52]), .Y(n108) );
  INVX1_HVT U76 ( .A(n49), .Y(n51) );
  NBUFFX2_HVT U77 ( .A(n160), .Y(n52) );
  INVX2_HVT U78 ( .A(in[123]), .Y(n465) );
  INVX1_HVT U79 ( .A(n149), .Y(n266) );
  NBUFFX16_HVT U80 ( .A(in[36]), .Y(n458) );
  INVX1_HVT U81 ( .A(in[72]), .Y(n472) );
  XOR3X2_HVT U82 ( .A1(n151), .A2(n368), .A3(n372), .Y(out[29]) );
  INVX1_HVT U83 ( .A(n151), .Y(n484) );
  INVX1_HVT U84 ( .A(n495), .Y(n290) );
  XOR2X2_HVT U85 ( .A1(n112), .A2(in[94]), .Y(n296) );
  INVX1_HVT U86 ( .A(in[82]), .Y(n399) );
  XOR2X2_HVT U87 ( .A1(n512), .A2(n552), .Y(n269) );
  INVX1_HVT U88 ( .A(in[90]), .Y(n409) );
  XOR2X2_HVT U89 ( .A1(in[57]), .A2(n311), .Y(n119) );
  INVX1_HVT U90 ( .A(in[49]), .Y(n55) );
  XOR2X2_HVT U91 ( .A1(in[121]), .A2(in[97]), .Y(n21) );
  XOR2X1_HVT U92 ( .A1(in[28]), .A2(n480), .Y(n479) );
  XOR2X1_HVT U93 ( .A1(n530), .A2(in[123]), .Y(n253) );
  INVX1_HVT U94 ( .A(in[50]), .Y(n352) );
  XOR3X2_HVT U95 ( .A1(n575), .A2(n379), .A3(n55), .Y(n390) );
  INVX1_HVT U96 ( .A(in[55]), .Y(n575) );
  IBUFFX16_HVT U97 ( .A(n533), .Y(n56) );
  XNOR2X2_HVT U98 ( .A1(n103), .A2(in[116]), .Y(n199) );
  INVX2_HVT U99 ( .A(n357), .Y(n473) );
  XOR3X2_HVT U100 ( .A1(n254), .A2(n255), .A3(n483), .Y(n96) );
  INVX1_HVT U101 ( .A(n83), .Y(n315) );
  XOR2X2_HVT U102 ( .A1(in[104]), .A2(n567), .Y(n208) );
  INVX2_HVT U103 ( .A(n274), .Y(n498) );
  XOR3X2_HVT U104 ( .A1(n184), .A2(n439), .A3(n179), .Y(out[109]) );
  IBUFFX2_HVT U105 ( .A(in[101]), .Y(n439) );
  INVX2_HVT U106 ( .A(n502), .Y(n520) );
  INVX2_HVT U107 ( .A(in[4]), .Y(n480) );
  XNOR2X2_HVT U108 ( .A1(n497), .A2(n567), .Y(n177) );
  NAND2X0_HVT U109 ( .A1(n389), .A2(n62), .Y(n68) );
  NAND2X0_HVT U110 ( .A1(n59), .A2(n370), .Y(n73) );
  NAND2X0_HVT U111 ( .A1(n68), .A2(n73), .Y(out[84]) );
  INVX1_HVT U112 ( .A(n389), .Y(n59) );
  INVX0_HVT U113 ( .A(n370), .Y(n62) );
  XOR3X2_HVT U114 ( .A1(n79), .A2(n378), .A3(n408), .Y(out[72]) );
  XNOR2X2_HVT U115 ( .A1(in[88]), .A2(n578), .Y(n79) );
  XOR2X1_HVT U116 ( .A1(in[62]), .A2(n555), .Y(n137) );
  INVX0_HVT U117 ( .A(n387), .Y(n166) );
  XOR2X2_HVT U118 ( .A1(in[84]), .A2(in[76]), .Y(n50) );
  XOR3X2_HVT U119 ( .A1(n268), .A2(n44), .A3(n45), .Y(out[89]) );
  INVX1_HVT U120 ( .A(n580), .Y(n303) );
  XOR2X1_HVT U121 ( .A1(in[32]), .A2(n1), .Y(n133) );
  INVX0_HVT U122 ( .A(in[52]), .Y(n537) );
  XOR3X1_HVT U123 ( .A1(n465), .A2(n496), .A3(n199), .Y(n221) );
  INVX0_HVT U124 ( .A(n522), .Y(n206) );
  IBUFFX2_HVT U125 ( .A(in[26]), .Y(n235) );
  INVX0_HVT U126 ( .A(n578), .Y(n82) );
  INVX2_HVT U127 ( .A(in[80]), .Y(n578) );
  INVX1_HVT U128 ( .A(n237), .Y(n107) );
  XOR2X2_HVT U129 ( .A1(n541), .A2(n367), .Y(n196) );
  INVX1_HVT U130 ( .A(in[3]), .Y(n427) );
  INVX1_HVT U131 ( .A(n427), .Y(n367) );
  XOR3X1_HVT U132 ( .A1(n547), .A2(n523), .A3(n172), .Y(n170) );
  NAND2X0_HVT U133 ( .A1(n80), .A2(n535), .Y(n97) );
  NAND2X0_HVT U134 ( .A1(n84), .A2(n85), .Y(n98) );
  NAND2X0_HVT U135 ( .A1(n97), .A2(n98), .Y(out[68]) );
  INVX0_HVT U136 ( .A(n80), .Y(n84) );
  INVX0_HVT U137 ( .A(n535), .Y(n85) );
  NBUFFX2_HVT U138 ( .A(in[127]), .Y(n571) );
  XNOR2X1_HVT U139 ( .A1(in[80]), .A2(in[72]), .Y(n411) );
  INVX0_HVT U140 ( .A(n82), .Y(n237) );
  INVX0_HVT U141 ( .A(in[25]), .Y(n331) );
  XNOR2X2_HVT U142 ( .A1(n424), .A2(n192), .Y(n423) );
  INVX1_HVT U143 ( .A(n527), .Y(n327) );
  INVX0_HVT U144 ( .A(n65), .Y(n579) );
  XOR3X2_HVT U145 ( .A1(n539), .A2(n507), .A3(n146), .Y(out[23]) );
  IBUFFX2_HVT U146 ( .A(in[12]), .Y(n384) );
  INVX0_HVT U147 ( .A(in[85]), .Y(n426) );
  INVX1_HVT U148 ( .A(in[106]), .Y(n516) );
  XNOR2X2_HVT U149 ( .A1(n107), .A2(n580), .Y(n47) );
  XOR3X1_HVT U150 ( .A1(n89), .A2(n437), .A3(n348), .Y(out[46]) );
  XOR2X2_HVT U151 ( .A1(in[68]), .A2(in[92]), .Y(n53) );
  XNOR2X2_HVT U152 ( .A1(n558), .A2(in[58]), .Y(n483) );
  INVX0_HVT U153 ( .A(n323), .Y(n110) );
  XNOR2X2_HVT U154 ( .A1(n576), .A2(n548), .Y(n174) );
  XOR2X2_HVT U156 ( .A1(n566), .A2(in[90]), .Y(n38) );
  INVX0_HVT U157 ( .A(n230), .Y(n228) );
  INVX0_HVT U158 ( .A(in[28]), .Y(n528) );
  XOR3X2_HVT U159 ( .A1(n214), .A2(in[19]), .A3(n109), .Y(n448) );
  IBUFFX16_HVT U160 ( .A(n381), .Y(n109) );
  XNOR2X2_HVT U161 ( .A1(n405), .A2(n110), .Y(n243) );
  INVX1_HVT U162 ( .A(n426), .Y(n112) );
  XOR3X2_HVT U163 ( .A1(n30), .A2(n113), .A3(n114), .Y(out[69]) );
  IBUFFX16_HVT U164 ( .A(n459), .Y(n113) );
  IBUFFX16_HVT U165 ( .A(n53), .Y(n114) );
  NAND2X0_HVT U166 ( .A1(n140), .A2(n463), .Y(n126) );
  NAND2X0_HVT U167 ( .A1(n120), .A2(n125), .Y(n127) );
  NAND2X0_HVT U168 ( .A1(n126), .A2(n127), .Y(out[36]) );
  INVX0_HVT U169 ( .A(n140), .Y(n120) );
  INVX1_HVT U170 ( .A(n463), .Y(n125) );
  INVX4_HVT U171 ( .A(n214), .Y(n350) );
  XOR3X2_HVT U172 ( .A1(n119), .A2(n105), .A3(n400), .Y(out[49]) );
  XOR2X1_HVT U173 ( .A1(in[96]), .A2(in[120]), .Y(n207) );
  NAND2X0_HVT U174 ( .A1(n139), .A2(n204), .Y(n132) );
  NAND2X0_HVT U175 ( .A1(n128), .A2(n131), .Y(n134) );
  NAND2X0_HVT U176 ( .A1(n132), .A2(n134), .Y(out[115]) );
  INVX1_HVT U177 ( .A(n139), .Y(n128) );
  INVX0_HVT U178 ( .A(n204), .Y(n131) );
  INVX1_HVT U179 ( .A(in[119]), .Y(n583) );
  INVX0_HVT U180 ( .A(n532), .Y(n252) );
  INVX2_HVT U181 ( .A(n529), .Y(n530) );
  XOR3X1_HVT U182 ( .A1(n561), .A2(n506), .A3(n70), .Y(n527) );
  XOR2X2_HVT U183 ( .A1(n351), .A2(n520), .Y(n70) );
  NAND2X0_HVT U184 ( .A1(n176), .A2(n173), .Y(n156) );
  NAND2X0_HVT U185 ( .A1(n142), .A2(n152), .Y(n161) );
  NAND2X0_HVT U186 ( .A1(n156), .A2(n161), .Y(out[12]) );
  INVX0_HVT U187 ( .A(n176), .Y(n142) );
  INVX0_HVT U188 ( .A(n173), .Y(n152) );
  XOR2X2_HVT U189 ( .A1(in[81]), .A2(n165), .Y(n267) );
  XOR3X2_HVT U190 ( .A1(n320), .A2(n164), .A3(n381), .Y(n318) );
  INVX0_HVT U191 ( .A(in[10]), .Y(n510) );
  XNOR2X2_HVT U192 ( .A1(in[62]), .A2(n391), .Y(n540) );
  XOR2X2_HVT U193 ( .A1(in[17]), .A2(in[9]), .Y(n168) );
  XOR3X2_HVT U194 ( .A1(n399), .A2(n166), .A3(n239), .Y(n213) );
  XOR2X1_HVT U195 ( .A1(in[62]), .A2(in[54]), .Y(n124) );
  XOR3X2_HVT U196 ( .A1(n567), .A2(n516), .A3(n496), .Y(n229) );
  INVX0_HVT U197 ( .A(n516), .Y(n517) );
  XOR3X2_HVT U198 ( .A1(n94), .A2(n171), .A3(n95), .Y(out[5]) );
  IBUFFX16_HVT U199 ( .A(in[13]), .Y(n171) );
  XOR3X2_HVT U200 ( .A1(n543), .A2(in[4]), .A3(n428), .Y(n173) );
  NBUFFX2_HVT U201 ( .A(in[127]), .Y(n570) );
  XOR3X2_HVT U202 ( .A1(n39), .A2(n399), .A3(n304), .Y(out[90]) );
  NAND2X0_HVT U203 ( .A1(n34), .A2(n349), .Y(n185) );
  NAND2X0_HVT U204 ( .A1(n175), .A2(n182), .Y(n191) );
  NAND2X0_HVT U205 ( .A1(n185), .A2(n191), .Y(out[92]) );
  INVX1_HVT U206 ( .A(n34), .Y(n175) );
  INVX0_HVT U207 ( .A(n349), .Y(n182) );
  INVX0_HVT U208 ( .A(n580), .Y(n192) );
  NAND2X0_HVT U209 ( .A1(n490), .A2(n515), .Y(n203) );
  NAND2X0_HVT U210 ( .A1(n194), .A2(n198), .Y(n205) );
  NAND2X0_HVT U211 ( .A1(n203), .A2(n205), .Y(out[44]) );
  INVX0_HVT U212 ( .A(n490), .Y(n194) );
  INVX1_HVT U213 ( .A(n515), .Y(n198) );
  XOR2X2_HVT U214 ( .A1(in[10]), .A2(n546), .Y(n210) );
  XNOR2X2_HVT U215 ( .A1(n36), .A2(n213), .Y(out[91]) );
  INVX2_HVT U216 ( .A(in[87]), .Y(n580) );
  NBUFFX2_HVT U217 ( .A(in[23]), .Y(n214) );
  INVX0_HVT U218 ( .A(n510), .Y(n216) );
  XOR2X2_HVT U219 ( .A1(in[17]), .A2(in[25]), .Y(n16) );
  XOR3X2_HVT U220 ( .A1(n464), .A2(in[19]), .A3(n154), .Y(n153) );
  XOR2X2_HVT U221 ( .A1(in[12]), .A2(in[20]), .Y(n118) );
  INVX2_HVT U222 ( .A(in[19]), .Y(n509) );
  XOR3X2_HVT U223 ( .A1(n509), .A2(n544), .A3(n216), .Y(n195) );
  INVX1_HVT U224 ( .A(n544), .Y(n454) );
  INVX1_HVT U226 ( .A(in[120]), .Y(n220) );
  INVX2_HVT U227 ( .A(n220), .Y(n222) );
  XNOR2X2_HVT U228 ( .A1(n223), .A2(n471), .Y(n334) );
  IBUFFX16_HVT U229 ( .A(n566), .Y(n223) );
  INVX1_HVT U230 ( .A(in[61]), .Y(n356) );
  XOR2X1_HVT U231 ( .A1(in[61]), .A2(n242), .Y(n138) );
  IBUFFX2_HVT U232 ( .A(n567), .Y(n238) );
  INVX0_HVT U233 ( .A(in[110]), .Y(n231) );
  XOR3X2_HVT U234 ( .A1(n224), .A2(n355), .A3(n147), .Y(out[22]) );
  XNOR2X1_HVT U235 ( .A1(in[30]), .A2(in[21]), .Y(n224) );
  INVX1_HVT U236 ( .A(n124), .Y(n574) );
  XNOR2X1_HVT U237 ( .A1(in[10]), .A2(in[2]), .Y(n158) );
  INVX1_HVT U238 ( .A(in[124]), .Y(n339) );
  XOR2X2_HVT U239 ( .A1(in[100]), .A2(in[124]), .Y(n202) );
  XOR2X2_HVT U240 ( .A1(in[116]), .A2(in[124]), .Y(n181) );
  XOR3X2_HVT U241 ( .A1(n21), .A2(n193), .A3(n225), .Y(out[113]) );
  XOR3X2_HVT U242 ( .A1(n568), .A2(n265), .A3(in[104]), .Y(n225) );
  INVX1_HVT U243 ( .A(n180), .Y(n310) );
  XOR3X1_HVT U244 ( .A1(n78), .A2(n462), .A3(n150), .Y(out[14]) );
  XNOR2X2_HVT U245 ( .A1(in[30]), .A2(in[22]), .Y(n78) );
  INVX0_HVT U246 ( .A(in[13]), .Y(n355) );
  XOR3X2_HVT U247 ( .A1(n178), .A2(n227), .A3(n209), .Y(out[111]) );
  IBUFFX16_HVT U248 ( .A(n572), .Y(n227) );
  XOR2X2_HVT U249 ( .A1(in[3]), .A2(n549), .Y(n157) );
  INVX0_HVT U250 ( .A(in[21]), .Y(n368) );
  XOR3X2_HVT U251 ( .A1(n159), .A2(n228), .A3(n538), .Y(out[0]) );
  XOR2X2_HVT U252 ( .A1(in[113]), .A2(in[121]), .Y(n189) );
  XOR3X2_HVT U253 ( .A1(n524), .A2(n520), .A3(n35), .Y(n34) );
  XOR2X2_HVT U254 ( .A1(in[76]), .A2(in[68]), .Y(n35) );
  XNOR2X2_HVT U255 ( .A1(n431), .A2(n229), .Y(out[107]) );
  XOR2X1_HVT U256 ( .A1(in[8]), .A2(n551), .Y(n162) );
  NBUFFX2_HVT U257 ( .A(in[16]), .Y(n230) );
  XOR2X2_HVT U258 ( .A1(n222), .A2(n569), .Y(n27) );
  XOR2X2_HVT U259 ( .A1(in[46]), .A2(in[38]), .Y(n87) );
  XNOR2X1_HVT U260 ( .A1(in[40]), .A2(n573), .Y(n145) );
  XOR3X2_HVT U261 ( .A1(n177), .A2(n231), .A3(n197), .Y(out[119]) );
  INVX0_HVT U262 ( .A(in[57]), .Y(n279) );
  XOR3X2_HVT U263 ( .A1(n46), .A2(n232), .A3(n47), .Y(out[88]) );
  IBUFFX16_HVT U264 ( .A(n584), .Y(n232) );
  INVX0_HVT U265 ( .A(in[0]), .Y(n246) );
  XOR3X2_HVT U266 ( .A1(n26), .A2(n233), .A3(n27), .Y(out[96]) );
  IBUFFX16_HVT U267 ( .A(n572), .Y(n233) );
  XNOR2X2_HVT U268 ( .A1(in[113]), .A2(in[105]), .Y(n24) );
  INVX0_HVT U269 ( .A(in[113]), .Y(n336) );
  INVX1_HVT U270 ( .A(n375), .Y(n376) );
  INVX1_HVT U271 ( .A(in[73]), .Y(n294) );
  XOR3X2_HVT U272 ( .A1(n162), .A2(n234), .A3(n163), .Y(out[24]) );
  IBUFFX16_HVT U273 ( .A(n577), .Y(n234) );
  INVX1_HVT U274 ( .A(n575), .Y(n254) );
  XOR3X2_HVT U275 ( .A1(n168), .A2(n235), .A3(n158), .Y(out[18]) );
  XOR3X2_HVT U276 ( .A1(n145), .A2(n236), .A3(n101), .Y(out[32]) );
  XNOR2X1_HVT U277 ( .A1(n568), .A2(n583), .Y(n404) );
  INVX0_HVT U278 ( .A(in[54]), .Y(n257) );
  XOR3X2_HVT U279 ( .A1(n217), .A2(n238), .A3(n23), .Y(out[104]) );
  IBUFFX16_HVT U280 ( .A(n460), .Y(n239) );
  XOR2X2_HVT U281 ( .A1(n61), .A2(n432), .Y(n240) );
  XOR2X2_HVT U282 ( .A1(n60), .A2(n240), .Y(out[80]) );
  XNOR2X1_HVT U283 ( .A1(in[88]), .A2(n580), .Y(n60) );
  IBUFFX2_HVT U284 ( .A(n584), .Y(n432) );
  XOR2X2_HVT U285 ( .A1(in[86]), .A2(in[94]), .Y(n65) );
  INVX2_HVT U286 ( .A(n555), .Y(n358) );
  INVX0_HVT U287 ( .A(in[42]), .Y(n375) );
  INVX0_HVT U288 ( .A(in[41]), .Y(n402) );
  XOR2X2_HVT U289 ( .A1(in[84]), .A2(in[92]), .Y(n32) );
  INVX0_HVT U290 ( .A(in[46]), .Y(n241) );
  INVX1_HVT U291 ( .A(n241), .Y(n242) );
  INVX1_HVT U292 ( .A(n289), .Y(n293) );
  INVX0_HVT U293 ( .A(n87), .Y(n289) );
  XOR3X1_HVT U294 ( .A1(n99), .A2(n263), .A3(n338), .Y(out[50]) );
  XNOR2X2_HVT U295 ( .A1(n243), .A2(n153), .Y(out[28]) );
  INVX0_HVT U296 ( .A(n492), .Y(n255) );
  INVX1_HVT U297 ( .A(n298), .Y(n244) );
  XOR3X2_HVT U298 ( .A1(n245), .A2(n553), .A3(n133), .Y(out[40]) );
  XNOR2X1_HVT U299 ( .A1(in[56]), .A2(n573), .Y(n245) );
  INVX0_HVT U300 ( .A(in[84]), .Y(n524) );
  XOR3X2_HVT U301 ( .A1(n541), .A2(n246), .A3(in[1]), .Y(n17) );
  INVX1_HVT U302 ( .A(n35), .Y(n247) );
  INVX1_HVT U303 ( .A(n247), .Y(n248) );
  NBUFFX2_HVT U304 ( .A(n543), .Y(n249) );
  INVX0_HVT U305 ( .A(in[98]), .Y(n250) );
  INVX1_HVT U306 ( .A(n250), .Y(n251) );
  NAND2X0_HVT U307 ( .A1(n556), .A2(n257), .Y(n258) );
  NAND2X0_HVT U308 ( .A1(n256), .A2(in[54]), .Y(n259) );
  NAND2X0_HVT U309 ( .A1(n259), .A2(n258), .Y(n106) );
  INVX1_HVT U310 ( .A(n556), .Y(n256) );
  XNOR2X2_HVT U311 ( .A1(n406), .A2(n498), .Y(n204) );
  INVX0_HVT U312 ( .A(in[79]), .Y(n260) );
  INVX0_HVT U313 ( .A(n260), .Y(n261) );
  INVX1_HVT U314 ( .A(in[58]), .Y(n262) );
  INVX1_HVT U315 ( .A(n262), .Y(n263) );
  XOR2X1_HVT U316 ( .A1(in[50]), .A2(in[58]), .Y(n130) );
  INVX1_HVT U317 ( .A(in[105]), .Y(n264) );
  INVX2_HVT U318 ( .A(in[48]), .Y(n573) );
  INVX2_HVT U319 ( .A(n438), .Y(n460) );
  XOR2X2_HVT U320 ( .A1(in[49]), .A2(n280), .Y(n100) );
  XOR2X2_HVT U321 ( .A1(n473), .A2(n493), .Y(n129) );
  XOR2X1_HVT U322 ( .A1(n557), .A2(n319), .Y(n104) );
  XOR3X2_HVT U323 ( .A1(n266), .A2(n299), .A3(n52), .Y(out[10]) );
  IBUFFX2_HVT U324 ( .A(in[67]), .Y(n394) );
  INVX0_HVT U325 ( .A(n518), .Y(n300) );
  NBUFFX2_HVT U326 ( .A(in[95]), .Y(n564) );
  XOR2X1_HVT U327 ( .A1(n558), .A2(in[59]), .Y(n143) );
  INVX0_HVT U328 ( .A(in[88]), .Y(n297) );
  INVX0_HVT U329 ( .A(n202), .Y(n301) );
  INVX1_HVT U330 ( .A(n387), .Y(n388) );
  INVX1_HVT U331 ( .A(in[67]), .Y(n438) );
  INVX0_HVT U332 ( .A(n424), .Y(n351) );
  XOR2X1_HVT U333 ( .A1(n542), .A2(n550), .Y(n136) );
  INVX0_HVT U334 ( .A(in[116]), .Y(n369) );
  INVX1_HVT U335 ( .A(in[112]), .Y(n582) );
  INVX1_HVT U336 ( .A(n505), .Y(n506) );
  INVX0_HVT U337 ( .A(n573), .Y(n379) );
  INVX0_HVT U338 ( .A(n89), .Y(n286) );
  INVX1_HVT U339 ( .A(n119), .Y(n377) );
  XOR2X1_HVT U340 ( .A1(n428), .A2(in[27]), .Y(n172) );
  INVX1_HVT U341 ( .A(in[24]), .Y(n344) );
  XNOR2X1_HVT U342 ( .A1(n5), .A2(n541), .Y(n538) );
  INVX1_HVT U343 ( .A(n546), .Y(n381) );
  INVX1_HVT U344 ( .A(in[107]), .Y(n274) );
  INVX1_HVT U345 ( .A(in[14]), .Y(n507) );
  INVX1_HVT U346 ( .A(n497), .Y(n572) );
  INVX1_HVT U347 ( .A(in[43]), .Y(n353) );
  XOR2X2_HVT U348 ( .A1(in[88]), .A2(n566), .Y(n268) );
  XOR2X2_HVT U349 ( .A1(n558), .A2(n254), .Y(n270) );
  XNOR2X2_HVT U350 ( .A1(in[0]), .A2(n542), .Y(n271) );
  INVX1_HVT U351 ( .A(in[59]), .Y(n357) );
  XOR2X2_HVT U352 ( .A1(n472), .A2(n563), .Y(n272) );
  INVX1_HVT U353 ( .A(in[64]), .Y(n584) );
  INVX1_HVT U354 ( .A(n552), .Y(n495) );
  XNOR2X2_HVT U355 ( .A1(in[118]), .A2(in[126]), .Y(n273) );
  INVX1_HVT U356 ( .A(in[122]), .Y(n307) );
  INVX0_HVT U357 ( .A(n201), .Y(n467) );
  INVX1_HVT U358 ( .A(in[75]), .Y(n387) );
  NAND2X0_HVT U359 ( .A1(n123), .A2(n325), .Y(n277) );
  NAND2X0_HVT U360 ( .A1(n275), .A2(n276), .Y(n278) );
  NAND2X0_HVT U361 ( .A1(n277), .A2(n278), .Y(out[47]) );
  INVX0_HVT U362 ( .A(n123), .Y(n275) );
  INVX0_HVT U363 ( .A(n325), .Y(n276) );
  XNOR2X2_HVT U364 ( .A1(n272), .A2(n295), .Y(n324) );
  INVX1_HVT U365 ( .A(n420), .Y(n319) );
  INVX1_HVT U366 ( .A(n279), .Y(n280) );
  XOR2X2_HVT U367 ( .A1(in[93]), .A2(in[78]), .Y(n76) );
  XOR3X2_HVT U368 ( .A1(n495), .A2(n7), .A3(n108), .Y(n140) );
  XOR3X2_HVT U369 ( .A1(n7), .A2(n458), .A3(n90), .Y(n515) );
  XOR3X2_HVT U370 ( .A1(n27), .A2(n190), .A3(n281), .Y(out[121]) );
  XOR3X2_HVT U371 ( .A1(n532), .A2(n337), .A3(n582), .Y(n281) );
  XOR2X1_HVT U372 ( .A1(n251), .A2(in[106]), .Y(n188) );
  INVX0_HVT U373 ( .A(n74), .Y(n408) );
  INVX1_HVT U374 ( .A(n130), .Y(n322) );
  XOR2X2_HVT U375 ( .A1(in[108]), .A2(in[100]), .Y(n184) );
  XOR3X2_HVT U376 ( .A1(n115), .A2(n401), .A3(n144), .Y(out[33]) );
  INVX0_HVT U377 ( .A(n115), .Y(n338) );
  NAND2X0_HVT U378 ( .A1(n54), .A2(n283), .Y(n284) );
  NAND2X0_HVT U379 ( .A1(n282), .A2(n419), .Y(n285) );
  NAND2X0_HVT U380 ( .A1(n284), .A2(n285), .Y(out[83]) );
  INVX0_HVT U381 ( .A(n54), .Y(n282) );
  INVX0_HVT U382 ( .A(n419), .Y(n283) );
  INVX1_HVT U383 ( .A(in[74]), .Y(n505) );
  XNOR2X2_HVT U384 ( .A1(in[87]), .A2(n564), .Y(n64) );
  XNOR2X2_HVT U385 ( .A1(n294), .A2(in[81]), .Y(n57) );
  INVX1_HVT U386 ( .A(n150), .Y(n372) );
  INVX1_HVT U387 ( .A(n286), .Y(n287) );
  XOR3X2_HVT U388 ( .A1(n23), .A2(n24), .A3(n288), .Y(out[97]) );
  XOR3X2_HVT U389 ( .A1(in[121]), .A2(n222), .A3(n569), .Y(n288) );
  NAND2X0_HVT U390 ( .A1(n293), .A2(n495), .Y(n291) );
  NAND2X0_HVT U391 ( .A1(n289), .A2(n290), .Y(n292) );
  NAND2X0_HVT U392 ( .A1(n291), .A2(n292), .Y(n325) );
  INVX1_HVT U393 ( .A(n294), .Y(n295) );
  XOR3X2_HVT U394 ( .A1(n443), .A2(n29), .A3(n296), .Y(out[86]) );
  XNOR2X2_HVT U395 ( .A1(n575), .A2(in[48]), .Y(n105) );
  INVX1_HVT U396 ( .A(in[68]), .Y(n534) );
  INVX0_HVT U397 ( .A(in[43]), .Y(n513) );
  XOR3X2_HVT U398 ( .A1(n566), .A2(n305), .A3(n297), .Y(n441) );
  INVX1_HVT U399 ( .A(n305), .Y(n306) );
  XOR3X2_HVT U400 ( .A1(n47), .A2(n58), .A3(n324), .Y(out[81]) );
  INVX0_HVT U401 ( .A(n532), .Y(n374) );
  INVX0_HVT U402 ( .A(n90), .Y(n321) );
  INVX1_HVT U403 ( .A(n394), .Y(n326) );
  INVX1_HVT U404 ( .A(in[2]), .Y(n298) );
  INVX1_HVT U405 ( .A(n298), .Y(n299) );
  INVX1_HVT U406 ( .A(n30), .Y(n418) );
  XOR3X2_HVT U407 ( .A1(n564), .A2(n424), .A3(n300), .Y(n349) );
  INVX1_HVT U408 ( .A(in[91]), .Y(n424) );
  IBUFFX2_HVT U409 ( .A(in[93]), .Y(n440) );
  XOR2X1_HVT U410 ( .A1(in[52]), .A2(in[60]), .Y(n90) );
  XOR3X1_HVT U411 ( .A1(n465), .A2(n307), .A3(n308), .Y(n413) );
  XOR2X2_HVT U412 ( .A1(n434), .A2(n570), .Y(n416) );
  INVX2_HVT U413 ( .A(n433), .Y(n434) );
  INVX0_HVT U414 ( .A(n242), .Y(n447) );
  XOR3X2_HVT U415 ( .A1(n579), .A2(n303), .A3(n28), .Y(out[95]) );
  XOR3X2_HVT U416 ( .A1(n180), .A2(n421), .A3(n273), .Y(out[110]) );
  XOR3X2_HVT U417 ( .A1(n169), .A2(n271), .A3(n168), .Y(out[1]) );
  IBUFFX2_HVT U418 ( .A(in[54]), .Y(n456) );
  INVX0_HVT U419 ( .A(n359), .Y(n302) );
  INVX1_HVT U420 ( .A(n69), .Y(n328) );
  XOR3X2_HVT U421 ( .A1(n303), .A2(in[81]), .A3(n578), .Y(n45) );
  INVX0_HVT U422 ( .A(n267), .Y(n304) );
  INVX0_HVT U423 ( .A(n472), .Y(n380) );
  XNOR2X1_HVT U424 ( .A1(in[30]), .A2(in[6]), .Y(n343) );
  XNOR2X2_HVT U425 ( .A1(in[14]), .A2(n462), .Y(n147) );
  XOR3X2_HVT U426 ( .A1(n452), .A2(n513), .A3(n111), .Y(n461) );
  XOR3X2_HVT U427 ( .A1(n340), .A2(n309), .A3(n310), .Y(out[117]) );
  NBUFFX2_HVT U428 ( .A(in[33]), .Y(n311) );
  NAND2X0_HVT U429 ( .A1(n519), .A2(n502), .Y(n313) );
  NAND2X0_HVT U430 ( .A1(n312), .A2(n51), .Y(n314) );
  NAND2X0_HVT U431 ( .A1(n313), .A2(n314), .Y(n81) );
  INVX0_HVT U432 ( .A(n519), .Y(n312) );
  NAND2X0_HVT U433 ( .A1(n83), .A2(in[90]), .Y(n316) );
  NAND2X0_HVT U434 ( .A1(n315), .A2(n409), .Y(n317) );
  NAND2X0_HVT U435 ( .A1(n316), .A2(n317), .Y(n519) );
  XNOR2X1_HVT U436 ( .A1(n357), .A2(n575), .Y(n385) );
  INVX1_HVT U437 ( .A(in[40]), .Y(n420) );
  XNOR2X2_HVT U438 ( .A1(in[74]), .A2(in[66]), .Y(n39) );
  INVX1_HVT U439 ( .A(in[51]), .Y(n492) );
  NBUFFX2_HVT U440 ( .A(in[9]), .Y(n320) );
  XOR2X2_HVT U441 ( .A1(in[1]), .A2(n320), .Y(n160) );
  XOR3X2_HVT U442 ( .A1(n377), .A2(n376), .A3(n322), .Y(out[34]) );
  XNOR2X2_HVT U443 ( .A1(in[77]), .A2(in[69]), .Y(n31) );
  IBUFFX2_HVT U444 ( .A(in[69]), .Y(n470) );
  INVX1_HVT U445 ( .A(n353), .Y(n333) );
  XOR3X2_HVT U446 ( .A1(n65), .A2(n422), .A3(n31), .Y(out[78]) );
  NBUFFX2_HVT U447 ( .A(in[103]), .Y(n497) );
  XOR3X2_HVT U448 ( .A1(n178), .A2(n342), .A3(n179), .Y(out[126]) );
  XNOR2X2_HVT U449 ( .A1(n345), .A2(in[125]), .Y(n179) );
  NBUFFX2_HVT U450 ( .A(in[27]), .Y(n323) );
  XOR3X2_HVT U451 ( .A1(n15), .A2(n508), .A3(n17), .Y(out[9]) );
  XOR3X2_HVT U452 ( .A1(n388), .A2(n505), .A3(n326), .Y(n419) );
  NAND2X0_HVT U453 ( .A1(n527), .A2(n69), .Y(n329) );
  NAND2X0_HVT U454 ( .A1(n327), .A2(n328), .Y(n330) );
  NAND2X0_HVT U455 ( .A1(n330), .A2(n329), .Y(out[75]) );
  IBUFFX2_HVT U456 ( .A(in[109]), .Y(n500) );
  XNOR3X1_HVT U457 ( .A1(n181), .A2(n345), .A3(n180), .Y(out[125]) );
  INVX1_HVT U458 ( .A(n331), .Y(n332) );
  XOR3X2_HVT U459 ( .A1(n555), .A2(n333), .A3(n495), .Y(n490) );
  INVX0_HVT U460 ( .A(in[44]), .Y(n451) );
  XOR2X2_HVT U461 ( .A1(in[36]), .A2(in[44]), .Y(n93) );
  XOR2X2_HVT U462 ( .A1(in[94]), .A2(n562), .Y(n75) );
  INVX1_HVT U463 ( .A(n513), .Y(n347) );
  XOR3X2_HVT U464 ( .A1(n28), .A2(in[78]), .A3(n334), .Y(out[87]) );
  XNOR2X2_HVT U465 ( .A1(n404), .A2(in[115]), .Y(n200) );
  XNOR2X2_HVT U466 ( .A1(n335), .A2(n183), .Y(out[124]) );
  XOR3X2_HVT U467 ( .A1(n570), .A2(in[123]), .A3(n435), .Y(n335) );
  INVX1_HVT U468 ( .A(n336), .Y(n337) );
  XOR3X2_HVT U469 ( .A1(n529), .A2(n571), .A3(n339), .Y(n450) );
  IBUFFX2_HVT U470 ( .A(in[118]), .Y(n341) );
  INVX1_HVT U471 ( .A(n341), .Y(n342) );
  XOR3X2_HVT U472 ( .A1(n147), .A2(n249), .A3(n405), .Y(out[15]) );
  XOR3X2_HVT U473 ( .A1(n343), .A2(n546), .A3(n63), .Y(out[7]) );
  XOR3X2_HVT U474 ( .A1(n549), .A2(n344), .A3(n332), .Y(n169) );
  NBUFFX2_HVT U475 ( .A(in[117]), .Y(n345) );
  XOR3X2_HVT U476 ( .A1(n94), .A2(n346), .A3(n147), .Y(out[30]) );
  XNOR2X2_HVT U477 ( .A1(in[41]), .A2(in[33]), .Y(n102) );
  XOR3X2_HVT U478 ( .A1(n347), .A2(n376), .A3(n7), .Y(n393) );
  NBUFFX2_HVT U479 ( .A(n124), .Y(n348) );
  XOR3X2_HVT U480 ( .A1(n384), .A2(n412), .A3(n479), .Y(n167) );
  XOR3X2_HVT U481 ( .A1(n78), .A2(n350), .A3(n146), .Y(out[31]) );
  XOR2X2_HVT U482 ( .A1(in[1]), .A2(in[25]), .Y(n148) );
  XNOR2X1_HVT U483 ( .A1(n494), .A2(n557), .Y(n123) );
  XNOR2X2_HVT U484 ( .A1(n222), .A2(n582), .Y(n217) );
  XNOR2X2_HVT U485 ( .A1(n354), .A2(n186), .Y(out[123]) );
  XOR3X2_HVT U486 ( .A1(in[122]), .A2(n435), .A3(n187), .Y(n354) );
  XOR3X2_HVT U487 ( .A1(n64), .A2(n410), .A3(n29), .Y(out[79]) );
  NBUFFX2_HVT U488 ( .A(in[47]), .Y(n555) );
  XOR3X2_HVT U489 ( .A1(n108), .A2(n356), .A3(n287), .Y(out[53]) );
  XNOR2X2_HVT U490 ( .A1(n290), .A2(n554), .Y(n86) );
  XOR3X2_HVT U491 ( .A1(n559), .A2(n584), .A3(in[65]), .Y(n72) );
  NBUFFX2_HVT U492 ( .A(in[95]), .Y(n565) );
  XOR3X2_HVT U493 ( .A1(n494), .A2(n492), .A3(n358), .Y(n491) );
  INVX1_HVT U494 ( .A(n492), .Y(n493) );
  IBUFFX2_HVT U495 ( .A(in[29]), .Y(n359) );
  INVX1_HVT U496 ( .A(n359), .Y(n360) );
  XOR2X2_HVT U497 ( .A1(n386), .A2(n556), .Y(n101) );
  NAND2X0_HVT U498 ( .A1(n530), .A2(n504), .Y(n362) );
  NAND2X0_HVT U499 ( .A1(n361), .A2(n251), .Y(n363) );
  NAND2X0_HVT U500 ( .A1(n362), .A2(n363), .Y(n215) );
  IBUFFX2_HVT U501 ( .A(n530), .Y(n361) );
  NBUFFX2_HVT U502 ( .A(in[71]), .Y(n559) );
  XNOR2X2_HVT U503 ( .A1(n364), .A2(n365), .Y(out[43]) );
  XOR3X1_HVT U504 ( .A1(n553), .A2(n375), .A3(n129), .Y(n364) );
  XNOR2X2_HVT U505 ( .A1(n96), .A2(n366), .Y(out[59]) );
  XOR3X2_HVT U506 ( .A1(n367), .A2(n542), .A3(n429), .Y(n116) );
  XOR3X2_HVT U507 ( .A1(n369), .A2(in[115]), .A3(n184), .Y(n183) );
  XOR3X2_HVT U508 ( .A1(in[76]), .A2(n371), .A3(n53), .Y(n370) );
  INVX1_HVT U509 ( .A(n387), .Y(n371) );
  XNOR2X2_HVT U510 ( .A1(n550), .A2(n10), .Y(n539) );
  NBUFFX2_HVT U511 ( .A(in[5]), .Y(n373) );
  XOR3X2_HVT U512 ( .A1(n273), .A2(n374), .A3(n177), .Y(out[127]) );
  XOR3X2_HVT U513 ( .A1(n86), .A2(n494), .A3(n574), .Y(out[63]) );
  XNOR2X2_HVT U514 ( .A1(n391), .A2(in[61]), .Y(n88) );
  INVX0_HVT U515 ( .A(n562), .Y(n378) );
  XOR3X2_HVT U516 ( .A1(n561), .A2(n387), .A3(n560), .Y(n66) );
  XOR3X2_HVT U517 ( .A1(n382), .A2(n501), .A3(n178), .Y(out[118]) );
  XNOR2X1_HVT U518 ( .A1(in[117]), .A2(in[126]), .Y(n382) );
  XOR3X2_HVT U519 ( .A1(n160), .A2(n159), .A3(n383), .Y(out[25]) );
  XOR3X2_HVT U520 ( .A1(n214), .A2(n230), .A3(in[17]), .Y(n383) );
  XOR3X2_HVT U521 ( .A1(n352), .A2(n358), .A3(n385), .Y(n392) );
  XOR3X2_HVT U522 ( .A1(n540), .A2(n474), .A3(n293), .Y(out[54]) );
  XOR3X2_HVT U523 ( .A1(n557), .A2(n386), .A3(n280), .Y(n144) );
  NBUFFX2_HVT U524 ( .A(in[79]), .Y(n561) );
  XOR3X2_HVT U525 ( .A1(n518), .A2(n51), .A3(n563), .Y(n389) );
  XOR3X2_HVT U526 ( .A1(n101), .A2(n102), .A3(n390), .Y(out[57]) );
  XOR3X2_HVT U527 ( .A1(n72), .A2(n61), .A3(n267), .Y(out[73]) );
  XNOR2X2_HVT U528 ( .A1(n392), .A2(n393), .Y(out[51]) );
  NAND2X0_HVT U529 ( .A1(n91), .A2(n396), .Y(n397) );
  NAND2X0_HVT U530 ( .A1(n395), .A2(n92), .Y(n398) );
  NAND2X0_HVT U531 ( .A1(n397), .A2(n398), .Y(out[60]) );
  INVX1_HVT U532 ( .A(n91), .Y(n395) );
  INVX0_HVT U533 ( .A(n92), .Y(n396) );
  XNOR2X2_HVT U534 ( .A1(n270), .A2(n473), .Y(n91) );
  XNOR2X2_HVT U535 ( .A1(n559), .A2(n563), .Y(n28) );
  XOR3X2_HVT U536 ( .A1(n554), .A2(n319), .A3(n403), .Y(n400) );
  INVX1_HVT U537 ( .A(n402), .Y(n403) );
  XOR2X2_HVT U538 ( .A1(in[49]), .A2(n403), .Y(n115) );
  INVX0_HVT U539 ( .A(in[104]), .Y(n414) );
  INVX0_HVT U540 ( .A(in[115]), .Y(n526) );
  INVX0_HVT U541 ( .A(n193), .Y(n415) );
  INVX1_HVT U542 ( .A(in[66]), .Y(n514) );
  XOR3X1_HVT U543 ( .A1(n560), .A2(n438), .A3(n50), .Y(n80) );
  INVX1_HVT U544 ( .A(in[6]), .Y(n462) );
  XNOR2X1_HVT U545 ( .A1(n576), .A2(in[16]), .Y(n455) );
  INVX0_HVT U546 ( .A(n551), .Y(n429) );
  INVX0_HVT U547 ( .A(n517), .Y(n417) );
  INVX0_HVT U548 ( .A(n581), .Y(n444) );
  INVX0_HVT U549 ( .A(n577), .Y(n446) );
  INVX0_HVT U550 ( .A(n94), .Y(n436) );
  INVX1_HVT U551 ( .A(in[18]), .Y(n523) );
  INVX0_HVT U552 ( .A(in[100]), .Y(n487) );
  XOR2X2_HVT U553 ( .A1(n547), .A2(n551), .Y(n405) );
  INVX1_HVT U554 ( .A(n532), .Y(n435) );
  XOR2X2_HVT U555 ( .A1(n568), .A2(in[106]), .Y(n406) );
  INVX0_HVT U556 ( .A(in[38]), .Y(n437) );
  INVX1_HVT U557 ( .A(in[83]), .Y(n502) );
  INVX1_HVT U558 ( .A(n560), .Y(n410) );
  INVX0_HVT U559 ( .A(in[70]), .Y(n422) );
  XOR3X2_HVT U560 ( .A1(n118), .A2(n360), .A3(n150), .Y(out[21]) );
  NAND2X0_HVT U561 ( .A1(n484), .A2(n381), .Y(n407) );
  XOR3X2_HVT U562 ( .A1(n39), .A2(n409), .A3(n57), .Y(out[82]) );
  XOR3X2_HVT U563 ( .A1(n149), .A2(n510), .A3(n148), .Y(out[2]) );
  XNOR2X2_HVT U564 ( .A1(in[65]), .A2(in[73]), .Y(n44) );
  XOR3X2_HVT U565 ( .A1(n411), .A2(n410), .A3(n268), .Y(out[64]) );
  XOR3X2_HVT U566 ( .A1(n78), .A2(n507), .A3(n77), .Y(out[6]) );
  XNOR2X2_HVT U567 ( .A1(n413), .A2(n19), .Y(out[99]) );
  XOR3X2_HVT U568 ( .A1(n16), .A2(n523), .A3(n158), .Y(out[26]) );
  XOR3X2_HVT U569 ( .A1(n416), .A2(n414), .A3(n415), .Y(out[120]) );
  XOR3X2_HVT U570 ( .A1(n22), .A2(n417), .A3(n21), .Y(out[98]) );
  XOR3X2_HVT U571 ( .A1(n248), .A2(n430), .A3(n418), .Y(out[77]) );
  IBUFFX2_HVT U572 ( .A(in[37]), .Y(n449) );
  XNOR2X2_HVT U573 ( .A1(n420), .A2(n553), .Y(n122) );
  INVX1_HVT U574 ( .A(n499), .Y(n421) );
  INVX1_HVT U575 ( .A(in[102]), .Y(n499) );
  XOR3X2_HVT U576 ( .A1(n64), .A2(n422), .A3(n75), .Y(out[71]) );
  XOR3X2_HVT U577 ( .A1(n189), .A2(n208), .A3(n425), .Y(out[105]) );
  XOR3X2_HVT U578 ( .A1(in[97]), .A2(n434), .A3(n497), .Y(n425) );
  XNOR2X2_HVT U579 ( .A1(in[85]), .A2(in[93]), .Y(n30) );
  XOR3X2_HVT U580 ( .A1(n31), .A2(n426), .A3(n32), .Y(out[93]) );
  INVX1_HVT U581 ( .A(n427), .Y(n428) );
  INVX1_HVT U582 ( .A(n470), .Y(n430) );
  XOR2X2_HVT U583 ( .A1(n565), .A2(n380), .Y(n46) );
  XNOR2X1_HVT U584 ( .A1(in[114]), .A2(in[122]), .Y(n22) );
  INVX1_HVT U585 ( .A(in[96]), .Y(n433) );
  XOR3X2_HVT U586 ( .A1(n207), .A2(n435), .A3(n208), .Y(out[112]) );
  XOR3X2_HVT U587 ( .A1(n436), .A2(n373), .A3(n154), .Y(out[13]) );
  XNOR2X1_HVT U588 ( .A1(n386), .A2(in[55]), .Y(n121) );
  XOR3X2_HVT U589 ( .A1(n137), .A2(n437), .A3(n123), .Y(out[39]) );
  XOR3X2_HVT U590 ( .A1(n202), .A2(n500), .A3(n179), .Y(out[101]) );
  XOR3X2_HVT U591 ( .A1(n273), .A2(n439), .A3(n219), .Y(out[102]) );
  XOR3X2_HVT U592 ( .A1(n31), .A2(n440), .A3(n50), .Y(out[85]) );
  XOR3X2_HVT U593 ( .A1(n57), .A2(n74), .A3(n441), .Y(out[65]) );
  XNOR2X2_HVT U594 ( .A1(n434), .A2(n496), .Y(n23) );
  XOR3X2_HVT U595 ( .A1(n442), .A2(n122), .A3(n100), .Y(out[41]) );
  XOR3X2_HVT U596 ( .A1(in[33]), .A2(in[32]), .A3(n290), .Y(n442) );
  INVX0_HVT U597 ( .A(n459), .Y(n443) );
  IBUFFX2_HVT U598 ( .A(in[45]), .Y(n474) );
  XOR3X2_HVT U599 ( .A1(n121), .A2(n444), .A3(n122), .Y(out[48]) );
  XNOR2X2_HVT U600 ( .A1(n81), .A2(n445), .Y(out[67]) );
  XOR3X2_HVT U601 ( .A1(n388), .A2(n559), .A3(n457), .Y(n445) );
  XOR3X2_HVT U602 ( .A1(n174), .A2(n446), .A3(n15), .Y(out[16]) );
  XOR3X2_HVT U603 ( .A1(n106), .A2(n447), .A3(n86), .Y(out[55]) );
  NBUFFX2_HVT U604 ( .A(in[7]), .Y(n541) );
  NBUFFX2_HVT U605 ( .A(in[47]), .Y(n554) );
  XOR2X2_HVT U606 ( .A1(n230), .A2(n548), .Y(n163) );
  XOR3X2_HVT U607 ( .A1(n138), .A2(n449), .A3(n574), .Y(out[38]) );
  IBUFFX2_HVT U608 ( .A(in[20]), .Y(n464) );
  INVX1_HVT U609 ( .A(n16), .Y(n508) );
  XNOR2X2_HVT U610 ( .A1(n221), .A2(n450), .Y(out[100]) );
  NBUFFX2_HVT U611 ( .A(in[103]), .Y(n496) );
  INVX1_HVT U612 ( .A(n451), .Y(n452) );
  NBUFFX2_HVT U613 ( .A(in[26]), .Y(n453) );
  XOR3X2_HVT U614 ( .A1(n455), .A2(n454), .A3(n271), .Y(out[8]) );
  XOR3X2_HVT U615 ( .A1(n87), .A2(n456), .A3(n88), .Y(out[62]) );
  XOR3X2_HVT U616 ( .A1(n93), .A2(n449), .A3(n88), .Y(out[45]) );
  INVX1_HVT U617 ( .A(n514), .Y(n457) );
  XNOR2X2_HVT U618 ( .A1(in[18]), .A2(in[26]), .Y(n149) );
  XOR3X2_HVT U619 ( .A1(n556), .A2(n476), .A3(n473), .Y(n463) );
  NAND2X0_HVT U620 ( .A1(n200), .A2(n467), .Y(n468) );
  NAND2X0_HVT U621 ( .A1(n466), .A2(n201), .Y(n469) );
  NAND2X0_HVT U622 ( .A1(n468), .A2(n469), .Y(out[116]) );
  INVX0_HVT U623 ( .A(n200), .Y(n466) );
  XOR3X2_HVT U624 ( .A1(n509), .A2(n523), .A3(n522), .Y(n477) );
  XOR2X2_HVT U625 ( .A1(n565), .A2(in[91]), .Y(n83) );
  XOR3X2_HVT U626 ( .A1(n76), .A2(n470), .A3(n579), .Y(out[70]) );
  XOR3X2_HVT U627 ( .A1(n29), .A2(n471), .A3(n30), .Y(out[94]) );
  XOR3X2_HVT U628 ( .A1(n111), .A2(n474), .A3(n88), .Y(out[37]) );
  AND2X1_HVT U629 ( .A1(n485), .A2(in[11]), .Y(n475) );
  NBUFFX2_HVT U630 ( .A(in[60]), .Y(n476) );
  INVX0_HVT U631 ( .A(n479), .Y(n95) );
  XNOR2X2_HVT U632 ( .A1(n155), .A2(n477), .Y(out[27]) );
  XOR3X2_HVT U633 ( .A1(n299), .A2(n323), .A3(n136), .Y(n478) );
  NAND2X0_HVT U634 ( .A1(n536), .A2(n412), .Y(n481) );
  NAND2X0_HVT U635 ( .A1(n475), .A2(n407), .Y(n482) );
  NAND2X0_HVT U636 ( .A1(n481), .A2(n482), .Y(n176) );
  XOR3X2_HVT U637 ( .A1(n99), .A2(n352), .A3(n100), .Y(out[58]) );
  NAND2X0_HVT U638 ( .A1(n151), .A2(n544), .Y(n485) );
  NAND2X0_HVT U639 ( .A1(n484), .A2(n381), .Y(n486) );
  NAND2X0_HVT U640 ( .A1(n486), .A2(n485), .Y(n536) );
  XOR3X2_HVT U641 ( .A1(n497), .A2(n487), .A3(n181), .Y(n212) );
  XOR3X2_HVT U642 ( .A1(n157), .A2(n350), .A3(n453), .Y(n155) );
  XOR2X2_HVT U643 ( .A1(n458), .A2(in[60]), .Y(n111) );
  INVX1_HVT U644 ( .A(n533), .Y(n488) );
  XNOR2X2_HVT U645 ( .A1(n489), .A2(n170), .Y(out[19]) );
  INVX0_HVT U646 ( .A(in[34]), .Y(n511) );
  XNOR2X2_HVT U647 ( .A1(n491), .A2(n461), .Y(out[52]) );
  NBUFFX2_HVT U648 ( .A(in[55]), .Y(n494) );
  XOR2X1_HVT U649 ( .A1(n4), .A2(n569), .Y(n187) );
  XOR3X2_HVT U650 ( .A1(n218), .A2(n499), .A3(n209), .Y(out[103]) );
  NBUFFX2_HVT U651 ( .A(in[111]), .Y(n567) );
  INVX1_HVT U652 ( .A(n500), .Y(n501) );
  XOR3X2_HVT U653 ( .A1(n24), .A2(n307), .A3(n188), .Y(out[114]) );
  XOR3X2_HVT U654 ( .A1(n38), .A2(n518), .A3(n502), .Y(n36) );
  XOR3X2_HVT U655 ( .A1(n189), .A2(n488), .A3(n188), .Y(out[122]) );
  INVX1_HVT U656 ( .A(in[114]), .Y(n533) );
  XOR3X2_HVT U657 ( .A1(n503), .A2(n568), .A3(n498), .Y(n211) );
  XOR3X2_HVT U658 ( .A1(n244), .A2(n323), .A3(n196), .Y(n531) );
  XOR2X2_HVT U659 ( .A1(n583), .A2(n570), .Y(n209) );
  XNOR2X2_HVT U660 ( .A1(in[112]), .A2(n583), .Y(n193) );
  XOR3X2_HVT U661 ( .A1(n522), .A2(n509), .A3(n453), .Y(n135) );
  XNOR2X2_HVT U662 ( .A1(n167), .A2(n448), .Y(out[20]) );
  INVX1_HVT U663 ( .A(n511), .Y(n512) );
  XNOR2X2_HVT U664 ( .A1(in[42]), .A2(n25), .Y(n99) );
  XOR3X2_HVT U665 ( .A1(n44), .A2(n514), .A3(n33), .Y(out[74]) );
  XOR3X2_HVT U666 ( .A1(n71), .A2(n506), .A3(n58), .Y(out[66]) );
  NBUFFX2_HVT U667 ( .A(in[87]), .Y(n518) );
  XNOR2X2_HVT U668 ( .A1(n141), .A2(n525), .Y(out[35]) );
  XOR3X2_HVT U669 ( .A1(n347), .A2(n552), .A3(n25), .Y(n525) );
  XOR3X2_HVT U670 ( .A1(n526), .A2(n533), .A3(n274), .Y(n186) );
  XOR3X2_HVT U671 ( .A1(in[115]), .A2(n498), .A3(n572), .Y(n19) );
  XNOR2X2_HVT U672 ( .A1(n531), .A2(n195), .Y(out[11]) );
  XOR3X2_HVT U673 ( .A1(n534), .A2(n460), .A3(n32), .Y(n67) );
  XOR3X2_HVT U674 ( .A1(in[92]), .A2(n564), .A3(n351), .Y(n535) );
  XOR2X2_HVT U675 ( .A1(in[20]), .A2(in[28]), .Y(n151) );
  XOR3X2_HVT U676 ( .A1(n537), .A2(n493), .A3(n93), .Y(n92) );
  XOR2X2_HVT U677 ( .A1(n545), .A2(n543), .Y(n146) );
  XNOR2X2_HVT U678 ( .A1(in[102]), .A2(in[110]), .Y(n178) );
  XNOR2X2_HVT U679 ( .A1(in[101]), .A2(in[109]), .Y(n180) );
  XOR2X2_HVT U680 ( .A1(in[13]), .A2(in[5]), .Y(n150) );
  XOR2X2_HVT U681 ( .A1(n306), .A2(in[65]), .Y(n58) );
  XOR2X2_HVT U682 ( .A1(in[64]), .A2(n560), .Y(n74) );
  XNOR2X2_HVT U683 ( .A1(in[45]), .A2(in[37]), .Y(n89) );
  XNOR2X2_HVT U684 ( .A1(in[21]), .A2(in[29]), .Y(n94) );
  XOR2X2_HVT U685 ( .A1(n380), .A2(n561), .Y(n61) );
  XNOR2X1_HVT U686 ( .A1(n548), .A2(n549), .Y(n63) );
  NBUFFX2_HVT U687 ( .A(in[39]), .Y(n552) );
  NBUFFX2_HVT U688 ( .A(in[15]), .Y(n546) );
  NBUFFX2_HVT U689 ( .A(in[15]), .Y(n545) );
  NBUFFX2_HVT U690 ( .A(in[63]), .Y(n558) );
  NBUFFX2_HVT U691 ( .A(in[95]), .Y(n566) );
  NBUFFX2_HVT U692 ( .A(in[111]), .Y(n568) );
  NBUFFX2_HVT U693 ( .A(in[23]), .Y(n548) );
  NBUFFX2_HVT U694 ( .A(in[31]), .Y(n551) );
  NBUFFX2_HVT U695 ( .A(n261), .Y(n563) );
  NBUFFX2_HVT U696 ( .A(in[71]), .Y(n560) );
  NBUFFX2_HVT U697 ( .A(in[7]), .Y(n543) );
  NBUFFX2_HVT U698 ( .A(in[63]), .Y(n557) );
  NBUFFX2_HVT U699 ( .A(in[7]), .Y(n542) );
  NBUFFX2_HVT U700 ( .A(n261), .Y(n562) );
  NBUFFX2_HVT U701 ( .A(in[63]), .Y(n556) );
  NBUFFX2_HVT U702 ( .A(in[31]), .Y(n550) );
  NBUFFX2_HVT U703 ( .A(in[23]), .Y(n547) );
  NBUFFX2_HVT U704 ( .A(in[15]), .Y(n544) );
  NBUFFX2_HVT U705 ( .A(in[127]), .Y(n569) );
  NBUFFX2_HVT U706 ( .A(in[31]), .Y(n549) );
  NBUFFX2_HVT U707 ( .A(in[47]), .Y(n553) );
  XOR2X1_HVT U708 ( .A1(n373), .A2(n302), .Y(n77) );
  INVX0_HVT U709 ( .A(in[0]), .Y(n577) );
  INVX0_HVT U710 ( .A(in[32]), .Y(n581) );
endmodule

