
module sbox_9 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n10, n17, n19, n23, n45, n46, n50, n51, n72, n73, n113, n114, n117,
         n118, n119, n170, n210, n211, n212, n213, n216, n217, n218, n219,
         n229, n231, n232, n235, n236, n238, n241, n249, n252, n253, n256,
         n258, n261, n264, n268, n273, n274, n275, n280, n282, n283, n285,
         n289, n293, n297, n301, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767;

  NAND2X0_HVT U4 ( .A1(n217), .A2(n765), .Y(n764) );
  NAND2X0_HVT U5 ( .A1(n312), .A2(n494), .Y(n762) );
  NAND2X0_HVT U15 ( .A1(n765), .A2(n231), .Y(n753) );
  NAND2X0_HVT U21 ( .A1(n497), .A2(n415), .Y(n749) );
  NAND2X0_HVT U24 ( .A1(n372), .A2(n446), .Y(n747) );
  NAND2X0_HVT U33 ( .A1(n540), .A2(n446), .Y(n738) );
  NAND2X0_HVT U35 ( .A1(n280), .A2(n383), .Y(n736) );
  NAND2X0_HVT U42 ( .A1(n268), .A2(n379), .Y(n729) );
  MUX41X1_HVT U51 ( .A1(n522), .A3(n544), .A2(n321), .A4(n524), .S0(n468), 
        .S1(n509), .Y(n724) );
  NAND2X0_HVT U53 ( .A1(n721), .A2(n728), .Y(n722) );
  NAND2X0_HVT U56 ( .A1(n498), .A2(n717), .Y(n718) );
  NAND2X0_HVT U58 ( .A1(n324), .A2(n347), .Y(n715) );
  NAND2X0_HVT U62 ( .A1(n415), .A2(n216), .Y(n711) );
  MUX41X1_HVT U63 ( .A1(n711), .A3(n526), .A2(n356), .A4(n525), .S0(n469), 
        .S1(n509), .Y(n710) );
  AO21X1_HVT U66 ( .A1(n557), .A2(n488), .A3(n559), .Y(n707) );
  NAND2X0_HVT U73 ( .A1(n702), .A2(n338), .Y(n703) );
  AND2X1_HVT U83 ( .A1(n361), .A2(n439), .Y(n691) );
  NAND2X0_HVT U85 ( .A1(n446), .A2(n342), .Y(n689) );
  MUX41X1_HVT U86 ( .A1(n552), .A3(n689), .A2(n473), .A4(n471), .S0(n386), 
        .S1(n466), .Y(n688) );
  AO21X1_HVT U93 ( .A1(n468), .A2(n681), .A3(n551), .Y(n682) );
  NAND2X0_HVT U101 ( .A1(n672), .A2(n671), .Y(n673) );
  MUX41X1_HVT U105 ( .A1(n550), .A3(n725), .A2(n668), .A4(n543), .S0(n386), 
        .S1(n466), .Y(n667) );
  NAND2X0_HVT U110 ( .A1(n500), .A2(n664), .Y(n665) );
  AND2X1_HVT U115 ( .A1(n268), .A2(n231), .Y(n662) );
  MUX41X1_HVT U116 ( .A1(n756), .A3(n662), .A2(n517), .A4(n740), .S0(n119), 
        .S1(n448), .Y(n661) );
  NAND2X0_HVT U123 ( .A1(n653), .A2(n652), .Y(n654) );
  MUX41X1_HVT U125 ( .A1(n749), .A3(n478), .A2(n528), .A4(n539), .S0(n119), 
        .S1(n432), .Y(n650) );
  MUX41X1_HVT U135 ( .A1(n531), .A3(n390), .A2(n762), .A4(n744), .S0(n485), 
        .S1(n469), .Y(n641) );
  MUX41X1_HVT U136 ( .A1(n471), .A3(n738), .A2(n521), .A4(n735), .S0(n380), 
        .S1(n469), .Y(n640) );
  AND2X1_HVT U140 ( .A1(n389), .A2(n353), .Y(n636) );
  MUX41X1_HVT U141 ( .A1(n746), .A3(n538), .A2(n636), .A4(n536), .S0(n485), 
        .S1(n448), .Y(n635) );
  MUX41X1_HVT U153 ( .A1(n665), .A3(n475), .A2(n216), .A4(n436), .S0(n380), 
        .S1(n399), .Y(n624) );
  AND2X1_HVT U154 ( .A1(n399), .A2(n372), .Y(n623) );
  NAND2X0_HVT U158 ( .A1(n268), .A2(n398), .Y(n619) );
  MUX41X1_HVT U159 ( .A1(n756), .A3(n231), .A2(n619), .A4(n560), .S0(n119), 
        .S1(n399), .Y(n618) );
  AND2X1_HVT U162 ( .A1(n229), .A2(n702), .Y(n615) );
  MUX41X1_HVT U163 ( .A1(n414), .A3(n615), .A2(n472), .A4(n616), .S0(n380), 
        .S1(n512), .Y(n614) );
  NAND2X0_HVT U166 ( .A1(n324), .A2(n717), .Y(n612) );
  NAND2X0_HVT U167 ( .A1(n520), .A2(n446), .Y(n611) );
  MUX41X1_HVT U168 ( .A1(n533), .A3(n338), .A2(n611), .A4(n612), .S0(n386), 
        .S1(n512), .Y(n610) );
  NAND2X0_HVT U177 ( .A1(n297), .A2(n280), .Y(n603) );
  MUX41X1_HVT U189 ( .A1(n592), .A3(n755), .A2(n593), .A4(n543), .S0(n432), 
        .S1(n17), .Y(n591) );
  MUX41X1_HVT U194 ( .A1(n730), .A3(n744), .A2(n531), .A4(n389), .S0(n448), 
        .S1(n485), .Y(n587) );
  MUX41X1_HVT U195 ( .A1(n229), .A3(n554), .A2(n503), .A4(n734), .S0(n119), 
        .S1(n343), .Y(n586) );
  NAND2X0_HVT U212 ( .A1(n312), .A2(n212), .Y(n717) );
  NAND2X0_HVT U214 ( .A1(n311), .A2(n383), .Y(n574) );
  NAND2X0_HVT U215 ( .A1(n664), .A2(n496), .Y(n573) );
  NAND2X0_HVT U218 ( .A1(n553), .A2(n453), .Y(n626) );
  NAND2X0_HVT U220 ( .A1(n514), .A2(n574), .Y(n694) );
  INVX0_HVT U241 ( .A(n747), .Y(n562) );
  INVX0_HVT U245 ( .A(n762), .Y(n560) );
  INVX0_HVT U250 ( .A(n758), .Y(n557) );
  INVX0_HVT U256 ( .A(n626), .Y(n551) );
  INVX0_HVT U268 ( .A(n749), .Y(n544) );
  INVX0_HVT U270 ( .A(n573), .Y(n543) );
  INVX0_HVT U273 ( .A(n681), .Y(n541) );
  INVX0_HVT U280 ( .A(n742), .Y(n535) );
  INVX0_HVT U289 ( .A(n671), .Y(n530) );
  INVX0_HVT U295 ( .A(n764), .Y(n527) );
  INVX0_HVT U296 ( .A(n753), .Y(n526) );
  INVX0_HVT U302 ( .A(n572), .Y(n522) );
  INVX0_HVT U306 ( .A(n611), .Y(n519) );
  INVX0_HVT U307 ( .A(n731), .Y(n518) );
  MUX21X1_HVT U1 ( .A1(n367), .A2(n405), .S0(n238), .Y(n416) );
  INVX1_HVT U2 ( .A(n114), .Y(n229) );
  INVX1_HVT U3 ( .A(n664), .Y(n542) );
  XOR2X1_HVT U6 ( .A1(n280), .A2(n504), .Y(n745) );
  INVX1_HVT U7 ( .A(n547), .Y(n439) );
  AND3X1_HVT U8 ( .A1(n500), .A2(n717), .A3(n694), .Y(n695) );
  MUX21X1_HVT U9 ( .A1(n457), .A2(n496), .S0(n368), .Y(n668) );
  OAI21X1_HVT U10 ( .A1(n441), .A2(n463), .A3(n416), .Y(n483) );
  MUX21X1_HVT U11 ( .A1(n609), .A2(n608), .S0(n17), .Y(n607) );
  INVX1_HVT U12 ( .A(n378), .Y(n737) );
  INVX1_HVT U13 ( .A(n339), .Y(n446) );
  INVX1_HVT U14 ( .A(n317), .Y(n212) );
  INVX1_HVT U16 ( .A(n507), .Y(n232) );
  INVX0_HVT U17 ( .A(in[1]), .Y(n418) );
  AND2X1_HVT U18 ( .A1(n377), .A2(n376), .Y(n10) );
  INVX1_HVT U19 ( .A(n547), .Y(n360) );
  INVX1_HVT U20 ( .A(n467), .Y(n761) );
  NAND2X0_HVT U22 ( .A1(n385), .A2(n17), .Y(n19) );
  NAND2X0_HVT U23 ( .A1(n556), .A2(n417), .Y(n23) );
  NAND2X0_HVT U25 ( .A1(n19), .A2(n23), .Y(n384) );
  INVX0_HVT U26 ( .A(n417), .Y(n17) );
  OA21X1_HVT U27 ( .A1(n476), .A2(n455), .A3(n740), .Y(n608) );
  OA21X1_HVT U28 ( .A1(n519), .A2(n455), .A3(n740), .Y(n632) );
  MUX21X1_HVT U29 ( .A1(n752), .A2(n536), .S0(n484), .Y(n645) );
  MUX21X1_HVT U30 ( .A1(n741), .A2(n550), .S0(n232), .Y(n648) );
  MUX41X1_HVT U31 ( .A1(n688), .A3(n692), .A2(n690), .A4(n693), .S0(n489), 
        .S1(n509), .Y(n687) );
  NAND2X0_HVT U32 ( .A1(n643), .A2(n386), .Y(n45) );
  NAND2X0_HVT U34 ( .A1(n516), .A2(n374), .Y(n46) );
  NAND2X0_HVT U36 ( .A1(n45), .A2(n46), .Y(n642) );
  MUX41X1_HVT U37 ( .A1(n533), .A3(n751), .A2(n718), .A4(n758), .S0(n468), 
        .S1(n509), .Y(n716) );
  INVX0_HVT U38 ( .A(n761), .Y(n114) );
  INVX0_HVT U39 ( .A(n502), .Y(n558) );
  MUX41X1_HVT U40 ( .A1(n631), .A3(n630), .A2(n635), .A4(n634), .S0(n428), 
        .S1(n489), .Y(n629) );
  MUX21X2_HVT U41 ( .A1(n458), .A2(n379), .S0(n453), .Y(n748) );
  INVX1_HVT U43 ( .A(n413), .Y(n396) );
  INVX0_HVT U44 ( .A(n558), .Y(n50) );
  OR2X1_HVT U45 ( .A1(n322), .A2(n490), .Y(n329) );
  NAND2X0_HVT U46 ( .A1(n495), .A2(n282), .Y(n51) );
  NAND2X0_HVT U47 ( .A1(n558), .A2(n238), .Y(n72) );
  NAND2X0_HVT U48 ( .A1(n51), .A2(n72), .Y(n758) );
  NAND2X0_HVT U49 ( .A1(n311), .A2(n446), .Y(n73) );
  NAND2X0_HVT U50 ( .A1(n492), .A2(n361), .Y(n113) );
  NAND2X0_HVT U52 ( .A1(n73), .A2(n113), .Y(n699) );
  MUX41X1_HVT U54 ( .A1(n529), .A3(n456), .A2(n542), .A4(n389), .S0(n484), 
        .S1(n468), .Y(n634) );
  INVX0_HVT U55 ( .A(n730), .Y(n523) );
  MUX21X2_HVT U57 ( .A1(n472), .A2(n454), .S0(n256), .Y(n646) );
  MUX21X2_HVT U59 ( .A1(n457), .A2(n464), .S0(n361), .Y(n679) );
  INVX1_HVT U60 ( .A(n484), .Y(n374) );
  MUX21X1_HVT U61 ( .A1(n436), .A2(n378), .S0(n256), .Y(n660) );
  INVX1_HVT U64 ( .A(n515), .Y(n512) );
  INVX1_HVT U65 ( .A(n507), .Y(n417) );
  MUX21X1_HVT U67 ( .A1(n503), .A2(n499), .S0(n383), .Y(n451) );
  INVX1_HVT U68 ( .A(n360), .Y(n280) );
  XNOR2X1_HVT U69 ( .A1(n398), .A2(n452), .Y(n473) );
  INVX1_HVT U70 ( .A(n212), .Y(n553) );
  OA21X1_HVT U71 ( .A1(n731), .A2(n455), .A3(n626), .Y(n627) );
  INVX0_HVT U72 ( .A(n502), .Y(n398) );
  NAND2X0_HVT U74 ( .A1(n541), .A2(n343), .Y(n345) );
  XNOR2X1_HVT U75 ( .A1(n311), .A2(n415), .Y(n727) );
  INVX1_HVT U76 ( .A(n574), .Y(n534) );
  INVX1_HVT U77 ( .A(n515), .Y(n466) );
  INVX1_HVT U78 ( .A(n589), .Y(n437) );
  NAND2X0_HVT U79 ( .A1(n722), .A2(n362), .Y(n258) );
  INVX1_HVT U80 ( .A(n374), .Y(n119) );
  NAND2X0_HVT U81 ( .A1(n659), .A2(n264), .Y(n309) );
  INVX1_HVT U82 ( .A(n417), .Y(n256) );
  INVX0_HVT U84 ( .A(n515), .Y(n513) );
  NBUFFX2_HVT U87 ( .A(n507), .Y(n484) );
  INVX1_HVT U88 ( .A(n487), .Y(n235) );
  INVX1_HVT U89 ( .A(n505), .Y(n452) );
  INVX0_HVT U90 ( .A(n513), .Y(n455) );
  INVX1_HVT U91 ( .A(n486), .Y(n348) );
  NBUFFX2_HVT U92 ( .A(n510), .Y(n488) );
  INVX1_HVT U94 ( .A(n369), .Y(n231) );
  INVX0_HVT U95 ( .A(n320), .Y(n330) );
  INVX0_HVT U96 ( .A(n553), .Y(n338) );
  INVX0_HVT U97 ( .A(n514), .Y(n426) );
  AND2X1_HVT U98 ( .A1(n273), .A2(n274), .Y(n117) );
  INVX0_HVT U99 ( .A(n367), .Y(n390) );
  INVX1_HVT U100 ( .A(n729), .Y(n561) );
  INVX0_HVT U102 ( .A(n559), .Y(n118) );
  INVX0_HVT U103 ( .A(n765), .Y(n397) );
  MUX41X1_HVT U104 ( .A1(n529), .A3(n229), .A2(n445), .A4(n691), .S0(n119), 
        .S1(n343), .Y(n690) );
  AND2X1_HVT U106 ( .A1(n315), .A2(n316), .Y(n170) );
  INVX1_HVT U107 ( .A(n452), .Y(n238) );
  MUX41X1_HVT U108 ( .A1(n595), .A3(n598), .A2(n591), .A4(n594), .S0(n487), 
        .S1(n427), .Y(n590) );
  MUX41X1_HVT U109 ( .A1(n756), .A3(n470), .A2(n527), .A4(n759), .S0(n469), 
        .S1(n417), .Y(n600) );
  INVX0_HVT U111 ( .A(n702), .Y(n559) );
  INVX0_HVT U112 ( .A(n506), .Y(n313) );
  MUX21X2_HVT U113 ( .A1(n500), .A2(n114), .S0(n361), .Y(n730) );
  INVX0_HVT U114 ( .A(n743), .Y(n550) );
  INVX1_HVT U117 ( .A(n745), .Y(n546) );
  INVX0_HVT U118 ( .A(n503), .Y(n342) );
  INVX0_HVT U119 ( .A(n447), .Y(n732) );
  MUX21X2_HVT U120 ( .A1(n423), .A2(n497), .S0(n339), .Y(n447) );
  AND2X1_HVT U121 ( .A1(n301), .A2(n303), .Y(n210) );
  MUX41X1_HVT U122 ( .A1(n638), .A3(n641), .A2(n640), .A4(n642), .S0(n489), 
        .S1(n488), .Y(n637) );
  INVX0_HVT U124 ( .A(n761), .Y(n456) );
  MUX41X1_HVT U126 ( .A1(n727), .A3(n749), .A2(n117), .A4(n549), .S0(n348), 
        .S1(n469), .Y(n613) );
  NAND2X0_HVT U127 ( .A1(n491), .A2(n493), .Y(n211) );
  INVX0_HVT U128 ( .A(n506), .Y(n504) );
  INVX1_HVT U129 ( .A(n458), .Y(n369) );
  MUX21X1_HVT U130 ( .A1(n439), .A2(n464), .S0(n383), .Y(n739) );
  INVX1_HVT U131 ( .A(n505), .Y(n383) );
  INVX1_HVT U132 ( .A(n428), .Y(n213) );
  INVX1_HVT U133 ( .A(n480), .Y(n216) );
  INVX1_HVT U134 ( .A(n500), .Y(n480) );
  INVX0_HVT U137 ( .A(n413), .Y(n735) );
  INVX0_HVT U138 ( .A(n540), .Y(n217) );
  MUX41X1_HVT U139 ( .A1(n552), .A3(n555), .A2(n517), .A4(n480), .S0(n374), 
        .S1(n512), .Y(n700) );
  MUX21X2_HVT U142 ( .A1(n447), .A2(n748), .S0(n408), .Y(n639) );
  INVX0_HVT U143 ( .A(n482), .Y(n663) );
  INVX0_HVT U144 ( .A(n317), .Y(n367) );
  NAND2X0_HVT U145 ( .A1(n405), .A2(n368), .Y(n218) );
  NAND2X0_HVT U146 ( .A1(n495), .A2(n313), .Y(n219) );
  NAND2X0_HVT U147 ( .A1(n218), .A2(n219), .Y(n757) );
  INVX1_HVT U148 ( .A(n506), .Y(n304) );
  INVX1_HVT U149 ( .A(n746), .Y(n517) );
  MUX21X2_HVT U150 ( .A1(n311), .A2(n520), .S0(n339), .Y(n746) );
  INVX1_HVT U151 ( .A(n490), .Y(n440) );
  NAND2X0_HVT U152 ( .A1(n313), .A2(n50), .Y(n702) );
  INVX1_HVT U155 ( .A(n342), .Y(n324) );
  MUX41X1_HVT U156 ( .A1(n556), .A3(n548), .A2(n347), .A4(n439), .S0(n232), 
        .S1(n426), .Y(n576) );
  MUX21X2_HVT U157 ( .A1(n337), .A2(n280), .S0(n465), .Y(n413) );
  INVX1_HVT U160 ( .A(n761), .Y(n458) );
  INVX0_HVT U161 ( .A(n445), .Y(n454) );
  NAND2X0_HVT U164 ( .A1(n361), .A2(n763), .Y(n664) );
  MUX41X1_HVT U165 ( .A1(n395), .A3(n483), .A2(n479), .A4(n384), .S0(n399), 
        .S1(n428), .Y(n482) );
  INVX1_HVT U169 ( .A(n455), .Y(n399) );
  INVX1_HVT U170 ( .A(n466), .Y(n236) );
  INVX1_HVT U171 ( .A(n740), .Y(n556) );
  INVX0_HVT U172 ( .A(n761), .Y(n457) );
  INVX1_HVT U173 ( .A(n512), .Y(n264) );
  XOR2X1_HVT U174 ( .A1(n513), .A2(n313), .Y(n477) );
  INVX0_HVT U175 ( .A(n506), .Y(n453) );
  INVX0_HVT U176 ( .A(n506), .Y(n312) );
  OA21X1_HVT U178 ( .A1(n737), .A2(n515), .A3(n529), .Y(n596) );
  MUX21X1_HVT U179 ( .A1(n597), .A2(n596), .S0(n232), .Y(n595) );
  INVX1_HVT U180 ( .A(n465), .Y(n297) );
  INVX1_HVT U181 ( .A(n717), .Y(n555) );
  MUX41X1_HVT U182 ( .A1(n670), .A3(n667), .A2(n674), .A4(n669), .S0(n427), 
        .S1(n487), .Y(n666) );
  NBUFFX2_HVT U183 ( .A(n440), .Y(n494) );
  MUX21X1_HVT U184 ( .A1(n379), .A2(n502), .S0(n452), .Y(n378) );
  AND3X1_HVT U185 ( .A1(n485), .A2(n353), .A3(n439), .Y(n647) );
  MUX41X1_HVT U186 ( .A1(n748), .A3(n378), .A2(n756), .A4(n718), .S0(n375), 
        .S1(n236), .Y(n577) );
  INVX1_HVT U187 ( .A(n232), .Y(n386) );
  MUX21X2_HVT U188 ( .A1(n210), .A2(n390), .S0(n488), .Y(n706) );
  INVX1_HVT U190 ( .A(n499), .Y(n520) );
  NAND2X0_HVT U191 ( .A1(n439), .A2(n238), .Y(n241) );
  NAND2X0_HVT U192 ( .A1(n494), .A2(n452), .Y(n249) );
  NAND2X0_HVT U193 ( .A1(n241), .A2(n249), .Y(n741) );
  INVX1_HVT U196 ( .A(n741), .Y(n549) );
  NAND2X0_HVT U197 ( .A1(n655), .A2(n362), .Y(n252) );
  NAND2X0_HVT U198 ( .A1(n654), .A2(n343), .Y(n253) );
  NAND2X0_HVT U199 ( .A1(n252), .A2(n253), .Y(n651) );
  MUX21X1_HVT U200 ( .A1(n537), .A2(n656), .S0(n485), .Y(n655) );
  NAND2X0_HVT U201 ( .A1(n723), .A2(n448), .Y(n261) );
  NAND2X0_HVT U202 ( .A1(n258), .A2(n261), .Y(n720) );
  MUX21X1_HVT U203 ( .A1(n492), .A2(n423), .S0(n417), .Y(n422) );
  INVX1_HVT U204 ( .A(n504), .Y(n368) );
  INVX1_HVT U205 ( .A(n490), .Y(n327) );
  MUX41X1_HVT U206 ( .A1(n554), .A3(n679), .A2(n562), .A4(n474), .S0(n119), 
        .S1(n264), .Y(n678) );
  INVX0_HVT U207 ( .A(n515), .Y(n514) );
  MUX21X1_HVT U208 ( .A1(n682), .A2(n683), .S0(n486), .Y(n680) );
  NAND2X0_HVT U209 ( .A1(n500), .A2(n268), .Y(n273) );
  NAND2X0_HVT U210 ( .A1(n389), .A2(n353), .Y(n274) );
  INVX0_HVT U211 ( .A(n465), .Y(n268) );
  INVX0_HVT U213 ( .A(n553), .Y(n389) );
  NBUFFX2_HVT U216 ( .A(n513), .Y(n469) );
  MUX41X1_HVT U217 ( .A1(n588), .A3(n586), .A2(n587), .A4(n583), .S0(n427), 
        .S1(n235), .Y(n582) );
  INVX1_HVT U219 ( .A(n327), .Y(n275) );
  NBUFFX2_HVT U221 ( .A(n322), .Y(n491) );
  INVX1_HVT U222 ( .A(n739), .Y(n536) );
  INVX0_HVT U223 ( .A(n757), .Y(n545) );
  NAND2X0_HVT U224 ( .A1(n405), .A2(n282), .Y(n283) );
  NAND2X0_HVT U225 ( .A1(n337), .A2(n453), .Y(n285) );
  NAND2X0_HVT U226 ( .A1(n283), .A2(n285), .Y(n681) );
  INVX0_HVT U227 ( .A(n504), .Y(n282) );
  NBUFFX2_HVT U228 ( .A(n767), .Y(n337) );
  MUX41X1_HVT U229 ( .A1(n624), .A3(n618), .A2(n625), .A4(n620), .S0(n427), 
        .S1(n213), .Y(n617) );
  INVX1_HVT U230 ( .A(n211), .Y(n464) );
  MUX41X1_HVT U231 ( .A1(n210), .A3(n347), .A2(n736), .A4(n535), .S0(n374), 
        .S1(n432), .Y(n669) );
  INVX0_HVT U232 ( .A(n321), .Y(n751) );
  AO21X1_HVT U233 ( .A1(n473), .A2(n399), .A3(n551), .Y(n584) );
  NAND2X0_HVT U234 ( .A1(n621), .A2(n348), .Y(n289) );
  NAND2X0_HVT U235 ( .A1(n622), .A2(n485), .Y(n293) );
  NAND2X0_HVT U236 ( .A1(n289), .A2(n293), .Y(n620) );
  INVX0_HVT U237 ( .A(n451), .Y(n744) );
  NAND2X0_HVT U238 ( .A1(n379), .A2(n297), .Y(n301) );
  NAND2X0_HVT U239 ( .A1(n498), .A2(n465), .Y(n303) );
  NAND2X0_HVT U240 ( .A1(n301), .A2(n303), .Y(n759) );
  NAND2X0_HVT U242 ( .A1(n456), .A2(n312), .Y(n305) );
  NAND2X0_HVT U243 ( .A1(n540), .A2(n506), .Y(n306) );
  NAND2X0_HVT U244 ( .A1(n305), .A2(n306), .Y(n463) );
  INVX0_HVT U246 ( .A(n405), .Y(n540) );
  INVX1_HVT U247 ( .A(in[1]), .Y(n506) );
  MUX41X1_HVT U248 ( .A1(n706), .A3(n528), .A2(n708), .A4(n707), .S0(n426), 
        .S1(n386), .Y(n705) );
  MUX21X1_HVT U249 ( .A1(n545), .A2(n446), .S0(n488), .Y(n708) );
  INVX0_HVT U251 ( .A(n760), .Y(n528) );
  INVX0_HVT U252 ( .A(n748), .Y(n529) );
  INVX1_HVT U253 ( .A(n494), .Y(n379) );
  NBUFFX2_HVT U254 ( .A(n327), .Y(n493) );
  INVX0_HVT U255 ( .A(n477), .Y(n402) );
  NAND2X0_HVT U257 ( .A1(n581), .A2(n486), .Y(n307) );
  NAND2X0_HVT U258 ( .A1(n580), .A2(n348), .Y(n308) );
  NAND2X0_HVT U259 ( .A1(n307), .A2(n308), .Y(n579) );
  INVX0_HVT U260 ( .A(n505), .Y(n465) );
  XNOR2X2_HVT U261 ( .A1(n497), .A2(n361), .Y(n472) );
  INVX1_HVT U262 ( .A(n418), .Y(n361) );
  NAND2X0_HVT U263 ( .A1(n660), .A2(n513), .Y(n310) );
  NAND2X0_HVT U264 ( .A1(n309), .A2(n310), .Y(n658) );
  AND2X1_HVT U265 ( .A1(n329), .A2(n328), .Y(n311) );
  INVX0_HVT U266 ( .A(n738), .Y(n537) );
  INVX1_HVT U267 ( .A(n571), .Y(n533) );
  MUX41X1_HVT U269 ( .A1(n715), .A3(n478), .A2(n416), .A4(n476), .S0(n408), 
        .S1(n509), .Y(n714) );
  MUX41X1_HVT U271 ( .A1(n743), .A3(n534), .A2(n548), .A4(n170), .S0(n512), 
        .S1(n256), .Y(n601) );
  NAND2X0_HVT U272 ( .A1(n496), .A2(n314), .Y(n315) );
  NAND2X0_HVT U274 ( .A1(n439), .A2(n368), .Y(n316) );
  INVX0_HVT U275 ( .A(n368), .Y(n314) );
  INVX1_HVT U276 ( .A(in[7]), .Y(n515) );
  AND2X1_HVT U277 ( .A1(n440), .A2(n360), .Y(n317) );
  INVX1_HVT U278 ( .A(in[2]), .Y(n508) );
  NBUFFX2_HVT U279 ( .A(in[3]), .Y(n490) );
  INVX0_HVT U281 ( .A(in[5]), .Y(n511) );
  NAND2X0_HVT U282 ( .A1(n496), .A2(n268), .Y(n318) );
  NAND2X0_HVT U283 ( .A1(n500), .A2(n282), .Y(n319) );
  NAND2X0_HVT U284 ( .A1(n318), .A2(n319), .Y(n754) );
  NBUFFX2_HVT U285 ( .A(n212), .Y(n496) );
  INVX0_HVT U286 ( .A(n754), .Y(n525) );
  INVX0_HVT U287 ( .A(in[4]), .Y(n322) );
  INVX0_HVT U288 ( .A(in[6]), .Y(n320) );
  NAND2X0_HVT U290 ( .A1(n352), .A2(n351), .Y(out[1]) );
  NAND2X0_HVT U291 ( .A1(n556), .A2(n348), .Y(n349) );
  MUX21X1_HVT U292 ( .A1(n495), .A2(n499), .S0(n465), .Y(n321) );
  INVX1_HVT U293 ( .A(n418), .Y(n505) );
  INVX0_HVT U294 ( .A(in[4]), .Y(n547) );
  INVX1_HVT U297 ( .A(n484), .Y(n441) );
  MUX21X1_HVT U298 ( .A1(n212), .A2(n280), .S0(n361), .Y(n704) );
  MUX21X1_HVT U299 ( .A1(n570), .A2(n324), .S0(n426), .Y(n323) );
  INVX0_HVT U300 ( .A(n570), .Y(n554) );
  MUX41X1_HVT U301 ( .A1(n602), .A3(n604), .A2(n600), .A4(n601), .S0(n487), 
        .S1(n427), .Y(n599) );
  INVX1_HVT U303 ( .A(n415), .Y(n339) );
  MUX21X1_HVT U304 ( .A1(n464), .A2(n520), .S0(n313), .Y(n605) );
  MUX41X1_HVT U305 ( .A1(n579), .A3(n578), .A2(n577), .A4(n576), .S0(n428), 
        .S1(n427), .Y(n575) );
  INVX0_HVT U308 ( .A(n455), .Y(n432) );
  INVX0_HVT U309 ( .A(n455), .Y(n343) );
  INVX1_HVT U310 ( .A(n372), .Y(n423) );
  NAND2X0_HVT U311 ( .A1(n367), .A2(n426), .Y(n325) );
  NAND2X0_HVT U312 ( .A1(n554), .A2(n343), .Y(n326) );
  NAND2X0_HVT U313 ( .A1(n326), .A2(n325), .Y(n609) );
  NAND2X0_HVT U314 ( .A1(n275), .A2(n547), .Y(n328) );
  NAND2X0_HVT U315 ( .A1(n328), .A2(n329), .Y(n467) );
  NAND2X0_HVT U316 ( .A1(n676), .A2(n330), .Y(n331) );
  NAND2X0_HVT U317 ( .A1(n666), .A2(n320), .Y(n332) );
  NAND2X0_HVT U318 ( .A1(n331), .A2(n332), .Y(out[2]) );
  INVX1_HVT U319 ( .A(n508), .Y(n507) );
  NAND2X0_HVT U320 ( .A1(n695), .A2(n486), .Y(n333) );
  NAND2X0_HVT U321 ( .A1(n696), .A2(n348), .Y(n334) );
  NAND2X0_HVT U322 ( .A1(n333), .A2(n334), .Y(n693) );
  NAND2X0_HVT U323 ( .A1(n439), .A2(n282), .Y(n335) );
  NAND2X0_HVT U324 ( .A1(n501), .A2(n297), .Y(n336) );
  NAND2X0_HVT U325 ( .A1(n335), .A2(n336), .Y(n750) );
  MUX21X1_HVT U326 ( .A1(n338), .A2(n750), .S0(n426), .Y(n696) );
  INVX1_HVT U327 ( .A(n750), .Y(n524) );
  MUX21X1_HVT U328 ( .A1(n573), .A2(n741), .S0(n408), .Y(n567) );
  MUX41X1_HVT U329 ( .A1(n704), .A3(n745), .A2(n703), .A4(n747), .S0(n386), 
        .S1(n512), .Y(n701) );
  INVX1_HVT U330 ( .A(n441), .Y(n380) );
  INVX1_HVT U331 ( .A(n564), .Y(n521) );
  INVX1_HVT U332 ( .A(n505), .Y(n415) );
  MUX41X1_HVT U333 ( .A1(n646), .A3(n648), .A2(n645), .A4(n647), .S0(n213), 
        .S1(n362), .Y(n644) );
  MUX21X2_HVT U334 ( .A1(n367), .A2(n502), .S0(n452), .Y(n740) );
  INVX0_HVT U335 ( .A(n411), .Y(n692) );
  MUX41X1_HVT U336 ( .A1(n605), .A3(n492), .A2(n755), .A4(n530), .S0(n264), 
        .S1(n256), .Y(n604) );
  NAND2X0_HVT U337 ( .A1(n712), .A2(n485), .Y(n340) );
  NAND2X0_HVT U338 ( .A1(n710), .A2(n441), .Y(n341) );
  NAND2X0_HVT U339 ( .A1(n340), .A2(n341), .Y(n709) );
  INVX1_HVT U340 ( .A(n514), .Y(n408) );
  NBUFFX2_HVT U341 ( .A(n211), .Y(n498) );
  INVX0_HVT U342 ( .A(n463), .Y(n734) );
  NAND2X0_HVT U343 ( .A1(n528), .A2(n432), .Y(n344) );
  AND2X1_HVT U344 ( .A1(n344), .A2(n538), .Y(n580) );
  INVX0_HVT U345 ( .A(n733), .Y(n538) );
  MUX21X1_HVT U346 ( .A1(n558), .A2(n464), .S0(n304), .Y(n733) );
  NAND2X0_HVT U347 ( .A1(n733), .A2(n426), .Y(n346) );
  NAND2X0_HVT U348 ( .A1(n345), .A2(n346), .Y(n621) );
  INVX0_HVT U349 ( .A(n414), .Y(n752) );
  INVX1_HVT U350 ( .A(n356), .Y(n756) );
  MUX41X1_HVT U351 ( .A1(n729), .A3(n686), .A2(n727), .A4(n522), .S0(n466), 
        .S1(n441), .Y(n685) );
  NBUFFX2_HVT U352 ( .A(n322), .Y(n492) );
  INVX1_HVT U353 ( .A(n397), .Y(n347) );
  NAND2X0_HVT U354 ( .A1(n504), .A2(n499), .Y(n765) );
  NAND2X0_HVT U355 ( .A1(n754), .A2(n485), .Y(n350) );
  NAND2X0_HVT U356 ( .A1(n349), .A2(n350), .Y(n675) );
  NAND2X0_HVT U357 ( .A1(n697), .A2(n330), .Y(n351) );
  NAND2X0_HVT U358 ( .A1(n687), .A2(n320), .Y(n352) );
  NAND2X0_HVT U359 ( .A1(n217), .A2(n353), .Y(n354) );
  NAND2X0_HVT U360 ( .A1(n389), .A2(n361), .Y(n355) );
  NAND2X0_HVT U361 ( .A1(n354), .A2(n355), .Y(n686) );
  INVX0_HVT U362 ( .A(n268), .Y(n353) );
  AND2X1_HVT U363 ( .A1(n755), .A2(n324), .Y(n356) );
  NAND2X0_HVT U364 ( .A1(n494), .A2(n357), .Y(n358) );
  NAND2X0_HVT U365 ( .A1(n367), .A2(n282), .Y(n359) );
  NAND2X0_HVT U366 ( .A1(n359), .A2(n358), .Y(n570) );
  INVX0_HVT U367 ( .A(n368), .Y(n357) );
  INVX0_HVT U368 ( .A(n665), .Y(n385) );
  NAND2X0_HVT U369 ( .A1(n561), .A2(n362), .Y(n363) );
  NAND2X0_HVT U370 ( .A1(n170), .A2(n469), .Y(n364) );
  NAND2X0_HVT U371 ( .A1(n363), .A2(n364), .Y(n585) );
  INVX0_HVT U372 ( .A(n514), .Y(n362) );
  NAND2X0_HVT U373 ( .A1(n584), .A2(n119), .Y(n365) );
  NAND2X0_HVT U374 ( .A1(n585), .A2(n374), .Y(n366) );
  NAND2X0_HVT U375 ( .A1(n365), .A2(n366), .Y(n583) );
  MUX41X1_HVT U376 ( .A1(n541), .A3(n759), .A2(n532), .A4(n699), .S0(n264), 
        .S1(n17), .Y(n698) );
  NAND2X0_HVT U377 ( .A1(n590), .A2(n320), .Y(n370) );
  NAND2X0_HVT U378 ( .A1(n599), .A2(in[6]), .Y(n371) );
  NAND2X0_HVT U379 ( .A1(n370), .A2(n371), .Y(out[6]) );
  MUX41X1_HVT U380 ( .A1(n603), .A3(n752), .A2(n733), .A4(n170), .S0(n375), 
        .S1(n466), .Y(n602) );
  MUX41X1_HVT U381 ( .A1(n700), .A3(n10), .A2(n698), .A4(n701), .S0(n489), 
        .S1(n235), .Y(n697) );
  NBUFFX2_HVT U382 ( .A(n275), .Y(n372) );
  MUX41X1_HVT U383 ( .A1(n447), .A3(n523), .A2(n498), .A4(n546), .S0(n386), 
        .S1(n468), .Y(n598) );
  MUX41X1_HVT U384 ( .A1(n314), .A3(n753), .A2(n555), .A4(n474), .S0(n386), 
        .S1(n362), .Y(n677) );
  MUX41X1_HVT U385 ( .A1(n685), .A3(n678), .A2(n680), .A4(n677), .S0(n427), 
        .S1(n428), .Y(n676) );
  NAND2X0_HVT U386 ( .A1(n486), .A2(n389), .Y(n373) );
  NAND2X0_HVT U387 ( .A1(n373), .A2(n456), .Y(n659) );
  NAND2X0_HVT U388 ( .A1(n442), .A2(n375), .Y(n376) );
  NAND2X0_HVT U389 ( .A1(n323), .A2(n380), .Y(n377) );
  INVX0_HVT U390 ( .A(n380), .Y(n375) );
  XNOR2X1_HVT U391 ( .A1(n451), .A2(n468), .Y(n442) );
  MUX41X1_HVT U392 ( .A1(n727), .A3(n118), .A2(n732), .A4(n474), .S0(n417), 
        .S1(n362), .Y(n594) );
  NAND2X0_HVT U393 ( .A1(n714), .A2(n348), .Y(n381) );
  NAND2X0_HVT U394 ( .A1(n716), .A2(n486), .Y(n382) );
  NAND2X0_HVT U395 ( .A1(n382), .A2(n381), .Y(n713) );
  MUX41X1_HVT U396 ( .A1(n739), .A3(n757), .A2(n518), .A4(n735), .S0(n374), 
        .S1(n408), .Y(n578) );
  INVX1_HVT U397 ( .A(n487), .Y(n428) );
  MUX41X1_HVT U398 ( .A1(n475), .A3(n414), .A2(n454), .A4(n231), .S0(n468), 
        .S1(n509), .Y(n712) );
  NAND2X0_HVT U399 ( .A1(n764), .A2(n386), .Y(n387) );
  NAND2X0_HVT U400 ( .A1(n639), .A2(n441), .Y(n388) );
  NAND2X0_HVT U401 ( .A1(n388), .A2(n387), .Y(n638) );
  INVX1_HVT U402 ( .A(n569), .Y(n552) );
  MUX21X1_HVT U403 ( .A1(n114), .A2(n342), .S0(n312), .Y(n760) );
  NAND2X0_HVT U404 ( .A1(n582), .A2(n330), .Y(n391) );
  NAND2X0_HVT U405 ( .A1(n575), .A2(n320), .Y(n392) );
  NAND2X0_HVT U406 ( .A1(n391), .A2(n392), .Y(out[7]) );
  MUX21X1_HVT U407 ( .A1(n372), .A2(n736), .S0(n488), .Y(n723) );
  MUX41X1_HVT U408 ( .A1(n727), .A3(n555), .A2(n118), .A4(n521), .S0(n348), 
        .S1(n236), .Y(n630) );
  NAND2X0_HVT U409 ( .A1(n724), .A2(n486), .Y(n393) );
  NAND2X0_HVT U410 ( .A1(n720), .A2(n375), .Y(n394) );
  NAND2X0_HVT U411 ( .A1(n393), .A2(n394), .Y(n719) );
  MUX41X1_HVT U412 ( .A1(n613), .A3(n607), .A2(n614), .A4(n610), .S0(n427), 
        .S1(n213), .Y(n606) );
  MUX21X1_HVT U413 ( .A1(n396), .A2(n397), .S0(n484), .Y(n395) );
  NAND2X0_HVT U414 ( .A1(n443), .A2(n444), .Y(out[4]) );
  INVX1_HVT U415 ( .A(n563), .Y(n548) );
  INVX1_HVT U416 ( .A(n567), .Y(n516) );
  AO21X1_HVT U417 ( .A1(n353), .A2(n390), .A3(n455), .Y(n672) );
  INVX1_HVT U418 ( .A(n565), .Y(n531) );
  NAND2X0_HVT U419 ( .A1(n623), .A2(n402), .Y(n400) );
  NAND2X0_HVT U420 ( .A1(n501), .A2(n477), .Y(n401) );
  NAND2X0_HVT U421 ( .A1(n400), .A2(n401), .Y(n622) );
  NAND2X0_HVT U422 ( .A1(n501), .A2(n402), .Y(n403) );
  NAND2X0_HVT U423 ( .A1(n684), .A2(n477), .Y(n404) );
  NAND2X0_HVT U424 ( .A1(n404), .A2(n403), .Y(n683) );
  NAND2X0_HVT U425 ( .A1(n491), .A2(n493), .Y(n405) );
  NAND2X0_HVT U426 ( .A1(n338), .A2(n399), .Y(n406) );
  NAND2X0_HVT U427 ( .A1(n539), .A2(n408), .Y(n407) );
  NAND2X0_HVT U428 ( .A1(n406), .A2(n407), .Y(n643) );
  MUX41X1_HVT U429 ( .A1(n709), .A3(n719), .A2(n705), .A4(n713), .S0(in[6]), 
        .S1(n427), .Y(out[0]) );
  NAND2X0_HVT U430 ( .A1(n264), .A2(n445), .Y(n409) );
  NAND2X0_HVT U431 ( .A1(n470), .A2(n432), .Y(n410) );
  NAND2X0_HVT U432 ( .A1(n409), .A2(n410), .Y(n581) );
  INVX1_HVT U433 ( .A(in[0]), .Y(n427) );
  MUX21X1_HVT U434 ( .A1(n494), .A2(n458), .S0(n282), .Y(n445) );
  MUX41X1_HVT U435 ( .A1(n412), .A3(n750), .A2(n747), .A4(n525), .S0(n380), 
        .S1(n466), .Y(n411) );
  XNOR2X1_HVT U436 ( .A1(n268), .A2(n553), .Y(n412) );
  MUX21X1_HVT U437 ( .A1(n212), .A2(n492), .S0(n383), .Y(n414) );
  MUX21X1_HVT U438 ( .A1(n689), .A2(n372), .S0(n514), .Y(n597) );
  INVX0_HVT U439 ( .A(n736), .Y(n436) );
  NAND2X0_HVT U440 ( .A1(n480), .A2(n419), .Y(n420) );
  NAND2X0_HVT U441 ( .A1(n422), .A2(n481), .Y(n421) );
  NAND2X0_HVT U442 ( .A1(n420), .A2(n421), .Y(n479) );
  INVX0_HVT U443 ( .A(n481), .Y(n419) );
  NAND2X0_HVT U444 ( .A1(n650), .A2(n428), .Y(n424) );
  NAND2X0_HVT U445 ( .A1(n651), .A2(n213), .Y(n425) );
  NAND2X0_HVT U446 ( .A1(n424), .A2(n425), .Y(n649) );
  INVX1_HVT U447 ( .A(n435), .Y(n588) );
  OR2X1_HVT U448 ( .A1(n383), .A2(n114), .Y(n755) );
  NAND2X0_HVT U449 ( .A1(n475), .A2(n429), .Y(n430) );
  NAND2X0_HVT U450 ( .A1(n675), .A2(n726), .Y(n431) );
  NAND2X0_HVT U451 ( .A1(n431), .A2(n430), .Y(n674) );
  INVX0_HVT U452 ( .A(n726), .Y(n429) );
  NAND2X0_HVT U453 ( .A1(n661), .A2(n213), .Y(n433) );
  NAND2X0_HVT U454 ( .A1(n658), .A2(n428), .Y(n434) );
  NAND2X0_HVT U455 ( .A1(n434), .A2(n433), .Y(n657) );
  MUX41X1_HVT U456 ( .A1(n438), .A3(n437), .A2(n561), .A4(n436), .S0(n485), 
        .S1(n236), .Y(n435) );
  XNOR2X1_HVT U457 ( .A1(n501), .A2(n304), .Y(n438) );
  OR2X1_HVT U458 ( .A1(n322), .A2(n440), .Y(n767) );
  NAND2X0_HVT U459 ( .A1(n461), .A2(n462), .Y(out[5]) );
  NAND2X0_HVT U460 ( .A1(n629), .A2(n320), .Y(n443) );
  NAND2X0_HVT U461 ( .A1(n637), .A2(in[6]), .Y(n444) );
  NAND2X0_HVT U462 ( .A1(n397), .A2(n448), .Y(n449) );
  NAND2X0_HVT U463 ( .A1(n742), .A2(n408), .Y(n450) );
  NAND2X0_HVT U464 ( .A1(n449), .A2(n450), .Y(n633) );
  INVX0_HVT U465 ( .A(n455), .Y(n448) );
  MUX21X1_HVT U466 ( .A1(n492), .A2(n464), .S0(n238), .Y(n742) );
  MUX21X1_HVT U467 ( .A1(n633), .A2(n632), .S0(n17), .Y(n631) );
  INVX1_HVT U468 ( .A(n566), .Y(n539) );
  NAND2X0_HVT U469 ( .A1(n627), .A2(n348), .Y(n459) );
  NAND2X0_HVT U470 ( .A1(n628), .A2(n486), .Y(n460) );
  NAND2X0_HVT U471 ( .A1(n459), .A2(n460), .Y(n625) );
  NAND2X0_HVT U472 ( .A1(n606), .A2(n320), .Y(n461) );
  NAND2X0_HVT U473 ( .A1(n617), .A2(in[6]), .Y(n462) );
  INVX1_HVT U474 ( .A(n568), .Y(n532) );
  INVX1_HVT U475 ( .A(n511), .Y(n510) );
  NBUFFX2_HVT U476 ( .A(n513), .Y(n468) );
  AND2X1_HVT U477 ( .A1(n231), .A2(n717), .Y(n470) );
  MUX21X1_HVT U478 ( .A1(n540), .A2(n342), .S0(n488), .Y(n721) );
  NBUFFX2_HVT U479 ( .A(n763), .Y(n497) );
  AND2X1_HVT U480 ( .A1(n216), .A2(n702), .Y(n471) );
  MUX21X1_HVT U481 ( .A1(n456), .A2(n280), .S0(n453), .Y(n671) );
  MUX21X1_HVT U482 ( .A1(n558), .A2(n457), .S0(n339), .Y(n616) );
  MUX21X1_HVT U483 ( .A1(n369), .A2(n553), .S0(n314), .Y(n565) );
  MUX21X1_HVT U484 ( .A1(n423), .A2(n311), .S0(n304), .Y(n568) );
  MUX21X1_HVT U485 ( .A1(n495), .A2(n520), .S0(n304), .Y(n731) );
  NAND2X0_HVT U486 ( .A1(n491), .A2(n493), .Y(n763) );
  MUX21X1_HVT U487 ( .A1(n540), .A2(n280), .S0(n313), .Y(n566) );
  NBUFFX2_HVT U488 ( .A(n766), .Y(n499) );
  MUX21X1_HVT U489 ( .A1(n492), .A2(n495), .S0(n304), .Y(n656) );
  NBUFFX2_HVT U490 ( .A(n766), .Y(n500) );
  MUX21X1_HVT U491 ( .A1(n501), .A2(n498), .S0(n357), .Y(n564) );
  XOR2X1_HVT U492 ( .A1(n486), .A2(n469), .Y(n726) );
  MUX21X1_HVT U493 ( .A1(n423), .A2(n492), .S0(n304), .Y(n589) );
  NBUFFX2_HVT U494 ( .A(n766), .Y(n501) );
  MUX21X1_HVT U495 ( .A1(n501), .A2(n492), .S0(n314), .Y(n572) );
  AND2X1_HVT U496 ( .A1(n339), .A2(n520), .Y(n474) );
  AND2X1_HVT U497 ( .A1(n337), .A2(n664), .Y(n475) );
  MUX21X1_HVT U498 ( .A1(n338), .A2(n324), .S0(n484), .Y(n653) );
  NBUFFX2_HVT U499 ( .A(n493), .Y(n495) );
  NBUFFX2_HVT U500 ( .A(n510), .Y(n487) );
  MUX21X1_HVT U501 ( .A1(n673), .A2(n516), .S0(n17), .Y(n670) );
  XOR2X1_HVT U502 ( .A1(n313), .A2(n379), .Y(n725) );
  MUX21X1_HVT U503 ( .A1(n532), .A2(n390), .S0(n514), .Y(n628) );
  AND2X1_HVT U504 ( .A1(n456), .A2(n415), .Y(n476) );
  NAND2X0_HVT U505 ( .A1(n547), .A2(n275), .Y(n766) );
  NBUFFX2_HVT U506 ( .A(n767), .Y(n502) );
  XOR2X1_HVT U507 ( .A1(n304), .A2(n487), .Y(n728) );
  MUX21X1_HVT U508 ( .A1(n347), .A2(n353), .S0(n486), .Y(n652) );
  MUX21X1_HVT U509 ( .A1(n372), .A2(n553), .S0(n453), .Y(n569) );
  MUX21X1_HVT U510 ( .A1(n372), .A2(n492), .S0(n514), .Y(n684) );
  NBUFFX2_HVT U511 ( .A(n767), .Y(n503) );
  AND2X1_HVT U512 ( .A1(n495), .A2(n383), .Y(n478) );
  NBUFFX2_HVT U513 ( .A(n510), .Y(n509) );
  MUX41X1_HVT U514 ( .A1(n644), .A3(n657), .A2(n649), .A4(n663), .S0(in[6]), 
        .S1(n489), .Y(out[3]) );
  MUX21X1_HVT U515 ( .A1(n423), .A2(n503), .S0(n297), .Y(n592) );
  MUX21X1_HVT U516 ( .A1(n337), .A2(n500), .S0(n297), .Y(n593) );
  MUX21X1_HVT U517 ( .A1(n439), .A2(n369), .S0(n357), .Y(n571) );
  MUX21X1_HVT U518 ( .A1(n337), .A2(n439), .S0(n312), .Y(n743) );
  MUX21X1_HVT U519 ( .A1(n439), .A2(n503), .S0(n453), .Y(n563) );
  NBUFFX2_HVT U520 ( .A(in[0]), .Y(n489) );
  NBUFFX2_HVT U521 ( .A(n507), .Y(n485) );
  NBUFFX2_HVT U522 ( .A(n507), .Y(n486) );
  XOR2X1_HVT U523 ( .A1(n312), .A2(n232), .Y(n481) );
endmodule

