
module inv_sbox_14 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n46, n177, n196, n197, n198, n199, n201, n202, n203, n205, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656;

  NAND2X0_HVT U1 ( .A1(in[3]), .A2(n359), .Y(n656) );
  NAND2X0_HVT U5 ( .A1(n653), .A2(n368), .Y(n652) );
  NAND2X0_HVT U7 ( .A1(n309), .A2(n371), .Y(n649) );
  NAND2X0_HVT U8 ( .A1(n377), .A2(n368), .Y(n648) );
  NAND2X0_HVT U9 ( .A1(n375), .A2(n648), .Y(n647) );
  NAND2X0_HVT U10 ( .A1(n374), .A2(n645), .Y(n646) );
  NAND2X0_HVT U11 ( .A1(n382), .A2(n373), .Y(n644) );
  NAND2X0_HVT U12 ( .A1(n377), .A2(n356), .Y(n643) );
  NAND2X0_HVT U13 ( .A1(n372), .A2(n648), .Y(n642) );
  NAND2X0_HVT U15 ( .A1(n367), .A2(n309), .Y(n640) );
  NAND2X0_HVT U19 ( .A1(n379), .A2(n448), .Y(n635) );
  NAND2X0_HVT U25 ( .A1(n334), .A2(n357), .Y(n651) );
  NAND2X0_HVT U32 ( .A1(n359), .A2(n382), .Y(n623) );
  NAND2X0_HVT U35 ( .A1(n648), .A2(n449), .Y(n620) );
  NAND2X0_HVT U38 ( .A1(n356), .A2(n382), .Y(n617) );
  OA21X1_HVT U53 ( .A1(n390), .A2(n606), .A3(n417), .Y(n604) );
  NAND2X0_HVT U55 ( .A1(n372), .A2(n653), .Y(n602) );
  MUX41X1_HVT U65 ( .A1(n408), .A3(n410), .A2(n409), .A4(n617), .S0(n349), 
        .S1(n325), .Y(n591) );
  NAND2X0_HVT U66 ( .A1(n379), .A2(n263), .Y(n590) );
  MUX41X1_HVT U67 ( .A1(n405), .A3(n431), .A2(n407), .A4(n590), .S0(n354), 
        .S1(n346), .Y(n589) );
  MUX41X1_HVT U68 ( .A1(n405), .A3(n327), .A2(n406), .A4(n375), .S0(n348), 
        .S1(n305), .Y(n588) );
  NAND2X0_HVT U72 ( .A1(n367), .A2(n649), .Y(n585) );
  MUX41X1_HVT U73 ( .A1(n628), .A3(n585), .A2(n240), .A4(n355), .S0(n295), 
        .S1(n345), .Y(n584) );
  MUX41X1_HVT U74 ( .A1(n646), .A3(n422), .A2(n421), .A4(n411), .S0(n349), 
        .S1(n325), .Y(n583) );
  MUX41X1_HVT U78 ( .A1(n580), .A3(n584), .A2(n583), .A4(n586), .S0(in[5]), 
        .S1(n328), .Y(n579) );
  NAND2X0_HVT U81 ( .A1(n373), .A2(n649), .Y(n576) );
  AND2X1_HVT U82 ( .A1(n650), .A2(n370), .Y(n575) );
  MUX41X1_HVT U83 ( .A1(n575), .A3(n419), .A2(n434), .A4(n576), .S0(n348), 
        .S1(n325), .Y(n574) );
  MUX41X1_HVT U84 ( .A1(n340), .A3(n418), .A2(n435), .A4(n630), .S0(n349), 
        .S1(n387), .Y(n573) );
  MUX41X1_HVT U85 ( .A1(n573), .A3(n577), .A2(n574), .A4(n578), .S0(n365), 
        .S1(n328), .Y(n572) );
  MUX41X1_HVT U88 ( .A1(n407), .A3(n393), .A2(n625), .A4(n610), .S0(n348), 
        .S1(n295), .Y(n570) );
  NAND2X0_HVT U89 ( .A1(n382), .A2(n446), .Y(n569) );
  MUX41X1_HVT U90 ( .A1(n343), .A3(n649), .A2(n609), .A4(n569), .S0(n348), 
        .S1(n387), .Y(n568) );
  MUX41X1_HVT U96 ( .A1(n431), .A3(n642), .A2(n416), .A4(n437), .S0(n349), 
        .S1(n385), .Y(n562) );
  MUX41X1_HVT U99 ( .A1(n623), .A3(n409), .A2(n608), .A4(n277), .S0(n387), 
        .S1(n346), .Y(n559) );
  NAND2X0_HVT U100 ( .A1(n382), .A2(n445), .Y(n558) );
  MUX41X1_HVT U101 ( .A1(n439), .A3(n643), .A2(n423), .A4(n558), .S0(n387), 
        .S1(n346), .Y(n557) );
  AND2X1_HVT U104 ( .A1(n649), .A2(n368), .Y(n555) );
  MUX41X1_HVT U105 ( .A1(n641), .A3(n440), .A2(n576), .A4(n555), .S0(n349), 
        .S1(n385), .Y(n554) );
  MUX41X1_HVT U107 ( .A1(n439), .A3(n370), .A2(n553), .A4(n238), .S0(n348), 
        .S1(n387), .Y(n552) );
  MUX41X1_HVT U108 ( .A1(n248), .A3(n277), .A2(n415), .A4(n373), .S0(n349), 
        .S1(n386), .Y(n551) );
  MUX41X1_HVT U109 ( .A1(n438), .A3(n393), .A2(n435), .A4(n429), .S0(n348), 
        .S1(n387), .Y(n550) );
  AO21X1_HVT U112 ( .A1(n426), .A2(n305), .A3(n631), .Y(n547) );
  NAND2X0_HVT U114 ( .A1(n375), .A2(n649), .Y(n545) );
  MUX41X1_HVT U115 ( .A1(n545), .A3(n644), .A2(n426), .A4(n370), .S0(n325), 
        .S1(n346), .Y(n544) );
  MUX41X1_HVT U116 ( .A1(n425), .A3(n418), .A2(n393), .A4(n640), .S0(n347), 
        .S1(n295), .Y(n543) );
  NAND2X0_HVT U118 ( .A1(n382), .A2(n327), .Y(n541) );
  MUX41X1_HVT U119 ( .A1(n441), .A3(n542), .A2(n618), .A4(n541), .S0(n347), 
        .S1(n325), .Y(n540) );
  MUX41X1_HVT U120 ( .A1(n540), .A3(n544), .A2(n543), .A4(n546), .S0(n365), 
        .S1(n363), .Y(n539) );
  MUX41X1_HVT U122 ( .A1(n430), .A3(n337), .A2(n610), .A4(n432), .S0(n347), 
        .S1(n386), .Y(n538) );
  MUX41X1_HVT U124 ( .A1(n338), .A3(n537), .A2(n632), .A4(n265), .S0(n353), 
        .S1(n347), .Y(n536) );
  AOI21X1_HVT U127 ( .A1(n352), .A2(n532), .A3(n399), .Y(n533) );
  NAND2X0_HVT U129 ( .A1(n351), .A2(n374), .Y(n530) );
  MUX41X1_HVT U130 ( .A1(n530), .A3(n531), .A2(n534), .A4(n533), .S0(n354), 
        .S1(n363), .Y(n529) );
  AND2X1_HVT U131 ( .A1(n263), .A2(n290), .Y(n528) );
  MUX41X1_HVT U132 ( .A1(n398), .A3(n528), .A2(n443), .A4(n405), .S0(n387), 
        .S1(n345), .Y(n527) );
  MUX41X1_HVT U133 ( .A1(n444), .A3(n342), .A2(n246), .A4(n235), .S0(n353), 
        .S1(n346), .Y(n526) );
  MUX41X1_HVT U136 ( .A1(n607), .A3(n558), .A2(n524), .A4(n403), .S0(n351), 
        .S1(n325), .Y(n523) );
  MUX41X1_HVT U137 ( .A1(n269), .A3(n626), .A2(n630), .A4(n437), .S0(n354), 
        .S1(n345), .Y(n522) );
  MUX41X1_HVT U139 ( .A1(n521), .A3(n525), .A2(n529), .A4(n535), .S0(n365), 
        .S1(n326), .Y(out[4]) );
  NAND2X0_HVT U141 ( .A1(n367), .A2(n382), .Y(n519) );
  MUX41X1_HVT U142 ( .A1(n519), .A3(n616), .A2(n442), .A4(n414), .S0(n352), 
        .S1(n385), .Y(n518) );
  MUX41X1_HVT U145 ( .A1(n624), .A3(n440), .A2(n516), .A4(n576), .S0(n352), 
        .S1(n387), .Y(n515) );
  MUX41X1_HVT U146 ( .A1(n515), .A3(n517), .A2(n518), .A4(n520), .S0(n362), 
        .S1(in[5]), .Y(n514) );
  MUX41X1_HVT U151 ( .A1(n434), .A3(n424), .A2(n412), .A4(n510), .S0(n353), 
        .S1(n345), .Y(n509) );
  MUX41X1_HVT U155 ( .A1(n414), .A3(n644), .A2(n636), .A4(n416), .S0(n350), 
        .S1(n386), .Y(n505) );
  NAND2X0_HVT U159 ( .A1(n501), .A2(n500), .Y(n502) );
  MUX41X1_HVT U162 ( .A1(n332), .A3(n410), .A2(n620), .A4(n498), .S0(n350), 
        .S1(n386), .Y(n497) );
  NAND2X0_HVT U163 ( .A1(n310), .A2(n446), .Y(n496) );
  MUX41X1_HVT U164 ( .A1(n647), .A3(n496), .A2(n618), .A4(n411), .S0(n347), 
        .S1(n385), .Y(n495) );
  NAND2X0_HVT U166 ( .A1(n645), .A2(n492), .Y(n493) );
  MUX41X1_HVT U170 ( .A1(n396), .A3(n336), .A2(n338), .A4(n489), .S0(n350), 
        .S1(n295), .Y(n488) );
  MUX41X1_HVT U172 ( .A1(n569), .A3(n487), .A2(n336), .A4(n633), .S0(n350), 
        .S1(n295), .Y(n486) );
  NAND2X0_HVT U177 ( .A1(n377), .A2(n327), .Y(n482) );
  AND2X1_HVT U179 ( .A1(n650), .A2(n369), .Y(n481) );
  MUX41X1_HVT U180 ( .A1(n623), .A3(n391), .A2(n481), .A4(n611), .S0(n350), 
        .S1(n386), .Y(n480) );
  AND2X1_HVT U185 ( .A1(n276), .A2(n290), .Y(n475) );
  OA21X1_HVT U189 ( .A1(n390), .A2(n418), .A3(n596), .Y(n471) );
  MUX41X1_HVT U190 ( .A1(n472), .A3(n473), .A2(n471), .A4(n474), .S0(n362), 
        .S1(n345), .Y(n470) );
  AND2X1_HVT U192 ( .A1(n422), .A2(n467), .Y(n468) );
  NAND2X0_HVT U194 ( .A1(n613), .A2(n467), .Y(n465) );
  NAND2X0_HVT U198 ( .A1(n379), .A2(n449), .Y(n645) );
  NAND2X0_HVT U200 ( .A1(n369), .A2(n382), .Y(n532) );
  NAND2X0_HVT U203 ( .A1(n448), .A2(n382), .Y(n463) );
  NAND2X0_HVT U207 ( .A1(n382), .A2(n343), .Y(n596) );
  INVX2_HVT U2 ( .A(n634), .Y(n411) );
  MUX21X1_HVT U3 ( .A1(n598), .A2(n597), .S0(n351), .Y(n595) );
  MUX21X1_HVT U4 ( .A1(n265), .A2(n602), .S0(n386), .Y(n598) );
  MUX21X1_HVT U6 ( .A1(n655), .A2(n266), .S0(n378), .Y(n265) );
  INVX1_HVT U14 ( .A(n381), .Y(n378) );
  NAND2X0_HVT U16 ( .A1(n502), .A2(n46), .Y(n177) );
  NAND2X0_HVT U17 ( .A1(n503), .A2(n352), .Y(n196) );
  NAND2X0_HVT U18 ( .A1(n177), .A2(n196), .Y(n499) );
  IBUFFX2_HVT U20 ( .A(n352), .Y(n46) );
  MUX21X1_HVT U21 ( .A1(n612), .A2(n432), .S0(n305), .Y(n503) );
  MUX41X1_HVT U22 ( .A1(n414), .A3(n644), .A2(n421), .A4(n339), .S0(n325), 
        .S1(n197), .Y(n520) );
  IBUFFX16_HVT U23 ( .A(n346), .Y(n197) );
  IBUFFX32_HVT U24 ( .A(n235), .Y(n650) );
  NOR2X4_HVT U26 ( .A1(n367), .A2(n235), .Y(n342) );
  INVX1_HVT U27 ( .A(n656), .Y(n343) );
  NAND2X0_HVT U28 ( .A1(n413), .A2(n198), .Y(n199) );
  NAND2X0_HVT U29 ( .A1(n600), .A2(n341), .Y(n201) );
  NAND2X0_HVT U30 ( .A1(n199), .A2(n201), .Y(n599) );
  IBUFFX2_HVT U31 ( .A(n341), .Y(n198) );
  NAND2X0_HVT U33 ( .A1(n360), .A2(n202), .Y(n203) );
  NAND2X0_HVT U34 ( .A1(n366), .A2(n250), .Y(n205) );
  NAND2X0_HVT U36 ( .A1(n203), .A2(n205), .Y(n630) );
  INVX0_HVT U37 ( .A(n250), .Y(n202) );
  MUX21X1_HVT U39 ( .A1(n414), .A2(n652), .S0(n352), .Y(n600) );
  DELLN1X2_HVT U40 ( .A(n333), .Y(n360) );
  INVX1_HVT U41 ( .A(n289), .Y(n250) );
  INVX1_HVT U42 ( .A(n630), .Y(n414) );
  MUX21X2_HVT U43 ( .A1(n367), .A2(n343), .S0(n309), .Y(n624) );
  NAND2X0_HVT U44 ( .A1(n604), .A2(n218), .Y(n219) );
  NAND2X0_HVT U45 ( .A1(n605), .A2(n271), .Y(n220) );
  NAND2X0_HVT U46 ( .A1(n219), .A2(n220), .Y(n603) );
  INVX0_HVT U47 ( .A(n271), .Y(n218) );
  MUX21X1_HVT U48 ( .A1(n236), .A2(n406), .S0(n354), .Y(n605) );
  IBUFFX2_HVT U49 ( .A(n351), .Y(n271) );
  NAND2X0_HVT U50 ( .A1(n355), .A2(n358), .Y(n329) );
  IBUFFX2_HVT U51 ( .A(n389), .Y(n387) );
  INVX0_HVT U52 ( .A(n389), .Y(n388) );
  INVX0_HVT U54 ( .A(n639), .Y(n449) );
  IBUFFX2_HVT U56 ( .A(n327), .Y(n266) );
  INVX1_HVT U57 ( .A(n296), .Y(n228) );
  INVX2_HVT U58 ( .A(n376), .Y(n382) );
  NAND2X0_HVT U59 ( .A1(n248), .A2(n221), .Y(n222) );
  NAND2X0_HVT U60 ( .A1(n593), .A2(n341), .Y(n223) );
  NAND2X0_HVT U61 ( .A1(n222), .A2(n223), .Y(n592) );
  INVX0_HVT U62 ( .A(n341), .Y(n221) );
  MUX21X1_HVT U63 ( .A1(n653), .A2(n412), .S0(n282), .Y(n593) );
  INVX0_HVT U64 ( .A(n633), .Y(n412) );
  MUX21X2_HVT U69 ( .A1(n507), .A2(n508), .S0(n352), .Y(n506) );
  INVX1_HVT U70 ( .A(n290), .Y(n376) );
  MUX41X1_HVT U71 ( .A1(n476), .A3(n464), .A2(n479), .A4(n470), .S0(n251), 
        .S1(n224), .Y(out[7]) );
  IBUFFX16_HVT U75 ( .A(n364), .Y(n224) );
  IBUFFX2_HVT U76 ( .A(n265), .Y(n632) );
  IBUFFX16_HVT U77 ( .A(n389), .Y(n305) );
  INVX0_HVT U79 ( .A(n325), .Y(n268) );
  IBUFFX16_HVT U80 ( .A(n389), .Y(n325) );
  OA21X1_HVT U86 ( .A1(n394), .A2(n390), .A3(n402), .Y(n507) );
  NAND2X0_HVT U87 ( .A1(n493), .A2(n225), .Y(n226) );
  NAND2X0_HVT U91 ( .A1(n494), .A2(n351), .Y(n227) );
  NAND2X0_HVT U92 ( .A1(n226), .A2(n227), .Y(n491) );
  IBUFFX2_HVT U93 ( .A(n351), .Y(n225) );
  MUX21X1_HVT U94 ( .A1(n629), .A2(n632), .S0(n353), .Y(n494) );
  MUX41X1_HVT U95 ( .A1(n506), .A3(n511), .A2(n505), .A4(n509), .S0(n365), 
        .S1(n228), .Y(n504) );
  MUX21X1_HVT U97 ( .A1(n374), .A2(n230), .S0(n380), .Y(n229) );
  IBUFFX16_HVT U98 ( .A(n229), .Y(n489) );
  IBUFFX16_HVT U102 ( .A(n448), .Y(n230) );
  NAND2X0_HVT U103 ( .A1(n376), .A2(n655), .Y(n653) );
  MUX41X1_HVT U106 ( .A1(n277), .A3(n267), .A2(n246), .A4(n415), .S0(n231), 
        .S1(n305), .Y(n601) );
  IBUFFX16_HVT U110 ( .A(n349), .Y(n231) );
  NAND2X0_HVT U111 ( .A1(n240), .A2(n232), .Y(n233) );
  NAND2X0_HVT U113 ( .A1(n614), .A2(n305), .Y(n234) );
  NAND2X0_HVT U117 ( .A1(n233), .A2(n234), .Y(n472) );
  INVX0_HVT U121 ( .A(n305), .Y(n232) );
  AND2X1_HVT U123 ( .A1(n289), .A2(n375), .Y(n235) );
  INVX0_HVT U125 ( .A(n628), .Y(n236) );
  INVX1_HVT U126 ( .A(n250), .Y(n237) );
  INVX0_HVT U128 ( .A(n628), .Y(n416) );
  INVX0_HVT U134 ( .A(n613), .Y(n238) );
  INVX1_HVT U135 ( .A(n342), .Y(n613) );
  INVX0_HVT U138 ( .A(n359), .Y(n241) );
  INVX1_HVT U140 ( .A(n245), .Y(n246) );
  INVX2_HVT U143 ( .A(n289), .Y(n290) );
  MUX21X2_HVT U144 ( .A1(n512), .A2(n513), .S0(n239), .Y(n511) );
  IBUFFX16_HVT U147 ( .A(n351), .Y(n239) );
  MUX21X1_HVT U148 ( .A1(n343), .A2(n446), .S0(n319), .Y(n627) );
  MUX21X1_HVT U149 ( .A1(n329), .A2(n241), .S0(n309), .Y(n240) );
  NAND2X0_HVT U150 ( .A1(n340), .A2(n242), .Y(n243) );
  NAND2X0_HVT U152 ( .A1(n608), .A2(n354), .Y(n244) );
  NAND2X0_HVT U153 ( .A1(n243), .A2(n244), .Y(n473) );
  IBUFFX2_HVT U154 ( .A(n354), .Y(n242) );
  NBUFFX4_HVT U156 ( .A(n388), .Y(n354) );
  INVX1_HVT U157 ( .A(n319), .Y(n288) );
  MUX21X2_HVT U158 ( .A1(n356), .A2(n367), .S0(n258), .Y(n634) );
  IBUFFX2_HVT U160 ( .A(n379), .Y(n258) );
  IBUFFX2_HVT U161 ( .A(n653), .Y(n397) );
  INVX0_HVT U165 ( .A(n602), .Y(n245) );
  INVX0_HVT U167 ( .A(n411), .Y(n247) );
  INVX0_HVT U168 ( .A(n247), .Y(n248) );
  NBUFFX2_HVT U169 ( .A(n639), .Y(n249) );
  NBUFFX2_HVT U171 ( .A(n249), .Y(n277) );
  IBUFFX16_HVT U173 ( .A(n278), .Y(n251) );
  NBUFFX4_HVT U174 ( .A(n447), .Y(n357) );
  MUX41X1_HVT U175 ( .A1(n495), .A3(n499), .A2(n491), .A4(n497), .S0(n252), 
        .S1(n253), .Y(n490) );
  IBUFFX16_HVT U176 ( .A(n364), .Y(n252) );
  IBUFFX16_HVT U178 ( .A(n328), .Y(n253) );
  MUX41X1_HVT U181 ( .A1(n411), .A3(n613), .A2(n427), .A4(n267), .S0(n254), 
        .S1(n274), .Y(n477) );
  IBUFFX16_HVT U182 ( .A(n273), .Y(n254) );
  MUX21X1_HVT U183 ( .A1(n432), .A2(n392), .S0(n354), .Y(n582) );
  OA21X1_HVT U184 ( .A1(n395), .A2(n390), .A3(n634), .Y(n581) );
  INVX0_HVT U186 ( .A(n358), .Y(n287) );
  NAND2X0_HVT U187 ( .A1(n340), .A2(n255), .Y(n256) );
  NAND2X0_HVT U188 ( .A1(n630), .A2(n261), .Y(n257) );
  NAND2X0_HVT U191 ( .A1(n256), .A2(n257), .Y(n508) );
  INVX0_HVT U193 ( .A(n261), .Y(n255) );
  IBUFFX2_HVT U195 ( .A(n305), .Y(n261) );
  INVX1_HVT U196 ( .A(n290), .Y(n310) );
  MUX41X1_HVT U197 ( .A1(n484), .A3(n485), .A2(n486), .A4(n488), .S0(n259), 
        .S1(n260), .Y(n483) );
  IBUFFX16_HVT U199 ( .A(n304), .Y(n259) );
  IBUFFX16_HVT U201 ( .A(n364), .Y(n260) );
  INVX0_HVT U202 ( .A(n334), .Y(n262) );
  INVX1_HVT U204 ( .A(n262), .Y(n263) );
  INVX0_HVT U205 ( .A(n333), .Y(n334) );
  OR2X2_HVT U206 ( .A1(n447), .A2(n333), .Y(n654) );
  MUX41X1_HVT U208 ( .A1(n343), .A3(n650), .A2(n401), .A4(n644), .S0(n264), 
        .S1(n305), .Y(n586) );
  IBUFFX16_HVT U209 ( .A(n348), .Y(n264) );
  MUX21X1_HVT U210 ( .A1(n602), .A2(n436), .S0(n317), .Y(n302) );
  INVX1_HVT U211 ( .A(n368), .Y(n446) );
  AO21X1_HVT U212 ( .A1(n249), .A2(n653), .A3(n390), .Y(n492) );
  MUX21X1_HVT U213 ( .A1(n651), .A2(n333), .S0(n290), .Y(n267) );
  MUX41X1_HVT U214 ( .A1(n652), .A3(n647), .A2(n267), .A4(n433), .S0(n272), 
        .S1(n268), .Y(n577) );
  INVX1_HVT U215 ( .A(n290), .Y(n380) );
  MUX21X2_HVT U216 ( .A1(n556), .A2(n563), .S0(n326), .Y(out[2]) );
  INVX1_HVT U217 ( .A(n307), .Y(n293) );
  MUX21X1_HVT U218 ( .A1(n375), .A2(n332), .S0(n308), .Y(n307) );
  MUX21X1_HVT U219 ( .A1(n369), .A2(n374), .S0(n377), .Y(n332) );
  IBUFFX2_HVT U220 ( .A(n297), .Y(n278) );
  INVX0_HVT U221 ( .A(n400), .Y(n269) );
  MUX41X1_HVT U222 ( .A1(n465), .A3(n469), .A2(n466), .A4(n468), .S0(n362), 
        .S1(n270), .Y(n464) );
  IBUFFX16_HVT U223 ( .A(n348), .Y(n270) );
  NAND2X1_HVT U224 ( .A1(n390), .A2(n404), .Y(n469) );
  INVX1_HVT U225 ( .A(n353), .Y(n273) );
  INVX0_HVT U226 ( .A(n286), .Y(n510) );
  IBUFFX16_HVT U227 ( .A(n348), .Y(n272) );
  MUX21X2_HVT U228 ( .A1(n539), .A2(n549), .S0(n326), .Y(out[3]) );
  IBUFFX16_HVT U229 ( .A(n345), .Y(n274) );
  MUX41X1_HVT U230 ( .A1(n599), .A3(n603), .A2(n595), .A4(n601), .S0(n365), 
        .S1(n275), .Y(n594) );
  IBUFFX16_HVT U231 ( .A(n328), .Y(n275) );
  INVX0_HVT U232 ( .A(n249), .Y(n276) );
  INVX0_HVT U233 ( .A(n619), .Y(n423) );
  MUX21X1_HVT U234 ( .A1(n582), .A2(n581), .S0(n352), .Y(n580) );
  INVX1_HVT U235 ( .A(n385), .Y(n284) );
  INVX1_HVT U236 ( .A(in[3]), .Y(n447) );
  NAND2X0_HVT U237 ( .A1(n371), .A2(n279), .Y(n280) );
  NAND2X0_HVT U238 ( .A1(n567), .A2(n285), .Y(n281) );
  NAND2X0_HVT U239 ( .A1(n280), .A2(n281), .Y(n566) );
  INVX0_HVT U240 ( .A(n285), .Y(n279) );
  NBUFFX4_HVT U241 ( .A(n654), .Y(n371) );
  IBUFFX2_HVT U242 ( .A(n380), .Y(n285) );
  IBUFFX16_HVT U243 ( .A(n351), .Y(n282) );
  MUX41X1_HVT U244 ( .A1(n627), .A3(n424), .A2(n438), .A4(n561), .S0(n283), 
        .S1(n284), .Y(n560) );
  IBUFFX16_HVT U245 ( .A(n349), .Y(n283) );
  MUX21X1_HVT U246 ( .A1(n368), .A2(n287), .S0(n288), .Y(n286) );
  INVX1_HVT U247 ( .A(in[6]), .Y(n333) );
  AO21X2_HVT U248 ( .A1(n377), .A2(n445), .A3(n389), .Y(n467) );
  IBUFFX2_HVT U249 ( .A(n388), .Y(n335) );
  IBUFFX2_HVT U250 ( .A(n447), .Y(n327) );
  INVX1_HVT U251 ( .A(n381), .Y(n289) );
  INVX1_HVT U252 ( .A(in[0]), .Y(n381) );
  INVX1_HVT U253 ( .A(n291), .Y(n614) );
  AO21X1_HVT U254 ( .A1(n354), .A2(n400), .A3(n445), .Y(n512) );
  XNOR2X1_HVT U255 ( .A1(n369), .A2(n380), .Y(n311) );
  MUX21X2_HVT U256 ( .A1(n302), .A2(n303), .S0(n295), .Y(n484) );
  MUX21X1_HVT U257 ( .A1(n333), .A2(n370), .S0(n380), .Y(n291) );
  INVX1_HVT U258 ( .A(n370), .Y(n448) );
  IBUFFX2_HVT U259 ( .A(n389), .Y(n386) );
  IBUFFX2_HVT U260 ( .A(n389), .Y(n385) );
  IBUFFX2_HVT U261 ( .A(n389), .Y(n295) );
  MUX21X1_HVT U262 ( .A1(n294), .A2(n293), .S0(n385), .Y(n292) );
  IBUFFX16_HVT U263 ( .A(n306), .Y(n294) );
  NBUFFX2_HVT U264 ( .A(in[7]), .Y(n326) );
  INVX0_HVT U265 ( .A(n362), .Y(n304) );
  INVX1_HVT U266 ( .A(n317), .Y(n308) );
  AO21X1_HVT U267 ( .A1(n596), .A2(n353), .A3(n634), .Y(n597) );
  INVX1_HVT U268 ( .A(n313), .Y(n296) );
  MUX41X1_HVT U269 ( .A1(n415), .A3(n436), .A2(n340), .A4(n397), .S0(n312), 
        .S1(n390), .Y(n571) );
  NAND2X0_HVT U270 ( .A1(n565), .A2(n312), .Y(n300) );
  INVX1_HVT U271 ( .A(n364), .Y(n365) );
  INVX1_HVT U272 ( .A(n318), .Y(n314) );
  INVX0_HVT U273 ( .A(n349), .Y(n312) );
  NBUFFX2_HVT U274 ( .A(n388), .Y(n353) );
  INVX0_HVT U275 ( .A(n326), .Y(n297) );
  INVX1_HVT U276 ( .A(n363), .Y(n313) );
  INVX0_HVT U277 ( .A(in[1]), .Y(n361) );
  INVX1_HVT U278 ( .A(n350), .Y(n317) );
  INVX1_HVT U279 ( .A(in[5]), .Y(n364) );
  INVX1_HVT U280 ( .A(n461), .Y(n432) );
  MUX41X1_HVT U281 ( .A1(n554), .A3(n551), .A2(n552), .A4(n550), .S0(n364), 
        .S1(n314), .Y(n549) );
  NAND2X0_HVT U282 ( .A1(n483), .A2(n297), .Y(n298) );
  NAND2X0_HVT U283 ( .A1(n490), .A2(n326), .Y(n299) );
  NAND2X0_HVT U284 ( .A1(n298), .A2(n299), .Y(out[6]) );
  INVX0_HVT U285 ( .A(n381), .Y(n379) );
  IBUFFX2_HVT U286 ( .A(n381), .Y(n377) );
  INVX1_HVT U287 ( .A(n311), .Y(n608) );
  MUX41X1_HVT U288 ( .A1(n564), .A3(n568), .A2(n570), .A4(n571), .S0(n328), 
        .S1(n365), .Y(n563) );
  NAND2X0_HVT U289 ( .A1(n566), .A2(n351), .Y(n301) );
  NAND2X0_HVT U290 ( .A1(n300), .A2(n301), .Y(n564) );
  INVX1_HVT U291 ( .A(in[4]), .Y(n389) );
  MUX21X1_HVT U292 ( .A1(n276), .A2(n444), .S0(n317), .Y(n303) );
  MUX21X1_HVT U293 ( .A1(n463), .A2(n344), .S0(n308), .Y(n306) );
  IBUFFX2_HVT U294 ( .A(n381), .Y(n309) );
  MUX41X1_HVT U295 ( .A1(n638), .A3(n420), .A2(n637), .A4(n418), .S0(n312), 
        .S1(n390), .Y(n578) );
  IBUFFX2_HVT U296 ( .A(n638), .Y(n407) );
  INVX1_HVT U297 ( .A(n626), .Y(n418) );
  NAND2X0_HVT U298 ( .A1(n480), .A2(n314), .Y(n315) );
  NAND2X0_HVT U299 ( .A1(n292), .A2(n318), .Y(n316) );
  NAND2X0_HVT U300 ( .A1(n315), .A2(n316), .Y(n479) );
  INVX0_HVT U301 ( .A(n313), .Y(n318) );
  AO21X2_HVT U302 ( .A1(n290), .A2(n374), .A3(n390), .Y(n500) );
  IBUFFX2_HVT U303 ( .A(n381), .Y(n319) );
  NAND2X0_HVT U304 ( .A1(n477), .A2(n320), .Y(n321) );
  NAND2X0_HVT U305 ( .A1(n478), .A2(n362), .Y(n322) );
  NAND2X0_HVT U306 ( .A1(n321), .A2(n322), .Y(n476) );
  IBUFFX2_HVT U307 ( .A(n362), .Y(n320) );
  INVX1_HVT U308 ( .A(n361), .Y(n362) );
  NAND2X0_HVT U309 ( .A1(n475), .A2(n390), .Y(n323) );
  NAND2X0_HVT U310 ( .A1(n433), .A2(n353), .Y(n324) );
  NAND2X0_HVT U311 ( .A1(n323), .A2(n324), .Y(n474) );
  INVX1_HVT U312 ( .A(n460), .Y(n433) );
  IBUFFX2_HVT U313 ( .A(in[4]), .Y(n390) );
  MUX21X2_HVT U314 ( .A1(n504), .A2(n514), .S0(n326), .Y(out[5]) );
  MUX41X1_HVT U315 ( .A1(n562), .A3(n559), .A2(n560), .A4(n557), .S0(n364), 
        .S1(n313), .Y(n556) );
  NBUFFX2_HVT U316 ( .A(n447), .Y(n355) );
  NAND2X0_HVT U317 ( .A1(n443), .A2(n335), .Y(n330) );
  MUX21X1_HVT U318 ( .A1(n358), .A2(n449), .S0(n319), .Y(n619) );
  INVX0_HVT U319 ( .A(n361), .Y(n328) );
  MUX41X1_HVT U320 ( .A1(n592), .A3(n589), .A2(n591), .A4(n588), .S0(n364), 
        .S1(n314), .Y(n587) );
  MUX41X1_HVT U321 ( .A1(n434), .A3(n397), .A2(n653), .A4(n342), .S0(n312), 
        .S1(n335), .Y(n478) );
  XNOR2X2_HVT U322 ( .A1(n358), .A2(n357), .Y(n639) );
  MUX21X1_HVT U323 ( .A1(n449), .A2(n445), .S0(n377), .Y(n633) );
  MUX41X1_HVT U324 ( .A1(n632), .A3(n635), .A2(n427), .A4(n446), .S0(n312), 
        .S1(n335), .Y(n517) );
  NAND2X0_HVT U325 ( .A1(n398), .A2(n353), .Y(n331) );
  NAND2X0_HVT U326 ( .A1(n330), .A2(n331), .Y(n513) );
  MUX41X1_HVT U327 ( .A1(n619), .A3(n373), .A2(n343), .A4(n375), .S0(n317), 
        .S1(n335), .Y(n485) );
  INVX0_HVT U328 ( .A(n463), .Y(n396) );
  MUX21X2_HVT U329 ( .A1(n587), .A2(n594), .S0(n326), .Y(out[0]) );
  MUX21X2_HVT U330 ( .A1(n572), .A2(n579), .S0(n326), .Y(out[1]) );
  MUX21X2_HVT U331 ( .A1(n522), .A2(n523), .S0(n362), .Y(n521) );
  MUX21X2_HVT U332 ( .A1(n526), .A2(n527), .S0(n363), .Y(n525) );
  INVX1_HVT U333 ( .A(n655), .Y(n445) );
  MUX21X1_HVT U334 ( .A1(n428), .A2(n338), .S0(n353), .Y(n466) );
  AND2X1_HVT U335 ( .A1(n650), .A2(n329), .Y(n336) );
  AND2X1_HVT U336 ( .A1(n329), .A2(n640), .Y(n337) );
  MUX21X1_HVT U337 ( .A1(n359), .A2(n445), .S0(n319), .Y(n629) );
  MUX21X1_HVT U338 ( .A1(n356), .A2(n448), .S0(n377), .Y(n612) );
  MUX21X1_HVT U339 ( .A1(n401), .A2(n249), .S0(n354), .Y(n565) );
  MUX21X1_HVT U340 ( .A1(n367), .A2(n360), .S0(n305), .Y(n567) );
  MUX21X1_HVT U341 ( .A1(n368), .A2(n371), .S0(n379), .Y(n498) );
  MUX21X1_HVT U342 ( .A1(n448), .A2(n356), .S0(n309), .Y(n461) );
  MUX21X1_HVT U343 ( .A1(n357), .A2(n445), .S0(n379), .Y(n625) );
  MUX21X1_HVT U344 ( .A1(n445), .A2(n448), .S0(n377), .Y(n606) );
  MUX21X1_HVT U345 ( .A1(n442), .A2(n339), .S0(n351), .Y(n534) );
  MUX21X1_HVT U346 ( .A1(n622), .A2(n337), .S0(n352), .Y(n531) );
  MUX21X1_HVT U347 ( .A1(n368), .A2(n373), .S0(n378), .Y(n451) );
  MUX21X1_HVT U348 ( .A1(n356), .A2(n329), .S0(n380), .Y(n460) );
  AND2X1_HVT U349 ( .A1(n310), .A2(n360), .Y(n338) );
  MUX21X1_HVT U350 ( .A1(n372), .A2(n329), .S0(n378), .Y(n637) );
  XNOR2X1_HVT U351 ( .A1(n329), .A2(n310), .Y(n339) );
  MUX21X1_HVT U352 ( .A1(n371), .A2(n357), .S0(n309), .Y(n636) );
  MUX21X1_HVT U353 ( .A1(n357), .A2(n359), .S0(n319), .Y(n611) );
  XOR2X1_HVT U354 ( .A1(n370), .A2(n319), .Y(n609) );
  MUX21X1_HVT U355 ( .A1(n355), .A2(n371), .S0(n309), .Y(n454) );
  NBUFFX2_HVT U356 ( .A(n651), .Y(n368) );
  NBUFFX2_HVT U357 ( .A(n654), .Y(n370) );
  AND2X1_HVT U358 ( .A1(n372), .A2(n382), .Y(n340) );
  MUX21X1_HVT U359 ( .A1(n536), .A2(n538), .S0(n362), .Y(n535) );
  MUX21X1_HVT U360 ( .A1(n372), .A2(n359), .S0(n380), .Y(n537) );
  MUX21X1_HVT U361 ( .A1(n329), .A2(n369), .S0(n319), .Y(n516) );
  NBUFFX2_HVT U362 ( .A(n654), .Y(n372) );
  MUX21X1_HVT U363 ( .A1(n547), .A2(n548), .S0(n352), .Y(n546) );
  MUX21X1_HVT U364 ( .A1(n399), .A2(n614), .S0(n354), .Y(n548) );
  NBUFFX2_HVT U365 ( .A(n651), .Y(n369) );
  NBUFFX2_HVT U366 ( .A(n447), .Y(n356) );
  NBUFFX2_HVT U367 ( .A(n384), .Y(n350) );
  NBUFFX2_HVT U368 ( .A(n383), .Y(n352) );
  NBUFFX2_HVT U369 ( .A(n383), .Y(n351) );
  XNOR2X1_HVT U370 ( .A1(n390), .A2(n347), .Y(n341) );
  NBUFFX2_HVT U371 ( .A(n384), .Y(n347) );
  NBUFFX2_HVT U372 ( .A(n383), .Y(n345) );
  NBUFFX2_HVT U373 ( .A(n384), .Y(n348) );
  NBUFFX2_HVT U374 ( .A(n384), .Y(n349) );
  NBUFFX2_HVT U375 ( .A(n383), .Y(n346) );
  INVX1_HVT U376 ( .A(n361), .Y(n363) );
  MUX21X1_HVT U377 ( .A1(n360), .A2(n327), .S0(n376), .Y(n628) );
  INVX0_HVT U378 ( .A(n482), .Y(n344) );
  MUX21X1_HVT U379 ( .A1(n375), .A2(n327), .S0(n379), .Y(n501) );
  MUX21X1_HVT U380 ( .A1(n368), .A2(n327), .S0(n310), .Y(n561) );
  MUX21X1_HVT U381 ( .A1(n327), .A2(n375), .S0(n319), .Y(n456) );
  MUX21X1_HVT U382 ( .A1(n448), .A2(n446), .S0(n237), .Y(n542) );
  MUX21X1_HVT U383 ( .A1(n327), .A2(n369), .S0(n380), .Y(n455) );
  NBUFFX2_HVT U384 ( .A(in[2]), .Y(n384) );
  NBUFFX2_HVT U385 ( .A(in[2]), .Y(n383) );
  XOR2X1_HVT U386 ( .A1(n366), .A2(n378), .Y(n610) );
  MUX21X1_HVT U387 ( .A1(n358), .A2(n373), .S0(n309), .Y(n553) );
  NBUFFX2_HVT U388 ( .A(n333), .Y(n358) );
  NBUFFX2_HVT U389 ( .A(n333), .Y(n359) );
  MUX21X1_HVT U390 ( .A1(n276), .A2(n360), .S0(n379), .Y(n452) );
  MUX21X1_HVT U391 ( .A1(n445), .A2(n449), .S0(n378), .Y(n622) );
  MUX21X1_HVT U392 ( .A1(n449), .A2(n357), .S0(n310), .Y(n616) );
  NBUFFX2_HVT U393 ( .A(n639), .Y(n366) );
  MUX21X1_HVT U394 ( .A1(n358), .A2(n249), .S0(n380), .Y(n615) );
  MUX21X1_HVT U395 ( .A1(n249), .A2(n446), .S0(n310), .Y(n621) );
  NBUFFX2_HVT U396 ( .A(n639), .Y(n367) );
  INVX1_HVT U397 ( .A(n459), .Y(n434) );
  NBUFFX2_HVT U398 ( .A(n655), .Y(n373) );
  NAND2X0_HVT U399 ( .A1(n355), .A2(n358), .Y(n655) );
  MUX21X1_HVT U400 ( .A1(n374), .A2(n373), .S0(n378), .Y(n641) );
  XOR2X1_HVT U401 ( .A1(n374), .A2(n376), .Y(n618) );
  MUX21X1_HVT U402 ( .A1(n343), .A2(n366), .S0(n309), .Y(n457) );
  MUX21X1_HVT U403 ( .A1(n343), .A2(n327), .S0(n378), .Y(n450) );
  MUX21X1_HVT U404 ( .A1(n343), .A2(n360), .S0(n377), .Y(n487) );
  MUX21X1_HVT U405 ( .A1(n355), .A2(n449), .S0(n310), .Y(n459) );
  MUX21X1_HVT U406 ( .A1(n445), .A2(n263), .S0(n310), .Y(n524) );
  XOR2X1_HVT U407 ( .A1(n319), .A2(n263), .Y(n607) );
  MUX21X1_HVT U408 ( .A1(n334), .A2(n343), .S0(n378), .Y(n631) );
  MUX21X1_HVT U409 ( .A1(n371), .A2(n263), .S0(n378), .Y(n458) );
  MUX21X1_HVT U410 ( .A1(n263), .A2(n372), .S0(n377), .Y(n462) );
  MUX21X1_HVT U411 ( .A1(n355), .A2(n263), .S0(n237), .Y(n453) );
  MUX21X1_HVT U412 ( .A1(n334), .A2(n374), .S0(n379), .Y(n638) );
  MUX21X1_HVT U413 ( .A1(n369), .A2(n334), .S0(n379), .Y(n626) );
  NBUFFX2_HVT U414 ( .A(n656), .Y(n375) );
  NBUFFX2_HVT U415 ( .A(n656), .Y(n374) );
  INVX0_HVT U416 ( .A(n644), .Y(n391) );
  INVX0_HVT U417 ( .A(n623), .Y(n392) );
  INVX0_HVT U418 ( .A(n617), .Y(n393) );
  INVX0_HVT U419 ( .A(n558), .Y(n394) );
  INVX0_HVT U420 ( .A(n519), .Y(n395) );
  INVX0_HVT U421 ( .A(n652), .Y(n398) );
  INVX0_HVT U422 ( .A(n649), .Y(n399) );
  INVX0_HVT U423 ( .A(n648), .Y(n400) );
  INVX0_HVT U424 ( .A(n620), .Y(n401) );
  INVX0_HVT U425 ( .A(n642), .Y(n402) );
  INVX0_HVT U426 ( .A(n647), .Y(n403) );
  INVX0_HVT U427 ( .A(n643), .Y(n404) );
  INVX0_HVT U428 ( .A(n641), .Y(n405) );
  INVX0_HVT U429 ( .A(n640), .Y(n406) );
  INVX0_HVT U430 ( .A(n637), .Y(n408) );
  INVX0_HVT U431 ( .A(n636), .Y(n409) );
  INVX0_HVT U432 ( .A(n635), .Y(n410) );
  INVX0_HVT U433 ( .A(n631), .Y(n413) );
  INVX0_HVT U434 ( .A(n629), .Y(n415) );
  INVX0_HVT U435 ( .A(n627), .Y(n417) );
  INVX0_HVT U436 ( .A(n625), .Y(n419) );
  INVX0_HVT U437 ( .A(n624), .Y(n420) );
  INVX0_HVT U438 ( .A(n622), .Y(n421) );
  INVX0_HVT U439 ( .A(n621), .Y(n422) );
  INVX0_HVT U440 ( .A(n618), .Y(n424) );
  INVX0_HVT U441 ( .A(n616), .Y(n425) );
  INVX0_HVT U442 ( .A(n615), .Y(n426) );
  INVX0_HVT U443 ( .A(n612), .Y(n427) );
  INVX0_HVT U444 ( .A(n611), .Y(n428) );
  INVX0_HVT U445 ( .A(n610), .Y(n429) );
  INVX0_HVT U446 ( .A(n646), .Y(n430) );
  INVX0_HVT U447 ( .A(n462), .Y(n431) );
  INVX0_HVT U448 ( .A(n458), .Y(n435) );
  INVX0_HVT U449 ( .A(n457), .Y(n436) );
  INVX0_HVT U450 ( .A(n456), .Y(n437) );
  INVX0_HVT U451 ( .A(n455), .Y(n438) );
  INVX0_HVT U452 ( .A(n454), .Y(n439) );
  INVX0_HVT U453 ( .A(n453), .Y(n440) );
  INVX0_HVT U454 ( .A(n501), .Y(n441) );
  INVX0_HVT U455 ( .A(n452), .Y(n442) );
  INVX0_HVT U456 ( .A(n451), .Y(n443) );
  INVX0_HVT U457 ( .A(n450), .Y(n444) );
endmodule

