
module keygen_0 ( round_num, keyin, keyout );
  input [0:3] round_num;
  input [0:127] keyin;
  output [0:127] keyout;
  wire   n1660, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n215, n216,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n520, n521, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n825, n826,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1128,
         n1129, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1334, n1335,
         n1336, n1337, n23, n49, n115, n130, n211, n212, n213, n214, n217,
         n218, n219, n220, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n328, n354, n398, n472, n516, n517, n518, n519, n522, n523, n524,
         n525, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n595, n596, n597, n598, n599, n600, n601, n603, n604,
         n605, n606, n607, n608, n609, n610, n633, n659, n822, n823, n824,
         n827, n828, n829, n830, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n938, n1083, n1125, n1126, n1127, n1130, n1131, n1132, n1133,
         n1134, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1277, n1333, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1389, n1390, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659;
  wire   [0:31] dummy;

  NAND2X0_HVT U4 ( .A1(n1355), .A2(n1233), .Y(n4) );
  NAND2X0_HVT U5 ( .A1(n1192), .A2(n1352), .Y(n5) );
  NAND2X0_HVT U6 ( .A1(n1231), .A2(n4), .Y(n6) );
  NAND2X0_HVT U15 ( .A1(n16), .A2(n1238), .Y(n15) );
  NAND2X0_HVT U17 ( .A1(n4), .A2(n1175), .Y(n18) );
  NAND2X0_HVT U21 ( .A1(n1230), .A2(n1357), .Y(n22) );
  NAND2X0_HVT U25 ( .A1(n1191), .A2(n1357), .Y(n26) );
  NAND2X0_HVT U33 ( .A1(n1357), .A2(n1589), .Y(n34) );
  NAND2X0_HVT U34 ( .A1(n1585), .A2(n1357), .Y(n35) );
  NAND2X0_HVT U39 ( .A1(n252), .A2(n1177), .Y(n40) );
  MUX41X1_HVT U50 ( .A1(n1571), .A3(n1528), .A2(n14), .A4(n1548), .S0(n854), 
        .S1(n1147), .Y(n51) );
  NAND2X0_HVT U52 ( .A1(n54), .A2(n43), .Y(n53) );
  MUX41X1_HVT U55 ( .A1(n871), .A3(n1547), .A2(n1546), .A4(n1174), .S0(n854), 
        .S1(n1148), .Y(n57) );
  NAND2X0_HVT U56 ( .A1(n1357), .A2(n1234), .Y(n58) );
  MUX41X1_HVT U57 ( .A1(n58), .A3(n1536), .A2(n1566), .A4(n1545), .S0(n854), 
        .S1(n1147), .Y(n59) );
  NAND2X0_HVT U59 ( .A1(n1231), .A2(n62), .Y(n61) );
  MUX41X1_HVT U60 ( .A1(n1572), .A3(n1544), .A2(n61), .A4(n11), .S0(n1363), 
        .S1(n1150), .Y(n63) );
  NAND2X0_HVT U61 ( .A1(n1238), .A2(n4), .Y(n64) );
  MUX41X1_HVT U62 ( .A1(n903), .A3(n64), .A2(n899), .A4(n1543), .S0(n1362), 
        .S1(n1147), .Y(n65) );
  AO21X1_HVT U65 ( .A1(n1541), .A2(n1152), .A3(n1565), .Y(n68) );
  MUX41X1_HVT U67 ( .A1(n1539), .A3(n68), .A2(n69), .A4(n67), .S0(n1359), .S1(
        n855), .Y(n70) );
  MUX41X1_HVT U69 ( .A1(n44), .A3(n1587), .A2(n26), .A4(n1573), .S0(n1149), 
        .S1(n254), .Y(n71) );
  NAND2X0_HVT U71 ( .A1(n1236), .A2(n74), .Y(n73) );
  AND3X1_HVT U75 ( .A1(n1234), .A2(n62), .A3(n79), .Y(n78) );
  MUX41X1_HVT U77 ( .A1(n46), .A3(n1529), .A2(n21), .A4(n1235), .S0(n1363), 
        .S1(n1147), .Y(n81) );
  MUX41X1_HVT U78 ( .A1(n81), .A3(n80), .A2(n76), .A4(n71), .S0(n272), .S1(
        n1195), .Y(n82) );
  MUX41X1_HVT U80 ( .A1(n83), .A3(n1574), .A2(n1575), .A4(n1550), .S0(n1150), 
        .S1(n855), .Y(n84) );
  MUX41X1_HVT U81 ( .A1(n10), .A3(n1567), .A2(n1576), .A4(n1588), .S0(n1150), 
        .S1(n254), .Y(n85) );
  AND2X1_HVT U82 ( .A1(n1355), .A2(n1194), .Y(n86) );
  NAND2X0_HVT U83 ( .A1(n1357), .A2(n1587), .Y(n87) );
  MUX41X1_HVT U84 ( .A1(n87), .A3(n247), .A2(n879), .A4(n86), .S0(n1150), .S1(
        n1361), .Y(n88) );
  MUX41X1_HVT U85 ( .A1(n1574), .A3(n1549), .A2(n890), .A4(n19), .S0(n1149), 
        .S1(n1363), .Y(n89) );
  MUX41X1_HVT U86 ( .A1(n89), .A3(n85), .A2(n88), .A4(n84), .S0(n1197), .S1(
        n271), .Y(n90) );
  AO21X1_HVT U93 ( .A1(n1155), .A2(n97), .A3(n1570), .Y(n96) );
  MUX41X1_HVT U94 ( .A1(n96), .A3(n94), .A2(n95), .A4(n92), .S0(n271), .S1(
        n1146), .Y(n98) );
  NAND2X0_HVT U97 ( .A1(n102), .A2(n103), .Y(n101) );
  MUX41X1_HVT U98 ( .A1(n101), .A3(n1555), .A2(n100), .A4(n99), .S0(n1359), 
        .S1(n1146), .Y(n104) );
  MUX41X1_HVT U102 ( .A1(n1567), .A3(n1529), .A2(n1355), .A4(n1573), .S0(n1149), .S1(n1361), .Y(n108) );
  MUX41X1_HVT U104 ( .A1(n48), .A3(n1569), .A2(n1540), .A4(n34), .S0(n1362), 
        .S1(n1148), .Y(n110) );
  MUX41X1_HVT U106 ( .A1(n1551), .A3(n4), .A2(n111), .A4(n1552), .S0(n1150), 
        .S1(n1363), .Y(n112) );
  NAND2X0_HVT U111 ( .A1(n1233), .A2(n117), .Y(n116) );
  NAND2X0_HVT U118 ( .A1(n125), .A2(n126), .Y(n124) );
  MUX41X1_HVT U120 ( .A1(n22), .A3(n903), .A2(n1539), .A4(n1578), .S0(n1359), 
        .S1(n1361), .Y(n128) );
  AO21X1_HVT U125 ( .A1(n1358), .A2(n1236), .A3(n247), .Y(n133) );
  AND3X1_HVT U129 ( .A1(n272), .A2(n1357), .A3(n1194), .Y(n137) );
  MUX41X1_HVT U132 ( .A1(n139), .A3(n137), .A2(n138), .A4(n136), .S0(n1149), 
        .S1(n1361), .Y(n140) );
  MUX41X1_HVT U133 ( .A1(n140), .A3(n135), .A2(n129), .A4(n121), .S0(n1196), 
        .S1(keyin[111]), .Y(dummy[4]) );
  MUX41X1_HVT U134 ( .A1(n1583), .A3(n27), .A2(n1578), .A4(n1235), .S0(n1362), 
        .S1(n1148), .Y(n141) );
  MUX41X1_HVT U137 ( .A1(n1174), .A3(n1561), .A2(n1235), .A4(n1556), .S0(n1149), .S1(n1362), .Y(n144) );
  AND2X1_HVT U138 ( .A1(n1237), .A2(n1356), .Y(n145) );
  MUX41X1_HVT U139 ( .A1(n1549), .A3(n1568), .A2(n25), .A4(n145), .S0(n1361), 
        .S1(n1146), .Y(n146) );
  MUX41X1_HVT U140 ( .A1(n146), .A3(n144), .A2(n143), .A4(n141), .S0(n272), 
        .S1(n1195), .Y(n147) );
  MUX41X1_HVT U143 ( .A1(n24), .A3(n879), .A2(n1560), .A4(n1580), .S0(n1150), 
        .S1(n855), .Y(n150) );
  NAND2X0_HVT U144 ( .A1(n1352), .A2(n1238), .Y(n74) );
  OA21X1_HVT U146 ( .A1(n1533), .A2(n1364), .A3(n30), .Y(n152) );
  MUX41X1_HVT U148 ( .A1(n1580), .A3(n1567), .A2(n29), .A4(n1535), .S0(n1363), 
        .S1(n1148), .Y(n154) );
  MUX41X1_HVT U149 ( .A1(n154), .A3(n150), .A2(n153), .A4(n149), .S0(n1197), 
        .S1(n272), .Y(n155) );
  MUX41X1_HVT U151 ( .A1(n871), .A3(n1530), .A2(n1575), .A4(n1583), .S0(n1363), 
        .S1(n1148), .Y(n156) );
  OA21X1_HVT U153 ( .A1(n41), .A2(n1364), .A3(n159), .Y(n158) );
  AND2X1_HVT U156 ( .A1(n247), .A2(n74), .Y(n162) );
  MUX41X1_HVT U158 ( .A1(n47), .A3(n162), .A2(n163), .A4(n161), .S0(n1153), 
        .S1(n1361), .Y(n164) );
  MUX41X1_HVT U159 ( .A1(n22), .A3(n1547), .A2(n1554), .A4(n893), .S0(n1149), 
        .S1(n1363), .Y(n165) );
  MUX41X1_HVT U160 ( .A1(n165), .A3(n164), .A2(n160), .A4(n156), .S0(n271), 
        .S1(n1195), .Y(n166) );
  AND2X1_HVT U161 ( .A1(n1155), .A2(n1192), .Y(n167) );
  NAND2X0_HVT U165 ( .A1(n1353), .A2(n1587), .Y(n171) );
  MUX41X1_HVT U166 ( .A1(n15), .A3(n39), .A2(n171), .A4(n1576), .S0(n1150), 
        .S1(n1362), .Y(n172) );
  NAND2X0_HVT U167 ( .A1(n1238), .A2(n62), .Y(n173) );
  OA21X1_HVT U169 ( .A1(n899), .A2(n1364), .A3(n30), .Y(n175) );
  NAND2X0_HVT U171 ( .A1(n1588), .A2(n1357), .Y(n177) );
  MUX41X1_HVT U172 ( .A1(n1235), .A3(n1573), .A2(n1572), .A4(n177), .S0(n1362), 
        .S1(n1148), .Y(n178) );
  NAND2X0_HVT U175 ( .A1(n1352), .A2(n8), .Y(n16) );
  NAND2X0_HVT U176 ( .A1(n253), .A2(n1589), .Y(n180) );
  MUX41X1_HVT U177 ( .A1(n180), .A3(n39), .A2(n1577), .A4(n16), .S0(n854), 
        .S1(n1146), .Y(n181) );
  MUX41X1_HVT U179 ( .A1(n20), .A3(n1589), .A2(n1581), .A4(n182), .S0(n1151), 
        .S1(n1362), .Y(n183) );
  MUX41X1_HVT U180 ( .A1(n87), .A3(n1192), .A2(n1564), .A4(n1532), .S0(n855), 
        .S1(n1146), .Y(n184) );
  MUX41X1_HVT U184 ( .A1(n187), .A3(n183), .A2(n184), .A4(n181), .S0(n1197), 
        .S1(n272), .Y(n188) );
  MUX41X1_HVT U185 ( .A1(n15), .A3(n1582), .A2(n874), .A4(n1581), .S0(n1151), 
        .S1(n1361), .Y(n189) );
  MUX41X1_HVT U186 ( .A1(n1537), .A3(n28), .A2(n10), .A4(n1534), .S0(n1151), 
        .S1(n855), .Y(n190) );
  MUX41X1_HVT U188 ( .A1(n191), .A3(n38), .A2(n1569), .A4(n47), .S0(n1149), 
        .S1(n855), .Y(n192) );
  MUX41X1_HVT U190 ( .A1(n193), .A3(n883), .A2(n16), .A4(n74), .S0(n1151), 
        .S1(n1363), .Y(n194) );
  MUX41X1_HVT U194 ( .A1(n1579), .A3(n34), .A2(n1235), .A4(n196), .S0(n1151), 
        .S1(n1362), .Y(n197) );
  MUX41X1_HVT U195 ( .A1(n42), .A3(n5), .A2(n27), .A4(n50), .S0(n1151), .S1(
        n1363), .Y(n198) );
  MUX41X1_HVT U196 ( .A1(n1563), .A3(n32), .A2(n19), .A4(n874), .S0(n1362), 
        .S1(n1150), .Y(n199) );
  OA21X1_HVT U198 ( .A1(n9), .A2(n1364), .A3(n1561), .Y(n201) );
  MUX41X1_HVT U200 ( .A1(n202), .A3(n198), .A2(n199), .A4(n197), .S0(n1197), 
        .S1(n1359), .Y(n203) );
  AO21X1_HVT U202 ( .A1(n890), .A2(n1154), .A3(n1570), .Y(n205) );
  MUX41X1_HVT U204 ( .A1(n1538), .A3(n247), .A2(n1581), .A4(n1), .S0(n1151), 
        .S1(n854), .Y(n207) );
  MUX41X1_HVT U205 ( .A1(n4), .A3(n15), .A2(n1553), .A4(n24), .S0(n1151), .S1(
        n854), .Y(n208) );
  MUX41X1_HVT U206 ( .A1(n1194), .A3(n61), .A2(n1582), .A4(n1557), .S0(n1151), 
        .S1(n1361), .Y(n209) );
  MUX41X1_HVT U207 ( .A1(n209), .A3(n207), .A2(n208), .A4(n206), .S0(n1196), 
        .S1(n272), .Y(n210) );
  NAND2X0_HVT U211 ( .A1(n1237), .A2(n1355), .Y(n62) );
  NAND2X0_HVT U212 ( .A1(n1353), .A2(n1230), .Y(n117) );
  NAND2X0_HVT U215 ( .A1(n247), .A2(n1357), .Y(n215) );
  NAND2X0_HVT U216 ( .A1(n1236), .A2(n117), .Y(n216) );
  AO21X1_HVT U218 ( .A1(n1357), .A2(n1583), .A3(n1364), .Y(n102) );
  NAND2X0_HVT U219 ( .A1(n253), .A2(n1583), .Y(n159) );
  NAND2X0_HVT U221 ( .A1(n1155), .A2(n215), .Y(n79) );
  NAND2X0_HVT U317 ( .A1(n1339), .A2(n1224), .Y(n309) );
  NAND2X0_HVT U318 ( .A1(n824), .A2(n1339), .Y(n310) );
  NAND2X0_HVT U319 ( .A1(n1222), .A2(n309), .Y(n311) );
  XOR2X2_HVT U320 ( .A1(n1172), .A2(n1187), .Y(n313) );
  NAND2X0_HVT U328 ( .A1(n321), .A2(n1229), .Y(n320) );
  NAND2X0_HVT U330 ( .A1(n309), .A2(n1171), .Y(n323) );
  NAND2X0_HVT U334 ( .A1(n1221), .A2(n1341), .Y(n327) );
  NAND2X0_HVT U338 ( .A1(n1186), .A2(n287), .Y(n331) );
  NAND2X0_HVT U346 ( .A1(n1341), .A2(n1526), .Y(n339) );
  NAND2X0_HVT U347 ( .A1(n1522), .A2(n287), .Y(n340) );
  NAND2X0_HVT U352 ( .A1(n1339), .A2(n1173), .Y(n345) );
  MUX41X1_HVT U363 ( .A1(n1508), .A3(n1466), .A2(n319), .A4(n1486), .S0(n1348), 
        .S1(n1345), .Y(n356) );
  NAND2X0_HVT U365 ( .A1(n359), .A2(n348), .Y(n358) );
  MUX41X1_HVT U368 ( .A1(n875), .A3(n1485), .A2(n1484), .A4(n1170), .S0(n1347), 
        .S1(n938), .Y(n362) );
  NAND2X0_HVT U369 ( .A1(n286), .A2(n1225), .Y(n363) );
  MUX41X1_HVT U370 ( .A1(n363), .A3(n1474), .A2(n1503), .A4(n1483), .S0(n259), 
        .S1(n1125), .Y(n364) );
  NAND2X0_HVT U372 ( .A1(n1222), .A2(n367), .Y(n366) );
  MUX41X1_HVT U373 ( .A1(n1509), .A3(n1482), .A2(n366), .A4(n316), .S0(n259), 
        .S1(n1345), .Y(n368) );
  NAND2X0_HVT U374 ( .A1(n1229), .A2(n309), .Y(n369) );
  MUX41X1_HVT U375 ( .A1(n904), .A3(n369), .A2(n901), .A4(n1481), .S0(n1347), 
        .S1(n1345), .Y(n370) );
  AO21X1_HVT U378 ( .A1(n1479), .A2(n1130), .A3(n1502), .Y(n373) );
  MUX41X1_HVT U380 ( .A1(n1477), .A3(n373), .A2(n374), .A4(n372), .S0(n1343), 
        .S1(n265), .Y(n375) );
  MUX41X1_HVT U382 ( .A1(n349), .A3(n1524), .A2(n331), .A4(n1510), .S0(n1125), 
        .S1(n1347), .Y(n376) );
  NAND2X0_HVT U384 ( .A1(n1227), .A2(n379), .Y(n378) );
  AND3X1_HVT U388 ( .A1(n1225), .A2(n367), .A3(n384), .Y(n383) );
  MUX41X1_HVT U390 ( .A1(n351), .A3(n1467), .A2(n326), .A4(n1226), .S0(n258), 
        .S1(n1126), .Y(n386) );
  MUX41X1_HVT U391 ( .A1(n386), .A3(n385), .A2(n381), .A4(n376), .S0(n1343), 
        .S1(n1189), .Y(n387) );
  MUX41X1_HVT U393 ( .A1(n388), .A3(n1511), .A2(n1512), .A4(n1488), .S0(n1126), 
        .S1(n1347), .Y(n389) );
  MUX41X1_HVT U394 ( .A1(n315), .A3(n1504), .A2(n1513), .A4(n1525), .S0(n1126), 
        .S1(n259), .Y(n390) );
  AND2X1_HVT U395 ( .A1(n1339), .A2(n1188), .Y(n391) );
  NAND2X0_HVT U396 ( .A1(n286), .A2(n1524), .Y(n392) );
  MUX41X1_HVT U397 ( .A1(n392), .A3(n313), .A2(n877), .A4(n391), .S0(n1126), 
        .S1(n1348), .Y(n393) );
  MUX41X1_HVT U398 ( .A1(n1511), .A3(n1487), .A2(n886), .A4(n324), .S0(n1125), 
        .S1(n1347), .Y(n394) );
  MUX41X1_HVT U399 ( .A1(n394), .A3(n390), .A2(n393), .A4(n389), .S0(n1190), 
        .S1(n1342), .Y(n395) );
  AO21X1_HVT U406 ( .A1(n1133), .A2(n402), .A3(n1507), .Y(n401) );
  NAND2X0_HVT U410 ( .A1(n407), .A2(n408), .Y(n406) );
  MUX41X1_HVT U415 ( .A1(n1504), .A3(n1467), .A2(n1339), .A4(n1510), .S0(n1125), .S1(n258), .Y(n413) );
  MUX41X1_HVT U417 ( .A1(n353), .A3(n1506), .A2(n1478), .A4(n339), .S0(n265), 
        .S1(n1083), .Y(n415) );
  MUX41X1_HVT U419 ( .A1(n1489), .A3(n309), .A2(n416), .A4(n1490), .S0(n1126), 
        .S1(n259), .Y(n417) );
  OA21X1_HVT U423 ( .A1(n1497), .A2(n1344), .A3(n1481), .Y(n420) );
  NAND2X0_HVT U424 ( .A1(n1224), .A2(n422), .Y(n421) );
  NAND2X0_HVT U431 ( .A1(n430), .A2(n431), .Y(n429) );
  MUX41X1_HVT U433 ( .A1(n327), .A3(n904), .A2(n1477), .A4(n1515), .S0(n1343), 
        .S1(n1349), .Y(n433) );
  AND2X1_HVT U435 ( .A1(n1339), .A2(n1170), .Y(n435) );
  MUX41X1_HVT U436 ( .A1(n320), .A3(n435), .A2(n1488), .A4(n335), .S0(n1343), 
        .S1(n1348), .Y(n436) );
  MUX41X1_HVT U445 ( .A1(n444), .A3(n442), .A2(n443), .A4(n441), .S0(n1125), 
        .S1(n1350), .Y(n445) );
  MUX41X1_HVT U447 ( .A1(n1520), .A3(n332), .A2(n1515), .A4(n1226), .S0(n258), 
        .S1(n1083), .Y(n446) );
  MUX41X1_HVT U450 ( .A1(n1170), .A3(n269), .A2(n1226), .A4(n1494), .S0(n1125), 
        .S1(n258), .Y(n449) );
  AND2X1_HVT U451 ( .A1(n1227), .A2(n286), .Y(n450) );
  MUX41X1_HVT U452 ( .A1(n1487), .A3(n1505), .A2(n330), .A4(n450), .S0(n259), 
        .S1(n938), .Y(n451) );
  MUX41X1_HVT U453 ( .A1(n451), .A3(n449), .A2(n448), .A4(n446), .S0(n1343), 
        .S1(n1189), .Y(n452) );
  MUX41X1_HVT U456 ( .A1(n329), .A3(n877), .A2(n1498), .A4(n1517), .S0(n1126), 
        .S1(n258), .Y(n455) );
  NAND2X0_HVT U457 ( .A1(n1339), .A2(n1229), .Y(n379) );
  MUX41X1_HVT U461 ( .A1(n1517), .A3(n1504), .A2(n334), .A4(n1473), .S0(n258), 
        .S1(n1083), .Y(n459) );
  MUX41X1_HVT U462 ( .A1(n459), .A3(n455), .A2(n458), .A4(n454), .S0(
        keyin[113]), .S1(n1343), .Y(n460) );
  MUX41X1_HVT U464 ( .A1(n875), .A3(n1468), .A2(n1512), .A4(n1520), .S0(n259), 
        .S1(n1083), .Y(n461) );
  AND2X1_HVT U469 ( .A1(n313), .A2(n379), .Y(n467) );
  MUX41X1_HVT U471 ( .A1(n352), .A3(n467), .A2(n468), .A4(n466), .S0(n1131), 
        .S1(n1347), .Y(n469) );
  MUX41X1_HVT U472 ( .A1(n327), .A3(n1485), .A2(n1492), .A4(n891), .S0(n1125), 
        .S1(n1348), .Y(n470) );
  MUX41X1_HVT U473 ( .A1(n470), .A3(n469), .A2(n465), .A4(n461), .S0(n1343), 
        .S1(n1189), .Y(n471) );
  NAND2X0_HVT U478 ( .A1(n1339), .A2(n1524), .Y(n476) );
  MUX41X1_HVT U479 ( .A1(n320), .A3(n344), .A2(n476), .A4(n1513), .S0(n1126), 
        .S1(n1350), .Y(n477) );
  NAND2X0_HVT U480 ( .A1(n1229), .A2(n367), .Y(n478) );
  NAND2X0_HVT U484 ( .A1(n1525), .A2(n1341), .Y(n482) );
  MUX41X1_HVT U485 ( .A1(n1226), .A3(n1510), .A2(n1509), .A4(n482), .S0(n259), 
        .S1(n1083), .Y(n483) );
  NAND2X0_HVT U488 ( .A1(n1339), .A2(n313), .Y(n321) );
  NAND2X0_HVT U489 ( .A1(n1339), .A2(n1526), .Y(n485) );
  MUX41X1_HVT U490 ( .A1(n485), .A3(n344), .A2(n1514), .A4(n321), .S0(n259), 
        .S1(n938), .Y(n486) );
  MUX41X1_HVT U492 ( .A1(n325), .A3(n1526), .A2(n1518), .A4(n487), .S0(n1127), 
        .S1(n258), .Y(n488) );
  MUX41X1_HVT U493 ( .A1(n392), .A3(n1186), .A2(n1501), .A4(n1470), .S0(n258), 
        .S1(n938), .Y(n489) );
  MUX41X1_HVT U498 ( .A1(n320), .A3(n1519), .A2(n872), .A4(n1518), .S0(n1127), 
        .S1(n259), .Y(n494) );
  MUX41X1_HVT U499 ( .A1(n1475), .A3(n333), .A2(n315), .A4(n1472), .S0(n1127), 
        .S1(n1348), .Y(n495) );
  MUX41X1_HVT U501 ( .A1(n496), .A3(n343), .A2(n1506), .A4(n352), .S0(n1125), 
        .S1(n1348), .Y(n497) );
  MUX41X1_HVT U503 ( .A1(n498), .A3(n884), .A2(n321), .A4(n379), .S0(n1127), 
        .S1(n258), .Y(n499) );
  MUX41X1_HVT U504 ( .A1(n499), .A3(n495), .A2(n497), .A4(n494), .S0(n1190), 
        .S1(n1342), .Y(n500) );
  MUX41X1_HVT U508 ( .A1(n347), .A3(n310), .A2(n332), .A4(n355), .S0(n1127), 
        .S1(n1348), .Y(n503) );
  MUX41X1_HVT U509 ( .A1(n1500), .A3(n337), .A2(n324), .A4(n872), .S0(n265), 
        .S1(n1126), .Y(n504) );
  AO21X1_HVT U515 ( .A1(n886), .A2(n266), .A3(n1507), .Y(n510) );
  MUX41X1_HVT U517 ( .A1(n1476), .A3(n313), .A2(n1518), .A4(n1228), .S0(n1127), 
        .S1(n1134), .Y(n512) );
  MUX41X1_HVT U518 ( .A1(n309), .A3(n320), .A2(n1491), .A4(n329), .S0(n1127), 
        .S1(n259), .Y(n513) );
  MUX41X1_HVT U519 ( .A1(n1188), .A3(n366), .A2(n1519), .A4(n1495), .S0(n1127), 
        .S1(n1348), .Y(n514) );
  NAND2X0_HVT U524 ( .A1(n1227), .A2(n1339), .Y(n367) );
  NAND2X0_HVT U525 ( .A1(n1339), .A2(n1221), .Y(n422) );
  NAND2X0_HVT U528 ( .A1(n313), .A2(n1341), .Y(n520) );
  NAND2X0_HVT U529 ( .A1(n1227), .A2(n422), .Y(n521) );
  NAND2X0_HVT U532 ( .A1(n1339), .A2(n1520), .Y(n464) );
  NAND2X0_HVT U534 ( .A1(n1350), .A2(n520), .Y(n384) );
  NAND2X0_HVT U631 ( .A1(n1183), .A2(n1243), .Y(n615) );
  NAND2X0_HVT U632 ( .A1(n1214), .A2(n614), .Y(n616) );
  XOR2X2_HVT U633 ( .A1(n1456), .A2(n1184), .Y(n618) );
  NAND2X0_HVT U641 ( .A1(n626), .A2(n1220), .Y(n625) );
  NAND2X0_HVT U643 ( .A1(n614), .A2(n1168), .Y(n628) );
  NAND2X0_HVT U647 ( .A1(n617), .A2(n1245), .Y(n632) );
  NAND2X0_HVT U651 ( .A1(n1182), .A2(n1245), .Y(n636) );
  NAND2X0_HVT U659 ( .A1(n1245), .A2(n1459), .Y(n644) );
  NAND2X0_HVT U660 ( .A1(n1455), .A2(n1245), .Y(n645) );
  NAND2X0_HVT U665 ( .A1(n1242), .A2(n1169), .Y(n650) );
  MUX41X1_HVT U676 ( .A1(n1441), .A3(n1398), .A2(n624), .A4(n1418), .S0(n608), 
        .S1(n1248), .Y(n661) );
  NAND2X0_HVT U678 ( .A1(n664), .A2(n653), .Y(n663) );
  MUX41X1_HVT U681 ( .A1(n876), .A3(n1417), .A2(n1416), .A4(n1167), .S0(n264), 
        .S1(n1248), .Y(n667) );
  NAND2X0_HVT U682 ( .A1(n1245), .A2(n1217), .Y(n668) );
  MUX41X1_HVT U683 ( .A1(n668), .A3(n1406), .A2(n1436), .A4(n1415), .S0(n913), 
        .S1(n908), .Y(n669) );
  NAND2X0_HVT U685 ( .A1(n1214), .A2(n672), .Y(n671) );
  MUX41X1_HVT U686 ( .A1(n1442), .A3(n1414), .A2(n671), .A4(n621), .S0(n1251), 
        .S1(n1248), .Y(n673) );
  NAND2X0_HVT U687 ( .A1(n1220), .A2(n614), .Y(n674) );
  MUX41X1_HVT U688 ( .A1(n905), .A3(n674), .A2(n902), .A4(n1413), .S0(n1252), 
        .S1(n909), .Y(n675) );
  AO21X1_HVT U691 ( .A1(n1411), .A2(n911), .A3(n1435), .Y(n678) );
  MUX41X1_HVT U693 ( .A1(n1409), .A3(n678), .A2(n679), .A4(n677), .S0(n288), 
        .S1(n608), .Y(n680) );
  MUX41X1_HVT U694 ( .A1(n680), .A3(n676), .A2(n670), .A4(n666), .S0(
        keyin[121]), .S1(keyin[127]), .Y(dummy[23]) );
  MUX41X1_HVT U695 ( .A1(n654), .A3(n1457), .A2(n636), .A4(n1443), .S0(n908), 
        .S1(n1251), .Y(n681) );
  NAND2X0_HVT U697 ( .A1(n1218), .A2(n684), .Y(n683) );
  AND3X1_HVT U701 ( .A1(n1217), .A2(n672), .A3(n689), .Y(n688) );
  MUX41X1_HVT U703 ( .A1(n656), .A3(n1399), .A2(n631), .A4(n1218), .S0(n264), 
        .S1(n910), .Y(n691) );
  MUX41X1_HVT U704 ( .A1(n691), .A3(n690), .A2(n686), .A4(n681), .S0(n251), 
        .S1(keyin[121]), .Y(n692) );
  MUX41X1_HVT U706 ( .A1(n693), .A3(n1444), .A2(n1445), .A4(n1420), .S0(n909), 
        .S1(n1252), .Y(n694) );
  MUX41X1_HVT U707 ( .A1(n620), .A3(n1437), .A2(n1446), .A4(n1458), .S0(n909), 
        .S1(n608), .Y(n695) );
  AND2X1_HVT U708 ( .A1(n1243), .A2(n1185), .Y(n696) );
  NAND2X0_HVT U709 ( .A1(n1245), .A2(n1457), .Y(n697) );
  MUX41X1_HVT U710 ( .A1(n697), .A3(n618), .A2(n878), .A4(n696), .S0(n909), 
        .S1(n607), .Y(n698) );
  MUX41X1_HVT U711 ( .A1(n1444), .A3(n1419), .A2(n887), .A4(n629), .S0(n908), 
        .S1(n1252), .Y(n699) );
  MUX41X1_HVT U712 ( .A1(n699), .A3(n695), .A2(n698), .A4(n694), .S0(
        keyin[121]), .S1(n251), .Y(n700) );
  AO21X1_HVT U719 ( .A1(n914), .A2(n707), .A3(n1440), .Y(n706) );
  MUX41X1_HVT U720 ( .A1(n706), .A3(n704), .A2(n705), .A4(n702), .S0(n288), 
        .S1(n1248), .Y(n708) );
  NAND2X0_HVT U723 ( .A1(n712), .A2(n713), .Y(n711) );
  MUX41X1_HVT U724 ( .A1(n711), .A3(n1425), .A2(n710), .A4(n709), .S0(n288), 
        .S1(n1248), .Y(n714) );
  MUX41X1_HVT U728 ( .A1(n1437), .A3(n1399), .A2(n1239), .A4(n1443), .S0(n908), 
        .S1(n608), .Y(n718) );
  MUX41X1_HVT U730 ( .A1(n658), .A3(n1439), .A2(n1410), .A4(n644), .S0(n1252), 
        .S1(n907), .Y(n720) );
  MUX41X1_HVT U732 ( .A1(n1421), .A3(n614), .A2(n721), .A4(n1422), .S0(n909), 
        .S1(n607), .Y(n722) );
  NAND2X0_HVT U737 ( .A1(n1216), .A2(n727), .Y(n726) );
  MUX41X1_HVT U741 ( .A1(n730), .A3(n724), .A2(n728), .A4(n725), .S0(n909), 
        .S1(n607), .Y(n731) );
  NAND2X0_HVT U744 ( .A1(n735), .A2(n736), .Y(n734) );
  MUX41X1_HVT U746 ( .A1(n632), .A3(n905), .A2(n1409), .A4(n1448), .S0(n288), 
        .S1(n608), .Y(n738) );
  AND2X1_HVT U748 ( .A1(n1243), .A2(n1167), .Y(n740) );
  MUX41X1_HVT U749 ( .A1(n625), .A3(n740), .A2(n1420), .A4(n640), .S0(n1246), 
        .S1(n607), .Y(n741) );
  MUX41X1_HVT U760 ( .A1(n1453), .A3(n637), .A2(n1448), .A4(n1219), .S0(n915), 
        .S1(n907), .Y(n751) );
  MUX41X1_HVT U763 ( .A1(n1167), .A3(n1431), .A2(n1218), .A4(n1426), .S0(n908), 
        .S1(n1251), .Y(n754) );
  AND2X1_HVT U764 ( .A1(n1219), .A2(n1244), .Y(n755) );
  MUX41X1_HVT U765 ( .A1(n1419), .A3(n1438), .A2(n635), .A4(n755), .S0(n264), 
        .S1(n1248), .Y(n756) );
  MUX41X1_HVT U766 ( .A1(n756), .A3(n754), .A2(n753), .A4(n751), .S0(n251), 
        .S1(keyin[121]), .Y(n757) );
  MUX41X1_HVT U769 ( .A1(n634), .A3(n878), .A2(n1430), .A4(n1450), .S0(n909), 
        .S1(n1251), .Y(n760) );
  NAND2X0_HVT U770 ( .A1(n1240), .A2(n1220), .Y(n684) );
  OA21X1_HVT U772 ( .A1(n1403), .A2(n1254), .A3(n640), .Y(n762) );
  MUX41X1_HVT U774 ( .A1(n1450), .A3(n1437), .A2(n639), .A4(n1405), .S0(n264), 
        .S1(n907), .Y(n764) );
  MUX41X1_HVT U775 ( .A1(n764), .A3(n760), .A2(n763), .A4(n759), .S0(
        keyin[121]), .S1(n251), .Y(n765) );
  MUX41X1_HVT U777 ( .A1(n876), .A3(n1400), .A2(n1445), .A4(n1453), .S0(n264), 
        .S1(n907), .Y(n766) );
  OA21X1_HVT U779 ( .A1(n651), .A2(n1254), .A3(n769), .Y(n768) );
  AND2X1_HVT U782 ( .A1(n618), .A2(n684), .Y(n772) );
  MUX41X1_HVT U784 ( .A1(n657), .A3(n772), .A2(n773), .A4(n771), .S0(n912), 
        .S1(n1251), .Y(n774) );
  MUX41X1_HVT U785 ( .A1(n632), .A3(n1417), .A2(n1424), .A4(n892), .S0(n908), 
        .S1(n1252), .Y(n775) );
  MUX41X1_HVT U786 ( .A1(n775), .A3(n774), .A2(n770), .A4(n766), .S0(n251), 
        .S1(keyin[121]), .Y(n776) );
  AND2X1_HVT U787 ( .A1(n915), .A2(n1183), .Y(n777) );
  NAND2X0_HVT U791 ( .A1(n213), .A2(n1457), .Y(n781) );
  MUX41X1_HVT U792 ( .A1(n625), .A3(n649), .A2(n781), .A4(n1446), .S0(n909), 
        .S1(n607), .Y(n782) );
  NAND2X0_HVT U793 ( .A1(n1220), .A2(n672), .Y(n783) );
  OA21X1_HVT U795 ( .A1(n902), .A2(n1254), .A3(n640), .Y(n785) );
  NAND2X0_HVT U797 ( .A1(n1458), .A2(n1245), .Y(n787) );
  MUX41X1_HVT U798 ( .A1(n1219), .A3(n1443), .A2(n1442), .A4(n787), .S0(n264), 
        .S1(n907), .Y(n788) );
  MUX41X1_HVT U799 ( .A1(n788), .A3(n782), .A2(n786), .A4(n780), .S0(
        keyin[121]), .S1(n251), .Y(n789) );
  NAND2X0_HVT U801 ( .A1(n1240), .A2(n618), .Y(n626) );
  NAND2X0_HVT U802 ( .A1(n1242), .A2(n1459), .Y(n790) );
  MUX41X1_HVT U803 ( .A1(n790), .A3(n649), .A2(n1447), .A4(n626), .S0(n914), 
        .S1(n1248), .Y(n791) );
  MUX41X1_HVT U805 ( .A1(n630), .A3(n1459), .A2(n1451), .A4(n792), .S0(n910), 
        .S1(n1252), .Y(n793) );
  MUX41X1_HVT U806 ( .A1(n697), .A3(n1183), .A2(n1434), .A4(n1402), .S0(n264), 
        .S1(n1249), .Y(n794) );
  OA21X1_HVT U808 ( .A1(n643), .A2(n1254), .A3(n1419), .Y(n796) );
  MUX41X1_HVT U810 ( .A1(n797), .A3(n793), .A2(n794), .A4(n791), .S0(
        keyin[121]), .S1(n288), .Y(n798) );
  MUX41X1_HVT U811 ( .A1(n625), .A3(n1452), .A2(n873), .A4(n1451), .S0(n910), 
        .S1(n1253), .Y(n799) );
  MUX41X1_HVT U812 ( .A1(n1407), .A3(n638), .A2(n620), .A4(n1404), .S0(n910), 
        .S1(n1252), .Y(n800) );
  MUX41X1_HVT U814 ( .A1(n801), .A3(n648), .A2(n1439), .A4(n657), .S0(n908), 
        .S1(n608), .Y(n802) );
  MUX41X1_HVT U816 ( .A1(n803), .A3(n885), .A2(n626), .A4(n684), .S0(n910), 
        .S1(n1252), .Y(n804) );
  MUX41X1_HVT U817 ( .A1(n804), .A3(n800), .A2(n802), .A4(n799), .S0(
        keyin[121]), .S1(n288), .Y(n805) );
  MUX41X1_HVT U820 ( .A1(n1449), .A3(n644), .A2(n1219), .A4(n806), .S0(n910), 
        .S1(n1251), .Y(n807) );
  MUX41X1_HVT U821 ( .A1(n652), .A3(n615), .A2(n637), .A4(n660), .S0(n910), 
        .S1(n1251), .Y(n808) );
  MUX41X1_HVT U822 ( .A1(n1433), .A3(n642), .A2(n629), .A4(n873), .S0(n607), 
        .S1(n1248), .Y(n809) );
  OA21X1_HVT U824 ( .A1(n619), .A2(n1254), .A3(n1431), .Y(n811) );
  MUX41X1_HVT U826 ( .A1(n812), .A3(n808), .A2(n809), .A4(n807), .S0(
        keyin[121]), .S1(n288), .Y(n813) );
  AO21X1_HVT U828 ( .A1(n887), .A2(n913), .A3(n1440), .Y(n815) );
  MUX41X1_HVT U830 ( .A1(n1408), .A3(n618), .A2(n1451), .A4(n611), .S0(n910), 
        .S1(n607), .Y(n817) );
  MUX41X1_HVT U831 ( .A1(n614), .A3(n625), .A2(n1423), .A4(n634), .S0(n910), 
        .S1(n1251), .Y(n818) );
  MUX41X1_HVT U832 ( .A1(n1185), .A3(n671), .A2(n1452), .A4(n1427), .S0(n910), 
        .S1(n607), .Y(n819) );
  NAND2X0_HVT U837 ( .A1(n1219), .A2(n1241), .Y(n672) );
  NAND2X0_HVT U838 ( .A1(n212), .A2(n617), .Y(n727) );
  NAND2X0_HVT U841 ( .A1(n618), .A2(n1245), .Y(n825) );
  NAND2X0_HVT U842 ( .A1(n1218), .A2(n727), .Y(n826) );
  AO21X1_HVT U844 ( .A1(n1245), .A2(n1453), .A3(n1254), .Y(n712) );
  NAND2X0_HVT U845 ( .A1(n212), .A2(n1453), .Y(n769) );
  NAND2X0_HVT U847 ( .A1(n915), .A2(n825), .Y(n689) );
  NAND2X0_HVT U942 ( .A1(n1367), .A2(n1206), .Y(n918) );
  NAND2X0_HVT U943 ( .A1(n1371), .A2(n1180), .Y(n920) );
  NAND2X0_HVT U944 ( .A1(n1201), .A2(n1366), .Y(n921) );
  NAND2X0_HVT U945 ( .A1(n1209), .A2(n918), .Y(n922) );
  NAND2X0_HVT U952 ( .A1(n929), .A2(n1213), .Y(n928) );
  NAND2X0_HVT U954 ( .A1(n918), .A2(n1178), .Y(n931) );
  NAND2X0_HVT U960 ( .A1(n1208), .A2(n1371), .Y(n937) );
  NAND2X0_HVT U963 ( .A1(n1200), .A2(n1371), .Y(n940) );
  NAND2X0_HVT U971 ( .A1(n1654), .A2(n1371), .Y(n949) );
  NAND2X0_HVT U977 ( .A1(n1365), .A2(n828), .Y(n955) );
  MUX41X1_HVT U990 ( .A1(n1641), .A3(n1599), .A2(n935), .A4(n1617), .S0(n1378), 
        .S1(n1162), .Y(n967) );
  NAND2X0_HVT U992 ( .A1(n970), .A2(n958), .Y(n969) );
  NAND2X0_HVT U995 ( .A1(n1209), .A2(n974), .Y(n973) );
  MUX41X1_HVT U996 ( .A1(n1642), .A3(n1616), .A2(n973), .A4(n926), .S0(n1164), 
        .S1(n1162), .Y(n975) );
  NAND2X0_HVT U997 ( .A1(n1213), .A2(n918), .Y(n976) );
  MUX41X1_HVT U998 ( .A1(n906), .A3(n976), .A2(n900), .A4(n1615), .S0(n1164), 
        .S1(n1162), .Y(n977) );
  MUX41X1_HVT U1000 ( .A1(n882), .A3(n1614), .A2(n1613), .A4(n1178), .S0(n1164), .S1(n1162), .Y(n979) );
  NAND2X0_HVT U1001 ( .A1(n1371), .A2(n1207), .Y(n980) );
  MUX41X1_HVT U1002 ( .A1(n980), .A3(n1605), .A2(n1636), .A4(n1612), .S0(n1164), .S1(n1161), .Y(n981) );
  AO21X1_HVT U1005 ( .A1(n1610), .A2(keyin[98]), .A3(n1635), .Y(n984) );
  MUX41X1_HVT U1007 ( .A1(n1608), .A3(n984), .A2(n985), .A4(n983), .S0(n1156), 
        .S1(n1376), .Y(n986) );
  MUX41X1_HVT U1008 ( .A1(n986), .A3(n978), .A2(n982), .A4(n972), .S0(n1204), 
        .S1(keyin[103]), .Y(dummy[31]) );
  NAND2X0_HVT U1012 ( .A1(n1211), .A2(n991), .Y(n990) );
  MUX41X1_HVT U1013 ( .A1(n989), .A3(n960), .A2(n990), .A4(n940), .S0(n1156), 
        .S1(n1376), .Y(n992) );
  MUX41X1_HVT U1014 ( .A1(n1639), .A3(n1644), .A2(n1657), .A4(n1619), .S0(
        n1156), .S1(n542), .Y(n993) );
  MUX41X1_HVT U1016 ( .A1(n925), .A3(n1646), .A2(n994), .A4(n1645), .S0(n1164), 
        .S1(n1372), .Y(n995) );
  AND3X1_HVT U1019 ( .A1(n974), .A2(n1206), .A3(n999), .Y(n998) );
  MUX41X1_HVT U1021 ( .A1(n961), .A3(n1617), .A2(n1600), .A4(n930), .S0(n1156), 
        .S1(n1376), .Y(n1001) );
  AND2X1_HVT U1022 ( .A1(n1366), .A2(n1203), .Y(n1002) );
  MUX41X1_HVT U1023 ( .A1(n1618), .A3(n942), .A2(n932), .A4(n1002), .S0(n1156), 
        .S1(n1376), .Y(n1003) );
  NAND2X0_HVT U1024 ( .A1(n1371), .A2(n1656), .Y(n1004) );
  MUX41X1_HVT U1025 ( .A1(n1644), .A3(n1004), .A2(n889), .A4(n881), .S0(n1157), 
        .S1(n1376), .Y(n1005) );
  MUX41X1_HVT U1026 ( .A1(n1005), .A3(n1001), .A2(n1003), .A4(n1000), .S0(
        n1198), .S1(n1162), .Y(n1006) );
  MUX41X1_HVT U1029 ( .A1(n962), .A3(n921), .A2(n1641), .A4(n1007), .S0(n1156), 
        .S1(n1377), .Y(n1008) );
  AO21X1_HVT U1032 ( .A1(n1166), .A2(n1012), .A3(n1640), .Y(n1011) );
  MUX41X1_HVT U1035 ( .A1(n1600), .A3(n894), .A2(n1643), .A4(n1014), .S0(n1158), .S1(n1377), .Y(n1015) );
  MUX41X1_HVT U1036 ( .A1(n1639), .A3(n894), .A2(n1367), .A4(n931), .S0(n1156), 
        .S1(n1376), .Y(n1016) );
  MUX41X1_HVT U1037 ( .A1(n1016), .A3(n1013), .A2(n1015), .A4(n1008), .S0(
        keyin[103]), .S1(n1161), .Y(n1017) );
  NAND2X0_HVT U1040 ( .A1(n1021), .A2(n1022), .Y(n1020) );
  MUX41X1_HVT U1042 ( .A1(n918), .A3(n1609), .A2(n1621), .A4(n920), .S0(n1156), 
        .S1(n542), .Y(n1024) );
  MUX41X1_HVT U1044 ( .A1(n1620), .A3(n964), .A2(n1025), .A4(n1638), .S0(n1156), .S1(n1376), .Y(n1026) );
  OA21X1_HVT U1048 ( .A1(n1628), .A2(n1374), .A3(n1615), .Y(n1029) );
  NAND2X0_HVT U1049 ( .A1(n1206), .A2(n1031), .Y(n1030) );
  MUX41X1_HVT U1053 ( .A1(n1034), .A3(n1028), .A2(n1032), .A4(n1029), .S0(
        keyin[98]), .S1(n542), .Y(n1035) );
  AND2X1_HVT U1054 ( .A1(n1368), .A2(n1658), .Y(n1036) );
  AO21X1_HVT U1057 ( .A1(n1160), .A2(n1210), .A3(n942), .Y(n1039) );
  NAND2X0_HVT U1062 ( .A1(n1045), .A2(n1046), .Y(n1044) );
  MUX41X1_HVT U1064 ( .A1(n937), .A3(n906), .A2(n1608), .A4(n1648), .S0(n1157), 
        .S1(n542), .Y(n1048) );
  AND3X1_HVT U1067 ( .A1(n1158), .A2(n1371), .A3(n1203), .Y(n1051) );
  MUX41X1_HVT U1070 ( .A1(n1053), .A3(n1051), .A2(n1052), .A4(n1050), .S0(
        keyin[98]), .S1(n1379), .Y(n1054) );
  MUX41X1_HVT U1071 ( .A1(n1054), .A3(n1041), .A2(n1049), .A4(n1035), .S0(
        n1204), .S1(n1198), .Y(dummy[28]) );
  MUX41X1_HVT U1074 ( .A1(n1649), .A3(n1653), .A2(n955), .A4(n943), .S0(n1158), 
        .S1(n1377), .Y(n1057) );
  MUX41X1_HVT U1075 ( .A1(n881), .A3(n949), .A2(n1650), .A4(n951), .S0(n1157), 
        .S1(n1378), .Y(n1058) );
  MUX41X1_HVT U1078 ( .A1(n1060), .A3(n1057), .A2(n1058), .A4(n1056), .S0(
        n1198), .S1(n1161), .Y(n1061) );
  AND2X1_HVT U1079 ( .A1(n1210), .A2(n1370), .Y(n1062) );
  MUX41X1_HVT U1081 ( .A1(n1618), .A3(n1658), .A2(n1637), .A4(n1210), .S0(
        n1157), .S1(n1378), .Y(n1064) );
  OA21X1_HVT U1083 ( .A1(n1602), .A2(n1380), .A3(n947), .Y(n1066) );
  NAND2X0_HVT U1085 ( .A1(n1365), .A2(n1213), .Y(n991) );
  MUX41X1_HVT U1086 ( .A1(n1650), .A3(n991), .A2(n1639), .A4(n962), .S0(n1158), 
        .S1(n1379), .Y(n1068) );
  MUX41X1_HVT U1087 ( .A1(n1068), .A3(n1064), .A2(n1067), .A4(n1063), .S0(
        keyin[103]), .S1(n1161), .Y(n1069) );
  OA21X1_HVT U1090 ( .A1(n956), .A2(n1380), .A3(n1072), .Y(n1071) );
  AND2X1_HVT U1093 ( .A1(n1166), .A2(n1200), .Y(n1075) );
  NAND2X0_HVT U1097 ( .A1(n282), .A2(n1656), .Y(n1079) );
  MUX41X1_HVT U1098 ( .A1(n928), .A3(n1658), .A2(n1079), .A4(n1631), .S0(n1158), .S1(n1377), .Y(n1080) );
  MUX41X1_HVT U1104 ( .A1(n937), .A3(n1622), .A2(n962), .A4(n1085), .S0(n1379), 
        .S1(n1372), .Y(n1086) );
  NAND2X0_HVT U1105 ( .A1(n1213), .A2(n974), .Y(n1087) );
  NAND2X0_HVT U1106 ( .A1(n1657), .A2(n1371), .Y(n1088) );
  MUX41X1_HVT U1107 ( .A1(n1642), .A3(n1210), .A2(n1088), .A4(n1087), .S0(
        n1373), .S1(n1376), .Y(n1089) );
  OA21X1_HVT U1109 ( .A1(n900), .A2(n1380), .A3(n947), .Y(n1091) );
  NAND2X0_HVT U1113 ( .A1(n282), .A2(n942), .Y(n929) );
  MUX41X1_HVT U1115 ( .A1(n1181), .A3(n1094), .A2(n1647), .A4(n929), .S0(n1379), .S1(n1373), .Y(n1095) );
  NAND2X0_HVT U1116 ( .A1(n1365), .A2(n1181), .Y(n1096) );
  MUX41X1_HVT U1117 ( .A1(n933), .A3(n1096), .A2(n1651), .A4(n953), .S0(n1373), 
        .S1(n1379), .Y(n1097) );
  MUX41X1_HVT U1118 ( .A1(n944), .A3(n1652), .A2(n1603), .A4(n1651), .S0(n1158), .S1(n1377), .Y(n1098) );
  MUX41X1_HVT U1119 ( .A1(n1606), .A3(n925), .A2(n928), .A4(n880), .S0(n1379), 
        .S1(n1372), .Y(n1099) );
  MUX41X1_HVT U1120 ( .A1(n1099), .A3(n1097), .A2(n1098), .A4(n1095), .S0(
        keyin[103]), .S1(n1163), .Y(n1100) );
  MUX41X1_HVT U1121 ( .A1(n1630), .A3(n1209), .A2(n1633), .A4(n1634), .S0(
        n1379), .S1(n1372), .Y(n1101) );
  OA21X1_HVT U1123 ( .A1(n950), .A2(n1380), .A3(n1618), .Y(n1103) );
  MUX41X1_HVT U1125 ( .A1(n894), .A3(n954), .A2(n991), .A4(n962), .S0(n1372), 
        .S1(n542), .Y(n1105) );
  MUX41X1_HVT U1128 ( .A1(n1107), .A3(n929), .A2(n1106), .A4(n1638), .S0(n1379), .S1(n1373), .Y(n1108) );
  MUX41X1_HVT U1132 ( .A1(n921), .A3(n920), .A2(n966), .A4(n1110), .S0(n1372), 
        .S1(n1377), .Y(n1111) );
  MUX41X1_HVT U1133 ( .A1(n957), .A3(n943), .A2(n1649), .A4(n1210), .S0(n1379), 
        .S1(n1373), .Y(n1112) );
  MUX41X1_HVT U1134 ( .A1(n942), .A3(n1643), .A2(n1212), .A4(n952), .S0(n1373), 
        .S1(n1377), .Y(n1113) );
  AO21X1_HVT U1136 ( .A1(n889), .A2(n1165), .A3(n1640), .Y(n1115) );
  OA21X1_HVT U1140 ( .A1(n924), .A2(n1380), .A3(n1629), .Y(n1119) );
  MUX41X1_HVT U1142 ( .A1(n951), .A3(n1632), .A2(n927), .A4(n948), .S0(n1373), 
        .S1(n542), .Y(n1121) );
  MUX41X1_HVT U1143 ( .A1(n973), .A3(n928), .A2(n1626), .A4(n939), .S0(n1372), 
        .S1(n542), .Y(n1122) );
  MUX41X1_HVT U1144 ( .A1(n1202), .A3(n918), .A2(n1652), .A4(n1624), .S0(n1372), .S1(n542), .Y(n1123) );
  NAND2X0_HVT U1147 ( .A1(n282), .A2(n1208), .Y(n1031) );
  NAND2X0_HVT U1150 ( .A1(n1211), .A2(n1366), .Y(n974) );
  NAND2X0_HVT U1152 ( .A1(n942), .A2(n1371), .Y(n1128) );
  NAND2X0_HVT U1153 ( .A1(n1211), .A2(n1031), .Y(n1129) );
  AO21X1_HVT U1154 ( .A1(n1370), .A2(n1653), .A3(n1380), .Y(n1021) );
  NAND2X0_HVT U1156 ( .A1(n1366), .A2(n1653), .Y(n1072) );
  NAND2X0_HVT U1159 ( .A1(n1165), .A2(n1128), .Y(n999) );
  XOR2X2_HVT U1317 ( .A1(keyin[3]), .A2(dummy[3]), .Y(n1257) );
  XOR2X2_HVT U1324 ( .A1(keyin[2]), .A2(dummy[2]), .Y(n1261) );
  XOR2X2_HVT U1326 ( .A1(keyin[1]), .A2(dummy[1]), .Y(n1262) );
  XNOR2X2_HVT U1343 ( .A1(keyin[23]), .A2(dummy[23]), .Y(n1318) );
  XNOR2X2_HVT U1345 ( .A1(dummy[22]), .A2(keyin[22]), .Y(n1319) );
  XNOR2X2_HVT U1347 ( .A1(dummy[21]), .A2(keyin[21]), .Y(n1320) );
  XNOR2X2_HVT U1351 ( .A1(dummy[19]), .A2(keyin[19]), .Y(n1322) );
  XNOR2X2_HVT U1353 ( .A1(dummy[18]), .A2(keyin[18]), .Y(n1323) );
  XNOR2X2_HVT U1355 ( .A1(dummy[17]), .A2(keyin[17]), .Y(n1324) );
  XNOR2X2_HVT U1357 ( .A1(keyin[16]), .A2(dummy[16]), .Y(n1325) );
  XNOR2X2_HVT U1359 ( .A1(dummy[15]), .A2(keyin[15]), .Y(n1326) );
  XNOR2X2_HVT U1365 ( .A1(dummy[12]), .A2(keyin[12]), .Y(n1329) );
  XNOR2X2_HVT U1367 ( .A1(keyin[11]), .A2(dummy[11]), .Y(n1330) );
  XNOR2X2_HVT U1369 ( .A1(dummy[10]), .A2(keyin[10]), .Y(n1331) );
  XNOR2X2_HVT U1371 ( .A1(keyin[9]), .A2(dummy[9]), .Y(n1299) );
  XNOR2X2_HVT U1373 ( .A1(dummy[8]), .A2(keyin[8]), .Y(n1300) );
  XOR2X2_HVT U1387 ( .A1(keyin[0]), .A2(dummy[0]), .Y(n1264) );
  XNOR3X1_HVT U1430 ( .A1(keyin[32]), .A2(keyin[64]), .A3(n1295), .Y(n1265) );
  NAND3X0_HVT U1431 ( .A1(n1305), .A2(n1306), .A3(n1307), .Y(n1301) );
  NAND4X0_HVT U1432 ( .A1(round_num[1]), .A2(round_num[3]), .A3(n1383), .A4(
        n1389), .Y(n1307) );
  AO21X1_HVT U1433 ( .A1(n1311), .A2(round_num[2]), .A3(n1386), .Y(n1308) );
  NAND4X0_HVT U1434 ( .A1(round_num[1]), .A2(round_num[2]), .A3(round_num[3]), 
        .A4(n1383), .Y(n1294) );
  XNOR3X1_HVT U1435 ( .A1(n1266), .A2(keyin[127]), .A3(n1309), .Y(keyout[127])
         );
  XNOR3X1_HVT U1436 ( .A1(n1267), .A2(n212), .A3(n1310), .Y(keyout[126]) );
  XNOR3X1_HVT U1440 ( .A1(n1271), .A2(n908), .A3(n1315), .Y(keyout[122]) );
  XNOR3X1_HVT U1444 ( .A1(n1275), .A2(n1255), .A3(n1319), .Y(keyout[118]) );
  XNOR3X1_HVT U1447 ( .A1(n1278), .A2(n1187), .A3(n1322), .Y(keyout[115]) );
  XNOR3X1_HVT U1448 ( .A1(n1279), .A2(n1125), .A3(n1323), .Y(keyout[114]) );
  XNOR3X1_HVT U1449 ( .A1(n1280), .A2(keyin[113]), .A3(n1324), .Y(keyout[113])
         );
  XNOR3X1_HVT U1451 ( .A1(n1282), .A2(keyin[111]), .A3(n1326), .Y(keyout[111])
         );
  XNOR3X1_HVT U1452 ( .A1(n1283), .A2(n1355), .A3(n1327), .Y(keyout[110]) );
  XNOR3X1_HVT U1454 ( .A1(n1285), .A2(n1192), .A3(n1329), .Y(keyout[108]) );
  XNOR3X1_HVT U1455 ( .A1(n1286), .A2(n1193), .A3(n1330), .Y(keyout[107]) );
  AND2X1_HVT U1461 ( .A1(n1306), .A2(n1334), .Y(n1291) );
  NAND3X0_HVT U1462 ( .A1(n1390), .A2(n1387), .A3(round_num[2]), .Y(n1334) );
  AND2X1_HVT U1464 ( .A1(n1305), .A2(n1336), .Y(n1297) );
  NAND4X0_HVT U1465 ( .A1(round_num[2]), .A2(round_num[3]), .A3(n1383), .A4(
        n1390), .Y(n1336) );
  NAND2X0_HVT U1466 ( .A1(round_num[2]), .A2(n1337), .Y(n1305) );
  AO21X1_HVT U1468 ( .A1(n1311), .A2(n1389), .A3(n1384), .Y(n1298) );
  NAND2X0_HVT U1469 ( .A1(round_num[0]), .A2(n1332), .Y(n1306) );
  AND3X1_HVT U1470 ( .A1(n1390), .A2(n1389), .A3(round_num[3]), .Y(n1332) );
  AND3X1_HVT U1471 ( .A1(n1383), .A2(n1387), .A3(round_num[1]), .Y(n1311) );
  NAND2X0_HVT U1472 ( .A1(n1337), .A2(n1389), .Y(n1295) );
  AND3X1_HVT U1473 ( .A1(n1390), .A2(n1387), .A3(round_num[0]), .Y(n1337) );
  INVX1_HVT U1 ( .A(n1290), .Y(n23) );
  NAND2X0_HVT U2 ( .A1(n90), .A2(n49), .Y(n115) );
  NAND2X0_HVT U3 ( .A1(n82), .A2(keyin[111]), .Y(n130) );
  NAND2X0_HVT U7 ( .A1(n115), .A2(n130), .Y(dummy[6]) );
  IBUFFX2_HVT U8 ( .A(keyin[111]), .Y(n49) );
  MUX21X2_HVT U9 ( .A1(n155), .A2(n147), .S0(n211), .Y(dummy[3]) );
  IBUFFX16_HVT U10 ( .A(n601), .Y(n211) );
  INVX4_HVT U11 ( .A(keyin[117]), .Y(n1344) );
  INVX2_HVT U12 ( .A(n1344), .Y(n1342) );
  XNOR3X2_HVT U13 ( .A1(n1276), .A2(n1343), .A3(n1320), .Y(keyout[117]) );
  INVX1_HVT U14 ( .A(n1318), .Y(keyout[23]) );
  IBUFFX2_HVT U16 ( .A(n1364), .Y(n855) );
  XNOR3X2_HVT U18 ( .A1(n1270), .A2(n1184), .A3(n1314), .Y(keyout[123]) );
  IBUFFX16_HVT U19 ( .A(n1364), .Y(n1361) );
  INVX2_HVT U20 ( .A(keyin[104]), .Y(n1364) );
  XOR2X1_HVT U22 ( .A1(n1256), .A2(n1257), .Y(keyout[35]) );
  XOR3X1_HVT U23 ( .A1(n600), .A2(n824), .A3(n1321), .Y(keyout[116]) );
  INVX1_HVT U24 ( .A(n1244), .Y(n212) );
  IBUFFX2_HVT U26 ( .A(n1244), .Y(n213) );
  IBUFFX2_HVT U27 ( .A(n1244), .Y(n1243) );
  MUX21X1_HVT U28 ( .A1(n815), .A2(n814), .S0(n911), .Y(n816) );
  IBUFFX2_HVT U29 ( .A(n634), .Y(n1419) );
  MUX21X2_HVT U30 ( .A1(n718), .A2(n717), .S0(n1246), .Y(n719) );
  MUX21X2_HVT U31 ( .A1(n628), .A2(n715), .S0(n912), .Y(n716) );
  IBUFFX16_HVT U32 ( .A(n1244), .Y(n1240) );
  INVX2_HVT U35 ( .A(keyin[126]), .Y(n1244) );
  NAND2X2_HVT U36 ( .A1(n757), .A2(n214), .Y(n217) );
  NAND2X0_HVT U37 ( .A1(n765), .A2(n220), .Y(n218) );
  NAND2X0_HVT U38 ( .A1(n217), .A2(n218), .Y(dummy[19]) );
  INVX1_HVT U40 ( .A(n220), .Y(n214) );
  IBUFFX2_HVT U41 ( .A(n604), .Y(n220) );
  INVX1_HVT U42 ( .A(n1320), .Y(keyout[21]) );
  MUX21X2_HVT U43 ( .A1(n885), .A2(n716), .S0(n913), .Y(n717) );
  MUX21X2_HVT U44 ( .A1(n798), .A2(n805), .S0(n219), .Y(dummy[17]) );
  IBUFFX16_HVT U45 ( .A(n604), .Y(n219) );
  MUX21X2_HVT U46 ( .A1(n761), .A2(n762), .S0(n912), .Y(n763) );
  MUX21X1_HVT U47 ( .A1(n336), .A2(n1489), .S0(n1344), .Y(n441) );
  INVX2_HVT U48 ( .A(n1319), .Y(keyout[22]) );
  XOR2X2_HVT U49 ( .A1(keyin[49]), .A2(keyout[17]), .Y(keyout[49]) );
  MUX21X1_HVT U51 ( .A1(n233), .A2(n833), .S0(n234), .Y(n232) );
  IBUFFX16_HVT U53 ( .A(n232), .Y(n814) );
  IBUFFX16_HVT U54 ( .A(n647), .Y(n233) );
  IBUFFX16_HVT U58 ( .A(n913), .Y(n234) );
  MUX41X1_HVT U63 ( .A1(n816), .A3(n818), .A2(n817), .A4(n819), .S0(n235), 
        .S1(n1247), .Y(n820) );
  IBUFFX16_HVT U64 ( .A(keyin[121]), .Y(n235) );
  INVX1_HVT U66 ( .A(n1247), .Y(n1246) );
  IBUFFX2_HVT U68 ( .A(n614), .Y(n1405) );
  NAND2X2_HVT U70 ( .A1(n1241), .A2(n1216), .Y(n614) );
  NAND2X0_HVT U72 ( .A1(n438), .A2(n236), .Y(n237) );
  NAND2X0_HVT U73 ( .A1(n437), .A2(n1133), .Y(n238) );
  NAND2X0_HVT U74 ( .A1(n237), .A2(n238), .Y(n439) );
  IBUFFX2_HVT U76 ( .A(n1133), .Y(n236) );
  NAND2X0_HVT U79 ( .A1(n436), .A2(n239), .Y(n240) );
  NAND2X0_HVT U87 ( .A1(n439), .A2(n244), .Y(n241) );
  NAND2X0_HVT U88 ( .A1(n240), .A2(n241), .Y(n440) );
  INVX0_HVT U89 ( .A(n244), .Y(n239) );
  XOR2X2_HVT U90 ( .A1(keyout[12]), .A2(n1285), .Y(keyout[76]) );
  NBUFFX4_HVT U91 ( .A(n1349), .Y(n1133) );
  IBUFFX2_HVT U92 ( .A(n1130), .Y(n244) );
  MUX21X2_HVT U95 ( .A1(n813), .A2(n820), .S0(n242), .Y(dummy[16]) );
  IBUFFX16_HVT U96 ( .A(n604), .Y(n242) );
  MUX21X2_HVT U99 ( .A1(n684), .A2(n657), .S0(n608), .Y(n761) );
  XOR2X2_HVT U100 ( .A1(keyin[55]), .A2(keyout[23]), .Y(keyout[55]) );
  MUX21X2_HVT U101 ( .A1(n428), .A2(n429), .S0(n243), .Y(n432) );
  IBUFFX16_HVT U103 ( .A(n538), .Y(n243) );
  INVX2_HVT U105 ( .A(n1325), .Y(keyout[16]) );
  INVX1_HVT U107 ( .A(n833), .Y(n1443) );
  MUX21X2_HVT U108 ( .A1(n433), .A2(n432), .S0(n1130), .Y(n434) );
  XOR3X2_HVT U109 ( .A1(n1274), .A2(n294), .A3(n1318), .Y(keyout[119]) );
  INVX1_HVT U110 ( .A(keyin[119]), .Y(n294) );
  MUX41X1_HVT U112 ( .A1(n749), .A3(n747), .A2(n748), .A4(n746), .S0(n297), 
        .S1(n245), .Y(n750) );
  IBUFFX16_HVT U113 ( .A(n296), .Y(n245) );
  INVX1_HVT U114 ( .A(n472), .Y(n297) );
  INVX1_HVT U115 ( .A(n8), .Y(n246) );
  INVX2_HVT U116 ( .A(n246), .Y(n247) );
  AO21X1_HVT U117 ( .A1(n249), .A2(keyin[104]), .A3(n250), .Y(n248) );
  IBUFFX16_HVT U119 ( .A(n248), .Y(n186) );
  IBUFFX16_HVT U121 ( .A(n33), .Y(n249) );
  IBUFFX16_HVT U122 ( .A(n1549), .Y(n250) );
  XNOR2X2_HVT U123 ( .A1(keyin[50]), .A2(n1323), .Y(keyout[50]) );
  INVX1_HVT U124 ( .A(n1323), .Y(keyout[18]) );
  XOR2X2_HVT U126 ( .A1(n1586), .A2(n1193), .Y(n8) );
  INVX0_HVT U127 ( .A(n8), .Y(n1584) );
  NBUFFX2_HVT U128 ( .A(n288), .Y(n251) );
  NBUFFX4_HVT U130 ( .A(keyin[125]), .Y(n288) );
  IBUFFX2_HVT U131 ( .A(n1356), .Y(n252) );
  IBUFFX2_HVT U135 ( .A(n1356), .Y(n253) );
  MUX21X1_HVT U136 ( .A1(n1245), .A2(n614), .S0(n1247), .Y(n736) );
  XNOR2X2_HVT U141 ( .A1(n1322), .A2(n1278), .Y(keyout[83]) );
  INVX1_HVT U142 ( .A(n1322), .Y(keyout[19]) );
  INVX1_HVT U145 ( .A(n599), .Y(n254) );
  MUX41X1_HVT U147 ( .A1(n189), .A3(n192), .A2(n190), .A4(n194), .S0(n255), 
        .S1(n256), .Y(n195) );
  IBUFFX16_HVT U150 ( .A(n1196), .Y(n255) );
  IBUFFX16_HVT U152 ( .A(n271), .Y(n256) );
  XOR2X2_HVT U154 ( .A1(n1319), .A2(n257), .Y(keyout[86]) );
  IBUFFX16_HVT U155 ( .A(n1275), .Y(n257) );
  INVX1_HVT U157 ( .A(n1351), .Y(n258) );
  INVX1_HVT U162 ( .A(n1351), .Y(n259) );
  MUX21X1_HVT U163 ( .A1(n262), .A2(n261), .S0(n263), .Y(n260) );
  IBUFFX16_HVT U164 ( .A(n260), .Y(n404) );
  IBUFFX16_HVT U168 ( .A(n322), .Y(n261) );
  IBUFFX16_HVT U170 ( .A(n875), .Y(n262) );
  IBUFFX16_HVT U173 ( .A(n1134), .Y(n263) );
  INVX1_HVT U174 ( .A(n1351), .Y(n1347) );
  XOR2X1_HVT U178 ( .A1(n1325), .A2(n270), .Y(keyout[80]) );
  INVX2_HVT U181 ( .A(n296), .Y(n264) );
  IBUFFX2_HVT U182 ( .A(n264), .Y(n587) );
  INVX1_HVT U183 ( .A(keyin[120]), .Y(n296) );
  INVX1_HVT U187 ( .A(n280), .Y(n265) );
  NBUFFX2_HVT U189 ( .A(n1132), .Y(n266) );
  INVX0_HVT U191 ( .A(n1347), .Y(n280) );
  IBUFFX16_HVT U192 ( .A(n1351), .Y(n1348) );
  INVX1_HVT U193 ( .A(n1340), .Y(n267) );
  INVX1_HVT U197 ( .A(n1340), .Y(n268) );
  MUX21X1_HVT U199 ( .A1(n312), .A2(n1228), .S0(n1341), .Y(n269) );
  IBUFFX16_HVT U201 ( .A(n269), .Y(n344) );
  IBUFFX16_HVT U203 ( .A(n1281), .Y(n270) );
  INVX0_HVT U208 ( .A(n1360), .Y(n271) );
  INVX1_HVT U209 ( .A(n1360), .Y(n272) );
  INVX0_HVT U210 ( .A(n1360), .Y(n1358) );
  MUX21X1_HVT U213 ( .A1(n1510), .A2(n342), .S0(n1132), .Y(n509) );
  MUX21X2_HVT U214 ( .A1(n738), .A2(n737), .S0(n273), .Y(n739) );
  IBUFFX16_HVT U217 ( .A(n289), .Y(n273) );
  MUX41X1_HVT U220 ( .A1(n739), .A3(n731), .A2(n750), .A4(n745), .S0(n274), 
        .S1(n354), .Y(dummy[20]) );
  IBUFFX16_HVT U222 ( .A(n328), .Y(n274) );
  XNOR2X2_HVT U223 ( .A1(keyin[53]), .A2(n1320), .Y(keyout[53]) );
  INVX1_HVT U224 ( .A(keyin[118]), .Y(n1340) );
  XNOR2X1_HVT U225 ( .A1(n275), .A2(n1351), .Y(n895) );
  IBUFFX16_HVT U226 ( .A(n287), .Y(n275) );
  NAND2X0_HVT U227 ( .A1(n593), .A2(n279), .Y(n276) );
  AND2X1_HVT U228 ( .A1(n276), .A2(n277), .Y(n399) );
  OR2X4_HVT U229 ( .A1(n278), .A2(n895), .Y(n277) );
  INVX1_HVT U230 ( .A(n586), .Y(n278) );
  AND2X1_HVT U231 ( .A1(n592), .A2(n586), .Y(n279) );
  IBUFFX4_HVT U232 ( .A(n1351), .Y(n1350) );
  XOR3X2_HVT U233 ( .A1(n1281), .A2(n280), .A3(n1325), .Y(keyout[112]) );
  XOR2X2_HVT U234 ( .A1(keyout[23]), .A2(n1274), .Y(keyout[87]) );
  XNOR2X2_HVT U235 ( .A1(keyin[44]), .A2(n1329), .Y(keyout[44]) );
  INVX1_HVT U236 ( .A(n1329), .Y(keyout[12]) );
  XNOR2X2_HVT U237 ( .A1(n1327), .A2(n1283), .Y(keyout[78]) );
  INVX0_HVT U238 ( .A(n1370), .Y(n281) );
  INVX0_HVT U239 ( .A(n1370), .Y(n282) );
  INVX0_HVT U240 ( .A(n1370), .Y(n1367) );
  MUX21X2_HVT U241 ( .A1(n880), .A2(n932), .S0(n283), .Y(n1118) );
  IBUFFX16_HVT U242 ( .A(n1164), .Y(n283) );
  MUX41X1_HVT U243 ( .A1(n1120), .A3(n1122), .A2(n1121), .A4(n1123), .S0(n284), 
        .S1(n285), .Y(n1124) );
  IBUFFX16_HVT U244 ( .A(n1198), .Y(n284) );
  IBUFFX16_HVT U245 ( .A(n1163), .Y(n285) );
  INVX1_HVT U246 ( .A(keyin[118]), .Y(n286) );
  INVX0_HVT U247 ( .A(keyin[118]), .Y(n287) );
  IBUFFX16_HVT U248 ( .A(n911), .Y(n289) );
  INVX1_HVT U249 ( .A(keyin[125]), .Y(n1247) );
  IBUFFX16_HVT U250 ( .A(n1370), .Y(n1366) );
  INVX0_HVT U251 ( .A(n287), .Y(n1339) );
  MUX41X1_HVT U252 ( .A1(n988), .A3(n993), .A2(n992), .A4(n995), .S0(n290), 
        .S1(n291), .Y(n996) );
  IBUFFX16_HVT U253 ( .A(n1198), .Y(n290) );
  IBUFFX16_HVT U254 ( .A(n1162), .Y(n291) );
  XOR2X2_HVT U255 ( .A1(keyout[15]), .A2(n1282), .Y(keyout[79]) );
  XNOR3X1_HVT U256 ( .A1(n1263), .A2(n1204), .A3(n1262), .Y(keyout[97]) );
  MUX21X2_HVT U257 ( .A1(n188), .A2(n195), .S0(n292), .Y(dummy[1]) );
  IBUFFX16_HVT U258 ( .A(keyin[111]), .Y(n292) );
  MUX41X1_HVT U259 ( .A1(n361), .A3(n365), .A2(n371), .A4(n375), .S0(n293), 
        .S1(n294), .Y(dummy[15]) );
  IBUFFX16_HVT U260 ( .A(n1190), .Y(n293) );
  INVX2_HVT U261 ( .A(n1370), .Y(n1368) );
  INVX2_HVT U262 ( .A(keyin[102]), .Y(n1370) );
  IBUFFX2_HVT U263 ( .A(n1254), .Y(n608) );
  MUX21X1_HVT U264 ( .A1(n733), .A2(n734), .S0(n608), .Y(n737) );
  INVX2_HVT U265 ( .A(n1351), .Y(n1349) );
  INVX2_HVT U266 ( .A(keyin[112]), .Y(n1351) );
  MUX21X1_HVT U267 ( .A1(n382), .A2(n383), .S0(n1131), .Y(n385) );
  MUX21X1_HVT U268 ( .A1(n1486), .A2(n322), .S0(n1133), .Y(n382) );
  INVX1_HVT U269 ( .A(n1244), .Y(n1239) );
  INVX1_HVT U270 ( .A(n1244), .Y(n1241) );
  INVX2_HVT U271 ( .A(n1244), .Y(n1242) );
  MUX21X1_HVT U272 ( .A1(n1426), .A2(n630), .S0(n1247), .Y(n749) );
  XNOR2X1_HVT U273 ( .A1(n1321), .A2(n295), .Y(keyout[84]) );
  IBUFFX16_HVT U274 ( .A(n600), .Y(n295) );
  IBUFFX2_HVT U275 ( .A(n1321), .Y(keyout[20]) );
  AND3X2_HVT U276 ( .A1(n1246), .A2(n1245), .A3(n1185), .Y(n747) );
  AO21X2_HVT U277 ( .A1(n1246), .A2(n1218), .A3(n618), .Y(n743) );
  NAND2X0_HVT U278 ( .A1(n741), .A2(n297), .Y(n298) );
  NAND2X0_HVT U279 ( .A1(n744), .A2(n472), .Y(n299) );
  NAND2X0_HVT U280 ( .A1(n299), .A2(n298), .Y(n745) );
  MUX21X1_HVT U281 ( .A1(n743), .A2(n742), .S0(n914), .Y(n744) );
  IBUFFX2_HVT U282 ( .A(n909), .Y(n472) );
  XOR2X2_HVT U283 ( .A1(keyin[47]), .A2(keyout[15]), .Y(keyout[47]) );
  MUX41X1_HVT U284 ( .A1(n304), .A3(n301), .A2(n303), .A4(n302), .S0(n1360), 
        .S1(n855), .Y(n300) );
  IBUFFX16_HVT U285 ( .A(n300), .Y(n131) );
  IBUFFX16_HVT U286 ( .A(n15), .Y(n301) );
  IBUFFX16_HVT U287 ( .A(n1550), .Y(n302) );
  IBUFFX16_HVT U288 ( .A(n30), .Y(n303) );
  NAND2X0_HVT U289 ( .A1(n1355), .A2(n1174), .Y(n304) );
  MUX21X2_HVT U290 ( .A1(n131), .A2(n134), .S0(n305), .Y(n135) );
  IBUFFX16_HVT U291 ( .A(n1152), .Y(n305) );
  IBUFFX16_HVT U292 ( .A(keyin[121]), .Y(n328) );
  IBUFFX16_HVT U293 ( .A(n604), .Y(n354) );
  XOR3X2_HVT U294 ( .A1(n1385), .A2(n605), .A3(n398), .Y(keyout[102]) );
  XNOR2X1_HVT U295 ( .A1(keyin[70]), .A2(n1369), .Y(n398) );
  XNOR3X1_HVT U296 ( .A1(n1382), .A2(n1335), .A3(n865), .Y(keyout[101]) );
  INVX4_HVT U297 ( .A(keyin[109]), .Y(n1360) );
  MUX41X1_HVT U298 ( .A1(n1625), .A3(n1062), .A2(n1629), .A4(n941), .S0(n516), 
        .S1(n1381), .Y(n1063) );
  IBUFFX16_HVT U299 ( .A(n1158), .Y(n516) );
  NAND2X0_HVT U300 ( .A1(keyin[32]), .A2(n518), .Y(n519) );
  NAND2X0_HVT U301 ( .A1(n517), .A2(keyout[0]), .Y(n522) );
  NAND2X0_HVT U302 ( .A1(n519), .A2(n522), .Y(keyout[32]) );
  IBUFFX2_HVT U303 ( .A(keyin[32]), .Y(n517) );
  INVX1_HVT U304 ( .A(keyout[0]), .Y(n518) );
  INVX2_HVT U305 ( .A(n1356), .Y(n1354) );
  INVX2_HVT U306 ( .A(keyin[110]), .Y(n1356) );
  XNOR2X2_HVT U307 ( .A1(n523), .A2(n1292), .Y(n606) );
  IBUFFX16_HVT U308 ( .A(n1293), .Y(n523) );
  IBUFFX2_HVT U309 ( .A(keyin[109]), .Y(n574) );
  INVX4_HVT U310 ( .A(n1381), .Y(n1378) );
  MUX21X1_HVT U311 ( .A1(n128), .A2(n127), .S0(n1152), .Y(n129) );
  NBUFFX2_HVT U312 ( .A(n1354), .Y(n524) );
  NBUFFX2_HVT U313 ( .A(n1354), .Y(n525) );
  NBUFFX2_HVT U314 ( .A(n1354), .Y(n537) );
  IBUFFX2_HVT U315 ( .A(n1356), .Y(n1353) );
  NAND2X0_HVT U316 ( .A1(n506), .A2(n1126), .Y(n583) );
  OA21X1_HVT U321 ( .A1(n314), .A2(n538), .A3(n269), .Y(n506) );
  MUX41X1_HVT U322 ( .A1(n1516), .A3(n339), .A2(n1226), .A4(n501), .S0(n1127), 
        .S1(n1347), .Y(n502) );
  NAND2X0_HVT U323 ( .A1(n491), .A2(n561), .Y(n540) );
  OA21X1_HVT U324 ( .A1(n338), .A2(n538), .A3(n1487), .Y(n491) );
  INVX1_HVT U325 ( .A(n1360), .Y(n1359) );
  INVX1_HVT U326 ( .A(n1380), .Y(n542) );
  IBUFFX2_HVT U327 ( .A(n1380), .Y(n1376) );
  INVX1_HVT U329 ( .A(keyin[13]), .Y(n572) );
  MUX21X1_HVT U331 ( .A1(n591), .A2(n1525), .S0(n895), .Y(n590) );
  OA21X1_HVT U332 ( .A1(n346), .A2(n538), .A3(n464), .Y(n463) );
  INVX1_HVT U333 ( .A(keyin[112]), .Y(n538) );
  NAND2X0_HVT U335 ( .A1(n508), .A2(n557), .Y(n596) );
  NAND2X0_HVT U336 ( .A1(n500), .A2(n597), .Y(n553) );
  NAND2X0_HVT U337 ( .A1(n1027), .A2(n580), .Y(n578) );
  INVX1_HVT U339 ( .A(n1315), .Y(keyout[26]) );
  INVX0_HVT U340 ( .A(n1269), .Y(n555) );
  INVX0_HVT U341 ( .A(n575), .Y(n573) );
  INVX1_HVT U342 ( .A(n1284), .Y(n575) );
  INVX1_HVT U343 ( .A(n1163), .Y(n545) );
  INVX1_HVT U344 ( .A(n938), .Y(n561) );
  INVX0_HVT U345 ( .A(n942), .Y(n1658) );
  INVX1_HVT U348 ( .A(n1198), .Y(n562) );
  INVX0_HVT U349 ( .A(n1157), .Y(n556) );
  INVX1_HVT U350 ( .A(keyin[97]), .Y(n580) );
  INVX0_HVT U351 ( .A(n580), .Y(n567) );
  INVX1_HVT U353 ( .A(keyin[119]), .Y(n597) );
  INVX0_HVT U354 ( .A(n597), .Y(n557) );
  INVX1_HVT U355 ( .A(n1344), .Y(n1343) );
  INVX0_HVT U356 ( .A(n1343), .Y(n560) );
  INVX1_HVT U357 ( .A(n1189), .Y(n598) );
  NBUFFX2_HVT U358 ( .A(n1349), .Y(n1134) );
  INVX1_HVT U359 ( .A(n855), .Y(n599) );
  INVX1_HVT U360 ( .A(n1300), .Y(keyout[8]) );
  MUX21X2_HVT U361 ( .A1(n1573), .A2(n37), .S0(n1154), .Y(n204) );
  XOR3X1_HVT U362 ( .A1(keyin[66]), .A2(n1260), .A3(n869), .Y(keyout[66]) );
  INVX2_HVT U364 ( .A(keyin[96]), .Y(n1381) );
  MUX21X1_HVT U366 ( .A1(n205), .A2(n204), .S0(n1152), .Y(n206) );
  MUX21X1_HVT U367 ( .A1(n352), .A2(n1508), .S0(n1134), .Y(n400) );
  MUX21X2_HVT U371 ( .A1(n510), .A2(n509), .S0(n938), .Y(n511) );
  XOR2X2_HVT U376 ( .A1(n539), .A2(dummy[14]), .Y(n1327) );
  IBUFFX16_HVT U377 ( .A(keyin[14]), .Y(n539) );
  INVX1_HVT U379 ( .A(n223), .Y(n1573) );
  MUX21X2_HVT U381 ( .A1(n210), .A2(n203), .S0(keyin[111]), .Y(dummy[0]) );
  MUX41X1_HVT U383 ( .A1(n400), .A3(n397), .A2(n401), .A4(n399), .S0(
        keyin[117]), .S1(n561), .Y(n403) );
  MUX41X1_HVT U385 ( .A1(n492), .A3(n489), .A2(n488), .A4(n486), .S0(n1343), 
        .S1(n1190), .Y(n493) );
  NAND2X0_HVT U386 ( .A1(n490), .A2(n1131), .Y(n541) );
  NAND2X0_HVT U387 ( .A1(n540), .A2(n541), .Y(n492) );
  XNOR2X1_HVT U389 ( .A1(dummy[6]), .A2(keyin[6]), .Y(n1290) );
  IBUFFX2_HVT U392 ( .A(n17), .Y(n1545) );
  MUX21X2_HVT U400 ( .A1(n1548), .A2(n17), .S0(n1155), .Y(n77) );
  MUX41X1_HVT U401 ( .A1(n1036), .A3(n947), .A2(n928), .A4(n1619), .S0(n1377), 
        .S1(n556), .Y(n1037) );
  INVX2_HVT U402 ( .A(n1380), .Y(n1377) );
  MUX21X1_HVT U403 ( .A1(n1040), .A2(n1037), .S0(n1375), .Y(n1041) );
  XOR2X2_HVT U404 ( .A1(n1313), .A2(n555), .Y(keyout[92]) );
  NAND2X0_HVT U405 ( .A1(n1100), .A2(n567), .Y(n543) );
  NAND2X0_HVT U407 ( .A1(n1109), .A2(n580), .Y(n544) );
  NAND2X0_HVT U408 ( .A1(n543), .A2(n544), .Y(dummy[25]) );
  MUX41X1_HVT U409 ( .A1(n1092), .A3(n1086), .A2(n1089), .A4(n1084), .S0(
        keyin[103]), .S1(n1161), .Y(n1093) );
  INVX2_HVT U411 ( .A(n1309), .Y(keyout[31]) );
  XNOR2X2_HVT U412 ( .A1(keyin[31]), .A2(dummy[31]), .Y(n1309) );
  MUX21X2_HVT U413 ( .A1(n971), .A2(n967), .S0(n1159), .Y(n972) );
  XNOR2X2_HVT U414 ( .A1(keyin[57]), .A2(n1316), .Y(keyout[57]) );
  XOR3X2_HVT U416 ( .A1(n1272), .A2(n860), .A3(n1316), .Y(keyout[121]) );
  XOR2X2_HVT U418 ( .A1(keyout[11]), .A2(n1286), .Y(keyout[75]) );
  MUX41X1_HVT U420 ( .A1(n1111), .A3(n1113), .A2(n1112), .A4(n1116), .S0(n562), 
        .S1(n545), .Y(n1117) );
  XNOR2X2_HVT U421 ( .A1(keyin[61]), .A2(n1312), .Y(keyout[61]) );
  INVX1_HVT U422 ( .A(n1312), .Y(keyout[29]) );
  XOR2X2_HVT U425 ( .A1(keyout[31]), .A2(n1266), .Y(keyout[95]) );
  MUX41X1_HVT U426 ( .A1(n511), .A3(n513), .A2(n512), .A4(n514), .S0(n598), 
        .S1(n1344), .Y(n515) );
  INVX0_HVT U427 ( .A(n1316), .Y(keyout[25]) );
  OR2X1_HVT U428 ( .A1(n1321), .A2(keyin[52]), .Y(n822) );
  AND3X2_HVT U429 ( .A1(n1342), .A2(n1341), .A3(n1188), .Y(n442) );
  AO21X2_HVT U430 ( .A1(n1342), .A2(n1227), .A3(n313), .Y(n438) );
  NAND2X0_HVT U432 ( .A1(n552), .A2(keyout[8]), .Y(n548) );
  NAND2X0_HVT U434 ( .A1(n546), .A2(n1300), .Y(n549) );
  NAND2X0_HVT U437 ( .A1(n548), .A2(n549), .Y(keyout[40]) );
  INVX1_HVT U438 ( .A(n552), .Y(n546) );
  IBUFFX2_HVT U439 ( .A(keyin[40]), .Y(n552) );
  XNOR3X1_HVT U440 ( .A1(n1269), .A2(n1183), .A3(n1313), .Y(keyout[124]) );
  NAND2X0_HVT U441 ( .A1(n866), .A2(n867), .Y(n475) );
  NAND2X1_HVT U442 ( .A1(n395), .A2(n597), .Y(n550) );
  NAND2X0_HVT U443 ( .A1(n387), .A2(n557), .Y(n551) );
  NAND2X0_HVT U444 ( .A1(n550), .A2(n551), .Y(dummy[14]) );
  XOR2X2_HVT U446 ( .A1(keyin[63]), .A2(keyout[31]), .Y(keyout[63]) );
  NAND2X0_HVT U448 ( .A1(n493), .A2(n557), .Y(n554) );
  NAND2X0_HVT U449 ( .A1(n553), .A2(n554), .Y(dummy[9]) );
  INVX1_HVT U454 ( .A(n1313), .Y(keyout[28]) );
  XOR2X2_HVT U455 ( .A1(keyout[9]), .A2(n1288), .Y(keyout[73]) );
  NAND2X0_HVT U458 ( .A1(n452), .A2(n557), .Y(n558) );
  NAND2X0_HVT U459 ( .A1(n460), .A2(n597), .Y(n559) );
  NAND2X0_HVT U460 ( .A1(n558), .A2(n559), .Y(dummy[11]) );
  MUX41X1_HVT U463 ( .A1(n404), .A3(n405), .A2(n1493), .A4(n406), .S0(n560), 
        .S1(n561), .Y(n409) );
  INVX1_HVT U465 ( .A(n531), .Y(n1493) );
  MUX41X1_HVT U466 ( .A1(n1101), .A3(n1104), .A2(n1105), .A4(n1108), .S0(n545), 
        .S1(n562), .Y(n1109) );
  NAND2X0_HVT U467 ( .A1(n480), .A2(n561), .Y(n563) );
  NAND2X0_HVT U468 ( .A1(n479), .A2(n1130), .Y(n564) );
  NAND2X0_HVT U470 ( .A1(n563), .A2(n564), .Y(n481) );
  NAND2X0_HVT U474 ( .A1(n317), .A2(n1134), .Y(n565) );
  NAND2X0_HVT U475 ( .A1(n341), .A2(n538), .Y(n566) );
  NAND2X0_HVT U476 ( .A1(n565), .A2(n566), .Y(n505) );
  MUX41X1_HVT U477 ( .A1(n507), .A3(n503), .A2(n504), .A4(n502), .S0(
        keyin[113]), .S1(n1343), .Y(n508) );
  NAND2X0_HVT U481 ( .A1(n1081), .A2(n567), .Y(n568) );
  NAND2X0_HVT U482 ( .A1(n1093), .A2(n580), .Y(n569) );
  NAND2X0_HVT U483 ( .A1(n568), .A2(n569), .Y(dummy[26]) );
  MUX41X1_HVT U486 ( .A1(n481), .A3(n475), .A2(n483), .A4(n477), .S0(n1190), 
        .S1(n560), .Y(n484) );
  NAND2X0_HVT U487 ( .A1(n1069), .A2(n580), .Y(n570) );
  NAND2X0_HVT U491 ( .A1(n1061), .A2(n567), .Y(n571) );
  NAND2X0_HVT U494 ( .A1(n570), .A2(n571), .Y(dummy[27]) );
  XOR2X2_HVT U495 ( .A1(n572), .A2(dummy[13]), .Y(n1328) );
  XOR3X2_HVT U496 ( .A1(n573), .A2(n574), .A3(n1328), .Y(keyout[109]) );
  NAND2X0_HVT U497 ( .A1(n1006), .A2(n580), .Y(n576) );
  NAND2X0_HVT U500 ( .A1(n996), .A2(n1204), .Y(n577) );
  NAND2X0_HVT U502 ( .A1(n576), .A2(n577), .Y(dummy[30]) );
  MUX41X1_HVT U505 ( .A1(n1080), .A3(n1074), .A2(n1078), .A4(n1073), .S0(
        keyin[103]), .S1(n1163), .Y(n1081) );
  NAND2X0_HVT U506 ( .A1(n1017), .A2(keyin[97]), .Y(n579) );
  NAND2X0_HVT U507 ( .A1(n578), .A2(n579), .Y(dummy[29]) );
  NAND2X0_HVT U510 ( .A1(n515), .A2(n597), .Y(n595) );
  NAND2X0_HVT U511 ( .A1(n1124), .A2(n580), .Y(n581) );
  NAND2X0_HVT U512 ( .A1(n1117), .A2(keyin[97]), .Y(n582) );
  NAND2X0_HVT U513 ( .A1(n581), .A2(n582), .Y(dummy[24]) );
  XNOR2X2_HVT U514 ( .A1(n1315), .A2(n1271), .Y(keyout[90]) );
  XOR2X2_HVT U516 ( .A1(n1265), .A2(n1264), .Y(keyout[64]) );
  XOR2X2_HVT U520 ( .A1(keyin[58]), .A2(keyout[26]), .Y(keyout[58]) );
  XNOR2X2_HVT U521 ( .A1(keyin[30]), .A2(dummy[30]), .Y(n1310) );
  NAND2X0_HVT U522 ( .A1(n505), .A2(n561), .Y(n584) );
  NAND2X0_HVT U523 ( .A1(n583), .A2(n584), .Y(n507) );
  XOR2X2_HVT U526 ( .A1(keyin[59]), .A2(keyout[27]), .Y(keyout[59]) );
  INVX2_HVT U527 ( .A(n1314), .Y(keyout[27]) );
  XOR3X2_HVT U530 ( .A1(n1288), .A2(n603), .A3(n1299), .Y(keyout[105]) );
  NAND2X0_HVT U531 ( .A1(n1223), .A2(n585), .Y(n586) );
  INVX0_HVT U533 ( .A(n895), .Y(n585) );
  XOR2X2_HVT U535 ( .A1(keyin[41]), .A2(keyout[9]), .Y(keyout[41]) );
  INVX2_HVT U536 ( .A(n1299), .Y(keyout[9]) );
  XOR2X2_HVT U537 ( .A1(keyin[46]), .A2(keyout[14]), .Y(keyout[46]) );
  XOR3X2_HVT U538 ( .A1(n1273), .A2(n587), .A3(n1317), .Y(keyout[120]) );
  NAND2X2_HVT U539 ( .A1(n471), .A2(n557), .Y(n588) );
  NAND2X0_HVT U540 ( .A1(n484), .A2(n597), .Y(n589) );
  NAND2X0_HVT U541 ( .A1(n589), .A2(n588), .Y(dummy[10]) );
  XOR2X2_HVT U542 ( .A1(keyin[43]), .A2(keyout[11]), .Y(keyout[43]) );
  INVX2_HVT U543 ( .A(n1330), .Y(keyout[11]) );
  MUX21X2_HVT U544 ( .A1(n311), .A2(n453), .S0(n1131), .Y(n454) );
  XOR2X2_HVT U545 ( .A1(keyin[62]), .A2(keyout[30]), .Y(keyout[62]) );
  INVX2_HVT U546 ( .A(n1310), .Y(keyout[30]) );
  XNOR2X2_HVT U547 ( .A1(n1331), .A2(n1287), .Y(keyout[74]) );
  IBUFFX2_HVT U548 ( .A(n1331), .Y(keyout[10]) );
  INVX1_HVT U549 ( .A(n590), .Y(n473) );
  NAND2X0_HVT U550 ( .A1(n1134), .A2(n824), .Y(n591) );
  INVX2_HVT U551 ( .A(n1317), .Y(keyout[24]) );
  XOR2X2_HVT U552 ( .A1(keyin[56]), .A2(keyout[24]), .Y(keyout[56]) );
  NAND2X0_HVT U553 ( .A1(n1186), .A2(n538), .Y(n592) );
  NAND2X0_HVT U554 ( .A1(n1526), .A2(n1134), .Y(n593) );
  XOR2X2_HVT U555 ( .A1(dummy[13]), .A2(keyin[13]), .Y(keyout[13]) );
  XNOR2X2_HVT U556 ( .A1(n1328), .A2(keyin[45]), .Y(keyout[45]) );
  XOR2X2_HVT U557 ( .A1(keyout[24]), .A2(n1273), .Y(keyout[88]) );
  XNOR2X2_HVT U558 ( .A1(keyin[24]), .A2(dummy[24]), .Y(n1317) );
  INVX2_HVT U559 ( .A(n1327), .Y(keyout[14]) );
  NAND2X0_HVT U560 ( .A1(n595), .A2(n596), .Y(dummy[8]) );
  MUX41X1_HVT U561 ( .A1(n403), .A3(n414), .A2(n409), .A4(n418), .S0(n597), 
        .S1(n598), .Y(dummy[13]) );
  XOR2X2_HVT U562 ( .A1(keyout[30]), .A2(n1267), .Y(keyout[94]) );
  MUX21X1_HVT U563 ( .A1(n122), .A2(n1531), .S0(n1360), .Y(n123) );
  MUX21X2_HVT U564 ( .A1(n124), .A2(n123), .S0(n599), .Y(n127) );
  XOR2X2_HVT U565 ( .A1(n1293), .A2(n1527), .Y(keyout[36]) );
  INVX1_HVT U566 ( .A(n1254), .Y(n1253) );
  XOR2X1_HVT U567 ( .A1(n618), .A2(n1242), .Y(n657) );
  INVX1_HVT U568 ( .A(keyin[120]), .Y(n1254) );
  INVX1_HVT U569 ( .A(n1082), .Y(n633) );
  INVX0_HVT U570 ( .A(n114), .Y(n843) );
  MUX21X1_HVT U571 ( .A1(n1551), .A2(n31), .S0(n1358), .Y(n136) );
  XOR2X1_HVT U572 ( .A1(n1373), .A2(n1369), .Y(n965) );
  INVX0_HVT U573 ( .A(keyin[42]), .Y(n856) );
  INVX1_HVT U574 ( .A(n829), .Y(n870) );
  INVX1_HVT U575 ( .A(n118), .Y(n844) );
  MUX21X1_HVT U576 ( .A1(n1530), .A2(n1557), .S0(n1358), .Y(n132) );
  NAND2X0_HVT U577 ( .A1(n474), .A2(n561), .Y(n866) );
  NAND2X0_HVT U578 ( .A1(n779), .A2(n862), .Y(n863) );
  INVX0_HVT U579 ( .A(n609), .Y(n1084) );
  INVX1_HVT U580 ( .A(n888), .Y(n610) );
  INVX1_HVT U581 ( .A(n1150), .Y(n845) );
  INVX1_HVT U582 ( .A(keyin[20]), .Y(n849) );
  INVX0_HVT U583 ( .A(keyin[121]), .Y(n860) );
  INVX0_HVT U584 ( .A(n1308), .Y(n858) );
  INVX0_HVT U585 ( .A(n1260), .Y(n859) );
  INVX1_HVT U586 ( .A(n1293), .Y(n847) );
  INVX1_HVT U587 ( .A(keyin[66]), .Y(n868) );
  INVX1_HVT U588 ( .A(n1256), .Y(n857) );
  INVX1_HVT U589 ( .A(keyin[101]), .Y(n1374) );
  INVX1_HVT U590 ( .A(n827), .Y(n604) );
  INVX1_HVT U591 ( .A(keyin[111]), .Y(n601) );
  XNOR2X2_HVT U592 ( .A1(keyin[52]), .A2(keyin[84]), .Y(n600) );
  INVX1_HVT U593 ( .A(n1173), .Y(n824) );
  INVX0_HVT U594 ( .A(n1201), .Y(n1655) );
  INVX0_HVT U595 ( .A(n1199), .Y(n828) );
  INVX1_HVT U596 ( .A(n1195), .Y(n603) );
  INVX1_HVT U597 ( .A(keyin[127]), .Y(n827) );
  MUX41X1_HVT U598 ( .A1(n60), .A3(n56), .A2(n70), .A4(n66), .S0(n1196), .S1(
        n601), .Y(dummy[7]) );
  XOR3X2_HVT U599 ( .A1(keyin[7]), .A2(n1332), .A3(dummy[7]), .Y(keyout[7]) );
  XNOR2X1_HVT U600 ( .A1(n1300), .A2(n1289), .Y(keyout[72]) );
  XOR3X2_HVT U601 ( .A1(n1162), .A2(n868), .A3(n1259), .Y(keyout[98]) );
  XOR3X2_HVT U602 ( .A1(keyin[70]), .A2(n23), .A3(n1303), .Y(keyout[70]) );
  INVX1_HVT U603 ( .A(n1303), .Y(n1385) );
  XNOR2X2_HVT U604 ( .A1(n1291), .A2(keyin[38]), .Y(n1303) );
  MUX41X1_HVT U605 ( .A1(n98), .A3(n109), .A2(n104), .A4(n113), .S0(n601), 
        .S1(n603), .Y(dummy[5]) );
  XOR3X2_HVT U606 ( .A1(n1287), .A2(n845), .A3(n1331), .Y(keyout[106]) );
  XOR3X2_HVT U607 ( .A1(keyin[71]), .A2(n562), .A3(n1302), .Y(keyout[103]) );
  INVX2_HVT U608 ( .A(keyin[96]), .Y(n1380) );
  XNOR2X2_HVT U609 ( .A1(n1294), .A2(n1262), .Y(keyout[1]) );
  XOR3X2_HVT U610 ( .A1(keyin[67]), .A2(n1257), .A3(n1256), .Y(keyout[67]) );
  XOR3X2_HVT U611 ( .A1(n1289), .A2(n599), .A3(n1300), .Y(keyout[104]) );
  XNOR2X2_HVT U612 ( .A1(n1660), .A2(keyin[39]), .Y(n1302) );
  XOR2X2_HVT U613 ( .A1(keyin[33]), .A2(keyout[1]), .Y(keyout[33]) );
  XOR2X2_HVT U614 ( .A1(keyin[54]), .A2(keyout[22]), .Y(keyout[54]) );
  INVX2_HVT U615 ( .A(n1324), .Y(keyout[17]) );
  XOR2X2_HVT U616 ( .A1(keyin[48]), .A2(keyout[16]), .Y(keyout[48]) );
  XOR2X2_HVT U617 ( .A1(keyin[51]), .A2(keyout[19]), .Y(keyout[51]) );
  MUX41X1_HVT U618 ( .A1(n1598), .A3(n1205), .A2(n882), .A4(n1030), .S0(n556), 
        .S1(n1381), .Y(n1074) );
  XOR2X2_HVT U619 ( .A1(dummy[6]), .A2(keyin[6]), .Y(n605) );
  XOR2X2_HVT U620 ( .A1(keyout[17]), .A2(n1280), .Y(keyout[81]) );
  XNOR2X2_HVT U621 ( .A1(n1295), .A2(n1264), .Y(keyout[0]) );
  XOR2X1_HVT U622 ( .A1(n1298), .A2(n1527), .Y(keyout[4]) );
  XOR2X2_HVT U623 ( .A1(keyin[71]), .A2(keyout[39]), .Y(keyout[71]) );
  XOR3X2_HVT U624 ( .A1(keyin[68]), .A2(n828), .A3(n606), .Y(keyout[100]) );
  IBUFFX2_HVT U625 ( .A(n1254), .Y(n607) );
  MUX41X1_HVT U626 ( .A1(n633), .A3(n610), .A2(n659), .A4(n933), .S0(n556), 
        .S1(n1381), .Y(n609) );
  NAND2X0_HVT U627 ( .A1(n942), .A2(n991), .Y(n659) );
  XNOR2X2_HVT U628 ( .A1(keyin[27]), .A2(dummy[27]), .Y(n1314) );
  XOR2X2_HVT U629 ( .A1(keyout[25]), .A2(n1272), .Y(keyout[89]) );
  XOR2X2_HVT U630 ( .A1(keyout[21]), .A2(n1276), .Y(keyout[85]) );
  MUX21X1_HVT U634 ( .A1(n732), .A2(n1401), .S0(n1247), .Y(n733) );
  XOR3X2_HVT U635 ( .A1(n1264), .A2(n1379), .A3(n1265), .Y(keyout[96]) );
  XNOR2X2_HVT U636 ( .A1(keyin[26]), .A2(dummy[26]), .Y(n1315) );
  OA21X2_HVT U637 ( .A1(n1429), .A2(n1247), .A3(n1413), .Y(n725) );
  MUX21X1_HVT U638 ( .A1(n669), .A2(n667), .S0(n1246), .Y(n670) );
  MUX21X1_HVT U639 ( .A1(n722), .A2(n720), .S0(n1246), .Y(n723) );
  XNOR3X2_HVT U640 ( .A1(n1268), .A2(n251), .A3(n1312), .Y(keyout[125]) );
  NAND2X0_HVT U642 ( .A1(keyin[52]), .A2(n1321), .Y(n823) );
  NAND2X0_HVT U644 ( .A1(n822), .A2(n823), .Y(keyout[52]) );
  MUX41X1_HVT U645 ( .A1(n426), .A3(n434), .A2(n440), .A4(n445), .S0(n598), 
        .S1(n597), .Y(dummy[12]) );
  MUX21X1_HVT U646 ( .A1(n1194), .A2(n1192), .S0(n1360), .Y(n119) );
  INVX1_HVT U648 ( .A(n120), .Y(n842) );
  INVX0_HVT U649 ( .A(n830), .Y(n121) );
  MUX21X1_HVT U650 ( .A1(n427), .A2(n1469), .S0(n1344), .Y(n428) );
  MUX41X1_HVT U652 ( .A1(n425), .A3(n419), .A2(n423), .A4(n420), .S0(n1126), 
        .S1(n1133), .Y(n426) );
  MUX21X1_HVT U653 ( .A1(n1185), .A2(n1183), .S0(n1247), .Y(n729) );
  MUX21X1_HVT U654 ( .A1(n729), .A2(n1216), .S0(n848), .Y(n730) );
  XOR2X1_HVT U655 ( .A1(n1360), .A2(n1356), .Y(n829) );
  MUX41X1_HVT U656 ( .A1(n846), .A3(n844), .A2(n843), .A4(n842), .S0(n845), 
        .S1(n599), .Y(n830) );
  OAI21X1_HVT U657 ( .A1(n1559), .A2(n1360), .A3(n1543), .Y(n846) );
  XOR3X2_HVT U658 ( .A1(keyin[68]), .A2(n847), .A3(n1292), .Y(keyout[68]) );
  XNOR2X2_HVT U661 ( .A1(dummy[25]), .A2(keyin[25]), .Y(n1316) );
  XNOR2X2_HVT U662 ( .A1(dummy[4]), .A2(keyin[4]), .Y(n1292) );
  MUX21X2_HVT U663 ( .A1(n1233), .A2(n119), .S0(n870), .Y(n120) );
  MUX21X1_HVT U664 ( .A1(n1188), .A2(n824), .S0(n1344), .Y(n424) );
  XOR2X1_HVT U666 ( .A1(n1247), .A2(n1244), .Y(n848) );
  XOR2X2_HVT U667 ( .A1(dummy[20]), .A2(n849), .Y(n1321) );
  NAND2X0_HVT U668 ( .A1(n1224), .A2(n850), .Y(n851) );
  NAND2X0_HVT U669 ( .A1(n424), .A2(n853), .Y(n852) );
  NAND2X0_HVT U670 ( .A1(n851), .A2(n852), .Y(n425) );
  INVX0_HVT U671 ( .A(n853), .Y(n850) );
  XNOR2X1_HVT U672 ( .A1(n1342), .A2(n1255), .Y(n853) );
  XOR2X1_HVT U673 ( .A1(n1374), .A2(n1381), .Y(n963) );
  MUX41X1_HVT U674 ( .A1(n1024), .A3(n1019), .A2(n1026), .A4(n1023), .S0(
        keyin[103]), .S1(n545), .Y(n1027) );
  XOR2X2_HVT U675 ( .A1(keyout[29]), .A2(n1268), .Y(keyout[93]) );
  XOR2X2_HVT U677 ( .A1(keyin[60]), .A2(keyout[28]), .Y(keyout[60]) );
  XNOR2X2_HVT U679 ( .A1(keyin[29]), .A2(dummy[29]), .Y(n1312) );
  XNOR2X2_HVT U680 ( .A1(dummy[28]), .A2(keyin[28]), .Y(n1313) );
  MUX21X2_HVT U684 ( .A1(n1033), .A2(n1207), .S0(n965), .Y(n1034) );
  XOR2X2_HVT U689 ( .A1(keyout[27]), .A2(n1270), .Y(keyout[91]) );
  MUX21X2_HVT U690 ( .A1(n882), .A2(n1018), .S0(n963), .Y(n1019) );
  MUX21X1_HVT U692 ( .A1(n1215), .A2(n703), .S0(n896), .Y(n704) );
  IBUFFX2_HVT U696 ( .A(n1364), .Y(n854) );
  IBUFFX2_HVT U698 ( .A(n1254), .Y(n1252) );
  IBUFFX2_HVT U699 ( .A(n1254), .Y(n1251) );
  XOR2X2_HVT U700 ( .A1(n856), .A2(n1331), .Y(keyout[42]) );
  XOR2X2_HVT U702 ( .A1(keyout[18]), .A2(n1279), .Y(keyout[82]) );
  XOR2X2_HVT U705 ( .A1(keyout[13]), .A2(n1284), .Y(keyout[77]) );
  XOR2X2_HVT U713 ( .A1(n1304), .A2(n861), .Y(keyout[37]) );
  AO21X2_HVT U714 ( .A1(n287), .A2(n1520), .A3(n538), .Y(n407) );
  OA21X2_HVT U715 ( .A1(n901), .A2(n538), .A3(n335), .Y(n480) );
  OA21X2_HVT U716 ( .A1(n1471), .A2(n538), .A3(n335), .Y(n457) );
  XOR3X2_HVT U717 ( .A1(n857), .A2(n1258), .A3(n1257), .Y(keyout[99]) );
  XNOR2X2_HVT U718 ( .A1(n859), .A2(n869), .Y(keyout[34]) );
  XNOR2X2_HVT U721 ( .A1(n858), .A2(n869), .Y(keyout[2]) );
  MUX41X1_HVT U722 ( .A1(n708), .A3(n719), .A2(n714), .A4(n723), .S0(n827), 
        .S1(n860), .Y(dummy[21]) );
  INVX1_HVT U725 ( .A(n1296), .Y(n861) );
  NAND2X0_HVT U726 ( .A1(n778), .A2(n912), .Y(n864) );
  NAND2X0_HVT U727 ( .A1(n863), .A2(n864), .Y(n780) );
  IBUFFX2_HVT U729 ( .A(n912), .Y(n862) );
  MUX21X1_HVT U731 ( .A1(n777), .A2(n1216), .S0(n896), .Y(n778) );
  XOR2X2_HVT U733 ( .A1(keyin[5]), .A2(dummy[5]), .Y(n865) );
  NAND2X0_HVT U734 ( .A1(n473), .A2(n1131), .Y(n867) );
  MUX21X2_HVT U735 ( .A1(n167), .A2(n1233), .S0(n897), .Y(n168) );
  XOR2X2_HVT U736 ( .A1(dummy[2]), .A2(keyin[2]), .Y(n869) );
  MUX41X1_HVT U738 ( .A1(n170), .A3(n176), .A2(n172), .A4(n178), .S0(n603), 
        .S1(n1360), .Y(n179) );
  MUX21X1_HVT U739 ( .A1(n1232), .A2(n93), .S0(n897), .Y(n94) );
  XNOR3X2_HVT U740 ( .A1(keyin[69]), .A2(n1382), .A3(n865), .Y(keyout[69]) );
  MUX21X2_HVT U742 ( .A1(n776), .A2(n789), .S0(n827), .Y(dummy[18]) );
  MUX21X2_HVT U743 ( .A1(n169), .A2(n168), .S0(n1153), .Y(n170) );
  MUX21X2_HVT U745 ( .A1(n179), .A2(n166), .S0(keyin[111]), .Y(dummy[2]) );
  XNOR2X2_HVT U747 ( .A1(n1260), .A2(n1261), .Y(n1259) );
  INVX1_HVT U750 ( .A(keyin[124]), .Y(n1456) );
  MUX21X2_HVT U751 ( .A1(n700), .A2(n692), .S0(n604), .Y(dummy[22]) );
  INVX0_HVT U752 ( .A(keyin[126]), .Y(n1245) );
  IBUFFX2_HVT U753 ( .A(n1356), .Y(n1352) );
  INVX1_HVT U754 ( .A(keyin[116]), .Y(n1523) );
  INVX0_HVT U755 ( .A(n1364), .Y(n1363) );
  INVX0_HVT U756 ( .A(keyin[118]), .Y(n1341) );
  MUX21X2_HVT U757 ( .A1(n55), .A2(n51), .S0(n271), .Y(n56) );
  MUX21X2_HVT U758 ( .A1(n112), .A2(n110), .S0(n1359), .Y(n113) );
  INVX0_HVT U759 ( .A(n1356), .Y(n1355) );
  XNOR2X2_HVT U761 ( .A1(keyin[5]), .A2(dummy[5]), .Y(n1296) );
  XOR3X2_HVT U762 ( .A1(keyin[7]), .A2(n1332), .A3(dummy[7]), .Y(n1660) );
  INVX1_HVT U767 ( .A(n923), .Y(n1654) );
  INVX1_HVT U768 ( .A(n7), .Y(n1585) );
  INVX1_HVT U771 ( .A(n312), .Y(n1522) );
  INVX1_HVT U773 ( .A(n617), .Y(n1455) );
  NBUFFX2_HVT U776 ( .A(n923), .Y(n1208) );
  NBUFFX2_HVT U778 ( .A(n923), .Y(n1209) );
  AND2X1_HVT U780 ( .A1(n1238), .A2(n117), .Y(n871) );
  MUX21X1_HVT U781 ( .A1(n875), .A2(n1491), .S0(n1132), .Y(n405) );
  MUX21X1_HVT U783 ( .A1(n876), .A2(n1423), .S0(n913), .Y(n710) );
  MUX21X1_HVT U788 ( .A1(n627), .A2(n876), .S0(n915), .Y(n709) );
  AND2X1_HVT U789 ( .A1(n1521), .A2(n367), .Y(n872) );
  AND2X1_HVT U790 ( .A1(n1454), .A2(n672), .Y(n873) );
  AND2X1_HVT U794 ( .A1(n1176), .A2(n62), .Y(n874) );
  AND2X1_HVT U796 ( .A1(n1229), .A2(n422), .Y(n875) );
  AND2X1_HVT U800 ( .A1(n1220), .A2(n727), .Y(n876) );
  AND2X1_HVT U804 ( .A1(n1224), .A2(n379), .Y(n877) );
  AND2X1_HVT U807 ( .A1(n1216), .A2(n684), .Y(n878) );
  MUX21X1_HVT U809 ( .A1(n871), .A2(n1553), .S0(n1154), .Y(n100) );
  MUX21X1_HVT U813 ( .A1(n17), .A2(n871), .S0(n1155), .Y(n99) );
  AND2X1_HVT U815 ( .A1(n1233), .A2(n74), .Y(n879) );
  MUX21X1_HVT U818 ( .A1(n1623), .A2(n1055), .S0(n1157), .Y(n1056) );
  MUX21X1_HVT U819 ( .A1(n1648), .A2(n1211), .S0(n1165), .Y(n1055) );
  MUX21X1_HVT U823 ( .A1(n1609), .A2(n1653), .S0(keyin[98]), .Y(n985) );
  AND2X1_HVT U825 ( .A1(n974), .A2(n1179), .Y(n880) );
  NBUFFX2_HVT U827 ( .A(n7), .Y(n1230) );
  AND2X1_HVT U829 ( .A1(n1206), .A2(n991), .Y(n881) );
  AND2X1_HVT U833 ( .A1(n1213), .A2(n1031), .Y(n882) );
  NBUFFX2_HVT U834 ( .A(n1584), .Y(n1175) );
  NBUFFX2_HVT U835 ( .A(n312), .Y(n1221) );
  NBUFFX2_HVT U836 ( .A(n1658), .Y(n1179) );
  NBUFFX2_HVT U839 ( .A(n1658), .Y(n1178) );
  NBUFFX2_HVT U840 ( .A(n7), .Y(n1231) );
  NBUFFX2_HVT U843 ( .A(n1521), .Y(n1170) );
  NBUFFX2_HVT U846 ( .A(n1454), .Y(n1167) );
  NBUFFX2_HVT U848 ( .A(n1584), .Y(n1174) );
  NBUFFX2_HVT U849 ( .A(n1521), .Y(n1171) );
  NBUFFX2_HVT U850 ( .A(n1454), .Y(n1168) );
  NBUFFX2_HVT U851 ( .A(n1584), .Y(n1176) );
  INVX1_HVT U852 ( .A(n1235), .Y(n1583) );
  INVX1_HVT U853 ( .A(n1226), .Y(n1520) );
  INVX1_HVT U854 ( .A(n612), .Y(n1453) );
  INVX1_HVT U855 ( .A(n1210), .Y(n1653) );
  INVX1_HVT U856 ( .A(n1228), .Y(n1524) );
  INVX1_HVT U857 ( .A(n611), .Y(n1457) );
  INVX1_HVT U858 ( .A(n1), .Y(n1587) );
  NAND2X0_HVT U859 ( .A1(n1180), .A2(n1655), .Y(n923) );
  NBUFFX2_HVT U860 ( .A(n617), .Y(n1214) );
  NBUFFX2_HVT U861 ( .A(n312), .Y(n1222) );
  INVX1_HVT U862 ( .A(n1212), .Y(n1656) );
  MUX21X1_HVT U863 ( .A1(n1170), .A2(n1499), .S0(n266), .Y(n474) );
  MUX21X1_HVT U864 ( .A1(n1167), .A2(n1432), .S0(n913), .Y(n779) );
  MUX21X1_HVT U865 ( .A1(n310), .A2(n396), .S0(n1132), .Y(n397) );
  MUX21X1_HVT U866 ( .A1(n657), .A2(n1441), .S0(n915), .Y(n705) );
  MUX21X1_HVT U867 ( .A1(n615), .A2(n701), .S0(n913), .Y(n702) );
  MUX21X1_HVT U868 ( .A1(n1174), .A2(n1562), .S0(n1154), .Y(n169) );
  MUX21X1_HVT U869 ( .A1(n53), .A2(n52), .S0(n1155), .Y(n55) );
  MUX21X1_HVT U870 ( .A1(n447), .A2(n1493), .S0(n1131), .Y(n448) );
  MUX21X1_HVT U871 ( .A1(n1516), .A2(n345), .S0(n1349), .Y(n447) );
  MUX21X1_HVT U872 ( .A1(n752), .A2(n1425), .S0(n912), .Y(n753) );
  MUX21X1_HVT U873 ( .A1(n1449), .A2(n650), .S0(n608), .Y(n752) );
  MUX21X1_HVT U874 ( .A1(n47), .A2(n1571), .S0(n1155), .Y(n95) );
  MUX21X1_HVT U875 ( .A1(n5), .A2(n91), .S0(n1154), .Y(n92) );
  MUX21X1_HVT U876 ( .A1(n65), .A2(n63), .S0(n1359), .Y(n66) );
  MUX21X1_HVT U877 ( .A1(n675), .A2(n673), .S0(n1246), .Y(n676) );
  MUX21X1_HVT U878 ( .A1(n360), .A2(n356), .S0(n1342), .Y(n361) );
  MUX21X1_HVT U879 ( .A1(n358), .A2(n357), .S0(n1133), .Y(n360) );
  MUX21X1_HVT U880 ( .A1(n665), .A2(n661), .S0(n1246), .Y(n666) );
  MUX21X1_HVT U881 ( .A1(n663), .A2(n662), .S0(n914), .Y(n665) );
  MUX21X1_HVT U882 ( .A1(n142), .A2(n1555), .S0(n1153), .Y(n143) );
  MUX21X1_HVT U883 ( .A1(n1579), .A2(n40), .S0(n1361), .Y(n142) );
  MUX21X1_HVT U884 ( .A1(n370), .A2(n368), .S0(n1342), .Y(n371) );
  MUX21X1_HVT U885 ( .A1(n133), .A2(n132), .S0(n1154), .Y(n134) );
  MUX21X1_HVT U886 ( .A1(n417), .A2(n415), .S0(n1343), .Y(n418) );
  XOR2X1_HVT U887 ( .A1(n1239), .A2(n1453), .Y(n656) );
  XOR2X1_HVT U888 ( .A1(n1255), .A2(n1520), .Y(n351) );
  XOR2X1_HVT U889 ( .A1(n1353), .A2(n1583), .Y(n46) );
  MUX21X1_HVT U890 ( .A1(n1624), .A2(n930), .S0(n1159), .Y(n1018) );
  MUX21X1_HVT U891 ( .A1(n1526), .A2(n1173), .S0(n1277), .Y(n427) );
  MUX21X1_HVT U892 ( .A1(n1459), .A2(n1169), .S0(n1239), .Y(n732) );
  MUX21X1_HVT U893 ( .A1(n1653), .A2(n1657), .S0(n1365), .Y(n1085) );
  MUX21X1_HVT U894 ( .A1(n1654), .A2(n1657), .S0(n1365), .Y(n1094) );
  MUX21X1_HVT U895 ( .A1(n1656), .A2(n1179), .S0(n1366), .Y(n1082) );
  MUX21X1_HVT U896 ( .A1(n1655), .A2(n1213), .S0(n282), .Y(n1107) );
  MUX21X1_HVT U897 ( .A1(n1212), .A2(n1206), .S0(n1368), .Y(n1106) );
  MUX21X1_HVT U898 ( .A1(n942), .A2(n1181), .S0(n1368), .Y(n994) );
  MUX21X1_HVT U899 ( .A1(n1589), .A2(n1177), .S0(n537), .Y(n122) );
  XOR2X1_HVT U900 ( .A1(n1205), .A2(n1369), .Y(n966) );
  MUX21X1_HVT U901 ( .A1(n1655), .A2(n1181), .S0(n1369), .Y(n1110) );
  MUX21X1_HVT U902 ( .A1(n336), .A2(n521), .S0(n1132), .Y(n531) );
  MUX21X1_HVT U903 ( .A1(n641), .A2(n826), .S0(n913), .Y(n836) );
  MUX21X1_HVT U904 ( .A1(n1228), .A2(n1225), .S0(n268), .Y(n496) );
  MUX21X1_HVT U905 ( .A1(n611), .A2(n1217), .S0(n213), .Y(n801) );
  MUX21X1_HVT U906 ( .A1(n1496), .A2(n309), .S0(n1342), .Y(n419) );
  MUX21X1_HVT U907 ( .A1(n1428), .A2(n614), .S0(n1246), .Y(n724) );
  MUX21X1_HVT U908 ( .A1(n687), .A2(n688), .S0(n912), .Y(n690) );
  MUX21X1_HVT U909 ( .A1(n1418), .A2(n627), .S0(n914), .Y(n687) );
  XOR2X1_HVT U910 ( .A1(n1215), .A2(n1242), .Y(n660) );
  XOR2X1_HVT U911 ( .A1(n1223), .A2(n1255), .Y(n355) );
  XOR2X1_HVT U912 ( .A1(n1232), .A2(n253), .Y(n50) );
  MUX21X1_HVT U913 ( .A1(n1520), .A2(n1525), .S0(n268), .Y(n468) );
  MUX21X1_HVT U914 ( .A1(n1524), .A2(n1171), .S0(n268), .Y(n466) );
  MUX21X1_HVT U915 ( .A1(n1453), .A2(n1458), .S0(n213), .Y(n773) );
  MUX21X1_HVT U916 ( .A1(n1457), .A2(n1168), .S0(n213), .Y(n771) );
  MUX21X1_HVT U917 ( .A1(n1), .A2(n1234), .S0(n525), .Y(n191) );
  MUX21X1_HVT U918 ( .A1(n1173), .A2(n1229), .S0(n267), .Y(n498) );
  MUX21X1_HVT U919 ( .A1(n1169), .A2(n1220), .S0(n1239), .Y(n803) );
  MUX21X1_HVT U920 ( .A1(n1179), .A2(n828), .S0(n1368), .Y(n932) );
  MUX21X1_HVT U921 ( .A1(n1177), .A2(n1587), .S0(n1354), .Y(n11) );
  MUX21X1_HVT U922 ( .A1(n1233), .A2(n1177), .S0(n1353), .Y(n14) );
  MUX21X1_HVT U923 ( .A1(n77), .A2(n78), .S0(n1153), .Y(n80) );
  MUX21X1_HVT U924 ( .A1(n997), .A2(n998), .S0(n1160), .Y(n1000) );
  MUX21X1_HVT U925 ( .A1(n936), .A2(n1211), .S0(n1165), .Y(n997) );
  MUX21X1_HVT U926 ( .A1(n335), .A2(n421), .S0(n1342), .Y(n423) );
  MUX21X1_HVT U927 ( .A1(n640), .A2(n726), .S0(n1246), .Y(n728) );
  MUX21X1_HVT U928 ( .A1(n884), .A2(n411), .S0(n266), .Y(n412) );
  MUX21X1_HVT U929 ( .A1(n323), .A2(n410), .S0(n1131), .Y(n411) );
  MUX21X1_HVT U930 ( .A1(n1171), .A2(n1522), .S0(n1277), .Y(n410) );
  MUX21X1_HVT U931 ( .A1(n1168), .A2(n1455), .S0(n1239), .Y(n715) );
  MUX21X1_HVT U932 ( .A1(n1583), .A2(n1588), .S0(n537), .Y(n163) );
  MUX21X1_HVT U933 ( .A1(n1587), .A2(n1175), .S0(n525), .Y(n161) );
  MUX21X1_HVT U934 ( .A1(n1177), .A2(n1238), .S0(n537), .Y(n193) );
  MUX21X1_HVT U935 ( .A1(n31), .A2(n216), .S0(n1154), .Y(n226) );
  MUX21X1_HVT U936 ( .A1(n1232), .A2(n1589), .S0(n525), .Y(n221) );
  AND2X1_HVT U937 ( .A1(n1355), .A2(n1588), .Y(n883) );
  AND2X1_HVT U938 ( .A1(n1339), .A2(n1525), .Y(n884) );
  AND2X1_HVT U939 ( .A1(n1241), .A2(n1458), .Y(n885) );
  MUX21X1_HVT U940 ( .A1(n1657), .A2(n1656), .S0(n1369), .Y(n943) );
  MUX21X1_HVT U941 ( .A1(n1212), .A2(n1211), .S0(n1366), .Y(n947) );
  MUX21X1_HVT U946 ( .A1(n1656), .A2(n1654), .S0(n282), .Y(n953) );
  MUX21X1_HVT U947 ( .A1(n1175), .A2(n1177), .S0(n253), .Y(n19) );
  MUX21X1_HVT U948 ( .A1(n1207), .A2(n1211), .S0(n282), .Y(n930) );
  MUX21X1_HVT U949 ( .A1(n1234), .A2(n1236), .S0(n252), .Y(n17) );
  MUX21X1_HVT U950 ( .A1(n1656), .A2(n828), .S0(n1368), .Y(n950) );
  MUX21X1_HVT U951 ( .A1(n1209), .A2(n1213), .S0(n1368), .Y(n1012) );
  MUX21X1_HVT U953 ( .A1(n828), .A2(n1657), .S0(n1369), .Y(n956) );
  MUX21X1_HVT U955 ( .A1(n1181), .A2(n1654), .S0(n282), .Y(n945) );
  MUX21X1_HVT U956 ( .A1(n1221), .A2(n313), .S0(n1338), .Y(n342) );
  MUX21X1_HVT U957 ( .A1(n1214), .A2(n618), .S0(n1243), .Y(n647) );
  MUX21X1_HVT U958 ( .A1(n1231), .A2(n1177), .S0(n1355), .Y(n12) );
  MUX21X1_HVT U959 ( .A1(n1558), .A2(n4), .S0(n1358), .Y(n114) );
  MUX21X1_HVT U961 ( .A1(n340), .A2(n341), .S0(n1133), .Y(n453) );
  MUX21X1_HVT U962 ( .A1(n616), .A2(n758), .S0(n912), .Y(n759) );
  MUX21X1_HVT U964 ( .A1(n645), .A2(n646), .S0(n914), .Y(n758) );
  MUX21X1_HVT U965 ( .A1(n1540), .A2(n1583), .S0(n1152), .Y(n69) );
  MUX21X1_HVT U966 ( .A1(n1114), .A2(n1115), .S0(n1159), .Y(n1116) );
  MUX21X1_HVT U967 ( .A1(n1607), .A2(n1651), .S0(n1165), .Y(n1114) );
  MUX21X1_HVT U968 ( .A1(n1227), .A2(n1173), .S0(n1277), .Y(n528) );
  MUX21X1_HVT U969 ( .A1(n1218), .A2(n1169), .S0(n1242), .Y(n833) );
  MUX21X1_HVT U970 ( .A1(n1039), .A2(n1038), .S0(n1165), .Y(n1040) );
  MUX21X1_HVT U972 ( .A1(n1598), .A2(n1626), .S0(n1157), .Y(n1038) );
  MUX21X1_HVT U973 ( .A1(n1059), .A2(n922), .S0(n1158), .Y(n1060) );
  MUX21X1_HVT U974 ( .A1(n939), .A2(n1630), .S0(n1166), .Y(n1059) );
  MUX21X1_HVT U975 ( .A1(n1043), .A2(n1044), .S0(n1166), .Y(n1047) );
  MUX21X1_HVT U976 ( .A1(n1601), .A2(n1042), .S0(n1160), .Y(n1043) );
  MUX21X1_HVT U978 ( .A1(n917), .A2(n1213), .S0(n1159), .Y(n1045) );
  MUX21X1_HVT U979 ( .A1(n883), .A2(n106), .S0(n1154), .Y(n107) );
  MUX21X1_HVT U980 ( .A1(n18), .A2(n105), .S0(n1153), .Y(n106) );
  MUX21X1_HVT U981 ( .A1(n1175), .A2(n1585), .S0(n525), .Y(n105) );
  MUX21X1_HVT U982 ( .A1(n1180), .A2(n828), .S0(n1365), .Y(n1042) );
  XOR2X1_HVT U983 ( .A1(n1367), .A2(n1653), .Y(n961) );
  MUX21X1_HVT U984 ( .A1(n1208), .A2(n1211), .S0(n1368), .Y(n1007) );
  MUX21X1_HVT U985 ( .A1(n1211), .A2(n828), .S0(n1367), .Y(n1137) );
  MUX21X1_HVT U986 ( .A1(n1654), .A2(n1180), .S0(n281), .Y(n1141) );
  MUX21X1_HVT U987 ( .A1(n828), .A2(n942), .S0(n1369), .Y(n1139) );
  MUX21X1_HVT U988 ( .A1(n946), .A2(n1129), .S0(n1164), .Y(n1140) );
  MUX21X1_HVT U989 ( .A1(n1583), .A2(n1585), .S0(n1353), .Y(n13) );
  MUX21X1_HVT U991 ( .A1(n1525), .A2(n1524), .S0(n268), .Y(n332) );
  MUX21X1_HVT U993 ( .A1(n1458), .A2(n1457), .S0(n213), .Y(n637) );
  MUX21X1_HVT U994 ( .A1(n1228), .A2(n1227), .S0(n1333), .Y(n335) );
  MUX21X1_HVT U999 ( .A1(n1220), .A2(n1218), .S0(n212), .Y(n640) );
  MUX21X1_HVT U1003 ( .A1(n1457), .A2(n1455), .S0(n213), .Y(n649) );
  MUX21X1_HVT U1004 ( .A1(n1587), .A2(n1585), .S0(n1353), .Y(n39) );
  MUX21X1_HVT U1006 ( .A1(n1225), .A2(n1227), .S0(n1277), .Y(n322) );
  MUX21X1_HVT U1009 ( .A1(n1217), .A2(n1218), .S0(n212), .Y(n627) );
  MUX21X1_HVT U1010 ( .A1(n1524), .A2(n1173), .S0(n1338), .Y(n338) );
  MUX21X1_HVT U1011 ( .A1(n1457), .A2(n1169), .S0(n1239), .Y(n643) );
  MUX21X1_HVT U1015 ( .A1(n1587), .A2(n1177), .S0(n524), .Y(n33) );
  MUX21X1_HVT U1017 ( .A1(n942), .A2(n1657), .S0(n1368), .Y(n941) );
  MUX21X1_HVT U1018 ( .A1(n1223), .A2(n1171), .S0(n1333), .Y(n347) );
  MUX21X1_HVT U1020 ( .A1(n1215), .A2(n1168), .S0(n1243), .Y(n652) );
  MUX21X1_HVT U1027 ( .A1(n1207), .A2(n1179), .S0(n1366), .Y(n957) );
  MUX21X1_HVT U1028 ( .A1(n1206), .A2(n828), .S0(n1365), .Y(n935) );
  MUX21X1_HVT U1030 ( .A1(n1224), .A2(n1173), .S0(n268), .Y(n319) );
  MUX21X1_HVT U1031 ( .A1(n1216), .A2(n1169), .S0(n212), .Y(n624) );
  MUX21X1_HVT U1033 ( .A1(n1208), .A2(n828), .S0(n281), .Y(n927) );
  MUX21X1_HVT U1034 ( .A1(n1209), .A2(n942), .S0(n1367), .Y(n952) );
  MUX21X1_HVT U1038 ( .A1(n1173), .A2(n1525), .S0(n267), .Y(n346) );
  MUX21X1_HVT U1039 ( .A1(n1169), .A2(n1458), .S0(n1240), .Y(n651) );
  MUX21X1_HVT U1041 ( .A1(n1230), .A2(n247), .S0(n1354), .Y(n37) );
  MUX21X1_HVT U1043 ( .A1(n1222), .A2(n1173), .S0(n267), .Y(n317) );
  MUX21X1_HVT U1045 ( .A1(n1214), .A2(n1169), .S0(n1242), .Y(n622) );
  MUX21X1_HVT U1046 ( .A1(n1178), .A2(n1181), .S0(n1367), .Y(n1022) );
  MUX21X1_HVT U1047 ( .A1(n1620), .A2(n946), .S0(n1157), .Y(n1050) );
  MUX21X1_HVT U1050 ( .A1(n977), .A2(n975), .S0(n1159), .Y(n978) );
  MUX21X1_HVT U1051 ( .A1(n6), .A2(n148), .S0(n1153), .Y(n149) );
  MUX21X1_HVT U1052 ( .A1(n35), .A2(n36), .S0(n1154), .Y(n148) );
  MUX21X1_HVT U1055 ( .A1(n30), .A2(n116), .S0(n1358), .Y(n118) );
  MUX21X1_HVT U1056 ( .A1(n1222), .A2(n1227), .S0(n1277), .Y(n396) );
  MUX21X1_HVT U1058 ( .A1(n1214), .A2(n1219), .S0(n1242), .Y(n701) );
  MUX21X1_HVT U1059 ( .A1(n1468), .A2(n1495), .S0(n1342), .Y(n437) );
  MUX21X1_HVT U1060 ( .A1(n1400), .A2(n1427), .S0(n1246), .Y(n742) );
  MUX21X1_HVT U1061 ( .A1(n1522), .A2(n1525), .S0(n1277), .Y(n487) );
  MUX21X1_HVT U1063 ( .A1(n1455), .A2(n1458), .S0(n1241), .Y(n792) );
  MUX21X1_HVT U1065 ( .A1(n1211), .A2(n1180), .S0(n1366), .Y(n989) );
  MUX21X1_HVT U1066 ( .A1(n1456), .A2(n1459), .S0(n1241), .Y(n806) );
  MUX21X1_HVT U1068 ( .A1(n1172), .A2(n1526), .S0(n1338), .Y(n501) );
  MUX21X1_HVT U1069 ( .A1(n1586), .A2(n1589), .S0(n524), .Y(n196) );
  MUX21X1_HVT U1072 ( .A1(n1179), .A2(n1654), .S0(n281), .Y(n1014) );
  MUX21X1_HVT U1073 ( .A1(n618), .A2(n1459), .S0(n1240), .Y(n693) );
  MUX21X1_HVT U1076 ( .A1(n313), .A2(n1526), .S0(n1333), .Y(n388) );
  MUX21X1_HVT U1077 ( .A1(n1236), .A2(n1177), .S0(n524), .Y(n223) );
  MUX21X1_HVT U1080 ( .A1(n942), .A2(n1653), .S0(n281), .Y(n1142) );
  MUX21X1_HVT U1082 ( .A1(n1205), .A2(n1180), .S0(n282), .Y(n1135) );
  MUX21X1_HVT U1084 ( .A1(n313), .A2(n1520), .S0(n268), .Y(n533) );
  MUX21X1_HVT U1088 ( .A1(n618), .A2(n1453), .S0(n1240), .Y(n838) );
  MUX21X1_HVT U1089 ( .A1(n1653), .A2(n1654), .S0(n1369), .Y(n934) );
  MUX21X1_HVT U1091 ( .A1(n1588), .A2(n1587), .S0(n252), .Y(n27) );
  MUX21X1_HVT U1092 ( .A1(n1), .A2(n1236), .S0(n537), .Y(n30) );
  MUX21X1_HVT U1094 ( .A1(n1171), .A2(n1173), .S0(n1333), .Y(n324) );
  MUX21X1_HVT U1095 ( .A1(n1168), .A2(n1169), .S0(n212), .Y(n629) );
  MUX21X1_HVT U1096 ( .A1(n1526), .A2(n1522), .S0(n267), .Y(n334) );
  MUX21X1_HVT U1099 ( .A1(n1459), .A2(n1455), .S0(n1243), .Y(n639) );
  MUX21X1_HVT U1100 ( .A1(n313), .A2(n1525), .S0(n267), .Y(n330) );
  MUX21X1_HVT U1101 ( .A1(n618), .A2(n1458), .S0(n1239), .Y(n635) );
  MUX21X1_HVT U1102 ( .A1(n1232), .A2(n1175), .S0(n525), .Y(n42) );
  MUX21X1_HVT U1103 ( .A1(n1173), .A2(n1524), .S0(n268), .Y(n316) );
  MUX21X1_HVT U1108 ( .A1(n1169), .A2(n1457), .S0(n1241), .Y(n621) );
  MUX21X1_HVT U1110 ( .A1(n1176), .A2(n1587), .S0(n253), .Y(n9) );
  MUX21X1_HVT U1111 ( .A1(n1170), .A2(n1524), .S0(n1338), .Y(n314) );
  MUX21X1_HVT U1112 ( .A1(n1167), .A2(n1457), .S0(n212), .Y(n619) );
  MUX21X1_HVT U1114 ( .A1(n1170), .A2(n1526), .S0(n1333), .Y(n408) );
  MUX21X1_HVT U1122 ( .A1(n1167), .A2(n1459), .S0(n1241), .Y(n713) );
  MUX21X1_HVT U1124 ( .A1(n1174), .A2(n1589), .S0(n537), .Y(n103) );
  MUX21X1_HVT U1126 ( .A1(n1453), .A2(n1455), .S0(n212), .Y(n623) );
  MUX21X1_HVT U1127 ( .A1(n1421), .A2(n641), .S0(n1246), .Y(n746) );
  MUX21X1_HVT U1129 ( .A1(n1478), .A2(n1520), .S0(n1130), .Y(n374) );
  MUX21X1_HVT U1130 ( .A1(n1410), .A2(n1453), .S0(n911), .Y(n679) );
  MUX21X1_HVT U1131 ( .A1(n891), .A2(n1484), .S0(n1342), .Y(n443) );
  MUX21X1_HVT U1135 ( .A1(n892), .A2(n1416), .S0(n1246), .Y(n748) );
  MUX21X1_HVT U1137 ( .A1(n325), .A2(n1494), .S0(n1342), .Y(n444) );
  MUX21X1_HVT U1138 ( .A1(n1223), .A2(n1526), .S0(n1338), .Y(n526) );
  MUX21X1_HVT U1139 ( .A1(n7), .A2(n1237), .S0(n252), .Y(n91) );
  MUX21X1_HVT U1141 ( .A1(n1456), .A2(n618), .S0(n1242), .Y(n835) );
  MUX21X1_HVT U1145 ( .A1(n1227), .A2(n1170), .S0(n268), .Y(n416) );
  MUX21X1_HVT U1146 ( .A1(n1218), .A2(n1167), .S0(n1243), .Y(n721) );
  MUX21X1_HVT U1148 ( .A1(n1585), .A2(n1587), .S0(n1152), .Y(n54) );
  MUX21X1_HVT U1149 ( .A1(n1585), .A2(n1588), .S0(n1354), .Y(n182) );
  MUX21X1_HVT U1151 ( .A1(n247), .A2(n1589), .S0(n524), .Y(n83) );
  XOR2X1_HVT U1155 ( .A1(n1148), .A2(n1352), .Y(n43) );
  MUX21X1_HVT U1157 ( .A1(n1172), .A2(n313), .S0(n268), .Y(n530) );
  MUX21X1_HVT U1158 ( .A1(n247), .A2(n1583), .S0(n537), .Y(n228) );
  MUX21X1_HVT U1160 ( .A1(n1215), .A2(n1459), .S0(n1240), .Y(n831) );
  MUX21X1_HVT U1161 ( .A1(n1520), .A2(n1522), .S0(n1277), .Y(n318) );
  MUX21X1_HVT U1162 ( .A1(n1589), .A2(n1585), .S0(n1355), .Y(n29) );
  MUX21X1_HVT U1163 ( .A1(n247), .A2(n1588), .S0(n1354), .Y(n25) );
  MUX21X1_HVT U1164 ( .A1(n1177), .A2(n1588), .S0(n253), .Y(n41) );
  MUX21X1_HVT U1165 ( .A1(n1236), .A2(n1176), .S0(n524), .Y(n111) );
  XOR2X1_HVT U1166 ( .A1(n942), .A2(n1365), .Y(n962) );
  XOR2X1_HVT U1167 ( .A1(n313), .A2(n1255), .Y(n352) );
  XOR2X1_HVT U1168 ( .A1(n1180), .A2(n1367), .Y(n960) );
  MUX21X1_HVT U1169 ( .A1(n1586), .A2(n247), .S0(n537), .Y(n225) );
  MUX21X1_HVT U1170 ( .A1(n1221), .A2(n1229), .S0(n1255), .Y(n402) );
  MUX21X1_HVT U1171 ( .A1(n1214), .A2(n1220), .S0(n1242), .Y(n707) );
  MUX21X1_HVT U1172 ( .A1(n1522), .A2(n1526), .S0(n1255), .Y(n532) );
  MUX21X1_HVT U1173 ( .A1(n893), .A2(n1546), .S0(n272), .Y(n138) );
  MUX21X1_HVT U1174 ( .A1(n20), .A2(n1556), .S0(n271), .Y(n139) );
  MUX21X1_HVT U1175 ( .A1(n1522), .A2(n1524), .S0(n1130), .Y(n359) );
  MUX21X1_HVT U1176 ( .A1(n1455), .A2(n1457), .S0(n911), .Y(n664) );
  XOR2X1_HVT U1177 ( .A1(n8), .A2(n1354), .Y(n47) );
  XNOR2X1_HVT U1178 ( .A1(n1228), .A2(n1255), .Y(n886) );
  XNOR2X1_HVT U1179 ( .A1(n611), .A2(n1242), .Y(n887) );
  MUX21X1_HVT U1180 ( .A1(n1654), .A2(n1656), .S0(keyin[98]), .Y(n970) );
  XOR2X1_HVT U1181 ( .A1(n281), .A2(n1163), .Y(n958) );
  MUX21X1_HVT U1182 ( .A1(n1455), .A2(n1459), .S0(n213), .Y(n837) );
  MUX21X1_HVT U1183 ( .A1(n1223), .A2(n1222), .S0(n1255), .Y(n534) );
  MUX21X1_HVT U1184 ( .A1(n1215), .A2(n1214), .S0(n1240), .Y(n839) );
  MUX21X1_HVT U1185 ( .A1(n1205), .A2(n1208), .S0(n281), .Y(n1143) );
  XNOR2X1_HVT U1186 ( .A1(n1208), .A2(n1368), .Y(n888) );
  XNOR2X1_HVT U1187 ( .A1(n1212), .A2(n282), .Y(n889) );
  XNOR2X1_HVT U1188 ( .A1(n1), .A2(n1353), .Y(n890) );
  MUX21X1_HVT U1189 ( .A1(n1231), .A2(n1238), .S0(n1353), .Y(n97) );
  MUX21X1_HVT U1190 ( .A1(n828), .A2(n1656), .S0(n281), .Y(n926) );
  MUX21X1_HVT U1191 ( .A1(n1178), .A2(n1656), .S0(n1365), .Y(n924) );
  NBUFFX2_HVT U1192 ( .A(n3), .Y(n1233) );
  XNOR2X1_HVT U1193 ( .A1(n1222), .A2(n1255), .Y(n891) );
  XNOR2X1_HVT U1194 ( .A1(n1214), .A2(n1243), .Y(n892) );
  XOR2X1_HVT U1195 ( .A1(n1083), .A2(n1255), .Y(n348) );
  XOR2X1_HVT U1196 ( .A1(n907), .A2(n1240), .Y(n653) );
  NAND2X0_HVT U1197 ( .A1(n1177), .A2(n1589), .Y(n7) );
  XNOR2X1_HVT U1198 ( .A1(n1231), .A2(n253), .Y(n893) );
  MUX21X1_HVT U1199 ( .A1(n1585), .A2(n1589), .S0(n1352), .Y(n227) );
  MUX21X1_HVT U1200 ( .A1(n1232), .A2(n1231), .S0(n1353), .Y(n229) );
  NBUFFX2_HVT U1201 ( .A(n308), .Y(n1224) );
  NBUFFX2_HVT U1202 ( .A(n613), .Y(n1216) );
  NBUFFX2_HVT U1203 ( .A(n3), .Y(n1234) );
  NAND2X0_HVT U1204 ( .A1(n1172), .A2(n1526), .Y(n312) );
  NAND2X0_HVT U1205 ( .A1(n1169), .A2(n1459), .Y(n617) );
  AND2X1_HVT U1206 ( .A1(n1657), .A2(n1369), .Y(n894) );
  NBUFFX2_HVT U1207 ( .A(n308), .Y(n1223) );
  NBUFFX2_HVT U1208 ( .A(n613), .Y(n1215) );
  NBUFFX2_HVT U1209 ( .A(n3), .Y(n1232) );
  INVX0_HVT U1210 ( .A(n313), .Y(n1521) );
  INVX0_HVT U1211 ( .A(n618), .Y(n1454) );
  NBUFFX2_HVT U1212 ( .A(n2), .Y(n1235) );
  NBUFFX2_HVT U1213 ( .A(n1523), .Y(n1172) );
  NBUFFX2_HVT U1214 ( .A(n308), .Y(n1225) );
  NBUFFX2_HVT U1215 ( .A(n613), .Y(n1217) );
  NBUFFX2_HVT U1216 ( .A(n306), .Y(n1228) );
  NBUFFX2_HVT U1217 ( .A(n307), .Y(n1226) );
  NBUFFX2_HVT U1218 ( .A(n917), .Y(n1210) );
  NBUFFX2_HVT U1219 ( .A(n2), .Y(n1236) );
  NBUFFX2_HVT U1220 ( .A(n919), .Y(n1205) );
  NBUFFX2_HVT U1221 ( .A(n916), .Y(n1212) );
  NBUFFX2_HVT U1222 ( .A(n1659), .Y(n1181) );
  NBUFFX2_HVT U1223 ( .A(n919), .Y(n1206) );
  NBUFFX2_HVT U1224 ( .A(n919), .Y(n1207) );
  NBUFFX2_HVT U1225 ( .A(n917), .Y(n1211) );
  NBUFFX2_HVT U1226 ( .A(n2), .Y(n1237) );
  NBUFFX2_HVT U1227 ( .A(n1378), .Y(n1166) );
  MUX21X1_HVT U1228 ( .A1(n1227), .A2(n1229), .S0(n1342), .Y(n430) );
  MUX21X1_HVT U1229 ( .A1(n1219), .A2(n1220), .S0(n1246), .Y(n735) );
  NBUFFX2_HVT U1230 ( .A(n307), .Y(n1227) );
  NBUFFX2_HVT U1231 ( .A(n612), .Y(n1218) );
  NBUFFX2_HVT U1232 ( .A(n612), .Y(n1219) );
  NBUFFX2_HVT U1233 ( .A(n611), .Y(n1220) );
  NBUFFX2_HVT U1234 ( .A(n306), .Y(n1229) );
  NBUFFX2_HVT U1235 ( .A(n1), .Y(n1238) );
  NBUFFX2_HVT U1236 ( .A(n1378), .Y(n1165) );
  NBUFFX2_HVT U1237 ( .A(n1378), .Y(n1164) );
  NBUFFX2_HVT U1238 ( .A(n916), .Y(n1213) );
  NBUFFX2_HVT U1239 ( .A(n1253), .Y(n915) );
  NBUFFX2_HVT U1240 ( .A(n1586), .Y(n1177) );
  MUX21X1_HVT U1241 ( .A1(n1237), .A2(n1238), .S0(n1358), .Y(n125) );
  NBUFFX2_HVT U1242 ( .A(keyin[104]), .Y(n1155) );
  NBUFFX2_HVT U1243 ( .A(n1253), .Y(n914) );
  NBUFFX2_HVT U1244 ( .A(n1349), .Y(n1132) );
  NBUFFX2_HVT U1245 ( .A(n1253), .Y(n913) );
  NBUFFX2_HVT U1246 ( .A(keyin[104]), .Y(n1154) );
  NBUFFX2_HVT U1247 ( .A(n1523), .Y(n1173) );
  NBUFFX2_HVT U1248 ( .A(n1456), .Y(n1169) );
  NBUFFX2_HVT U1249 ( .A(n1659), .Y(n1180) );
  NBUFFX2_HVT U1250 ( .A(n1375), .Y(n1163) );
  NBUFFX2_HVT U1251 ( .A(keyin[101]), .Y(n1157) );
  NBUFFX2_HVT U1252 ( .A(keyin[101]), .Y(n1160) );
  NBUFFX2_HVT U1253 ( .A(keyin[101]), .Y(n1159) );
  NBUFFX2_HVT U1254 ( .A(keyin[101]), .Y(n1158) );
  NBUFFX2_HVT U1255 ( .A(n1375), .Y(n1162) );
  NBUFFX2_HVT U1256 ( .A(n1163), .Y(n1161) );
  NBUFFX2_HVT U1257 ( .A(keyin[101]), .Y(n1156) );
  MUX21X1_HVT U1258 ( .A1(n1182), .A2(n1459), .S0(n915), .Y(n703) );
  XNOR2X1_HVT U1259 ( .A1(n1244), .A2(n1253), .Y(n896) );
  XNOR2X1_HVT U1260 ( .A1(n1356), .A2(n854), .Y(n897) );
  MUX21X1_HVT U1261 ( .A1(n1191), .A2(n1589), .S0(n1155), .Y(n93) );
  MUX21X1_HVT U1262 ( .A1(n456), .A2(n457), .S0(n1131), .Y(n458) );
  MUX21X1_HVT U1263 ( .A1(n379), .A2(n352), .S0(n1349), .Y(n456) );
  MUX21X1_HVT U1264 ( .A1(n462), .A2(n463), .S0(n1130), .Y(n465) );
  MUX21X1_HVT U1265 ( .A1(n421), .A2(n1225), .S0(n1349), .Y(n462) );
  MUX21X1_HVT U1266 ( .A1(n767), .A2(n768), .S0(n911), .Y(n770) );
  MUX21X1_HVT U1267 ( .A1(n726), .A2(n1217), .S0(n1253), .Y(n767) );
  MUX21X1_HVT U1268 ( .A1(n151), .A2(n152), .S0(n1153), .Y(n153) );
  MUX21X1_HVT U1269 ( .A1(n74), .A2(n47), .S0(n855), .Y(n151) );
  MUX21X1_HVT U1270 ( .A1(n157), .A2(n158), .S0(n1152), .Y(n160) );
  MUX21X1_HVT U1271 ( .A1(n116), .A2(n1234), .S0(n854), .Y(n157) );
  XOR2X1_HVT U1272 ( .A1(n1296), .A2(n1297), .Y(keyout[5]) );
  XOR2X1_HVT U1273 ( .A1(n1301), .A2(n1257), .Y(keyout[3]) );
  XOR2X1_HVT U1274 ( .A1(n1303), .A2(n605), .Y(keyout[38]) );
  XNOR2X1_HVT U1275 ( .A1(n1263), .A2(n1262), .Y(keyout[65]) );
  XOR2X1_HVT U1276 ( .A1(n1290), .A2(n1291), .Y(keyout[6]) );
  MUX21X1_HVT U1277 ( .A1(n1200), .A2(n1203), .S0(n1160), .Y(n1033) );
  MUX21X1_HVT U1278 ( .A1(n1627), .A2(n918), .S0(n1160), .Y(n1028) );
  MUX21X1_HVT U1279 ( .A1(n947), .A2(n1030), .S0(n1157), .Y(n1032) );
  MUX21X1_HVT U1280 ( .A1(n969), .A2(n968), .S0(n1164), .Y(n971) );
  MUX21X1_HVT U1281 ( .A1(n1200), .A2(n920), .S0(n1375), .Y(n968) );
  MUX21X1_HVT U1282 ( .A1(n888), .A2(n1613), .S0(n1160), .Y(n1052) );
  MUX21X1_HVT U1283 ( .A1(n933), .A2(n1625), .S0(n1158), .Y(n1053) );
  MUX21X1_HVT U1284 ( .A1(n1203), .A2(n1207), .S0(n1365), .Y(n936) );
  MUX21X1_HVT U1285 ( .A1(n1119), .A2(n1118), .S0(n1159), .Y(n1120) );
  MUX21X1_HVT U1286 ( .A1(n307), .A2(n478), .S0(n1134), .Y(n479) );
  MUX21X1_HVT U1287 ( .A1(n785), .A2(n784), .S0(n911), .Y(n786) );
  MUX21X1_HVT U1288 ( .A1(n1219), .A2(n783), .S0(n915), .Y(n784) );
  MUX21X1_HVT U1289 ( .A1(n685), .A2(n655), .S0(n911), .Y(n686) );
  XOR2X1_HVT U1290 ( .A1(n1254), .A2(n637), .Y(n655) );
  MUX21X1_HVT U1291 ( .A1(n682), .A2(n683), .S0(n914), .Y(n685) );
  MUX21X1_HVT U1292 ( .A1(n1219), .A2(n1459), .S0(n1241), .Y(n682) );
  MUX21X1_HVT U1293 ( .A1(n380), .A2(n350), .S0(n1130), .Y(n381) );
  XOR2X1_HVT U1294 ( .A1(n538), .A2(n332), .Y(n350) );
  MUX21X1_HVT U1295 ( .A1(n377), .A2(n378), .S0(n1133), .Y(n380) );
  MUX21X1_HVT U1296 ( .A1(n1227), .A2(n1526), .S0(n1338), .Y(n377) );
  MUX21X1_HVT U1297 ( .A1(n309), .A2(n286), .S0(n1342), .Y(n431) );
  MUX21X1_HVT U1298 ( .A1(n1230), .A2(n1192), .S0(n252), .Y(n10) );
  MUX21X1_HVT U1299 ( .A1(n1194), .A2(n1583), .S0(n253), .Y(n20) );
  MUX21X1_HVT U1300 ( .A1(n1178), .A2(n1201), .S0(n281), .Y(n939) );
  MUX21X1_HVT U1301 ( .A1(n1188), .A2(n1524), .S0(n1338), .Y(n341) );
  MUX21X1_HVT U1302 ( .A1(n1185), .A2(n1457), .S0(n213), .Y(n646) );
  MUX21X1_HVT U1303 ( .A1(n828), .A2(n1203), .S0(n281), .Y(n946) );
  MUX21X1_HVT U1304 ( .A1(n1201), .A2(n1654), .S0(n1367), .Y(n954) );
  MUX21X1_HVT U1305 ( .A1(n1654), .A2(n1203), .S0(n1367), .Y(n948) );
  MUX21X1_HVT U1306 ( .A1(n1194), .A2(n1234), .S0(n1355), .Y(n21) );
  MUX21X1_HVT U1307 ( .A1(n1020), .A2(n1623), .S0(n1158), .Y(n1023) );
  MUX21X1_HVT U1308 ( .A1(n1011), .A2(n1010), .S0(n1160), .Y(n1013) );
  MUX21X1_HVT U1309 ( .A1(n1205), .A2(n1009), .S0(n898), .Y(n1010) );
  MUX21X1_HVT U1310 ( .A1(n1201), .A2(n1180), .S0(n1166), .Y(n1009) );
  MUX21X1_HVT U1311 ( .A1(n1071), .A2(n1070), .S0(n1156), .Y(n1073) );
  MUX21X1_HVT U1312 ( .A1(n1645), .A2(n1653), .S0(n1166), .Y(n1070) );
  MUX21X1_HVT U1313 ( .A1(n175), .A2(n174), .S0(n1152), .Y(n176) );
  MUX21X1_HVT U1314 ( .A1(n1237), .A2(n173), .S0(n1155), .Y(n174) );
  MUX21X1_HVT U1315 ( .A1(n1103), .A2(n1102), .S0(n1160), .Y(n1104) );
  MUX21X1_HVT U1316 ( .A1(n1004), .A2(n1200), .S0(n1165), .Y(n1102) );
  MUX21X1_HVT U1318 ( .A1(n959), .A2(n987), .S0(n1159), .Y(n988) );
  MUX21X1_HVT U1319 ( .A1(n1656), .A2(n1643), .S0(n1166), .Y(n987) );
  XOR2X1_HVT U1320 ( .A1(n1380), .A2(n943), .Y(n959) );
  MUX21X1_HVT U1321 ( .A1(n1542), .A2(n1357), .S0(n1152), .Y(n67) );
  MUX21X1_HVT U1322 ( .A1(n1090), .A2(n1091), .S0(n1156), .Y(n1092) );
  MUX21X1_HVT U1323 ( .A1(n917), .A2(n1643), .S0(n1166), .Y(n1090) );
  MUX21X1_HVT U1325 ( .A1(n1065), .A2(n1066), .S0(n1158), .Y(n1067) );
  MUX21X1_HVT U1327 ( .A1(n945), .A2(n1604), .S0(n1165), .Y(n1065) );
  MUX21X1_HVT U1328 ( .A1(n1077), .A2(n1076), .S0(n1160), .Y(n1078) );
  MUX21X1_HVT U1329 ( .A1(n1075), .A2(n1207), .S0(n898), .Y(n1076) );
  MUX21X1_HVT U1330 ( .A1(n953), .A2(n1646), .S0(n1165), .Y(n1077) );
  MUX21X1_HVT U1331 ( .A1(n75), .A2(n45), .S0(n1152), .Y(n76) );
  XOR2X1_HVT U1332 ( .A1(n1364), .A2(n27), .Y(n45) );
  MUX21X1_HVT U1333 ( .A1(n72), .A2(n73), .S0(n1154), .Y(n75) );
  MUX21X1_HVT U1334 ( .A1(n1237), .A2(n1589), .S0(n1352), .Y(n72) );
  MUX21X1_HVT U1335 ( .A1(n1192), .A2(n34), .S0(n1153), .Y(n52) );
  MUX21X1_HVT U1336 ( .A1(n4), .A2(n1357), .S0(n1358), .Y(n126) );
  MUX21X1_HVT U1337 ( .A1(n1203), .A2(n1211), .S0(n1365), .Y(n1144) );
  MUX21X1_HVT U1338 ( .A1(n1194), .A2(n247), .S0(n525), .Y(n222) );
  INVX1_HVT U1339 ( .A(n1340), .Y(n1333) );
  INVX1_HVT U1340 ( .A(n1340), .Y(n1277) );
  NBUFFX2_HVT U1341 ( .A(keyin[106]), .Y(n1153) );
  MUX21X1_HVT U1342 ( .A1(n1203), .A2(n1656), .S0(n282), .Y(n951) );
  MUX21X1_HVT U1344 ( .A1(n1209), .A2(n1200), .S0(n281), .Y(n925) );
  MUX21X1_HVT U1346 ( .A1(n1203), .A2(n1653), .S0(n1369), .Y(n933) );
  MUX21X1_HVT U1348 ( .A1(n1194), .A2(n1587), .S0(n252), .Y(n36) );
  MUX21X1_HVT U1349 ( .A1(n1188), .A2(n1225), .S0(n267), .Y(n326) );
  MUX21X1_HVT U1350 ( .A1(n1185), .A2(n1217), .S0(n1239), .Y(n631) );
  MUX21X1_HVT U1352 ( .A1(n1186), .A2(n1522), .S0(n1333), .Y(n343) );
  MUX21X1_HVT U1354 ( .A1(n1182), .A2(n1455), .S0(n213), .Y(n648) );
  MUX21X1_HVT U1356 ( .A1(n1191), .A2(n1585), .S0(n1352), .Y(n38) );
  MUX21X1_HVT U1358 ( .A1(n1213), .A2(n1203), .S0(n1366), .Y(n944) );
  MUX21X1_HVT U1360 ( .A1(n1498), .A2(n1221), .S0(n1133), .Y(n490) );
  MUX21X1_HVT U1361 ( .A1(n796), .A2(n795), .S0(n912), .Y(n797) );
  MUX21X1_HVT U1362 ( .A1(n1430), .A2(n617), .S0(n914), .Y(n795) );
  MUX21X1_HVT U1363 ( .A1(n186), .A2(n185), .S0(n1153), .Y(n187) );
  MUX21X1_HVT U1364 ( .A1(n1560), .A2(n1230), .S0(n1155), .Y(n185) );
  MUX21X1_HVT U1366 ( .A1(n1611), .A2(n1370), .S0(keyin[98]), .Y(n983) );
  MUX21X1_HVT U1368 ( .A1(n810), .A2(n811), .S0(n912), .Y(n812) );
  MUX21X1_HVT U1370 ( .A1(n646), .A2(n622), .S0(n915), .Y(n810) );
  MUX21X1_HVT U1372 ( .A1(n200), .A2(n201), .S0(n1153), .Y(n202) );
  MUX21X1_HVT U1374 ( .A1(n36), .A2(n12), .S0(n1155), .Y(n200) );
  XOR2X1_HVT U1375 ( .A1(n1199), .A2(n282), .Y(n964) );
  MUX21X1_HVT U1376 ( .A1(n1211), .A2(n1178), .S0(n1367), .Y(n1025) );
  MUX21X1_HVT U1377 ( .A1(n1188), .A2(n1227), .S0(n1338), .Y(n535) );
  MUX21X1_HVT U1378 ( .A1(n1185), .A2(n1219), .S0(n213), .Y(n840) );
  MUX21X1_HVT U1379 ( .A1(n1194), .A2(n1237), .S0(n524), .Y(n230) );
  MUX21X1_HVT U1380 ( .A1(n1201), .A2(n1653), .S0(n1369), .Y(n1138) );
  MUX21X1_HVT U1381 ( .A1(n1186), .A2(n1520), .S0(n267), .Y(n529) );
  MUX21X1_HVT U1382 ( .A1(n1182), .A2(n1453), .S0(n1241), .Y(n834) );
  MUX21X1_HVT U1383 ( .A1(n1203), .A2(n942), .S0(n1366), .Y(n1136) );
  INVX1_HVT U1384 ( .A(n1340), .Y(n1338) );
  MUX21X1_HVT U1385 ( .A1(n1170), .A2(n1186), .S0(n1277), .Y(n329) );
  MUX21X1_HVT U1386 ( .A1(n1167), .A2(n1182), .S0(n1239), .Y(n634) );
  MUX21X1_HVT U1388 ( .A1(n1176), .A2(n1191), .S0(n252), .Y(n24) );
  MUX21X1_HVT U1389 ( .A1(n1221), .A2(n824), .S0(n1333), .Y(n315) );
  MUX21X1_HVT U1390 ( .A1(n617), .A2(n1183), .S0(n1243), .Y(n620) );
  MUX21X1_HVT U1391 ( .A1(n1188), .A2(n1520), .S0(n1333), .Y(n325) );
  MUX21X1_HVT U1392 ( .A1(n1185), .A2(n1453), .S0(n1243), .Y(n630) );
  MUX21X1_HVT U1393 ( .A1(n1173), .A2(n1188), .S0(n1338), .Y(n336) );
  MUX21X1_HVT U1394 ( .A1(n1169), .A2(n1185), .S0(n212), .Y(n641) );
  MUX21X1_HVT U1395 ( .A1(n1522), .A2(n1188), .S0(n1333), .Y(n337) );
  MUX21X1_HVT U1396 ( .A1(n1455), .A2(n1185), .S0(n212), .Y(n642) );
  MUX21X1_HVT U1397 ( .A1(n1585), .A2(n1194), .S0(n252), .Y(n32) );
  MUX21X1_HVT U1398 ( .A1(n1229), .A2(n1188), .S0(n267), .Y(n333) );
  MUX21X1_HVT U1399 ( .A1(n1220), .A2(n1185), .S0(n1241), .Y(n638) );
  MUX21X1_HVT U1400 ( .A1(n1238), .A2(n1194), .S0(n1352), .Y(n28) );
  MUX21X1_HVT U1401 ( .A1(n1480), .A2(n286), .S0(n1130), .Y(n372) );
  MUX21X1_HVT U1402 ( .A1(n1412), .A2(n1245), .S0(n911), .Y(n677) );
  XNOR2X1_HVT U1403 ( .A1(n1380), .A2(n1368), .Y(n898) );
  MUX21X1_HVT U1404 ( .A1(n1188), .A2(n313), .S0(n1277), .Y(n527) );
  MUX21X1_HVT U1405 ( .A1(n1185), .A2(n618), .S0(n1240), .Y(n832) );
  INVX1_HVT U1406 ( .A(n1370), .Y(n1365) );
  NBUFFX2_HVT U1407 ( .A(keyin[106]), .Y(n1152) );
  MUX21X1_HVT U1408 ( .A1(n1177), .A2(n1194), .S0(n1352), .Y(n31) );
  MUX21X1_HVT U1409 ( .A1(n824), .A2(n339), .S0(n1131), .Y(n357) );
  MUX21X1_HVT U1410 ( .A1(n1183), .A2(n644), .S0(n912), .Y(n662) );
  MUX21X1_HVT U1411 ( .A1(n1191), .A2(n1583), .S0(n525), .Y(n224) );
  INVX1_HVT U1412 ( .A(n286), .Y(n1255) );
  NBUFFX2_HVT U1413 ( .A(keyin[114]), .Y(n1131) );
  NBUFFX2_HVT U1414 ( .A(n1250), .Y(n912) );
  MUX21X1_HVT U1415 ( .A1(n1188), .A2(n1229), .S0(n1255), .Y(n536) );
  MUX21X1_HVT U1416 ( .A1(n1185), .A2(n1220), .S0(n1240), .Y(n841) );
  MUX21X1_HVT U1417 ( .A1(n1194), .A2(n1238), .S0(n252), .Y(n231) );
  MUX21X1_HVT U1418 ( .A1(n1203), .A2(n1213), .S0(n1366), .Y(n1145) );
  INVX1_HVT U1419 ( .A(n1370), .Y(n1369) );
  INVX1_HVT U1420 ( .A(n1364), .Y(n1362) );
  NBUFFX2_HVT U1421 ( .A(keyin[114]), .Y(n1130) );
  NBUFFX2_HVT U1422 ( .A(n1250), .Y(n911) );
  MUX21X1_HVT U1423 ( .A1(n918), .A2(n1371), .S0(n1159), .Y(n1046) );
  XOR2X1_HVT U1424 ( .A1(n1186), .A2(n1255), .Y(n353) );
  XOR2X1_HVT U1425 ( .A1(n1183), .A2(n1239), .Y(n658) );
  NAND2X0_HVT U1426 ( .A1(n1589), .A2(n1192), .Y(n3) );
  INVX1_HVT U1427 ( .A(keyin[107]), .Y(n1589) );
  XOR2X1_HVT U1428 ( .A1(n1192), .A2(n253), .Y(n48) );
  INVX1_HVT U1429 ( .A(keyin[108]), .Y(n1586) );
  XOR2X1_HVT U1437 ( .A1(n1659), .A2(n1199), .Y(n942) );
  NAND2X0_HVT U1438 ( .A1(n1526), .A2(n1186), .Y(n308) );
  NAND2X0_HVT U1439 ( .A1(n1459), .A2(n1183), .Y(n613) );
  INVX1_HVT U1441 ( .A(keyin[115]), .Y(n1526) );
  INVX1_HVT U1442 ( .A(keyin[123]), .Y(n1459) );
  INVX1_HVT U1443 ( .A(n1202), .Y(n1659) );
  NBUFFX2_HVT U1445 ( .A(n1345), .Y(n1127) );
  NBUFFX2_HVT U1446 ( .A(n1250), .Y(n910) );
  NBUFFX2_HVT U1450 ( .A(n1147), .Y(n1151) );
  NAND2X0_HVT U1453 ( .A1(n1193), .A2(n1586), .Y(n2) );
  AND2X1_HVT U1456 ( .A1(n1176), .A2(n1357), .Y(n899) );
  NAND2X0_HVT U1457 ( .A1(n1187), .A2(n1186), .Y(n306) );
  NAND2X0_HVT U1458 ( .A1(n1184), .A2(n1182), .Y(n611) );
  NAND2X0_HVT U1459 ( .A1(n1193), .A2(n1191), .Y(n1) );
  NAND2X0_HVT U1460 ( .A1(n1187), .A2(n1172), .Y(n307) );
  NAND2X0_HVT U1463 ( .A1(n1184), .A2(n1456), .Y(n612) );
  NAND2X0_HVT U1467 ( .A1(n1655), .A2(n1202), .Y(n917) );
  AND2X1_HVT U1474 ( .A1(n1178), .A2(n1371), .Y(n900) );
  AND2X1_HVT U1475 ( .A1(n1521), .A2(n1341), .Y(n901) );
  AND2X1_HVT U1476 ( .A1(n1454), .A2(n1245), .Y(n902) );
  NAND2X0_HVT U1477 ( .A1(n1199), .A2(n1202), .Y(n916) );
  NAND2X0_HVT U1478 ( .A1(n1199), .A2(n1181), .Y(n919) );
  AND2X1_HVT U1479 ( .A1(n1357), .A2(n1177), .Y(n903) );
  XOR2X1_HVT U1480 ( .A1(n286), .A2(n1187), .Y(n349) );
  XOR2X1_HVT U1481 ( .A1(n1245), .A2(n1184), .Y(n654) );
  INVX1_HVT U1482 ( .A(n1381), .Y(n1379) );
  XOR2X1_HVT U1483 ( .A1(n1357), .A2(n1193), .Y(n44) );
  AND2X1_HVT U1484 ( .A1(n287), .A2(n1173), .Y(n904) );
  AND2X1_HVT U1485 ( .A1(n1245), .A2(n1169), .Y(n905) );
  NBUFFX2_HVT U1486 ( .A(keyin[106]), .Y(n1148) );
  AND2X1_HVT U1487 ( .A1(n828), .A2(n1371), .Y(n906) );
  NBUFFX2_HVT U1488 ( .A(keyin[106]), .Y(n1147) );
  NBUFFX2_HVT U1489 ( .A(n1346), .Y(n1083) );
  NBUFFX2_HVT U1490 ( .A(n1249), .Y(n907) );
  NBUFFX2_HVT U1491 ( .A(n1346), .Y(n1125) );
  NBUFFX2_HVT U1492 ( .A(n1249), .Y(n908) );
  NBUFFX2_HVT U1493 ( .A(keyin[98]), .Y(n1375) );
  NBUFFX2_HVT U1494 ( .A(n1346), .Y(n1126) );
  NBUFFX2_HVT U1495 ( .A(n1249), .Y(n909) );
  NBUFFX2_HVT U1496 ( .A(keyin[106]), .Y(n1149) );
  INVX1_HVT U1497 ( .A(n1374), .Y(n1372) );
  NBUFFX2_HVT U1498 ( .A(n1345), .Y(n938) );
  NBUFFX2_HVT U1499 ( .A(n1149), .Y(n1146) );
  NBUFFX2_HVT U1500 ( .A(keyin[106]), .Y(n1150) );
  INVX1_HVT U1501 ( .A(n1374), .Y(n1373) );
  MUX21X1_HVT U1502 ( .A1(n413), .A2(n412), .S0(n1343), .Y(n414) );
  XOR2X1_HVT U1503 ( .A1(keyin[69]), .A2(n1372), .Y(n1335) );
  MUX21X1_HVT U1504 ( .A1(n59), .A2(n57), .S0(n1359), .Y(n60) );
  MUX21X1_HVT U1505 ( .A1(n108), .A2(n107), .S0(n271), .Y(n109) );
  XNOR2X1_HVT U1506 ( .A1(keyin[67]), .A2(n1202), .Y(n1258) );
  MUX21X1_HVT U1507 ( .A1(n364), .A2(n362), .S0(n1343), .Y(n365) );
  MUX21X1_HVT U1508 ( .A1(n1048), .A2(n1047), .S0(keyin[98]), .Y(n1049) );
  MUX21X1_HVT U1509 ( .A1(n981), .A2(n979), .S0(n1159), .Y(n982) );
  XOR2X1_HVT U1510 ( .A1(n1298), .A2(keyin[36]), .Y(n1293) );
  XOR2X1_HVT U1511 ( .A1(n1301), .A2(keyin[35]), .Y(n1256) );
  XOR2X1_HVT U1512 ( .A1(n1308), .A2(keyin[34]), .Y(n1260) );
  XNOR2X1_HVT U1513 ( .A1(n1297), .A2(keyin[37]), .Y(n1304) );
  XOR3X1_HVT U1514 ( .A1(keyin[65]), .A2(keyin[33]), .A3(n1294), .Y(n1263) );
  NBUFFX2_HVT U1515 ( .A(keyin[122]), .Y(n1250) );
  NBUFFX2_HVT U1516 ( .A(keyin[107]), .Y(n1193) );
  NBUFFX2_HVT U1517 ( .A(keyin[99]), .Y(n1202) );
  NBUFFX2_HVT U1518 ( .A(keyin[100]), .Y(n1199) );
  NBUFFX2_HVT U1519 ( .A(keyin[115]), .Y(n1187) );
  NBUFFX2_HVT U1520 ( .A(keyin[123]), .Y(n1184) );
  NBUFFX2_HVT U1521 ( .A(keyin[124]), .Y(n1182) );
  NBUFFX2_HVT U1522 ( .A(keyin[116]), .Y(n1186) );
  NBUFFX2_HVT U1523 ( .A(keyin[108]), .Y(n1191) );
  NBUFFX2_HVT U1524 ( .A(keyin[100]), .Y(n1201) );
  INVX0_HVT U1525 ( .A(keyin[110]), .Y(n1357) );
  NBUFFX2_HVT U1526 ( .A(keyin[108]), .Y(n1192) );
  NBUFFX2_HVT U1527 ( .A(keyin[124]), .Y(n1183) );
  INVX0_HVT U1528 ( .A(keyin[102]), .Y(n1371) );
  NBUFFX2_HVT U1529 ( .A(keyin[107]), .Y(n1194) );
  NBUFFX2_HVT U1530 ( .A(keyin[99]), .Y(n1203) );
  NBUFFX2_HVT U1531 ( .A(keyin[100]), .Y(n1200) );
  NBUFFX2_HVT U1532 ( .A(keyin[123]), .Y(n1185) );
  NBUFFX2_HVT U1533 ( .A(keyin[115]), .Y(n1188) );
  NBUFFX2_HVT U1534 ( .A(keyin[114]), .Y(n1346) );
  NBUFFX2_HVT U1535 ( .A(keyin[122]), .Y(n1249) );
  NBUFFX2_HVT U1536 ( .A(keyin[114]), .Y(n1345) );
  NBUFFX2_HVT U1537 ( .A(keyin[122]), .Y(n1248) );
  NBUFFX2_HVT U1538 ( .A(keyin[105]), .Y(n1196) );
  NBUFFX2_HVT U1539 ( .A(keyin[103]), .Y(n1198) );
  NBUFFX2_HVT U1540 ( .A(keyin[113]), .Y(n1189) );
  NBUFFX2_HVT U1541 ( .A(keyin[113]), .Y(n1190) );
  NBUFFX2_HVT U1542 ( .A(keyin[105]), .Y(n1197) );
  NBUFFX2_HVT U1543 ( .A(keyin[105]), .Y(n1195) );
  NBUFFX2_HVT U1544 ( .A(keyin[97]), .Y(n1204) );
  XOR2X1_HVT U1545 ( .A1(keyin[55]), .A2(keyin[87]), .Y(n1274) );
  XOR2X1_HVT U1546 ( .A1(keyin[47]), .A2(keyin[79]), .Y(n1282) );
  XOR2X1_HVT U1547 ( .A1(keyin[41]), .A2(keyin[73]), .Y(n1288) );
  XOR2X1_HVT U1548 ( .A1(keyin[49]), .A2(keyin[81]), .Y(n1280) );
  XOR2X1_HVT U1549 ( .A1(keyin[42]), .A2(keyin[74]), .Y(n1287) );
  XOR2X1_HVT U1550 ( .A1(keyin[50]), .A2(keyin[82]), .Y(n1279) );
  XOR2X1_HVT U1551 ( .A1(keyin[63]), .A2(keyin[95]), .Y(n1266) );
  XOR2X1_HVT U1552 ( .A1(keyin[51]), .A2(keyin[83]), .Y(n1278) );
  XOR2X1_HVT U1553 ( .A1(keyin[43]), .A2(keyin[75]), .Y(n1286) );
  XOR2X1_HVT U1554 ( .A1(keyin[44]), .A2(keyin[76]), .Y(n1285) );
  XOR2X1_HVT U1555 ( .A1(keyin[57]), .A2(keyin[89]), .Y(n1272) );
  XOR2X1_HVT U1556 ( .A1(keyin[46]), .A2(keyin[78]), .Y(n1283) );
  XOR2X1_HVT U1557 ( .A1(keyin[54]), .A2(keyin[86]), .Y(n1275) );
  XOR2X1_HVT U1558 ( .A1(keyin[58]), .A2(keyin[90]), .Y(n1271) );
  XOR2X1_HVT U1559 ( .A1(keyin[45]), .A2(keyin[77]), .Y(n1284) );
  XOR2X1_HVT U1560 ( .A1(keyin[53]), .A2(keyin[85]), .Y(n1276) );
  XOR2X1_HVT U1561 ( .A1(keyin[60]), .A2(keyin[92]), .Y(n1269) );
  XOR2X1_HVT U1562 ( .A1(keyin[59]), .A2(keyin[91]), .Y(n1270) );
  XOR2X1_HVT U1563 ( .A1(keyin[40]), .A2(keyin[72]), .Y(n1289) );
  XOR2X1_HVT U1564 ( .A1(keyin[48]), .A2(keyin[80]), .Y(n1281) );
  XOR2X1_HVT U1565 ( .A1(keyin[62]), .A2(keyin[94]), .Y(n1267) );
  XOR2X1_HVT U1566 ( .A1(keyin[61]), .A2(keyin[93]), .Y(n1268) );
  XOR2X1_HVT U1567 ( .A1(keyin[56]), .A2(keyin[88]), .Y(n1273) );
  INVX0_HVT U1568 ( .A(n1304), .Y(n1382) );
  INVX0_HVT U1569 ( .A(round_num[0]), .Y(n1383) );
  INVX0_HVT U1570 ( .A(n1306), .Y(n1384) );
  INVX0_HVT U1571 ( .A(n1305), .Y(n1386) );
  INVX0_HVT U1572 ( .A(round_num[3]), .Y(n1387) );
  INVX0_HVT U1573 ( .A(n1302), .Y(keyout[39]) );
  INVX0_HVT U1574 ( .A(round_num[2]), .Y(n1389) );
  INVX0_HVT U1575 ( .A(round_num[1]), .Y(n1390) );
  INVX0_HVT U1576 ( .A(n632), .Y(n1398) );
  INVX0_HVT U1577 ( .A(n636), .Y(n1399) );
  INVX0_HVT U1578 ( .A(n644), .Y(n1400) );
  INVX0_HVT U1579 ( .A(n645), .Y(n1401) );
  INVX0_HVT U1580 ( .A(n654), .Y(n1402) );
  INVX0_HVT U1581 ( .A(n787), .Y(n1403) );
  INVX0_HVT U1582 ( .A(n825), .Y(n1404) );
  INVX0_HVT U1583 ( .A(n628), .Y(n1406) );
  INVX0_HVT U1584 ( .A(n616), .Y(n1407) );
  INVX0_HVT U1585 ( .A(n615), .Y(n1408) );
  INVX0_HVT U1586 ( .A(n619), .Y(n1409) );
  INVX0_HVT U1587 ( .A(n620), .Y(n1410) );
  INVX0_HVT U1588 ( .A(n621), .Y(n1411) );
  INVX0_HVT U1589 ( .A(n622), .Y(n1412) );
  INVX0_HVT U1590 ( .A(n623), .Y(n1413) );
  INVX0_HVT U1591 ( .A(n624), .Y(n1414) );
  INVX0_HVT U1592 ( .A(n627), .Y(n1415) );
  INVX0_HVT U1593 ( .A(n629), .Y(n1416) );
  INVX0_HVT U1594 ( .A(n630), .Y(n1417) );
  INVX0_HVT U1595 ( .A(n631), .Y(n1418) );
  INVX0_HVT U1596 ( .A(n635), .Y(n1420) );
  INVX0_HVT U1597 ( .A(n638), .Y(n1421) );
  INVX0_HVT U1598 ( .A(n639), .Y(n1422) );
  INVX0_HVT U1599 ( .A(n640), .Y(n1423) );
  INVX0_HVT U1600 ( .A(n641), .Y(n1424) );
  INVX0_HVT U1601 ( .A(n836), .Y(n1425) );
  INVX0_HVT U1602 ( .A(n642), .Y(n1426) );
  INVX0_HVT U1603 ( .A(n643), .Y(n1427) );
  INVX0_HVT U1604 ( .A(n646), .Y(n1428) );
  INVX0_HVT U1605 ( .A(n647), .Y(n1429) );
  INVX0_HVT U1606 ( .A(n648), .Y(n1430) );
  INVX0_HVT U1607 ( .A(n649), .Y(n1431) );
  INVX0_HVT U1608 ( .A(n650), .Y(n1432) );
  INVX0_HVT U1609 ( .A(n651), .Y(n1433) );
  INVX0_HVT U1610 ( .A(n652), .Y(n1434) );
  INVX0_HVT U1611 ( .A(n684), .Y(n1435) );
  INVX0_HVT U1612 ( .A(n625), .Y(n1436) );
  INVX0_HVT U1613 ( .A(n672), .Y(n1437) );
  INVX0_HVT U1614 ( .A(n727), .Y(n1438) );
  INVX0_HVT U1615 ( .A(n826), .Y(n1439) );
  INVX0_HVT U1616 ( .A(n769), .Y(n1440) );
  INVX0_HVT U1617 ( .A(n831), .Y(n1441) );
  INVX0_HVT U1618 ( .A(n832), .Y(n1442) );
  INVX0_HVT U1619 ( .A(n834), .Y(n1444) );
  INVX0_HVT U1620 ( .A(n835), .Y(n1445) );
  INVX0_HVT U1621 ( .A(n707), .Y(n1446) );
  INVX0_HVT U1622 ( .A(n713), .Y(n1447) );
  INVX0_HVT U1623 ( .A(n837), .Y(n1448) );
  INVX0_HVT U1624 ( .A(n838), .Y(n1449) );
  INVX0_HVT U1625 ( .A(n839), .Y(n1450) );
  INVX0_HVT U1626 ( .A(n840), .Y(n1451) );
  INVX0_HVT U1627 ( .A(n841), .Y(n1452) );
  INVX0_HVT U1628 ( .A(n1215), .Y(n1458) );
  INVX0_HVT U1629 ( .A(n1326), .Y(keyout[15]) );
  INVX0_HVT U1630 ( .A(n327), .Y(n1466) );
  INVX0_HVT U1631 ( .A(n331), .Y(n1467) );
  INVX0_HVT U1632 ( .A(n339), .Y(n1468) );
  INVX0_HVT U1633 ( .A(n340), .Y(n1469) );
  INVX0_HVT U1634 ( .A(n349), .Y(n1470) );
  INVX0_HVT U1635 ( .A(n482), .Y(n1471) );
  INVX0_HVT U1636 ( .A(n520), .Y(n1472) );
  INVX0_HVT U1637 ( .A(n309), .Y(n1473) );
  INVX0_HVT U1638 ( .A(n323), .Y(n1474) );
  INVX0_HVT U1639 ( .A(n311), .Y(n1475) );
  INVX0_HVT U1640 ( .A(n310), .Y(n1476) );
  INVX0_HVT U1641 ( .A(n314), .Y(n1477) );
  INVX0_HVT U1642 ( .A(n315), .Y(n1478) );
  INVX0_HVT U1643 ( .A(n316), .Y(n1479) );
  INVX0_HVT U1644 ( .A(n317), .Y(n1480) );
  INVX0_HVT U1645 ( .A(n318), .Y(n1481) );
  INVX0_HVT U1646 ( .A(n319), .Y(n1482) );
  INVX0_HVT U1647 ( .A(n322), .Y(n1483) );
  INVX0_HVT U1648 ( .A(n324), .Y(n1484) );
  INVX0_HVT U1649 ( .A(n325), .Y(n1485) );
  INVX0_HVT U1650 ( .A(n326), .Y(n1486) );
  INVX0_HVT U1651 ( .A(n329), .Y(n1487) );
  INVX0_HVT U1652 ( .A(n330), .Y(n1488) );
  INVX0_HVT U1653 ( .A(n333), .Y(n1489) );
  INVX0_HVT U1654 ( .A(n334), .Y(n1490) );
  INVX0_HVT U1655 ( .A(n335), .Y(n1491) );
  INVX0_HVT U1656 ( .A(n336), .Y(n1492) );
  INVX0_HVT U1657 ( .A(n337), .Y(n1494) );
  INVX0_HVT U1658 ( .A(n338), .Y(n1495) );
  INVX0_HVT U1659 ( .A(n341), .Y(n1496) );
  INVX0_HVT U1660 ( .A(n342), .Y(n1497) );
  INVX0_HVT U1661 ( .A(n343), .Y(n1498) );
  INVX0_HVT U1662 ( .A(n345), .Y(n1499) );
  INVX0_HVT U1663 ( .A(n346), .Y(n1500) );
  INVX0_HVT U1664 ( .A(n347), .Y(n1501) );
  INVX0_HVT U1665 ( .A(n379), .Y(n1502) );
  INVX0_HVT U1666 ( .A(n320), .Y(n1503) );
  INVX0_HVT U1667 ( .A(n367), .Y(n1504) );
  INVX0_HVT U1668 ( .A(n422), .Y(n1505) );
  INVX0_HVT U1669 ( .A(n521), .Y(n1506) );
  INVX0_HVT U1670 ( .A(n464), .Y(n1507) );
  INVX0_HVT U1671 ( .A(n526), .Y(n1508) );
  INVX0_HVT U1672 ( .A(n527), .Y(n1509) );
  INVX0_HVT U1673 ( .A(n528), .Y(n1510) );
  INVX0_HVT U1674 ( .A(n529), .Y(n1511) );
  INVX0_HVT U1675 ( .A(n530), .Y(n1512) );
  INVX0_HVT U1676 ( .A(n402), .Y(n1513) );
  INVX0_HVT U1677 ( .A(n408), .Y(n1514) );
  INVX0_HVT U1678 ( .A(n532), .Y(n1515) );
  INVX0_HVT U1679 ( .A(n533), .Y(n1516) );
  INVX0_HVT U1680 ( .A(n534), .Y(n1517) );
  INVX0_HVT U1681 ( .A(n535), .Y(n1518) );
  INVX0_HVT U1682 ( .A(n536), .Y(n1519) );
  INVX0_HVT U1683 ( .A(n1223), .Y(n1525) );
  INVX0_HVT U1684 ( .A(n1292), .Y(n1527) );
  INVX0_HVT U1685 ( .A(n22), .Y(n1528) );
  INVX0_HVT U1686 ( .A(n26), .Y(n1529) );
  INVX0_HVT U1687 ( .A(n34), .Y(n1530) );
  INVX0_HVT U1688 ( .A(n35), .Y(n1531) );
  INVX0_HVT U1689 ( .A(n44), .Y(n1532) );
  INVX0_HVT U1690 ( .A(n177), .Y(n1533) );
  INVX0_HVT U1691 ( .A(n215), .Y(n1534) );
  INVX0_HVT U1692 ( .A(n4), .Y(n1535) );
  INVX0_HVT U1693 ( .A(n18), .Y(n1536) );
  INVX0_HVT U1694 ( .A(n6), .Y(n1537) );
  INVX0_HVT U1695 ( .A(n5), .Y(n1538) );
  INVX0_HVT U1696 ( .A(n9), .Y(n1539) );
  INVX0_HVT U1697 ( .A(n10), .Y(n1540) );
  INVX0_HVT U1698 ( .A(n11), .Y(n1541) );
  INVX0_HVT U1699 ( .A(n12), .Y(n1542) );
  INVX0_HVT U1700 ( .A(n13), .Y(n1543) );
  INVX0_HVT U1701 ( .A(n14), .Y(n1544) );
  INVX0_HVT U1702 ( .A(n19), .Y(n1546) );
  INVX0_HVT U1703 ( .A(n20), .Y(n1547) );
  INVX0_HVT U1704 ( .A(n21), .Y(n1548) );
  INVX0_HVT U1705 ( .A(n24), .Y(n1549) );
  INVX0_HVT U1706 ( .A(n25), .Y(n1550) );
  INVX0_HVT U1707 ( .A(n28), .Y(n1551) );
  INVX0_HVT U1708 ( .A(n29), .Y(n1552) );
  INVX0_HVT U1709 ( .A(n30), .Y(n1553) );
  INVX0_HVT U1710 ( .A(n31), .Y(n1554) );
  INVX0_HVT U1711 ( .A(n226), .Y(n1555) );
  INVX0_HVT U1712 ( .A(n32), .Y(n1556) );
  INVX0_HVT U1713 ( .A(n33), .Y(n1557) );
  INVX0_HVT U1714 ( .A(n36), .Y(n1558) );
  INVX0_HVT U1715 ( .A(n37), .Y(n1559) );
  INVX0_HVT U1716 ( .A(n38), .Y(n1560) );
  INVX0_HVT U1717 ( .A(n39), .Y(n1561) );
  INVX0_HVT U1718 ( .A(n40), .Y(n1562) );
  INVX0_HVT U1719 ( .A(n41), .Y(n1563) );
  INVX0_HVT U1720 ( .A(n42), .Y(n1564) );
  INVX0_HVT U1721 ( .A(n74), .Y(n1565) );
  INVX0_HVT U1722 ( .A(n15), .Y(n1566) );
  INVX0_HVT U1723 ( .A(n62), .Y(n1567) );
  INVX0_HVT U1724 ( .A(n117), .Y(n1568) );
  INVX0_HVT U1725 ( .A(n216), .Y(n1569) );
  INVX0_HVT U1726 ( .A(n159), .Y(n1570) );
  INVX0_HVT U1727 ( .A(n221), .Y(n1571) );
  INVX0_HVT U1728 ( .A(n222), .Y(n1572) );
  INVX0_HVT U1729 ( .A(n224), .Y(n1574) );
  INVX0_HVT U1730 ( .A(n225), .Y(n1575) );
  INVX0_HVT U1731 ( .A(n97), .Y(n1576) );
  INVX0_HVT U1732 ( .A(n103), .Y(n1577) );
  INVX0_HVT U1733 ( .A(n227), .Y(n1578) );
  INVX0_HVT U1734 ( .A(n228), .Y(n1579) );
  INVX0_HVT U1735 ( .A(n229), .Y(n1580) );
  INVX0_HVT U1736 ( .A(n230), .Y(n1581) );
  INVX0_HVT U1737 ( .A(n231), .Y(n1582) );
  INVX0_HVT U1738 ( .A(n1232), .Y(n1588) );
  INVX0_HVT U1739 ( .A(n920), .Y(n1598) );
  INVX0_HVT U1740 ( .A(n937), .Y(n1599) );
  INVX0_HVT U1741 ( .A(n940), .Y(n1600) );
  INVX0_HVT U1742 ( .A(n949), .Y(n1601) );
  INVX0_HVT U1743 ( .A(n1088), .Y(n1602) );
  INVX0_HVT U1744 ( .A(n1128), .Y(n1603) );
  INVX0_HVT U1745 ( .A(n918), .Y(n1604) );
  INVX0_HVT U1746 ( .A(n931), .Y(n1605) );
  INVX0_HVT U1747 ( .A(n922), .Y(n1606) );
  INVX0_HVT U1748 ( .A(n921), .Y(n1607) );
  INVX0_HVT U1749 ( .A(n924), .Y(n1608) );
  INVX0_HVT U1750 ( .A(n925), .Y(n1609) );
  INVX0_HVT U1751 ( .A(n926), .Y(n1610) );
  INVX0_HVT U1752 ( .A(n927), .Y(n1611) );
  INVX0_HVT U1753 ( .A(n930), .Y(n1612) );
  INVX0_HVT U1754 ( .A(n932), .Y(n1613) );
  INVX0_HVT U1755 ( .A(n933), .Y(n1614) );
  INVX0_HVT U1756 ( .A(n934), .Y(n1615) );
  INVX0_HVT U1757 ( .A(n935), .Y(n1616) );
  INVX0_HVT U1758 ( .A(n936), .Y(n1617) );
  INVX0_HVT U1759 ( .A(n939), .Y(n1618) );
  INVX0_HVT U1760 ( .A(n941), .Y(n1619) );
  INVX0_HVT U1761 ( .A(n944), .Y(n1620) );
  INVX0_HVT U1762 ( .A(n945), .Y(n1621) );
  INVX0_HVT U1763 ( .A(n946), .Y(n1622) );
  INVX0_HVT U1764 ( .A(n1140), .Y(n1623) );
  INVX0_HVT U1765 ( .A(n947), .Y(n1624) );
  INVX0_HVT U1766 ( .A(n948), .Y(n1625) );
  INVX0_HVT U1767 ( .A(n950), .Y(n1626) );
  INVX0_HVT U1768 ( .A(n951), .Y(n1627) );
  INVX0_HVT U1769 ( .A(n952), .Y(n1628) );
  INVX0_HVT U1770 ( .A(n953), .Y(n1629) );
  INVX0_HVT U1771 ( .A(n954), .Y(n1630) );
  INVX0_HVT U1772 ( .A(n955), .Y(n1631) );
  INVX0_HVT U1773 ( .A(n956), .Y(n1632) );
  INVX0_HVT U1774 ( .A(n957), .Y(n1633) );
  INVX0_HVT U1775 ( .A(n960), .Y(n1634) );
  INVX0_HVT U1776 ( .A(n991), .Y(n1635) );
  INVX0_HVT U1777 ( .A(n928), .Y(n1636) );
  INVX0_HVT U1778 ( .A(n1031), .Y(n1637) );
  INVX0_HVT U1779 ( .A(n1129), .Y(n1638) );
  INVX0_HVT U1780 ( .A(n974), .Y(n1639) );
  INVX0_HVT U1781 ( .A(n1072), .Y(n1640) );
  INVX0_HVT U1782 ( .A(n1135), .Y(n1641) );
  INVX0_HVT U1783 ( .A(n1136), .Y(n1642) );
  INVX0_HVT U1784 ( .A(n1137), .Y(n1643) );
  INVX0_HVT U1785 ( .A(n1138), .Y(n1644) );
  INVX0_HVT U1786 ( .A(n1139), .Y(n1645) );
  INVX0_HVT U1787 ( .A(n1012), .Y(n1646) );
  INVX0_HVT U1788 ( .A(n1022), .Y(n1647) );
  INVX0_HVT U1789 ( .A(n1141), .Y(n1648) );
  INVX0_HVT U1790 ( .A(n1142), .Y(n1649) );
  INVX0_HVT U1791 ( .A(n1143), .Y(n1650) );
  INVX0_HVT U1792 ( .A(n1144), .Y(n1651) );
  INVX0_HVT U1793 ( .A(n1145), .Y(n1652) );
  INVX0_HVT U1794 ( .A(n1205), .Y(n1657) );
endmodule

