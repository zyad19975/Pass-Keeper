
module sbox_19 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n39, n45, n46, n48, n50, n72, n87, n142, n147, n160, n210, n211,
         n212, n213, n216, n217, n218, n219, n231, n232, n236, n238, n239,
         n240, n243, n246, n249, n251, n252, n257, n261, n264, n269, n275,
         n282, n283, n285, n289, n291, n293, n296, n297, n300, n301, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718;

  NAND2X0_HVT U4 ( .A1(n714), .A2(n301), .Y(n715) );
  NAND2X0_HVT U5 ( .A1(n297), .A2(n435), .Y(n713) );
  NAND2X0_HVT U15 ( .A1(n301), .A2(n355), .Y(n703) );
  NAND2X0_HVT U21 ( .A1(n438), .A2(n216), .Y(n697) );
  NAND2X0_HVT U24 ( .A1(n330), .A2(n377), .Y(n695) );
  NAND2X0_HVT U33 ( .A1(n315), .A2(n307), .Y(n686) );
  NAND2X0_HVT U35 ( .A1(n432), .A2(n450), .Y(n684) );
  NAND2X0_HVT U42 ( .A1(n240), .A2(n330), .Y(n678) );
  MUX41X1_HVT U51 ( .A1(n466), .A3(n490), .A2(n219), .A4(n359), .S0(n456), 
        .S1(n425), .Y(n673) );
  NAND2X0_HVT U53 ( .A1(n670), .A2(n677), .Y(n671) );
  NAND2X0_HVT U56 ( .A1(n438), .A2(n666), .Y(n667) );
  MUX41X1_HVT U57 ( .A1(n477), .A3(n699), .A2(n667), .A4(n708), .S0(n456), 
        .S1(n425), .Y(n665) );
  NAND2X0_HVT U58 ( .A1(n442), .A2(n301), .Y(n664) );
  MUX41X1_HVT U59 ( .A1(n416), .A3(n664), .A2(n415), .A4(n480), .S0(n458), 
        .S1(n425), .Y(n663) );
  MUX41X1_HVT U61 ( .A1(n410), .A3(n339), .A2(n329), .A4(n355), .S0(n458), 
        .S1(n425), .Y(n661) );
  NAND2X0_HVT U62 ( .A1(n239), .A2(n87), .Y(n660) );
  AO21X1_HVT U66 ( .A1(n502), .A2(n426), .A3(n311), .Y(n656) );
  NAND2X0_HVT U73 ( .A1(n285), .A2(n650), .Y(n651) );
  MUX41X1_HVT U75 ( .A1(n501), .A3(n499), .A2(n72), .A4(n399), .S0(n422), .S1(
        n391), .Y(n648) );
  NAND2X0_HVT U85 ( .A1(n377), .A2(n236), .Y(n638) );
  MUX41X1_HVT U86 ( .A1(n499), .A3(n638), .A2(n412), .A4(n408), .S0(n419), 
        .S1(n459), .Y(n637) );
  MUX41X1_HVT U90 ( .A1(n676), .A3(n678), .A2(n466), .A4(n635), .S0(n282), 
        .S1(n391), .Y(n634) );
  MUX41X1_HVT U97 ( .A1(n501), .A3(n413), .A2(n444), .A4(n703), .S0(n419), 
        .S1(n391), .Y(n626) );
  NAND2X0_HVT U101 ( .A1(n621), .A2(n620), .Y(n622) );
  MUX41X1_HVT U103 ( .A1(n301), .A3(n492), .A2(n481), .A4(n684), .S0(n282), 
        .S1(n458), .Y(n618) );
  OA21X1_HVT U109 ( .A1(n479), .A2(n453), .A3(n480), .Y(n613) );
  NAND2X0_HVT U110 ( .A1(n45), .A2(n611), .Y(n612) );
  AND2X1_HVT U115 ( .A1(n447), .A2(n355), .Y(n606) );
  MUX41X1_HVT U116 ( .A1(n706), .A3(n606), .A2(n399), .A4(n688), .S0(n308), 
        .S1(n457), .Y(n605) );
  NAND2X0_HVT U123 ( .A1(n597), .A2(n596), .Y(n598) );
  MUX41X1_HVT U131 ( .A1(n589), .A3(n591), .A2(n590), .A4(n592), .S0(n426), 
        .S1(n459), .Y(n588) );
  MUX41X1_HVT U132 ( .A1(n588), .A3(n601), .A2(n593), .A4(n607), .S0(n309), 
        .S1(n429), .Y(out[3]) );
  MUX41X1_HVT U136 ( .A1(n408), .A3(n686), .A2(n465), .A4(n683), .S0(n282), 
        .S1(n459), .Y(n585) );
  MUX41X1_HVT U139 ( .A1(n583), .A3(n257), .A2(n585), .A4(n586), .S0(n429), 
        .S1(n424), .Y(n582) );
  MUX41X1_HVT U147 ( .A1(n465), .A3(n650), .A2(n501), .A4(n676), .S0(n282), 
        .S1(n366), .Y(n576) );
  NAND2X0_HVT U158 ( .A1(n240), .A2(n236), .Y(n566) );
  MUX41X1_HVT U159 ( .A1(n706), .A3(n474), .A2(n566), .A4(n504), .S0(n418), 
        .S1(n251), .Y(n565) );
  AND2X1_HVT U162 ( .A1(n352), .A2(n650), .Y(n562) );
  MUX41X1_HVT U163 ( .A1(n339), .A3(n562), .A2(n411), .A4(n563), .S0(n418), 
        .S1(n457), .Y(n561) );
  NAND2X0_HVT U166 ( .A1(n442), .A2(n666), .Y(n558) );
  NAND2X0_HVT U167 ( .A1(n336), .A2(n216), .Y(n557) );
  MUX41X1_HVT U168 ( .A1(n477), .A3(n289), .A2(n557), .A4(n558), .S0(n418), 
        .S1(n456), .Y(n556) );
  MUX41X1_HVT U176 ( .A1(n232), .A3(n551), .A2(n473), .A4(n705), .S0(n458), 
        .S1(n421), .Y(n550) );
  NAND2X0_HVT U177 ( .A1(n369), .A2(n232), .Y(n549) );
  MUX41X1_HVT U178 ( .A1(n701), .A3(n549), .A2(n496), .A4(n400), .S0(n282), 
        .S1(n459), .Y(n548) );
  MUX41X1_HVT U179 ( .A1(n691), .A3(n495), .A2(n478), .A4(n496), .S0(n418), 
        .S1(n365), .Y(n547) );
  MUX41X1_HVT U180 ( .A1(n470), .A3(n710), .A2(n706), .A4(n409), .S0(n366), 
        .S1(n308), .Y(n546) );
  MUX41X1_HVT U189 ( .A1(n538), .A3(n705), .A2(n539), .A4(n489), .S0(n365), 
        .S1(n423), .Y(n537) );
  MUX41X1_HVT U190 ( .A1(n537), .A3(n540), .A2(n541), .A4(n544), .S0(n424), 
        .S1(n429), .Y(n536) );
  MUX41X1_HVT U193 ( .A1(n678), .A3(n684), .A2(n674), .A4(n535), .S0(n418), 
        .S1(n456), .Y(n534) );
  MUX41X1_HVT U194 ( .A1(n679), .A3(n692), .A2(n475), .A4(n291), .S0(n456), 
        .S1(n308), .Y(n533) );
  MUX41X1_HVT U195 ( .A1(n352), .A3(n500), .A2(n441), .A4(n682), .S0(n418), 
        .S1(n391), .Y(n532) );
  AO21X1_HVT U197 ( .A1(n412), .A2(n427), .A3(n498), .Y(n530) );
  MUX41X1_HVT U199 ( .A1(n529), .A3(n533), .A2(n532), .A4(n534), .S0(n429), 
        .S1(n160), .Y(n528) );
  MUX41X1_HVT U203 ( .A1(n683), .A3(n463), .A2(n707), .A4(n687), .S0(n418), 
        .S1(n456), .Y(n524) );
  MUX41X1_HVT U204 ( .A1(n667), .A3(n706), .A2(n503), .A4(n696), .S0(n418), 
        .S1(n458), .Y(n523) );
  MUX41X1_HVT U205 ( .A1(n325), .A3(n301), .A2(n495), .A4(n381), .S0(n418), 
        .S1(n459), .Y(n522) );
  NAND2X0_HVT U208 ( .A1(n240), .A2(n438), .Y(n611) );
  NAND2X0_HVT U212 ( .A1(n240), .A2(n285), .Y(n666) );
  NAND2X0_HVT U214 ( .A1(n353), .A2(n450), .Y(n520) );
  NAND2X0_HVT U215 ( .A1(n611), .A2(n289), .Y(n519) );
  NAND2X0_HVT U218 ( .A1(n293), .A2(n446), .Y(n572) );
  NAND2X0_HVT U220 ( .A1(n427), .A2(n520), .Y(n642) );
  INVX0_HVT U241 ( .A(n695), .Y(n507) );
  INVX0_HVT U242 ( .A(n678), .Y(n506) );
  INVX0_HVT U245 ( .A(n713), .Y(n504) );
  INVX0_HVT U250 ( .A(n708), .Y(n502) );
  INVX0_HVT U252 ( .A(n666), .Y(n501) );
  INVX0_HVT U255 ( .A(n515), .Y(n499) );
  INVX0_HVT U256 ( .A(n572), .Y(n498) );
  INVX0_HVT U261 ( .A(n509), .Y(n496) );
  INVX0_HVT U262 ( .A(n508), .Y(n495) );
  INVX0_HVT U267 ( .A(n707), .Y(n491) );
  INVX0_HVT U268 ( .A(n697), .Y(n490) );
  INVX0_HVT U270 ( .A(n519), .Y(n489) );
  INVX0_HVT U271 ( .A(n611), .Y(n488) );
  INVX0_HVT U273 ( .A(n630), .Y(n487) );
  INVX0_HVT U281 ( .A(n700), .Y(n480) );
  INVX0_HVT U282 ( .A(n682), .Y(n479) );
  INVX0_HVT U284 ( .A(n520), .Y(n478) );
  INVX0_HVT U285 ( .A(n517), .Y(n477) );
  INVX0_HVT U289 ( .A(n620), .Y(n473) );
  INVX0_HVT U295 ( .A(n715), .Y(n470) );
  INVX0_HVT U296 ( .A(n703), .Y(n469) );
  INVX0_HVT U300 ( .A(n679), .Y(n467) );
  INVX0_HVT U303 ( .A(n510), .Y(n465) );
  INVX0_HVT U306 ( .A(n557), .Y(n464) );
  INVX1_HVT U1 ( .A(n356), .Y(n357) );
  MUX21X1_HVT U2 ( .A1(n236), .A2(n357), .S0(n307), .Y(n711) );
  INVX1_HVT U3 ( .A(n714), .Y(n315) );
  MUX21X1_HVT U6 ( .A1(n326), .A2(n432), .S0(n447), .Y(n296) );
  MUX21X1_HVT U7 ( .A1(n45), .A2(n633), .S0(n414), .Y(n632) );
  INVX1_HVT U8 ( .A(n435), .Y(n330) );
  INVX1_HVT U9 ( .A(n417), .Y(n418) );
  MUX21X1_HVT U10 ( .A1(n526), .A2(n527), .S0(n421), .Y(n525) );
  XOR2X1_HVT U11 ( .A1(n307), .A2(n422), .Y(n347) );
  INVX1_HVT U12 ( .A(n329), .Y(n702) );
  AO21X1_HVT U13 ( .A1(n423), .A2(n285), .A3(n353), .Y(n603) );
  INVX1_HVT U14 ( .A(n46), .Y(n647) );
  AND3X1_HVT U16 ( .A1(n87), .A2(n666), .A3(n642), .Y(n643) );
  INVX1_HVT U17 ( .A(n704), .Y(n468) );
  INVX1_HVT U18 ( .A(n453), .Y(n452) );
  XNOR2X1_HVT U19 ( .A1(n444), .A2(n291), .Y(n23) );
  INVX1_HVT U20 ( .A(in[0]), .Y(n39) );
  NBUFFX2_HVT U22 ( .A(n87), .Y(n440) );
  MUX41X1_HVT U23 ( .A1(n524), .A3(n522), .A2(n525), .A4(n523), .S0(n39), .S1(
        n160), .Y(n521) );
  INVX0_HVT U25 ( .A(n72), .Y(n45) );
  MUX21X1_HVT U26 ( .A1(n673), .A2(n669), .S0(n378), .Y(n668) );
  MUX41X1_HVT U27 ( .A1(n619), .A3(n623), .A2(n616), .A4(n618), .S0(n424), 
        .S1(n39), .Y(n615) );
  MUX41X1_HVT U28 ( .A1(n497), .A3(n617), .A2(n675), .A4(n489), .S0(n391), 
        .S1(n452), .Y(n616) );
  XOR2X1_HVT U29 ( .A1(n371), .A2(n330), .Y(n675) );
  MUX21X2_HVT U30 ( .A1(n353), .A2(n336), .S0(n297), .Y(n694) );
  INVX1_HVT U31 ( .A(n474), .Y(n353) );
  MUX21X2_HVT U32 ( .A1(n354), .A2(n330), .S0(n310), .Y(n329) );
  INVX0_HVT U34 ( .A(n430), .Y(n505) );
  MUX41X1_HVT U36 ( .A1(n359), .A3(n23), .A2(n704), .A4(n507), .S0(n362), .S1(
        n458), .Y(n640) );
  INVX1_HVT U37 ( .A(n712), .Y(n351) );
  INVX0_HVT U38 ( .A(n306), .Y(n303) );
  INVX1_HVT U39 ( .A(n518), .Y(n466) );
  MUX21X1_HVT U40 ( .A1(n351), .A2(n325), .S0(n370), .Y(n46) );
  MUX41X1_HVT U41 ( .A1(n646), .A3(n649), .A2(n648), .A4(n653), .S0(n429), 
        .S1(n425), .Y(n645) );
  INVX0_HVT U43 ( .A(n351), .Y(n352) );
  MUX21X1_HVT U44 ( .A1(n395), .A2(n394), .S0(n323), .Y(n639) );
  INVX1_HVT U45 ( .A(n451), .Y(n417) );
  INVX1_HVT U46 ( .A(in[7]), .Y(n460) );
  INVX1_HVT U47 ( .A(in[7]), .Y(n461) );
  INVX1_HVT U48 ( .A(n461), .Y(n391) );
  MUX21X1_HVT U49 ( .A1(n439), .A2(n328), .S0(n239), .Y(n698) );
  INVX1_HVT U50 ( .A(n511), .Y(n475) );
  NAND2X0_HVT U52 ( .A1(n542), .A2(n321), .Y(n349) );
  OA21X1_HVT U54 ( .A1(n685), .A2(n460), .A3(n472), .Y(n542) );
  INVX1_HVT U55 ( .A(n461), .Y(n458) );
  INVX1_HVT U60 ( .A(n461), .Y(n456) );
  MUX21X1_HVT U63 ( .A1(n578), .A2(n579), .S0(n378), .Y(n577) );
  INVX1_HVT U64 ( .A(n420), .Y(n312) );
  INVX1_HVT U65 ( .A(n461), .Y(n459) );
  MUX21X1_HVT U67 ( .A1(n701), .A2(n482), .S0(n282), .Y(n589) );
  AND3X1_HVT U68 ( .A1(n422), .A2(n216), .A3(n325), .Y(n591) );
  INVX1_HVT U69 ( .A(n321), .Y(n308) );
  MUX21X1_HVT U70 ( .A1(n599), .A2(n598), .S0(n457), .Y(n595) );
  NAND2X0_HVT U71 ( .A1(n483), .A2(n378), .Y(n379) );
  MUX21X1_HVT U72 ( .A1(n275), .A2(n716), .S0(n419), .Y(n614) );
  NAND2X0_HVT U74 ( .A1(n536), .A2(n348), .Y(n396) );
  MUX21X1_HVT U76 ( .A1(n330), .A2(n432), .S0(n428), .Y(n633) );
  AO21X1_HVT U77 ( .A1(n456), .A2(n630), .A3(n498), .Y(n631) );
  MUX21X1_HVT U78 ( .A1(n431), .A2(n486), .S0(n446), .Y(n628) );
  AO21X1_HVT U79 ( .A1(n239), .A2(n261), .A3(n460), .Y(n621) );
  INVX1_HVT U80 ( .A(n690), .Y(n481) );
  MUX21X1_HVT U81 ( .A1(n486), .A2(n336), .S0(n369), .Y(n551) );
  INVX1_HVT U82 ( .A(n328), .Y(n232) );
  INVX1_HVT U83 ( .A(n147), .Y(n574) );
  MUX21X1_HVT U84 ( .A1(n530), .A2(n531), .S0(n321), .Y(n529) );
  MUX21X1_HVT U87 ( .A1(n506), .A2(n496), .S0(n427), .Y(n531) );
  OA21X1_HVT U88 ( .A1(n464), .A2(n460), .A3(n688), .Y(n578) );
  INVX1_HVT U89 ( .A(n311), .Y(n650) );
  INVX1_HVT U91 ( .A(n275), .Y(n683) );
  NBUFFX2_HVT U92 ( .A(n452), .Y(n420) );
  INVX1_HVT U93 ( .A(n342), .Y(n706) );
  MUX21X1_HVT U94 ( .A1(n503), .A2(n493), .S0(n362), .Y(n604) );
  INVX0_HVT U95 ( .A(n420), .Y(n362) );
  INVX1_HVT U96 ( .A(n327), .Y(n693) );
  INVX1_HVT U98 ( .A(n219), .Y(n699) );
  NAND2X0_HVT U99 ( .A1(n671), .A2(n323), .Y(n363) );
  OA21X1_HVT U100 ( .A1(n415), .A2(n460), .A3(n688), .Y(n554) );
  MUX21X1_HVT U102 ( .A1(n595), .A2(n594), .S0(n210), .Y(n593) );
  INVX0_HVT U104 ( .A(n420), .Y(n321) );
  INVX1_HVT U105 ( .A(n456), .Y(n346) );
  INVX1_HVT U106 ( .A(n460), .Y(n457) );
  INVX0_HVT U107 ( .A(n455), .Y(n160) );
  INVX0_HVT U108 ( .A(in[5]), .Y(n455) );
  INVX1_HVT U111 ( .A(n377), .Y(n297) );
  INVX0_HVT U112 ( .A(n424), .Y(n210) );
  INVX1_HVT U113 ( .A(n376), .Y(n371) );
  INVX1_HVT U114 ( .A(n371), .Y(n307) );
  INVX0_HVT U117 ( .A(n709), .Y(n283) );
  INVX1_HVT U118 ( .A(n448), .Y(n239) );
  INVX0_HVT U119 ( .A(n711), .Y(n471) );
  INVX0_HVT U120 ( .A(n339), .Y(n701) );
  INVX1_HVT U121 ( .A(n433), .Y(n328) );
  MUX21X1_HVT U122 ( .A1(n486), .A2(n328), .S0(n445), .Y(n687) );
  INVX0_HVT U124 ( .A(n291), .Y(n261) );
  INVX1_HVT U125 ( .A(n376), .Y(n448) );
  INVX0_HVT U126 ( .A(n211), .Y(n216) );
  INVX1_HVT U127 ( .A(n310), .Y(n450) );
  NBUFFX2_HVT U128 ( .A(n454), .Y(n426) );
  MUX41X1_HVT U129 ( .A1(n639), .A3(n641), .A2(n637), .A4(n640), .S0(n429), 
        .S1(n210), .Y(n636) );
  INVX0_HVT U130 ( .A(n331), .Y(n395) );
  INVX0_HVT U133 ( .A(n689), .Y(n48) );
  INVX1_HVT U134 ( .A(n48), .Y(n50) );
  MUX21X1_HVT U135 ( .A1(n50), .A2(n497), .S0(n312), .Y(n592) );
  MUX21X1_HVT U137 ( .A1(n492), .A2(n293), .S0(n426), .Y(n655) );
  INVX0_HVT U138 ( .A(n710), .Y(n492) );
  MUX41X1_HVT U140 ( .A1(n656), .A3(n471), .A2(n657), .A4(n655), .S0(n362), 
        .S1(n428), .Y(n654) );
  MUX41X1_HVT U141 ( .A1(n559), .A3(n553), .A2(n561), .A4(n556), .S0(n39), 
        .S1(n424), .Y(n552) );
  NBUFFX2_HVT U142 ( .A(n505), .Y(n434) );
  MUX21X1_HVT U143 ( .A1(n491), .A2(n450), .S0(n426), .Y(n657) );
  INVX0_HVT U144 ( .A(n717), .Y(n72) );
  INVX1_HVT U145 ( .A(n72), .Y(n87) );
  MUX21X1_HVT U146 ( .A1(n336), .A2(n261), .S0(n450), .Y(n560) );
  INVX0_HVT U148 ( .A(n702), .Y(n142) );
  MUX21X1_HVT U149 ( .A1(n437), .A2(n514), .S0(n249), .Y(n147) );
  MUX41X1_HVT U150 ( .A1(n570), .A3(n565), .A2(n571), .A4(n567), .S0(n39), 
        .S1(n160), .Y(n564) );
  MUX41X1_HVT U151 ( .A1(n550), .A3(n547), .A2(n548), .A4(n546), .S0(n39), 
        .S1(n210), .Y(n545) );
  INVX1_HVT U152 ( .A(n354), .Y(n355) );
  NBUFFX2_HVT U153 ( .A(n494), .Y(n433) );
  INVX0_HVT U154 ( .A(n449), .Y(n211) );
  INVX1_HVT U155 ( .A(n449), .Y(n445) );
  INVX0_HVT U156 ( .A(n448), .Y(n449) );
  MUX21X2_HVT U157 ( .A1(n644), .A2(n643), .S0(n423), .Y(n641) );
  NAND2X0_HVT U160 ( .A1(n573), .A2(n378), .Y(n212) );
  NAND2X0_HVT U161 ( .A1(n574), .A2(n423), .Y(n213) );
  NAND2X0_HVT U164 ( .A1(n212), .A2(n213), .Y(n571) );
  NAND2X0_HVT U165 ( .A1(n434), .A2(n216), .Y(n217) );
  NAND2X0_HVT U169 ( .A1(n352), .A2(n446), .Y(n218) );
  NAND2X0_HVT U170 ( .A1(n217), .A2(n218), .Y(n514) );
  INVX0_HVT U171 ( .A(n449), .Y(n446) );
  INVX0_HVT U172 ( .A(n514), .Y(n476) );
  INVX0_HVT U173 ( .A(n698), .Y(n359) );
  MUX21X1_HVT U174 ( .A1(n439), .A2(n436), .S0(n445), .Y(n219) );
  OA21X1_HVT U175 ( .A1(n680), .A2(n460), .A3(n572), .Y(n573) );
  MUX41X1_HVT U181 ( .A1(n627), .A3(n626), .A2(n634), .A4(n629), .S0(n210), 
        .S1(n429), .Y(n625) );
  MUX41X1_HVT U182 ( .A1(n560), .A3(n676), .A2(n48), .A4(n697), .S0(n346), 
        .S1(n417), .Y(n559) );
  MUX41X1_HVT U183 ( .A1(n476), .A3(n647), .A2(n487), .A4(n710), .S0(n323), 
        .S1(n453), .Y(n646) );
  MUX21X1_HVT U184 ( .A1(n554), .A2(n555), .S0(n378), .Y(n553) );
  INVX1_HVT U185 ( .A(in[2]), .Y(n453) );
  INVX1_HVT U186 ( .A(n516), .Y(n500) );
  INVX0_HVT U187 ( .A(n712), .Y(n474) );
  INVX1_HVT U188 ( .A(n430), .Y(n306) );
  NAND2X0_HVT U191 ( .A1(n433), .A2(n505), .Y(n231) );
  INVX0_HVT U192 ( .A(n351), .Y(n354) );
  NBUFFX2_HVT U196 ( .A(n714), .Y(n438) );
  INVX1_HVT U198 ( .A(n385), .Y(n400) );
  OA21X1_HVT U200 ( .A1(n460), .A2(n711), .A3(n385), .Y(n526) );
  INVX0_HVT U201 ( .A(n398), .Y(n581) );
  INVX1_HVT U202 ( .A(n318), .Y(n692) );
  MUX41X1_HVT U206 ( .A1(n576), .A3(n580), .A2(n577), .A4(n581), .S0(n429), 
        .S1(n424), .Y(n575) );
  INVX0_HVT U207 ( .A(n442), .Y(n236) );
  INVX1_HVT U209 ( .A(n252), .Y(n238) );
  INVX1_HVT U210 ( .A(n494), .Y(n252) );
  MUX21X1_HVT U211 ( .A1(n443), .A2(n432), .S0(n450), .Y(n275) );
  NAND2X0_HVT U213 ( .A1(n238), .A2(n306), .Y(n714) );
  MUX21X1_HVT U216 ( .A1(n689), .A2(n519), .S0(n366), .Y(n513) );
  INVX0_HVT U217 ( .A(n441), .Y(n382) );
  INVX1_HVT U219 ( .A(n296), .Y(n689) );
  MUX21X1_HVT U221 ( .A1(n353), .A2(n714), .S0(n450), .Y(n682) );
  IBUFFX2_HVT U222 ( .A(n449), .Y(n370) );
  NBUFFX2_HVT U223 ( .A(n310), .Y(n240) );
  IBUFFX2_HVT U224 ( .A(n376), .Y(n310) );
  INVX1_HVT U225 ( .A(n319), .Y(n653) );
  INVX1_HVT U226 ( .A(in[4]), .Y(n494) );
  INVX0_HVT U227 ( .A(n239), .Y(n447) );
  INVX0_HVT U228 ( .A(n448), .Y(n377) );
  INVX0_HVT U229 ( .A(n324), .Y(n600) );
  INVX1_HVT U230 ( .A(n449), .Y(n369) );
  INVX0_HVT U231 ( .A(n694), .Y(n399) );
  NBUFFX2_HVT U232 ( .A(n306), .Y(n436) );
  NAND2X0_HVT U233 ( .A1(n603), .A2(n323), .Y(n243) );
  NAND2X0_HVT U234 ( .A1(n604), .A2(n427), .Y(n246) );
  NAND2X0_HVT U235 ( .A1(n243), .A2(n246), .Y(n602) );
  INVX0_HVT U236 ( .A(n388), .Y(n249) );
  INVX1_HVT U237 ( .A(n249), .Y(n251) );
  INVX0_HVT U238 ( .A(n461), .Y(n388) );
  MUX21X1_HVT U239 ( .A1(n432), .A2(n437), .S0(n371), .Y(n339) );
  INVX1_HVT U240 ( .A(n685), .Y(n503) );
  MUX21X1_HVT U243 ( .A1(n622), .A2(n462), .S0(n422), .Y(n619) );
  MUX41X1_HVT U244 ( .A1(n713), .A3(n692), .A2(n475), .A4(n261), .S0(n421), 
        .S1(n460), .Y(n257) );
  MUX21X1_HVT U246 ( .A1(n352), .A2(n293), .S0(n211), .Y(n511) );
  INVX1_HVT U247 ( .A(in[1]), .Y(n376) );
  MUX21X1_HVT U248 ( .A1(n431), .A2(n326), .S0(n447), .Y(n696) );
  MUX21X1_HVT U249 ( .A1(n432), .A2(n486), .S0(n297), .Y(n690) );
  NAND2X0_HVT U251 ( .A1(n715), .A2(n308), .Y(n264) );
  NAND2X0_HVT U253 ( .A1(n584), .A2(n312), .Y(n269) );
  NAND2X0_HVT U254 ( .A1(n264), .A2(n269), .Y(n583) );
  MUX21X1_HVT U257 ( .A1(n381), .A2(n704), .S0(n423), .Y(n624) );
  MUX21X2_HVT U258 ( .A1(n437), .A2(n440), .S0(n239), .Y(n704) );
  MUX41X1_HVT U259 ( .A1(n351), .A3(n472), .A2(n289), .A4(n488), .S0(n321), 
        .S1(n457), .Y(n580) );
  MUX21X1_HVT U260 ( .A1(n328), .A2(n443), .S0(n450), .Y(n691) );
  NBUFFX2_HVT U263 ( .A(n452), .Y(n282) );
  INVX0_HVT U264 ( .A(n283), .Y(n285) );
  INVX0_HVT U265 ( .A(n283), .Y(n289) );
  INVX0_HVT U266 ( .A(n283), .Y(n291) );
  INVX1_HVT U269 ( .A(n437), .Y(n293) );
  NBUFFX2_HVT U272 ( .A(in[3]), .Y(n430) );
  NBUFFX2_HVT U274 ( .A(n494), .Y(n432) );
  INVX0_HVT U275 ( .A(n716), .Y(n300) );
  INVX1_HVT U276 ( .A(n300), .Y(n301) );
  NAND2X0_HVT U277 ( .A1(n444), .A2(n87), .Y(n716) );
  INVX0_HVT U278 ( .A(n680), .Y(n463) );
  MUX41X1_HVT U279 ( .A1(n658), .A3(n654), .A2(n668), .A4(n662), .S0(n39), 
        .S1(n309), .Y(out[0]) );
  MUX21X2_HVT U280 ( .A1(n661), .A2(n659), .S0(n378), .Y(n658) );
  INVX1_HVT U283 ( .A(n439), .Y(n336) );
  NAND2X0_HVT U286 ( .A1(n433), .A2(n505), .Y(n304) );
  NAND2X0_HVT U287 ( .A1(n252), .A2(n303), .Y(n305) );
  NAND2X0_HVT U288 ( .A1(n305), .A2(n231), .Y(n712) );
  INVX1_HVT U290 ( .A(n696), .Y(n472) );
  MUX21X1_HVT U291 ( .A1(n377), .A2(n716), .S0(n312), .Y(n596) );
  MUX41X1_HVT U292 ( .A1(n697), .A3(n416), .A2(n471), .A4(n485), .S0(n308), 
        .S1(n391), .Y(n594) );
  INVX1_HVT U293 ( .A(n348), .Y(n309) );
  INVX1_HVT U294 ( .A(in[6]), .Y(n348) );
  NOR2X0_HVT U297 ( .A1(n307), .A2(n382), .Y(n311) );
  INVX1_HVT U298 ( .A(n691), .Y(n497) );
  NAND2X0_HVT U299 ( .A1(n300), .A2(n365), .Y(n313) );
  NAND2X0_HVT U301 ( .A1(n690), .A2(n323), .Y(n314) );
  NAND2X0_HVT U302 ( .A1(n313), .A2(n314), .Y(n579) );
  INVX1_HVT U304 ( .A(n687), .Y(n482) );
  NAND2X0_HVT U305 ( .A1(n484), .A2(n365), .Y(n316) );
  NAND2X0_HVT U307 ( .A1(n696), .A2(n323), .Y(n317) );
  NAND2X0_HVT U308 ( .A1(n316), .A2(n317), .Y(n584) );
  INVX1_HVT U309 ( .A(n681), .Y(n484) );
  MUX21X1_HVT U310 ( .A1(n87), .A2(n443), .S0(n444), .Y(n318) );
  MUX21X1_HVT U311 ( .A1(n320), .A2(n338), .S0(n421), .Y(n319) );
  XOR2X2_HVT U312 ( .A1(n251), .A2(n692), .Y(n320) );
  INVX0_HVT U313 ( .A(n432), .Y(n325) );
  INVX1_HVT U314 ( .A(n304), .Y(n486) );
  MUX21X1_HVT U315 ( .A1(n289), .A2(n500), .S0(n428), .Y(n555) );
  INVX1_HVT U316 ( .A(n365), .Y(n323) );
  INVX0_HVT U317 ( .A(n322), .Y(n394) );
  INVX1_HVT U318 ( .A(n436), .Y(n326) );
  MUX21X1_HVT U319 ( .A1(n351), .A2(n696), .S0(n312), .Y(n322) );
  INVX1_HVT U320 ( .A(n376), .Y(n444) );
  MUX41X1_HVT U321 ( .A1(n507), .A3(n413), .A2(n500), .A4(n628), .S0(n419), 
        .S1(n459), .Y(n627) );
  MUX21X1_HVT U322 ( .A1(n325), .A2(n326), .S0(n369), .Y(n324) );
  XNOR2X1_HVT U323 ( .A1(n328), .A2(n307), .Y(n327) );
  MUX41X1_HVT U324 ( .A1(n467), .A3(n327), .A2(n484), .A4(n304), .S0(n251), 
        .S1(n417), .Y(n544) );
  MUX21X1_HVT U325 ( .A1(n329), .A2(n332), .S0(n419), .Y(n331) );
  NAND2X0_HVT U326 ( .A1(n444), .A2(n325), .Y(n332) );
  NAND2X0_HVT U327 ( .A1(n142), .A2(n423), .Y(n333) );
  NAND2X0_HVT U328 ( .A1(n411), .A2(n312), .Y(n334) );
  NAND2X0_HVT U329 ( .A1(n333), .A2(n334), .Y(n590) );
  INVX1_HVT U330 ( .A(n512), .Y(n485) );
  INVX1_HVT U331 ( .A(n335), .Y(n569) );
  MUX21X1_HVT U332 ( .A1(n337), .A2(n336), .S0(n414), .Y(n335) );
  NAND2X0_HVT U333 ( .A1(n365), .A2(n330), .Y(n337) );
  MUX41X1_HVT U334 ( .A1(n693), .A3(n652), .A2(n695), .A4(n651), .S0(n362), 
        .S1(n366), .Y(n649) );
  MUX21X1_HVT U335 ( .A1(n441), .A2(n516), .S0(n427), .Y(n338) );
  MUX21X1_HVT U336 ( .A1(n289), .A2(n432), .S0(n370), .Y(n652) );
  NBUFFX2_HVT U337 ( .A(n709), .Y(n437) );
  MUX21X1_HVT U338 ( .A1(n436), .A2(n438), .S0(n377), .Y(n707) );
  NAND2X0_HVT U339 ( .A1(n688), .A2(n378), .Y(n340) );
  NAND2X0_HVT U340 ( .A1(n612), .A2(n423), .Y(n341) );
  NAND2X0_HVT U341 ( .A1(n341), .A2(n340), .Y(n610) );
  MUX21X2_HVT U342 ( .A1(n564), .A2(n552), .S0(n348), .Y(out[5]) );
  NAND2X0_HVT U343 ( .A1(n521), .A2(n348), .Y(n360) );
  INVX0_HVT U344 ( .A(n358), .Y(n644) );
  OR2X1_HVT U345 ( .A1(n239), .A2(n351), .Y(n705) );
  AND2X1_HVT U346 ( .A1(n705), .A2(n442), .Y(n342) );
  MUX41X1_HVT U347 ( .A1(n608), .A3(n610), .A2(n614), .A4(n613), .S0(n427), 
        .S1(n426), .Y(n607) );
  NAND2X0_HVT U348 ( .A1(n45), .A2(n343), .Y(n344) );
  NAND2X0_HVT U349 ( .A1(n609), .A2(n347), .Y(n345) );
  NAND2X0_HVT U350 ( .A1(n344), .A2(n345), .Y(n608) );
  INVX0_HVT U351 ( .A(n347), .Y(n343) );
  MUX41X1_HVT U352 ( .A1(n469), .A3(n660), .A2(n468), .A4(n342), .S0(n346), 
        .S1(n425), .Y(n659) );
  XOR2X2_HVT U353 ( .A1(n353), .A2(n371), .Y(n676) );
  MUX21X2_HVT U354 ( .A1(n645), .A2(n636), .S0(n348), .Y(out[1]) );
  NAND2X0_HVT U355 ( .A1(n543), .A2(n421), .Y(n350) );
  NAND2X0_HVT U356 ( .A1(n349), .A2(n350), .Y(n541) );
  MUX21X1_HVT U357 ( .A1(n638), .A2(n326), .S0(n427), .Y(n543) );
  INVX1_HVT U358 ( .A(n431), .Y(n356) );
  MUX21X1_HVT U359 ( .A1(n359), .A2(n261), .S0(n251), .Y(n358) );
  NAND2X0_HVT U360 ( .A1(n528), .A2(n309), .Y(n361) );
  NAND2X0_HVT U361 ( .A1(n360), .A2(n361), .Y(out[7]) );
  NAND2X0_HVT U362 ( .A1(n615), .A2(n348), .Y(n402) );
  MUX41X1_HVT U363 ( .A1(n410), .A3(n612), .A2(n493), .A4(n439), .S0(n362), 
        .S1(n251), .Y(n570) );
  INVX0_HVT U364 ( .A(n686), .Y(n483) );
  NAND2X0_HVT U365 ( .A1(n672), .A2(n366), .Y(n364) );
  NAND2X0_HVT U366 ( .A1(n363), .A2(n364), .Y(n669) );
  MUX21X1_HVT U367 ( .A1(n330), .A2(n684), .S0(n426), .Y(n672) );
  INVX0_HVT U368 ( .A(n684), .Y(n493) );
  NBUFFX2_HVT U369 ( .A(n388), .Y(n365) );
  NBUFFX2_HVT U370 ( .A(n388), .Y(n366) );
  NAND2X0_HVT U371 ( .A1(n587), .A2(n419), .Y(n367) );
  NAND2X0_HVT U372 ( .A1(n378), .A2(n462), .Y(n368) );
  NAND2X0_HVT U373 ( .A1(n367), .A2(n368), .Y(n586) );
  INVX1_HVT U374 ( .A(n513), .Y(n462) );
  NAND2X0_HVT U375 ( .A1(n582), .A2(n309), .Y(n387) );
  NAND2X0_HVT U376 ( .A1(n702), .A2(n323), .Y(n372) );
  NAND2X0_HVT U377 ( .A1(n409), .A2(n366), .Y(n373) );
  NAND2X0_HVT U378 ( .A1(n372), .A2(n373), .Y(n527) );
  NAND2X0_HVT U379 ( .A1(n631), .A2(n362), .Y(n374) );
  NAND2X0_HVT U380 ( .A1(n632), .A2(n423), .Y(n375) );
  NAND2X0_HVT U381 ( .A1(n375), .A2(n374), .Y(n629) );
  INVX1_HVT U382 ( .A(n381), .Y(n688) );
  NAND2X0_HVT U383 ( .A1(n600), .A2(n419), .Y(n380) );
  NAND2X0_HVT U384 ( .A1(n379), .A2(n380), .Y(n599) );
  INVX0_HVT U385 ( .A(n420), .Y(n378) );
  MUX21X1_HVT U386 ( .A1(n382), .A2(n293), .S0(n445), .Y(n381) );
  NAND2X0_HVT U387 ( .A1(n569), .A2(n423), .Y(n383) );
  NAND2X0_HVT U388 ( .A1(n568), .A2(n362), .Y(n384) );
  NAND2X0_HVT U389 ( .A1(n383), .A2(n384), .Y(n567) );
  MUX21X1_HVT U390 ( .A1(n441), .A2(n304), .S0(n445), .Y(n385) );
  MUX21X1_HVT U391 ( .A1(n400), .A2(n487), .S0(n251), .Y(n568) );
  NAND2X0_HVT U392 ( .A1(n575), .A2(n348), .Y(n386) );
  NAND2X0_HVT U393 ( .A1(n386), .A2(n387), .Y(out[4]) );
  NAND2X0_HVT U394 ( .A1(n663), .A2(n312), .Y(n389) );
  NAND2X0_HVT U395 ( .A1(n665), .A2(n421), .Y(n390) );
  NAND2X0_HVT U396 ( .A1(n389), .A2(n390), .Y(n662) );
  NAND2X0_HVT U397 ( .A1(n602), .A2(n210), .Y(n392) );
  NAND2X0_HVT U398 ( .A1(n605), .A2(n426), .Y(n393) );
  NAND2X0_HVT U399 ( .A1(n392), .A2(n393), .Y(n601) );
  NAND2X0_HVT U400 ( .A1(n545), .A2(n309), .Y(n397) );
  NAND2X0_HVT U401 ( .A1(n396), .A2(n397), .Y(out[6]) );
  MUX41X1_HVT U402 ( .A1(n681), .A3(n413), .A2(n676), .A4(n650), .S0(n417), 
        .S1(n458), .Y(n540) );
  XNOR2X1_HVT U403 ( .A1(n421), .A2(n427), .Y(n407) );
  NAND2X0_HVT U404 ( .A1(n625), .A2(n309), .Y(n403) );
  MUX41X1_HVT U405 ( .A1(n401), .A3(n687), .A2(n399), .A4(n400), .S0(n282), 
        .S1(n460), .Y(n398) );
  NAND2X0_HVT U406 ( .A1(n291), .A2(n216), .Y(n401) );
  NAND2X0_HVT U407 ( .A1(n403), .A2(n402), .Y(out[2]) );
  NAND2X0_HVT U408 ( .A1(n624), .A2(n404), .Y(n405) );
  NAND2X0_HVT U409 ( .A1(n410), .A2(n407), .Y(n406) );
  NAND2X0_HVT U410 ( .A1(n405), .A2(n406), .Y(n623) );
  INVX0_HVT U411 ( .A(n407), .Y(n404) );
  INVX1_HVT U412 ( .A(n455), .Y(n454) );
  MUX21X1_HVT U413 ( .A1(n485), .A2(n289), .S0(n365), .Y(n587) );
  AND2X1_HVT U414 ( .A1(n45), .A2(n650), .Y(n408) );
  AND2X1_HVT U415 ( .A1(n355), .A2(n666), .Y(n409) );
  AND2X1_HVT U416 ( .A1(n442), .A2(n611), .Y(n410) );
  NBUFFX2_HVT U417 ( .A(n474), .Y(n431) );
  MUX21X1_HVT U418 ( .A1(n289), .A2(n443), .S0(n422), .Y(n597) );
  MUX21X1_HVT U419 ( .A1(n382), .A2(n435), .S0(n369), .Y(n685) );
  MUX21X1_HVT U420 ( .A1(n45), .A2(n357), .S0(n211), .Y(n679) );
  MUX21X1_HVT U421 ( .A1(n436), .A2(n236), .S0(n371), .Y(n708) );
  MUX21X1_HVT U422 ( .A1(n436), .A2(n336), .S0(n446), .Y(n680) );
  MUX21X1_HVT U423 ( .A1(n236), .A2(n355), .S0(n370), .Y(n563) );
  XOR2X1_HVT U424 ( .A1(n45), .A2(n371), .Y(n674) );
  MUX21X1_HVT U425 ( .A1(n434), .A2(n232), .S0(n370), .Y(n535) );
  MUX21X1_HVT U426 ( .A1(n438), .A2(n291), .S0(n445), .Y(n635) );
  MUX21X1_HVT U427 ( .A1(n285), .A2(n435), .S0(n370), .Y(n516) );
  MUX21X1_HVT U428 ( .A1(n293), .A2(n315), .S0(n297), .Y(n700) );
  MUX21X1_HVT U429 ( .A1(n357), .A2(n232), .S0(n369), .Y(n620) );
  MUX21X1_HVT U430 ( .A1(n434), .A2(n443), .S0(n446), .Y(n538) );
  MUX21X1_HVT U431 ( .A1(n441), .A2(n440), .S0(n446), .Y(n539) );
  MUX21X1_HVT U432 ( .A1(n440), .A2(n232), .S0(n211), .Y(n518) );
  MUX21X1_HVT U433 ( .A1(n304), .A2(n443), .S0(n444), .Y(n630) );
  MUX21X1_HVT U434 ( .A1(n486), .A2(n232), .S0(n240), .Y(n512) );
  XNOR2X1_HVT U435 ( .A1(n304), .A2(n444), .Y(n411) );
  MUX21X1_HVT U436 ( .A1(n440), .A2(n438), .S0(n444), .Y(n510) );
  MUX21X1_HVT U437 ( .A1(n315), .A2(n236), .S0(n426), .Y(n670) );
  XOR2X1_HVT U438 ( .A1(n211), .A2(n160), .Y(n677) );
  XNOR2X1_HVT U439 ( .A1(n441), .A2(n369), .Y(n412) );
  AND2X1_HVT U440 ( .A1(n240), .A2(n336), .Y(n413) );
  NBUFFX2_HVT U441 ( .A(n718), .Y(n441) );
  NBUFFX2_HVT U442 ( .A(n306), .Y(n435) );
  NBUFFX2_HVT U443 ( .A(n717), .Y(n439) );
  NBUFFX2_HVT U444 ( .A(n718), .Y(n443) );
  NBUFFX2_HVT U445 ( .A(n718), .Y(n442) );
  NBUFFX2_HVT U446 ( .A(n388), .Y(n428) );
  NBUFFX2_HVT U447 ( .A(n388), .Y(n427) );
  NBUFFX2_HVT U448 ( .A(n451), .Y(n423) );
  NBUFFX2_HVT U449 ( .A(n454), .Y(n425) );
  NBUFFX2_HVT U450 ( .A(n452), .Y(n422) );
  NBUFFX2_HVT U451 ( .A(n451), .Y(n421) );
  NBUFFX2_HVT U452 ( .A(n452), .Y(n419) );
  NBUFFX2_HVT U453 ( .A(n160), .Y(n424) );
  MUX21X1_HVT U454 ( .A1(n714), .A2(n326), .S0(n297), .Y(n710) );
  MUX21X1_HVT U455 ( .A1(n330), .A2(n315), .S0(n211), .Y(n681) );
  MUX21X1_HVT U456 ( .A1(n328), .A2(n285), .S0(n369), .Y(n509) );
  MUX21X1_HVT U457 ( .A1(n285), .A2(n431), .S0(n445), .Y(n617) );
  MUX21X1_HVT U458 ( .A1(n328), .A2(n442), .S0(n446), .Y(n508) );
  MUX21X1_HVT U459 ( .A1(n330), .A2(n293), .S0(n369), .Y(n515) );
  MUX21X1_HVT U460 ( .A1(n325), .A2(n352), .S0(n211), .Y(n517) );
  XNOR2X1_HVT U461 ( .A1(n461), .A2(n240), .Y(n414) );
  MUX21X1_HVT U462 ( .A1(n326), .A2(n328), .S0(n420), .Y(n609) );
  NAND2X0_HVT U463 ( .A1(n252), .A2(n505), .Y(n709) );
  NAND2X0_HVT U464 ( .A1(n430), .A2(n252), .Y(n718) );
  AND2X1_HVT U465 ( .A1(n357), .A2(n377), .Y(n415) );
  NAND2X0_HVT U466 ( .A1(n238), .A2(n303), .Y(n717) );
  AND2X1_HVT U467 ( .A1(n436), .A2(n239), .Y(n416) );
  INVX1_HVT U468 ( .A(n453), .Y(n451) );
  NBUFFX2_HVT U469 ( .A(in[0]), .Y(n429) );
endmodule

