
module sbox_10 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n5, n9, n18, n19, n23, n35, n50, n114, n119, n210, n211, n212, n213,
         n216, n217, n218, n219, n221, n224, n226, n227, n229, n231, n232,
         n236, n238, n241, n242, n249, n252, n253, n258, n261, n264, n267,
         n272, n273, n274, n277, n278, n279, n280, n282, n283, n284, n289,
         n293, n297, n299, n301, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754;

  NAND2X0_HVT U4 ( .A1(n19), .A2(n752), .Y(n751) );
  NAND2X0_HVT U5 ( .A1(n490), .A2(n481), .Y(n750) );
  NAND2X0_HVT U13 ( .A1(n743), .A2(n488), .Y(n744) );
  NAND2X0_HVT U15 ( .A1(n752), .A2(n477), .Y(n741) );
  NAND2X0_HVT U21 ( .A1(n19), .A2(n412), .Y(n737) );
  NAND2X0_HVT U33 ( .A1(n523), .A2(n410), .Y(n726) );
  NAND2X0_HVT U35 ( .A1(n479), .A2(n410), .Y(n725) );
  NAND2X0_HVT U42 ( .A1(n489), .A2(n414), .Y(n718) );
  NAND2X0_HVT U53 ( .A1(n707), .A2(n717), .Y(n708) );
  NAND2X0_HVT U56 ( .A1(n19), .A2(n703), .Y(n704) );
  MUX41X1_HVT U57 ( .A1(n18), .A3(n739), .A2(n704), .A4(n746), .S0(n447), .S1(
        n469), .Y(n702) );
  MUX41X1_HVT U61 ( .A1(n453), .A3(n391), .A2(n515), .A4(n475), .S0(n447), 
        .S1(n469), .Y(n698) );
  NAND2X0_HVT U62 ( .A1(n412), .A2(n361), .Y(n697) );
  AO21X1_HVT U66 ( .A1(n338), .A2(n470), .A3(n542), .Y(n693) );
  NAND2X0_HVT U73 ( .A1(n389), .A2(n686), .Y(n687) );
  MUX41X1_HVT U75 ( .A1(n539), .A3(n536), .A2(n365), .A4(n504), .S0(n349), 
        .S1(n500), .Y(n684) );
  MUX41X1_HVT U77 ( .A1(n114), .A3(n524), .A2(n683), .A4(n437), .S0(n471), 
        .S1(n495), .Y(n682) );
  AND2X1_HVT U83 ( .A1(n394), .A2(n423), .Y(n675) );
  MUX41X1_HVT U84 ( .A1(n5), .A3(n427), .A2(n740), .A4(n675), .S0(n465), .S1(
        n501), .Y(n674) );
  NAND2X0_HVT U85 ( .A1(n410), .A2(n387), .Y(n673) );
  MUX41X1_HVT U90 ( .A1(n714), .A3(n718), .A2(n508), .A4(n670), .S0(n349), 
        .S1(n499), .Y(n669) );
  AO21X1_HVT U93 ( .A1(n472), .A2(n665), .A3(n535), .Y(n666) );
  MUX41X1_HVT U97 ( .A1(n539), .A3(n452), .A2(n336), .A4(n741), .S0(n349), 
        .S1(n390), .Y(n661) );
  MUX41X1_HVT U98 ( .A1(n661), .A3(n664), .A2(n662), .A4(n669), .S0(n473), 
        .S1(n468), .Y(n660) );
  NAND2X0_HVT U101 ( .A1(n656), .A2(n655), .Y(n657) );
  MUX41X1_HVT U103 ( .A1(n752), .A3(n312), .A2(n422), .A4(n725), .S0(n430), 
        .S1(n390), .Y(n653) );
  MUX41X1_HVT U105 ( .A1(n534), .A3(n712), .A2(n652), .A4(n526), .S0(n465), 
        .S1(n500), .Y(n651) );
  NAND2X0_HVT U110 ( .A1(n361), .A2(n647), .Y(n648) );
  AND2X1_HVT U115 ( .A1(n341), .A2(n475), .Y(n643) );
  NAND2X0_HVT U123 ( .A1(n634), .A2(n633), .Y(n635) );
  MUX41X1_HVT U125 ( .A1(n737), .A3(n456), .A2(n514), .A4(n416), .S0(n465), 
        .S1(n446), .Y(n631) );
  AND2X1_HVT U140 ( .A1(n389), .A2(n392), .Y(n617) );
  MUX41X1_HVT U141 ( .A1(n734), .A3(n521), .A2(n617), .A4(n519), .S0(n350), 
        .S1(n445), .Y(n616) );
  MUX41X1_HVT U142 ( .A1(n5), .A3(n475), .A2(n525), .A4(n389), .S0(n349), .S1(
        n445), .Y(n615) );
  AND2X1_HVT U154 ( .A1(n472), .A2(n339), .Y(n604) );
  NAND2X0_HVT U158 ( .A1(n489), .A2(n387), .Y(n600) );
  MUX41X1_HVT U159 ( .A1(n744), .A3(n475), .A2(n600), .A4(n543), .S0(n494), 
        .S1(n348), .Y(n599) );
  AND2X1_HVT U162 ( .A1(n427), .A2(n686), .Y(n596) );
  NAND2X0_HVT U167 ( .A1(n365), .A2(n410), .Y(n591) );
  NAND2X0_HVT U174 ( .A1(n749), .A2(n490), .Y(n743) );
  MUX41X1_HVT U176 ( .A1(n479), .A3(n585), .A2(n516), .A4(n743), .S0(n447), 
        .S1(n350), .Y(n584) );
  NAND2X0_HVT U177 ( .A1(n489), .A2(n478), .Y(n583) );
  MUX41X1_HVT U180 ( .A1(n513), .A3(n114), .A2(n216), .A4(n448), .S0(n471), 
        .S1(n407), .Y(n580) );
  MUX41X1_HVT U182 ( .A1(n522), .A3(n19), .A2(n509), .A4(n529), .S0(n446), 
        .S1(n495), .Y(n578) );
  MUX41X1_HVT U189 ( .A1(n572), .A3(n355), .A2(n573), .A4(n526), .S0(n471), 
        .S1(n407), .Y(n571) );
  AO21X1_HVT U197 ( .A1(n451), .A2(n500), .A3(n535), .Y(n564) );
  MUX41X1_HVT U205 ( .A1(n423), .A3(n752), .A2(n532), .A4(n540), .S0(n350), 
        .S1(n348), .Y(n556) );
  NAND2X0_HVT U208 ( .A1(n249), .A2(n485), .Y(n647) );
  NAND2X0_HVT U212 ( .A1(n490), .A2(n483), .Y(n703) );
  NAND2X0_HVT U214 ( .A1(n345), .A2(n410), .Y(n554) );
  NAND2X0_HVT U215 ( .A1(n647), .A2(n484), .Y(n553) );
  NAND2X0_HVT U218 ( .A1(n537), .A2(n418), .Y(n607) );
  NAND2X0_HVT U220 ( .A1(n471), .A2(n554), .Y(n678) );
  INVX0_HVT U242 ( .A(n718), .Y(n545) );
  INVX0_HVT U245 ( .A(n750), .Y(n543) );
  INVX0_HVT U256 ( .A(n607), .Y(n535) );
  INVX0_HVT U259 ( .A(n729), .Y(n533) );
  INVX0_HVT U262 ( .A(n547), .Y(n532) );
  INVX0_HVT U264 ( .A(n725), .Y(n530) );
  INVX0_HVT U265 ( .A(n733), .Y(n529) );
  INVX0_HVT U268 ( .A(n737), .Y(n527) );
  INVX0_HVT U270 ( .A(n553), .Y(n526) );
  INVX0_HVT U271 ( .A(n647), .Y(n525) );
  INVX0_HVT U277 ( .A(n722), .Y(n521) );
  INVX0_HVT U278 ( .A(n726), .Y(n520) );
  INVX0_HVT U284 ( .A(n554), .Y(n517) );
  INVX0_HVT U289 ( .A(n655), .Y(n516) );
  INVX0_HVT U295 ( .A(n751), .Y(n513) );
  INVX0_HVT U296 ( .A(n741), .Y(n512) );
  INVX0_HVT U302 ( .A(n552), .Y(n508) );
  INVX0_HVT U306 ( .A(n591), .Y(n505) );
  MUX21X1_HVT U1 ( .A1(n479), .A2(n487), .S0(n418), .Y(n340) );
  MUX21X1_HVT U2 ( .A1(n486), .A2(n483), .S0(n336), .Y(n728) );
  NAND2X0_HVT U3 ( .A1(n491), .A2(n486), .Y(n686) );
  MUX21X1_HVT U6 ( .A1(n438), .A2(n444), .S0(n394), .Y(n437) );
  XOR2X1_HVT U7 ( .A1(n732), .A2(n404), .Y(n716) );
  MUX21X1_HVT U8 ( .A1(n340), .A2(n752), .S0(n494), .Y(n649) );
  MUX21X1_HVT U9 ( .A1(n728), .A2(n648), .S0(n350), .Y(n646) );
  INVX1_HVT U10 ( .A(n548), .Y(n507) );
  OA21X1_HVT U11 ( .A1(n505), .A2(n419), .A3(n728), .Y(n613) );
  INVX1_HVT U12 ( .A(n482), .Y(n537) );
  MUX21X1_HVT U14 ( .A1(n417), .A2(n388), .S0(n249), .Y(n307) );
  INVX1_HVT U16 ( .A(n719), .Y(n509) );
  XOR2X1_HVT U17 ( .A1(n362), .A2(n490), .Y(n711) );
  MUX21X1_HVT U18 ( .A1(n484), .A2(n479), .S0(n418), .Y(n688) );
  INVX1_HVT U19 ( .A(n469), .Y(n35) );
  MUX21X1_HVT U20 ( .A1(n680), .A2(n679), .S0(n467), .Y(n677) );
  OA21X1_HVT U22 ( .A1(n454), .A2(n419), .A3(n728), .Y(n588) );
  AND2X1_HVT U23 ( .A1(n353), .A2(n354), .Y(n5) );
  INVX0_HVT U24 ( .A(n753), .Y(n506) );
  INVX1_HVT U25 ( .A(in[0]), .Y(n23) );
  AND2X1_HVT U26 ( .A1(n370), .A2(n371), .Y(n9) );
  AND2X1_HVT U27 ( .A1(n355), .A2(n385), .Y(n18) );
  INVX1_HVT U28 ( .A(n236), .Y(n752) );
  MUX21X1_HVT U29 ( .A1(n478), .A2(n480), .S0(n229), .Y(n569) );
  INVX1_HVT U30 ( .A(n459), .Y(n361) );
  MUX21X2_HVT U31 ( .A1(n673), .A2(n339), .S0(n445), .Y(n577) );
  INVX1_HVT U32 ( .A(n393), .Y(n401) );
  MUX41X1_HVT U34 ( .A1(n451), .A3(n536), .A2(n449), .A4(n673), .S0(n404), 
        .S1(n119), .Y(n672) );
  MUX21X2_HVT U36 ( .A1(n476), .A2(n541), .S0(n336), .Y(n748) );
  INVX1_HVT U37 ( .A(n388), .Y(n389) );
  MUX41X1_HVT U38 ( .A1(n719), .A3(n732), .A2(n375), .A4(n389), .S0(n446), 
        .S1(n467), .Y(n567) );
  MUX21X2_HVT U39 ( .A1(n361), .A2(n476), .S0(n401), .Y(n719) );
  MUX21X1_HVT U40 ( .A1(n311), .A2(n426), .S0(n319), .Y(n375) );
  INVX1_HVT U41 ( .A(n372), .Y(n19) );
  INVX1_HVT U43 ( .A(n372), .Y(n386) );
  INVX0_HVT U44 ( .A(n727), .Y(n519) );
  MUX41X1_HVT U45 ( .A1(n689), .A3(n684), .A2(n685), .A4(n682), .S0(n23), .S1(
        n35), .Y(n681) );
  INVX1_HVT U46 ( .A(n325), .Y(n392) );
  INVX1_HVT U47 ( .A(n735), .Y(n546) );
  AO21X1_HVT U48 ( .A1(n467), .A2(n389), .A3(n427), .Y(n640) );
  INVX1_HVT U49 ( .A(n399), .Y(n400) );
  INVX1_HVT U50 ( .A(n400), .Y(n499) );
  NBUFFX2_HVT U51 ( .A(n399), .Y(n472) );
  NBUFFX2_HVT U52 ( .A(n482), .Y(n484) );
  INVX1_HVT U54 ( .A(n466), .Y(n381) );
  INVX1_HVT U55 ( .A(n745), .Y(n528) );
  MUX21X1_HVT U58 ( .A1(n339), .A2(n487), .S0(n489), .Y(n338) );
  NAND2X0_HVT U59 ( .A1(n690), .A2(n430), .Y(n431) );
  MUX21X1_HVT U60 ( .A1(n667), .A2(n666), .S0(n420), .Y(n664) );
  INVX1_HVT U63 ( .A(n703), .Y(n539) );
  INVX1_HVT U64 ( .A(n393), .Y(n337) );
  INVX1_HVT U65 ( .A(n344), .Y(n345) );
  INVX1_HVT U67 ( .A(n393), .Y(n489) );
  INVX1_HVT U68 ( .A(n380), .Y(n238) );
  INVX1_HVT U69 ( .A(n386), .Y(n523) );
  INVX1_HVT U70 ( .A(n447), .Y(n436) );
  INVX1_HVT U71 ( .A(n466), .Y(n366) );
  INVX1_HVT U72 ( .A(n465), .Y(n322) );
  INVX1_HVT U74 ( .A(n400), .Y(n500) );
  INVX1_HVT U76 ( .A(n346), .Y(n119) );
  INVX1_HVT U78 ( .A(n350), .Y(n346) );
  INVX1_HVT U79 ( .A(n349), .Y(n420) );
  NAND2X0_HVT U80 ( .A1(n641), .A2(n348), .Y(n313) );
  NOR3X0_HVT U81 ( .A1(n346), .A2(n369), .A3(n478), .Y(n628) );
  MUX21X1_HVT U82 ( .A1(n522), .A2(n736), .S0(n404), .Y(n620) );
  INVX1_HVT U86 ( .A(n496), .Y(n494) );
  INVX1_HVT U87 ( .A(n400), .Y(n348) );
  MUX21X1_HVT U88 ( .A1(n608), .A2(n609), .S0(n467), .Y(n606) );
  MUX21X1_HVT U89 ( .A1(n437), .A2(n537), .S0(n447), .Y(n609) );
  MUX21X1_HVT U91 ( .A1(n589), .A2(n588), .S0(n430), .Y(n587) );
  INVX0_HVT U92 ( .A(n337), .Y(n280) );
  INVX1_HVT U94 ( .A(n401), .Y(n380) );
  INVX1_HVT U95 ( .A(n496), .Y(n495) );
  INVX0_HVT U96 ( .A(n392), .Y(n418) );
  INVX1_HVT U99 ( .A(n249), .Y(n347) );
  INVX0_HVT U100 ( .A(in[1]), .Y(n493) );
  INVX1_HVT U102 ( .A(n493), .Y(n325) );
  INVX0_HVT U104 ( .A(n497), .Y(n252) );
  NBUFFX2_HVT U106 ( .A(n497), .Y(n469) );
  INVX1_HVT U107 ( .A(n447), .Y(n421) );
  INVX0_HVT U108 ( .A(n229), .Y(n491) );
  INVX0_HVT U109 ( .A(n470), .Y(n326) );
  INVX0_HVT U111 ( .A(n491), .Y(n415) );
  AND2X1_HVT U112 ( .A1(n289), .A2(n293), .Y(n50) );
  INVX1_HVT U113 ( .A(n506), .Y(n363) );
  INVX0_HVT U114 ( .A(n734), .Y(n504) );
  INVX0_HVT U116 ( .A(n742), .Y(n511) );
  MUX21X1_HVT U117 ( .A1(n364), .A2(n483), .S0(n418), .Y(n742) );
  INVX0_HVT U118 ( .A(n445), .Y(n318) );
  NBUFFX2_HVT U119 ( .A(n386), .Y(n485) );
  INVX0_HVT U120 ( .A(n472), .Y(n404) );
  NAND2X0_HVT U121 ( .A1(n320), .A2(n321), .Y(n114) );
  INVX1_HVT U122 ( .A(n488), .Y(n387) );
  INVX1_HVT U124 ( .A(n728), .Y(n540) );
  AND2X1_HVT U126 ( .A1(n241), .A2(n242), .Y(n210) );
  MUX21X1_HVT U127 ( .A1(n311), .A2(n426), .S0(n347), .Y(n211) );
  MUX41X1_HVT U128 ( .A1(n578), .A3(n575), .A2(n574), .A4(n571), .S0(n326), 
        .S1(n23), .Y(n570) );
  INVX1_HVT U129 ( .A(n388), .Y(n311) );
  INVX1_HVT U130 ( .A(n392), .Y(n341) );
  MUX21X1_HVT U131 ( .A1(n19), .A2(n480), .S0(n394), .Y(n745) );
  INVX1_HVT U132 ( .A(n531), .Y(n212) );
  INVX1_HVT U133 ( .A(n212), .Y(n213) );
  INVX0_HVT U134 ( .A(n518), .Y(n216) );
  MUX41X1_HVT U135 ( .A1(n619), .A3(n622), .A2(n621), .A4(n623), .S0(n473), 
        .S1(n468), .Y(n618) );
  NBUFFX2_HVT U136 ( .A(n487), .Y(n217) );
  MUX21X1_HVT U137 ( .A1(n312), .A2(n537), .S0(n497), .Y(n692) );
  INVX1_HVT U138 ( .A(n721), .Y(n522) );
  INVX1_HVT U139 ( .A(n550), .Y(n536) );
  OAI21X1_HVT U143 ( .A1(n434), .A2(n496), .A3(n50), .Y(n464) );
  INVX0_HVT U144 ( .A(n340), .Y(n724) );
  MUX41X1_HVT U145 ( .A1(n584), .A3(n581), .A2(n582), .A4(n580), .S0(n23), 
        .S1(n252), .Y(n579) );
  MUX41X1_HVT U146 ( .A1(n744), .A3(n704), .A2(n736), .A4(n413), .S0(n308), 
        .S1(n499), .Y(n557) );
  NAND2X0_HVT U147 ( .A1(n305), .A2(n410), .Y(n218) );
  NAND2X0_HVT U148 ( .A1(n365), .A2(n337), .Y(n219) );
  NAND2X0_HVT U149 ( .A1(n218), .A2(n219), .Y(n734) );
  MUX41X1_HVT U150 ( .A1(n510), .A3(n715), .A2(n742), .A4(n546), .S0(n420), 
        .S1(n499), .Y(n676) );
  NAND2X0_HVT U151 ( .A1(n729), .A2(n407), .Y(n221) );
  NAND2X0_HVT U152 ( .A1(n534), .A2(n366), .Y(n224) );
  NAND2X0_HVT U153 ( .A1(n221), .A2(n224), .Y(n629) );
  INVX0_HVT U155 ( .A(n731), .Y(n534) );
  MUX21X2_HVT U156 ( .A1(n576), .A2(n577), .S0(n466), .Y(n575) );
  INVX0_HVT U157 ( .A(n749), .Y(n426) );
  MUX21X1_HVT U160 ( .A1(n417), .A2(n486), .S0(n229), .Y(n731) );
  NBUFFX2_HVT U161 ( .A(n495), .Y(n467) );
  INVX0_HVT U163 ( .A(n753), .Y(n365) );
  INVX1_HVT U164 ( .A(n744), .Y(n518) );
  MUX41X1_HVT U165 ( .A1(n692), .A3(n694), .A2(n514), .A4(n693), .S0(n333), 
        .S1(n419), .Y(n691) );
  INVX0_HVT U166 ( .A(n455), .Y(n358) );
  NBUFFX2_HVT U168 ( .A(n747), .Y(n482) );
  INVX0_HVT U169 ( .A(n491), .Y(n319) );
  NAND2X0_HVT U170 ( .A1(n365), .A2(n347), .Y(n226) );
  NAND2X0_HVT U171 ( .A1(n541), .A2(n341), .Y(n227) );
  NAND2X0_HVT U172 ( .A1(n226), .A2(n227), .Y(n732) );
  INVX0_HVT U173 ( .A(n486), .Y(n541) );
  INVX1_HVT U175 ( .A(n325), .Y(n229) );
  MUX41X1_HVT U178 ( .A1(n629), .A3(n628), .A2(n627), .A4(n626), .S0(n404), 
        .S1(n252), .Y(n625) );
  NBUFFX2_HVT U179 ( .A(n501), .Y(n446) );
  NAND2X0_HVT U181 ( .A1(n519), .A2(n407), .Y(n408) );
  MUX21X1_HVT U183 ( .A1(n448), .A2(n740), .S0(n419), .Y(n561) );
  NAND2X0_HVT U184 ( .A1(n702), .A2(n430), .Y(n231) );
  NAND2X0_HVT U185 ( .A1(n700), .A2(n433), .Y(n232) );
  NAND2X0_HVT U186 ( .A1(n231), .A2(n232), .Y(n699) );
  INVX0_HVT U187 ( .A(in[1]), .Y(n393) );
  OR2X1_HVT U188 ( .A1(n306), .A2(n474), .Y(n267) );
  MUX41X1_HVT U190 ( .A1(n558), .A3(n559), .A2(n556), .A4(n557), .S0(n470), 
        .S1(n23), .Y(n555) );
  INVX0_HVT U191 ( .A(n338), .Y(n746) );
  XOR2X1_HVT U192 ( .A1(n319), .A2(n311), .Y(n715) );
  INVX1_HVT U193 ( .A(n531), .Y(n317) );
  AND2X1_HVT U194 ( .A1(n401), .A2(n362), .Y(n236) );
  INVX0_HVT U195 ( .A(n665), .Y(n524) );
  NAND2X0_HVT U196 ( .A1(n414), .A2(n337), .Y(n241) );
  NAND2X0_HVT U198 ( .A1(n488), .A2(n415), .Y(n242) );
  NAND2X0_HVT U199 ( .A1(n242), .A2(n241), .Y(n413) );
  MUX21X1_HVT U200 ( .A1(n481), .A2(n364), .S0(n412), .Y(n411) );
  NAND2X0_HVT U201 ( .A1(n379), .A2(n415), .Y(n735) );
  INVX0_HVT U202 ( .A(n394), .Y(n412) );
  MUX21X1_HVT U203 ( .A1(n365), .A2(n537), .S0(n280), .Y(n594) );
  MUX41X1_HVT U204 ( .A1(n594), .A3(n714), .A2(n533), .A4(n737), .S0(n318), 
        .S1(n433), .Y(n593) );
  NBUFFX2_HVT U206 ( .A(n501), .Y(n390) );
  INVX1_HVT U207 ( .A(n502), .Y(n501) );
  NBUFFX2_HVT U209 ( .A(n325), .Y(n249) );
  MUX41X1_HVT U210 ( .A1(n644), .A3(n638), .A2(n630), .A4(n625), .S0(n23), 
        .S1(n439), .Y(out[3]) );
  MUX21X1_HVT U211 ( .A1(n541), .A2(n523), .S0(n341), .Y(n722) );
  MUX41X1_HVT U213 ( .A1(n688), .A3(n687), .A2(n733), .A4(n735), .S0(n348), 
        .S1(n467), .Y(n685) );
  NAND2X0_HVT U216 ( .A1(n706), .A2(n322), .Y(n253) );
  NAND2X0_HVT U217 ( .A1(n710), .A2(n333), .Y(n258) );
  NAND2X0_HVT U219 ( .A1(n253), .A2(n258), .Y(n705) );
  INVX0_HVT U221 ( .A(n393), .Y(n490) );
  INVX1_HVT U222 ( .A(n393), .Y(n336) );
  MUX21X1_HVT U223 ( .A1(n545), .A2(n9), .S0(n501), .Y(n565) );
  NAND2X0_HVT U224 ( .A1(n264), .A2(n267), .Y(n261) );
  INVX0_HVT U225 ( .A(n344), .Y(n305) );
  INVX1_HVT U226 ( .A(n478), .Y(n417) );
  INVX0_HVT U227 ( .A(n740), .Y(n515) );
  INVX0_HVT U228 ( .A(in[5]), .Y(n498) );
  MUX21X1_HVT U229 ( .A1(n752), .A2(n392), .S0(n466), .Y(n633) );
  INVX1_HVT U230 ( .A(n749), .Y(n344) );
  MUX21X1_HVT U231 ( .A1(n477), .A2(n523), .S0(n249), .Y(n663) );
  INVX0_HVT U232 ( .A(n307), .Y(n391) );
  INVX0_HVT U233 ( .A(n480), .Y(n438) );
  MUX41X1_HVT U234 ( .A1(n583), .A3(n307), .A2(n722), .A4(n9), .S0(n420), .S1(
        n390), .Y(n582) );
  INVX0_HVT U235 ( .A(n480), .Y(n414) );
  INVX1_HVT U236 ( .A(in[4]), .Y(n531) );
  NAND2X0_HVT U237 ( .A1(n306), .A2(n474), .Y(n264) );
  NAND2X0_HVT U238 ( .A1(n264), .A2(n267), .Y(n444) );
  INVX0_HVT U239 ( .A(n444), .Y(n749) );
  NAND2X0_HVT U240 ( .A1(n476), .A2(n418), .Y(n272) );
  NAND2X0_HVT U241 ( .A1(n435), .A2(n392), .Y(n273) );
  NAND2X0_HVT U243 ( .A1(n272), .A2(n273), .Y(n434) );
  NBUFFX2_HVT U244 ( .A(n261), .Y(n476) );
  INVX0_HVT U246 ( .A(in[3]), .Y(n544) );
  INVX0_HVT U247 ( .A(n394), .Y(n410) );
  INVX0_HVT U248 ( .A(n461), .Y(n644) );
  INVX0_HVT U249 ( .A(n434), .Y(n723) );
  INVX0_HVT U250 ( .A(n482), .Y(n388) );
  INVX1_HVT U251 ( .A(in[2]), .Y(n496) );
  NAND2X0_HVT U252 ( .A1(n478), .A2(n337), .Y(n274) );
  NAND2X0_HVT U253 ( .A1(n475), .A2(n280), .Y(n277) );
  NAND2X0_HVT U254 ( .A1(n274), .A2(n277), .Y(n655) );
  NAND2X0_HVT U255 ( .A1(n650), .A2(n439), .Y(n278) );
  NAND2X0_HVT U257 ( .A1(n660), .A2(n304), .Y(n279) );
  NAND2X0_HVT U258 ( .A1(n278), .A2(n279), .Y(out[2]) );
  INVX1_HVT U260 ( .A(n229), .Y(n492) );
  NAND2X0_HVT U261 ( .A1(n453), .A2(n282), .Y(n283) );
  NAND2X0_HVT U263 ( .A1(n659), .A2(n713), .Y(n284) );
  NAND2X0_HVT U266 ( .A1(n283), .A2(n284), .Y(n658) );
  INVX0_HVT U267 ( .A(n713), .Y(n282) );
  MUX41X1_HVT U269 ( .A1(n452), .A3(n546), .A2(n663), .A4(n538), .S0(n420), 
        .S1(n500), .Y(n662) );
  NAND2X0_HVT U272 ( .A1(n537), .A2(n280), .Y(n289) );
  NAND2X0_HVT U273 ( .A1(n523), .A2(n336), .Y(n293) );
  NAND2X0_HVT U274 ( .A1(n696), .A2(n322), .Y(n297) );
  NAND2X0_HVT U275 ( .A1(n698), .A2(n430), .Y(n299) );
  NAND2X0_HVT U276 ( .A1(n297), .A2(n299), .Y(n695) );
  INVX1_HVT U279 ( .A(n380), .Y(n369) );
  MUX21X1_HVT U280 ( .A1(n657), .A2(n503), .S0(n333), .Y(n654) );
  NAND2X0_HVT U281 ( .A1(n345), .A2(n280), .Y(n301) );
  NAND2X0_HVT U282 ( .A1(n479), .A2(n401), .Y(n303) );
  NAND2X0_HVT U283 ( .A1(n301), .A2(n303), .Y(n683) );
  INVX1_HVT U285 ( .A(n551), .Y(n538) );
  INVX1_HVT U286 ( .A(n439), .Y(n304) );
  INVX1_HVT U287 ( .A(in[6]), .Y(n439) );
  NAND2X0_HVT U288 ( .A1(n488), .A2(n703), .Y(n592) );
  NBUFFX2_HVT U290 ( .A(in[3]), .Y(n474) );
  INVX1_HVT U291 ( .A(n317), .Y(n306) );
  MUX21X1_HVT U292 ( .A1(n729), .A2(n553), .S0(n499), .Y(n549) );
  MUX21X1_HVT U293 ( .A1(n488), .A2(n19), .S0(n415), .Y(n665) );
  OR2X1_HVT U294 ( .A1(n387), .A2(n236), .Y(n701) );
  INVX0_HVT U297 ( .A(n481), .Y(n379) );
  INVX0_HVT U298 ( .A(n481), .Y(n339) );
  INVX0_HVT U299 ( .A(n411), .Y(n739) );
  INVX1_HVT U300 ( .A(n493), .Y(n394) );
  NAND2X0_HVT U301 ( .A1(n450), .A2(n308), .Y(n309) );
  NAND2X0_HVT U303 ( .A1(n515), .A2(n349), .Y(n310) );
  NAND2X0_HVT U304 ( .A1(n309), .A2(n310), .Y(n627) );
  INVX0_HVT U305 ( .A(n349), .Y(n308) );
  XNOR2X1_HVT U307 ( .A1(n485), .A2(n249), .Y(n450) );
  AND2X1_HVT U308 ( .A1(n320), .A2(n321), .Y(n312) );
  INVX1_HVT U309 ( .A(n426), .Y(n427) );
  NAND2X0_HVT U310 ( .A1(n640), .A2(n318), .Y(n314) );
  NAND2X0_HVT U311 ( .A1(n313), .A2(n314), .Y(n639) );
  NAND2X0_HVT U312 ( .A1(n642), .A2(n468), .Y(n315) );
  NAND2X0_HVT U313 ( .A1(n639), .A2(n326), .Y(n316) );
  NAND2X0_HVT U314 ( .A1(n315), .A2(n316), .Y(n638) );
  MUX21X1_HVT U315 ( .A1(n530), .A2(n413), .S0(n465), .Y(n641) );
  OA21X1_HVT U316 ( .A1(n748), .A2(n421), .A3(n521), .Y(n560) );
  MUX41X1_HVT U317 ( .A1(n728), .A3(n504), .A2(n643), .A4(n744), .S0(n420), 
        .S1(n421), .Y(n642) );
  MUX41X1_HVT U318 ( .A1(n676), .A3(n677), .A2(n672), .A4(n674), .S0(n468), 
        .S1(n23), .Y(n671) );
  INVX0_HVT U319 ( .A(n422), .Y(n730) );
  MUX41X1_HVT U320 ( .A1(n537), .A3(n732), .A2(n211), .A4(n750), .S0(n501), 
        .S1(n381), .Y(n622) );
  MUX21X1_HVT U321 ( .A1(n523), .A2(n423), .S0(n394), .Y(n727) );
  NAND2X0_HVT U322 ( .A1(n485), .A2(n319), .Y(n320) );
  NAND2X0_HVT U323 ( .A1(n379), .A2(n238), .Y(n321) );
  NBUFFX2_HVT U324 ( .A(n261), .Y(n477) );
  MUX41X1_HVT U325 ( .A1(n538), .A3(n427), .A2(n723), .A4(n488), .S0(n322), 
        .S1(n390), .Y(n566) );
  NAND2X0_HVT U326 ( .A1(n598), .A2(n304), .Y(n323) );
  NAND2X0_HVT U327 ( .A1(n586), .A2(n439), .Y(n324) );
  NAND2X0_HVT U328 ( .A1(n324), .A2(n323), .Y(out[5]) );
  INVX1_HVT U329 ( .A(n459), .Y(n362) );
  MUX21X1_HVT U330 ( .A1(n541), .A2(n477), .S0(n492), .Y(n597) );
  NBUFFX2_HVT U331 ( .A(n399), .Y(n471) );
  NAND2X0_HVT U332 ( .A1(n570), .A2(n439), .Y(n327) );
  NAND2X0_HVT U333 ( .A1(n579), .A2(n304), .Y(n328) );
  NAND2X0_HVT U334 ( .A1(n327), .A2(n328), .Y(out[6]) );
  MUX41X1_HVT U335 ( .A1(n596), .A3(n391), .A2(n597), .A4(n450), .S0(n366), 
        .S1(n348), .Y(n595) );
  MUX41X1_HVT U336 ( .A1(n727), .A3(n745), .A2(n378), .A4(n724), .S0(n308), 
        .S1(n436), .Y(n558) );
  INVX0_HVT U337 ( .A(n485), .Y(n435) );
  INVX0_HVT U338 ( .A(n466), .Y(n433) );
  NAND2X0_HVT U339 ( .A1(n560), .A2(n366), .Y(n329) );
  NAND2X0_HVT U340 ( .A1(n561), .A2(n466), .Y(n330) );
  NAND2X0_HVT U341 ( .A1(n329), .A2(n330), .Y(n559) );
  MUX41X1_HVT U342 ( .A1(n453), .A3(n648), .A2(n530), .A4(n363), .S0(n381), 
        .S1(n501), .Y(n605) );
  NAND2X0_HVT U343 ( .A1(n708), .A2(n318), .Y(n331) );
  NAND2X0_HVT U344 ( .A1(n709), .A2(n471), .Y(n332) );
  NAND2X0_HVT U345 ( .A1(n332), .A2(n331), .Y(n706) );
  NAND2X0_HVT U346 ( .A1(n624), .A2(n333), .Y(n334) );
  NAND2X0_HVT U347 ( .A1(n346), .A2(n503), .Y(n335) );
  NAND2X0_HVT U348 ( .A1(n334), .A2(n335), .Y(n623) );
  INVX0_HVT U349 ( .A(n366), .Y(n333) );
  XNOR2X2_HVT U350 ( .A1(n345), .A2(n347), .Y(n714) );
  MUX41X1_HVT U351 ( .A1(n449), .A3(n726), .A2(n507), .A4(n724), .S0(n465), 
        .S1(n446), .Y(n621) );
  INVX0_HVT U352 ( .A(n378), .Y(n720) );
  MUX41X1_HVT U353 ( .A1(n593), .A3(n587), .A2(n595), .A4(n590), .S0(n23), 
        .S1(n468), .Y(n586) );
  MUX41X1_HVT U354 ( .A1(n612), .A3(n611), .A2(n616), .A4(n615), .S0(n326), 
        .S1(n473), .Y(n610) );
  NAND2X0_HVT U355 ( .A1(n730), .A2(n404), .Y(n342) );
  NAND2X0_HVT U356 ( .A1(n236), .A2(n472), .Y(n343) );
  NAND2X0_HVT U357 ( .A1(n342), .A2(n343), .Y(n614) );
  MUX21X1_HVT U358 ( .A1(n614), .A2(n613), .S0(n407), .Y(n612) );
  INVX0_HVT U359 ( .A(n748), .Y(n514) );
  NBUFFX2_HVT U360 ( .A(n497), .Y(n470) );
  MUX41X1_HVT U361 ( .A1(n691), .A3(n699), .A2(n695), .A4(n705), .S0(n304), 
        .S1(n473), .Y(out[0]) );
  MUX41X1_HVT U362 ( .A1(n411), .A3(n510), .A2(n508), .A4(n527), .S0(n446), 
        .S1(n252), .Y(n710) );
  NBUFFX2_HVT U363 ( .A(n213), .Y(n479) );
  INVX1_HVT U364 ( .A(n479), .Y(n423) );
  MUX41X1_HVT U365 ( .A1(n721), .A3(n714), .A2(n452), .A4(n686), .S0(n500), 
        .S1(n322), .Y(n574) );
  MUX41X1_HVT U366 ( .A1(n697), .A3(n512), .A2(n518), .A4(n511), .S0(n446), 
        .S1(n469), .Y(n696) );
  NBUFFX2_HVT U367 ( .A(n494), .Y(n349) );
  NBUFFX2_HVT U368 ( .A(n494), .Y(n350) );
  NBUFFX2_HVT U369 ( .A(n494), .Y(n465) );
  INVX1_HVT U370 ( .A(in[7]), .Y(n502) );
  NAND2X0_HVT U371 ( .A1(n751), .A2(n465), .Y(n351) );
  NAND2X0_HVT U372 ( .A1(n620), .A2(n420), .Y(n352) );
  NAND2X0_HVT U373 ( .A1(n351), .A2(n352), .Y(n619) );
  NAND2X0_HVT U374 ( .A1(n414), .A2(n491), .Y(n353) );
  NAND2X0_HVT U375 ( .A1(n476), .A2(n347), .Y(n354) );
  NAND2X0_HVT U376 ( .A1(n353), .A2(n354), .Y(n736) );
  MUX41X1_HVT U377 ( .A1(n18), .A3(n389), .A2(n591), .A4(n592), .S0(n407), 
        .S1(n348), .Y(n590) );
  NAND2X0_HVT U378 ( .A1(n427), .A2(n492), .Y(n355) );
  NAND2X0_HVT U379 ( .A1(n414), .A2(n318), .Y(n356) );
  NAND2X0_HVT U380 ( .A1(n479), .A2(n472), .Y(n357) );
  NAND2X0_HVT U381 ( .A1(n356), .A2(n357), .Y(n668) );
  NAND2X0_HVT U382 ( .A1(n361), .A2(n358), .Y(n359) );
  NAND2X0_HVT U383 ( .A1(n668), .A2(n455), .Y(n360) );
  NAND2X0_HVT U384 ( .A1(n359), .A2(n360), .Y(n667) );
  XNOR2X1_HVT U385 ( .A1(n400), .A2(n394), .Y(n455) );
  INVX0_HVT U386 ( .A(n506), .Y(n364) );
  INVX1_HVT U387 ( .A(n753), .Y(n459) );
  MUX41X1_HVT U388 ( .A1(n567), .A3(n563), .A2(n568), .A4(n566), .S0(n23), 
        .S1(n470), .Y(n562) );
  MUX41X1_HVT U389 ( .A1(n725), .A3(n718), .A2(n569), .A4(n711), .S0(n366), 
        .S1(n500), .Y(n568) );
  INVX0_HVT U390 ( .A(n686), .Y(n542) );
  NAND2X0_HVT U391 ( .A1(n564), .A2(n407), .Y(n367) );
  NAND2X0_HVT U392 ( .A1(n565), .A2(n381), .Y(n368) );
  NAND2X0_HVT U393 ( .A1(n367), .A2(n368), .Y(n563) );
  NAND2X0_HVT U394 ( .A1(n483), .A2(n369), .Y(n370) );
  NAND2X0_HVT U395 ( .A1(n423), .A2(n380), .Y(n371) );
  AND2X1_HVT U396 ( .A1(n213), .A2(n544), .Y(n372) );
  NAND2X0_HVT U397 ( .A1(n481), .A2(n491), .Y(n373) );
  NAND2X0_HVT U398 ( .A1(n477), .A2(n410), .Y(n374) );
  NAND2X0_HVT U399 ( .A1(n373), .A2(n374), .Y(n740) );
  NAND2X0_HVT U400 ( .A1(n480), .A2(n280), .Y(n376) );
  NAND2X0_HVT U401 ( .A1(n423), .A2(n401), .Y(n377) );
  NAND2X0_HVT U402 ( .A1(n376), .A2(n377), .Y(n729) );
  MUX21X1_HVT U403 ( .A1(n364), .A2(n379), .S0(n380), .Y(n378) );
  MUX21X1_HVT U404 ( .A1(n484), .A2(n416), .S0(n318), .Y(n624) );
  NAND2X0_HVT U405 ( .A1(n484), .A2(n447), .Y(n382) );
  NAND2X0_HVT U406 ( .A1(n738), .A2(n421), .Y(n383) );
  NAND2X0_HVT U407 ( .A1(n382), .A2(n383), .Y(n680) );
  NAND2X0_HVT U408 ( .A1(n364), .A2(n341), .Y(n384) );
  NAND2X0_HVT U409 ( .A1(n417), .A2(n415), .Y(n385) );
  NAND2X0_HVT U410 ( .A1(n384), .A2(n385), .Y(n738) );
  NBUFFX2_HVT U411 ( .A(n754), .Y(n487) );
  AO21X1_HVT U412 ( .A1(n392), .A2(n537), .A3(n421), .Y(n656) );
  NAND2X0_HVT U413 ( .A1(n604), .A2(n358), .Y(n395) );
  NAND2X0_HVT U414 ( .A1(n363), .A2(n455), .Y(n396) );
  NAND2X0_HVT U415 ( .A1(n395), .A2(n396), .Y(n603) );
  NAND2X0_HVT U416 ( .A1(n602), .A2(n346), .Y(n397) );
  NAND2X0_HVT U417 ( .A1(n603), .A2(n119), .Y(n398) );
  NAND2X0_HVT U418 ( .A1(n397), .A2(n398), .Y(n601) );
  MUX21X1_HVT U419 ( .A1(n722), .A2(n524), .S0(n471), .Y(n602) );
  INVX1_HVT U420 ( .A(n549), .Y(n503) );
  INVX1_HVT U421 ( .A(n502), .Y(n399) );
  INVX1_HVT U422 ( .A(n471), .Y(n419) );
  MUX21X1_HVT U423 ( .A1(n19), .A2(n417), .S0(n492), .Y(n416) );
  MUX41X1_HVT U424 ( .A1(n653), .A3(n658), .A2(n651), .A4(n654), .S0(n473), 
        .S1(n326), .Y(n650) );
  NAND2X0_HVT U425 ( .A1(n631), .A2(n326), .Y(n402) );
  NAND2X0_HVT U426 ( .A1(n632), .A2(n468), .Y(n403) );
  NAND2X0_HVT U427 ( .A1(n402), .A2(n403), .Y(n630) );
  MUX21X1_HVT U428 ( .A1(n365), .A2(n458), .S0(n460), .Y(n457) );
  INVX1_HVT U429 ( .A(n645), .Y(n458) );
  INVX0_HVT U430 ( .A(n738), .Y(n510) );
  NAND2X0_HVT U431 ( .A1(n429), .A2(n428), .Y(out[4]) );
  NAND2X0_HVT U432 ( .A1(n636), .A2(n436), .Y(n405) );
  NAND2X0_HVT U433 ( .A1(n635), .A2(n472), .Y(n406) );
  NAND2X0_HVT U434 ( .A1(n405), .A2(n406), .Y(n632) );
  MUX21X1_HVT U435 ( .A1(n520), .A2(n637), .S0(n349), .Y(n636) );
  NAND2X0_HVT U436 ( .A1(n307), .A2(n346), .Y(n409) );
  NAND2X0_HVT U437 ( .A1(n408), .A2(n409), .Y(n626) );
  INVX0_HVT U438 ( .A(n496), .Y(n407) );
  MUX41X1_HVT U439 ( .A1(n601), .A3(n606), .A2(n599), .A4(n605), .S0(n473), 
        .S1(n326), .Y(n598) );
  NBUFFX2_HVT U440 ( .A(n754), .Y(n488) );
  MUX41X1_HVT U441 ( .A1(n50), .A3(n454), .A2(n701), .A4(n456), .S0(n318), 
        .S1(n252), .Y(n700) );
  MUX21X1_HVT U442 ( .A1(n423), .A2(n386), .S0(n337), .Y(n422) );
  NAND2X0_HVT U443 ( .A1(n540), .A2(n322), .Y(n424) );
  NAND2X0_HVT U444 ( .A1(n742), .A2(n467), .Y(n425) );
  NAND2X0_HVT U445 ( .A1(n424), .A2(n425), .Y(n659) );
  AND3X1_HVT U446 ( .A1(n363), .A2(n703), .A3(n678), .Y(n679) );
  NAND2X0_HVT U447 ( .A1(n441), .A2(n440), .Y(out[1]) );
  OA21X1_HVT U448 ( .A1(n720), .A2(n421), .A3(n607), .Y(n608) );
  NAND2X0_HVT U449 ( .A1(n618), .A2(n304), .Y(n428) );
  NAND2X0_HVT U450 ( .A1(n610), .A2(n439), .Y(n429) );
  NAND2X0_HVT U451 ( .A1(n716), .A2(n433), .Y(n432) );
  NAND2X0_HVT U452 ( .A1(n431), .A2(n432), .Y(n689) );
  INVX1_HVT U453 ( .A(n433), .Y(n430) );
  OA21X1_HVT U454 ( .A1(n210), .A2(n421), .A3(n5), .Y(n576) );
  MUX41X1_HVT U455 ( .A1(n9), .A3(n517), .A2(n532), .A4(n731), .S0(n366), .S1(
        n436), .Y(n581) );
  MUX41X1_HVT U456 ( .A1(n714), .A3(n539), .A2(n686), .A4(n507), .S0(n381), 
        .S1(n436), .Y(n611) );
  NBUFFX2_HVT U457 ( .A(n476), .Y(n475) );
  NAND2X0_HVT U458 ( .A1(n671), .A2(n439), .Y(n440) );
  NAND2X0_HVT U459 ( .A1(n681), .A2(n304), .Y(n441) );
  NAND2X0_HVT U460 ( .A1(n555), .A2(n439), .Y(n442) );
  NAND2X0_HVT U461 ( .A1(n562), .A2(n304), .Y(n443) );
  NAND2X0_HVT U462 ( .A1(n442), .A2(n443), .Y(out[7]) );
  INVX1_HVT U463 ( .A(n646), .Y(n463) );
  INVX1_HVT U464 ( .A(n498), .Y(n497) );
  MUX41X1_HVT U465 ( .A1(n457), .A3(n462), .A2(n463), .A4(n464), .S0(n468), 
        .S1(n499), .Y(n461) );
  NBUFFX2_HVT U466 ( .A(n399), .Y(n445) );
  NBUFFX2_HVT U467 ( .A(n399), .Y(n447) );
  AND2X1_HVT U468 ( .A1(n477), .A2(n703), .Y(n448) );
  MUX21X1_HVT U469 ( .A1(n523), .A2(n387), .S0(n497), .Y(n707) );
  AND2X1_HVT U470 ( .A1(n363), .A2(n686), .Y(n449) );
  MUX21X1_HVT U471 ( .A1(n523), .A2(n365), .S0(n238), .Y(n585) );
  MUX21X1_HVT U472 ( .A1(n479), .A2(n480), .S0(n369), .Y(n637) );
  MUX21X1_HVT U473 ( .A1(n485), .A2(n484), .S0(n336), .Y(n670) );
  MUX21X1_HVT U474 ( .A1(n363), .A2(n485), .S0(n341), .Y(n548) );
  MUX21X1_HVT U475 ( .A1(n361), .A2(n478), .S0(n369), .Y(n552) );
  XNOR2X1_HVT U476 ( .A1(n487), .A2(n492), .Y(n451) );
  AND2X1_HVT U477 ( .A1(n401), .A2(n365), .Y(n452) );
  MUX21X1_HVT U478 ( .A1(n483), .A2(n481), .S0(n492), .Y(n551) );
  AND2X1_HVT U479 ( .A1(n217), .A2(n647), .Y(n453) );
  MUX21X1_HVT U480 ( .A1(n389), .A2(n217), .S0(n407), .Y(n634) );
  XOR2X1_HVT U481 ( .A1(n478), .A2(n337), .Y(n733) );
  NBUFFX2_HVT U482 ( .A(n544), .Y(n480) );
  NBUFFX2_HVT U483 ( .A(n544), .Y(n481) );
  NBUFFX2_HVT U484 ( .A(in[5]), .Y(n468) );
  MUX21X1_HVT U485 ( .A1(n484), .A2(n538), .S0(n472), .Y(n589) );
  XOR2X1_HVT U486 ( .A1(n341), .A2(n379), .Y(n712) );
  MUX21X1_HVT U487 ( .A1(n389), .A2(n426), .S0(n336), .Y(n652) );
  AND2X1_HVT U488 ( .A1(n477), .A2(n412), .Y(n454) );
  MUX21X1_HVT U489 ( .A1(n414), .A2(n523), .S0(n238), .Y(n721) );
  MUX21X1_HVT U490 ( .A1(n387), .A2(n538), .S0(n472), .Y(n690) );
  NAND2X0_HVT U491 ( .A1(n306), .A2(n474), .Y(n753) );
  INVX1_HVT U492 ( .A(n649), .Y(n462) );
  MUX21X1_HVT U493 ( .A1(n414), .A2(n725), .S0(n497), .Y(n709) );
  XOR2X1_HVT U494 ( .A1(n337), .A2(n470), .Y(n717) );
  NBUFFX2_HVT U495 ( .A(n754), .Y(n486) );
  MUX21X1_HVT U496 ( .A1(n379), .A2(n537), .S0(n489), .Y(n550) );
  MUX21X1_HVT U497 ( .A1(n528), .A2(n415), .S0(n497), .Y(n694) );
  NBUFFX2_HVT U498 ( .A(n747), .Y(n483) );
  NBUFFX2_HVT U499 ( .A(n531), .Y(n478) );
  AND2X1_HVT U500 ( .A1(n481), .A2(n280), .Y(n456) );
  MUX21X1_HVT U501 ( .A1(n480), .A2(n217), .S0(n341), .Y(n572) );
  MUX21X1_HVT U502 ( .A1(n487), .A2(n363), .S0(n490), .Y(n573) );
  NAND2X0_HVT U503 ( .A1(n474), .A2(n317), .Y(n754) );
  NAND2X0_HVT U504 ( .A1(n544), .A2(n317), .Y(n747) );
  MUX21X1_HVT U505 ( .A1(n417), .A2(n488), .S0(n489), .Y(n547) );
  MUX21X1_HVT U506 ( .A1(n438), .A2(n417), .S0(n494), .Y(n645) );
  NBUFFX2_HVT U507 ( .A(in[0]), .Y(n473) );
  NBUFFX2_HVT U508 ( .A(n495), .Y(n466) );
  XOR2X1_HVT U509 ( .A1(n490), .A2(n496), .Y(n460) );
  XOR2X1_HVT U510 ( .A1(n495), .A2(n445), .Y(n713) );
endmodule

