
module keygen_1 ( round_num, keyin, keyout );
  input [0:3] round_num;
  input [0:127] keyin;
  output [0:127] keyout;
  wire   n23, n49, n152, n211, n212, n213, n214, n217, n218, n219, n220, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n242, n243, n244,
         n245, n246, n247, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n293, n294, n295, n296, n297, n298, n300, n301, n302,
         n303, n304, n305, n328, n354, n457, n516, n517, n519, n522, n523,
         n524, n525, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n609, n610, n633, n659, n821, n822, n823, n824, n827,
         n828, n829, n830, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n938,
         n965, n1125, n1126, n1130, n1131, n1132, n1133, n1134, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1259, n1333,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700;
  wire   [0:31] dummy;

  NAND2X0_HVT U4 ( .A1(n1443), .A2(n1405), .Y(n2697) );
  NAND2X0_HVT U5 ( .A1(n1368), .A2(n1441), .Y(n2696) );
  NAND2X0_HVT U6 ( .A1(n1403), .A2(n2697), .Y(n2695) );
  NAND2X0_HVT U15 ( .A1(n2685), .A2(n1410), .Y(n2686) );
  NAND2X0_HVT U17 ( .A1(n2697), .A2(n273), .Y(n2683) );
  NAND2X0_HVT U21 ( .A1(n1402), .A2(n1446), .Y(n2679) );
  NAND2X0_HVT U25 ( .A1(n1368), .A2(n1446), .Y(n2676) );
  NAND2X0_HVT U33 ( .A1(n1446), .A2(n1674), .Y(n2668) );
  NAND2X0_HVT U34 ( .A1(n1670), .A2(n1446), .Y(n2667) );
  NAND2X0_HVT U39 ( .A1(n1440), .A2(n234), .Y(n2662) );
  MUX41X1_HVT U50 ( .A1(n1656), .A3(n1614), .A2(n2687), .A4(n1633), .S0(n1452), 
        .S1(n1239), .Y(n2652) );
  NAND2X0_HVT U52 ( .A1(n2649), .A2(n2659), .Y(n2650) );
  MUX41X1_HVT U55 ( .A1(n1189), .A3(n1632), .A2(n1631), .A4(n238), .S0(n517), 
        .S1(n1450), .Y(n2646) );
  NAND2X0_HVT U56 ( .A1(n1446), .A2(n1406), .Y(n2645) );
  MUX41X1_HVT U57 ( .A1(n2645), .A3(n1621), .A2(n1651), .A4(n1630), .S0(n870), 
        .S1(n1450), .Y(n2644) );
  NAND2X0_HVT U59 ( .A1(n1403), .A2(n2641), .Y(n2642) );
  MUX41X1_HVT U60 ( .A1(n1657), .A3(n1629), .A2(n2642), .A4(n2690), .S0(n1245), 
        .S1(n1450), .Y(n2640) );
  NAND2X0_HVT U61 ( .A1(n1410), .A2(n2697), .Y(n2639) );
  MUX41X1_HVT U62 ( .A1(n1217), .A3(n2639), .A2(n1214), .A4(n1628), .S0(n1452), 
        .S1(n1239), .Y(n2638) );
  AO21X1_HVT U65 ( .A1(n1626), .A2(n1242), .A3(n1650), .Y(n2635) );
  MUX41X1_HVT U67 ( .A1(n1624), .A3(n2635), .A2(n2634), .A4(n2636), .S0(n1448), 
        .S1(n892), .Y(n2633) );
  MUX41X1_HVT U68 ( .A1(n2633), .A3(n2637), .A2(n2643), .A4(n2647), .S0(
        keyin[105]), .S1(n1366), .Y(dummy[7]) );
  MUX41X1_HVT U69 ( .A1(n2658), .A3(n1672), .A2(n2676), .A4(n1658), .S0(n1239), 
        .S1(n1452), .Y(n2632) );
  NAND2X0_HVT U71 ( .A1(n1408), .A2(n2629), .Y(n2630) );
  AND3X1_HVT U75 ( .A1(n1406), .A2(n2641), .A3(n2624), .Y(n2625) );
  MUX41X1_HVT U77 ( .A1(n2656), .A3(n1615), .A2(n2680), .A4(n1407), .S0(n892), 
        .S1(n1243), .Y(n2622) );
  MUX41X1_HVT U80 ( .A1(n2620), .A3(n1659), .A2(n1660), .A4(n1635), .S0(n1240), 
        .S1(n870), .Y(n2619) );
  MUX41X1_HVT U81 ( .A1(n2691), .A3(n1652), .A2(n1661), .A4(n1673), .S0(n1240), 
        .S1(n517), .Y(n2618) );
  AND2X1_HVT U82 ( .A1(n1444), .A2(n1370), .Y(n2617) );
  NAND2X0_HVT U83 ( .A1(n1446), .A2(n1672), .Y(n2616) );
  MUX41X1_HVT U84 ( .A1(n2616), .A3(n2693), .A2(n1191), .A4(n2617), .S0(n1240), 
        .S1(n1452), .Y(n2615) );
  MUX41X1_HVT U85 ( .A1(n1659), .A3(n1634), .A2(n1204), .A4(n2682), .S0(n1239), 
        .S1(n870), .Y(n2614) );
  AO21X1_HVT U93 ( .A1(n1245), .A2(n2606), .A3(n1655), .Y(n2607) );
  MUX41X1_HVT U94 ( .A1(n2607), .A3(n2609), .A2(n2608), .A4(n2611), .S0(n298), 
        .S1(n1241), .Y(n2605) );
  NAND2X0_HVT U97 ( .A1(n2601), .A2(n2600), .Y(n2602) );
  MUX41X1_HVT U98 ( .A1(n2602), .A3(n1640), .A2(n2603), .A4(n2604), .S0(n1448), 
        .S1(n1240), .Y(n2599) );
  MUX41X1_HVT U102 ( .A1(n1652), .A3(n1615), .A2(n1440), .A4(n1658), .S0(n1239), .S1(n1244), .Y(n2595) );
  MUX41X1_HVT U104 ( .A1(n2654), .A3(n1654), .A2(n1625), .A4(n2668), .S0(n517), 
        .S1(n1238), .Y(n2593) );
  OA21X1_HVT U110 ( .A1(n1644), .A2(n1449), .A3(n1628), .Y(n2588) );
  NAND2X0_HVT U111 ( .A1(n1405), .A2(n2586), .Y(n2587) );
  NAND2X0_HVT U118 ( .A1(n2578), .A2(n2577), .Y(n2579) );
  MUX41X1_HVT U120 ( .A1(n2679), .A3(n1217), .A2(n1624), .A4(n1663), .S0(n1448), .S1(n1452), .Y(n2575) );
  AND2X1_HVT U122 ( .A1(n1440), .A2(n238), .Y(n2573) );
  MUX41X1_HVT U123 ( .A1(n2686), .A3(n2573), .A2(n1635), .A4(n2672), .S0(n298), 
        .S1(n870), .Y(n2572) );
  AO21X1_HVT U125 ( .A1(n298), .A2(n1408), .A3(n2693), .Y(n2570) );
  AND3X1_HVT U129 ( .A1(n297), .A2(n1446), .A3(n237), .Y(n2566) );
  MUX41X1_HVT U132 ( .A1(n2564), .A3(n2566), .A2(n2565), .A4(n2567), .S0(n1239), .S1(n1452), .Y(n2563) );
  MUX41X1_HVT U134 ( .A1(n1668), .A3(n2675), .A2(n1663), .A4(n1407), .S0(n517), 
        .S1(n1238), .Y(n2562) );
  AND2X1_HVT U138 ( .A1(n2699), .A2(n1445), .Y(n2558) );
  MUX41X1_HVT U139 ( .A1(n1634), .A3(n1653), .A2(n2677), .A4(n2558), .S0(n517), 
        .S1(n1240), .Y(n2557) );
  MUX41X1_HVT U140 ( .A1(n2557), .A3(n2559), .A2(n2560), .A4(n2562), .S0(n1448), .S1(keyin[105]), .Y(n2556) );
  MUX41X1_HVT U143 ( .A1(n2678), .A3(n1191), .A2(n1645), .A4(n1665), .S0(n1240), .S1(n1451), .Y(n2553) );
  NAND2X0_HVT U144 ( .A1(n1444), .A2(n1410), .Y(n2629) );
  MUX41X1_HVT U148 ( .A1(n1665), .A3(n1652), .A2(n2673), .A4(n1620), .S0(n1452), .S1(n1238), .Y(n2550) );
  MUX41X1_HVT U151 ( .A1(n1189), .A3(n1616), .A2(n1660), .A4(n1668), .S0(n892), 
        .S1(n1238), .Y(n2548) );
  AND2X1_HVT U156 ( .A1(n2693), .A2(n2629), .Y(n2542) );
  MUX41X1_HVT U158 ( .A1(n2655), .A3(n2542), .A2(n2541), .A4(n2543), .S0(n1243), .S1(n1451), .Y(n2540) );
  MUX41X1_HVT U159 ( .A1(n2679), .A3(n1632), .A2(n1639), .A4(n1206), .S0(n1239), .S1(n870), .Y(n2539) );
  AND2X1_HVT U161 ( .A1(n1451), .A2(n1368), .Y(n2537) );
  NAND2X0_HVT U165 ( .A1(n1440), .A2(n1672), .Y(n2533) );
  MUX41X1_HVT U166 ( .A1(n2686), .A3(n2663), .A2(n2533), .A4(n1661), .S0(n1240), .S1(n892), .Y(n2532) );
  NAND2X0_HVT U167 ( .A1(n1410), .A2(n2641), .Y(n2531) );
  NAND2X0_HVT U171 ( .A1(n1673), .A2(n1446), .Y(n2527) );
  NAND2X0_HVT U175 ( .A1(n1442), .A2(n2693), .Y(n2685) );
  NAND2X0_HVT U176 ( .A1(n1442), .A2(n1674), .Y(n2524) );
  MUX41X1_HVT U179 ( .A1(n2681), .A3(n1674), .A2(n1666), .A4(n2522), .S0(n1241), .S1(n870), .Y(n2521) );
  MUX41X1_HVT U180 ( .A1(n2616), .A3(n233), .A2(n1649), .A4(n1617), .S0(n1452), 
        .S1(keyin[106]), .Y(n2520) );
  MUX41X1_HVT U184 ( .A1(n2517), .A3(n2521), .A2(n2520), .A4(n2523), .S0(
        keyin[105]), .S1(n1448), .Y(n2516) );
  MUX41X1_HVT U185 ( .A1(n2686), .A3(n1667), .A2(n1190), .A4(n1666), .S0(n1241), .S1(n1245), .Y(n2515) );
  MUX41X1_HVT U186 ( .A1(n1622), .A3(n2674), .A2(n2691), .A4(n1619), .S0(n1241), .S1(n892), .Y(n2514) );
  MUX41X1_HVT U188 ( .A1(n2513), .A3(n2664), .A2(n1654), .A4(n2655), .S0(n1239), .S1(n1244), .Y(n2512) );
  MUX41X1_HVT U190 ( .A1(n2511), .A3(n1197), .A2(n2685), .A4(n2629), .S0(n1241), .S1(n892), .Y(n2510) );
  MUX41X1_HVT U191 ( .A1(n2510), .A3(n2514), .A2(n2512), .A4(n2515), .S0(
        keyin[105]), .S1(n297), .Y(n2509) );
  MUX41X1_HVT U194 ( .A1(n1664), .A3(n2668), .A2(n1407), .A4(n2508), .S0(n1241), .S1(n892), .Y(n2507) );
  MUX41X1_HVT U195 ( .A1(n2660), .A3(n2696), .A2(n2675), .A4(n2653), .S0(n1241), .S1(n1452), .Y(n2506) );
  AO21X1_HVT U202 ( .A1(n1204), .A2(n1244), .A3(n1655), .Y(n2499) );
  MUX41X1_HVT U204 ( .A1(n1623), .A3(n2693), .A2(n1666), .A4(n1409), .S0(n1241), .S1(n892), .Y(n2497) );
  MUX41X1_HVT U205 ( .A1(n2697), .A3(n2686), .A2(n1638), .A4(n2678), .S0(n1241), .S1(n1452), .Y(n2496) );
  MUX41X1_HVT U206 ( .A1(n237), .A3(n2642), .A2(n1667), .A4(n1642), .S0(n1241), 
        .S1(n870), .Y(n2495) );
  MUX41X1_HVT U207 ( .A1(n2495), .A3(n2497), .A2(n2496), .A4(n2498), .S0(
        keyin[105]), .S1(n297), .Y(n2494) );
  NAND2X0_HVT U211 ( .A1(n1408), .A2(n1444), .Y(n2641) );
  NAND2X0_HVT U212 ( .A1(n1441), .A2(n1402), .Y(n2586) );
  NAND2X0_HVT U215 ( .A1(n2693), .A2(n1446), .Y(n2493) );
  NAND2X0_HVT U216 ( .A1(n1408), .A2(n2586), .Y(n2492) );
  NAND2X0_HVT U219 ( .A1(n1444), .A2(n1668), .Y(n2545) );
  NAND2X0_HVT U221 ( .A1(n1452), .A2(n2493), .Y(n2624) );
  NAND2X0_HVT U317 ( .A1(n1428), .A2(n1397), .Y(n2477) );
  NAND2X0_HVT U318 ( .A1(n1362), .A2(n1427), .Y(n2476) );
  NAND2X0_HVT U319 ( .A1(n1395), .A2(n2477), .Y(n2475) );
  XOR2X2_HVT U320 ( .A1(n1608), .A2(n1363), .Y(n2473) );
  NAND2X0_HVT U328 ( .A1(n2465), .A2(n1401), .Y(n2466) );
  NAND2X0_HVT U330 ( .A1(n2477), .A2(n1343), .Y(n2463) );
  NAND2X0_HVT U334 ( .A1(n2474), .A2(n1432), .Y(n2459) );
  NAND2X0_HVT U338 ( .A1(n1361), .A2(n1432), .Y(n2456) );
  NAND2X0_HVT U346 ( .A1(n1432), .A2(n1611), .Y(n2448) );
  NAND2X0_HVT U347 ( .A1(n1607), .A2(n1432), .Y(n2447) );
  NAND2X0_HVT U352 ( .A1(n1427), .A2(n1344), .Y(n2442) );
  MUX41X1_HVT U363 ( .A1(n1593), .A3(n1550), .A2(n2467), .A4(n1570), .S0(n251), 
        .S1(n1434), .Y(n2432) );
  NAND2X0_HVT U365 ( .A1(n2429), .A2(n2439), .Y(n2430) );
  MUX41X1_HVT U368 ( .A1(n1183), .A3(n1569), .A2(n1568), .A4(n1342), .S0(n1437), .S1(n1229), .Y(n2426) );
  NAND2X0_HVT U369 ( .A1(n1432), .A2(n1398), .Y(n2425) );
  MUX41X1_HVT U370 ( .A1(n2425), .A3(n1558), .A2(n1588), .A4(n1567), .S0(n250), 
        .S1(n1435), .Y(n2424) );
  NAND2X0_HVT U372 ( .A1(n1395), .A2(n2421), .Y(n2422) );
  MUX41X1_HVT U373 ( .A1(n1594), .A3(n1566), .A2(n2422), .A4(n2470), .S0(n251), 
        .S1(n1229), .Y(n2420) );
  NAND2X0_HVT U374 ( .A1(n1401), .A2(n2477), .Y(n2419) );
  MUX41X1_HVT U375 ( .A1(n1215), .A3(n2419), .A2(n1211), .A4(n1565), .S0(n247), 
        .S1(n1229), .Y(n2418) );
  AO21X1_HVT U378 ( .A1(n1563), .A2(n1233), .A3(n1587), .Y(n2415) );
  MUX41X1_HVT U380 ( .A1(n1561), .A3(n2415), .A2(n2414), .A4(n2416), .S0(n516), 
        .S1(n1437), .Y(n2413) );
  MUX41X1_HVT U382 ( .A1(n2438), .A3(n1609), .A2(n2456), .A4(n1595), .S0(n1231), .S1(n1437), .Y(n2412) );
  NAND2X0_HVT U384 ( .A1(n1400), .A2(n2409), .Y(n2410) );
  AND3X1_HVT U388 ( .A1(n1398), .A2(n2421), .A3(n2404), .Y(n2405) );
  MUX41X1_HVT U390 ( .A1(n2436), .A3(n1551), .A2(n2460), .A4(n1399), .S0(n1235), .S1(n1232), .Y(n2402) );
  MUX41X1_HVT U393 ( .A1(n2400), .A3(n1596), .A2(n1597), .A4(n1572), .S0(n1434), .S1(n251), .Y(n2399) );
  MUX41X1_HVT U394 ( .A1(n2471), .A3(n1589), .A2(n1598), .A4(n1610), .S0(n1434), .S1(n842), .Y(n2398) );
  AND2X1_HVT U395 ( .A1(n1427), .A2(n1365), .Y(n2397) );
  NAND2X0_HVT U396 ( .A1(n1432), .A2(n1609), .Y(n2396) );
  MUX41X1_HVT U397 ( .A1(n2396), .A3(n242), .A2(n1185), .A4(n2397), .S0(n1434), 
        .S1(n842), .Y(n2395) );
  MUX41X1_HVT U398 ( .A1(n1596), .A3(n1571), .A2(n1200), .A4(n2462), .S0(n1231), .S1(n830), .Y(n2394) );
  MUX41X1_HVT U399 ( .A1(n2394), .A3(n2398), .A2(n2395), .A4(n2399), .S0(
        keyin[113]), .S1(n516), .Y(n2393) );
  AO21X1_HVT U406 ( .A1(n247), .A2(n2386), .A3(n1592), .Y(n2387) );
  NAND2X0_HVT U410 ( .A1(n2381), .A2(n2380), .Y(n2382) );
  MUX41X1_HVT U411 ( .A1(n2382), .A3(n1577), .A2(n2383), .A4(n2384), .S0(n516), 
        .S1(n1228), .Y(n2379) );
  MUX41X1_HVT U415 ( .A1(n1589), .A3(n1551), .A2(n1426), .A4(n1595), .S0(n1231), .S1(n1437), .Y(n2375) );
  MUX41X1_HVT U417 ( .A1(n2434), .A3(n1591), .A2(n1562), .A4(n2448), .S0(n247), 
        .S1(n1230), .Y(n2373) );
  MUX41X1_HVT U419 ( .A1(n1573), .A3(n2477), .A2(n2372), .A4(n1574), .S0(n1228), .S1(n251), .Y(n2371) );
  OA21X1_HVT U423 ( .A1(n1581), .A2(n1433), .A3(n1565), .Y(n2368) );
  NAND2X0_HVT U424 ( .A1(n1397), .A2(n2366), .Y(n2367) );
  NAND2X0_HVT U431 ( .A1(n2358), .A2(n2357), .Y(n2359) );
  AND2X1_HVT U435 ( .A1(n1430), .A2(n1342), .Y(n2353) );
  MUX41X1_HVT U436 ( .A1(n2466), .A3(n2353), .A2(n1572), .A4(n2452), .S0(n516), 
        .S1(n842), .Y(n2352) );
  AO21X1_HVT U438 ( .A1(n245), .A2(n1400), .A3(n242), .Y(n2350) );
  AND3X1_HVT U442 ( .A1(n245), .A2(n1432), .A3(n1364), .Y(n2346) );
  MUX41X1_HVT U447 ( .A1(n1605), .A3(n2455), .A2(n1600), .A4(n1399), .S0(n251), 
        .S1(n1230), .Y(n2342) );
  MUX41X1_HVT U450 ( .A1(n1342), .A3(n1583), .A2(n1399), .A4(n1578), .S0(n1231), .S1(n1235), .Y(n2339) );
  AND2X1_HVT U451 ( .A1(n2479), .A2(n1431), .Y(n2338) );
  MUX41X1_HVT U452 ( .A1(n1571), .A3(n1590), .A2(n2457), .A4(n2338), .S0(n1235), .S1(n1228), .Y(n2337) );
  MUX41X1_HVT U453 ( .A1(n2337), .A3(n2339), .A2(n2340), .A4(n2342), .S0(n516), 
        .S1(keyin[113]), .Y(n2336) );
  MUX41X1_HVT U456 ( .A1(n2458), .A3(n1185), .A2(n1582), .A4(n1602), .S0(n1229), .S1(n250), .Y(n2333) );
  NAND2X0_HVT U457 ( .A1(n1429), .A2(n1401), .Y(n2409) );
  MUX41X1_HVT U461 ( .A1(n1602), .A3(n1589), .A2(n2453), .A4(n1557), .S0(
        keyin[112]), .S1(n1230), .Y(n2330) );
  MUX41X1_HVT U464 ( .A1(n1183), .A3(n1552), .A2(n1597), .A4(n1605), .S0(
        keyin[112]), .S1(n1230), .Y(n2328) );
  AND2X1_HVT U469 ( .A1(n242), .A2(n2409), .Y(n2322) );
  MUX41X1_HVT U471 ( .A1(n2435), .A3(n2322), .A2(n2321), .A4(n2323), .S0(n1234), .S1(n842), .Y(n2320) );
  MUX41X1_HVT U472 ( .A1(n2459), .A3(n1569), .A2(n1576), .A4(n1202), .S0(n1231), .S1(n830), .Y(n2319) );
  MUX41X1_HVT U473 ( .A1(n2319), .A3(n2320), .A2(n2324), .A4(n2328), .S0(n516), 
        .S1(keyin[113]), .Y(n2318) );
  AND2X1_HVT U474 ( .A1(n1235), .A2(n1362), .Y(n2317) );
  NAND2X0_HVT U478 ( .A1(n1427), .A2(n1609), .Y(n2313) );
  MUX41X1_HVT U479 ( .A1(n2466), .A3(n2443), .A2(n2313), .A4(n1598), .S0(n1231), .S1(n250), .Y(n2312) );
  NAND2X0_HVT U480 ( .A1(n1401), .A2(n2421), .Y(n2311) );
  NAND2X0_HVT U484 ( .A1(n1610), .A2(n1432), .Y(n2307) );
  MUX41X1_HVT U485 ( .A1(n1399), .A3(n1595), .A2(n1594), .A4(n2307), .S0(
        keyin[112]), .S1(n1230), .Y(n2306) );
  NAND2X0_HVT U488 ( .A1(n1430), .A2(n242), .Y(n2465) );
  NAND2X0_HVT U489 ( .A1(n1426), .A2(n1611), .Y(n2304) );
  MUX41X1_HVT U490 ( .A1(n2304), .A3(n2443), .A2(n1599), .A4(n2465), .S0(n247), 
        .S1(n1228), .Y(n2303) );
  MUX41X1_HVT U492 ( .A1(n2461), .A3(n1611), .A2(n1603), .A4(n2302), .S0(n1232), .S1(n830), .Y(n2301) );
  MUX41X1_HVT U493 ( .A1(n2396), .A3(n1360), .A2(n1586), .A4(n1554), .S0(n1235), .S1(n1228), .Y(n2300) );
  MUX41X1_HVT U498 ( .A1(n2466), .A3(n1604), .A2(n1187), .A4(n1603), .S0(n1232), .S1(n1437), .Y(n2295) );
  MUX41X1_HVT U499 ( .A1(n1559), .A3(n2454), .A2(n2471), .A4(n1556), .S0(n1232), .S1(n247), .Y(n2294) );
  MUX41X1_HVT U501 ( .A1(n2293), .A3(n2444), .A2(n1591), .A4(n2435), .S0(n1231), .S1(n1437), .Y(n2292) );
  MUX41X1_HVT U503 ( .A1(n2291), .A3(n1195), .A2(n2465), .A4(n2409), .S0(n1232), .S1(n251), .Y(n2290) );
  MUX41X1_HVT U504 ( .A1(n2290), .A3(n2294), .A2(n2292), .A4(n2295), .S0(
        keyin[113]), .S1(n516), .Y(n2289) );
  MUX41X1_HVT U507 ( .A1(n1601), .A3(n2448), .A2(n1399), .A4(n2288), .S0(n1232), .S1(n830), .Y(n2287) );
  MUX41X1_HVT U508 ( .A1(n2440), .A3(n2476), .A2(n2455), .A4(n2433), .S0(n1232), .S1(n842), .Y(n2286) );
  MUX41X1_HVT U509 ( .A1(n1585), .A3(n2450), .A2(n2462), .A4(n1187), .S0(n1235), .S1(n1229), .Y(n2285) );
  MUX41X1_HVT U513 ( .A1(n2282), .A3(n2286), .A2(n2285), .A4(n2287), .S0(
        keyin[113]), .S1(n516), .Y(n2281) );
  AO21X1_HVT U515 ( .A1(n1200), .A2(n1237), .A3(n1592), .Y(n2279) );
  MUX41X1_HVT U517 ( .A1(n1560), .A3(n242), .A2(n1603), .A4(n2480), .S0(n1232), 
        .S1(n247), .Y(n2277) );
  MUX41X1_HVT U518 ( .A1(n2477), .A3(n2466), .A2(n1575), .A4(n2458), .S0(n1232), .S1(n830), .Y(n2276) );
  MUX41X1_HVT U519 ( .A1(n1364), .A3(n2422), .A2(n1604), .A4(n1579), .S0(n1232), .S1(n250), .Y(n2275) );
  NAND2X0_HVT U524 ( .A1(n1400), .A2(n1430), .Y(n2421) );
  NAND2X0_HVT U525 ( .A1(n1427), .A2(n2474), .Y(n2366) );
  NAND2X0_HVT U528 ( .A1(n242), .A2(n1432), .Y(n2273) );
  NAND2X0_HVT U529 ( .A1(n1400), .A2(n2366), .Y(n2272) );
  NAND2X0_HVT U532 ( .A1(n1429), .A2(n1605), .Y(n2325) );
  NAND2X0_HVT U534 ( .A1(n1235), .A2(n2273), .Y(n2404) );
  NAND2X0_HVT U630 ( .A1(n1414), .A2(n1389), .Y(n2257) );
  NAND2X0_HVT U631 ( .A1(n1357), .A2(n1413), .Y(n2256) );
  NAND2X0_HVT U632 ( .A1(n1387), .A2(n2257), .Y(n2255) );
  NAND2X0_HVT U641 ( .A1(n2245), .A2(n1393), .Y(n2246) );
  NAND2X0_HVT U643 ( .A1(n2257), .A2(n1339), .Y(n2243) );
  NAND2X0_HVT U647 ( .A1(n1386), .A2(n1417), .Y(n2239) );
  NAND2X0_HVT U651 ( .A1(n1357), .A2(n1417), .Y(n2236) );
  NAND2X0_HVT U659 ( .A1(n1417), .A2(n1542), .Y(n2228) );
  NAND2X0_HVT U660 ( .A1(n1538), .A2(n1417), .Y(n2227) );
  NAND2X0_HVT U665 ( .A1(n1411), .A2(n1341), .Y(n2222) );
  MUX41X1_HVT U676 ( .A1(n1525), .A3(n1484), .A2(n2247), .A4(n1504), .S0(n279), 
        .S1(n1219), .Y(n2212) );
  NAND2X0_HVT U678 ( .A1(n2209), .A2(n2219), .Y(n2210) );
  MUX41X1_HVT U681 ( .A1(n1184), .A3(n1503), .A2(n1502), .A4(n1338), .S0(n256), 
        .S1(n1220), .Y(n2206) );
  NAND2X0_HVT U682 ( .A1(n1417), .A2(n1390), .Y(n2205) );
  MUX41X1_HVT U683 ( .A1(n2205), .A3(n1492), .A2(n1520), .A4(n1501), .S0(n279), 
        .S1(n1219), .Y(n2204) );
  NAND2X0_HVT U685 ( .A1(n1387), .A2(n2201), .Y(n2202) );
  MUX41X1_HVT U686 ( .A1(n1526), .A3(n1500), .A2(n2202), .A4(n2250), .S0(n597), 
        .S1(n1220), .Y(n2200) );
  NAND2X0_HVT U687 ( .A1(n1393), .A2(n2257), .Y(n2199) );
  MUX41X1_HVT U688 ( .A1(n1216), .A3(n2199), .A2(n1212), .A4(n1499), .S0(n828), 
        .S1(n1219), .Y(n2198) );
  AO21X1_HVT U691 ( .A1(n1497), .A2(n1225), .A3(n1519), .Y(n2195) );
  MUX41X1_HVT U693 ( .A1(n1495), .A3(n2195), .A2(n2194), .A4(n2196), .S0(n289), 
        .S1(n597), .Y(n2193) );
  MUX41X1_HVT U695 ( .A1(n2218), .A3(n219), .A2(n2236), .A4(n1527), .S0(n1222), 
        .S1(n279), .Y(n2192) );
  NAND2X0_HVT U697 ( .A1(n1392), .A2(n2189), .Y(n2190) );
  AND3X1_HVT U701 ( .A1(n1390), .A2(n2201), .A3(n2184), .Y(n2185) );
  MUX41X1_HVT U703 ( .A1(n2216), .A3(n1485), .A2(n2240), .A4(n1391), .S0(n597), 
        .S1(n1219), .Y(n2182) );
  MUX41X1_HVT U704 ( .A1(n2182), .A3(n2183), .A2(n2187), .A4(n2192), .S0(n289), 
        .S1(keyin[121]), .Y(n2181) );
  MUX41X1_HVT U706 ( .A1(n2180), .A3(n1528), .A2(n1529), .A4(n1506), .S0(n1223), .S1(n1423), .Y(n2179) );
  MUX41X1_HVT U707 ( .A1(n2251), .A3(n1521), .A2(n1530), .A4(n1541), .S0(n1223), .S1(n1423), .Y(n2178) );
  AND2X1_HVT U708 ( .A1(n1413), .A2(n1358), .Y(n2177) );
  NAND2X0_HVT U709 ( .A1(n1417), .A2(n219), .Y(n2176) );
  MUX41X1_HVT U710 ( .A1(n2176), .A3(n2253), .A2(n1186), .A4(n2177), .S0(n1223), .S1(n596), .Y(n2175) );
  MUX41X1_HVT U711 ( .A1(n1528), .A3(n1505), .A2(n1201), .A4(n2242), .S0(n1222), .S1(n256), .Y(n2174) );
  AO21X1_HVT U719 ( .A1(n597), .A2(n2166), .A3(n1524), .Y(n2167) );
  NAND2X0_HVT U723 ( .A1(n2161), .A2(n2160), .Y(n2162) );
  MUX41X1_HVT U724 ( .A1(n2162), .A3(n1510), .A2(n2163), .A4(n2164), .S0(n289), 
        .S1(n1222), .Y(n2159) );
  MUX41X1_HVT U730 ( .A1(n2214), .A3(n1523), .A2(n1496), .A4(n2228), .S0(n828), 
        .S1(n1221), .Y(n2153) );
  NAND2X0_HVT U737 ( .A1(n1389), .A2(n2146), .Y(n2147) );
  MUX41X1_HVT U741 ( .A1(n2143), .A3(n2149), .A2(n2145), .A4(n2148), .S0(n1223), .S1(n828), .Y(n2142) );
  NAND2X0_HVT U744 ( .A1(n2138), .A2(n2137), .Y(n2139) );
  MUX41X1_HVT U746 ( .A1(n2239), .A3(n1216), .A2(n1495), .A4(n1532), .S0(n289), 
        .S1(n279), .Y(n2135) );
  AND2X1_HVT U748 ( .A1(n1411), .A2(n1338), .Y(n2133) );
  MUX41X1_HVT U749 ( .A1(n2246), .A3(n2133), .A2(n1506), .A4(n2232), .S0(n290), 
        .S1(n1423), .Y(n2132) );
  AO21X1_HVT U751 ( .A1(n289), .A2(n1392), .A3(n2253), .Y(n2130) );
  AND3X1_HVT U755 ( .A1(n1418), .A2(n1417), .A3(n1358), .Y(n2126) );
  MUX41X1_HVT U760 ( .A1(n1537), .A3(n2235), .A2(n1532), .A4(n1391), .S0(n279), 
        .S1(n1221), .Y(n2122) );
  AND2X1_HVT U764 ( .A1(n2259), .A2(n1416), .Y(n2118) );
  NAND2X0_HVT U770 ( .A1(n1412), .A2(n1394), .Y(n2189) );
  MUX41X1_HVT U777 ( .A1(n1184), .A3(n1486), .A2(n1529), .A4(n1537), .S0(n828), 
        .S1(n1221), .Y(n2107) );
  AND2X1_HVT U782 ( .A1(n2253), .A2(n2189), .Y(n2101) );
  MUX41X1_HVT U784 ( .A1(n2215), .A3(n2101), .A2(n2100), .A4(n2102), .S0(n1226), .S1(n279), .Y(n2099) );
  MUX41X1_HVT U785 ( .A1(n2239), .A3(n1503), .A2(n1509), .A4(n1203), .S0(n1222), .S1(n597), .Y(n2098) );
  AND2X1_HVT U787 ( .A1(n1424), .A2(n1357), .Y(n2096) );
  NAND2X0_HVT U791 ( .A1(n1411), .A2(n219), .Y(n2092) );
  MUX41X1_HVT U792 ( .A1(n2246), .A3(n2223), .A2(n2092), .A4(n1530), .S0(n1223), .S1(n256), .Y(n2091) );
  NAND2X0_HVT U793 ( .A1(n1393), .A2(n2201), .Y(n2090) );
  NAND2X0_HVT U797 ( .A1(n1541), .A2(n1417), .Y(n2086) );
  MUX41X1_HVT U798 ( .A1(n1391), .A3(n1527), .A2(n1526), .A4(n2086), .S0(n597), 
        .S1(n1221), .Y(n2085) );
  MUX41X1_HVT U799 ( .A1(n2085), .A3(n2091), .A2(n2087), .A4(n2093), .S0(n1359), .S1(n290), .Y(n2084) );
  NAND2X0_HVT U801 ( .A1(n1411), .A2(n2253), .Y(n2245) );
  NAND2X0_HVT U802 ( .A1(n1413), .A2(n1542), .Y(n2083) );
  MUX41X1_HVT U803 ( .A1(n2083), .A3(n2223), .A2(n1531), .A4(n2245), .S0(n596), 
        .S1(n1420), .Y(n2082) );
  MUX41X1_HVT U805 ( .A1(n2241), .A3(n1542), .A2(n1535), .A4(n2081), .S0(n1224), .S1(n279), .Y(n2080) );
  MUX41X1_HVT U806 ( .A1(n2176), .A3(keyin[124]), .A2(n1518), .A4(n1488), .S0(
        n279), .S1(n1223), .Y(n2079) );
  MUX41X1_HVT U810 ( .A1(n2076), .A3(n2080), .A2(n2079), .A4(n2082), .S0(
        keyin[121]), .S1(n1418), .Y(n2075) );
  MUX41X1_HVT U811 ( .A1(n2246), .A3(n1536), .A2(n1188), .A4(n1535), .S0(n1224), .S1(n1423), .Y(n2074) );
  MUX41X1_HVT U812 ( .A1(n1493), .A3(n2234), .A2(n2251), .A4(n1490), .S0(n1224), .S1(n596), .Y(n2073) );
  MUX41X1_HVT U814 ( .A1(n2072), .A3(n2224), .A2(n1523), .A4(n2215), .S0(n1222), .S1(n828), .Y(n2071) );
  MUX41X1_HVT U820 ( .A1(n1533), .A3(n2228), .A2(n1391), .A4(n2067), .S0(n1224), .S1(n596), .Y(n2066) );
  MUX41X1_HVT U821 ( .A1(n2220), .A3(n2256), .A2(n2235), .A4(n2213), .S0(n1224), .S1(n256), .Y(n2065) );
  MUX41X1_HVT U822 ( .A1(n1517), .A3(n2230), .A2(n2242), .A4(n1188), .S0(n256), 
        .S1(n1220), .Y(n2064) );
  MUX41X1_HVT U826 ( .A1(n2061), .A3(n2065), .A2(n2064), .A4(n2066), .S0(
        keyin[121]), .S1(n290), .Y(n2060) );
  AO21X1_HVT U828 ( .A1(n1201), .A2(n1227), .A3(n1524), .Y(n2058) );
  MUX41X1_HVT U830 ( .A1(n1494), .A3(n2253), .A2(n1535), .A4(n1393), .S0(n1224), .S1(n279), .Y(n2056) );
  MUX41X1_HVT U831 ( .A1(n2257), .A3(n2246), .A2(n545), .A4(n2238), .S0(n1224), 
        .S1(n596), .Y(n2055) );
  MUX41X1_HVT U832 ( .A1(n1358), .A3(n2202), .A2(n1536), .A4(n1512), .S0(n1224), .S1(n1423), .Y(n2054) );
  NAND2X0_HVT U837 ( .A1(n1392), .A2(n1413), .Y(n2201) );
  NAND2X0_HVT U838 ( .A1(n1414), .A2(n1386), .Y(n2146) );
  NAND2X0_HVT U841 ( .A1(n2253), .A2(n1417), .Y(n2052) );
  NAND2X0_HVT U842 ( .A1(n1392), .A2(n2146), .Y(n2051) );
  NAND2X0_HVT U845 ( .A1(n1412), .A2(n1537), .Y(n2104) );
  NAND2X0_HVT U847 ( .A1(n256), .A2(n2052), .Y(n2184) );
  NAND2X0_HVT U942 ( .A1(n301), .A2(n1378), .Y(n2037) );
  NAND2X0_HVT U943 ( .A1(n1459), .A2(n1354), .Y(n2035) );
  NAND2X0_HVT U944 ( .A1(n1372), .A2(n1457), .Y(n2034) );
  NAND2X0_HVT U945 ( .A1(n1381), .A2(n2037), .Y(n2033) );
  NAND2X0_HVT U952 ( .A1(n2026), .A2(n1384), .Y(n2027) );
  NAND2X0_HVT U954 ( .A1(n2037), .A2(n1351), .Y(n2024) );
  NAND2X0_HVT U960 ( .A1(n1381), .A2(n1459), .Y(n2018) );
  NAND2X0_HVT U963 ( .A1(n1372), .A2(n1459), .Y(n2016) );
  NAND2X0_HVT U971 ( .A1(n1735), .A2(n1459), .Y(n2007) );
  NAND2X0_HVT U977 ( .A1(n300), .A2(n1349), .Y(n2001) );
  MUX41X1_HVT U990 ( .A1(n1722), .A3(n1680), .A2(n2020), .A4(n1698), .S0(n305), 
        .S1(n1463), .Y(n1991) );
  NAND2X0_HVT U992 ( .A1(n1988), .A2(n1998), .Y(n1989) );
  NAND2X0_HVT U995 ( .A1(n1381), .A2(n1984), .Y(n1985) );
  MUX41X1_HVT U996 ( .A1(n1723), .A3(n1697), .A2(n1985), .A4(n2029), .S0(n1255), .S1(n1463), .Y(n1983) );
  NAND2X0_HVT U997 ( .A1(n1384), .A2(n2037), .Y(n1982) );
  MUX41X1_HVT U1000 ( .A1(n1193), .A3(n1695), .A2(n1694), .A4(n1353), .S0(
        n1255), .S1(n1463), .Y(n1979) );
  NAND2X0_HVT U1001 ( .A1(n1459), .A2(n1379), .Y(n1978) );
  MUX41X1_HVT U1002 ( .A1(n1978), .A3(n1686), .A2(n1717), .A4(n1693), .S0(
        n1255), .S1(n1252), .Y(n1977) );
  AO21X1_HVT U1005 ( .A1(n1691), .A2(n1254), .A3(n1716), .Y(n1974) );
  MUX41X1_HVT U1007 ( .A1(n1689), .A3(n1974), .A2(n1973), .A4(n1975), .S0(
        n1246), .S1(n1465), .Y(n1972) );
  NAND2X0_HVT U1012 ( .A1(n1383), .A2(n1967), .Y(n1968) );
  MUX41X1_HVT U1013 ( .A1(n1969), .A3(n1996), .A2(n1968), .A4(n2016), .S0(
        n1246), .S1(n1465), .Y(n1966) );
  MUX41X1_HVT U1014 ( .A1(n1720), .A3(n1725), .A2(n1738), .A4(n1700), .S0(
        n1246), .S1(n1464), .Y(n1965) );
  MUX41X1_HVT U1016 ( .A1(n2030), .A3(n1727), .A2(n1964), .A4(n1726), .S0(
        n1255), .S1(n1460), .Y(n1963) );
  MUX41X1_HVT U1017 ( .A1(n1963), .A3(n1966), .A2(n1965), .A4(n1970), .S0(
        n1371), .S1(n1463), .Y(n1962) );
  AND3X1_HVT U1019 ( .A1(n1984), .A2(n1378), .A3(n1959), .Y(n1960) );
  MUX41X1_HVT U1021 ( .A1(n1995), .A3(n1698), .A2(n1681), .A4(n2025), .S0(
        n1246), .S1(n293), .Y(n1957) );
  AND2X1_HVT U1022 ( .A1(n1456), .A2(n1375), .Y(n1956) );
  MUX41X1_HVT U1023 ( .A1(n1699), .A3(n524), .A2(n2023), .A4(n1956), .S0(n1246), .S1(n293), .Y(n1955) );
  NAND2X0_HVT U1024 ( .A1(n1459), .A2(n1737), .Y(n1954) );
  MUX41X1_HVT U1025 ( .A1(n1725), .A3(n1954), .A2(n1199), .A4(n1194), .S0(
        n1247), .S1(n293), .Y(n1953) );
  MUX41X1_HVT U1026 ( .A1(n1953), .A3(n1957), .A2(n1955), .A4(n1958), .S0(
        n1371), .S1(n1463), .Y(n1952) );
  AO21X1_HVT U1032 ( .A1(n1333), .A2(n1946), .A3(n1721), .Y(n1947) );
  MUX41X1_HVT U1035 ( .A1(n1681), .A3(n1205), .A2(n1724), .A4(n1944), .S0(
        n1248), .S1(n1464), .Y(n1943) );
  MUX41X1_HVT U1036 ( .A1(n1720), .A3(n1205), .A2(n276), .A4(n2024), .S0(n1246), .S1(n1464), .Y(n1942) );
  NAND2X0_HVT U1040 ( .A1(n1937), .A2(n1936), .Y(n1938) );
  MUX41X1_HVT U1042 ( .A1(n2037), .A3(n1690), .A2(n1702), .A4(n2035), .S0(
        n1246), .S1(n293), .Y(n1934) );
  MUX41X1_HVT U1044 ( .A1(n1701), .A3(n1993), .A2(n1933), .A4(n1719), .S0(
        n1246), .S1(n1464), .Y(n1932) );
  OA21X1_HVT U1048 ( .A1(n1709), .A2(n1462), .A3(n1696), .Y(n1929) );
  NAND2X0_HVT U1049 ( .A1(n1378), .A2(n1927), .Y(n1928) );
  MUX41X1_HVT U1053 ( .A1(n1924), .A3(n1930), .A2(n1926), .A4(n1929), .S0(
        n1254), .S1(n1464), .Y(n1923) );
  AND2X1_HVT U1054 ( .A1(n827), .A2(n1353), .Y(n1922) );
  MUX41X1_HVT U1055 ( .A1(n2027), .A3(n1922), .A2(n1700), .A4(n2009), .S0(
        n1247), .S1(n1465), .Y(n1921) );
  AO21X1_HVT U1057 ( .A1(n1251), .A2(n1382), .A3(n524), .Y(n1919) );
  NAND2X0_HVT U1062 ( .A1(n1913), .A2(n1912), .Y(n1914) );
  MUX41X1_HVT U1064 ( .A1(n2018), .A3(n1218), .A2(n1689), .A4(n1729), .S0(
        n1247), .S1(n1465), .Y(n1910) );
  AND3X1_HVT U1067 ( .A1(n1250), .A2(n1459), .A3(n1376), .Y(n1907) );
  MUX41X1_HVT U1070 ( .A1(n1905), .A3(n1907), .A2(n1906), .A4(n1908), .S0(
        n1254), .S1(n305), .Y(n1904) );
  MUX41X1_HVT U1074 ( .A1(n1730), .A3(n152), .A2(n2001), .A4(n2013), .S0(n1248), .S1(n1465), .Y(n1901) );
  MUX41X1_HVT U1075 ( .A1(n1194), .A3(n2007), .A2(n1731), .A4(n2005), .S0(
        n1247), .S1(n304), .Y(n1900) );
  MUX41X1_HVT U1078 ( .A1(n1898), .A3(n1901), .A2(n1900), .A4(n1902), .S0(
        n1371), .S1(n1252), .Y(n1897) );
  AND2X1_HVT U1079 ( .A1(n1382), .A2(n1458), .Y(n1896) );
  MUX41X1_HVT U1080 ( .A1(n2015), .A3(n1710), .A2(n1896), .A4(n1706), .S0(
        n1248), .S1(n304), .Y(n1895) );
  MUX41X1_HVT U1081 ( .A1(n1699), .A3(n1351), .A2(n1718), .A4(n1382), .S0(
        n1247), .S1(n305), .Y(n1894) );
  NAND2X0_HVT U1085 ( .A1(n1456), .A2(n1385), .Y(n1967) );
  MUX41X1_HVT U1086 ( .A1(n1731), .A3(n1967), .A2(n1720), .A4(n1994), .S0(
        n1248), .S1(n305), .Y(n1890) );
  MUX41X1_HVT U1087 ( .A1(n1890), .A3(n1894), .A2(n1891), .A4(n1895), .S0(
        keyin[103]), .S1(n1252), .Y(n1889) );
  MUX41X1_HVT U1092 ( .A1(n1928), .A3(n1193), .A2(n1377), .A4(n1679), .S0(
        n1247), .S1(n1466), .Y(n1884) );
  AND2X1_HVT U1093 ( .A1(n1333), .A2(n1372), .Y(n1883) );
  NAND2X0_HVT U1097 ( .A1(n301), .A2(n1737), .Y(n1879) );
  MUX41X1_HVT U1098 ( .A1(n2027), .A3(n1353), .A2(n1879), .A4(n1712), .S0(
        n1248), .S1(n1465), .Y(n1878) );
  AND2X1_HVT U1101 ( .A1(n524), .A2(n1967), .Y(n1875) );
  MUX41X1_HVT U1102 ( .A1(n1695), .A3(n1875), .A2(n1198), .A4(n1876), .S0(
        n1460), .S1(n304), .Y(n1874) );
  MUX41X1_HVT U1104 ( .A1(n2018), .A3(n1703), .A2(n1994), .A4(n1873), .S0(
        n1466), .S1(n1460), .Y(n1872) );
  NAND2X0_HVT U1105 ( .A1(n1384), .A2(n1984), .Y(n1871) );
  NAND2X0_HVT U1106 ( .A1(n1738), .A2(n1459), .Y(n1870) );
  MUX41X1_HVT U1107 ( .A1(n1723), .A3(n1382), .A2(n1870), .A4(n1871), .S0(
        n1249), .S1(n843), .Y(n1869) );
  MUX41X1_HVT U1111 ( .A1(n1866), .A3(n1872), .A2(n1869), .A4(n1874), .S0(
        n1371), .S1(n1253), .Y(n1865) );
  MUX21X2_HVT U1112 ( .A1(n1865), .A2(n1877), .S0(keyin[97]), .Y(dummy[26]) );
  NAND2X0_HVT U1113 ( .A1(n300), .A2(n2014), .Y(n2026) );
  MUX41X1_HVT U1115 ( .A1(n1355), .A3(n1864), .A2(n1728), .A4(n2026), .S0(n304), .S1(n1460), .Y(n1863) );
  NAND2X0_HVT U1116 ( .A1(n276), .A2(n1355), .Y(n1862) );
  MUX41X1_HVT U1117 ( .A1(n2022), .A3(n1862), .A2(n1732), .A4(n2003), .S0(
        n1250), .S1(n1466), .Y(n1861) );
  MUX41X1_HVT U1118 ( .A1(n2012), .A3(n1733), .A2(n1684), .A4(n1732), .S0(
        n1248), .S1(n293), .Y(n1860) );
  MUX41X1_HVT U1119 ( .A1(n1687), .A3(n2030), .A2(n2027), .A4(n1192), .S0(
        n1466), .S1(n1460), .Y(n1859) );
  MUX41X1_HVT U1120 ( .A1(n1859), .A3(n1861), .A2(n1860), .A4(n1863), .S0(
        keyin[103]), .S1(n1253), .Y(n1858) );
  MUX41X1_HVT U1121 ( .A1(n1711), .A3(n1380), .A2(n1714), .A4(n1715), .S0(
        n1466), .S1(n1460), .Y(n1857) );
  MUX41X1_HVT U1128 ( .A1(n1851), .A3(n2026), .A2(n1852), .A4(n1719), .S0(n304), .S1(n1460), .Y(n1850) );
  MUX41X1_HVT U1129 ( .A1(n1850), .A3(n1853), .A2(n1854), .A4(n1857), .S0(
        n1253), .S1(n1371), .Y(n1849) );
  MUX41X1_HVT U1132 ( .A1(n2034), .A3(n2035), .A2(n1992), .A4(n1848), .S0(
        n1460), .S1(n843), .Y(n1847) );
  MUX41X1_HVT U1133 ( .A1(n1999), .A3(n2013), .A2(n1730), .A4(n1382), .S0(n305), .S1(n1460), .Y(n1846) );
  MUX41X1_HVT U1134 ( .A1(n524), .A3(n1724), .A2(n1385), .A4(n2004), .S0(n1250), .S1(n843), .Y(n1845) );
  AO21X1_HVT U1136 ( .A1(n1199), .A2(n1259), .A3(n1721), .Y(n1843) );
  MUX41X1_HVT U1142 ( .A1(n2005), .A3(n1713), .A2(n2028), .A4(n2008), .S0(
        n1249), .S1(n843), .Y(n1837) );
  MUX41X1_HVT U1143 ( .A1(n1985), .A3(n2027), .A2(n1707), .A4(n2017), .S0(
        n1251), .S1(n843), .Y(n1836) );
  MUX41X1_HVT U1144 ( .A1(n288), .A3(n2037), .A2(n1733), .A4(n1705), .S0(n1249), .S1(n843), .Y(n1835) );
  MUX41X1_HVT U1145 ( .A1(n1835), .A3(n1837), .A2(n1836), .A4(n1838), .S0(
        n1371), .S1(n1253), .Y(n1834) );
  NAND2X0_HVT U1147 ( .A1(n827), .A2(n1381), .Y(n1927) );
  NAND2X0_HVT U1150 ( .A1(n1383), .A2(n300), .Y(n1984) );
  NAND2X0_HVT U1152 ( .A1(n524), .A2(n1459), .Y(n1833) );
  NAND2X0_HVT U1153 ( .A1(n1383), .A2(n1927), .Y(n1832) );
  NAND2X0_HVT U1156 ( .A1(n824), .A2(n1734), .Y(n1886) );
  NAND2X0_HVT U1159 ( .A1(n1259), .A2(n1833), .Y(n1959) );
  XOR2X2_HVT U1258 ( .A1(keyout[28]), .A2(n1808), .Y(keyout[92]) );
  XOR2X2_HVT U1260 ( .A1(keyout[26]), .A2(n1806), .Y(keyout[90]) );
  XOR2X2_HVT U1279 ( .A1(keyout[39]), .A2(keyin[71]), .Y(keyout[71]) );
  XOR3X2_HVT U1281 ( .A1(keyin[67]), .A2(n1820), .A3(n1819), .Y(keyout[67]) );
  XOR3X2_HVT U1282 ( .A1(keyin[66]), .A2(n1817), .A3(n1816), .Y(keyout[66]) );
  XOR2X2_HVT U1301 ( .A1(n1779), .A2(n1613), .Y(keyout[4]) );
  XOR2X2_HVT U1304 ( .A1(keyin[47]), .A2(n829), .Y(keyout[47]) );
  XOR2X2_HVT U1315 ( .A1(n1784), .A2(n1613), .Y(keyout[36]) );
  XOR2X2_HVT U1317 ( .A1(keyin[3]), .A2(dummy[3]), .Y(n1819) );
  XOR2X2_HVT U1322 ( .A1(keyin[32]), .A2(keyout[0]), .Y(keyout[32]) );
  XNOR2X2_HVT U1325 ( .A1(n1815), .A2(n1783), .Y(keyout[1]) );
  XOR2X2_HVT U1326 ( .A1(dummy[1]), .A2(keyin[1]), .Y(n1815) );
  XNOR2X2_HVT U1327 ( .A1(keyin[31]), .A2(dummy[31]), .Y(n1768) );
  XNOR2X2_HVT U1329 ( .A1(keyin[30]), .A2(dummy[30]), .Y(n1767) );
  XNOR2X2_HVT U1333 ( .A1(dummy[28]), .A2(keyin[28]), .Y(n1764) );
  XNOR2X2_HVT U1339 ( .A1(keyin[25]), .A2(dummy[25]), .Y(n1761) );
  XNOR2X2_HVT U1343 ( .A1(dummy[23]), .A2(keyin[23]), .Y(n1759) );
  XNOR2X2_HVT U1347 ( .A1(dummy[21]), .A2(keyin[21]), .Y(n1757) );
  XNOR2X2_HVT U1349 ( .A1(dummy[20]), .A2(keyin[20]), .Y(n1756) );
  XNOR2X2_HVT U1351 ( .A1(dummy[19]), .A2(keyin[19]), .Y(n1755) );
  XNOR2X2_HVT U1353 ( .A1(dummy[18]), .A2(keyin[18]), .Y(n1754) );
  XNOR2X2_HVT U1355 ( .A1(dummy[17]), .A2(keyin[17]), .Y(n1753) );
  XNOR2X2_HVT U1357 ( .A1(dummy[16]), .A2(keyin[16]), .Y(n1752) );
  XNOR2X2_HVT U1361 ( .A1(dummy[14]), .A2(keyin[14]), .Y(n1750) );
  XNOR2X2_HVT U1363 ( .A1(dummy[13]), .A2(keyin[13]), .Y(n1749) );
  XNOR2X2_HVT U1365 ( .A1(dummy[12]), .A2(keyin[12]), .Y(n1748) );
  XNOR2X2_HVT U1367 ( .A1(dummy[11]), .A2(keyin[11]), .Y(n1747) );
  XNOR2X2_HVT U1369 ( .A1(keyin[10]), .A2(dummy[10]), .Y(n1746) );
  XNOR2X2_HVT U1371 ( .A1(dummy[9]), .A2(keyin[9]), .Y(n1778) );
  XNOR2X2_HVT U1373 ( .A1(dummy[8]), .A2(keyin[8]), .Y(n1777) );
  XNOR2X2_HVT U1375 ( .A1(keyout[7]), .A2(keyin[39]), .Y(n1775) );
  XNOR2X2_HVT U1378 ( .A1(dummy[6]), .A2(keyin[6]), .Y(n1787) );
  XNOR2X2_HVT U1386 ( .A1(n1813), .A2(n1782), .Y(keyout[0]) );
  XOR2X2_HVT U1387 ( .A1(dummy[0]), .A2(keyin[0]), .Y(n1813) );
  XNOR3X1_HVT U1430 ( .A1(keyin[32]), .A2(keyin[64]), .A3(n1782), .Y(n1812) );
  NAND3X0_HVT U1431 ( .A1(n1772), .A2(n1771), .A3(n1770), .Y(n1776) );
  NAND4X0_HVT U1432 ( .A1(round_num[1]), .A2(round_num[3]), .A3(n1475), .A4(
        n1477), .Y(n1770) );
  AO21X1_HVT U1433 ( .A1(n1766), .A2(round_num[2]), .A3(n1470), .Y(n1769) );
  NAND4X0_HVT U1434 ( .A1(round_num[1]), .A2(round_num[2]), .A3(round_num[3]), 
        .A4(n1475), .Y(n1783) );
  XNOR3X1_HVT U1435 ( .A1(n1811), .A2(n1356), .A3(n1768), .Y(keyout[127]) );
  XNOR3X1_HVT U1436 ( .A1(n1810), .A2(n1413), .A3(n1767), .Y(keyout[126]) );
  XNOR3X1_HVT U1438 ( .A1(n1808), .A2(keyin[124]), .A3(n1764), .Y(keyout[124])
         );
  XNOR3X1_HVT U1439 ( .A1(n1807), .A2(n1358), .A3(n1763), .Y(keyout[123]) );
  XNOR3X1_HVT U1440 ( .A1(n1806), .A2(n1222), .A3(n1762), .Y(keyout[122]) );
  XNOR3X1_HVT U1441 ( .A1(n1805), .A2(keyin[121]), .A3(n212), .Y(keyout[121])
         );
  XNOR3X1_HVT U1443 ( .A1(n1803), .A2(keyin[119]), .A3(n1759), .Y(keyout[119])
         );
  XNOR3X1_HVT U1444 ( .A1(n1802), .A2(n1429), .A3(n1758), .Y(keyout[118]) );
  XNOR3X1_HVT U1446 ( .A1(n1800), .A2(n1360), .A3(n1756), .Y(keyout[116]) );
  XNOR3X1_HVT U1447 ( .A1(n1799), .A2(n1363), .A3(n610), .Y(keyout[115]) );
  XNOR3X1_HVT U1448 ( .A1(n1798), .A2(n1231), .A3(n1754), .Y(keyout[114]) );
  XNOR3X1_HVT U1449 ( .A1(n1797), .A2(keyin[113]), .A3(n1753), .Y(keyout[113])
         );
  XNOR3X1_HVT U1451 ( .A1(n1795), .A2(n1366), .A3(n1751), .Y(keyout[111]) );
  XNOR3X1_HVT U1452 ( .A1(n1794), .A2(n1440), .A3(n1750), .Y(keyout[110]) );
  XNOR3X1_HVT U1454 ( .A1(n1792), .A2(n233), .A3(n1748), .Y(keyout[108]) );
  XNOR3X1_HVT U1455 ( .A1(n1791), .A2(n1370), .A3(n1747), .Y(keyout[107]) );
  XNOR3X1_HVT U1456 ( .A1(n1790), .A2(n1239), .A3(n1746), .Y(keyout[106]) );
  XNOR3X1_HVT U1459 ( .A1(keyin[71]), .A2(keyin[103]), .A3(n1775), .Y(
        keyout[103]) );
  AND2X1_HVT U1461 ( .A1(n1771), .A2(n1744), .Y(n1786) );
  NAND3X0_HVT U1462 ( .A1(n1474), .A2(n1476), .A3(round_num[2]), .Y(n1744) );
  XNOR3X1_HVT U1463 ( .A1(n1471), .A2(n1743), .A3(n887), .Y(keyout[101]) );
  AND2X1_HVT U1464 ( .A1(n1772), .A2(n1742), .Y(n1780) );
  NAND4X0_HVT U1465 ( .A1(round_num[2]), .A2(round_num[3]), .A3(n1475), .A4(
        n1474), .Y(n1742) );
  NAND2X0_HVT U1466 ( .A1(round_num[2]), .A2(n1741), .Y(n1772) );
  AO21X1_HVT U1468 ( .A1(n1766), .A2(n1477), .A3(n1472), .Y(n1779) );
  NAND2X0_HVT U1469 ( .A1(round_num[0]), .A2(n1745), .Y(n1771) );
  AND3X1_HVT U1470 ( .A1(n1474), .A2(n1477), .A3(round_num[3]), .Y(n1745) );
  AND3X1_HVT U1471 ( .A1(n1475), .A2(n1476), .A3(round_num[1]), .Y(n1766) );
  NAND2X0_HVT U1472 ( .A1(n1741), .A2(n1477), .Y(n1782) );
  AND3X1_HVT U1473 ( .A1(n1474), .A2(n1476), .A3(round_num[0]), .Y(n1741) );
  INVX0_HVT U1 ( .A(n2254), .Y(n1538) );
  INVX2_HVT U2 ( .A(n609), .Y(n610) );
  NAND2X0_HVT U3 ( .A1(n855), .A2(n856), .Y(n23) );
  INVX0_HVT U7 ( .A(n1763), .Y(n49) );
  XNOR2X2_HVT U8 ( .A1(n23), .A2(keyin[27]), .Y(n1763) );
  NBUFFX2_HVT U9 ( .A(n1734), .Y(n152) );
  INVX0_HVT U10 ( .A(n1761), .Y(n211) );
  INVX1_HVT U11 ( .A(n211), .Y(n212) );
  AO21X1_HVT U12 ( .A1(n1458), .A2(n152), .A3(n1468), .Y(n1937) );
  XNOR2X1_HVT U13 ( .A1(n212), .A2(n1805), .Y(keyout[89]) );
  MUX21X1_HVT U14 ( .A1(n214), .A2(n2254), .S0(n1411), .Y(n213) );
  IBUFFX16_HVT U16 ( .A(n213), .Y(n2224) );
  IBUFFX16_HVT U18 ( .A(n1357), .Y(n214) );
  MUX21X2_HVT U19 ( .A1(n2078), .A2(n2077), .S0(n217), .Y(n2076) );
  IBUFFX16_HVT U20 ( .A(n1226), .Y(n217) );
  INVX0_HVT U22 ( .A(n1540), .Y(n218) );
  INVX1_HVT U23 ( .A(n218), .Y(n219) );
  INVX1_HVT U24 ( .A(n1394), .Y(n546) );
  INVX1_HVT U26 ( .A(n1416), .Y(n1414) );
  INVX1_HVT U27 ( .A(n1404), .Y(n1673) );
  XOR2X2_HVT U28 ( .A1(n862), .A2(n2675), .Y(n2657) );
  MUX21X1_HVT U29 ( .A1(n1388), .A2(n2170), .S0(n1208), .Y(n2169) );
  INVX1_HVT U30 ( .A(n1755), .Y(n609) );
  OR2X1_HVT U31 ( .A1(n220), .A2(n1365), .Y(n2474) );
  IBUFFX16_HVT U32 ( .A(n1344), .Y(n220) );
  MUX21X2_HVT U35 ( .A1(n2377), .A2(n1195), .S0(n232), .Y(n2376) );
  IBUFFX16_HVT U36 ( .A(n1235), .Y(n232) );
  INVX2_HVT U37 ( .A(keyin[123]), .Y(n1542) );
  INVX0_HVT U38 ( .A(n1671), .Y(n233) );
  INVX1_HVT U40 ( .A(n233), .Y(n234) );
  MUX41X1_HVT U41 ( .A1(n2554), .A3(n2551), .A2(n2553), .A4(n2550), .S0(n235), 
        .S1(n236), .Y(n2549) );
  IBUFFX16_HVT U42 ( .A(keyin[105]), .Y(n235) );
  IBUFFX16_HVT U43 ( .A(n298), .Y(n236) );
  XNOR2X1_HVT U44 ( .A1(dummy[26]), .A2(keyin[26]), .Y(n1762) );
  INVX1_HVT U45 ( .A(n1388), .Y(n1541) );
  NBUFFX2_HVT U46 ( .A(keyin[107]), .Y(n237) );
  INVX1_HVT U47 ( .A(n271), .Y(n238) );
  INVX1_HVT U48 ( .A(n1669), .Y(n271) );
  MUX21X2_HVT U49 ( .A1(n2111), .A2(n2112), .S0(n239), .Y(n2110) );
  IBUFFX16_HVT U51 ( .A(n1226), .Y(n239) );
  MUX41X1_HVT U53 ( .A1(n2110), .A3(n2114), .A2(n2109), .A4(n2113), .S0(
        keyin[121]), .S1(n240), .Y(n2108) );
  IBUFFX16_HVT U54 ( .A(keyin[125]), .Y(n240) );
  XOR2X2_HVT U58 ( .A1(dummy[27]), .A2(keyin[27]), .Y(keyout[27]) );
  XNOR2X2_HVT U63 ( .A1(n1767), .A2(n1810), .Y(keyout[94]) );
  NBUFFX2_HVT U64 ( .A(n2473), .Y(n242) );
  MUX41X1_HVT U66 ( .A1(n2278), .A3(n2276), .A2(n2277), .A4(n2275), .S0(n243), 
        .S1(n244), .Y(n2274) );
  IBUFFX16_HVT U70 ( .A(keyin[113]), .Y(n243) );
  IBUFFX16_HVT U72 ( .A(n516), .Y(n244) );
  NBUFFX2_HVT U73 ( .A(keyin[117]), .Y(n245) );
  MUX21X1_HVT U74 ( .A1(n2367), .A2(n2452), .S0(n246), .Y(n2365) );
  IBUFFX16_HVT U76 ( .A(n245), .Y(n246) );
  INVX1_HVT U78 ( .A(keyin[117]), .Y(n1433) );
  MUX21X1_HVT U79 ( .A1(n2371), .A2(n2373), .S0(n245), .Y(n2370) );
  INVX2_HVT U86 ( .A(n549), .Y(n247) );
  MUX21X2_HVT U87 ( .A1(n2446), .A2(n2447), .S0(n891), .Y(n2335) );
  INVX1_HVT U88 ( .A(n1236), .Y(n549) );
  INVX1_HVT U89 ( .A(n1236), .Y(n891) );
  XOR2X2_HVT U90 ( .A1(dummy[26]), .A2(keyin[26]), .Y(keyout[26]) );
  INVX1_HVT U91 ( .A(keyin[104]), .Y(n249) );
  MUX21X1_HVT U92 ( .A1(n1609), .A2(n1342), .S0(n263), .Y(n2472) );
  OA21X1_HVT U95 ( .A1(n2472), .A2(n1439), .A3(n1583), .Y(n2283) );
  INVX0_HVT U96 ( .A(n1439), .Y(n250) );
  INVX0_HVT U99 ( .A(n1439), .Y(n251) );
  MUX21X1_HVT U100 ( .A1(n255), .A2(n253), .S0(n254), .Y(n252) );
  IBUFFX16_HVT U101 ( .A(n252), .Y(n2331) );
  IBUFFX16_HVT U103 ( .A(n2332), .Y(n253) );
  IBUFFX16_HVT U105 ( .A(n1234), .Y(n254) );
  OAI21X2_HVT U106 ( .A1(n1555), .A2(n1439), .A3(n2452), .Y(n255) );
  IBUFFX2_HVT U107 ( .A(n1439), .Y(n1437) );
  XNOR2X1_HVT U108 ( .A1(keyin[58]), .A2(n1762), .Y(keyout[58]) );
  INVX0_HVT U109 ( .A(n1425), .Y(n256) );
  INVX2_HVT U112 ( .A(keyin[120]), .Y(n1425) );
  OA21X1_HVT U113 ( .A1(n1683), .A2(n1468), .A3(n2009), .Y(n1892) );
  MUX21X1_HVT U114 ( .A1(n1918), .A2(n1921), .S0(n1254), .Y(n1917) );
  IBUFFX2_HVT U115 ( .A(n251), .Y(n270) );
  MUX21X2_HVT U116 ( .A1(n2405), .A2(n2406), .S0(n257), .Y(n2403) );
  IBUFFX16_HVT U117 ( .A(n1234), .Y(n257) );
  MUX41X1_HVT U119 ( .A1(n2403), .A3(n2402), .A2(n2412), .A4(n2407), .S0(n258), 
        .S1(keyin[113]), .Y(n2401) );
  IBUFFX16_HVT U121 ( .A(n516), .Y(n258) );
  INVX2_HVT U124 ( .A(keyin[102]), .Y(n1458) );
  INVX0_HVT U126 ( .A(n1458), .Y(n1455) );
  INVX0_HVT U127 ( .A(n1458), .Y(n824) );
  INVX0_HVT U128 ( .A(n1458), .Y(n1457) );
  INVX0_HVT U130 ( .A(n1458), .Y(n1456) );
  MUX41X1_HVT U131 ( .A1(n2171), .A3(n2168), .A2(n2169), .A4(n2167), .S0(n259), 
        .S1(n260), .Y(n2165) );
  IBUFFX16_HVT U133 ( .A(n1418), .Y(n259) );
  IBUFFX16_HVT U135 ( .A(n1220), .Y(n260) );
  XOR2X1_HVT U136 ( .A1(n523), .A2(n827), .Y(n261) );
  IBUFFX16_HVT U137 ( .A(n261), .Y(n1994) );
  MUX41X1_HVT U141 ( .A1(n2002), .A3(n1205), .A2(n1994), .A4(n1967), .S0(n262), 
        .S1(n293), .Y(n1853) );
  IBUFFX16_HVT U142 ( .A(n1248), .Y(n262) );
  INVX1_HVT U145 ( .A(n1462), .Y(n1461) );
  INVX2_HVT U146 ( .A(n1462), .Y(n1460) );
  INVX2_HVT U147 ( .A(keyin[101]), .Y(n1462) );
  NAND2X0_HVT U149 ( .A1(n1839), .A2(n554), .Y(n555) );
  IBUFFX16_HVT U150 ( .A(n1426), .Y(n263) );
  MUX21X2_HVT U152 ( .A1(n2283), .A2(n2284), .S0(n264), .Y(n2282) );
  IBUFFX16_HVT U153 ( .A(n1234), .Y(n264) );
  XOR2X2_HVT U154 ( .A1(keyin[124]), .A2(keyin[123]), .Y(n265) );
  INVX8_HVT U155 ( .A(n265), .Y(n2253) );
  INVX0_HVT U157 ( .A(keyin[124]), .Y(n1539) );
  XOR2X1_HVT U160 ( .A1(n1462), .A2(n267), .Y(n266) );
  IBUFFX16_HVT U162 ( .A(n266), .Y(n1178) );
  IBUFFX16_HVT U163 ( .A(n1466), .Y(n267) );
  INVX1_HVT U164 ( .A(n1377), .Y(n1738) );
  MUX21X2_HVT U168 ( .A1(n1706), .A2(n2022), .S0(n268), .Y(n1905) );
  IBUFFX16_HVT U169 ( .A(n1248), .Y(n268) );
  MUX21X1_HVT U170 ( .A1(n2477), .A2(n1580), .S0(n1433), .Y(n2369) );
  MUX41X1_HVT U172 ( .A1(n2368), .A3(n2365), .A2(n2369), .A4(n2363), .S0(n269), 
        .S1(n270), .Y(n2362) );
  IBUFFX16_HVT U173 ( .A(n1434), .Y(n269) );
  INVX1_HVT U174 ( .A(n271), .Y(n272) );
  INVX0_HVT U177 ( .A(n271), .Y(n273) );
  MUX41X1_HVT U178 ( .A1(n2334), .A3(n2331), .A2(n2333), .A4(n2330), .S0(n274), 
        .S1(n275), .Y(n2329) );
  IBUFFX16_HVT U181 ( .A(keyin[113]), .Y(n274) );
  IBUFFX16_HVT U182 ( .A(n516), .Y(n275) );
  NBUFFX2_HVT U183 ( .A(keyin[102]), .Y(n276) );
  MUX41X1_HVT U187 ( .A1(n1885), .A3(n1880), .A2(n1884), .A4(n1878), .S0(n277), 
        .S1(n278), .Y(n1877) );
  IBUFFX16_HVT U189 ( .A(keyin[103]), .Y(n277) );
  IBUFFX16_HVT U192 ( .A(n1252), .Y(n278) );
  NBUFFX4_HVT U193 ( .A(keyin[120]), .Y(n279) );
  INVX1_HVT U196 ( .A(keyin[120]), .Y(n866) );
  MUX41X1_HVT U197 ( .A1(n2391), .A3(n2388), .A2(n2389), .A4(n2387), .S0(n280), 
        .S1(n281), .Y(n2385) );
  IBUFFX16_HVT U198 ( .A(n516), .Y(n280) );
  IBUFFX16_HVT U199 ( .A(n1229), .Y(n281) );
  MUX41X1_HVT U200 ( .A1(n1939), .A3(n1934), .A2(n1935), .A4(n1932), .S0(n282), 
        .S1(n283), .Y(n1931) );
  IBUFFX16_HVT U201 ( .A(keyin[103]), .Y(n282) );
  IBUFFX16_HVT U203 ( .A(n1252), .Y(n283) );
  INVX0_HVT U208 ( .A(keyin[99]), .Y(n284) );
  INVX0_HVT U209 ( .A(n284), .Y(n285) );
  MUX21X2_HVT U210 ( .A1(n1882), .A2(n1881), .S0(n286), .Y(n1880) );
  IBUFFX16_HVT U213 ( .A(n1251), .Y(n286) );
  XNOR2X2_HVT U214 ( .A1(n554), .A2(n287), .Y(n1179) );
  IBUFFX16_HVT U217 ( .A(n827), .Y(n287) );
  XOR2X2_HVT U218 ( .A1(n1671), .A2(n1369), .Y(n2693) );
  NBUFFX2_HVT U220 ( .A(n285), .Y(n288) );
  XNOR2X1_HVT U222 ( .A1(n1765), .A2(n1809), .Y(keyout[93]) );
  INVX0_HVT U223 ( .A(n1250), .Y(n554) );
  INVX0_HVT U224 ( .A(n1419), .Y(n289) );
  INVX1_HVT U225 ( .A(n1419), .Y(n290) );
  MUX41X1_HVT U226 ( .A1(n2203), .A3(n2207), .A2(n2193), .A4(n2197), .S0(n291), 
        .S1(n295), .Y(dummy[23]) );
  IBUFFX16_HVT U227 ( .A(n294), .Y(n291) );
  INVX0_HVT U228 ( .A(n1419), .Y(n589) );
  XOR2X2_HVT U229 ( .A1(keyin[31]), .A2(dummy[31]), .Y(keyout[31]) );
  INVX1_HVT U230 ( .A(n1468), .Y(n293) );
  INVX1_HVT U231 ( .A(n1468), .Y(n1464) );
  MUX21X1_HVT U232 ( .A1(n2256), .A2(n2172), .S0(n1227), .Y(n2171) );
  XOR2X2_HVT U233 ( .A1(keyin[57]), .A2(keyout[25]), .Y(keyout[57]) );
  INVX2_HVT U234 ( .A(n1761), .Y(keyout[25]) );
  MUX21X2_HVT U235 ( .A1(n1911), .A2(n1910), .S0(n850), .Y(n1909) );
  IBUFFX16_HVT U236 ( .A(n1359), .Y(n294) );
  IBUFFX16_HVT U237 ( .A(n1356), .Y(n295) );
  MUX21X1_HVT U238 ( .A1(n2198), .A2(n2200), .S0(n289), .Y(n2197) );
  XOR2X2_HVT U239 ( .A1(keyin[61]), .A2(keyout[29]), .Y(keyout[61]) );
  NAND2X0_HVT U240 ( .A1(n900), .A2(n901), .Y(n296) );
  INVX1_HVT U241 ( .A(n1449), .Y(n297) );
  INVX1_HVT U242 ( .A(n1449), .Y(n298) );
  INVX0_HVT U243 ( .A(n1449), .Y(n1447) );
  MUX21X1_HVT U244 ( .A1(n2575), .A2(n2576), .S0(keyin[106]), .Y(n2574) );
  XOR2X2_HVT U245 ( .A1(n296), .A2(keyin[18]), .Y(keyout[18]) );
  XNOR2X2_HVT U246 ( .A1(keyin[62]), .A2(n1767), .Y(keyout[62]) );
  INVX0_HVT U247 ( .A(n1458), .Y(n300) );
  INVX0_HVT U248 ( .A(n1458), .Y(n1454) );
  MUX41X1_HVT U249 ( .A1(n1407), .A3(n1658), .A2(n1657), .A4(n2527), .S0(n892), 
        .S1(n1238), .Y(n2526) );
  NBUFFX2_HVT U250 ( .A(keyin[102]), .Y(n301) );
  MUX41X1_HVT U251 ( .A1(n1696), .A3(n1213), .A2(n1982), .A4(n1218), .S0(n302), 
        .S1(n303), .Y(n1981) );
  IBUFFX16_HVT U252 ( .A(n1255), .Y(n302) );
  IBUFFX16_HVT U253 ( .A(n1463), .Y(n303) );
  INVX1_HVT U254 ( .A(n1469), .Y(n304) );
  INVX1_HVT U255 ( .A(n1469), .Y(n305) );
  MUX21X2_HVT U256 ( .A1(n1991), .A2(n1987), .S0(n328), .Y(n1986) );
  IBUFFX16_HVT U257 ( .A(n1249), .Y(n328) );
  INVX0_HVT U258 ( .A(n1469), .Y(n1467) );
  MUX21X1_HVT U259 ( .A1(n1352), .A2(n1372), .S0(n300), .Y(n2017) );
  INVX0_HVT U260 ( .A(n249), .Y(n354) );
  INVX1_HVT U261 ( .A(n354), .Y(n457) );
  INVX1_HVT U262 ( .A(keyin[104]), .Y(n862) );
  NBUFFX4_HVT U263 ( .A(keyin[117]), .Y(n516) );
  XNOR2X2_HVT U264 ( .A1(keyin[44]), .A2(n1748), .Y(keyout[44]) );
  NBUFFX2_HVT U265 ( .A(n870), .Y(n517) );
  NBUFFX2_HVT U266 ( .A(keyin[104]), .Y(n870) );
  INVX0_HVT U267 ( .A(n290), .Y(n563) );
  XOR2X2_HVT U268 ( .A1(dummy[20]), .A2(keyin[20]), .Y(keyout[20]) );
  MUX21X2_HVT U269 ( .A1(n2130), .A2(n2131), .S0(n828), .Y(n2129) );
  XNOR2X1_HVT U270 ( .A1(keyin[52]), .A2(n1756), .Y(keyout[52]) );
  XOR2X2_HVT U271 ( .A1(n1817), .A2(n1168), .Y(keyout[34]) );
  MUX41X1_HVT U272 ( .A1(n2539), .A3(n2540), .A2(n2544), .A4(n2548), .S0(n298), 
        .S1(n519), .Y(n2538) );
  IBUFFX16_HVT U273 ( .A(n1160), .Y(n519) );
  MUX41X1_HVT U274 ( .A1(n2594), .A3(n2605), .A2(n2590), .A4(n2599), .S0(n1366), .S1(n522), .Y(n882) );
  IBUFFX16_HVT U275 ( .A(keyin[105]), .Y(n522) );
  INVX1_HVT U276 ( .A(n2014), .Y(n523) );
  INVX2_HVT U277 ( .A(n523), .Y(n524) );
  MUX41X1_HVT U278 ( .A1(n1986), .A3(n1976), .A2(n1980), .A4(n1972), .S0(n525), 
        .S1(n537), .Y(dummy[31]) );
  IBUFFX16_HVT U279 ( .A(keyin[97]), .Y(n525) );
  IBUFFX16_HVT U280 ( .A(keyin[103]), .Y(n537) );
  XNOR2X1_HVT U281 ( .A1(n882), .A2(keyin[5]), .Y(n1781) );
  XOR3X2_HVT U282 ( .A1(keyin[7]), .A2(n1745), .A3(dummy[7]), .Y(keyout[7]) );
  INVX0_HVT U283 ( .A(n2014), .Y(n1739) );
  XOR2X2_HVT U284 ( .A1(keyin[63]), .A2(keyout[31]), .Y(keyout[63]) );
  MUX21X2_HVT U285 ( .A1(n2595), .A2(n2596), .S0(keyin[109]), .Y(n2594) );
  XOR2X2_HVT U286 ( .A1(n1812), .A2(n884), .Y(keyout[64]) );
  XOR2X2_HVT U287 ( .A1(n1820), .A2(n1819), .Y(keyout[35]) );
  MUX41X1_HVT U288 ( .A1(n2502), .A3(n2506), .A2(n2505), .A4(n2507), .S0(n540), 
        .S1(n538), .Y(n2501) );
  IBUFFX16_HVT U289 ( .A(n541), .Y(n538) );
  XOR2X2_HVT U290 ( .A1(n1774), .A2(n1612), .Y(keyout[38]) );
  OAI21X2_HVT U291 ( .A1(n1618), .A2(n862), .A3(n2672), .Y(n1155) );
  OA21X1_HVT U292 ( .A1(n2692), .A2(n249), .A3(n1646), .Y(n2503) );
  OA21X1_HVT U293 ( .A1(n2669), .A2(n249), .A3(n1634), .Y(n2518) );
  OA21X1_HVT U294 ( .A1(n2661), .A2(n249), .A3(n2545), .Y(n2546) );
  XOR3X2_HVT U295 ( .A1(n1774), .A2(n1787), .A3(n539), .Y(keyout[102]) );
  XNOR2X1_HVT U296 ( .A1(keyin[70]), .A2(n1456), .Y(n539) );
  INVX0_HVT U297 ( .A(n1774), .Y(n1473) );
  XNOR2X2_HVT U298 ( .A1(n1786), .A2(keyin[38]), .Y(n1774) );
  INVX1_HVT U299 ( .A(n1787), .Y(n1612) );
  IBUFFX16_HVT U300 ( .A(n1160), .Y(n540) );
  IBUFFX16_HVT U301 ( .A(keyin[109]), .Y(n541) );
  IBUFFX16_HVT U302 ( .A(n1445), .Y(n1441) );
  INVX1_HVT U303 ( .A(n1416), .Y(n1413) );
  INVX0_HVT U304 ( .A(n1416), .Y(n1412) );
  INVX1_HVT U305 ( .A(n1416), .Y(n1411) );
  MUX21X2_HVT U306 ( .A1(n2106), .A2(n2105), .S0(n542), .Y(n2103) );
  IBUFFX16_HVT U307 ( .A(n544), .Y(n542) );
  INVX2_HVT U308 ( .A(n1453), .Y(n1451) );
  INVX1_HVT U309 ( .A(keyin[104]), .Y(n1453) );
  MUX21X2_HVT U310 ( .A1(n1711), .A2(n2017), .S0(n543), .Y(n1899) );
  IBUFFX16_HVT U311 ( .A(n1333), .Y(n543) );
  XOR2X2_HVT U312 ( .A1(n49), .A2(n1807), .Y(keyout[91]) );
  IBUFFX16_HVT U313 ( .A(n1225), .Y(n544) );
  INVX2_HVT U314 ( .A(keyin[125]), .Y(n1419) );
  INVX1_HVT U315 ( .A(n545), .Y(n2232) );
  IBUFFX2_HVT U316 ( .A(n589), .Y(n548) );
  MUX21X1_HVT U321 ( .A1(n546), .A2(n547), .S0(n1415), .Y(n545) );
  IBUFFX16_HVT U322 ( .A(n1392), .Y(n547) );
  MUX21X2_HVT U323 ( .A1(n2147), .A2(n2232), .S0(n548), .Y(n2145) );
  NBUFFX2_HVT U324 ( .A(n1739), .Y(n1352) );
  OA21X1_HVT U325 ( .A1(n1212), .A2(n866), .A3(n2232), .Y(n2088) );
  XOR2X2_HVT U326 ( .A1(keyin[55]), .A2(n1478), .Y(keyout[55]) );
  IBUFFX2_HVT U327 ( .A(n2250), .Y(n1497) );
  MUX21X2_HVT U329 ( .A1(n2279), .A2(n2280), .S0(n1233), .Y(n2278) );
  MUX21X2_HVT U331 ( .A1(n1595), .A2(n2445), .S0(n1237), .Y(n2280) );
  NAND2X0_HVT U332 ( .A1(n1570), .A2(n549), .Y(n550) );
  NAND2X0_HVT U333 ( .A1(n2464), .A2(n247), .Y(n551) );
  NAND2X0_HVT U335 ( .A1(n550), .A2(n551), .Y(n2406) );
  XNOR2X2_HVT U336 ( .A1(n610), .A2(n1799), .Y(keyout[83]) );
  MUX41X1_HVT U337 ( .A1(n1508), .A3(n2152), .A2(n2257), .A4(n1507), .S0(n552), 
        .S1(n1425), .Y(n2151) );
  IBUFFX16_HVT U339 ( .A(n1223), .Y(n552) );
  XOR2X2_HVT U340 ( .A1(keyin[24]), .A2(dummy[24]), .Y(keyout[24]) );
  NAND2X0_HVT U341 ( .A1(n1840), .A2(n1250), .Y(n556) );
  NAND2X0_HVT U342 ( .A1(n555), .A2(n556), .Y(n1838) );
  MUX21X1_HVT U343 ( .A1(n2023), .A2(n1192), .S0(n1255), .Y(n1840) );
  IBUFFX2_HVT U344 ( .A(n1431), .Y(n1429) );
  INVX2_HVT U345 ( .A(n1445), .Y(n1443) );
  MUX41X1_HVT U348 ( .A1(n2159), .A3(n2150), .A2(n2165), .A4(n2154), .S0(n557), 
        .S1(keyin[121]), .Y(dummy[21]) );
  IBUFFX16_HVT U349 ( .A(n1356), .Y(n557) );
  OA21X1_HVT U350 ( .A1(n1489), .A2(n866), .A3(n2232), .Y(n2111) );
  MUX41X1_HVT U351 ( .A1(n2534), .A3(n2532), .A2(n2528), .A4(n2526), .S0(n1449), .S1(n1160), .Y(n2525) );
  NAND2X1_HVT U353 ( .A1(n2535), .A2(n558), .Y(n559) );
  NAND2X0_HVT U354 ( .A1(n2536), .A2(n1243), .Y(n560) );
  NAND2X0_HVT U355 ( .A1(n560), .A2(n559), .Y(n2534) );
  IBUFFX2_HVT U356 ( .A(n1243), .Y(n558) );
  INVX0_HVT U357 ( .A(keyin[105]), .Y(n1160) );
  MUX21X1_HVT U358 ( .A1(n2537), .A2(n1405), .S0(n1209), .Y(n2536) );
  MUX21X2_HVT U359 ( .A1(n1899), .A2(n2033), .S0(n1248), .Y(n1898) );
  MUX21X1_HVT U360 ( .A1(n2538), .A2(n2525), .S0(n878), .Y(n881) );
  INVX2_HVT U361 ( .A(n1419), .Y(n1418) );
  INVX2_HVT U362 ( .A(keyin[110]), .Y(n1445) );
  MUX21X2_HVT U364 ( .A1(n2626), .A2(n2625), .S0(n1243), .Y(n2623) );
  MUX21X2_HVT U366 ( .A1(n1184), .A2(n2244), .S0(n1425), .Y(n2164) );
  IBUFFX2_HVT U367 ( .A(n1425), .Y(n596) );
  MUX21X2_HVT U371 ( .A1(n1633), .A2(n2684), .S0(n1245), .Y(n2626) );
  IBUFFX2_HVT U376 ( .A(n2244), .Y(n1501) );
  MUX41X1_HVT U377 ( .A1(n2128), .A3(n2142), .A2(n2123), .A4(n2134), .S0(n561), 
        .S1(n562), .Y(dummy[20]) );
  IBUFFX16_HVT U379 ( .A(n1132), .Y(n561) );
  IBUFFX16_HVT U381 ( .A(n1359), .Y(n562) );
  MUX41X1_HVT U383 ( .A1(n2099), .A3(n2098), .A2(n2107), .A4(n2103), .S0(n563), 
        .S1(n1359), .Y(n2097) );
  XNOR2X1_HVT U385 ( .A1(n1754), .A2(n1798), .Y(keyout[82]) );
  NBUFFX2_HVT U386 ( .A(n1443), .Y(n564) );
  NBUFFX4_HVT U387 ( .A(n1443), .Y(n565) );
  IBUFFX2_HVT U389 ( .A(n1445), .Y(n1442) );
  NBUFFX2_HVT U391 ( .A(n1428), .Y(n566) );
  NBUFFX2_HVT U392 ( .A(n1428), .Y(n567) );
  NBUFFX2_HVT U400 ( .A(n1428), .Y(n568) );
  IBUFFX2_HVT U401 ( .A(n1431), .Y(n1427) );
  NBUFFX2_HVT U402 ( .A(n1414), .Y(n569) );
  NBUFFX2_HVT U403 ( .A(n1414), .Y(n570) );
  NAND2X0_HVT U404 ( .A1(n605), .A2(n606), .Y(n2354) );
  INVX1_HVT U405 ( .A(n849), .Y(n598) );
  INVX1_HVT U407 ( .A(n1431), .Y(n1428) );
  OA21X1_HVT U408 ( .A1(n866), .A2(n2221), .A3(n2104), .Y(n2105) );
  OA21X1_HVT U409 ( .A1(n2006), .A2(n1468), .A3(n1699), .Y(n1855) );
  OA21X1_HVT U412 ( .A1(n2000), .A2(n1468), .A3(n1886), .Y(n1887) );
  INVX1_HVT U413 ( .A(keyin[96]), .Y(n1469) );
  INVX0_HVT U414 ( .A(n1227), .Y(n580) );
  NBUFFX2_HVT U416 ( .A(n1461), .Y(n1249) );
  XOR2X2_HVT U418 ( .A1(keyin[70]), .A2(n1473), .Y(n571) );
  XNOR3X1_HVT U420 ( .A1(n1801), .A2(n516), .A3(n1757), .Y(keyout[117]) );
  INVX0_HVT U421 ( .A(n1249), .Y(n581) );
  XNOR2X2_HVT U422 ( .A1(n1750), .A2(n1794), .Y(keyout[78]) );
  INVX1_HVT U425 ( .A(n1453), .Y(n892) );
  INVX1_HVT U426 ( .A(keyin[103]), .Y(n588) );
  INVX1_HVT U427 ( .A(keyin[97]), .Y(n587) );
  XNOR2X2_HVT U428 ( .A1(n1751), .A2(n1795), .Y(keyout[79]) );
  INVX0_HVT U429 ( .A(n898), .Y(n592) );
  INVX1_HVT U430 ( .A(keyin[119]), .Y(n898) );
  INVX1_HVT U432 ( .A(keyin[119]), .Y(n584) );
  INVX0_HVT U433 ( .A(n898), .Y(n604) );
  INVX1_HVT U434 ( .A(n1425), .Y(n597) );
  INVX1_HVT U437 ( .A(n1242), .Y(n1164) );
  INVX0_HVT U439 ( .A(n1233), .Y(n601) );
  NAND2X0_HVT U440 ( .A1(n2281), .A2(n575), .Y(n576) );
  NAND2X0_HVT U441 ( .A1(n2274), .A2(n584), .Y(n577) );
  NAND2X0_HVT U443 ( .A1(n576), .A2(n577), .Y(dummy[8]) );
  INVX1_HVT U444 ( .A(n584), .Y(n575) );
  MUX21X1_HVT U445 ( .A1(n2155), .A2(n2156), .S0(n290), .Y(n2154) );
  MUX41X1_HVT U446 ( .A1(n1521), .A3(n1485), .A2(n1415), .A4(n1527), .S0(n1222), .S1(n597), .Y(n2155) );
  INVX1_HVT U448 ( .A(n2048), .Y(n1527) );
  NAND2X0_HVT U449 ( .A1(n2243), .A2(n823), .Y(n578) );
  NAND2X0_HVT U454 ( .A1(n2158), .A2(n1226), .Y(n579) );
  NAND2X0_HVT U455 ( .A1(n578), .A2(n579), .Y(n2157) );
  MUX21X2_HVT U458 ( .A1(n2157), .A2(n1196), .S0(n580), .Y(n2156) );
  NAND2X0_HVT U459 ( .A1(n1977), .A2(n581), .Y(n582) );
  NAND2X0_HVT U460 ( .A1(n1979), .A2(n1249), .Y(n583) );
  NAND2X0_HVT U462 ( .A1(n582), .A2(n583), .Y(n1976) );
  XOR2X2_HVT U463 ( .A1(keyout[31]), .A2(n1811), .Y(keyout[95]) );
  NAND2X0_HVT U465 ( .A1(n2289), .A2(n584), .Y(n585) );
  NAND2X0_HVT U466 ( .A1(n2296), .A2(n592), .Y(n586) );
  NAND2X0_HVT U467 ( .A1(n585), .A2(n586), .Y(dummy[9]) );
  IBUFFX2_HVT U468 ( .A(keyin[126]), .Y(n1417) );
  MUX41X1_HVT U470 ( .A1(n1923), .A3(n1909), .A2(n1917), .A4(n1904), .S0(n587), 
        .S1(n588), .Y(dummy[28]) );
  MUX21X2_HVT U475 ( .A1(n2129), .A2(n2132), .S0(n1225), .Y(n2128) );
  NAND2X0_HVT U476 ( .A1(n2153), .A2(n289), .Y(n590) );
  NAND2X0_HVT U477 ( .A1(n2151), .A2(n1419), .Y(n591) );
  NAND2X0_HVT U481 ( .A1(n590), .A2(n591), .Y(n2150) );
  NAND2X0_HVT U482 ( .A1(n2408), .A2(n601), .Y(n593) );
  NAND2X0_HVT U483 ( .A1(n2437), .A2(n1233), .Y(n594) );
  NAND2X0_HVT U486 ( .A1(n593), .A2(n594), .Y(n2407) );
  MUX21X1_HVT U487 ( .A1(n2411), .A2(n2410), .S0(n1236), .Y(n2408) );
  XOR2X1_HVT U491 ( .A1(n1439), .A2(n2455), .Y(n2437) );
  NAND2X0_HVT U494 ( .A1(n859), .A2(n860), .Y(n595) );
  XOR2X2_HVT U495 ( .A1(keyin[56]), .A2(n844), .Y(keyout[56]) );
  IBUFFX2_HVT U496 ( .A(keyin[118]), .Y(n1432) );
  MUX21X1_HVT U497 ( .A1(n1610), .A2(n1609), .S0(n1430), .Y(n2455) );
  INVX2_HVT U500 ( .A(keyin[118]), .Y(n1431) );
  IBUFFX2_HVT U502 ( .A(n1431), .Y(n1430) );
  MUX41X1_HVT U505 ( .A1(n2300), .A3(n2303), .A2(n2297), .A4(n2301), .S0(
        keyin[113]), .S1(n1433), .Y(n2296) );
  XNOR2X2_HVT U506 ( .A1(keyin[51]), .A2(n610), .Y(keyout[51]) );
  IBUFFX2_HVT U510 ( .A(n1755), .Y(keyout[19]) );
  MUX21X2_HVT U511 ( .A1(n2227), .A2(n2226), .S0(n597), .Y(n2115) );
  MUX41X1_HVT U512 ( .A1(n2348), .A3(n2362), .A2(n2343), .A4(n2354), .S0(n604), 
        .S1(n848), .Y(dummy[12]) );
  MUX41X1_HVT U514 ( .A1(n2238), .A3(n1186), .A2(n213), .A4(n1534), .S0(n1223), 
        .S1(n596), .Y(n2113) );
  XOR2X2_HVT U516 ( .A1(n1478), .A2(n1803), .Y(keyout[87]) );
  INVX2_HVT U520 ( .A(keyin[126]), .Y(n1416) );
  IBUFFX2_HVT U521 ( .A(n1416), .Y(n1415) );
  MUX41X1_HVT U522 ( .A1(n1534), .A3(n1521), .A2(n2233), .A4(n1491), .S0(n597), 
        .S1(n598), .Y(n2109) );
  NAND2X0_HVT U523 ( .A1(n2255), .A2(n823), .Y(n599) );
  NAND2X0_HVT U526 ( .A1(n2115), .A2(n1226), .Y(n600) );
  NAND2X0_HVT U527 ( .A1(n599), .A2(n600), .Y(n2114) );
  MUX41X1_HVT U530 ( .A1(n1600), .A3(n1561), .A2(n1215), .A4(n2459), .S0(n1433), .S1(n891), .Y(n2355) );
  NAND2X0_HVT U531 ( .A1(n2349), .A2(n601), .Y(n602) );
  NAND2X0_HVT U533 ( .A1(n2352), .A2(n1233), .Y(n603) );
  NAND2X0_HVT U535 ( .A1(n602), .A2(n603), .Y(n2348) );
  MUX41X1_HVT U536 ( .A1(n2344), .A3(n2346), .A2(n2345), .A4(n2347), .S0(n1231), .S1(n250), .Y(n2343) );
  NAND2X0_HVT U537 ( .A1(n2356), .A2(n1228), .Y(n605) );
  NAND2X0_HVT U538 ( .A1(n2355), .A2(n601), .Y(n606) );
  MUX21X1_HVT U539 ( .A1(n2359), .A2(n2360), .S0(n891), .Y(n2356) );
  XOR2X2_HVT U540 ( .A1(dummy[15]), .A2(keyin[15]), .Y(keyout[15]) );
  MUX41X1_HVT U541 ( .A1(n2413), .A3(n2423), .A2(n2417), .A4(n2427), .S0(n575), 
        .S1(keyin[113]), .Y(dummy[15]) );
  MUX21X1_HVT U542 ( .A1(n2424), .A2(n2426), .S0(n245), .Y(n2423) );
  MUX21X1_HVT U543 ( .A1(n2428), .A2(n2432), .S0(n245), .Y(n2427) );
  XOR2X1_HVT U544 ( .A1(dummy[15]), .A2(keyin[15]), .Y(n829) );
  INVX1_HVT U545 ( .A(n1439), .Y(n1438) );
  OA21X1_HVT U546 ( .A1(n2449), .A2(n1439), .A3(n1571), .Y(n2298) );
  INVX1_HVT U547 ( .A(keyin[112]), .Y(n1439) );
  INVX1_HVT U548 ( .A(n1469), .Y(n1466) );
  INVX1_HVT U549 ( .A(n1449), .Y(n1448) );
  INVX2_HVT U550 ( .A(keyin[109]), .Y(n1449) );
  INVX1_HVT U551 ( .A(keyin[29]), .Y(n845) );
  OA21X1_HVT U552 ( .A1(n2441), .A2(n1439), .A3(n2325), .Y(n2326) );
  NAND2X0_HVT U553 ( .A1(n2315), .A2(n601), .Y(n851) );
  MUX21X1_HVT U554 ( .A1(n1395), .A2(n1344), .S0(n1427), .Y(n2469) );
  INVX1_HVT U555 ( .A(n861), .Y(n1180) );
  MUX21X1_HVT U556 ( .A1(n1398), .A2(n1400), .S0(n1429), .Y(n2464) );
  INVX0_HVT U557 ( .A(n1153), .Y(n2551) );
  INVX1_HVT U558 ( .A(keyin[4]), .Y(n907) );
  INVX1_HVT U559 ( .A(n1366), .Y(n906) );
  INVX1_HVT U560 ( .A(keyin[68]), .Y(n1134) );
  NAND2X0_HVT U561 ( .A1(n1889), .A2(n587), .Y(n855) );
  XNOR3X1_HVT U562 ( .A1(n1814), .A2(keyin[97]), .A3(n1815), .Y(keyout[97]) );
  INVX2_HVT U563 ( .A(n1767), .Y(keyout[30]) );
  INVX0_HVT U564 ( .A(n1167), .Y(n822) );
  INVX0_HVT U565 ( .A(n1793), .Y(n1167) );
  INVX0_HVT U566 ( .A(n633), .Y(n2580) );
  INVX1_HVT U567 ( .A(n2581), .Y(n659) );
  INVX1_HVT U568 ( .A(n2552), .Y(n1154) );
  MUX21X1_HVT U569 ( .A1(n1640), .A2(n2561), .S0(n1164), .Y(n2560) );
  MUX21X1_HVT U570 ( .A1(n2096), .A2(n1389), .S0(n1208), .Y(n2095) );
  INVX1_HVT U571 ( .A(n2640), .Y(n1150) );
  INVX0_HVT U572 ( .A(n1132), .Y(n867) );
  MUX21X1_HVT U573 ( .A1(n1989), .A2(n1990), .S0(n1255), .Y(n1987) );
  OA21X1_HVT U574 ( .A1(n1213), .A2(n1468), .A3(n2009), .Y(n1867) );
  MUX21X1_HVT U575 ( .A1(n2420), .A2(n2418), .S0(n1433), .Y(n2417) );
  INVX1_HVT U576 ( .A(keyin[22]), .Y(n877) );
  MUX21X1_HVT U577 ( .A1(n2204), .A2(n2206), .S0(n1418), .Y(n2203) );
  NAND2X0_HVT U578 ( .A1(n2318), .A2(n592), .Y(n1176) );
  INVX0_HVT U579 ( .A(keyin[69]), .Y(n875) );
  INVX1_HVT U580 ( .A(n1820), .Y(n1133) );
  INVX1_HVT U581 ( .A(n821), .Y(keyout[105]) );
  INVX1_HVT U582 ( .A(n1784), .Y(n1130) );
  INVX0_HVT U583 ( .A(n1776), .Y(n1159) );
  INVX0_HVT U584 ( .A(n1752), .Y(keyout[16]) );
  INVX1_HVT U585 ( .A(n1758), .Y(keyout[22]) );
  INVX1_HVT U586 ( .A(n1764), .Y(keyout[28]) );
  INVX0_HVT U587 ( .A(keyin[33]), .Y(n888) );
  INVX1_HVT U588 ( .A(n1420), .Y(n823) );
  INVX1_HVT U589 ( .A(n1221), .Y(n849) );
  INVX1_HVT U590 ( .A(n1367), .Y(n878) );
  INVX1_HVT U591 ( .A(n1359), .Y(n1131) );
  INVX1_HVT U592 ( .A(keyin[127]), .Y(n876) );
  INVX1_HVT U593 ( .A(keyin[113]), .Y(n848) );
  XNOR2X2_HVT U594 ( .A1(n1753), .A2(n1797), .Y(keyout[81]) );
  INVX0_HVT U595 ( .A(n1361), .Y(n847) );
  INVX1_HVT U596 ( .A(n1453), .Y(n1452) );
  INVX0_HVT U597 ( .A(n1373), .Y(n1146) );
  INVX1_HVT U598 ( .A(n1425), .Y(n1424) );
  INVX1_HVT U599 ( .A(n1425), .Y(n828) );
  XNOR2X1_HVT U600 ( .A1(n1431), .A2(n1237), .Y(n1207) );
  INVX0_HVT U601 ( .A(n1253), .Y(n850) );
  NBUFFX2_HVT U602 ( .A(n1436), .Y(n1234) );
  INVX1_HVT U603 ( .A(n1746), .Y(keyout[10]) );
  INVX1_HVT U604 ( .A(n1747), .Y(keyout[11]) );
  MUX21X1_HVT U605 ( .A1(n659), .A2(n2667), .S0(n1449), .Y(n633) );
  XOR2X2_HVT U606 ( .A1(n1740), .A2(n1374), .Y(n2014) );
  XOR3X2_HVT U607 ( .A1(n1788), .A2(n862), .A3(n1777), .Y(keyout[104]) );
  XOR3X2_HVT U608 ( .A1(n1789), .A2(keyin[105]), .A3(n1778), .Y(n821) );
  MUX21X1_HVT U609 ( .A1(n1387), .A2(n1341), .S0(n1413), .Y(n2249) );
  MUX21X1_HVT U610 ( .A1(n1390), .A2(n1392), .S0(n1414), .Y(n2244) );
  INVX1_HVT U611 ( .A(n1749), .Y(keyout[13]) );
  XNOR2X2_HVT U612 ( .A1(n1749), .A2(n822), .Y(keyout[77]) );
  XNOR3X1_HVT U613 ( .A1(n1793), .A2(n297), .A3(n1749), .Y(keyout[109]) );
  MUX41X1_HVT U614 ( .A1(n2118), .A3(n2237), .A2(n1522), .A4(n1505), .S0(n866), 
        .S1(n823), .Y(n2117) );
  MUX41X1_HVT U615 ( .A1(n2120), .A3(n2122), .A2(n2117), .A4(n2119), .S0(
        keyin[125]), .S1(n1131), .Y(n2116) );
  XNOR2X1_HVT U616 ( .A1(n1747), .A2(n1791), .Y(keyout[75]) );
  IBUFFX2_HVT U617 ( .A(n1468), .Y(n843) );
  XNOR2X1_HVT U618 ( .A1(dummy[15]), .A2(keyin[15]), .Y(n1751) );
  IBUFFX2_HVT U619 ( .A(n1468), .Y(n1465) );
  INVX1_HVT U620 ( .A(n1748), .Y(keyout[12]) );
  INVX0_HVT U621 ( .A(n1458), .Y(n827) );
  MUX21X1_HVT U622 ( .A1(n1738), .A2(n1737), .S0(n1454), .Y(n2013) );
  XOR2X2_HVT U623 ( .A1(n1468), .A2(n2013), .Y(n1997) );
  XNOR2X1_HVT U624 ( .A1(keyin[24]), .A2(n595), .Y(n1760) );
  OA21X1_HVT U625 ( .A1(n2031), .A2(n1468), .A3(n1710), .Y(n1839) );
  XNOR2X2_HVT U626 ( .A1(n1758), .A2(n1802), .Y(keyout[86]) );
  XNOR2X2_HVT U627 ( .A1(n1754), .A2(keyin[50]), .Y(keyout[50]) );
  XNOR2X1_HVT U628 ( .A1(keyin[49]), .A2(n1753), .Y(keyout[49]) );
  IBUFFX2_HVT U629 ( .A(n1753), .Y(keyout[17]) );
  MUX41X1_HVT U633 ( .A1(n1511), .A3(n1391), .A2(n1515), .A4(n1338), .S0(n823), 
        .S1(n866), .Y(n2119) );
  IBUFFX2_HVT U634 ( .A(n1439), .Y(n830) );
  IBUFFX2_HVT U635 ( .A(n1439), .Y(n842) );
  XNOR2X1_HVT U636 ( .A1(n1777), .A2(n1788), .Y(keyout[72]) );
  INVX1_HVT U637 ( .A(n846), .Y(n2390) );
  XOR2X2_HVT U638 ( .A1(keyin[24]), .A2(dummy[24]), .Y(n844) );
  XOR2X2_HVT U639 ( .A1(dummy[29]), .A2(n845), .Y(n1765) );
  MUX21X1_HVT U640 ( .A1(n847), .A2(n1365), .S0(n1237), .Y(n846) );
  MUX41X1_HVT U642 ( .A1(n2385), .A3(n2374), .A2(n2379), .A4(n2370), .S0(n898), 
        .S1(n848), .Y(dummy[13]) );
  IBUFFX2_HVT U644 ( .A(n1425), .Y(n1423) );
  XOR2X1_HVT U645 ( .A1(n844), .A2(n1804), .Y(keyout[88]) );
  MUX21X2_HVT U646 ( .A1(n2309), .A2(n2310), .S0(n1233), .Y(n2308) );
  IBUFFX2_HVT U648 ( .A(n1750), .Y(keyout[14]) );
  INVX0_HVT U649 ( .A(n1207), .Y(n1173) );
  XNOR2X1_HVT U650 ( .A1(keyin[59]), .A2(n1763), .Y(keyout[59]) );
  INVX2_HVT U652 ( .A(n1765), .Y(keyout[29]) );
  XNOR3X1_HVT U653 ( .A1(n1809), .A2(n1418), .A3(n1765), .Y(keyout[125]) );
  XNOR3X1_HVT U654 ( .A1(n1804), .A2(n828), .A3(n1760), .Y(keyout[120]) );
  MUX41X1_HVT U655 ( .A1(n2034), .A3(n1994), .A2(n1951), .A4(n1722), .S0(n581), 
        .S1(n1464), .Y(n1950) );
  MUX41X1_HVT U656 ( .A1(n1943), .A3(n1950), .A2(n1942), .A4(n1945), .S0(
        keyin[103]), .S1(n850), .Y(n1941) );
  MUX41X1_HVT U657 ( .A1(n1847), .A3(n1845), .A2(n1846), .A4(n1842), .S0(n588), 
        .S1(n850), .Y(n1841) );
  MUX41X1_HVT U658 ( .A1(n2189), .A3(n2245), .A2(n1196), .A4(n2070), .S0(n823), 
        .S1(n866), .Y(n2069) );
  XNOR2X2_HVT U661 ( .A1(n1747), .A2(keyin[43]), .Y(keyout[43]) );
  NAND2X0_HVT U662 ( .A1(n2401), .A2(n592), .Y(n889) );
  NAND2X0_HVT U663 ( .A1(n2316), .A2(n1234), .Y(n852) );
  NAND2X0_HVT U664 ( .A1(n851), .A2(n852), .Y(n2314) );
  NAND2X0_HVT U666 ( .A1(n1941), .A2(keyin[97]), .Y(n902) );
  XNOR2X2_HVT U667 ( .A1(n1752), .A2(n1796), .Y(keyout[80]) );
  NAND2X0_HVT U668 ( .A1(n2075), .A2(n899), .Y(n871) );
  NAND2X0_HVT U669 ( .A1(n1952), .A2(n587), .Y(n853) );
  NAND2X0_HVT U670 ( .A1(n1962), .A2(keyin[97]), .Y(n854) );
  NAND2X0_HVT U671 ( .A1(n853), .A2(n854), .Y(dummy[30]) );
  NAND2X0_HVT U672 ( .A1(n2116), .A2(n867), .Y(n868) );
  NAND2X0_HVT U673 ( .A1(n1897), .A2(keyin[97]), .Y(n856) );
  NAND2X0_HVT U674 ( .A1(n855), .A2(n856), .Y(dummy[27]) );
  NAND2X0_HVT U675 ( .A1(n1858), .A2(keyin[97]), .Y(n857) );
  NAND2X0_HVT U677 ( .A1(n1849), .A2(n587), .Y(n858) );
  NAND2X0_HVT U679 ( .A1(n857), .A2(n858), .Y(dummy[25]) );
  MUX41X1_HVT U680 ( .A1(n2055), .A3(n2057), .A2(n2054), .A4(n2056), .S0(n1359), .S1(n1419), .Y(n2053) );
  OA21X1_HVT U684 ( .A1(n2229), .A2(n866), .A3(n1505), .Y(n2077) );
  NAND2X0_HVT U689 ( .A1(n1834), .A2(n587), .Y(n859) );
  NAND2X0_HVT U690 ( .A1(n1841), .A2(keyin[97]), .Y(n860) );
  NAND2X0_HVT U692 ( .A1(n859), .A2(n860), .Y(dummy[24]) );
  XOR2X1_HVT U694 ( .A1(n1433), .A2(n1431), .Y(n861) );
  IBUFFX2_HVT U696 ( .A(n1431), .Y(n1426) );
  XNOR2X1_HVT U698 ( .A1(n571), .A2(n1612), .Y(keyout[70]) );
  MUX21X1_HVT U699 ( .A1(n2657), .A2(n2628), .S0(n1164), .Y(n2627) );
  NAND2X0_HVT U700 ( .A1(n1404), .A2(n863), .Y(n864) );
  NAND2X0_HVT U702 ( .A1(n2610), .A2(n1209), .Y(n865) );
  NAND2X0_HVT U705 ( .A1(n864), .A2(n865), .Y(n2609) );
  INVX0_HVT U712 ( .A(n1209), .Y(n863) );
  MUX41X1_HVT U713 ( .A1(n2124), .A3(n2126), .A2(n2125), .A4(n2127), .S0(n1222), .S1(n279), .Y(n2123) );
  INVX2_HVT U714 ( .A(keyin[96]), .Y(n1468) );
  MUX41X1_HVT U715 ( .A1(n2074), .A3(n2071), .A2(n2073), .A4(n2069), .S0(n1131), .S1(n1419), .Y(n2068) );
  NAND2X0_HVT U716 ( .A1(n2108), .A2(n1132), .Y(n869) );
  NAND2X0_HVT U717 ( .A1(n868), .A2(n869), .Y(dummy[19]) );
  AO21X2_HVT U718 ( .A1(n1417), .A2(n1537), .A3(n866), .Y(n2161) );
  OA21X2_HVT U720 ( .A1(n2252), .A2(n866), .A3(n1515), .Y(n2062) );
  NAND2X0_HVT U721 ( .A1(n2068), .A2(n876), .Y(n872) );
  NAND2X0_HVT U722 ( .A1(n871), .A2(n872), .Y(dummy[17]) );
  NAND2X0_HVT U725 ( .A1(n2499), .A2(n1164), .Y(n873) );
  NAND2X0_HVT U726 ( .A1(n2500), .A2(n1242), .Y(n874) );
  NAND2X0_HVT U727 ( .A1(n873), .A2(n874), .Y(n2498) );
  INVX0_HVT U728 ( .A(n1813), .Y(n883) );
  MUX41X1_HVT U729 ( .A1(n2618), .A3(n2614), .A2(n2619), .A4(n2615), .S0(n1160), .S1(n298), .Y(n2613) );
  XOR3X2_HVT U731 ( .A1(n875), .A2(n1471), .A3(n887), .Y(keyout[69]) );
  XNOR2X1_HVT U732 ( .A1(keyin[54]), .A2(n1758), .Y(keyout[54]) );
  XNOR2X1_HVT U733 ( .A1(keyin[48]), .A2(n1752), .Y(keyout[48]) );
  MUX41X1_HVT U734 ( .A1(n1637), .A3(n2592), .A2(n2697), .A4(n1636), .S0(n1164), .S1(n457), .Y(n2591) );
  MUX21X1_HVT U735 ( .A1(n1365), .A2(n1362), .S0(n1433), .Y(n2364) );
  XOR2X2_HVT U736 ( .A1(dummy[22]), .A2(n877), .Y(n1758) );
  MUX41X1_HVT U738 ( .A1(n2632), .A3(n2627), .A2(n2623), .A4(n2622), .S0(n1161), .S1(n1160), .Y(n2621) );
  INVX1_HVT U739 ( .A(n1447), .Y(n1161) );
  NAND2X0_HVT U740 ( .A1(n2097), .A2(n899), .Y(n900) );
  MUX41X1_HVT U742 ( .A1(n2174), .A3(n2175), .A2(n2178), .A4(n2179), .S0(
        keyin[125]), .S1(keyin[121]), .Y(n2173) );
  XOR2X2_HVT U743 ( .A1(n1773), .A2(n887), .Y(keyout[37]) );
  NAND2X0_HVT U745 ( .A1(n2525), .A2(n878), .Y(n879) );
  NAND2X0_HVT U747 ( .A1(n2538), .A2(n1367), .Y(n880) );
  NAND2X0_HVT U750 ( .A1(n879), .A2(n880), .Y(dummy[2]) );
  XNOR2X2_HVT U752 ( .A1(n1815), .A2(n1814), .Y(keyout[65]) );
  INVX1_HVT U753 ( .A(n883), .Y(n884) );
  NAND2X0_HVT U754 ( .A1(n2494), .A2(n878), .Y(n885) );
  NAND2X0_HVT U756 ( .A1(n2501), .A2(n1367), .Y(n886) );
  NAND2X0_HVT U757 ( .A1(n885), .A2(n886), .Y(dummy[0]) );
  XOR2X2_HVT U758 ( .A1(n882), .A2(keyin[5]), .Y(n887) );
  NAND2X0_HVT U759 ( .A1(n2613), .A2(n878), .Y(n904) );
  XNOR2X2_HVT U761 ( .A1(keyout[1]), .A2(n888), .Y(keyout[33]) );
  NAND2X0_HVT U762 ( .A1(n2509), .A2(n878), .Y(n1151) );
  MUX21X1_HVT U763 ( .A1(n2361), .A2(n1553), .S0(n1433), .Y(n2360) );
  NAND2X0_HVT U765 ( .A1(n2393), .A2(n898), .Y(n890) );
  NAND2X0_HVT U766 ( .A1(n890), .A2(n889), .Y(dummy[14]) );
  XNOR2X2_HVT U767 ( .A1(n1778), .A2(n1789), .Y(keyout[73]) );
  IBUFFX2_HVT U768 ( .A(n1778), .Y(keyout[9]) );
  IBUFFX2_HVT U769 ( .A(n1777), .Y(keyout[8]) );
  XNOR2X2_HVT U771 ( .A1(n1161), .A2(n1446), .Y(n1182) );
  INVX1_HVT U772 ( .A(n1785), .Y(n1613) );
  NAND2X0_HVT U773 ( .A1(n2579), .A2(n892), .Y(n893) );
  NAND2X0_HVT U774 ( .A1(n2580), .A2(n249), .Y(n894) );
  NAND2X0_HVT U775 ( .A1(n893), .A2(n894), .Y(n2576) );
  NAND2X0_HVT U776 ( .A1(n1397), .A2(n861), .Y(n895) );
  NAND2X0_HVT U778 ( .A1(n2364), .A2(n1180), .Y(n896) );
  NAND2X0_HVT U779 ( .A1(n895), .A2(n896), .Y(n2363) );
  XNOR2X2_HVT U780 ( .A1(n1756), .A2(n1800), .Y(keyout[84]) );
  XNOR2X2_HVT U781 ( .A1(keyin[46]), .A2(n1750), .Y(keyout[46]) );
  XNOR2X2_HVT U783 ( .A1(keyin[40]), .A2(n1777), .Y(keyout[40]) );
  NAND2X0_HVT U786 ( .A1(n2084), .A2(n876), .Y(n901) );
  NAND2X0_HVT U788 ( .A1(n900), .A2(n901), .Y(dummy[18]) );
  INVX0_HVT U789 ( .A(n876), .Y(n899) );
  XNOR2X2_HVT U790 ( .A1(n1757), .A2(n1801), .Y(keyout[85]) );
  IBUFFX2_HVT U794 ( .A(n1757), .Y(keyout[21]) );
  NAND2X0_HVT U795 ( .A1(n1931), .A2(n587), .Y(n903) );
  NAND2X0_HVT U796 ( .A1(n902), .A2(n903), .Y(dummy[29]) );
  MUX41X1_HVT U800 ( .A1(n2685), .A3(n1662), .A2(n2663), .A4(n2524), .S0(n457), 
        .S1(n1164), .Y(n2523) );
  XOR2X2_HVT U804 ( .A1(n1781), .A2(n1780), .Y(keyout[5]) );
  INVX1_HVT U807 ( .A(n1148), .Y(n2637) );
  NAND2X0_HVT U808 ( .A1(n2621), .A2(n1367), .Y(n905) );
  NAND2X0_HVT U809 ( .A1(n904), .A2(n905), .Y(dummy[6]) );
  XNOR2X2_HVT U813 ( .A1(n1748), .A2(n1792), .Y(keyout[76]) );
  MUX21X1_HVT U815 ( .A1(n237), .A2(n1368), .S0(n1449), .Y(n2584) );
  MUX41X1_HVT U816 ( .A1(n2574), .A3(n2582), .A2(n2563), .A4(n2568), .S0(
        keyin[105]), .S1(n906), .Y(dummy[4]) );
  XOR3X1_HVT U817 ( .A1(n1134), .A2(n1146), .A3(n1147), .Y(keyout[100]) );
  XNOR2X2_HVT U818 ( .A1(n1784), .A2(n1785), .Y(n1147) );
  XOR2X2_HVT U819 ( .A1(dummy[4]), .A2(n907), .Y(n1785) );
  MUX21X1_HVT U823 ( .A1(n1358), .A2(n1357), .S0(n1419), .Y(n2144) );
  NAND2X0_HVT U824 ( .A1(n2135), .A2(n849), .Y(n908) );
  NAND2X0_HVT U825 ( .A1(n2136), .A2(n1225), .Y(n909) );
  NAND2X0_HVT U827 ( .A1(n908), .A2(n909), .Y(n2134) );
  MUX21X1_HVT U829 ( .A1(n2140), .A2(n2139), .S0(n1423), .Y(n2136) );
  MUX41X1_HVT U833 ( .A1(n1190), .A3(n2682), .A2(n2670), .A4(n1648), .S0(n457), 
        .S1(n1164), .Y(n2505) );
  NAND2X0_HVT U834 ( .A1(n2053), .A2(n876), .Y(n910) );
  NAND2X0_HVT U835 ( .A1(n2060), .A2(n867), .Y(n911) );
  NAND2X0_HVT U836 ( .A1(n910), .A2(n911), .Y(dummy[16]) );
  NAND2X0_HVT U839 ( .A1(n2181), .A2(n867), .Y(n912) );
  NAND2X0_HVT U840 ( .A1(n2173), .A2(n1132), .Y(n913) );
  NAND2X0_HVT U843 ( .A1(n912), .A2(n913), .Y(dummy[22]) );
  INVX1_HVT U844 ( .A(n1356), .Y(n1132) );
  MUX41X1_HVT U846 ( .A1(n2583), .A3(n2585), .A2(n2589), .A4(n2588), .S0(n517), 
        .S1(n1240), .Y(n2582) );
  NAND2X0_HVT U848 ( .A1(n1405), .A2(n914), .Y(n915) );
  NAND2X0_HVT U849 ( .A1(n2584), .A2(n1182), .Y(n938) );
  NAND2X0_HVT U850 ( .A1(n938), .A2(n915), .Y(n2583) );
  INVX0_HVT U851 ( .A(n1182), .Y(n914) );
  XNOR3X1_HVT U852 ( .A1(n1796), .A2(keyin[112]), .A3(n1752), .Y(keyout[112])
         );
  IBUFFX2_HVT U853 ( .A(n1759), .Y(keyout[23]) );
  INVX1_HVT U854 ( .A(n1759), .Y(n1478) );
  NAND2X0_HVT U855 ( .A1(n1389), .A2(n965), .Y(n1125) );
  NAND2X0_HVT U856 ( .A1(n2144), .A2(n1181), .Y(n1126) );
  NAND2X0_HVT U857 ( .A1(n1125), .A2(n1126), .Y(n2143) );
  INVX0_HVT U858 ( .A(n1181), .Y(n965) );
  OA21X1_HVT U859 ( .A1(n1514), .A2(n1419), .A3(n1499), .Y(n2148) );
  MUX41X1_HVT U860 ( .A1(n1641), .A3(n1407), .A2(n1646), .A4(n238), .S0(n1164), 
        .S1(n862), .Y(n2559) );
  XOR2X2_HVT U861 ( .A1(keyout[7]), .A2(keyin[39]), .Y(keyout[39]) );
  XOR3X2_HVT U862 ( .A1(n1134), .A2(n1130), .A3(n1613), .Y(keyout[68]) );
  XOR3X2_HVT U863 ( .A1(n1133), .A2(n1819), .A3(n1818), .Y(keyout[99]) );
  INVX1_HVT U864 ( .A(n2638), .Y(n1149) );
  XOR3X2_HVT U865 ( .A1(n884), .A2(n304), .A3(n1812), .Y(keyout[96]) );
  MUX21X1_HVT U866 ( .A1(n1150), .A2(n1149), .S0(n1449), .Y(n1148) );
  XNOR2X2_HVT U867 ( .A1(keyin[60]), .A2(n1764), .Y(keyout[60]) );
  MUX21X1_HVT U868 ( .A1(n1406), .A2(n2587), .S0(n862), .Y(n2547) );
  XOR2X1_HVT U869 ( .A1(keyin[2]), .A2(n881), .Y(n1816) );
  NAND2X0_HVT U870 ( .A1(n2516), .A2(n1367), .Y(n1152) );
  NAND2X0_HVT U871 ( .A1(n1151), .A2(n1152), .Y(dummy[1]) );
  MUX21X1_HVT U872 ( .A1(n2655), .A2(n2629), .S0(n249), .Y(n2552) );
  MUX21X1_HVT U873 ( .A1(n1155), .A2(n1154), .S0(n1164), .Y(n1153) );
  AO21X2_HVT U874 ( .A1(n1446), .A2(n1668), .A3(n457), .Y(n2601) );
  OA21X2_HVT U875 ( .A1(n1214), .A2(n249), .A3(n2672), .Y(n2529) );
  NAND2X0_HVT U876 ( .A1(n2569), .A2(n1164), .Y(n1156) );
  NAND2X0_HVT U877 ( .A1(n2572), .A2(n1242), .Y(n1157) );
  NAND2X0_HVT U878 ( .A1(n1156), .A2(n1157), .Y(n2568) );
  MUX21X1_HVT U879 ( .A1(n2662), .A2(n1664), .S0(n249), .Y(n2561) );
  XOR3X2_HVT U880 ( .A1(n1253), .A2(keyin[66]), .A3(n1158), .Y(keyout[98]) );
  XOR2X2_HVT U881 ( .A1(n1168), .A2(n1817), .Y(n1158) );
  XNOR2X2_HVT U882 ( .A1(n1159), .A2(n1819), .Y(keyout[3]) );
  NAND2X0_HVT U883 ( .A1(n2648), .A2(n1161), .Y(n1162) );
  NAND2X0_HVT U884 ( .A1(n2652), .A2(n297), .Y(n1163) );
  NAND2X0_HVT U885 ( .A1(n1162), .A2(n1163), .Y(n2647) );
  MUX21X1_HVT U886 ( .A1(n2650), .A2(n2651), .S0(n1245), .Y(n2648) );
  MUX21X2_HVT U887 ( .A1(n2546), .A2(n2547), .S0(n1164), .Y(n2544) );
  NAND2X0_HVT U888 ( .A1(n2549), .A2(n878), .Y(n1165) );
  NAND2X0_HVT U889 ( .A1(n2556), .A2(n1367), .Y(n1166) );
  NAND2X0_HVT U890 ( .A1(n1165), .A2(n1166), .Y(dummy[3]) );
  XNOR2X2_HVT U891 ( .A1(keyin[41]), .A2(n1778), .Y(keyout[41]) );
  OA21X2_HVT U892 ( .A1(n1211), .A2(n1439), .A3(n2452), .Y(n2309) );
  AO21X2_HVT U893 ( .A1(n1432), .A2(n1605), .A3(n1439), .Y(n2381) );
  XNOR2X1_HVT U894 ( .A1(n1440), .A2(n862), .Y(n1209) );
  IBUFFX2_HVT U895 ( .A(n1445), .Y(n1444) );
  XOR2X2_HVT U896 ( .A1(keyin[2]), .A2(dummy[2]), .Y(n1168) );
  MUX41X1_HVT U897 ( .A1(n2314), .A3(n2312), .A2(n2308), .A4(n2306), .S0(n1433), .S1(n848), .Y(n2305) );
  NAND2X0_HVT U898 ( .A1(n2317), .A2(n1173), .Y(n1169) );
  NAND2X0_HVT U899 ( .A1(n1397), .A2(n1207), .Y(n1170) );
  NAND2X0_HVT U900 ( .A1(n1169), .A2(n1170), .Y(n2316) );
  NAND2X0_HVT U901 ( .A1(n2329), .A2(n898), .Y(n1171) );
  NAND2X0_HVT U902 ( .A1(n2336), .A2(n604), .Y(n1172) );
  NAND2X0_HVT U903 ( .A1(n1171), .A2(n1172), .Y(dummy[11]) );
  NAND2X0_HVT U904 ( .A1(n1396), .A2(n1173), .Y(n1174) );
  NAND2X0_HVT U905 ( .A1(n2390), .A2(n1207), .Y(n1175) );
  NAND2X0_HVT U906 ( .A1(n1174), .A2(n1175), .Y(n2389) );
  NAND2X0_HVT U907 ( .A1(n2305), .A2(n898), .Y(n1177) );
  NAND2X0_HVT U908 ( .A1(n1177), .A2(n1176), .Y(dummy[10]) );
  XNOR2X2_HVT U909 ( .A1(keyin[53]), .A2(n1757), .Y(keyout[53]) );
  XNOR2X2_HVT U910 ( .A1(keyin[45]), .A2(n1749), .Y(keyout[45]) );
  MUX21X2_HVT U911 ( .A1(n2094), .A2(n2095), .S0(n1226), .Y(n2093) );
  XNOR2X1_HVT U912 ( .A1(keyin[42]), .A2(n1746), .Y(keyout[42]) );
  XOR2X2_HVT U913 ( .A1(keyout[10]), .A2(n1790), .Y(keyout[74]) );
  MUX21X1_HVT U914 ( .A1(n2208), .A2(n2212), .S0(n1418), .Y(n2207) );
  MUX21X1_HVT U915 ( .A1(n1573), .A2(n2451), .S0(n245), .Y(n2347) );
  MUX21X1_HVT U916 ( .A1(n1507), .A2(n2231), .S0(n589), .Y(n2127) );
  MUX21X1_HVT U917 ( .A1(n1552), .A2(n1579), .S0(n245), .Y(n2351) );
  MUX21X1_HVT U918 ( .A1(n1486), .A2(n1512), .S0(n589), .Y(n2131) );
  MUX21X1_HVT U919 ( .A1(n1202), .A2(n1568), .S0(n245), .Y(n2345) );
  MUX21X1_HVT U920 ( .A1(n1203), .A2(n1502), .S0(n290), .Y(n2125) );
  MUX21X2_HVT U921 ( .A1(n1379), .A2(n1925), .S0(n1179), .Y(n1924) );
  MUX21X2_HVT U922 ( .A1(n2591), .A2(n2593), .S0(n1448), .Y(n2590) );
  XOR2X1_HVT U923 ( .A1(n1779), .A2(keyin[36]), .Y(n1784) );
  XOR2X1_HVT U924 ( .A1(keyin[40]), .A2(keyin[72]), .Y(n1788) );
  XOR2X1_HVT U925 ( .A1(keyin[41]), .A2(keyin[73]), .Y(n1789) );
  XOR2X1_HVT U926 ( .A1(keyin[42]), .A2(keyin[74]), .Y(n1790) );
  XOR2X1_HVT U927 ( .A1(keyin[43]), .A2(keyin[75]), .Y(n1791) );
  XOR2X1_HVT U928 ( .A1(keyin[44]), .A2(keyin[76]), .Y(n1792) );
  XOR2X1_HVT U929 ( .A1(keyin[45]), .A2(keyin[77]), .Y(n1793) );
  XOR2X1_HVT U930 ( .A1(keyin[46]), .A2(keyin[78]), .Y(n1794) );
  XOR2X1_HVT U931 ( .A1(keyin[47]), .A2(keyin[79]), .Y(n1795) );
  XOR2X1_HVT U932 ( .A1(keyin[48]), .A2(keyin[80]), .Y(n1796) );
  XOR2X1_HVT U933 ( .A1(keyin[49]), .A2(keyin[81]), .Y(n1797) );
  XOR2X1_HVT U934 ( .A1(keyin[50]), .A2(keyin[82]), .Y(n1798) );
  XOR2X1_HVT U935 ( .A1(keyin[51]), .A2(keyin[83]), .Y(n1799) );
  XOR2X1_HVT U936 ( .A1(keyin[52]), .A2(keyin[84]), .Y(n1800) );
  XOR2X1_HVT U937 ( .A1(keyin[53]), .A2(keyin[85]), .Y(n1801) );
  XOR2X1_HVT U938 ( .A1(keyin[54]), .A2(keyin[86]), .Y(n1802) );
  XOR2X1_HVT U939 ( .A1(keyin[55]), .A2(keyin[87]), .Y(n1803) );
  XOR2X1_HVT U940 ( .A1(keyin[56]), .A2(keyin[88]), .Y(n1804) );
  XOR2X1_HVT U941 ( .A1(keyin[57]), .A2(keyin[89]), .Y(n1805) );
  XOR2X1_HVT U946 ( .A1(keyin[58]), .A2(keyin[90]), .Y(n1806) );
  MUX21X2_HVT U947 ( .A1(n1940), .A2(n1193), .S0(n1178), .Y(n1939) );
  INVX0_HVT U948 ( .A(n2693), .Y(n1669) );
  XNOR2X1_HVT U949 ( .A1(n589), .A2(n1415), .Y(n1181) );
  XOR2X2_HVT U950 ( .A1(n1769), .A2(keyin[34]), .Y(n1817) );
  XOR3X2_HVT U951 ( .A1(keyin[65]), .A2(keyin[33]), .A3(n1783), .Y(n1814) );
  XOR2X2_HVT U953 ( .A1(keyin[60]), .A2(keyin[92]), .Y(n1808) );
  XOR2X2_HVT U955 ( .A1(keyin[61]), .A2(keyin[93]), .Y(n1809) );
  XOR2X2_HVT U956 ( .A1(keyin[62]), .A2(keyin[94]), .Y(n1810) );
  XOR2X2_HVT U957 ( .A1(keyin[63]), .A2(keyin[95]), .Y(n1811) );
  XOR2X2_HVT U958 ( .A1(keyin[59]), .A2(keyin[91]), .Y(n1807) );
  INVX1_HVT U959 ( .A(n1380), .Y(n1735) );
  INVX1_HVT U961 ( .A(n2474), .Y(n1607) );
  INVX1_HVT U962 ( .A(n2694), .Y(n1670) );
  NBUFFX2_HVT U964 ( .A(n2032), .Y(n1380) );
  NBUFFX2_HVT U965 ( .A(n2032), .Y(n1381) );
  AND2X1_HVT U966 ( .A1(n1401), .A2(n2366), .Y(n1183) );
  MUX21X1_HVT U967 ( .A1(n1183), .A2(n1575), .S0(n1237), .Y(n2383) );
  MUX21X1_HVT U968 ( .A1(n1184), .A2(n545), .S0(n1227), .Y(n2163) );
  MUX21X1_HVT U969 ( .A1(n2464), .A2(n1183), .S0(n1237), .Y(n2384) );
  AND2X1_HVT U970 ( .A1(n1393), .A2(n2146), .Y(n1184) );
  AND2X1_HVT U972 ( .A1(n1397), .A2(n2409), .Y(n1185) );
  AND2X1_HVT U973 ( .A1(n1389), .A2(n2189), .Y(n1186) );
  AND2X1_HVT U974 ( .A1(n1606), .A2(n2421), .Y(n1187) );
  AND2X1_HVT U975 ( .A1(n1340), .A2(n2201), .Y(n1188) );
  AND2X1_HVT U976 ( .A1(n1410), .A2(n2586), .Y(n1189) );
  MUX21X1_HVT U978 ( .A1(n1704), .A2(n1903), .S0(n1247), .Y(n1902) );
  MUX21X1_HVT U979 ( .A1(n1729), .A2(n1383), .S0(n1259), .Y(n1903) );
  AND2X1_HVT U980 ( .A1(n272), .A2(n2641), .Y(n1190) );
  MUX21X1_HVT U981 ( .A1(n1690), .A2(n1734), .S0(n1254), .Y(n1973) );
  MUX21X1_HVT U982 ( .A1(n2684), .A2(n1189), .S0(n1451), .Y(n2604) );
  AND2X1_HVT U983 ( .A1(n1405), .A2(n2629), .Y(n1191) );
  MUX21X1_HVT U984 ( .A1(n1189), .A2(n1638), .S0(n1244), .Y(n2603) );
  AND2X1_HVT U985 ( .A1(n1984), .A2(n1351), .Y(n1192) );
  AND2X1_HVT U986 ( .A1(n1384), .A2(n1927), .Y(n1193) );
  AND2X1_HVT U987 ( .A1(n1378), .A2(n1967), .Y(n1194) );
  NBUFFX2_HVT U988 ( .A(n1739), .Y(n1353) );
  NBUFFX2_HVT U989 ( .A(n2254), .Y(n1386) );
  NBUFFX2_HVT U991 ( .A(n1739), .Y(n1351) );
  NBUFFX2_HVT U993 ( .A(n1606), .Y(n1342) );
  NBUFFX2_HVT U994 ( .A(n265), .Y(n1338) );
  NBUFFX2_HVT U998 ( .A(n1606), .Y(n1343) );
  NBUFFX2_HVT U999 ( .A(n265), .Y(n1340) );
  NBUFFX2_HVT U1003 ( .A(n265), .Y(n1339) );
  INVX1_HVT U1004 ( .A(n1399), .Y(n1605) );
  INVX1_HVT U1006 ( .A(n1391), .Y(n1537) );
  NBUFFX2_HVT U1008 ( .A(n2694), .Y(n1402) );
  NBUFFX2_HVT U1009 ( .A(n1669), .Y(n1347) );
  INVX1_HVT U1010 ( .A(n1382), .Y(n1734) );
  INVX1_HVT U1011 ( .A(n2480), .Y(n1609) );
  INVX1_HVT U1015 ( .A(n2260), .Y(n1540) );
  NAND2X0_HVT U1018 ( .A1(n1354), .A2(n1350), .Y(n2032) );
  NBUFFX2_HVT U1020 ( .A(n2474), .Y(n1395) );
  NBUFFX2_HVT U1027 ( .A(n2254), .Y(n1387) );
  INVX1_HVT U1028 ( .A(n2039), .Y(n1737) );
  NBUFFX2_HVT U1029 ( .A(n2694), .Y(n1403) );
  NBUFFX2_HVT U1030 ( .A(n1669), .Y(n1346) );
  INVX1_HVT U1031 ( .A(n1407), .Y(n1668) );
  INVX1_HVT U1033 ( .A(n1409), .Y(n1672) );
  MUX21X1_HVT U1034 ( .A1(n1342), .A2(n1584), .S0(n1235), .Y(n2315) );
  MUX21X1_HVT U1037 ( .A1(n1338), .A2(n1516), .S0(n1424), .Y(n2094) );
  MUX21X1_HVT U1038 ( .A1(n2435), .A2(n1593), .S0(n1237), .Y(n2388) );
  MUX21X1_HVT U1039 ( .A1(n2476), .A2(n2392), .S0(n1237), .Y(n2391) );
  MUX21X1_HVT U1041 ( .A1(n2215), .A2(n1525), .S0(n256), .Y(n2168) );
  MUX21X1_HVT U1043 ( .A1(n2341), .A2(n1577), .S0(n1234), .Y(n2340) );
  MUX21X1_HVT U1045 ( .A1(n1601), .A2(n2442), .S0(n830), .Y(n2341) );
  MUX21X1_HVT U1046 ( .A1(n2121), .A2(n1510), .S0(n1226), .Y(n2120) );
  MUX21X1_HVT U1047 ( .A1(n1533), .A2(n2222), .S0(n1424), .Y(n2121) );
  MUX21X1_HVT U1050 ( .A1(n2350), .A2(n2351), .S0(n247), .Y(n2349) );
  MUX21X1_HVT U1051 ( .A1(n238), .A2(n1647), .S0(n1244), .Y(n2535) );
  MUX21X1_HVT U1052 ( .A1(n2430), .A2(n2431), .S0(n247), .Y(n2428) );
  MUX21X1_HVT U1056 ( .A1(n2210), .A2(n2211), .S0(n256), .Y(n2208) );
  MUX21X1_HVT U1058 ( .A1(n2655), .A2(n1656), .S0(n892), .Y(n2608) );
  MUX21X1_HVT U1059 ( .A1(n2696), .A2(n2612), .S0(n1244), .Y(n2611) );
  XOR2X1_HVT U1060 ( .A1(n1426), .A2(n1605), .Y(n2436) );
  XOR2X1_HVT U1061 ( .A1(n1413), .A2(n1537), .Y(n2216) );
  MUX21X1_HVT U1063 ( .A1(n2570), .A2(n2571), .S0(n1245), .Y(n2569) );
  XOR2X1_HVT U1065 ( .A1(n1442), .A2(n1668), .Y(n2656) );
  MUX21X1_HVT U1066 ( .A1(n1705), .A2(n2025), .S0(n1250), .Y(n1940) );
  MUX21X1_HVT U1068 ( .A1(n1611), .A2(n1344), .S0(n566), .Y(n2361) );
  MUX21X1_HVT U1069 ( .A1(n1487), .A2(n2141), .S0(n589), .Y(n2140) );
  MUX21X1_HVT U1071 ( .A1(n1542), .A2(n1341), .S0(n569), .Y(n2141) );
  MUX21X1_HVT U1072 ( .A1(n1734), .A2(n1738), .S0(n1455), .Y(n1873) );
  MUX21X1_HVT U1073 ( .A1(n1735), .A2(n1738), .S0(n276), .Y(n1864) );
  MUX21X1_HVT U1076 ( .A1(n1349), .A2(n1385), .S0(n300), .Y(n1851) );
  MUX21X1_HVT U1077 ( .A1(n1384), .A2(n1378), .S0(n301), .Y(n1852) );
  MUX21X1_HVT U1082 ( .A1(n524), .A2(n1355), .S0(n1455), .Y(n1964) );
  MUX21X1_HVT U1083 ( .A1(n1737), .A2(n1352), .S0(n824), .Y(n1876) );
  XOR2X1_HVT U1084 ( .A1(n1377), .A2(n1457), .Y(n1992) );
  MUX21X1_HVT U1088 ( .A1(n1146), .A2(n1355), .S0(n824), .Y(n1848) );
  MUX21X1_HVT U1089 ( .A1(n1674), .A2(n234), .S0(n1444), .Y(n2581) );
  MUX21X1_HVT U1090 ( .A1(n2451), .A2(n2272), .S0(n1235), .Y(n2266) );
  MUX21X1_HVT U1091 ( .A1(n2231), .A2(n2051), .S0(n1227), .Y(n2045) );
  MUX21X1_HVT U1094 ( .A1(n1605), .A2(n1610), .S0(n567), .Y(n2321) );
  MUX21X1_HVT U1095 ( .A1(n1609), .A2(n1343), .S0(n568), .Y(n2323) );
  MUX21X1_HVT U1096 ( .A1(n1537), .A2(n1541), .S0(n570), .Y(n2100) );
  MUX21X1_HVT U1099 ( .A1(n219), .A2(n1339), .S0(n569), .Y(n2102) );
  MUX21X1_HVT U1100 ( .A1(n1401), .A2(n1398), .S0(n567), .Y(n2293) );
  MUX21X1_HVT U1103 ( .A1(n1393), .A2(n1390), .S0(n570), .Y(n2072) );
  MUX21X1_HVT U1108 ( .A1(n1513), .A2(n2257), .S0(n589), .Y(n2149) );
  MUX21X1_HVT U1109 ( .A1(n2186), .A2(n2185), .S0(n1226), .Y(n2183) );
  MUX21X1_HVT U1110 ( .A1(n1504), .A2(n2244), .S0(n1423), .Y(n2186) );
  MUX21X1_HVT U1114 ( .A1(n2463), .A2(n2378), .S0(n1234), .Y(n2377) );
  MUX21X1_HVT U1122 ( .A1(n1343), .A2(n1607), .S0(n566), .Y(n2378) );
  MUX21X1_HVT U1123 ( .A1(n1339), .A2(n1538), .S0(n569), .Y(n2158) );
  XOR2X1_HVT U1124 ( .A1(n1396), .A2(n1426), .Y(n2433) );
  XOR2X1_HVT U1125 ( .A1(n1388), .A2(n1415), .Y(n2213) );
  MUX21X1_HVT U1126 ( .A1(n1345), .A2(n1401), .S0(n568), .Y(n2291) );
  MUX21X1_HVT U1127 ( .A1(n1341), .A2(n1393), .S0(n569), .Y(n2070) );
  AND2X1_HVT U1130 ( .A1(n1430), .A2(n1610), .Y(n1195) );
  AND2X1_HVT U1131 ( .A1(n1413), .A2(n1541), .Y(n1196) );
  MUX21X1_HVT U1135 ( .A1(n1384), .A2(n1383), .S0(n1454), .Y(n2009) );
  MUX21X1_HVT U1137 ( .A1(n1379), .A2(n1383), .S0(n301), .Y(n2025) );
  MUX21X1_HVT U1138 ( .A1(n1352), .A2(n1350), .S0(n1455), .Y(n2023) );
  MUX21X1_HVT U1139 ( .A1(n2058), .A2(n2059), .S0(n1225), .Y(n2057) );
  MUX21X1_HVT U1140 ( .A1(n1527), .A2(n2225), .S0(n1227), .Y(n2059) );
  MUX21X1_HVT U1141 ( .A1(n1961), .A2(n1960), .S0(n1251), .Y(n1958) );
  MUX21X1_HVT U1146 ( .A1(n2019), .A2(n1383), .S0(n1259), .Y(n1961) );
  MUX21X1_HVT U1148 ( .A1(n2480), .A2(n1400), .S0(n1428), .Y(n2452) );
  MUX21X1_HVT U1149 ( .A1(n1737), .A2(n1735), .S0(n276), .Y(n2003) );
  MUX21X1_HVT U1151 ( .A1(n1737), .A2(n1350), .S0(n1455), .Y(n2006) );
  MUX21X1_HVT U1154 ( .A1(n524), .A2(n1738), .S0(n827), .Y(n2015) );
  MUX21X1_HVT U1155 ( .A1(n1380), .A2(n1385), .S0(n1457), .Y(n1946) );
  MUX21X1_HVT U1157 ( .A1(n1378), .A2(n1349), .S0(n1454), .Y(n2020) );
  MUX21X1_HVT U1158 ( .A1(n1381), .A2(n1349), .S0(n301), .Y(n2028) );
  MUX21X1_HVT U1160 ( .A1(n1381), .A2(n524), .S0(n300), .Y(n2004) );
  MUX21X1_HVT U1161 ( .A1(n1349), .A2(n1738), .S0(n276), .Y(n2000) );
  MUX21X1_HVT U1162 ( .A1(n1355), .A2(n1735), .S0(n1457), .Y(n2011) );
  MUX21X1_HVT U1163 ( .A1(n1395), .A2(n242), .S0(n1428), .Y(n2445) );
  MUX21X1_HVT U1164 ( .A1(n1386), .A2(n2253), .S0(n1412), .Y(n2225) );
  MUX21X1_HVT U1165 ( .A1(n1735), .A2(n1354), .S0(n301), .Y(n1825) );
  MUX21X1_HVT U1166 ( .A1(n1701), .A2(n2010), .S0(n1247), .Y(n1908) );
  MUX21X1_HVT U1167 ( .A1(n2475), .A2(n2335), .S0(n1234), .Y(n2334) );
  MUX21X1_HVT U1168 ( .A1(n1844), .A2(n1843), .S0(n1249), .Y(n1842) );
  MUX21X1_HVT U1169 ( .A1(n1688), .A2(n1732), .S0(n1259), .Y(n1844) );
  MUX21X1_HVT U1170 ( .A1(n1400), .A2(n1345), .S0(n566), .Y(n2269) );
  MUX21X1_HVT U1171 ( .A1(n1392), .A2(n1341), .S0(n569), .Y(n2048) );
  MUX21X1_HVT U1172 ( .A1(n1919), .A2(n1920), .S0(n1259), .Y(n1918) );
  MUX21X1_HVT U1173 ( .A1(n1679), .A2(n1707), .S0(n1247), .Y(n1920) );
  MUX21X1_HVT U1174 ( .A1(n1915), .A2(n1914), .S0(n1333), .Y(n1911) );
  MUX21X1_HVT U1175 ( .A1(n1682), .A2(n1916), .S0(n1251), .Y(n1915) );
  MUX21X1_HVT U1176 ( .A1(n1382), .A2(n1385), .S0(n1249), .Y(n1913) );
  MUX21X1_HVT U1177 ( .A1(n1354), .A2(n1349), .S0(n1455), .Y(n1916) );
  XOR2X1_HVT U1178 ( .A1(n300), .A2(n152), .Y(n1995) );
  MUX21X1_HVT U1179 ( .A1(n1383), .A2(n1354), .S0(n1456), .Y(n1969) );
  MUX21X1_HVT U1180 ( .A1(n1381), .A2(n1383), .S0(n1456), .Y(n1951) );
  MUX21X1_HVT U1181 ( .A1(n1351), .A2(n1735), .S0(n1455), .Y(n1944) );
  MUX21X1_HVT U1182 ( .A1(n1383), .A2(n1350), .S0(n276), .Y(n1829) );
  MUX21X1_HVT U1183 ( .A1(n1146), .A2(n524), .S0(n1457), .Y(n1827) );
  MUX21X1_HVT U1184 ( .A1(n2010), .A2(n1832), .S0(n1255), .Y(n1826) );
  MUX21X1_HVT U1185 ( .A1(n1541), .A2(n1540), .S0(n1415), .Y(n2235) );
  MUX21X1_HVT U1186 ( .A1(n1609), .A2(n1607), .S0(n1427), .Y(n2443) );
  MUX21X1_HVT U1187 ( .A1(n219), .A2(n1538), .S0(n1414), .Y(n2223) );
  MUX21X1_HVT U1188 ( .A1(n1343), .A2(n1344), .S0(n1427), .Y(n2462) );
  MUX21X1_HVT U1189 ( .A1(n1339), .A2(n1341), .S0(n1411), .Y(n2242) );
  MUX21X1_HVT U1190 ( .A1(n1609), .A2(n1345), .S0(n1430), .Y(n2449) );
  MUX21X1_HVT U1191 ( .A1(n1540), .A2(n1341), .S0(n1414), .Y(n2229) );
  MUX21X1_HVT U1192 ( .A1(n242), .A2(n1610), .S0(n1427), .Y(n2457) );
  MUX21X1_HVT U1193 ( .A1(n2253), .A2(n1541), .S0(n1412), .Y(n2237) );
  MUX21X1_HVT U1194 ( .A1(n1396), .A2(n1343), .S0(n1430), .Y(n2440) );
  MUX21X1_HVT U1195 ( .A1(n1388), .A2(n1339), .S0(n1412), .Y(n2220) );
  MUX21X1_HVT U1196 ( .A1(n1344), .A2(n1609), .S0(n1430), .Y(n2470) );
  MUX21X1_HVT U1197 ( .A1(n1341), .A2(n1540), .S0(n1414), .Y(n2250) );
  MUX21X1_HVT U1198 ( .A1(n1379), .A2(n1351), .S0(n276), .Y(n1999) );
  MUX21X1_HVT U1199 ( .A1(n1397), .A2(n1345), .S0(n1428), .Y(n2467) );
  MUX21X1_HVT U1200 ( .A1(n1389), .A2(n1341), .S0(n1412), .Y(n2247) );
  MUX21X1_HVT U1201 ( .A1(n1344), .A2(n1610), .S0(n1429), .Y(n2441) );
  MUX21X1_HVT U1202 ( .A1(n1341), .A2(n1541), .S0(n1414), .Y(n2221) );
  MUX21X1_HVT U1203 ( .A1(n1340), .A2(n219), .S0(n1413), .Y(n2252) );
  MUX21X1_HVT U1204 ( .A1(n1351), .A2(n1355), .S0(n1457), .Y(n1936) );
  MUX21X1_HVT U1205 ( .A1(n1981), .A2(n1983), .S0(n1249), .Y(n1980) );
  MUX21X1_HVT U1206 ( .A1(n1377), .A2(n1354), .S0(n1456), .Y(n1831) );
  MUX21X1_HVT U1207 ( .A1(n1395), .A2(n1400), .S0(n1428), .Y(n2392) );
  MUX21X1_HVT U1208 ( .A1(n1387), .A2(n1392), .S0(n1412), .Y(n2172) );
  MUX21X1_HVT U1209 ( .A1(n1539), .A2(n2253), .S0(n570), .Y(n2046) );
  MUX21X1_HVT U1210 ( .A1(n1400), .A2(n1342), .S0(n1428), .Y(n2372) );
  MUX21X1_HVT U1211 ( .A1(n1392), .A2(n1340), .S0(n1411), .Y(n2152) );
  XOR2X1_HVT U1212 ( .A1(n1404), .A2(n1443), .Y(n2653) );
  MUX21X1_HVT U1213 ( .A1(n1607), .A2(n1610), .S0(n1429), .Y(n2302) );
  MUX21X1_HVT U1214 ( .A1(n1538), .A2(n1541), .S0(n1415), .Y(n2081) );
  MUX21X1_HVT U1215 ( .A1(n1409), .A2(n1406), .S0(n1440), .Y(n2513) );
  MUX21X1_HVT U1216 ( .A1(n1345), .A2(n1611), .S0(n1426), .Y(n2288) );
  MUX21X1_HVT U1217 ( .A1(n1539), .A2(n1542), .S0(n1412), .Y(n2067) );
  MUX21X1_HVT U1218 ( .A1(n242), .A2(n1611), .S0(n567), .Y(n2400) );
  MUX21X1_HVT U1219 ( .A1(n2253), .A2(n1542), .S0(n570), .Y(n2180) );
  MUX21X1_HVT U1220 ( .A1(n524), .A2(n1734), .S0(n301), .Y(n1824) );
  MUX21X1_HVT U1221 ( .A1(n1345), .A2(n242), .S0(n568), .Y(n2267) );
  MUX21X1_HVT U1222 ( .A1(n2671), .A2(n2492), .S0(n1244), .Y(n2486) );
  MUX21X1_HVT U1223 ( .A1(n242), .A2(n1605), .S0(n568), .Y(n2264) );
  MUX21X1_HVT U1224 ( .A1(n2253), .A2(n1537), .S0(n569), .Y(n2043) );
  MUX21X1_HVT U1225 ( .A1(n1396), .A2(n1611), .S0(n567), .Y(n2271) );
  MUX21X1_HVT U1226 ( .A1(n1388), .A2(n1542), .S0(n569), .Y(n2050) );
  MUX21X1_HVT U1227 ( .A1(n1734), .A2(n1735), .S0(n827), .Y(n2021) );
  AND2X1_HVT U1228 ( .A1(n1440), .A2(n1673), .Y(n1197) );
  MUX21X1_HVT U1229 ( .A1(n1611), .A2(n1607), .S0(n1426), .Y(n2453) );
  MUX21X1_HVT U1230 ( .A1(n1542), .A2(n1538), .S0(n1413), .Y(n2233) );
  MUX21X1_HVT U1231 ( .A1(n1342), .A2(n1611), .S0(n567), .Y(n2380) );
  MUX21X1_HVT U1232 ( .A1(n1338), .A2(n1542), .S0(n570), .Y(n2160) );
  MUX21X1_HVT U1233 ( .A1(n1537), .A2(n1538), .S0(n1413), .Y(n2248) );
  MUX21X1_HVT U1234 ( .A1(n1658), .A2(n2665), .S0(n1244), .Y(n2500) );
  MUX21X1_HVT U1235 ( .A1(n1562), .A2(n1605), .S0(n1233), .Y(n2414) );
  MUX21X1_HVT U1236 ( .A1(n1496), .A2(n1537), .S0(n1225), .Y(n2194) );
  MUX21X1_HVT U1237 ( .A1(n2461), .A2(n1578), .S0(n245), .Y(n2344) );
  MUX21X1_HVT U1238 ( .A1(n2241), .A2(n1511), .S0(n289), .Y(n2124) );
  MUX21X1_HVT U1239 ( .A1(n1607), .A2(n1609), .S0(n1233), .Y(n2429) );
  MUX21X1_HVT U1240 ( .A1(n1538), .A2(n219), .S0(n1225), .Y(n2209) );
  MUX21X1_HVT U1241 ( .A1(n1668), .A2(n1673), .S0(n1442), .Y(n2541) );
  MUX21X1_HVT U1242 ( .A1(n1672), .A2(n1347), .S0(n1441), .Y(n2543) );
  MUX21X1_HVT U1243 ( .A1(n234), .A2(n1410), .S0(n1442), .Y(n2511) );
  MUX21X1_HVT U1244 ( .A1(n1605), .A2(n1607), .S0(n1429), .Y(n2468) );
  MUX21X1_HVT U1245 ( .A1(n1348), .A2(n1672), .S0(n1443), .Y(n2690) );
  MUX21X1_HVT U1246 ( .A1(n1405), .A2(n1348), .S0(n564), .Y(n2687) );
  MUX21X1_HVT U1247 ( .A1(n1643), .A2(n2697), .S0(n1447), .Y(n2589) );
  MUX21X1_HVT U1248 ( .A1(n1404), .A2(n1674), .S0(n1441), .Y(n2491) );
  MUX21X1_HVT U1249 ( .A1(n1197), .A2(n2597), .S0(n1244), .Y(n2596) );
  MUX21X1_HVT U1250 ( .A1(n2683), .A2(n2598), .S0(n1243), .Y(n2597) );
  MUX21X1_HVT U1251 ( .A1(n1347), .A2(n1670), .S0(n1444), .Y(n2598) );
  XOR2X1_HVT U1252 ( .A1(n2473), .A2(n1428), .Y(n2435) );
  XOR2X1_HVT U1253 ( .A1(n2253), .A2(n1414), .Y(n2215) );
  XOR2X1_HVT U1254 ( .A1(n1355), .A2(n301), .Y(n1996) );
  MUX21X1_HVT U1255 ( .A1(n1668), .A2(n1670), .S0(n1443), .Y(n2688) );
  XNOR2X1_HVT U1256 ( .A1(n1380), .A2(n1455), .Y(n1198) );
  XNOR2X1_HVT U1257 ( .A1(n1385), .A2(n1456), .Y(n1199) );
  MUX21X1_HVT U1259 ( .A1(n1673), .A2(n1672), .S0(n564), .Y(n2675) );
  MUX21X1_HVT U1261 ( .A1(n1672), .A2(n1670), .S0(n565), .Y(n2663) );
  MUX21X1_HVT U1262 ( .A1(n1347), .A2(n234), .S0(n1442), .Y(n2682) );
  MUX21X1_HVT U1263 ( .A1(n1406), .A2(n1408), .S0(n1443), .Y(n2684) );
  MUX21X1_HVT U1264 ( .A1(n1672), .A2(n234), .S0(n564), .Y(n2669) );
  MUX21X1_HVT U1265 ( .A1(n1395), .A2(n1401), .S0(n1430), .Y(n2386) );
  MUX21X1_HVT U1266 ( .A1(n1386), .A2(n1394), .S0(n1415), .Y(n2166) );
  MUX21X1_HVT U1267 ( .A1(n1353), .A2(n1737), .S0(n824), .Y(n2031) );
  MUX21X1_HVT U1268 ( .A1(n1402), .A2(n2693), .S0(n565), .Y(n2665) );
  MUX21X1_HVT U1269 ( .A1(n1403), .A2(n1348), .S0(n1443), .Y(n2689) );
  MUX21X1_HVT U1270 ( .A1(n1607), .A2(n1611), .S0(n1430), .Y(n2265) );
  MUX21X1_HVT U1271 ( .A1(n2695), .A2(n2555), .S0(n1243), .Y(n2554) );
  MUX21X1_HVT U1272 ( .A1(n2667), .A2(n2666), .S0(n1245), .Y(n2555) );
  MUX21X1_HVT U1273 ( .A1(n1625), .A2(n1668), .S0(n1242), .Y(n2634) );
  MUX21X1_HVT U1274 ( .A1(n2672), .A2(n2587), .S0(n1447), .Y(n2585) );
  MUX21X1_HVT U1275 ( .A1(n1396), .A2(n1395), .S0(n1429), .Y(n2263) );
  MUX21X1_HVT U1276 ( .A1(n1388), .A2(n1387), .S0(n1412), .Y(n2042) );
  MUX21X1_HVT U1277 ( .A1(n1377), .A2(n1381), .S0(n827), .Y(n1823) );
  MUX21X1_HVT U1278 ( .A1(n1408), .A2(n234), .S0(n1440), .Y(n2489) );
  MUX21X1_HVT U1280 ( .A1(n1670), .A2(n1672), .S0(n1242), .Y(n2649) );
  MUX21X1_HVT U1283 ( .A1(n1670), .A2(n1673), .S0(n565), .Y(n2522) );
  MUX21X1_HVT U1284 ( .A1(n1348), .A2(n1674), .S0(n565), .Y(n2508) );
  XNOR2X1_HVT U1285 ( .A1(n2480), .A2(n1429), .Y(n1200) );
  XNOR2X1_HVT U1286 ( .A1(n1393), .A2(n1411), .Y(n1201) );
  XOR2X1_HVT U1287 ( .A1(n1230), .A2(n1426), .Y(n2439) );
  XOR2X1_HVT U1288 ( .A1(n1221), .A2(n1412), .Y(n2219) );
  MUX21X1_HVT U1289 ( .A1(n1735), .A2(n1737), .S0(n1254), .Y(n1988) );
  XOR2X1_HVT U1290 ( .A1(n1457), .A2(n1253), .Y(n1998) );
  MUX21X1_HVT U1291 ( .A1(n1538), .A2(n1542), .S0(n1412), .Y(n2044) );
  XNOR2X1_HVT U1292 ( .A1(n1395), .A2(n1430), .Y(n1202) );
  XNOR2X1_HVT U1293 ( .A1(n1387), .A2(n1413), .Y(n1203) );
  MUX21X1_HVT U1294 ( .A1(n1409), .A2(n1408), .S0(n564), .Y(n2672) );
  MUX21X1_HVT U1295 ( .A1(n1404), .A2(n273), .S0(n565), .Y(n2660) );
  MUX21X1_HVT U1296 ( .A1(n1349), .A2(n1737), .S0(n1454), .Y(n2029) );
  MUX21X1_HVT U1297 ( .A1(n1348), .A2(n1673), .S0(n564), .Y(n2661) );
  MUX21X1_HVT U1298 ( .A1(n272), .A2(n1672), .S0(n1440), .Y(n2692) );
  MUX21X1_HVT U1299 ( .A1(n1346), .A2(n1674), .S0(n1442), .Y(n2600) );
  MUX21X1_HVT U1300 ( .A1(n2693), .A2(n1668), .S0(n1444), .Y(n2484) );
  MUX21X1_HVT U1302 ( .A1(n1616), .A2(n1642), .S0(n1447), .Y(n2571) );
  MUX21X1_HVT U1303 ( .A1(n2693), .A2(n1674), .S0(n1444), .Y(n2620) );
  MUX21X1_HVT U1305 ( .A1(n1674), .A2(n1670), .S0(n1440), .Y(n2673) );
  MUX21X1_HVT U1306 ( .A1(n2693), .A2(n1673), .S0(n1442), .Y(n2677) );
  MUX21X1_HVT U1307 ( .A1(n1636), .A2(n2671), .S0(n1447), .Y(n2567) );
  MUX21X1_HVT U1308 ( .A1(n1402), .A2(n1408), .S0(n565), .Y(n2612) );
  MUX21X1_HVT U1309 ( .A1(n1671), .A2(n2693), .S0(n1444), .Y(n2487) );
  MUX21X1_HVT U1310 ( .A1(n1408), .A2(n272), .S0(n565), .Y(n2592) );
  NBUFFX2_HVT U1311 ( .A(n2478), .Y(n1397) );
  NBUFFX2_HVT U1312 ( .A(n2258), .Y(n1389) );
  XOR2X1_HVT U1313 ( .A1(n1238), .A2(n1444), .Y(n2659) );
  NBUFFX2_HVT U1314 ( .A(n2478), .Y(n1396) );
  NBUFFX2_HVT U1316 ( .A(n2258), .Y(n1388) );
  NAND2X0_HVT U1318 ( .A1(n1341), .A2(n1542), .Y(n2254) );
  INVX0_HVT U1319 ( .A(n2473), .Y(n1606) );
  MUX21X1_HVT U1320 ( .A1(n1206), .A2(n1631), .S0(n1448), .Y(n2565) );
  MUX21X1_HVT U1321 ( .A1(n2681), .A2(n1641), .S0(n297), .Y(n2564) );
  NBUFFX2_HVT U1323 ( .A(n2698), .Y(n1405) );
  NBUFFX2_HVT U1324 ( .A(n2478), .Y(n1398) );
  NBUFFX2_HVT U1328 ( .A(n2258), .Y(n1390) );
  XOR2X1_HVT U1330 ( .A1(n2693), .A2(n1443), .Y(n2655) );
  XNOR2X1_HVT U1331 ( .A1(n1409), .A2(n1441), .Y(n1204) );
  AND2X1_HVT U1332 ( .A1(n1738), .A2(n300), .Y(n1205) );
  NBUFFX2_HVT U1334 ( .A(n2479), .Y(n1399) );
  NBUFFX2_HVT U1335 ( .A(n2259), .Y(n1391) );
  MUX21X1_HVT U1336 ( .A1(n1403), .A2(n1410), .S0(n1440), .Y(n2606) );
  MUX21X1_HVT U1337 ( .A1(n1404), .A2(n1403), .S0(n1441), .Y(n2483) );
  MUX21X1_HVT U1338 ( .A1(n2479), .A2(n1401), .S0(n245), .Y(n2358) );
  MUX21X1_HVT U1340 ( .A1(n2259), .A2(n1394), .S0(n1418), .Y(n2138) );
  NAND2X0_HVT U1341 ( .A1(n1348), .A2(n1674), .Y(n2694) );
  NBUFFX2_HVT U1342 ( .A(n2038), .Y(n1382) );
  MUX21X1_HVT U1344 ( .A1(n1670), .A2(n1674), .S0(n1441), .Y(n2485) );
  XNOR2X1_HVT U1345 ( .A1(n1402), .A2(n1440), .Y(n1206) );
  NBUFFX2_HVT U1346 ( .A(n2036), .Y(n1377) );
  NBUFFX2_HVT U1348 ( .A(n1740), .Y(n1355) );
  NBUFFX2_HVT U1350 ( .A(n2036), .Y(n1378) );
  NBUFFX2_HVT U1352 ( .A(n2698), .Y(n1406) );
  NBUFFX2_HVT U1354 ( .A(n2698), .Y(n1404) );
  NBUFFX2_HVT U1356 ( .A(n2699), .Y(n1407) );
  NBUFFX2_HVT U1358 ( .A(n2036), .Y(n1379) );
  NBUFFX2_HVT U1359 ( .A(n2479), .Y(n1400) );
  NBUFFX2_HVT U1360 ( .A(n2259), .Y(n1392) );
  NBUFFX2_HVT U1362 ( .A(n2038), .Y(n1383) );
  NBUFFX2_HVT U1364 ( .A(n1438), .Y(n1237) );
  NBUFFX2_HVT U1366 ( .A(n2480), .Y(n1401) );
  NBUFFX2_HVT U1368 ( .A(n2260), .Y(n1394) );
  NBUFFX2_HVT U1370 ( .A(n2039), .Y(n1385) );
  NBUFFX2_HVT U1372 ( .A(keyin[112]), .Y(n1236) );
  NBUFFX2_HVT U1374 ( .A(n1438), .Y(n1235) );
  NBUFFX2_HVT U1376 ( .A(n1424), .Y(n1227) );
  NBUFFX2_HVT U1377 ( .A(keyin[98]), .Y(n1254) );
  NBUFFX2_HVT U1379 ( .A(n2700), .Y(n1409) );
  NBUFFX2_HVT U1380 ( .A(n1467), .Y(n1333) );
  NBUFFX2_HVT U1381 ( .A(n1467), .Y(n1259) );
  MUX21X1_HVT U1382 ( .A1(n2699), .A2(n1410), .S0(n298), .Y(n2578) );
  NBUFFX2_HVT U1383 ( .A(n2260), .Y(n1393) );
  NBUFFX2_HVT U1384 ( .A(n1736), .Y(n1350) );
  NBUFFX2_HVT U1385 ( .A(keyin[98]), .Y(n1253) );
  NBUFFX2_HVT U1388 ( .A(n1467), .Y(n1255) );
  NBUFFX2_HVT U1389 ( .A(n1461), .Y(n1247) );
  NBUFFX2_HVT U1390 ( .A(n1736), .Y(n1349) );
  NBUFFX2_HVT U1391 ( .A(n2699), .Y(n1408) );
  NBUFFX2_HVT U1392 ( .A(n2039), .Y(n1384) );
  NBUFFX2_HVT U1393 ( .A(n1461), .Y(n1251) );
  NBUFFX2_HVT U1394 ( .A(n1608), .Y(n1344) );
  NBUFFX2_HVT U1395 ( .A(n1539), .Y(n1341) );
  NBUFFX2_HVT U1396 ( .A(n1608), .Y(n1345) );
  NBUFFX2_HVT U1397 ( .A(n1740), .Y(n1354) );
  NBUFFX2_HVT U1398 ( .A(n2700), .Y(n1410) );
  NBUFFX2_HVT U1399 ( .A(n1451), .Y(n1245) );
  NBUFFX2_HVT U1400 ( .A(n1461), .Y(n1250) );
  NBUFFX2_HVT U1401 ( .A(n1461), .Y(n1248) );
  NBUFFX2_HVT U1402 ( .A(n1463), .Y(n1252) );
  NBUFFX2_HVT U1403 ( .A(n1451), .Y(n1244) );
  NBUFFX2_HVT U1404 ( .A(n1251), .Y(n1246) );
  NBUFFX2_HVT U1405 ( .A(n1671), .Y(n1348) );
  XNOR2X1_HVT U1406 ( .A1(n1416), .A2(n1424), .Y(n1208) );
  MUX21X1_HVT U1407 ( .A1(n1357), .A2(n1542), .S0(n1424), .Y(n2170) );
  MUX21X1_HVT U1408 ( .A1(n2409), .A2(n2435), .S0(n842), .Y(n2332) );
  MUX21X1_HVT U1409 ( .A1(n2189), .A2(n2215), .S0(n1424), .Y(n2112) );
  MUX21X1_HVT U1410 ( .A1(n2327), .A2(n2326), .S0(n1233), .Y(n2324) );
  MUX21X1_HVT U1411 ( .A1(n2367), .A2(n1398), .S0(n250), .Y(n2327) );
  MUX21X1_HVT U1412 ( .A1(n2147), .A2(n1390), .S0(n1424), .Y(n2106) );
  MUX21X1_HVT U1413 ( .A1(n1368), .A2(n1674), .S0(n1451), .Y(n2610) );
  XOR2X1_HVT U1414 ( .A1(n1769), .A2(n1168), .Y(keyout[2]) );
  XOR2X1_HVT U1415 ( .A1(n1787), .A2(n1786), .Y(keyout[6]) );
  MUX21X1_HVT U1416 ( .A1(n1372), .A2(n1375), .S0(n1251), .Y(n1925) );
  MUX21X1_HVT U1417 ( .A1(n1708), .A2(n2037), .S0(n1251), .Y(n1930) );
  MUX21X1_HVT U1418 ( .A1(n2009), .A2(n1928), .S0(n1247), .Y(n1926) );
  MUX21X1_HVT U1419 ( .A1(n1372), .A2(n2035), .S0(n1254), .Y(n1990) );
  MUX21X1_HVT U1420 ( .A1(n1198), .A2(n1694), .S0(n1250), .Y(n1906) );
  MUX21X1_HVT U1421 ( .A1(n2479), .A2(n2311), .S0(n1237), .Y(n2310) );
  MUX21X1_HVT U1422 ( .A1(n2088), .A2(n2089), .S0(n1225), .Y(n2087) );
  MUX21X1_HVT U1423 ( .A1(n1392), .A2(n2090), .S0(n828), .Y(n2089) );
  MUX21X1_HVT U1424 ( .A1(n288), .A2(n1379), .S0(n1454), .Y(n2019) );
  MUX21X1_HVT U1425 ( .A1(n1997), .A2(n1971), .S0(n1249), .Y(n1970) );
  MUX21X1_HVT U1426 ( .A1(n1737), .A2(n1724), .S0(n1333), .Y(n1971) );
  MUX21X1_HVT U1427 ( .A1(n1400), .A2(n1611), .S0(n1430), .Y(n2411) );
  MUX21X1_HVT U1428 ( .A1(n2188), .A2(n2217), .S0(n1225), .Y(n2187) );
  XOR2X1_HVT U1429 ( .A1(n866), .A2(n2235), .Y(n2217) );
  MUX21X1_HVT U1437 ( .A1(n2191), .A2(n2190), .S0(n596), .Y(n2188) );
  MUX21X1_HVT U1442 ( .A1(n1392), .A2(n1542), .S0(n1411), .Y(n2191) );
  MUX21X1_HVT U1445 ( .A1(n2477), .A2(n1432), .S0(n245), .Y(n2357) );
  MUX21X1_HVT U1450 ( .A1(n2257), .A2(n1417), .S0(n290), .Y(n2137) );
  MUX21X1_HVT U1453 ( .A1(n1376), .A2(n1737), .S0(n824), .Y(n2005) );
  MUX21X1_HVT U1457 ( .A1(n1381), .A2(n1372), .S0(n1454), .Y(n2030) );
  MUX21X1_HVT U1458 ( .A1(n1364), .A2(n1609), .S0(n1428), .Y(n2446) );
  MUX21X1_HVT U1460 ( .A1(n1358), .A2(n1540), .S0(n1411), .Y(n2226) );
  MUX21X1_HVT U1467 ( .A1(n1350), .A2(n1375), .S0(n824), .Y(n2010) );
  MUX21X1_HVT U1474 ( .A1(n1373), .A2(n1735), .S0(n276), .Y(n2002) );
  MUX21X1_HVT U1475 ( .A1(n1735), .A2(n288), .S0(n1456), .Y(n2008) );
  MUX21X1_HVT U1476 ( .A1(n1938), .A2(n1704), .S0(n1250), .Y(n1935) );
  MUX21X1_HVT U1477 ( .A1(n1947), .A2(n1948), .S0(n1250), .Y(n1945) );
  MUX21X1_HVT U1478 ( .A1(n1377), .A2(n1949), .S0(n1210), .Y(n1948) );
  MUX21X1_HVT U1479 ( .A1(n1373), .A2(n1354), .S0(n1333), .Y(n1949) );
  MUX21X1_HVT U1480 ( .A1(n1887), .A2(n1888), .S0(n1250), .Y(n1885) );
  MUX21X1_HVT U1481 ( .A1(n1726), .A2(n152), .S0(n1333), .Y(n1888) );
  MUX21X1_HVT U1482 ( .A1(n1855), .A2(n1856), .S0(n1251), .Y(n1854) );
  MUX21X1_HVT U1483 ( .A1(n1954), .A2(n1373), .S0(n1259), .Y(n1856) );
  MUX21X1_HVT U1484 ( .A1(n2446), .A2(n2469), .S0(n1237), .Y(n2284) );
  MUX21X1_HVT U1485 ( .A1(n2063), .A2(n2062), .S0(n1226), .Y(n2061) );
  MUX21X1_HVT U1486 ( .A1(n2226), .A2(n2249), .S0(n828), .Y(n2063) );
  MUX21X1_HVT U1487 ( .A1(n1868), .A2(n1867), .S0(n1250), .Y(n1866) );
  MUX21X1_HVT U1488 ( .A1(n1383), .A2(n1724), .S0(n1333), .Y(n1868) );
  MUX21X1_HVT U1489 ( .A1(n1893), .A2(n1892), .S0(n1248), .Y(n1891) );
  MUX21X1_HVT U1490 ( .A1(n2011), .A2(n1685), .S0(n1259), .Y(n1893) );
  MUX21X1_HVT U1491 ( .A1(n1883), .A2(n1379), .S0(n1210), .Y(n1882) );
  MUX21X1_HVT U1492 ( .A1(n2003), .A2(n1727), .S0(n1259), .Y(n1881) );
  MUX21X1_HVT U1493 ( .A1(n1376), .A2(n1383), .S0(n1457), .Y(n1822) );
  MUX21X1_HVT U1494 ( .A1(n1342), .A2(n1361), .S0(n1429), .Y(n2458) );
  MUX21X1_HVT U1495 ( .A1(n1340), .A2(n1357), .S0(n1412), .Y(n2238) );
  MUX21X1_HVT U1496 ( .A1(n2474), .A2(n1362), .S0(n1426), .Y(n2471) );
  MUX21X1_HVT U1497 ( .A1(n1386), .A2(n1357), .S0(n1415), .Y(n2251) );
  MUX21X1_HVT U1498 ( .A1(n1376), .A2(n1734), .S0(n301), .Y(n2022) );
  MUX21X1_HVT U1499 ( .A1(n1365), .A2(n1398), .S0(n1426), .Y(n2460) );
  MUX21X1_HVT U1500 ( .A1(n1358), .A2(n1390), .S0(n1413), .Y(n2240) );
  MUX21X1_HVT U1501 ( .A1(n1361), .A2(n1607), .S0(n1429), .Y(n2444) );
  MUX21X1_HVT U1502 ( .A1(n1401), .A2(n1364), .S0(n1429), .Y(n2454) );
  MUX21X1_HVT U1503 ( .A1(n1394), .A2(n1358), .S0(n1415), .Y(n2234) );
  MUX21X1_HVT U1504 ( .A1(n1385), .A2(n288), .S0(n301), .Y(n2012) );
  MUX21X1_HVT U1505 ( .A1(n1373), .A2(n152), .S0(n300), .Y(n1828) );
  MUX21X1_HVT U1506 ( .A1(n2298), .A2(n2299), .S0(n1234), .Y(n2297) );
  MUX21X1_HVT U1507 ( .A1(n1582), .A2(n2474), .S0(n1236), .Y(n2299) );
  MUX21X1_HVT U1508 ( .A1(n213), .A2(n1386), .S0(n256), .Y(n2078) );
  MUX21X1_HVT U1509 ( .A1(n1692), .A2(n1458), .S0(n1254), .Y(n1975) );
  MUX21X1_HVT U1510 ( .A1(n1364), .A2(n1400), .S0(n568), .Y(n2262) );
  MUX21X1_HVT U1511 ( .A1(n1358), .A2(n1392), .S0(n570), .Y(n2041) );
  MUX21X1_HVT U1512 ( .A1(n1361), .A2(n1605), .S0(n568), .Y(n2268) );
  MUX21X1_HVT U1513 ( .A1(n1362), .A2(n2448), .S0(n1234), .Y(n2431) );
  MUX21X1_HVT U1514 ( .A1(n1357), .A2(n2228), .S0(n1226), .Y(n2211) );
  XOR2X1_HVT U1515 ( .A1(n1373), .A2(n824), .Y(n1993) );
  MUX21X1_HVT U1516 ( .A1(n1383), .A2(n1353), .S0(n827), .Y(n1933) );
  MUX21X1_HVT U1517 ( .A1(n1357), .A2(n1537), .S0(n570), .Y(n2047) );
  MUX21X1_HVT U1518 ( .A1(n1375), .A2(n524), .S0(n824), .Y(n1830) );
  NBUFFX2_HVT U1519 ( .A(n1422), .Y(n1226) );
  MUX21X1_HVT U1520 ( .A1(n1364), .A2(n1605), .S0(n1427), .Y(n2461) );
  MUX21X1_HVT U1521 ( .A1(n1358), .A2(n1537), .S0(n1411), .Y(n2241) );
  MUX21X1_HVT U1522 ( .A1(n1345), .A2(n1365), .S0(n1427), .Y(n2451) );
  MUX21X1_HVT U1523 ( .A1(n1341), .A2(n1358), .S0(n1414), .Y(n2231) );
  MUX21X1_HVT U1524 ( .A1(n1607), .A2(n1364), .S0(n1427), .Y(n2450) );
  MUX21X1_HVT U1525 ( .A1(n1538), .A2(n1358), .S0(n1415), .Y(n2230) );
  MUX21X1_HVT U1526 ( .A1(n2529), .A2(n2530), .S0(n1242), .Y(n2528) );
  MUX21X1_HVT U1527 ( .A1(n1408), .A2(n2531), .S0(n1451), .Y(n2530) );
  MUX21X1_HVT U1528 ( .A1(n1564), .A2(n1432), .S0(n1233), .Y(n2416) );
  MUX21X1_HVT U1529 ( .A1(n1498), .A2(n1417), .S0(n1225), .Y(n2196) );
  XNOR2X1_HVT U1530 ( .A1(n1468), .A2(n1454), .Y(n1210) );
  MUX21X1_HVT U1531 ( .A1(n1365), .A2(n242), .S0(n567), .Y(n2270) );
  MUX21X1_HVT U1532 ( .A1(n1358), .A2(n2253), .S0(n570), .Y(n2049) );
  NBUFFX2_HVT U1533 ( .A(n1436), .Y(n1233) );
  NBUFFX2_HVT U1534 ( .A(n1422), .Y(n1225) );
  MUX21X1_HVT U1535 ( .A1(n237), .A2(n1406), .S0(n1441), .Y(n2680) );
  MUX21X1_HVT U1536 ( .A1(n288), .A2(n1384), .S0(n276), .Y(n1821) );
  MUX21X1_HVT U1537 ( .A1(n1368), .A2(n2668), .S0(n1243), .Y(n2651) );
  MUX21X1_HVT U1538 ( .A1(n2697), .A2(n1446), .S0(n1447), .Y(n2577) );
  MUX21X1_HVT U1539 ( .A1(n237), .A2(n2693), .S0(n1442), .Y(n2490) );
  NBUFFX2_HVT U1540 ( .A(n1450), .Y(n1243) );
  MUX21X1_HVT U1541 ( .A1(n1402), .A2(n1368), .S0(n1441), .Y(n2691) );
  MUX21X1_HVT U1542 ( .A1(n237), .A2(n1668), .S0(n1441), .Y(n2681) );
  MUX21X1_HVT U1543 ( .A1(n1370), .A2(n1672), .S0(n564), .Y(n2666) );
  MUX21X1_HVT U1544 ( .A1(n1368), .A2(n1670), .S0(n565), .Y(n2664) );
  MUX21X1_HVT U1545 ( .A1(n2518), .A2(n2519), .S0(n1243), .Y(n2517) );
  MUX21X1_HVT U1546 ( .A1(n1645), .A2(n1402), .S0(n1245), .Y(n2519) );
  MUX21X1_HVT U1547 ( .A1(n1627), .A2(n1446), .S0(n1242), .Y(n2636) );
  MUX21X1_HVT U1548 ( .A1(n2631), .A2(n2630), .S0(n1245), .Y(n2628) );
  MUX21X1_HVT U1549 ( .A1(n1408), .A2(n1674), .S0(n564), .Y(n2631) );
  MUX21X1_HVT U1550 ( .A1(n2504), .A2(n2503), .S0(n1243), .Y(n2502) );
  MUX21X1_HVT U1551 ( .A1(n2666), .A2(n2689), .S0(n1451), .Y(n2504) );
  XOR2X1_HVT U1552 ( .A1(n1360), .A2(n1426), .Y(n2434) );
  XOR2X1_HVT U1553 ( .A1(keyin[124]), .A2(n1411), .Y(n2214) );
  MUX21X1_HVT U1554 ( .A1(n237), .A2(n1408), .S0(n1442), .Y(n2482) );
  MUX21X1_HVT U1555 ( .A1(n1365), .A2(n1401), .S0(n1426), .Y(n2261) );
  MUX21X1_HVT U1556 ( .A1(n1358), .A2(n1394), .S0(n1415), .Y(n2040) );
  NBUFFX2_HVT U1557 ( .A(keyin[106]), .Y(n1242) );
  MUX21X1_HVT U1558 ( .A1(n1346), .A2(n1368), .S0(n1441), .Y(n2678) );
  MUX21X1_HVT U1559 ( .A1(n1670), .A2(n237), .S0(n1441), .Y(n2670) );
  MUX21X1_HVT U1560 ( .A1(n1410), .A2(n1370), .S0(n1442), .Y(n2674) );
  MUX21X1_HVT U1561 ( .A1(n2037), .A2(n1459), .S0(n1249), .Y(n1912) );
  INVX1_HVT U1562 ( .A(keyin[99]), .Y(n1740) );
  NBUFFX2_HVT U1563 ( .A(n1436), .Y(n1232) );
  NBUFFX2_HVT U1564 ( .A(n1422), .Y(n1224) );
  MUX21X1_HVT U1565 ( .A1(n1348), .A2(n1370), .S0(n1443), .Y(n2671) );
  MUX21X1_HVT U1566 ( .A1(n1368), .A2(n1668), .S0(n1442), .Y(n2488) );
  NAND2X0_HVT U1567 ( .A1(n1611), .A2(n1362), .Y(n2478) );
  NAND2X0_HVT U1568 ( .A1(n1542), .A2(n1357), .Y(n2258) );
  INVX1_HVT U1569 ( .A(n1365), .Y(n1611) );
  INVX1_HVT U1570 ( .A(n1445), .Y(n1440) );
  INVX1_HVT U1571 ( .A(n1360), .Y(n1608) );
  MUX21X1_HVT U1572 ( .A1(n1370), .A2(n1410), .S0(n1444), .Y(n2481) );
  NAND2X0_HVT U1573 ( .A1(n1674), .A2(n1368), .Y(n2698) );
  NAND2X0_HVT U1574 ( .A1(n1363), .A2(n847), .Y(n2479) );
  NAND2X0_HVT U1575 ( .A1(keyin[123]), .A2(n1539), .Y(n2259) );
  INVX1_HVT U1576 ( .A(keyin[107]), .Y(n1674) );
  NAND2X0_HVT U1577 ( .A1(n1363), .A2(n1361), .Y(n2480) );
  NAND2X0_HVT U1578 ( .A1(keyin[123]), .A2(n1357), .Y(n2260) );
  NAND2X0_HVT U1579 ( .A1(n1375), .A2(n1736), .Y(n2038) );
  AND2X1_HVT U1580 ( .A1(n1606), .A2(n1432), .Y(n1211) );
  AND2X1_HVT U1581 ( .A1(n1340), .A2(n1417), .Y(n1212) );
  AND2X1_HVT U1582 ( .A1(n1353), .A2(n1459), .Y(n1213) );
  INVX1_HVT U1583 ( .A(keyin[108]), .Y(n1671) );
  INVX1_HVT U1584 ( .A(n1374), .Y(n1736) );
  NBUFFX2_HVT U1585 ( .A(n1450), .Y(n1241) );
  XOR2X1_HVT U1586 ( .A1(n233), .A2(n1444), .Y(n2654) );
  NAND2X0_HVT U1587 ( .A1(n1372), .A2(n1376), .Y(n2039) );
  NAND2X0_HVT U1588 ( .A1(n1373), .A2(n1355), .Y(n2036) );
  NAND2X0_HVT U1589 ( .A1(n1370), .A2(n1671), .Y(n2699) );
  AND2X1_HVT U1590 ( .A1(n272), .A2(n1446), .Y(n1214) );
  XOR2X1_HVT U1591 ( .A1(n1432), .A2(n1363), .Y(n2438) );
  XOR2X1_HVT U1592 ( .A1(n1417), .A2(n1358), .Y(n2218) );
  NAND2X0_HVT U1593 ( .A1(n237), .A2(n1368), .Y(n2700) );
  AND2X1_HVT U1594 ( .A1(n1432), .A2(n1345), .Y(n1215) );
  AND2X1_HVT U1595 ( .A1(n1417), .A2(n1341), .Y(n1216) );
  AND2X1_HVT U1596 ( .A1(n1446), .A2(n234), .Y(n1217) );
  NBUFFX2_HVT U1597 ( .A(n1435), .Y(n1230) );
  NBUFFX2_HVT U1598 ( .A(n1421), .Y(n1221) );
  NBUFFX2_HVT U1599 ( .A(keyin[98]), .Y(n1463) );
  XOR2X1_HVT U1600 ( .A1(n1446), .A2(n1370), .Y(n2658) );
  NBUFFX2_HVT U1601 ( .A(n1435), .Y(n1231) );
  NBUFFX2_HVT U1602 ( .A(n1421), .Y(n1222) );
  AND2X1_HVT U1603 ( .A1(n1350), .A2(n1459), .Y(n1218) );
  NBUFFX2_HVT U1604 ( .A(n1450), .Y(n1238) );
  NBUFFX2_HVT U1605 ( .A(n1421), .Y(n1223) );
  NBUFFX2_HVT U1606 ( .A(n1434), .Y(n1228) );
  NBUFFX2_HVT U1607 ( .A(n1434), .Y(n1229) );
  NBUFFX2_HVT U1608 ( .A(n1420), .Y(n1220) );
  NBUFFX2_HVT U1609 ( .A(n1420), .Y(n1219) );
  NBUFFX2_HVT U1610 ( .A(n1450), .Y(n1239) );
  NBUFFX2_HVT U1611 ( .A(n1450), .Y(n1240) );
  MUX21X1_HVT U1612 ( .A1(n2375), .A2(n2376), .S0(n245), .Y(n2374) );
  XOR2X1_HVT U1613 ( .A1(keyin[69]), .A2(n1461), .Y(n1743) );
  MUX21X1_HVT U1614 ( .A1(n2644), .A2(n2646), .S0(n297), .Y(n2643) );
  XNOR2X1_HVT U1615 ( .A1(keyin[67]), .A2(n1375), .Y(n1818) );
  NBUFFX2_HVT U1616 ( .A(keyin[114]), .Y(n1436) );
  NBUFFX2_HVT U1617 ( .A(keyin[122]), .Y(n1422) );
  NBUFFX2_HVT U1618 ( .A(keyin[100]), .Y(n1372) );
  NBUFFX2_HVT U1619 ( .A(keyin[115]), .Y(n1365) );
  NBUFFX2_HVT U1620 ( .A(keyin[116]), .Y(n1360) );
  NBUFFX2_HVT U1621 ( .A(keyin[115]), .Y(n1363) );
  NBUFFX2_HVT U1622 ( .A(keyin[116]), .Y(n1361) );
  NBUFFX2_HVT U1623 ( .A(keyin[124]), .Y(n1357) );
  NBUFFX2_HVT U1624 ( .A(keyin[100]), .Y(n1374) );
  NBUFFX2_HVT U1625 ( .A(keyin[107]), .Y(n1369) );
  NBUFFX2_HVT U1626 ( .A(keyin[116]), .Y(n1362) );
  NBUFFX2_HVT U1627 ( .A(keyin[108]), .Y(n1368) );
  INVX0_HVT U1628 ( .A(keyin[110]), .Y(n1446) );
  INVX0_HVT U1629 ( .A(keyin[102]), .Y(n1459) );
  NBUFFX2_HVT U1630 ( .A(keyin[99]), .Y(n1375) );
  NBUFFX2_HVT U1631 ( .A(n285), .Y(n1376) );
  NBUFFX2_HVT U1632 ( .A(keyin[115]), .Y(n1364) );
  NBUFFX2_HVT U1633 ( .A(keyin[123]), .Y(n1358) );
  NBUFFX2_HVT U1634 ( .A(keyin[114]), .Y(n1435) );
  NBUFFX2_HVT U1635 ( .A(keyin[122]), .Y(n1421) );
  NBUFFX2_HVT U1636 ( .A(keyin[100]), .Y(n1373) );
  NBUFFX2_HVT U1637 ( .A(keyin[106]), .Y(n1450) );
  NBUFFX2_HVT U1638 ( .A(keyin[107]), .Y(n1370) );
  NBUFFX2_HVT U1639 ( .A(keyin[114]), .Y(n1434) );
  NBUFFX2_HVT U1640 ( .A(keyin[122]), .Y(n1420) );
  NBUFFX2_HVT U1641 ( .A(keyin[103]), .Y(n1371) );
  NBUFFX2_HVT U1642 ( .A(keyin[121]), .Y(n1359) );
  NBUFFX2_HVT U1643 ( .A(keyin[127]), .Y(n1356) );
  NBUFFX2_HVT U1644 ( .A(keyin[111]), .Y(n1366) );
  NBUFFX2_HVT U1645 ( .A(keyin[111]), .Y(n1367) );
  XOR2X1_HVT U1646 ( .A1(n1776), .A2(keyin[35]), .Y(n1820) );
  XNOR2X1_HVT U1647 ( .A1(n1780), .A2(keyin[37]), .Y(n1773) );
  INVX0_HVT U1648 ( .A(n1772), .Y(n1470) );
  INVX0_HVT U1649 ( .A(n1773), .Y(n1471) );
  INVX0_HVT U1650 ( .A(n1771), .Y(n1472) );
  INVX0_HVT U1651 ( .A(round_num[1]), .Y(n1474) );
  INVX0_HVT U1652 ( .A(round_num[0]), .Y(n1475) );
  INVX0_HVT U1653 ( .A(round_num[3]), .Y(n1476) );
  INVX0_HVT U1654 ( .A(round_num[2]), .Y(n1477) );
  INVX0_HVT U1655 ( .A(n2239), .Y(n1484) );
  INVX0_HVT U1656 ( .A(n2236), .Y(n1485) );
  INVX0_HVT U1657 ( .A(n2228), .Y(n1486) );
  INVX0_HVT U1658 ( .A(n2227), .Y(n1487) );
  INVX0_HVT U1659 ( .A(n2218), .Y(n1488) );
  INVX0_HVT U1660 ( .A(n2086), .Y(n1489) );
  INVX0_HVT U1661 ( .A(n2052), .Y(n1490) );
  INVX0_HVT U1662 ( .A(n2257), .Y(n1491) );
  INVX0_HVT U1663 ( .A(n2243), .Y(n1492) );
  INVX0_HVT U1664 ( .A(n2255), .Y(n1493) );
  INVX0_HVT U1665 ( .A(n2256), .Y(n1494) );
  INVX0_HVT U1666 ( .A(n2252), .Y(n1495) );
  INVX0_HVT U1667 ( .A(n2251), .Y(n1496) );
  INVX0_HVT U1668 ( .A(n2249), .Y(n1498) );
  INVX0_HVT U1669 ( .A(n2248), .Y(n1499) );
  INVX0_HVT U1670 ( .A(n2247), .Y(n1500) );
  INVX0_HVT U1671 ( .A(n2242), .Y(n1502) );
  INVX0_HVT U1672 ( .A(n2241), .Y(n1503) );
  INVX0_HVT U1673 ( .A(n2240), .Y(n1504) );
  INVX0_HVT U1674 ( .A(n2238), .Y(n1505) );
  INVX0_HVT U1675 ( .A(n2237), .Y(n1506) );
  INVX0_HVT U1676 ( .A(n2234), .Y(n1507) );
  INVX0_HVT U1677 ( .A(n2233), .Y(n1508) );
  INVX0_HVT U1678 ( .A(n2231), .Y(n1509) );
  INVX0_HVT U1679 ( .A(n2045), .Y(n1510) );
  INVX0_HVT U1680 ( .A(n2230), .Y(n1511) );
  INVX0_HVT U1681 ( .A(n2229), .Y(n1512) );
  INVX0_HVT U1682 ( .A(n2226), .Y(n1513) );
  INVX0_HVT U1683 ( .A(n2225), .Y(n1514) );
  INVX0_HVT U1684 ( .A(n2223), .Y(n1515) );
  INVX0_HVT U1685 ( .A(n2222), .Y(n1516) );
  INVX0_HVT U1686 ( .A(n2221), .Y(n1517) );
  INVX0_HVT U1687 ( .A(n2220), .Y(n1518) );
  INVX0_HVT U1688 ( .A(n2189), .Y(n1519) );
  INVX0_HVT U1689 ( .A(n2246), .Y(n1520) );
  INVX0_HVT U1690 ( .A(n2201), .Y(n1521) );
  INVX0_HVT U1691 ( .A(n2146), .Y(n1522) );
  INVX0_HVT U1692 ( .A(n2051), .Y(n1523) );
  INVX0_HVT U1693 ( .A(n2104), .Y(n1524) );
  INVX0_HVT U1694 ( .A(n2050), .Y(n1525) );
  INVX0_HVT U1695 ( .A(n2049), .Y(n1526) );
  INVX0_HVT U1696 ( .A(n2047), .Y(n1528) );
  INVX0_HVT U1697 ( .A(n2046), .Y(n1529) );
  INVX0_HVT U1698 ( .A(n2166), .Y(n1530) );
  INVX0_HVT U1699 ( .A(n2160), .Y(n1531) );
  INVX0_HVT U1700 ( .A(n2044), .Y(n1532) );
  INVX0_HVT U1701 ( .A(n2043), .Y(n1533) );
  INVX0_HVT U1702 ( .A(n2042), .Y(n1534) );
  INVX0_HVT U1703 ( .A(n2041), .Y(n1535) );
  INVX0_HVT U1704 ( .A(n2040), .Y(n1536) );
  INVX0_HVT U1705 ( .A(n2459), .Y(n1550) );
  INVX0_HVT U1706 ( .A(n2456), .Y(n1551) );
  INVX0_HVT U1707 ( .A(n2448), .Y(n1552) );
  INVX0_HVT U1708 ( .A(n2447), .Y(n1553) );
  INVX0_HVT U1709 ( .A(n2438), .Y(n1554) );
  INVX0_HVT U1710 ( .A(n2307), .Y(n1555) );
  INVX0_HVT U1711 ( .A(n2273), .Y(n1556) );
  INVX0_HVT U1712 ( .A(n2477), .Y(n1557) );
  INVX0_HVT U1713 ( .A(n2463), .Y(n1558) );
  INVX0_HVT U1714 ( .A(n2475), .Y(n1559) );
  INVX0_HVT U1715 ( .A(n2476), .Y(n1560) );
  INVX0_HVT U1716 ( .A(n2472), .Y(n1561) );
  INVX0_HVT U1717 ( .A(n2471), .Y(n1562) );
  INVX0_HVT U1718 ( .A(n2470), .Y(n1563) );
  INVX0_HVT U1719 ( .A(n2469), .Y(n1564) );
  INVX0_HVT U1720 ( .A(n2468), .Y(n1565) );
  INVX0_HVT U1721 ( .A(n2467), .Y(n1566) );
  INVX0_HVT U1722 ( .A(n2464), .Y(n1567) );
  INVX0_HVT U1723 ( .A(n2462), .Y(n1568) );
  INVX0_HVT U1724 ( .A(n2461), .Y(n1569) );
  INVX0_HVT U1725 ( .A(n2460), .Y(n1570) );
  INVX0_HVT U1726 ( .A(n2458), .Y(n1571) );
  INVX0_HVT U1727 ( .A(n2457), .Y(n1572) );
  INVX0_HVT U1728 ( .A(n2454), .Y(n1573) );
  INVX0_HVT U1729 ( .A(n2453), .Y(n1574) );
  INVX0_HVT U1730 ( .A(n2452), .Y(n1575) );
  INVX0_HVT U1731 ( .A(n2451), .Y(n1576) );
  INVX0_HVT U1732 ( .A(n2266), .Y(n1577) );
  INVX0_HVT U1733 ( .A(n2450), .Y(n1578) );
  INVX0_HVT U1734 ( .A(n2449), .Y(n1579) );
  INVX0_HVT U1735 ( .A(n2446), .Y(n1580) );
  INVX0_HVT U1736 ( .A(n2445), .Y(n1581) );
  INVX0_HVT U1737 ( .A(n2444), .Y(n1582) );
  INVX0_HVT U1738 ( .A(n2443), .Y(n1583) );
  INVX0_HVT U1739 ( .A(n2442), .Y(n1584) );
  INVX0_HVT U1740 ( .A(n2441), .Y(n1585) );
  INVX0_HVT U1741 ( .A(n2440), .Y(n1586) );
  INVX0_HVT U1742 ( .A(n2409), .Y(n1587) );
  INVX0_HVT U1743 ( .A(n2466), .Y(n1588) );
  INVX0_HVT U1744 ( .A(n2421), .Y(n1589) );
  INVX0_HVT U1745 ( .A(n2366), .Y(n1590) );
  INVX0_HVT U1746 ( .A(n2272), .Y(n1591) );
  INVX0_HVT U1747 ( .A(n2325), .Y(n1592) );
  INVX0_HVT U1748 ( .A(n2271), .Y(n1593) );
  INVX0_HVT U1749 ( .A(n2270), .Y(n1594) );
  INVX0_HVT U1750 ( .A(n2269), .Y(n1595) );
  INVX0_HVT U1751 ( .A(n2268), .Y(n1596) );
  INVX0_HVT U1752 ( .A(n2267), .Y(n1597) );
  INVX0_HVT U1753 ( .A(n2386), .Y(n1598) );
  INVX0_HVT U1754 ( .A(n2380), .Y(n1599) );
  INVX0_HVT U1755 ( .A(n2265), .Y(n1600) );
  INVX0_HVT U1756 ( .A(n2264), .Y(n1601) );
  INVX0_HVT U1757 ( .A(n2263), .Y(n1602) );
  INVX0_HVT U1758 ( .A(n2262), .Y(n1603) );
  INVX0_HVT U1759 ( .A(n2261), .Y(n1604) );
  INVX0_HVT U1760 ( .A(n1396), .Y(n1610) );
  INVX0_HVT U1761 ( .A(n2679), .Y(n1614) );
  INVX0_HVT U1762 ( .A(n2676), .Y(n1615) );
  INVX0_HVT U1763 ( .A(n2668), .Y(n1616) );
  INVX0_HVT U1764 ( .A(n2658), .Y(n1617) );
  INVX0_HVT U1765 ( .A(n2527), .Y(n1618) );
  INVX0_HVT U1766 ( .A(n2493), .Y(n1619) );
  INVX0_HVT U1767 ( .A(n2697), .Y(n1620) );
  INVX0_HVT U1768 ( .A(n2683), .Y(n1621) );
  INVX0_HVT U1769 ( .A(n2695), .Y(n1622) );
  INVX0_HVT U1770 ( .A(n2696), .Y(n1623) );
  INVX0_HVT U1771 ( .A(n2692), .Y(n1624) );
  INVX0_HVT U1772 ( .A(n2691), .Y(n1625) );
  INVX0_HVT U1773 ( .A(n2690), .Y(n1626) );
  INVX0_HVT U1774 ( .A(n2689), .Y(n1627) );
  INVX0_HVT U1775 ( .A(n2688), .Y(n1628) );
  INVX0_HVT U1776 ( .A(n2687), .Y(n1629) );
  INVX0_HVT U1777 ( .A(n2684), .Y(n1630) );
  INVX0_HVT U1778 ( .A(n2682), .Y(n1631) );
  INVX0_HVT U1779 ( .A(n2681), .Y(n1632) );
  INVX0_HVT U1780 ( .A(n2680), .Y(n1633) );
  INVX0_HVT U1781 ( .A(n2678), .Y(n1634) );
  INVX0_HVT U1782 ( .A(n2677), .Y(n1635) );
  INVX0_HVT U1783 ( .A(n2674), .Y(n1636) );
  INVX0_HVT U1784 ( .A(n2673), .Y(n1637) );
  INVX0_HVT U1785 ( .A(n2672), .Y(n1638) );
  INVX0_HVT U1786 ( .A(n2671), .Y(n1639) );
  INVX0_HVT U1787 ( .A(n2486), .Y(n1640) );
  INVX0_HVT U1788 ( .A(n2670), .Y(n1641) );
  INVX0_HVT U1789 ( .A(n2669), .Y(n1642) );
  INVX0_HVT U1790 ( .A(n2666), .Y(n1643) );
  INVX0_HVT U1791 ( .A(n2665), .Y(n1644) );
  INVX0_HVT U1792 ( .A(n2664), .Y(n1645) );
  INVX0_HVT U1793 ( .A(n2663), .Y(n1646) );
  INVX0_HVT U1794 ( .A(n2662), .Y(n1647) );
  INVX0_HVT U1795 ( .A(n2661), .Y(n1648) );
  INVX0_HVT U1796 ( .A(n2660), .Y(n1649) );
  INVX0_HVT U1797 ( .A(n2629), .Y(n1650) );
  INVX0_HVT U1798 ( .A(n2686), .Y(n1651) );
  INVX0_HVT U1799 ( .A(n2641), .Y(n1652) );
  INVX0_HVT U1800 ( .A(n2586), .Y(n1653) );
  INVX0_HVT U1801 ( .A(n2492), .Y(n1654) );
  INVX0_HVT U1802 ( .A(n2545), .Y(n1655) );
  INVX0_HVT U1803 ( .A(n2491), .Y(n1656) );
  INVX0_HVT U1804 ( .A(n2490), .Y(n1657) );
  INVX0_HVT U1805 ( .A(n2489), .Y(n1658) );
  INVX0_HVT U1806 ( .A(n2488), .Y(n1659) );
  INVX0_HVT U1807 ( .A(n2487), .Y(n1660) );
  INVX0_HVT U1808 ( .A(n2606), .Y(n1661) );
  INVX0_HVT U1809 ( .A(n2600), .Y(n1662) );
  INVX0_HVT U1810 ( .A(n2485), .Y(n1663) );
  INVX0_HVT U1811 ( .A(n2484), .Y(n1664) );
  INVX0_HVT U1812 ( .A(n2483), .Y(n1665) );
  INVX0_HVT U1813 ( .A(n2482), .Y(n1666) );
  INVX0_HVT U1814 ( .A(n2481), .Y(n1667) );
  INVX0_HVT U1815 ( .A(n2035), .Y(n1679) );
  INVX0_HVT U1816 ( .A(n2018), .Y(n1680) );
  INVX0_HVT U1817 ( .A(n2016), .Y(n1681) );
  INVX0_HVT U1818 ( .A(n2007), .Y(n1682) );
  INVX0_HVT U1819 ( .A(n1870), .Y(n1683) );
  INVX0_HVT U1820 ( .A(n1833), .Y(n1684) );
  INVX0_HVT U1821 ( .A(n2037), .Y(n1685) );
  INVX0_HVT U1822 ( .A(n2024), .Y(n1686) );
  INVX0_HVT U1823 ( .A(n2033), .Y(n1687) );
  INVX0_HVT U1824 ( .A(n2034), .Y(n1688) );
  INVX0_HVT U1825 ( .A(n2031), .Y(n1689) );
  INVX0_HVT U1826 ( .A(n2030), .Y(n1690) );
  INVX0_HVT U1827 ( .A(n2029), .Y(n1691) );
  INVX0_HVT U1828 ( .A(n2028), .Y(n1692) );
  INVX0_HVT U1829 ( .A(n2025), .Y(n1693) );
  INVX0_HVT U1830 ( .A(n2023), .Y(n1694) );
  INVX0_HVT U1831 ( .A(n2022), .Y(n1695) );
  INVX0_HVT U1832 ( .A(n2021), .Y(n1696) );
  INVX0_HVT U1833 ( .A(n2020), .Y(n1697) );
  INVX0_HVT U1834 ( .A(n2019), .Y(n1698) );
  INVX0_HVT U1835 ( .A(n2017), .Y(n1699) );
  INVX0_HVT U1836 ( .A(n2015), .Y(n1700) );
  INVX0_HVT U1837 ( .A(n2012), .Y(n1701) );
  INVX0_HVT U1838 ( .A(n2011), .Y(n1702) );
  INVX0_HVT U1839 ( .A(n2010), .Y(n1703) );
  INVX0_HVT U1840 ( .A(n1826), .Y(n1704) );
  INVX0_HVT U1841 ( .A(n2009), .Y(n1705) );
  INVX0_HVT U1842 ( .A(n2008), .Y(n1706) );
  INVX0_HVT U1843 ( .A(n2006), .Y(n1707) );
  INVX0_HVT U1844 ( .A(n2005), .Y(n1708) );
  INVX0_HVT U1845 ( .A(n2004), .Y(n1709) );
  INVX0_HVT U1846 ( .A(n2003), .Y(n1710) );
  INVX0_HVT U1847 ( .A(n2002), .Y(n1711) );
  INVX0_HVT U1848 ( .A(n2001), .Y(n1712) );
  INVX0_HVT U1849 ( .A(n2000), .Y(n1713) );
  INVX0_HVT U1850 ( .A(n1999), .Y(n1714) );
  INVX0_HVT U1851 ( .A(n1996), .Y(n1715) );
  INVX0_HVT U1852 ( .A(n1967), .Y(n1716) );
  INVX0_HVT U1853 ( .A(n2027), .Y(n1717) );
  INVX0_HVT U1854 ( .A(n1927), .Y(n1718) );
  INVX0_HVT U1855 ( .A(n1832), .Y(n1719) );
  INVX0_HVT U1856 ( .A(n1984), .Y(n1720) );
  INVX0_HVT U1857 ( .A(n1886), .Y(n1721) );
  INVX0_HVT U1858 ( .A(n1831), .Y(n1722) );
  INVX0_HVT U1859 ( .A(n1830), .Y(n1723) );
  INVX0_HVT U1860 ( .A(n1829), .Y(n1724) );
  INVX0_HVT U1861 ( .A(n1828), .Y(n1725) );
  INVX0_HVT U1862 ( .A(n1827), .Y(n1726) );
  INVX0_HVT U1863 ( .A(n1946), .Y(n1727) );
  INVX0_HVT U1864 ( .A(n1936), .Y(n1728) );
  INVX0_HVT U1865 ( .A(n1825), .Y(n1729) );
  INVX0_HVT U1866 ( .A(n1824), .Y(n1730) );
  INVX0_HVT U1867 ( .A(n1823), .Y(n1731) );
  INVX0_HVT U1868 ( .A(n1822), .Y(n1732) );
  INVX0_HVT U1869 ( .A(n1821), .Y(n1733) );
endmodule

