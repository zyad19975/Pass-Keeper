
module inv_sbox_13 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n24, n196, n197, n198, n199, n200, n201, n202, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643;

  NAND2X0_HVT U3 ( .A1(n309), .A2(n319), .Y(n641) );
  NAND2X0_HVT U5 ( .A1(n640), .A2(n353), .Y(n639) );
  NAND2X0_HVT U7 ( .A1(n277), .A2(n354), .Y(n636) );
  NAND2X0_HVT U8 ( .A1(n363), .A2(n353), .Y(n635) );
  NAND2X0_HVT U9 ( .A1(n312), .A2(n635), .Y(n634) );
  NAND2X0_HVT U10 ( .A1(n313), .A2(n632), .Y(n633) );
  NAND2X0_HVT U11 ( .A1(n226), .A2(n359), .Y(n631) );
  NAND2X0_HVT U12 ( .A1(n363), .A2(n341), .Y(n630) );
  NAND2X0_HVT U13 ( .A1(n355), .A2(n267), .Y(n629) );
  NAND2X0_HVT U15 ( .A1(n350), .A2(n365), .Y(n627) );
  NAND2X0_HVT U19 ( .A1(n362), .A2(n432), .Y(n622) );
  NAND2X0_HVT U32 ( .A1(n342), .A2(n282), .Y(n611) );
  NAND2X0_HVT U35 ( .A1(n635), .A2(n433), .Y(n608) );
  NAND2X0_HVT U38 ( .A1(n341), .A2(n226), .Y(n605) );
  NAND2X0_HVT U42 ( .A1(n315), .A2(n433), .Y(n601) );
  OA21X1_HVT U53 ( .A1(n372), .A2(n593), .A3(n399), .Y(n591) );
  NAND2X0_HVT U55 ( .A1(n355), .A2(n640), .Y(n589) );
  MUX41X1_HVT U56 ( .A1(n412), .A3(n626), .A2(n397), .A4(n589), .S0(n334), 
        .S1(n369), .Y(n588) );
  AO21X1_HVT U60 ( .A1(n583), .A2(n337), .A3(n621), .Y(n584) );
  MUX41X1_HVT U62 ( .A1(n582), .A3(n588), .A2(n586), .A4(n590), .S0(n349), 
        .S1(n345), .Y(n581) );
  MUX41X1_HVT U65 ( .A1(n391), .A3(n393), .A2(n392), .A4(n605), .S0(n334), 
        .S1(n369), .Y(n578) );
  NAND2X0_HVT U66 ( .A1(n227), .A2(n327), .Y(n577) );
  MUX41X1_HVT U67 ( .A1(n388), .A3(n413), .A2(n390), .A4(n577), .S0(n339), 
        .S1(n331), .Y(n576) );
  MUX41X1_HVT U68 ( .A1(n388), .A3(n309), .A2(n389), .A4(n313), .S0(n333), 
        .S1(n283), .Y(n575) );
  MUX41X1_HVT U69 ( .A1(n575), .A3(n578), .A2(n576), .A4(n579), .S0(n349), 
        .S1(n345), .Y(n574) );
  NAND2X0_HVT U72 ( .A1(n351), .A2(n636), .Y(n572) );
  MUX41X1_HVT U73 ( .A1(n616), .A3(n572), .A2(n414), .A4(n340), .S0(n338), 
        .S1(n330), .Y(n571) );
  MUX41X1_HVT U74 ( .A1(n633), .A3(n404), .A2(n403), .A4(n394), .S0(n334), 
        .S1(n369), .Y(n570) );
  MUX41X1_HVT U78 ( .A1(n567), .A3(n571), .A2(n570), .A4(n573), .S0(n349), 
        .S1(n345), .Y(n566) );
  NAND2X0_HVT U81 ( .A1(n359), .A2(n636), .Y(n563) );
  AND2X1_HVT U82 ( .A1(n315), .A2(n355), .Y(n562) );
  MUX41X1_HVT U84 ( .A1(n325), .A3(n400), .A2(n418), .A4(n618), .S0(n334), 
        .S1(n283), .Y(n560) );
  MUX41X1_HVT U85 ( .A1(n560), .A3(n564), .A2(n561), .A4(n565), .S0(n349), 
        .S1(n345), .Y(n559) );
  MUX41X1_HVT U87 ( .A1(n378), .A3(n325), .A2(n419), .A4(n397), .S0(n332), 
        .S1(n369), .Y(n558) );
  MUX41X1_HVT U88 ( .A1(n390), .A3(n375), .A2(n613), .A4(n597), .S0(n333), 
        .S1(n235), .Y(n557) );
  NAND2X0_HVT U89 ( .A1(n282), .A2(n429), .Y(n556) );
  MUX41X1_HVT U96 ( .A1(n413), .A3(n629), .A2(n398), .A4(n420), .S0(n334), 
        .S1(n296), .Y(n549) );
  MUX41X1_HVT U99 ( .A1(n611), .A3(n392), .A2(n595), .A4(n626), .S0(n283), 
        .S1(n331), .Y(n546) );
  NAND2X0_HVT U100 ( .A1(n247), .A2(n428), .Y(n545) );
  MUX41X1_HVT U101 ( .A1(n422), .A3(n630), .A2(n310), .A4(n545), .S0(n283), 
        .S1(n330), .Y(n544) );
  AND2X1_HVT U104 ( .A1(n636), .A2(n352), .Y(n542) );
  MUX41X1_HVT U105 ( .A1(n628), .A3(n423), .A2(n563), .A4(n542), .S0(n334), 
        .S1(n235), .Y(n541) );
  MUX41X1_HVT U107 ( .A1(n422), .A3(n356), .A2(n540), .A4(n381), .S0(n333), 
        .S1(n235), .Y(n539) );
  MUX41X1_HVT U108 ( .A1(n394), .A3(n626), .A2(n397), .A4(n357), .S0(n334), 
        .S1(n235), .Y(n538) );
  MUX41X1_HVT U109 ( .A1(n421), .A3(n375), .A2(n418), .A4(n410), .S0(n333), 
        .S1(n368), .Y(n537) );
  AO21X1_HVT U112 ( .A1(n407), .A2(n338), .A3(n619), .Y(n534) );
  NAND2X0_HVT U114 ( .A1(n312), .A2(n636), .Y(n532) );
  MUX41X1_HVT U115 ( .A1(n532), .A3(n631), .A2(n407), .A4(n356), .S0(n283), 
        .S1(n331), .Y(n531) );
  NAND2X0_HVT U118 ( .A1(n226), .A2(n309), .Y(n528) );
  MUX41X1_HVT U119 ( .A1(n424), .A3(n529), .A2(n606), .A4(n528), .S0(n332), 
        .S1(n296), .Y(n527) );
  MUX41X1_HVT U122 ( .A1(n411), .A3(n321), .A2(n597), .A4(n415), .S0(n332), 
        .S1(n369), .Y(n525) );
  MUX41X1_HVT U124 ( .A1(n323), .A3(n524), .A2(n620), .A4(n306), .S0(n337), 
        .S1(n332), .Y(n523) );
  AOI21X1_HVT U127 ( .A1(n336), .A2(n519), .A3(n382), .Y(n520) );
  NAND2X0_HVT U129 ( .A1(n330), .A2(n312), .Y(n517) );
  MUX41X1_HVT U130 ( .A1(n517), .A3(n518), .A2(n521), .A4(n520), .S0(n339), 
        .S1(n347), .Y(n516) );
  AND2X1_HVT U131 ( .A1(n327), .A2(n366), .Y(n515) );
  MUX41X1_HVT U132 ( .A1(n379), .A3(n515), .A2(n426), .A4(n388), .S0(n338), 
        .S1(n336), .Y(n514) );
  MUX41X1_HVT U133 ( .A1(n427), .A3(n381), .A2(n589), .A4(n380), .S0(n337), 
        .S1(n330), .Y(n513) );
  MUX41X1_HVT U136 ( .A1(n594), .A3(n545), .A2(n511), .A4(n386), .S0(n335), 
        .S1(n296), .Y(n510) );
  MUX41X1_HVT U137 ( .A1(n267), .A3(n199), .A2(n618), .A4(n420), .S0(n339), 
        .S1(n330), .Y(n509) );
  MUX41X1_HVT U139 ( .A1(n508), .A3(n512), .A2(n516), .A4(n522), .S0(n349), 
        .S1(n307), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n403), .A3(n322), .A2(n396), .A4(n631), .S0(n338), 
        .S1(n331), .Y(n507) );
  NAND2X0_HVT U141 ( .A1(n350), .A2(n276), .Y(n506) );
  MUX41X1_HVT U142 ( .A1(n506), .A3(n604), .A2(n425), .A4(n396), .S0(n336), 
        .S1(n296), .Y(n505) );
  MUX41X1_HVT U143 ( .A1(n429), .A3(n408), .A2(n622), .A4(n620), .S0(n335), 
        .S1(n368), .Y(n504) );
  MUX41X1_HVT U145 ( .A1(n612), .A3(n423), .A2(n503), .A4(n563), .S0(n336), 
        .S1(n296), .Y(n502) );
  MUX41X1_HVT U146 ( .A1(n502), .A3(n504), .A2(n505), .A4(n507), .S0(n346), 
        .S1(n349), .Y(n501) );
  AO21X1_HVT U148 ( .A1(n339), .A2(n383), .A3(n428), .Y(n499) );
  MUX41X1_HVT U155 ( .A1(n396), .A3(n631), .A2(n623), .A4(n398), .S0(n335), 
        .S1(n272), .Y(n492) );
  NAND2X0_HVT U159 ( .A1(n488), .A2(n487), .Y(n489) );
  MUX41X1_HVT U162 ( .A1(n255), .A3(n393), .A2(n608), .A4(n485), .S0(n335), 
        .S1(n272), .Y(n484) );
  NAND2X0_HVT U163 ( .A1(n278), .A2(n429), .Y(n483) );
  MUX41X1_HVT U164 ( .A1(n634), .A3(n483), .A2(n606), .A4(n394), .S0(n332), 
        .S1(n369), .Y(n482) );
  NAND2X0_HVT U166 ( .A1(n632), .A2(n479), .Y(n480) );
  MUX41X1_HVT U172 ( .A1(n556), .A3(n474), .A2(n320), .A4(n258), .S0(n335), 
        .S1(n296), .Y(n473) );
  MUX41X1_HVT U173 ( .A1(n312), .A3(n431), .A2(n357), .A4(n607), .S0(n335), 
        .S1(n235), .Y(n472) );
  NAND2X0_HVT U177 ( .A1(n362), .A2(n309), .Y(n469) );
  AND2X1_HVT U179 ( .A1(n315), .A2(n352), .Y(n467) );
  MUX41X1_HVT U180 ( .A1(n611), .A3(n373), .A2(n467), .A4(n598), .S0(n335), 
        .S1(n368), .Y(n466) );
  MUX41X1_HVT U182 ( .A1(n381), .A3(n640), .A2(n378), .A4(n417), .S0(n332), 
        .S1(n283), .Y(n464) );
  MUX41X1_HVT U183 ( .A1(n408), .A3(n412), .A2(n394), .A4(n601), .S0(n337), 
        .S1(n331), .Y(n463) );
  AND2X1_HVT U185 ( .A1(n433), .A2(n366), .Y(n461) );
  NAND2X0_HVT U191 ( .A1(n372), .A2(n387), .Y(n455) );
  AND2X1_HVT U192 ( .A1(n404), .A2(n453), .Y(n454) );
  NAND2X0_HVT U194 ( .A1(n601), .A2(n453), .Y(n451) );
  MUX41X1_HVT U195 ( .A1(n452), .A3(n451), .A2(n454), .A4(n455), .S0(n333), 
        .S1(n346), .Y(n450) );
  NAND2X0_HVT U198 ( .A1(n361), .A2(n433), .Y(n632) );
  NAND2X0_HVT U200 ( .A1(n353), .A2(n247), .Y(n519) );
  NAND2X0_HVT U207 ( .A1(n282), .A2(n314), .Y(n583) );
  MUX41X1_HVT U1 ( .A1(n456), .A3(n450), .A2(n465), .A4(n462), .S0(n261), .S1(
        n240), .Y(out[7]) );
  NAND2X0_HVT U2 ( .A1(n325), .A2(n24), .Y(n196) );
  NAND2X0_HVT U4 ( .A1(n595), .A2(n339), .Y(n197) );
  NAND2X0_HVT U6 ( .A1(n196), .A2(n197), .Y(n459) );
  IBUFFX2_HVT U14 ( .A(n339), .Y(n24) );
  IBUFFX2_HVT U16 ( .A(n308), .Y(n240) );
  XOR2X1_HVT U17 ( .A1(n352), .A2(n365), .Y(n595) );
  OA21X1_HVT U18 ( .A1(n400), .A2(n371), .A3(n583), .Y(n457) );
  INVX0_HVT U20 ( .A(n614), .Y(n198) );
  INVX0_HVT U21 ( .A(n198), .Y(n199) );
  INVX1_HVT U22 ( .A(n444), .Y(n417) );
  INVX1_HVT U23 ( .A(n297), .Y(n247) );
  INVX1_HVT U24 ( .A(n366), .Y(n297) );
  MUX21X1_HVT U25 ( .A1(n325), .A2(n618), .S0(n299), .Y(n495) );
  MUX21X2_HVT U26 ( .A1(n351), .A2(n342), .S0(n364), .Y(n618) );
  INVX0_HVT U27 ( .A(n600), .Y(n408) );
  OR2X1_HVT U28 ( .A1(n200), .A2(n311), .Y(n637) );
  IBUFFX16_HVT U29 ( .A(n298), .Y(n200) );
  NAND2X0_HVT U30 ( .A1(n356), .A2(n201), .Y(n202) );
  NAND2X0_HVT U31 ( .A1(n342), .A2(n298), .Y(n218) );
  NAND2X0_HVT U33 ( .A1(n202), .A2(n218), .Y(n524) );
  IBUFFX2_HVT U34 ( .A(n298), .Y(n201) );
  NAND2X0_HVT U36 ( .A1(n525), .A2(n219), .Y(n220) );
  NAND2X0_HVT U37 ( .A1(n523), .A2(n224), .Y(n221) );
  NAND2X0_HVT U39 ( .A1(n220), .A2(n221), .Y(n522) );
  INVX0_HVT U40 ( .A(n224), .Y(n219) );
  NBUFFX4_HVT U41 ( .A(n434), .Y(n343) );
  INVX0_HVT U43 ( .A(n366), .Y(n298) );
  IBUFFX2_HVT U44 ( .A(n346), .Y(n224) );
  INVX1_HVT U45 ( .A(n371), .Y(n368) );
  IBUFFX2_HVT U46 ( .A(n371), .Y(n369) );
  INVX1_HVT U47 ( .A(n299), .Y(n272) );
  INVX0_HVT U48 ( .A(in[4]), .Y(n371) );
  INVX1_HVT U49 ( .A(n287), .Y(n261) );
  NBUFFX2_HVT U50 ( .A(n434), .Y(n222) );
  INVX0_HVT U51 ( .A(in[6]), .Y(n434) );
  NBUFFX2_HVT U52 ( .A(n434), .Y(n342) );
  INVX1_HVT U54 ( .A(n222), .Y(n319) );
  INVX0_HVT U57 ( .A(n364), .Y(n282) );
  INVX0_HVT U58 ( .A(n366), .Y(n361) );
  MUX41X1_HVT U59 ( .A1(n401), .A3(n562), .A2(n563), .A4(n417), .S0(n223), 
        .S1(n369), .Y(n561) );
  IBUFFX16_HVT U61 ( .A(n333), .Y(n223) );
  INVX1_HVT U63 ( .A(n366), .Y(n363) );
  MUX21X2_HVT U64 ( .A1(n400), .A2(n406), .S0(n271), .Y(n269) );
  MUX21X1_HVT U70 ( .A1(n316), .A2(n640), .S0(n330), .Y(n580) );
  AO21X1_HVT U71 ( .A1(n351), .A2(n640), .A3(n372), .Y(n479) );
  INVX1_HVT U75 ( .A(n366), .Y(n362) );
  INVX1_HVT U76 ( .A(in[5]), .Y(n230) );
  INVX1_HVT U77 ( .A(n348), .Y(n228) );
  XOR2X2_HVT U79 ( .A1(n343), .A2(n236), .Y(n626) );
  MUX41X1_HVT U80 ( .A1(n459), .A3(n458), .A2(n460), .A4(n457), .S0(n304), 
        .S1(n225), .Y(n456) );
  IBUFFX16_HVT U83 ( .A(n305), .Y(n225) );
  INVX1_HVT U86 ( .A(n298), .Y(n226) );
  INVX2_HVT U90 ( .A(n226), .Y(n227) );
  MUX41X1_HVT U91 ( .A1(n551), .A3(n557), .A2(n555), .A4(n558), .S0(n228), 
        .S1(n229), .Y(n550) );
  IBUFFX16_HVT U92 ( .A(n304), .Y(n229) );
  INVX1_HVT U93 ( .A(n621), .Y(n394) );
  INVX0_HVT U94 ( .A(n258), .Y(n316) );
  MUX41X1_HVT U95 ( .A1(n533), .A3(n530), .A2(n531), .A4(n527), .S0(n230), 
        .S1(n231), .Y(n526) );
  IBUFFX16_HVT U97 ( .A(n347), .Y(n231) );
  INVX0_HVT U98 ( .A(n366), .Y(n364) );
  MUX21X1_HVT U102 ( .A1(n382), .A2(n602), .S0(n339), .Y(n535) );
  NAND2X0_HVT U103 ( .A1(n568), .A2(n232), .Y(n233) );
  NAND2X0_HVT U106 ( .A1(n569), .A2(n245), .Y(n234) );
  NAND2X0_HVT U110 ( .A1(n233), .A2(n234), .Y(n567) );
  INVX0_HVT U111 ( .A(n245), .Y(n232) );
  IBUFFX2_HVT U113 ( .A(n336), .Y(n245) );
  NBUFFX2_HVT U116 ( .A(n368), .Y(n235) );
  AO21X2_HVT U117 ( .A1(n366), .A2(n313), .A3(n372), .Y(n487) );
  INVX1_HVT U120 ( .A(n430), .Y(n236) );
  INVX1_HVT U121 ( .A(n643), .Y(n311) );
  NAND2X0_HVT U123 ( .A1(n574), .A2(n237), .Y(n238) );
  NAND2X0_HVT U125 ( .A1(n581), .A2(n307), .Y(n239) );
  NAND2X0_HVT U126 ( .A1(n238), .A2(n239), .Y(out[0]) );
  IBUFFX2_HVT U128 ( .A(n307), .Y(n237) );
  NAND2X0_HVT U134 ( .A1(n489), .A2(n241), .Y(n242) );
  NAND2X0_HVT U135 ( .A1(n490), .A2(n336), .Y(n243) );
  NAND2X0_HVT U138 ( .A1(n242), .A2(n243), .Y(n486) );
  IBUFFX2_HVT U144 ( .A(n336), .Y(n241) );
  MUX21X1_HVT U147 ( .A1(n600), .A2(n415), .S0(n338), .Y(n490) );
  MUX21X1_HVT U149 ( .A1(n340), .A2(n432), .S0(n361), .Y(n600) );
  NAND2X1_HVT U150 ( .A1(n501), .A2(in[7]), .Y(n300) );
  MUX21X2_HVT U151 ( .A1(n591), .A2(n592), .S0(n244), .Y(n590) );
  IBUFFX16_HVT U152 ( .A(n335), .Y(n244) );
  INVX2_HVT U153 ( .A(n337), .Y(n299) );
  OA21X2_HVT U154 ( .A1(n376), .A2(n372), .A3(n385), .Y(n494) );
  OA21X2_HVT U156 ( .A1(n377), .A2(n372), .A3(n621), .Y(n568) );
  AO21X2_HVT U157 ( .A1(n361), .A2(n428), .A3(n371), .Y(n453) );
  INVX0_HVT U158 ( .A(n350), .Y(n259) );
  INVX0_HVT U160 ( .A(n341), .Y(n246) );
  NBUFFX4_HVT U161 ( .A(n430), .Y(n341) );
  INVX0_HVT U165 ( .A(n357), .Y(n260) );
  IBUFFX4_HVT U167 ( .A(n337), .Y(n256) );
  OR2X1_HVT U168 ( .A1(n343), .A2(n246), .Y(n638) );
  IBUFFX2_HVT U169 ( .A(n343), .Y(n327) );
  MUX21X1_HVT U170 ( .A1(n327), .A2(n353), .S0(n247), .Y(n614) );
  INVX2_HVT U171 ( .A(n276), .Y(n278) );
  MUX21X2_HVT U174 ( .A1(n514), .A2(n513), .S0(n248), .Y(n512) );
  IBUFFX16_HVT U175 ( .A(n347), .Y(n248) );
  NAND2X0_HVT U176 ( .A1(n363), .A2(n358), .Y(n640) );
  NAND2X0_HVT U178 ( .A1(n480), .A2(n249), .Y(n250) );
  NAND2X0_HVT U181 ( .A1(n481), .A2(n331), .Y(n251) );
  NAND2X0_HVT U184 ( .A1(n250), .A2(n251), .Y(n478) );
  IBUFFX2_HVT U186 ( .A(n331), .Y(n249) );
  MUX21X1_HVT U187 ( .A1(n617), .A2(n620), .S0(n337), .Y(n481) );
  INVX1_HVT U188 ( .A(n617), .Y(n397) );
  MUX21X2_HVT U189 ( .A1(n536), .A2(n526), .S0(n252), .Y(out[3]) );
  IBUFFX16_HVT U190 ( .A(n307), .Y(n252) );
  INVX1_HVT U193 ( .A(n348), .Y(n287) );
  INVX1_HVT U196 ( .A(n446), .Y(n415) );
  MUX41X1_HVT U197 ( .A1(n484), .A3(n486), .A2(n478), .A4(n482), .S0(n253), 
        .S1(n254), .Y(n477) );
  IBUFFX16_HVT U199 ( .A(n293), .Y(n253) );
  IBUFFX16_HVT U201 ( .A(n349), .Y(n254) );
  INVX1_HVT U202 ( .A(n449), .Y(n412) );
  INVX2_HVT U203 ( .A(n430), .Y(n309) );
  INVX1_HVT U204 ( .A(in[3]), .Y(n430) );
  INVX1_HVT U205 ( .A(n354), .Y(n432) );
  MUX21X1_HVT U206 ( .A1(n353), .A2(n360), .S0(n298), .Y(n255) );
  IBUFFX16_HVT U208 ( .A(n255), .Y(n599) );
  MUX41X1_HVT U209 ( .A1(n497), .A3(n316), .A2(n405), .A4(n417), .S0(n256), 
        .S1(n257), .Y(n496) );
  IBUFFX16_HVT U210 ( .A(n330), .Y(n257) );
  IBUFFX2_HVT U211 ( .A(n371), .Y(n296) );
  MUX21X1_HVT U212 ( .A1(n259), .A2(n260), .S0(n362), .Y(n258) );
  MUX21X1_HVT U213 ( .A1(n509), .A2(n510), .S0(n346), .Y(n508) );
  MUX21X2_HVT U214 ( .A1(n494), .A2(n495), .S0(n336), .Y(n493) );
  MUX21X2_HVT U215 ( .A1(n584), .A2(n585), .S0(n262), .Y(n582) );
  IBUFFX16_HVT U216 ( .A(n335), .Y(n262) );
  NAND2X0_HVT U217 ( .A1(n543), .A2(n263), .Y(n264) );
  NAND2X0_HVT U218 ( .A1(n550), .A2(n307), .Y(n265) );
  NAND2X0_HVT U219 ( .A1(n264), .A2(n265), .Y(out[2]) );
  IBUFFX2_HVT U220 ( .A(n307), .Y(n263) );
  INVX0_HVT U221 ( .A(n635), .Y(n266) );
  INVX1_HVT U222 ( .A(n266), .Y(n267) );
  MUX41X1_HVT U223 ( .A1(n469), .A3(n324), .A2(n599), .A4(n314), .S0(n268), 
        .S1(n283), .Y(n468) );
  IBUFFX16_HVT U224 ( .A(n335), .Y(n268) );
  IBUFFX2_HVT U225 ( .A(n366), .Y(n365) );
  INVX0_HVT U226 ( .A(n640), .Y(n378) );
  MUX21X2_HVT U227 ( .A1(n306), .A2(n589), .S0(n338), .Y(n585) );
  MUX21X2_HVT U228 ( .A1(n534), .A2(n535), .S0(n336), .Y(n533) );
  MUX21X1_HVT U229 ( .A1(n627), .A2(n375), .S0(n271), .Y(n270) );
  MUX21X1_HVT U230 ( .A1(n269), .A2(n270), .S0(n296), .Y(n530) );
  IBUFFX2_HVT U231 ( .A(n332), .Y(n271) );
  NAND2X0_HVT U232 ( .A1(n379), .A2(n272), .Y(n273) );
  NAND2X0_HVT U233 ( .A1(n426), .A2(n299), .Y(n274) );
  NAND2X0_HVT U234 ( .A1(n273), .A2(n274), .Y(n500) );
  MUX21X2_HVT U235 ( .A1(n500), .A2(n499), .S0(n275), .Y(n498) );
  IBUFFX16_HVT U236 ( .A(n305), .Y(n275) );
  INVX1_HVT U237 ( .A(n436), .Y(n426) );
  INVX1_HVT U238 ( .A(n297), .Y(n276) );
  INVX1_HVT U239 ( .A(n276), .Y(n277) );
  NAND2X0_HVT U240 ( .A1(n355), .A2(n279), .Y(n280) );
  NAND2X0_HVT U241 ( .A1(n554), .A2(n282), .Y(n281) );
  NAND2X0_HVT U242 ( .A1(n280), .A2(n281), .Y(n553) );
  INVX0_HVT U243 ( .A(n282), .Y(n279) );
  MUX21X2_HVT U244 ( .A1(n552), .A2(n553), .S0(n331), .Y(n551) );
  INVX0_HVT U245 ( .A(n371), .Y(n370) );
  NBUFFX2_HVT U246 ( .A(n368), .Y(n286) );
  INVX1_HVT U247 ( .A(n371), .Y(n283) );
  INVX1_HVT U248 ( .A(in[4]), .Y(n372) );
  MUX21X2_HVT U249 ( .A1(n566), .A2(n559), .S0(n284), .Y(out[1]) );
  IBUFFX16_HVT U250 ( .A(n307), .Y(n284) );
  MUX41X1_HVT U251 ( .A1(n615), .A3(n405), .A2(n421), .A4(n548), .S0(n285), 
        .S1(n299), .Y(n547) );
  IBUFFX16_HVT U252 ( .A(n334), .Y(n285) );
  MUX41X1_HVT U253 ( .A1(n541), .A3(n538), .A2(n539), .A4(n537), .S0(n288), 
        .S1(n289), .Y(n536) );
  IBUFFX16_HVT U254 ( .A(n349), .Y(n288) );
  IBUFFX16_HVT U255 ( .A(n347), .Y(n289) );
  INVX1_HVT U256 ( .A(n345), .Y(n290) );
  INVX0_HVT U257 ( .A(n618), .Y(n396) );
  INVX1_HVT U258 ( .A(in[5]), .Y(n348) );
  INVX1_HVT U259 ( .A(n348), .Y(n349) );
  INVX1_HVT U260 ( .A(n346), .Y(n304) );
  INVX1_HVT U261 ( .A(n347), .Y(n293) );
  INVX1_HVT U262 ( .A(n333), .Y(n305) );
  MUX41X1_HVT U263 ( .A1(n549), .A3(n546), .A2(n547), .A4(n544), .S0(n348), 
        .S1(n290), .Y(n543) );
  NAND2X0_HVT U264 ( .A1(n470), .A2(n308), .Y(n291) );
  NAND2X0_HVT U265 ( .A1(n477), .A2(n307), .Y(n292) );
  NAND2X0_HVT U266 ( .A1(n291), .A2(n292), .Y(out[6]) );
  MUX41X1_HVT U267 ( .A1(n589), .A3(n419), .A2(n433), .A4(n427), .S0(n305), 
        .S1(n368), .Y(n471) );
  NAND2X0_HVT U268 ( .A1(n466), .A2(n293), .Y(n294) );
  NAND2X0_HVT U269 ( .A1(n468), .A2(n347), .Y(n295) );
  NAND2X0_HVT U270 ( .A1(n294), .A2(n295), .Y(n465) );
  MUX41X1_HVT U271 ( .A1(n556), .A3(n596), .A2(n636), .A4(n311), .S0(n305), 
        .S1(n372), .Y(n555) );
  NAND2X0_HVT U272 ( .A1(n491), .A2(n308), .Y(n301) );
  NAND2X0_HVT U273 ( .A1(n300), .A2(n301), .Y(out[5]) );
  NAND2X0_HVT U274 ( .A1(n414), .A2(n299), .Y(n302) );
  NAND2X0_HVT U275 ( .A1(n602), .A2(n338), .Y(n303) );
  NAND2X0_HVT U276 ( .A1(n302), .A2(n303), .Y(n458) );
  INVX1_HVT U277 ( .A(n614), .Y(n400) );
  INVX1_HVT U278 ( .A(n447), .Y(n414) );
  MUX41X1_HVT U279 ( .A1(n639), .A3(n634), .A2(n412), .A4(n416), .S0(n305), 
        .S1(n372), .Y(n564) );
  MUX21X1_HVT U280 ( .A1(n428), .A2(n222), .S0(n226), .Y(n617) );
  INVX1_HVT U281 ( .A(n306), .Y(n620) );
  MUX41X1_HVT U282 ( .A1(n493), .A3(n498), .A2(n492), .A4(n496), .S0(in[5]), 
        .S1(n293), .Y(n491) );
  MUX21X1_HVT U283 ( .A1(n642), .A2(n340), .S0(n297), .Y(n306) );
  INVX0_HVT U284 ( .A(n642), .Y(n428) );
  INVX1_HVT U285 ( .A(in[0]), .Y(n366) );
  NBUFFX2_HVT U286 ( .A(in[7]), .Y(n307) );
  MUX41X1_HVT U287 ( .A1(n384), .A3(n631), .A2(n431), .A4(n315), .S0(n305), 
        .S1(n372), .Y(n573) );
  INVX0_HVT U288 ( .A(in[7]), .Y(n308) );
  INVX1_HVT U289 ( .A(n318), .Y(n474) );
  INVX0_HVT U290 ( .A(n310), .Y(n607) );
  INVX0_HVT U291 ( .A(n317), .Y(n476) );
  INVX1_HVT U292 ( .A(n360), .Y(n431) );
  MUX41X1_HVT U293 ( .A1(n625), .A3(n402), .A2(n624), .A4(n400), .S0(n305), 
        .S1(n372), .Y(n565) );
  INVX1_HVT U294 ( .A(n344), .Y(n346) );
  NBUFFX2_HVT U295 ( .A(n430), .Y(n340) );
  MUX21X1_HVT U296 ( .A1(n351), .A2(n319), .S0(n226), .Y(n310) );
  INVX1_HVT U297 ( .A(n311), .Y(n312) );
  INVX1_HVT U298 ( .A(n311), .Y(n313) );
  INVX1_HVT U299 ( .A(n360), .Y(n314) );
  INVX1_HVT U300 ( .A(n380), .Y(n315) );
  MUX21X1_HVT U301 ( .A1(n356), .A2(n312), .S0(n282), .Y(n317) );
  MUX21X1_HVT U302 ( .A1(n312), .A2(n319), .S0(n362), .Y(n318) );
  MUX41X1_HVT U303 ( .A1(n475), .A3(n473), .A2(n472), .A4(n471), .S0(n344), 
        .S1(n348), .Y(n470) );
  INVX0_HVT U304 ( .A(in[1]), .Y(n344) );
  INVX1_HVT U305 ( .A(n352), .Y(n429) );
  NBUFFX2_HVT U306 ( .A(n642), .Y(n357) );
  NBUFFX2_HVT U307 ( .A(n638), .Y(n352) );
  NBUFFX2_HVT U308 ( .A(n357), .Y(n359) );
  NBUFFX2_HVT U309 ( .A(n642), .Y(n358) );
  NBUFFX2_HVT U310 ( .A(n638), .Y(n353) );
  AND2X1_HVT U311 ( .A1(n637), .A2(n358), .Y(n320) );
  AND2X1_HVT U312 ( .A1(n358), .A2(n627), .Y(n321) );
  NAND2X0_HVT U313 ( .A1(n340), .A2(n342), .Y(n642) );
  MUX21X1_HVT U314 ( .A1(n428), .A2(n433), .S0(n361), .Y(n610) );
  MUX21X1_HVT U315 ( .A1(n222), .A2(n429), .S0(n365), .Y(n497) );
  MUX41X1_HVT U316 ( .A1(n324), .A3(n320), .A2(n323), .A4(n476), .S0(n335), 
        .S1(n286), .Y(n475) );
  MUX21X1_HVT U317 ( .A1(n314), .A2(n429), .S0(n361), .Y(n615) );
  MUX21X1_HVT U318 ( .A1(n341), .A2(n428), .S0(n278), .Y(n613) );
  MUX21X1_HVT U319 ( .A1(n394), .A2(n580), .S0(n326), .Y(n579) );
  MUX21X1_HVT U320 ( .A1(n431), .A2(n351), .S0(n227), .Y(n442) );
  MUX21X1_HVT U321 ( .A1(n610), .A2(n321), .S0(n336), .Y(n518) );
  MUX21X1_HVT U322 ( .A1(n341), .A2(n433), .S0(n361), .Y(n444) );
  MUX21X1_HVT U323 ( .A1(n352), .A2(n355), .S0(n277), .Y(n485) );
  MUX21X1_HVT U324 ( .A1(n425), .A2(n322), .S0(n331), .Y(n521) );
  INVX1_HVT U325 ( .A(n626), .Y(n433) );
  MUX21X1_HVT U326 ( .A1(n350), .A2(n341), .S0(n365), .Y(n621) );
  MUX21X1_HVT U327 ( .A1(n433), .A2(n340), .S0(n361), .Y(n604) );
  MUX21X1_HVT U328 ( .A1(n350), .A2(n431), .S0(n227), .Y(n612) );
  MUX21X1_HVT U329 ( .A1(n428), .A2(n432), .S0(n277), .Y(n593) );
  MUX21X1_HVT U330 ( .A1(n357), .A2(n353), .S0(n278), .Y(n503) );
  XOR2X1_HVT U331 ( .A1(n356), .A2(n278), .Y(n596) );
  XNOR2X1_HVT U332 ( .A1(n357), .A2(n365), .Y(n322) );
  MUX21X1_HVT U333 ( .A1(n432), .A2(n340), .S0(n297), .Y(n446) );
  MUX21X1_HVT U334 ( .A1(n351), .A2(n429), .S0(n364), .Y(n609) );
  MUX21X1_HVT U335 ( .A1(n433), .A2(n222), .S0(n278), .Y(n437) );
  MUX21X1_HVT U336 ( .A1(n352), .A2(n359), .S0(n362), .Y(n436) );
  MUX21X1_HVT U337 ( .A1(n384), .A2(n350), .S0(n339), .Y(n552) );
  MUX21X1_HVT U338 ( .A1(n350), .A2(n222), .S0(n338), .Y(n554) );
  MUX21X1_HVT U339 ( .A1(n340), .A2(n358), .S0(n277), .Y(n445) );
  MUX21X1_HVT U340 ( .A1(n355), .A2(n358), .S0(n365), .Y(n624) );
  MUX21X1_HVT U341 ( .A1(n313), .A2(n359), .S0(n364), .Y(n628) );
  MUX21X1_HVT U342 ( .A1(n342), .A2(n359), .S0(n364), .Y(n540) );
  XOR2X1_HVT U343 ( .A1(n351), .A2(n297), .Y(n597) );
  MUX21X1_HVT U344 ( .A1(n356), .A2(n340), .S0(n227), .Y(n623) );
  MUX21X1_HVT U345 ( .A1(n395), .A2(n587), .S0(n326), .Y(n586) );
  MUX21X1_HVT U346 ( .A1(n396), .A2(n639), .S0(n336), .Y(n587) );
  XOR2X1_HVT U347 ( .A1(n313), .A2(n362), .Y(n606) );
  MUX21X1_HVT U348 ( .A1(n222), .A2(n351), .S0(n278), .Y(n603) );
  MUX21X1_HVT U349 ( .A1(n341), .A2(n356), .S0(n364), .Y(n439) );
  NBUFFX2_HVT U350 ( .A(n370), .Y(n338) );
  NBUFFX2_HVT U351 ( .A(n370), .Y(n337) );
  NBUFFX2_HVT U352 ( .A(n370), .Y(n339) );
  AND2X1_HVT U353 ( .A1(n361), .A2(n342), .Y(n323) );
  MUX21X1_HVT U354 ( .A1(n461), .A2(n416), .S0(n337), .Y(n460) );
  NBUFFX2_HVT U355 ( .A(n643), .Y(n360) );
  MUX21X1_HVT U356 ( .A1(n409), .A2(n323), .S0(n337), .Y(n452) );
  NBUFFX2_HVT U357 ( .A(n626), .Y(n350) );
  AND2X1_HVT U358 ( .A1(n432), .A2(n247), .Y(n324) );
  MUX21X1_HVT U359 ( .A1(n398), .A2(n389), .S0(n339), .Y(n592) );
  NBUFFX2_HVT U360 ( .A(n641), .Y(n354) );
  NBUFFX2_HVT U361 ( .A(n626), .Y(n351) );
  AND2X1_HVT U362 ( .A1(n356), .A2(n247), .Y(n325) );
  MUX21X1_HVT U363 ( .A1(n415), .A2(n374), .S0(n339), .Y(n569) );
  NBUFFX2_HVT U364 ( .A(n641), .Y(n356) );
  NBUFFX2_HVT U365 ( .A(n641), .Y(n355) );
  NBUFFX2_HVT U366 ( .A(n367), .Y(n335) );
  NBUFFX2_HVT U367 ( .A(n367), .Y(n336) );
  XNOR2X1_HVT U368 ( .A1(n371), .A2(n332), .Y(n326) );
  NBUFFX2_HVT U369 ( .A(n333), .Y(n334) );
  NBUFFX2_HVT U370 ( .A(n367), .Y(n332) );
  NBUFFX2_HVT U371 ( .A(in[2]), .Y(n333) );
  NBUFFX2_HVT U372 ( .A(n367), .Y(n331) );
  NBUFFX2_HVT U373 ( .A(n367), .Y(n330) );
  INVX1_HVT U374 ( .A(n344), .Y(n347) );
  INVX1_HVT U375 ( .A(n344), .Y(n345) );
  NAND2X0_HVT U376 ( .A1(n309), .A2(n342), .Y(n643) );
  MUX21X1_HVT U377 ( .A1(n353), .A2(n309), .S0(n365), .Y(n548) );
  MUX21X1_HVT U378 ( .A1(n431), .A2(n309), .S0(n362), .Y(n435) );
  MUX21X1_HVT U379 ( .A1(n432), .A2(n429), .S0(n227), .Y(n529) );
  MUX21X1_HVT U380 ( .A1(n309), .A2(n353), .S0(n363), .Y(n440) );
  MUX21X1_HVT U381 ( .A1(n312), .A2(n309), .S0(n362), .Y(n488) );
  MUX21X1_HVT U382 ( .A1(n309), .A2(n313), .S0(n363), .Y(n441) );
  MUX21X1_HVT U383 ( .A1(n222), .A2(n309), .S0(n363), .Y(n616) );
  NBUFFX2_HVT U384 ( .A(in[2]), .Y(n367) );
  MUX21X1_HVT U385 ( .A1(n341), .A2(n222), .S0(n297), .Y(n598) );
  MUX21X1_HVT U386 ( .A1(n428), .A2(n342), .S0(n363), .Y(n447) );
  NAND2X0_HVT U387 ( .A1(n463), .A2(n293), .Y(n328) );
  NAND2X0_HVT U388 ( .A1(n464), .A2(n346), .Y(n329) );
  NAND2X0_HVT U389 ( .A1(n328), .A2(n329), .Y(n462) );
  MUX21X1_HVT U390 ( .A1(n428), .A2(n327), .S0(n364), .Y(n511) );
  XOR2X1_HVT U391 ( .A1(n363), .A2(n327), .Y(n594) );
  MUX21X1_HVT U392 ( .A1(n327), .A2(n314), .S0(n364), .Y(n619) );
  MUX21X1_HVT U393 ( .A1(n355), .A2(n327), .S0(n363), .Y(n443) );
  MUX21X1_HVT U394 ( .A1(n327), .A2(n355), .S0(n365), .Y(n448) );
  MUX21X1_HVT U395 ( .A1(n340), .A2(n327), .S0(n227), .Y(n438) );
  MUX21X1_HVT U396 ( .A1(n327), .A2(n312), .S0(n362), .Y(n625) );
  MUX21X1_HVT U397 ( .A1(n327), .A2(n429), .S0(n361), .Y(n449) );
  MUX21X1_HVT U398 ( .A1(n327), .A2(n432), .S0(n297), .Y(n602) );
  INVX0_HVT U399 ( .A(n631), .Y(n373) );
  INVX0_HVT U400 ( .A(n611), .Y(n374) );
  INVX0_HVT U401 ( .A(n605), .Y(n375) );
  INVX0_HVT U402 ( .A(n545), .Y(n376) );
  INVX0_HVT U403 ( .A(n506), .Y(n377) );
  INVX0_HVT U404 ( .A(n639), .Y(n379) );
  INVX0_HVT U405 ( .A(n637), .Y(n380) );
  INVX0_HVT U406 ( .A(n601), .Y(n381) );
  INVX0_HVT U407 ( .A(n636), .Y(n382) );
  INVX0_HVT U408 ( .A(n267), .Y(n383) );
  INVX0_HVT U409 ( .A(n608), .Y(n384) );
  INVX0_HVT U410 ( .A(n629), .Y(n385) );
  INVX0_HVT U411 ( .A(n634), .Y(n386) );
  INVX0_HVT U412 ( .A(n630), .Y(n387) );
  INVX0_HVT U413 ( .A(n628), .Y(n388) );
  INVX0_HVT U414 ( .A(n627), .Y(n389) );
  INVX0_HVT U415 ( .A(n625), .Y(n390) );
  INVX0_HVT U416 ( .A(n624), .Y(n391) );
  INVX0_HVT U417 ( .A(n623), .Y(n392) );
  INVX0_HVT U418 ( .A(n622), .Y(n393) );
  INVX0_HVT U419 ( .A(n619), .Y(n395) );
  INVX0_HVT U420 ( .A(n616), .Y(n398) );
  INVX0_HVT U421 ( .A(n615), .Y(n399) );
  INVX0_HVT U422 ( .A(n613), .Y(n401) );
  INVX0_HVT U423 ( .A(n612), .Y(n402) );
  INVX0_HVT U424 ( .A(n610), .Y(n403) );
  INVX0_HVT U425 ( .A(n609), .Y(n404) );
  INVX0_HVT U426 ( .A(n606), .Y(n405) );
  INVX0_HVT U427 ( .A(n604), .Y(n406) );
  INVX0_HVT U428 ( .A(n603), .Y(n407) );
  INVX0_HVT U429 ( .A(n598), .Y(n409) );
  INVX0_HVT U430 ( .A(n597), .Y(n410) );
  INVX0_HVT U431 ( .A(n633), .Y(n411) );
  INVX0_HVT U432 ( .A(n448), .Y(n413) );
  INVX0_HVT U433 ( .A(n445), .Y(n416) );
  INVX0_HVT U434 ( .A(n443), .Y(n418) );
  INVX0_HVT U435 ( .A(n442), .Y(n419) );
  INVX0_HVT U436 ( .A(n441), .Y(n420) );
  INVX0_HVT U437 ( .A(n440), .Y(n421) );
  INVX0_HVT U438 ( .A(n439), .Y(n422) );
  INVX0_HVT U439 ( .A(n438), .Y(n423) );
  INVX0_HVT U440 ( .A(n488), .Y(n424) );
  INVX0_HVT U441 ( .A(n437), .Y(n425) );
  INVX0_HVT U442 ( .A(n435), .Y(n427) );
endmodule

