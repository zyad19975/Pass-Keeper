
module cde ( clk, rst, cam_start, pass, start_dec, start_enc, master_key, 
        account, data_flash, flash_pass_reg, flash_acc_reg, flash_or_acc_reg, 
        flash_or_acc_sel, pass_enc_reg, new_old_pass_sel, plain_reg, 
        local_master_reg, local_master_sel, out_reg, write_en, write_add, 
        boot_lood, match, dec_done, ready_encryption, write_data_flash, 
        add_flash, final_output );
  input [127:0] pass;
  input [127:0] master_key;
  input [127:0] account;
  input [255:0] data_flash;
  input [3:0] write_add;
  output [255:0] write_data_flash;
  output [3:0] add_flash;
  output [127:0] final_output;
  input clk, rst, cam_start, start_dec, start_enc, flash_pass_reg,
         flash_acc_reg, flash_or_acc_reg, flash_or_acc_sel, pass_enc_reg,
         new_old_pass_sel, plain_reg, local_master_reg, local_master_sel,
         out_reg, write_en, boot_lood;
  output match, dec_done, ready_encryption;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306;
  wire   [127:0] out_flash_or_acc_sel;
  wire   [3:0] match_add;
  wire   [127:0] out_new_old_pass_sel;
  wire   [127:0] out_decry;
  wire   [127:0] out_local_master_sel;
  wire   [127:0] out_reg_flash_or_acc;
  wire   [127:0] out_encryption;
  wire   [127:0] out_reg_pass_enc;
  wire   [127:0] out_reg_plain_reg;
  wire   [127:0] out_local_master_reg;

  AO22X1_HVT U6 ( .A1(out_decry[99]), .A2(n267), .A3(pass[99]), .A4(n73), .Y(
        out_new_old_pass_sel[99]) );
  AO22X1_HVT U7 ( .A1(out_decry[98]), .A2(n137), .A3(pass[98]), .A4(n73), .Y(
        out_new_old_pass_sel[98]) );
  AO22X1_HVT U8 ( .A1(out_decry[97]), .A2(n268), .A3(pass[97]), .A4(n280), .Y(
        out_new_old_pass_sel[97]) );
  AO22X1_HVT U9 ( .A1(out_decry[96]), .A2(n268), .A3(pass[96]), .A4(n19), .Y(
        out_new_old_pass_sel[96]) );
  AO22X1_HVT U10 ( .A1(out_decry[95]), .A2(n210), .A3(pass[95]), .A4(n278), 
        .Y(out_new_old_pass_sel[95]) );
  AO22X1_HVT U11 ( .A1(out_decry[94]), .A2(n267), .A3(pass[94]), .A4(n280), 
        .Y(out_new_old_pass_sel[94]) );
  AO22X1_HVT U12 ( .A1(out_decry[93]), .A2(n269), .A3(pass[93]), .A4(n278), 
        .Y(out_new_old_pass_sel[93]) );
  AO22X1_HVT U13 ( .A1(out_decry[92]), .A2(n269), .A3(pass[92]), .A4(n73), .Y(
        out_new_old_pass_sel[92]) );
  AO22X1_HVT U14 ( .A1(out_decry[91]), .A2(n237), .A3(pass[91]), .A4(n11), .Y(
        out_new_old_pass_sel[91]) );
  AO22X1_HVT U15 ( .A1(out_decry[90]), .A2(n268), .A3(pass[90]), .A4(n19), .Y(
        out_new_old_pass_sel[90]) );
  AO22X1_HVT U17 ( .A1(out_decry[89]), .A2(n269), .A3(pass[89]), .A4(n42), .Y(
        out_new_old_pass_sel[89]) );
  AO22X1_HVT U18 ( .A1(out_decry[88]), .A2(n210), .A3(pass[88]), .A4(n42), .Y(
        out_new_old_pass_sel[88]) );
  AO22X1_HVT U19 ( .A1(out_decry[87]), .A2(n63), .A3(pass[87]), .A4(n192), .Y(
        out_new_old_pass_sel[87]) );
  AO22X1_HVT U20 ( .A1(out_decry[86]), .A2(n236), .A3(pass[86]), .A4(n42), .Y(
        out_new_old_pass_sel[86]) );
  AO22X1_HVT U21 ( .A1(out_decry[85]), .A2(n236), .A3(pass[85]), .A4(n192), 
        .Y(out_new_old_pass_sel[85]) );
  AO22X1_HVT U22 ( .A1(out_decry[84]), .A2(n237), .A3(pass[84]), .A4(n192), 
        .Y(out_new_old_pass_sel[84]) );
  AO22X1_HVT U23 ( .A1(out_decry[83]), .A2(n267), .A3(pass[83]), .A4(n27), .Y(
        out_new_old_pass_sel[83]) );
  AO22X1_HVT U24 ( .A1(out_decry[82]), .A2(n9), .A3(pass[82]), .A4(n27), .Y(
        out_new_old_pass_sel[82]) );
  AO22X1_HVT U25 ( .A1(out_decry[81]), .A2(n138), .A3(pass[81]), .A4(n27), .Y(
        out_new_old_pass_sel[81]) );
  AO22X1_HVT U26 ( .A1(out_decry[80]), .A2(n137), .A3(pass[80]), .A4(n277), 
        .Y(out_new_old_pass_sel[80]) );
  AO22X1_HVT U28 ( .A1(out_decry[79]), .A2(n9), .A3(pass[79]), .A4(n282), .Y(
        out_new_old_pass_sel[79]) );
  AO22X1_HVT U29 ( .A1(out_decry[78]), .A2(n17), .A3(pass[78]), .A4(n66), .Y(
        out_new_old_pass_sel[78]) );
  AO22X1_HVT U30 ( .A1(out_decry[77]), .A2(n266), .A3(pass[77]), .A4(n276), 
        .Y(out_new_old_pass_sel[77]) );
  AO22X1_HVT U31 ( .A1(out_decry[76]), .A2(n138), .A3(pass[76]), .A4(n27), .Y(
        out_new_old_pass_sel[76]) );
  AO22X1_HVT U32 ( .A1(out_decry[75]), .A2(n17), .A3(pass[75]), .A4(n56), .Y(
        out_new_old_pass_sel[75]) );
  AO22X1_HVT U33 ( .A1(out_decry[74]), .A2(n266), .A3(pass[74]), .A4(n276), 
        .Y(out_new_old_pass_sel[74]) );
  AO22X1_HVT U34 ( .A1(out_decry[73]), .A2(n137), .A3(pass[73]), .A4(n281), 
        .Y(out_new_old_pass_sel[73]) );
  AO22X1_HVT U35 ( .A1(out_decry[72]), .A2(n266), .A3(pass[72]), .A4(n66), .Y(
        out_new_old_pass_sel[72]) );
  AO22X1_HVT U36 ( .A1(out_decry[71]), .A2(n9), .A3(pass[71]), .A4(n73), .Y(
        out_new_old_pass_sel[71]) );
  AO22X1_HVT U37 ( .A1(out_decry[70]), .A2(n138), .A3(pass[70]), .A4(n282), 
        .Y(out_new_old_pass_sel[70]) );
  AO22X1_HVT U39 ( .A1(out_decry[69]), .A2(n9), .A3(pass[69]), .A4(n280), .Y(
        out_new_old_pass_sel[69]) );
  AO22X1_HVT U40 ( .A1(out_decry[68]), .A2(n138), .A3(pass[68]), .A4(n11), .Y(
        out_new_old_pass_sel[68]) );
  AO22X1_HVT U41 ( .A1(out_decry[67]), .A2(n191), .A3(pass[67]), .A4(n11), .Y(
        out_new_old_pass_sel[67]) );
  AO22X1_HVT U42 ( .A1(out_decry[66]), .A2(n17), .A3(pass[66]), .A4(n281), .Y(
        out_new_old_pass_sel[66]) );
  AO22X1_HVT U43 ( .A1(out_decry[65]), .A2(n137), .A3(pass[65]), .A4(n276), 
        .Y(out_new_old_pass_sel[65]) );
  AO22X1_HVT U44 ( .A1(out_decry[64]), .A2(n237), .A3(pass[64]), .A4(n280), 
        .Y(out_new_old_pass_sel[64]) );
  AO22X1_HVT U45 ( .A1(out_decry[63]), .A2(n267), .A3(pass[63]), .A4(n280), 
        .Y(out_new_old_pass_sel[63]) );
  AO22X1_HVT U46 ( .A1(out_decry[62]), .A2(n210), .A3(pass[62]), .A4(n11), .Y(
        out_new_old_pass_sel[62]) );
  AO22X1_HVT U47 ( .A1(out_decry[61]), .A2(n210), .A3(pass[61]), .A4(n42), .Y(
        out_new_old_pass_sel[61]) );
  AO22X1_HVT U48 ( .A1(out_decry[60]), .A2(n237), .A3(pass[60]), .A4(n277), 
        .Y(out_new_old_pass_sel[60]) );
  AO22X1_HVT U49 ( .A1(out_decry[5]), .A2(n236), .A3(pass[5]), .A4(n280), .Y(
        out_new_old_pass_sel[5]) );
  AO22X1_HVT U50 ( .A1(out_decry[59]), .A2(n236), .A3(pass[59]), .A4(n275), 
        .Y(out_new_old_pass_sel[59]) );
  AO22X1_HVT U51 ( .A1(out_decry[58]), .A2(n269), .A3(pass[58]), .A4(n279), 
        .Y(out_new_old_pass_sel[58]) );
  AO22X1_HVT U52 ( .A1(out_decry[57]), .A2(n63), .A3(pass[57]), .A4(n11), .Y(
        out_new_old_pass_sel[57]) );
  AO22X1_HVT U53 ( .A1(out_decry[56]), .A2(n236), .A3(pass[56]), .A4(n42), .Y(
        out_new_old_pass_sel[56]) );
  AO22X1_HVT U54 ( .A1(out_decry[55]), .A2(n237), .A3(pass[55]), .A4(n11), .Y(
        out_new_old_pass_sel[55]) );
  AO22X1_HVT U55 ( .A1(out_decry[54]), .A2(n268), .A3(pass[54]), .A4(n282), 
        .Y(out_new_old_pass_sel[54]) );
  AO22X1_HVT U56 ( .A1(out_decry[53]), .A2(n137), .A3(pass[53]), .A4(n276), 
        .Y(out_new_old_pass_sel[53]) );
  AO22X1_HVT U57 ( .A1(out_decry[52]), .A2(n268), .A3(pass[52]), .A4(n27), .Y(
        out_new_old_pass_sel[52]) );
  AO22X1_HVT U59 ( .A1(out_decry[50]), .A2(n269), .A3(pass[50]), .A4(n77), .Y(
        out_new_old_pass_sel[50]) );
  AO22X1_HVT U61 ( .A1(out_decry[49]), .A2(n237), .A3(pass[49]), .A4(n27), .Y(
        out_new_old_pass_sel[49]) );
  AO22X1_HVT U62 ( .A1(out_decry[48]), .A2(n236), .A3(pass[48]), .A4(n281), 
        .Y(out_new_old_pass_sel[48]) );
  AO22X1_HVT U68 ( .A1(out_decry[42]), .A2(n273), .A3(pass[42]), .A4(n56), .Y(
        out_new_old_pass_sel[42]) );
  AO22X1_HVT U69 ( .A1(out_decry[41]), .A2(n239), .A3(pass[41]), .A4(n56), .Y(
        out_new_old_pass_sel[41]) );
  AO22X1_HVT U70 ( .A1(out_decry[40]), .A2(n272), .A3(pass[40]), .A4(n281), 
        .Y(out_new_old_pass_sel[40]) );
  AO22X1_HVT U72 ( .A1(out_decry[39]), .A2(n270), .A3(pass[39]), .A4(n56), .Y(
        out_new_old_pass_sel[39]) );
  AO22X1_HVT U73 ( .A1(out_decry[38]), .A2(n271), .A3(pass[38]), .A4(n42), .Y(
        out_new_old_pass_sel[38]) );
  AO22X1_HVT U74 ( .A1(out_decry[37]), .A2(n271), .A3(pass[37]), .A4(n277), 
        .Y(out_new_old_pass_sel[37]) );
  AO22X1_HVT U75 ( .A1(out_decry[36]), .A2(n238), .A3(pass[36]), .A4(n281), 
        .Y(out_new_old_pass_sel[36]) );
  AO22X1_HVT U76 ( .A1(out_decry[35]), .A2(n148), .A3(pass[35]), .A4(n56), .Y(
        out_new_old_pass_sel[35]) );
  AO22X1_HVT U77 ( .A1(out_decry[34]), .A2(n10), .A3(pass[34]), .A4(n209), .Y(
        out_new_old_pass_sel[34]) );
  AO22X1_HVT U78 ( .A1(out_decry[33]), .A2(n272), .A3(pass[33]), .A4(n18), .Y(
        out_new_old_pass_sel[33]) );
  AO22X1_HVT U79 ( .A1(out_decry[32]), .A2(n10), .A3(pass[32]), .A4(n209), .Y(
        out_new_old_pass_sel[32]) );
  AO22X1_HVT U80 ( .A1(out_decry[31]), .A2(n147), .A3(pass[31]), .A4(n209), 
        .Y(out_new_old_pass_sel[31]) );
  AO22X1_HVT U81 ( .A1(out_decry[30]), .A2(n273), .A3(pass[30]), .A4(n209), 
        .Y(out_new_old_pass_sel[30]) );
  AO22X1_HVT U82 ( .A1(out_decry[2]), .A2(n148), .A3(pass[2]), .A4(n209), .Y(
        out_new_old_pass_sel[2]) );
  AO22X1_HVT U83 ( .A1(out_decry[29]), .A2(n270), .A3(pass[29]), .A4(n68), .Y(
        out_new_old_pass_sel[29]) );
  AO22X1_HVT U84 ( .A1(out_decry[28]), .A2(n239), .A3(pass[28]), .A4(n68), .Y(
        out_new_old_pass_sel[28]) );
  AO22X1_HVT U85 ( .A1(out_decry[27]), .A2(n147), .A3(pass[27]), .A4(n68), .Y(
        out_new_old_pass_sel[27]) );
  AO22X1_HVT U86 ( .A1(out_decry[26]), .A2(n273), .A3(pass[26]), .A4(n68), .Y(
        out_new_old_pass_sel[26]) );
  AO22X1_HVT U87 ( .A1(out_decry[25]), .A2(n239), .A3(pass[25]), .A4(n281), 
        .Y(out_new_old_pass_sel[25]) );
  AO22X1_HVT U88 ( .A1(out_decry[24]), .A2(n272), .A3(pass[24]), .A4(n56), .Y(
        out_new_old_pass_sel[24]) );
  AO22X1_HVT U90 ( .A1(out_decry[22]), .A2(n148), .A3(pass[22]), .A4(n66), .Y(
        out_new_old_pass_sel[22]) );
  AO22X1_HVT U91 ( .A1(out_decry[21]), .A2(n148), .A3(pass[21]), .A4(n66), .Y(
        out_new_old_pass_sel[21]) );
  AO22X1_HVT U92 ( .A1(out_decry[20]), .A2(n271), .A3(pass[20]), .A4(n277), 
        .Y(out_new_old_pass_sel[20]) );
  AO22X1_HVT U94 ( .A1(out_decry[19]), .A2(n148), .A3(pass[19]), .A4(n282), 
        .Y(out_new_old_pass_sel[19]) );
  AO22X1_HVT U96 ( .A1(out_decry[17]), .A2(n271), .A3(pass[17]), .A4(n66), .Y(
        out_new_old_pass_sel[17]) );
  AO22X1_HVT U97 ( .A1(out_decry[16]), .A2(n273), .A3(pass[16]), .A4(n278), 
        .Y(out_new_old_pass_sel[16]) );
  AO22X1_HVT U98 ( .A1(out_decry[15]), .A2(n10), .A3(pass[15]), .A4(n11), .Y(
        out_new_old_pass_sel[15]) );
  AO22X1_HVT U99 ( .A1(out_decry[14]), .A2(n239), .A3(pass[14]), .A4(n282), 
        .Y(out_new_old_pass_sel[14]) );
  AO22X1_HVT U100 ( .A1(out_decry[13]), .A2(n271), .A3(pass[13]), .A4(n277), 
        .Y(out_new_old_pass_sel[13]) );
  AO22X1_HVT U101 ( .A1(out_decry[12]), .A2(n271), .A3(pass[12]), .A4(n280), 
        .Y(out_new_old_pass_sel[12]) );
  AO22X1_HVT U102 ( .A1(out_decry[127]), .A2(n239), .A3(pass[127]), .A4(n279), 
        .Y(out_new_old_pass_sel[127]) );
  AO22X1_HVT U103 ( .A1(out_decry[126]), .A2(n270), .A3(pass[126]), .A4(n19), 
        .Y(out_new_old_pass_sel[126]) );
  AO22X1_HVT U104 ( .A1(out_decry[125]), .A2(n239), .A3(pass[125]), .A4(n19), 
        .Y(out_new_old_pass_sel[125]) );
  AO22X1_HVT U105 ( .A1(out_decry[124]), .A2(n238), .A3(pass[124]), .A4(n73), 
        .Y(out_new_old_pass_sel[124]) );
  AO22X1_HVT U106 ( .A1(out_decry[123]), .A2(n270), .A3(pass[123]), .A4(n73), 
        .Y(out_new_old_pass_sel[123]) );
  AO22X1_HVT U107 ( .A1(out_decry[122]), .A2(n271), .A3(pass[122]), .A4(n280), 
        .Y(out_new_old_pass_sel[122]) );
  AO22X1_HVT U108 ( .A1(out_decry[121]), .A2(n238), .A3(pass[121]), .A4(n281), 
        .Y(out_new_old_pass_sel[121]) );
  AO22X1_HVT U109 ( .A1(out_decry[120]), .A2(n238), .A3(pass[120]), .A4(n56), 
        .Y(out_new_old_pass_sel[120]) );
  AO22X1_HVT U110 ( .A1(out_decry[11]), .A2(n270), .A3(pass[11]), .A4(n278), 
        .Y(out_new_old_pass_sel[11]) );
  AO22X1_HVT U111 ( .A1(out_decry[119]), .A2(n272), .A3(pass[119]), .A4(n73), 
        .Y(out_new_old_pass_sel[119]) );
  AO22X1_HVT U112 ( .A1(out_decry[118]), .A2(n270), .A3(pass[118]), .A4(n277), 
        .Y(out_new_old_pass_sel[118]) );
  AO22X1_HVT U113 ( .A1(out_decry[117]), .A2(n238), .A3(pass[117]), .A4(n16), 
        .Y(out_new_old_pass_sel[117]) );
  AO22X1_HVT U114 ( .A1(out_decry[116]), .A2(n10), .A3(pass[116]), .A4(n16), 
        .Y(out_new_old_pass_sel[116]) );
  AO22X1_HVT U115 ( .A1(out_decry[115]), .A2(n239), .A3(pass[115]), .A4(n16), 
        .Y(out_new_old_pass_sel[115]) );
  AO22X1_HVT U116 ( .A1(out_decry[114]), .A2(n273), .A3(pass[114]), .A4(n16), 
        .Y(out_new_old_pass_sel[114]) );
  AO22X1_HVT U117 ( .A1(out_decry[113]), .A2(n271), .A3(pass[113]), .A4(n208), 
        .Y(out_new_old_pass_sel[113]) );
  AO22X1_HVT U118 ( .A1(out_decry[112]), .A2(n10), .A3(pass[112]), .A4(n208), 
        .Y(out_new_old_pass_sel[112]) );
  AO22X1_HVT U119 ( .A1(out_decry[111]), .A2(n238), .A3(pass[111]), .A4(n283), 
        .Y(out_new_old_pass_sel[111]) );
  AO22X1_HVT U120 ( .A1(out_decry[110]), .A2(n148), .A3(pass[110]), .A4(n283), 
        .Y(out_new_old_pass_sel[110]) );
  AO22X1_HVT U121 ( .A1(out_decry[10]), .A2(n272), .A3(pass[10]), .A4(n283), 
        .Y(out_new_old_pass_sel[10]) );
  AO22X1_HVT U122 ( .A1(out_decry[109]), .A2(n272), .A3(pass[109]), .A4(n283), 
        .Y(out_new_old_pass_sel[109]) );
  AO22X1_HVT U123 ( .A1(out_decry[108]), .A2(n10), .A3(pass[108]), .A4(n283), 
        .Y(out_new_old_pass_sel[108]) );
  AO22X1_HVT U124 ( .A1(out_decry[107]), .A2(n273), .A3(pass[107]), .A4(n283), 
        .Y(out_new_old_pass_sel[107]) );
  AO22X1_HVT U125 ( .A1(out_decry[106]), .A2(n273), .A3(pass[106]), .A4(n284), 
        .Y(out_new_old_pass_sel[106]) );
  AO22X1_HVT U126 ( .A1(out_decry[105]), .A2(n272), .A3(pass[105]), .A4(n284), 
        .Y(out_new_old_pass_sel[105]) );
  AO22X1_HVT U127 ( .A1(out_decry[104]), .A2(n239), .A3(pass[104]), .A4(n284), 
        .Y(out_new_old_pass_sel[104]) );
  AO22X1_HVT U128 ( .A1(out_decry[103]), .A2(n210), .A3(pass[103]), .A4(n284), 
        .Y(out_new_old_pass_sel[103]) );
  AO22X1_HVT U129 ( .A1(out_decry[102]), .A2(n268), .A3(pass[102]), .A4(n284), 
        .Y(out_new_old_pass_sel[102]) );
  AO22X1_HVT U130 ( .A1(out_decry[101]), .A2(n269), .A3(pass[101]), .A4(n284), 
        .Y(out_new_old_pass_sel[101]) );
  AO22X1_HVT U131 ( .A1(out_decry[100]), .A2(n191), .A3(pass[100]), .A4(n284), 
        .Y(out_new_old_pass_sel[100]) );
  AND2X1_HVT U133 ( .A1(master_key[9]), .A2(n122), .Y(out_local_master_sel[9])
         );
  AND2X1_HVT U134 ( .A1(master_key[99]), .A2(n123), .Y(
        out_local_master_sel[99]) );
  AND2X1_HVT U135 ( .A1(master_key[98]), .A2(n123), .Y(
        out_local_master_sel[98]) );
  AND2X1_HVT U136 ( .A1(master_key[97]), .A2(n122), .Y(
        out_local_master_sel[97]) );
  AND2X1_HVT U137 ( .A1(master_key[96]), .A2(n253), .Y(
        out_local_master_sel[96]) );
  AND2X1_HVT U138 ( .A1(master_key[95]), .A2(n260), .Y(
        out_local_master_sel[95]) );
  AND2X1_HVT U139 ( .A1(master_key[94]), .A2(n260), .Y(
        out_local_master_sel[94]) );
  AND2X1_HVT U140 ( .A1(master_key[93]), .A2(n263), .Y(
        out_local_master_sel[93]) );
  AND2X1_HVT U141 ( .A1(master_key[92]), .A2(n259), .Y(
        out_local_master_sel[92]) );
  AND2X1_HVT U142 ( .A1(master_key[91]), .A2(n262), .Y(
        out_local_master_sel[91]) );
  AND2X1_HVT U143 ( .A1(master_key[90]), .A2(n259), .Y(
        out_local_master_sel[90]) );
  AND2X1_HVT U144 ( .A1(master_key[8]), .A2(n164), .Y(out_local_master_sel[8])
         );
  AND2X1_HVT U145 ( .A1(master_key[89]), .A2(n164), .Y(
        out_local_master_sel[89]) );
  AND2X1_HVT U146 ( .A1(master_key[88]), .A2(n259), .Y(
        out_local_master_sel[88]) );
  AND2X1_HVT U147 ( .A1(master_key[87]), .A2(n164), .Y(
        out_local_master_sel[87]) );
  AND2X1_HVT U148 ( .A1(master_key[86]), .A2(n259), .Y(
        out_local_master_sel[86]) );
  AND2X1_HVT U149 ( .A1(master_key[85]), .A2(n163), .Y(
        out_local_master_sel[85]) );
  AND2X1_HVT U150 ( .A1(master_key[84]), .A2(n164), .Y(
        out_local_master_sel[84]) );
  AND2X1_HVT U151 ( .A1(master_key[83]), .A2(n163), .Y(
        out_local_master_sel[83]) );
  AND2X1_HVT U152 ( .A1(master_key[82]), .A2(n262), .Y(
        out_local_master_sel[82]) );
  AND2X1_HVT U153 ( .A1(master_key[81]), .A2(n161), .Y(
        out_local_master_sel[81]) );
  AND2X1_HVT U154 ( .A1(master_key[80]), .A2(n254), .Y(
        out_local_master_sel[80]) );
  AND2X1_HVT U155 ( .A1(master_key[7]), .A2(n261), .Y(out_local_master_sel[7])
         );
  AND2X1_HVT U156 ( .A1(master_key[79]), .A2(n162), .Y(
        out_local_master_sel[79]) );
  AND2X1_HVT U157 ( .A1(master_key[78]), .A2(n161), .Y(
        out_local_master_sel[78]) );
  AND2X1_HVT U158 ( .A1(master_key[77]), .A2(n254), .Y(
        out_local_master_sel[77]) );
  AND2X1_HVT U159 ( .A1(master_key[76]), .A2(n162), .Y(
        out_local_master_sel[76]) );
  AND2X1_HVT U160 ( .A1(master_key[75]), .A2(n161), .Y(
        out_local_master_sel[75]) );
  AND2X1_HVT U161 ( .A1(master_key[74]), .A2(n254), .Y(
        out_local_master_sel[74]) );
  AND2X1_HVT U162 ( .A1(master_key[73]), .A2(n162), .Y(
        out_local_master_sel[73]) );
  AND2X1_HVT U163 ( .A1(master_key[72]), .A2(n161), .Y(
        out_local_master_sel[72]) );
  AND2X1_HVT U164 ( .A1(master_key[71]), .A2(n254), .Y(
        out_local_master_sel[71]) );
  AND2X1_HVT U165 ( .A1(master_key[70]), .A2(n263), .Y(
        out_local_master_sel[70]) );
  AND2X1_HVT U166 ( .A1(master_key[6]), .A2(n260), .Y(out_local_master_sel[6])
         );
  AND2X1_HVT U167 ( .A1(master_key[69]), .A2(n260), .Y(
        out_local_master_sel[69]) );
  AND2X1_HVT U168 ( .A1(master_key[68]), .A2(n263), .Y(
        out_local_master_sel[68]) );
  AND2X1_HVT U169 ( .A1(master_key[67]), .A2(n122), .Y(
        out_local_master_sel[67]) );
  AND2X1_HVT U170 ( .A1(master_key[66]), .A2(n122), .Y(
        out_local_master_sel[66]) );
  AND2X1_HVT U171 ( .A1(master_key[65]), .A2(n253), .Y(
        out_local_master_sel[65]) );
  AND2X1_HVT U172 ( .A1(master_key[64]), .A2(n123), .Y(
        out_local_master_sel[64]) );
  AND2X1_HVT U173 ( .A1(master_key[63]), .A2(n123), .Y(
        out_local_master_sel[63]) );
  AND2X1_HVT U174 ( .A1(master_key[62]), .A2(n253), .Y(
        out_local_master_sel[62]) );
  AND2X1_HVT U175 ( .A1(master_key[61]), .A2(n263), .Y(
        out_local_master_sel[61]) );
  AND2X1_HVT U176 ( .A1(master_key[60]), .A2(n260), .Y(
        out_local_master_sel[60]) );
  AND2X1_HVT U177 ( .A1(master_key[5]), .A2(n262), .Y(out_local_master_sel[5])
         );
  AND2X1_HVT U178 ( .A1(master_key[59]), .A2(n164), .Y(
        out_local_master_sel[59]) );
  AND2X1_HVT U179 ( .A1(master_key[58]), .A2(n259), .Y(
        out_local_master_sel[58]) );
  AND2X1_HVT U180 ( .A1(master_key[57]), .A2(n262), .Y(
        out_local_master_sel[57]) );
  AND2X1_HVT U181 ( .A1(master_key[56]), .A2(n163), .Y(
        out_local_master_sel[56]) );
  AND2X1_HVT U182 ( .A1(master_key[55]), .A2(n163), .Y(
        out_local_master_sel[55]) );
  AND2X1_HVT U183 ( .A1(master_key[54]), .A2(n262), .Y(
        out_local_master_sel[54]) );
  AND2X1_HVT U184 ( .A1(master_key[53]), .A2(n259), .Y(
        out_local_master_sel[53]) );
  AND2X1_HVT U185 ( .A1(master_key[52]), .A2(n262), .Y(
        out_local_master_sel[52]) );
  AND2X1_HVT U186 ( .A1(master_key[51]), .A2(n163), .Y(
        out_local_master_sel[51]) );
  AND2X1_HVT U187 ( .A1(master_key[50]), .A2(n163), .Y(
        out_local_master_sel[50]) );
  AND2X1_HVT U188 ( .A1(master_key[4]), .A2(n164), .Y(out_local_master_sel[4])
         );
  AND2X1_HVT U189 ( .A1(master_key[49]), .A2(n160), .Y(
        out_local_master_sel[49]) );
  AND2X1_HVT U190 ( .A1(master_key[48]), .A2(n159), .Y(
        out_local_master_sel[48]) );
  AND2X1_HVT U191 ( .A1(master_key[47]), .A2(n258), .Y(
        out_local_master_sel[47]) );
  AND2X1_HVT U192 ( .A1(master_key[46]), .A2(n256), .Y(
        out_local_master_sel[46]) );
  AND2X1_HVT U193 ( .A1(master_key[45]), .A2(n160), .Y(
        out_local_master_sel[45]) );
  AND2X1_HVT U194 ( .A1(master_key[44]), .A2(n159), .Y(
        out_local_master_sel[44]) );
  AND2X1_HVT U195 ( .A1(master_key[43]), .A2(n258), .Y(
        out_local_master_sel[43]) );
  AND2X1_HVT U196 ( .A1(master_key[42]), .A2(n256), .Y(
        out_local_master_sel[42]) );
  AND2X1_HVT U197 ( .A1(master_key[41]), .A2(n160), .Y(
        out_local_master_sel[41]) );
  AND2X1_HVT U198 ( .A1(master_key[40]), .A2(n159), .Y(
        out_local_master_sel[40]) );
  AND2X1_HVT U199 ( .A1(master_key[3]), .A2(n258), .Y(out_local_master_sel[3])
         );
  AND2X1_HVT U200 ( .A1(master_key[39]), .A2(n256), .Y(
        out_local_master_sel[39]) );
  AND2X1_HVT U201 ( .A1(master_key[38]), .A2(n257), .Y(
        out_local_master_sel[38]) );
  AND2X1_HVT U202 ( .A1(master_key[37]), .A2(n257), .Y(
        out_local_master_sel[37]) );
  AND2X1_HVT U203 ( .A1(master_key[36]), .A2(n257), .Y(
        out_local_master_sel[36]) );
  AND2X1_HVT U204 ( .A1(master_key[35]), .A2(n257), .Y(
        out_local_master_sel[35]) );
  AND2X1_HVT U205 ( .A1(master_key[34]), .A2(n257), .Y(
        out_local_master_sel[34]) );
  AND2X1_HVT U206 ( .A1(master_key[33]), .A2(n257), .Y(
        out_local_master_sel[33]) );
  AND2X1_HVT U207 ( .A1(master_key[32]), .A2(n257), .Y(
        out_local_master_sel[32]) );
  AND2X1_HVT U208 ( .A1(master_key[31]), .A2(n262), .Y(
        out_local_master_sel[31]) );
  AND2X1_HVT U209 ( .A1(master_key[30]), .A2(n164), .Y(
        out_local_master_sel[30]) );
  AND2X1_HVT U210 ( .A1(master_key[2]), .A2(n259), .Y(out_local_master_sel[2])
         );
  AND2X1_HVT U211 ( .A1(master_key[29]), .A2(n262), .Y(
        out_local_master_sel[29]) );
  AND2X1_HVT U212 ( .A1(master_key[28]), .A2(n163), .Y(
        out_local_master_sel[28]) );
  AND2X1_HVT U213 ( .A1(master_key[27]), .A2(n160), .Y(
        out_local_master_sel[27]) );
  AND2X1_HVT U214 ( .A1(master_key[26]), .A2(n159), .Y(
        out_local_master_sel[26]) );
  AND2X1_HVT U215 ( .A1(master_key[25]), .A2(n258), .Y(
        out_local_master_sel[25]) );
  AND2X1_HVT U216 ( .A1(master_key[24]), .A2(n256), .Y(
        out_local_master_sel[24]) );
  AND2X1_HVT U217 ( .A1(master_key[23]), .A2(n160), .Y(
        out_local_master_sel[23]) );
  AND2X1_HVT U218 ( .A1(master_key[22]), .A2(n159), .Y(
        out_local_master_sel[22]) );
  AND2X1_HVT U219 ( .A1(master_key[21]), .A2(n258), .Y(
        out_local_master_sel[21]) );
  AND2X1_HVT U220 ( .A1(master_key[20]), .A2(n256), .Y(
        out_local_master_sel[20]) );
  AND2X1_HVT U221 ( .A1(master_key[1]), .A2(n160), .Y(out_local_master_sel[1])
         );
  AND2X1_HVT U222 ( .A1(master_key[19]), .A2(n159), .Y(
        out_local_master_sel[19]) );
  AND2X1_HVT U223 ( .A1(master_key[18]), .A2(n258), .Y(
        out_local_master_sel[18]) );
  AND2X1_HVT U224 ( .A1(master_key[17]), .A2(n256), .Y(
        out_local_master_sel[17]) );
  AND2X1_HVT U225 ( .A1(master_key[16]), .A2(n255), .Y(
        out_local_master_sel[16]) );
  AND2X1_HVT U226 ( .A1(master_key[15]), .A2(n160), .Y(
        out_local_master_sel[15]) );
  AND2X1_HVT U227 ( .A1(master_key[14]), .A2(n159), .Y(
        out_local_master_sel[14]) );
  AND2X1_HVT U228 ( .A1(master_key[13]), .A2(n258), .Y(
        out_local_master_sel[13]) );
  AND2X1_HVT U229 ( .A1(master_key[12]), .A2(n256), .Y(
        out_local_master_sel[12]) );
  AND2X1_HVT U230 ( .A1(master_key[127]), .A2(n255), .Y(
        out_local_master_sel[127]) );
  AND2X1_HVT U231 ( .A1(master_key[126]), .A2(n255), .Y(
        out_local_master_sel[126]) );
  AND2X1_HVT U232 ( .A1(master_key[125]), .A2(n255), .Y(
        out_local_master_sel[125]) );
  AND2X1_HVT U233 ( .A1(master_key[124]), .A2(n255), .Y(
        out_local_master_sel[124]) );
  AND2X1_HVT U234 ( .A1(master_key[123]), .A2(n255), .Y(
        out_local_master_sel[123]) );
  AND2X1_HVT U235 ( .A1(master_key[122]), .A2(n255), .Y(
        out_local_master_sel[122]) );
  AND2X1_HVT U236 ( .A1(master_key[121]), .A2(n255), .Y(
        out_local_master_sel[121]) );
  AND2X1_HVT U237 ( .A1(master_key[120]), .A2(n261), .Y(
        out_local_master_sel[120]) );
  AND2X1_HVT U238 ( .A1(master_key[11]), .A2(n261), .Y(
        out_local_master_sel[11]) );
  AND2X1_HVT U239 ( .A1(master_key[119]), .A2(n261), .Y(
        out_local_master_sel[119]) );
  AND2X1_HVT U240 ( .A1(master_key[118]), .A2(n261), .Y(
        out_local_master_sel[118]) );
  AND2X1_HVT U241 ( .A1(master_key[117]), .A2(n261), .Y(
        out_local_master_sel[117]) );
  AND2X1_HVT U242 ( .A1(master_key[116]), .A2(n162), .Y(
        out_local_master_sel[116]) );
  AND2X1_HVT U243 ( .A1(master_key[115]), .A2(n161), .Y(
        out_local_master_sel[115]) );
  AND2X1_HVT U244 ( .A1(master_key[114]), .A2(n254), .Y(
        out_local_master_sel[114]) );
  AND2X1_HVT U245 ( .A1(master_key[113]), .A2(n162), .Y(
        out_local_master_sel[113]) );
  AND2X1_HVT U246 ( .A1(master_key[112]), .A2(n161), .Y(
        out_local_master_sel[112]) );
  AND2X1_HVT U247 ( .A1(master_key[111]), .A2(n254), .Y(
        out_local_master_sel[111]) );
  AND2X1_HVT U248 ( .A1(master_key[110]), .A2(n162), .Y(
        out_local_master_sel[110]) );
  AND2X1_HVT U249 ( .A1(master_key[10]), .A2(n260), .Y(
        out_local_master_sel[10]) );
  AND2X1_HVT U250 ( .A1(master_key[109]), .A2(n263), .Y(
        out_local_master_sel[109]) );
  AND2X1_HVT U251 ( .A1(master_key[108]), .A2(n122), .Y(
        out_local_master_sel[108]) );
  AND2X1_HVT U252 ( .A1(master_key[107]), .A2(n123), .Y(
        out_local_master_sel[107]) );
  AND2X1_HVT U253 ( .A1(master_key[106]), .A2(n253), .Y(
        out_local_master_sel[106]) );
  AND2X1_HVT U254 ( .A1(master_key[105]), .A2(n260), .Y(
        out_local_master_sel[105]) );
  AND2X1_HVT U255 ( .A1(master_key[104]), .A2(n263), .Y(
        out_local_master_sel[104]) );
  AND2X1_HVT U256 ( .A1(master_key[103]), .A2(n122), .Y(
        out_local_master_sel[103]) );
  AND2X1_HVT U257 ( .A1(master_key[102]), .A2(n123), .Y(
        out_local_master_sel[102]) );
  AND2X1_HVT U258 ( .A1(master_key[101]), .A2(n253), .Y(
        out_local_master_sel[101]) );
  AND2X1_HVT U259 ( .A1(master_key[100]), .A2(n253), .Y(
        out_local_master_sel[100]) );
  AND2X1_HVT U260 ( .A1(master_key[0]), .A2(n253), .Y(out_local_master_sel[0])
         );
  AO22X1_HVT U263 ( .A1(data_flash[226]), .A2(n297), .A3(account[98]), .A4(
        n289), .Y(out_flash_or_acc_sel[98]) );
  AO22X1_HVT U264 ( .A1(data_flash[225]), .A2(n220), .A3(account[97]), .A4(
        n288), .Y(out_flash_or_acc_sel[97]) );
  AO22X1_HVT U265 ( .A1(data_flash[224]), .A2(n221), .A3(account[96]), .A4(
        n288), .Y(out_flash_or_acc_sel[96]) );
  AO22X1_HVT U269 ( .A1(data_flash[220]), .A2(n221), .A3(account[92]), .A4(
        n176), .Y(out_flash_or_acc_sel[92]) );
  AO22X1_HVT U273 ( .A1(data_flash[217]), .A2(n302), .A3(account[89]), .A4(
        n290), .Y(out_flash_or_acc_sel[89]) );
  AO22X1_HVT U274 ( .A1(data_flash[216]), .A2(n298), .A3(account[88]), .A4(
        n113), .Y(out_flash_or_acc_sel[88]) );
  AO22X1_HVT U275 ( .A1(data_flash[215]), .A2(n25), .A3(account[87]), .A4(n290), .Y(out_flash_or_acc_sel[87]) );
  AO22X1_HVT U276 ( .A1(data_flash[214]), .A2(n223), .A3(account[86]), .A4(
        n167), .Y(out_flash_or_acc_sel[86]) );
  AO22X1_HVT U278 ( .A1(data_flash[212]), .A2(n25), .A3(account[84]), .A4(n184), .Y(out_flash_or_acc_sel[84]) );
  AO22X1_HVT U279 ( .A1(data_flash[211]), .A2(n221), .A3(account[83]), .A4(
        n176), .Y(out_flash_or_acc_sel[83]) );
  AO22X1_HVT U280 ( .A1(data_flash[210]), .A2(n222), .A3(account[82]), .A4(
        n184), .Y(out_flash_or_acc_sel[82]) );
  AO22X1_HVT U281 ( .A1(data_flash[209]), .A2(n296), .A3(account[81]), .A4(n45), .Y(out_flash_or_acc_sel[81]) );
  AO22X1_HVT U282 ( .A1(data_flash[208]), .A2(n299), .A3(account[80]), .A4(
        n113), .Y(out_flash_or_acc_sel[80]) );
  AO22X1_HVT U283 ( .A1(data_flash[135]), .A2(n36), .A3(account[7]), .A4(n45), 
        .Y(out_flash_or_acc_sel[7]) );
  AO22X1_HVT U284 ( .A1(data_flash[207]), .A2(n52), .A3(account[79]), .A4(n45), 
        .Y(out_flash_or_acc_sel[79]) );
  AO22X1_HVT U287 ( .A1(data_flash[204]), .A2(n221), .A3(account[76]), .A4(n45), .Y(out_flash_or_acc_sel[76]) );
  AO22X1_HVT U288 ( .A1(data_flash[203]), .A2(n298), .A3(account[75]), .A4(n45), .Y(out_flash_or_acc_sel[75]) );
  AO22X1_HVT U291 ( .A1(data_flash[200]), .A2(n303), .A3(account[72]), .A4(n45), .Y(out_flash_or_acc_sel[72]) );
  AO22X1_HVT U292 ( .A1(data_flash[199]), .A2(n302), .A3(account[71]), .A4(n45), .Y(out_flash_or_acc_sel[71]) );
  AO22X1_HVT U293 ( .A1(data_flash[198]), .A2(n222), .A3(account[70]), .A4(n62), .Y(out_flash_or_acc_sel[70]) );
  AO22X1_HVT U294 ( .A1(data_flash[134]), .A2(n52), .A3(account[6]), .A4(n78), 
        .Y(out_flash_or_acc_sel[6]) );
  AO22X1_HVT U295 ( .A1(data_flash[197]), .A2(n25), .A3(account[69]), .A4(n288), .Y(out_flash_or_acc_sel[69]) );
  AO22X1_HVT U296 ( .A1(data_flash[196]), .A2(n303), .A3(account[68]), .A4(n62), .Y(out_flash_or_acc_sel[68]) );
  AO22X1_HVT U297 ( .A1(data_flash[195]), .A2(n297), .A3(account[67]), .A4(
        n184), .Y(out_flash_or_acc_sel[67]) );
  AO22X1_HVT U298 ( .A1(data_flash[194]), .A2(n294), .A3(account[66]), .A4(
        n288), .Y(out_flash_or_acc_sel[66]) );
  AO22X1_HVT U302 ( .A1(data_flash[190]), .A2(n220), .A3(account[62]), .A4(
        n289), .Y(out_flash_or_acc_sel[62]) );
  AO22X1_HVT U303 ( .A1(data_flash[189]), .A2(n301), .A3(account[61]), .A4(
        n289), .Y(out_flash_or_acc_sel[61]) );
  AO22X1_HVT U304 ( .A1(data_flash[188]), .A2(n303), .A3(account[60]), .A4(
        n288), .Y(out_flash_or_acc_sel[60]) );
  AO22X1_HVT U306 ( .A1(data_flash[187]), .A2(n298), .A3(account[59]), .A4(
        n291), .Y(out_flash_or_acc_sel[59]) );
  AO22X1_HVT U307 ( .A1(data_flash[186]), .A2(n251), .A3(account[58]), .A4(
        n286), .Y(out_flash_or_acc_sel[58]) );
  AO22X1_HVT U308 ( .A1(data_flash[185]), .A2(n302), .A3(account[57]), .A4(n69), .Y(out_flash_or_acc_sel[57]) );
  AO22X1_HVT U309 ( .A1(data_flash[184]), .A2(n36), .A3(account[56]), .A4(n290), .Y(out_flash_or_acc_sel[56]) );
  AO22X1_HVT U311 ( .A1(data_flash[182]), .A2(n223), .A3(account[54]), .A4(
        n167), .Y(out_flash_or_acc_sel[54]) );
  AO22X1_HVT U312 ( .A1(data_flash[181]), .A2(n297), .A3(account[53]), .A4(
        n290), .Y(out_flash_or_acc_sel[53]) );
  AO22X1_HVT U313 ( .A1(data_flash[180]), .A2(n251), .A3(account[52]), .A4(n62), .Y(out_flash_or_acc_sel[52]) );
  AO22X1_HVT U314 ( .A1(data_flash[179]), .A2(n223), .A3(account[51]), .A4(n69), .Y(out_flash_or_acc_sel[51]) );
  AO22X1_HVT U315 ( .A1(data_flash[178]), .A2(n223), .A3(account[50]), .A4(
        n168), .Y(out_flash_or_acc_sel[50]) );
  AO22X1_HVT U316 ( .A1(data_flash[132]), .A2(n220), .A3(account[4]), .A4(n168), .Y(out_flash_or_acc_sel[4]) );
  AO22X1_HVT U318 ( .A1(data_flash[176]), .A2(n303), .A3(account[48]), .A4(
        n168), .Y(out_flash_or_acc_sel[48]) );
  AO22X1_HVT U319 ( .A1(data_flash[175]), .A2(n220), .A3(account[47]), .A4(n62), .Y(out_flash_or_acc_sel[47]) );
  AO22X1_HVT U320 ( .A1(data_flash[174]), .A2(n297), .A3(account[46]), .A4(n69), .Y(out_flash_or_acc_sel[46]) );
  AO22X1_HVT U321 ( .A1(data_flash[173]), .A2(n52), .A3(account[45]), .A4(n291), .Y(out_flash_or_acc_sel[45]) );
  AO22X1_HVT U322 ( .A1(data_flash[172]), .A2(n301), .A3(account[44]), .A4(
        n290), .Y(out_flash_or_acc_sel[44]) );
  AO22X1_HVT U323 ( .A1(data_flash[171]), .A2(n303), .A3(account[43]), .A4(
        n286), .Y(out_flash_or_acc_sel[43]) );
  AO22X1_HVT U324 ( .A1(data_flash[170]), .A2(n12), .A3(account[42]), .A4(n291), .Y(out_flash_or_acc_sel[42]) );
  AO22X1_HVT U327 ( .A1(data_flash[131]), .A2(n251), .A3(account[3]), .A4(n167), .Y(out_flash_or_acc_sel[3]) );
  AO22X1_HVT U328 ( .A1(data_flash[167]), .A2(n296), .A3(account[39]), .A4(n62), .Y(out_flash_or_acc_sel[39]) );
  AO22X1_HVT U329 ( .A1(data_flash[166]), .A2(n296), .A3(account[38]), .A4(
        n286), .Y(out_flash_or_acc_sel[38]) );
  AO22X1_HVT U332 ( .A1(data_flash[163]), .A2(n299), .A3(account[35]), .A4(
        n291), .Y(out_flash_or_acc_sel[35]) );
  AO22X1_HVT U333 ( .A1(data_flash[162]), .A2(n251), .A3(account[34]), .A4(
        n291), .Y(out_flash_or_acc_sel[34]) );
  AO22X1_HVT U336 ( .A1(data_flash[159]), .A2(n301), .A3(account[31]), .A4(
        n286), .Y(out_flash_or_acc_sel[31]) );
  AO22X1_HVT U337 ( .A1(data_flash[158]), .A2(n301), .A3(account[30]), .A4(
        n168), .Y(out_flash_or_acc_sel[30]) );
  AO22X1_HVT U340 ( .A1(data_flash[156]), .A2(n222), .A3(account[28]), .A4(
        n119), .Y(out_flash_or_acc_sel[28]) );
  AO22X1_HVT U341 ( .A1(data_flash[155]), .A2(n297), .A3(account[27]), .A4(n78), .Y(out_flash_or_acc_sel[27]) );
  AO22X1_HVT U343 ( .A1(data_flash[153]), .A2(n296), .A3(account[25]), .A4(n78), .Y(out_flash_or_acc_sel[25]) );
  AO22X1_HVT U344 ( .A1(data_flash[152]), .A2(n36), .A3(account[24]), .A4(n155), .Y(out_flash_or_acc_sel[24]) );
  AO22X1_HVT U345 ( .A1(data_flash[151]), .A2(n156), .A3(account[23]), .A4(n78), .Y(out_flash_or_acc_sel[23]) );
  AO22X1_HVT U346 ( .A1(data_flash[150]), .A2(n156), .A3(account[22]), .A4(
        n184), .Y(out_flash_or_acc_sel[22]) );
  AO22X1_HVT U348 ( .A1(data_flash[148]), .A2(n299), .A3(account[20]), .A4(n78), .Y(out_flash_or_acc_sel[20]) );
  AO22X1_HVT U351 ( .A1(data_flash[146]), .A2(n223), .A3(account[18]), .A4(
        n289), .Y(out_flash_or_acc_sel[18]) );
  AO22X1_HVT U352 ( .A1(data_flash[145]), .A2(n297), .A3(account[17]), .A4(
        n288), .Y(out_flash_or_acc_sel[17]) );
  AO22X1_HVT U353 ( .A1(n36), .A2(data_flash[144]), .A3(account[16]), .A4(n289), .Y(out_flash_or_acc_sel[16]) );
  AO22X1_HVT U354 ( .A1(data_flash[143]), .A2(n12), .A3(account[15]), .A4(n289), .Y(out_flash_or_acc_sel[15]) );
  AO22X1_HVT U355 ( .A1(data_flash[142]), .A2(n296), .A3(account[14]), .A4(n78), .Y(out_flash_or_acc_sel[14]) );
  AO22X1_HVT U359 ( .A1(data_flash[254]), .A2(n12), .A3(account[126]), .A4(n62), .Y(out_flash_or_acc_sel[126]) );
  AO22X1_HVT U362 ( .A1(data_flash[251]), .A2(n301), .A3(account[123]), .A4(
        n184), .Y(out_flash_or_acc_sel[123]) );
  AO22X1_HVT U363 ( .A1(data_flash[250]), .A2(n299), .A3(account[122]), .A4(
        n184), .Y(out_flash_or_acc_sel[122]) );
  AO22X1_HVT U364 ( .A1(data_flash[249]), .A2(n223), .A3(account[121]), .A4(
        n62), .Y(out_flash_or_acc_sel[121]) );
  AO22X1_HVT U367 ( .A1(data_flash[247]), .A2(n301), .A3(account[119]), .A4(
        n291), .Y(out_flash_or_acc_sel[119]) );
  AO22X1_HVT U368 ( .A1(data_flash[246]), .A2(n296), .A3(account[118]), .A4(
        n167), .Y(out_flash_or_acc_sel[118]) );
  AO22X1_HVT U369 ( .A1(data_flash[245]), .A2(n25), .A3(account[117]), .A4(
        n290), .Y(out_flash_or_acc_sel[117]) );
  AO22X1_HVT U373 ( .A1(data_flash[241]), .A2(n302), .A3(account[113]), .A4(
        n168), .Y(out_flash_or_acc_sel[113]) );
  AO22X1_HVT U374 ( .A1(data_flash[240]), .A2(n298), .A3(account[112]), .A4(
        n167), .Y(out_flash_or_acc_sel[112]) );
  AO22X1_HVT U375 ( .A1(data_flash[239]), .A2(n52), .A3(account[111]), .A4(
        n290), .Y(out_flash_or_acc_sel[111]) );
  AO22X1_HVT U377 ( .A1(data_flash[138]), .A2(n25), .A3(account[10]), .A4(n167), .Y(out_flash_or_acc_sel[10]) );
  AO22X1_HVT U379 ( .A1(data_flash[236]), .A2(n294), .A3(account[108]), .A4(
        n286), .Y(out_flash_or_acc_sel[108]) );
  AO22X1_HVT U380 ( .A1(data_flash[235]), .A2(n303), .A3(account[107]), .A4(
        n69), .Y(out_flash_or_acc_sel[107]) );
  AO22X1_HVT U381 ( .A1(data_flash[234]), .A2(n221), .A3(account[106]), .A4(
        n286), .Y(out_flash_or_acc_sel[106]) );
  AO22X1_HVT U383 ( .A1(data_flash[232]), .A2(n52), .A3(account[104]), .A4(
        n168), .Y(out_flash_or_acc_sel[104]) );
  AO22X1_HVT U384 ( .A1(data_flash[231]), .A2(n298), .A3(account[103]), .A4(
        n168), .Y(out_flash_or_acc_sel[103]) );
  AO22X1_HVT U385 ( .A1(data_flash[230]), .A2(n294), .A3(account[102]), .A4(
        n168), .Y(out_flash_or_acc_sel[102]) );
  AO22X1_HVT U386 ( .A1(data_flash[229]), .A2(n302), .A3(account[101]), .A4(
        n290), .Y(out_flash_or_acc_sel[101]) );
  AO22X1_HVT U387 ( .A1(data_flash[228]), .A2(n25), .A3(account[100]), .A4(n69), .Y(out_flash_or_acc_sel[100]) );
  AO22X1_HVT U388 ( .A1(data_flash[128]), .A2(n298), .A3(account[0]), .A4(n69), 
        .Y(out_flash_or_acc_sel[0]) );
  AO22X1_HVT U391 ( .A1(n244), .A2(match_add[1]), .A3(n228), .A4(write_add[1]), 
        .Y(add_flash[1]) );
  AO22X1_HVT U392 ( .A1(boot_lood), .A2(match_add[0]), .A3(n306), .A4(
        write_add[0]), .Y(add_flash[0]) );
  reg_D_0 reg_flash_or_acc ( .clk(clk), .rst(n304), .enable(flash_or_acc_reg), 
        .in({out_flash_or_acc_sel[127:65], n216, out_flash_or_acc_sel[63:56], 
        n175, out_flash_or_acc_sel[54:34], n183, out_flash_or_acc_sel[32:14], 
        n118, out_flash_or_acc_sel[12:0]}), .out(out_reg_flash_or_acc) );
  reg_D_6 reg_flash_account ( .clk(clk), .rst(n304), .enable(flash_acc_reg), 
        .in(out_reg_flash_or_acc), .out(write_data_flash[255:128]) );
  reg_D_5 reg_flash_pass ( .clk(clk), .rst(n304), .enable(flash_pass_reg), 
        .in(out_encryption), .out(write_data_flash[127:0]) );
  reg_D_4 reg_pass_enc ( .clk(clk), .rst(n304), .enable(pass_enc_reg), .in(
        data_flash[127:0]), .out(out_reg_pass_enc) );
  reg_D_3 reg_plain_reg ( .clk(clk), .rst(n304), .enable(plain_reg), .in({
        out_new_old_pass_sel[127:44], n39, out_new_old_pass_sel[42:9], n55, 
        out_new_old_pass_sel[7:2], n26, out_new_old_pass_sel[0]}), .out(
        out_reg_plain_reg) );
  reg_D_2 reg_local_master ( .clk(clk), .rst(n304), .enable(local_master_reg), 
        .in(out_local_master_sel), .out(out_local_master_reg) );
  reg_D_1 reg_out_reg ( .clk(clk), .rst(n304), .enable(out_reg), .in(
        out_encryption), .out(final_output) );
  cam_DATA_WIDTH128_ADDR_WIDTH4 cam_inst ( .clk(clk), .rst(n304), .start(
        cam_start), .write_enable(write_en), .din({
        out_reg_flash_or_acc[127:125], n80, out_reg_flash_or_acc[123:121], n81, 
        out_reg_flash_or_acc[119:117], n82, out_reg_flash_or_acc[115:113], n83, 
        out_reg_flash_or_acc[111:109], n84, out_reg_flash_or_acc[107:105], n85, 
        out_reg_flash_or_acc[103:101], n86, out_reg_flash_or_acc[99:97], n87, 
        out_reg_flash_or_acc[95:93], n88, out_reg_flash_or_acc[91:89], n89, 
        out_reg_flash_or_acc[87:85], n90, out_reg_flash_or_acc[83:81], n91, 
        out_reg_flash_or_acc[79:77], n92, out_reg_flash_or_acc[75:73], n93, 
        out_reg_flash_or_acc[71:69], n94, out_reg_flash_or_acc[67:65], n95, 
        out_reg_flash_or_acc[63:61], n96, out_reg_flash_or_acc[59:57], n97, 
        out_reg_flash_or_acc[55:53], n98, out_reg_flash_or_acc[51:49], n99, 
        out_reg_flash_or_acc[47:45], n100, out_reg_flash_or_acc[43:41], n101, 
        out_reg_flash_or_acc[39:37], n102, out_reg_flash_or_acc[35:33], n103, 
        out_reg_flash_or_acc[31:29], n104, out_reg_flash_or_acc[27:25], n105, 
        out_reg_flash_or_acc[23:21], n106, out_reg_flash_or_acc[19:17], n107, 
        out_reg_flash_or_acc[15:13], n108, out_reg_flash_or_acc[11:9], n109, 
        out_reg_flash_or_acc[7:5], n110, out_reg_flash_or_acc[3:1], n79}), 
        .write_addr(write_add), .match(match), .match_addr(match_add) );
  aes ENC ( .plaintext(out_reg_plain_reg), .key(out_local_master_reg), .clk(
        clk), .reset(n304), .start(start_enc), .cipher_text(out_encryption), 
        .ready(ready_encryption) );
  inv_aes DEC ( .clk(clk), .rest(n304), .start(start_dec), .plaintext1(
        out_reg_pass_enc), .local_key({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cipher_text(out_decry), .done(dec_done) );
  NAND2X0_HVT U2 ( .A1(data_flash[223]), .A2(n222), .Y(n1) );
  NAND2X0_HVT U3 ( .A1(account[95]), .A2(n289), .Y(n2) );
  NAND2X0_HVT U4 ( .A1(n1), .A2(n2), .Y(out_flash_or_acc_sel[95]) );
  INVX0_HVT U5 ( .A(n245), .Y(n217) );
  NAND2X0_HVT U16 ( .A1(data_flash[227]), .A2(n52), .Y(n3) );
  NAND2X0_HVT U27 ( .A1(account[99]), .A2(n62), .Y(n4) );
  NAND2X0_HVT U38 ( .A1(n3), .A2(n4), .Y(out_flash_or_acc_sel[99]) );
  NAND2X0_HVT U58 ( .A1(data_flash[244]), .A2(n302), .Y(n5) );
  NAND2X0_HVT U60 ( .A1(account[116]), .A2(n62), .Y(n6) );
  NAND2X0_HVT U63 ( .A1(n5), .A2(n6), .Y(out_flash_or_acc_sel[116]) );
  NAND2X0_HVT U64 ( .A1(data_flash[191]), .A2(n294), .Y(n7) );
  NAND2X0_HVT U65 ( .A1(account[63]), .A2(n78), .Y(n8) );
  NAND2X0_HVT U66 ( .A1(n7), .A2(n8), .Y(out_flash_or_acc_sel[63]) );
  INVX0_HVT U67 ( .A(n186), .Y(n262) );
  INVX1_HVT U71 ( .A(n203), .Y(n196) );
  INVX0_HVT U89 ( .A(n18), .Y(n9) );
  INVX0_HVT U93 ( .A(n17), .Y(n18) );
  IBUFFX2_HVT U95 ( .A(n67), .Y(n10) );
  NBUFFX2_HVT U132 ( .A(n203), .Y(n11) );
  INVX0_HVT U261 ( .A(n227), .Y(n302) );
  NBUFFX2_HVT U262 ( .A(n20), .Y(n25) );
  INVX0_HVT U266 ( .A(n136), .Y(n12) );
  INVX0_HVT U267 ( .A(n226), .Y(n13) );
  INVX0_HVT U268 ( .A(n13), .Y(n14) );
  INVX0_HVT U270 ( .A(n208), .Y(n15) );
  INVX0_HVT U271 ( .A(n15), .Y(n16) );
  INVX0_HVT U272 ( .A(n192), .Y(n17) );
  NBUFFX2_HVT U277 ( .A(n20), .Y(n52) );
  NBUFFX2_HVT U285 ( .A(n278), .Y(n19) );
  INVX0_HVT U286 ( .A(n14), .Y(n20) );
  INVX0_HVT U289 ( .A(n285), .Y(n227) );
  INVX0_HVT U290 ( .A(n267), .Y(n278) );
  INVX0_HVT U299 ( .A(n227), .Y(n303) );
  NBUFFX2_HVT U300 ( .A(flash_or_acc_sel), .Y(n113) );
  INVX0_HVT U301 ( .A(n33), .Y(n301) );
  INVX0_HVT U305 ( .A(n33), .Y(n297) );
  NAND2X0_HVT U310 ( .A1(data_flash[141]), .A2(n202), .Y(n21) );
  NAND2X0_HVT U317 ( .A1(account[13]), .A2(n119), .Y(n22) );
  NAND2X0_HVT U325 ( .A1(n21), .A2(n22), .Y(n118) );
  IBUFFX2_HVT U326 ( .A(n294), .Y(n119) );
  NAND2X0_HVT U330 ( .A1(data_flash[164]), .A2(n223), .Y(n23) );
  NAND2X0_HVT U331 ( .A1(account[36]), .A2(n291), .Y(n24) );
  NAND2X0_HVT U334 ( .A1(n23), .A2(n24), .Y(out_flash_or_acc_sel[36]) );
  INVX0_HVT U335 ( .A(n33), .Y(n223) );
  INVX0_HVT U338 ( .A(n249), .Y(n228) );
  INVX0_HVT U339 ( .A(local_master_sel), .Y(n264) );
  INVX0_HVT U342 ( .A(n77), .Y(n210) );
  INVX0_HVT U347 ( .A(n76), .Y(n282) );
  INVX0_HVT U349 ( .A(n224), .Y(n280) );
  INVX0_HVT U350 ( .A(n33), .Y(n296) );
  INVX0_HVT U356 ( .A(n252), .Y(n291) );
  AO22X1_HVT U357 ( .A1(out_decry[1]), .A2(n138), .A3(pass[1]), .A4(n209), .Y(
        n26) );
  INVX0_HVT U358 ( .A(n202), .Y(n78) );
  INVX0_HVT U360 ( .A(n75), .Y(n27) );
  NBUFFX2_HVT U361 ( .A(n224), .Y(n75) );
  INVX0_HVT U365 ( .A(n113), .Y(n252) );
  NAND2X0_HVT U366 ( .A1(data_flash[243]), .A2(n303), .Y(n28) );
  NAND2X0_HVT U370 ( .A1(account[115]), .A2(n167), .Y(n29) );
  NAND2X0_HVT U371 ( .A1(n28), .A2(n29), .Y(out_flash_or_acc_sel[115]) );
  IBUFFX2_HVT U372 ( .A(n252), .Y(n167) );
  NAND2X0_HVT U376 ( .A1(data_flash[133]), .A2(n221), .Y(n30) );
  NAND2X0_HVT U378 ( .A1(account[5]), .A2(n167), .Y(n31) );
  NAND2X0_HVT U382 ( .A1(n30), .A2(n31), .Y(out_flash_or_acc_sel[5]) );
  INVX0_HVT U389 ( .A(n227), .Y(n221) );
  INVX0_HVT U390 ( .A(n226), .Y(n32) );
  INVX1_HVT U393 ( .A(n32), .Y(n33) );
  NAND2X0_HVT U394 ( .A1(data_flash[177]), .A2(n294), .Y(n34) );
  NAND2X0_HVT U395 ( .A1(account[49]), .A2(n69), .Y(n35) );
  NAND2X0_HVT U396 ( .A1(n34), .A2(n35), .Y(out_flash_or_acc_sel[49]) );
  INVX0_HVT U397 ( .A(n227), .Y(n294) );
  IBUFFX2_HVT U398 ( .A(n136), .Y(n251) );
  INVX0_HVT U399 ( .A(n136), .Y(n299) );
  NBUFFX2_HVT U400 ( .A(n300), .Y(n36) );
  NAND2X0_HVT U401 ( .A1(data_flash[157]), .A2(n297), .Y(n37) );
  NAND2X0_HVT U402 ( .A1(account[29]), .A2(n69), .Y(n38) );
  NAND2X0_HVT U403 ( .A1(n37), .A2(n38), .Y(out_flash_or_acc_sel[29]) );
  INVX0_HVT U404 ( .A(n32), .Y(n69) );
  INVX1_HVT U405 ( .A(n300), .Y(n136) );
  AO22X1_HVT U406 ( .A1(out_decry[43]), .A2(n266), .A3(pass[43]), .A4(n68), 
        .Y(n39) );
  IBUFFX2_HVT U407 ( .A(n274), .Y(n147) );
  INVX0_HVT U408 ( .A(n224), .Y(n284) );
  NAND2X0_HVT U409 ( .A1(data_flash[160]), .A2(n220), .Y(n40) );
  NAND2X0_HVT U410 ( .A1(account[32]), .A2(n286), .Y(n41) );
  NAND2X0_HVT U411 ( .A1(n40), .A2(n41), .Y(out_flash_or_acc_sel[32]) );
  INVX0_HVT U412 ( .A(n252), .Y(n168) );
  INVX0_HVT U413 ( .A(n75), .Y(n42) );
  NAND2X0_HVT U414 ( .A1(data_flash[161]), .A2(n202), .Y(n43) );
  NAND2X0_HVT U415 ( .A1(account[33]), .A2(n184), .Y(n44) );
  NAND2X0_HVT U416 ( .A1(n43), .A2(n44), .Y(n183) );
  INVX0_HVT U417 ( .A(n244), .Y(n245) );
  NBUFFX2_HVT U418 ( .A(n155), .Y(n45) );
  INVX1_HVT U419 ( .A(n295), .Y(n292) );
  INVX0_HVT U420 ( .A(n196), .Y(n192) );
  IBUFFX2_HVT U421 ( .A(n227), .Y(n298) );
  INVX0_HVT U422 ( .A(n225), .Y(n295) );
  INVX0_HVT U423 ( .A(n295), .Y(n184) );
  NAND2X0_HVT U424 ( .A1(data_flash[255]), .A2(n12), .Y(n46) );
  NAND2X0_HVT U425 ( .A1(account[127]), .A2(n288), .Y(n47) );
  NAND2X0_HVT U426 ( .A1(n46), .A2(n47), .Y(out_flash_or_acc_sel[127]) );
  NAND2X0_HVT U427 ( .A1(data_flash[136]), .A2(n220), .Y(n48) );
  NAND2X0_HVT U428 ( .A1(account[8]), .A2(n184), .Y(n49) );
  NAND2X0_HVT U429 ( .A1(n48), .A2(n49), .Y(out_flash_or_acc_sel[8]) );
  IBUFFX2_HVT U430 ( .A(n196), .Y(n73) );
  NAND2X0_HVT U431 ( .A1(n217), .A2(match_add[3]), .Y(n50) );
  NAND2X0_HVT U432 ( .A1(write_add[3]), .A2(n228), .Y(n51) );
  NAND2X0_HVT U433 ( .A1(n50), .A2(n51), .Y(add_flash[3]) );
  INVX0_HVT U434 ( .A(n250), .Y(n244) );
  NAND2X0_HVT U435 ( .A1(data_flash[222]), .A2(n301), .Y(n53) );
  NAND2X0_HVT U436 ( .A1(account[94]), .A2(n184), .Y(n54) );
  NAND2X0_HVT U437 ( .A1(n53), .A2(n54), .Y(out_flash_or_acc_sel[94]) );
  INVX0_HVT U438 ( .A(n121), .Y(n224) );
  INVX1_HVT U439 ( .A(out_decry[6]), .Y(n72) );
  INVX1_HVT U440 ( .A(out_decry[7]), .Y(n234) );
  INVX1_HVT U441 ( .A(out_decry[18]), .Y(n60) );
  INVX1_HVT U442 ( .A(out_decry[44]), .Y(n198) );
  INVX1_HVT U443 ( .A(out_decry[45]), .Y(n212) );
  INVX1_HVT U444 ( .A(out_decry[46]), .Y(n194) );
  INVX0_HVT U445 ( .A(n267), .Y(n209) );
  INVX0_HVT U446 ( .A(n76), .Y(n277) );
  INVX0_HVT U447 ( .A(local_master_sel), .Y(n186) );
  INVX0_HVT U448 ( .A(n137), .Y(n68) );
  INVX0_HVT U449 ( .A(n77), .Y(n269) );
  INVX1_HVT U450 ( .A(account[21]), .Y(n126) );
  INVX1_HVT U451 ( .A(account[41]), .Y(n70) );
  INVX1_HVT U452 ( .A(account[65]), .Y(n129) );
  INVX0_HVT U453 ( .A(n136), .Y(n220) );
  INVX1_HVT U454 ( .A(account[105]), .Y(n241) );
  INVX1_HVT U455 ( .A(pass[3]), .Y(n150) );
  INVX1_HVT U456 ( .A(out_decry[3]), .Y(n149) );
  INVX1_HVT U457 ( .A(pass[4]), .Y(n201) );
  INVX1_HVT U458 ( .A(out_decry[4]), .Y(n200) );
  INVX0_HVT U459 ( .A(n71), .Y(out_new_old_pass_sel[6]) );
  INVX1_HVT U460 ( .A(pass[6]), .Y(n74) );
  INVX1_HVT U461 ( .A(pass[7]), .Y(n235) );
  INVX1_HVT U462 ( .A(pass[9]), .Y(n65) );
  INVX1_HVT U463 ( .A(out_decry[9]), .Y(n64) );
  INVX0_HVT U464 ( .A(n59), .Y(out_new_old_pass_sel[18]) );
  INVX1_HVT U465 ( .A(pass[18]), .Y(n61) );
  INVX1_HVT U466 ( .A(pass[23]), .Y(n58) );
  INVX1_HVT U467 ( .A(out_decry[23]), .Y(n57) );
  INVX1_HVT U468 ( .A(pass[44]), .Y(n199) );
  INVX1_HVT U469 ( .A(pass[45]), .Y(n213) );
  INVX0_HVT U470 ( .A(n193), .Y(out_new_old_pass_sel[46]) );
  INVX1_HVT U471 ( .A(pass[46]), .Y(n195) );
  INVX1_HVT U472 ( .A(pass[47]), .Y(n190) );
  INVX1_HVT U473 ( .A(out_decry[47]), .Y(n189) );
  INVX1_HVT U474 ( .A(pass[51]), .Y(n182) );
  INVX1_HVT U475 ( .A(out_decry[51]), .Y(n181) );
  INVX1_HVT U476 ( .A(account[1]), .Y(n243) );
  INVX1_HVT U477 ( .A(account[37]), .Y(n158) );
  INVX1_HVT U478 ( .A(account[124]), .Y(n128) );
  INVX0_HVT U479 ( .A(n202), .Y(n288) );
  INVX0_HVT U480 ( .A(n75), .Y(n281) );
  INVX0_HVT U481 ( .A(n32), .Y(n290) );
  AO22X1_HVT U482 ( .A1(out_decry[8]), .A2(n137), .A3(pass[8]), .A4(n27), .Y(
        n55) );
  INVX0_HVT U483 ( .A(n67), .Y(n148) );
  INVX0_HVT U484 ( .A(n75), .Y(n56) );
  OAI22X1_HVT U485 ( .A1(n57), .A2(n77), .A3(n58), .A4(n63), .Y(
        out_new_old_pass_sel[23]) );
  OA22X1_HVT U486 ( .A1(n60), .A2(n276), .A3(n61), .A4(n63), .Y(n59) );
  INVX0_HVT U487 ( .A(n275), .Y(n191) );
  NBUFFX2_HVT U488 ( .A(n113), .Y(n62) );
  INVX0_HVT U489 ( .A(n279), .Y(n63) );
  INVX0_HVT U490 ( .A(n252), .Y(n286) );
  OAI22X1_HVT U491 ( .A1(n64), .A2(n279), .A3(n65), .A4(n63), .Y(
        out_new_old_pass_sel[9]) );
  INVX0_HVT U492 ( .A(n266), .Y(n66) );
  NBUFFX2_HVT U493 ( .A(n274), .Y(n67) );
  IBUFFX2_HVT U494 ( .A(new_old_pass_sel), .Y(n274) );
  INVX0_HVT U495 ( .A(n76), .Y(n279) );
  INVX0_HVT U496 ( .A(n266), .Y(n276) );
  IBUFFX2_HVT U497 ( .A(n121), .Y(n137) );
  IBUFFX2_HVT U498 ( .A(n32), .Y(n287) );
  OR2X2_HVT U499 ( .A1(n70), .A2(n156), .Y(n180) );
  OA22X1_HVT U500 ( .A1(n72), .A2(n279), .A3(n74), .A4(n196), .Y(n71) );
  NBUFFX2_HVT U501 ( .A(n225), .Y(n226) );
  INVX0_HVT U502 ( .A(n197), .Y(out_new_old_pass_sel[44]) );
  OA22X1_HVT U503 ( .A1(n198), .A2(n66), .A3(n199), .A4(n17), .Y(n197) );
  NBUFFX2_HVT U504 ( .A(n120), .Y(n76) );
  INVX0_HVT U505 ( .A(n147), .Y(n77) );
  NBUFFX2_HVT U506 ( .A(out_reg_flash_or_acc[116]), .Y(n82) );
  NBUFFX2_HVT U507 ( .A(out_reg_flash_or_acc[108]), .Y(n84) );
  NBUFFX2_HVT U508 ( .A(out_reg_flash_or_acc[100]), .Y(n86) );
  NBUFFX2_HVT U509 ( .A(out_reg_flash_or_acc[68]), .Y(n94) );
  NBUFFX2_HVT U510 ( .A(out_reg_flash_or_acc[64]), .Y(n95) );
  NBUFFX2_HVT U511 ( .A(out_reg_flash_or_acc[52]), .Y(n98) );
  NBUFFX2_HVT U512 ( .A(out_reg_flash_or_acc[44]), .Y(n100) );
  NBUFFX2_HVT U513 ( .A(out_reg_flash_or_acc[24]), .Y(n105) );
  NBUFFX2_HVT U514 ( .A(out_reg_flash_or_acc[20]), .Y(n106) );
  INVX0_HVT U515 ( .A(new_old_pass_sel), .Y(n246) );
  NBUFFX2_HVT U516 ( .A(out_reg_flash_or_acc[0]), .Y(n79) );
  NBUFFX2_HVT U517 ( .A(out_reg_flash_or_acc[124]), .Y(n80) );
  NBUFFX2_HVT U518 ( .A(out_reg_flash_or_acc[120]), .Y(n81) );
  NBUFFX2_HVT U519 ( .A(out_reg_flash_or_acc[112]), .Y(n83) );
  NBUFFX2_HVT U520 ( .A(out_reg_flash_or_acc[104]), .Y(n85) );
  NBUFFX2_HVT U521 ( .A(out_reg_flash_or_acc[96]), .Y(n87) );
  NBUFFX2_HVT U522 ( .A(out_reg_flash_or_acc[92]), .Y(n88) );
  NBUFFX2_HVT U523 ( .A(out_reg_flash_or_acc[88]), .Y(n89) );
  NBUFFX2_HVT U524 ( .A(out_reg_flash_or_acc[84]), .Y(n90) );
  NBUFFX2_HVT U525 ( .A(out_reg_flash_or_acc[80]), .Y(n91) );
  NBUFFX2_HVT U526 ( .A(out_reg_flash_or_acc[76]), .Y(n92) );
  NBUFFX2_HVT U527 ( .A(out_reg_flash_or_acc[72]), .Y(n93) );
  NBUFFX2_HVT U528 ( .A(out_reg_flash_or_acc[60]), .Y(n96) );
  NBUFFX2_HVT U529 ( .A(out_reg_flash_or_acc[56]), .Y(n97) );
  NBUFFX2_HVT U530 ( .A(out_reg_flash_or_acc[48]), .Y(n99) );
  NBUFFX2_HVT U531 ( .A(out_reg_flash_or_acc[40]), .Y(n101) );
  NBUFFX2_HVT U532 ( .A(out_reg_flash_or_acc[36]), .Y(n102) );
  NBUFFX2_HVT U533 ( .A(out_reg_flash_or_acc[32]), .Y(n103) );
  NBUFFX2_HVT U534 ( .A(out_reg_flash_or_acc[28]), .Y(n104) );
  NBUFFX2_HVT U535 ( .A(out_reg_flash_or_acc[16]), .Y(n107) );
  NBUFFX2_HVT U536 ( .A(out_reg_flash_or_acc[12]), .Y(n108) );
  NBUFFX2_HVT U537 ( .A(out_reg_flash_or_acc[8]), .Y(n109) );
  NBUFFX2_HVT U538 ( .A(out_reg_flash_or_acc[4]), .Y(n110) );
  IBUFFX2_HVT U539 ( .A(n202), .Y(n293) );
  NBUFFX2_HVT U540 ( .A(n295), .Y(n202) );
  NAND2X0_HVT U541 ( .A1(data_flash[140]), .A2(n296), .Y(n111) );
  NAND2X0_HVT U542 ( .A1(account[12]), .A2(n293), .Y(n112) );
  NAND2X0_HVT U543 ( .A1(n111), .A2(n112), .Y(out_flash_or_acc_sel[12]) );
  NAND2X0_HVT U544 ( .A1(data_flash[213]), .A2(n223), .Y(n114) );
  NAND2X0_HVT U545 ( .A1(account[85]), .A2(n287), .Y(n115) );
  NAND2X0_HVT U546 ( .A1(n114), .A2(n115), .Y(out_flash_or_acc_sel[85]) );
  NAND2X0_HVT U547 ( .A1(data_flash[192]), .A2(n302), .Y(n116) );
  NAND2X0_HVT U548 ( .A1(account[64]), .A2(n227), .Y(n117) );
  NAND2X0_HVT U549 ( .A1(n116), .A2(n117), .Y(n216) );
  INVX0_HVT U550 ( .A(n246), .Y(n120) );
  INVX0_HVT U551 ( .A(n120), .Y(n121) );
  INVX0_HVT U552 ( .A(n185), .Y(n122) );
  INVX0_HVT U553 ( .A(n185), .Y(n123) );
  NAND2X0_HVT U554 ( .A1(data_flash[154]), .A2(n156), .Y(n124) );
  NAND2X0_HVT U555 ( .A1(account[26]), .A2(n293), .Y(n125) );
  NAND2X0_HVT U556 ( .A1(n124), .A2(n125), .Y(out_flash_or_acc_sel[26]) );
  INVX0_HVT U557 ( .A(n202), .Y(n289) );
  IBUFFX2_HVT U558 ( .A(n121), .Y(n138) );
  OR2X1_HVT U559 ( .A1(n126), .A2(n296), .Y(n166) );
  INVX0_HVT U560 ( .A(data_flash[252]), .Y(n127) );
  NAND2X0_HVT U561 ( .A1(data_flash[253]), .A2(n12), .Y(n134) );
  OAI22X1_HVT U562 ( .A1(n292), .A2(n127), .A3(n128), .A4(n156), .Y(
        out_flash_or_acc_sel[124]) );
  OR2X1_HVT U563 ( .A1(n129), .A2(n156), .Y(n178) );
  NAND2X0_HVT U564 ( .A1(data_flash[168]), .A2(n301), .Y(n130) );
  NAND2X0_HVT U565 ( .A1(account[40]), .A2(n287), .Y(n131) );
  NAND2X0_HVT U566 ( .A1(n130), .A2(n131), .Y(out_flash_or_acc_sel[40]) );
  NAND2X0_HVT U567 ( .A1(n217), .A2(match_add[2]), .Y(n132) );
  NAND2X0_HVT U568 ( .A1(write_add[2]), .A2(n245), .Y(n133) );
  NAND2X0_HVT U569 ( .A1(n133), .A2(n132), .Y(add_flash[2]) );
  NAND2X0_HVT U570 ( .A1(account[125]), .A2(n293), .Y(n135) );
  NAND2X0_HVT U571 ( .A1(n134), .A2(n135), .Y(out_flash_or_acc_sel[125]) );
  INVX0_HVT U572 ( .A(n136), .Y(n222) );
  INVX0_HVT U573 ( .A(n14), .Y(n300) );
  IBUFFX2_HVT U574 ( .A(n246), .Y(n267) );
  IBUFFX2_HVT U575 ( .A(n120), .Y(n203) );
  IBUFFX2_HVT U576 ( .A(n274), .Y(n271) );
  NAND2X0_HVT U577 ( .A1(data_flash[237]), .A2(n303), .Y(n139) );
  NAND2X0_HVT U578 ( .A1(account[109]), .A2(n287), .Y(n140) );
  NAND2X0_HVT U579 ( .A1(n139), .A2(n140), .Y(out_flash_or_acc_sel[109]) );
  IBUFFX2_HVT U580 ( .A(n246), .Y(n266) );
  NAND2X0_HVT U581 ( .A1(data_flash[205]), .A2(n294), .Y(n141) );
  NAND2X0_HVT U582 ( .A1(account[77]), .A2(n155), .Y(n142) );
  NAND2X0_HVT U583 ( .A1(n141), .A2(n142), .Y(out_flash_or_acc_sel[77]) );
  NAND2X0_HVT U584 ( .A1(data_flash[248]), .A2(n299), .Y(n143) );
  NAND2X0_HVT U585 ( .A1(account[120]), .A2(n286), .Y(n144) );
  NAND2X0_HVT U586 ( .A1(n143), .A2(n144), .Y(out_flash_or_acc_sel[120]) );
  NAND2X0_HVT U587 ( .A1(data_flash[147]), .A2(n156), .Y(n145) );
  NAND2X0_HVT U588 ( .A1(account[19]), .A2(n293), .Y(n146) );
  NAND2X0_HVT U589 ( .A1(n145), .A2(n146), .Y(out_flash_or_acc_sel[19]) );
  OAI22X1_HVT U590 ( .A1(n149), .A2(n282), .A3(n150), .A4(n191), .Y(
        out_new_old_pass_sel[3]) );
  NAND2X0_HVT U591 ( .A1(data_flash[238]), .A2(n221), .Y(n151) );
  NAND2X0_HVT U592 ( .A1(account[110]), .A2(n287), .Y(n152) );
  NAND2X0_HVT U593 ( .A1(n151), .A2(n152), .Y(out_flash_or_acc_sel[110]) );
  NAND2X0_HVT U594 ( .A1(data_flash[218]), .A2(n297), .Y(n153) );
  NAND2X0_HVT U595 ( .A1(account[90]), .A2(n287), .Y(n154) );
  NAND2X0_HVT U596 ( .A1(n153), .A2(n154), .Y(out_flash_or_acc_sel[90]) );
  NBUFFX2_HVT U597 ( .A(n292), .Y(n155) );
  INVX0_HVT U598 ( .A(data_flash[165]), .Y(n157) );
  NBUFFX2_HVT U599 ( .A(n300), .Y(n156) );
  OAI22X1_HVT U600 ( .A1(n157), .A2(n176), .A3(n158), .A4(n221), .Y(
        out_flash_or_acc_sel[37]) );
  INVX0_HVT U601 ( .A(n52), .Y(n176) );
  INVX0_HVT U602 ( .A(n264), .Y(n159) );
  INVX0_HVT U603 ( .A(n264), .Y(n160) );
  INVX0_HVT U604 ( .A(n265), .Y(n161) );
  INVX0_HVT U605 ( .A(n265), .Y(n162) );
  IBUFFX2_HVT U606 ( .A(n172), .Y(n265) );
  INVX0_HVT U607 ( .A(n265), .Y(n261) );
  INVX0_HVT U608 ( .A(n186), .Y(n163) );
  INVX0_HVT U609 ( .A(n186), .Y(n164) );
  INVX0_HVT U610 ( .A(n186), .Y(n257) );
  INVX0_HVT U611 ( .A(n264), .Y(n256) );
  INVX0_HVT U612 ( .A(n264), .Y(n255) );
  NAND2X0_HVT U613 ( .A1(data_flash[149]), .A2(n156), .Y(n165) );
  NAND2X0_HVT U614 ( .A1(n165), .A2(n166), .Y(out_flash_or_acc_sel[21]) );
  NAND2X0_HVT U615 ( .A1(n36), .A2(data_flash[139]), .Y(n169) );
  NAND2X0_HVT U616 ( .A1(account[11]), .A2(n287), .Y(n170) );
  NAND2X0_HVT U617 ( .A1(n169), .A2(n170), .Y(out_flash_or_acc_sel[11]) );
  INVX0_HVT U618 ( .A(n185), .Y(n253) );
  INVX0_HVT U619 ( .A(n185), .Y(n260) );
  IBUFFX2_HVT U620 ( .A(n185), .Y(n263) );
  INVX0_HVT U621 ( .A(local_master_sel), .Y(n171) );
  INVX0_HVT U622 ( .A(n171), .Y(n172) );
  NAND2X0_HVT U623 ( .A1(data_flash[242]), .A2(n25), .Y(n173) );
  NAND2X0_HVT U624 ( .A1(account[114]), .A2(n287), .Y(n174) );
  NAND2X0_HVT U625 ( .A1(n173), .A2(n174), .Y(out_flash_or_acc_sel[114]) );
  AO22X1_HVT U626 ( .A1(n294), .A2(data_flash[183]), .A3(account[55]), .A4(
        n176), .Y(n175) );
  NAND2X0_HVT U627 ( .A1(data_flash[193]), .A2(n298), .Y(n177) );
  NAND2X0_HVT U628 ( .A1(n177), .A2(n178), .Y(out_flash_or_acc_sel[65]) );
  NAND2X0_HVT U629 ( .A1(data_flash[169]), .A2(n251), .Y(n179) );
  NAND2X0_HVT U630 ( .A1(n179), .A2(n180), .Y(out_flash_or_acc_sel[41]) );
  OAI22X1_HVT U631 ( .A1(n181), .A2(n282), .A3(n182), .A4(n191), .Y(
        out_new_old_pass_sel[51]) );
  IBUFFX2_HVT U632 ( .A(n275), .Y(n268) );
  OA22X2_HVT U633 ( .A1(n234), .A2(n77), .A3(n235), .A4(n266), .Y(n233) );
  INVX0_HVT U634 ( .A(n172), .Y(n185) );
  INVX0_HVT U635 ( .A(n264), .Y(n258) );
  NAND2X0_HVT U636 ( .A1(data_flash[202]), .A2(n12), .Y(n187) );
  NAND2X0_HVT U637 ( .A1(account[74]), .A2(n292), .Y(n188) );
  NAND2X0_HVT U638 ( .A1(n187), .A2(n188), .Y(out_flash_or_acc_sel[74]) );
  OAI22X1_HVT U639 ( .A1(n189), .A2(n277), .A3(n190), .A4(n191), .Y(
        out_new_old_pass_sel[47]) );
  OA22X1_HVT U640 ( .A1(n194), .A2(n209), .A3(n195), .A4(n196), .Y(n193) );
  OAI22X1_HVT U641 ( .A1(n200), .A2(n276), .A3(n201), .A4(n148), .Y(
        out_new_old_pass_sel[4]) );
  INVX0_HVT U642 ( .A(n147), .Y(n275) );
  INVX0_HVT U643 ( .A(n285), .Y(n225) );
  NAND2X0_HVT U644 ( .A1(data_flash[130]), .A2(n299), .Y(n204) );
  NAND2X0_HVT U645 ( .A1(account[2]), .A2(n291), .Y(n205) );
  NAND2X0_HVT U646 ( .A1(n204), .A2(n205), .Y(out_flash_or_acc_sel[2]) );
  INVX0_HVT U647 ( .A(n211), .Y(out_new_old_pass_sel[45]) );
  NAND2X0_HVT U648 ( .A1(data_flash[201]), .A2(n222), .Y(n206) );
  NAND2X0_HVT U649 ( .A1(account[73]), .A2(n292), .Y(n207) );
  NAND2X0_HVT U650 ( .A1(n206), .A2(n207), .Y(out_flash_or_acc_sel[73]) );
  NBUFFX2_HVT U651 ( .A(n279), .Y(n208) );
  OA22X1_HVT U652 ( .A1(n212), .A2(n42), .A3(n213), .A4(n147), .Y(n211) );
  NAND2X0_HVT U653 ( .A1(out_decry[0]), .A2(n210), .Y(n214) );
  NAND2X0_HVT U654 ( .A1(pass[0]), .A2(n284), .Y(n215) );
  NAND2X0_HVT U655 ( .A1(n214), .A2(n215), .Y(out_new_old_pass_sel[0]) );
  IBUFFX2_HVT U656 ( .A(n275), .Y(n236) );
  IBUFFX2_HVT U657 ( .A(n275), .Y(n237) );
  INVX0_HVT U658 ( .A(n233), .Y(out_new_old_pass_sel[7]) );
  INVX0_HVT U659 ( .A(n250), .Y(n249) );
  NAND2X0_HVT U660 ( .A1(data_flash[206]), .A2(n299), .Y(n218) );
  NAND2X0_HVT U661 ( .A1(account[78]), .A2(n292), .Y(n219) );
  NAND2X0_HVT U662 ( .A1(n218), .A2(n219), .Y(out_flash_or_acc_sel[78]) );
  IBUFFX2_HVT U663 ( .A(n67), .Y(n270) );
  IBUFFX2_HVT U664 ( .A(n67), .Y(n273) );
  IBUFFX2_HVT U665 ( .A(n67), .Y(n238) );
  IBUFFX2_HVT U666 ( .A(n274), .Y(n239) );
  INVX0_HVT U667 ( .A(flash_or_acc_sel), .Y(n285) );
  NAND2X0_HVT U668 ( .A1(data_flash[137]), .A2(n251), .Y(n229) );
  NAND2X0_HVT U669 ( .A1(n293), .A2(account[9]), .Y(n230) );
  NAND2X0_HVT U670 ( .A1(n229), .A2(n230), .Y(out_flash_or_acc_sel[9]) );
  NAND2X0_HVT U671 ( .A1(data_flash[221]), .A2(n52), .Y(n231) );
  NAND2X0_HVT U672 ( .A1(account[93]), .A2(n293), .Y(n232) );
  NAND2X0_HVT U673 ( .A1(n231), .A2(n232), .Y(out_flash_or_acc_sel[93]) );
  INVX0_HVT U674 ( .A(data_flash[233]), .Y(n240) );
  INVX0_HVT U675 ( .A(data_flash[129]), .Y(n242) );
  OAI22X1_HVT U676 ( .A1(n136), .A2(n240), .A3(n241), .A4(n302), .Y(
        out_flash_or_acc_sel[105]) );
  OAI22X1_HVT U677 ( .A1(n293), .A2(n242), .A3(n243), .A4(n25), .Y(
        out_flash_or_acc_sel[1]) );
  IBUFFX2_HVT U678 ( .A(n67), .Y(n272) );
  NAND2X0_HVT U679 ( .A1(data_flash[219]), .A2(n222), .Y(n247) );
  NAND2X0_HVT U680 ( .A1(account[91]), .A2(n287), .Y(n248) );
  NAND2X0_HVT U681 ( .A1(n247), .A2(n248), .Y(out_flash_or_acc_sel[91]) );
  NBUFFX2_HVT U682 ( .A(n306), .Y(n250) );
  INVX0_HVT U683 ( .A(n138), .Y(n283) );
  INVX1_HVT U684 ( .A(n186), .Y(n259) );
  INVX1_HVT U685 ( .A(n265), .Y(n254) );
  INVX1_HVT U686 ( .A(n305), .Y(n304) );
  INVX1_HVT U687 ( .A(rst), .Y(n305) );
  INVX0_HVT U688 ( .A(boot_lood), .Y(n306) );
endmodule

