
module inv_shift_rows ( in, out );
  input [127:0] in;
  output [127:0] out;

  assign out[127] = in[127];
  assign out[126] = in[126];
  assign out[125] = in[125];
  assign out[124] = in[124];
  assign out[123] = in[123];
  assign out[122] = in[122];
  assign out[121] = in[121];
  assign out[120] = in[120];
  assign out[119] = in[23];
  assign out[118] = in[22];
  assign out[117] = in[21];
  assign out[116] = in[20];
  assign out[115] = in[19];
  assign out[114] = in[18];
  assign out[113] = in[17];
  assign out[112] = in[16];
  assign out[111] = in[47];
  assign out[110] = in[46];
  assign out[109] = in[45];
  assign out[108] = in[44];
  assign out[107] = in[43];
  assign out[106] = in[42];
  assign out[105] = in[41];
  assign out[104] = in[40];
  assign out[103] = in[71];
  assign out[102] = in[70];
  assign out[101] = in[69];
  assign out[100] = in[68];
  assign out[99] = in[67];
  assign out[98] = in[66];
  assign out[97] = in[65];
  assign out[96] = in[64];
  assign out[95] = in[95];
  assign out[94] = in[94];
  assign out[93] = in[93];
  assign out[92] = in[92];
  assign out[91] = in[91];
  assign out[90] = in[90];
  assign out[89] = in[89];
  assign out[88] = in[88];
  assign out[87] = in[119];
  assign out[86] = in[118];
  assign out[85] = in[117];
  assign out[84] = in[116];
  assign out[83] = in[115];
  assign out[82] = in[114];
  assign out[81] = in[113];
  assign out[80] = in[112];
  assign out[79] = in[15];
  assign out[78] = in[14];
  assign out[77] = in[13];
  assign out[76] = in[12];
  assign out[75] = in[11];
  assign out[74] = in[10];
  assign out[73] = in[9];
  assign out[72] = in[8];
  assign out[71] = in[39];
  assign out[70] = in[38];
  assign out[69] = in[37];
  assign out[68] = in[36];
  assign out[67] = in[35];
  assign out[66] = in[34];
  assign out[65] = in[33];
  assign out[64] = in[32];
  assign out[63] = in[63];
  assign out[62] = in[62];
  assign out[61] = in[61];
  assign out[60] = in[60];
  assign out[59] = in[59];
  assign out[58] = in[58];
  assign out[57] = in[57];
  assign out[56] = in[56];
  assign out[55] = in[87];
  assign out[54] = in[86];
  assign out[53] = in[85];
  assign out[52] = in[84];
  assign out[51] = in[83];
  assign out[50] = in[82];
  assign out[49] = in[81];
  assign out[48] = in[80];
  assign out[47] = in[111];
  assign out[46] = in[110];
  assign out[45] = in[109];
  assign out[44] = in[108];
  assign out[43] = in[107];
  assign out[42] = in[106];
  assign out[41] = in[105];
  assign out[40] = in[104];
  assign out[39] = in[7];
  assign out[38] = in[6];
  assign out[37] = in[5];
  assign out[36] = in[4];
  assign out[35] = in[3];
  assign out[34] = in[2];
  assign out[33] = in[1];
  assign out[32] = in[0];
  assign out[31] = in[31];
  assign out[30] = in[30];
  assign out[29] = in[29];
  assign out[28] = in[28];
  assign out[27] = in[27];
  assign out[26] = in[26];
  assign out[25] = in[25];
  assign out[24] = in[24];
  assign out[23] = in[55];
  assign out[22] = in[54];
  assign out[21] = in[53];
  assign out[20] = in[52];
  assign out[19] = in[51];
  assign out[18] = in[50];
  assign out[17] = in[49];
  assign out[16] = in[48];
  assign out[15] = in[79];
  assign out[14] = in[78];
  assign out[13] = in[77];
  assign out[12] = in[76];
  assign out[11] = in[75];
  assign out[10] = in[74];
  assign out[9] = in[73];
  assign out[8] = in[72];
  assign out[7] = in[103];
  assign out[6] = in[102];
  assign out[5] = in[101];
  assign out[4] = in[100];
  assign out[3] = in[99];
  assign out[2] = in[98];
  assign out[1] = in[97];
  assign out[0] = in[96];

endmodule

