
module keygen ( round_num, keyin, keyout );
  input [0:3] round_num;
  input [0:127] keyin;
  output [0:127] keyout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479;

  XNOR3X1_HVT U1 ( .A1(n1), .A2(keyin[67]), .A3(keyout[35]), .Y(keyout[99]) );
  XNOR2X1_HVT U2 ( .A1(keyout[66]), .A2(n2), .Y(keyout[98]) );
  XOR2X1_HVT U3 ( .A1(keyin[97]), .A2(keyout[65]), .Y(keyout[97]) );
  XNOR2X1_HVT U4 ( .A1(n3), .A2(keyout[64]), .Y(keyout[96]) );
  INVX0_HVT U5 ( .A(n4), .Y(keyout[83]) );
  INVX0_HVT U6 ( .A(n5), .Y(keyout[75]) );
  XOR2X1_HVT U7 ( .A1(keyout[38]), .A2(keyin[70]), .Y(keyout[70]) );
  XNOR2X1_HVT U8 ( .A1(n6), .A2(n7), .Y(keyout[6]) );
  XOR2X1_HVT U9 ( .A1(keyin[69]), .A2(keyout[37]), .Y(keyout[69]) );
  XNOR2X1_HVT U10 ( .A1(keyin[67]), .A2(n8), .Y(keyout[67]) );
  XOR2X1_HVT U11 ( .A1(keyout[34]), .A2(keyin[66]), .Y(keyout[66]) );
  XOR3X1_HVT U12 ( .A1(n9), .A2(n10), .A3(n11), .Y(keyout[65]) );
  XOR2X1_HVT U13 ( .A1(keyin[65]), .A2(keyin[33]), .Y(n10) );
  XOR3X1_HVT U14 ( .A1(n12), .A2(n13), .A3(n14), .Y(keyout[64]) );
  XOR2X1_HVT U15 ( .A1(keyin[64]), .A2(keyin[32]), .Y(n13) );
  XOR2X1_HVT U16 ( .A1(keyin[63]), .A2(keyout[31]), .Y(keyout[63]) );
  XOR2X1_HVT U17 ( .A1(keyout[30]), .A2(keyin[62]), .Y(keyout[62]) );
  XOR2X1_HVT U18 ( .A1(keyin[61]), .A2(keyout[29]), .Y(keyout[61]) );
  XOR2X1_HVT U19 ( .A1(keyin[60]), .A2(keyout[28]), .Y(keyout[60]) );
  XNOR2X1_HVT U20 ( .A1(n15), .A2(n16), .Y(keyout[5]) );
  XOR2X1_HVT U21 ( .A1(keyout[27]), .A2(keyin[59]), .Y(keyout[59]) );
  XOR2X1_HVT U22 ( .A1(keyin[58]), .A2(keyout[26]), .Y(keyout[58]) );
  XOR2X1_HVT U23 ( .A1(keyout[25]), .A2(keyin[57]), .Y(keyout[57]) );
  XOR2X1_HVT U24 ( .A1(keyout[24]), .A2(keyin[56]), .Y(keyout[56]) );
  XNOR2X1_HVT U25 ( .A1(keyin[55]), .A2(n17), .Y(keyout[55]) );
  XOR2X1_HVT U26 ( .A1(keyin[54]), .A2(keyout[22]), .Y(keyout[54]) );
  XOR2X1_HVT U27 ( .A1(keyout[21]), .A2(keyin[53]), .Y(keyout[53]) );
  XOR2X1_HVT U28 ( .A1(keyout[20]), .A2(keyin[52]), .Y(keyout[52]) );
  XOR2X1_HVT U29 ( .A1(keyin[51]), .A2(keyout[19]), .Y(keyout[51]) );
  XOR2X1_HVT U30 ( .A1(keyin[50]), .A2(keyout[18]), .Y(keyout[50]) );
  XNOR2X1_HVT U31 ( .A1(n18), .A2(n19), .Y(keyout[4]) );
  XOR2X1_HVT U32 ( .A1(keyin[49]), .A2(keyout[17]), .Y(keyout[49]) );
  XOR2X1_HVT U33 ( .A1(keyin[48]), .A2(keyout[16]), .Y(keyout[48]) );
  XNOR2X1_HVT U34 ( .A1(keyin[47]), .A2(n20), .Y(keyout[47]) );
  XOR2X1_HVT U35 ( .A1(keyin[46]), .A2(keyout[14]), .Y(keyout[46]) );
  XOR2X1_HVT U36 ( .A1(keyout[13]), .A2(keyin[45]), .Y(keyout[45]) );
  XOR2X1_HVT U37 ( .A1(keyout[12]), .A2(keyin[44]), .Y(keyout[44]) );
  XOR2X1_HVT U38 ( .A1(keyin[43]), .A2(keyout[11]), .Y(keyout[43]) );
  XOR2X1_HVT U39 ( .A1(keyin[42]), .A2(keyout[10]), .Y(keyout[42]) );
  XOR2X1_HVT U40 ( .A1(keyin[41]), .A2(keyout[9]), .Y(keyout[41]) );
  XOR2X1_HVT U41 ( .A1(keyin[40]), .A2(keyout[8]), .Y(keyout[40]) );
  XOR2X1_HVT U42 ( .A1(n21), .A2(n22), .Y(keyout[3]) );
  INVX0_HVT U43 ( .A(n8), .Y(keyout[35]) );
  XNOR3X1_HVT U44 ( .A1(n21), .A2(keyin[35]), .A3(n22), .Y(n8) );
  XOR2X1_HVT U45 ( .A1(n23), .A2(keyin[3]), .Y(n22) );
  MUX21X1_HVT U46 ( .A1(n24), .A2(n25), .S0(n26), .Y(n23) );
  AO221X1_HVT U47 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .A5(n31), .Y(n25)
         );
  AO22X1_HVT U48 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .Y(n31) );
  AO222X1_HVT U49 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .A5(n40), .A6(n41), 
        .Y(n35) );
  NAND2X0_HVT U50 ( .A1(n42), .A2(n43), .Y(n38) );
  NAND3X0_HVT U51 ( .A1(keyin[106]), .A2(n44), .A3(n45), .Y(n43) );
  AO221X1_HVT U52 ( .A1(n46), .A2(n47), .A3(n48), .A4(n36), .A5(n49), .Y(n33)
         );
  AO22X1_HVT U53 ( .A1(n50), .A2(n40), .A3(n51), .A4(n52), .Y(n49) );
  AO222X1_HVT U54 ( .A1(n46), .A2(n53), .A3(n54), .A4(n55), .A5(n52), .A6(n56), 
        .Y(n30) );
  AO221X1_HVT U55 ( .A1(n57), .A2(n46), .A3(n36), .A4(n58), .A5(n59), .Y(n28)
         );
  AO22X1_HVT U56 ( .A1(n60), .A2(n40), .A3(n48), .A4(n52), .Y(n59) );
  AND2X1_HVT U57 ( .A1(n61), .A2(n62), .Y(n48) );
  AND2X1_HVT U58 ( .A1(n37), .A2(n63), .Y(n57) );
  AO221X1_HVT U59 ( .A1(n36), .A2(n64), .A3(n40), .A4(n65), .A5(n66), .Y(n24)
         );
  AO221X1_HVT U60 ( .A1(n52), .A2(n67), .A3(n46), .A4(n68), .A5(n69), .Y(n66)
         );
  AND3X1_HVT U61 ( .A1(n70), .A2(n27), .A3(keyin[106]), .Y(n69) );
  AO222X1_HVT U62 ( .A1(n29), .A2(n71), .A3(n72), .A4(n34), .A5(n32), .A6(n73), 
        .Y(n68) );
  INVX0_HVT U63 ( .A(n74), .Y(n71) );
  AO22X1_HVT U64 ( .A1(n34), .A2(n75), .A3(n76), .A4(n77), .Y(n67) );
  AO21X1_HVT U65 ( .A1(n32), .A2(n44), .A3(n29), .Y(n76) );
  INVX0_HVT U66 ( .A(n78), .Y(n75) );
  AO221X1_HVT U67 ( .A1(n34), .A2(n77), .A3(n29), .A4(n79), .A5(n80), .Y(n65)
         );
  AO22X1_HVT U68 ( .A1(n27), .A2(n81), .A3(n82), .A4(n32), .Y(n80) );
  INVX0_HVT U69 ( .A(n62), .Y(n82) );
  AO221X1_HVT U70 ( .A1(n83), .A2(n32), .A3(n84), .A4(n27), .A5(n85), .Y(n64)
         );
  AO22X1_HVT U71 ( .A1(n86), .A2(n29), .A3(n87), .A4(n34), .Y(n85) );
  NAND2X0_HVT U72 ( .A1(n88), .A2(n89), .Y(n21) );
  MUX21X1_HVT U73 ( .A1(n90), .A2(n91), .S0(n92), .Y(n88) );
  NAND3X0_HVT U74 ( .A1(round_num[3]), .A2(n93), .A3(round_num[1]), .Y(n91) );
  XNOR3X1_HVT U75 ( .A1(n94), .A2(keyin[34]), .A3(n95), .Y(keyout[34]) );
  XOR2X1_HVT U76 ( .A1(keyin[33]), .A2(keyout[1]), .Y(keyout[33]) );
  XOR2X1_HVT U77 ( .A1(keyin[32]), .A2(keyout[0]), .Y(keyout[32]) );
  XNOR2X1_HVT U78 ( .A1(n95), .A2(n94), .Y(keyout[2]) );
  AO21X1_HVT U79 ( .A1(n96), .A2(round_num[2]), .A3(n97), .Y(n94) );
  XNOR2X1_HVT U80 ( .A1(keyin[2]), .A2(n98), .Y(n95) );
  MUX21X1_HVT U81 ( .A1(n99), .A2(n100), .S0(n26), .Y(n98) );
  AO221X1_HVT U82 ( .A1(n32), .A2(n101), .A3(n27), .A4(n102), .A5(n103), .Y(
        n100) );
  AO22X1_HVT U83 ( .A1(n34), .A2(n104), .A3(n29), .A4(n105), .Y(n103) );
  OAI221X1_HVT U84 ( .A1(n106), .A2(n81), .A3(n107), .A4(n108), .A5(n109), .Y(
        n105) );
  MUX21X1_HVT U85 ( .A1(n110), .A2(n111), .S0(n112), .Y(n109) );
  NAND2X0_HVT U86 ( .A1(keyin[106]), .A2(n63), .Y(n111) );
  NAND2X0_HVT U87 ( .A1(keyin[108]), .A2(n52), .Y(n110) );
  AO222X1_HVT U88 ( .A1(n113), .A2(n39), .A3(n52), .A4(n114), .A5(n46), .A6(
        n77), .Y(n104) );
  NAND2X0_HVT U89 ( .A1(n115), .A2(n116), .Y(n114) );
  OAI21X1_HVT U90 ( .A1(n117), .A2(keyin[106]), .A3(n108), .Y(n113) );
  AO221X1_HVT U91 ( .A1(n36), .A2(n118), .A3(n119), .A4(n52), .A5(n120), .Y(
        n102) );
  AO22X1_HVT U92 ( .A1(n46), .A2(n121), .A3(n40), .A4(n122), .Y(n120) );
  AO221X1_HVT U93 ( .A1(n52), .A2(n123), .A3(n124), .A4(n46), .A5(n125), .Y(
        n101) );
  AO22X1_HVT U94 ( .A1(n126), .A2(n40), .A3(n36), .A4(n77), .Y(n125) );
  INVX0_HVT U95 ( .A(n127), .Y(n124) );
  NAND2X0_HVT U96 ( .A1(n45), .A2(n44), .Y(n123) );
  AO221X1_HVT U97 ( .A1(n29), .A2(n128), .A3(n32), .A4(n129), .A5(n130), .Y(
        n99) );
  AO22X1_HVT U98 ( .A1(n27), .A2(n131), .A3(n34), .A4(n132), .Y(n130) );
  AO221X1_HVT U99 ( .A1(n133), .A2(n37), .A3(n36), .A4(n41), .A5(n134), .Y(
        n132) );
  AO22X1_HVT U100 ( .A1(n40), .A2(n135), .A3(n52), .A4(n136), .Y(n134) );
  NAND2X0_HVT U101 ( .A1(n137), .A2(n138), .Y(n136) );
  NAND2X0_HVT U102 ( .A1(n139), .A2(n140), .Y(n135) );
  AO222X1_HVT U103 ( .A1(n36), .A2(n141), .A3(n142), .A4(n143), .A5(n40), .A6(
        n63), .Y(n131) );
  AO21X1_HVT U104 ( .A1(keyin[106]), .A2(n144), .A3(n46), .Y(n142) );
  NAND2X0_HVT U105 ( .A1(n145), .A2(n139), .Y(n144) );
  AO221X1_HVT U106 ( .A1(n146), .A2(n52), .A3(n147), .A4(n40), .A5(n148), .Y(
        n129) );
  AO22X1_HVT U107 ( .A1(n36), .A2(n149), .A3(n150), .A4(n46), .Y(n148) );
  INVX0_HVT U108 ( .A(n151), .Y(n146) );
  AO221X1_HVT U109 ( .A1(n152), .A2(n46), .A3(n153), .A4(n36), .A5(n154), .Y(
        n128) );
  AO22X1_HVT U110 ( .A1(n155), .A2(n40), .A3(n86), .A4(n52), .Y(n154) );
  INVX0_HVT U111 ( .A(n17), .Y(keyout[23]) );
  XOR2X1_HVT U112 ( .A1(n11), .A2(n9), .Y(keyout[1]) );
  NAND2X0_HVT U113 ( .A1(n156), .A2(round_num[1]), .Y(n9) );
  XNOR2X1_HVT U114 ( .A1(keyin[1]), .A2(n157), .Y(n11) );
  MUX21X1_HVT U115 ( .A1(n158), .A2(n159), .S0(n26), .Y(n157) );
  AO221X1_HVT U116 ( .A1(n34), .A2(n160), .A3(n32), .A4(n161), .A5(n162), .Y(
        n159) );
  OAI22X1_HVT U117 ( .A1(n163), .A2(n164), .A3(n165), .A4(n166), .Y(n162) );
  OA221X1_HVT U118 ( .A1(n167), .A2(n168), .A3(n169), .A4(n108), .A5(n170), 
        .Y(n165) );
  OA22X1_HVT U119 ( .A1(n106), .A2(n171), .A3(n42), .A4(n172), .Y(n170) );
  NAND2X0_HVT U120 ( .A1(n87), .A2(n115), .Y(n171) );
  OA221X1_HVT U121 ( .A1(n167), .A2(n173), .A3(n108), .A4(n54), .A5(n174), .Y(
        n163) );
  AOI22X1_HVT U122 ( .A1(n175), .A2(n46), .A3(n176), .A4(n40), .Y(n174) );
  NAND2X0_HVT U123 ( .A1(n177), .A2(n178), .Y(n54) );
  AO221X1_HVT U124 ( .A1(n52), .A2(n37), .A3(n40), .A4(n179), .A5(n180), .Y(
        n161) );
  AO22X1_HVT U125 ( .A1(n181), .A2(n46), .A3(n36), .A4(n182), .Y(n180) );
  NAND2X0_HVT U126 ( .A1(n37), .A2(n145), .Y(n182) );
  AO221X1_HVT U127 ( .A1(n36), .A2(n183), .A3(n46), .A4(n184), .A5(n185), .Y(
        n160) );
  AO22X1_HVT U128 ( .A1(n186), .A2(n40), .A3(n52), .A4(n41), .Y(n185) );
  NAND2X0_HVT U129 ( .A1(n177), .A2(n187), .Y(n183) );
  AO221X1_HVT U130 ( .A1(n29), .A2(n188), .A3(n27), .A4(n189), .A5(n190), .Y(
        n158) );
  AO22X1_HVT U131 ( .A1(n34), .A2(n191), .A3(n32), .A4(n192), .Y(n190) );
  AO222X1_HVT U132 ( .A1(n60), .A2(n46), .A3(n83), .A4(n193), .A5(n52), .A6(
        n178), .Y(n192) );
  AO21X1_HVT U133 ( .A1(n194), .A2(n55), .A3(n36), .Y(n193) );
  INVX0_HVT U134 ( .A(n184), .Y(n60) );
  NAND2X0_HVT U135 ( .A1(n195), .A2(n196), .Y(n184) );
  AO221X1_HVT U136 ( .A1(n36), .A2(n138), .A3(n197), .A4(n46), .A5(n198), .Y(
        n191) );
  OAI22X1_HVT U137 ( .A1(n106), .A2(n199), .A3(n200), .A4(n167), .Y(n198) );
  INVX0_HVT U138 ( .A(n201), .Y(n197) );
  AO221X1_HVT U139 ( .A1(n36), .A2(n202), .A3(n203), .A4(n40), .A5(n204), .Y(
        n189) );
  AO22X1_HVT U140 ( .A1(n46), .A2(n205), .A3(n52), .A4(n206), .Y(n204) );
  NAND2X0_HVT U141 ( .A1(n53), .A2(n139), .Y(n206) );
  AO221X1_HVT U142 ( .A1(n52), .A2(n179), .A3(n40), .A4(n121), .A5(n207), .Y(
        n188) );
  AO21X1_HVT U143 ( .A1(n208), .A2(n209), .A3(n210), .Y(n207) );
  INVX0_HVT U144 ( .A(n20), .Y(keyout[15]) );
  XNOR2X1_HVT U145 ( .A1(n211), .A2(keyout[95]), .Y(keyout[127]) );
  XOR3X1_HVT U146 ( .A1(keyin[63]), .A2(keyin[95]), .A3(keyout[31]), .Y(
        keyout[95]) );
  XOR2X1_HVT U147 ( .A1(keyin[31]), .A2(n212), .Y(keyout[31]) );
  MUX41X1_HVT U148 ( .A1(n213), .A3(n214), .A2(n215), .A4(n216), .S0(n217), 
        .S1(keyin[97]), .Y(n212) );
  MUX21X1_HVT U149 ( .A1(n218), .A2(n219), .S0(n2), .Y(n216) );
  NAND4X0_HVT U150 ( .A1(n220), .A2(n221), .A3(n222), .A4(n223), .Y(n219) );
  OA22X1_HVT U151 ( .A1(n224), .A2(n225), .A3(n226), .A4(n227), .Y(n223) );
  NAND2X0_HVT U152 ( .A1(n228), .A2(n229), .Y(n222) );
  AO221X1_HVT U153 ( .A1(n229), .A2(n230), .A3(n231), .A4(n232), .A5(n233), 
        .Y(n218) );
  AO22X1_HVT U154 ( .A1(n234), .A2(n235), .A3(n236), .A4(n237), .Y(n233) );
  NAND2X0_HVT U155 ( .A1(n238), .A2(n239), .Y(n232) );
  NAND2X0_HVT U156 ( .A1(n240), .A2(n241), .Y(n230) );
  MUX21X1_HVT U157 ( .A1(n242), .A2(n243), .S0(n2), .Y(n215) );
  AO221X1_HVT U158 ( .A1(n244), .A2(n229), .A3(n235), .A4(keyin[100]), .A5(
        n245), .Y(n243) );
  AO21X1_HVT U159 ( .A1(n237), .A2(n246), .A3(n247), .Y(n245) );
  AO221X1_HVT U160 ( .A1(n237), .A2(n248), .A3(n229), .A4(n225), .A5(n249), 
        .Y(n242) );
  AO22X1_HVT U161 ( .A1(n235), .A2(n250), .A3(n231), .A4(n251), .Y(n249) );
  NAND2X0_HVT U162 ( .A1(n252), .A2(n253), .Y(n225) );
  AO221X1_HVT U163 ( .A1(n254), .A2(n231), .A3(n255), .A4(n237), .A5(n256), 
        .Y(n214) );
  AO21X1_HVT U164 ( .A1(n257), .A2(n229), .A3(n258), .Y(n256) );
  MUX21X1_HVT U165 ( .A1(n259), .A2(n260), .S0(n2), .Y(n258) );
  OAI22X1_HVT U166 ( .A1(n261), .A2(n227), .A3(n262), .A4(n224), .Y(n260) );
  OAI222X1_HVT U167 ( .A1(n224), .A2(keyin[102]), .A3(n263), .A4(n264), .A5(
        n265), .A6(n227), .Y(n259) );
  INVX0_HVT U168 ( .A(n266), .Y(n254) );
  MUX21X1_HVT U169 ( .A1(n267), .A2(n268), .S0(n2), .Y(n213) );
  AO221X1_HVT U170 ( .A1(n269), .A2(n270), .A3(n237), .A4(n253), .A5(n271), 
        .Y(n268) );
  AO22X1_HVT U171 ( .A1(n272), .A2(n231), .A3(n273), .A4(n229), .Y(n271) );
  INVX0_HVT U172 ( .A(n274), .Y(n272) );
  AND2X1_HVT U173 ( .A1(n235), .A2(n275), .Y(n269) );
  AO221X1_HVT U174 ( .A1(n276), .A2(n237), .A3(n277), .A4(n229), .A5(n278), 
        .Y(n267) );
  AO22X1_HVT U175 ( .A1(n279), .A2(n235), .A3(n270), .A4(n231), .Y(n278) );
  XNOR2X1_HVT U176 ( .A1(keyout[94]), .A2(n280), .Y(keyout[126]) );
  XOR3X1_HVT U177 ( .A1(keyin[62]), .A2(keyin[94]), .A3(keyout[30]), .Y(
        keyout[94]) );
  MUX21X1_HVT U178 ( .A1(n281), .A2(n282), .S0(keyin[97]), .Y(keyout[30]) );
  XOR2X1_HVT U179 ( .A1(n283), .A2(keyin[30]), .Y(n282) );
  AO221X1_HVT U180 ( .A1(n284), .A2(n285), .A3(n286), .A4(n287), .A5(n288), 
        .Y(n283) );
  AO22X1_HVT U181 ( .A1(n289), .A2(n290), .A3(n291), .A4(n292), .Y(n288) );
  AO221X1_HVT U182 ( .A1(n293), .A2(n231), .A3(n294), .A4(n235), .A5(n295), 
        .Y(n292) );
  OAI21X1_HVT U183 ( .A1(n296), .A2(n297), .A3(n298), .Y(n295) );
  AO221X1_HVT U184 ( .A1(n229), .A2(n299), .A3(n300), .A4(n231), .A5(n301), 
        .Y(n290) );
  MUX21X1_HVT U185 ( .A1(n237), .A2(n235), .S0(n302), .Y(n301) );
  AO221X1_HVT U186 ( .A1(n303), .A2(n231), .A3(n304), .A4(n235), .A5(n305), 
        .Y(n287) );
  AO22X1_HVT U187 ( .A1(n237), .A2(n261), .A3(n229), .A4(n306), .Y(n305) );
  NAND2X0_HVT U188 ( .A1(n307), .A2(n308), .Y(n306) );
  INVX0_HVT U189 ( .A(n309), .Y(n304) );
  NAND3X0_HVT U190 ( .A1(n310), .A2(n311), .A3(n312), .Y(n285) );
  AOI222X1_HVT U191 ( .A1(n231), .A2(n313), .A3(n237), .A4(n314), .A5(n229), 
        .A6(n315), .Y(n312) );
  NAND2X0_HVT U192 ( .A1(n308), .A2(n316), .Y(n314) );
  NAND2X0_HVT U193 ( .A1(n257), .A2(n235), .Y(n311) );
  INVX0_HVT U194 ( .A(n317), .Y(n257) );
  XNOR2X1_HVT U195 ( .A1(keyin[30]), .A2(n318), .Y(n281) );
  OA221X1_HVT U196 ( .A1(n319), .A2(n320), .A3(n321), .A4(n322), .A5(n323), 
        .Y(n318) );
  OA22X1_HVT U197 ( .A1(n324), .A2(n325), .A3(n326), .A4(n327), .Y(n323) );
  OA221X1_HVT U198 ( .A1(n277), .A2(n227), .A3(n270), .A4(n297), .A5(n328), 
        .Y(n326) );
  OA21X1_HVT U199 ( .A1(n224), .A2(n329), .A3(n330), .Y(n328) );
  OA221X1_HVT U200 ( .A1(n331), .A2(n227), .A3(n251), .A4(n332), .A5(n333), 
        .Y(n324) );
  NAND3X0_HVT U201 ( .A1(n334), .A2(n241), .A3(n335), .Y(n333) );
  AO21X1_HVT U202 ( .A1(n336), .A2(keyin[101]), .A3(n229), .Y(n335) );
  INVX0_HVT U203 ( .A(n337), .Y(n251) );
  OA221X1_HVT U204 ( .A1(n279), .A2(n224), .A3(n297), .A4(n337), .A5(n338), 
        .Y(n321) );
  OA221X1_HVT U205 ( .A1(n227), .A2(n263), .A3(n332), .A4(n339), .A5(n298), 
        .Y(n338) );
  NAND2X0_HVT U206 ( .A1(n275), .A2(n340), .Y(n337) );
  INVX0_HVT U207 ( .A(n341), .Y(n279) );
  OA221X1_HVT U208 ( .A1(n227), .A2(n342), .A3(n332), .A4(n296), .A5(n343), 
        .Y(n319) );
  OA22X1_HVT U209 ( .A1(n224), .A2(n344), .A3(n345), .A4(n297), .Y(n343) );
  INVX0_HVT U210 ( .A(n248), .Y(n345) );
  NAND2X0_HVT U211 ( .A1(n317), .A2(n334), .Y(n344) );
  NAND2X0_HVT U212 ( .A1(n346), .A2(n263), .Y(n296) );
  XNOR2X1_HVT U213 ( .A1(n347), .A2(keyout[93]), .Y(keyout[125]) );
  XOR3X1_HVT U214 ( .A1(keyin[61]), .A2(keyin[93]), .A3(keyout[29]), .Y(
        keyout[93]) );
  XOR2X1_HVT U215 ( .A1(keyin[29]), .A2(n348), .Y(keyout[29]) );
  MUX21X1_HVT U216 ( .A1(n349), .A2(n350), .S0(keyin[97]), .Y(n348) );
  AO221X1_HVT U217 ( .A1(n286), .A2(n351), .A3(n289), .A4(n352), .A5(n353), 
        .Y(n350) );
  AO22X1_HVT U218 ( .A1(n291), .A2(n354), .A3(n284), .A4(n355), .Y(n353) );
  AO221X1_HVT U219 ( .A1(n235), .A2(n309), .A3(n356), .A4(n264), .A5(n357), 
        .Y(n355) );
  MUX21X1_HVT U220 ( .A1(n358), .A2(n359), .S0(n360), .Y(n357) );
  AO22X1_HVT U221 ( .A1(n231), .A2(n1), .A3(n229), .A4(keyin[100]), .Y(n359)
         );
  AND2X1_HVT U222 ( .A1(keyin[101]), .A2(n334), .Y(n358) );
  NAND3X0_HVT U223 ( .A1(n361), .A2(n362), .A3(n363), .Y(n354) );
  OA22X1_HVT U224 ( .A1(n332), .A2(n263), .A3(n227), .A4(n364), .Y(n363) );
  AO21X1_HVT U225 ( .A1(n246), .A2(n365), .A3(n224), .Y(n361) );
  AO221X1_HVT U226 ( .A1(n366), .A2(n231), .A3(n244), .A4(n235), .A5(n367), 
        .Y(n352) );
  AO221X1_HVT U227 ( .A1(n237), .A2(n368), .A3(n229), .A4(n262), .A5(n247), 
        .Y(n367) );
  AND2X1_HVT U228 ( .A1(n253), .A2(n308), .Y(n244) );
  NAND4X0_HVT U229 ( .A1(n369), .A2(n362), .A3(n370), .A4(n298), .Y(n351) );
  NAND2X0_HVT U230 ( .A1(n371), .A2(n229), .Y(n362) );
  AO21X1_HVT U231 ( .A1(n270), .A2(n275), .A3(n224), .Y(n369) );
  AO221X1_HVT U232 ( .A1(n291), .A2(n372), .A3(n286), .A4(n373), .A5(n374), 
        .Y(n349) );
  AO22X1_HVT U233 ( .A1(n284), .A2(n375), .A3(n376), .A4(n289), .Y(n374) );
  MUX21X1_HVT U234 ( .A1(n377), .A2(n273), .S0(n378), .Y(n376) );
  AND2X1_HVT U235 ( .A1(n227), .A2(n297), .Y(n378) );
  MUX21X1_HVT U236 ( .A1(n341), .A2(n379), .S0(n264), .Y(n377) );
  NAND2X0_HVT U237 ( .A1(n241), .A2(n253), .Y(n341) );
  AO221X1_HVT U238 ( .A1(n380), .A2(n229), .A3(n235), .A4(n265), .A5(n381), 
        .Y(n375) );
  AO21X1_HVT U239 ( .A1(n382), .A2(n264), .A3(n383), .Y(n381) );
  AO221X1_HVT U240 ( .A1(n235), .A2(n384), .A3(n385), .A4(n237), .A5(n386), 
        .Y(n373) );
  AO21X1_HVT U241 ( .A1(n229), .A2(n387), .A3(n383), .Y(n386) );
  INVX0_HVT U242 ( .A(n388), .Y(n383) );
  NAND2X0_HVT U243 ( .A1(n252), .A2(n263), .Y(n387) );
  INVX0_HVT U244 ( .A(n389), .Y(n385) );
  NAND2X0_HVT U245 ( .A1(n390), .A2(n316), .Y(n384) );
  AO221X1_HVT U246 ( .A1(n235), .A2(n391), .A3(n237), .A4(n275), .A5(n392), 
        .Y(n372) );
  AO22X1_HVT U247 ( .A1(n231), .A2(n250), .A3(n393), .A4(n229), .Y(n392) );
  NAND2X0_HVT U248 ( .A1(n340), .A2(n394), .Y(n391) );
  XNOR2X1_HVT U249 ( .A1(n395), .A2(keyout[92]), .Y(keyout[124]) );
  XOR3X1_HVT U250 ( .A1(keyin[60]), .A2(keyin[92]), .A3(keyout[28]), .Y(
        keyout[92]) );
  XOR2X1_HVT U251 ( .A1(keyin[28]), .A2(n396), .Y(keyout[28]) );
  MUX21X1_HVT U252 ( .A1(n397), .A2(n398), .S0(keyin[97]), .Y(n396) );
  MUX41X1_HVT U253 ( .A1(n399), .A3(n400), .A2(n401), .A4(n402), .S0(n217), 
        .S1(keyin[98]), .Y(n398) );
  AO221X1_HVT U254 ( .A1(n403), .A2(n229), .A3(n237), .A4(n404), .A5(n405), 
        .Y(n402) );
  AO22X1_HVT U255 ( .A1(n293), .A2(n235), .A3(n231), .A4(n406), .Y(n405) );
  INVX0_HVT U256 ( .A(n407), .Y(n293) );
  INVX0_HVT U257 ( .A(n390), .Y(n403) );
  AO222X1_HVT U258 ( .A1(n408), .A2(n237), .A3(n234), .A4(n409), .A5(n229), 
        .A6(n275), .Y(n401) );
  AO21X1_HVT U259 ( .A1(keyin[96]), .A2(n410), .A3(n235), .Y(n409) );
  NAND2X0_HVT U260 ( .A1(n266), .A2(n390), .Y(n410) );
  AND2X1_HVT U261 ( .A1(n246), .A2(n339), .Y(n234) );
  INVX0_HVT U262 ( .A(n411), .Y(n408) );
  AO221X1_HVT U263 ( .A1(n412), .A2(n235), .A3(n413), .A4(n3), .A5(n414), .Y(
        n400) );
  AO22X1_HVT U264 ( .A1(n415), .A2(n231), .A3(n229), .A4(n265), .Y(n414) );
  AO221X1_HVT U265 ( .A1(n231), .A2(n416), .A3(n235), .A4(n406), .A5(n417), 
        .Y(n399) );
  MUX21X1_HVT U266 ( .A1(n418), .A2(n419), .S0(n420), .Y(n417) );
  AND2X1_HVT U267 ( .A1(n334), .A2(n3), .Y(n419) );
  AO22X1_HVT U268 ( .A1(n229), .A2(keyin[99]), .A3(n237), .A4(keyin[100]), .Y(
        n418) );
  MUX41X1_HVT U269 ( .A1(n421), .A3(n422), .A2(n423), .A4(n424), .S0(n217), 
        .S1(keyin[98]), .Y(n397) );
  OAI222X1_HVT U270 ( .A1(n224), .A2(n380), .A3(n340), .A4(n297), .A5(n389), 
        .A6(n227), .Y(n424) );
  NAND3X0_HVT U271 ( .A1(n425), .A2(n310), .A3(n426), .Y(n423) );
  OA221X1_HVT U272 ( .A1(n264), .A2(n252), .A3(n332), .A4(n266), .A5(n220), 
        .Y(n426) );
  OA22X1_HVT U273 ( .A1(n265), .A2(n227), .A3(n224), .A4(n427), .Y(n310) );
  OA22X1_HVT U274 ( .A1(n297), .A2(n250), .A3(n226), .A4(n224), .Y(n425) );
  AO221X1_HVT U275 ( .A1(n277), .A2(n231), .A3(n428), .A4(n235), .A5(n429), 
        .Y(n422) );
  AO22X1_HVT U276 ( .A1(n430), .A2(n229), .A3(n237), .A4(n274), .Y(n429) );
  INVX0_HVT U277 ( .A(n431), .Y(n428) );
  INVX0_HVT U278 ( .A(n432), .Y(n277) );
  AO221X1_HVT U279 ( .A1(n433), .A2(n231), .A3(n255), .A4(n235), .A5(n434), 
        .Y(n421) );
  AO22X1_HVT U280 ( .A1(n237), .A2(n435), .A3(n436), .A4(n229), .Y(n434) );
  INVX0_HVT U281 ( .A(n437), .Y(n255) );
  XNOR2X1_HVT U282 ( .A1(keyout[91]), .A2(n438), .Y(keyout[123]) );
  XOR3X1_HVT U283 ( .A1(keyin[59]), .A2(keyin[91]), .A3(keyout[27]), .Y(
        keyout[91]) );
  MUX21X1_HVT U284 ( .A1(n439), .A2(n440), .S0(keyin[97]), .Y(keyout[27]) );
  XOR2X1_HVT U285 ( .A1(n441), .A2(keyin[27]), .Y(n440) );
  AO221X1_HVT U286 ( .A1(n286), .A2(n442), .A3(n289), .A4(n443), .A5(n444), 
        .Y(n441) );
  AO22X1_HVT U287 ( .A1(n291), .A2(n445), .A3(n284), .A4(n446), .Y(n444) );
  AO221X1_HVT U288 ( .A1(n235), .A2(n252), .A3(n447), .A4(n237), .A5(n448), 
        .Y(n446) );
  AO22X1_HVT U289 ( .A1(n231), .A2(n302), .A3(n331), .A4(n229), .Y(n448) );
  AO221X1_HVT U290 ( .A1(n231), .A2(n411), .A3(n449), .A4(n235), .A5(n450), 
        .Y(n445) );
  AO22X1_HVT U291 ( .A1(n229), .A2(n266), .A3(n451), .A4(n237), .Y(n450) );
  AND2X1_HVT U292 ( .A1(n317), .A2(n334), .Y(n451) );
  AO221X1_HVT U293 ( .A1(n433), .A2(n229), .A3(n452), .A4(n235), .A5(n453), 
        .Y(n443) );
  AO21X1_HVT U294 ( .A1(n380), .A2(n237), .A3(n454), .Y(n453) );
  AND2X1_HVT U295 ( .A1(n266), .A2(n308), .Y(n433) );
  AO222X1_HVT U296 ( .A1(n237), .A2(n455), .A3(keyin[101]), .A4(n456), .A5(
        n457), .A6(n235), .Y(n442) );
  NAND2X0_HVT U297 ( .A1(n275), .A2(n240), .Y(n456) );
  XOR2X1_HVT U298 ( .A1(n458), .A2(keyin[27]), .Y(n439) );
  AO221X1_HVT U299 ( .A1(n289), .A2(n459), .A3(n291), .A4(n460), .A5(n461), 
        .Y(n458) );
  AO22X1_HVT U300 ( .A1(n286), .A2(n462), .A3(n284), .A4(n463), .Y(n461) );
  NAND3X0_HVT U301 ( .A1(n464), .A2(n330), .A3(n465), .Y(n463) );
  OA22X1_HVT U302 ( .A1(n227), .A2(n394), .A3(n297), .A4(n413), .Y(n465) );
  AO221X1_HVT U303 ( .A1(n449), .A2(n237), .A3(n229), .A4(n317), .A5(n466), 
        .Y(n462) );
  AO22X1_HVT U304 ( .A1(n366), .A2(n235), .A3(n231), .A4(n368), .Y(n466) );
  AND2X1_HVT U305 ( .A1(n253), .A2(n394), .Y(n449) );
  AO221X1_HVT U306 ( .A1(n237), .A2(n467), .A3(n468), .A4(n406), .A5(n469), 
        .Y(n460) );
  INVX0_HVT U307 ( .A(n220), .Y(n469) );
  OR2X1_HVT U308 ( .A1(n275), .A2(n227), .Y(n220) );
  NAND2X0_HVT U309 ( .A1(n297), .A2(n470), .Y(n468) );
  NAND3X0_HVT U310 ( .A1(keyin[101]), .A2(n427), .A3(n294), .Y(n470) );
  NAND2X0_HVT U311 ( .A1(n250), .A2(n246), .Y(n467) );
  AO221X1_HVT U312 ( .A1(n471), .A2(n235), .A3(n237), .A4(n407), .A5(n472), 
        .Y(n459) );
  AO22X1_HVT U313 ( .A1(n430), .A2(n231), .A3(n473), .A4(n229), .Y(n472) );
  INVX0_HVT U314 ( .A(n474), .Y(n430) );
  NAND2X0_HVT U315 ( .A1(n307), .A2(n475), .Y(n407) );
  INVX0_HVT U316 ( .A(n316), .Y(n471) );
  XNOR2X1_HVT U317 ( .A1(n476), .A2(keyout[90]), .Y(keyout[122]) );
  XOR3X1_HVT U318 ( .A1(keyin[58]), .A2(keyin[90]), .A3(keyout[26]), .Y(
        keyout[90]) );
  XOR2X1_HVT U319 ( .A1(keyin[26]), .A2(n477), .Y(keyout[26]) );
  MUX21X1_HVT U320 ( .A1(n478), .A2(n479), .S0(keyin[97]), .Y(n477) );
  AO221X1_HVT U321 ( .A1(n286), .A2(n480), .A3(n289), .A4(n481), .A5(n482), 
        .Y(n479) );
  AO22X1_HVT U322 ( .A1(n284), .A2(n483), .A3(n291), .A4(n484), .Y(n482) );
  OAI221X1_HVT U323 ( .A1(n473), .A2(n332), .A3(n227), .A4(n309), .A5(n485), 
        .Y(n484) );
  MUX21X1_HVT U324 ( .A1(n486), .A2(n487), .S0(n360), .Y(n485) );
  XNOR2X1_HVT U325 ( .A1(n3), .A2(keyin[102]), .Y(n360) );
  NAND2X0_HVT U326 ( .A1(keyin[101]), .A2(n334), .Y(n487) );
  NAND2X0_HVT U327 ( .A1(n231), .A2(keyin[100]), .Y(n486) );
  NAND2X0_HVT U328 ( .A1(n317), .A2(n435), .Y(n309) );
  AO221X1_HVT U329 ( .A1(n237), .A2(n416), .A3(n273), .A4(n229), .A5(n488), 
        .Y(n483) );
  AO22X1_HVT U330 ( .A1(n235), .A2(n334), .A3(n412), .A4(n231), .Y(n488) );
  INVX0_HVT U331 ( .A(n250), .Y(n412) );
  AND2X1_HVT U332 ( .A1(n226), .A2(n394), .Y(n273) );
  NAND2X0_HVT U333 ( .A1(n334), .A2(n394), .Y(n416) );
  AO222X1_HVT U334 ( .A1(n303), .A2(n229), .A3(n489), .A4(n346), .A5(n331), 
        .A6(n231), .Y(n481) );
  AO21X1_HVT U335 ( .A1(n490), .A2(n264), .A3(n237), .Y(n489) );
  NAND2X0_HVT U336 ( .A1(n475), .A2(n239), .Y(n490) );
  AND2X1_HVT U337 ( .A1(n491), .A2(n239), .Y(n303) );
  AO221X1_HVT U338 ( .A1(n235), .A2(n238), .A3(n492), .A4(n231), .A5(n493), 
        .Y(n480) );
  AO22X1_HVT U339 ( .A1(n270), .A2(n229), .A3(n237), .A4(n404), .Y(n493) );
  INVX0_HVT U340 ( .A(n252), .Y(n492) );
  AO221X1_HVT U341 ( .A1(n291), .A2(n494), .A3(n289), .A4(n495), .A5(n496), 
        .Y(n478) );
  AO22X1_HVT U342 ( .A1(n284), .A2(n497), .A3(n286), .A4(n498), .Y(n496) );
  AO222X1_HVT U343 ( .A1(n237), .A2(n265), .A3(n499), .A4(n406), .A5(n300), 
        .A6(n235), .Y(n498) );
  AO21X1_HVT U344 ( .A1(n236), .A2(keyin[101]), .A3(n229), .Y(n499) );
  INVX0_HVT U345 ( .A(n365), .Y(n236) );
  AO221X1_HVT U346 ( .A1(n231), .A2(n500), .A3(n237), .A4(n435), .A5(n501), 
        .Y(n497) );
  AO22X1_HVT U347 ( .A1(n380), .A2(n235), .A3(n229), .A4(n368), .Y(n501) );
  AND2X1_HVT U348 ( .A1(n329), .A2(n239), .Y(n380) );
  NAND2X0_HVT U349 ( .A1(n475), .A2(n339), .Y(n500) );
  NAND2X0_HVT U350 ( .A1(n331), .A2(n427), .Y(n339) );
  NAND3X0_HVT U351 ( .A1(n502), .A2(n503), .A3(n504), .Y(n495) );
  OA22X1_HVT U352 ( .A1(n332), .A2(n274), .A3(n227), .A4(n431), .Y(n504) );
  NAND2X0_HVT U353 ( .A1(n435), .A2(n246), .Y(n431) );
  NAND3X0_HVT U354 ( .A1(n317), .A2(n413), .A3(n229), .Y(n503) );
  AO21X1_HVT U355 ( .A1(n248), .A2(n390), .A3(n224), .Y(n502) );
  AO221X1_HVT U356 ( .A1(n229), .A2(n265), .A3(n235), .A4(n334), .A5(n505), 
        .Y(n494) );
  AO221X1_HVT U357 ( .A1(n231), .A2(n506), .A3(n228), .A4(n237), .A5(n507), 
        .Y(n505) );
  INVX0_HVT U358 ( .A(n370), .Y(n507) );
  NAND2X0_HVT U359 ( .A1(n235), .A2(keyin[102]), .Y(n370) );
  AND2X1_HVT U360 ( .A1(n491), .A2(n340), .Y(n228) );
  NAND2X0_HVT U361 ( .A1(n226), .A2(n241), .Y(n506) );
  XNOR2X1_HVT U362 ( .A1(keyout[89]), .A2(n508), .Y(keyout[121]) );
  XOR3X1_HVT U363 ( .A1(keyin[57]), .A2(keyin[89]), .A3(keyout[25]), .Y(
        keyout[89]) );
  MUX21X1_HVT U364 ( .A1(n509), .A2(n510), .S0(keyin[97]), .Y(keyout[25]) );
  XOR2X1_HVT U365 ( .A1(n511), .A2(keyin[25]), .Y(n510) );
  AO221X1_HVT U366 ( .A1(n291), .A2(n512), .A3(n286), .A4(n513), .A5(n514), 
        .Y(n511) );
  AO22X1_HVT U367 ( .A1(n289), .A2(n515), .A3(n284), .A4(n516), .Y(n514) );
  AO221X1_HVT U368 ( .A1(n231), .A2(n517), .A3(n518), .A4(n235), .A5(n519), 
        .Y(n516) );
  AO22X1_HVT U369 ( .A1(n237), .A2(n274), .A3(n229), .A4(n308), .Y(n519) );
  NAND2X0_HVT U370 ( .A1(n346), .A2(n340), .Y(n274) );
  AO221X1_HVT U371 ( .A1(n235), .A2(n520), .A3(n229), .A4(n382), .A5(n521), 
        .Y(n515) );
  AO22X1_HVT U372 ( .A1(n231), .A2(n491), .A3(n237), .A4(n1), .Y(n521) );
  NAND2X0_HVT U373 ( .A1(n329), .A2(n307), .Y(n382) );
  NAND2X0_HVT U374 ( .A1(n266), .A2(n475), .Y(n520) );
  NAND3X0_HVT U375 ( .A1(n522), .A2(n523), .A3(n524), .Y(n513) );
  OA22X1_HVT U376 ( .A1(n276), .A2(n297), .A3(n393), .A4(n227), .Y(n524) );
  INVX0_HVT U377 ( .A(n261), .Y(n393) );
  NAND2X0_HVT U378 ( .A1(n262), .A2(n435), .Y(n261) );
  NAND3X0_HVT U379 ( .A1(n275), .A2(n240), .A3(n237), .Y(n522) );
  AO221X1_HVT U380 ( .A1(n525), .A2(n229), .A3(n518), .A4(n231), .A5(n526), 
        .Y(n512) );
  AO22X1_HVT U381 ( .A1(n237), .A2(n389), .A3(n336), .A4(n235), .Y(n526) );
  INVX0_HVT U382 ( .A(n307), .Y(n336) );
  NAND2X0_HVT U383 ( .A1(n329), .A2(n527), .Y(n389) );
  XOR2X1_HVT U384 ( .A1(n528), .A2(keyin[25]), .Y(n509) );
  AO221X1_HVT U385 ( .A1(n284), .A2(n529), .A3(n286), .A4(n530), .A5(n531), 
        .Y(n528) );
  AO22X1_HVT U386 ( .A1(n289), .A2(n532), .A3(n291), .A4(n533), .Y(n531) );
  AO221X1_HVT U387 ( .A1(n371), .A2(n237), .A3(n229), .A4(n534), .A5(n535), 
        .Y(n533) );
  AO22X1_HVT U388 ( .A1(n235), .A2(n317), .A3(n231), .A4(n368), .Y(n535) );
  NAND2X0_HVT U389 ( .A1(n307), .A2(n390), .Y(n368) );
  INVX0_HVT U390 ( .A(n475), .Y(n371) );
  AO221X1_HVT U391 ( .A1(n457), .A2(n237), .A3(n536), .A4(n229), .A5(n537), 
        .Y(n532) );
  OAI22X1_HVT U392 ( .A1(n227), .A2(n538), .A3(n315), .A4(n224), .Y(n537) );
  NAND2X0_HVT U393 ( .A1(n250), .A2(n329), .Y(n315) );
  INVX0_HVT U394 ( .A(n539), .Y(n536) );
  INVX0_HVT U395 ( .A(n534), .Y(n457) );
  NAND2X0_HVT U396 ( .A1(n246), .A2(n263), .Y(n534) );
  NAND4X0_HVT U397 ( .A1(n221), .A2(n388), .A3(n540), .A4(n541), .Y(n530) );
  OA22X1_HVT U398 ( .A1(n297), .A2(n275), .A3(n542), .A4(n227), .Y(n541) );
  NAND3X0_HVT U399 ( .A1(n226), .A2(n3), .A3(n420), .Y(n540) );
  XNOR2X1_HVT U400 ( .A1(n264), .A2(keyin[102]), .Y(n420) );
  NAND2X0_HVT U401 ( .A1(n452), .A2(n231), .Y(n388) );
  AND2X1_HVT U402 ( .A1(n265), .A2(n394), .Y(n452) );
  NAND2X0_HVT U403 ( .A1(keyin[102]), .A2(n240), .Y(n394) );
  NAND2X0_HVT U404 ( .A1(n436), .A2(n237), .Y(n221) );
  INVX0_HVT U405 ( .A(n239), .Y(n436) );
  AO221X1_HVT U406 ( .A1(n229), .A2(n248), .A3(n231), .A4(keyin[100]), .A5(
        n543), .Y(n529) );
  OAI21X1_HVT U407 ( .A1(n415), .A2(keyin[101]), .A3(n330), .Y(n543) );
  OR2X1_HVT U408 ( .A1(n455), .A2(n332), .Y(n330) );
  XNOR2X1_HVT U409 ( .A1(keyout[88]), .A2(n544), .Y(keyout[120]) );
  XOR3X1_HVT U410 ( .A1(keyin[56]), .A2(keyin[88]), .A3(keyout[24]), .Y(
        keyout[88]) );
  MUX21X1_HVT U411 ( .A1(n545), .A2(n546), .S0(keyin[97]), .Y(keyout[24]) );
  XOR2X1_HVT U412 ( .A1(n547), .A2(keyin[24]), .Y(n546) );
  AO221X1_HVT U413 ( .A1(n284), .A2(n548), .A3(n286), .A4(n549), .A5(n550), 
        .Y(n547) );
  AO22X1_HVT U414 ( .A1(n289), .A2(n551), .A3(n291), .A4(n552), .Y(n550) );
  AO221X1_HVT U415 ( .A1(n542), .A2(n231), .A3(n235), .A4(n226), .A5(n553), 
        .Y(n552) );
  AO221X1_HVT U416 ( .A1(n237), .A2(n413), .A3(n300), .A4(n229), .A5(n247), 
        .Y(n553) );
  NOR2X0_HVT U417 ( .A1(n435), .A2(n224), .Y(n247) );
  INVX0_HVT U418 ( .A(n364), .Y(n300) );
  NAND2X0_HVT U419 ( .A1(n252), .A2(n316), .Y(n364) );
  NAND2X0_HVT U420 ( .A1(n265), .A2(n427), .Y(n316) );
  INVX0_HVT U421 ( .A(n491), .Y(n542) );
  AO221X1_HVT U422 ( .A1(n231), .A2(n554), .A3(n235), .A4(n555), .A5(n556), 
        .Y(n551) );
  AO22X1_HVT U423 ( .A1(n229), .A2(n250), .A3(n237), .A4(n262), .Y(n556) );
  NAND2X0_HVT U424 ( .A1(n1), .A2(n427), .Y(n250) );
  NAND2X0_HVT U425 ( .A1(n253), .A2(n475), .Y(n555) );
  NAND2X0_HVT U426 ( .A1(n294), .A2(keyin[102]), .Y(n475) );
  INVX0_HVT U427 ( .A(n334), .Y(n294) );
  NAND2X0_HVT U428 ( .A1(n308), .A2(n239), .Y(n554) );
  NAND2X0_HVT U429 ( .A1(n313), .A2(n427), .Y(n239) );
  NAND2X0_HVT U430 ( .A1(keyin[102]), .A2(n1), .Y(n308) );
  AO221X1_HVT U431 ( .A1(n518), .A2(n235), .A3(n356), .A4(keyin[101]), .A5(
        n557), .Y(n549) );
  OAI22X1_HVT U432 ( .A1(n342), .A2(n224), .A3(n262), .A4(n332), .Y(n557) );
  NAND2X0_HVT U433 ( .A1(n238), .A2(n527), .Y(n342) );
  INVX0_HVT U434 ( .A(n346), .Y(n356) );
  AND2X1_HVT U435 ( .A1(n241), .A2(n340), .Y(n518) );
  AO221X1_HVT U436 ( .A1(n447), .A2(n229), .A3(n235), .A4(n302), .A5(n558), 
        .Y(n548) );
  AO21X1_HVT U437 ( .A1(n237), .A2(n539), .A3(n454), .Y(n558) );
  INVX0_HVT U438 ( .A(n464), .Y(n454) );
  NAND2X0_HVT U439 ( .A1(n231), .A2(n265), .Y(n464) );
  NAND2X0_HVT U440 ( .A1(n253), .A2(n390), .Y(n539) );
  NAND2X0_HVT U441 ( .A1(n270), .A2(keyin[102]), .Y(n390) );
  NAND2X0_HVT U442 ( .A1(n334), .A2(n427), .Y(n253) );
  OAI21X1_HVT U443 ( .A1(n334), .A2(keyin[102]), .A3(n238), .Y(n302) );
  AND2X1_HVT U444 ( .A1(n346), .A2(n307), .Y(n447) );
  NAND2X0_HVT U445 ( .A1(n413), .A2(n427), .Y(n307) );
  NAND2X0_HVT U446 ( .A1(n331), .A2(keyin[102]), .Y(n346) );
  INVX0_HVT U447 ( .A(n265), .Y(n331) );
  XOR2X1_HVT U448 ( .A1(n559), .A2(keyin[24]), .Y(n545) );
  AO221X1_HVT U449 ( .A1(n284), .A2(n560), .A3(n291), .A4(n561), .A5(n562), 
        .Y(n559) );
  AO22X1_HVT U450 ( .A1(n289), .A2(n563), .A3(n286), .A4(n564), .Y(n562) );
  AO221X1_HVT U451 ( .A1(n379), .A2(n231), .A3(n525), .A4(n235), .A5(n565), 
        .Y(n564) );
  AO22X1_HVT U452 ( .A1(n229), .A2(n275), .A3(n237), .A4(keyin[99]), .Y(n565)
         );
  AND2X1_HVT U453 ( .A1(n317), .A2(n340), .Y(n525) );
  NAND2X0_HVT U454 ( .A1(keyin[102]), .A2(n226), .Y(n317) );
  INVX0_HVT U455 ( .A(n406), .Y(n379) );
  NAND2X0_HVT U456 ( .A1(n241), .A2(n527), .Y(n406) );
  NAND2X0_HVT U457 ( .A1(n226), .A2(n427), .Y(n527) );
  INVX0_HVT U458 ( .A(n320), .Y(n286) );
  NAND2X0_HVT U459 ( .A1(n217), .A2(n2), .Y(n320) );
  AO221X1_HVT U460 ( .A1(n473), .A2(n566), .A3(n229), .A4(n432), .A5(n567), 
        .Y(n563) );
  INVX0_HVT U461 ( .A(n523), .Y(n567) );
  NAND3X0_HVT U462 ( .A1(n231), .A2(n241), .A3(n270), .Y(n523) );
  NAND2X0_HVT U463 ( .A1(n252), .A2(n365), .Y(n432) );
  AO21X1_HVT U464 ( .A1(n437), .A2(n264), .A3(n237), .Y(n566) );
  NAND2X0_HVT U465 ( .A1(n238), .A2(n365), .Y(n437) );
  INVX0_HVT U466 ( .A(n517), .Y(n473) );
  NAND2X0_HVT U467 ( .A1(n248), .A2(n246), .Y(n517) );
  NAND2X0_HVT U468 ( .A1(n538), .A2(keyin[102]), .Y(n246) );
  INVX0_HVT U469 ( .A(n325), .Y(n289) );
  NAND2X0_HVT U470 ( .A1(keyin[103]), .A2(keyin[98]), .Y(n325) );
  AO221X1_HVT U471 ( .A1(n231), .A2(n455), .A3(n415), .A4(n235), .A5(n568), 
        .Y(n561) );
  OAI221X1_HVT U472 ( .A1(n240), .A2(n332), .A3(n297), .A4(n276), .A5(n298), 
        .Y(n568) );
  NAND2X0_HVT U473 ( .A1(n366), .A2(n237), .Y(n298) );
  INVX0_HVT U474 ( .A(n241), .Y(n366) );
  NAND2X0_HVT U475 ( .A1(keyin[102]), .A2(n265), .Y(n241) );
  NAND2X0_HVT U476 ( .A1(keyin[99]), .A2(n313), .Y(n265) );
  INVX0_HVT U477 ( .A(n404), .Y(n276) );
  NAND2X0_HVT U478 ( .A1(n226), .A2(n491), .Y(n404) );
  NAND2X0_HVT U479 ( .A1(keyin[102]), .A2(n413), .Y(n491) );
  AND2X1_HVT U480 ( .A1(n248), .A2(n252), .Y(n415) );
  NAND2X0_HVT U481 ( .A1(n299), .A2(n427), .Y(n248) );
  NAND2X0_HVT U482 ( .A1(n262), .A2(n365), .Y(n455) );
  NAND2X0_HVT U483 ( .A1(n270), .A2(n427), .Y(n365) );
  INVX0_HVT U484 ( .A(n413), .Y(n270) );
  NAND2X0_HVT U485 ( .A1(n226), .A2(n240), .Y(n413) );
  NAND2X0_HVT U486 ( .A1(keyin[102]), .A2(keyin[100]), .Y(n262) );
  INVX0_HVT U487 ( .A(n327), .Y(n291) );
  NAND2X0_HVT U488 ( .A1(keyin[98]), .A2(n217), .Y(n327) );
  AO221X1_HVT U489 ( .A1(n229), .A2(n569), .A3(n235), .A4(n570), .A5(n571), 
        .Y(n560) );
  AO22X1_HVT U490 ( .A1(n231), .A2(n474), .A3(n237), .A4(n411), .Y(n571) );
  NAND2X0_HVT U491 ( .A1(n340), .A2(n238), .Y(n411) );
  NAND2X0_HVT U492 ( .A1(keyin[102]), .A2(n299), .Y(n238) );
  INVX0_HVT U493 ( .A(n226), .Y(n299) );
  NAND2X0_HVT U494 ( .A1(keyin[100]), .A2(keyin[99]), .Y(n226) );
  NAND2X0_HVT U495 ( .A1(keyin[99]), .A2(n427), .Y(n340) );
  INVX0_HVT U496 ( .A(n332), .Y(n237) );
  NAND2X0_HVT U497 ( .A1(n264), .A2(n3), .Y(n332) );
  NAND2X0_HVT U498 ( .A1(n329), .A2(n266), .Y(n474) );
  NAND2X0_HVT U499 ( .A1(n538), .A2(n427), .Y(n266) );
  INVX0_HVT U500 ( .A(n240), .Y(n538) );
  NAND2X0_HVT U501 ( .A1(keyin[102]), .A2(keyin[99]), .Y(n329) );
  INVX0_HVT U502 ( .A(n224), .Y(n231) );
  NAND2X0_HVT U503 ( .A1(keyin[101]), .A2(keyin[96]), .Y(n224) );
  NAND2X0_HVT U504 ( .A1(n435), .A2(n252), .Y(n570) );
  NAND2X0_HVT U505 ( .A1(keyin[102]), .A2(n313), .Y(n252) );
  NAND2X0_HVT U506 ( .A1(n427), .A2(n240), .Y(n435) );
  NAND2X0_HVT U507 ( .A1(n1), .A2(n313), .Y(n240) );
  INVX0_HVT U508 ( .A(n227), .Y(n235) );
  NAND2X0_HVT U509 ( .A1(keyin[96]), .A2(n264), .Y(n227) );
  NAND2X0_HVT U510 ( .A1(n275), .A2(n263), .Y(n569) );
  NAND2X0_HVT U511 ( .A1(keyin[100]), .A2(n427), .Y(n263) );
  NAND2X0_HVT U512 ( .A1(keyin[102]), .A2(n334), .Y(n275) );
  NAND2X0_HVT U513 ( .A1(keyin[100]), .A2(n1), .Y(n334) );
  INVX0_HVT U514 ( .A(keyin[99]), .Y(n1) );
  INVX0_HVT U515 ( .A(n297), .Y(n229) );
  NAND2X0_HVT U516 ( .A1(keyin[101]), .A2(n3), .Y(n297) );
  INVX0_HVT U517 ( .A(keyin[96]), .Y(n3) );
  INVX0_HVT U518 ( .A(n322), .Y(n284) );
  NAND2X0_HVT U519 ( .A1(keyin[103]), .A2(n2), .Y(n322) );
  INVX0_HVT U520 ( .A(keyin[98]), .Y(n2) );
  XNOR2X1_HVT U521 ( .A1(keyout[87]), .A2(n572), .Y(keyout[119]) );
  XNOR3X1_HVT U522 ( .A1(keyin[87]), .A2(keyin[55]), .A3(n17), .Y(keyout[87])
         );
  XNOR2X1_HVT U523 ( .A1(n573), .A2(keyin[23]), .Y(n17) );
  AO221X1_HVT U524 ( .A1(n574), .A2(n575), .A3(n576), .A4(n577), .A5(n578), 
        .Y(n573) );
  AO22X1_HVT U525 ( .A1(n579), .A2(n580), .A3(n581), .A4(n582), .Y(n578) );
  NAND2X0_HVT U526 ( .A1(n583), .A2(n584), .Y(n582) );
  OA222X1_HVT U527 ( .A1(n585), .A2(n586), .A3(n587), .A4(n588), .A5(
        keyin[125]), .A6(n589), .Y(n584) );
  OA22X1_HVT U528 ( .A1(n590), .A2(n591), .A3(n592), .A4(n593), .Y(n589) );
  OA21X1_HVT U529 ( .A1(n594), .A2(n595), .A3(n596), .Y(n587) );
  OA222X1_HVT U530 ( .A1(n597), .A2(n598), .A3(n599), .A4(n600), .A5(n601), 
        .A6(n602), .Y(n583) );
  NAND3X0_HVT U531 ( .A1(n603), .A2(n604), .A3(n605), .Y(n580) );
  OA222X1_HVT U532 ( .A1(n395), .A2(n595), .A3(n597), .A4(n606), .A5(n596), 
        .A6(n607), .Y(n605) );
  OA22X1_HVT U533 ( .A1(n585), .A2(n608), .A3(keyin[125]), .A4(n609), .Y(n604)
         );
  OA221X1_HVT U534 ( .A1(n610), .A2(n591), .A3(n611), .A4(n592), .A5(n612), 
        .Y(n609) );
  AOI22X1_HVT U535 ( .A1(n613), .A2(n614), .A3(n615), .A4(n616), .Y(n603) );
  NAND4X0_HVT U536 ( .A1(n617), .A2(n618), .A3(n619), .A4(n620), .Y(n577) );
  OA221X1_HVT U537 ( .A1(n621), .A2(n599), .A3(n622), .A4(n623), .A5(n624), 
        .Y(n620) );
  OA22X1_HVT U538 ( .A1(n601), .A2(n625), .A3(n597), .A4(n613), .Y(n624) );
  NAND2X0_HVT U539 ( .A1(n626), .A2(n627), .Y(n613) );
  OA22X1_HVT U540 ( .A1(n628), .A2(n629), .A3(n630), .A4(n585), .Y(n619) );
  AO21X1_HVT U541 ( .A1(n629), .A2(n631), .A3(n596), .Y(n618) );
  AO21X1_HVT U542 ( .A1(n632), .A2(n633), .A3(n595), .Y(n617) );
  AO221X1_HVT U543 ( .A1(n616), .A2(n634), .A3(n635), .A4(n636), .A5(n637), 
        .Y(n575) );
  AO222X1_HVT U544 ( .A1(n638), .A2(n280), .A3(n639), .A4(n640), .A5(n641), 
        .A6(n642), .Y(n637) );
  INVX0_HVT U545 ( .A(n643), .Y(n640) );
  AOI21X1_HVT U546 ( .A1(n644), .A2(keyin[125]), .A3(keyin[120]), .Y(n639) );
  AO21X1_HVT U547 ( .A1(keyin[125]), .A2(n645), .A3(n646), .Y(n638) );
  AO22X1_HVT U548 ( .A1(keyin[122]), .A2(keyin[124]), .A3(keyin[120]), .A4(
        n610), .Y(n645) );
  INVX0_HVT U549 ( .A(n647), .Y(n636) );
  XNOR2X1_HVT U550 ( .A1(n648), .A2(keyout[86]), .Y(keyout[118]) );
  XOR3X1_HVT U551 ( .A1(keyin[54]), .A2(keyin[86]), .A3(keyout[22]), .Y(
        keyout[86]) );
  XOR2X1_HVT U552 ( .A1(keyin[22]), .A2(n649), .Y(keyout[22]) );
  MUX21X1_HVT U553 ( .A1(n650), .A2(n651), .S0(n211), .Y(n649) );
  AO221X1_HVT U554 ( .A1(n652), .A2(n653), .A3(n654), .A4(n655), .A5(n656), 
        .Y(n651) );
  AO22X1_HVT U555 ( .A1(n657), .A2(n658), .A3(n659), .A4(n660), .Y(n656) );
  AO221X1_HVT U556 ( .A1(n661), .A2(n662), .A3(n663), .A4(n664), .A5(n665), 
        .Y(n660) );
  AO22X1_HVT U557 ( .A1(n666), .A2(n667), .A3(n668), .A4(n600), .Y(n665) );
  AO221X1_HVT U558 ( .A1(n669), .A2(n668), .A3(n670), .A4(n667), .A5(n671), 
        .Y(n658) );
  AO22X1_HVT U559 ( .A1(n664), .A2(n647), .A3(n672), .A4(n662), .Y(n671) );
  AO221X1_HVT U560 ( .A1(n673), .A2(n668), .A3(n674), .A4(n667), .A5(n675), 
        .Y(n655) );
  AO22X1_HVT U561 ( .A1(n663), .A2(n662), .A3(n664), .A4(n676), .Y(n675) );
  NAND2X0_HVT U562 ( .A1(n677), .A2(n678), .Y(n676) );
  AND2X1_HVT U563 ( .A1(n679), .A2(n680), .Y(n663) );
  NAND3X0_HVT U564 ( .A1(n681), .A2(n682), .A3(n683), .Y(n653) );
  OA22X1_HVT U565 ( .A1(n684), .A2(n685), .A3(n611), .A4(n591), .Y(n683) );
  INVX0_HVT U566 ( .A(n686), .Y(n611) );
  NAND3X0_HVT U567 ( .A1(n687), .A2(n644), .A3(n667), .Y(n681) );
  AO221X1_HVT U568 ( .A1(n652), .A2(n688), .A3(n654), .A4(n689), .A5(n690), 
        .Y(n650) );
  AO22X1_HVT U569 ( .A1(n657), .A2(n691), .A3(n659), .A4(n692), .Y(n690) );
  AO221X1_HVT U570 ( .A1(n664), .A2(n693), .A3(n694), .A4(n667), .A5(n695), 
        .Y(n692) );
  AO22X1_HVT U571 ( .A1(n668), .A2(n696), .A3(n662), .A4(n607), .Y(n695) );
  INVX0_HVT U572 ( .A(n680), .Y(n694) );
  NAND2X0_HVT U573 ( .A1(n697), .A2(n698), .Y(n693) );
  AO221X1_HVT U574 ( .A1(n664), .A2(n699), .A3(n667), .A4(n700), .A5(n701), 
        .Y(n691) );
  MUX21X1_HVT U575 ( .A1(n662), .A2(n668), .S0(n702), .Y(n701) );
  NAND2X0_HVT U576 ( .A1(n696), .A2(n644), .Y(n700) );
  NAND2X0_HVT U577 ( .A1(n677), .A2(n703), .Y(n699) );
  AO221X1_HVT U578 ( .A1(n664), .A2(n704), .A3(n705), .A4(n668), .A5(n706), 
        .Y(n689) );
  AO22X1_HVT U579 ( .A1(n662), .A2(n707), .A3(n667), .A4(n680), .Y(n706) );
  AO222X1_HVT U580 ( .A1(n708), .A2(n664), .A3(n709), .A4(n710), .A5(n667), 
        .A6(n602), .Y(n688) );
  OAI21X1_HVT U581 ( .A1(n678), .A2(n476), .A3(n592), .Y(n710) );
  AND2X1_HVT U582 ( .A1(n697), .A2(n687), .Y(n709) );
  INVX0_HVT U583 ( .A(n607), .Y(n708) );
  NAND2X0_HVT U584 ( .A1(n633), .A2(n711), .Y(n607) );
  XNOR2X1_HVT U585 ( .A1(keyout[85]), .A2(n712), .Y(keyout[117]) );
  XOR3X1_HVT U586 ( .A1(keyin[53]), .A2(keyin[85]), .A3(keyout[21]), .Y(
        keyout[85]) );
  XOR2X1_HVT U587 ( .A1(n713), .A2(keyin[21]), .Y(keyout[21]) );
  AO221X1_HVT U588 ( .A1(n581), .A2(n714), .A3(n579), .A4(n715), .A5(n716), 
        .Y(n713) );
  AO22X1_HVT U589 ( .A1(n576), .A2(n717), .A3(n574), .A4(n718), .Y(n716) );
  NAND4X0_HVT U590 ( .A1(n719), .A2(n720), .A3(n721), .A4(n722), .Y(n718) );
  OA221X1_HVT U591 ( .A1(n601), .A2(n723), .A3(n647), .A4(n599), .A5(n724), 
        .Y(n722) );
  OA22X1_HVT U592 ( .A1(n597), .A2(n725), .A3(n726), .A4(n596), .Y(n724) );
  OA22X1_HVT U593 ( .A1(n628), .A2(n727), .A3(n594), .A4(n622), .Y(n721) );
  AO21X1_HVT U594 ( .A1(n626), .A2(n680), .A3(n585), .Y(n720) );
  AO21X1_HVT U595 ( .A1(n728), .A2(n703), .A3(n595), .Y(n719) );
  NAND4X0_HVT U596 ( .A1(n729), .A2(n730), .A3(n731), .A4(n732), .Y(n717) );
  OA222X1_HVT U597 ( .A1(n280), .A2(n595), .A3(n622), .A4(n680), .A5(n601), 
        .A6(n733), .Y(n732) );
  OA22X1_HVT U598 ( .A1(n734), .A2(n596), .A3(n628), .A4(n697), .Y(n731) );
  AND2X1_HVT U599 ( .A1(n735), .A2(n623), .Y(n734) );
  NAND3X0_HVT U600 ( .A1(keyin[125]), .A2(n544), .A3(n736), .Y(n730) );
  AO21X1_HVT U601 ( .A1(n737), .A2(n633), .A3(n597), .Y(n729) );
  NAND4X0_HVT U602 ( .A1(n738), .A2(n739), .A3(n740), .A4(n741), .Y(n715) );
  OA221X1_HVT U603 ( .A1(n670), .A2(n595), .A3(n596), .A4(n697), .A5(n742), 
        .Y(n741) );
  MUX21X1_HVT U604 ( .A1(n743), .A2(n679), .S0(n347), .Y(n742) );
  OA21X1_HVT U605 ( .A1(n476), .A2(n606), .A3(n744), .Y(n743) );
  MUX21X1_HVT U606 ( .A1(n745), .A2(n746), .S0(n747), .Y(n744) );
  NAND2X0_HVT U607 ( .A1(n664), .A2(keyin[124]), .Y(n746) );
  NAND2X0_HVT U608 ( .A1(n687), .A2(n476), .Y(n745) );
  OA22X1_HVT U609 ( .A1(n642), .A2(n599), .A3(n601), .A4(n608), .Y(n740) );
  NAND2X0_HVT U610 ( .A1(n627), .A2(n677), .Y(n608) );
  NAND3X0_HVT U611 ( .A1(n747), .A2(n438), .A3(n641), .Y(n739) );
  NAND2X0_HVT U612 ( .A1(n748), .A2(n749), .Y(n738) );
  INVX0_HVT U613 ( .A(n622), .Y(n748) );
  AO221X1_HVT U614 ( .A1(n614), .A2(n602), .A3(n750), .A4(n616), .A5(n751), 
        .Y(n714) );
  AO222X1_HVT U615 ( .A1(n752), .A2(n476), .A3(n753), .A4(n754), .A5(n635), 
        .A6(n698), .Y(n751) );
  NAND2X0_HVT U616 ( .A1(n596), .A2(n622), .Y(n754) );
  MUX21X1_HVT U617 ( .A1(n755), .A2(n756), .S0(n347), .Y(n752) );
  INVX0_HVT U618 ( .A(n601), .Y(n616) );
  NAND2X0_HVT U619 ( .A1(n697), .A2(n627), .Y(n602) );
  XNOR2X1_HVT U620 ( .A1(keyout[84]), .A2(n757), .Y(keyout[116]) );
  XOR3X1_HVT U621 ( .A1(keyin[52]), .A2(keyin[84]), .A3(keyout[20]), .Y(
        keyout[84]) );
  XOR2X1_HVT U622 ( .A1(n758), .A2(keyin[20]), .Y(keyout[20]) );
  AO221X1_HVT U623 ( .A1(n574), .A2(n759), .A3(n576), .A4(n760), .A5(n761), 
        .Y(n758) );
  AO22X1_HVT U624 ( .A1(n579), .A2(n762), .A3(n581), .A4(n763), .Y(n761) );
  NAND4X0_HVT U625 ( .A1(n764), .A2(n765), .A3(n766), .A4(n767), .Y(n763) );
  OA221X1_HVT U626 ( .A1(n643), .A2(n595), .A3(n597), .A4(n768), .A5(n769), 
        .Y(n767) );
  AOI22X1_HVT U627 ( .A1(n770), .A2(n646), .A3(n614), .A4(n726), .Y(n769) );
  INVX0_HVT U628 ( .A(n596), .Y(n646) );
  OA22X1_HVT U629 ( .A1(n771), .A2(n628), .A3(n622), .A4(n772), .Y(n766) );
  INVX0_HVT U630 ( .A(n606), .Y(n771) );
  NAND3X0_HVT U631 ( .A1(n773), .A2(n395), .A3(keyin[125]), .Y(n765) );
  AO21X1_HVT U632 ( .A1(keyin[122]), .A2(keyin[126]), .A3(n774), .Y(n773) );
  AO21X1_HVT U633 ( .A1(n696), .A2(n633), .A3(n601), .Y(n764) );
  AND2X1_HVT U634 ( .A1(keyin[127]), .A2(n508), .Y(n581) );
  NAND3X0_HVT U635 ( .A1(n775), .A2(n776), .A3(n777), .Y(n762) );
  AOI222X1_HVT U636 ( .A1(n778), .A2(n635), .A3(n779), .A4(n641), .A5(n633), 
        .A6(n614), .Y(n777) );
  INVX0_HVT U637 ( .A(n599), .Y(n614) );
  INVX0_HVT U638 ( .A(n597), .Y(n641) );
  INVX0_HVT U639 ( .A(n595), .Y(n635) );
  AO21X1_HVT U640 ( .A1(n601), .A2(n780), .A3(n625), .Y(n776) );
  NAND2X0_HVT U641 ( .A1(n735), .A2(n698), .Y(n625) );
  AO21X1_HVT U642 ( .A1(n728), .A2(n772), .A3(n684), .Y(n780) );
  OA22X1_HVT U643 ( .A1(n591), .A2(n781), .A3(n622), .A4(n782), .Y(n775) );
  MUX21X1_HVT U644 ( .A1(n783), .A2(n669), .S0(n784), .Y(n781) );
  XNOR2X1_HVT U645 ( .A1(n280), .A2(keyin[125]), .Y(n784) );
  MUX21X1_HVT U646 ( .A1(n438), .A2(n395), .S0(n347), .Y(n783) );
  AND2X1_HVT U647 ( .A1(keyin[127]), .A2(keyin[121]), .Y(n579) );
  NAND4X0_HVT U648 ( .A1(n785), .A2(n786), .A3(n787), .A4(n788), .Y(n760) );
  OA22X1_HVT U649 ( .A1(n634), .A2(n585), .A3(n789), .A4(n622), .Y(n788) );
  NAND2X0_HVT U650 ( .A1(n662), .A2(n347), .Y(n622) );
  OA22X1_HVT U651 ( .A1(n599), .A2(n728), .A3(n601), .A4(n790), .Y(n787) );
  OA22X1_HVT U652 ( .A1(n597), .A2(n791), .A3(n750), .A4(n596), .Y(n786) );
  OA22X1_HVT U653 ( .A1(n595), .A2(n615), .A3(n737), .A4(n591), .Y(n785) );
  AND2X1_HVT U654 ( .A1(keyin[121]), .A2(n211), .Y(n576) );
  NAND3X0_HVT U655 ( .A1(n792), .A2(n793), .A3(n794), .Y(n759) );
  OA222X1_HVT U656 ( .A1(n595), .A2(n795), .A3(n597), .A4(n600), .A5(n796), 
        .A6(n596), .Y(n794) );
  NAND2X0_HVT U657 ( .A1(n668), .A2(keyin[125]), .Y(n596) );
  NAND2X0_HVT U658 ( .A1(n667), .A2(keyin[125]), .Y(n597) );
  NAND2X0_HVT U659 ( .A1(n667), .A2(n347), .Y(n595) );
  OA22X1_HVT U660 ( .A1(n797), .A2(n628), .A3(n585), .A4(n798), .Y(n793) );
  NAND2X0_HVT U661 ( .A1(n664), .A2(keyin[125]), .Y(n585) );
  NAND2X0_HVT U662 ( .A1(n664), .A2(n347), .Y(n628) );
  OA22X1_HVT U663 ( .A1(n599), .A2(n711), .A3(n601), .A4(n727), .Y(n792) );
  NAND2X0_HVT U664 ( .A1(n668), .A2(n347), .Y(n601) );
  NAND2X0_HVT U665 ( .A1(n662), .A2(keyin[125]), .Y(n599) );
  AND2X1_HVT U666 ( .A1(n508), .A2(n211), .Y(n574) );
  XNOR2X1_HVT U667 ( .A1(keyin[115]), .A2(n4), .Y(keyout[115]) );
  XNOR3X1_HVT U668 ( .A1(keyin[83]), .A2(keyin[51]), .A3(keyout[19]), .Y(n4)
         );
  XNOR2X1_HVT U669 ( .A1(n799), .A2(keyin[19]), .Y(keyout[19]) );
  MUX21X1_HVT U670 ( .A1(n800), .A2(n801), .S0(n211), .Y(n799) );
  AOI221X1_HVT U671 ( .A1(n657), .A2(n802), .A3(n654), .A4(n803), .A5(n804), 
        .Y(n801) );
  AO22X1_HVT U672 ( .A1(n659), .A2(n805), .A3(n652), .A4(n806), .Y(n804) );
  AO222X1_HVT U673 ( .A1(n664), .A2(n644), .A3(n807), .A4(n778), .A5(n667), 
        .A6(n749), .Y(n806) );
  NAND2X0_HVT U674 ( .A1(n592), .A2(n808), .Y(n807) );
  NAND3X0_HVT U675 ( .A1(keyin[122]), .A2(n280), .A3(n669), .Y(n808) );
  AO221X1_HVT U676 ( .A1(n662), .A2(n723), .A3(n809), .A4(n664), .A5(n810), 
        .Y(n805) );
  AO22X1_HVT U677 ( .A1(n672), .A2(n667), .A3(n594), .A4(n668), .Y(n810) );
  INVX0_HVT U678 ( .A(n633), .Y(n594) );
  INVX0_HVT U679 ( .A(n697), .Y(n672) );
  NAND2X0_HVT U680 ( .A1(n615), .A2(n735), .Y(n723) );
  AO222X1_HVT U681 ( .A1(n662), .A2(n772), .A3(n811), .A4(n476), .A5(n668), 
        .A6(n782), .Y(n803) );
  AO221X1_HVT U682 ( .A1(n812), .A2(n662), .A3(n664), .A4(n813), .A5(n814), 
        .Y(n802) );
  AO22X1_HVT U683 ( .A1(n815), .A2(n667), .A3(n809), .A4(n668), .Y(n814) );
  AND2X1_HVT U684 ( .A1(n627), .A2(n816), .Y(n809) );
  AND2X1_HVT U685 ( .A1(n687), .A2(n644), .Y(n812) );
  OA221X1_HVT U686 ( .A1(n817), .A2(n818), .A3(n819), .A4(n591), .A5(n820), 
        .Y(n800) );
  OA221X1_HVT U687 ( .A1(n821), .A2(n592), .A3(n822), .A4(n684), .A5(n823), 
        .Y(n820) );
  NAND3X0_HVT U688 ( .A1(n657), .A2(keyin[122]), .A3(n755), .Y(n823) );
  MUX21X1_HVT U689 ( .A1(n824), .A2(n796), .S0(n544), .Y(n755) );
  OA22X1_HVT U690 ( .A1(n634), .A2(n825), .A3(n826), .A4(n798), .Y(n822) );
  OA21X1_HVT U691 ( .A1(keyin[126]), .A2(n827), .A3(n828), .Y(n825) );
  OA222X1_HVT U692 ( .A1(n673), .A2(n827), .A3(n826), .A4(n829), .A5(n828), 
        .A6(n768), .Y(n821) );
  NAND2X0_HVT U693 ( .A1(n677), .A2(n772), .Y(n768) );
  INVX0_HVT U694 ( .A(n790), .Y(n673) );
  NAND2X0_HVT U695 ( .A1(n678), .A2(n830), .Y(n790) );
  OA221X1_HVT U696 ( .A1(n831), .A2(n832), .A3(n827), .A4(n813), .A5(n833), 
        .Y(n819) );
  OA22X1_HVT U697 ( .A1(n588), .A2(n826), .A3(n696), .A4(n828), .Y(n833) );
  OA221X1_HVT U698 ( .A1(n834), .A2(n828), .A3(n634), .A4(n826), .A5(n835), 
        .Y(n817) );
  OA22X1_HVT U699 ( .A1(n827), .A2(n816), .A3(n836), .A4(n831), .Y(n835) );
  INVX0_HVT U700 ( .A(n626), .Y(n836) );
  XNOR2X1_HVT U701 ( .A1(n837), .A2(keyout[82]), .Y(keyout[114]) );
  XOR3X1_HVT U702 ( .A1(keyin[50]), .A2(keyin[82]), .A3(keyout[18]), .Y(
        keyout[82]) );
  XOR2X1_HVT U703 ( .A1(keyin[18]), .A2(n838), .Y(keyout[18]) );
  MUX21X1_HVT U704 ( .A1(n839), .A2(n840), .S0(n211), .Y(n838) );
  AO221X1_HVT U705 ( .A1(n659), .A2(n841), .A3(n657), .A4(n842), .A5(n843), 
        .Y(n840) );
  AO22X1_HVT U706 ( .A1(n652), .A2(n844), .A3(n654), .A4(n845), .Y(n843) );
  OAI221X1_HVT U707 ( .A1(n818), .A2(n626), .A3(n588), .A4(n591), .A5(n846), 
        .Y(n845) );
  MUX21X1_HVT U708 ( .A1(n847), .A2(n848), .S0(n747), .Y(n846) );
  XNOR2X1_HVT U709 ( .A1(n544), .A2(keyin[126]), .Y(n747) );
  NAND2X0_HVT U710 ( .A1(keyin[122]), .A2(n687), .Y(n848) );
  NAND2X0_HVT U711 ( .A1(n668), .A2(keyin[124]), .Y(n847) );
  AO222X1_HVT U712 ( .A1(n849), .A2(n778), .A3(n668), .A4(n850), .A5(n662), 
        .A6(n696), .Y(n844) );
  NAND2X0_HVT U713 ( .A1(n697), .A2(n632), .Y(n850) );
  OAI21X1_HVT U714 ( .A1(n623), .A2(keyin[122]), .A3(n591), .Y(n849) );
  AO221X1_HVT U715 ( .A1(n664), .A2(n593), .A3(n670), .A4(n668), .A5(n851), 
        .Y(n842) );
  AO22X1_HVT U716 ( .A1(n662), .A2(n829), .A3(n667), .A4(n631), .Y(n851) );
  AND2X1_HVT U717 ( .A1(n644), .A2(n606), .Y(n670) );
  AO221X1_HVT U718 ( .A1(n668), .A2(n852), .A3(n662), .A4(n853), .A5(n854), 
        .Y(n841) );
  AO22X1_HVT U719 ( .A1(n705), .A2(n667), .A3(n664), .A4(n696), .Y(n854) );
  INVX0_HVT U720 ( .A(n630), .Y(n853) );
  NAND2X0_HVT U721 ( .A1(n855), .A2(n711), .Y(n630) );
  NAND2X0_HVT U722 ( .A1(n669), .A2(n280), .Y(n852) );
  AO221X1_HVT U723 ( .A1(n654), .A2(n856), .A3(n659), .A4(n857), .A5(n858), 
        .Y(n839) );
  AO22X1_HVT U724 ( .A1(n657), .A2(n859), .A3(n652), .A4(n860), .Y(n858) );
  AO221X1_HVT U725 ( .A1(n861), .A2(n644), .A3(n664), .A4(n749), .A5(n862), 
        .Y(n860) );
  AO22X1_HVT U726 ( .A1(n667), .A2(n863), .A3(n668), .A4(n864), .Y(n862) );
  NAND2X0_HVT U727 ( .A1(n686), .A2(n728), .Y(n864) );
  NAND2X0_HVT U728 ( .A1(n830), .A2(n698), .Y(n863) );
  NAND2X0_HVT U729 ( .A1(n634), .A2(n280), .Y(n698) );
  AO222X1_HVT U730 ( .A1(n664), .A2(n779), .A3(n865), .A4(n679), .A5(n667), 
        .A6(n687), .Y(n859) );
  AO21X1_HVT U731 ( .A1(keyin[122]), .A2(n866), .A3(n662), .Y(n865) );
  NAND2X0_HVT U732 ( .A1(n629), .A2(n830), .Y(n866) );
  NAND2X0_HVT U733 ( .A1(n687), .A2(n816), .Y(n779) );
  AO221X1_HVT U734 ( .A1(n867), .A2(n668), .A3(n796), .A4(n667), .A5(n868), 
        .Y(n857) );
  AO22X1_HVT U735 ( .A1(n664), .A2(n606), .A3(n797), .A4(n662), .Y(n868) );
  INVX0_HVT U736 ( .A(n598), .Y(n797) );
  AND2X1_HVT U737 ( .A1(n629), .A2(n685), .Y(n796) );
  INVX0_HVT U738 ( .A(n795), .Y(n867) );
  NAND2X0_HVT U739 ( .A1(n606), .A2(n735), .Y(n795) );
  AO221X1_HVT U740 ( .A1(n674), .A2(n662), .A3(n753), .A4(n664), .A5(n869), 
        .Y(n856) );
  AO22X1_HVT U741 ( .A1(n726), .A2(n667), .A3(n634), .A4(n668), .Y(n869) );
  INVX0_HVT U742 ( .A(n615), .Y(n726) );
  INVX0_HVT U743 ( .A(n586), .Y(n753) );
  NAND2X0_HVT U744 ( .A1(n632), .A2(n816), .Y(n586) );
  AND2X1_HVT U745 ( .A1(n855), .A2(n629), .Y(n674) );
  XNOR2X1_HVT U746 ( .A1(n870), .A2(keyout[81]), .Y(keyout[113]) );
  XOR3X1_HVT U747 ( .A1(keyin[49]), .A2(keyin[81]), .A3(keyout[17]), .Y(
        keyout[81]) );
  XOR2X1_HVT U748 ( .A1(keyin[17]), .A2(n871), .Y(keyout[17]) );
  MUX21X1_HVT U749 ( .A1(n872), .A2(n873), .S0(n211), .Y(n871) );
  AO221X1_HVT U750 ( .A1(n652), .A2(n874), .A3(n659), .A4(n875), .A5(n876), 
        .Y(n873) );
  OAI22X1_HVT U751 ( .A1(n877), .A2(n831), .A3(n878), .A4(n828), .Y(n876) );
  OA221X1_HVT U752 ( .A1(n684), .A2(n879), .A3(n789), .A4(n591), .A5(n880), 
        .Y(n878) );
  OA22X1_HVT U753 ( .A1(n818), .A2(n881), .A3(n592), .A4(n882), .Y(n880) );
  NAND2X0_HVT U754 ( .A1(n737), .A2(n697), .Y(n881) );
  INVX0_HVT U755 ( .A(n593), .Y(n789) );
  OA221X1_HVT U756 ( .A1(n684), .A2(n678), .A3(n591), .A4(n811), .A5(n883), 
        .Y(n877) );
  AOI22X1_HVT U757 ( .A1(n727), .A2(n662), .A3(n647), .A4(n667), .Y(n883) );
  NAND2X0_HVT U758 ( .A1(n606), .A2(n884), .Y(n647) );
  NAND2X0_HVT U759 ( .A1(n770), .A2(n685), .Y(n727) );
  NAND2X0_HVT U760 ( .A1(n633), .A2(n885), .Y(n811) );
  AO221X1_HVT U761 ( .A1(n668), .A2(n644), .A3(n667), .A4(n855), .A5(n886), 
        .Y(n875) );
  AO22X1_HVT U762 ( .A1(n736), .A2(n662), .A3(n664), .A4(n887), .Y(n886) );
  NAND2X0_HVT U763 ( .A1(n644), .A2(n629), .Y(n887) );
  AO221X1_HVT U764 ( .A1(n664), .A2(n888), .A3(n662), .A4(n889), .A5(n890), 
        .Y(n874) );
  AO22X1_HVT U765 ( .A1(n824), .A2(n667), .A3(n668), .A4(n749), .Y(n890) );
  NAND2X0_HVT U766 ( .A1(n728), .A2(n678), .Y(n749) );
  INVX0_HVT U767 ( .A(n725), .Y(n824) );
  NAND2X0_HVT U768 ( .A1(n696), .A2(n816), .Y(n725) );
  NAND2X0_HVT U769 ( .A1(keyin[126]), .A2(n885), .Y(n816) );
  NAND2X0_HVT U770 ( .A1(n633), .A2(n770), .Y(n888) );
  AO221X1_HVT U771 ( .A1(n654), .A2(n891), .A3(n657), .A4(n892), .A5(n893), 
        .Y(n872) );
  AO22X1_HVT U772 ( .A1(n652), .A2(n894), .A3(n659), .A4(n895), .Y(n893) );
  AO222X1_HVT U773 ( .A1(n815), .A2(n662), .A3(n661), .A4(n896), .A5(n668), 
        .A6(n885), .Y(n895) );
  AO21X1_HVT U774 ( .A1(n791), .A2(n476), .A3(n664), .Y(n896) );
  INVX0_HVT U775 ( .A(n813), .Y(n661) );
  INVX0_HVT U776 ( .A(n889), .Y(n815) );
  NAND2X0_HVT U777 ( .A1(n735), .A2(n680), .Y(n889) );
  AO221X1_HVT U778 ( .A1(n664), .A2(n686), .A3(n897), .A4(n662), .A5(n898), 
        .Y(n894) );
  OAI22X1_HVT U779 ( .A1(n818), .A2(n395), .A3(n704), .A4(n684), .Y(n898) );
  NAND2X0_HVT U780 ( .A1(n615), .A2(n685), .Y(n704) );
  INVX0_HVT U781 ( .A(n899), .Y(n897) );
  AO221X1_HVT U782 ( .A1(n664), .A2(n598), .A3(n900), .A4(n667), .A5(n901), 
        .Y(n892) );
  AO22X1_HVT U783 ( .A1(n662), .A2(n438), .A3(n668), .A4(n902), .Y(n901) );
  NAND2X0_HVT U784 ( .A1(n772), .A2(n830), .Y(n902) );
  NAND2X0_HVT U785 ( .A1(n679), .A2(n711), .Y(n598) );
  AO221X1_HVT U786 ( .A1(n668), .A2(n855), .A3(n667), .A4(n829), .A5(n903), 
        .Y(n891) );
  AO21X1_HVT U787 ( .A1(n756), .A2(n544), .A3(n774), .Y(n903) );
  INVX0_HVT U788 ( .A(n612), .Y(n774) );
  NAND2X0_HVT U789 ( .A1(n664), .A2(n280), .Y(n612) );
  NAND2X0_HVT U790 ( .A1(n685), .A2(n678), .Y(n756) );
  XNOR2X1_HVT U791 ( .A1(n904), .A2(keyout[80]), .Y(keyout[112]) );
  XOR3X1_HVT U792 ( .A1(keyin[48]), .A2(keyin[80]), .A3(keyout[16]), .Y(
        keyout[80]) );
  XOR2X1_HVT U793 ( .A1(keyin[16]), .A2(n905), .Y(keyout[16]) );
  MUX21X1_HVT U794 ( .A1(n906), .A2(n907), .S0(n211), .Y(n905) );
  INVX0_HVT U795 ( .A(keyin[127]), .Y(n211) );
  AO221X1_HVT U796 ( .A1(n652), .A2(n908), .A3(n657), .A4(n909), .A5(n910), 
        .Y(n907) );
  AO22X1_HVT U797 ( .A1(n659), .A2(n911), .A3(n654), .A4(n912), .Y(n910) );
  AO221X1_HVT U798 ( .A1(n668), .A2(n913), .A3(n705), .A4(n662), .A5(n914), 
        .Y(n912) );
  AO22X1_HVT U799 ( .A1(n915), .A2(n476), .A3(n666), .A4(n667), .Y(n914) );
  AND2X1_HVT U800 ( .A1(n631), .A2(n770), .Y(n666) );
  INVX0_HVT U801 ( .A(n679), .Y(n915) );
  INVX0_HVT U802 ( .A(n733), .Y(n705) );
  NAND2X0_HVT U803 ( .A1(n626), .A2(n703), .Y(n733) );
  NAND2X0_HVT U804 ( .A1(n696), .A2(n280), .Y(n703) );
  NAND2X0_HVT U805 ( .A1(n855), .A2(n606), .Y(n913) );
  OAI221X1_HVT U806 ( .A1(n791), .A2(n684), .A3(n882), .A4(n818), .A5(n916), 
        .Y(n911) );
  OA22X1_HVT U807 ( .A1(n591), .A2(n438), .A3(n592), .A4(n621), .Y(n916) );
  AND2X1_HVT U808 ( .A1(n885), .A2(n697), .Y(n621) );
  NAND2X0_HVT U809 ( .A1(n644), .A2(n711), .Y(n882) );
  NAND2X0_HVT U810 ( .A1(keyin[126]), .A2(n632), .Y(n644) );
  NAND2X0_HVT U811 ( .A1(n686), .A2(n626), .Y(n791) );
  AO221X1_HVT U812 ( .A1(n668), .A2(n632), .A3(n900), .A4(n667), .A5(n917), 
        .Y(n909) );
  AO21X1_HVT U813 ( .A1(n664), .A2(n642), .A3(n861), .Y(n917) );
  INVX0_HVT U814 ( .A(n682), .Y(n861) );
  NAND2X0_HVT U815 ( .A1(n662), .A2(n588), .Y(n682) );
  INVX0_HVT U816 ( .A(n884), .Y(n642) );
  INVX0_HVT U817 ( .A(n879), .Y(n900) );
  NAND2X0_HVT U818 ( .A1(n697), .A2(n711), .Y(n879) );
  AO221X1_HVT U819 ( .A1(n662), .A2(n593), .A3(n664), .A4(n633), .A5(n918), 
        .Y(n908) );
  AO22X1_HVT U820 ( .A1(n750), .A2(n667), .A3(n668), .A4(n813), .Y(n918) );
  NAND2X0_HVT U821 ( .A1(n884), .A2(n623), .Y(n813) );
  INVX0_HVT U822 ( .A(n778), .Y(n750) );
  NAND2X0_HVT U823 ( .A1(n697), .A2(n770), .Y(n778) );
  NAND2X0_HVT U824 ( .A1(n632), .A2(n280), .Y(n770) );
  NAND2X0_HVT U825 ( .A1(n632), .A2(n855), .Y(n593) );
  NAND2X0_HVT U826 ( .A1(keyin[126]), .A2(n588), .Y(n855) );
  AO221X1_HVT U827 ( .A1(n659), .A2(n919), .A3(n657), .A4(n920), .A5(n921), 
        .Y(n906) );
  AO22X1_HVT U828 ( .A1(n654), .A2(n922), .A3(n652), .A4(n923), .Y(n921) );
  NAND3X0_HVT U829 ( .A1(n924), .A2(n925), .A3(n926), .Y(n923) );
  AOI22X1_HVT U830 ( .A1(n600), .A2(n662), .A3(n798), .A4(n667), .Y(n926) );
  NAND2X0_HVT U831 ( .A1(n772), .A2(n685), .Y(n798) );
  NAND2X0_HVT U832 ( .A1(keyin[126]), .A2(keyin[123]), .Y(n685) );
  NAND2X0_HVT U833 ( .A1(n610), .A2(n280), .Y(n772) );
  NAND2X0_HVT U834 ( .A1(n626), .A2(n623), .Y(n600) );
  NAND3X0_HVT U835 ( .A1(n737), .A2(n697), .A3(n668), .Y(n925) );
  NAND2X0_HVT U836 ( .A1(keyin[126]), .A2(n696), .Y(n697) );
  AO21X1_HVT U837 ( .A1(n633), .A2(n680), .A3(n591), .Y(n924) );
  NAND2X0_HVT U838 ( .A1(keyin[124]), .A2(n280), .Y(n680) );
  NAND2X0_HVT U839 ( .A1(keyin[126]), .A2(n687), .Y(n633) );
  INVX0_HVT U840 ( .A(n826), .Y(n652) );
  NAND2X0_HVT U841 ( .A1(keyin[125]), .A2(n508), .Y(n826) );
  AO221X1_HVT U842 ( .A1(n927), .A2(n664), .A3(n667), .A4(n696), .A5(n928), 
        .Y(n922) );
  AO22X1_HVT U843 ( .A1(n662), .A2(n615), .A3(n668), .A4(n929), .Y(n928) );
  NAND2X0_HVT U844 ( .A1(n629), .A2(n677), .Y(n929) );
  NAND2X0_HVT U845 ( .A1(keyin[126]), .A2(n438), .Y(n677) );
  NAND2X0_HVT U846 ( .A1(n395), .A2(n280), .Y(n629) );
  NAND2X0_HVT U847 ( .A1(n280), .A2(n438), .Y(n615) );
  INVX0_HVT U848 ( .A(n832), .Y(n927) );
  NAND2X0_HVT U849 ( .A1(n679), .A2(n678), .Y(n832) );
  NAND2X0_HVT U850 ( .A1(n588), .A2(n280), .Y(n678) );
  NAND2X0_HVT U851 ( .A1(n634), .A2(keyin[126]), .Y(n679) );
  INVX0_HVT U852 ( .A(n696), .Y(n634) );
  NAND2X0_HVT U853 ( .A1(keyin[123]), .A2(n395), .Y(n696) );
  INVX0_HVT U854 ( .A(n828), .Y(n654) );
  NAND2X0_HVT U855 ( .A1(keyin[121]), .A2(keyin[125]), .Y(n828) );
  AO221X1_HVT U856 ( .A1(n664), .A2(n899), .A3(n667), .A4(n702), .A5(n930), 
        .Y(n920) );
  AO222X1_HVT U857 ( .A1(n662), .A2(n884), .A3(n736), .A4(n668), .A5(n590), 
        .A6(keyin[122]), .Y(n930) );
  INVX0_HVT U858 ( .A(n627), .Y(n590) );
  INVX0_HVT U859 ( .A(n684), .Y(n668) );
  NAND2X0_HVT U860 ( .A1(keyin[122]), .A2(keyin[120]), .Y(n684) );
  INVX0_HVT U861 ( .A(n830), .Y(n736) );
  NAND2X0_HVT U862 ( .A1(n669), .A2(keyin[126]), .Y(n830) );
  INVX0_HVT U863 ( .A(n687), .Y(n669) );
  NAND2X0_HVT U864 ( .A1(keyin[126]), .A2(keyin[124]), .Y(n884) );
  INVX0_HVT U865 ( .A(n834), .Y(n702) );
  OA21X1_HVT U866 ( .A1(n687), .A2(keyin[126]), .A3(n631), .Y(n834) );
  NAND2X0_HVT U867 ( .A1(n627), .A2(n728), .Y(n899) );
  NAND2X0_HVT U868 ( .A1(n737), .A2(keyin[126]), .Y(n728) );
  NAND2X0_HVT U869 ( .A1(n687), .A2(n280), .Y(n627) );
  NAND2X0_HVT U870 ( .A1(keyin[124]), .A2(n438), .Y(n687) );
  INVX0_HVT U871 ( .A(n831), .Y(n657) );
  NAND2X0_HVT U872 ( .A1(keyin[121]), .A2(n347), .Y(n831) );
  AO222X1_HVT U873 ( .A1(n931), .A2(n932), .A3(n667), .A4(n933), .A5(n664), 
        .A6(n782), .Y(n919) );
  NAND2X0_HVT U874 ( .A1(n711), .A2(n631), .Y(n782) );
  NAND2X0_HVT U875 ( .A1(keyin[123]), .A2(n280), .Y(n711) );
  INVX0_HVT U876 ( .A(n591), .Y(n664) );
  NAND2X0_HVT U877 ( .A1(n544), .A2(n476), .Y(n591) );
  NAND2X0_HVT U878 ( .A1(n606), .A2(n626), .Y(n933) );
  NAND2X0_HVT U879 ( .A1(keyin[126]), .A2(n395), .Y(n626) );
  NAND2X0_HVT U880 ( .A1(n280), .A2(n885), .Y(n606) );
  INVX0_HVT U881 ( .A(n818), .Y(n667) );
  NAND2X0_HVT U882 ( .A1(keyin[120]), .A2(n476), .Y(n818) );
  INVX0_HVT U883 ( .A(keyin[122]), .Y(n476) );
  AO21X1_HVT U884 ( .A1(keyin[122]), .A2(n643), .A3(n662), .Y(n932) );
  INVX0_HVT U885 ( .A(n592), .Y(n662) );
  NAND2X0_HVT U886 ( .A1(keyin[122]), .A2(n544), .Y(n592) );
  INVX0_HVT U887 ( .A(keyin[120]), .Y(n544) );
  NAND2X0_HVT U888 ( .A1(n631), .A2(n623), .Y(n643) );
  NAND2X0_HVT U889 ( .A1(n737), .A2(n280), .Y(n623) );
  INVX0_HVT U890 ( .A(n588), .Y(n737) );
  NAND2X0_HVT U891 ( .A1(n885), .A2(n632), .Y(n588) );
  NAND2X0_HVT U892 ( .A1(n707), .A2(keyin[126]), .Y(n631) );
  INVX0_HVT U893 ( .A(n829), .Y(n931) );
  NAND2X0_HVT U894 ( .A1(n686), .A2(n735), .Y(n829) );
  NAND2X0_HVT U895 ( .A1(n610), .A2(keyin[126]), .Y(n735) );
  INVX0_HVT U896 ( .A(n885), .Y(n610) );
  NAND2X0_HVT U897 ( .A1(n395), .A2(n438), .Y(n885) );
  INVX0_HVT U898 ( .A(keyin[123]), .Y(n438) );
  INVX0_HVT U899 ( .A(keyin[124]), .Y(n395) );
  NAND2X0_HVT U900 ( .A1(n707), .A2(n280), .Y(n686) );
  INVX0_HVT U901 ( .A(keyin[126]), .Y(n280) );
  INVX0_HVT U902 ( .A(n632), .Y(n707) );
  NAND2X0_HVT U903 ( .A1(keyin[124]), .A2(keyin[123]), .Y(n632) );
  INVX0_HVT U904 ( .A(n827), .Y(n659) );
  NAND2X0_HVT U905 ( .A1(n508), .A2(n347), .Y(n827) );
  INVX0_HVT U906 ( .A(keyin[125]), .Y(n347) );
  INVX0_HVT U907 ( .A(keyin[121]), .Y(n508) );
  XNOR2X1_HVT U908 ( .A1(keyout[79]), .A2(n26), .Y(keyout[111]) );
  XNOR3X1_HVT U909 ( .A1(keyin[79]), .A2(keyin[47]), .A3(n20), .Y(keyout[79])
         );
  XNOR2X1_HVT U910 ( .A1(n934), .A2(keyin[15]), .Y(n20) );
  AO221X1_HVT U911 ( .A1(n935), .A2(n936), .A3(n937), .A4(n938), .A5(n939), 
        .Y(n934) );
  AO22X1_HVT U912 ( .A1(n940), .A2(n941), .A3(n942), .A4(n943), .Y(n939) );
  NAND2X0_HVT U913 ( .A1(n944), .A2(n945), .Y(n943) );
  OA222X1_HVT U914 ( .A1(n946), .A2(n947), .A3(n948), .A4(n949), .A5(
        keyin[117]), .A6(n950), .Y(n945) );
  OA22X1_HVT U915 ( .A1(n951), .A2(n952), .A3(n953), .A4(n954), .Y(n950) );
  OA21X1_HVT U916 ( .A1(n955), .A2(n956), .A3(n957), .Y(n948) );
  OA222X1_HVT U917 ( .A1(n958), .A2(n959), .A3(n960), .A4(n961), .A5(n962), 
        .A6(n963), .Y(n944) );
  NAND3X0_HVT U918 ( .A1(n964), .A2(n965), .A3(n966), .Y(n941) );
  OA222X1_HVT U919 ( .A1(n757), .A2(n956), .A3(n958), .A4(n967), .A5(n957), 
        .A6(n968), .Y(n966) );
  OA22X1_HVT U920 ( .A1(n946), .A2(n969), .A3(keyin[117]), .A4(n970), .Y(n965)
         );
  OA221X1_HVT U921 ( .A1(n971), .A2(n952), .A3(n972), .A4(n953), .A5(n973), 
        .Y(n970) );
  AOI22X1_HVT U922 ( .A1(n974), .A2(n975), .A3(n976), .A4(n977), .Y(n964) );
  NAND4X0_HVT U923 ( .A1(n978), .A2(n979), .A3(n980), .A4(n981), .Y(n938) );
  OA221X1_HVT U924 ( .A1(n982), .A2(n960), .A3(n983), .A4(n984), .A5(n985), 
        .Y(n981) );
  OA22X1_HVT U925 ( .A1(n962), .A2(n986), .A3(n958), .A4(n974), .Y(n985) );
  NAND2X0_HVT U926 ( .A1(n987), .A2(n988), .Y(n974) );
  OA22X1_HVT U927 ( .A1(n989), .A2(n990), .A3(n991), .A4(n946), .Y(n980) );
  AO21X1_HVT U928 ( .A1(n990), .A2(n992), .A3(n957), .Y(n979) );
  AO21X1_HVT U929 ( .A1(n993), .A2(n994), .A3(n956), .Y(n978) );
  AO221X1_HVT U930 ( .A1(n977), .A2(n995), .A3(n996), .A4(n997), .A5(n998), 
        .Y(n936) );
  AO221X1_HVT U931 ( .A1(n999), .A2(n648), .A3(n1000), .A4(n1001), .A5(n1002), 
        .Y(n998) );
  AND3X1_HVT U932 ( .A1(n1003), .A2(n904), .A3(n1004), .Y(n1002) );
  NAND2X0_HVT U933 ( .A1(keyin[117]), .A2(n1005), .Y(n1004) );
  INVX0_HVT U934 ( .A(n1006), .Y(n1003) );
  AO21X1_HVT U935 ( .A1(keyin[117]), .A2(n1007), .A3(n1008), .Y(n999) );
  AO22X1_HVT U936 ( .A1(keyin[114]), .A2(keyin[116]), .A3(keyin[112]), .A4(
        n971), .Y(n1007) );
  INVX0_HVT U937 ( .A(n1009), .Y(n997) );
  XNOR2X1_HVT U938 ( .A1(n44), .A2(keyout[78]), .Y(keyout[110]) );
  XOR3X1_HVT U939 ( .A1(keyin[46]), .A2(keyin[78]), .A3(keyout[14]), .Y(
        keyout[78]) );
  XOR2X1_HVT U940 ( .A1(keyin[14]), .A2(n1010), .Y(keyout[14]) );
  MUX21X1_HVT U941 ( .A1(n1011), .A2(n1012), .S0(n572), .Y(n1010) );
  AO221X1_HVT U942 ( .A1(n1013), .A2(n1014), .A3(n1015), .A4(n1016), .A5(n1017), .Y(n1012) );
  AO22X1_HVT U943 ( .A1(n1018), .A2(n1019), .A3(n1020), .A4(n1021), .Y(n1017)
         );
  AO221X1_HVT U944 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .A5(n1026), .Y(n1021) );
  AO22X1_HVT U945 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n961), .Y(n1026)
         );
  AO221X1_HVT U946 ( .A1(n1030), .A2(n1029), .A3(n1031), .A4(n1028), .A5(n1032), .Y(n1019) );
  AO22X1_HVT U947 ( .A1(n1025), .A2(n1009), .A3(n1033), .A4(n1022), .Y(n1032)
         );
  AO221X1_HVT U948 ( .A1(n1034), .A2(n1029), .A3(n1035), .A4(n1028), .A5(n1036), .Y(n1016) );
  AO22X1_HVT U949 ( .A1(n1024), .A2(n1022), .A3(n1025), .A4(n1037), .Y(n1036)
         );
  NAND2X0_HVT U950 ( .A1(n1038), .A2(n1039), .Y(n1037) );
  AND2X1_HVT U951 ( .A1(n1040), .A2(n1041), .Y(n1024) );
  NAND3X0_HVT U952 ( .A1(n1042), .A2(n1043), .A3(n1044), .Y(n1014) );
  OA22X1_HVT U953 ( .A1(n1045), .A2(n1046), .A3(n972), .A4(n952), .Y(n1044) );
  INVX0_HVT U954 ( .A(n1047), .Y(n972) );
  NAND3X0_HVT U955 ( .A1(n1048), .A2(n1005), .A3(n1028), .Y(n1042) );
  AO221X1_HVT U956 ( .A1(n1013), .A2(n1049), .A3(n1015), .A4(n1050), .A5(n1051), .Y(n1011) );
  AO22X1_HVT U957 ( .A1(n1018), .A2(n1052), .A3(n1020), .A4(n1053), .Y(n1051)
         );
  AO221X1_HVT U958 ( .A1(n1025), .A2(n1054), .A3(n1055), .A4(n1028), .A5(n1056), .Y(n1053) );
  AO22X1_HVT U959 ( .A1(n1029), .A2(n1057), .A3(n1022), .A4(n968), .Y(n1056)
         );
  INVX0_HVT U960 ( .A(n1041), .Y(n1055) );
  NAND2X0_HVT U961 ( .A1(n1058), .A2(n1059), .Y(n1054) );
  AO221X1_HVT U962 ( .A1(n1025), .A2(n1060), .A3(n1028), .A4(n1061), .A5(n1062), .Y(n1052) );
  MUX21X1_HVT U963 ( .A1(n1022), .A2(n1029), .S0(n1063), .Y(n1062) );
  NAND2X0_HVT U964 ( .A1(n1057), .A2(n1005), .Y(n1061) );
  NAND2X0_HVT U965 ( .A1(n1038), .A2(n1064), .Y(n1060) );
  AO221X1_HVT U966 ( .A1(n1025), .A2(n1065), .A3(n1066), .A4(n1029), .A5(n1067), .Y(n1050) );
  AO22X1_HVT U967 ( .A1(n1022), .A2(n1068), .A3(n1028), .A4(n1041), .Y(n1067)
         );
  AO222X1_HVT U968 ( .A1(n1069), .A2(n1025), .A3(n1070), .A4(n1071), .A5(n1028), .A6(n963), .Y(n1049) );
  OAI21X1_HVT U969 ( .A1(n1039), .A2(n837), .A3(n953), .Y(n1071) );
  AND2X1_HVT U970 ( .A1(n1058), .A2(n1048), .Y(n1070) );
  INVX0_HVT U971 ( .A(n968), .Y(n1069) );
  NAND2X0_HVT U972 ( .A1(n994), .A2(n1072), .Y(n968) );
  XNOR2X1_HVT U973 ( .A1(keyout[77]), .A2(n1073), .Y(keyout[109]) );
  XOR3X1_HVT U974 ( .A1(keyin[45]), .A2(keyin[77]), .A3(keyout[13]), .Y(
        keyout[77]) );
  XOR2X1_HVT U975 ( .A1(n1074), .A2(keyin[13]), .Y(keyout[13]) );
  AO221X1_HVT U976 ( .A1(n942), .A2(n1075), .A3(n940), .A4(n1076), .A5(n1077), 
        .Y(n1074) );
  AO22X1_HVT U977 ( .A1(n937), .A2(n1078), .A3(n935), .A4(n1079), .Y(n1077) );
  NAND4X0_HVT U978 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .Y(n1079)
         );
  OA221X1_HVT U979 ( .A1(n1084), .A2(n957), .A3(n1085), .A4(n958), .A5(n1086), 
        .Y(n1083) );
  OA22X1_HVT U980 ( .A1(n1009), .A2(n960), .A3(n962), .A4(n1087), .Y(n1086) );
  OA22X1_HVT U981 ( .A1(n989), .A2(n1088), .A3(n955), .A4(n983), .Y(n1082) );
  AO21X1_HVT U982 ( .A1(n987), .A2(n1041), .A3(n946), .Y(n1081) );
  AO21X1_HVT U983 ( .A1(n1089), .A2(n1064), .A3(n956), .Y(n1080) );
  NAND4X0_HVT U984 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .Y(n1078)
         );
  OA222X1_HVT U985 ( .A1(n648), .A2(n956), .A3(n983), .A4(n1041), .A5(n1094), 
        .A6(n962), .Y(n1093) );
  OA22X1_HVT U986 ( .A1(n1095), .A2(n957), .A3(n989), .A4(n1058), .Y(n1092) );
  AND2X1_HVT U987 ( .A1(n1096), .A2(n984), .Y(n1095) );
  NAND3X0_HVT U988 ( .A1(keyin[117]), .A2(n904), .A3(n1097), .Y(n1091) );
  AO21X1_HVT U989 ( .A1(n1098), .A2(n994), .A3(n958), .Y(n1090) );
  NAND4X0_HVT U990 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .Y(n1076)
         );
  OA221X1_HVT U991 ( .A1(n1031), .A2(n956), .A3(n957), .A4(n1058), .A5(n1103), 
        .Y(n1102) );
  MUX21X1_HVT U992 ( .A1(n1104), .A2(n1040), .S0(n712), .Y(n1103) );
  OA21X1_HVT U993 ( .A1(n837), .A2(n967), .A3(n1105), .Y(n1104) );
  MUX21X1_HVT U994 ( .A1(n1106), .A2(n1107), .S0(n1108), .Y(n1105) );
  NAND2X0_HVT U995 ( .A1(n1025), .A2(keyin[116]), .Y(n1107) );
  NAND2X0_HVT U996 ( .A1(n1048), .A2(n837), .Y(n1106) );
  OA22X1_HVT U997 ( .A1(n1001), .A2(n960), .A3(n962), .A4(n969), .Y(n1101) );
  NAND2X0_HVT U998 ( .A1(n988), .A2(n1038), .Y(n969) );
  NAND3X0_HVT U999 ( .A1(n1108), .A2(n1109), .A3(n1000), .Y(n1100) );
  NAND2X0_HVT U1000 ( .A1(n1110), .A2(n1111), .Y(n1099) );
  INVX0_HVT U1001 ( .A(n983), .Y(n1110) );
  AO221X1_HVT U1002 ( .A1(n975), .A2(n963), .A3(n977), .A4(n1112), .A5(n1113), 
        .Y(n1075) );
  AO222X1_HVT U1003 ( .A1(n1114), .A2(n837), .A3(n1115), .A4(n1116), .A5(n996), 
        .A6(n1059), .Y(n1113) );
  NAND2X0_HVT U1004 ( .A1(n957), .A2(n983), .Y(n1116) );
  MUX21X1_HVT U1005 ( .A1(n1117), .A2(n1118), .S0(n712), .Y(n1114) );
  INVX0_HVT U1006 ( .A(n962), .Y(n977) );
  NAND2X0_HVT U1007 ( .A1(n1058), .A2(n988), .Y(n963) );
  XNOR2X1_HVT U1008 ( .A1(keyout[76]), .A2(n199), .Y(keyout[108]) );
  XOR3X1_HVT U1009 ( .A1(keyin[44]), .A2(keyin[76]), .A3(keyout[12]), .Y(
        keyout[76]) );
  XOR2X1_HVT U1010 ( .A1(n1119), .A2(keyin[12]), .Y(keyout[12]) );
  AO221X1_HVT U1011 ( .A1(n935), .A2(n1120), .A3(n937), .A4(n1121), .A5(n1122), 
        .Y(n1119) );
  AO22X1_HVT U1012 ( .A1(n940), .A2(n1123), .A3(n942), .A4(n1124), .Y(n1122)
         );
  NAND4X0_HVT U1013 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .Y(n1124) );
  OA221X1_HVT U1014 ( .A1(n1006), .A2(n956), .A3(n958), .A4(n1129), .A5(n1130), 
        .Y(n1128) );
  AOI22X1_HVT U1015 ( .A1(n1131), .A2(n1008), .A3(n975), .A4(n1084), .Y(n1130)
         );
  INVX0_HVT U1016 ( .A(n957), .Y(n1008) );
  OA22X1_HVT U1017 ( .A1(n1132), .A2(n989), .A3(n983), .A4(n1133), .Y(n1127)
         );
  INVX0_HVT U1018 ( .A(n967), .Y(n1132) );
  NAND3X0_HVT U1019 ( .A1(n1134), .A2(n757), .A3(keyin[117]), .Y(n1126) );
  AO21X1_HVT U1020 ( .A1(keyin[114]), .A2(keyin[118]), .A3(n1135), .Y(n1134)
         );
  AO21X1_HVT U1021 ( .A1(n1057), .A2(n994), .A3(n962), .Y(n1125) );
  AND2X1_HVT U1022 ( .A1(keyin[119]), .A2(n870), .Y(n942) );
  NAND3X0_HVT U1023 ( .A1(n1136), .A2(n1137), .A3(n1138), .Y(n1123) );
  AOI222X1_HVT U1024 ( .A1(n1139), .A2(n996), .A3(n1140), .A4(n1000), .A5(n994), .A6(n975), .Y(n1138) );
  INVX0_HVT U1025 ( .A(n960), .Y(n975) );
  INVX0_HVT U1026 ( .A(n958), .Y(n1000) );
  INVX0_HVT U1027 ( .A(n956), .Y(n996) );
  AO21X1_HVT U1028 ( .A1(n962), .A2(n1141), .A3(n986), .Y(n1137) );
  NAND2X0_HVT U1029 ( .A1(n1096), .A2(n1059), .Y(n986) );
  AO21X1_HVT U1030 ( .A1(n1089), .A2(n1133), .A3(n1045), .Y(n1141) );
  OA22X1_HVT U1031 ( .A1(n952), .A2(n1142), .A3(n983), .A4(n1143), .Y(n1136)
         );
  MUX21X1_HVT U1032 ( .A1(n1144), .A2(n1030), .S0(n1145), .Y(n1142) );
  XNOR2X1_HVT U1033 ( .A1(n648), .A2(keyin[117]), .Y(n1145) );
  MUX21X1_HVT U1034 ( .A1(n1109), .A2(n757), .S0(n712), .Y(n1144) );
  AND2X1_HVT U1035 ( .A1(keyin[119]), .A2(keyin[113]), .Y(n940) );
  NAND4X0_HVT U1036 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .Y(n1121) );
  OA22X1_HVT U1037 ( .A1(n995), .A2(n946), .A3(n1150), .A4(n983), .Y(n1149) );
  NAND2X0_HVT U1038 ( .A1(n1022), .A2(n712), .Y(n983) );
  OA22X1_HVT U1039 ( .A1(n960), .A2(n1089), .A3(n962), .A4(n1151), .Y(n1148)
         );
  OA22X1_HVT U1040 ( .A1(n1152), .A2(n958), .A3(n1112), .A4(n957), .Y(n1147)
         );
  OA22X1_HVT U1041 ( .A1(n956), .A2(n976), .A3(n1098), .A4(n952), .Y(n1146) );
  AND2X1_HVT U1042 ( .A1(keyin[113]), .A2(n572), .Y(n937) );
  NAND3X0_HVT U1043 ( .A1(n1153), .A2(n1154), .A3(n1155), .Y(n1120) );
  OA222X1_HVT U1044 ( .A1(n956), .A2(n1156), .A3(n958), .A4(n961), .A5(n1157), 
        .A6(n957), .Y(n1155) );
  NAND2X0_HVT U1045 ( .A1(keyin[117]), .A2(n1029), .Y(n957) );
  NAND2X0_HVT U1046 ( .A1(n1028), .A2(keyin[117]), .Y(n958) );
  NAND2X0_HVT U1047 ( .A1(n1028), .A2(n712), .Y(n956) );
  OA22X1_HVT U1048 ( .A1(n1158), .A2(n989), .A3(n946), .A4(n1159), .Y(n1154)
         );
  NAND2X0_HVT U1049 ( .A1(n1025), .A2(keyin[117]), .Y(n946) );
  NAND2X0_HVT U1050 ( .A1(n1025), .A2(n712), .Y(n989) );
  OA22X1_HVT U1051 ( .A1(n960), .A2(n1072), .A3(n962), .A4(n1088), .Y(n1153)
         );
  NAND2X0_HVT U1052 ( .A1(n1029), .A2(n712), .Y(n962) );
  NAND2X0_HVT U1053 ( .A1(keyin[117]), .A2(n1022), .Y(n960) );
  AND2X1_HVT U1054 ( .A1(n870), .A2(n572), .Y(n935) );
  XNOR2X1_HVT U1055 ( .A1(keyin[107]), .A2(n5), .Y(keyout[107]) );
  XNOR3X1_HVT U1056 ( .A1(keyin[75]), .A2(keyin[43]), .A3(keyout[11]), .Y(n5)
         );
  XNOR2X1_HVT U1057 ( .A1(n1160), .A2(keyin[11]), .Y(keyout[11]) );
  MUX21X1_HVT U1058 ( .A1(n1161), .A2(n1162), .S0(n572), .Y(n1160) );
  AOI221X1_HVT U1059 ( .A1(n1018), .A2(n1163), .A3(n1015), .A4(n1164), .A5(
        n1165), .Y(n1162) );
  AO22X1_HVT U1060 ( .A1(n1020), .A2(n1166), .A3(n1013), .A4(n1167), .Y(n1165)
         );
  AO222X1_HVT U1061 ( .A1(n1025), .A2(n1005), .A3(n1168), .A4(n1139), .A5(
        n1028), .A6(n1111), .Y(n1167) );
  NAND2X0_HVT U1062 ( .A1(n953), .A2(n1169), .Y(n1168) );
  NAND3X0_HVT U1063 ( .A1(keyin[114]), .A2(n648), .A3(n1030), .Y(n1169) );
  AO221X1_HVT U1064 ( .A1(n1022), .A2(n1087), .A3(n1170), .A4(n1025), .A5(
        n1171), .Y(n1166) );
  AO22X1_HVT U1065 ( .A1(n1033), .A2(n1028), .A3(n955), .A4(n1029), .Y(n1171)
         );
  INVX0_HVT U1066 ( .A(n994), .Y(n955) );
  INVX0_HVT U1067 ( .A(n1058), .Y(n1033) );
  NAND2X0_HVT U1068 ( .A1(n976), .A2(n1096), .Y(n1087) );
  AO222X1_HVT U1069 ( .A1(n1022), .A2(n1133), .A3(n1172), .A4(n837), .A5(n1029), .A6(n1143), .Y(n1164) );
  AO221X1_HVT U1070 ( .A1(n1173), .A2(n1022), .A3(n1025), .A4(n1174), .A5(
        n1175), .Y(n1163) );
  AO22X1_HVT U1071 ( .A1(n1028), .A2(n1176), .A3(n1170), .A4(n1029), .Y(n1175)
         );
  AND2X1_HVT U1072 ( .A1(n988), .A2(n1177), .Y(n1170) );
  AND2X1_HVT U1073 ( .A1(n1048), .A2(n1005), .Y(n1173) );
  OA221X1_HVT U1074 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n952), .A5(n1181), .Y(n1161) );
  OA221X1_HVT U1075 ( .A1(n1182), .A2(n953), .A3(n1183), .A4(n1045), .A5(n1184), .Y(n1181) );
  NAND3X0_HVT U1076 ( .A1(n1018), .A2(keyin[114]), .A3(n1117), .Y(n1184) );
  MUX21X1_HVT U1077 ( .A1(n1185), .A2(n1157), .S0(n904), .Y(n1117) );
  OA22X1_HVT U1078 ( .A1(n995), .A2(n1186), .A3(n1187), .A4(n1159), .Y(n1183)
         );
  OA21X1_HVT U1079 ( .A1(keyin[118]), .A2(n1188), .A3(n1189), .Y(n1186) );
  OA222X1_HVT U1080 ( .A1(n1034), .A2(n1188), .A3(n1187), .A4(n1190), .A5(
        n1189), .A6(n1129), .Y(n1182) );
  NAND2X0_HVT U1081 ( .A1(n1038), .A2(n1133), .Y(n1129) );
  INVX0_HVT U1082 ( .A(n1151), .Y(n1034) );
  NAND2X0_HVT U1083 ( .A1(n1039), .A2(n1191), .Y(n1151) );
  OA221X1_HVT U1084 ( .A1(n1192), .A2(n1193), .A3(n1174), .A4(n1188), .A5(
        n1194), .Y(n1180) );
  OA22X1_HVT U1085 ( .A1(n949), .A2(n1187), .A3(n1189), .A4(n1057), .Y(n1194)
         );
  OA221X1_HVT U1086 ( .A1(n1195), .A2(n1189), .A3(n995), .A4(n1187), .A5(n1196), .Y(n1178) );
  OA22X1_HVT U1087 ( .A1(n1188), .A2(n1177), .A3(n1197), .A4(n1192), .Y(n1196)
         );
  INVX0_HVT U1088 ( .A(n987), .Y(n1197) );
  XNOR2X1_HVT U1089 ( .A1(n55), .A2(keyout[74]), .Y(keyout[106]) );
  XOR3X1_HVT U1090 ( .A1(keyin[42]), .A2(keyin[74]), .A3(keyout[10]), .Y(
        keyout[74]) );
  XOR2X1_HVT U1091 ( .A1(keyin[10]), .A2(n1198), .Y(keyout[10]) );
  MUX21X1_HVT U1092 ( .A1(n1199), .A2(n1200), .S0(n572), .Y(n1198) );
  AO221X1_HVT U1093 ( .A1(n1020), .A2(n1201), .A3(n1018), .A4(n1202), .A5(
        n1203), .Y(n1200) );
  AO22X1_HVT U1094 ( .A1(n1013), .A2(n1204), .A3(n1015), .A4(n1205), .Y(n1203)
         );
  OAI221X1_HVT U1095 ( .A1(n1179), .A2(n987), .A3(n949), .A4(n952), .A5(n1206), 
        .Y(n1205) );
  MUX21X1_HVT U1096 ( .A1(n1207), .A2(n1208), .S0(n1108), .Y(n1206) );
  XNOR2X1_HVT U1097 ( .A1(n904), .A2(keyin[118]), .Y(n1108) );
  NAND2X0_HVT U1098 ( .A1(keyin[114]), .A2(n1048), .Y(n1208) );
  NAND2X0_HVT U1099 ( .A1(n1029), .A2(keyin[116]), .Y(n1207) );
  AO222X1_HVT U1100 ( .A1(n1209), .A2(n1139), .A3(n1029), .A4(n1210), .A5(
        n1022), .A6(n1057), .Y(n1204) );
  NAND2X0_HVT U1101 ( .A1(n1058), .A2(n993), .Y(n1210) );
  OAI21X1_HVT U1102 ( .A1(n984), .A2(keyin[114]), .A3(n952), .Y(n1209) );
  AO221X1_HVT U1103 ( .A1(n1025), .A2(n954), .A3(n1031), .A4(n1029), .A5(n1211), .Y(n1202) );
  AO22X1_HVT U1104 ( .A1(n1022), .A2(n1190), .A3(n1028), .A4(n992), .Y(n1211)
         );
  AND2X1_HVT U1105 ( .A1(n1005), .A2(n967), .Y(n1031) );
  AO221X1_HVT U1106 ( .A1(n1029), .A2(n1212), .A3(n1213), .A4(n1022), .A5(
        n1214), .Y(n1201) );
  AO22X1_HVT U1107 ( .A1(n1066), .A2(n1028), .A3(n1025), .A4(n1057), .Y(n1214)
         );
  INVX0_HVT U1108 ( .A(n991), .Y(n1213) );
  NAND2X0_HVT U1109 ( .A1(n1215), .A2(n1072), .Y(n991) );
  NAND2X0_HVT U1110 ( .A1(n1030), .A2(n648), .Y(n1212) );
  AO221X1_HVT U1111 ( .A1(n1015), .A2(n1216), .A3(n1020), .A4(n1217), .A5(
        n1218), .Y(n1199) );
  AO22X1_HVT U1112 ( .A1(n1018), .A2(n1219), .A3(n1013), .A4(n1220), .Y(n1218)
         );
  AO221X1_HVT U1113 ( .A1(n1221), .A2(n1005), .A3(n1025), .A4(n1111), .A5(
        n1222), .Y(n1220) );
  AO22X1_HVT U1114 ( .A1(n1028), .A2(n1223), .A3(n1029), .A4(n1224), .Y(n1222)
         );
  NAND2X0_HVT U1115 ( .A1(n1047), .A2(n1089), .Y(n1224) );
  NAND2X0_HVT U1116 ( .A1(n1191), .A2(n1059), .Y(n1223) );
  NAND2X0_HVT U1117 ( .A1(n995), .A2(n648), .Y(n1059) );
  AO222X1_HVT U1118 ( .A1(n1025), .A2(n1140), .A3(n1225), .A4(n1040), .A5(
        n1028), .A6(n1048), .Y(n1219) );
  AO21X1_HVT U1119 ( .A1(keyin[114]), .A2(n1226), .A3(n1022), .Y(n1225) );
  NAND2X0_HVT U1120 ( .A1(n990), .A2(n1191), .Y(n1226) );
  NAND2X0_HVT U1121 ( .A1(n1048), .A2(n1177), .Y(n1140) );
  AO221X1_HVT U1122 ( .A1(n1227), .A2(n1029), .A3(n1157), .A4(n1028), .A5(
        n1228), .Y(n1217) );
  AO22X1_HVT U1123 ( .A1(n1025), .A2(n967), .A3(n1158), .A4(n1022), .Y(n1228)
         );
  INVX0_HVT U1124 ( .A(n959), .Y(n1158) );
  AND2X1_HVT U1125 ( .A1(n990), .A2(n1046), .Y(n1157) );
  INVX0_HVT U1126 ( .A(n1156), .Y(n1227) );
  NAND2X0_HVT U1127 ( .A1(n967), .A2(n1096), .Y(n1156) );
  AO221X1_HVT U1128 ( .A1(n1035), .A2(n1022), .A3(n1115), .A4(n1025), .A5(
        n1229), .Y(n1216) );
  AO22X1_HVT U1129 ( .A1(n1084), .A2(n1028), .A3(n995), .A4(n1029), .Y(n1229)
         );
  INVX0_HVT U1130 ( .A(n976), .Y(n1084) );
  INVX0_HVT U1131 ( .A(n947), .Y(n1115) );
  NAND2X0_HVT U1132 ( .A1(n993), .A2(n1177), .Y(n947) );
  AND2X1_HVT U1133 ( .A1(n1215), .A2(n990), .Y(n1035) );
  XNOR2X1_HVT U1134 ( .A1(n1230), .A2(keyout[73]), .Y(keyout[105]) );
  XOR3X1_HVT U1135 ( .A1(keyin[41]), .A2(keyin[73]), .A3(keyout[9]), .Y(
        keyout[73]) );
  XOR2X1_HVT U1136 ( .A1(keyin[9]), .A2(n1231), .Y(keyout[9]) );
  MUX21X1_HVT U1137 ( .A1(n1232), .A2(n1233), .S0(n572), .Y(n1231) );
  AO221X1_HVT U1138 ( .A1(n1013), .A2(n1234), .A3(n1020), .A4(n1235), .A5(
        n1236), .Y(n1233) );
  OAI22X1_HVT U1139 ( .A1(n1237), .A2(n1192), .A3(n1238), .A4(n1189), .Y(n1236) );
  OA221X1_HVT U1140 ( .A1(n1045), .A2(n1239), .A3(n1150), .A4(n952), .A5(n1240), .Y(n1238) );
  OA22X1_HVT U1141 ( .A1(n1179), .A2(n1241), .A3(n953), .A4(n1242), .Y(n1240)
         );
  NAND2X0_HVT U1142 ( .A1(n1098), .A2(n1058), .Y(n1241) );
  INVX0_HVT U1143 ( .A(n954), .Y(n1150) );
  OA221X1_HVT U1144 ( .A1(n1045), .A2(n1039), .A3(n952), .A4(n1172), .A5(n1243), .Y(n1237) );
  AOI22X1_HVT U1145 ( .A1(n1088), .A2(n1022), .A3(n1009), .A4(n1028), .Y(n1243) );
  NAND2X0_HVT U1146 ( .A1(n967), .A2(n1244), .Y(n1009) );
  NAND2X0_HVT U1147 ( .A1(n1131), .A2(n1046), .Y(n1088) );
  NAND2X0_HVT U1148 ( .A1(n1245), .A2(n994), .Y(n1172) );
  AO221X1_HVT U1149 ( .A1(n1029), .A2(n1005), .A3(n1028), .A4(n1215), .A5(
        n1246), .Y(n1235) );
  AO22X1_HVT U1150 ( .A1(n1097), .A2(n1022), .A3(n1025), .A4(n1247), .Y(n1246)
         );
  NAND2X0_HVT U1151 ( .A1(n1005), .A2(n990), .Y(n1247) );
  AO221X1_HVT U1152 ( .A1(n1025), .A2(n1248), .A3(n1022), .A4(n1249), .A5(
        n1250), .Y(n1234) );
  AO22X1_HVT U1153 ( .A1(n1185), .A2(n1028), .A3(n1029), .A4(n1111), .Y(n1250)
         );
  NAND2X0_HVT U1154 ( .A1(n1089), .A2(n1039), .Y(n1111) );
  INVX0_HVT U1155 ( .A(n1085), .Y(n1185) );
  NAND2X0_HVT U1156 ( .A1(n1057), .A2(n1177), .Y(n1085) );
  NAND2X0_HVT U1157 ( .A1(keyin[118]), .A2(n1245), .Y(n1177) );
  NAND2X0_HVT U1158 ( .A1(n994), .A2(n1131), .Y(n1248) );
  AO221X1_HVT U1159 ( .A1(n1015), .A2(n1251), .A3(n1018), .A4(n1252), .A5(
        n1253), .Y(n1232) );
  AO22X1_HVT U1160 ( .A1(n1013), .A2(n1254), .A3(n1020), .A4(n1255), .Y(n1253)
         );
  AO222X1_HVT U1161 ( .A1(n1022), .A2(n1176), .A3(n1023), .A4(n1256), .A5(
        n1029), .A6(n1245), .Y(n1255) );
  AO21X1_HVT U1162 ( .A1(n1152), .A2(n837), .A3(n1025), .Y(n1256) );
  INVX0_HVT U1163 ( .A(n1174), .Y(n1023) );
  INVX0_HVT U1164 ( .A(n1249), .Y(n1176) );
  NAND2X0_HVT U1165 ( .A1(n1096), .A2(n1041), .Y(n1249) );
  AO221X1_HVT U1166 ( .A1(n1025), .A2(n1047), .A3(n1257), .A4(n1022), .A5(
        n1258), .Y(n1254) );
  OAI22X1_HVT U1167 ( .A1(n1179), .A2(n757), .A3(n1065), .A4(n1045), .Y(n1258)
         );
  NAND2X0_HVT U1168 ( .A1(n976), .A2(n1046), .Y(n1065) );
  INVX0_HVT U1169 ( .A(n1259), .Y(n1257) );
  AO221X1_HVT U1170 ( .A1(n1025), .A2(n959), .A3(n1260), .A4(n1028), .A5(n1261), .Y(n1252) );
  AO22X1_HVT U1171 ( .A1(n1022), .A2(n1109), .A3(n1029), .A4(n1262), .Y(n1261)
         );
  NAND2X0_HVT U1172 ( .A1(n1133), .A2(n1191), .Y(n1262) );
  NAND2X0_HVT U1173 ( .A1(n1040), .A2(n1072), .Y(n959) );
  AO221X1_HVT U1174 ( .A1(n1029), .A2(n1215), .A3(n1028), .A4(n1190), .A5(
        n1263), .Y(n1251) );
  AO21X1_HVT U1175 ( .A1(n1118), .A2(n904), .A3(n1135), .Y(n1263) );
  INVX0_HVT U1176 ( .A(n973), .Y(n1135) );
  NAND2X0_HVT U1177 ( .A1(n1025), .A2(n648), .Y(n973) );
  NAND2X0_HVT U1178 ( .A1(n1046), .A2(n1039), .Y(n1118) );
  XNOR2X1_HVT U1179 ( .A1(n209), .A2(keyout[72]), .Y(keyout[104]) );
  XOR3X1_HVT U1180 ( .A1(keyin[40]), .A2(keyin[72]), .A3(keyout[8]), .Y(
        keyout[72]) );
  XOR2X1_HVT U1181 ( .A1(keyin[8]), .A2(n1264), .Y(keyout[8]) );
  MUX21X1_HVT U1182 ( .A1(n1265), .A2(n1266), .S0(n572), .Y(n1264) );
  INVX0_HVT U1183 ( .A(keyin[119]), .Y(n572) );
  AO221X1_HVT U1184 ( .A1(n1013), .A2(n1267), .A3(n1018), .A4(n1268), .A5(
        n1269), .Y(n1266) );
  AO22X1_HVT U1185 ( .A1(n1020), .A2(n1270), .A3(n1015), .A4(n1271), .Y(n1269)
         );
  AO221X1_HVT U1186 ( .A1(n1029), .A2(n1272), .A3(n1066), .A4(n1022), .A5(
        n1273), .Y(n1271) );
  AO22X1_HVT U1187 ( .A1(n1274), .A2(n837), .A3(n1027), .A4(n1028), .Y(n1273)
         );
  AND2X1_HVT U1188 ( .A1(n992), .A2(n1131), .Y(n1027) );
  INVX0_HVT U1189 ( .A(n1040), .Y(n1274) );
  INVX0_HVT U1190 ( .A(n1094), .Y(n1066) );
  NAND2X0_HVT U1191 ( .A1(n987), .A2(n1064), .Y(n1094) );
  NAND2X0_HVT U1192 ( .A1(n1057), .A2(n648), .Y(n1064) );
  NAND2X0_HVT U1193 ( .A1(n1215), .A2(n967), .Y(n1272) );
  OAI221X1_HVT U1194 ( .A1(n1152), .A2(n1045), .A3(n1242), .A4(n1179), .A5(
        n1275), .Y(n1270) );
  OA22X1_HVT U1195 ( .A1(n952), .A2(n1109), .A3(n953), .A4(n982), .Y(n1275) );
  AND2X1_HVT U1196 ( .A1(n1245), .A2(n1058), .Y(n982) );
  NAND2X0_HVT U1197 ( .A1(n1005), .A2(n1072), .Y(n1242) );
  NAND2X0_HVT U1198 ( .A1(keyin[118]), .A2(n993), .Y(n1005) );
  NAND2X0_HVT U1199 ( .A1(n1047), .A2(n987), .Y(n1152) );
  AO221X1_HVT U1200 ( .A1(n1029), .A2(n993), .A3(n1260), .A4(n1028), .A5(n1276), .Y(n1268) );
  AO21X1_HVT U1201 ( .A1(n1001), .A2(n1025), .A3(n1221), .Y(n1276) );
  INVX0_HVT U1202 ( .A(n1043), .Y(n1221) );
  NAND2X0_HVT U1203 ( .A1(n1022), .A2(n949), .Y(n1043) );
  INVX0_HVT U1204 ( .A(n1244), .Y(n1001) );
  INVX0_HVT U1205 ( .A(n1239), .Y(n1260) );
  NAND2X0_HVT U1206 ( .A1(n1058), .A2(n1072), .Y(n1239) );
  AO221X1_HVT U1207 ( .A1(n1022), .A2(n954), .A3(n1025), .A4(n994), .A5(n1277), 
        .Y(n1267) );
  AO22X1_HVT U1208 ( .A1(n1112), .A2(n1028), .A3(n1029), .A4(n1174), .Y(n1277)
         );
  NAND2X0_HVT U1209 ( .A1(n1244), .A2(n984), .Y(n1174) );
  INVX0_HVT U1210 ( .A(n1139), .Y(n1112) );
  NAND2X0_HVT U1211 ( .A1(n1058), .A2(n1131), .Y(n1139) );
  NAND2X0_HVT U1212 ( .A1(n993), .A2(n648), .Y(n1131) );
  NAND2X0_HVT U1213 ( .A1(n993), .A2(n1215), .Y(n954) );
  NAND2X0_HVT U1214 ( .A1(keyin[118]), .A2(n949), .Y(n1215) );
  AO221X1_HVT U1215 ( .A1(n1020), .A2(n1278), .A3(n1018), .A4(n1279), .A5(
        n1280), .Y(n1265) );
  AO22X1_HVT U1216 ( .A1(n1015), .A2(n1281), .A3(n1013), .A4(n1282), .Y(n1280)
         );
  NAND3X0_HVT U1217 ( .A1(n1283), .A2(n1284), .A3(n1285), .Y(n1282) );
  AOI22X1_HVT U1218 ( .A1(n961), .A2(n1022), .A3(n1159), .A4(n1028), .Y(n1285)
         );
  NAND2X0_HVT U1219 ( .A1(n1133), .A2(n1046), .Y(n1159) );
  NAND2X0_HVT U1220 ( .A1(keyin[118]), .A2(keyin[115]), .Y(n1046) );
  NAND2X0_HVT U1221 ( .A1(n971), .A2(n648), .Y(n1133) );
  NAND2X0_HVT U1222 ( .A1(n987), .A2(n984), .Y(n961) );
  NAND3X0_HVT U1223 ( .A1(n1098), .A2(n1058), .A3(n1029), .Y(n1284) );
  NAND2X0_HVT U1224 ( .A1(keyin[118]), .A2(n1057), .Y(n1058) );
  AO21X1_HVT U1225 ( .A1(n994), .A2(n1041), .A3(n952), .Y(n1283) );
  NAND2X0_HVT U1226 ( .A1(keyin[116]), .A2(n648), .Y(n1041) );
  NAND2X0_HVT U1227 ( .A1(keyin[118]), .A2(n1048), .Y(n994) );
  INVX0_HVT U1228 ( .A(n1187), .Y(n1013) );
  NAND2X0_HVT U1229 ( .A1(keyin[117]), .A2(n870), .Y(n1187) );
  AO221X1_HVT U1230 ( .A1(n1286), .A2(n1025), .A3(n1028), .A4(n1057), .A5(
        n1287), .Y(n1281) );
  AO22X1_HVT U1231 ( .A1(n1022), .A2(n976), .A3(n1029), .A4(n1288), .Y(n1287)
         );
  NAND2X0_HVT U1232 ( .A1(n990), .A2(n1038), .Y(n1288) );
  NAND2X0_HVT U1233 ( .A1(keyin[118]), .A2(n1109), .Y(n1038) );
  NAND2X0_HVT U1234 ( .A1(n757), .A2(n648), .Y(n990) );
  NAND2X0_HVT U1235 ( .A1(n648), .A2(n1109), .Y(n976) );
  INVX0_HVT U1236 ( .A(n1193), .Y(n1286) );
  NAND2X0_HVT U1237 ( .A1(n1040), .A2(n1039), .Y(n1193) );
  NAND2X0_HVT U1238 ( .A1(n949), .A2(n648), .Y(n1039) );
  NAND2X0_HVT U1239 ( .A1(n995), .A2(keyin[118]), .Y(n1040) );
  INVX0_HVT U1240 ( .A(n1057), .Y(n995) );
  NAND2X0_HVT U1241 ( .A1(keyin[115]), .A2(n757), .Y(n1057) );
  INVX0_HVT U1242 ( .A(n1189), .Y(n1015) );
  NAND2X0_HVT U1243 ( .A1(keyin[113]), .A2(keyin[117]), .Y(n1189) );
  AO221X1_HVT U1244 ( .A1(n1025), .A2(n1259), .A3(n1028), .A4(n1063), .A5(
        n1289), .Y(n1279) );
  AO222X1_HVT U1245 ( .A1(n1022), .A2(n1244), .A3(n1097), .A4(n1029), .A5(n951), .A6(keyin[114]), .Y(n1289) );
  INVX0_HVT U1246 ( .A(n988), .Y(n951) );
  INVX0_HVT U1247 ( .A(n1045), .Y(n1029) );
  NAND2X0_HVT U1248 ( .A1(keyin[112]), .A2(keyin[114]), .Y(n1045) );
  INVX0_HVT U1249 ( .A(n1191), .Y(n1097) );
  NAND2X0_HVT U1250 ( .A1(n1030), .A2(keyin[118]), .Y(n1191) );
  INVX0_HVT U1251 ( .A(n1048), .Y(n1030) );
  NAND2X0_HVT U1252 ( .A1(keyin[118]), .A2(keyin[116]), .Y(n1244) );
  INVX0_HVT U1253 ( .A(n1195), .Y(n1063) );
  OA21X1_HVT U1254 ( .A1(n1048), .A2(keyin[118]), .A3(n992), .Y(n1195) );
  NAND2X0_HVT U1255 ( .A1(n988), .A2(n1089), .Y(n1259) );
  NAND2X0_HVT U1256 ( .A1(keyin[118]), .A2(n1098), .Y(n1089) );
  NAND2X0_HVT U1257 ( .A1(n1048), .A2(n648), .Y(n988) );
  NAND2X0_HVT U1258 ( .A1(keyin[116]), .A2(n1109), .Y(n1048) );
  INVX0_HVT U1259 ( .A(n1192), .Y(n1018) );
  NAND2X0_HVT U1260 ( .A1(keyin[113]), .A2(n712), .Y(n1192) );
  AO222X1_HVT U1261 ( .A1(n1290), .A2(n1291), .A3(n1028), .A4(n1292), .A5(
        n1025), .A6(n1143), .Y(n1278) );
  NAND2X0_HVT U1262 ( .A1(n1072), .A2(n992), .Y(n1143) );
  NAND2X0_HVT U1263 ( .A1(keyin[115]), .A2(n648), .Y(n1072) );
  INVX0_HVT U1264 ( .A(n952), .Y(n1025) );
  NAND2X0_HVT U1265 ( .A1(n904), .A2(n837), .Y(n952) );
  NAND2X0_HVT U1266 ( .A1(n967), .A2(n987), .Y(n1292) );
  NAND2X0_HVT U1267 ( .A1(keyin[118]), .A2(n757), .Y(n987) );
  NAND2X0_HVT U1268 ( .A1(n648), .A2(n1245), .Y(n967) );
  INVX0_HVT U1269 ( .A(n1179), .Y(n1028) );
  NAND2X0_HVT U1270 ( .A1(keyin[112]), .A2(n837), .Y(n1179) );
  INVX0_HVT U1271 ( .A(keyin[114]), .Y(n837) );
  AO21X1_HVT U1272 ( .A1(keyin[114]), .A2(n1006), .A3(n1022), .Y(n1291) );
  INVX0_HVT U1273 ( .A(n953), .Y(n1022) );
  NAND2X0_HVT U1274 ( .A1(keyin[114]), .A2(n904), .Y(n953) );
  INVX0_HVT U1275 ( .A(keyin[112]), .Y(n904) );
  NAND2X0_HVT U1276 ( .A1(n992), .A2(n984), .Y(n1006) );
  NAND2X0_HVT U1277 ( .A1(n1098), .A2(n648), .Y(n984) );
  INVX0_HVT U1278 ( .A(n949), .Y(n1098) );
  NAND2X0_HVT U1279 ( .A1(n1245), .A2(n993), .Y(n949) );
  NAND2X0_HVT U1280 ( .A1(n1068), .A2(keyin[118]), .Y(n992) );
  INVX0_HVT U1281 ( .A(n1190), .Y(n1290) );
  NAND2X0_HVT U1282 ( .A1(n1047), .A2(n1096), .Y(n1190) );
  NAND2X0_HVT U1283 ( .A1(n971), .A2(keyin[118]), .Y(n1096) );
  INVX0_HVT U1284 ( .A(n1245), .Y(n971) );
  NAND2X0_HVT U1285 ( .A1(n757), .A2(n1109), .Y(n1245) );
  INVX0_HVT U1286 ( .A(keyin[115]), .Y(n1109) );
  INVX0_HVT U1287 ( .A(keyin[116]), .Y(n757) );
  NAND2X0_HVT U1288 ( .A1(n1068), .A2(n648), .Y(n1047) );
  INVX0_HVT U1289 ( .A(keyin[118]), .Y(n648) );
  INVX0_HVT U1290 ( .A(n993), .Y(n1068) );
  NAND2X0_HVT U1291 ( .A1(keyin[116]), .A2(keyin[115]), .Y(n993) );
  INVX0_HVT U1292 ( .A(n1188), .Y(n1020) );
  NAND2X0_HVT U1293 ( .A1(n870), .A2(n712), .Y(n1188) );
  INVX0_HVT U1294 ( .A(keyin[117]), .Y(n712) );
  INVX0_HVT U1295 ( .A(keyin[113]), .Y(n870) );
  XNOR2X1_HVT U1296 ( .A1(keyout[71]), .A2(n217), .Y(keyout[103]) );
  INVX0_HVT U1297 ( .A(keyin[103]), .Y(n217) );
  XOR2X1_HVT U1298 ( .A1(keyout[39]), .A2(keyin[71]), .Y(keyout[71]) );
  XOR2X1_HVT U1299 ( .A1(keyout[7]), .A2(keyin[39]), .Y(keyout[39]) );
  XNOR3X1_HVT U1300 ( .A1(n90), .A2(keyin[7]), .A3(n1293), .Y(keyout[7]) );
  AO221X1_HVT U1301 ( .A1(n1294), .A2(n1295), .A3(n1296), .A4(n1297), .A5(
        n1298), .Y(n1293) );
  AO22X1_HVT U1302 ( .A1(n1299), .A2(n1300), .A3(n1301), .A4(n1302), .Y(n1298)
         );
  AO221X1_HVT U1303 ( .A1(n1303), .A2(n86), .A3(n1304), .A4(n1305), .A5(n1306), 
        .Y(n1302) );
  AO221X1_HVT U1304 ( .A1(n1307), .A2(n44), .A3(n1308), .A4(n1309), .A5(n1310), 
        .Y(n1306) );
  AND3X1_HVT U1305 ( .A1(n1311), .A2(n209), .A3(n1312), .Y(n1310) );
  NAND2X0_HVT U1306 ( .A1(keyin[109]), .A2(n37), .Y(n1312) );
  INVX0_HVT U1307 ( .A(n1313), .Y(n1311) );
  AO21X1_HVT U1308 ( .A1(keyin[109]), .A2(n1314), .A3(n1315), .Y(n1307) );
  AO22X1_HVT U1309 ( .A1(keyin[108]), .A2(keyin[106]), .A3(n1316), .A4(
        keyin[104]), .Y(n1314) );
  INVX0_HVT U1310 ( .A(n176), .Y(n1305) );
  NAND4X0_HVT U1311 ( .A1(n1317), .A2(n1318), .A3(n1319), .A4(n1320), .Y(n1300) );
  OA221X1_HVT U1312 ( .A1(n1321), .A2(n1322), .A3(n117), .A4(n1323), .A5(n1324), .Y(n1320) );
  OA22X1_HVT U1313 ( .A1(n1325), .A2(n1326), .A3(n1327), .A4(n1328), .Y(n1324)
         );
  OA22X1_HVT U1314 ( .A1(n1329), .A2(n145), .A3(n127), .A4(n1330), .Y(n1319)
         );
  NAND2X0_HVT U1315 ( .A1(n179), .A2(n1331), .Y(n127) );
  AO21X1_HVT U1316 ( .A1(n145), .A2(n122), .A3(n1332), .Y(n1318) );
  AO21X1_HVT U1317 ( .A1(n116), .A2(n177), .A3(n1333), .Y(n1317) );
  NAND3X0_HVT U1318 ( .A1(n1334), .A2(n1335), .A3(n1336), .Y(n1297) );
  OA222X1_HVT U1319 ( .A1(n199), .A2(n1333), .A3(n1327), .A4(n149), .A5(n1332), 
        .A6(n1337), .Y(n1336) );
  OA22X1_HVT U1320 ( .A1(n1330), .A2(n1338), .A3(keyin[109]), .A4(n1339), .Y(
        n1335) );
  OA221X1_HVT U1321 ( .A1(n1316), .A2(n108), .A3(n1340), .A4(n42), .A5(n1341), 
        .Y(n1339) );
  AOI22X1_HVT U1322 ( .A1(n1328), .A2(n1342), .A3(n1343), .A4(n1303), .Y(n1334) );
  NAND2X0_HVT U1323 ( .A1(n81), .A2(n61), .Y(n1328) );
  NAND2X0_HVT U1324 ( .A1(n1344), .A2(n1345), .Y(n1295) );
  OA222X1_HVT U1325 ( .A1(n1346), .A2(n1330), .A3(n1347), .A4(n107), .A5(
        keyin[109]), .A6(n1348), .Y(n1345) );
  OA22X1_HVT U1326 ( .A1(n1349), .A2(n108), .A3(n42), .A4(n118), .Y(n1348) );
  OA21X1_HVT U1327 ( .A1(n51), .A2(n1333), .A3(n1332), .Y(n1347) );
  OA222X1_HVT U1328 ( .A1(n202), .A2(n1327), .A3(n1322), .A4(n1350), .A5(n1325), .A6(n1351), .Y(n1344) );
  XNOR3X1_HVT U1329 ( .A1(keyin[70]), .A2(n427), .A3(keyout[38]), .Y(
        keyout[102]) );
  XNOR3X1_HVT U1330 ( .A1(n7), .A2(keyin[38]), .A3(n6), .Y(keyout[38]) );
  XNOR2X1_HVT U1331 ( .A1(keyin[6]), .A2(n1352), .Y(n6) );
  MUX21X1_HVT U1332 ( .A1(n1353), .A2(n1354), .S0(n26), .Y(n1352) );
  AO221X1_HVT U1333 ( .A1(n34), .A2(n1355), .A3(n29), .A4(n1356), .A5(n1357), 
        .Y(n1354) );
  AO22X1_HVT U1334 ( .A1(n27), .A2(n1358), .A3(n32), .A4(n1359), .Y(n1357) );
  AO221X1_HVT U1335 ( .A1(n83), .A2(n46), .A3(n1360), .A4(n36), .A5(n1361), 
        .Y(n1359) );
  AO22X1_HVT U1336 ( .A1(n1362), .A2(n40), .A3(n52), .A4(n1350), .Y(n1361) );
  INVX0_HVT U1337 ( .A(n58), .Y(n83) );
  AO221X1_HVT U1338 ( .A1(n45), .A2(n52), .A3(n119), .A4(n40), .A5(n1363), .Y(
        n1358) );
  AO22X1_HVT U1339 ( .A1(n36), .A2(n176), .A3(n50), .A4(n46), .Y(n1363) );
  INVX0_HVT U1340 ( .A(n115), .Y(n50) );
  AO221X1_HVT U1341 ( .A1(n1364), .A2(n52), .A3(n152), .A4(n40), .A5(n1365), 
        .Y(n1356) );
  AO22X1_HVT U1342 ( .A1(n1360), .A2(n46), .A3(n36), .A4(n1366), .Y(n1365) );
  NAND2X0_HVT U1343 ( .A1(n1367), .A2(n173), .Y(n1366) );
  AND2X1_HVT U1344 ( .A1(n143), .A2(n196), .Y(n1360) );
  AND2X1_HVT U1345 ( .A1(n179), .A2(n145), .Y(n152) );
  INVX0_HVT U1346 ( .A(n73), .Y(n1364) );
  NAND3X0_HVT U1347 ( .A1(n1368), .A2(n1369), .A3(n1370), .Y(n1355) );
  OA22X1_HVT U1348 ( .A1(n1340), .A2(n108), .A3(n167), .A4(n1371), .Y(n1370)
         );
  INVX0_HVT U1349 ( .A(n138), .Y(n1340) );
  NAND3X0_HVT U1350 ( .A1(n37), .A2(n63), .A3(n40), .Y(n1368) );
  AO221X1_HVT U1351 ( .A1(n34), .A2(n1372), .A3(n29), .A4(n1373), .A5(n1374), 
        .Y(n1353) );
  AO22X1_HVT U1352 ( .A1(n27), .A2(n1375), .A3(n32), .A4(n1376), .Y(n1374) );
  AO221X1_HVT U1353 ( .A1(n36), .A2(n1377), .A3(n1378), .A4(n40), .A5(n1379), 
        .Y(n1376) );
  AO22X1_HVT U1354 ( .A1(n52), .A2(n77), .A3(n46), .A4(n1337), .Y(n1379) );
  INVX0_HVT U1355 ( .A(n196), .Y(n1378) );
  NAND2X0_HVT U1356 ( .A1(n115), .A2(n140), .Y(n1377) );
  AO221X1_HVT U1357 ( .A1(n36), .A2(n1380), .A3(n40), .A4(n1381), .A5(n1382), 
        .Y(n1375) );
  MUX21X1_HVT U1358 ( .A1(n46), .A2(n52), .S0(n79), .Y(n1382) );
  NAND2X0_HVT U1359 ( .A1(n77), .A2(n37), .Y(n1381) );
  NAND2X0_HVT U1360 ( .A1(n1367), .A2(n1383), .Y(n1380) );
  AO221X1_HVT U1361 ( .A1(n36), .A2(n200), .A3(n126), .A4(n52), .A5(n1384), 
        .Y(n1373) );
  AO22X1_HVT U1362 ( .A1(n46), .A2(n1385), .A3(n40), .A4(n196), .Y(n1384) );
  NAND2X0_HVT U1363 ( .A1(n1343), .A2(n1371), .Y(n200) );
  AO222X1_HVT U1364 ( .A1(n1386), .A2(n36), .A3(n1387), .A4(n1388), .A5(n40), 
        .A6(n1351), .Y(n1372) );
  OAI21X1_HVT U1365 ( .A1(n173), .A2(n55), .A3(n42), .Y(n1388) );
  AND2X1_HVT U1366 ( .A1(n115), .A2(n63), .Y(n1387) );
  INVX0_HVT U1367 ( .A(n1337), .Y(n1386) );
  NAND2X0_HVT U1368 ( .A1(n177), .A2(n1331), .Y(n1337) );
  AO21X1_HVT U1369 ( .A1(n1389), .A2(round_num[0]), .A3(n1390), .Y(n7) );
  INVX0_HVT U1370 ( .A(keyin[102]), .Y(n427) );
  XNOR3X1_HVT U1371 ( .A1(keyin[69]), .A2(n264), .A3(keyout[37]), .Y(
        keyout[101]) );
  XNOR3X1_HVT U1372 ( .A1(n15), .A2(keyin[37]), .A3(n16), .Y(keyout[37]) );
  XNOR2X1_HVT U1373 ( .A1(n1391), .A2(keyin[5]), .Y(n16) );
  AO221X1_HVT U1374 ( .A1(n1294), .A2(n1392), .A3(n1296), .A4(n1393), .A5(
        n1394), .Y(n1391) );
  AO22X1_HVT U1375 ( .A1(n1299), .A2(n1395), .A3(n1301), .A4(n1396), .Y(n1394)
         );
  NAND4X0_HVT U1376 ( .A1(n1397), .A2(n1398), .A3(n1399), .A4(n1400), .Y(n1396) );
  OA221X1_HVT U1377 ( .A1(n155), .A2(n1332), .A3(n1401), .A4(n1327), .A5(n1402), .Y(n1400) );
  OA22X1_HVT U1378 ( .A1(n176), .A2(n1322), .A3(n1325), .A4(n47), .Y(n1402) );
  NAND2X0_HVT U1379 ( .A1(n1343), .A2(n195), .Y(n47) );
  NAND2X0_HVT U1380 ( .A1(n149), .A2(n1403), .Y(n176) );
  OA22X1_HVT U1381 ( .A1(n1329), .A2(n175), .A3(n51), .A4(n1323), .Y(n1399) );
  INVX0_HVT U1382 ( .A(n177), .Y(n51) );
  AO21X1_HVT U1383 ( .A1(n81), .A2(n196), .A3(n1330), .Y(n1398) );
  AO21X1_HVT U1384 ( .A1(n137), .A2(n1383), .A3(n1333), .Y(n1397) );
  NAND4X0_HVT U1385 ( .A1(n1404), .A2(n1405), .A3(n1406), .A4(n1407), .Y(n1395) );
  OA222X1_HVT U1386 ( .A1(n44), .A2(n1333), .A3(n1323), .A4(n196), .A5(n1408), 
        .A6(n1325), .Y(n1407) );
  OA22X1_HVT U1387 ( .A1(n1409), .A2(n1332), .A3(n115), .A4(n1329), .Y(n1406)
         );
  AND2X1_HVT U1388 ( .A1(n195), .A2(n117), .Y(n1409) );
  NAND3X0_HVT U1389 ( .A1(keyin[109]), .A2(n209), .A3(n181), .Y(n1405) );
  AO21X1_HVT U1390 ( .A1(n87), .A2(n177), .A3(n1327), .Y(n1404) );
  NAND4X0_HVT U1391 ( .A1(n1410), .A2(n1411), .A3(n1412), .A4(n1413), .Y(n1393) );
  OA221X1_HVT U1392 ( .A1(n119), .A2(n1333), .A3(n115), .A4(n1332), .A5(n1414), 
        .Y(n1413) );
  MUX21X1_HVT U1393 ( .A1(n1415), .A2(n143), .S0(n1073), .Y(n1414) );
  OA21X1_HVT U1394 ( .A1(n55), .A2(n149), .A3(n1416), .Y(n1415) );
  MUX21X1_HVT U1395 ( .A1(n1417), .A2(n1418), .S0(n112), .Y(n1416) );
  NAND2X0_HVT U1396 ( .A1(n36), .A2(keyin[108]), .Y(n1418) );
  NAND2X0_HVT U1397 ( .A1(n63), .A2(n55), .Y(n1417) );
  AND2X1_HVT U1398 ( .A1(n149), .A2(n37), .Y(n119) );
  OA22X1_HVT U1399 ( .A1(n1309), .A2(n1322), .A3(n1325), .A4(n1338), .Y(n1412)
         );
  NAND2X0_HVT U1400 ( .A1(n61), .A2(n1367), .Y(n1338) );
  NAND3X0_HVT U1401 ( .A1(n112), .A2(n205), .A3(n1308), .Y(n1411) );
  XNOR2X1_HVT U1402 ( .A1(n209), .A2(keyin[110]), .Y(n112) );
  NAND2X0_HVT U1403 ( .A1(n1419), .A2(n41), .Y(n1410) );
  NAND2X0_HVT U1404 ( .A1(n137), .A2(n173), .Y(n41) );
  INVX0_HVT U1405 ( .A(n1323), .Y(n1419) );
  AO221X1_HVT U1406 ( .A1(n1342), .A2(n1351), .A3(n1303), .A4(n1420), .A5(
        n1421), .Y(n1392) );
  AO222X1_HVT U1407 ( .A1(n1422), .A2(n55), .A3(n153), .A4(n1423), .A5(n1304), 
        .A6(n140), .Y(n1421) );
  NAND2X0_HVT U1408 ( .A1(n1332), .A2(n1323), .Y(n1423) );
  INVX0_HVT U1409 ( .A(n1346), .Y(n153) );
  NAND2X0_HVT U1410 ( .A1(n116), .A2(n62), .Y(n1346) );
  MUX21X1_HVT U1411 ( .A1(n70), .A2(n208), .S0(n1073), .Y(n1422) );
  NAND2X0_HVT U1412 ( .A1(n1371), .A2(n173), .Y(n208) );
  MUX21X1_HVT U1413 ( .A1(n186), .A2(n147), .S0(n209), .Y(n70) );
  INVX0_HVT U1414 ( .A(n1401), .Y(n186) );
  NAND2X0_HVT U1415 ( .A1(n77), .A2(n62), .Y(n1401) );
  INVX0_HVT U1416 ( .A(n1325), .Y(n1303) );
  NAND2X0_HVT U1417 ( .A1(n115), .A2(n61), .Y(n1351) );
  AO21X1_HVT U1418 ( .A1(n156), .A2(n1424), .A3(n97), .Y(n15) );
  INVX0_HVT U1419 ( .A(n89), .Y(n97) );
  NAND2X0_HVT U1420 ( .A1(round_num[0]), .A2(n1390), .Y(n89) );
  AND3X1_HVT U1421 ( .A1(n1424), .A2(n1425), .A3(round_num[2]), .Y(n1390) );
  AND3X1_HVT U1422 ( .A1(round_num[2]), .A2(n92), .A3(round_num[3]), .Y(n156)
         );
  INVX0_HVT U1423 ( .A(keyin[101]), .Y(n264) );
  XNOR2X1_HVT U1424 ( .A1(n313), .A2(keyout[68]), .Y(keyout[100]) );
  XOR2X1_HVT U1425 ( .A1(keyout[36]), .A2(keyin[68]), .Y(keyout[68]) );
  XNOR3X1_HVT U1426 ( .A1(n18), .A2(keyin[36]), .A3(n19), .Y(keyout[36]) );
  XNOR2X1_HVT U1427 ( .A1(n1426), .A2(keyin[4]), .Y(n19) );
  AO221X1_HVT U1428 ( .A1(n1301), .A2(n1427), .A3(n1299), .A4(n1428), .A5(
        n1429), .Y(n1426) );
  AO22X1_HVT U1429 ( .A1(n1296), .A2(n1430), .A3(n1294), .A4(n1431), .Y(n1429)
         );
  NAND4X0_HVT U1430 ( .A1(n1432), .A2(n1433), .A3(n1434), .A4(n1435), .Y(n1431) );
  OA221X1_HVT U1431 ( .A1(n1313), .A2(n1333), .A3(n74), .A4(n1327), .A5(n1436), 
        .Y(n1435) );
  AOI22X1_HVT U1432 ( .A1(n187), .A2(n1315), .A3(n155), .A4(n1342), .Y(n1436)
         );
  INVX0_HVT U1433 ( .A(n1343), .Y(n155) );
  INVX0_HVT U1434 ( .A(n1332), .Y(n1315) );
  NAND2X0_HVT U1435 ( .A1(n1367), .A2(n53), .Y(n74) );
  OA22X1_HVT U1436 ( .A1(n1437), .A2(n1329), .A3(n1323), .A4(n53), .Y(n1434)
         );
  INVX0_HVT U1437 ( .A(n149), .Y(n1437) );
  NAND3X0_HVT U1438 ( .A1(n1438), .A2(n199), .A3(keyin[109]), .Y(n1433) );
  AO21X1_HVT U1439 ( .A1(keyin[106]), .A2(keyin[110]), .A3(n210), .Y(n1438) );
  INVX0_HVT U1440 ( .A(n1341), .Y(n210) );
  NAND2X0_HVT U1441 ( .A1(n36), .A2(n44), .Y(n1341) );
  AO21X1_HVT U1442 ( .A1(n77), .A2(n177), .A3(n1325), .Y(n1432) );
  AND2X1_HVT U1443 ( .A1(keyin[111]), .A2(n1230), .Y(n1294) );
  NAND3X0_HVT U1444 ( .A1(n1439), .A2(n1440), .A3(n1441), .Y(n1430) );
  AOI222X1_HVT U1445 ( .A1(n39), .A2(n1304), .A3(n141), .A4(n1308), .A5(n177), 
        .A6(n1342), .Y(n1441) );
  INVX0_HVT U1446 ( .A(n1322), .Y(n1342) );
  INVX0_HVT U1447 ( .A(n1327), .Y(n1308) );
  NAND2X0_HVT U1448 ( .A1(n63), .A2(n62), .Y(n141) );
  NAND2X0_HVT U1449 ( .A1(keyin[110]), .A2(n178), .Y(n62) );
  INVX0_HVT U1450 ( .A(n1333), .Y(n1304) );
  AO21X1_HVT U1451 ( .A1(n1325), .A2(n1442), .A3(n1326), .Y(n1440) );
  NAND2X0_HVT U1452 ( .A1(n195), .A2(n140), .Y(n1326) );
  NAND2X0_HVT U1453 ( .A1(n86), .A2(n44), .Y(n140) );
  AO21X1_HVT U1454 ( .A1(n137), .A2(n53), .A3(n167), .Y(n1442) );
  OA22X1_HVT U1455 ( .A1(n108), .A2(n1443), .A3(n1323), .A4(n56), .Y(n1439) );
  MUX21X1_HVT U1456 ( .A1(n1444), .A2(n45), .S0(n1445), .Y(n1443) );
  XNOR2X1_HVT U1457 ( .A1(n44), .A2(keyin[109]), .Y(n1445) );
  MUX21X1_HVT U1458 ( .A1(n205), .A2(n199), .S0(n1073), .Y(n1444) );
  AND2X1_HVT U1459 ( .A1(keyin[111]), .A2(keyin[105]), .Y(n1296) );
  NAND4X0_HVT U1460 ( .A1(n1446), .A2(n1447), .A3(n1448), .A4(n1449), .Y(n1428) );
  OA22X1_HVT U1461 ( .A1(n86), .A2(n1330), .A3(n169), .A4(n1323), .Y(n1449) );
  NAND2X0_HVT U1462 ( .A1(n46), .A2(n1073), .Y(n1323) );
  INVX0_HVT U1463 ( .A(n118), .Y(n169) );
  OA22X1_HVT U1464 ( .A1(n1322), .A2(n137), .A3(n1325), .A4(n73), .Y(n1448) );
  NAND2X0_HVT U1465 ( .A1(n173), .A2(n139), .Y(n73) );
  OA22X1_HVT U1466 ( .A1(n194), .A2(n1327), .A3(n1420), .A4(n1332), .Y(n1447)
         );
  OA22X1_HVT U1467 ( .A1(n1343), .A2(n1333), .A3(n87), .A4(n108), .Y(n1446) );
  AND2X1_HVT U1468 ( .A1(keyin[105]), .A2(n26), .Y(n1299) );
  NAND3X0_HVT U1469 ( .A1(n1450), .A2(n1451), .A3(n1452), .Y(n1427) );
  OA222X1_HVT U1470 ( .A1(n151), .A2(n1333), .A3(n1327), .A4(n1350), .A5(n147), 
        .A6(n1332), .Y(n1452) );
  NAND2X0_HVT U1471 ( .A1(n52), .A2(keyin[109]), .Y(n1332) );
  AND2X1_HVT U1472 ( .A1(n145), .A2(n1371), .Y(n147) );
  NAND2X0_HVT U1473 ( .A1(n40), .A2(keyin[109]), .Y(n1327) );
  NAND2X0_HVT U1474 ( .A1(n40), .A2(n1073), .Y(n1333) );
  NAND2X0_HVT U1475 ( .A1(n149), .A2(n195), .Y(n151) );
  OA22X1_HVT U1476 ( .A1(n150), .A2(n1329), .A3(n78), .A4(n1330), .Y(n1451) );
  NAND2X0_HVT U1477 ( .A1(n36), .A2(keyin[109]), .Y(n1330) );
  NAND2X0_HVT U1478 ( .A1(n36), .A2(n1073), .Y(n1329) );
  INVX0_HVT U1479 ( .A(n202), .Y(n150) );
  NAND2X0_HVT U1480 ( .A1(n143), .A2(n1331), .Y(n202) );
  OA22X1_HVT U1481 ( .A1(n1322), .A2(n1331), .A3(n1325), .A4(n175), .Y(n1450)
         );
  NAND2X0_HVT U1482 ( .A1(n187), .A2(n1371), .Y(n175) );
  NAND2X0_HVT U1483 ( .A1(n52), .A2(n1073), .Y(n1325) );
  NAND2X0_HVT U1484 ( .A1(n46), .A2(keyin[109]), .Y(n1322) );
  AND2X1_HVT U1485 ( .A1(n1230), .A2(n26), .Y(n1301) );
  AO22X1_HVT U1486 ( .A1(n1389), .A2(round_num[0]), .A3(n96), .A4(n93), .Y(n18) );
  AND3X1_HVT U1487 ( .A1(n92), .A2(n1425), .A3(round_num[1]), .Y(n96) );
  INVX0_HVT U1488 ( .A(round_num[0]), .Y(n92) );
  INVX0_HVT U1489 ( .A(n90), .Y(n1389) );
  NAND3X0_HVT U1490 ( .A1(n1424), .A2(n93), .A3(round_num[3]), .Y(n90) );
  INVX0_HVT U1491 ( .A(keyin[100]), .Y(n313) );
  XOR2X1_HVT U1492 ( .A1(n14), .A2(n12), .Y(keyout[0]) );
  NAND4X0_HVT U1493 ( .A1(round_num[0]), .A2(n1424), .A3(n93), .A4(n1425), .Y(
        n12) );
  INVX0_HVT U1494 ( .A(round_num[3]), .Y(n1425) );
  INVX0_HVT U1495 ( .A(round_num[2]), .Y(n93) );
  INVX0_HVT U1496 ( .A(round_num[1]), .Y(n1424) );
  XNOR2X1_HVT U1497 ( .A1(keyin[0]), .A2(n1453), .Y(n14) );
  MUX21X1_HVT U1498 ( .A1(n1454), .A2(n1455), .S0(n26), .Y(n1453) );
  INVX0_HVT U1499 ( .A(keyin[111]), .Y(n26) );
  AO221X1_HVT U1500 ( .A1(n34), .A2(n1456), .A3(n27), .A4(n1457), .A5(n1458), 
        .Y(n1455) );
  AO22X1_HVT U1501 ( .A1(n32), .A2(n1459), .A3(n29), .A4(n1460), .Y(n1458) );
  AO221X1_HVT U1502 ( .A1(n52), .A2(n1461), .A3(n126), .A4(n46), .A5(n1462), 
        .Y(n1460) );
  AO22X1_HVT U1503 ( .A1(n1463), .A2(n55), .A3(n1362), .A4(n40), .Y(n1462) );
  AND2X1_HVT U1504 ( .A1(n122), .A2(n187), .Y(n1362) );
  INVX0_HVT U1505 ( .A(n143), .Y(n1463) );
  INVX0_HVT U1506 ( .A(n1408), .Y(n126) );
  NAND2X0_HVT U1507 ( .A1(n81), .A2(n1383), .Y(n1408) );
  NAND2X0_HVT U1508 ( .A1(n77), .A2(n44), .Y(n1383) );
  NAND2X0_HVT U1509 ( .A1(n179), .A2(n149), .Y(n1461) );
  OAI221X1_HVT U1510 ( .A1(n194), .A2(n167), .A3(n172), .A4(n106), .A5(n1464), 
        .Y(n1459) );
  OA22X1_HVT U1511 ( .A1(n108), .A2(n205), .A3(n42), .A4(n1321), .Y(n1464) );
  AND2X1_HVT U1512 ( .A1(n178), .A2(n115), .Y(n1321) );
  NAND2X0_HVT U1513 ( .A1(n37), .A2(n1331), .Y(n172) );
  NAND2X0_HVT U1514 ( .A1(keyin[110]), .A2(n116), .Y(n37) );
  NAND2X0_HVT U1515 ( .A1(n81), .A2(n138), .Y(n194) );
  AO221X1_HVT U1516 ( .A1(n52), .A2(n116), .A3(n203), .A4(n40), .A5(n1465), 
        .Y(n1457) );
  AO21X1_HVT U1517 ( .A1(n1309), .A2(n36), .A3(n133), .Y(n1465) );
  INVX0_HVT U1518 ( .A(n1369), .Y(n133) );
  NAND2X0_HVT U1519 ( .A1(n46), .A2(n107), .Y(n1369) );
  INVX0_HVT U1520 ( .A(n1403), .Y(n1309) );
  INVX0_HVT U1521 ( .A(n168), .Y(n203) );
  NAND2X0_HVT U1522 ( .A1(n115), .A2(n1331), .Y(n168) );
  AO221X1_HVT U1523 ( .A1(n46), .A2(n118), .A3(n36), .A4(n177), .A5(n1466), 
        .Y(n1456) );
  AO22X1_HVT U1524 ( .A1(n1420), .A2(n40), .A3(n52), .A4(n58), .Y(n1466) );
  NAND2X0_HVT U1525 ( .A1(n1403), .A2(n117), .Y(n58) );
  INVX0_HVT U1526 ( .A(n39), .Y(n1420) );
  NAND2X0_HVT U1527 ( .A1(n115), .A2(n187), .Y(n39) );
  NAND2X0_HVT U1528 ( .A1(n116), .A2(n44), .Y(n187) );
  NAND2X0_HVT U1529 ( .A1(n116), .A2(n179), .Y(n118) );
  NAND2X0_HVT U1530 ( .A1(keyin[110]), .A2(n107), .Y(n179) );
  AO221X1_HVT U1531 ( .A1(n32), .A2(n1467), .A3(n27), .A4(n1468), .A5(n1469), 
        .Y(n1454) );
  AO22X1_HVT U1532 ( .A1(n29), .A2(n1470), .A3(n34), .A4(n1471), .Y(n1469) );
  NAND3X0_HVT U1533 ( .A1(n1472), .A2(n1473), .A3(n1474), .Y(n1471) );
  AOI22X1_HVT U1534 ( .A1(n1350), .A2(n46), .A3(n78), .A4(n40), .Y(n1474) );
  NAND2X0_HVT U1535 ( .A1(n53), .A2(n1371), .Y(n78) );
  NAND2X0_HVT U1536 ( .A1(keyin[107]), .A2(keyin[110]), .Y(n1371) );
  NAND2X0_HVT U1537 ( .A1(n1316), .A2(n44), .Y(n53) );
  NAND2X0_HVT U1538 ( .A1(n81), .A2(n117), .Y(n1350) );
  NAND3X0_HVT U1539 ( .A1(n52), .A2(n115), .A3(n87), .Y(n1473) );
  NAND2X0_HVT U1540 ( .A1(keyin[110]), .A2(n77), .Y(n115) );
  AO21X1_HVT U1541 ( .A1(n177), .A2(n196), .A3(n108), .Y(n1472) );
  NAND2X0_HVT U1542 ( .A1(keyin[108]), .A2(n44), .Y(n196) );
  NAND2X0_HVT U1543 ( .A1(keyin[110]), .A2(n63), .Y(n177) );
  AND2X1_HVT U1544 ( .A1(keyin[109]), .A2(n1230), .Y(n34) );
  AO221X1_HVT U1545 ( .A1(n36), .A2(n84), .A3(n40), .A4(n77), .A5(n1475), .Y(
        n1470) );
  AO22X1_HVT U1546 ( .A1(n46), .A2(n1343), .A3(n52), .A4(n1476), .Y(n1475) );
  NAND2X0_HVT U1547 ( .A1(n145), .A2(n1367), .Y(n1476) );
  NAND2X0_HVT U1548 ( .A1(keyin[110]), .A2(n205), .Y(n1367) );
  NAND2X0_HVT U1549 ( .A1(n199), .A2(n44), .Y(n145) );
  NAND2X0_HVT U1550 ( .A1(n44), .A2(n205), .Y(n1343) );
  AND2X1_HVT U1551 ( .A1(n143), .A2(n173), .Y(n84) );
  NAND2X0_HVT U1552 ( .A1(n107), .A2(n44), .Y(n173) );
  NAND2X0_HVT U1553 ( .A1(n86), .A2(keyin[110]), .Y(n143) );
  INVX0_HVT U1554 ( .A(n77), .Y(n86) );
  NAND2X0_HVT U1555 ( .A1(keyin[107]), .A2(n199), .Y(n77) );
  INVX0_HVT U1556 ( .A(n166), .Y(n29) );
  NAND2X0_HVT U1557 ( .A1(keyin[109]), .A2(keyin[105]), .Y(n166) );
  AO221X1_HVT U1558 ( .A1(n36), .A2(n201), .A3(n40), .A4(n79), .A5(n1477), .Y(
        n1468) );
  AO222X1_HVT U1559 ( .A1(n46), .A2(n1403), .A3(n181), .A4(n52), .A5(n1349), 
        .A6(keyin[106]), .Y(n1477) );
  INVX0_HVT U1560 ( .A(n61), .Y(n1349) );
  INVX0_HVT U1561 ( .A(n167), .Y(n52) );
  NAND2X0_HVT U1562 ( .A1(keyin[106]), .A2(keyin[104]), .Y(n167) );
  INVX0_HVT U1563 ( .A(n139), .Y(n181) );
  NAND2X0_HVT U1564 ( .A1(n45), .A2(keyin[110]), .Y(n139) );
  INVX0_HVT U1565 ( .A(n63), .Y(n45) );
  NAND2X0_HVT U1566 ( .A1(keyin[108]), .A2(keyin[110]), .Y(n1403) );
  OAI21X1_HVT U1567 ( .A1(n63), .A2(keyin[110]), .A3(n122), .Y(n79) );
  NAND2X0_HVT U1568 ( .A1(n61), .A2(n137), .Y(n201) );
  NAND2X0_HVT U1569 ( .A1(n87), .A2(keyin[110]), .Y(n137) );
  NAND2X0_HVT U1570 ( .A1(n63), .A2(n44), .Y(n61) );
  NAND2X0_HVT U1571 ( .A1(keyin[108]), .A2(n205), .Y(n63) );
  INVX0_HVT U1572 ( .A(n164), .Y(n27) );
  NAND2X0_HVT U1573 ( .A1(keyin[105]), .A2(n1073), .Y(n164) );
  AO222X1_HVT U1574 ( .A1(n72), .A2(n1478), .A3(n40), .A4(n1479), .A5(n36), 
        .A6(n56), .Y(n1467) );
  NAND2X0_HVT U1575 ( .A1(n1331), .A2(n122), .Y(n56) );
  NAND2X0_HVT U1576 ( .A1(keyin[107]), .A2(n44), .Y(n1331) );
  INVX0_HVT U1577 ( .A(n108), .Y(n36) );
  NAND2X0_HVT U1578 ( .A1(n209), .A2(n55), .Y(n108) );
  NAND2X0_HVT U1579 ( .A1(n149), .A2(n81), .Y(n1479) );
  NAND2X0_HVT U1580 ( .A1(keyin[110]), .A2(n199), .Y(n81) );
  NAND2X0_HVT U1581 ( .A1(n44), .A2(n178), .Y(n149) );
  INVX0_HVT U1582 ( .A(n106), .Y(n40) );
  NAND2X0_HVT U1583 ( .A1(keyin[104]), .A2(n55), .Y(n106) );
  INVX0_HVT U1584 ( .A(keyin[106]), .Y(n55) );
  AO21X1_HVT U1585 ( .A1(keyin[106]), .A2(n1313), .A3(n46), .Y(n1478) );
  INVX0_HVT U1586 ( .A(n42), .Y(n46) );
  NAND2X0_HVT U1587 ( .A1(keyin[106]), .A2(n209), .Y(n42) );
  INVX0_HVT U1588 ( .A(keyin[104]), .Y(n209) );
  NAND2X0_HVT U1589 ( .A1(n122), .A2(n117), .Y(n1313) );
  NAND2X0_HVT U1590 ( .A1(n87), .A2(n44), .Y(n117) );
  INVX0_HVT U1591 ( .A(n107), .Y(n87) );
  NAND2X0_HVT U1592 ( .A1(n178), .A2(n116), .Y(n107) );
  NAND2X0_HVT U1593 ( .A1(n1385), .A2(keyin[110]), .Y(n122) );
  INVX0_HVT U1594 ( .A(n121), .Y(n72) );
  NAND2X0_HVT U1595 ( .A1(n195), .A2(n138), .Y(n121) );
  NAND2X0_HVT U1596 ( .A1(n1385), .A2(n44), .Y(n138) );
  INVX0_HVT U1597 ( .A(keyin[110]), .Y(n44) );
  INVX0_HVT U1598 ( .A(n116), .Y(n1385) );
  NAND2X0_HVT U1599 ( .A1(keyin[108]), .A2(keyin[107]), .Y(n116) );
  NAND2X0_HVT U1600 ( .A1(n1316), .A2(keyin[110]), .Y(n195) );
  INVX0_HVT U1601 ( .A(n178), .Y(n1316) );
  NAND2X0_HVT U1602 ( .A1(n199), .A2(n205), .Y(n178) );
  INVX0_HVT U1603 ( .A(keyin[107]), .Y(n205) );
  INVX0_HVT U1604 ( .A(keyin[108]), .Y(n199) );
  AND2X1_HVT U1605 ( .A1(n1230), .A2(n1073), .Y(n32) );
  INVX0_HVT U1606 ( .A(keyin[109]), .Y(n1073) );
  INVX0_HVT U1607 ( .A(keyin[105]), .Y(n1230) );
endmodule

