
module inv_sbox_2 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n33, n184, n185, n196, n197, n198, n199, n200, n201, n202, n206, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644;

  NAND2X0_HVT U1 ( .A1(n263), .A2(n353), .Y(n644) );
  NAND2X0_HVT U7 ( .A1(n276), .A2(n361), .Y(n637) );
  NAND2X0_HVT U8 ( .A1(n367), .A2(n244), .Y(n636) );
  NAND2X0_HVT U9 ( .A1(n366), .A2(n636), .Y(n635) );
  NAND2X0_HVT U10 ( .A1(n365), .A2(n633), .Y(n634) );
  NAND2X0_HVT U11 ( .A1(n289), .A2(n323), .Y(n632) );
  NAND2X0_HVT U12 ( .A1(n370), .A2(n351), .Y(n631) );
  NAND2X0_HVT U13 ( .A1(n363), .A2(n636), .Y(n630) );
  NAND2X0_HVT U15 ( .A1(n359), .A2(n369), .Y(n628) );
  NAND2X0_HVT U19 ( .A1(n276), .A2(n436), .Y(n623) );
  NAND2X0_HVT U32 ( .A1(n353), .A2(n289), .Y(n612) );
  NAND2X0_HVT U38 ( .A1(n351), .A2(n291), .Y(n606) );
  NAND2X0_HVT U42 ( .A1(n638), .A2(n437), .Y(n602) );
  OA21X1_HVT U53 ( .A1(n381), .A2(n594), .A3(n407), .Y(n592) );
  MUX41X1_HVT U56 ( .A1(n419), .A3(n360), .A2(n405), .A4(n590), .S0(n374), 
        .S1(n378), .Y(n589) );
  AO21X1_HVT U60 ( .A1(n584), .A2(n347), .A3(n622), .Y(n585) );
  NAND2X0_HVT U66 ( .A1(n276), .A2(n338), .Y(n578) );
  MUX41X1_HVT U67 ( .A1(n395), .A3(n420), .A2(n397), .A4(n578), .S0(n349), 
        .S1(n342), .Y(n577) );
  MUX41X1_HVT U68 ( .A1(n395), .A3(n310), .A2(n396), .A4(n366), .S0(n344), 
        .S1(n349), .Y(n576) );
  MUX41X1_HVT U69 ( .A1(n576), .A3(n579), .A2(n577), .A4(n580), .S0(n358), 
        .S1(n355), .Y(n575) );
  NAND2X0_HVT U72 ( .A1(n360), .A2(n281), .Y(n573) );
  MUX41X1_HVT U73 ( .A1(n616), .A3(n573), .A2(n421), .A4(n350), .S0(n348), 
        .S1(n341), .Y(n572) );
  MUX41X1_HVT U74 ( .A1(n634), .A3(n411), .A2(n410), .A4(n401), .S0(n344), 
        .S1(n378), .Y(n571) );
  MUX41X1_HVT U80 ( .A1(n422), .A3(n419), .A2(n635), .A4(n640), .S0(n344), 
        .S1(n378), .Y(n565) );
  NAND2X0_HVT U81 ( .A1(n323), .A2(n637), .Y(n564) );
  AND2X1_HVT U82 ( .A1(n294), .A2(n362), .Y(n563) );
  MUX41X1_HVT U83 ( .A1(n563), .A3(n409), .A2(n423), .A4(n564), .S0(n344), 
        .S1(n378), .Y(n562) );
  MUX41X1_HVT U84 ( .A1(n335), .A3(n231), .A2(n424), .A4(n314), .S0(n341), 
        .S1(n378), .Y(n561) );
  MUX41X1_HVT U85 ( .A1(n561), .A3(n565), .A2(n562), .A4(n566), .S0(n358), 
        .S1(n355), .Y(n560) );
  MUX41X1_HVT U88 ( .A1(n397), .A3(n384), .A2(n613), .A4(n598), .S0(n344), 
        .S1(n377), .Y(n558) );
  NAND2X0_HVT U89 ( .A1(n290), .A2(n434), .Y(n557) );
  MUX41X1_HVT U90 ( .A1(n317), .A3(n281), .A2(n597), .A4(n557), .S0(n344), 
        .S1(n378), .Y(n556) );
  MUX41X1_HVT U96 ( .A1(n420), .A3(n630), .A2(n406), .A4(n426), .S0(n340), 
        .S1(n377), .Y(n550) );
  MUX41X1_HVT U99 ( .A1(n612), .A3(n399), .A2(n596), .A4(n360), .S0(n378), 
        .S1(n342), .Y(n547) );
  MUX41X1_HVT U101 ( .A1(n428), .A3(n631), .A2(n238), .A4(n546), .S0(n349), 
        .S1(n340), .Y(n545) );
  MUX41X1_HVT U102 ( .A1(n545), .A3(n548), .A2(n547), .A4(n550), .S0(in[5]), 
        .S1(n355), .Y(n544) );
  AND2X1_HVT U104 ( .A1(n281), .A2(n322), .Y(n543) );
  MUX41X1_HVT U105 ( .A1(n629), .A3(n429), .A2(n564), .A4(n543), .S0(n346), 
        .S1(n377), .Y(n542) );
  MUX41X1_HVT U107 ( .A1(n428), .A3(n362), .A2(n541), .A4(n389), .S0(n344), 
        .S1(n377), .Y(n540) );
  MUX41X1_HVT U108 ( .A1(n401), .A3(n360), .A2(n405), .A4(n321), .S0(n374), 
        .S1(n377), .Y(n539) );
  MUX41X1_HVT U109 ( .A1(n427), .A3(n384), .A2(n424), .A4(n417), .S0(n344), 
        .S1(n309), .Y(n538) );
  MUX41X1_HVT U110 ( .A1(n538), .A3(n540), .A2(n539), .A4(n542), .S0(n358), 
        .S1(n356), .Y(n537) );
  NAND2X0_HVT U114 ( .A1(n365), .A2(n281), .Y(n533) );
  MUX41X1_HVT U115 ( .A1(n533), .A3(n632), .A2(n414), .A4(n363), .S0(n265), 
        .S1(n342), .Y(n532) );
  MUX41X1_HVT U116 ( .A1(n413), .A3(n237), .A2(n384), .A4(n628), .S0(n343), 
        .S1(n377), .Y(n531) );
  NAND2X0_HVT U118 ( .A1(n290), .A2(n310), .Y(n529) );
  MUX41X1_HVT U119 ( .A1(n430), .A3(n530), .A2(n243), .A4(n529), .S0(n343), 
        .S1(n377), .Y(n528) );
  MUX41X1_HVT U120 ( .A1(n528), .A3(n532), .A2(n531), .A4(n534), .S0(in[5]), 
        .S1(n355), .Y(n527) );
  MUX41X1_HVT U122 ( .A1(n418), .A3(n332), .A2(n598), .A4(n272), .S0(n343), 
        .S1(n309), .Y(n526) );
  MUX41X1_HVT U124 ( .A1(n334), .A3(n525), .A2(n620), .A4(n402), .S0(n347), 
        .S1(n343), .Y(n524) );
  AOI21X1_HVT U127 ( .A1(n345), .A2(n520), .A3(n390), .Y(n521) );
  NAND2X0_HVT U129 ( .A1(n346), .A2(n365), .Y(n518) );
  MUX41X1_HVT U130 ( .A1(n518), .A3(n519), .A2(n522), .A4(n521), .S0(n349), 
        .S1(n356), .Y(n517) );
  AND2X1_HVT U131 ( .A1(n338), .A2(n291), .Y(n516) );
  MUX41X1_HVT U132 ( .A1(n324), .A3(n516), .A2(n432), .A4(n395), .S0(n348), 
        .S1(n341), .Y(n515) );
  MUX41X1_HVT U133 ( .A1(n433), .A3(n389), .A2(n590), .A4(n388), .S0(n347), 
        .S1(n340), .Y(n514) );
  MUX41X1_HVT U136 ( .A1(n595), .A3(n546), .A2(n512), .A4(n393), .S0(n346), 
        .S1(n309), .Y(n511) );
  MUX41X1_HVT U137 ( .A1(n315), .A3(n614), .A2(n314), .A4(n426), .S0(n349), 
        .S1(n340), .Y(n510) );
  MUX41X1_HVT U140 ( .A1(n410), .A3(n333), .A2(n404), .A4(n632), .S0(n348), 
        .S1(n342), .Y(n508) );
  NAND2X0_HVT U141 ( .A1(n359), .A2(n291), .Y(n507) );
  MUX41X1_HVT U142 ( .A1(n507), .A3(n605), .A2(n431), .A4(n404), .S0(n374), 
        .S1(n309), .Y(n506) );
  MUX41X1_HVT U145 ( .A1(n316), .A3(n429), .A2(n504), .A4(n564), .S0(n345), 
        .S1(n271), .Y(n503) );
  MUX41X1_HVT U146 ( .A1(n503), .A3(n505), .A2(n506), .A4(n508), .S0(n356), 
        .S1(n358), .Y(n502) );
  AO21X1_HVT U148 ( .A1(n349), .A2(n391), .A3(n326), .Y(n500) );
  MUX41X1_HVT U151 ( .A1(n423), .A3(n412), .A2(n250), .A4(n498), .S0(n347), 
        .S1(n340), .Y(n497) );
  MUX41X1_HVT U155 ( .A1(n404), .A3(n632), .A2(n624), .A4(n406), .S0(n345), 
        .S1(n271), .Y(n493) );
  NAND2X0_HVT U159 ( .A1(n489), .A2(n488), .Y(n490) );
  NAND2X0_HVT U163 ( .A1(n367), .A2(n434), .Y(n484) );
  MUX41X1_HVT U164 ( .A1(n635), .A3(n484), .A2(n243), .A4(n401), .S0(n343), 
        .S1(n271), .Y(n483) );
  NAND2X0_HVT U166 ( .A1(n633), .A2(n480), .Y(n481) );
  MUX41X1_HVT U174 ( .A1(n425), .A3(n590), .A2(n433), .A4(n437), .S0(n345), 
        .S1(n271), .Y(n472) );
  NAND2X0_HVT U177 ( .A1(n370), .A2(n310), .Y(n470) );
  AND2X1_HVT U179 ( .A1(n294), .A2(n244), .Y(n468) );
  MUX41X1_HVT U180 ( .A1(n612), .A3(n382), .A2(n468), .A4(n599), .S0(n345), 
        .S1(n376), .Y(n467) );
  MUX41X1_HVT U183 ( .A1(n415), .A3(n419), .A2(n401), .A4(n602), .S0(n347), 
        .S1(n341), .Y(n464) );
  NAND2X0_HVT U191 ( .A1(n381), .A2(n394), .Y(n458) );
  AND2X1_HVT U192 ( .A1(n411), .A2(n456), .Y(n457) );
  NAND2X0_HVT U194 ( .A1(n456), .A2(n602), .Y(n454) );
  MUX41X1_HVT U195 ( .A1(n455), .A3(n454), .A2(n457), .A4(n458), .S0(n344), 
        .S1(n356), .Y(n453) );
  NAND2X0_HVT U198 ( .A1(n277), .A2(n437), .Y(n633) );
  NAND2X0_HVT U200 ( .A1(n244), .A2(n290), .Y(n520) );
  NAND2X0_HVT U207 ( .A1(n291), .A2(n317), .Y(n584) );
  MUX21X1_HVT U2 ( .A1(n321), .A2(n361), .S0(n373), .Y(n625) );
  IBUFFX2_HVT U3 ( .A(n372), .Y(n367) );
  MUX41X1_HVT U4 ( .A1(n466), .A3(n463), .A2(n459), .A4(n453), .S0(n357), .S1(
        n33), .Y(out[7]) );
  IBUFFX16_HVT U5 ( .A(n292), .Y(n33) );
  MUX21X2_HVT U6 ( .A1(n338), .A2(n366), .S0(n247), .Y(n626) );
  INVX1_HVT U14 ( .A(n381), .Y(n201) );
  NAND2X0_HVT U16 ( .A1(n360), .A2(n184), .Y(n185) );
  NAND2X0_HVT U17 ( .A1(n317), .A2(n367), .Y(n196) );
  NAND2X0_HVT U18 ( .A1(n185), .A2(n196), .Y(n316) );
  IBUFFX2_HVT U20 ( .A(n367), .Y(n184) );
  NAND2X0_HVT U21 ( .A1(n492), .A2(n197), .Y(n198) );
  NAND2X0_HVT U22 ( .A1(n502), .A2(n206), .Y(n199) );
  NAND2X0_HVT U23 ( .A1(n198), .A2(n199), .Y(out[5]) );
  INVX0_HVT U24 ( .A(n206), .Y(n197) );
  IBUFFX2_HVT U25 ( .A(n295), .Y(n206) );
  MUX21X2_HVT U26 ( .A1(n627), .A2(n251), .S0(n370), .Y(n250) );
  MUX21X1_HVT U27 ( .A1(n279), .A2(n359), .S0(n349), .Y(n553) );
  NBUFFX4_HVT U28 ( .A(n435), .Y(n350) );
  INVX1_HVT U29 ( .A(n329), .Y(n321) );
  MUX21X2_HVT U30 ( .A1(n317), .A2(n360), .S0(n368), .Y(n446) );
  MUX21X2_HVT U31 ( .A1(n422), .A2(n219), .S0(n220), .Y(n218) );
  MUX41X1_HVT U33 ( .A1(n408), .A3(n625), .A2(n319), .A4(n626), .S0(n200), 
        .S1(n201), .Y(n566) );
  IBUFFX16_HVT U34 ( .A(n293), .Y(n200) );
  INVX1_HVT U35 ( .A(n371), .Y(n373) );
  IBUFFX2_HVT U36 ( .A(n325), .Y(n600) );
  INVX1_HVT U37 ( .A(n446), .Y(n425) );
  MUX21X2_HVT U39 ( .A1(n592), .A2(n593), .S0(n202), .Y(n591) );
  IBUFFX16_HVT U40 ( .A(n346), .Y(n202) );
  INVX1_HVT U41 ( .A(n627), .Y(n437) );
  IBUFFX16_HVT U43 ( .A(n298), .Y(n219) );
  IBUFFX16_HVT U44 ( .A(n347), .Y(n220) );
  INVX1_HVT U45 ( .A(n449), .Y(n422) );
  MUX21X1_HVT U46 ( .A1(n366), .A2(n222), .S0(n369), .Y(n221) );
  IBUFFX16_HVT U47 ( .A(n221), .Y(n475) );
  IBUFFX16_HVT U48 ( .A(n354), .Y(n222) );
  MUX41X1_HVT U49 ( .A1(n621), .A3(n331), .A2(n475), .A4(n557), .S0(n223), 
        .S1(n224), .Y(n474) );
  IBUFFX16_HVT U50 ( .A(n345), .Y(n223) );
  IBUFFX16_HVT U51 ( .A(n271), .Y(n224) );
  INVX0_HVT U52 ( .A(n316), .Y(n319) );
  MUX41X1_HVT U54 ( .A1(n218), .A3(n460), .A2(n462), .A4(n461), .S0(n225), 
        .S1(n226), .Y(n459) );
  IBUFFX16_HVT U55 ( .A(n356), .Y(n225) );
  IBUFFX16_HVT U57 ( .A(n341), .Y(n226) );
  MUX41X1_HVT U58 ( .A1(n279), .A3(n632), .A2(n317), .A4(n294), .S0(n227), 
        .S1(n262), .Y(n574) );
  IBUFFX16_HVT U59 ( .A(n344), .Y(n227) );
  IBUFFX2_HVT U61 ( .A(n380), .Y(n378) );
  INVX2_HVT U62 ( .A(n376), .Y(n262) );
  AO21X1_HVT U63 ( .A1(n291), .A2(n366), .A3(n381), .Y(n488) );
  INVX0_HVT U64 ( .A(n598), .Y(n417) );
  INVX1_HVT U65 ( .A(in[6]), .Y(n438) );
  NBUFFX2_HVT U70 ( .A(n438), .Y(n352) );
  NBUFFX2_HVT U71 ( .A(n438), .Y(n354) );
  INVX0_HVT U75 ( .A(n250), .Y(n621) );
  MUX21X2_HVT U76 ( .A1(n365), .A2(n322), .S0(n289), .Y(n325) );
  MUX41X1_HVT U77 ( .A1(n591), .A3(n587), .A2(n589), .A4(n583), .S0(n357), 
        .S1(n330), .Y(n582) );
  IBUFFX2_HVT U78 ( .A(n330), .Y(n355) );
  INVX0_HVT U79 ( .A(n347), .Y(n278) );
  INVX0_HVT U86 ( .A(n347), .Y(n253) );
  MUX41X1_HVT U87 ( .A1(n568), .A3(n571), .A2(n572), .A4(n574), .S0(n355), 
        .S1(n358), .Y(n567) );
  NAND2X0_HVT U91 ( .A1(n569), .A2(n228), .Y(n229) );
  NAND2X0_HVT U92 ( .A1(n570), .A2(n249), .Y(n230) );
  NAND2X0_HVT U93 ( .A1(n229), .A2(n230), .Y(n568) );
  INVX0_HVT U94 ( .A(n249), .Y(n228) );
  INVX1_HVT U95 ( .A(n357), .Y(n358) );
  IBUFFX2_HVT U97 ( .A(n345), .Y(n249) );
  INVX0_HVT U98 ( .A(n326), .Y(n251) );
  INVX0_HVT U100 ( .A(n372), .Y(n369) );
  INVX0_HVT U103 ( .A(n236), .Y(n231) );
  INVX1_HVT U106 ( .A(n408), .Y(n236) );
  MUX21X2_HVT U111 ( .A1(n510), .A2(n511), .S0(n356), .Y(n509) );
  MUX21X2_HVT U112 ( .A1(n403), .A2(n588), .S0(n337), .Y(n587) );
  XOR2X2_HVT U113 ( .A1(n352), .A2(n263), .Y(n627) );
  NAND2X0_HVT U117 ( .A1(n544), .A2(n232), .Y(n233) );
  NAND2X0_HVT U121 ( .A1(n551), .A2(in[7]), .Y(n234) );
  NAND2X0_HVT U123 ( .A1(n233), .A2(n234), .Y(out[2]) );
  IBUFFX2_HVT U125 ( .A(in[7]), .Y(n232) );
  MUX21X2_HVT U126 ( .A1(n537), .A2(n527), .S0(n235), .Y(out[3]) );
  IBUFFX16_HVT U128 ( .A(in[7]), .Y(n235) );
  INVX0_HVT U134 ( .A(n236), .Y(n237) );
  MUX21X1_HVT U135 ( .A1(n322), .A2(n363), .S0(n277), .Y(n486) );
  AO21X2_HVT U138 ( .A1(n414), .A2(n348), .A3(n619), .Y(n535) );
  INVX1_HVT U139 ( .A(n238), .Y(n608) );
  MUX21X1_HVT U143 ( .A1(n239), .A2(n627), .S0(n277), .Y(n238) );
  IBUFFX16_HVT U144 ( .A(n352), .Y(n239) );
  MUX41X1_HVT U147 ( .A1(n608), .A3(n364), .A2(n317), .A4(n365), .S0(n240), 
        .S1(n241), .Y(n473) );
  IBUFFX16_HVT U149 ( .A(n345), .Y(n240) );
  IBUFFX16_HVT U150 ( .A(n376), .Y(n241) );
  INVX1_HVT U152 ( .A(n607), .Y(n242) );
  INVX1_HVT U153 ( .A(n242), .Y(n243) );
  NBUFFX2_HVT U154 ( .A(n639), .Y(n244) );
  NAND2X0_HVT U156 ( .A1(in[6]), .A2(n351), .Y(n639) );
  NBUFFX4_HVT U157 ( .A(n435), .Y(n351) );
  XNOR2X1_HVT U158 ( .A1(n245), .A2(n247), .Y(n607) );
  IBUFFX16_HVT U160 ( .A(n365), .Y(n245) );
  MUX21X2_HVT U161 ( .A1(n554), .A2(n553), .S0(n246), .Y(n552) );
  IBUFFX16_HVT U162 ( .A(n346), .Y(n246) );
  INVX1_HVT U165 ( .A(n366), .Y(n317) );
  INVX0_HVT U167 ( .A(n639), .Y(n434) );
  IBUFFX2_HVT U168 ( .A(n372), .Y(n247) );
  MUX21X2_HVT U169 ( .A1(n390), .A2(n603), .S0(n349), .Y(n536) );
  INVX1_HVT U170 ( .A(n607), .Y(n412) );
  MUX41X1_HVT U171 ( .A1(n400), .A3(n325), .A2(n486), .A4(n609), .S0(n248), 
        .S1(n271), .Y(n485) );
  IBUFFX16_HVT U172 ( .A(n345), .Y(n248) );
  INVX0_HVT U173 ( .A(n279), .Y(n609) );
  XOR2X2_HVT U175 ( .A1(n322), .A2(n368), .Y(n596) );
  XOR2X2_HVT U176 ( .A1(n360), .A2(n276), .Y(n598) );
  INVX1_HVT U178 ( .A(n372), .Y(n371) );
  MUX21X2_HVT U181 ( .A1(n320), .A2(n250), .S0(n252), .Y(n581) );
  IBUFFX16_HVT U182 ( .A(n346), .Y(n252) );
  MUX21X1_HVT U184 ( .A1(n353), .A2(n350), .S0(n373), .Y(n599) );
  MUX21X2_HVT U185 ( .A1(n272), .A2(n601), .S0(n301), .Y(n491) );
  INVX1_HVT U186 ( .A(n259), .Y(n272) );
  NAND2X0_HVT U187 ( .A1(n617), .A2(n253), .Y(n254) );
  NAND2X0_HVT U188 ( .A1(n620), .A2(n347), .Y(n255) );
  NAND2X0_HVT U189 ( .A1(n254), .A2(n255), .Y(n482) );
  NBUFFX4_HVT U190 ( .A(n379), .Y(n347) );
  INVX0_HVT U193 ( .A(n620), .Y(n402) );
  MUX21X2_HVT U196 ( .A1(n401), .A2(n581), .S0(n337), .Y(n580) );
  INVX1_HVT U197 ( .A(n372), .Y(n370) );
  INVX1_HVT U199 ( .A(n614), .Y(n408) );
  OA21X1_HVT U201 ( .A1(n381), .A2(n408), .A3(n584), .Y(n460) );
  MUX21X1_HVT U202 ( .A1(n351), .A2(n321), .S0(n277), .Y(n449) );
  INVX0_HVT U203 ( .A(n369), .Y(n269) );
  MUX21X1_HVT U204 ( .A1(n322), .A2(n310), .S0(n276), .Y(n549) );
  NAND2X0_HVT U205 ( .A1(n490), .A2(n256), .Y(n257) );
  NAND2X0_HVT U206 ( .A1(n491), .A2(n340), .Y(n258) );
  NAND2X0_HVT U208 ( .A1(n257), .A2(n258), .Y(n487) );
  IBUFFX2_HVT U209 ( .A(n340), .Y(n256) );
  MUX21X1_HVT U210 ( .A1(n260), .A2(n351), .S0(n370), .Y(n259) );
  IBUFFX16_HVT U211 ( .A(n361), .Y(n260) );
  MUX41X1_HVT U212 ( .A1(n423), .A3(n387), .A2(n320), .A4(n389), .S0(n261), 
        .S1(n262), .Y(n465) );
  IBUFFX16_HVT U213 ( .A(n343), .Y(n261) );
  INVX2_HVT U214 ( .A(n347), .Y(n311) );
  INVX0_HVT U215 ( .A(n349), .Y(n286) );
  INVX1_HVT U216 ( .A(n380), .Y(n379) );
  INVX2_HVT U217 ( .A(n311), .Y(n309) );
  NBUFFX2_HVT U218 ( .A(in[3]), .Y(n263) );
  OR2X1_HVT U219 ( .A1(n435), .A2(n354), .Y(n642) );
  IBUFFX2_HVT U220 ( .A(n435), .Y(n310) );
  INVX1_HVT U221 ( .A(n354), .Y(n338) );
  INVX0_HVT U222 ( .A(n601), .Y(n415) );
  INVX0_HVT U223 ( .A(n377), .Y(n264) );
  INVX1_HVT U224 ( .A(n264), .Y(n265) );
  IBUFFX4_HVT U225 ( .A(n380), .Y(n377) );
  NAND2X0_HVT U226 ( .A1(n560), .A2(n266), .Y(n267) );
  NAND2X0_HVT U227 ( .A1(n567), .A2(in[7]), .Y(n268) );
  NAND2X0_HVT U228 ( .A1(n267), .A2(n268), .Y(out[1]) );
  IBUFFX2_HVT U229 ( .A(in[7]), .Y(n266) );
  OA21X2_HVT U230 ( .A1(n385), .A2(n381), .A3(n392), .Y(n495) );
  AO21X2_HVT U231 ( .A1(n360), .A2(n320), .A3(n381), .Y(n480) );
  MUX21X1_HVT U232 ( .A1(n272), .A2(n383), .S0(n349), .Y(n570) );
  MUX21X2_HVT U233 ( .A1(n535), .A2(n536), .S0(n342), .Y(n534) );
  MUX21X1_HVT U234 ( .A1(n353), .A2(n363), .S0(n269), .Y(n525) );
  MUX21X2_HVT U235 ( .A1(n526), .A2(n524), .S0(n270), .Y(n523) );
  IBUFFX16_HVT U236 ( .A(n356), .Y(n270) );
  NBUFFX16_HVT U237 ( .A(n379), .Y(n349) );
  MUX21X2_HVT U238 ( .A1(n351), .A2(n436), .S0(n277), .Y(n601) );
  NBUFFX2_HVT U239 ( .A(n376), .Y(n271) );
  INVX1_HVT U240 ( .A(n380), .Y(n376) );
  MUX21X1_HVT U241 ( .A1(n406), .A2(n396), .S0(n349), .Y(n593) );
  INVX1_HVT U242 ( .A(n363), .Y(n285) );
  INVX1_HVT U243 ( .A(n361), .Y(n436) );
  NAND2X0_HVT U244 ( .A1(n585), .A2(n273), .Y(n274) );
  NAND2X0_HVT U245 ( .A1(n586), .A2(n293), .Y(n275) );
  NAND2X0_HVT U246 ( .A1(n274), .A2(n275), .Y(n583) );
  IBUFFX2_HVT U247 ( .A(n293), .Y(n273) );
  IBUFFX2_HVT U248 ( .A(n372), .Y(n276) );
  INVX1_HVT U249 ( .A(n372), .Y(n277) );
  MUX21X1_HVT U250 ( .A1(n402), .A2(n590), .S0(n348), .Y(n586) );
  MUX21X2_HVT U251 ( .A1(n334), .A2(n416), .S0(n278), .Y(n455) );
  INVX1_HVT U252 ( .A(n622), .Y(n401) );
  OA21X1_HVT U253 ( .A1(n386), .A2(n381), .A3(n622), .Y(n569) );
  AND2X1_HVT U254 ( .A1(n636), .A2(n437), .Y(n279) );
  MUX41X1_HVT U255 ( .A1(n487), .A3(n485), .A2(n483), .A4(n479), .S0(n280), 
        .S1(n357), .Y(n478) );
  IBUFFX16_HVT U256 ( .A(n355), .Y(n280) );
  INVX1_HVT U257 ( .A(n390), .Y(n281) );
  INVX1_HVT U258 ( .A(n637), .Y(n390) );
  NAND2X0_HVT U259 ( .A1(n481), .A2(n282), .Y(n283) );
  NAND2X0_HVT U260 ( .A1(n482), .A2(n346), .Y(n284) );
  NAND2X0_HVT U261 ( .A1(n283), .A2(n284), .Y(n479) );
  IBUFFX2_HVT U262 ( .A(n346), .Y(n282) );
  MUX21X1_HVT U263 ( .A1(n329), .A2(n310), .S0(n369), .Y(n620) );
  OR2X1_HVT U264 ( .A1(n285), .A2(n387), .Y(n590) );
  INVX0_HVT U265 ( .A(n387), .Y(n320) );
  IBUFFX2_HVT U266 ( .A(n636), .Y(n391) );
  NAND2X0_HVT U267 ( .A1(n335), .A2(n286), .Y(n287) );
  NAND2X0_HVT U268 ( .A1(n596), .A2(n349), .Y(n288) );
  NAND2X0_HVT U269 ( .A1(n287), .A2(n288), .Y(n462) );
  INVX1_HVT U270 ( .A(in[0]), .Y(n372) );
  NBUFFX2_HVT U271 ( .A(n373), .Y(n289) );
  NBUFFX2_HVT U272 ( .A(n373), .Y(n290) );
  NBUFFX2_HVT U273 ( .A(n373), .Y(n291) );
  INVX1_HVT U274 ( .A(n330), .Y(n356) );
  INVX1_HVT U275 ( .A(n295), .Y(n292) );
  INVX0_HVT U276 ( .A(n643), .Y(n326) );
  INVX1_HVT U277 ( .A(in[7]), .Y(n295) );
  INVX1_HVT U278 ( .A(in[1]), .Y(n330) );
  INVX1_HVT U279 ( .A(in[5]), .Y(n357) );
  INVX1_HVT U280 ( .A(n374), .Y(n293) );
  INVX0_HVT U281 ( .A(n348), .Y(n301) );
  MUX41X1_HVT U282 ( .A1(n387), .A3(n335), .A2(n425), .A4(n405), .S0(n343), 
        .S1(n378), .Y(n559) );
  MUX41X1_HVT U283 ( .A1(n552), .A3(n556), .A2(n558), .A4(n559), .S0(n355), 
        .S1(n358), .Y(n551) );
  MUX41X1_HVT U284 ( .A1(n427), .A3(n549), .A2(n615), .A4(n412), .S0(n293), 
        .S1(n377), .Y(n548) );
  INVX1_HVT U285 ( .A(n388), .Y(n294) );
  INVX0_HVT U286 ( .A(n638), .Y(n388) );
  IBUFFX2_HVT U287 ( .A(n615), .Y(n407) );
  NAND2X0_HVT U288 ( .A1(n471), .A2(n295), .Y(n296) );
  NAND2X0_HVT U289 ( .A1(n370), .A2(n366), .Y(n638) );
  NAND2X0_HVT U290 ( .A1(n478), .A2(in[7]), .Y(n297) );
  NAND2X0_HVT U291 ( .A1(n296), .A2(n297), .Y(out[6]) );
  INVX1_HVT U292 ( .A(n602), .Y(n389) );
  MUX41X1_HVT U293 ( .A1(n472), .A3(n473), .A2(n474), .A4(n476), .S0(n356), 
        .S1(n358), .Y(n471) );
  NAND2X0_HVT U294 ( .A1(n437), .A2(n290), .Y(n298) );
  NAND2X0_HVT U295 ( .A1(n464), .A2(n330), .Y(n299) );
  NAND2X0_HVT U296 ( .A1(n465), .A2(n356), .Y(n300) );
  NAND2X0_HVT U297 ( .A1(n299), .A2(n300), .Y(n463) );
  IBUFFX2_HVT U298 ( .A(n372), .Y(n368) );
  NAND2X0_HVT U299 ( .A1(n421), .A2(n301), .Y(n302) );
  NAND2X0_HVT U300 ( .A1(n603), .A2(n348), .Y(n303) );
  NAND2X0_HVT U301 ( .A1(n302), .A2(n303), .Y(n461) );
  NAND2X0_HVT U302 ( .A1(n469), .A2(n304), .Y(n305) );
  NAND2X0_HVT U303 ( .A1(n467), .A2(n330), .Y(n306) );
  NAND2X0_HVT U304 ( .A1(n305), .A2(n306), .Y(n466) );
  INVX0_HVT U305 ( .A(n330), .Y(n304) );
  NAND2X0_HVT U306 ( .A1(n575), .A2(n295), .Y(n307) );
  NAND2X0_HVT U307 ( .A1(n582), .A2(in[7]), .Y(n308) );
  NAND2X0_HVT U308 ( .A1(n308), .A2(n307), .Y(out[0]) );
  INVX0_HVT U309 ( .A(n327), .Y(n498) );
  INVX0_HVT U310 ( .A(n352), .Y(n328) );
  MUX21X1_HVT U311 ( .A1(n324), .A2(n432), .S0(n311), .Y(n501) );
  INVX0_HVT U312 ( .A(n369), .Y(n318) );
  MUX21X1_HVT U313 ( .A1(n359), .A2(n351), .S0(n277), .Y(n622) );
  INVX0_HVT U314 ( .A(in[3]), .Y(n435) );
  INVX0_HVT U315 ( .A(n324), .Y(n640) );
  INVX1_HVT U316 ( .A(in[4]), .Y(n381) );
  MUX41X1_HVT U317 ( .A1(n606), .A3(n399), .A2(n400), .A4(n398), .S0(n293), 
        .S1(n381), .Y(n579) );
  AO21X2_HVT U318 ( .A1(n368), .A2(n326), .A3(n381), .Y(n456) );
  MUX41X1_HVT U319 ( .A1(n509), .A3(n513), .A2(n517), .A4(n523), .S0(in[5]), 
        .S1(in[7]), .Y(out[4]) );
  MUX21X1_HVT U320 ( .A1(n354), .A2(n627), .S0(n372), .Y(n618) );
  NAND2X0_HVT U321 ( .A1(n514), .A2(n330), .Y(n312) );
  NAND2X0_HVT U322 ( .A1(n515), .A2(n355), .Y(n313) );
  NAND2X0_HVT U323 ( .A1(n312), .A2(n313), .Y(n513) );
  NBUFFX2_HVT U324 ( .A(n618), .Y(n314) );
  INVX0_HVT U325 ( .A(n391), .Y(n315) );
  XOR2X2_HVT U326 ( .A1(n364), .A2(n318), .Y(n333) );
  NAND2X0_HVT U327 ( .A1(n368), .A2(n364), .Y(n641) );
  NBUFFX2_HVT U328 ( .A(n639), .Y(n322) );
  INVX1_HVT U329 ( .A(n440), .Y(n432) );
  MUX21X1_HVT U330 ( .A1(n323), .A2(n244), .S0(n289), .Y(n440) );
  INVX1_HVT U331 ( .A(n452), .Y(n419) );
  NBUFFX2_HVT U332 ( .A(n643), .Y(n323) );
  AND2X1_HVT U333 ( .A1(n641), .A2(n244), .Y(n324) );
  MUX21X1_HVT U334 ( .A1(n244), .A2(n328), .S0(n290), .Y(n327) );
  AND2X1_HVT U335 ( .A1(n350), .A2(n352), .Y(n329) );
  INVX1_HVT U336 ( .A(n611), .Y(n410) );
  MUX41X1_HVT U337 ( .A1(n499), .A3(n494), .A2(n497), .A4(n493), .S0(n357), 
        .S1(n330), .Y(n492) );
  MUX41X1_HVT U338 ( .A1(n623), .A3(n620), .A2(n434), .A4(n415), .S0(n345), 
        .S1(n311), .Y(n505) );
  MUX41X1_HVT U339 ( .A1(n600), .A3(n317), .A2(n470), .A4(n336), .S0(n293), 
        .S1(n311), .Y(n469) );
  INVX1_HVT U340 ( .A(n450), .Y(n421) );
  MUX21X2_HVT U341 ( .A1(n501), .A2(n500), .S0(n346), .Y(n499) );
  INVX0_HVT U342 ( .A(n339), .Y(n477) );
  NBUFFX2_HVT U343 ( .A(n643), .Y(n364) );
  AND2X1_HVT U344 ( .A1(n294), .A2(n321), .Y(n331) );
  AND2X1_HVT U345 ( .A1(n364), .A2(n628), .Y(n332) );
  NAND2X0_HVT U346 ( .A1(n350), .A2(n352), .Y(n643) );
  MUX21X1_HVT U347 ( .A1(n437), .A2(n350), .S0(n370), .Y(n605) );
  MUX21X1_HVT U348 ( .A1(n323), .A2(n322), .S0(n367), .Y(n504) );
  MUX21X1_HVT U349 ( .A1(n437), .A2(n354), .S0(n370), .Y(n441) );
  MUX21X1_HVT U350 ( .A1(n317), .A2(n434), .S0(n369), .Y(n615) );
  MUX21X1_HVT U351 ( .A1(n350), .A2(n326), .S0(n247), .Y(n613) );
  MUX21X1_HVT U352 ( .A1(n326), .A2(n436), .S0(n369), .Y(n594) );
  MUX21X1_HVT U353 ( .A1(n359), .A2(n434), .S0(n368), .Y(n610) );
  MUX21X1_HVT U354 ( .A1(n555), .A2(n363), .S0(n369), .Y(n554) );
  MUX21X1_HVT U355 ( .A1(n359), .A2(n354), .S0(n348), .Y(n555) );
  MUX21X1_HVT U356 ( .A1(n431), .A2(n333), .S0(n346), .Y(n522) );
  XOR2X1_HVT U357 ( .A1(n362), .A2(n368), .Y(n597) );
  INVX0_HVT U358 ( .A(n605), .Y(n413) );
  MUX21X1_HVT U359 ( .A1(n363), .A2(n350), .S0(n247), .Y(n624) );
  MUX21X1_HVT U360 ( .A1(n404), .A2(n640), .S0(n341), .Y(n588) );
  MUX21X1_HVT U361 ( .A1(n352), .A2(n321), .S0(n371), .Y(n541) );
  MUX21X1_HVT U362 ( .A1(n365), .A2(n321), .S0(n371), .Y(n629) );
  MUX21X1_HVT U363 ( .A1(n352), .A2(n360), .S0(n367), .Y(n604) );
  MUX21X1_HVT U364 ( .A1(n350), .A2(n362), .S0(n371), .Y(n443) );
  AND2X1_HVT U365 ( .A1(n367), .A2(n354), .Y(n334) );
  NBUFFX2_HVT U366 ( .A(n379), .Y(n348) );
  MUX21X1_HVT U367 ( .A1(n495), .A2(n496), .S0(n340), .Y(n494) );
  MUX21X1_HVT U368 ( .A1(n618), .A2(n335), .S0(n348), .Y(n496) );
  NAND2X0_HVT U369 ( .A1(n290), .A2(n329), .Y(n546) );
  NBUFFX2_HVT U370 ( .A(n644), .Y(n365) );
  NBUFFX2_HVT U371 ( .A(n627), .Y(n360) );
  AND2X1_HVT U372 ( .A1(n363), .A2(n372), .Y(n335) );
  AND2X1_HVT U373 ( .A1(n436), .A2(n291), .Y(n336) );
  NBUFFX2_HVT U374 ( .A(n642), .Y(n361) );
  NBUFFX2_HVT U375 ( .A(n642), .Y(n363) );
  NBUFFX2_HVT U376 ( .A(n627), .Y(n359) );
  NBUFFX2_HVT U377 ( .A(n642), .Y(n362) );
  NBUFFX2_HVT U378 ( .A(n644), .Y(n366) );
  NBUFFX2_HVT U379 ( .A(n375), .Y(n345) );
  NBUFFX2_HVT U380 ( .A(n375), .Y(n346) );
  NBUFFX2_HVT U381 ( .A(n438), .Y(n353) );
  XNOR2X1_HVT U382 ( .A1(n381), .A2(n343), .Y(n337) );
  NBUFFX2_HVT U383 ( .A(n375), .Y(n343) );
  NBUFFX2_HVT U384 ( .A(n374), .Y(n342) );
  NBUFFX2_HVT U385 ( .A(n374), .Y(n340) );
  NBUFFX2_HVT U386 ( .A(n374), .Y(n344) );
  NBUFFX2_HVT U387 ( .A(n374), .Y(n341) );
  MUX21X1_HVT U388 ( .A1(n317), .A2(n310), .S0(n247), .Y(n439) );
  MUX21X1_HVT U389 ( .A1(n436), .A2(n434), .S0(n277), .Y(n530) );
  MUX21X1_HVT U390 ( .A1(n366), .A2(n310), .S0(n371), .Y(n489) );
  MUX21X1_HVT U391 ( .A1(n310), .A2(n244), .S0(n247), .Y(n444) );
  MUX21X1_HVT U392 ( .A1(n310), .A2(n365), .S0(n370), .Y(n445) );
  MUX21X1_HVT U393 ( .A1(n354), .A2(n310), .S0(n247), .Y(n616) );
  NBUFFX2_HVT U394 ( .A(in[2]), .Y(n375) );
  NBUFFX2_HVT U395 ( .A(in[2]), .Y(n374) );
  MUX21X1_HVT U396 ( .A1(n611), .A2(n332), .S0(n342), .Y(n519) );
  MUX21X1_HVT U397 ( .A1(n329), .A2(n437), .S0(n276), .Y(n611) );
  MUX21X1_HVT U398 ( .A1(n350), .A2(n437), .S0(n370), .Y(n448) );
  MUX21X1_HVT U399 ( .A1(n362), .A2(n366), .S0(n291), .Y(n339) );
  MUX41X1_HVT U400 ( .A1(n477), .A3(n334), .A2(n331), .A4(n336), .S0(n293), 
        .S1(n311), .Y(n476) );
  MUX21X1_HVT U401 ( .A1(n326), .A2(n338), .S0(n277), .Y(n512) );
  XOR2X1_HVT U402 ( .A1(n276), .A2(n338), .Y(n595) );
  MUX21X1_HVT U403 ( .A1(n338), .A2(n317), .S0(n369), .Y(n619) );
  MUX21X1_HVT U404 ( .A1(n338), .A2(n362), .S0(n367), .Y(n451) );
  MUX21X1_HVT U405 ( .A1(n362), .A2(n338), .S0(n371), .Y(n447) );
  MUX21X1_HVT U406 ( .A1(n244), .A2(n338), .S0(n367), .Y(n614) );
  MUX21X1_HVT U407 ( .A1(n338), .A2(n434), .S0(n247), .Y(n452) );
  MUX21X1_HVT U408 ( .A1(n353), .A2(n329), .S0(n276), .Y(n617) );
  MUX21X1_HVT U409 ( .A1(n329), .A2(n353), .S0(n276), .Y(n450) );
  INVX1_HVT U410 ( .A(n448), .Y(n423) );
  MUX21X1_HVT U411 ( .A1(n350), .A2(n338), .S0(n368), .Y(n442) );
  MUX21X1_HVT U412 ( .A1(n338), .A2(n436), .S0(n368), .Y(n603) );
  INVX1_HVT U413 ( .A(in[4]), .Y(n380) );
  INVX0_HVT U414 ( .A(n632), .Y(n382) );
  INVX0_HVT U415 ( .A(n612), .Y(n383) );
  INVX0_HVT U416 ( .A(n606), .Y(n384) );
  INVX0_HVT U417 ( .A(n546), .Y(n385) );
  INVX0_HVT U418 ( .A(n507), .Y(n386) );
  INVX0_HVT U419 ( .A(n641), .Y(n387) );
  INVX0_HVT U420 ( .A(n630), .Y(n392) );
  INVX0_HVT U421 ( .A(n635), .Y(n393) );
  INVX0_HVT U422 ( .A(n631), .Y(n394) );
  INVX0_HVT U423 ( .A(n629), .Y(n395) );
  INVX0_HVT U424 ( .A(n628), .Y(n396) );
  INVX0_HVT U425 ( .A(n626), .Y(n397) );
  INVX0_HVT U426 ( .A(n625), .Y(n398) );
  INVX0_HVT U427 ( .A(n624), .Y(n399) );
  INVX0_HVT U428 ( .A(n623), .Y(n400) );
  INVX0_HVT U429 ( .A(n619), .Y(n403) );
  INVX0_HVT U430 ( .A(n618), .Y(n404) );
  INVX0_HVT U431 ( .A(n617), .Y(n405) );
  INVX0_HVT U432 ( .A(n616), .Y(n406) );
  INVX0_HVT U433 ( .A(n613), .Y(n409) );
  INVX0_HVT U434 ( .A(n610), .Y(n411) );
  INVX0_HVT U435 ( .A(n604), .Y(n414) );
  INVX0_HVT U436 ( .A(n599), .Y(n416) );
  INVX0_HVT U437 ( .A(n634), .Y(n418) );
  INVX0_HVT U438 ( .A(n451), .Y(n420) );
  INVX0_HVT U439 ( .A(n447), .Y(n424) );
  INVX0_HVT U440 ( .A(n445), .Y(n426) );
  INVX0_HVT U441 ( .A(n444), .Y(n427) );
  INVX0_HVT U442 ( .A(n443), .Y(n428) );
  INVX0_HVT U443 ( .A(n442), .Y(n429) );
  INVX0_HVT U444 ( .A(n489), .Y(n430) );
  INVX0_HVT U445 ( .A(n441), .Y(n431) );
  INVX0_HVT U446 ( .A(n439), .Y(n433) );
endmodule

