
module sbox_7 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n50, n99, n210, n211, n212, n213, n216, n217, n218, n219,
         n229, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674;

  NAND2X0_HVT U4 ( .A1(n293), .A2(n672), .Y(n671) );
  NAND2X0_HVT U5 ( .A1(n390), .A2(n372), .Y(n669) );
  NAND2X0_HVT U13 ( .A1(n661), .A2(n388), .Y(n662) );
  NAND2X0_HVT U15 ( .A1(n672), .A2(n374), .Y(n659) );
  NAND2X0_HVT U21 ( .A1(n294), .A2(n395), .Y(n653) );
  NAND2X0_HVT U24 ( .A1(n379), .A2(n395), .Y(n651) );
  NAND2X0_HVT U33 ( .A1(n291), .A2(n395), .Y(n642) );
  NAND2X0_HVT U35 ( .A1(n377), .A2(n395), .Y(n640) );
  NAND2X0_HVT U42 ( .A1(n391), .A2(n379), .Y(n633) );
  MUX41X1_HVT U51 ( .A1(n441), .A3(n405), .A2(n421), .A4(n219), .S0(n404), 
        .S1(n400), .Y(n626) );
  NAND2X0_HVT U53 ( .A1(n623), .A2(n632), .Y(n624) );
  NAND2X0_HVT U56 ( .A1(n293), .A2(n619), .Y(n620) );
  MUX41X1_HVT U57 ( .A1(n442), .A3(n655), .A2(n620), .A4(n664), .S0(n404), 
        .S1(n400), .Y(n618) );
  NAND2X0_HVT U58 ( .A1(n388), .A2(n672), .Y(n617) );
  NAND2X0_HVT U62 ( .A1(n395), .A2(n386), .Y(n613) );
  MUX41X1_HVT U63 ( .A1(n613), .A3(n412), .A2(n436), .A4(n333), .S0(n404), 
        .S1(n400), .Y(n612) );
  AO21X1_HVT U66 ( .A1(n285), .A2(n368), .A3(n435), .Y(n609) );
  MUX41X1_HVT U68 ( .A1(n415), .A3(n609), .A2(n608), .A4(n610), .S0(n367), 
        .S1(n403), .Y(n607) );
  MUX41X1_HVT U69 ( .A1(n607), .A3(n615), .A2(n611), .A4(n621), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n381), .A2(n602), .Y(n603) );
  MUX41X1_HVT U74 ( .A1(n604), .A3(n649), .A2(n603), .A4(n651), .S0(n365), 
        .S1(n402), .Y(n601) );
  AND3X1_HVT U80 ( .A1(n385), .A2(n619), .A3(n594), .Y(n595) );
  MUX41X1_HVT U82 ( .A1(n630), .A3(n219), .A2(n406), .A4(n660), .S0(in[2]), 
        .S1(n402), .Y(n592) );
  AND2X1_HVT U83 ( .A1(n389), .A2(n236), .Y(n591) );
  MUX41X1_HVT U84 ( .A1(n422), .A3(n308), .A2(n658), .A4(n591), .S0(n367), 
        .S1(n351), .Y(n590) );
  NAND2X0_HVT U85 ( .A1(n395), .A2(n455), .Y(n589) );
  MUX41X1_HVT U86 ( .A1(n444), .A3(n589), .A2(n358), .A4(n356), .S0(n366), 
        .S1(n402), .Y(n588) );
  AO21X1_HVT U93 ( .A1(n371), .A2(n581), .A3(n440), .Y(n582) );
  MUX41X1_HVT U97 ( .A1(n439), .A3(n359), .A2(n392), .A4(n659), .S0(n366), 
        .S1(n403), .Y(n578) );
  NAND2X0_HVT U101 ( .A1(n573), .A2(n572), .Y(n574) );
  MUX41X1_HVT U103 ( .A1(n672), .A3(n416), .A2(n265), .A4(n640), .S0(n398), 
        .S1(n403), .Y(n570) );
  MUX41X1_HVT U105 ( .A1(n424), .A3(n628), .A2(n569), .A4(n438), .S0(n367), 
        .S1(n402), .Y(n568) );
  MUX41X1_HVT U106 ( .A1(n568), .A3(n571), .A2(n570), .A4(n575), .S0(in[0]), 
        .S1(n400), .Y(n567) );
  OA21X1_HVT U109 ( .A1(n431), .A2(n399), .A3(n420), .Y(n565) );
  NAND2X0_HVT U110 ( .A1(n385), .A2(n563), .Y(n564) );
  MUX41X1_HVT U114 ( .A1(n560), .A3(n566), .A2(n562), .A4(n565), .S0(n368), 
        .S1(n351), .Y(n559) );
  AND2X1_HVT U115 ( .A1(n393), .A2(n374), .Y(n558) );
  MUX41X1_HVT U116 ( .A1(n662), .A3(n558), .A2(n316), .A4(n644), .S0(n364), 
        .S1(n404), .Y(n557) );
  AO21X1_HVT U118 ( .A1(n398), .A2(n380), .A3(n308), .Y(n555) );
  NAND2X0_HVT U123 ( .A1(n549), .A2(n548), .Y(n550) );
  MUX41X1_HVT U135 ( .A1(n449), .A3(n453), .A2(n669), .A4(n648), .S0(n365), 
        .S1(n351), .Y(n537) );
  MUX41X1_HVT U136 ( .A1(n356), .A3(n642), .A2(n450), .A4(n245), .S0(n364), 
        .S1(n404), .Y(n536) );
  MUX41X1_HVT U139 ( .A1(n534), .A3(n537), .A2(n536), .A4(n538), .S0(in[0]), 
        .S1(in[5]), .Y(n533) );
  AND2X1_HVT U140 ( .A1(n380), .A2(n394), .Y(n532) );
  NAND2X0_HVT U146 ( .A1(n390), .A2(n388), .Y(n602) );
  OA21X1_HVT U151 ( .A1(n341), .A2(n635), .A3(n522), .Y(n523) );
  MUX41X1_HVT U153 ( .A1(n564), .A3(n360), .A2(n386), .A4(n408), .S0(n364), 
        .S1(n403), .Y(n520) );
  AND2X1_HVT U154 ( .A1(n371), .A2(n379), .Y(n519) );
  NAND2X0_HVT U158 ( .A1(n314), .A2(n455), .Y(n515) );
  MUX41X1_HVT U159 ( .A1(n327), .A3(n375), .A2(n515), .A4(n414), .S0(n397), 
        .S1(n351), .Y(n514) );
  MUX41X1_HVT U160 ( .A1(n514), .A3(n520), .A2(n516), .A4(n521), .S0(in[0]), 
        .S1(in[5]), .Y(n513) );
  AND2X1_HVT U162 ( .A1(n308), .A2(n602), .Y(n511) );
  MUX41X1_HVT U163 ( .A1(n419), .A3(n511), .A2(n357), .A4(n512), .S0(n397), 
        .S1(n351), .Y(n510) );
  NAND2X0_HVT U166 ( .A1(n388), .A2(n619), .Y(n507) );
  NAND2X0_HVT U167 ( .A1(n456), .A2(n395), .Y(n506) );
  MUX41X1_HVT U168 ( .A1(n442), .A3(n380), .A2(n506), .A4(n507), .S0(n397), 
        .S1(n351), .Y(n505) );
  NAND2X0_HVT U174 ( .A1(n390), .A2(n668), .Y(n661) );
  MUX41X1_HVT U176 ( .A1(n324), .A3(n500), .A2(n447), .A4(n661), .S0(n404), 
        .S1(n397), .Y(n499) );
  NAND2X0_HVT U177 ( .A1(n393), .A2(n377), .Y(n498) );
  MUX41X1_HVT U178 ( .A1(n657), .A3(n498), .A2(n234), .A4(n637), .S0(n365), 
        .S1(n403), .Y(n497) );
  MUX41X1_HVT U179 ( .A1(n647), .A3(n451), .A2(n410), .A4(n234), .S0(n398), 
        .S1(n402), .Y(n496) );
  MUX41X1_HVT U180 ( .A1(n413), .A3(n666), .A2(n327), .A4(n355), .S0(n369), 
        .S1(n397), .Y(n495) );
  MUX41X1_HVT U181 ( .A1(n495), .A3(n497), .A2(n496), .A4(n499), .S0(in[0]), 
        .S1(in[5]), .Y(n494) );
  MUX41X1_HVT U182 ( .A1(n432), .A3(n294), .A2(n434), .A4(n423), .S0(n404), 
        .S1(n398), .Y(n493) );
  OA21X1_HVT U184 ( .A1(n641), .A2(n341), .A3(n422), .Y(n491) );
  MUX41X1_HVT U189 ( .A1(n487), .A3(n661), .A2(n488), .A4(n438), .S0(n369), 
        .S1(n398), .Y(n486) );
  MUX41X1_HVT U190 ( .A1(n486), .A3(n489), .A2(n490), .A4(n493), .S0(in[5]), 
        .S1(in[0]), .Y(n485) );
  MUX41X1_HVT U194 ( .A1(n634), .A3(n648), .A2(n449), .A4(n380), .S0(n369), 
        .S1(n398), .Y(n482) );
  AO21X1_HVT U197 ( .A1(n358), .A2(n370), .A3(n440), .Y(n479) );
  OA21X1_HVT U201 ( .A1(n667), .A2(n341), .A3(n258), .Y(n475) );
  MUX41X1_HVT U204 ( .A1(n620), .A3(n662), .A2(n429), .A4(n652), .S0(n398), 
        .S1(n402), .Y(n472) );
  MUX41X1_HVT U205 ( .A1(n236), .A3(n672), .A2(n451), .A4(n427), .S0(n397), 
        .S1(n403), .Y(n471) );
  NAND2X0_HVT U208 ( .A1(n389), .A2(n293), .Y(n563) );
  NAND2X0_HVT U212 ( .A1(n389), .A2(n381), .Y(n619) );
  NAND2X0_HVT U214 ( .A1(n308), .A2(n395), .Y(n469) );
  NAND2X0_HVT U215 ( .A1(n563), .A2(n382), .Y(n468) );
  NAND2X0_HVT U218 ( .A1(n453), .A2(n314), .Y(n522) );
  NAND2X0_HVT U220 ( .A1(n370), .A2(n469), .Y(n594) );
  IBUFFX2_HVT U1 ( .A(n389), .Y(n266) );
  INVX2_HVT U2 ( .A(n394), .Y(n389) );
  XOR2X1_HVT U3 ( .A1(n668), .A2(n392), .Y(n629) );
  IBUFFX2_HVT U6 ( .A(n394), .Y(n392) );
  AO21X2_HVT U7 ( .A1(n394), .A2(n453), .A3(n341), .Y(n573) );
  MUX21X1_HVT U8 ( .A1(n297), .A2(n387), .S0(n394), .Y(n296) );
  IBUFFX2_HVT U9 ( .A(n394), .Y(n390) );
  IBUFFX2_HVT U10 ( .A(n394), .Y(n393) );
  MUX41X2_HVT U11 ( .A1(n653), .A3(n363), .A2(n415), .A4(n448), .S0(n364), 
        .S1(n404), .Y(n546) );
  NAND2X0_HVT U12 ( .A1(n256), .A2(n257), .Y(out[1]) );
  OR2X1_HVT U14 ( .A1(n395), .A2(n23), .Y(n672) );
  IBUFFX16_HVT U16 ( .A(n384), .Y(n23) );
  IBUFFX2_HVT U17 ( .A(n390), .Y(n301) );
  NAND2X0_HVT U18 ( .A1(n554), .A2(n48), .Y(n50) );
  NAND2X0_HVT U19 ( .A1(n557), .A2(n243), .Y(n99) );
  NAND2X0_HVT U20 ( .A1(n50), .A2(n99), .Y(n553) );
  INVX0_HVT U22 ( .A(n243), .Y(n48) );
  INVX1_HVT U23 ( .A(n328), .Y(n243) );
  MUX21X1_HVT U25 ( .A1(n216), .A2(n633), .S0(n218), .Y(n217) );
  INVX1_HVT U26 ( .A(n216), .Y(n234) );
  INVX1_HVT U27 ( .A(n217), .Y(n480) );
  MUX41X1_HVT U28 ( .A1(n473), .A3(n474), .A2(n471), .A4(n472), .S0(n210), 
        .S1(n211), .Y(n470) );
  IBUFFX16_HVT U29 ( .A(n338), .Y(n210) );
  IBUFFX16_HVT U30 ( .A(n336), .Y(n211) );
  MUX41X1_HVT U31 ( .A1(n527), .A3(n526), .A2(n531), .A4(n530), .S0(n322), 
        .S1(n318), .Y(n525) );
  MUX41X2_HVT U32 ( .A1(n422), .A3(n375), .A2(n437), .A4(n380), .S0(n364), 
        .S1(n403), .Y(n530) );
  INVX1_HVT U34 ( .A(n321), .Y(n318) );
  IBUFFX2_HVT U36 ( .A(n400), .Y(n322) );
  MUX21X1_HVT U37 ( .A1(n539), .A2(n426), .S0(n260), .Y(n538) );
  MUX21X1_HVT U38 ( .A1(n386), .A2(n387), .S0(n313), .Y(n488) );
  INVX1_HVT U39 ( .A(n313), .Y(n314) );
  INVX0_HVT U40 ( .A(n258), .Y(n637) );
  MUX21X2_HVT U41 ( .A1(n645), .A2(n468), .S0(n369), .Y(n462) );
  MUX21X2_HVT U43 ( .A1(n427), .A2(n660), .S0(n365), .Y(n576) );
  MUX41X1_HVT U44 ( .A1(n433), .A3(n639), .A2(n643), .A4(n663), .S0(n212), 
        .S1(n213), .Y(n473) );
  IBUFFX16_HVT U45 ( .A(n397), .Y(n212) );
  IBUFFX16_HVT U46 ( .A(n320), .Y(n213) );
  OA21X2_HVT U47 ( .A1(n409), .A2(n341), .A3(n644), .Y(n528) );
  MUX21X1_HVT U48 ( .A1(n323), .A2(n381), .S0(n391), .Y(n216) );
  IBUFFX16_HVT U49 ( .A(n370), .Y(n218) );
  MUX21X2_HVT U50 ( .A1(n407), .A2(n552), .S0(n365), .Y(n551) );
  MUX21X1_HVT U52 ( .A1(n229), .A2(n324), .S0(n395), .Y(n219) );
  IBUFFX16_HVT U54 ( .A(n219), .Y(n654) );
  IBUFFX16_HVT U55 ( .A(n386), .Y(n229) );
  IBUFFX2_HVT U59 ( .A(n351), .Y(n238) );
  INVX1_HVT U60 ( .A(n320), .Y(n351) );
  OA21X2_HVT U61 ( .A1(n361), .A2(n341), .A3(n644), .Y(n503) );
  MUX21X2_HVT U64 ( .A1(n550), .A2(n551), .S0(n341), .Y(n547) );
  MUX21X1_HVT U65 ( .A1(n456), .A2(n455), .S0(n393), .Y(n648) );
  MUX21X2_HVT U67 ( .A1(n546), .A2(n547), .S0(n368), .Y(n545) );
  IBUFFX2_HVT U70 ( .A(n320), .Y(n403) );
  NAND2X0_HVT U71 ( .A1(n479), .A2(n231), .Y(n232) );
  NAND2X0_HVT U72 ( .A1(n480), .A2(n343), .Y(n233) );
  NAND2X0_HVT U75 ( .A1(n232), .A2(n233), .Y(n478) );
  IBUFFX2_HVT U76 ( .A(n343), .Y(n231) );
  IBUFFX2_HVT U77 ( .A(n643), .Y(n428) );
  MUX21X2_HVT U78 ( .A1(n382), .A2(n654), .S0(n278), .Y(n596) );
  IBUFFX2_HVT U79 ( .A(n389), .Y(n311) );
  MUX21X1_HVT U81 ( .A1(n350), .A2(n385), .S0(n389), .Y(n316) );
  MUX21X1_HVT U87 ( .A1(n373), .A2(n456), .S0(n389), .Y(n635) );
  MUX41X1_HVT U88 ( .A1(n545), .A3(n559), .A2(n540), .A4(n553), .S0(n235), 
        .S1(n346), .Y(out[3]) );
  IBUFFX16_HVT U89 ( .A(n352), .Y(n235) );
  INVX1_HVT U90 ( .A(n324), .Y(n236) );
  MUX21X2_HVT U91 ( .A1(n513), .A2(n501), .S0(n237), .Y(out[5]) );
  IBUFFX16_HVT U92 ( .A(in[6]), .Y(n237) );
  INVX0_HVT U94 ( .A(n316), .Y(n650) );
  MUX21X2_HVT U95 ( .A1(n523), .A2(n524), .S0(n366), .Y(n521) );
  NBUFFX2_HVT U96 ( .A(n673), .Y(n384) );
  MUX21X1_HVT U98 ( .A1(n582), .A2(n583), .S0(n366), .Y(n580) );
  INVX1_HVT U99 ( .A(n281), .Y(n584) );
  INVX0_HVT U100 ( .A(n639), .Y(n430) );
  MUX21X1_HVT U102 ( .A1(n374), .A2(n373), .S0(n393), .Y(n658) );
  MUX41X1_HVT U104 ( .A1(n627), .A3(n484), .A2(n633), .A4(n640), .S0(n398), 
        .S1(n238), .Y(n483) );
  INVX0_HVT U107 ( .A(n341), .Y(n329) );
  MUX21X2_HVT U108 ( .A1(n355), .A2(n658), .S0(n239), .Y(n476) );
  IBUFFX16_HVT U111 ( .A(n369), .Y(n239) );
  NAND2X0_HVT U112 ( .A1(n616), .A2(n240), .Y(n241) );
  NAND2X0_HVT U113 ( .A1(n618), .A2(n366), .Y(n242) );
  NAND2X0_HVT U117 ( .A1(n241), .A2(n242), .Y(n615) );
  IBUFFX2_HVT U119 ( .A(n366), .Y(n240) );
  INVX1_HVT U120 ( .A(n384), .Y(n456) );
  INVX1_HVT U121 ( .A(n670), .Y(n292) );
  MUX41X1_HVT U122 ( .A1(n316), .A3(n456), .A2(n444), .A4(n439), .S0(n244), 
        .S1(n320), .Y(n600) );
  IBUFFX16_HVT U124 ( .A(n366), .Y(n244) );
  INVX0_HVT U125 ( .A(n430), .Y(n245) );
  MUX41X1_HVT U126 ( .A1(n605), .A3(n600), .A2(n601), .A4(n598), .S0(n246), 
        .S1(n247), .Y(n597) );
  IBUFFX16_HVT U127 ( .A(in[0]), .Y(n246) );
  IBUFFX16_HVT U128 ( .A(n401), .Y(n247) );
  NBUFFX2_HVT U129 ( .A(n648), .Y(n248) );
  NAND2X0_HVT U130 ( .A1(n533), .A2(n249), .Y(n250) );
  NAND2X0_HVT U131 ( .A1(n525), .A2(n332), .Y(n251) );
  NAND2X0_HVT U132 ( .A1(n250), .A2(n251), .Y(out[4]) );
  INVX1_HVT U133 ( .A(n332), .Y(n249) );
  IBUFFX2_HVT U134 ( .A(in[6]), .Y(n332) );
  NAND2X0_HVT U137 ( .A1(n567), .A2(n252), .Y(n253) );
  NAND2X0_HVT U138 ( .A1(n577), .A2(in[6]), .Y(n254) );
  NAND2X0_HVT U141 ( .A1(n253), .A2(n254), .Y(out[2]) );
  IBUFFX2_HVT U142 ( .A(in[6]), .Y(n252) );
  NAND2X0_HVT U143 ( .A1(n587), .A2(n255), .Y(n256) );
  NAND2X0_HVT U144 ( .A1(n597), .A2(in[6]), .Y(n257) );
  IBUFFX2_HVT U145 ( .A(in[6]), .Y(n255) );
  IBUFFX2_HVT U147 ( .A(n563), .Y(n437) );
  MUX21X1_HVT U148 ( .A1(n387), .A2(n288), .S0(n391), .Y(n258) );
  INVX0_HVT U149 ( .A(n288), .Y(n290) );
  MUX21X2_HVT U150 ( .A1(n395), .A2(n417), .S0(n259), .Y(n610) );
  IBUFFX16_HVT U152 ( .A(n368), .Y(n259) );
  INVX0_HVT U155 ( .A(n461), .Y(n448) );
  IBUFFX16_HVT U156 ( .A(n367), .Y(n260) );
  IBUFFX16_HVT U157 ( .A(n394), .Y(n391) );
  INVX1_HVT U161 ( .A(n462), .Y(n426) );
  MUX21X2_HVT U164 ( .A1(n596), .A2(n595), .S0(n365), .Y(n593) );
  MUX21X1_HVT U165 ( .A1(n446), .A2(n637), .S0(n261), .Y(n517) );
  IBUFFX16_HVT U169 ( .A(n369), .Y(n261) );
  INVX1_HVT U170 ( .A(n262), .Y(n539) );
  MUX21X1_HVT U171 ( .A1(n263), .A2(n461), .S0(n264), .Y(n262) );
  IBUFFX16_HVT U172 ( .A(n382), .Y(n263) );
  IBUFFX16_HVT U173 ( .A(n370), .Y(n264) );
  INVX1_HVT U175 ( .A(n296), .Y(n641) );
  INVX0_HVT U183 ( .A(n658), .Y(n418) );
  MUX21X1_HVT U185 ( .A1(n288), .A2(n323), .S0(n266), .Y(n265) );
  INVX8_HVT U186 ( .A(n265), .Y(n646) );
  NAND2X0_HVT U187 ( .A1(n606), .A2(n267), .Y(n268) );
  NAND2X0_HVT U188 ( .A1(n631), .A2(n276), .Y(n269) );
  NAND2X0_HVT U191 ( .A1(n268), .A2(n269), .Y(n605) );
  INVX0_HVT U192 ( .A(n276), .Y(n267) );
  XOR2X1_HVT U193 ( .A1(n248), .A2(n341), .Y(n631) );
  IBUFFX2_HVT U195 ( .A(n366), .Y(n276) );
  NAND2X0_HVT U196 ( .A1(n671), .A2(n270), .Y(n271) );
  NAND2X0_HVT U198 ( .A1(n535), .A2(n284), .Y(n272) );
  NAND2X0_HVT U199 ( .A1(n271), .A2(n272), .Y(n534) );
  INVX0_HVT U200 ( .A(n284), .Y(n270) );
  NAND2X0_HVT U202 ( .A1(n379), .A2(n273), .Y(n274) );
  NAND2X0_HVT U203 ( .A1(n375), .A2(n280), .Y(n275) );
  NAND2X0_HVT U206 ( .A1(n274), .A2(n275), .Y(n652) );
  IBUFFX4_HVT U207 ( .A(n280), .Y(n273) );
  IBUFFX2_HVT U209 ( .A(n398), .Y(n284) );
  IBUFFX2_HVT U210 ( .A(n389), .Y(n280) );
  INVX0_HVT U211 ( .A(n652), .Y(n422) );
  MUX21X2_HVT U213 ( .A1(n646), .A2(n411), .S0(n371), .Y(n529) );
  INVX1_HVT U216 ( .A(n309), .Y(n599) );
  MUX21X2_HVT U217 ( .A1(n529), .A2(n528), .S0(n367), .Y(n527) );
  MUX21X2_HVT U219 ( .A1(n518), .A2(n517), .S0(n277), .Y(n516) );
  IBUFFX16_HVT U221 ( .A(n367), .Y(n277) );
  IBUFFX16_HVT U222 ( .A(n371), .Y(n278) );
  MUX21X2_HVT U223 ( .A1(n432), .A2(n652), .S0(n279), .Y(n535) );
  IBUFFX16_HVT U224 ( .A(n370), .Y(n279) );
  INVX0_HVT U225 ( .A(n392), .Y(n287) );
  INVX1_HVT U226 ( .A(n285), .Y(n664) );
  MUX21X1_HVT U227 ( .A1(n323), .A2(n282), .S0(n283), .Y(n281) );
  IBUFFX16_HVT U228 ( .A(n379), .Y(n282) );
  IBUFFX16_HVT U229 ( .A(n371), .Y(n283) );
  INVX1_HVT U230 ( .A(n323), .Y(n324) );
  IBUFFX2_HVT U231 ( .A(n672), .Y(n411) );
  MUX21X2_HVT U232 ( .A1(n574), .A2(n426), .S0(n367), .Y(n571) );
  MUX21X1_HVT U233 ( .A1(n387), .A2(n286), .S0(n287), .Y(n285) );
  IBUFFX16_HVT U234 ( .A(n373), .Y(n286) );
  INVX2_HVT U235 ( .A(n292), .Y(n293) );
  INVX1_HVT U236 ( .A(n452), .Y(n288) );
  INVX0_HVT U237 ( .A(n452), .Y(n289) );
  INVX1_HVT U238 ( .A(n289), .Y(n291) );
  INVX1_HVT U239 ( .A(n292), .Y(n294) );
  MUX21X2_HVT U240 ( .A1(n386), .A2(n584), .S0(n362), .Y(n583) );
  IBUFFX2_HVT U241 ( .A(n324), .Y(n310) );
  MUX41X1_HVT U242 ( .A1(n420), .A3(n361), .A2(n617), .A4(n363), .S0(n320), 
        .S1(n295), .Y(n616) );
  IBUFFX16_HVT U243 ( .A(n400), .Y(n295) );
  IBUFFX2_HVT U244 ( .A(n320), .Y(n404) );
  INVX1_HVT U245 ( .A(n656), .Y(n420) );
  INVX1_HVT U246 ( .A(n302), .Y(n579) );
  INVX0_HVT U247 ( .A(n381), .Y(n335) );
  INVX0_HVT U248 ( .A(n333), .Y(n660) );
  IBUFFX16_HVT U249 ( .A(n372), .Y(n297) );
  MUX21X2_HVT U250 ( .A1(n492), .A2(n491), .S0(n298), .Y(n490) );
  IBUFFX16_HVT U251 ( .A(n366), .Y(n298) );
  MUX21X1_HVT U252 ( .A1(n293), .A2(n300), .S0(n301), .Y(n299) );
  IBUFFX16_HVT U253 ( .A(n374), .Y(n300) );
  MUX41X1_HVT U254 ( .A1(n299), .A3(n305), .A2(n304), .A4(n303), .S0(n306), 
        .S1(n312), .Y(n302) );
  IBUFFX16_HVT U255 ( .A(n406), .Y(n303) );
  IBUFFX16_HVT U256 ( .A(n359), .Y(n304) );
  IBUFFX16_HVT U257 ( .A(n443), .Y(n305) );
  IBUFFX16_HVT U258 ( .A(in[2]), .Y(n306) );
  INVX2_HVT U259 ( .A(n312), .Y(n402) );
  INVX0_HVT U260 ( .A(n369), .Y(n312) );
  INVX0_HVT U261 ( .A(n668), .Y(n307) );
  INVX1_HVT U262 ( .A(n307), .Y(n308) );
  INVX1_HVT U263 ( .A(n350), .Y(n668) );
  MUX21X1_HVT U264 ( .A1(n310), .A2(n350), .S0(n311), .Y(n309) );
  MUX41X1_HVT U265 ( .A1(n445), .A3(n599), .A2(n446), .A4(n666), .S0(n312), 
        .S1(n399), .Y(n598) );
  INVX0_HVT U266 ( .A(in[7]), .Y(n320) );
  INVX0_HVT U267 ( .A(n380), .Y(n453) );
  INVX0_HVT U268 ( .A(n389), .Y(n313) );
  INVX0_HVT U269 ( .A(n384), .Y(n334) );
  MUX41X1_HVT U270 ( .A1(n544), .A3(n542), .A2(n543), .A4(n541), .S0(n315), 
        .S1(n312), .Y(n540) );
  IBUFFX16_HVT U271 ( .A(n368), .Y(n315) );
  MUX41X1_HVT U272 ( .A1(n428), .A3(n532), .A2(n258), .A4(n650), .S0(n317), 
        .S1(n341), .Y(n531) );
  IBUFFX16_HVT U273 ( .A(n365), .Y(n317) );
  MUX41X1_HVT U274 ( .A1(n629), .A3(n439), .A2(n602), .A4(n450), .S0(n319), 
        .S1(n320), .Y(n526) );
  IBUFFX16_HVT U275 ( .A(n365), .Y(n319) );
  IBUFFX16_HVT U276 ( .A(in[0]), .Y(n321) );
  INVX1_HVT U277 ( .A(n377), .Y(n323) );
  INVX1_HVT U278 ( .A(n383), .Y(n452) );
  MUX41X1_HVT U279 ( .A1(n441), .A3(n586), .A2(n629), .A4(n633), .S0(n364), 
        .S1(n312), .Y(n585) );
  MUX41X1_HVT U280 ( .A1(n585), .A3(n579), .A2(n580), .A4(n578), .S0(n325), 
        .S1(n326), .Y(n577) );
  IBUFFX16_HVT U281 ( .A(in[0]), .Y(n325) );
  IBUFFX16_HVT U282 ( .A(n401), .Y(n326) );
  INVX0_HVT U283 ( .A(n436), .Y(n327) );
  IBUFFX16_HVT U284 ( .A(n368), .Y(n328) );
  MUX41X1_HVT U285 ( .A1(n636), .A3(n359), .A2(n629), .A4(n602), .S0(n399), 
        .S1(n329), .Y(n489) );
  MUX41X1_HVT U286 ( .A1(n510), .A3(n505), .A2(n508), .A4(n502), .S0(n330), 
        .S1(n331), .Y(n501) );
  IBUFFX16_HVT U287 ( .A(in[0]), .Y(n330) );
  IBUFFX16_HVT U288 ( .A(n400), .Y(n331) );
  MUX21X1_HVT U289 ( .A1(n335), .A2(n334), .S0(n395), .Y(n333) );
  IBUFFX16_HVT U290 ( .A(n346), .Y(n336) );
  INVX2_HVT U291 ( .A(in[1]), .Y(n394) );
  MUX41X1_HVT U292 ( .A1(n629), .A3(n509), .A2(n653), .A4(n425), .S0(n404), 
        .S1(n337), .Y(n508) );
  IBUFFX16_HVT U293 ( .A(n398), .Y(n337) );
  NAND2X0_HVT U294 ( .A1(n349), .A2(n348), .Y(out[7]) );
  INVX0_HVT U295 ( .A(n352), .Y(n347) );
  MUX21X1_HVT U296 ( .A1(n375), .A2(n455), .S0(n393), .Y(n667) );
  NBUFFX2_HVT U297 ( .A(n396), .Y(n364) );
  INVX1_HVT U298 ( .A(in[0]), .Y(n346) );
  INVX1_HVT U299 ( .A(n371), .Y(n341) );
  NBUFFX2_HVT U300 ( .A(n350), .Y(n374) );
  INVX1_HVT U301 ( .A(n400), .Y(n338) );
  INVX0_HVT U302 ( .A(n366), .Y(n343) );
  INVX1_HVT U303 ( .A(n399), .Y(n396) );
  MUX41X1_HVT U304 ( .A1(n593), .A3(n590), .A2(n592), .A4(n588), .S0(n346), 
        .S1(n338), .Y(n587) );
  IBUFFX2_HVT U305 ( .A(in[1]), .Y(n395) );
  NAND2X0_HVT U306 ( .A1(n614), .A2(n366), .Y(n339) );
  NAND2X0_HVT U307 ( .A1(n612), .A2(n343), .Y(n340) );
  NAND2X0_HVT U308 ( .A1(n339), .A2(n340), .Y(n611) );
  MUX41X1_HVT U309 ( .A1(n360), .A3(n419), .A2(n418), .A4(n374), .S0(n404), 
        .S1(in[5]), .Y(n614) );
  INVX1_HVT U310 ( .A(n463), .Y(n445) );
  INVX1_HVT U311 ( .A(n342), .Y(n524) );
  MUX21X1_HVT U312 ( .A1(n380), .A2(n463), .S0(n341), .Y(n342) );
  NAND2X0_HVT U313 ( .A1(n475), .A2(n343), .Y(n344) );
  NAND2X0_HVT U314 ( .A1(n476), .A2(n366), .Y(n345) );
  NAND2X0_HVT U315 ( .A1(n344), .A2(n345), .Y(n474) );
  NAND2X0_HVT U316 ( .A1(n477), .A2(n347), .Y(n348) );
  NAND2X0_HVT U317 ( .A1(n470), .A2(n352), .Y(n349) );
  INVX0_HVT U318 ( .A(in[6]), .Y(n352) );
  XNOR2X2_HVT U319 ( .A1(n457), .A2(n378), .Y(n350) );
  INVX1_HVT U320 ( .A(in[2]), .Y(n399) );
  XNOR2X1_HVT U321 ( .A1(n397), .A2(n351), .Y(n353) );
  MUX21X1_HVT U322 ( .A1(n385), .A2(n561), .S0(n354), .Y(n560) );
  MUX41X1_HVT U323 ( .A1(n443), .A3(n308), .A2(n638), .A4(n387), .S0(n399), 
        .S1(n402), .Y(n481) );
  IBUFFX2_HVT U324 ( .A(n399), .Y(n398) );
  AND3X2_HVT U325 ( .A1(n367), .A2(n395), .A3(n236), .Y(n543) );
  XNOR2X1_HVT U326 ( .A1(n314), .A2(n396), .Y(n354) );
  MUX41X1_HVT U327 ( .A1(n483), .A3(n481), .A2(n482), .A4(n478), .S0(n346), 
        .S1(n338), .Y(n477) );
  MUX21X2_HVT U328 ( .A1(n576), .A2(n360), .S0(n353), .Y(n575) );
  INVX0_HVT U329 ( .A(n378), .Y(n454) );
  MUX21X2_HVT U330 ( .A1(n485), .A2(n494), .S0(in[6]), .Y(out[6]) );
  MUX21X2_HVT U331 ( .A1(n622), .A2(n626), .S0(n367), .Y(n621) );
  INVX0_HVT U332 ( .A(n399), .Y(n397) );
  NBUFFX2_HVT U333 ( .A(n350), .Y(n375) );
  MUX21X1_HVT U334 ( .A1(n357), .A2(n418), .S0(n364), .Y(n542) );
  AND2X1_HVT U335 ( .A1(n375), .A2(n619), .Y(n355) );
  NBUFFX2_HVT U336 ( .A(n670), .Y(n383) );
  MUX21X1_HVT U337 ( .A1(n290), .A2(n455), .S0(n368), .Y(n623) );
  MUX21X1_HVT U338 ( .A1(n644), .A2(n564), .S0(n364), .Y(n562) );
  MUX21X1_HVT U339 ( .A1(n416), .A2(n453), .S0(n368), .Y(n608) );
  AND2X1_HVT U340 ( .A1(n385), .A2(n602), .Y(n356) );
  MUX21X1_HVT U341 ( .A1(n386), .A2(n374), .S0(n391), .Y(n634) );
  MUX21X1_HVT U342 ( .A1(n294), .A2(n668), .S0(n393), .Y(n638) );
  MUX21X1_HVT U343 ( .A1(n375), .A2(n377), .S0(n389), .Y(n572) );
  MUX21X1_HVT U344 ( .A1(n290), .A2(n456), .S0(n392), .Y(n500) );
  NAND2X0_HVT U345 ( .A1(n376), .A2(n454), .Y(n670) );
  MUX21X1_HVT U346 ( .A1(n308), .A2(n453), .S0(n393), .Y(n460) );
  MUX21X1_HVT U347 ( .A1(n455), .A2(n374), .S0(n314), .Y(n512) );
  MUX21X1_HVT U348 ( .A1(n294), .A2(n382), .S0(n390), .Y(n586) );
  INVX1_HVT U349 ( .A(n387), .Y(n455) );
  MUX21X1_HVT U350 ( .A1(n555), .A2(n556), .S0(n370), .Y(n554) );
  MUX21X1_HVT U351 ( .A1(n408), .A2(n429), .S0(n364), .Y(n556) );
  NBUFFX2_HVT U352 ( .A(n384), .Y(n385) );
  MUX21X1_HVT U353 ( .A1(n372), .A2(n377), .S0(n392), .Y(n484) );
  XOR2X1_HVT U354 ( .A1(n385), .A2(n392), .Y(n627) );
  MUX21X1_HVT U355 ( .A1(n291), .A2(n324), .S0(n391), .Y(n461) );
  MUX21X1_HVT U356 ( .A1(n373), .A2(n668), .S0(n391), .Y(n463) );
  MUX21X1_HVT U357 ( .A1(n293), .A2(n372), .S0(n393), .Y(n663) );
  MUX21X1_HVT U358 ( .A1(n377), .A2(n373), .S0(n391), .Y(n552) );
  MUX21X1_HVT U359 ( .A1(n372), .A2(n388), .S0(n391), .Y(n487) );
  MUX21X1_HVT U360 ( .A1(n335), .A2(n291), .S0(n392), .Y(n656) );
  MUX21X1_HVT U361 ( .A1(n387), .A2(n381), .S0(n390), .Y(n644) );
  MUX21X1_HVT U362 ( .A1(n294), .A2(n388), .S0(n392), .Y(n581) );
  NBUFFX2_HVT U363 ( .A(n673), .Y(n386) );
  XOR2X1_HVT U364 ( .A1(n314), .A2(n335), .Y(n630) );
  XNOR2X1_HVT U365 ( .A1(n293), .A2(n390), .Y(n357) );
  XNOR2X1_HVT U366 ( .A1(n387), .A2(n390), .Y(n358) );
  AND2X1_HVT U367 ( .A1(n391), .A2(n456), .Y(n359) );
  MUX21X1_HVT U368 ( .A1(n381), .A2(n372), .S0(n389), .Y(n465) );
  MUX21X1_HVT U369 ( .A1(n386), .A2(n324), .S0(n390), .Y(n467) );
  MUX21X1_HVT U370 ( .A1(n386), .A2(n294), .S0(n392), .Y(n459) );
  AND2X1_HVT U371 ( .A1(n388), .A2(n563), .Y(n360) );
  MUX21X1_HVT U372 ( .A1(n382), .A2(n377), .S0(n390), .Y(n604) );
  MUX21X1_HVT U373 ( .A1(n382), .A2(n388), .S0(n367), .Y(n549) );
  XOR2X1_HVT U374 ( .A1(n377), .A2(n393), .Y(n649) );
  NBUFFX2_HVT U375 ( .A(in[7]), .Y(n370) );
  NBUFFX2_HVT U376 ( .A(in[7]), .Y(n369) );
  NBUFFX2_HVT U377 ( .A(in[7]), .Y(n371) );
  NBUFFX2_HVT U378 ( .A(n454), .Y(n373) );
  NBUFFX2_HVT U379 ( .A(n454), .Y(n372) );
  NBUFFX2_HVT U380 ( .A(n401), .Y(n368) );
  NBUFFX2_HVT U381 ( .A(n396), .Y(n366) );
  NBUFFX2_HVT U382 ( .A(n396), .Y(n365) );
  NBUFFX2_HVT U383 ( .A(n396), .Y(n367) );
  MUX21X1_HVT U384 ( .A1(n589), .A2(n379), .S0(n370), .Y(n492) );
  XOR2X1_HVT U385 ( .A1(n392), .A2(n378), .Y(n628) );
  MUX21X1_HVT U386 ( .A1(n381), .A2(n375), .S0(n314), .Y(n569) );
  NAND2X0_HVT U387 ( .A1(n378), .A2(n376), .Y(n673) );
  NBUFFX2_HVT U388 ( .A(n376), .Y(n377) );
  AND2X1_HVT U389 ( .A1(n375), .A2(n395), .Y(n361) );
  NBUFFX2_HVT U390 ( .A(n674), .Y(n387) );
  NBUFFX2_HVT U391 ( .A(n665), .Y(n380) );
  MUX21X1_HVT U392 ( .A1(n379), .A2(n291), .S0(n393), .Y(n636) );
  MUX21X1_HVT U393 ( .A1(n455), .A2(n443), .S0(n371), .Y(n606) );
  MUX21X1_HVT U394 ( .A1(n504), .A2(n503), .S0(n367), .Y(n502) );
  MUX21X1_HVT U395 ( .A1(n382), .A2(n443), .S0(n371), .Y(n504) );
  MUX21X1_HVT U396 ( .A1(n334), .A2(n379), .S0(n391), .Y(n655) );
  MUX21X1_HVT U397 ( .A1(n430), .A2(n672), .S0(n365), .Y(n566) );
  MUX21X1_HVT U398 ( .A1(n657), .A2(n428), .S0(n365), .Y(n541) );
  MUX21X1_HVT U399 ( .A1(n672), .A2(n394), .S0(n366), .Y(n548) );
  MUX21X1_HVT U400 ( .A1(n453), .A2(n456), .S0(n390), .Y(n509) );
  NBUFFX2_HVT U401 ( .A(n665), .Y(n381) );
  MUX21X1_HVT U402 ( .A1(n519), .A2(n385), .S0(n362), .Y(n518) );
  MUX21X1_HVT U403 ( .A1(n624), .A2(n625), .S0(n369), .Y(n622) );
  MUX21X1_HVT U404 ( .A1(n379), .A2(n640), .S0(n368), .Y(n625) );
  XOR2X1_HVT U405 ( .A1(n389), .A2(n401), .Y(n632) );
  MUX21X1_HVT U406 ( .A1(n379), .A2(n335), .S0(n393), .Y(n464) );
  NBUFFX2_HVT U407 ( .A(n674), .Y(n388) );
  MUX21X1_HVT U408 ( .A1(n293), .A2(n379), .S0(n390), .Y(n666) );
  MUX21X1_HVT U409 ( .A1(n424), .A2(n645), .S0(n365), .Y(n544) );
  NBUFFX2_HVT U410 ( .A(n457), .Y(n376) );
  NBUFFX2_HVT U411 ( .A(n665), .Y(n382) );
  XNOR2X1_HVT U412 ( .A1(n341), .A2(n392), .Y(n362) );
  AND2X1_HVT U413 ( .A1(n373), .A2(n395), .Y(n363) );
  NBUFFX2_HVT U414 ( .A(in[5]), .Y(n401) );
  NBUFFX2_HVT U415 ( .A(in[5]), .Y(n400) );
  INVX0_HVT U416 ( .A(in[4]), .Y(n457) );
  MUX21X1_HVT U417 ( .A1(n290), .A2(n236), .S0(n391), .Y(n643) );
  NAND2X0_HVT U418 ( .A1(in[4]), .A2(n454), .Y(n665) );
  NAND2X0_HVT U419 ( .A1(n378), .A2(in[4]), .Y(n674) );
  MUX21X1_HVT U420 ( .A1(n236), .A2(n455), .S0(n393), .Y(n639) );
  MUX21X1_HVT U421 ( .A1(n236), .A2(n668), .S0(n391), .Y(n466) );
  MUX21X1_HVT U422 ( .A1(n236), .A2(n335), .S0(n389), .Y(n657) );
  MUX21X1_HVT U423 ( .A1(n236), .A2(n388), .S0(n314), .Y(n458) );
  MUX21X1_HVT U424 ( .A1(n388), .A2(n236), .S0(n392), .Y(n647) );
  MUX21X1_HVT U425 ( .A1(n379), .A2(n236), .S0(n364), .Y(n561) );
  MUX21X1_HVT U426 ( .A1(n372), .A2(n236), .S0(n391), .Y(n645) );
  NBUFFX2_HVT U427 ( .A(in[3]), .Y(n378) );
  NBUFFX2_HVT U428 ( .A(in[3]), .Y(n379) );
  INVX0_HVT U429 ( .A(n653), .Y(n405) );
  INVX0_HVT U430 ( .A(n651), .Y(n406) );
  INVX0_HVT U431 ( .A(n642), .Y(n407) );
  INVX0_HVT U432 ( .A(n640), .Y(n408) );
  INVX0_HVT U433 ( .A(n506), .Y(n409) );
  INVX0_HVT U434 ( .A(n469), .Y(n410) );
  INVX0_HVT U435 ( .A(n659), .Y(n412) );
  INVX0_HVT U436 ( .A(n671), .Y(n413) );
  INVX0_HVT U437 ( .A(n669), .Y(n414) );
  INVX0_HVT U438 ( .A(n667), .Y(n415) );
  INVX0_HVT U439 ( .A(n666), .Y(n416) );
  INVX0_HVT U440 ( .A(n663), .Y(n417) );
  INVX0_HVT U441 ( .A(n657), .Y(n419) );
  INVX0_HVT U442 ( .A(n655), .Y(n421) );
  INVX0_HVT U443 ( .A(n649), .Y(n423) );
  INVX0_HVT U444 ( .A(n647), .Y(n424) );
  INVX0_HVT U445 ( .A(n645), .Y(n425) );
  INVX0_HVT U446 ( .A(n644), .Y(n427) );
  INVX0_HVT U447 ( .A(n641), .Y(n429) );
  INVX0_HVT U448 ( .A(n638), .Y(n431) );
  INVX0_HVT U449 ( .A(n636), .Y(n432) );
  INVX0_HVT U450 ( .A(n635), .Y(n433) );
  INVX0_HVT U451 ( .A(n634), .Y(n434) );
  INVX0_HVT U452 ( .A(n602), .Y(n435) );
  INVX0_HVT U453 ( .A(n662), .Y(n436) );
  INVX0_HVT U454 ( .A(n468), .Y(n438) );
  INVX0_HVT U455 ( .A(n619), .Y(n439) );
  INVX0_HVT U456 ( .A(n522), .Y(n440) );
  INVX0_HVT U457 ( .A(n467), .Y(n441) );
  INVX0_HVT U458 ( .A(n466), .Y(n442) );
  INVX0_HVT U459 ( .A(n465), .Y(n443) );
  INVX0_HVT U460 ( .A(n464), .Y(n444) );
  INVX0_HVT U461 ( .A(n581), .Y(n446) );
  INVX0_HVT U462 ( .A(n572), .Y(n447) );
  INVX0_HVT U463 ( .A(n460), .Y(n449) );
  INVX0_HVT U464 ( .A(n459), .Y(n450) );
  INVX0_HVT U465 ( .A(n458), .Y(n451) );
endmodule

