
module sbox_6 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n5, n23, n28, n47, n50, n114, n117, n118, n119, n210, n211, n212,
         n213, n216, n217, n218, n219, n224, n226, n227, n228, n229, n231,
         n232, n236, n238, n241, n252, n253, n259, n261, n264, n267, n274,
         n275, n276, n278, n279, n280, n282, n283, n284, n289, n290, n293,
         n295, n296, n297, n299, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790;

  NAND2X0_HVT U4 ( .A1(n409), .A2(n788), .Y(n787) );
  NAND2X0_HVT U5 ( .A1(n306), .A2(n520), .Y(n786) );
  NAND2X0_HVT U15 ( .A1(n788), .A2(n373), .Y(n776) );
  NAND2X0_HVT U21 ( .A1(n409), .A2(n391), .Y(n770) );
  NAND2X0_HVT U24 ( .A1(n456), .A2(n391), .Y(n768) );
  NAND2X0_HVT U33 ( .A1(n331), .A2(n391), .Y(n760) );
  NAND2X0_HVT U42 ( .A1(n306), .A2(n456), .Y(n751) );
  MUX41X1_HVT U51 ( .A1(n542), .A3(n561), .A2(n539), .A4(n544), .S0(n489), 
        .S1(n508), .Y(n744) );
  NAND2X0_HVT U53 ( .A1(n741), .A2(n750), .Y(n742) );
  NAND2X0_HVT U56 ( .A1(n409), .A2(n737), .Y(n738) );
  NAND2X0_HVT U58 ( .A1(n334), .A2(n788), .Y(n735) );
  MUX41X1_HVT U59 ( .A1(n498), .A3(n735), .A2(n496), .A4(n551), .S0(n488), 
        .S1(n508), .Y(n734) );
  MUX41X1_HVT U61 ( .A1(n492), .A3(n569), .A2(n548), .A4(n382), .S0(n488), 
        .S1(n508), .Y(n732) );
  NAND2X0_HVT U62 ( .A1(n450), .A2(n310), .Y(n731) );
  AO21X1_HVT U66 ( .A1(n576), .A2(n531), .A3(n578), .Y(n727) );
  NAND2X0_HVT U73 ( .A1(n386), .A2(n720), .Y(n721) );
  MUX41X1_HVT U74 ( .A1(n722), .A3(n766), .A2(n721), .A4(n768), .S0(n259), 
        .S1(n321), .Y(n719) );
  MUX41X1_HVT U77 ( .A1(n783), .A3(n558), .A2(n717), .A4(n47), .S0(n511), .S1(
        n507), .Y(n716) );
  MUX41X1_HVT U82 ( .A1(n748), .A3(n544), .A2(n582), .A4(n777), .S0(n259), 
        .S1(n489), .Y(n710) );
  AND2X1_HVT U83 ( .A1(n526), .A2(n411), .Y(n709) );
  MUX41X1_HVT U84 ( .A1(n5), .A3(n390), .A2(n775), .A4(n709), .S0(n259), .S1(
        n535), .Y(n708) );
  NAND2X0_HVT U85 ( .A1(n328), .A2(n449), .Y(n707) );
  MUX41X1_HVT U96 ( .A1(n582), .A3(n495), .A2(n573), .A4(n697), .S0(n401), 
        .S1(n485), .Y(n696) );
  NAND2X0_HVT U101 ( .A1(n690), .A2(n689), .Y(n691) );
  MUX41X1_HVT U103 ( .A1(n788), .A3(n562), .A2(n552), .A4(n758), .S0(n363), 
        .S1(n512), .Y(n687) );
  MUX41X1_HVT U105 ( .A1(n568), .A3(n746), .A2(n686), .A4(n560), .S0(n363), 
        .S1(n485), .Y(n685) );
  NAND2X0_HVT U110 ( .A1(n524), .A2(n681), .Y(n682) );
  AND2X1_HVT U115 ( .A1(n347), .A2(n373), .Y(n679) );
  NAND2X0_HVT U123 ( .A1(n670), .A2(n669), .Y(n671) );
  MUX41X1_HVT U131 ( .A1(n662), .A3(n664), .A2(n663), .A4(n665), .S0(n509), 
        .S1(n488), .Y(n661) );
  MUX41X1_HVT U135 ( .A1(n23), .A3(n315), .A2(n786), .A4(n427), .S0(n264), 
        .S1(n487), .Y(n658) );
  MUX41X1_HVT U136 ( .A1(n491), .A3(n760), .A2(n28), .A4(n757), .S0(n264), 
        .S1(n488), .Y(n657) );
  AND2X1_HVT U140 ( .A1(n359), .A2(n328), .Y(n653) );
  MUX41X1_HVT U141 ( .A1(n767), .A3(n555), .A2(n653), .A4(n553), .S0(n264), 
        .S1(n487), .Y(n652) );
  MUX41X1_HVT U142 ( .A1(n5), .A3(n382), .A2(n559), .A4(n359), .S0(n416), .S1(
        n487), .Y(n651) );
  MUX41X1_HVT U153 ( .A1(n682), .A3(n492), .A2(n310), .A4(n564), .S0(n335), 
        .S1(n536), .Y(n641) );
  AND2X1_HVT U154 ( .A1(n512), .A2(n407), .Y(n640) );
  NAND2X0_HVT U158 ( .A1(n413), .A2(n449), .Y(n636) );
  MUX41X1_HVT U159 ( .A1(n779), .A3(n373), .A2(n636), .A4(n579), .S0(n264), 
        .S1(n535), .Y(n635) );
  AND2X1_HVT U162 ( .A1(n785), .A2(n720), .Y(n632) );
  MUX41X1_HVT U165 ( .A1(n770), .A3(n567), .A2(n398), .A4(n630), .S0(n489), 
        .S1(n506), .Y(n629) );
  NAND2X0_HVT U166 ( .A1(n336), .A2(n737), .Y(n628) );
  NAND2X0_HVT U167 ( .A1(n311), .A2(n328), .Y(n627) );
  MUX41X1_HVT U168 ( .A1(n550), .A3(n386), .A2(n627), .A4(n628), .S0(n416), 
        .S1(n535), .Y(n626) );
  NAND2X0_HVT U174 ( .A1(n452), .A2(n403), .Y(n778) );
  MUX41X1_HVT U176 ( .A1(n397), .A3(n621), .A2(n549), .A4(n327), .S0(n489), 
        .S1(n435), .Y(n620) );
  NAND2X0_HVT U177 ( .A1(n392), .A2(n519), .Y(n619) );
  MUX41X1_HVT U182 ( .A1(n556), .A3(n523), .A2(n543), .A4(n563), .S0(n489), 
        .S1(n507), .Y(n614) );
  MUX41X1_HVT U189 ( .A1(n608), .A3(n327), .A2(n609), .A4(n560), .S0(n510), 
        .S1(n335), .Y(n607) );
  AO21X1_HVT U197 ( .A1(n494), .A2(n511), .A3(n570), .Y(n600) );
  MUX41X1_HVT U205 ( .A1(n411), .A3(n788), .A2(n566), .A4(n575), .S0(n506), 
        .S1(n536), .Y(n592) );
  NAND2X0_HVT U208 ( .A1(n527), .A2(n313), .Y(n681) );
  NAND2X0_HVT U215 ( .A1(n681), .A2(n412), .Y(n589) );
  NAND2X0_HVT U218 ( .A1(n314), .A2(n527), .Y(n643) );
  NAND2X0_HVT U220 ( .A1(n510), .A2(n590), .Y(n712) );
  INVX0_HVT U241 ( .A(n768), .Y(n582) );
  INVX0_HVT U242 ( .A(n751), .Y(n581) );
  INVX0_HVT U245 ( .A(n786), .Y(n579) );
  INVX0_HVT U256 ( .A(n643), .Y(n570) );
  INVX0_HVT U265 ( .A(n766), .Y(n563) );
  INVX0_HVT U268 ( .A(n770), .Y(n561) );
  INVX0_HVT U276 ( .A(n754), .Y(n556) );
  INVX0_HVT U278 ( .A(n760), .Y(n554) );
  INVX0_HVT U295 ( .A(n787), .Y(n546) );
  INVX0_HVT U302 ( .A(n588), .Y(n542) );
  INVX0_HVT U306 ( .A(n627), .Y(n541) );
  NBUFFX2_HVT U1 ( .A(in[3]), .Y(n515) );
  XNOR2X1_HVT U2 ( .A1(n473), .A2(n227), .Y(n497) );
  INVX0_HVT U3 ( .A(n764), .Y(n552) );
  OAI21X1_HVT U6 ( .A1(n530), .A2(n480), .A3(n551), .Y(n505) );
  INVX1_HVT U7 ( .A(n441), .Y(n457) );
  OA21X1_HVT U8 ( .A1(n496), .A2(n422), .A3(n762), .Y(n624) );
  XOR2X1_HVT U9 ( .A1(n408), .A2(n457), .Y(n766) );
  MUX21X1_HVT U10 ( .A1(n211), .A2(n518), .S0(n227), .Y(n717) );
  MUX21X1_HVT U11 ( .A1(n548), .A2(n493), .S0(n445), .Y(n663) );
  MUX21X1_HVT U12 ( .A1(n676), .A2(n677), .S0(n536), .Y(n675) );
  INVX1_HVT U13 ( .A(n441), .Y(n458) );
  INVX1_HVT U14 ( .A(n401), .Y(n445) );
  INVX0_HVT U16 ( .A(n529), .Y(n469) );
  INVX1_HVT U17 ( .A(n469), .Y(n451) );
  AND2X1_HVT U18 ( .A1(n388), .A2(n389), .Y(n5) );
  AND2X1_HVT U19 ( .A1(n378), .A2(n379), .Y(n23) );
  AND2X1_HVT U20 ( .A1(n114), .A2(n117), .Y(n28) );
  AND2X1_HVT U22 ( .A1(n217), .A2(n218), .Y(n47) );
  INVX1_HVT U23 ( .A(n517), .Y(n423) );
  INVX1_HVT U25 ( .A(n316), .Y(n402) );
  IBUFFX2_HVT U26 ( .A(n483), .Y(n753) );
  OR2X1_HVT U27 ( .A1(n316), .A2(n515), .Y(n313) );
  INVX1_HVT U28 ( .A(n515), .Y(n454) );
  INVX1_HVT U29 ( .A(n515), .Y(n406) );
  INVX1_HVT U30 ( .A(n385), .Y(n779) );
  MUX41X1_HVT U31 ( .A1(n574), .A3(n28), .A2(n398), .A4(n228), .S0(n421), .S1(
        n506), .Y(n647) );
  MUX41X1_HVT U32 ( .A1(n648), .A3(n647), .A2(n652), .A4(n651), .S0(n438), 
        .S1(n514), .Y(n646) );
  INVX1_HVT U34 ( .A(n755), .Y(n555) );
  NAND2X0_HVT U35 ( .A1(n409), .A2(n50), .Y(n114) );
  NAND2X0_HVT U36 ( .A1(n524), .A2(n216), .Y(n117) );
  INVX0_HVT U37 ( .A(n216), .Y(n50) );
  MUX41X1_HVT U38 ( .A1(n655), .A3(n657), .A2(n658), .A4(n659), .S0(n532), 
        .S1(n513), .Y(n654) );
  NAND2X0_HVT U39 ( .A1(n455), .A2(n517), .Y(n118) );
  MUX21X1_HVT U40 ( .A1(n361), .A2(n702), .S0(n497), .Y(n701) );
  INVX1_HVT U41 ( .A(n737), .Y(n574) );
  NBUFFX2_HVT U43 ( .A(n362), .Y(n489) );
  INVX1_HVT U44 ( .A(n525), .Y(n391) );
  NBUFFX2_HVT U45 ( .A(n565), .Y(n517) );
  INVX1_HVT U46 ( .A(n449), .Y(n334) );
  INVX1_HVT U47 ( .A(n296), .Y(n590) );
  NBUFFX2_HVT U48 ( .A(n532), .Y(n508) );
  INVX1_HVT U49 ( .A(n585), .Y(n571) );
  MUX21X1_HVT U50 ( .A1(n313), .A2(n474), .S0(n354), .Y(n405) );
  INVX1_HVT U52 ( .A(n259), .Y(n446) );
  INVX1_HVT U54 ( .A(n338), .Y(n759) );
  INVX1_HVT U55 ( .A(n477), .Y(n259) );
  INVX1_HVT U57 ( .A(n537), .Y(n534) );
  MUX21X1_HVT U60 ( .A1(n346), .A2(n577), .S0(n413), .Y(n784) );
  NBUFFX2_HVT U63 ( .A(n402), .Y(n397) );
  MUX21X1_HVT U64 ( .A1(n700), .A2(n701), .S0(n507), .Y(n698) );
  MUX21X1_HVT U65 ( .A1(n788), .A2(n345), .S0(n477), .Y(n683) );
  MUX21X1_HVT U67 ( .A1(n640), .A2(n310), .S0(n497), .Y(n639) );
  NBUFFX2_HVT U68 ( .A(n402), .Y(n519) );
  INVX1_HVT U69 ( .A(n341), .Y(n535) );
  NAND2X0_HVT U70 ( .A1(n338), .A2(n290), .Y(n293) );
  INVX1_HVT U71 ( .A(n387), .Y(n788) );
  MUX21X1_HVT U72 ( .A1(n568), .A2(n763), .S0(n451), .Y(n665) );
  AO21X1_HVT U75 ( .A1(n401), .A2(n522), .A3(n390), .Y(n676) );
  NBUFFX2_HVT U76 ( .A(n534), .Y(n362) );
  INVX0_HVT U78 ( .A(n362), .Y(n473) );
  INVX1_HVT U79 ( .A(n414), .Y(n347) );
  INVX1_HVT U80 ( .A(n445), .Y(n416) );
  NBUFFX2_HVT U81 ( .A(n529), .Y(n507) );
  INVX1_HVT U86 ( .A(n354), .Y(n414) );
  INVX1_HVT U87 ( .A(n414), .Y(n527) );
  INVX1_HVT U88 ( .A(n261), .Y(n450) );
  INVX1_HVT U89 ( .A(n451), .Y(n290) );
  INVX1_HVT U90 ( .A(n511), .Y(n422) );
  INVX0_HVT U91 ( .A(n341), .Y(n536) );
  INVX1_HVT U92 ( .A(n509), .Y(n438) );
  INVX1_HVT U93 ( .A(n765), .Y(n568) );
  INVX1_HVT U94 ( .A(n312), .Y(n360) );
  NBUFFX2_HVT U95 ( .A(n790), .Y(n329) );
  INVX1_HVT U97 ( .A(n790), .Y(n449) );
  INVX0_HVT U98 ( .A(n767), .Y(n540) );
  MUX21X1_HVT U99 ( .A1(n314), .A2(n562), .S0(n289), .Y(n726) );
  INVX0_HVT U100 ( .A(n772), .Y(n539) );
  MUX41X1_HVT U102 ( .A1(n745), .A3(n751), .A2(n605), .A4(n758), .S0(n504), 
        .S1(n451), .Y(n604) );
  INVX0_HVT U104 ( .A(n580), .Y(n456) );
  INVX1_HVT U106 ( .A(n119), .Y(n424) );
  MUX41X1_HVT U107 ( .A1(n783), .A3(n546), .A2(n490), .A4(n482), .S0(n447), 
        .S1(n451), .Y(n616) );
  INVX1_HVT U108 ( .A(n313), .Y(n481) );
  MUX21X1_HVT U109 ( .A1(n456), .A2(n523), .S0(n458), .Y(n783) );
  INVX0_HVT U111 ( .A(n776), .Y(n545) );
  INVX0_HVT U112 ( .A(n528), .Y(n525) );
  INVX0_HVT U113 ( .A(n528), .Y(n227) );
  INVX1_HVT U114 ( .A(n477), .Y(n335) );
  INVX0_HVT U116 ( .A(n528), .Y(n413) );
  INVX0_HVT U117 ( .A(n227), .Y(n241) );
  MUX41X1_HVT U118 ( .A1(n716), .A3(n718), .A2(n719), .A4(n723), .S0(n508), 
        .S1(n513), .Y(n715) );
  INVX0_HVT U119 ( .A(n454), .Y(n119) );
  INVX0_HVT U120 ( .A(n454), .Y(n455) );
  INVX0_HVT U121 ( .A(n515), .Y(n580) );
  MUX21X1_HVT U122 ( .A1(n774), .A2(n553), .S0(n435), .Y(n662) );
  INVX0_HVT U124 ( .A(in[1]), .Y(n528) );
  MUX41X1_HVT U125 ( .A1(n482), .A3(n540), .A2(n679), .A4(n762), .S0(n488), 
        .S1(n335), .Y(n678) );
  MUX21X2_HVT U126 ( .A1(n226), .A2(n484), .S0(n457), .Y(n483) );
  INVX1_HVT U127 ( .A(n330), .Y(n210) );
  INVX1_HVT U128 ( .A(n210), .Y(n211) );
  INVX1_HVT U129 ( .A(n284), .Y(n728) );
  AO21X1_HVT U130 ( .A1(n512), .A2(n699), .A3(n570), .Y(n700) );
  INVX1_HVT U132 ( .A(n565), .Y(n316) );
  NAND2X0_HVT U133 ( .A1(n644), .A2(n381), .Y(n212) );
  NAND2X0_HVT U134 ( .A1(n645), .A2(n507), .Y(n213) );
  NAND2X0_HVT U137 ( .A1(n212), .A2(n213), .Y(n642) );
  NAND2X0_HVT U138 ( .A1(n520), .A2(n216), .Y(n217) );
  NAND2X0_HVT U139 ( .A1(n211), .A2(n403), .Y(n218) );
  INVX0_HVT U143 ( .A(n525), .Y(n216) );
  MUX21X1_HVT U144 ( .A1(n314), .A2(n47), .S0(n473), .Y(n645) );
  INVX1_HVT U145 ( .A(n530), .Y(n529) );
  INVX0_HVT U146 ( .A(in[2]), .Y(n530) );
  INVX0_HVT U147 ( .A(n459), .Y(n777) );
  MUX21X1_HVT U148 ( .A1(n763), .A2(n589), .S0(n511), .Y(n584) );
  INVX1_HVT U149 ( .A(n514), .Y(n324) );
  NAND2X0_HVT U150 ( .A1(n357), .A2(n358), .Y(n219) );
  MUX41X1_HVT U151 ( .A1(n594), .A3(n595), .A2(n592), .A4(n593), .S0(n509), 
        .S1(n324), .Y(n591) );
  INVX0_HVT U152 ( .A(n789), .Y(n224) );
  INVX1_HVT U155 ( .A(n224), .Y(n226) );
  INVX0_HVT U156 ( .A(n762), .Y(n575) );
  INVX1_HVT U157 ( .A(n470), .Y(n321) );
  INVX0_HVT U160 ( .A(n345), .Y(n757) );
  INVX0_HVT U161 ( .A(n385), .Y(n482) );
  MUX21X2_HVT U163 ( .A1(n412), .A2(n405), .S0(n473), .Y(n660) );
  INVX0_HVT U164 ( .A(n578), .Y(n228) );
  INVX1_HVT U169 ( .A(n720), .Y(n578) );
  NAND2X0_HVT U170 ( .A1(n347), .A2(n415), .Y(n720) );
  MUX21X1_HVT U171 ( .A1(n481), .A2(n275), .S0(n458), .Y(n697) );
  INVX1_HVT U172 ( .A(n439), .Y(n390) );
  NAND2X0_HVT U173 ( .A1(n460), .A2(n229), .Y(n231) );
  NAND2X0_HVT U175 ( .A1(n410), .A2(n501), .Y(n232) );
  NAND2X0_HVT U178 ( .A1(n231), .A2(n232), .Y(n499) );
  INVX0_HVT U179 ( .A(n501), .Y(n229) );
  INVX0_HVT U180 ( .A(n361), .Y(n460) );
  XNOR2X1_HVT U181 ( .A1(n392), .A2(n529), .Y(n501) );
  MUX41X1_HVT U183 ( .A1(n687), .A3(n685), .A2(n692), .A4(n688), .S0(n438), 
        .S1(n514), .Y(n684) );
  INVX1_HVT U184 ( .A(n330), .Y(n439) );
  INVX1_HVT U185 ( .A(n440), .Y(n441) );
  INVX1_HVT U186 ( .A(in[4]), .Y(n565) );
  INVX1_HVT U187 ( .A(n368), .Y(n403) );
  NBUFFX2_HVT U188 ( .A(n313), .Y(n523) );
  NAND2X0_HVT U190 ( .A1(n490), .A2(n511), .Y(n236) );
  NAND2X0_HVT U191 ( .A1(n775), .A2(n470), .Y(n238) );
  NAND2X0_HVT U192 ( .A1(n236), .A2(n238), .Y(n597) );
  MUX21X1_HVT U193 ( .A1(n226), .A2(n275), .S0(n227), .Y(n752) );
  MUX41X1_HVT U194 ( .A1(n495), .A3(n574), .A2(n776), .A4(n403), .S0(n381), 
        .S1(n488), .Y(n695) );
  INVX0_HVT U195 ( .A(n360), .Y(n361) );
  INVX0_HVT U196 ( .A(n460), .Y(n310) );
  OR2X1_HVT U198 ( .A1(n474), .A2(n261), .Y(n758) );
  MUX41X1_HVT U199 ( .A1(n703), .A3(n696), .A2(n698), .A4(n695), .S0(n324), 
        .S1(n289), .Y(n694) );
  MUX21X1_HVT U200 ( .A1(n484), .A2(n500), .S0(n450), .Y(n772) );
  MUX41X1_HVT U201 ( .A1(n772), .A3(n550), .A2(n781), .A4(n738), .S0(n470), 
        .S1(n508), .Y(n736) );
  INVX0_HVT U202 ( .A(n528), .Y(n526) );
  MUX41X1_HVT U203 ( .A1(n491), .A3(n707), .A2(n494), .A4(n571), .S0(n447), 
        .S1(n290), .Y(n706) );
  INVX1_HVT U204 ( .A(n531), .Y(n289) );
  MUX21X1_HVT U206 ( .A1(n516), .A2(n449), .S0(n457), .Y(n633) );
  MUX41X1_HVT U207 ( .A1(n633), .A3(n493), .A2(n632), .A4(n569), .S0(n446), 
        .S1(n447), .Y(n631) );
  INVX0_HVT U209 ( .A(n783), .Y(n562) );
  INVX1_HVT U210 ( .A(n784), .Y(n547) );
  INVX1_HVT U211 ( .A(n341), .Y(n485) );
  INVX0_HVT U212 ( .A(n789), .Y(n311) );
  NBUFFX2_HVT U213 ( .A(n532), .Y(n509) );
  XNOR2X2_HVT U214 ( .A1(n346), .A2(n261), .Y(n398) );
  INVX1_HVT U216 ( .A(n391), .Y(n392) );
  INVX1_HVT U217 ( .A(n440), .Y(n354) );
  INVX1_HVT U219 ( .A(n587), .Y(n550) );
  NAND2X0_HVT U221 ( .A1(n241), .A2(n211), .Y(n252) );
  NAND2X0_HVT U222 ( .A1(n360), .A2(n526), .Y(n253) );
  NAND2X0_HVT U223 ( .A1(n253), .A2(n252), .Y(n767) );
  MUX41X1_HVT U224 ( .A1(n765), .A3(n566), .A2(n296), .A4(n434), .S0(n259), 
        .S1(n485), .Y(n617) );
  NBUFFX2_HVT U225 ( .A(n441), .Y(n261) );
  NAND2X0_HVT U226 ( .A1(n724), .A2(n264), .Y(n267) );
  NAND2X0_HVT U227 ( .A1(n749), .A2(n446), .Y(n274) );
  NAND2X0_HVT U228 ( .A1(n267), .A2(n274), .Y(n723) );
  INVX0_HVT U229 ( .A(n477), .Y(n264) );
  XNOR2X1_HVT U230 ( .A1(n448), .A2(n321), .Y(n749) );
  MUX41X1_HVT U231 ( .A1(n725), .A3(n733), .A2(n729), .A4(n739), .S0(in[6]), 
        .S1(n513), .Y(out[0]) );
  NAND2X0_HVT U232 ( .A1(n118), .A2(n426), .Y(n275) );
  MUX41X1_HVT U233 ( .A1(n571), .A3(n574), .A2(n540), .A4(n460), .S0(n445), 
        .S1(n321), .Y(n718) );
  MUX21X1_HVT U234 ( .A1(n572), .A2(n481), .S0(n526), .Y(n773) );
  NAND2X0_HVT U235 ( .A1(n449), .A2(n422), .Y(n276) );
  NAND2X0_HVT U236 ( .A1(n573), .A2(n512), .Y(n278) );
  NAND2X0_HVT U237 ( .A1(n276), .A2(n278), .Y(n724) );
  NAND2X0_HVT U238 ( .A1(n625), .A2(n290), .Y(n279) );
  NAND2X0_HVT U239 ( .A1(n624), .A2(n506), .Y(n280) );
  NAND2X0_HVT U240 ( .A1(n279), .A2(n280), .Y(n623) );
  MUX21X1_HVT U243 ( .A1(n359), .A2(n573), .S0(n512), .Y(n625) );
  INVX1_HVT U244 ( .A(n297), .Y(n314) );
  XOR2X2_HVT U246 ( .A1(n403), .A2(n453), .Y(n748) );
  MUX41X1_HVT U247 ( .A1(n626), .A3(n623), .A2(n631), .A4(n629), .S0(n438), 
        .S1(n514), .Y(n622) );
  INVX0_HVT U248 ( .A(in[1]), .Y(n440) );
  NAND2X0_HVT U249 ( .A1(n434), .A2(n512), .Y(n282) );
  NAND2X0_HVT U250 ( .A1(n581), .A2(n470), .Y(n283) );
  NAND2X0_HVT U251 ( .A1(n282), .A2(n283), .Y(n601) );
  MUX41X1_HVT U252 ( .A1(n710), .A3(n706), .A2(n711), .A4(n708), .S0(n324), 
        .S1(n509), .Y(n705) );
  INVX1_HVT U253 ( .A(n397), .Y(n411) );
  AND3X1_HVT U254 ( .A1(n310), .A2(n737), .A3(n712), .Y(n713) );
  MUX21X1_HVT U255 ( .A1(n306), .A2(n780), .S0(n289), .Y(n284) );
  MUX41X1_HVT U257 ( .A1(n728), .A3(n726), .A2(n727), .A4(n547), .S0(n381), 
        .S1(n341), .Y(n725) );
  MUX41X1_HVT U258 ( .A1(n573), .A3(n390), .A2(n756), .A4(n415), .S0(n381), 
        .S1(n535), .Y(n602) );
  NAND2X0_HVT U259 ( .A1(n769), .A2(n451), .Y(n295) );
  NAND2X0_HVT U260 ( .A1(n293), .A2(n295), .Y(n463) );
  AND2X1_HVT U261 ( .A1(n785), .A2(n457), .Y(n296) );
  MUX21X1_HVT U262 ( .A1(n415), .A2(n782), .S0(n525), .Y(n762) );
  NAND2X0_HVT U263 ( .A1(n684), .A2(n464), .Y(n395) );
  MUX41X1_HVT U264 ( .A1(n610), .A3(n614), .A2(n607), .A4(n611), .S0(n513), 
        .S1(n438), .Y(n606) );
  INVX0_HVT U266 ( .A(n313), .Y(n557) );
  INVX1_HVT U267 ( .A(n572), .Y(n297) );
  MUX21X2_HVT U269 ( .A1(n650), .A2(n649), .S0(n506), .Y(n648) );
  NAND2X0_HVT U270 ( .A1(n740), .A2(n446), .Y(n299) );
  NAND2X0_HVT U271 ( .A1(n744), .A2(n363), .Y(n303) );
  NAND2X0_HVT U272 ( .A1(n303), .A2(n299), .Y(n739) );
  INVX1_HVT U273 ( .A(n381), .Y(n363) );
  INVX0_HVT U274 ( .A(n480), .Y(n756) );
  MUX21X1_HVT U275 ( .A1(n481), .A2(n516), .S0(n347), .Y(n480) );
  OA21X1_HVT U277 ( .A1(n784), .A2(n447), .A3(n555), .Y(n596) );
  NAND2X0_HVT U279 ( .A1(n787), .A2(n259), .Y(n304) );
  NAND2X0_HVT U280 ( .A1(n656), .A2(n446), .Y(n305) );
  NAND2X0_HVT U281 ( .A1(n304), .A2(n305), .Y(n655) );
  MUX21X1_HVT U282 ( .A1(n769), .A2(n556), .S0(n511), .Y(n656) );
  MUX41X1_HVT U283 ( .A1(n618), .A3(n620), .A2(n616), .A4(n617), .S0(n509), 
        .S1(n324), .Y(n615) );
  NAND2X0_HVT U284 ( .A1(n518), .A2(n306), .Y(n307) );
  NAND2X0_HVT U285 ( .A1(n216), .A2(n275), .Y(n308) );
  NAND2X0_HVT U286 ( .A1(n307), .A2(n308), .Y(n689) );
  INVX0_HVT U287 ( .A(n216), .Y(n306) );
  NAND2X0_HVT U288 ( .A1(n407), .A2(n518), .Y(n309) );
  INVX0_HVT U289 ( .A(n401), .Y(n477) );
  INVX0_HVT U290 ( .A(n435), .Y(n381) );
  INVX1_HVT U291 ( .A(n311), .Y(n312) );
  INVX0_HVT U292 ( .A(n380), .Y(n315) );
  INVX0_HVT U293 ( .A(n752), .Y(n543) );
  NBUFFX2_HVT U294 ( .A(n565), .Y(n518) );
  INVX0_HVT U296 ( .A(in[5]), .Y(n533) );
  NAND2X0_HVT U297 ( .A1(n518), .A2(n241), .Y(n317) );
  NAND2X0_HVT U298 ( .A1(n315), .A2(n50), .Y(n318) );
  NAND2X0_HVT U299 ( .A1(n317), .A2(n318), .Y(n434) );
  MUX21X1_HVT U300 ( .A1(n329), .A2(n411), .S0(n450), .Y(n583) );
  MUX21X2_HVT U301 ( .A1(n564), .A2(n338), .S0(n435), .Y(n677) );
  MUX21X1_HVT U303 ( .A1(n500), .A2(n481), .S0(n458), .Y(n621) );
  MUX21X1_HVT U304 ( .A1(n397), .A2(n406), .S0(n469), .Y(n410) );
  INVX1_HVT U305 ( .A(n583), .Y(n566) );
  NAND2X0_HVT U307 ( .A1(n423), .A2(n424), .Y(n319) );
  NAND2X0_HVT U308 ( .A1(n423), .A2(n424), .Y(n320) );
  MUX21X1_HVT U309 ( .A1(n336), .A2(n521), .S0(n241), .Y(n608) );
  NAND2X0_HVT U310 ( .A1(n713), .A2(n451), .Y(n322) );
  NAND2X0_HVT U311 ( .A1(n714), .A2(n290), .Y(n323) );
  NAND2X0_HVT U312 ( .A1(n322), .A2(n323), .Y(n711) );
  MUX21X1_HVT U313 ( .A1(n386), .A2(n771), .S0(n422), .Y(n714) );
  INVX0_HVT U314 ( .A(n689), .Y(n549) );
  XNOR2X2_HVT U315 ( .A1(n334), .A2(n413), .Y(n494) );
  NAND2X0_HVT U316 ( .A1(n743), .A2(n489), .Y(n325) );
  NAND2X0_HVT U317 ( .A1(n742), .A2(n422), .Y(n326) );
  NAND2X0_HVT U318 ( .A1(n325), .A2(n326), .Y(n740) );
  INVX0_HVT U319 ( .A(n380), .Y(n572) );
  INVX0_HVT U320 ( .A(n461), .Y(n412) );
  NAND2X0_HVT U321 ( .A1(n403), .A2(n452), .Y(n327) );
  NBUFFX2_HVT U322 ( .A(n580), .Y(n521) );
  INVX0_HVT U323 ( .A(n761), .Y(n553) );
  INVX0_HVT U324 ( .A(n413), .Y(n328) );
  INVX0_HVT U325 ( .A(n510), .Y(n470) );
  AND2X1_HVT U326 ( .A1(n118), .A2(n320), .Y(n330) );
  NAND2X0_HVT U327 ( .A1(n523), .A2(n413), .Y(n332) );
  NAND2X0_HVT U328 ( .A1(n331), .A2(n328), .Y(n333) );
  NAND2X0_HVT U329 ( .A1(n332), .A2(n333), .Y(n493) );
  INVX0_HVT U330 ( .A(n523), .Y(n331) );
  INVX0_HVT U331 ( .A(n309), .Y(n500) );
  INVX1_HVT U332 ( .A(n502), .Y(n680) );
  MUX21X1_HVT U333 ( .A1(n474), .A2(n557), .S0(n414), .Y(n761) );
  INVX1_HVT U334 ( .A(n775), .Y(n548) );
  INVX0_HVT U335 ( .A(n758), .Y(n564) );
  NBUFFX2_HVT U336 ( .A(n401), .Y(n435) );
  OR2X1_HVT U337 ( .A1(n406), .A2(n402), .Y(n336) );
  INVX1_HVT U338 ( .A(n336), .Y(n577) );
  AND2X1_HVT U339 ( .A1(n241), .A2(n411), .Y(n337) );
  AND2X1_HVT U340 ( .A1(n337), .A2(n506), .Y(n664) );
  NBUFFX2_HVT U341 ( .A(n529), .Y(n506) );
  AND2X1_HVT U342 ( .A1(n369), .A2(n370), .Y(n338) );
  OA21X1_HVT U343 ( .A1(n759), .A2(n447), .A3(n5), .Y(n612) );
  NAND2X0_HVT U344 ( .A1(n520), .A2(n391), .Y(n339) );
  NAND2X0_HVT U345 ( .A1(n474), .A2(n527), .Y(n340) );
  NAND2X0_HVT U346 ( .A1(n339), .A2(n340), .Y(n763) );
  INVX1_HVT U347 ( .A(n517), .Y(n474) );
  INVX0_HVT U348 ( .A(n763), .Y(n567) );
  MUX21X1_HVT U349 ( .A1(n314), .A2(n311), .S0(n391), .Y(n459) );
  INVX1_HVT U350 ( .A(n534), .Y(n341) );
  NBUFFX2_HVT U351 ( .A(n534), .Y(n510) );
  INVX0_HVT U352 ( .A(n682), .Y(n351) );
  INVX0_HVT U353 ( .A(n681), .Y(n559) );
  INVX1_HVT U354 ( .A(in[7]), .Y(n537) );
  INVX1_HVT U355 ( .A(n683), .Y(n503) );
  NAND2X0_HVT U356 ( .A1(n478), .A2(n479), .Y(out[4]) );
  NAND2X0_HVT U357 ( .A1(n538), .A2(n381), .Y(n342) );
  NAND2X0_HVT U358 ( .A1(n660), .A2(n335), .Y(n343) );
  NAND2X0_HVT U359 ( .A1(n343), .A2(n342), .Y(n659) );
  INVX0_HVT U360 ( .A(n519), .Y(n408) );
  INVX1_HVT U361 ( .A(n464), .Y(n344) );
  INVX0_HVT U362 ( .A(in[6]), .Y(n464) );
  MUX41X1_HVT U363 ( .A1(n604), .A3(n602), .A2(n603), .A4(n599), .S0(n324), 
        .S1(n438), .Y(n598) );
  MUX21X1_HVT U364 ( .A1(n790), .A2(n397), .S0(n368), .Y(n345) );
  NAND2X0_HVT U365 ( .A1(n118), .A2(n426), .Y(n346) );
  INVX0_HVT U366 ( .A(n785), .Y(n382) );
  MUX41X1_HVT U367 ( .A1(n757), .A3(n219), .A2(n483), .A4(n761), .S0(n485), 
        .S1(n507), .Y(n594) );
  NBUFFX2_HVT U368 ( .A(in[2]), .Y(n401) );
  NAND2X0_HVT U369 ( .A1(n360), .A2(n392), .Y(n348) );
  NAND2X0_HVT U370 ( .A1(n314), .A2(n414), .Y(n349) );
  NAND2X0_HVT U371 ( .A1(n348), .A2(n349), .Y(n630) );
  MUX21X1_HVT U372 ( .A1(n575), .A2(n351), .S0(n506), .Y(n350) );
  NAND2X0_HVT U373 ( .A1(n764), .A2(n470), .Y(n352) );
  NAND2X0_HVT U374 ( .A1(n387), .A2(n512), .Y(n353) );
  NAND2X0_HVT U375 ( .A1(n352), .A2(n353), .Y(n650) );
  MUX21X1_HVT U376 ( .A1(n557), .A2(n518), .S0(n458), .Y(n764) );
  MUX21X1_HVT U377 ( .A1(n575), .A2(n777), .S0(n507), .Y(n693) );
  MUX41X1_HVT U378 ( .A1(n637), .A3(n635), .A2(n642), .A4(n641), .S0(n438), 
        .S1(n513), .Y(n634) );
  INVX0_HVT U379 ( .A(n589), .Y(n560) );
  NAND2X0_HVT U380 ( .A1(n672), .A2(n447), .Y(n355) );
  NAND2X0_HVT U381 ( .A1(n671), .A2(n512), .Y(n356) );
  NAND2X0_HVT U382 ( .A1(n355), .A2(n356), .Y(n668) );
  NAND2X0_HVT U383 ( .A1(n409), .A2(n241), .Y(n357) );
  NAND2X0_HVT U384 ( .A1(n521), .A2(n306), .Y(n358) );
  NAND2X0_HVT U385 ( .A1(n358), .A2(n357), .Y(n780) );
  INVX1_HVT U386 ( .A(n481), .Y(n409) );
  NBUFFX2_HVT U387 ( .A(n532), .Y(n531) );
  INVX0_HVT U388 ( .A(n461), .Y(n359) );
  MUX41X1_HVT U389 ( .A1(n545), .A3(n731), .A2(n459), .A4(n385), .S0(n422), 
        .S1(n508), .Y(n730) );
  INVX0_HVT U390 ( .A(n781), .Y(n576) );
  INVX1_HVT U391 ( .A(n390), .Y(n373) );
  NBUFFX2_HVT U392 ( .A(n362), .Y(n512) );
  NAND2X0_HVT U393 ( .A1(n600), .A2(n363), .Y(n364) );
  NAND2X0_HVT U394 ( .A1(n601), .A2(n381), .Y(n365) );
  NAND2X0_HVT U395 ( .A1(n364), .A2(n365), .Y(n599) );
  NAND2X0_HVT U396 ( .A1(n462), .A2(n422), .Y(n366) );
  NAND2X0_HVT U397 ( .A1(n463), .A2(n536), .Y(n367) );
  NAND2X0_HVT U398 ( .A1(n366), .A2(n367), .Y(n593) );
  NAND2X0_HVT U399 ( .A1(n577), .A2(n368), .Y(n369) );
  NAND2X0_HVT U400 ( .A1(n520), .A2(n527), .Y(n370) );
  INVX0_HVT U401 ( .A(n354), .Y(n368) );
  INVX1_HVT U402 ( .A(n404), .Y(n702) );
  INVX1_HVT U403 ( .A(n485), .Y(n447) );
  MUX21X1_HVT U404 ( .A1(n577), .A2(n557), .S0(n413), .Y(n755) );
  NAND2X0_HVT U405 ( .A1(n606), .A2(n464), .Y(n371) );
  NAND2X0_HVT U406 ( .A1(n615), .A2(n344), .Y(n372) );
  NAND2X0_HVT U407 ( .A1(n372), .A2(n371), .Y(out[6]) );
  NAND2X0_HVT U408 ( .A1(n639), .A2(n264), .Y(n374) );
  NAND2X0_HVT U409 ( .A1(n638), .A2(n446), .Y(n375) );
  NAND2X0_HVT U410 ( .A1(n374), .A2(n375), .Y(n637) );
  MUX21X1_HVT U411 ( .A1(n558), .A2(n755), .S0(n422), .Y(n638) );
  NAND2X0_HVT U412 ( .A1(n678), .A2(n531), .Y(n376) );
  NAND2X0_HVT U413 ( .A1(n675), .A2(n438), .Y(n377) );
  NAND2X0_HVT U414 ( .A1(n376), .A2(n377), .Y(n674) );
  MUX41X1_HVT U415 ( .A1(n666), .A3(n661), .A2(n680), .A4(n674), .S0(n324), 
        .S1(in[6]), .Y(out[3]) );
  OR2X1_HVT U416 ( .A1(n406), .A2(n402), .Y(n790) );
  INVX1_HVT U417 ( .A(n406), .Y(n407) );
  NAND2X0_HVT U418 ( .A1(n452), .A2(n328), .Y(n378) );
  NAND2X0_HVT U419 ( .A1(n315), .A2(n403), .Y(n379) );
  NAND2X0_HVT U420 ( .A1(n423), .A2(n580), .Y(n380) );
  INVX1_HVT U421 ( .A(n439), .Y(n785) );
  MUX21X1_HVT U422 ( .A1(n520), .A2(n486), .S0(n457), .Y(n775) );
  XOR2X1_HVT U423 ( .A1(n261), .A2(n456), .Y(n746) );
  NAND2X0_HVT U424 ( .A1(n734), .A2(n530), .Y(n383) );
  NAND2X0_HVT U425 ( .A1(n736), .A2(n401), .Y(n384) );
  NAND2X0_HVT U426 ( .A1(n384), .A2(n383), .Y(n733) );
  AND2X1_HVT U427 ( .A1(n778), .A2(n336), .Y(n385) );
  XOR2X2_HVT U428 ( .A1(n312), .A2(n526), .Y(n745) );
  NAND2X0_HVT U429 ( .A1(n715), .A2(n344), .Y(n436) );
  INVX0_HVT U430 ( .A(n535), .Y(n421) );
  INVX0_HVT U431 ( .A(n315), .Y(n386) );
  AND2X1_HVT U432 ( .A1(n526), .A2(n309), .Y(n387) );
  NAND2X0_HVT U433 ( .A1(n275), .A2(n216), .Y(n388) );
  NAND2X0_HVT U434 ( .A1(n456), .A2(n403), .Y(n389) );
  NAND2X0_HVT U435 ( .A1(n388), .A2(n389), .Y(n769) );
  NAND2X0_HVT U436 ( .A1(n622), .A2(n464), .Y(n393) );
  NAND2X0_HVT U437 ( .A1(n634), .A2(n344), .Y(n394) );
  NAND2X0_HVT U438 ( .A1(n393), .A2(n394), .Y(out[5]) );
  INVX0_HVT U439 ( .A(n521), .Y(n484) );
  NAND2X0_HVT U440 ( .A1(n694), .A2(n344), .Y(n396) );
  NAND2X0_HVT U441 ( .A1(n396), .A2(n395), .Y(out[2]) );
  MUX21X1_HVT U442 ( .A1(n474), .A2(n226), .S0(n347), .Y(n771) );
  NAND2X0_HVT U443 ( .A1(n779), .A2(n416), .Y(n399) );
  NAND2X0_HVT U444 ( .A1(n738), .A2(n469), .Y(n400) );
  NAND2X0_HVT U445 ( .A1(n399), .A2(n400), .Y(n462) );
  MUX21X1_HVT U446 ( .A1(n408), .A2(n520), .S0(n473), .Y(n404) );
  INVX1_HVT U447 ( .A(n586), .Y(n573) );
  INVX0_HVT U448 ( .A(n782), .Y(n461) );
  NAND2X0_HVT U449 ( .A1(n455), .A2(n316), .Y(n415) );
  NAND2X0_HVT U450 ( .A1(n613), .A2(n416), .Y(n417) );
  NAND2X0_HVT U451 ( .A1(n612), .A2(n445), .Y(n418) );
  NAND2X0_HVT U452 ( .A1(n417), .A2(n418), .Y(n611) );
  NAND2X0_HVT U453 ( .A1(n691), .A2(n446), .Y(n419) );
  NAND2X0_HVT U454 ( .A1(n264), .A2(n538), .Y(n420) );
  NAND2X0_HVT U455 ( .A1(n419), .A2(n420), .Y(n688) );
  INVX1_HVT U456 ( .A(n584), .Y(n538) );
  MUX41X1_HVT U457 ( .A1(n398), .A3(n228), .A2(n754), .A4(n495), .S0(n446), 
        .S1(n421), .Y(n610) );
  INVX1_HVT U458 ( .A(n522), .Y(n453) );
  NAND2X0_HVT U459 ( .A1(n455), .A2(n517), .Y(n425) );
  NAND2X0_HVT U460 ( .A1(n423), .A2(n424), .Y(n426) );
  NAND2X0_HVT U461 ( .A1(n425), .A2(n319), .Y(n486) );
  NBUFFX2_HVT U462 ( .A(n486), .Y(n516) );
  NAND2X0_HVT U463 ( .A1(n430), .A2(n431), .Y(n427) );
  MUX41X1_HVT U464 ( .A1(n619), .A3(n755), .A2(n774), .A4(n434), .S0(n536), 
        .S1(n445), .Y(n618) );
  NAND2X0_HVT U465 ( .A1(n474), .A2(n241), .Y(n428) );
  NAND2X0_HVT U466 ( .A1(n461), .A2(n347), .Y(n429) );
  NAND2X0_HVT U467 ( .A1(n428), .A2(n429), .Y(n774) );
  INVX0_HVT U468 ( .A(n699), .Y(n558) );
  INVX0_HVT U469 ( .A(n774), .Y(n569) );
  MUX41X1_HVT U470 ( .A1(n704), .A3(n542), .A2(n751), .A4(n398), .S0(n290), 
        .S1(n421), .Y(n703) );
  MUX41X1_HVT U471 ( .A1(n752), .A3(n23), .A2(n427), .A4(n386), .S0(n416), 
        .S1(n510), .Y(n603) );
  NAND2X0_HVT U472 ( .A1(n577), .A2(n227), .Y(n430) );
  NAND2X0_HVT U473 ( .A1(n500), .A2(n450), .Y(n431) );
  NAND2X0_HVT U474 ( .A1(n431), .A2(n430), .Y(n448) );
  MUX41X1_HVT U475 ( .A1(n505), .A3(n350), .A2(n503), .A4(n499), .S0(n289), 
        .S1(n504), .Y(n502) );
  NAND2X0_HVT U476 ( .A1(n596), .A2(n290), .Y(n432) );
  NAND2X0_HVT U477 ( .A1(n597), .A2(n401), .Y(n433) );
  NAND2X0_HVT U478 ( .A1(n432), .A2(n433), .Y(n595) );
  OR2X1_HVT U479 ( .A1(n457), .A2(n572), .Y(n737) );
  NAND2X0_HVT U480 ( .A1(n705), .A2(n464), .Y(n437) );
  NAND2X0_HVT U481 ( .A1(n437), .A2(n436), .Y(out[1]) );
  MUX21X2_HVT U482 ( .A1(n412), .A2(n409), .S0(n450), .Y(n704) );
  MUX21X1_HVT U483 ( .A1(n407), .A2(n557), .S0(n347), .Y(n754) );
  NAND2X0_HVT U484 ( .A1(n492), .A2(n442), .Y(n443) );
  NAND2X0_HVT U485 ( .A1(n693), .A2(n747), .Y(n444) );
  NAND2X0_HVT U486 ( .A1(n443), .A2(n444), .Y(n692) );
  INVX0_HVT U487 ( .A(n747), .Y(n442) );
  OA21X1_HVT U488 ( .A1(n541), .A2(n422), .A3(n762), .Y(n649) );
  MUX21X1_HVT U489 ( .A1(n554), .A2(n673), .S0(n335), .Y(n672) );
  MUX21X1_HVT U490 ( .A1(n415), .A2(n313), .S0(n458), .Y(n699) );
  INVX0_HVT U491 ( .A(n771), .Y(n544) );
  INVX1_HVT U492 ( .A(n516), .Y(n452) );
  INVX1_HVT U493 ( .A(n773), .Y(n551) );
  AO21X1_HVT U494 ( .A1(n241), .A2(n453), .A3(n421), .Y(n690) );
  NBUFFX2_HVT U495 ( .A(n782), .Y(n522) );
  OA21X1_HVT U496 ( .A1(n753), .A2(n422), .A3(n643), .Y(n644) );
  NAND2X0_HVT U497 ( .A1(n591), .A2(n464), .Y(n465) );
  NAND2X0_HVT U498 ( .A1(n598), .A2(n344), .Y(n466) );
  NAND2X0_HVT U499 ( .A1(n466), .A2(n465), .Y(out[7]) );
  NAND2X0_HVT U500 ( .A1(n484), .A2(n289), .Y(n467) );
  NAND2X0_HVT U501 ( .A1(n758), .A2(in[5]), .Y(n468) );
  NAND2X0_HVT U502 ( .A1(n467), .A2(n468), .Y(n743) );
  MUX21X1_HVT U503 ( .A1(n707), .A2(n407), .S0(n510), .Y(n613) );
  MUX21X1_HVT U504 ( .A1(n519), .A2(n521), .S0(n458), .Y(n605) );
  NAND2X0_HVT U505 ( .A1(n667), .A2(n438), .Y(n471) );
  NAND2X0_HVT U506 ( .A1(n668), .A2(n532), .Y(n472) );
  NAND2X0_HVT U507 ( .A1(n471), .A2(n472), .Y(n666) );
  MUX41X1_HVT U508 ( .A1(n770), .A3(n498), .A2(n547), .A4(n405), .S0(n416), 
        .S1(n489), .Y(n667) );
  NAND2X0_HVT U509 ( .A1(n732), .A2(n264), .Y(n475) );
  NAND2X0_HVT U510 ( .A1(n730), .A2(n477), .Y(n476) );
  NAND2X0_HVT U511 ( .A1(n475), .A2(n476), .Y(n729) );
  NAND2X0_HVT U512 ( .A1(n646), .A2(n464), .Y(n478) );
  NAND2X0_HVT U513 ( .A1(n654), .A2(in[6]), .Y(n479) );
  INVX1_HVT U514 ( .A(n533), .Y(n532) );
  INVX0_HVT U515 ( .A(n536), .Y(n504) );
  NBUFFX2_HVT U516 ( .A(n510), .Y(n487) );
  NBUFFX2_HVT U517 ( .A(n362), .Y(n488) );
  AND2X1_HVT U518 ( .A1(n382), .A2(n737), .Y(n490) );
  MUX21X1_HVT U519 ( .A1(n331), .A2(n577), .S0(n531), .Y(n741) );
  AND2X1_HVT U520 ( .A1(n361), .A2(n720), .Y(n491) );
  MUX21X1_HVT U521 ( .A1(n329), .A2(n524), .S0(n526), .Y(n609) );
  MUX21X1_HVT U522 ( .A1(n521), .A2(n449), .S0(n527), .Y(n781) );
  MUX21X1_HVT U523 ( .A1(n397), .A2(n521), .S0(n392), .Y(n673) );
  NBUFFX2_HVT U524 ( .A(n309), .Y(n524) );
  MUX21X1_HVT U525 ( .A1(n226), .A2(n519), .S0(n392), .Y(n588) );
  AND2X1_HVT U526 ( .A1(n329), .A2(n681), .Y(n492) );
  AND2X1_HVT U527 ( .A1(n403), .A2(n360), .Y(n495) );
  MUX21X1_HVT U528 ( .A1(n297), .A2(n520), .S0(n261), .Y(n586) );
  MUX21X1_HVT U529 ( .A1(n412), .A2(n518), .S0(n527), .Y(n722) );
  MUX21X1_HVT U530 ( .A1(n386), .A2(n329), .S0(n506), .Y(n670) );
  NBUFFX2_HVT U531 ( .A(n580), .Y(n520) );
  NBUFFX2_HVT U532 ( .A(n534), .Y(n511) );
  MUX21X1_HVT U533 ( .A1(n359), .A2(n439), .S0(n526), .Y(n686) );
  AND2X1_HVT U534 ( .A1(n373), .A2(n391), .Y(n496) );
  NAND2X0_HVT U535 ( .A1(n407), .A2(n518), .Y(n789) );
  XOR2X1_HVT U536 ( .A1(n306), .A2(n509), .Y(n750) );
  MUX21X1_HVT U537 ( .A1(n456), .A2(n315), .S0(n413), .Y(n585) );
  MUX21X1_HVT U538 ( .A1(n788), .A2(n216), .S0(n401), .Y(n669) );
  AND2X1_HVT U539 ( .A1(n521), .A2(n457), .Y(n498) );
  MUX21X1_HVT U540 ( .A1(n474), .A2(n785), .S0(n50), .Y(n587) );
  NAND2X0_HVT U541 ( .A1(n580), .A2(n316), .Y(n782) );
  MUX21X1_HVT U542 ( .A1(n790), .A2(n474), .S0(n525), .Y(n765) );
  NBUFFX2_HVT U543 ( .A(in[0]), .Y(n514) );
  NBUFFX2_HVT U544 ( .A(in[0]), .Y(n513) );
  XOR2X1_HVT U545 ( .A1(n507), .A2(n487), .Y(n747) );
endmodule

