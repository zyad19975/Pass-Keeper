
module inv_sbox_14 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n24, n160, n178, n196, n197, n198, n199, n200, n201, n202, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599;

  NAND2X0_HVT U1 ( .A1(n264), .A2(n315), .Y(n599) );
  NAND2X0_HVT U3 ( .A1(n264), .A2(n282), .Y(n597) );
  NAND2X0_HVT U5 ( .A1(n596), .A2(n277), .Y(n595) );
  NAND2X0_HVT U6 ( .A1(n327), .A2(n297), .Y(n593) );
  NAND2X0_HVT U7 ( .A1(n244), .A2(n325), .Y(n592) );
  NAND2X0_HVT U8 ( .A1(n261), .A2(n277), .Y(n591) );
  NAND2X0_HVT U9 ( .A1(n300), .A2(n591), .Y(n590) );
  NAND2X0_HVT U10 ( .A1(n297), .A2(n588), .Y(n589) );
  NAND2X0_HVT U11 ( .A1(n273), .A2(n286), .Y(n587) );
  NAND2X0_HVT U12 ( .A1(n330), .A2(n313), .Y(n586) );
  NAND2X0_HVT U13 ( .A1(n326), .A2(n591), .Y(n585) );
  NAND2X0_HVT U15 ( .A1(n322), .A2(n244), .Y(n583) );
  NAND2X0_HVT U19 ( .A1(n261), .A2(n229), .Y(n578) );
  NAND2X0_HVT U25 ( .A1(n282), .A2(n312), .Y(n594) );
  NAND2X0_HVT U32 ( .A1(n315), .A2(n273), .Y(n567) );
  NAND2X0_HVT U35 ( .A1(n591), .A2(n392), .Y(n564) );
  NAND2X0_HVT U38 ( .A1(n313), .A2(n273), .Y(n561) );
  NAND2X0_HVT U42 ( .A1(n593), .A2(n392), .Y(n557) );
  OA21X1_HVT U53 ( .A1(n256), .A2(n549), .A3(n361), .Y(n547) );
  NAND2X0_HVT U55 ( .A1(n326), .A2(n596), .Y(n545) );
  MUX41X1_HVT U56 ( .A1(n373), .A3(n582), .A2(n359), .A4(n545), .S0(n303), 
        .S1(n260), .Y(n544) );
  AO21X1_HVT U60 ( .A1(n539), .A2(n309), .A3(n577), .Y(n540) );
  MUX41X1_HVT U62 ( .A1(n538), .A3(n544), .A2(n542), .A4(n546), .S0(n321), 
        .S1(n318), .Y(n537) );
  MUX41X1_HVT U65 ( .A1(n353), .A3(n355), .A2(n354), .A4(n561), .S0(n305), 
        .S1(n334), .Y(n534) );
  NAND2X0_HVT U66 ( .A1(n262), .A2(n251), .Y(n533) );
  MUX41X1_HVT U67 ( .A1(n350), .A3(n374), .A2(n352), .A4(n533), .S0(n311), 
        .S1(n303), .Y(n532) );
  MUX41X1_HVT U68 ( .A1(n350), .A3(n264), .A2(n351), .A4(n300), .S0(n305), 
        .S1(n334), .Y(n531) );
  MUX41X1_HVT U69 ( .A1(n531), .A3(n534), .A2(n532), .A4(n535), .S0(n321), 
        .S1(n318), .Y(n530) );
  MUX41X1_HVT U71 ( .A1(n593), .A3(n299), .A2(n587), .A4(n346), .S0(n305), 
        .S1(n335), .Y(n529) );
  NAND2X0_HVT U72 ( .A1(n322), .A2(n592), .Y(n528) );
  MUX41X1_HVT U73 ( .A1(n572), .A3(n528), .A2(n375), .A4(n312), .S0(n310), 
        .S1(n302), .Y(n527) );
  MUX41X1_HVT U74 ( .A1(n589), .A3(n366), .A2(n365), .A4(n356), .S0(n305), 
        .S1(n259), .Y(n526) );
  OA21X1_HVT U76 ( .A1(n339), .A2(n336), .A3(n577), .Y(n524) );
  MUX41X1_HVT U78 ( .A1(n523), .A3(n527), .A2(n526), .A4(n529), .S0(n321), 
        .S1(n318), .Y(n522) );
  MUX41X1_HVT U80 ( .A1(n377), .A3(n373), .A2(n590), .A4(n201), .S0(n305), 
        .S1(n260), .Y(n520) );
  NAND2X0_HVT U81 ( .A1(n286), .A2(n592), .Y(n519) );
  AND2X1_HVT U82 ( .A1(n593), .A2(n324), .Y(n518) );
  MUX41X1_HVT U83 ( .A1(n518), .A3(n363), .A2(n378), .A4(n519), .S0(n305), 
        .S1(n259), .Y(n517) );
  MUX41X1_HVT U84 ( .A1(n295), .A3(n362), .A2(n379), .A4(n574), .S0(n303), 
        .S1(n241), .Y(n516) );
  MUX41X1_HVT U85 ( .A1(n516), .A3(n520), .A2(n517), .A4(n521), .S0(n321), 
        .S1(n318), .Y(n515) );
  MUX41X1_HVT U87 ( .A1(n340), .A3(n295), .A2(n380), .A4(n359), .S0(n304), 
        .S1(n242), .Y(n514) );
  MUX41X1_HVT U88 ( .A1(n352), .A3(n337), .A2(n569), .A4(n553), .S0(n305), 
        .S1(n241), .Y(n513) );
  NAND2X0_HVT U89 ( .A1(n273), .A2(n279), .Y(n512) );
  MUX41X1_HVT U98 ( .A1(n504), .A3(n382), .A2(n367), .A4(n571), .S0(n302), 
        .S1(n334), .Y(n503) );
  MUX41X1_HVT U99 ( .A1(n567), .A3(n354), .A2(n551), .A4(n322), .S0(n260), 
        .S1(n303), .Y(n502) );
  NAND2X0_HVT U100 ( .A1(n273), .A2(n389), .Y(n501) );
  MUX41X1_HVT U101 ( .A1(n383), .A3(n586), .A2(n272), .A4(n501), .S0(n241), 
        .S1(n302), .Y(n500) );
  MUX41X1_HVT U102 ( .A1(n500), .A3(n503), .A2(n502), .A4(n505), .S0(in[5]), 
        .S1(n318), .Y(n499) );
  AND2X1_HVT U104 ( .A1(n592), .A2(n277), .Y(n498) );
  MUX41X1_HVT U105 ( .A1(n584), .A3(n384), .A2(n519), .A4(n498), .S0(n303), 
        .S1(n241), .Y(n497) );
  MUX41X1_HVT U107 ( .A1(n383), .A3(n324), .A2(n496), .A4(n343), .S0(n305), 
        .S1(n259), .Y(n495) );
  MUX41X1_HVT U108 ( .A1(n356), .A3(n266), .A2(n359), .A4(n285), .S0(n302), 
        .S1(n260), .Y(n494) );
  MUX41X1_HVT U109 ( .A1(n382), .A3(n337), .A2(n379), .A4(n371), .S0(n305), 
        .S1(n335), .Y(n493) );
  MUX41X1_HVT U110 ( .A1(n493), .A3(n495), .A2(n494), .A4(n497), .S0(n321), 
        .S1(n271), .Y(n492) );
  AO21X1_HVT U112 ( .A1(n369), .A2(n310), .A3(n575), .Y(n490) );
  NAND2X0_HVT U114 ( .A1(n301), .A2(n592), .Y(n488) );
  MUX41X1_HVT U115 ( .A1(n488), .A3(n587), .A2(n369), .A4(n324), .S0(n334), 
        .S1(n303), .Y(n487) );
  MUX41X1_HVT U116 ( .A1(n368), .A3(n362), .A2(n337), .A4(n583), .S0(n304), 
        .S1(n334), .Y(n486) );
  NAND2X0_HVT U118 ( .A1(n273), .A2(n264), .Y(n484) );
  MUX41X1_HVT U119 ( .A1(n385), .A3(n485), .A2(n562), .A4(n484), .S0(n304), 
        .S1(n259), .Y(n483) );
  MUX41X1_HVT U120 ( .A1(n483), .A3(n487), .A2(n486), .A4(n489), .S0(in[5]), 
        .S1(n271), .Y(n482) );
  MUX41X1_HVT U122 ( .A1(n372), .A3(n291), .A2(n553), .A4(n376), .S0(n304), 
        .S1(n335), .Y(n481) );
  MUX41X1_HVT U124 ( .A1(n293), .A3(n480), .A2(n576), .A4(n280), .S0(n309), 
        .S1(n304), .Y(n479) );
  AOI21X1_HVT U127 ( .A1(n308), .A2(n475), .A3(n344), .Y(n476) );
  NAND2X0_HVT U129 ( .A1(n307), .A2(n300), .Y(n473) );
  MUX41X1_HVT U130 ( .A1(n473), .A3(n474), .A2(n477), .A4(n476), .S0(n311), 
        .S1(n271), .Y(n472) );
  AND2X1_HVT U131 ( .A1(n251), .A2(n252), .Y(n471) );
  MUX41X1_HVT U132 ( .A1(n341), .A3(n471), .A2(n387), .A4(n350), .S0(n310), 
        .S1(n302), .Y(n470) );
  MUX41X1_HVT U133 ( .A1(n388), .A3(n343), .A2(n545), .A4(n342), .S0(n309), 
        .S1(n308), .Y(n469) );
  MUX41X1_HVT U136 ( .A1(n550), .A3(n501), .A2(n467), .A4(n348), .S0(n307), 
        .S1(n242), .Y(n466) );
  MUX41X1_HVT U137 ( .A1(n591), .A3(n570), .A2(n574), .A4(n381), .S0(n311), 
        .S1(n305), .Y(n465) );
  MUX41X1_HVT U139 ( .A1(n464), .A3(n468), .A2(n472), .A4(n478), .S0(n321), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n365), .A3(n292), .A2(n358), .A4(n587), .S0(n310), 
        .S1(n303), .Y(n463) );
  NAND2X0_HVT U141 ( .A1(n322), .A2(n273), .Y(n462) );
  MUX41X1_HVT U142 ( .A1(n462), .A3(n560), .A2(n386), .A4(n358), .S0(n308), 
        .S1(n242), .Y(n461) );
  MUX41X1_HVT U143 ( .A1(n279), .A3(n274), .A2(n578), .A4(n576), .S0(n306), 
        .S1(n242), .Y(n460) );
  MUX41X1_HVT U145 ( .A1(n568), .A3(n384), .A2(n459), .A4(n519), .S0(n308), 
        .S1(n335), .Y(n458) );
  MUX41X1_HVT U146 ( .A1(n458), .A3(n460), .A2(n461), .A4(n463), .S0(n319), 
        .S1(n321), .Y(n457) );
  AO21X1_HVT U148 ( .A1(n311), .A2(n345), .A3(n389), .Y(n455) );
  MUX41X1_HVT U151 ( .A1(n378), .A3(n367), .A2(n287), .A4(n453), .S0(n309), 
        .S1(n303), .Y(n452) );
  OA21X1_HVT U153 ( .A1(n338), .A2(n289), .A3(n347), .Y(n450) );
  MUX41X1_HVT U155 ( .A1(n358), .A3(n587), .A2(n579), .A4(n360), .S0(n306), 
        .S1(n242), .Y(n448) );
  NAND2X0_HVT U159 ( .A1(n444), .A2(n443), .Y(n445) );
  NAND2X0_HVT U163 ( .A1(n262), .A2(n279), .Y(n440) );
  MUX41X1_HVT U164 ( .A1(n590), .A3(n440), .A2(n562), .A4(n356), .S0(n304), 
        .S1(n335), .Y(n439) );
  NAND2X0_HVT U166 ( .A1(n588), .A2(n436), .Y(n437) );
  MUX41X1_HVT U172 ( .A1(n512), .A3(n431), .A2(n290), .A4(n223), .S0(n306), 
        .S1(n260), .Y(n430) );
  NAND2X0_HVT U177 ( .A1(n262), .A2(n264), .Y(n426) );
  MUX41X1_HVT U178 ( .A1(n294), .A3(n426), .A2(n299), .A4(n555), .S0(n306), 
        .S1(n259), .Y(n425) );
  MUX41X1_HVT U182 ( .A1(n343), .A3(n596), .A2(n340), .A4(n378), .S0(n304), 
        .S1(n241), .Y(n422) );
  MUX41X1_HVT U183 ( .A1(n221), .A3(n373), .A2(n356), .A4(n557), .S0(n309), 
        .S1(n302), .Y(n421) );
  AND2X1_HVT U185 ( .A1(n392), .A2(n252), .Y(n419) );
  MUX41X1_HVT U190 ( .A1(n416), .A3(n417), .A2(n415), .A4(n418), .S0(n319), 
        .S1(n302), .Y(n414) );
  NAND2X0_HVT U191 ( .A1(n256), .A2(n349), .Y(n413) );
  AND2X1_HVT U192 ( .A1(n366), .A2(n411), .Y(n412) );
  NAND2X0_HVT U194 ( .A1(n557), .A2(n411), .Y(n409) );
  MUX41X1_HVT U195 ( .A1(n410), .A3(n409), .A2(n412), .A4(n413), .S0(n305), 
        .S1(n319), .Y(n408) );
  NAND2X0_HVT U198 ( .A1(n329), .A2(n392), .Y(n588) );
  NAND2X0_HVT U200 ( .A1(n278), .A2(n252), .Y(n475) );
  AO21X1_HVT U204 ( .A1(n322), .A2(n596), .A3(n289), .Y(n436) );
  AO21X1_HVT U205 ( .A1(n252), .A2(n300), .A3(n289), .Y(n443) );
  NAND2X0_HVT U207 ( .A1(n252), .A2(n298), .Y(n539) );
  MUX21X2_HVT U2 ( .A1(n344), .A2(n558), .S0(n311), .Y(n491) );
  MUX21X2_HVT U4 ( .A1(n375), .A2(n558), .S0(n310), .Y(n416) );
  INVX1_HVT U14 ( .A(n324), .Y(n391) );
  INVX1_HVT U16 ( .A(n582), .Y(n224) );
  MUX41X1_HVT U17 ( .A1(n449), .A3(n454), .A2(n448), .A4(n452), .S0(n321), 
        .S1(n317), .Y(n447) );
  IBUFFX2_HVT U18 ( .A(n317), .Y(n271) );
  INVX1_HVT U20 ( .A(n394), .Y(n387) );
  INVX2_HVT U21 ( .A(n320), .Y(n321) );
  MUX21X1_HVT U22 ( .A1(n280), .A2(n545), .S0(n310), .Y(n541) );
  MUX21X2_HVT U23 ( .A1(n424), .A2(n425), .S0(n271), .Y(n423) );
  MUX21X2_HVT U24 ( .A1(n525), .A2(n524), .S0(n308), .Y(n523) );
  MUX21X2_HVT U26 ( .A1(n376), .A2(n254), .S0(n311), .Y(n525) );
  NAND2X0_HVT U27 ( .A1(n325), .A2(n24), .Y(n160) );
  NAND2X0_HVT U28 ( .A1(n510), .A2(n228), .Y(n178) );
  NAND2X0_HVT U29 ( .A1(n160), .A2(n178), .Y(n509) );
  INVX0_HVT U30 ( .A(n228), .Y(n24) );
  MUX21X1_HVT U31 ( .A1(n323), .A2(n316), .S0(n310), .Y(n510) );
  IBUFFX2_HVT U33 ( .A(n262), .Y(n228) );
  NBUFFX2_HVT U34 ( .A(n258), .Y(n310) );
  MUX21X1_HVT U36 ( .A1(n446), .A2(n445), .S0(n233), .Y(n442) );
  MUX21X1_HVT U37 ( .A1(n325), .A2(n275), .S0(n273), .Y(n274) );
  MUX21X2_HVT U39 ( .A1(n387), .A2(n341), .S0(n309), .Y(n456) );
  INVX2_HVT U40 ( .A(n390), .Y(n301) );
  NAND2X1_HVT U41 ( .A1(n530), .A2(n196), .Y(n197) );
  NAND2X0_HVT U43 ( .A1(n537), .A2(in[7]), .Y(n198) );
  NAND2X0_HVT U44 ( .A1(n197), .A2(n198), .Y(out[0]) );
  IBUFFX2_HVT U45 ( .A(in[7]), .Y(n196) );
  MUX21X1_HVT U46 ( .A1(n313), .A2(n265), .S0(n252), .Y(n280) );
  INVX1_HVT U47 ( .A(n261), .Y(n252) );
  INVX0_HVT U48 ( .A(n223), .Y(n287) );
  MUX21X2_HVT U49 ( .A1(n541), .A2(n540), .S0(n307), .Y(n538) );
  MUX41X1_HVT U50 ( .A1(n420), .A3(n423), .A2(n408), .A4(n414), .S0(in[5]), 
        .S1(n199), .Y(out[7]) );
  IBUFFX16_HVT U51 ( .A(in[7]), .Y(n199) );
  MUX21X2_HVT U52 ( .A1(n499), .A2(n506), .S0(n200), .Y(out[2]) );
  IBUFFX16_HVT U54 ( .A(n240), .Y(n200) );
  NBUFFX2_HVT U57 ( .A(n595), .Y(n201) );
  NAND2X2_HVT U58 ( .A1(n262), .A2(n265), .Y(n596) );
  MUX21X2_HVT U59 ( .A1(n456), .A2(n455), .S0(n307), .Y(n454) );
  MUX21X1_HVT U61 ( .A1(n287), .A2(n596), .S0(n307), .Y(n536) );
  NAND2X0_HVT U63 ( .A1(n295), .A2(n202), .Y(n218) );
  NAND2X0_HVT U64 ( .A1(n551), .A2(n311), .Y(n219) );
  NAND2X0_HVT U70 ( .A1(n218), .A2(n219), .Y(n417) );
  IBUFFX2_HVT U75 ( .A(n311), .Y(n202) );
  XOR2X1_HVT U77 ( .A1(n278), .A2(n245), .Y(n551) );
  MUX21X1_HVT U79 ( .A1(n419), .A2(n377), .S0(n309), .Y(n418) );
  IBUFFX2_HVT U86 ( .A(n331), .Y(n245) );
  INVX1_HVT U90 ( .A(n555), .Y(n370) );
  MUX21X2_HVT U91 ( .A1(n279), .A2(n299), .S0(n330), .Y(n555) );
  MUX41X1_HVT U92 ( .A1(n513), .A3(n507), .A2(n514), .A4(n511), .S0(n320), 
        .S1(n220), .Y(n506) );
  IBUFFX16_HVT U93 ( .A(n317), .Y(n220) );
  INVX0_HVT U94 ( .A(n556), .Y(n221) );
  MUX21X2_HVT U95 ( .A1(n492), .A2(n482), .S0(n222), .Y(out[3]) );
  IBUFFX16_HVT U96 ( .A(in[7]), .Y(n222) );
  MUX21X1_HVT U97 ( .A1(n282), .A2(n391), .S0(n244), .Y(n558) );
  MUX21X1_HVT U103 ( .A1(n224), .A2(n225), .S0(n329), .Y(n223) );
  IBUFFX16_HVT U106 ( .A(n265), .Y(n225) );
  INVX2_HVT U111 ( .A(n309), .Y(n256) );
  OA21X1_HVT U113 ( .A1(n362), .A2(n256), .A3(n539), .Y(n415) );
  IBUFFX2_HVT U117 ( .A(n331), .Y(n244) );
  AO21X2_HVT U121 ( .A1(n329), .A2(n389), .A3(n256), .Y(n411) );
  INVX0_HVT U123 ( .A(n310), .Y(n230) );
  IBUFFX2_HVT U125 ( .A(n331), .Y(n329) );
  IBUFFX2_HVT U126 ( .A(n390), .Y(n226) );
  INVX1_HVT U128 ( .A(n226), .Y(n227) );
  INVX0_HVT U134 ( .A(n324), .Y(n229) );
  INVX2_HVT U135 ( .A(n263), .Y(n264) );
  INVX1_HVT U138 ( .A(n331), .Y(n328) );
  NAND2X1_HVT U144 ( .A1(n556), .A2(n230), .Y(n231) );
  NAND2X0_HVT U147 ( .A1(n376), .A2(n310), .Y(n232) );
  NAND2X0_HVT U149 ( .A1(n231), .A2(n232), .Y(n446) );
  IBUFFX16_HVT U150 ( .A(n308), .Y(n233) );
  NAND2X0_HVT U152 ( .A1(n427), .A2(n234), .Y(n235) );
  NAND2X0_HVT U154 ( .A1(n434), .A2(in[7]), .Y(n236) );
  NAND2X0_HVT U156 ( .A1(n235), .A2(n236), .Y(out[6]) );
  IBUFFX2_HVT U157 ( .A(in[7]), .Y(n234) );
  INVX1_HVT U158 ( .A(n331), .Y(n262) );
  NAND2X1_HVT U160 ( .A1(n508), .A2(n237), .Y(n238) );
  NAND2X0_HVT U161 ( .A1(n509), .A2(n307), .Y(n239) );
  NAND2X0_HVT U162 ( .A1(n238), .A2(n239), .Y(n507) );
  IBUFFX2_HVT U165 ( .A(n307), .Y(n237) );
  IBUFFX16_HVT U167 ( .A(in[7]), .Y(n240) );
  MUX21X1_HVT U168 ( .A1(n346), .A2(n322), .S0(n311), .Y(n508) );
  INVX0_HVT U169 ( .A(n331), .Y(n261) );
  INVX0_HVT U170 ( .A(n331), .Y(n327) );
  XNOR2X1_HVT U171 ( .A1(n314), .A2(n263), .Y(n582) );
  INVX1_HVT U173 ( .A(n258), .Y(n289) );
  INVX1_HVT U174 ( .A(n336), .Y(n241) );
  INVX1_HVT U175 ( .A(n336), .Y(n242) );
  MUX41X1_HVT U176 ( .A1(n290), .A3(n294), .A2(n433), .A4(n293), .S0(n243), 
        .S1(n334), .Y(n432) );
  IBUFFX16_HVT U179 ( .A(n306), .Y(n243) );
  INVX1_HVT U180 ( .A(in[4]), .Y(n336) );
  NAND2X0_HVT U181 ( .A1(n421), .A2(n246), .Y(n247) );
  NAND2X0_HVT U184 ( .A1(n422), .A2(n319), .Y(n248) );
  NAND2X0_HVT U186 ( .A1(n247), .A2(n248), .Y(n420) );
  IBUFFX2_HVT U187 ( .A(n319), .Y(n246) );
  INVX1_HVT U188 ( .A(n336), .Y(n334) );
  INVX1_HVT U189 ( .A(n336), .Y(n259) );
  INVX0_HVT U193 ( .A(in[7]), .Y(n249) );
  INVX0_HVT U196 ( .A(n317), .Y(n318) );
  INVX1_HVT U197 ( .A(in[1]), .Y(n317) );
  INVX0_HVT U199 ( .A(n272), .Y(n563) );
  INVX0_HVT U201 ( .A(in[5]), .Y(n320) );
  INVX1_HVT U202 ( .A(n598), .Y(n389) );
  INVX1_HVT U203 ( .A(n599), .Y(n390) );
  IBUFFX2_HVT U206 ( .A(n593), .Y(n342) );
  IBUFFX2_HVT U208 ( .A(n571), .Y(n361) );
  MUX21X2_HVT U209 ( .A1(n457), .A2(n447), .S0(n249), .Y(out[5]) );
  IBUFFX2_HVT U210 ( .A(n596), .Y(n340) );
  INVX1_HVT U211 ( .A(n594), .Y(n279) );
  INVX0_HVT U212 ( .A(n574), .Y(n358) );
  INVX0_HVT U213 ( .A(n253), .Y(n424) );
  INVX1_HVT U214 ( .A(n306), .Y(n288) );
  INVX1_HVT U215 ( .A(n390), .Y(n297) );
  INVX1_HVT U216 ( .A(n261), .Y(n273) );
  INVX1_HVT U217 ( .A(n577), .Y(n356) );
  INVX1_HVT U218 ( .A(n554), .Y(n255) );
  INVX1_HVT U219 ( .A(n301), .Y(n299) );
  INVX1_HVT U220 ( .A(in[3]), .Y(n263) );
  INVX0_HVT U221 ( .A(n567), .Y(n254) );
  INVX1_HVT U222 ( .A(n276), .Y(n278) );
  INVX1_HVT U223 ( .A(n282), .Y(n250) );
  INVX2_HVT U224 ( .A(n250), .Y(n251) );
  INVX1_HVT U225 ( .A(n281), .Y(n282) );
  MUX41X1_HVT U226 ( .A1(n255), .A3(n257), .A2(n587), .A4(n254), .S0(n288), 
        .S1(n256), .Y(n253) );
  NAND2X0_HVT U227 ( .A1(n593), .A2(n278), .Y(n257) );
  INVX1_HVT U228 ( .A(in[0]), .Y(n331) );
  MUX21X1_HVT U229 ( .A1(n389), .A2(n315), .S0(n252), .Y(n573) );
  XOR2X1_HVT U230 ( .A1(n300), .A2(n330), .Y(n562) );
  MUX41X1_HVT U231 ( .A1(n430), .A3(n432), .A2(n428), .A4(n429), .S0(n271), 
        .S1(n320), .Y(n427) );
  INVX0_HVT U232 ( .A(n274), .Y(n556) );
  NBUFFX2_HVT U233 ( .A(in[4]), .Y(n258) );
  MUX21X1_HVT U234 ( .A1(n574), .A2(n295), .S0(n310), .Y(n451) );
  IBUFFX2_HVT U235 ( .A(n336), .Y(n260) );
  IBUFFX2_HVT U236 ( .A(n336), .Y(n335) );
  MUX21X1_HVT U237 ( .A1(n298), .A2(n316), .S0(n328), .Y(n431) );
  MUX41X1_HVT U238 ( .A1(n512), .A3(n552), .A2(n592), .A4(n227), .S0(n288), 
        .S1(n336), .Y(n511) );
  MUX21X1_HVT U239 ( .A1(n229), .A2(n227), .S0(n252), .Y(n433) );
  INVX0_HVT U240 ( .A(n331), .Y(n330) );
  MUX41X1_HVT U241 ( .A1(n381), .A3(n360), .A2(n585), .A4(n374), .S0(n288), 
        .S1(n256), .Y(n505) );
  MUX41X1_HVT U242 ( .A1(n581), .A3(n364), .A2(n580), .A4(n362), .S0(n288), 
        .S1(n289), .Y(n521) );
  MUX21X2_HVT U243 ( .A1(n515), .A2(n522), .S0(in[7]), .Y(out[1]) );
  NAND2X0_HVT U244 ( .A1(n312), .A2(n283), .Y(n265) );
  INVX0_HVT U245 ( .A(n598), .Y(n284) );
  MUX21X2_HVT U246 ( .A1(n360), .A2(n351), .S0(n311), .Y(n548) );
  INVX0_HVT U247 ( .A(n270), .Y(n266) );
  INVX0_HVT U248 ( .A(n313), .Y(n275) );
  MUX21X1_HVT U249 ( .A1(n278), .A2(n326), .S0(n262), .Y(n267) );
  NAND2X0_HVT U250 ( .A1(n437), .A2(n288), .Y(n268) );
  NAND2X0_HVT U251 ( .A1(n438), .A2(n307), .Y(n269) );
  NAND2X0_HVT U252 ( .A1(n268), .A2(n269), .Y(n435) );
  MUX21X1_HVT U253 ( .A1(n576), .A2(n573), .S0(n289), .Y(n438) );
  INVX0_HVT U254 ( .A(n594), .Y(n276) );
  NBUFFX2_HVT U255 ( .A(n392), .Y(n270) );
  INVX0_HVT U256 ( .A(n582), .Y(n392) );
  MUX41X1_HVT U257 ( .A1(n564), .A3(n267), .A2(n370), .A4(n355), .S0(n306), 
        .S1(n289), .Y(n441) );
  MUX41X1_HVT U258 ( .A1(n545), .A3(n380), .A2(n270), .A4(n388), .S0(n288), 
        .S1(n258), .Y(n428) );
  MUX21X1_HVT U259 ( .A1(n251), .A2(n323), .S0(n327), .Y(n272) );
  INVX1_HVT U260 ( .A(n400), .Y(n380) );
  MUX41X1_HVT U261 ( .A1(n439), .A3(n442), .A2(n435), .A4(n441), .S0(n321), 
        .S1(n317), .Y(n434) );
  MUX21X1_HVT U262 ( .A1(n313), .A2(n582), .S0(n252), .Y(n577) );
  INVX1_HVT U263 ( .A(n404), .Y(n376) );
  IBUFFX2_HVT U264 ( .A(n573), .Y(n359) );
  INVX0_HVT U265 ( .A(n280), .Y(n576) );
  INVX1_HVT U266 ( .A(n276), .Y(n277) );
  MUX21X1_HVT U267 ( .A1(n323), .A2(n316), .S0(n261), .Y(n574) );
  INVX0_HVT U268 ( .A(in[6]), .Y(n281) );
  NBUFFX2_HVT U269 ( .A(n281), .Y(n283) );
  MUX41X1_HVT U270 ( .A1(n563), .A3(n298), .A2(n286), .A4(n300), .S0(n289), 
        .S1(n288), .Y(n429) );
  INVX0_HVT U271 ( .A(n284), .Y(n285) );
  INVX0_HVT U272 ( .A(n284), .Y(n286) );
  INVX1_HVT U273 ( .A(n402), .Y(n378) );
  MUX21X2_HVT U274 ( .A1(n450), .A2(n451), .S0(n308), .Y(n449) );
  MUX21X2_HVT U275 ( .A1(n548), .A2(n547), .S0(n307), .Y(n546) );
  AND2X1_HVT U276 ( .A1(n593), .A2(n598), .Y(n290) );
  AND2X1_HVT U277 ( .A1(n285), .A2(n583), .Y(n291) );
  MUX21X1_HVT U278 ( .A1(n255), .A2(n293), .S0(n309), .Y(n410) );
  MUX21X1_HVT U279 ( .A1(n356), .A2(n536), .S0(n296), .Y(n535) );
  MUX21X1_HVT U280 ( .A1(n284), .A2(n392), .S0(n329), .Y(n566) );
  MUX21X1_HVT U281 ( .A1(n270), .A2(n316), .S0(n329), .Y(n395) );
  MUX21X1_HVT U282 ( .A1(n284), .A2(n315), .S0(n262), .Y(n405) );
  MUX21X1_HVT U283 ( .A1(n283), .A2(n279), .S0(n327), .Y(n453) );
  NAND2X0_HVT U284 ( .A1(n312), .A2(n283), .Y(n598) );
  MUX21X1_HVT U285 ( .A1(n270), .A2(n313), .S0(n328), .Y(n560) );
  MUX21X1_HVT U286 ( .A1(n298), .A2(n323), .S0(n245), .Y(n400) );
  MUX21X1_HVT U287 ( .A1(n313), .A2(n389), .S0(n262), .Y(n569) );
  MUX21X1_HVT U288 ( .A1(n386), .A2(n292), .S0(n307), .Y(n477) );
  MUX21X1_HVT U289 ( .A1(n566), .A2(n291), .S0(n308), .Y(n474) );
  MUX21X1_HVT U290 ( .A1(n322), .A2(n298), .S0(n245), .Y(n568) );
  MUX21X1_HVT U291 ( .A1(n389), .A2(n391), .S0(n244), .Y(n549) );
  MUX21X1_HVT U292 ( .A1(n283), .A2(n265), .S0(n245), .Y(n496) );
  XOR2X1_HVT U293 ( .A1(n323), .A2(n245), .Y(n553) );
  MUX21X1_HVT U294 ( .A1(n391), .A2(n313), .S0(n245), .Y(n404) );
  MUX21X1_HVT U295 ( .A1(n322), .A2(n279), .S0(n330), .Y(n565) );
  MUX21X1_HVT U296 ( .A1(n326), .A2(n286), .S0(n244), .Y(n580) );
  MUX21X1_HVT U297 ( .A1(n313), .A2(n285), .S0(n328), .Y(n403) );
  XNOR2X1_HVT U298 ( .A1(n286), .A2(n329), .Y(n292) );
  MUX21X1_HVT U299 ( .A1(n277), .A2(n285), .S0(n329), .Y(n394) );
  MUX21X1_HVT U300 ( .A1(n283), .A2(n322), .S0(n328), .Y(n559) );
  MUX21X1_HVT U301 ( .A1(n299), .A2(n279), .S0(n244), .Y(n571) );
  MUX21X1_HVT U302 ( .A1(n301), .A2(n286), .S0(n244), .Y(n584) );
  MUX21X1_HVT U303 ( .A1(n325), .A2(n313), .S0(n330), .Y(n579) );
  MUX21X1_HVT U304 ( .A1(n313), .A2(n315), .S0(n328), .Y(n554) );
  XOR2X1_HVT U305 ( .A1(n324), .A2(n327), .Y(n552) );
  AND2X1_HVT U306 ( .A1(n327), .A2(n316), .Y(n293) );
  MUX21X1_HVT U307 ( .A1(n312), .A2(n325), .S0(n330), .Y(n397) );
  NBUFFX2_HVT U308 ( .A(n258), .Y(n311) );
  NBUFFX2_HVT U309 ( .A(n258), .Y(n309) );
  NBUFFX2_HVT U310 ( .A(n281), .Y(n314) );
  NBUFFX2_HVT U311 ( .A(n582), .Y(n322) );
  NBUFFX2_HVT U312 ( .A(n582), .Y(n323) );
  NBUFFX2_HVT U313 ( .A(n314), .Y(n315) );
  MUX21X1_HVT U314 ( .A1(n479), .A2(n481), .S0(n319), .Y(n478) );
  MUX21X1_HVT U315 ( .A1(n326), .A2(n315), .S0(n261), .Y(n480) );
  MUX21X1_HVT U316 ( .A1(n357), .A2(n543), .S0(n296), .Y(n542) );
  MUX21X1_HVT U317 ( .A1(n358), .A2(n595), .S0(n308), .Y(n543) );
  AND2X1_HVT U318 ( .A1(n229), .A2(n273), .Y(n294) );
  MUX21X1_HVT U319 ( .A1(n285), .A2(n277), .S0(n245), .Y(n459) );
  NBUFFX2_HVT U320 ( .A(n597), .Y(n324) );
  AND2X1_HVT U321 ( .A1(n326), .A2(n273), .Y(n295) );
  MUX21X1_HVT U322 ( .A1(n490), .A2(n491), .S0(n308), .Y(n489) );
  NBUFFX2_HVT U323 ( .A(n597), .Y(n326) );
  NBUFFX2_HVT U324 ( .A(n597), .Y(n325) );
  NBUFFX2_HVT U325 ( .A(n283), .Y(n316) );
  NBUFFX2_HVT U326 ( .A(n263), .Y(n312) );
  NBUFFX2_HVT U327 ( .A(n263), .Y(n313) );
  NBUFFX2_HVT U328 ( .A(n332), .Y(n306) );
  NBUFFX2_HVT U329 ( .A(n333), .Y(n308) );
  NBUFFX2_HVT U330 ( .A(n333), .Y(n307) );
  XNOR2X1_HVT U331 ( .A1(n289), .A2(n304), .Y(n296) );
  NBUFFX2_HVT U332 ( .A(n333), .Y(n304) );
  NBUFFX2_HVT U333 ( .A(n333), .Y(n305) );
  NBUFFX2_HVT U334 ( .A(n332), .Y(n302) );
  NBUFFX2_HVT U335 ( .A(n332), .Y(n303) );
  INVX1_HVT U336 ( .A(n317), .Y(n319) );
  MUX21X1_HVT U337 ( .A1(n465), .A2(n466), .S0(n319), .Y(n464) );
  MUX21X1_HVT U338 ( .A1(n469), .A2(n470), .S0(n271), .Y(n468) );
  MUX21X1_HVT U339 ( .A1(n299), .A2(n264), .S0(n328), .Y(n393) );
  MUX21X1_HVT U340 ( .A1(n301), .A2(n264), .S0(n329), .Y(n444) );
  MUX21X1_HVT U341 ( .A1(n277), .A2(n264), .S0(n244), .Y(n504) );
  MUX21X1_HVT U342 ( .A1(n316), .A2(n264), .S0(n330), .Y(n572) );
  MUX21X1_HVT U343 ( .A1(n229), .A2(n279), .S0(n328), .Y(n485) );
  MUX21X1_HVT U344 ( .A1(n264), .A2(n300), .S0(n329), .Y(n399) );
  MUX21X1_HVT U345 ( .A1(n264), .A2(n278), .S0(n244), .Y(n398) );
  NBUFFX2_HVT U346 ( .A(in[2]), .Y(n333) );
  NBUFFX2_HVT U347 ( .A(in[2]), .Y(n332) );
  MUX21X1_HVT U348 ( .A1(n389), .A2(n251), .S0(n327), .Y(n467) );
  XOR2X1_HVT U349 ( .A1(n245), .A2(n251), .Y(n550) );
  MUX21X1_HVT U350 ( .A1(n251), .A2(n298), .S0(n245), .Y(n575) );
  MUX21X1_HVT U351 ( .A1(n325), .A2(n251), .S0(n328), .Y(n401) );
  MUX21X1_HVT U352 ( .A1(n282), .A2(n326), .S0(n327), .Y(n406) );
  MUX21X1_HVT U353 ( .A1(n312), .A2(n251), .S0(n327), .Y(n396) );
  MUX21X1_HVT U354 ( .A1(n251), .A2(n301), .S0(n330), .Y(n581) );
  MUX21X1_HVT U355 ( .A1(n278), .A2(n282), .S0(n328), .Y(n570) );
  MUX21X1_HVT U356 ( .A1(n282), .A2(n279), .S0(n262), .Y(n407) );
  MUX21X1_HVT U357 ( .A1(n312), .A2(n392), .S0(n327), .Y(n402) );
  INVX1_HVT U358 ( .A(n297), .Y(n298) );
  INVX0_HVT U359 ( .A(n390), .Y(n300) );
  INVX0_HVT U360 ( .A(n561), .Y(n337) );
  INVX0_HVT U361 ( .A(n501), .Y(n338) );
  INVX0_HVT U362 ( .A(n462), .Y(n339) );
  INVX0_HVT U363 ( .A(n595), .Y(n341) );
  INVX0_HVT U364 ( .A(n557), .Y(n343) );
  INVX0_HVT U365 ( .A(n592), .Y(n344) );
  INVX0_HVT U366 ( .A(n591), .Y(n345) );
  INVX0_HVT U367 ( .A(n564), .Y(n346) );
  INVX0_HVT U368 ( .A(n585), .Y(n347) );
  INVX0_HVT U369 ( .A(n590), .Y(n348) );
  INVX0_HVT U370 ( .A(n586), .Y(n349) );
  INVX0_HVT U371 ( .A(n584), .Y(n350) );
  INVX0_HVT U372 ( .A(n583), .Y(n351) );
  INVX0_HVT U373 ( .A(n581), .Y(n352) );
  INVX0_HVT U374 ( .A(n580), .Y(n353) );
  INVX0_HVT U375 ( .A(n579), .Y(n354) );
  INVX0_HVT U376 ( .A(n578), .Y(n355) );
  INVX0_HVT U377 ( .A(n575), .Y(n357) );
  INVX0_HVT U378 ( .A(n572), .Y(n360) );
  INVX0_HVT U379 ( .A(n570), .Y(n362) );
  INVX0_HVT U380 ( .A(n569), .Y(n363) );
  INVX0_HVT U381 ( .A(n568), .Y(n364) );
  INVX0_HVT U382 ( .A(n566), .Y(n365) );
  INVX0_HVT U383 ( .A(n565), .Y(n366) );
  INVX0_HVT U384 ( .A(n562), .Y(n367) );
  INVX0_HVT U385 ( .A(n560), .Y(n368) );
  INVX0_HVT U386 ( .A(n559), .Y(n369) );
  INVX0_HVT U387 ( .A(n553), .Y(n371) );
  INVX0_HVT U388 ( .A(n589), .Y(n372) );
  INVX0_HVT U389 ( .A(n407), .Y(n373) );
  INVX0_HVT U390 ( .A(n406), .Y(n374) );
  INVX0_HVT U391 ( .A(n405), .Y(n375) );
  INVX0_HVT U392 ( .A(n403), .Y(n377) );
  INVX0_HVT U393 ( .A(n401), .Y(n379) );
  INVX0_HVT U394 ( .A(n399), .Y(n381) );
  INVX0_HVT U395 ( .A(n398), .Y(n382) );
  INVX0_HVT U396 ( .A(n397), .Y(n383) );
  INVX0_HVT U397 ( .A(n396), .Y(n384) );
  INVX0_HVT U398 ( .A(n444), .Y(n385) );
  INVX0_HVT U399 ( .A(n395), .Y(n386) );
  INVX0_HVT U400 ( .A(n393), .Y(n388) );
endmodule

