
module sbox_3 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n10, n23, n38, n50, n65, n113, n114, n117, n118, n119, n210, n211,
         n212, n213, n216, n217, n218, n219, n222, n224, n225, n229, n231,
         n232, n236, n238, n240, n245, n246, n252, n253, n256, n259, n261,
         n264, n271, n274, n275, n278, n280, n282, n283, n288, n290, n293,
         n297, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748;

  NAND2X0_HVT U4 ( .A1(n375), .A2(n306), .Y(n745) );
  NAND2X0_HVT U5 ( .A1(n393), .A2(n390), .Y(n743) );
  NAND2X0_HVT U15 ( .A1(n746), .A2(n364), .Y(n734) );
  NAND2X0_HVT U21 ( .A1(n375), .A2(n486), .Y(n728) );
  NAND2X0_HVT U42 ( .A1(n484), .A2(n417), .Y(n709) );
  MUX41X1_HVT U51 ( .A1(n500), .A3(n522), .A2(n494), .A4(n502), .S0(n474), 
        .S1(n347), .Y(n701) );
  NAND2X0_HVT U53 ( .A1(n698), .A2(n708), .Y(n699) );
  NAND2X0_HVT U56 ( .A1(n374), .A2(n694), .Y(n695) );
  NAND2X0_HVT U58 ( .A1(n245), .A2(n746), .Y(n692) );
  MUX41X1_HVT U61 ( .A1(n459), .A3(n529), .A2(n506), .A4(n259), .S0(n491), 
        .S1(n402), .Y(n689) );
  AO21X1_HVT U66 ( .A1(n534), .A2(n470), .A3(n536), .Y(n685) );
  MUX41X1_HVT U68 ( .A1(n505), .A3(n685), .A2(n684), .A4(n686), .S0(n468), 
        .S1(n437), .Y(n683) );
  NAND2X0_HVT U73 ( .A1(n409), .A2(n678), .Y(n679) );
  MUX41X1_HVT U74 ( .A1(n680), .A3(n724), .A2(n679), .A4(n726), .S0(n325), 
        .S1(n240), .Y(n677) );
  AND2X1_HVT U83 ( .A1(n483), .A2(n408), .Y(n667) );
  MUX41X1_HVT U84 ( .A1(n507), .A3(n312), .A2(n733), .A4(n667), .S0(n380), 
        .S1(n490), .Y(n666) );
  NAND2X0_HVT U85 ( .A1(n486), .A2(n382), .Y(n665) );
  NAND2X0_HVT U101 ( .A1(n648), .A2(n647), .Y(n649) );
  MUX41X1_HVT U103 ( .A1(n306), .A3(n523), .A2(n513), .A4(n715), .S0(n379), 
        .S1(n449), .Y(n645) );
  NAND2X0_HVT U110 ( .A1(n481), .A2(n640), .Y(n641) );
  AND2X1_HVT U115 ( .A1(n393), .A2(n364), .Y(n638) );
  NAND2X0_HVT U123 ( .A1(n628), .A2(n629), .Y(n630) );
  MUX41X1_HVT U125 ( .A1(n728), .A3(n463), .A2(n505), .A4(n517), .S0(n325), 
        .S1(n449), .Y(n626) );
  MUX41X1_HVT U136 ( .A1(n456), .A3(n717), .A2(n499), .A4(n714), .S0(n380), 
        .S1(n437), .Y(n616) );
  AND2X1_HVT U140 ( .A1(n414), .A2(n422), .Y(n612) );
  MUX41X1_HVT U141 ( .A1(n725), .A3(n515), .A2(n612), .A4(n305), .S0(n314), 
        .S1(n473), .Y(n611) );
  MUX41X1_HVT U142 ( .A1(n507), .A3(n259), .A2(n520), .A4(n414), .S0(n469), 
        .S1(n491), .Y(n610) );
  NAND2X0_HVT U146 ( .A1(n117), .A2(n311), .Y(n678) );
  AND2X1_HVT U154 ( .A1(n473), .A2(n400), .Y(n599) );
  NAND2X0_HVT U158 ( .A1(n484), .A2(n346), .Y(n595) );
  MUX41X1_HVT U159 ( .A1(n737), .A3(n364), .A2(n595), .A4(n537), .S0(n469), 
        .S1(n240), .Y(n594) );
  AND2X1_HVT U162 ( .A1(n312), .A2(n678), .Y(n591) );
  NAND2X0_HVT U166 ( .A1(n341), .A2(n322), .Y(n587) );
  NAND2X0_HVT U167 ( .A1(n308), .A2(n486), .Y(n586) );
  MUX41X1_HVT U168 ( .A1(n510), .A3(n414), .A2(n586), .A4(n587), .S0(n380), 
        .S1(n437), .Y(n585) );
  MUX41X1_HVT U172 ( .A1(n582), .A3(n588), .A2(n585), .A4(n590), .S0(in[0]), 
        .S1(n470), .Y(n581) );
  MUX41X1_HVT U176 ( .A1(n479), .A3(n580), .A2(n508), .A4(n736), .S0(n449), 
        .S1(n395), .Y(n579) );
  NAND2X0_HVT U177 ( .A1(n399), .A2(n478), .Y(n578) );
  MUX41X1_HVT U178 ( .A1(n732), .A3(n578), .A2(n324), .A4(n713), .S0(n314), 
        .S1(n240), .Y(n577) );
  MUX41X1_HVT U182 ( .A1(n516), .A3(n374), .A2(n501), .A4(n524), .S0(n474), 
        .S1(n333), .Y(n573) );
  MUX41X1_HVT U189 ( .A1(n567), .A3(n736), .A2(n568), .A4(n521), .S0(n449), 
        .S1(n333), .Y(n566) );
  MUX41X1_HVT U194 ( .A1(n710), .A3(n723), .A2(n509), .A4(n410), .S0(n449), 
        .S1(n395), .Y(n562) );
  AO21X1_HVT U197 ( .A1(n460), .A2(n449), .A3(n530), .Y(n559) );
  MUX41X1_HVT U203 ( .A1(n714), .A3(n496), .A2(n738), .A4(n718), .S0(n395), 
        .S1(n490), .Y(n553) );
  NAND2X0_HVT U208 ( .A1(n425), .A2(n375), .Y(n640) );
  NAND2X0_HVT U212 ( .A1(n482), .A2(n409), .Y(n694) );
  NAND2X0_HVT U214 ( .A1(n312), .A2(n486), .Y(n549) );
  NAND2X0_HVT U215 ( .A1(n640), .A2(n416), .Y(n548) );
  NAND2X0_HVT U218 ( .A1(n412), .A2(n399), .Y(n602) );
  NAND2X0_HVT U220 ( .A1(n474), .A2(n549), .Y(n670) );
  INVX0_HVT U245 ( .A(n743), .Y(n537) );
  INVX0_HVT U255 ( .A(n545), .Y(n531) );
  INVX0_HVT U256 ( .A(n602), .Y(n530) );
  INVX0_HVT U262 ( .A(n541), .Y(n526) );
  INVX0_HVT U265 ( .A(n724), .Y(n524) );
  INVX0_HVT U268 ( .A(n728), .Y(n522) );
  INVX0_HVT U270 ( .A(n548), .Y(n521) );
  INVX0_HVT U271 ( .A(n640), .Y(n520) );
  INVX0_HVT U278 ( .A(n717), .Y(n514) );
  INVX0_HVT U280 ( .A(n721), .Y(n513) );
  INVX0_HVT U284 ( .A(n549), .Y(n511) );
  INVX0_HVT U289 ( .A(n647), .Y(n508) );
  INVX0_HVT U293 ( .A(n733), .Y(n506) );
  INVX0_HVT U294 ( .A(n741), .Y(n505) );
  INVX0_HVT U295 ( .A(n745), .Y(n504) );
  INVX0_HVT U297 ( .A(n746), .Y(n503) );
  INVX0_HVT U303 ( .A(n542), .Y(n499) );
  INVX0_HVT U306 ( .A(n586), .Y(n497) );
  INVX0_HVT U309 ( .A(n730), .Y(n494) );
  MUX21X1_HVT U1 ( .A1(n409), .A2(n479), .S0(n393), .Y(n680) );
  AO21X1_HVT U2 ( .A1(n333), .A2(n414), .A3(n312), .Y(n635) );
  MUX21X1_HVT U3 ( .A1(n403), .A2(n535), .S0(n468), .Y(n636) );
  INVX1_HVT U6 ( .A(n423), .Y(n482) );
  AND3X1_HVT U7 ( .A1(n469), .A2(n486), .A3(n408), .Y(n623) );
  NBUFFX2_HVT U8 ( .A(in[5]), .Y(n470) );
  INVX1_HVT U9 ( .A(n219), .Y(n742) );
  AND2X1_HVT U10 ( .A1(n404), .A2(n318), .Y(n10) );
  AND2X1_HVT U11 ( .A1(n486), .A2(n481), .Y(n23) );
  AND2X1_HVT U12 ( .A1(n351), .A2(n252), .Y(n38) );
  INVX1_HVT U13 ( .A(in[7]), .Y(n493) );
  INVX1_HVT U14 ( .A(n472), .Y(n433) );
  INVX1_HVT U16 ( .A(n490), .Y(n429) );
  INVX1_HVT U17 ( .A(n311), .Y(n382) );
  MUX21X2_HVT U18 ( .A1(n476), .A2(n372), .S0(n399), .Y(n655) );
  MUX21X1_HVT U19 ( .A1(n503), .A2(n714), .S0(n222), .Y(n50) );
  NBUFFX2_HVT U20 ( .A(n525), .Y(n381) );
  MUX21X2_HVT U22 ( .A1(n404), .A2(n368), .S0(n394), .Y(n714) );
  XOR2X2_HVT U23 ( .A1(n518), .A2(n405), .Y(n457) );
  MUX21X2_HVT U24 ( .A1(n65), .A2(n619), .S0(n469), .Y(n618) );
  INVX1_HVT U25 ( .A(n400), .Y(n224) );
  AND3X1_HVT U26 ( .A1(n481), .A2(n322), .A3(n670), .Y(n671) );
  INVX1_HVT U27 ( .A(n726), .Y(n540) );
  MUX21X1_HVT U28 ( .A1(n721), .A2(n503), .S0(n449), .Y(n609) );
  MUX21X1_HVT U29 ( .A1(n416), .A2(n517), .S0(n450), .Y(n619) );
  NOR2X0_HVT U30 ( .A1(n404), .A2(n117), .Y(n403) );
  INVX1_HVT U31 ( .A(n493), .Y(n492) );
  INVX1_HVT U32 ( .A(n403), .Y(n715) );
  INVX1_HVT U33 ( .A(n489), .Y(n395) );
  INVX1_HVT U34 ( .A(n428), .Y(n333) );
  INVX1_HVT U35 ( .A(n238), .Y(n491) );
  XNOR2X1_HVT U36 ( .A1(n450), .A2(n218), .Y(n462) );
  INVX1_HVT U37 ( .A(n483), .Y(n485) );
  INVX1_HVT U38 ( .A(in[2]), .Y(n489) );
  AO21X1_HVT U39 ( .A1(n119), .A2(n413), .A3(n450), .Y(n648) );
  MUX21X1_HVT U40 ( .A1(n584), .A2(n583), .S0(n469), .Y(n582) );
  INVX1_HVT U41 ( .A(n709), .Y(n539) );
  INVX1_HVT U43 ( .A(n314), .Y(n447) );
  INVX1_HVT U44 ( .A(n488), .Y(n222) );
  MUX21X1_HVT U45 ( .A1(n498), .A2(n417), .S0(n394), .Y(n730) );
  INVX1_HVT U46 ( .A(n678), .Y(n536) );
  MUX21X1_HVT U47 ( .A1(n414), .A2(n729), .S0(n278), .Y(n672) );
  INVX1_HVT U48 ( .A(n379), .Y(n283) );
  INVX1_HVT U49 ( .A(n428), .Y(n314) );
  OA21X1_HVT U50 ( .A1(n497), .A2(n450), .A3(n719), .Y(n608) );
  MUX21X1_HVT U52 ( .A1(n745), .A2(n615), .S0(n283), .Y(n614) );
  INVX1_HVT U54 ( .A(n238), .Y(n240) );
  INVX1_HVT U55 ( .A(n710), .Y(n501) );
  INVX1_HVT U57 ( .A(n469), .Y(n430) );
  MUX21X1_HVT U59 ( .A1(n571), .A2(n572), .S0(n314), .Y(n570) );
  INVX1_HVT U60 ( .A(n380), .Y(n441) );
  MUX21X1_HVT U62 ( .A1(n457), .A2(n506), .S0(n380), .Y(n622) );
  NAND2X0_HVT U63 ( .A1(n388), .A2(n389), .Y(n464) );
  MUX21X1_HVT U64 ( .A1(n370), .A2(n498), .S0(n399), .Y(n580) );
  INVX0_HVT U65 ( .A(n493), .Y(n490) );
  INVX1_HVT U67 ( .A(n213), .Y(n347) );
  INVX0_HVT U69 ( .A(n238), .Y(n437) );
  INVX1_HVT U70 ( .A(n471), .Y(n213) );
  INVX1_HVT U71 ( .A(n472), .Y(n278) );
  INVX1_HVT U72 ( .A(n424), .Y(n238) );
  INVX1_HVT U75 ( .A(n471), .Y(n261) );
  INVX0_HVT U76 ( .A(n393), .Y(n119) );
  INVX0_HVT U77 ( .A(n394), .Y(n438) );
  INVX1_HVT U78 ( .A(n485), .Y(n406) );
  INVX0_HVT U79 ( .A(n483), .Y(n448) );
  INVX0_HVT U80 ( .A(n438), .Y(n218) );
  INVX0_HVT U81 ( .A(n485), .Y(n425) );
  INVX1_HVT U82 ( .A(n470), .Y(n354) );
  AND2X1_HVT U86 ( .A1(n339), .A2(n340), .Y(n65) );
  INVX0_HVT U87 ( .A(n408), .Y(n212) );
  INVX1_HVT U88 ( .A(n401), .Y(n113) );
  INVX1_HVT U89 ( .A(n113), .Y(n114) );
  MUX21X1_HVT U90 ( .A1(n479), .A2(n224), .S0(n246), .Y(n632) );
  INVX0_HVT U91 ( .A(n744), .Y(n518) );
  INVX0_HVT U92 ( .A(n744), .Y(n373) );
  MUX41X1_HVT U93 ( .A1(n607), .A3(n611), .A2(n606), .A4(n610), .S0(n475), 
        .S1(n261), .Y(n605) );
  INVX0_HVT U94 ( .A(n422), .Y(n407) );
  INVX1_HVT U95 ( .A(n485), .Y(n256) );
  INVX0_HVT U96 ( .A(n720), .Y(n527) );
  INVX1_HVT U97 ( .A(n518), .Y(n371) );
  MUX41X1_HVT U98 ( .A1(n730), .A3(n510), .A2(n739), .A4(n695), .S0(n429), 
        .S1(n470), .Y(n693) );
  INVX1_HVT U99 ( .A(n307), .Y(n564) );
  MUX41X1_HVT U100 ( .A1(n38), .A3(n312), .A2(n336), .A4(n748), .S0(n430), 
        .S1(n490), .Y(n561) );
  MUX41X1_HVT U102 ( .A1(n740), .A3(n504), .A2(n455), .A4(n737), .S0(n433), 
        .S1(n395), .Y(n575) );
  MUX21X1_HVT U104 ( .A1(n375), .A2(n417), .S0(n482), .Y(n740) );
  INVX0_HVT U105 ( .A(n740), .Y(n523) );
  INVX0_HVT U106 ( .A(n454), .Y(n365) );
  INVX0_HVT U107 ( .A(n489), .Y(n488) );
  NBUFFX2_HVT U108 ( .A(n483), .Y(n117) );
  XOR2X1_HVT U109 ( .A1(n478), .A2(n484), .Y(n724) );
  OA21X1_HVT U111 ( .A1(n461), .A2(n450), .A3(n719), .Y(n583) );
  INVX0_HVT U112 ( .A(n416), .Y(n118) );
  INVX0_HVT U113 ( .A(n411), .Y(n412) );
  INVX1_HVT U114 ( .A(n10), .Y(n416) );
  INVX1_HVT U116 ( .A(n444), .Y(n336) );
  INVX1_HVT U117 ( .A(n479), .Y(n408) );
  INVX1_HVT U118 ( .A(n381), .Y(n376) );
  INVX1_HVT U119 ( .A(n422), .Y(n484) );
  NAND2X0_HVT U120 ( .A1(n736), .A2(n245), .Y(n737) );
  INVX1_HVT U121 ( .A(n225), .Y(n245) );
  INVX0_HVT U122 ( .A(n345), .Y(n688) );
  MUX21X1_HVT U124 ( .A1(n411), .A2(n38), .S0(n474), .Y(n584) );
  INVX1_HVT U126 ( .A(n10), .Y(n411) );
  NBUFFX2_HVT U127 ( .A(n525), .Y(n477) );
  MUX41X1_HVT U128 ( .A1(n562), .A3(n558), .A2(n563), .A4(n561), .S0(n313), 
        .S1(n470), .Y(n557) );
  MUX21X2_HVT U129 ( .A1(n480), .A2(n476), .S0(n406), .Y(n710) );
  MUX21X1_HVT U130 ( .A1(n413), .A2(n370), .S0(n482), .Y(n731) );
  XOR2X1_HVT U131 ( .A1(n480), .A2(n482), .Y(n702) );
  MUX21X1_HVT U132 ( .A1(n409), .A2(n454), .S0(n482), .Y(n644) );
  MUX21X1_HVT U133 ( .A1(n375), .A2(n411), .S0(n482), .Y(n662) );
  MUX21X2_HVT U134 ( .A1(n631), .A2(n630), .S0(n474), .Y(n627) );
  MUX41X1_HVT U135 ( .A1(n705), .A3(n712), .A2(n678), .A4(n458), .S0(n278), 
        .S1(n430), .Y(n569) );
  MUX41X1_HVT U137 ( .A1(n719), .A3(n495), .A2(n638), .A4(n737), .S0(n430), 
        .S1(n433), .Y(n637) );
  INVX1_HVT U138 ( .A(n117), .Y(n486) );
  OR2X1_HVT U139 ( .A1(n448), .A2(n454), .Y(n736) );
  INVX1_HVT U143 ( .A(n742), .Y(n364) );
  NAND2X0_HVT U144 ( .A1(n382), .A2(n119), .Y(n210) );
  NAND2X0_HVT U145 ( .A1(n364), .A2(n393), .Y(n211) );
  NAND2X0_HVT U147 ( .A1(n210), .A2(n211), .Y(n592) );
  MUX21X2_HVT U148 ( .A1(n528), .A2(n720), .S0(n468), .Y(n624) );
  MUX21X1_HVT U149 ( .A1(n225), .A2(n370), .S0(n407), .Y(n713) );
  MUX21X2_HVT U150 ( .A1(n514), .A2(n632), .S0(n379), .Y(n631) );
  MUX21X1_HVT U151 ( .A1(n371), .A2(n479), .S0(n394), .Y(n305) );
  INVX1_HVT U152 ( .A(n478), .Y(n436) );
  MUX41X1_HVT U153 ( .A1(n622), .A3(n621), .A2(n624), .A4(n623), .S0(n433), 
        .S1(n402), .Y(n620) );
  INVX0_HVT U155 ( .A(n311), .Y(n368) );
  MUX41X1_HVT U156 ( .A1(n552), .A3(n551), .A2(n554), .A4(n553), .S0(n261), 
        .S1(n475), .Y(n550) );
  INVX1_HVT U157 ( .A(in[1]), .Y(n423) );
  NAND2X0_HVT U160 ( .A1(n732), .A2(n222), .Y(n216) );
  NAND2X0_HVT U161 ( .A1(n305), .A2(n379), .Y(n217) );
  NAND2X0_HVT U163 ( .A1(n216), .A2(n217), .Y(n621) );
  INVX0_HVT U164 ( .A(n466), .Y(n639) );
  OA21X1_HVT U165 ( .A1(n716), .A2(n450), .A3(n507), .Y(n571) );
  INVX1_HVT U169 ( .A(n544), .Y(n517) );
  INVX1_HVT U170 ( .A(n485), .Y(n405) );
  XNOR2X2_HVT U171 ( .A1(n477), .A2(n229), .Y(n219) );
  INVX0_HVT U173 ( .A(n719), .Y(n533) );
  MUX41X1_HVT U174 ( .A1(n746), .A3(n408), .A2(n533), .A4(n526), .S0(n222), 
        .S1(n491), .Y(n551) );
  INVX0_HVT U175 ( .A(n423), .Y(n394) );
  MUX41X1_HVT U179 ( .A1(n502), .A3(n735), .A2(n706), .A4(n540), .S0(n437), 
        .S1(n283), .Y(n668) );
  NBUFFX2_HVT U180 ( .A(n492), .Y(n449) );
  NBUFFX2_HVT U181 ( .A(n492), .Y(n472) );
  INVX1_HVT U183 ( .A(n373), .Y(n375) );
  OR2X1_HVT U184 ( .A1(n224), .A2(n218), .Y(n726) );
  NBUFFX2_HVT U185 ( .A(n492), .Y(n474) );
  INVX0_HVT U186 ( .A(n371), .Y(n372) );
  AND2X1_HVT U187 ( .A1(n114), .A2(n376), .Y(n225) );
  INVX1_HVT U188 ( .A(n538), .Y(n229) );
  INVX1_HVT U190 ( .A(in[3]), .Y(n538) );
  MUX41X1_HVT U191 ( .A1(n661), .A3(n656), .A2(n654), .A4(n653), .S0(n354), 
        .S1(n313), .Y(n652) );
  MUX41X1_HVT U192 ( .A1(n641), .A3(n459), .A2(n481), .A4(n403), .S0(n380), 
        .S1(n240), .Y(n600) );
  MUX41X1_HVT U193 ( .A1(n596), .A3(n601), .A2(n594), .A4(n600), .S0(n475), 
        .S1(n354), .Y(n593) );
  NAND2X0_HVT U195 ( .A1(n599), .A2(n231), .Y(n232) );
  NAND2X0_HVT U196 ( .A1(n481), .A2(n462), .Y(n236) );
  NAND2X0_HVT U198 ( .A1(n232), .A2(n236), .Y(n598) );
  INVX0_HVT U199 ( .A(n462), .Y(n231) );
  INVX0_HVT U200 ( .A(n489), .Y(n487) );
  MUX21X1_HVT U201 ( .A1(n479), .A2(n113), .S0(n428), .Y(n344) );
  MUX21X2_HVT U202 ( .A1(n480), .A2(n416), .S0(n407), .Y(n735) );
  NBUFFX2_HVT U204 ( .A(n219), .Y(n476) );
  INVX0_HVT U205 ( .A(n725), .Y(n495) );
  INVX0_HVT U206 ( .A(n493), .Y(n424) );
  INVX1_HVT U207 ( .A(n448), .Y(n246) );
  NAND2X0_HVT U209 ( .A1(n224), .A2(n246), .Y(n252) );
  NAND2X0_HVT U210 ( .A1(n219), .A2(n448), .Y(n253) );
  NAND2X0_HVT U211 ( .A1(n252), .A2(n253), .Y(n733) );
  MUX21X1_HVT U213 ( .A1(n455), .A2(n733), .S0(n433), .Y(n556) );
  INVX1_HVT U216 ( .A(n722), .Y(n528) );
  INVX0_HVT U217 ( .A(in[1]), .Y(n422) );
  INVX0_HVT U219 ( .A(n365), .Y(n259) );
  INVX0_HVT U221 ( .A(n305), .Y(n718) );
  MUX41X1_HVT U222 ( .A1(n579), .A3(n576), .A2(n577), .A4(n575), .S0(n313), 
        .S1(n261), .Y(n574) );
  INVX1_HVT U223 ( .A(in[0]), .Y(n313) );
  MUX21X1_HVT U224 ( .A1(n212), .A2(n364), .S0(n438), .Y(n647) );
  NAND2X0_HVT U225 ( .A1(n603), .A2(n447), .Y(n264) );
  NAND2X0_HVT U226 ( .A1(n604), .A2(n325), .Y(n271) );
  NAND2X0_HVT U227 ( .A1(n264), .A2(n271), .Y(n601) );
  NAND2X0_HVT U228 ( .A1(n400), .A2(n119), .Y(n274) );
  NAND2X0_HVT U229 ( .A1(n476), .A2(n406), .Y(n275) );
  NAND2X0_HVT U230 ( .A1(n274), .A2(n275), .Y(n323) );
  OA21X1_HVT U231 ( .A1(n450), .A2(n711), .A3(n602), .Y(n603) );
  MUX21X1_HVT U232 ( .A1(n323), .A2(n412), .S0(n474), .Y(n604) );
  INVX0_HVT U233 ( .A(n390), .Y(n400) );
  OR2X1_HVT U234 ( .A1(n369), .A2(n425), .Y(n717) );
  INVX1_HVT U235 ( .A(n369), .Y(n370) );
  INVX1_HVT U236 ( .A(n423), .Y(n399) );
  MUX41X1_HVT U237 ( .A1(n643), .A3(n645), .A2(n646), .A4(n650), .S0(n470), 
        .S1(n475), .Y(n642) );
  NAND2X0_HVT U238 ( .A1(n727), .A2(n278), .Y(n280) );
  NAND2X0_HVT U239 ( .A1(n516), .A2(n472), .Y(n282) );
  NAND2X0_HVT U240 ( .A1(n280), .A2(n282), .Y(n615) );
  INVX0_HVT U241 ( .A(n712), .Y(n516) );
  NBUFFX2_HVT U242 ( .A(n401), .Y(n417) );
  NAND2X0_HVT U243 ( .A1(n348), .A2(n349), .Y(n681) );
  XOR2X2_HVT U244 ( .A1(n406), .A2(n742), .Y(n705) );
  MUX41X1_HVT U246 ( .A1(n519), .A3(n740), .A2(n323), .A4(n675), .S0(n429), 
        .S1(n488), .Y(n674) );
  INVX0_HVT U247 ( .A(n422), .Y(n393) );
  NAND2X0_HVT U248 ( .A1(n401), .A2(n478), .Y(n288) );
  INVX0_HVT U249 ( .A(n657), .Y(n519) );
  NAND2X0_HVT U250 ( .A1(n581), .A2(n451), .Y(n352) );
  INVX1_HVT U251 ( .A(n213), .Y(n402) );
  MUX41X1_HVT U252 ( .A1(n705), .A3(n500), .A2(n709), .A4(n662), .S0(n240), 
        .S1(n488), .Y(n661) );
  MUX41X1_HVT U253 ( .A1(n531), .A3(n532), .A2(n495), .A4(n308), .S0(n441), 
        .S1(n240), .Y(n676) );
  NAND2X0_HVT U254 ( .A1(n539), .A2(n278), .Y(n290) );
  NAND2X0_HVT U257 ( .A1(n324), .A2(n472), .Y(n293) );
  NAND2X0_HVT U258 ( .A1(n290), .A2(n293), .Y(n560) );
  NAND2X0_HVT U259 ( .A1(n559), .A2(n333), .Y(n297) );
  NAND2X0_HVT U260 ( .A1(n560), .A2(n441), .Y(n302) );
  NAND2X0_HVT U261 ( .A1(n297), .A2(n302), .Y(n558) );
  MUX41X1_HVT U263 ( .A1(n618), .A3(n616), .A2(n617), .A4(n614), .S0(n313), 
        .S1(n261), .Y(n613) );
  NAND2X0_HVT U264 ( .A1(n365), .A2(n119), .Y(n303) );
  NAND2X0_HVT U266 ( .A1(n212), .A2(n406), .Y(n304) );
  NAND2X0_HVT U267 ( .A1(n303), .A2(n304), .Y(n675) );
  INVX1_HVT U269 ( .A(n398), .Y(n723) );
  MUX41X1_HVT U272 ( .A1(n690), .A3(n683), .A2(n696), .A4(n687), .S0(n451), 
        .S1(n475), .Y(out[0]) );
  INVX1_HVT U273 ( .A(n503), .Y(n306) );
  MUX21X1_HVT U274 ( .A1(n400), .A2(n404), .S0(n256), .Y(n307) );
  INVX1_HVT U275 ( .A(n317), .Y(n324) );
  INVX1_HVT U276 ( .A(n412), .Y(n414) );
  INVX1_HVT U277 ( .A(n410), .Y(n415) );
  INVX0_HVT U279 ( .A(n411), .Y(n413) );
  INVX0_HVT U281 ( .A(n288), .Y(n308) );
  INVX0_HVT U282 ( .A(n288), .Y(n498) );
  MUX21X1_HVT U283 ( .A1(n436), .A2(n118), .S0(n399), .Y(n732) );
  INVX1_HVT U285 ( .A(n547), .Y(n500) );
  NAND2X0_HVT U286 ( .A1(n117), .A2(n288), .Y(n746) );
  NAND2X0_HVT U287 ( .A1(n245), .A2(n256), .Y(n309) );
  NAND2X0_HVT U288 ( .A1(n225), .A2(n350), .Y(n310) );
  NAND2X0_HVT U290 ( .A1(n309), .A2(n310), .Y(n460) );
  NAND2X0_HVT U291 ( .A1(n376), .A2(n401), .Y(n311) );
  INVX1_HVT U292 ( .A(n538), .Y(n401) );
  NBUFFX2_HVT U296 ( .A(n365), .Y(n312) );
  NBUFFX2_HVT U298 ( .A(n525), .Y(n478) );
  NAND2X0_HVT U299 ( .A1(n659), .A2(n314), .Y(n315) );
  NAND2X0_HVT U300 ( .A1(n658), .A2(n447), .Y(n316) );
  NAND2X0_HVT U301 ( .A1(n315), .A2(n316), .Y(n656) );
  MUX21X1_HVT U302 ( .A1(n408), .A2(n411), .S0(n484), .Y(n317) );
  NBUFFX2_HVT U304 ( .A(n538), .Y(n318) );
  NAND2X0_HVT U305 ( .A1(n598), .A2(n314), .Y(n319) );
  NAND2X0_HVT U307 ( .A1(n597), .A2(n447), .Y(n320) );
  NAND2X0_HVT U308 ( .A1(n319), .A2(n320), .Y(n596) );
  INVX1_HVT U310 ( .A(n451), .Y(n321) );
  INVX1_HVT U311 ( .A(in[6]), .Y(n451) );
  INVX1_HVT U312 ( .A(n532), .Y(n322) );
  INVX1_HVT U313 ( .A(n694), .Y(n532) );
  INVX1_HVT U314 ( .A(n732), .Y(n529) );
  NAND2X0_HVT U315 ( .A1(n671), .A2(n325), .Y(n326) );
  NAND2X0_HVT U316 ( .A1(n672), .A2(n430), .Y(n327) );
  NAND2X0_HVT U317 ( .A1(n326), .A2(n327), .Y(n669) );
  INVX0_HVT U318 ( .A(n283), .Y(n325) );
  NAND2X0_HVT U319 ( .A1(n498), .A2(n218), .Y(n328) );
  NAND2X0_HVT U320 ( .A1(n365), .A2(n438), .Y(n329) );
  NAND2X0_HVT U321 ( .A1(n329), .A2(n328), .Y(n725) );
  MUX21X1_HVT U322 ( .A1(n311), .A2(n410), .S0(n405), .Y(n719) );
  INVX1_HVT U323 ( .A(n423), .Y(n483) );
  INVX0_HVT U324 ( .A(n407), .Y(n350) );
  NAND2X0_HVT U325 ( .A1(n459), .A2(n330), .Y(n331) );
  NAND2X0_HVT U326 ( .A1(n651), .A2(n704), .Y(n332) );
  NAND2X0_HVT U327 ( .A1(n331), .A2(n332), .Y(n650) );
  INVX0_HVT U328 ( .A(n704), .Y(n330) );
  NAND2X0_HVT U329 ( .A1(n359), .A2(n333), .Y(n334) );
  NAND2X0_HVT U330 ( .A1(n533), .A2(n428), .Y(n335) );
  NAND2X0_HVT U331 ( .A1(n334), .A2(n335), .Y(n358) );
  INVX1_HVT U332 ( .A(n468), .Y(n428) );
  INVX0_HVT U333 ( .A(n373), .Y(n369) );
  MUX21X1_HVT U334 ( .A1(n374), .A2(n748), .S0(n117), .Y(n657) );
  AO21X1_HVT U335 ( .A1(n336), .A2(n380), .A3(n731), .Y(n467) );
  NAND2X0_HVT U336 ( .A1(n649), .A2(n222), .Y(n337) );
  NAND2X0_HVT U337 ( .A1(n65), .A2(n469), .Y(n338) );
  NAND2X0_HVT U338 ( .A1(n337), .A2(n338), .Y(n646) );
  NAND2X0_HVT U339 ( .A1(n720), .A2(n433), .Y(n339) );
  NAND2X0_HVT U340 ( .A1(n548), .A2(n473), .Y(n340) );
  NBUFFX2_HVT U341 ( .A(n492), .Y(n473) );
  NBUFFX2_HVT U342 ( .A(n748), .Y(n341) );
  NAND2X0_HVT U343 ( .A1(n635), .A2(n238), .Y(n342) );
  NAND2X0_HVT U344 ( .A1(n636), .A2(n473), .Y(n343) );
  NAND2X0_HVT U345 ( .A1(n342), .A2(n343), .Y(n634) );
  MUX41X1_HVT U346 ( .A1(n218), .A3(n532), .A2(n734), .A4(n458), .S0(n429), 
        .S1(n395), .Y(n653) );
  INVX1_HVT U347 ( .A(n716), .Y(n535) );
  MUX41X1_HVT U348 ( .A1(n464), .A3(n358), .A2(n50), .A4(n467), .S0(n473), 
        .S1(n471), .Y(n466) );
  NAND2X0_HVT U349 ( .A1(n699), .A2(n493), .Y(n360) );
  INVX0_HVT U350 ( .A(n641), .Y(n359) );
  MUX41X1_HVT U351 ( .A1(n734), .A3(n23), .A2(n735), .A4(n737), .S0(n429), 
        .S1(n347), .Y(n345) );
  NBUFFX2_HVT U352 ( .A(n538), .Y(n390) );
  INVX1_HVT U353 ( .A(n357), .Y(n686) );
  NBUFFX2_HVT U354 ( .A(n382), .Y(n346) );
  MUX21X1_HVT U355 ( .A1(n390), .A2(n382), .S0(n422), .Y(n716) );
  MUX41X1_HVT U356 ( .A1(n665), .A3(n531), .A2(n456), .A4(n460), .S0(n430), 
        .S1(n490), .Y(n664) );
  MUX21X1_HVT U357 ( .A1(n390), .A2(n374), .S0(n422), .Y(n738) );
  MUX41X1_HVT U358 ( .A1(n528), .A3(n644), .A2(n703), .A4(n521), .S0(n473), 
        .S1(n379), .Y(n643) );
  NAND2X0_HVT U359 ( .A1(n392), .A2(n391), .Y(out[6]) );
  MUX41X1_HVT U360 ( .A1(n674), .A3(n677), .A2(n676), .A4(n681), .S0(n475), 
        .S1(n347), .Y(n673) );
  NAND2X0_HVT U361 ( .A1(n682), .A2(n333), .Y(n348) );
  NAND2X0_HVT U362 ( .A1(n707), .A2(n441), .Y(n349) );
  NAND2X0_HVT U363 ( .A1(n409), .A2(n350), .Y(n351) );
  MUX21X1_HVT U364 ( .A1(n346), .A2(n38), .S0(n472), .Y(n682) );
  INVX0_HVT U365 ( .A(n729), .Y(n502) );
  MUX21X1_HVT U366 ( .A1(n436), .A2(n480), .S0(n407), .Y(n729) );
  XNOR2X1_HVT U367 ( .A1(n350), .A2(n417), .Y(n703) );
  MUX41X1_HVT U368 ( .A1(n668), .A3(n664), .A2(n669), .A4(n666), .S0(n313), 
        .S1(n470), .Y(n663) );
  NAND2X0_HVT U369 ( .A1(n593), .A2(n321), .Y(n353) );
  NAND2X0_HVT U370 ( .A1(n352), .A2(n353), .Y(out[5]) );
  NAND2X0_HVT U371 ( .A1(n354), .A2(n523), .Y(n355) );
  NAND2X0_HVT U372 ( .A1(n412), .A2(n470), .Y(n356) );
  NAND2X0_HVT U373 ( .A1(n355), .A2(n356), .Y(n684) );
  MUX21X1_HVT U374 ( .A1(n218), .A2(n738), .S0(n213), .Y(n357) );
  MUX21X1_HVT U375 ( .A1(n519), .A2(n713), .S0(n278), .Y(n597) );
  MUX41X1_HVT U376 ( .A1(n458), .A3(n540), .A2(n655), .A4(n38), .S0(n283), 
        .S1(n437), .Y(n654) );
  NAND2X0_HVT U377 ( .A1(n700), .A2(n449), .Y(n361) );
  NAND2X0_HVT U378 ( .A1(n361), .A2(n360), .Y(n697) );
  INVX1_HVT U379 ( .A(in[4]), .Y(n525) );
  NAND2X0_HVT U380 ( .A1(n454), .A2(n350), .Y(n362) );
  NAND2X0_HVT U381 ( .A1(n417), .A2(n407), .Y(n363) );
  NAND2X0_HVT U382 ( .A1(n362), .A2(n363), .Y(n727) );
  INVX0_HVT U383 ( .A(n727), .Y(n507) );
  NAND2X0_HVT U384 ( .A1(n533), .A2(n222), .Y(n366) );
  NAND2X0_HVT U385 ( .A1(n488), .A2(n735), .Y(n367) );
  NAND2X0_HVT U386 ( .A1(n366), .A2(n367), .Y(n651) );
  MUX41X1_HVT U387 ( .A1(n509), .A3(n743), .A2(n413), .A4(n723), .S0(n491), 
        .S1(n380), .Y(n617) );
  INVX0_HVT U388 ( .A(n739), .Y(n534) );
  MUX41X1_HVT U389 ( .A1(n705), .A3(n589), .A2(n728), .A4(n527), .S0(n437), 
        .S1(n283), .Y(n588) );
  INVX1_HVT U390 ( .A(n373), .Y(n374) );
  NAND2X0_HVT U391 ( .A1(n689), .A2(n325), .Y(n377) );
  NAND2X0_HVT U392 ( .A1(n688), .A2(n441), .Y(n378) );
  NAND2X0_HVT U393 ( .A1(n377), .A2(n378), .Y(n687) );
  MUX41X1_HVT U394 ( .A1(n591), .A3(n529), .A2(n592), .A4(n457), .S0(n441), 
        .S1(n491), .Y(n590) );
  NBUFFX2_HVT U395 ( .A(n487), .Y(n379) );
  NBUFFX2_HVT U396 ( .A(n487), .Y(n380) );
  NBUFFX2_HVT U397 ( .A(n487), .Y(n468) );
  NAND2X0_HVT U398 ( .A1(n701), .A2(n395), .Y(n383) );
  NAND2X0_HVT U399 ( .A1(n697), .A2(n283), .Y(n384) );
  NAND2X0_HVT U400 ( .A1(n384), .A2(n383), .Y(n696) );
  NAND2X0_HVT U401 ( .A1(n691), .A2(n441), .Y(n385) );
  NAND2X0_HVT U402 ( .A1(n693), .A2(n325), .Y(n386) );
  NAND2X0_HVT U403 ( .A1(n386), .A2(n385), .Y(n690) );
  NAND2X0_HVT U404 ( .A1(n308), .A2(n387), .Y(n388) );
  NAND2X0_HVT U405 ( .A1(n344), .A2(n465), .Y(n389) );
  INVX0_HVT U406 ( .A(n465), .Y(n387) );
  INVX0_HVT U407 ( .A(n713), .Y(n515) );
  MUX21X1_HVT U408 ( .A1(n417), .A2(n715), .S0(n402), .Y(n700) );
  MUX41X1_HVT U409 ( .A1(n512), .A3(n461), .A2(n692), .A4(n463), .S0(n493), 
        .S1(n261), .Y(n691) );
  NAND2X0_HVT U410 ( .A1(n574), .A2(n321), .Y(n391) );
  NAND2X0_HVT U411 ( .A1(n565), .A2(n451), .Y(n392) );
  OA21X1_HVT U412 ( .A1(n741), .A2(n450), .A3(n515), .Y(n555) );
  INVX1_HVT U413 ( .A(n543), .Y(n509) );
  NAND2X0_HVT U414 ( .A1(n450), .A2(n398), .Y(n396) );
  NAND2X0_HVT U415 ( .A1(n473), .A2(n723), .Y(n397) );
  NAND2X0_HVT U416 ( .A1(n396), .A2(n397), .Y(n707) );
  MUX21X1_HVT U417 ( .A1(n288), .A2(n245), .S0(n393), .Y(n398) );
  NBUFFX2_HVT U418 ( .A(n238), .Y(n450) );
  INVX0_HVT U419 ( .A(n381), .Y(n404) );
  MUX41X1_HVT U420 ( .A1(n566), .A3(n569), .A2(n570), .A4(n573), .S0(n402), 
        .S1(n475), .Y(n565) );
  INVX0_HVT U421 ( .A(n711), .Y(n496) );
  NAND2X0_HVT U422 ( .A1(n436), .A2(n390), .Y(n409) );
  NAND2X0_HVT U423 ( .A1(n436), .A2(n390), .Y(n410) );
  INVX1_HVT U424 ( .A(n731), .Y(n512) );
  NAND2X0_HVT U425 ( .A1(n608), .A2(n325), .Y(n418) );
  NAND2X0_HVT U426 ( .A1(n609), .A2(n222), .Y(n419) );
  NAND2X0_HVT U427 ( .A1(n418), .A2(n419), .Y(n607) );
  INVX1_HVT U428 ( .A(n546), .Y(n510) );
  NAND2X0_HVT U429 ( .A1(n550), .A2(n451), .Y(n420) );
  NAND2X0_HVT U430 ( .A1(n557), .A2(n321), .Y(n421) );
  NAND2X0_HVT U431 ( .A1(n421), .A2(n420), .Y(out[7]) );
  MUX41X1_HVT U432 ( .A1(n625), .A3(n639), .A2(n620), .A4(n633), .S0(n321), 
        .S1(n313), .Y(out[3]) );
  MUX21X1_HVT U433 ( .A1(n113), .A2(n368), .S0(n425), .Y(n739) );
  AO21X1_HVT U434 ( .A1(n657), .A2(n473), .A3(n530), .Y(n658) );
  MUX41X1_HVT U435 ( .A1(n324), .A3(n511), .A2(n526), .A4(n722), .S0(n428), 
        .S1(n278), .Y(n576) );
  NAND2X0_HVT U436 ( .A1(n446), .A2(n445), .Y(out[2]) );
  NAND2X0_HVT U437 ( .A1(n626), .A2(n354), .Y(n426) );
  NAND2X0_HVT U438 ( .A1(n627), .A2(n402), .Y(n427) );
  NAND2X0_HVT U439 ( .A1(n427), .A2(n426), .Y(n625) );
  MUX41X1_HVT U440 ( .A1(n737), .A3(n695), .A2(n727), .A4(n535), .S0(n447), 
        .S1(n491), .Y(n552) );
  NAND2X0_HVT U441 ( .A1(n555), .A2(n428), .Y(n431) );
  NAND2X0_HVT U442 ( .A1(n556), .A2(n469), .Y(n432) );
  NAND2X0_HVT U443 ( .A1(n431), .A2(n432), .Y(n554) );
  MUX21X1_HVT U444 ( .A1(n476), .A2(n382), .S0(n394), .Y(n741) );
  NAND2X0_HVT U445 ( .A1(n440), .A2(n439), .Y(out[1]) );
  NAND2X0_HVT U446 ( .A1(n634), .A2(n354), .Y(n434) );
  NAND2X0_HVT U447 ( .A1(n637), .A2(n402), .Y(n435) );
  NAND2X0_HVT U448 ( .A1(n435), .A2(n434), .Y(n633) );
  MUX41X1_HVT U449 ( .A1(n678), .A3(n499), .A2(n705), .A4(n532), .S0(n441), 
        .S1(n474), .Y(n606) );
  NAND2X0_HVT U450 ( .A1(n663), .A2(n451), .Y(n439) );
  NAND2X0_HVT U451 ( .A1(n673), .A2(n321), .Y(n440) );
  NAND2X0_HVT U452 ( .A1(n453), .A2(n452), .Y(out[4]) );
  MUX41X1_HVT U453 ( .A1(n564), .A3(n702), .A2(n715), .A4(n709), .S0(n441), 
        .S1(n429), .Y(n563) );
  NAND2X0_HVT U454 ( .A1(n481), .A2(n231), .Y(n442) );
  NAND2X0_HVT U455 ( .A1(n660), .A2(n462), .Y(n443) );
  NAND2X0_HVT U456 ( .A1(n442), .A2(n443), .Y(n659) );
  MUX21X1_HVT U457 ( .A1(n417), .A2(n212), .S0(n472), .Y(n660) );
  MUX21X1_HVT U458 ( .A1(n370), .A2(n454), .S0(n484), .Y(n444) );
  NAND2X0_HVT U459 ( .A1(n642), .A2(n451), .Y(n445) );
  NAND2X0_HVT U460 ( .A1(n652), .A2(n321), .Y(n446) );
  NBUFFX2_HVT U461 ( .A(n525), .Y(n479) );
  NAND2X0_HVT U462 ( .A1(n605), .A2(n451), .Y(n452) );
  NAND2X0_HVT U463 ( .A1(n613), .A2(n321), .Y(n453) );
  XNOR2X2_HVT U464 ( .A1(n477), .A2(n229), .Y(n454) );
  AND2X1_HVT U465 ( .A1(n364), .A2(n694), .Y(n455) );
  MUX21X1_HVT U466 ( .A1(n372), .A2(n346), .S0(n402), .Y(n698) );
  AND2X1_HVT U467 ( .A1(n481), .A2(n678), .Y(n456) );
  MUX21X1_HVT U468 ( .A1(n365), .A2(n118), .S0(n399), .Y(n543) );
  MUX21X1_HVT U469 ( .A1(n479), .A2(n372), .S0(n256), .Y(n721) );
  NAND2X0_HVT U470 ( .A1(n381), .A2(n318), .Y(n744) );
  MUX21X1_HVT U471 ( .A1(n372), .A2(n478), .S0(n425), .Y(n544) );
  MUX21X1_HVT U472 ( .A1(n113), .A2(n498), .S0(n246), .Y(n711) );
  NBUFFX2_HVT U473 ( .A(n747), .Y(n480) );
  MUX21X1_HVT U474 ( .A1(n480), .A2(n374), .S0(n246), .Y(n542) );
  MUX21X1_HVT U475 ( .A1(n224), .A2(n341), .S0(n406), .Y(n567) );
  MUX21X1_HVT U476 ( .A1(n245), .A2(n481), .S0(n405), .Y(n568) );
  XOR2X1_HVT U477 ( .A1(n484), .A2(n415), .Y(n706) );
  NBUFFX2_HVT U478 ( .A(n747), .Y(n481) );
  MUX21X1_HVT U479 ( .A1(n480), .A2(n212), .S0(n256), .Y(n547) );
  AND2X1_HVT U480 ( .A1(n394), .A2(n308), .Y(n458) );
  AND2X1_HVT U481 ( .A1(n341), .A2(n640), .Y(n459) );
  MUX21X1_HVT U482 ( .A1(n414), .A2(n341), .S0(n469), .Y(n629) );
  NBUFFX2_HVT U483 ( .A(n487), .Y(n469) );
  NBUFFX2_HVT U484 ( .A(in[5]), .Y(n471) );
  MUX21X1_HVT U485 ( .A1(n665), .A2(n417), .S0(n474), .Y(n572) );
  MUX21X1_HVT U486 ( .A1(n417), .A2(n370), .S0(n406), .Y(n712) );
  NAND2X0_HVT U487 ( .A1(n401), .A2(n381), .Y(n747) );
  AND2X1_HVT U488 ( .A1(n259), .A2(n486), .Y(n461) );
  MUX21X1_HVT U489 ( .A1(n415), .A2(n498), .S0(n256), .Y(n589) );
  XOR2X1_HVT U490 ( .A1(n246), .A2(n471), .Y(n708) );
  MUX21X1_HVT U491 ( .A1(n306), .A2(n119), .S0(n395), .Y(n628) );
  MUX21X1_HVT U492 ( .A1(n400), .A2(n118), .S0(n399), .Y(n545) );
  AND2X1_HVT U493 ( .A1(n113), .A2(n486), .Y(n463) );
  MUX21X1_HVT U494 ( .A1(n408), .A2(n742), .S0(n393), .Y(n546) );
  NAND2X0_HVT U495 ( .A1(n114), .A2(n376), .Y(n748) );
  MUX21X1_HVT U496 ( .A1(n748), .A2(n408), .S0(n425), .Y(n722) );
  MUX21X1_HVT U497 ( .A1(n408), .A2(n748), .S0(n117), .Y(n541) );
  MUX21X1_HVT U498 ( .A1(n390), .A2(n436), .S0(n405), .Y(n720) );
  NBUFFX2_HVT U499 ( .A(in[0]), .Y(n475) );
  XOR2X1_HVT U500 ( .A1(n488), .A2(n472), .Y(n704) );
  XNOR2X1_HVT U501 ( .A1(n399), .A2(n488), .Y(n465) );
endmodule

