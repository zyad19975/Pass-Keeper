
module sbox_18 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n46, n48, n210, n211, n212, n213, n216, n217, n218, n219, n224,
         n231, n232, n236, n238, n240, n243, n252, n256, n261, n264, n271,
         n278, n280, n282, n283, n284, n290, n293, n297, n301, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716;

  NAND2X0_HVT U4 ( .A1(n424), .A2(n714), .Y(n713) );
  NAND2X0_HVT U5 ( .A1(n428), .A2(n419), .Y(n711) );
  NAND2X0_HVT U13 ( .A1(n703), .A2(n307), .Y(n704) );
  NAND2X0_HVT U15 ( .A1(n714), .A2(n353), .Y(n701) );
  NAND2X0_HVT U21 ( .A1(n424), .A2(n212), .Y(n695) );
  NAND2X0_HVT U24 ( .A1(n414), .A2(n312), .Y(n693) );
  NAND2X0_HVT U33 ( .A1(n473), .A2(n433), .Y(n684) );
  NAND2X0_HVT U42 ( .A1(n252), .A2(n414), .Y(n675) );
  MUX41X1_HVT U51 ( .A1(n453), .A3(n477), .A2(n309), .A4(n455), .S0(n445), 
        .S1(n438), .Y(n668) );
  NAND2X0_HVT U53 ( .A1(n665), .A2(n674), .Y(n666) );
  NAND2X0_HVT U56 ( .A1(n424), .A2(n661), .Y(n662) );
  NAND2X0_HVT U58 ( .A1(n716), .A2(n271), .Y(n659) );
  MUX41X1_HVT U59 ( .A1(n402), .A3(n659), .A2(n401), .A4(n467), .S0(n445), 
        .S1(n438), .Y(n658) );
  MUX41X1_HVT U61 ( .A1(n396), .A3(n486), .A2(n460), .A4(n359), .S0(n445), 
        .S1(n438), .Y(n656) );
  NAND2X0_HVT U62 ( .A1(n212), .A2(n427), .Y(n655) );
  MUX41X1_HVT U63 ( .A1(n655), .A3(n457), .A2(n465), .A4(n331), .S0(n411), 
        .S1(n438), .Y(n654) );
  AO21X1_HVT U66 ( .A1(n492), .A2(n409), .A3(n494), .Y(n651) );
  MUX41X1_HVT U69 ( .A1(n649), .A3(n657), .A2(n653), .A4(n663), .S0(in[6]), 
        .S1(n413), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n421), .A2(n644), .Y(n645) );
  MUX41X1_HVT U75 ( .A1(n491), .A3(n488), .A2(n451), .A4(n448), .S0(n435), 
        .S1(n442), .Y(n642) );
  MUX41X1_HVT U77 ( .A1(n708), .A3(n474), .A2(n641), .A4(n340), .S0(n410), 
        .S1(n405), .Y(n640) );
  AND2X1_HVT U83 ( .A1(n430), .A2(n416), .Y(n633) );
  MUX41X1_HVT U84 ( .A1(n264), .A3(n358), .A2(n700), .A4(n633), .S0(n435), 
        .S1(n444), .Y(n632) );
  NAND2X0_HVT U85 ( .A1(n432), .A2(n304), .Y(n631) );
  MUX41X1_HVT U90 ( .A1(n672), .A3(n675), .A2(n453), .A4(n628), .S0(n406), 
        .S1(n410), .Y(n627) );
  NAND2X0_HVT U101 ( .A1(n614), .A2(n613), .Y(n615) );
  MUX41X1_HVT U103 ( .A1(n271), .A3(n479), .A2(n468), .A4(n682), .S0(n408), 
        .S1(n410), .Y(n611) );
  NAND2X0_HVT U110 ( .A1(n426), .A2(n604), .Y(n605) );
  AND2X1_HVT U115 ( .A1(n428), .A2(n359), .Y(n599) );
  AO21X1_HVT U118 ( .A1(n408), .A2(n240), .A3(n355), .Y(n596) );
  NAND2X0_HVT U123 ( .A1(n590), .A2(n589), .Y(n591) );
  MUX41X1_HVT U135 ( .A1(n462), .A3(n489), .A2(n711), .A4(n690), .S0(n408), 
        .S1(n445), .Y(n578) );
  MUX41X1_HVT U136 ( .A1(n394), .A3(n684), .A2(n452), .A4(n681), .S0(n434), 
        .S1(n445), .Y(n577) );
  AND2X1_HVT U140 ( .A1(n240), .A2(n243), .Y(n573) );
  MUX41X1_HVT U142 ( .A1(n264), .A3(n353), .A2(n475), .A4(n240), .S0(n316), 
        .S1(n444), .Y(n571) );
  MUX41X1_HVT U147 ( .A1(n452), .A3(n644), .A2(n491), .A4(n672), .S0(n435), 
        .S1(n444), .Y(n567) );
  MUX41X1_HVT U153 ( .A1(n605), .A3(n396), .A2(n283), .A4(n297), .S0(n316), 
        .S1(n445), .Y(n561) );
  AND2X1_HVT U154 ( .A1(n412), .A2(n414), .Y(n560) );
  NAND2X0_HVT U158 ( .A1(n430), .A2(n303), .Y(n556) );
  MUX41X1_HVT U159 ( .A1(n704), .A3(n359), .A2(n556), .A4(n495), .S0(n405), 
        .S1(n375), .Y(n555) );
  AND2X1_HVT U162 ( .A1(n355), .A2(n644), .Y(n552) );
  MUX41X1_HVT U163 ( .A1(n486), .A3(n552), .A2(n397), .A4(n553), .S0(n405), 
        .S1(n445), .Y(n551) );
  NAND2X0_HVT U166 ( .A1(n306), .A2(n661), .Y(n548) );
  NAND2X0_HVT U167 ( .A1(n451), .A2(n212), .Y(n547) );
  MUX41X1_HVT U168 ( .A1(n463), .A3(n240), .A2(n547), .A4(n548), .S0(n405), 
        .S1(n442), .Y(n546) );
  NAND2X0_HVT U174 ( .A1(n429), .A2(n355), .Y(n703) );
  MUX41X1_HVT U176 ( .A1(n418), .A3(n541), .A2(n461), .A4(n703), .S0(n411), 
        .S1(n404), .Y(n540) );
  NAND2X0_HVT U177 ( .A1(n430), .A2(n417), .Y(n539) );
  MUX41X1_HVT U189 ( .A1(n528), .A3(n703), .A2(n529), .A4(n476), .S0(n410), 
        .S1(n404), .Y(n527) );
  MUX41X1_HVT U194 ( .A1(n676), .A3(n690), .A2(n462), .A4(n240), .S0(n410), 
        .S1(n404), .Y(n523) );
  MUX41X1_HVT U195 ( .A1(n355), .A3(n490), .A2(n307), .A4(n680), .S0(n405), 
        .S1(n442), .Y(n522) );
  MUX21X2_HVT U196 ( .A1(n497), .A2(n483), .S0(n411), .Y(n521) );
  AO21X1_HVT U197 ( .A1(n398), .A2(n411), .A3(n487), .Y(n520) );
  MUX41X1_HVT U199 ( .A1(n519), .A3(n523), .A2(n522), .A4(n524), .S0(n413), 
        .S1(n440), .Y(n518) );
  NAND2X0_HVT U208 ( .A1(n428), .A2(n423), .Y(n604) );
  NAND2X0_HVT U212 ( .A1(n362), .A2(n421), .Y(n661) );
  NAND2X0_HVT U214 ( .A1(n358), .A2(n212), .Y(n510) );
  NAND2X0_HVT U215 ( .A1(n604), .A2(n422), .Y(n509) );
  NAND2X0_HVT U218 ( .A1(n489), .A2(n430), .Y(n563) );
  NAND2X0_HVT U220 ( .A1(n411), .A2(n510), .Y(n636) );
  INVX0_HVT U241 ( .A(n693), .Y(n498) );
  INVX0_HVT U242 ( .A(n675), .Y(n497) );
  INVX0_HVT U245 ( .A(n711), .Y(n495) );
  INVX0_HVT U247 ( .A(n644), .Y(n494) );
  INVX0_HVT U250 ( .A(n706), .Y(n492) );
  INVX0_HVT U255 ( .A(n505), .Y(n488) );
  INVX0_HVT U256 ( .A(n563), .Y(n487) );
  INVX0_HVT U259 ( .A(n687), .Y(n484) );
  INVX0_HVT U265 ( .A(n691), .Y(n480) );
  INVX0_HVT U266 ( .A(n708), .Y(n479) );
  INVX0_HVT U268 ( .A(n695), .Y(n477) );
  INVX0_HVT U270 ( .A(n509), .Y(n476) );
  INVX0_HVT U271 ( .A(n604), .Y(n475) );
  INVX0_HVT U281 ( .A(n698), .Y(n467) );
  INVX0_HVT U283 ( .A(n704), .Y(n465) );
  INVX0_HVT U284 ( .A(n510), .Y(n464) );
  INVX0_HVT U285 ( .A(n507), .Y(n463) );
  INVX0_HVT U289 ( .A(n613), .Y(n461) );
  INVX0_HVT U295 ( .A(n713), .Y(n458) );
  INVX0_HVT U297 ( .A(n714), .Y(n456) );
  INVX0_HVT U300 ( .A(n676), .Y(n454) );
  INVX0_HVT U302 ( .A(n508), .Y(n453) );
  INVX0_HVT U303 ( .A(n501), .Y(n452) );
  INVX0_HVT U306 ( .A(n547), .Y(n450) );
  INVX0_HVT U307 ( .A(n677), .Y(n449) );
  MUX21X1_HVT U1 ( .A1(n303), .A2(n238), .S0(n379), .Y(n351) );
  INVX1_HVT U2 ( .A(n415), .Y(n481) );
  MUX21X1_HVT U3 ( .A1(n573), .A2(n378), .S0(n408), .Y(n386) );
  INVX1_HVT U6 ( .A(n433), .Y(n338) );
  XNOR2X1_HVT U7 ( .A1(n404), .A2(n411), .Y(n393) );
  INVX1_HVT U8 ( .A(n380), .Y(n339) );
  INVX1_HVT U9 ( .A(in[1]), .Y(n380) );
  INVX1_HVT U10 ( .A(n432), .Y(n379) );
  MUX21X1_HVT U11 ( .A1(n533), .A2(n532), .S0(n23), .Y(n531) );
  OA21X1_HVT U12 ( .A1(n683), .A2(n261), .A3(n264), .Y(n532) );
  INVX1_HVT U14 ( .A(n403), .Y(n404) );
  INVX1_HVT U16 ( .A(n256), .Y(n442) );
  OA21X1_HVT U17 ( .A1(n677), .A2(n256), .A3(n563), .Y(n564) );
  OA21X1_HVT U18 ( .A1(n450), .A2(n256), .A3(n686), .Y(n569) );
  INVX1_HVT U19 ( .A(in[7]), .Y(n256) );
  MUX21X1_HVT U20 ( .A1(n284), .A2(n271), .S0(n408), .Y(n607) );
  AND3X1_HVT U22 ( .A1(n407), .A2(n212), .A3(n416), .Y(n584) );
  MUX21X1_HVT U23 ( .A1(n485), .A2(n687), .S0(n408), .Y(n585) );
  MUX21X1_HVT U25 ( .A1(n637), .A2(n638), .S0(n210), .Y(n635) );
  INVX1_HVT U26 ( .A(in[3]), .Y(n496) );
  INVX1_HVT U27 ( .A(in[7]), .Y(n261) );
  INVX1_HVT U28 ( .A(n406), .Y(n23) );
  MUX21X1_HVT U29 ( .A1(n351), .A2(n702), .S0(n408), .Y(n617) );
  AO21X1_HVT U30 ( .A1(n212), .A2(n489), .A3(n213), .Y(n614) );
  MUX21X1_HVT U31 ( .A1(n615), .A2(n447), .S0(n407), .Y(n612) );
  MUX21X1_HVT U32 ( .A1(n520), .A2(n521), .S0(n23), .Y(n519) );
  MUX21X1_HVT U34 ( .A1(n395), .A2(n700), .S0(n213), .Y(n517) );
  INVX1_HVT U35 ( .A(n500), .Y(n483) );
  INVX0_HVT U36 ( .A(n351), .Y(n686) );
  INVX1_HVT U37 ( .A(in[3]), .Y(n308) );
  INVX0_HVT U38 ( .A(n380), .Y(n362) );
  INVX1_HVT U39 ( .A(n380), .Y(n430) );
  MUX21X1_HVT U40 ( .A1(n496), .A2(n353), .S0(n312), .Y(n700) );
  INVX0_HVT U41 ( .A(n380), .Y(n428) );
  INVX1_HVT U43 ( .A(n380), .Y(n431) );
  INVX1_HVT U44 ( .A(n689), .Y(n485) );
  MUX21X1_HVT U45 ( .A1(n418), .A2(n473), .S0(n339), .Y(n688) );
  MUX21X1_HVT U46 ( .A1(n426), .A2(n416), .S0(n433), .Y(n696) );
  INVX1_HVT U47 ( .A(n412), .Y(n369) );
  INVX1_HVT U48 ( .A(n425), .Y(n451) );
  INVX1_HVT U49 ( .A(n684), .Y(n469) );
  INVX1_HVT U50 ( .A(n420), .Y(n489) );
  NBUFFX2_HVT U52 ( .A(n436), .Y(n408) );
  NAND2X0_HVT U54 ( .A1(n427), .A2(n352), .Y(n290) );
  MUX21X1_HVT U55 ( .A1(n473), .A2(n451), .S0(n338), .Y(n541) );
  INVX1_HVT U57 ( .A(n679), .Y(n470) );
  INVX1_HVT U60 ( .A(n356), .Y(n357) );
  MUX21X1_HVT U64 ( .A1(n427), .A2(n419), .S0(n339), .Y(n309) );
  INVX1_HVT U65 ( .A(n405), .Y(n374) );
  XOR2X1_HVT U67 ( .A1(n312), .A2(n403), .Y(n670) );
  MUX21X1_HVT U68 ( .A1(n496), .A2(n416), .S0(n431), .Y(n687) );
  INVX1_HVT U70 ( .A(n434), .Y(n403) );
  INVX1_HVT U71 ( .A(n405), .Y(n337) );
  OA21X1_HVT U72 ( .A1(n401), .A2(n261), .A3(n686), .Y(n544) );
  INVX1_HVT U74 ( .A(n282), .Y(n283) );
  MUX21X1_HVT U76 ( .A1(n558), .A2(n559), .S0(n408), .Y(n557) );
  MUX21X1_HVT U78 ( .A1(n474), .A2(n679), .S0(n213), .Y(n558) );
  MUX21X1_HVT U79 ( .A1(n456), .A2(n688), .S0(n213), .Y(n570) );
  INVX1_HVT U80 ( .A(n284), .Y(n681) );
  XOR2X1_HVT U81 ( .A1(n339), .A2(n414), .Y(n671) );
  INVX1_HVT U82 ( .A(n688), .Y(n468) );
  INVX1_HVT U86 ( .A(n435), .Y(n210) );
  MUX21X1_HVT U87 ( .A1(n422), .A2(n696), .S0(n369), .Y(n638) );
  AND3X1_HVT U88 ( .A1(n426), .A2(n661), .A3(n636), .Y(n637) );
  INVX1_HVT U89 ( .A(n496), .Y(n341) );
  MUX21X1_HVT U91 ( .A1(n489), .A2(n479), .S0(n441), .Y(n650) );
  OA21X1_HVT U92 ( .A1(n466), .A2(n437), .A3(n467), .Y(n606) );
  INVX0_HVT U93 ( .A(n680), .Y(n466) );
  MUX21X1_HVT U94 ( .A1(n605), .A2(n686), .S0(n23), .Y(n603) );
  NAND2X0_HVT U95 ( .A1(n591), .A2(n375), .Y(n349) );
  MUX21X1_HVT U96 ( .A1(n469), .A2(n593), .S0(n435), .Y(n592) );
  MUX21X1_HVT U97 ( .A1(n596), .A2(n597), .S0(n411), .Y(n595) );
  MUX21X1_HVT U98 ( .A1(n624), .A2(n625), .S0(n408), .Y(n622) );
  INVX0_HVT U99 ( .A(n437), .Y(n435) );
  INVX1_HVT U100 ( .A(n23), .Y(n316) );
  INVX1_HVT U102 ( .A(n412), .Y(n213) );
  INVX1_HVT U104 ( .A(n261), .Y(n375) );
  INVX1_HVT U105 ( .A(n440), .Y(n211) );
  NBUFFX2_HVT U106 ( .A(n443), .Y(n412) );
  INVX1_HVT U107 ( .A(n716), .Y(n305) );
  INVX0_HVT U108 ( .A(n446), .Y(n444) );
  NBUFFX2_HVT U109 ( .A(n439), .Y(n409) );
  INVX1_HVT U111 ( .A(in[6]), .Y(n344) );
  INVX1_HVT U112 ( .A(n431), .Y(n243) );
  INVX1_HVT U113 ( .A(n710), .Y(n354) );
  INVX0_HVT U114 ( .A(n378), .Y(n685) );
  MUX21X1_HVT U116 ( .A1(n417), .A2(n423), .S0(n312), .Y(n378) );
  INVX0_HVT U117 ( .A(in[7]), .Y(n446) );
  MUX21X1_HVT U119 ( .A1(n307), .A2(n283), .S0(n432), .Y(n325) );
  INVX0_HVT U120 ( .A(n325), .Y(n690) );
  INVX0_HVT U121 ( .A(n415), .Y(n46) );
  INVX0_HVT U122 ( .A(n46), .Y(n48) );
  MUX21X1_HVT U124 ( .A1(n423), .A2(n414), .S0(n362), .Y(n708) );
  XNOR2X2_HVT U125 ( .A1(n319), .A2(n325), .Y(n673) );
  MUX41X1_HVT U126 ( .A1(n691), .A3(n646), .A2(n693), .A4(n645), .S0(n210), 
        .S1(n443), .Y(n643) );
  MUX41X1_HVT U127 ( .A1(n643), .A3(n647), .A2(n640), .A4(n642), .S0(n438), 
        .S1(n387), .Y(n639) );
  INVX1_HVT U128 ( .A(n696), .Y(n455) );
  MUX41X1_HVT U129 ( .A1(n423), .A3(n471), .A2(n480), .A4(n454), .S0(n336), 
        .S1(n404), .Y(n534) );
  MUX41X1_HVT U130 ( .A1(n611), .A3(n616), .A2(n609), .A4(n612), .S0(n413), 
        .S1(n211), .Y(n608) );
  MUX41X1_HVT U131 ( .A1(n650), .A3(n652), .A2(n459), .A4(n651), .S0(n436), 
        .S1(n256), .Y(n649) );
  MUX41X1_HVT U132 ( .A1(n708), .A3(n458), .A2(n395), .A4(n326), .S0(n319), 
        .S1(n434), .Y(n536) );
  MUX41X1_HVT U133 ( .A1(n536), .A3(n538), .A2(n537), .A4(n540), .S0(n413), 
        .S1(n439), .Y(n535) );
  MUX41X1_HVT U134 ( .A1(n546), .A3(n551), .A2(n543), .A4(n549), .S0(n413), 
        .S1(n211), .Y(n542) );
  INVX0_HVT U137 ( .A(n709), .Y(n459) );
  MUX41X1_HVT U138 ( .A1(n271), .A3(n351), .A2(n416), .A4(n482), .S0(n442), 
        .S1(n403), .Y(n512) );
  MUX21X1_HVT U139 ( .A1(n354), .A2(n304), .S0(n428), .Y(n709) );
  INVX0_HVT U141 ( .A(n700), .Y(n460) );
  MUX21X2_HVT U143 ( .A1(n397), .A2(n460), .S0(n407), .Y(n583) );
  MUX41X1_HVT U144 ( .A1(n515), .A3(n513), .A2(n514), .A4(n512), .S0(n387), 
        .S1(n211), .Y(n511) );
  INVX1_HVT U145 ( .A(in[2]), .Y(n437) );
  MUX41X1_HVT U146 ( .A1(n601), .A3(n607), .A2(n603), .A4(n606), .S0(n439), 
        .S1(n375), .Y(n600) );
  INVX1_HVT U148 ( .A(n710), .Y(n353) );
  INVX1_HVT U149 ( .A(in[1]), .Y(n433) );
  AO21X1_HVT U150 ( .A1(n412), .A2(n623), .A3(n487), .Y(n624) );
  INVX1_HVT U151 ( .A(n692), .Y(n448) );
  MUX21X1_HVT U152 ( .A1(n451), .A2(n358), .S0(n243), .Y(n692) );
  MUX21X1_HVT U155 ( .A1(n473), .A2(n304), .S0(n433), .Y(n679) );
  MUX41X1_HVT U156 ( .A1(n585), .A3(n583), .A2(n584), .A4(n582), .S0(n211), 
        .S1(n261), .Y(n581) );
  MUX41X1_HVT U157 ( .A1(n476), .A3(n610), .A2(n671), .A4(n485), .S0(n337), 
        .S1(n336), .Y(n609) );
  INVX0_HVT U160 ( .A(n623), .Y(n474) );
  MUX41X1_HVT U161 ( .A1(n685), .A3(n705), .A2(n449), .A4(n681), .S0(n337), 
        .S1(n256), .Y(n514) );
  MUX21X2_HVT U164 ( .A1(n516), .A2(n517), .S0(n406), .Y(n515) );
  MUX41X1_HVT U165 ( .A1(n600), .A3(n594), .A2(n586), .A4(n581), .S0(n387), 
        .S1(n344), .Y(out[3]) );
  INVX1_HVT U169 ( .A(n297), .Y(n682) );
  MUX21X1_HVT U170 ( .A1(n666), .A2(n667), .S0(n410), .Y(n664) );
  INVX0_HVT U171 ( .A(n444), .Y(n336) );
  INVX0_HVT U172 ( .A(in[1]), .Y(n432) );
  INVX1_HVT U173 ( .A(n354), .Y(n355) );
  NBUFFX2_HVT U175 ( .A(n433), .Y(n212) );
  INVX1_HVT U178 ( .A(n358), .Y(n359) );
  OR2X1_HVT U179 ( .A1(n496), .A2(n243), .Y(n363) );
  NAND2X0_HVT U180 ( .A1(n447), .A2(n374), .Y(n216) );
  NAND2X0_HVT U181 ( .A1(n580), .A2(n407), .Y(n217) );
  NAND2X0_HVT U182 ( .A1(n216), .A2(n217), .Y(n579) );
  MUX21X1_HVT U183 ( .A1(n422), .A2(n472), .S0(n369), .Y(n580) );
  NAND2X0_HVT U184 ( .A1(n692), .A2(n210), .Y(n218) );
  NAND2X0_HVT U185 ( .A1(n470), .A2(n435), .Y(n219) );
  NAND2X0_HVT U186 ( .A1(n218), .A2(n219), .Y(n385) );
  OR2X1_HVT U187 ( .A1(n243), .A2(n304), .Y(n644) );
  NAND2X0_HVT U188 ( .A1(n713), .A2(n407), .Y(n224) );
  NAND2X0_HVT U190 ( .A1(n576), .A2(n210), .Y(n231) );
  NAND2X0_HVT U191 ( .A1(n224), .A2(n231), .Y(n575) );
  NAND2X0_HVT U192 ( .A1(n473), .A2(n430), .Y(n232) );
  NAND2X0_HVT U193 ( .A1(n414), .A2(n243), .Y(n236) );
  NAND2X0_HVT U198 ( .A1(n232), .A2(n236), .Y(n678) );
  INVX0_HVT U200 ( .A(n678), .Y(n471) );
  MUX21X1_HVT U201 ( .A1(n509), .A2(n687), .S0(n213), .Y(n504) );
  INVX1_HVT U202 ( .A(n712), .Y(n473) );
  INVX1_HVT U203 ( .A(n420), .Y(n238) );
  INVX1_HVT U204 ( .A(n238), .Y(n240) );
  INVX1_HVT U205 ( .A(n502), .Y(n462) );
  NBUFFX2_HVT U206 ( .A(n481), .Y(n418) );
  INVX1_HVT U207 ( .A(n417), .Y(n301) );
  INVX1_HVT U209 ( .A(n431), .Y(n312) );
  INVX1_HVT U210 ( .A(n243), .Y(n252) );
  INVX1_HVT U211 ( .A(n504), .Y(n447) );
  IBUFFX2_HVT U213 ( .A(n380), .Y(n429) );
  AND2X1_HVT U216 ( .A1(n364), .A2(n363), .Y(n264) );
  INVX1_HVT U217 ( .A(n456), .Y(n271) );
  NAND2X0_HVT U219 ( .A1(n212), .A2(n440), .Y(n278) );
  NAND2X0_HVT U221 ( .A1(n478), .A2(n441), .Y(n280) );
  NAND2X0_HVT U222 ( .A1(n278), .A2(n280), .Y(n652) );
  INVX1_HVT U223 ( .A(n705), .Y(n478) );
  INVX1_HVT U224 ( .A(n425), .Y(n282) );
  INVX0_HVT U225 ( .A(n661), .Y(n491) );
  MUX21X1_HVT U226 ( .A1(n414), .A2(n682), .S0(n409), .Y(n667) );
  MUX21X1_HVT U227 ( .A1(n414), .A2(n418), .S0(n412), .Y(n626) );
  INVX0_HVT U228 ( .A(n309), .Y(n697) );
  MUX41X1_HVT U229 ( .A1(n498), .A3(n399), .A2(n490), .A4(n621), .S0(n435), 
        .S1(n444), .Y(n620) );
  INVX1_HVT U230 ( .A(n315), .Y(n621) );
  NAND2X0_HVT U231 ( .A1(n471), .A2(n375), .Y(n360) );
  XNOR2X1_HVT U232 ( .A1(n710), .A2(n433), .Y(n672) );
  MUX21X1_HVT U233 ( .A1(n418), .A2(n716), .S0(n430), .Y(n284) );
  MUX41X1_HVT U234 ( .A1(n622), .A3(n627), .A2(n619), .A4(n620), .S0(n438), 
        .S1(n387), .Y(n618) );
  NAND2X0_HVT U235 ( .A1(n626), .A2(n400), .Y(n293) );
  NAND2X0_HVT U236 ( .A1(n290), .A2(n293), .Y(n625) );
  NAND2X0_HVT U237 ( .A1(n428), .A2(n426), .Y(n714) );
  INVX1_HVT U238 ( .A(n499), .Y(n482) );
  MUX41X1_HVT U239 ( .A1(n568), .A3(n567), .A2(n572), .A4(n571), .S0(n211), 
        .S1(n413), .Y(n566) );
  NOR2X0_HVT U240 ( .A1(n301), .A2(n379), .Y(n297) );
  MUX41X1_HVT U243 ( .A1(n482), .A3(n689), .A2(n483), .A4(n464), .S0(n337), 
        .S1(n442), .Y(n537) );
  MUX41X1_HVT U244 ( .A1(n539), .A3(n699), .A2(n679), .A4(n483), .S0(n374), 
        .S1(n442), .Y(n538) );
  INVX1_HVT U246 ( .A(n352), .Y(n400) );
  MUX21X1_HVT U248 ( .A1(n424), .A2(n356), .S0(n362), .Y(n680) );
  MUX21X1_HVT U249 ( .A1(n341), .A2(n354), .S0(n379), .Y(n340) );
  MUX21X1_HVT U251 ( .A1(n212), .A2(n271), .S0(n23), .Y(n589) );
  INVX1_HVT U252 ( .A(n335), .Y(n550) );
  NBUFFX2_HVT U253 ( .A(n415), .Y(n416) );
  INVX1_HVT U254 ( .A(n716), .Y(n303) );
  INVX1_HVT U257 ( .A(n716), .Y(n304) );
  INVX1_HVT U258 ( .A(n305), .Y(n306) );
  INVX1_HVT U260 ( .A(n305), .Y(n307) );
  INVX0_HVT U261 ( .A(n702), .Y(n331) );
  INVX1_HVT U262 ( .A(n455), .Y(n330) );
  XNOR2X2_HVT U263 ( .A1(n481), .A2(n308), .Y(n710) );
  MUX41X1_HVT U264 ( .A1(n706), .A3(n662), .A2(n697), .A4(n463), .S0(n336), 
        .S1(n441), .Y(n660) );
  INVX0_HVT U267 ( .A(n701), .Y(n457) );
  INVX1_HVT U269 ( .A(n444), .Y(n319) );
  NAND2X0_HVT U272 ( .A1(n565), .A2(n407), .Y(n310) );
  NAND2X0_HVT U273 ( .A1(n564), .A2(n374), .Y(n311) );
  NAND2X0_HVT U274 ( .A1(n310), .A2(n311), .Y(n562) );
  NAND2X0_HVT U275 ( .A1(n419), .A2(n312), .Y(n313) );
  NAND2X0_HVT U276 ( .A1(n451), .A2(n428), .Y(n314) );
  NAND2X0_HVT U277 ( .A1(n313), .A2(n314), .Y(n677) );
  NBUFFX2_HVT U278 ( .A(n496), .Y(n419) );
  MUX21X1_HVT U279 ( .A1(n355), .A2(n423), .S0(n362), .Y(n315) );
  INVX0_HVT U280 ( .A(n707), .Y(n327) );
  NAND2X0_HVT U282 ( .A1(n378), .A2(n316), .Y(n317) );
  NAND2X0_HVT U286 ( .A1(n699), .A2(n210), .Y(n318) );
  NAND2X0_HVT U287 ( .A1(n317), .A2(n318), .Y(n582) );
  MUX21X1_HVT U288 ( .A1(n416), .A2(n327), .S0(n429), .Y(n699) );
  MUX41X1_HVT U290 ( .A1(n701), .A3(n428), .A2(n399), .A4(n491), .S0(n374), 
        .S1(n319), .Y(n619) );
  INVX0_HVT U291 ( .A(n699), .Y(n486) );
  NAND2X0_HVT U292 ( .A1(n654), .A2(n23), .Y(n365) );
  NAND2X0_HVT U293 ( .A1(n664), .A2(n337), .Y(n320) );
  NAND2X0_HVT U294 ( .A1(n668), .A2(n407), .Y(n321) );
  NAND2X0_HVT U296 ( .A1(n320), .A2(n321), .Y(n663) );
  NAND2X0_HVT U298 ( .A1(n602), .A2(n322), .Y(n323) );
  NAND2X0_HVT U299 ( .A1(n427), .A2(n670), .Y(n324) );
  NAND2X0_HVT U301 ( .A1(n323), .A2(n324), .Y(n601) );
  INVX0_HVT U304 ( .A(n670), .Y(n322) );
  MUX41X1_HVT U305 ( .A1(n579), .A3(n577), .A2(n578), .A4(n575), .S0(n387), 
        .S1(n211), .Y(n574) );
  MUX41X1_HVT U308 ( .A1(n557), .A3(n562), .A2(n555), .A4(n561), .S0(n413), 
        .S1(n211), .Y(n554) );
  NAND2X0_HVT U309 ( .A1(n703), .A2(n306), .Y(n326) );
  INVX0_HVT U310 ( .A(n327), .Y(n328) );
  INVX1_HVT U311 ( .A(n403), .Y(n405) );
  MUX41X1_HVT U312 ( .A1(n694), .A3(n493), .A2(n704), .A4(n662), .S0(n337), 
        .S1(n256), .Y(n513) );
  MUX21X1_HVT U313 ( .A1(n587), .A2(n588), .S0(n409), .Y(n586) );
  INVX1_HVT U314 ( .A(n329), .Y(n634) );
  MUX41X1_HVT U315 ( .A1(n488), .A3(n631), .A2(n398), .A4(n394), .S0(n435), 
        .S1(n410), .Y(n630) );
  MUX41X1_HVT U316 ( .A1(n693), .A3(n331), .A2(n332), .A4(n330), .S0(n435), 
        .S1(n369), .Y(n329) );
  XNOR2X1_HVT U317 ( .A1(n252), .A2(n489), .Y(n332) );
  NAND2X0_HVT U318 ( .A1(n595), .A2(n211), .Y(n333) );
  NAND2X0_HVT U319 ( .A1(n598), .A2(n409), .Y(n334) );
  NAND2X0_HVT U320 ( .A1(n333), .A2(n334), .Y(n594) );
  INVX1_HVT U321 ( .A(n503), .Y(n472) );
  MUX21X1_HVT U322 ( .A1(n283), .A2(n240), .S0(n212), .Y(n335) );
  MUX41X1_HVT U323 ( .A1(n484), .A3(n695), .A2(n550), .A4(n672), .S0(n336), 
        .S1(n404), .Y(n549) );
  MUX21X1_HVT U324 ( .A1(n340), .A2(n489), .S0(n411), .Y(n565) );
  MUX21X1_HVT U325 ( .A1(n427), .A2(n421), .S0(n339), .Y(n702) );
  NAND2X0_HVT U326 ( .A1(n673), .A2(n374), .Y(n342) );
  NAND2X0_HVT U327 ( .A1(n648), .A2(n406), .Y(n343) );
  NAND2X0_HVT U328 ( .A1(n342), .A2(n343), .Y(n647) );
  NAND2X0_HVT U329 ( .A1(n629), .A2(n344), .Y(n345) );
  NAND2X0_HVT U330 ( .A1(n639), .A2(in[6]), .Y(n346) );
  NAND2X0_HVT U331 ( .A1(n345), .A2(n346), .Y(out[1]) );
  MUX21X1_HVT U332 ( .A1(n304), .A2(n490), .S0(n412), .Y(n648) );
  NAND2X0_HVT U333 ( .A1(n526), .A2(n344), .Y(n347) );
  NAND2X0_HVT U334 ( .A1(n535), .A2(in[6]), .Y(n348) );
  NAND2X0_HVT U335 ( .A1(n347), .A2(n348), .Y(out[6]) );
  NAND2X0_HVT U336 ( .A1(n592), .A2(n369), .Y(n350) );
  NAND2X0_HVT U337 ( .A1(n349), .A2(n350), .Y(n588) );
  XOR2X1_HVT U338 ( .A1(in[7]), .A2(n433), .Y(n352) );
  INVX1_HVT U339 ( .A(n353), .Y(n356) );
  INVX1_HVT U340 ( .A(n354), .Y(n358) );
  NAND2X0_HVT U341 ( .A1(n694), .A2(n336), .Y(n361) );
  NAND2X0_HVT U342 ( .A1(n360), .A2(n361), .Y(n576) );
  NAND2X0_HVT U343 ( .A1(n353), .A2(n432), .Y(n364) );
  NAND2X0_HVT U344 ( .A1(n363), .A2(n364), .Y(n694) );
  NAND2X0_HVT U345 ( .A1(n656), .A2(n406), .Y(n366) );
  NAND2X0_HVT U346 ( .A1(n365), .A2(n366), .Y(n653) );
  OA21X1_HVT U347 ( .A1(n256), .A2(n709), .A3(n470), .Y(n516) );
  MUX41X1_HVT U348 ( .A1(n695), .A3(n402), .A2(n459), .A4(n472), .S0(n316), 
        .S1(n375), .Y(n587) );
  MUX41X1_HVT U349 ( .A1(n635), .A3(n634), .A2(n632), .A4(n630), .S0(n211), 
        .S1(n387), .Y(n629) );
  NAND2X0_HVT U350 ( .A1(n658), .A2(n337), .Y(n367) );
  NAND2X0_HVT U351 ( .A1(n660), .A2(n406), .Y(n368) );
  NAND2X0_HVT U352 ( .A1(n367), .A2(n368), .Y(n657) );
  NAND2X0_HVT U353 ( .A1(n570), .A2(n337), .Y(n370) );
  NAND2X0_HVT U354 ( .A1(n569), .A2(n407), .Y(n371) );
  NAND2X0_HVT U355 ( .A1(n370), .A2(n371), .Y(n568) );
  NAND2X0_HVT U356 ( .A1(n566), .A2(n344), .Y(n372) );
  NAND2X0_HVT U357 ( .A1(n574), .A2(in[6]), .Y(n373) );
  NAND2X0_HVT U358 ( .A1(n373), .A2(n372), .Y(out[4]) );
  INVX1_HVT U359 ( .A(n506), .Y(n490) );
  MUX41X1_HVT U360 ( .A1(n672), .A3(n644), .A2(n678), .A4(n399), .S0(n374), 
        .S1(n261), .Y(n530) );
  NAND2X0_HVT U361 ( .A1(n386), .A2(n375), .Y(n376) );
  NAND2X0_HVT U362 ( .A1(n385), .A2(n319), .Y(n377) );
  NAND2X0_HVT U363 ( .A1(n377), .A2(n376), .Y(n572) );
  MUX41X1_HVT U364 ( .A1(n686), .A3(n448), .A2(n599), .A4(n326), .S0(n374), 
        .S1(n319), .Y(n598) );
  MUX41X1_HVT U365 ( .A1(n527), .A3(n530), .A2(n531), .A4(n534), .S0(n439), 
        .S1(n413), .Y(n526) );
  NAND2X0_HVT U366 ( .A1(n518), .A2(in[6]), .Y(n381) );
  NAND2X0_HVT U367 ( .A1(n511), .A2(n344), .Y(n382) );
  NAND2X0_HVT U368 ( .A1(n381), .A2(n382), .Y(out[7]) );
  INVX0_HVT U369 ( .A(n683), .Y(n493) );
  MUX21X1_HVT U370 ( .A1(n297), .A2(n493), .S0(n406), .Y(n597) );
  INVX0_HVT U371 ( .A(n446), .Y(n443) );
  INVX1_HVT U372 ( .A(n446), .Y(n445) );
  MUX41X1_HVT U373 ( .A1(n525), .A3(n669), .A2(n682), .A4(n675), .S0(n403), 
        .S1(n261), .Y(n524) );
  NAND2X0_HVT U374 ( .A1(n554), .A2(in[6]), .Y(n383) );
  NAND2X0_HVT U375 ( .A1(n542), .A2(n344), .Y(n384) );
  NAND2X0_HVT U376 ( .A1(n383), .A2(n384), .Y(out[5]) );
  INVX1_HVT U377 ( .A(in[0]), .Y(n387) );
  NAND2X0_HVT U378 ( .A1(n618), .A2(in[6]), .Y(n389) );
  NAND2X0_HVT U379 ( .A1(n608), .A2(n344), .Y(n388) );
  NAND2X0_HVT U380 ( .A1(n389), .A2(n388), .Y(out[2]) );
  NAND2X0_HVT U381 ( .A1(n617), .A2(n390), .Y(n391) );
  NAND2X0_HVT U382 ( .A1(n396), .A2(n393), .Y(n392) );
  NAND2X0_HVT U383 ( .A1(n391), .A2(n392), .Y(n616) );
  INVX0_HVT U384 ( .A(n393), .Y(n390) );
  INVX1_HVT U385 ( .A(n441), .Y(n440) );
  INVX0_HVT U386 ( .A(n437), .Y(n436) );
  INVX1_HVT U387 ( .A(in[5]), .Y(n441) );
  NBUFFX2_HVT U388 ( .A(n712), .Y(n423) );
  NBUFFX2_HVT U389 ( .A(n712), .Y(n424) );
  AND2X1_HVT U390 ( .A1(n426), .A2(n644), .Y(n394) );
  AND2X1_HVT U391 ( .A1(n359), .A2(n661), .Y(n395) );
  AND2X1_HVT U392 ( .A1(n307), .A2(n604), .Y(n396) );
  NAND2X0_HVT U393 ( .A1(n481), .A2(n308), .Y(n712) );
  MUX21X1_HVT U394 ( .A1(n422), .A2(n307), .S0(n407), .Y(n590) );
  MUX21X1_HVT U395 ( .A1(n303), .A2(n496), .S0(n429), .Y(n683) );
  MUX21X1_HVT U396 ( .A1(n426), .A2(n357), .S0(n338), .Y(n676) );
  MUX21X1_HVT U397 ( .A1(n419), .A2(n304), .S0(n429), .Y(n706) );
  MUX21X1_HVT U398 ( .A1(n424), .A2(n419), .S0(n252), .Y(n705) );
  MUX21X1_HVT U399 ( .A1(n303), .A2(n357), .S0(n338), .Y(n553) );
  XOR2X1_HVT U400 ( .A1(n283), .A2(n362), .Y(n669) );
  MUX21X1_HVT U401 ( .A1(n496), .A2(n417), .S0(n429), .Y(n525) );
  MUX21X1_HVT U402 ( .A1(n418), .A2(n419), .S0(n339), .Y(n593) );
  MUX21X1_HVT U403 ( .A1(n424), .A2(n422), .S0(n362), .Y(n628) );
  MUX21X1_HVT U404 ( .A1(n421), .A2(n496), .S0(n339), .Y(n506) );
  MUX21X1_HVT U405 ( .A1(n327), .A2(n473), .S0(n252), .Y(n698) );
  MUX21X1_HVT U406 ( .A1(n359), .A2(n418), .S0(n379), .Y(n613) );
  MUX21X1_HVT U407 ( .A1(n422), .A2(n417), .S0(n379), .Y(n646) );
  MUX21X1_HVT U408 ( .A1(n356), .A2(n418), .S0(n379), .Y(n641) );
  MUX21X1_HVT U409 ( .A1(n419), .A2(n306), .S0(n338), .Y(n528) );
  MUX21X1_HVT U410 ( .A1(n307), .A2(n427), .S0(n428), .Y(n529) );
  MUX21X1_HVT U411 ( .A1(n283), .A2(n417), .S0(n362), .Y(n508) );
  MUX21X1_HVT U412 ( .A1(n358), .A2(n489), .S0(n379), .Y(n502) );
  MUX21X1_HVT U413 ( .A1(n424), .A2(n306), .S0(n431), .Y(n623) );
  MUX21X1_HVT U414 ( .A1(n473), .A2(n417), .S0(n428), .Y(n503) );
  MUX21X1_HVT U415 ( .A1(n283), .A2(n423), .S0(n430), .Y(n501) );
  XOR2X1_HVT U416 ( .A1(n417), .A2(n429), .Y(n691) );
  XNOR2X1_HVT U417 ( .A1(n423), .A2(n431), .Y(n397) );
  MUX21X1_HVT U418 ( .A1(n473), .A2(n303), .S0(n409), .Y(n665) );
  XOR2X1_HVT U419 ( .A1(n430), .A2(n439), .Y(n674) );
  XNOR2X1_HVT U420 ( .A1(n306), .A2(n429), .Y(n398) );
  AND2X1_HVT U421 ( .A1(n252), .A2(n451), .Y(n399) );
  NBUFFX2_HVT U422 ( .A(n707), .Y(n420) );
  NBUFFX2_HVT U423 ( .A(n328), .Y(n421) );
  NBUFFX2_HVT U424 ( .A(n715), .Y(n425) );
  NBUFFX2_HVT U425 ( .A(n328), .Y(n422) );
  NBUFFX2_HVT U426 ( .A(n715), .Y(n426) );
  NBUFFX2_HVT U427 ( .A(n715), .Y(n427) );
  NBUFFX2_HVT U428 ( .A(n481), .Y(n417) );
  NBUFFX2_HVT U429 ( .A(n443), .Y(n411) );
  NBUFFX2_HVT U430 ( .A(n443), .Y(n410) );
  NBUFFX2_HVT U431 ( .A(n436), .Y(n407) );
  NBUFFX2_HVT U432 ( .A(n436), .Y(n406) );
  MUX21X1_HVT U433 ( .A1(n560), .A2(n427), .S0(n400), .Y(n559) );
  MUX21X1_HVT U434 ( .A1(n545), .A2(n544), .S0(n407), .Y(n543) );
  MUX21X1_HVT U435 ( .A1(n422), .A2(n490), .S0(n412), .Y(n545) );
  MUX21X1_HVT U436 ( .A1(n416), .A2(n421), .S0(n338), .Y(n500) );
  MUX21X1_HVT U437 ( .A1(n631), .A2(n414), .S0(n411), .Y(n533) );
  MUX21X1_HVT U438 ( .A1(n307), .A2(n416), .S0(n430), .Y(n689) );
  MUX21X1_HVT U439 ( .A1(n421), .A2(n357), .S0(n338), .Y(n610) );
  MUX21X1_HVT U440 ( .A1(n416), .A2(n306), .S0(n379), .Y(n499) );
  MUX21X1_HVT U441 ( .A1(n414), .A2(n489), .S0(n338), .Y(n505) );
  MUX21X1_HVT U442 ( .A1(n416), .A2(n355), .S0(n339), .Y(n507) );
  MUX21X1_HVT U443 ( .A1(n414), .A2(n416), .S0(n406), .Y(n602) );
  NAND2X0_HVT U444 ( .A1(n48), .A2(n308), .Y(n707) );
  NAND2X0_HVT U445 ( .A1(in[3]), .A2(n48), .Y(n716) );
  AND2X1_HVT U446 ( .A1(n357), .A2(n312), .Y(n401) );
  NAND2X0_HVT U447 ( .A1(in[3]), .A2(n481), .Y(n715) );
  AND2X1_HVT U448 ( .A1(n419), .A2(n212), .Y(n402) );
  INVX1_HVT U449 ( .A(n437), .Y(n434) );
  NBUFFX2_HVT U450 ( .A(n440), .Y(n439) );
  NBUFFX2_HVT U451 ( .A(n440), .Y(n438) );
  NBUFFX2_HVT U452 ( .A(in[3]), .Y(n414) );
  NBUFFX2_HVT U453 ( .A(in[4]), .Y(n415) );
  NBUFFX2_HVT U454 ( .A(in[0]), .Y(n413) );
endmodule

