
module sbox_15 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n38, n47, n50, n113, n114, n117, n118, n119, n127, n204, n210,
         n211, n212, n213, n216, n217, n218, n219, n222, n224, n227, n229,
         n231, n232, n236, n238, n241, n242, n245, n246, n252, n253, n257,
         n258, n259, n261, n263, n264, n270, n271, n273, n274, n275, n278,
         n279, n280, n282, n283, n285, n289, n293, n296, n297, n300, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757;

  NAND2X0_HVT U4 ( .A1(n216), .A2(n755), .Y(n754) );
  NAND2X0_HVT U5 ( .A1(n293), .A2(n493), .Y(n752) );
  NAND2X0_HVT U15 ( .A1(n755), .A2(n236), .Y(n742) );
  NAND2X0_HVT U21 ( .A1(n216), .A2(n451), .Y(n736) );
  NAND2X0_HVT U24 ( .A1(n453), .A2(n353), .Y(n734) );
  NAND2X0_HVT U33 ( .A1(n333), .A2(n353), .Y(n725) );
  NAND2X0_HVT U42 ( .A1(n439), .A2(n331), .Y(n717) );
  MUX41X1_HVT U51 ( .A1(n516), .A3(n534), .A2(n512), .A4(n518), .S0(n462), 
        .S1(n483), .Y(n710) );
  NAND2X0_HVT U53 ( .A1(n707), .A2(n716), .Y(n708) );
  NAND2X0_HVT U56 ( .A1(n216), .A2(n703), .Y(n704) );
  MUX41X1_HVT U57 ( .A1(n525), .A3(n738), .A2(n704), .A4(n747), .S0(n462), 
        .S1(n483), .Y(n702) );
  MUX41X1_HVT U61 ( .A1(n467), .A3(n540), .A2(n452), .A4(n236), .S0(n461), 
        .S1(n483), .Y(n698) );
  NAND2X0_HVT U62 ( .A1(n451), .A2(n497), .Y(n697) );
  AO21X1_HVT U66 ( .A1(n407), .A2(n506), .A3(n546), .Y(n693) );
  NAND2X0_HVT U73 ( .A1(n428), .A2(n686), .Y(n687) );
  MUX41X1_HVT U77 ( .A1(n749), .A3(n532), .A2(n683), .A4(n448), .S0(n484), 
        .S1(n473), .Y(n682) );
  MUX41X1_HVT U82 ( .A1(n714), .A3(n518), .A2(n550), .A4(n743), .S0(n473), 
        .S1(n462), .Y(n676) );
  AND2X1_HVT U83 ( .A1(n438), .A2(n406), .Y(n675) );
  MUX41X1_HVT U84 ( .A1(n523), .A3(n332), .A2(n741), .A4(n675), .S0(n503), 
        .S1(n390), .Y(n674) );
  NAND2X0_HVT U85 ( .A1(n451), .A2(n545), .Y(n673) );
  NAND2X0_HVT U101 ( .A1(n656), .A2(n655), .Y(n657) );
  MUX41X1_HVT U103 ( .A1(n755), .A3(n339), .A2(n527), .A4(n723), .S0(n379), 
        .S1(n245), .Y(n653) );
  NAND2X0_HVT U110 ( .A1(n257), .A2(n648), .Y(n649) );
  AND2X1_HVT U115 ( .A1(n439), .A2(n236), .Y(n646) );
  NAND2X0_HVT U123 ( .A1(n638), .A2(n637), .Y(n639) );
  MUX41X1_HVT U125 ( .A1(n736), .A3(n471), .A2(n522), .A4(n530), .S0(n340), 
        .S1(n485), .Y(n635) );
  MUX41X1_HVT U135 ( .A1(n38), .A3(n425), .A2(n752), .A4(n313), .S0(n335), 
        .S1(n461), .Y(n626) );
  MUX41X1_HVT U136 ( .A1(n464), .A3(n725), .A2(n515), .A4(n722), .S0(n480), 
        .S1(n461), .Y(n625) );
  AND2X1_HVT U140 ( .A1(n428), .A2(n451), .Y(n621) );
  MUX41X1_HVT U153 ( .A1(n649), .A3(n467), .A2(n257), .A4(n535), .S0(n319), 
        .S1(n390), .Y(n609) );
  AND2X1_HVT U154 ( .A1(n486), .A2(n408), .Y(n608) );
  NAND2X0_HVT U158 ( .A1(n440), .A2(n545), .Y(n604) );
  MUX41X1_HVT U159 ( .A1(n329), .A3(n489), .A2(n604), .A4(n547), .S0(n472), 
        .S1(n507), .Y(n603) );
  AND2X1_HVT U162 ( .A1(n332), .A2(n270), .Y(n600) );
  MUX41X1_HVT U165 ( .A1(n736), .A3(n538), .A2(n113), .A4(n598), .S0(n461), 
        .S1(n473), .Y(n597) );
  NAND2X0_HVT U166 ( .A1(n499), .A2(n703), .Y(n596) );
  NAND2X0_HVT U167 ( .A1(n410), .A2(n451), .Y(n595) );
  MUX41X1_HVT U168 ( .A1(n525), .A3(n422), .A2(n595), .A4(n596), .S0(n472), 
        .S1(n229), .Y(n594) );
  MUX41X1_HVT U172 ( .A1(n591), .A3(n597), .A2(n594), .A4(n599), .S0(n488), 
        .S1(n482), .Y(n590) );
  NAND2X0_HVT U177 ( .A1(n119), .A2(n490), .Y(n587) );
  MUX41X1_HVT U178 ( .A1(n740), .A3(n587), .A2(n419), .A4(n721), .S0(n319), 
        .S1(n507), .Y(n586) );
  MUX41X1_HVT U179 ( .A1(n730), .A3(n537), .A2(n526), .A4(n419), .S0(n472), 
        .S1(n229), .Y(n585) );
  MUX41X1_HVT U180 ( .A1(n521), .A3(n749), .A2(n329), .A4(n463), .S0(n484), 
        .S1(n472), .Y(n584) );
  MUX41X1_HVT U186 ( .A1(n466), .A3(n720), .A2(n270), .A4(n113), .S0(n472), 
        .S1(n461), .Y(n578) );
  MUX41X1_HVT U189 ( .A1(n576), .A3(n744), .A2(n577), .A4(n533), .S0(n484), 
        .S1(n472), .Y(n575) );
  MUX41X1_HVT U190 ( .A1(n575), .A3(n578), .A2(n579), .A4(n582), .S0(n505), 
        .S1(n488), .Y(n574) );
  AO21X1_HVT U197 ( .A1(n468), .A2(n485), .A3(n541), .Y(n568) );
  NAND2X0_HVT U208 ( .A1(n434), .A2(n495), .Y(n648) );
  NAND2X0_HVT U212 ( .A1(n119), .A2(n400), .Y(n703) );
  NAND2X0_HVT U214 ( .A1(n372), .A2(n353), .Y(n559) );
  NAND2X0_HVT U215 ( .A1(n648), .A2(n428), .Y(n558) );
  NAND2X0_HVT U218 ( .A1(n424), .A2(n441), .Y(n611) );
  NAND2X0_HVT U220 ( .A1(n485), .A2(n559), .Y(n678) );
  INVX0_HVT U241 ( .A(n734), .Y(n550) );
  INVX0_HVT U242 ( .A(n717), .Y(n549) );
  INVX0_HVT U245 ( .A(n752), .Y(n547) );
  INVX0_HVT U251 ( .A(n727), .Y(n544) );
  INVX0_HVT U252 ( .A(n703), .Y(n543) );
  INVX0_HVT U256 ( .A(n611), .Y(n541) );
  INVX0_HVT U264 ( .A(n723), .Y(n535) );
  INVX0_HVT U268 ( .A(n736), .Y(n534) );
  INVX0_HVT U284 ( .A(n559), .Y(n526) );
  INVX0_HVT U289 ( .A(n655), .Y(n524) );
  INVX0_HVT U295 ( .A(n754), .Y(n521) );
  INVX0_HVT U302 ( .A(n557), .Y(n516) );
  INVX0_HVT U306 ( .A(n595), .Y(n514) );
  INVX0_HVT U307 ( .A(n719), .Y(n513) );
  INVX0_HVT U309 ( .A(n738), .Y(n512) );
  XNOR2X1_HVT U1 ( .A1(n450), .A2(n385), .Y(n470) );
  NBUFFX2_HVT U2 ( .A(n211), .Y(n492) );
  INVX1_HVT U3 ( .A(n502), .Y(n459) );
  AND3X1_HVT U6 ( .A1(n497), .A2(n703), .A3(n678), .Y(n679) );
  INVX1_HVT U7 ( .A(n735), .Y(n523) );
  MUX21X1_HVT U8 ( .A1(n242), .A2(n400), .S0(n431), .Y(n727) );
  INVX1_HVT U9 ( .A(n442), .Y(n433) );
  OA21X1_HVT U10 ( .A1(n432), .A2(n719), .A3(n611), .Y(n612) );
  MUX21X1_HVT U11 ( .A1(n497), .A2(n421), .S0(n441), .Y(n718) );
  MUX21X1_HVT U12 ( .A1(n330), .A2(n395), .S0(n506), .Y(n694) );
  XOR2X1_HVT U13 ( .A1(n731), .A2(n432), .Y(n715) );
  INVX1_HVT U14 ( .A(n416), .Y(n340) );
  INVX1_HVT U16 ( .A(n504), .Y(n503) );
  AND2X1_HVT U17 ( .A1(n212), .A2(n213), .Y(n23) );
  AND2X1_HVT U18 ( .A1(n241), .A2(n238), .Y(n38) );
  AND2X1_HVT U19 ( .A1(n300), .A2(n303), .Y(n47) );
  AND2X1_HVT U20 ( .A1(n252), .A2(n253), .Y(n50) );
  AND2X1_HVT U22 ( .A1(n252), .A2(n253), .Y(n113) );
  INVX1_HVT U23 ( .A(n487), .Y(n114) );
  NBUFFX2_HVT U25 ( .A(n536), .Y(n491) );
  INVX1_HVT U26 ( .A(in[4]), .Y(n536) );
  NOR2X1_HVT U27 ( .A1(n459), .A2(n421), .Y(n458) );
  MUX41X1_HVT U28 ( .A1(n745), .A3(n704), .A2(n735), .A4(n327), .S0(n368), 
        .S1(n508), .Y(n562) );
  MUX21X1_HVT U29 ( .A1(n318), .A2(n460), .S0(n459), .Y(n735) );
  INVX1_HVT U30 ( .A(n117), .Y(n548) );
  MUX21X1_HVT U31 ( .A1(n465), .A2(n452), .S0(n340), .Y(n631) );
  INVX0_HVT U32 ( .A(n477), .Y(n647) );
  MUX41X1_HVT U34 ( .A1(n564), .A3(n563), .A2(n562), .A4(n561), .S0(n307), 
        .S1(n114), .Y(n560) );
  XOR2X2_HVT U35 ( .A1(n441), .A2(n423), .Y(n714) );
  MUX21X2_HVT U36 ( .A1(n545), .A2(n328), .S0(n486), .Y(n690) );
  INVX0_HVT U37 ( .A(n351), .Y(n117) );
  INVX1_HVT U38 ( .A(n460), .Y(n420) );
  XOR2X1_HVT U39 ( .A1(n433), .A2(n504), .Y(n476) );
  INVX1_HVT U40 ( .A(n338), .Y(n335) );
  INVX1_HVT U41 ( .A(n400), .Y(n427) );
  INVX1_HVT U43 ( .A(n481), .Y(n334) );
  INVX1_HVT U44 ( .A(n490), .Y(n342) );
  INVX1_HVT U45 ( .A(n510), .Y(n508) );
  INVX1_HVT U46 ( .A(n338), .Y(n379) );
  INVX1_HVT U47 ( .A(n508), .Y(n457) );
  INVX1_HVT U48 ( .A(n422), .Y(n423) );
  INVX1_HVT U49 ( .A(n558), .Y(n533) );
  INVX1_HVT U50 ( .A(n510), .Y(n507) );
  INVX1_HVT U52 ( .A(n504), .Y(n472) );
  INVX1_HVT U54 ( .A(in[2]), .Y(n504) );
  MUX21X1_HVT U55 ( .A1(n497), .A2(n668), .S0(n470), .Y(n667) );
  MUX21X1_HVT U58 ( .A1(n490), .A2(n495), .S0(n430), .Y(n429) );
  OA21X1_HVT U59 ( .A1(n514), .A2(n432), .A3(n727), .Y(n617) );
  MUX21X1_HVT U60 ( .A1(n424), .A2(n553), .S0(n412), .Y(n411) );
  MUX21X1_HVT U63 ( .A1(n529), .A2(n735), .S0(n412), .Y(n624) );
  INVX1_HVT U64 ( .A(n429), .Y(n726) );
  INVX1_HVT U65 ( .A(n743), .Y(n519) );
  MUX21X1_HVT U67 ( .A1(n339), .A2(n425), .S0(n506), .Y(n692) );
  INVX1_HVT U68 ( .A(n443), .Y(n438) );
  MUX21X1_HVT U69 ( .A1(n426), .A2(n216), .S0(n395), .Y(n670) );
  NAND2X0_HVT U70 ( .A1(n643), .A2(n275), .Y(n127) );
  MUX21X1_HVT U71 ( .A1(n640), .A2(n639), .S0(n486), .Y(n636) );
  AND3X1_HVT U72 ( .A1(n480), .A2(n395), .A3(n342), .Y(n632) );
  INVX1_HVT U74 ( .A(n728), .Y(n538) );
  MUX21X1_HVT U75 ( .A1(n612), .A2(n613), .S0(n319), .Y(n610) );
  MUX21X1_HVT U76 ( .A1(n607), .A2(n606), .S0(n334), .Y(n605) );
  XOR2X1_HVT U78 ( .A1(n342), .A2(n433), .Y(n341) );
  XOR2X1_HVT U79 ( .A1(n498), .A2(n369), .Y(n711) );
  MUX21X1_HVT U80 ( .A1(n426), .A2(n737), .S0(n450), .Y(n680) );
  XNOR2X1_HVT U81 ( .A1(n353), .A2(n408), .Y(n712) );
  INVX1_HVT U86 ( .A(n729), .Y(n527) );
  MUX21X1_HVT U87 ( .A1(n657), .A2(n511), .S0(n480), .Y(n654) );
  AO21X1_HVT U88 ( .A1(n442), .A2(n423), .A3(n432), .Y(n656) );
  INVX1_HVT U89 ( .A(n338), .Y(n319) );
  INVX1_HVT U90 ( .A(n457), .Y(n229) );
  INVX1_HVT U91 ( .A(n450), .Y(n390) );
  INVX1_HVT U92 ( .A(n479), .Y(n416) );
  INVX1_HVT U93 ( .A(n432), .Y(n245) );
  INVX1_HVT U94 ( .A(in[7]), .Y(n510) );
  INVX1_HVT U95 ( .A(n501), .Y(n430) );
  INVX1_HVT U96 ( .A(n395), .Y(n385) );
  INVX1_HVT U97 ( .A(n441), .Y(n323) );
  INVX0_HVT U98 ( .A(n441), .Y(n395) );
  INVX0_HVT U99 ( .A(n442), .Y(n434) );
  INVX1_HVT U100 ( .A(n494), .Y(n408) );
  INVX1_HVT U102 ( .A(n498), .Y(n410) );
  INVX1_HVT U104 ( .A(n497), .Y(n475) );
  INVX1_HVT U105 ( .A(n499), .Y(n118) );
  MUX21X1_HVT U106 ( .A1(n399), .A2(n423), .S0(n439), .Y(n740) );
  INVX0_HVT U107 ( .A(n750), .Y(n522) );
  INVX0_HVT U108 ( .A(n737), .Y(n518) );
  INVX1_HVT U109 ( .A(n449), .Y(n362) );
  INVX1_HVT U111 ( .A(n323), .Y(n293) );
  INVX1_HVT U112 ( .A(n351), .Y(n352) );
  INVX0_HVT U113 ( .A(n407), .Y(n747) );
  INVX0_HVT U114 ( .A(n742), .Y(n520) );
  OR2X1_HVT U116 ( .A1(n118), .A2(n397), .Y(n701) );
  INVX1_HVT U117 ( .A(n397), .Y(n755) );
  INVX1_HVT U118 ( .A(n739), .Y(n289) );
  MUX21X2_HVT U119 ( .A1(n493), .A2(n399), .S0(n501), .Y(n728) );
  MUX41X1_HVT U120 ( .A1(n571), .A3(n572), .A2(n567), .A4(n570), .S0(n482), 
        .S1(n114), .Y(n566) );
  INVX0_HVT U121 ( .A(n372), .Y(n236) );
  INVX1_HVT U122 ( .A(n377), .Y(n119) );
  INVX0_HVT U124 ( .A(n456), .Y(n381) );
  MUX21X1_HVT U126 ( .A1(n539), .A2(n728), .S0(n480), .Y(n633) );
  IBUFFX2_HVT U127 ( .A(n377), .Y(n369) );
  INVX1_HVT U128 ( .A(in[3]), .Y(n351) );
  INVX1_HVT U129 ( .A(n375), .Y(n372) );
  IBUFFX2_HVT U130 ( .A(n502), .Y(n353) );
  INVX1_HVT U131 ( .A(n504), .Y(n473) );
  NAND2X0_HVT U132 ( .A1(n644), .A2(n485), .Y(n204) );
  NAND2X0_HVT U133 ( .A1(n127), .A2(n204), .Y(n642) );
  AO21X1_HVT U134 ( .A1(n481), .A2(n426), .A3(n332), .Y(n643) );
  INVX0_HVT U137 ( .A(n473), .Y(n368) );
  INVX1_HVT U138 ( .A(n536), .Y(n210) );
  INVX1_HVT U139 ( .A(n210), .Y(n211) );
  MUX41X1_HVT U141 ( .A1(n409), .A3(n697), .A2(n519), .A4(n520), .S0(n307), 
        .S1(n462), .Y(n696) );
  INVX1_HVT U142 ( .A(n509), .Y(n275) );
  MUX41X1_HVT U143 ( .A1(n629), .A3(n634), .A2(n641), .A4(n647), .S0(n488), 
        .S1(n326), .Y(out[3]) );
  NAND2X0_HVT U144 ( .A1(n456), .A2(n218), .Y(n212) );
  NAND2X0_HVT U145 ( .A1(n375), .A2(n385), .Y(n213) );
  INVX0_HVT U146 ( .A(n496), .Y(n456) );
  INVX0_HVT U147 ( .A(n420), .Y(n375) );
  MUX21X1_HVT U148 ( .A1(n545), .A2(n375), .S0(n218), .Y(n750) );
  MUX41X1_HVT U149 ( .A1(n735), .A3(n332), .A2(n648), .A4(n427), .S0(n379), 
        .S1(n462), .Y(n376) );
  INVX1_HVT U150 ( .A(in[1]), .Y(n377) );
  INVX0_HVT U151 ( .A(n377), .Y(n441) );
  INVX0_HVT U152 ( .A(n333), .Y(n216) );
  MUX41X1_HVT U155 ( .A1(n513), .A3(n271), .A2(n726), .A4(n746), .S0(n384), 
        .S1(n507), .Y(n563) );
  MUX41X1_HVT U156 ( .A1(n524), .A3(n744), .A2(n304), .A4(n589), .S0(n462), 
        .S1(n334), .Y(n588) );
  NAND2X0_HVT U157 ( .A1(n363), .A2(n364), .Y(n217) );
  MUX21X1_HVT U160 ( .A1(n531), .A2(n410), .S0(n431), .Y(n589) );
  NAND2X0_HVT U161 ( .A1(n475), .A2(n218), .Y(n219) );
  NAND2X0_HVT U163 ( .A1(n408), .A2(n438), .Y(n222) );
  NAND2X0_HVT U164 ( .A1(n219), .A2(n222), .Y(n738) );
  INVX0_HVT U169 ( .A(n438), .Y(n218) );
  MUX41X1_HVT U170 ( .A1(n623), .A3(n625), .A2(n626), .A4(n627), .S0(n482), 
        .S1(n488), .Y(n622) );
  INVX1_HVT U171 ( .A(n721), .Y(n528) );
  MUX41X1_HVT U173 ( .A1(n584), .A3(n585), .A2(n586), .A4(n588), .S0(n505), 
        .S1(n487), .Y(n583) );
  INVX1_HVT U174 ( .A(n377), .Y(n502) );
  INVX0_HVT U175 ( .A(n718), .Y(n517) );
  INVX0_HVT U176 ( .A(n726), .Y(n224) );
  MUX41X1_HVT U181 ( .A1(n672), .A3(n676), .A2(n674), .A4(n677), .S0(n488), 
        .S1(n482), .Y(n671) );
  OR2X1_HVT U182 ( .A1(n227), .A2(n379), .Y(n417) );
  NAND2X0_HVT U183 ( .A1(n231), .A2(n528), .Y(n227) );
  NAND2X0_HVT U184 ( .A1(n522), .A2(n229), .Y(n231) );
  MUX21X1_HVT U185 ( .A1(n408), .A2(n399), .S0(n430), .Y(n232) );
  INVX1_HVT U187 ( .A(n342), .Y(n304) );
  INVX1_HVT U188 ( .A(n443), .Y(n439) );
  NAND2X0_HVT U191 ( .A1(n423), .A2(n501), .Y(n238) );
  NAND2X0_HVT U192 ( .A1(n420), .A2(n323), .Y(n241) );
  INVX1_HVT U193 ( .A(n496), .Y(n531) );
  INVX1_HVT U194 ( .A(n420), .Y(n421) );
  NAND2X0_HVT U195 ( .A1(n318), .A2(n210), .Y(n242) );
  MUX41X1_HVT U196 ( .A1(n471), .A3(n701), .A2(n469), .A4(n289), .S0(n245), 
        .S1(n483), .Y(n700) );
  NAND2X0_HVT U198 ( .A1(n369), .A2(n751), .Y(n252) );
  NAND2X0_HVT U199 ( .A1(n246), .A2(n451), .Y(n253) );
  INVX0_HVT U200 ( .A(n751), .Y(n246) );
  MUX21X1_HVT U201 ( .A1(n531), .A2(n246), .S0(n353), .Y(n663) );
  MUX41X1_HVT U202 ( .A1(n682), .A3(n685), .A2(n684), .A4(n689), .S0(n487), 
        .S1(n506), .Y(n681) );
  INVX1_HVT U203 ( .A(n410), .Y(n257) );
  MUX41X1_HVT U204 ( .A1(n711), .A3(n573), .A2(n717), .A4(n723), .S0(n379), 
        .S1(n457), .Y(n572) );
  OR2X1_HVT U205 ( .A1(n406), .A2(n501), .Y(n723) );
  NBUFFX2_HVT U206 ( .A(n745), .Y(n329) );
  INVX1_HVT U207 ( .A(n730), .Y(n539) );
  MUX21X1_HVT U209 ( .A1(n331), .A2(n456), .S0(n430), .Y(n330) );
  INVX0_HVT U210 ( .A(n489), .Y(n258) );
  MUX21X1_HVT U211 ( .A1(n495), .A2(n498), .S0(n459), .Y(n552) );
  OA21X1_HVT U213 ( .A1(n469), .A2(n432), .A3(n727), .Y(n592) );
  NAND2X0_HVT U216 ( .A1(n569), .A2(n416), .Y(n259) );
  NAND2X0_HVT U217 ( .A1(n568), .A2(n379), .Y(n261) );
  NAND2X0_HVT U219 ( .A1(n259), .A2(n261), .Y(n567) );
  MUX41X1_HVT U221 ( .A1(n401), .A3(n542), .A2(n410), .A4(n543), .S0(n275), 
        .S1(n334), .Y(n684) );
  NAND2X0_HVT U222 ( .A1(n453), .A2(n438), .Y(n263) );
  NAND2X0_HVT U223 ( .A1(n430), .A2(n751), .Y(n264) );
  NAND2X0_HVT U224 ( .A1(n263), .A2(n264), .Y(n452) );
  INVX1_HVT U225 ( .A(n546), .Y(n270) );
  INVX1_HVT U226 ( .A(n686), .Y(n546) );
  NAND2X0_HVT U227 ( .A1(n439), .A2(n242), .Y(n686) );
  NAND2X0_HVT U228 ( .A1(n354), .A2(n355), .Y(n271) );
  INVX1_HVT U229 ( .A(n552), .Y(n515) );
  NAND2X0_HVT U230 ( .A1(n224), .A2(n481), .Y(n273) );
  NAND2X0_HVT U231 ( .A1(n740), .A2(n334), .Y(n274) );
  NAND2X0_HVT U232 ( .A1(n273), .A2(n274), .Y(n630) );
  INVX0_HVT U233 ( .A(n452), .Y(n741) );
  MUX41X1_HVT U234 ( .A1(n694), .A3(n692), .A2(n693), .A4(n522), .S0(n396), 
        .S1(n275), .Y(n691) );
  INVX1_HVT U235 ( .A(n330), .Y(n746) );
  NAND2X0_HVT U236 ( .A1(n532), .A2(n461), .Y(n278) );
  NAND2X0_HVT U237 ( .A1(n275), .A2(n721), .Y(n279) );
  NAND2X0_HVT U238 ( .A1(n278), .A2(n279), .Y(n606) );
  MUX21X1_HVT U239 ( .A1(n545), .A2(n531), .S0(n362), .Y(n721) );
  MUX21X1_HVT U240 ( .A1(n271), .A2(n397), .S0(n335), .Y(n280) );
  INVX0_HVT U243 ( .A(n748), .Y(n424) );
  MUX21X1_HVT U244 ( .A1(n428), .A2(n246), .S0(n434), .Y(n652) );
  MUX21X1_HVT U246 ( .A1(n492), .A2(n531), .S0(n440), .Y(n729) );
  NAND2X0_HVT U247 ( .A1(n617), .A2(n379), .Y(n282) );
  NAND2X0_HVT U248 ( .A1(n618), .A2(n396), .Y(n283) );
  NAND2X0_HVT U249 ( .A1(n282), .A2(n283), .Y(n616) );
  INVX0_HVT U250 ( .A(n665), .Y(n532) );
  INVX1_HVT U253 ( .A(n376), .Y(n619) );
  INVX0_HVT U254 ( .A(n470), .Y(n310) );
  MUX41X1_HVT U255 ( .A1(n691), .A3(n699), .A2(n695), .A4(n705), .S0(n326), 
        .S1(n487), .Y(out[0]) );
  INVX1_HVT U257 ( .A(n757), .Y(n545) );
  NAND2X0_HVT U258 ( .A1(n23), .A2(n340), .Y(n285) );
  NAND2X0_HVT U259 ( .A1(n285), .A2(n289), .Y(n478) );
  MUX41X1_HVT U260 ( .A1(n328), .A3(n258), .A2(n23), .A4(n500), .S0(n396), 
        .S1(n507), .Y(n570) );
  NAND2X0_HVT U261 ( .A1(n408), .A2(n293), .Y(n296) );
  NAND2X0_HVT U262 ( .A1(n500), .A2(n451), .Y(n297) );
  NAND2X0_HVT U263 ( .A1(n296), .A2(n297), .Y(n327) );
  MUX21X1_HVT U265 ( .A1(n535), .A2(n327), .S0(n472), .Y(n644) );
  INVX1_HVT U266 ( .A(n556), .Y(n525) );
  NAND2X0_HVT U267 ( .A1(n727), .A2(n334), .Y(n300) );
  NAND2X0_HVT U269 ( .A1(n649), .A2(n480), .Y(n303) );
  MUX41X1_HVT U270 ( .A1(n600), .A3(n540), .A2(n601), .A4(n465), .S0(n384), 
        .S1(n507), .Y(n599) );
  XNOR2X2_HVT U271 ( .A1(n381), .A2(n369), .Y(n465) );
  INVX1_HVT U272 ( .A(n401), .Y(n733) );
  NAND2X0_HVT U273 ( .A1(n706), .A2(n334), .Y(n305) );
  NAND2X0_HVT U274 ( .A1(n710), .A2(n480), .Y(n306) );
  NAND2X0_HVT U275 ( .A1(n305), .A2(n306), .Y(n705) );
  INVX1_HVT U276 ( .A(n322), .Y(n688) );
  INVX0_HVT U277 ( .A(n341), .Y(n732) );
  MUX41X1_HVT U278 ( .A1(n474), .A3(n47), .A2(n280), .A4(n478), .S0(n390), 
        .S1(n505), .Y(n477) );
  MUX41X1_HVT U279 ( .A1(n651), .A3(n653), .A2(n654), .A4(n658), .S0(n482), 
        .S1(n488), .Y(n650) );
  MUX41X1_HVT U280 ( .A1(n652), .A3(n539), .A2(n533), .A4(n712), .S0(n275), 
        .S1(n319), .Y(n651) );
  MUX21X1_HVT U281 ( .A1(n399), .A2(n378), .S0(n440), .Y(n737) );
  NAND2X0_HVT U282 ( .A1(n331), .A2(n307), .Y(n308) );
  NAND2X0_HVT U283 ( .A1(n723), .A2(n506), .Y(n309) );
  NAND2X0_HVT U285 ( .A1(n308), .A2(n309), .Y(n709) );
  INVX0_HVT U286 ( .A(n506), .Y(n307) );
  INVX0_HVT U287 ( .A(n494), .Y(n331) );
  MUX21X1_HVT U288 ( .A1(n708), .A2(n709), .S0(n484), .Y(n706) );
  NAND2X0_HVT U290 ( .A1(n608), .A2(n310), .Y(n311) );
  NAND2X0_HVT U291 ( .A1(n257), .A2(n470), .Y(n312) );
  NAND2X0_HVT U292 ( .A1(n311), .A2(n312), .Y(n607) );
  MUX41X1_HVT U293 ( .A1(n216), .A3(n529), .A2(n341), .A4(n517), .S0(n457), 
        .S1(n473), .Y(n582) );
  NAND2X0_HVT U294 ( .A1(n371), .A2(n370), .Y(n313) );
  MUX21X1_HVT U296 ( .A1(n460), .A2(n378), .S0(n431), .Y(n401) );
  NAND2X0_HVT U297 ( .A1(n628), .A2(n379), .Y(n314) );
  NAND2X0_HVT U298 ( .A1(n511), .A2(n368), .Y(n315) );
  NAND2X0_HVT U299 ( .A1(n314), .A2(n315), .Y(n627) );
  MUX41X1_HVT U300 ( .A1(n605), .A3(n603), .A2(n610), .A4(n609), .S0(n307), 
        .S1(n487), .Y(n602) );
  NAND2X0_HVT U301 ( .A1(n423), .A2(n245), .Y(n316) );
  NAND2X0_HVT U303 ( .A1(n217), .A2(n275), .Y(n317) );
  NAND2X0_HVT U304 ( .A1(n316), .A2(n317), .Y(n613) );
  MUX21X1_HVT U305 ( .A1(n545), .A2(n375), .S0(n433), .Y(n601) );
  NAND2X0_HVT U308 ( .A1(n590), .A2(n365), .Y(n366) );
  MUX21X1_HVT U310 ( .A1(n593), .A2(n592), .S0(n480), .Y(n591) );
  MUX21X2_HVT U311 ( .A1(n453), .A2(n425), .S0(n459), .Y(n328) );
  INVX0_HVT U312 ( .A(n351), .Y(n318) );
  INVX1_HVT U313 ( .A(n458), .Y(n744) );
  INVX0_HVT U314 ( .A(n740), .Y(n540) );
  MUX41X1_HVT U315 ( .A1(n661), .A3(n662), .A2(n664), .A4(n669), .S0(n482), 
        .S1(n487), .Y(n660) );
  AO21X1_HVT U316 ( .A1(n486), .A2(n665), .A3(n541), .Y(n666) );
  INVX1_HVT U317 ( .A(n427), .Y(n428) );
  INVX0_HVT U318 ( .A(n246), .Y(n332) );
  MUX41X1_HVT U319 ( .A1(n466), .A3(n550), .A2(n663), .A4(n328), .S0(n396), 
        .S1(n245), .Y(n662) );
  INVX0_HVT U320 ( .A(n327), .Y(n724) );
  NAND2X0_HVT U321 ( .A1(n489), .A2(n395), .Y(n320) );
  NAND2X0_HVT U322 ( .A1(n492), .A2(n434), .Y(n321) );
  NAND2X0_HVT U323 ( .A1(n320), .A2(n321), .Y(n655) );
  MUX41X1_HVT U324 ( .A1(n433), .A3(n742), .A2(n543), .A4(n466), .S0(n340), 
        .S1(n275), .Y(n661) );
  INVX0_HVT U325 ( .A(n493), .Y(n453) );
  MUX21X1_HVT U326 ( .A1(n741), .A2(n463), .S0(n484), .Y(n565) );
  MUX21X1_HVT U327 ( .A1(n427), .A2(n342), .S0(n362), .Y(n322) );
  NAND2X0_HVT U328 ( .A1(n378), .A2(n323), .Y(n324) );
  NAND2X0_HVT U329 ( .A1(n426), .A2(n293), .Y(n325) );
  NAND2X0_HVT U330 ( .A1(n324), .A2(n325), .Y(n743) );
  MUX41X1_HVT U331 ( .A1(n468), .A3(n464), .A2(n542), .A4(n673), .S0(n319), 
        .S1(n457), .Y(n672) );
  INVX1_HVT U332 ( .A(n555), .Y(n542) );
  INVX1_HVT U333 ( .A(n365), .Y(n326) );
  INVX0_HVT U334 ( .A(in[6]), .Y(n365) );
  NAND2X0_HVT U335 ( .A1(n671), .A2(n365), .Y(n444) );
  NAND2X0_HVT U336 ( .A1(n389), .A2(n388), .Y(out[6]) );
  NAND2X0_HVT U337 ( .A1(n347), .A2(n346), .Y(out[2]) );
  INVX0_HVT U338 ( .A(in[1]), .Y(n443) );
  MUX41X1_HVT U339 ( .A1(n50), .A3(n543), .A2(n270), .A4(n515), .S0(n396), 
        .S1(n412), .Y(n615) );
  INVX1_HVT U340 ( .A(n425), .Y(n426) );
  MUX21X1_HVT U341 ( .A1(n304), .A2(n494), .S0(n416), .Y(n380) );
  INVX0_HVT U342 ( .A(n443), .Y(n431) );
  INVX0_HVT U343 ( .A(n339), .Y(n749) );
  INVX0_HVT U344 ( .A(n495), .Y(n333) );
  NAND2X0_HVT U345 ( .A1(n442), .A2(n335), .Y(n336) );
  NAND2X0_HVT U346 ( .A1(n755), .A2(n338), .Y(n337) );
  NAND2X0_HVT U347 ( .A1(n336), .A2(n337), .Y(n637) );
  INVX1_HVT U348 ( .A(n479), .Y(n338) );
  MUX41X1_HVT U349 ( .A1(n631), .A3(n633), .A2(n630), .A4(n632), .S0(n482), 
        .S1(n275), .Y(n629) );
  AND2X1_HVT U350 ( .A1(n356), .A2(n357), .Y(n339) );
  NAND2X0_HVT U351 ( .A1(n467), .A2(n343), .Y(n344) );
  NAND2X0_HVT U352 ( .A1(n659), .A2(n713), .Y(n345) );
  NAND2X0_HVT U353 ( .A1(n344), .A2(n345), .Y(n658) );
  INVX0_HVT U354 ( .A(n713), .Y(n343) );
  NAND2X0_HVT U355 ( .A1(n650), .A2(n365), .Y(n346) );
  NAND2X0_HVT U356 ( .A1(n660), .A2(n326), .Y(n347) );
  MUX21X1_HVT U357 ( .A1(n544), .A2(n743), .S0(n481), .Y(n659) );
  XOR2X1_HVT U358 ( .A1(n473), .A2(n508), .Y(n713) );
  NAND2X0_HVT U359 ( .A1(n666), .A2(n368), .Y(n348) );
  NAND2X0_HVT U360 ( .A1(n667), .A2(n481), .Y(n349) );
  NAND2X0_HVT U361 ( .A1(n348), .A2(n349), .Y(n664) );
  MUX41X1_HVT U362 ( .A1(n516), .A3(n113), .A2(n670), .A4(n717), .S0(n412), 
        .S1(n340), .Y(n669) );
  INVX0_HVT U363 ( .A(n460), .Y(n751) );
  INVX1_HVT U364 ( .A(n411), .Y(n628) );
  INVX0_HVT U365 ( .A(n510), .Y(n509) );
  NBUFFX2_HVT U366 ( .A(n509), .Y(n486) );
  NBUFFX2_HVT U367 ( .A(n509), .Y(n484) );
  INVX1_HVT U368 ( .A(n502), .Y(n442) );
  INVX0_HVT U369 ( .A(n350), .Y(n640) );
  MUX21X1_HVT U370 ( .A1(n725), .A2(n232), .S0(n335), .Y(n350) );
  INVX0_HVT U371 ( .A(n502), .Y(n451) );
  NAND2X0_HVT U372 ( .A1(n406), .A2(n353), .Y(n354) );
  NAND2X0_HVT U373 ( .A1(n545), .A2(n119), .Y(n355) );
  NAND2X0_HVT U374 ( .A1(n354), .A2(n355), .Y(n722) );
  INVX0_HVT U375 ( .A(n500), .Y(n435) );
  MUX21X1_HVT U376 ( .A1(n549), .A2(n419), .S0(n485), .Y(n569) );
  OR2X1_HVT U377 ( .A1(n118), .A2(n458), .Y(n745) );
  NAND2X0_HVT U378 ( .A1(n495), .A2(n323), .Y(n356) );
  NAND2X0_HVT U379 ( .A1(n331), .A2(n440), .Y(n357) );
  MUX21X1_HVT U380 ( .A1(n427), .A2(n333), .S0(n434), .Y(n739) );
  INVX0_HVT U381 ( .A(n553), .Y(n530) );
  INVX1_HVT U382 ( .A(n377), .Y(n440) );
  INVX0_HVT U383 ( .A(n473), .Y(n384) );
  INVX1_HVT U384 ( .A(n476), .Y(n413) );
  NAND2X0_HVT U385 ( .A1(n754), .A2(n319), .Y(n358) );
  NAND2X0_HVT U386 ( .A1(n624), .A2(n396), .Y(n359) );
  NAND2X0_HVT U387 ( .A1(n359), .A2(n358), .Y(n623) );
  NAND2X0_HVT U388 ( .A1(n453), .A2(n323), .Y(n360) );
  NAND2X0_HVT U389 ( .A1(n531), .A2(n440), .Y(n361) );
  NAND2X0_HVT U390 ( .A1(n360), .A2(n361), .Y(n720) );
  INVX1_HVT U391 ( .A(n481), .Y(n396) );
  INVX0_HVT U392 ( .A(n720), .Y(n529) );
  NAND2X0_HVT U393 ( .A1(n246), .A2(n362), .Y(n363) );
  NAND2X0_HVT U394 ( .A1(n318), .A2(n449), .Y(n364) );
  NAND2X0_HVT U395 ( .A1(n363), .A2(n364), .Y(n448) );
  NAND2X0_HVT U396 ( .A1(n602), .A2(n326), .Y(n367) );
  NAND2X0_HVT U397 ( .A1(n367), .A2(n366), .Y(out[5]) );
  INVX0_HVT U398 ( .A(n119), .Y(n449) );
  INVX1_HVT U399 ( .A(n424), .Y(n400) );
  INVX1_HVT U400 ( .A(n486), .Y(n450) );
  MUX41X1_HVT U401 ( .A1(n732), .A3(n688), .A2(n734), .A4(n687), .S0(n368), 
        .S1(n507), .Y(n685) );
  NAND2X0_HVT U402 ( .A1(n446), .A2(n447), .Y(out[4]) );
  NBUFFX2_HVT U403 ( .A(in[5]), .Y(n506) );
  NAND2X0_HVT U404 ( .A1(n545), .A2(n119), .Y(n370) );
  NAND2X0_HVT U405 ( .A1(n410), .A2(n218), .Y(n371) );
  NAND2X0_HVT U406 ( .A1(n370), .A2(n371), .Y(n731) );
  NAND2X0_HVT U407 ( .A1(n679), .A2(n379), .Y(n373) );
  NAND2X0_HVT U408 ( .A1(n680), .A2(n396), .Y(n374) );
  NAND2X0_HVT U409 ( .A1(n374), .A2(n373), .Y(n677) );
  INVX0_HVT U410 ( .A(n492), .Y(n406) );
  NAND2X0_HVT U411 ( .A1(n318), .A2(n492), .Y(n378) );
  NAND2X0_HVT U412 ( .A1(n690), .A2(n379), .Y(n382) );
  NAND2X0_HVT U413 ( .A1(n715), .A2(n368), .Y(n383) );
  NAND2X0_HVT U414 ( .A1(n382), .A2(n383), .Y(n689) );
  MUX41X1_HVT U415 ( .A1(n718), .A3(n38), .A2(n313), .A4(n428), .S0(n473), 
        .S1(n484), .Y(n571) );
  INVX1_HVT U416 ( .A(n490), .Y(n399) );
  MUX41X1_HVT U417 ( .A1(n544), .A3(n537), .A2(n755), .A4(n406), .S0(n384), 
        .S1(n432), .Y(n561) );
  NAND2X0_HVT U418 ( .A1(n304), .A2(n385), .Y(n386) );
  NAND2X0_HVT U419 ( .A1(n258), .A2(n395), .Y(n387) );
  NAND2X0_HVT U420 ( .A1(n386), .A2(n387), .Y(n683) );
  NAND2X0_HVT U421 ( .A1(n574), .A2(n365), .Y(n388) );
  NAND2X0_HVT U422 ( .A1(n583), .A2(n326), .Y(n389) );
  MUX41X1_HVT U423 ( .A1(n616), .A3(n615), .A2(n620), .A4(n619), .S0(n307), 
        .S1(n488), .Y(n614) );
  NAND2X0_HVT U424 ( .A1(n390), .A2(n397), .Y(n391) );
  NAND2X0_HVT U425 ( .A1(n729), .A2(n450), .Y(n392) );
  NAND2X0_HVT U426 ( .A1(n391), .A2(n392), .Y(n618) );
  NAND2X0_HVT U427 ( .A1(n700), .A2(n396), .Y(n393) );
  NAND2X0_HVT U428 ( .A1(n702), .A2(n379), .Y(n394) );
  NAND2X0_HVT U429 ( .A1(n394), .A2(n393), .Y(n699) );
  INVX1_HVT U430 ( .A(n398), .Y(n419) );
  OA21X1_HVT U431 ( .A1(n724), .A2(n432), .A3(n523), .Y(n580) );
  AND2X1_HVT U432 ( .A1(n369), .A2(n378), .Y(n397) );
  NAND2X0_HVT U433 ( .A1(n403), .A2(n402), .Y(out[7]) );
  MUX21X1_HVT U434 ( .A1(n399), .A2(n400), .S0(n439), .Y(n398) );
  NAND2X0_HVT U435 ( .A1(n560), .A2(n365), .Y(n402) );
  NAND2X0_HVT U436 ( .A1(n566), .A2(n326), .Y(n403) );
  MUX41X1_HVT U437 ( .A1(n733), .A3(n621), .A2(n528), .A4(n429), .S0(n484), 
        .S1(n335), .Y(n620) );
  NAND2X0_HVT U438 ( .A1(n645), .A2(n482), .Y(n404) );
  NAND2X0_HVT U439 ( .A1(n642), .A2(n307), .Y(n405) );
  NAND2X0_HVT U440 ( .A1(n404), .A2(n405), .Y(n641) );
  XNOR2X2_HVT U441 ( .A1(n491), .A2(n352), .Y(n460) );
  INVX0_HVT U442 ( .A(n485), .Y(n412) );
  NBUFFX2_HVT U443 ( .A(n211), .Y(n490) );
  MUX21X1_HVT U444 ( .A1(n500), .A2(n408), .S0(n459), .Y(n407) );
  AND2X1_HVT U445 ( .A1(n744), .A2(n499), .Y(n409) );
  NAND2X0_HVT U446 ( .A1(n475), .A2(n413), .Y(n414) );
  NAND2X0_HVT U447 ( .A1(n380), .A2(n476), .Y(n415) );
  NAND2X0_HVT U448 ( .A1(n415), .A2(n414), .Y(n474) );
  NAND2X0_HVT U449 ( .A1(n565), .A2(n479), .Y(n418) );
  NAND2X0_HVT U450 ( .A1(n417), .A2(n418), .Y(n564) );
  INVX1_HVT U451 ( .A(n551), .Y(n537) );
  INVX1_HVT U452 ( .A(n554), .Y(n511) );
  NBUFFX2_HVT U453 ( .A(n748), .Y(n422) );
  INVX1_HVT U454 ( .A(n422), .Y(n425) );
  INVX1_HVT U455 ( .A(n508), .Y(n432) );
  XNOR2X1_HVT U456 ( .A1(n435), .A2(n442), .Y(n468) );
  NAND2X0_HVT U457 ( .A1(n698), .A2(n319), .Y(n436) );
  NAND2X0_HVT U458 ( .A1(n696), .A2(n396), .Y(n437) );
  NAND2X0_HVT U459 ( .A1(n437), .A2(n436), .Y(n695) );
  INVX0_HVT U460 ( .A(n443), .Y(n501) );
  NAND2X0_HVT U461 ( .A1(n681), .A2(n326), .Y(n445) );
  NAND2X0_HVT U462 ( .A1(n444), .A2(n445), .Y(out[1]) );
  NAND2X0_HVT U463 ( .A1(n622), .A2(n326), .Y(n446) );
  NAND2X0_HVT U464 ( .A1(n614), .A2(n365), .Y(n447) );
  NAND2X0_HVT U465 ( .A1(n635), .A2(n307), .Y(n454) );
  NAND2X0_HVT U466 ( .A1(n636), .A2(n482), .Y(n455) );
  NAND2X0_HVT U467 ( .A1(n454), .A2(n455), .Y(n634) );
  NBUFFX2_HVT U468 ( .A(n421), .Y(n489) );
  MUX41X1_HVT U469 ( .A1(n401), .A3(n727), .A2(n745), .A4(n646), .S0(n472), 
        .S1(n457), .Y(n645) );
  NBUFFX2_HVT U470 ( .A(n508), .Y(n461) );
  NBUFFX2_HVT U471 ( .A(n508), .Y(n462) );
  AND2X1_HVT U472 ( .A1(n236), .A2(n703), .Y(n463) );
  NBUFFX2_HVT U473 ( .A(n753), .Y(n495) );
  MUX21X1_HVT U474 ( .A1(n333), .A2(n545), .S0(n506), .Y(n707) );
  NBUFFX2_HVT U475 ( .A(n753), .Y(n496) );
  AND2X1_HVT U476 ( .A1(n257), .A2(n686), .Y(n464) );
  MUX21X1_HVT U477 ( .A1(n494), .A2(n475), .S0(n119), .Y(n719) );
  NAND2X0_HVT U478 ( .A1(n491), .A2(n548), .Y(n753) );
  MUX21X1_HVT U479 ( .A1(n531), .A2(n304), .S0(n369), .Y(n553) );
  NBUFFX2_HVT U480 ( .A(n756), .Y(n497) );
  NBUFFX2_HVT U481 ( .A(n756), .Y(n498) );
  MUX21X1_HVT U482 ( .A1(n493), .A2(n304), .S0(n439), .Y(n573) );
  MUX21X1_HVT U483 ( .A1(n493), .A2(n500), .S0(n440), .Y(n576) );
  MUX21X1_HVT U484 ( .A1(n500), .A2(n497), .S0(n439), .Y(n577) );
  MUX21X1_HVT U485 ( .A1(n381), .A2(n500), .S0(n293), .Y(n665) );
  MUX21X1_HVT U486 ( .A1(n497), .A2(n492), .S0(n440), .Y(n557) );
  AND2X1_HVT U487 ( .A1(n431), .A2(n410), .Y(n466) );
  AND2X1_HVT U488 ( .A1(n499), .A2(n648), .Y(n467) );
  MUX21X1_HVT U489 ( .A1(n428), .A2(n500), .S0(n480), .Y(n638) );
  NBUFFX2_HVT U490 ( .A(n548), .Y(n493) );
  NBUFFX2_HVT U491 ( .A(n548), .Y(n494) );
  NBUFFX2_HVT U492 ( .A(n509), .Y(n485) );
  NBUFFX2_HVT U493 ( .A(n503), .Y(n480) );
  NBUFFX2_HVT U494 ( .A(n503), .Y(n481) );
  NBUFFX2_HVT U495 ( .A(n503), .Y(n479) );
  NBUFFX2_HVT U496 ( .A(n505), .Y(n483) );
  NBUFFX2_HVT U497 ( .A(n505), .Y(n482) );
  MUX21X1_HVT U498 ( .A1(n580), .A2(n581), .S0(n479), .Y(n579) );
  MUX21X1_HVT U499 ( .A1(n673), .A2(n331), .S0(n485), .Y(n581) );
  MUX21X1_HVT U500 ( .A1(n426), .A2(n328), .S0(n486), .Y(n593) );
  AND2X1_HVT U501 ( .A1(n489), .A2(n451), .Y(n469) );
  MUX21X1_HVT U502 ( .A1(n427), .A2(n475), .S0(n369), .Y(n598) );
  NAND2X0_HVT U503 ( .A1(n318), .A2(n491), .Y(n756) );
  XOR2X1_HVT U504 ( .A1(n438), .A2(n505), .Y(n716) );
  MUX21X1_HVT U505 ( .A1(n408), .A2(n427), .S0(n119), .Y(n555) );
  MUX21X1_HVT U506 ( .A1(n728), .A2(n558), .S0(n484), .Y(n554) );
  MUX21X1_HVT U507 ( .A1(n453), .A2(n304), .S0(n486), .Y(n668) );
  NBUFFX2_HVT U508 ( .A(n757), .Y(n500) );
  NBUFFX2_HVT U509 ( .A(n242), .Y(n499) );
  AND2X1_HVT U510 ( .A1(n494), .A2(n353), .Y(n471) );
  NBUFFX2_HVT U511 ( .A(in[5]), .Y(n505) );
  NAND2X0_HVT U512 ( .A1(n210), .A2(n352), .Y(n757) );
  MUX21X1_HVT U513 ( .A1(n399), .A2(n372), .S0(n431), .Y(n556) );
  NAND2X0_HVT U514 ( .A1(n210), .A2(n548), .Y(n748) );
  MUX21X1_HVT U515 ( .A1(n242), .A2(n406), .S0(n438), .Y(n730) );
  MUX21X1_HVT U516 ( .A1(n406), .A2(n499), .S0(n438), .Y(n551) );
  NBUFFX2_HVT U517 ( .A(in[0]), .Y(n487) );
  NBUFFX2_HVT U518 ( .A(in[0]), .Y(n488) );
endmodule

