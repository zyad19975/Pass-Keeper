
module sbox_2 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n12, n15, n19, n23, n32, n37, n50, n118, n119, n204, n210, n211, n212,
         n213, n216, n217, n218, n219, n227, n231, n232, n236, n238, n242,
         n243, n249, n252, n256, n259, n261, n264, n268, n272, n273, n279,
         n280, n282, n283, n286, n290, n291, n293, n296, n297, n301, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789;

  NAND2X0_HVT U4 ( .A1(n513), .A2(n787), .Y(n786) );
  NAND2X0_HVT U5 ( .A1(n521), .A2(n511), .Y(n784) );
  NAND2X0_HVT U13 ( .A1(n777), .A2(n312), .Y(n778) );
  NAND2X0_HVT U15 ( .A1(n787), .A2(n356), .Y(n776) );
  NAND2X0_HVT U21 ( .A1(n513), .A2(n523), .Y(n771) );
  NAND2X0_HVT U24 ( .A1(n324), .A2(n523), .Y(n769) );
  NAND2X0_HVT U33 ( .A1(n346), .A2(n523), .Y(n761) );
  MUX41X1_HVT U51 ( .A1(n538), .A3(n559), .A2(n454), .A4(n405), .S0(n484), 
        .S1(n528), .Y(n745) );
  NAND2X0_HVT U53 ( .A1(n742), .A2(n752), .Y(n743) );
  NAND2X0_HVT U56 ( .A1(n515), .A2(n738), .Y(n739) );
  MUX41X1_HVT U57 ( .A1(n547), .A3(n773), .A2(n739), .A4(n779), .S0(n531), 
        .S1(n527), .Y(n737) );
  NAND2X0_HVT U58 ( .A1(n517), .A2(n787), .Y(n736) );
  MUX41X1_HVT U61 ( .A1(n490), .A3(n441), .A2(n543), .A4(n462), .S0(n329), 
        .S1(n527), .Y(n733) );
  NAND2X0_HVT U62 ( .A1(n523), .A2(n232), .Y(n732) );
  AO21X1_HVT U66 ( .A1(n436), .A2(n505), .A3(n574), .Y(n728) );
  NAND2X0_HVT U73 ( .A1(n404), .A2(n297), .Y(n722) );
  MUX41X1_HVT U74 ( .A1(n723), .A3(n767), .A2(n722), .A4(n769), .S0(n500), 
        .S1(n484), .Y(n720) );
  AND2X1_HVT U83 ( .A1(n316), .A2(n342), .Y(n710) );
  MUX41X1_HVT U84 ( .A1(n544), .A3(n218), .A2(n351), .A4(n710), .S0(n264), 
        .S1(n529), .Y(n709) );
  NAND2X0_HVT U85 ( .A1(n523), .A2(n367), .Y(n708) );
  NAND2X0_HVT U101 ( .A1(n691), .A2(n690), .Y(n692) );
  MUX41X1_HVT U103 ( .A1(n357), .A3(n560), .A2(n442), .A4(n759), .S0(n470), 
        .S1(n473), .Y(n688) );
  MUX41X1_HVT U105 ( .A1(n566), .A3(n747), .A2(n687), .A4(n558), .S0(n377), 
        .S1(n529), .Y(n686) );
  NAND2X0_HVT U110 ( .A1(n417), .A2(n681), .Y(n682) );
  AND2X1_HVT U115 ( .A1(n336), .A2(n463), .Y(n678) );
  MUX41X1_HVT U116 ( .A1(n778), .A3(n678), .A2(n534), .A4(n212), .S0(n470), 
        .S1(n529), .Y(n677) );
  AND2X1_HVT U140 ( .A1(n512), .A2(n433), .Y(n652) );
  MUX41X1_HVT U153 ( .A1(n682), .A3(n490), .A2(n417), .A4(n341), .S0(n502), 
        .S1(n531), .Y(n640) );
  AND2X1_HVT U154 ( .A1(n486), .A2(n50), .Y(n639) );
  NAND2X0_HVT U158 ( .A1(n518), .A2(n367), .Y(n635) );
  MUX41X1_HVT U159 ( .A1(n211), .A3(n463), .A2(n635), .A4(n575), .S0(n498), 
        .S1(n529), .Y(n634) );
  AND2X1_HVT U162 ( .A1(n218), .A2(n19), .Y(n631) );
  NAND2X0_HVT U166 ( .A1(n312), .A2(n738), .Y(n627) );
  NAND2X0_HVT U167 ( .A1(n414), .A2(n523), .Y(n626) );
  MUX41X1_HVT U168 ( .A1(n547), .A3(n401), .A2(n626), .A4(n627), .S0(n498), 
        .S1(n368), .Y(n625) );
  NAND2X0_HVT U177 ( .A1(n316), .A2(n466), .Y(n618) );
  MUX41X1_HVT U178 ( .A1(n774), .A3(n618), .A2(n564), .A4(n757), .S0(n500), 
        .S1(n484), .Y(n617) );
  MUX41X1_HVT U180 ( .A1(n542), .A3(n781), .A2(n211), .A4(n487), .S0(n507), 
        .S1(n498), .Y(n615) );
  MUX41X1_HVT U182 ( .A1(n430), .A3(n515), .A2(n539), .A4(n561), .S0(n531), 
        .S1(n497), .Y(n613) );
  MUX41X1_HVT U189 ( .A1(n607), .A3(n777), .A2(n608), .A4(n558), .S0(n486), 
        .S1(n498), .Y(n606) );
  NAND2X0_HVT U208 ( .A1(n268), .A2(n514), .Y(n681) );
  NAND2X0_HVT U212 ( .A1(n440), .A2(n399), .Y(n738) );
  NAND2X0_HVT U214 ( .A1(n218), .A2(n523), .Y(n590) );
  NAND2X0_HVT U215 ( .A1(n681), .A2(n404), .Y(n589) );
  NAND2X0_HVT U218 ( .A1(n569), .A2(n256), .Y(n642) );
  NAND2X0_HVT U220 ( .A1(n486), .A2(n590), .Y(n713) );
  INVX0_HVT U241 ( .A(n769), .Y(n578) );
  INVX0_HVT U245 ( .A(n784), .Y(n575) );
  INVX0_HVT U256 ( .A(n642), .Y(n567) );
  INVX0_HVT U265 ( .A(n767), .Y(n561) );
  INVX0_HVT U268 ( .A(n771), .Y(n559) );
  INVX0_HVT U270 ( .A(n589), .Y(n558) );
  INVX0_HVT U278 ( .A(n761), .Y(n552) );
  INVX0_HVT U284 ( .A(n590), .Y(n548) );
  INVX0_HVT U289 ( .A(n690), .Y(n545) );
  INVX0_HVT U295 ( .A(n786), .Y(n542) );
  INVX0_HVT U296 ( .A(n776), .Y(n541) );
  INVX0_HVT U297 ( .A(n787), .Y(n540) );
  INVX0_HVT U306 ( .A(n626), .Y(n536) );
  MUX21X1_HVT U1 ( .A1(n312), .A2(n345), .S0(n321), .Y(n436) );
  NBUFFX2_HVT U2 ( .A(n335), .Y(n481) );
  MUX21X1_HVT U3 ( .A1(n415), .A2(n517), .S0(n339), .Y(n376) );
  INVX1_HVT U6 ( .A(n481), .Y(n380) );
  MUX21X1_HVT U7 ( .A1(n560), .A2(n400), .S0(n505), .Y(n727) );
  MUX21X1_HVT U8 ( .A1(n459), .A2(n340), .S0(n336), .Y(n718) );
  INVX1_HVT U9 ( .A(n481), .Y(n523) );
  INVX1_HVT U10 ( .A(n217), .Y(n231) );
  INVX1_HVT U11 ( .A(n758), .Y(n550) );
  INVX1_HVT U12 ( .A(n522), .Y(n518) );
  MUX21X1_HVT U14 ( .A1(n573), .A2(n463), .S0(n519), .Y(n632) );
  AND3X1_HVT U16 ( .A1(n500), .A2(n523), .A3(n485), .Y(n663) );
  MUX21X1_HVT U17 ( .A1(n643), .A2(n644), .S0(n377), .Y(n641) );
  MUX21X1_HVT U18 ( .A1(n546), .A2(n403), .S0(n507), .Y(n644) );
  INVX0_HVT U19 ( .A(n532), .Y(n530) );
  INVX0_HVT U20 ( .A(n439), .Y(n23) );
  MUX21X1_HVT U22 ( .A1(n462), .A2(n573), .S0(n518), .Y(n782) );
  AND2X1_HVT U23 ( .A1(n322), .A2(n323), .Y(n12) );
  AND2X1_HVT U25 ( .A1(n420), .A2(n419), .Y(n15) );
  NAND2X0_HVT U26 ( .A1(n268), .A2(n314), .Y(n19) );
  INVX1_HVT U27 ( .A(n327), .Y(n314) );
  INVX1_HVT U28 ( .A(n460), .Y(n462) );
  INVX1_HVT U29 ( .A(n458), .Y(n461) );
  NAND2X0_HVT U30 ( .A1(n466), .A2(n23), .Y(n32) );
  NAND2X0_HVT U31 ( .A1(n374), .A2(n439), .Y(n37) );
  NAND2X0_HVT U32 ( .A1(n32), .A2(n37), .Y(n405) );
  INVX1_HVT U34 ( .A(n389), .Y(n362) );
  INVX1_HVT U35 ( .A(n700), .Y(n556) );
  INVX1_HVT U36 ( .A(n789), .Y(n327) );
  MUX41X1_HVT U37 ( .A1(n578), .A3(n361), .A2(n750), .A4(n405), .S0(n502), 
        .S1(n317), .Y(n711) );
  INVX1_HVT U38 ( .A(in[1]), .Y(n433) );
  INVX1_HVT U39 ( .A(n518), .Y(n390) );
  INVX0_HVT U40 ( .A(n518), .Y(n413) );
  INVX0_HVT U41 ( .A(n789), .Y(n573) );
  INVX1_HVT U42 ( .A(n204), .Y(n210) );
  INVX1_HVT U43 ( .A(n338), .Y(n291) );
  NAND2X0_HVT U44 ( .A1(n283), .A2(n576), .Y(n118) );
  NAND2X0_HVT U45 ( .A1(n355), .A2(n50), .Y(n119) );
  NAND2X0_HVT U46 ( .A1(n118), .A2(n119), .Y(n783) );
  INVX0_HVT U47 ( .A(n576), .Y(n50) );
  INVX0_HVT U48 ( .A(n785), .Y(n204) );
  INVX1_HVT U49 ( .A(n344), .Y(n391) );
  MUX41X1_HVT U50 ( .A1(n718), .A3(n546), .A2(n781), .A4(n556), .S0(n282), 
        .S1(n526), .Y(n717) );
  AO21X1_HVT U52 ( .A1(n502), .A2(n404), .A3(n218), .Y(n675) );
  INVX1_HVT U54 ( .A(n763), .Y(n565) );
  NOR2X0_HVT U55 ( .A1(n342), .A2(n268), .Y(n341) );
  INVX1_HVT U59 ( .A(n330), .Y(n529) );
  INVX1_HVT U60 ( .A(n324), .Y(n375) );
  INVX1_HVT U63 ( .A(n501), .Y(n457) );
  MUX21X1_HVT U64 ( .A1(n460), .A2(n374), .S0(n520), .Y(n768) );
  INVX1_HVT U65 ( .A(n355), .Y(n283) );
  AND3X1_HVT U67 ( .A1(n232), .A2(n738), .A3(n713), .Y(n714) );
  MUX21X1_HVT U68 ( .A1(n401), .A2(n466), .S0(n336), .Y(n723) );
  MUX21X1_HVT U69 ( .A1(n344), .A2(n523), .S0(n505), .Y(n729) );
  MUX21X1_HVT U70 ( .A1(n12), .A2(n361), .S0(n502), .Y(n694) );
  MUX21X1_HVT U71 ( .A1(n515), .A2(n401), .S0(n521), .Y(n705) );
  INVX1_HVT U72 ( .A(n738), .Y(n571) );
  NAND2X0_HVT U75 ( .A1(n675), .A2(n383), .Y(n384) );
  MUX21X1_HVT U76 ( .A1(n556), .A2(n757), .S0(n272), .Y(n637) );
  MUX21X1_HVT U77 ( .A1(n624), .A2(n623), .S0(n377), .Y(n622) );
  XNOR2X1_HVT U78 ( .A1(n459), .A2(n321), .Y(n749) );
  INVX1_HVT U79 ( .A(n496), .Y(n498) );
  INVX1_HVT U80 ( .A(n532), .Y(n484) );
  INVX1_HVT U81 ( .A(n753), .Y(n577) );
  INVX1_HVT U82 ( .A(n530), .Y(n418) );
  INVX1_HVT U86 ( .A(in[7]), .Y(n532) );
  MUX21X1_HVT U87 ( .A1(n692), .A2(n533), .S0(n470), .Y(n689) );
  MUX21X1_HVT U88 ( .A1(n401), .A2(n356), .S0(n336), .Y(n687) );
  XOR2X1_HVT U89 ( .A1(n339), .A2(n324), .Y(n747) );
  MUX21X1_HVT U90 ( .A1(n611), .A2(n612), .S0(n377), .Y(n610) );
  MUX21X1_HVT U91 ( .A1(n708), .A2(n324), .S0(n473), .Y(n612) );
  INVX1_HVT U92 ( .A(n501), .Y(n443) );
  NBUFFX2_HVT U93 ( .A(in[5]), .Y(n527) );
  INVX1_HVT U94 ( .A(n506), .Y(n429) );
  INVX1_HVT U95 ( .A(n427), .Y(n282) );
  INVX0_HVT U96 ( .A(n506), .Y(n386) );
  INVX1_HVT U97 ( .A(n429), .Y(n368) );
  INVX1_HVT U98 ( .A(n484), .Y(n272) );
  NBUFFX2_HVT U99 ( .A(n524), .Y(n500) );
  INVX1_HVT U100 ( .A(n500), .Y(n304) );
  INVX1_HVT U102 ( .A(n506), .Y(n421) );
  INVX1_HVT U104 ( .A(n338), .Y(n268) );
  INVX0_HVT U106 ( .A(n330), .Y(n531) );
  INVX0_HVT U107 ( .A(n507), .Y(n383) );
  INVX1_HVT U108 ( .A(n338), .Y(n339) );
  INVX1_HVT U109 ( .A(n522), .Y(n521) );
  NBUFFX2_HVT U111 ( .A(n530), .Y(n506) );
  INVX1_HVT U112 ( .A(n335), .Y(n522) );
  INVX1_HVT U113 ( .A(n390), .Y(n256) );
  INVX0_HVT U114 ( .A(n516), .Y(n414) );
  NBUFFX2_HVT U117 ( .A(n528), .Y(n505) );
  INVX0_HVT U118 ( .A(n506), .Y(n427) );
  INVX1_HVT U119 ( .A(n380), .Y(n309) );
  INVX1_HVT U120 ( .A(n320), .Y(n315) );
  INVX1_HVT U121 ( .A(n503), .Y(n480) );
  INVX0_HVT U122 ( .A(n524), .Y(n496) );
  INVX1_HVT U123 ( .A(n337), .Y(n460) );
  INVX0_HVT U124 ( .A(n512), .Y(n569) );
  INVX0_HVT U125 ( .A(n486), .Y(n317) );
  INVX0_HVT U126 ( .A(n465), .Y(n342) );
  INVX1_HVT U127 ( .A(n573), .Y(n312) );
  NAND2X0_HVT U128 ( .A1(n777), .A2(n312), .Y(n211) );
  INVX1_HVT U129 ( .A(n768), .Y(n534) );
  INVX1_HVT U130 ( .A(n781), .Y(n560) );
  INVX1_HVT U131 ( .A(n782), .Y(n280) );
  XNOR2X2_HVT U132 ( .A1(n516), .A2(n413), .Y(n746) );
  INVX0_HVT U133 ( .A(n436), .Y(n779) );
  INVX0_HVT U134 ( .A(n517), .Y(n367) );
  MUX21X1_HVT U135 ( .A1(n463), .A2(n555), .S0(n309), .Y(n698) );
  MUX41X1_HVT U136 ( .A1(n680), .A3(n683), .A2(n15), .A4(n684), .S0(n504), 
        .S1(n427), .Y(n679) );
  INVX1_HVT U137 ( .A(n331), .Y(n313) );
  MUX41X1_HVT U138 ( .A1(n686), .A3(n689), .A2(n688), .A4(n693), .S0(in[0]), 
        .S1(n503), .Y(n685) );
  INVX0_HVT U139 ( .A(n12), .Y(n212) );
  INVX0_HVT U141 ( .A(n457), .Y(n264) );
  INVX1_HVT U142 ( .A(n460), .Y(n356) );
  INVX0_HVT U143 ( .A(n783), .Y(n458) );
  INVX0_HVT U144 ( .A(n757), .Y(n553) );
  NAND2X0_HVT U145 ( .A1(n415), .A2(n23), .Y(n213) );
  NAND2X0_HVT U146 ( .A1(n462), .A2(n313), .Y(n216) );
  NAND2X0_HVT U147 ( .A1(n213), .A2(n216), .Y(n754) );
  INVX1_HVT U148 ( .A(n754), .Y(n539) );
  MUX21X1_HVT U149 ( .A1(n517), .A2(n485), .S0(n380), .Y(n579) );
  MUX41X1_HVT U150 ( .A1(n342), .A3(n563), .A2(n357), .A4(n12), .S0(n282), 
        .S1(n524), .Y(n592) );
  NBUFFX2_HVT U151 ( .A(in[0]), .Y(n508) );
  INVX0_HVT U152 ( .A(in[3]), .Y(n389) );
  MUX21X1_HVT U155 ( .A1(n327), .A2(n342), .S0(n331), .Y(n217) );
  INVX0_HVT U156 ( .A(n433), .Y(n439) );
  NBUFFX2_HVT U157 ( .A(n461), .Y(n218) );
  NAND2X0_HVT U160 ( .A1(n714), .A2(n500), .Y(n219) );
  NAND2X0_HVT U161 ( .A1(n715), .A2(n457), .Y(n227) );
  NAND2X0_HVT U163 ( .A1(n219), .A2(n227), .Y(n712) );
  MUX41X1_HVT U164 ( .A1(n717), .A3(n719), .A2(n720), .A4(n724), .S0(n527), 
        .S1(n508), .Y(n716) );
  INVX0_HVT U165 ( .A(n783), .Y(n337) );
  INVX1_HVT U169 ( .A(n376), .Y(n766) );
  MUX21X1_HVT U170 ( .A1(n512), .A2(n772), .S0(n421), .Y(n715) );
  INVX0_HVT U171 ( .A(n414), .Y(n232) );
  XOR2X2_HVT U172 ( .A1(n316), .A2(n402), .Y(n750) );
  NAND2X0_HVT U173 ( .A1(n356), .A2(n23), .Y(n236) );
  NAND2X0_HVT U174 ( .A1(n431), .A2(n519), .Y(n238) );
  NAND2X0_HVT U175 ( .A1(n236), .A2(n238), .Y(n351) );
  NAND2X0_HVT U176 ( .A1(n280), .A2(n282), .Y(n242) );
  NAND2X0_HVT U179 ( .A1(n242), .A2(n243), .Y(n472) );
  AND2X1_HVT U181 ( .A1(n443), .A2(n553), .Y(n243) );
  MUX41X1_HVT U183 ( .A1(n592), .A3(n594), .A2(n593), .A4(n595), .S0(n508), 
        .S1(n503), .Y(n591) );
  MUX41X1_HVT U184 ( .A1(n651), .A3(n647), .A2(n650), .A4(n646), .S0(n476), 
        .S1(n480), .Y(n645) );
  MUX41X1_HVT U185 ( .A1(n753), .A3(n366), .A2(n705), .A4(n538), .S0(n452), 
        .S1(n531), .Y(n704) );
  MUX41X1_HVT U186 ( .A1(n628), .A3(n630), .A2(n622), .A4(n625), .S0(n503), 
        .S1(n388), .Y(n621) );
  NBUFFX2_HVT U187 ( .A(n562), .Y(n509) );
  MUX41X1_HVT U188 ( .A1(n641), .A3(n640), .A2(n636), .A4(n634), .S0(n480), 
        .S1(n388), .Y(n633) );
  INVX1_HVT U190 ( .A(n508), .Y(n388) );
  INVX1_HVT U191 ( .A(n522), .Y(n520) );
  NAND2X0_HVT U192 ( .A1(n430), .A2(n368), .Y(n249) );
  NAND2X0_HVT U193 ( .A1(n328), .A2(n317), .Y(n252) );
  NAND2X0_HVT U194 ( .A1(n249), .A2(n252), .Y(n655) );
  NAND2X0_HVT U195 ( .A1(n467), .A2(n256), .Y(n259) );
  NAND2X0_HVT U196 ( .A1(n337), .A2(n390), .Y(n261) );
  NAND2X0_HVT U197 ( .A1(n259), .A2(n261), .Y(n770) );
  MUX21X1_HVT U198 ( .A1(n431), .A2(n515), .S0(n439), .Y(n430) );
  INVX0_HVT U199 ( .A(n544), .Y(n328) );
  INVX0_HVT U200 ( .A(n770), .Y(n544) );
  OA21X1_HVT U201 ( .A1(n536), .A2(n427), .A3(n212), .Y(n648) );
  INVX1_HVT U202 ( .A(n588), .Y(n538) );
  MUX41X1_HVT U203 ( .A1(n489), .A3(n632), .A2(n441), .A4(n631), .S0(n264), 
        .S1(n330), .Y(n630) );
  INVX0_HVT U204 ( .A(n749), .Y(n365) );
  MUX21X1_HVT U205 ( .A1(n788), .A2(n431), .S0(n519), .Y(n454) );
  INVX1_HVT U206 ( .A(n430), .Y(n756) );
  MUX41X1_HVT U207 ( .A1(n734), .A3(n740), .A2(n726), .A4(n730), .S0(n508), 
        .S1(n424), .Y(out[0]) );
  INVX1_HVT U209 ( .A(n440), .Y(n338) );
  INVX1_HVT U210 ( .A(n522), .Y(n336) );
  MUX21X1_HVT U211 ( .A1(n540), .A2(n764), .S0(n386), .Y(n649) );
  INVX0_HVT U213 ( .A(n421), .Y(n455) );
  MUX41X1_HVT U216 ( .A1(n729), .A3(n727), .A2(n728), .A4(n280), .S0(n387), 
        .S1(n272), .Y(n726) );
  INVX1_HVT U217 ( .A(n520), .Y(n428) );
  NAND2X0_HVT U219 ( .A1(n741), .A2(n304), .Y(n273) );
  NAND2X0_HVT U221 ( .A1(n745), .A2(n264), .Y(n279) );
  NAND2X0_HVT U222 ( .A1(n279), .A2(n273), .Y(n740) );
  INVX1_HVT U223 ( .A(n405), .Y(n772) );
  INVX0_HVT U224 ( .A(n532), .Y(n329) );
  MUX41X1_HVT U225 ( .A1(n602), .A3(n598), .A2(n603), .A4(n601), .S0(n388), 
        .S1(n504), .Y(n597) );
  NAND2X0_HVT U226 ( .A1(n408), .A2(n409), .Y(n658) );
  INVX1_HVT U227 ( .A(n496), .Y(n497) );
  INVX1_HVT U228 ( .A(n562), .Y(n355) );
  INVX0_HVT U229 ( .A(n433), .Y(n519) );
  NAND2X0_HVT U230 ( .A1(n763), .A2(n502), .Y(n286) );
  NAND2X0_HVT U231 ( .A1(n566), .A2(n304), .Y(n290) );
  NAND2X0_HVT U232 ( .A1(n286), .A2(n290), .Y(n664) );
  NAND2X0_HVT U233 ( .A1(n485), .A2(n291), .Y(n293) );
  NAND2X0_HVT U234 ( .A1(n314), .A2(n338), .Y(n296) );
  NAND2X0_HVT U235 ( .A1(n293), .A2(n296), .Y(n765) );
  INVX0_HVT U236 ( .A(n765), .Y(n566) );
  INVX1_HVT U237 ( .A(n342), .Y(n340) );
  MUX41X1_HVT U238 ( .A1(n217), .A3(n537), .A2(n761), .A4(n488), .S0(n343), 
        .S1(n272), .Y(n656) );
  INVX1_HVT U239 ( .A(n574), .Y(n297) );
  INVX0_HVT U240 ( .A(n19), .Y(n574) );
  MUX41X1_HVT U242 ( .A1(n654), .A3(n656), .A2(n657), .A4(n658), .S0(n503), 
        .S1(n508), .Y(n653) );
  INVX1_HVT U243 ( .A(n519), .Y(n321) );
  INVX0_HVT U244 ( .A(n775), .Y(n543) );
  NAND2X0_HVT U246 ( .A1(n787), .A2(n500), .Y(n301) );
  NAND2X0_HVT U247 ( .A1(n231), .A2(n304), .Y(n303) );
  NAND2X0_HVT U248 ( .A1(n301), .A2(n303), .Y(n684) );
  MUX41X1_HVT U249 ( .A1(n280), .A3(n554), .A2(n771), .A4(n495), .S0(n470), 
        .S1(n421), .Y(n666) );
  NAND2X0_HVT U250 ( .A1(n774), .A2(n304), .Y(n305) );
  NAND2X0_HVT U251 ( .A1(n551), .A2(n500), .Y(n306) );
  NAND2X0_HVT U252 ( .A1(n305), .A2(n306), .Y(n661) );
  NAND2X0_HVT U253 ( .A1(n485), .A2(n309), .Y(n307) );
  NAND2X0_HVT U254 ( .A1(n555), .A2(n413), .Y(n308) );
  NAND2X0_HVT U255 ( .A1(n307), .A2(n308), .Y(n762) );
  INVX0_HVT U257 ( .A(n514), .Y(n555) );
  INVX0_HVT U258 ( .A(n762), .Y(n551) );
  NAND2X0_HVT U259 ( .A1(n672), .A2(n500), .Y(n310) );
  NAND2X0_HVT U260 ( .A1(n552), .A2(n304), .Y(n311) );
  NAND2X0_HVT U261 ( .A1(n310), .A2(n311), .Y(n671) );
  MUX21X1_HVT U262 ( .A1(n670), .A2(n671), .S0(n427), .Y(n667) );
  MUX41X1_HVT U263 ( .A1(n491), .A3(n571), .A2(n776), .A4(n291), .S0(n452), 
        .S1(n529), .Y(n696) );
  MUX41X1_HVT U264 ( .A1(n771), .A3(n565), .A2(n366), .A4(n629), .S0(n282), 
        .S1(n497), .Y(n628) );
  INVX1_HVT U266 ( .A(n454), .Y(n773) );
  INVX1_HVT U267 ( .A(n440), .Y(n331) );
  INVX0_HVT U269 ( .A(n465), .Y(n485) );
  INVX1_HVT U271 ( .A(n526), .Y(n525) );
  MUX41X1_HVT U272 ( .A1(n704), .A3(n699), .A2(n697), .A4(n696), .S0(n480), 
        .S1(n388), .Y(n695) );
  MUX21X2_HVT U273 ( .A1(n345), .A2(n346), .S0(n380), .Y(n344) );
  INVX1_HVT U274 ( .A(n514), .Y(n346) );
  INVX1_HVT U275 ( .A(n362), .Y(n320) );
  MUX21X1_HVT U276 ( .A1(n466), .A2(n398), .S0(n439), .Y(n441) );
  INVX1_HVT U277 ( .A(n331), .Y(n316) );
  NAND2X0_HVT U279 ( .A1(n511), .A2(n380), .Y(n318) );
  NAND2X0_HVT U280 ( .A1(n485), .A2(n313), .Y(n319) );
  NAND2X0_HVT U281 ( .A1(n318), .A2(n319), .Y(n763) );
  AO21X1_HVT U282 ( .A1(n433), .A2(n400), .A3(n386), .Y(n691) );
  INVX1_HVT U283 ( .A(n399), .Y(n400) );
  NAND2X0_HVT U285 ( .A1(n517), .A2(n321), .Y(n322) );
  NAND2X0_HVT U286 ( .A1(n780), .A2(n316), .Y(n323) );
  INVX0_HVT U287 ( .A(n374), .Y(n415) );
  INVX0_HVT U288 ( .A(n788), .Y(n416) );
  XNOR2X1_HVT U290 ( .A1(n314), .A2(n521), .Y(n492) );
  INVX1_HVT U291 ( .A(n579), .Y(n563) );
  INVX1_HVT U292 ( .A(n431), .Y(n324) );
  INVX1_HVT U293 ( .A(n467), .Y(n431) );
  NAND2X0_HVT U294 ( .A1(n564), .A2(n368), .Y(n325) );
  NAND2X0_HVT U298 ( .A1(n577), .A2(n418), .Y(n326) );
  NAND2X0_HVT U299 ( .A1(n325), .A2(n326), .Y(n600) );
  NBUFFX2_HVT U300 ( .A(n315), .Y(n467) );
  AO21X1_HVT U301 ( .A1(n486), .A2(n700), .A3(n567), .Y(n701) );
  NBUFFX2_HVT U302 ( .A(n562), .Y(n465) );
  MUX21X1_HVT U303 ( .A1(n514), .A2(n467), .S0(n313), .Y(n781) );
  NAND2X0_HVT U304 ( .A1(n520), .A2(n345), .Y(n753) );
  MUX41X1_HVT U305 ( .A1(n770), .A3(n572), .A2(n211), .A4(n739), .S0(n343), 
        .S1(n532), .Y(n593) );
  INVX1_HVT U307 ( .A(n334), .Y(n335) );
  NAND2X0_HVT U308 ( .A1(n518), .A2(n788), .Y(n787) );
  INVX1_HVT U309 ( .A(n329), .Y(n330) );
  INVX1_HVT U310 ( .A(n760), .Y(n572) );
  NAND2X0_HVT U311 ( .A1(n513), .A2(n331), .Y(n332) );
  NAND2X0_HVT U312 ( .A1(n461), .A2(n440), .Y(n333) );
  NAND2X0_HVT U313 ( .A1(n332), .A2(n333), .Y(n758) );
  INVX0_HVT U314 ( .A(in[1]), .Y(n334) );
  MUX41X1_HVT U315 ( .A1(n604), .A3(n759), .A2(n746), .A4(n753), .S0(n383), 
        .S1(n452), .Y(n603) );
  INVX1_HVT U316 ( .A(n341), .Y(n759) );
  INVX1_HVT U317 ( .A(n497), .Y(n452) );
  OR2X1_HVT U318 ( .A1(n390), .A2(n458), .Y(n777) );
  INVX0_HVT U319 ( .A(n498), .Y(n343) );
  INVX1_HVT U320 ( .A(n526), .Y(n524) );
  INVX0_HVT U321 ( .A(n433), .Y(n440) );
  MUX41X1_HVT U322 ( .A1(n754), .A3(n766), .A2(n456), .A4(n404), .S0(n455), 
        .S1(n525), .Y(n602) );
  INVX0_HVT U323 ( .A(n540), .Y(n357) );
  AO21X1_HVT U324 ( .A1(n492), .A2(n455), .A3(n567), .Y(n599) );
  INVX0_HVT U325 ( .A(n511), .Y(n345) );
  INVX0_HVT U326 ( .A(in[3]), .Y(n576) );
  INVX1_HVT U327 ( .A(n424), .Y(n347) );
  INVX1_HVT U328 ( .A(in[6]), .Y(n424) );
  NAND2X0_HVT U329 ( .A1(n653), .A2(n347), .Y(n348) );
  NAND2X0_HVT U330 ( .A1(n645), .A2(n424), .Y(n349) );
  NAND2X0_HVT U331 ( .A1(n349), .A2(n348), .Y(out[4]) );
  NAND2X0_HVT U332 ( .A1(n450), .A2(n451), .Y(out[6]) );
  NBUFFX2_HVT U333 ( .A(n530), .Y(n507) );
  MUX21X1_HVT U334 ( .A1(n403), .A2(n374), .S0(n413), .Y(n350) );
  NAND2X0_HVT U335 ( .A1(n489), .A2(n457), .Y(n468) );
  MUX41X1_HVT U336 ( .A1(n491), .A3(n578), .A2(n698), .A4(n570), .S0(n343), 
        .S1(n484), .Y(n697) );
  MUX41X1_HVT U337 ( .A1(n568), .A3(n708), .A2(n492), .A4(n488), .S0(n264), 
        .S1(n455), .Y(n707) );
  NAND2X0_HVT U338 ( .A1(n268), .A2(n314), .Y(n721) );
  MUX21X1_HVT U339 ( .A1(n337), .A2(n511), .S0(n339), .Y(n775) );
  NBUFFX2_HVT U340 ( .A(n210), .Y(n515) );
  MUX21X1_HVT U341 ( .A1(n573), .A2(n555), .S0(n521), .Y(n757) );
  NAND2X0_HVT U342 ( .A1(n516), .A2(n352), .Y(n353) );
  NAND2X0_HVT U343 ( .A1(n703), .A2(n494), .Y(n354) );
  NAND2X0_HVT U344 ( .A1(n353), .A2(n354), .Y(n702) );
  INVX0_HVT U345 ( .A(n494), .Y(n352) );
  MUX41X1_HVT U346 ( .A1(n665), .A3(n660), .A2(n679), .A4(n673), .S0(n476), 
        .S1(in[6]), .Y(out[3]) );
  NAND2X0_HVT U347 ( .A1(n490), .A2(n358), .Y(n359) );
  NAND2X0_HVT U348 ( .A1(n694), .A2(n748), .Y(n360) );
  NAND2X0_HVT U349 ( .A1(n359), .A2(n360), .Y(n693) );
  INVX0_HVT U350 ( .A(n748), .Y(n358) );
  INVX0_HVT U351 ( .A(n350), .Y(n361) );
  MUX41X1_HVT U352 ( .A1(n777), .A3(n545), .A2(n620), .A4(n340), .S0(n317), 
        .S1(n343), .Y(n619) );
  INVX0_HVT U353 ( .A(n442), .Y(n764) );
  MUX41X1_HVT U354 ( .A1(n568), .A3(n571), .A2(n534), .A4(n414), .S0(n443), 
        .S1(n507), .Y(n719) );
  XNOR2X1_HVT U355 ( .A1(n502), .A2(n418), .Y(n748) );
  INVX1_HVT U356 ( .A(in[2]), .Y(n526) );
  INVX0_HVT U357 ( .A(n681), .Y(n557) );
  INVX0_HVT U358 ( .A(n585), .Y(n568) );
  INVX1_HVT U359 ( .A(n412), .Y(n499) );
  INVX0_HVT U360 ( .A(n509), .Y(n464) );
  NAND2X0_HVT U361 ( .A1(n737), .A2(n264), .Y(n363) );
  NAND2X0_HVT U362 ( .A1(n735), .A2(n443), .Y(n364) );
  NAND2X0_HVT U363 ( .A1(n363), .A2(n364), .Y(n734) );
  MUX41X1_HVT U364 ( .A1(n610), .A3(n613), .A2(n606), .A4(n609), .S0(n504), 
        .S1(n476), .Y(n605) );
  INVX1_HVT U365 ( .A(n365), .Y(n366) );
  INVX0_HVT U366 ( .A(n498), .Y(n387) );
  NAND2X0_HVT U367 ( .A1(n744), .A2(n368), .Y(n369) );
  NAND2X0_HVT U368 ( .A1(n743), .A2(n383), .Y(n370) );
  NAND2X0_HVT U369 ( .A1(n369), .A2(n370), .Y(n741) );
  INVX0_HVT U370 ( .A(n755), .Y(n535) );
  NAND2X0_HVT U371 ( .A1(n786), .A2(n377), .Y(n371) );
  NAND2X0_HVT U372 ( .A1(n655), .A2(n443), .Y(n372) );
  NAND2X0_HVT U373 ( .A1(n372), .A2(n371), .Y(n654) );
  INVX1_HVT U374 ( .A(n403), .Y(n404) );
  MUX41X1_HVT U375 ( .A1(n711), .A3(n707), .A2(n712), .A4(n709), .S0(n476), 
        .S1(n503), .Y(n706) );
  INVX1_HVT U376 ( .A(n373), .Y(n456) );
  MUX21X1_HVT U377 ( .A1(n459), .A2(n402), .S0(n268), .Y(n373) );
  AND2X1_HVT U378 ( .A1(n315), .A2(n465), .Y(n374) );
  MUX41X1_HVT U379 ( .A1(n652), .A3(n551), .A2(n768), .A4(n553), .S0(n500), 
        .S1(n418), .Y(n651) );
  OR2X1_HVT U380 ( .A1(n375), .A2(n527), .Y(n392) );
  MUX41X1_HVT U381 ( .A1(n297), .A3(n537), .A2(n749), .A4(n571), .S0(n443), 
        .S1(n530), .Y(n646) );
  NAND2X0_HVT U382 ( .A1(n725), .A2(n377), .Y(n378) );
  NAND2X0_HVT U383 ( .A1(n751), .A2(n443), .Y(n379) );
  NAND2X0_HVT U384 ( .A1(n378), .A2(n379), .Y(n724) );
  INVX0_HVT U385 ( .A(n457), .Y(n377) );
  NAND2X0_HVT U386 ( .A1(n478), .A2(n479), .Y(out[1]) );
  MUX21X1_HVT U387 ( .A1(n367), .A2(n570), .S0(n486), .Y(n725) );
  MUX41X1_HVT U388 ( .A1(n617), .A3(n619), .A2(n615), .A4(n616), .S0(n504), 
        .S1(n476), .Y(n614) );
  INVX1_HVT U389 ( .A(n508), .Y(n476) );
  NBUFFX2_HVT U390 ( .A(n525), .Y(n501) );
  NAND2X0_HVT U391 ( .A1(n427), .A2(n376), .Y(n381) );
  NAND2X0_HVT U392 ( .A1(n368), .A2(n766), .Y(n382) );
  NAND2X0_HVT U393 ( .A1(n381), .A2(n382), .Y(n751) );
  NAND2X0_HVT U394 ( .A1(n676), .A2(n507), .Y(n385) );
  NAND2X0_HVT U395 ( .A1(n384), .A2(n385), .Y(n674) );
  MUX21X1_HVT U396 ( .A1(n511), .A2(n374), .S0(n291), .Y(n755) );
  NAND2X0_HVT U397 ( .A1(n669), .A2(n668), .Y(n670) );
  MUX41X1_HVT U398 ( .A1(n662), .A3(n664), .A2(n661), .A4(n663), .S0(n527), 
        .S1(n386), .Y(n660) );
  MUX41X1_HVT U399 ( .A1(n570), .A3(n218), .A2(n758), .A4(n517), .S0(n387), 
        .S1(n484), .Y(n601) );
  INVX1_HVT U400 ( .A(in[4]), .Y(n562) );
  INVX0_HVT U401 ( .A(n778), .Y(n549) );
  INVX1_HVT U402 ( .A(n581), .Y(n537) );
  NAND2X0_HVT U403 ( .A1(n759), .A2(n505), .Y(n393) );
  NAND2X0_HVT U404 ( .A1(n393), .A2(n392), .Y(n744) );
  NAND2X0_HVT U405 ( .A1(n638), .A2(n470), .Y(n394) );
  NAND2X0_HVT U406 ( .A1(n637), .A2(n387), .Y(n395) );
  NAND2X0_HVT U407 ( .A1(n394), .A2(n395), .Y(n636) );
  NAND2X0_HVT U408 ( .A1(n621), .A2(n424), .Y(n396) );
  NAND2X0_HVT U409 ( .A1(n633), .A2(n347), .Y(n397) );
  NAND2X0_HVT U410 ( .A1(n396), .A2(n397), .Y(out[5]) );
  MUX21X1_HVT U411 ( .A1(n639), .A2(n232), .S0(n494), .Y(n638) );
  NAND2X0_HVT U412 ( .A1(n464), .A2(n510), .Y(n398) );
  NAND2X0_HVT U413 ( .A1(n464), .A2(n320), .Y(n399) );
  INVX1_HVT U414 ( .A(n400), .Y(n401) );
  INVX0_HVT U415 ( .A(n398), .Y(n402) );
  INVX0_HVT U416 ( .A(n780), .Y(n403) );
  INVX1_HVT U417 ( .A(n441), .Y(n774) );
  NAND2X0_HVT U418 ( .A1(n599), .A2(n502), .Y(n406) );
  NAND2X0_HVT U419 ( .A1(n600), .A2(n443), .Y(n407) );
  NAND2X0_HVT U420 ( .A1(n406), .A2(n407), .Y(n598) );
  NAND2X0_HVT U421 ( .A1(n659), .A2(n377), .Y(n408) );
  NAND2X0_HVT U422 ( .A1(n533), .A2(n387), .Y(n409) );
  NAND2X0_HVT U423 ( .A1(n666), .A2(n480), .Y(n410) );
  NAND2X0_HVT U424 ( .A1(n667), .A2(n503), .Y(n411) );
  NAND2X0_HVT U425 ( .A1(n411), .A2(n410), .Y(n665) );
  XNOR2X1_HVT U426 ( .A1(n520), .A2(n496), .Y(n412) );
  MUX21X1_HVT U427 ( .A1(n398), .A2(n485), .S0(n413), .Y(n580) );
  INVX1_HVT U428 ( .A(n416), .Y(n417) );
  MUX41X1_HVT U429 ( .A1(n766), .A3(n784), .A2(n569), .A4(n456), .S0(n304), 
        .S1(n418), .Y(n657) );
  NAND2X0_HVT U430 ( .A1(n414), .A2(n412), .Y(n419) );
  NAND2X0_HVT U431 ( .A1(n432), .A2(n499), .Y(n420) );
  OA21X1_HVT U432 ( .A1(n755), .A2(n386), .A3(n642), .Y(n643) );
  NAND2X0_HVT U433 ( .A1(n701), .A2(n443), .Y(n422) );
  NAND2X0_HVT U434 ( .A1(n702), .A2(n502), .Y(n423) );
  NAND2X0_HVT U435 ( .A1(n422), .A2(n423), .Y(n699) );
  NAND2X0_HVT U436 ( .A1(n685), .A2(n424), .Y(n425) );
  NAND2X0_HVT U437 ( .A1(n695), .A2(n347), .Y(n426) );
  NAND2X0_HVT U438 ( .A1(n425), .A2(n426), .Y(out[2]) );
  INVX1_HVT U439 ( .A(n584), .Y(n546) );
  MUX41X1_HVT U440 ( .A1(n557), .A3(n512), .A2(n544), .A4(n356), .S0(n470), 
        .S1(n429), .Y(n650) );
  MUX21X1_HVT U441 ( .A1(n416), .A2(n403), .S0(n428), .Y(n629) );
  MUX21X1_HVT U442 ( .A1(n431), .A2(n466), .S0(n525), .Y(n432) );
  INVX1_HVT U443 ( .A(n580), .Y(n564) );
  NAND2X0_HVT U444 ( .A1(n648), .A2(n377), .Y(n434) );
  NAND2X0_HVT U445 ( .A1(n649), .A2(n443), .Y(n435) );
  NAND2X0_HVT U446 ( .A1(n434), .A2(n435), .Y(n647) );
  NAND2X0_HVT U447 ( .A1(n512), .A2(n531), .Y(n437) );
  NAND2X0_HVT U448 ( .A1(n554), .A2(n383), .Y(n438) );
  NAND2X0_HVT U449 ( .A1(n437), .A2(n438), .Y(n659) );
  INVX1_HVT U450 ( .A(n587), .Y(n547) );
  MUX21X1_HVT U451 ( .A1(n513), .A2(n464), .S0(n428), .Y(n442) );
  NAND2X0_HVT U452 ( .A1(n731), .A2(n443), .Y(n444) );
  NAND2X0_HVT U453 ( .A1(n733), .A2(n501), .Y(n445) );
  NAND2X0_HVT U454 ( .A1(n444), .A2(n445), .Y(n730) );
  NAND2X0_HVT U455 ( .A1(n682), .A2(n264), .Y(n446) );
  NAND2X0_HVT U456 ( .A1(n212), .A2(n457), .Y(n447) );
  NAND2X0_HVT U457 ( .A1(n446), .A2(n447), .Y(n680) );
  NAND2X0_HVT U458 ( .A1(n591), .A2(n424), .Y(n448) );
  NAND2X0_HVT U459 ( .A1(n597), .A2(n347), .Y(n449) );
  NAND2X0_HVT U460 ( .A1(n449), .A2(n448), .Y(out[7]) );
  NAND2X0_HVT U461 ( .A1(n605), .A2(n424), .Y(n450) );
  NAND2X0_HVT U462 ( .A1(n614), .A2(n347), .Y(n451) );
  OA21X1_HVT U463 ( .A1(n493), .A2(n427), .A3(n212), .Y(n623) );
  MUX21X1_HVT U464 ( .A1(n780), .A2(n513), .S0(n256), .Y(n453) );
  INVX1_HVT U465 ( .A(n583), .Y(n533) );
  INVX1_HVT U466 ( .A(n582), .Y(n554) );
  OA21X1_HVT U467 ( .A1(n760), .A2(n386), .A3(n544), .Y(n611) );
  MUX41X1_HVT U468 ( .A1(n736), .A3(n495), .A2(n453), .A4(n493), .S0(n383), 
        .S1(n528), .Y(n735) );
  MUX41X1_HVT U469 ( .A1(n563), .A3(n765), .A2(n564), .A4(n548), .S0(n387), 
        .S1(n531), .Y(n616) );
  MUX41X1_HVT U470 ( .A1(n749), .A3(n297), .A2(n756), .A4(n491), .S0(n496), 
        .S1(n429), .Y(n609) );
  INVX1_HVT U471 ( .A(n337), .Y(n459) );
  INVX1_HVT U472 ( .A(n461), .Y(n463) );
  NBUFFX2_HVT U473 ( .A(n283), .Y(n466) );
  NAND2X0_HVT U474 ( .A1(n543), .A2(n264), .Y(n469) );
  NAND2X0_HVT U475 ( .A1(n468), .A2(n469), .Y(n662) );
  NAND2X0_HVT U476 ( .A1(n596), .A2(n470), .Y(n471) );
  NAND2X0_HVT U477 ( .A1(n472), .A2(n471), .Y(n595) );
  INVX0_HVT U478 ( .A(n457), .Y(n470) );
  NAND2X0_HVT U479 ( .A1(n487), .A2(n473), .Y(n474) );
  NAND2X0_HVT U480 ( .A1(n775), .A2(n317), .Y(n475) );
  NAND2X0_HVT U481 ( .A1(n475), .A2(n474), .Y(n596) );
  INVX0_HVT U482 ( .A(n421), .Y(n473) );
  INVX0_HVT U483 ( .A(n504), .Y(n477) );
  XNOR2X1_HVT U484 ( .A1(n330), .A2(n521), .Y(n494) );
  MUX41X1_HVT U485 ( .A1(n350), .A3(n549), .A2(n541), .A4(n732), .S0(n383), 
        .S1(n477), .Y(n731) );
  NAND2X0_HVT U486 ( .A1(n706), .A2(n424), .Y(n478) );
  NAND2X0_HVT U487 ( .A1(n716), .A2(n347), .Y(n479) );
  INVX1_HVT U488 ( .A(n586), .Y(n570) );
  MUX41X1_HVT U489 ( .A1(n391), .A3(n762), .A2(n217), .A4(n535), .S0(n497), 
        .S1(n418), .Y(n594) );
  NAND2X0_HVT U490 ( .A1(n674), .A2(n480), .Y(n482) );
  NAND2X0_HVT U491 ( .A1(n677), .A2(n505), .Y(n483) );
  NAND2X0_HVT U492 ( .A1(n482), .A2(n483), .Y(n673) );
  NBUFFX2_HVT U493 ( .A(n530), .Y(n486) );
  AND2X1_HVT U494 ( .A1(n356), .A2(n738), .Y(n487) );
  NBUFFX2_HVT U495 ( .A(n210), .Y(n513) );
  MUX21X1_HVT U496 ( .A1(n555), .A2(n367), .S0(n505), .Y(n742) );
  NBUFFX2_HVT U497 ( .A(n785), .Y(n514) );
  AND2X1_HVT U498 ( .A1(n417), .A2(n721), .Y(n488) );
  MUX21X1_HVT U499 ( .A1(n463), .A2(n466), .S0(n336), .Y(n690) );
  MUX21X1_HVT U500 ( .A1(n555), .A2(n416), .S0(n439), .Y(n620) );
  NAND2X0_HVT U501 ( .A1(n509), .A2(n320), .Y(n785) );
  MUX21X1_HVT U502 ( .A1(n555), .A2(n340), .S0(n309), .Y(n582) );
  MUX21X1_HVT U503 ( .A1(n510), .A2(n461), .S0(n291), .Y(n584) );
  NBUFFX2_HVT U504 ( .A(n788), .Y(n516) );
  MUX21X1_HVT U505 ( .A1(n341), .A2(n572), .S0(n502), .Y(n676) );
  MUX21X1_HVT U506 ( .A1(n573), .A2(n510), .S0(n521), .Y(n760) );
  MUX21X1_HVT U507 ( .A1(n340), .A2(n510), .S0(n256), .Y(n672) );
  MUX21X1_HVT U508 ( .A1(n510), .A2(n314), .S0(n336), .Y(n607) );
  MUX21X1_HVT U509 ( .A1(n314), .A2(n417), .S0(n520), .Y(n608) );
  MUX21X1_HVT U510 ( .A1(n513), .A2(n517), .S0(n268), .Y(n700) );
  MUX21X1_HVT U511 ( .A1(n511), .A2(n340), .S0(n519), .Y(n604) );
  MUX21X1_HVT U512 ( .A1(n516), .A2(n515), .S0(n339), .Y(n581) );
  XNOR2X1_HVT U513 ( .A1(n515), .A2(n309), .Y(n489) );
  MUX21X1_HVT U514 ( .A1(n417), .A2(n466), .S0(n316), .Y(n588) );
  AND2X1_HVT U515 ( .A1(n312), .A2(n681), .Y(n490) );
  AND2X1_HVT U516 ( .A1(n520), .A2(n416), .Y(n491) );
  MUX21X1_HVT U517 ( .A1(n398), .A2(n511), .S0(n519), .Y(n586) );
  MUX21X1_HVT U518 ( .A1(n404), .A2(n314), .S0(n497), .Y(n669) );
  XOR2X1_HVT U519 ( .A1(n466), .A2(n439), .Y(n767) );
  NBUFFX2_HVT U520 ( .A(n389), .Y(n510) );
  NBUFFX2_HVT U521 ( .A(n576), .Y(n511) );
  NBUFFX2_HVT U522 ( .A(n528), .Y(n504) );
  NBUFFX2_HVT U523 ( .A(n525), .Y(n502) );
  NBUFFX2_HVT U524 ( .A(n527), .Y(n503) );
  MUX21X1_HVT U525 ( .A1(n512), .A2(n570), .S0(n507), .Y(n624) );
  NAND2X0_HVT U526 ( .A1(n315), .A2(n509), .Y(n788) );
  AND2X1_HVT U527 ( .A1(n462), .A2(n523), .Y(n493) );
  OA21X1_HVT U528 ( .A1(n550), .A2(n526), .A3(n453), .Y(n683) );
  NBUFFX2_HVT U529 ( .A(n780), .Y(n512) );
  XOR2X1_HVT U530 ( .A1(n309), .A2(n504), .Y(n752) );
  MUX21X1_HVT U531 ( .A1(n763), .A2(n589), .S0(n486), .Y(n583) );
  MUX21X1_HVT U532 ( .A1(n345), .A2(n400), .S0(n309), .Y(n585) );
  MUX21X1_HVT U533 ( .A1(n787), .A2(n428), .S0(n501), .Y(n668) );
  MUX21X1_HVT U534 ( .A1(n324), .A2(n340), .S0(n506), .Y(n703) );
  NBUFFX2_HVT U535 ( .A(n789), .Y(n517) );
  AND2X1_HVT U536 ( .A1(n375), .A2(n523), .Y(n495) );
  NBUFFX2_HVT U537 ( .A(in[5]), .Y(n528) );
  NAND2X0_HVT U538 ( .A1(n362), .A2(n355), .Y(n789) );
  NAND2X0_HVT U539 ( .A1(n464), .A2(n510), .Y(n780) );
  MUX21X1_HVT U540 ( .A1(n485), .A2(n218), .S0(n256), .Y(n587) );
endmodule

