
module sbox_9 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n7, n23, n210, n211, n212, n213, n216, n217, n218, n219, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580;

  NAND2X0_HVT U4 ( .A1(n289), .A2(n578), .Y(n577) );
  NAND2X0_HVT U5 ( .A1(n219), .A2(n280), .Y(n575) );
  NAND2X0_HVT U13 ( .A1(n568), .A2(n292), .Y(n569) );
  NAND2X0_HVT U15 ( .A1(n578), .A2(n282), .Y(n566) );
  NAND2X0_HVT U21 ( .A1(n289), .A2(n299), .Y(n560) );
  NAND2X0_HVT U24 ( .A1(n286), .A2(n299), .Y(n558) );
  NAND2X0_HVT U33 ( .A1(n356), .A2(n299), .Y(n549) );
  NAND2X0_HVT U35 ( .A1(n284), .A2(n299), .Y(n547) );
  NAND2X0_HVT U42 ( .A1(n297), .A2(n285), .Y(n540) );
  MUX41X1_HVT U51 ( .A1(n345), .A3(n305), .A2(n322), .A4(n323), .S0(n246), 
        .S1(n300), .Y(n531) );
  NAND2X0_HVT U53 ( .A1(n528), .A2(n539), .Y(n529) );
  NAND2X0_HVT U56 ( .A1(n289), .A2(n524), .Y(n525) );
  MUX41X1_HVT U57 ( .A1(n346), .A3(n562), .A2(n525), .A4(n571), .S0(n246), 
        .S1(n300), .Y(n523) );
  NAND2X0_HVT U58 ( .A1(n292), .A2(n578), .Y(n522) );
  MUX41X1_HVT U59 ( .A1(n270), .A3(n522), .A2(n268), .A4(n321), .S0(n246), 
        .S1(n300), .Y(n521) );
  MUX41X1_HVT U61 ( .A1(n267), .A3(n320), .A2(n239), .A4(n281), .S0(n246), 
        .S1(in[5]), .Y(n519) );
  NAND2X0_HVT U62 ( .A1(n299), .A2(n579), .Y(n518) );
  MUX41X1_HVT U63 ( .A1(n518), .A3(n312), .A2(n340), .A4(n319), .S0(n246), 
        .S1(n300), .Y(n517) );
  AO21X1_HVT U66 ( .A1(n317), .A2(in[5]), .A3(n339), .Y(n514) );
  MUX41X1_HVT U68 ( .A1(n315), .A3(n514), .A2(n513), .A4(n515), .S0(n271), 
        .S1(n249), .Y(n512) );
  MUX41X1_HVT U69 ( .A1(n512), .A3(n520), .A2(n516), .A4(n526), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n287), .A2(n507), .Y(n508) );
  MUX41X1_HVT U74 ( .A1(n509), .A3(n556), .A2(n508), .A4(n558), .S0(n273), 
        .S1(n302), .Y(n506) );
  MUX41X1_HVT U75 ( .A1(n343), .A3(n348), .A2(n232), .A4(n254), .S0(n271), 
        .S1(n210), .Y(n505) );
  MUX41X1_HVT U77 ( .A1(n573), .A3(n350), .A2(n504), .A4(n349), .S0(n277), 
        .S1(n273), .Y(n503) );
  MUX41X1_HVT U78 ( .A1(n503), .A3(n506), .A2(n505), .A4(n510), .S0(in[0]), 
        .S1(n301), .Y(n502) );
  AND3X1_HVT U80 ( .A1(n290), .A2(n524), .A3(n499), .Y(n500) );
  MUX41X1_HVT U82 ( .A1(n537), .A3(n323), .A2(n306), .A4(n567), .S0(n271), 
        .S1(n210), .Y(n497) );
  AND2X1_HVT U83 ( .A1(n294), .A2(n245), .Y(n496) );
  MUX41X1_HVT U84 ( .A1(n324), .A3(n240), .A2(n565), .A4(n496), .S0(n271), 
        .S1(n210), .Y(n495) );
  NAND2X0_HVT U85 ( .A1(n299), .A2(n359), .Y(n494) );
  AO21X1_HVT U93 ( .A1(n279), .A2(n486), .A3(n344), .Y(n487) );
  MUX41X1_HVT U96 ( .A1(n306), .A3(n266), .A2(n347), .A4(n484), .S0(n271), 
        .S1(n210), .Y(n483) );
  MUX41X1_HVT U97 ( .A1(n343), .A3(n266), .A2(n231), .A4(n566), .S0(n271), 
        .S1(n304), .Y(n482) );
  MUX41X1_HVT U98 ( .A1(n482), .A3(n485), .A2(n483), .A4(n490), .S0(in[0]), 
        .S1(n301), .Y(n481) );
  NAND2X0_HVT U101 ( .A1(n477), .A2(n476), .Y(n478) );
  MUX41X1_HVT U103 ( .A1(n578), .A3(n316), .A2(n244), .A4(n547), .S0(n271), 
        .S1(n304), .Y(n474) );
  MUX41X1_HVT U105 ( .A1(n326), .A3(n534), .A2(n473), .A4(n342), .S0(n271), 
        .S1(n304), .Y(n472) );
  NAND2X0_HVT U110 ( .A1(n290), .A2(n467), .Y(n468) );
  AND2X1_HVT U115 ( .A1(n296), .A2(n281), .Y(n462) );
  MUX41X1_HVT U116 ( .A1(n569), .A3(n462), .A2(n254), .A4(n551), .S0(n272), 
        .S1(n302), .Y(n461) );
  AO21X1_HVT U118 ( .A1(n275), .A2(n572), .A3(n240), .Y(n459) );
  NAND2X0_HVT U123 ( .A1(n453), .A2(n452), .Y(n454) );
  MUX41X1_HVT U125 ( .A1(n560), .A3(n270), .A2(n315), .A4(n352), .S0(n272), 
        .S1(n302), .Y(n450) );
  MUX41X1_HVT U131 ( .A1(n445), .A3(n447), .A2(n446), .A4(n448), .S0(in[5]), 
        .S1(n246), .Y(n444) );
  MUX41X1_HVT U135 ( .A1(n353), .A3(n357), .A2(n575), .A4(n555), .S0(n274), 
        .S1(n249), .Y(n441) );
  MUX41X1_HVT U136 ( .A1(n263), .A3(n549), .A2(n354), .A4(n546), .S0(n272), 
        .S1(n249), .Y(n440) );
  AND2X1_HVT U140 ( .A1(n572), .A2(n299), .Y(n436) );
  MUX41X1_HVT U141 ( .A1(n557), .A3(n334), .A2(n436), .A4(n330), .S0(n271), 
        .S1(n304), .Y(n435) );
  MUX41X1_HVT U142 ( .A1(n324), .A3(n281), .A2(n341), .A4(n572), .S0(n272), 
        .S1(n302), .Y(n434) );
  NAND2X0_HVT U146 ( .A1(n297), .A2(n292), .Y(n507) );
  MUX41X1_HVT U148 ( .A1(n430), .A3(n434), .A2(n431), .A4(n435), .S0(in[0]), 
        .S1(n300), .Y(n429) );
  MUX41X1_HVT U153 ( .A1(n468), .A3(n267), .A2(n579), .A4(n308), .S0(n272), 
        .S1(n302), .Y(n424) );
  AND2X1_HVT U154 ( .A1(n279), .A2(n286), .Y(n423) );
  NAND2X0_HVT U158 ( .A1(n294), .A2(n359), .Y(n419) );
  MUX41X1_HVT U159 ( .A1(n569), .A3(n281), .A2(n419), .A4(n314), .S0(n271), 
        .S1(n304), .Y(n418) );
  MUX41X1_HVT U160 ( .A1(n418), .A3(n424), .A2(n420), .A4(n425), .S0(in[0]), 
        .S1(n276), .Y(n417) );
  AND2X1_HVT U162 ( .A1(n240), .A2(n507), .Y(n415) );
  MUX41X1_HVT U163 ( .A1(n320), .A3(n415), .A2(n264), .A4(n416), .S0(n274), 
        .S1(n304), .Y(n414) );
  NAND2X0_HVT U166 ( .A1(n292), .A2(n524), .Y(n411) );
  NAND2X0_HVT U167 ( .A1(n232), .A2(n299), .Y(n410) );
  MUX41X1_HVT U168 ( .A1(n346), .A3(n572), .A2(n410), .A4(n411), .S0(n273), 
        .S1(n249), .Y(n409) );
  MUX41X1_HVT U172 ( .A1(n406), .A3(n412), .A2(n409), .A4(n414), .S0(in[0]), 
        .S1(n276), .Y(n405) );
  NAND2X0_HVT U174 ( .A1(n231), .A2(n240), .Y(n568) );
  NAND2X0_HVT U177 ( .A1(n294), .A2(n283), .Y(n402) );
  MUX41X1_HVT U178 ( .A1(n564), .A3(n402), .A2(n242), .A4(n544), .S0(n275), 
        .S1(n249), .Y(n401) );
  MUX41X1_HVT U179 ( .A1(n554), .A3(n355), .A2(n310), .A4(n242), .S0(n275), 
        .S1(n249), .Y(n400) );
  MUX41X1_HVT U180 ( .A1(n313), .A3(n573), .A2(n569), .A4(n262), .S0(n277), 
        .S1(n275), .Y(n399) );
  MUX41X1_HVT U181 ( .A1(n399), .A3(n401), .A2(n400), .A4(n403), .S0(in[0]), 
        .S1(n276), .Y(n398) );
  MUX41X1_HVT U186 ( .A1(n266), .A3(n543), .A2(n507), .A4(n536), .S0(n275), 
        .S1(n302), .Y(n393) );
  MUX41X1_HVT U189 ( .A1(n391), .A3(n568), .A2(n392), .A4(n342), .S0(n277), 
        .S1(n274), .Y(n390) );
  AO21X1_HVT U197 ( .A1(n265), .A2(n278), .A3(n344), .Y(n383) );
  MUX41X1_HVT U203 ( .A1(n546), .A3(n336), .A2(n570), .A4(n550), .S0(n271), 
        .S1(n304), .Y(n377) );
  MUX41X1_HVT U205 ( .A1(n245), .A3(n578), .A2(n355), .A4(n329), .S0(n274), 
        .S1(n210), .Y(n375) );
  NAND2X0_HVT U208 ( .A1(n218), .A2(n289), .Y(n467) );
  NAND2X0_HVT U212 ( .A1(n293), .A2(n287), .Y(n524) );
  NAND2X0_HVT U214 ( .A1(n240), .A2(n299), .Y(n373) );
  NAND2X0_HVT U215 ( .A1(n467), .A2(n287), .Y(n372) );
  NAND2X0_HVT U218 ( .A1(n357), .A2(n296), .Y(n426) );
  NAND2X0_HVT U220 ( .A1(n278), .A2(n373), .Y(n499) );
  NAND2X0_HVT U1 ( .A1(n251), .A2(n252), .Y(out[4]) );
  MUX21X1_HVT U2 ( .A1(n379), .A2(n380), .S0(n273), .Y(n378) );
  INVX2_HVT U3 ( .A(in[1]), .Y(n299) );
  IBUFFX2_HVT U6 ( .A(n210), .Y(n212) );
  MUX21X1_HVT U7 ( .A1(n500), .A2(n501), .S0(n255), .Y(n498) );
  MUX41X1_HVT U8 ( .A1(n442), .A3(n440), .A2(n441), .A4(n438), .S0(n7), .S1(
        n23), .Y(n437) );
  IBUFFX16_HVT U9 ( .A(in[0]), .Y(n7) );
  IBUFFX16_HVT U10 ( .A(n276), .Y(n23) );
  INVX1_HVT U11 ( .A(n248), .Y(n210) );
  MUX41X1_HVT U12 ( .A1(n263), .A3(n265), .A2(n494), .A4(n348), .S0(n211), 
        .S1(n212), .Y(n493) );
  IBUFFX16_HVT U14 ( .A(n271), .Y(n211) );
  INVX0_HVT U16 ( .A(n248), .Y(n303) );
  INVX2_HVT U17 ( .A(n298), .Y(n293) );
  INVX2_HVT U18 ( .A(in[1]), .Y(n298) );
  XOR2X1_HVT U19 ( .A1(n253), .A2(n555), .Y(n538) );
  MUX21X1_HVT U20 ( .A1(n232), .A2(n359), .S0(n293), .Y(n555) );
  MUX41X1_HVT U22 ( .A1(n498), .A3(n495), .A2(n497), .A4(n493), .S0(n213), 
        .S1(n216), .Y(n492) );
  IBUFFX16_HVT U23 ( .A(in[0]), .Y(n213) );
  IBUFFX16_HVT U25 ( .A(n300), .Y(n216) );
  MUX21X2_HVT U26 ( .A1(n328), .A2(n443), .S0(n217), .Y(n442) );
  IBUFFX16_HVT U27 ( .A(n255), .Y(n217) );
  INVX1_HVT U28 ( .A(n365), .Y(n352) );
  NAND2X1_HVT U29 ( .A1(n294), .A2(n290), .Y(n578) );
  NBUFFX2_HVT U30 ( .A(n293), .Y(n218) );
  NBUFFX2_HVT U31 ( .A(n293), .Y(n219) );
  NBUFFX2_HVT U32 ( .A(n293), .Y(n231) );
  IBUFFX2_HVT U34 ( .A(n298), .Y(n295) );
  MUX21X1_HVT U36 ( .A1(n359), .A2(n347), .S0(n279), .Y(n511) );
  INVX1_HVT U37 ( .A(n248), .Y(n304) );
  INVX0_HVT U38 ( .A(n569), .Y(n340) );
  OA21X1_HVT U39 ( .A1(n548), .A2(n253), .A3(n324), .Y(n395) );
  XOR2X1_HVT U40 ( .A1(n240), .A2(n293), .Y(n536) );
  OA21X1_HVT U41 ( .A1(n542), .A2(n253), .A3(n426), .Y(n427) );
  INVX2_HVT U43 ( .A(in[7]), .Y(n248) );
  INVX1_HVT U44 ( .A(n278), .Y(n257) );
  INVX1_HVT U45 ( .A(in[0]), .Y(n247) );
  INVX1_HVT U46 ( .A(n579), .Y(n232) );
  XNOR2X1_HVT U47 ( .A1(n360), .A2(in[3]), .Y(n256) );
  INVX1_HVT U48 ( .A(n282), .Y(n240) );
  INVX1_HVT U49 ( .A(n284), .Y(n245) );
  INVX1_HVT U50 ( .A(in[4]), .Y(n360) );
  INVX1_HVT U52 ( .A(n279), .Y(n233) );
  INVX1_HVT U54 ( .A(n303), .Y(n253) );
  NBUFFX2_HVT U55 ( .A(n301), .Y(n276) );
  INVX0_HVT U60 ( .A(n300), .Y(n243) );
  INVX1_HVT U64 ( .A(in[2]), .Y(n255) );
  INVX1_HVT U65 ( .A(n272), .Y(n241) );
  INVX1_HVT U67 ( .A(n298), .Y(n296) );
  MUX21X2_HVT U70 ( .A1(n389), .A2(n398), .S0(in[6]), .Y(out[6]) );
  INVX2_HVT U71 ( .A(n298), .Y(n294) );
  MUX21X1_HVT U72 ( .A1(n565), .A2(n262), .S0(n277), .Y(n380) );
  XOR2X1_HVT U76 ( .A1(n299), .A2(n241), .Y(n533) );
  MUX21X2_HVT U79 ( .A1(n372), .A2(n552), .S0(n253), .Y(n366) );
  XNOR2X1_HVT U81 ( .A1(n232), .A2(n295), .Y(n532) );
  MUX41X1_HVT U86 ( .A1(n291), .A3(n545), .A2(n240), .A4(n347), .S0(n275), 
        .S1(n257), .Y(n385) );
  IBUFFX2_HVT U87 ( .A(n248), .Y(n302) );
  IBUFFX2_HVT U88 ( .A(n545), .Y(n333) );
  MUX21X2_HVT U89 ( .A1(n384), .A2(n383), .S0(n273), .Y(n382) );
  IBUFFX2_HVT U90 ( .A(n552), .Y(n327) );
  INVX0_HVT U91 ( .A(n561), .Y(n323) );
  MUX21X2_HVT U92 ( .A1(n577), .A2(n439), .S0(n255), .Y(n438) );
  INVX1_HVT U94 ( .A(n559), .Y(n324) );
  MUX21X2_HVT U95 ( .A1(n287), .A2(n561), .S0(n233), .Y(n501) );
  INVX0_HVT U99 ( .A(n254), .Y(n557) );
  MUX21X1_HVT U100 ( .A1(n579), .A2(n256), .S0(n299), .Y(n254) );
  NAND2X0_HVT U102 ( .A1(n553), .A2(n233), .Y(n234) );
  NAND2X0_HVT U104 ( .A1(n311), .A2(n279), .Y(n235) );
  NAND2X0_HVT U106 ( .A1(n234), .A2(n235), .Y(n433) );
  NBUFFX4_HVT U107 ( .A(n303), .Y(n279) );
  MUX21X1_HVT U108 ( .A1(n433), .A2(n432), .S0(n274), .Y(n431) );
  NAND2X0_HVT U109 ( .A1(n290), .A2(n236), .Y(n237) );
  NAND2X0_HVT U111 ( .A1(n489), .A2(n269), .Y(n238) );
  NAND2X0_HVT U112 ( .A1(n237), .A2(n238), .Y(n488) );
  INVX0_HVT U113 ( .A(n269), .Y(n236) );
  MUX21X1_HVT U114 ( .A1(n487), .A2(n488), .S0(n275), .Y(n485) );
  INVX1_HVT U117 ( .A(n366), .Y(n328) );
  MUX21X2_HVT U119 ( .A1(n405), .A2(n417), .S0(in[6]), .Y(out[5]) );
  MUX21X2_HVT U120 ( .A1(n421), .A2(n422), .S0(n275), .Y(n420) );
  OA21X1_HVT U121 ( .A1(n574), .A2(n233), .A3(n334), .Y(n379) );
  INVX0_HVT U122 ( .A(n239), .Y(n565) );
  MUX21X1_HVT U124 ( .A1(n240), .A2(n285), .S0(n296), .Y(n239) );
  MUX21X2_HVT U126 ( .A1(n381), .A2(n374), .S0(n258), .Y(out[7]) );
  INVX0_HVT U127 ( .A(n244), .Y(n553) );
  MUX21X1_HVT U128 ( .A1(n338), .A2(n242), .S0(n278), .Y(n384) );
  MUX41X1_HVT U129 ( .A1(n491), .A3(n345), .A2(n540), .A4(n536), .S0(n241), 
        .S1(n257), .Y(n490) );
  OA21X1_HVT U130 ( .A1(n309), .A2(n253), .A3(n551), .Y(n432) );
  IBUFFX2_HVT U132 ( .A(n298), .Y(n297) );
  INVX1_HVT U133 ( .A(n362), .Y(n242) );
  MUX41X1_HVT U134 ( .A1(n547), .A3(n540), .A2(n388), .A4(n532), .S0(n255), 
        .S1(n249), .Y(n387) );
  MUX41X1_HVT U137 ( .A1(n474), .A3(n479), .A2(n472), .A4(n475), .S0(in[0]), 
        .S1(n243), .Y(n471) );
  MUX21X1_HVT U138 ( .A1(n245), .A2(n288), .S0(n295), .Y(n244) );
  MUX21X2_HVT U139 ( .A1(n427), .A2(n428), .S0(n275), .Y(n425) );
  MUX21X2_HVT U143 ( .A1(n538), .A2(n511), .S0(n273), .Y(n510) );
  INVX1_HVT U144 ( .A(n369), .Y(n347) );
  IBUFFX2_HVT U145 ( .A(n253), .Y(n246) );
  MUX41X1_HVT U147 ( .A1(n378), .A3(n377), .A2(n376), .A4(n375), .S0(n243), 
        .S1(n247), .Y(n374) );
  MUX41X1_HVT U149 ( .A1(n331), .A3(n559), .A2(n525), .A4(n569), .S0(in[2]), 
        .S1(n233), .Y(n376) );
  INVX1_HVT U150 ( .A(n248), .Y(n249) );
  NAND2X0_HVT U151 ( .A1(n437), .A2(n250), .Y(n251) );
  NAND2X0_HVT U152 ( .A1(n429), .A2(n258), .Y(n252) );
  INVX1_HVT U155 ( .A(n258), .Y(n250) );
  INVX1_HVT U156 ( .A(n367), .Y(n349) );
  MUX21X2_HVT U157 ( .A1(n492), .A2(n502), .S0(in[6]), .Y(out[1]) );
  AND3X2_HVT U161 ( .A1(n274), .A2(n299), .A3(n245), .Y(n447) );
  OA21X2_HVT U164 ( .A1(n268), .A2(n233), .A3(n551), .Y(n407) );
  AO21X2_HVT U165 ( .A1(n299), .A2(n357), .A3(n253), .Y(n477) );
  MUX41X1_HVT U169 ( .A1(n536), .A3(n343), .A2(n507), .A4(n354), .S0(n255), 
        .S1(n248), .Y(n430) );
  INVX0_HVT U170 ( .A(in[6]), .Y(n258) );
  MUX41X1_HVT U171 ( .A1(n572), .A3(n353), .A2(n555), .A4(n541), .S0(n257), 
        .S1(n241), .Y(n386) );
  OA21X2_HVT U173 ( .A1(n333), .A2(n255), .A3(n321), .Y(n469) );
  MUX21X2_HVT U175 ( .A1(n335), .A2(n559), .S0(n257), .Y(n439) );
  NBUFFX2_HVT U176 ( .A(n256), .Y(n282) );
  MUX41X1_HVT U182 ( .A1(n568), .A3(n351), .A2(n404), .A4(n283), .S0(n233), 
        .S1(n255), .Y(n403) );
  MUX41X1_HVT U183 ( .A1(n325), .A3(n337), .A2(n288), .A4(n335), .S0(n253), 
        .S1(n241), .Y(n397) );
  MUX41X1_HVT U184 ( .A1(n394), .A3(n397), .A2(n390), .A4(n393), .S0(n276), 
        .S1(n247), .Y(n389) );
  MUX41X1_HVT U185 ( .A1(n463), .A3(n449), .A2(n457), .A4(n444), .S0(n258), 
        .S1(n247), .Y(out[3]) );
  MUX41X1_HVT U187 ( .A1(n413), .A3(n536), .A2(n327), .A4(n560), .S0(n233), 
        .S1(n241), .Y(n412) );
  XOR2X1_HVT U188 ( .A1(n255), .A2(n257), .Y(n535) );
  MUX41X1_HVT U190 ( .A1(n386), .A3(n387), .A2(n382), .A4(n385), .S0(n300), 
        .S1(n247), .Y(n381) );
  MUX41X1_HVT U191 ( .A1(n464), .A3(n466), .A2(n470), .A4(n469), .S0(n210), 
        .S1(n301), .Y(n463) );
  NAND2X0_HVT U192 ( .A1(n465), .A2(n259), .Y(n260) );
  NAND2X0_HVT U193 ( .A1(n579), .A2(n533), .Y(n261) );
  NAND2X0_HVT U194 ( .A1(n260), .A2(n261), .Y(n464) );
  INVX0_HVT U195 ( .A(n533), .Y(n259) );
  MUX21X2_HVT U196 ( .A1(n471), .A2(n481), .S0(in[6]), .Y(out[2]) );
  INVX0_HVT U198 ( .A(in[3]), .Y(n358) );
  MUX21X2_HVT U199 ( .A1(n267), .A2(n480), .S0(n535), .Y(n479) );
  MUX21X2_HVT U200 ( .A1(n329), .A2(n567), .S0(n275), .Y(n480) );
  INVX1_HVT U201 ( .A(n288), .Y(n356) );
  MUX21X1_HVT U202 ( .A1(n264), .A2(n239), .S0(n272), .Y(n446) );
  NBUFFX2_HVT U204 ( .A(n256), .Y(n281) );
  AND2X1_HVT U206 ( .A1(n281), .A2(n524), .Y(n262) );
  NBUFFX2_HVT U207 ( .A(n576), .Y(n288) );
  MUX21X1_HVT U209 ( .A1(n356), .A2(n359), .S0(in[5]), .Y(n528) );
  NBUFFX2_HVT U210 ( .A(n576), .Y(n289) );
  MUX21X1_HVT U211 ( .A1(n551), .A2(n468), .S0(n272), .Y(n466) );
  MUX21X1_HVT U213 ( .A1(n316), .A2(n357), .S0(in[5]), .Y(n513) );
  AND2X1_HVT U216 ( .A1(n290), .A2(n507), .Y(n263) );
  MUX21X1_HVT U217 ( .A1(n281), .A2(n359), .S0(n295), .Y(n574) );
  MUX21X1_HVT U219 ( .A1(n450), .A2(n451), .S0(in[5]), .Y(n449) );
  MUX21X1_HVT U221 ( .A1(n455), .A2(n454), .S0(n279), .Y(n451) );
  MUX21X1_HVT U222 ( .A1(n290), .A2(n282), .S0(n297), .Y(n541) );
  MUX21X1_HVT U223 ( .A1(n281), .A2(n284), .S0(n294), .Y(n476) );
  MUX21X1_HVT U224 ( .A1(n356), .A2(n232), .S0(n294), .Y(n404) );
  MUX21X1_HVT U225 ( .A1(n289), .A2(n240), .S0(n293), .Y(n545) );
  MUX21X1_HVT U226 ( .A1(n359), .A2(n282), .S0(n219), .Y(n416) );
  MUX21X1_HVT U227 ( .A1(n282), .A2(n356), .S0(n297), .Y(n484) );
  MUX21X1_HVT U228 ( .A1(n240), .A2(n357), .S0(n231), .Y(n364) );
  MUX21X1_HVT U229 ( .A1(n240), .A2(n284), .S0(n296), .Y(n504) );
  MUX21X1_HVT U230 ( .A1(n280), .A2(n240), .S0(n295), .Y(n367) );
  MUX21X1_HVT U231 ( .A1(n359), .A2(n356), .S0(n297), .Y(n544) );
  MUX21X1_HVT U232 ( .A1(n359), .A2(n280), .S0(n295), .Y(n548) );
  MUX21X1_HVT U233 ( .A1(n280), .A2(n232), .S0(n296), .Y(n542) );
  MUX21X1_HVT U234 ( .A1(n352), .A2(n287), .S0(n278), .Y(n443) );
  MUX21X1_HVT U235 ( .A1(n459), .A2(n460), .S0(n278), .Y(n458) );
  MUX21X1_HVT U236 ( .A1(n308), .A2(n331), .S0(n272), .Y(n460) );
  MUX21X1_HVT U237 ( .A1(n289), .A2(n287), .S0(n297), .Y(n491) );
  NAND2X0_HVT U238 ( .A1(n283), .A2(n358), .Y(n576) );
  MUX21X1_HVT U239 ( .A1(n356), .A2(n283), .S0(n296), .Y(n365) );
  INVX1_HVT U240 ( .A(n572), .Y(n357) );
  INVX1_HVT U241 ( .A(n291), .Y(n359) );
  MUX21X1_HVT U242 ( .A1(n307), .A2(n456), .S0(n274), .Y(n455) );
  MUX21X1_HVT U243 ( .A1(n283), .A2(n280), .S0(n295), .Y(n456) );
  NBUFFX2_HVT U244 ( .A(n579), .Y(n290) );
  MUX21X1_HVT U245 ( .A1(n358), .A2(n292), .S0(n297), .Y(n391) );
  MUX21X1_HVT U246 ( .A1(n291), .A2(n290), .S0(n231), .Y(n392) );
  XOR2X1_HVT U247 ( .A1(n295), .A2(n357), .Y(n537) );
  MUX21X1_HVT U248 ( .A1(n357), .A2(n356), .S0(n219), .Y(n563) );
  MUX21X1_HVT U249 ( .A1(n290), .A2(n287), .S0(n293), .Y(n567) );
  MUX21X1_HVT U250 ( .A1(n288), .A2(n292), .S0(n218), .Y(n486) );
  MUX21X1_HVT U251 ( .A1(n280), .A2(n359), .S0(n294), .Y(n571) );
  MUX21X1_HVT U252 ( .A1(n289), .A2(n280), .S0(n294), .Y(n570) );
  MUX21X1_HVT U253 ( .A1(n280), .A2(n284), .S0(n219), .Y(n388) );
  XNOR2X1_HVT U254 ( .A1(n288), .A2(n296), .Y(n264) );
  MUX21X1_HVT U255 ( .A1(n291), .A2(n287), .S0(n294), .Y(n551) );
  MUX21X1_HVT U256 ( .A1(n579), .A2(n283), .S0(n295), .Y(n371) );
  MUX21X1_HVT U257 ( .A1(n579), .A2(n289), .S0(n297), .Y(n363) );
  XNOR2X1_HVT U258 ( .A1(n291), .A2(n294), .Y(n265) );
  AND2X1_HVT U259 ( .A1(n296), .A2(n232), .Y(n266) );
  MUX21X1_HVT U260 ( .A1(n287), .A2(n280), .S0(n297), .Y(n369) );
  AND2X1_HVT U261 ( .A1(n292), .A2(n467), .Y(n267) );
  MUX21X1_HVT U262 ( .A1(n287), .A2(n283), .S0(n296), .Y(n509) );
  MUX21X1_HVT U263 ( .A1(n572), .A2(n292), .S0(n274), .Y(n453) );
  XOR2X1_HVT U264 ( .A1(n283), .A2(n296), .Y(n556) );
  NBUFFX2_HVT U265 ( .A(n303), .Y(n277) );
  NBUFFX2_HVT U266 ( .A(n303), .Y(n278) );
  NBUFFX2_HVT U267 ( .A(n358), .Y(n280) );
  NBUFFX2_HVT U268 ( .A(in[2]), .Y(n272) );
  NBUFFX2_HVT U269 ( .A(in[2]), .Y(n274) );
  NBUFFX2_HVT U270 ( .A(in[2]), .Y(n275) );
  NBUFFX2_HVT U271 ( .A(in[2]), .Y(n273) );
  NBUFFX2_HVT U272 ( .A(in[2]), .Y(n271) );
  MUX21X1_HVT U273 ( .A1(n281), .A2(n286), .S0(n293), .Y(n559) );
  MUX21X1_HVT U274 ( .A1(n478), .A2(n328), .S0(n274), .Y(n475) );
  MUX21X1_HVT U275 ( .A1(n395), .A2(n396), .S0(n273), .Y(n394) );
  MUX21X1_HVT U276 ( .A1(n494), .A2(n285), .S0(n278), .Y(n396) );
  MUX21X1_HVT U277 ( .A1(n517), .A2(n519), .S0(n273), .Y(n516) );
  XOR2X1_HVT U278 ( .A1(n294), .A2(n285), .Y(n534) );
  MUX21X1_HVT U279 ( .A1(n287), .A2(n282), .S0(n295), .Y(n473) );
  MUX21X1_HVT U280 ( .A1(n349), .A2(n357), .S0(n278), .Y(n428) );
  MUX21X1_HVT U281 ( .A1(n408), .A2(n407), .S0(n274), .Y(n406) );
  MUX21X1_HVT U282 ( .A1(n572), .A2(n347), .S0(n279), .Y(n408) );
  AND2X1_HVT U283 ( .A1(n282), .A2(n299), .Y(n268) );
  MUX21X1_HVT U284 ( .A1(n285), .A2(n356), .S0(n296), .Y(n543) );
  MUX21X1_HVT U285 ( .A1(n564), .A2(n330), .S0(n275), .Y(n445) );
  MUX21X1_HVT U286 ( .A1(n357), .A2(n232), .S0(n219), .Y(n413) );
  NAND2X0_HVT U287 ( .A1(n285), .A2(n284), .Y(n579) );
  NBUFFX2_HVT U288 ( .A(n360), .Y(n284) );
  NBUFFX2_HVT U289 ( .A(n580), .Y(n291) );
  MUX21X1_HVT U290 ( .A1(n232), .A2(n285), .S0(n231), .Y(n562) );
  MUX21X1_HVT U291 ( .A1(n332), .A2(n578), .S0(n273), .Y(n470) );
  MUX21X1_HVT U292 ( .A1(n423), .A2(n290), .S0(n269), .Y(n422) );
  MUX21X1_HVT U293 ( .A1(n544), .A2(n350), .S0(n277), .Y(n421) );
  MUX21X1_HVT U294 ( .A1(n578), .A2(n299), .S0(n273), .Y(n452) );
  MUX21X1_HVT U295 ( .A1(n529), .A2(n530), .S0(n277), .Y(n527) );
  MUX21X1_HVT U296 ( .A1(n286), .A2(n547), .S0(n301), .Y(n530) );
  XOR2X1_HVT U297 ( .A1(n219), .A2(n276), .Y(n539) );
  NBUFFX2_HVT U298 ( .A(n572), .Y(n287) );
  MUX21X1_HVT U299 ( .A1(n285), .A2(n357), .S0(n295), .Y(n368) );
  MUX21X1_HVT U300 ( .A1(n289), .A2(n286), .S0(n297), .Y(n573) );
  MUX21X1_HVT U301 ( .A1(n326), .A2(n552), .S0(n273), .Y(n448) );
  MUX21X1_HVT U302 ( .A1(n318), .A2(n299), .S0(in[5]), .Y(n515) );
  MUX21X1_HVT U303 ( .A1(n285), .A2(n283), .S0(n279), .Y(n489) );
  NBUFFX2_HVT U304 ( .A(n580), .Y(n292) );
  NBUFFX2_HVT U305 ( .A(n360), .Y(n283) );
  XNOR2X1_HVT U306 ( .A1(n253), .A2(n293), .Y(n269) );
  AND2X1_HVT U307 ( .A1(n280), .A2(n299), .Y(n270) );
  NBUFFX2_HVT U308 ( .A(in[5]), .Y(n301) );
  NBUFFX2_HVT U309 ( .A(in[5]), .Y(n300) );
  MUX21X1_HVT U310 ( .A1(n458), .A2(n461), .S0(n300), .Y(n457) );
  MUX21X1_HVT U311 ( .A1(n527), .A2(n531), .S0(n274), .Y(n526) );
  MUX21X1_HVT U312 ( .A1(n521), .A2(n523), .S0(n273), .Y(n520) );
  MUX21X1_HVT U313 ( .A1(n356), .A2(n245), .S0(n293), .Y(n550) );
  MUX21X1_HVT U314 ( .A1(n245), .A2(n240), .S0(n294), .Y(n370) );
  NAND2X0_HVT U315 ( .A1(in[4]), .A2(n358), .Y(n572) );
  NAND2X0_HVT U316 ( .A1(n286), .A2(in[4]), .Y(n580) );
  MUX21X1_HVT U317 ( .A1(n245), .A2(n359), .S0(n297), .Y(n546) );
  MUX21X1_HVT U318 ( .A1(n245), .A2(n357), .S0(n231), .Y(n564) );
  MUX21X1_HVT U319 ( .A1(n245), .A2(n290), .S0(n296), .Y(n561) );
  MUX21X1_HVT U320 ( .A1(n245), .A2(n287), .S0(n293), .Y(n362) );
  MUX21X1_HVT U321 ( .A1(n292), .A2(n245), .S0(n295), .Y(n554) );
  MUX21X1_HVT U322 ( .A1(n286), .A2(n245), .S0(n272), .Y(n465) );
  MUX21X1_HVT U323 ( .A1(n245), .A2(n292), .S0(n297), .Y(n361) );
  MUX21X1_HVT U324 ( .A1(n280), .A2(n245), .S0(n218), .Y(n552) );
  NBUFFX2_HVT U325 ( .A(in[3]), .Y(n285) );
  NBUFFX2_HVT U326 ( .A(in[3]), .Y(n286) );
  INVX0_HVT U327 ( .A(n560), .Y(n305) );
  INVX0_HVT U328 ( .A(n558), .Y(n306) );
  INVX0_HVT U329 ( .A(n549), .Y(n307) );
  INVX0_HVT U330 ( .A(n547), .Y(n308) );
  INVX0_HVT U331 ( .A(n410), .Y(n309) );
  INVX0_HVT U332 ( .A(n373), .Y(n310) );
  INVX0_HVT U333 ( .A(n578), .Y(n311) );
  INVX0_HVT U334 ( .A(n566), .Y(n312) );
  INVX0_HVT U335 ( .A(n577), .Y(n313) );
  INVX0_HVT U336 ( .A(n575), .Y(n314) );
  INVX0_HVT U337 ( .A(n574), .Y(n315) );
  INVX0_HVT U338 ( .A(n573), .Y(n316) );
  INVX0_HVT U339 ( .A(n571), .Y(n317) );
  INVX0_HVT U340 ( .A(n570), .Y(n318) );
  INVX0_HVT U341 ( .A(n567), .Y(n319) );
  INVX0_HVT U342 ( .A(n564), .Y(n320) );
  INVX0_HVT U343 ( .A(n563), .Y(n321) );
  INVX0_HVT U344 ( .A(n562), .Y(n322) );
  INVX0_HVT U345 ( .A(n556), .Y(n325) );
  INVX0_HVT U346 ( .A(n554), .Y(n326) );
  INVX0_HVT U347 ( .A(n551), .Y(n329) );
  INVX0_HVT U348 ( .A(n550), .Y(n330) );
  INVX0_HVT U349 ( .A(n548), .Y(n331) );
  INVX0_HVT U350 ( .A(n546), .Y(n332) );
  INVX0_HVT U351 ( .A(n544), .Y(n334) );
  INVX0_HVT U352 ( .A(n543), .Y(n335) );
  INVX0_HVT U353 ( .A(n542), .Y(n336) );
  INVX0_HVT U354 ( .A(n541), .Y(n337) );
  INVX0_HVT U355 ( .A(n540), .Y(n338) );
  INVX0_HVT U356 ( .A(n507), .Y(n339) );
  INVX0_HVT U357 ( .A(n467), .Y(n341) );
  INVX0_HVT U358 ( .A(n372), .Y(n342) );
  INVX0_HVT U359 ( .A(n524), .Y(n343) );
  INVX0_HVT U360 ( .A(n426), .Y(n344) );
  INVX0_HVT U361 ( .A(n371), .Y(n345) );
  INVX0_HVT U362 ( .A(n370), .Y(n346) );
  INVX0_HVT U363 ( .A(n368), .Y(n348) );
  INVX0_HVT U364 ( .A(n486), .Y(n350) );
  INVX0_HVT U365 ( .A(n476), .Y(n351) );
  INVX0_HVT U366 ( .A(n364), .Y(n353) );
  INVX0_HVT U367 ( .A(n363), .Y(n354) );
  INVX0_HVT U368 ( .A(n361), .Y(n355) );
endmodule

