
module Mix_Column ( in, out );
  input [127:0] in;
  output [127:0] out;
  wire   n3, n6, n8, n11, n12, n14, n15, n16, n18, n21, n22, n24, n25, n27,
         n28, n29, n30, n31, n32, n35, n37, n38, n39, n40, n42, n43, n44, n46,
         n48, n50, n52, n53, n54, n58, n60, n61, n63, n64, n66, n68, n69, n71,
         n74, n75, n77, n78, n80, n82, n84, n85, n86, n88, n89, n90, n92, n93,
         n94, n95, n96, n99, n100, n101, n102, n104, n105, n106, n108, n109,
         n111, n113, n115, n118, n119, n121, n122, n123, n126, n127, n130,
         n134, n140, n141, n144, n146, n147, n148, n149, n150, n151, n152,
         n154, n158, n159, n160, n162, n163, n168, n171, n176, n177, n178,
         n179, n180, n181, n183, n184, n186, n188, n189, n191, n193, n194,
         n199, n200, n202, n208, n210, n217, n218, n220, n1, n2, n4, n5, n7,
         n9, n10, n13, n17, n19, n20, n23, n26, n33, n34, n36, n41, n45, n47,
         n49, n51, n55, n56, n57, n59, n62, n65, n67, n70, n72, n73, n76, n79,
         n81, n83, n87, n91, n97, n98, n103, n107, n110, n112, n114, n116,
         n117, n120, n124, n125, n128, n129, n131, n132, n133, n135, n136,
         n137, n138, n139, n142, n143, n145, n153, n155, n156, n157, n161,
         n164, n165, n166, n167, n169, n170, n172, n174, n175, n182, n185,
         n187, n190, n192, n195, n196, n197, n198, n201, n203, n204, n205,
         n206, n207, n209, n211, n212, n213, n214, n215, n216, n219, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070;

  XNOR2X2_HVT U95 ( .A1(n409), .A2(n594), .Y(n101) );
  XNOR2X1_HVT U1 ( .A1(n681), .A2(n230), .Y(n236) );
  NBUFFX2_HVT U2 ( .A(n461), .Y(n1064) );
  INVX1_HVT U3 ( .A(in[43]), .Y(n1056) );
  NBUFFX2_HVT U4 ( .A(n1012), .Y(n779) );
  INVX1_HVT U5 ( .A(in[91]), .Y(n756) );
  INVX1_HVT U6 ( .A(in[115]), .Y(n701) );
  INVX1_HVT U7 ( .A(in[107]), .Y(n1040) );
  INVX1_HVT U8 ( .A(n498), .Y(n916) );
  NBUFFX2_HVT U9 ( .A(n417), .Y(n1062) );
  INVX1_HVT U10 ( .A(n964), .Y(n230) );
  INVX1_HVT U11 ( .A(n817), .Y(n429) );
  INVX1_HVT U12 ( .A(in[96]), .Y(n690) );
  INVX1_HVT U13 ( .A(n690), .Y(n450) );
  INVX1_HVT U14 ( .A(n117), .Y(n939) );
  INVX1_HVT U15 ( .A(n42), .Y(n960) );
  INVX0_HVT U16 ( .A(n56), .Y(n604) );
  INVX1_HVT U17 ( .A(n946), .Y(n947) );
  INVX0_HVT U18 ( .A(n101), .Y(n378) );
  INVX1_HVT U19 ( .A(n51), .Y(n964) );
  XOR2X1_HVT U20 ( .A1(n728), .A2(n739), .Y(n713) );
  XNOR2X1_HVT U21 ( .A1(n19), .A2(n439), .Y(n99) );
  INVX1_HVT U22 ( .A(n882), .Y(n259) );
  INVX1_HVT U23 ( .A(n972), .Y(n284) );
  INVX1_HVT U24 ( .A(n971), .Y(n821) );
  INVX1_HVT U25 ( .A(n318), .Y(n298) );
  INVX0_HVT U26 ( .A(n193), .Y(n677) );
  INVX0_HVT U27 ( .A(n181), .Y(n864) );
  XOR3X1_HVT U28 ( .A1(n27), .A2(n934), .A3(n504), .Y(out[96]) );
  INVX1_HVT U29 ( .A(n701), .Y(n702) );
  INVX0_HVT U30 ( .A(n11), .Y(n329) );
  INVX1_HVT U31 ( .A(in[48]), .Y(n11) );
  INVX1_HVT U32 ( .A(n524), .Y(n512) );
  INVX1_HVT U33 ( .A(n777), .Y(n778) );
  INVX1_HVT U34 ( .A(n832), .Y(n833) );
  AND2X1_HVT U35 ( .A1(n469), .A2(n142), .Y(n1) );
  INVX0_HVT U36 ( .A(n444), .Y(n1001) );
  AND2X1_HVT U37 ( .A1(n522), .A2(n523), .Y(n2) );
  AND2X1_HVT U38 ( .A1(n234), .A2(n233), .Y(n4) );
  AND2X1_HVT U39 ( .A1(n398), .A2(n399), .Y(n5) );
  INVX1_HVT U40 ( .A(in[45]), .Y(n406) );
  INVX1_HVT U41 ( .A(n871), .Y(n740) );
  INVX1_HVT U42 ( .A(in[122]), .Y(n977) );
  INVX1_HVT U43 ( .A(n1070), .Y(n45) );
  INVX1_HVT U44 ( .A(in[28]), .Y(n792) );
  INVX1_HVT U45 ( .A(in[121]), .Y(n1004) );
  INVX1_HVT U46 ( .A(n1003), .Y(n465) );
  INVX1_HVT U47 ( .A(n413), .Y(n244) );
  INVX1_HVT U48 ( .A(in[80]), .Y(n858) );
  INVX1_HVT U49 ( .A(n667), .Y(n855) );
  INVX1_HVT U50 ( .A(in[76]), .Y(n435) );
  INVX0_HVT U51 ( .A(n938), .Y(n432) );
  INVX1_HVT U52 ( .A(n436), .Y(n1052) );
  NAND2X0_HVT U53 ( .A1(n565), .A2(n970), .Y(n10) );
  NAND2X0_HVT U54 ( .A1(n7), .A2(n9), .Y(n13) );
  NAND2X0_HVT U55 ( .A1(n10), .A2(n13), .Y(n38) );
  INVX0_HVT U56 ( .A(n565), .Y(n7) );
  INVX0_HVT U57 ( .A(n87), .Y(n9) );
  AND2X1_HVT U58 ( .A1(n47), .A2(n49), .Y(n17) );
  XOR3X1_HVT U59 ( .A1(n17), .A2(n821), .A3(n229), .Y(out[111]) );
  INVX1_HVT U60 ( .A(n658), .Y(n917) );
  INVX1_HVT U61 ( .A(n507), .Y(n490) );
  INVX0_HVT U62 ( .A(in[47]), .Y(n379) );
  INVX1_HVT U63 ( .A(in[7]), .Y(n416) );
  INVX1_HVT U64 ( .A(n962), .Y(n825) );
  XOR3X2_HVT U65 ( .A1(n587), .A2(n928), .A3(n35), .Y(n919) );
  INVX1_HVT U66 ( .A(n658), .Y(n642) );
  INVX1_HVT U67 ( .A(in[94]), .Y(n424) );
  INVX1_HVT U68 ( .A(n667), .Y(n19) );
  XOR3X2_HVT U69 ( .A1(n129), .A2(n231), .A3(n515), .Y(out[58]) );
  INVX1_HVT U70 ( .A(in[11]), .Y(n968) );
  INVX1_HVT U71 ( .A(in[3]), .Y(n719) );
  INVX1_HVT U72 ( .A(in[97]), .Y(n619) );
  XNOR2X2_HVT U73 ( .A1(n426), .A2(n776), .Y(n160) );
  INVX0_HVT U74 ( .A(n426), .Y(n339) );
  INVX1_HVT U75 ( .A(in[9]), .Y(n426) );
  NAND2X0_HVT U76 ( .A1(n389), .A2(n23), .Y(n26) );
  NAND2X0_HVT U77 ( .A1(n20), .A2(n377), .Y(n33) );
  NAND2X0_HVT U78 ( .A1(n26), .A2(n33), .Y(n936) );
  INVX0_HVT U79 ( .A(n389), .Y(n20) );
  INVX0_HVT U80 ( .A(n377), .Y(n23) );
  NAND2X0_HVT U81 ( .A1(n421), .A2(n466), .Y(n34) );
  NAND2X0_HVT U82 ( .A1(n420), .A2(n465), .Y(n36) );
  NAND2X0_HVT U83 ( .A1(n34), .A2(n36), .Y(n40) );
  NAND2X0_HVT U84 ( .A1(n112), .A2(n1070), .Y(n47) );
  NAND2X0_HVT U85 ( .A1(n41), .A2(n45), .Y(n49) );
  INVX1_HVT U86 ( .A(n112), .Y(n41) );
  INVX0_HVT U87 ( .A(n962), .Y(n112) );
  INVX0_HVT U88 ( .A(n424), .Y(n389) );
  XOR3X2_HVT U89 ( .A1(n488), .A2(n883), .A3(n277), .Y(n1009) );
  INVX0_HVT U90 ( .A(n883), .Y(n601) );
  INVX1_HVT U91 ( .A(in[41]), .Y(n883) );
  XNOR2X2_HVT U92 ( .A1(n51), .A2(n371), .Y(n122) );
  OR2X1_HVT U93 ( .A1(n582), .A2(n926), .Y(n878) );
  INVX1_HVT U94 ( .A(in[83]), .Y(n870) );
  INVX1_HVT U96 ( .A(n902), .Y(n1034) );
  INVX1_HVT U97 ( .A(in[59]), .Y(n908) );
  INVX1_HVT U98 ( .A(in[79]), .Y(n830) );
  INVX0_HVT U99 ( .A(n601), .Y(n264) );
  XOR3X2_HVT U100 ( .A1(n277), .A2(n1060), .A3(n759), .Y(n922) );
  INVX1_HVT U101 ( .A(in[73]), .Y(n643) );
  INVX1_HVT U102 ( .A(n777), .Y(n594) );
  INVX0_HVT U103 ( .A(n962), .Y(n745) );
  INVX1_HVT U104 ( .A(n664), .Y(n117) );
  INVX0_HVT U105 ( .A(n379), .Y(n51) );
  INVX0_HVT U106 ( .A(n420), .Y(n55) );
  INVX1_HVT U107 ( .A(in[52]), .Y(n926) );
  INVX1_HVT U108 ( .A(in[19]), .Y(n924) );
  INVX1_HVT U109 ( .A(n127), .Y(n812) );
  INVX1_HVT U110 ( .A(n825), .Y(n1014) );
  INVX1_HVT U111 ( .A(in[112]), .Y(n3) );
  INVX0_HVT U112 ( .A(in[2]), .Y(n857) );
  INVX0_HVT U113 ( .A(n1065), .Y(n682) );
  INVX1_HVT U114 ( .A(in[85]), .Y(n676) );
  NAND2X0_HVT U115 ( .A1(n301), .A2(n302), .Y(n56) );
  INVX1_HVT U116 ( .A(in[81]), .Y(n420) );
  XOR3X2_HVT U117 ( .A1(n619), .A2(n690), .A3(n355), .Y(n839) );
  INVX1_HVT U118 ( .A(n670), .Y(n624) );
  INVX1_HVT U119 ( .A(in[15]), .Y(n930) );
  INVX1_HVT U120 ( .A(in[11]), .Y(n1042) );
  INVX1_HVT U121 ( .A(in[32]), .Y(n12) );
  INVX1_HVT U122 ( .A(n669), .Y(n664) );
  NAND2X0_HVT U123 ( .A1(n473), .A2(n248), .Y(n59) );
  NAND2X0_HVT U124 ( .A1(n57), .A2(n598), .Y(n62) );
  NAND2X0_HVT U125 ( .A1(n59), .A2(n62), .Y(n163) );
  INVX0_HVT U126 ( .A(n473), .Y(n57) );
  INVX0_HVT U127 ( .A(n163), .Y(n946) );
  INVX1_HVT U128 ( .A(in[16]), .Y(n286) );
  INVX1_HVT U129 ( .A(n926), .Y(n927) );
  NBUFFX2_HVT U130 ( .A(in[127]), .Y(n65) );
  INVX1_HVT U131 ( .A(in[35]), .Y(n1012) );
  INVX1_HVT U132 ( .A(n811), .Y(n707) );
  INVX1_HVT U133 ( .A(n917), .Y(n114) );
  INVX1_HVT U134 ( .A(in[39]), .Y(n658) );
  INVX1_HVT U135 ( .A(in[40]), .Y(n488) );
  XNOR2X2_HVT U136 ( .A1(n1053), .A2(n444), .Y(n53) );
  INVX1_HVT U137 ( .A(in[72]), .Y(n691) );
  XOR3X2_HVT U138 ( .A1(n627), .A2(n722), .A3(n67), .Y(n126) );
  AND2X1_HVT U139 ( .A1(n878), .A2(n879), .Y(n67) );
  INVX1_HVT U140 ( .A(in[123]), .Y(n669) );
  INVX1_HVT U141 ( .A(in[57]), .Y(n757) );
  INVX1_HVT U142 ( .A(in[119]), .Y(n962) );
  INVX1_HVT U143 ( .A(n938), .Y(n817) );
  INVX1_HVT U144 ( .A(n745), .Y(n746) );
  INVX1_HVT U145 ( .A(n1041), .Y(n891) );
  XOR2X1_HVT U146 ( .A1(n7), .A2(n422), .Y(n71) );
  INVX1_HVT U147 ( .A(n801), .Y(n966) );
  INVX0_HVT U148 ( .A(n1062), .Y(n629) );
  INVX1_HVT U149 ( .A(n629), .Y(n506) );
  INVX1_HVT U150 ( .A(n313), .Y(n979) );
  INVX1_HVT U151 ( .A(in[99]), .Y(n623) );
  XNOR2X1_HVT U152 ( .A1(n707), .A2(n521), .Y(n63) );
  INVX1_HVT U153 ( .A(n974), .Y(n550) );
  INVX1_HVT U154 ( .A(n1056), .Y(n1057) );
  INVX1_HVT U155 ( .A(n728), .Y(n546) );
  INVX1_HVT U156 ( .A(in[70]), .Y(n809) );
  INVX1_HVT U157 ( .A(in[93]), .Y(n941) );
  INVX1_HVT U158 ( .A(n312), .Y(n245) );
  INVX1_HVT U159 ( .A(n420), .Y(n421) );
  XNOR2X1_HVT U160 ( .A1(n455), .A2(n740), .Y(n39) );
  INVX1_HVT U161 ( .A(n932), .Y(n686) );
  INVX0_HVT U162 ( .A(n354), .Y(n136) );
  INVX1_HVT U163 ( .A(n446), .Y(n785) );
  INVX1_HVT U164 ( .A(n1014), .Y(n818) );
  INVX0_HVT U165 ( .A(n605), .Y(n973) );
  INVX1_HVT U166 ( .A(n100), .Y(n515) );
  XOR3X1_HVT U167 ( .A1(n53), .A2(n245), .A3(n161), .Y(out[69]) );
  XOR2X1_HVT U168 ( .A1(n476), .A2(in[88]), .Y(n920) );
  INVX1_HVT U169 ( .A(n133), .Y(n489) );
  INVX1_HVT U170 ( .A(n348), .Y(n294) );
  INVX1_HVT U171 ( .A(n29), .Y(n395) );
  INVX1_HVT U172 ( .A(n50), .Y(n716) );
  XNOR2X1_HVT U173 ( .A1(n460), .A2(n628), .Y(n15) );
  INVX0_HVT U174 ( .A(in[38]), .Y(n978) );
  INVX0_HVT U175 ( .A(n978), .Y(n828) );
  INVX0_HVT U176 ( .A(in[110]), .Y(n782) );
  INVX0_HVT U177 ( .A(n977), .Y(n732) );
  INVX1_HVT U178 ( .A(n447), .Y(n356) );
  INVX0_HVT U179 ( .A(n974), .Y(n411) );
  INVX1_HVT U180 ( .A(n107), .Y(n945) );
  INVX0_HVT U181 ( .A(n213), .Y(n107) );
  INVX1_HVT U182 ( .A(n788), .Y(n780) );
  INVX0_HVT U183 ( .A(n908), .Y(n798) );
  INVX1_HVT U184 ( .A(n287), .Y(n473) );
  INVX0_HVT U185 ( .A(n331), .Y(n1035) );
  INVX0_HVT U186 ( .A(n211), .Y(n212) );
  INVX1_HVT U187 ( .A(n292), .Y(n293) );
  INVX0_HVT U188 ( .A(n858), .Y(n476) );
  INVX0_HVT U189 ( .A(n435), .Y(n436) );
  INVX0_HVT U190 ( .A(n858), .Y(n70) );
  INVX1_HVT U191 ( .A(n70), .Y(n72) );
  INVX0_HVT U192 ( .A(n1004), .Y(n97) );
  INVX0_HVT U193 ( .A(in[104]), .Y(n491) );
  NBUFFX2_HVT U194 ( .A(in[47]), .Y(n277) );
  XOR3X2_HVT U195 ( .A1(n277), .A2(n819), .A3(n820), .Y(n127) );
  INVX0_HVT U196 ( .A(n39), .Y(n575) );
  INVX1_HVT U197 ( .A(n133), .Y(n492) );
  INVX1_HVT U198 ( .A(n76), .Y(n934) );
  INVX1_HVT U199 ( .A(n821), .Y(n76) );
  INVX0_HVT U200 ( .A(n877), .Y(n880) );
  NAND2X0_HVT U201 ( .A1(n205), .A2(n1004), .Y(n73) );
  NAND2X0_HVT U202 ( .A1(n308), .A2(n309), .Y(n79) );
  INVX0_HVT U203 ( .A(n786), .Y(n787) );
  INVX1_HVT U204 ( .A(n956), .Y(n531) );
  INVX0_HVT U205 ( .A(n782), .Y(n318) );
  INVX1_HVT U206 ( .A(n1011), .Y(n508) );
  NAND2X0_HVT U207 ( .A1(n337), .A2(n785), .Y(n697) );
  INVX1_HVT U208 ( .A(n340), .Y(n314) );
  INVX1_HVT U209 ( .A(n582), .Y(n877) );
  INVX1_HVT U210 ( .A(n337), .Y(n153) );
  INVX0_HVT U211 ( .A(in[53]), .Y(n728) );
  XOR3X2_HVT U212 ( .A1(n108), .A2(n739), .A3(n227), .Y(out[53]) );
  OR2X1_HVT U213 ( .A1(n995), .A2(n214), .Y(n737) );
  INVX1_HVT U214 ( .A(n214), .Y(n6) );
  INVX1_HVT U215 ( .A(n434), .Y(n187) );
  INVX0_HVT U216 ( .A(n612), .Y(n952) );
  INVX0_HVT U217 ( .A(n748), .Y(n612) );
  INVX1_HVT U218 ( .A(in[6]), .Y(n81) );
  INVX1_HVT U219 ( .A(n902), .Y(n956) );
  INVX1_HVT U220 ( .A(n211), .Y(n87) );
  INVX1_HVT U221 ( .A(in[125]), .Y(n261) );
  INVX0_HVT U222 ( .A(n671), .Y(n451) );
  INVX0_HVT U223 ( .A(n501), .Y(n459) );
  INVX0_HVT U224 ( .A(n454), .Y(n455) );
  XOR3X2_HVT U225 ( .A1(n180), .A2(n686), .A3(n215), .Y(out[110]) );
  INVX0_HVT U226 ( .A(n534), .Y(n535) );
  INVX1_HVT U227 ( .A(n534), .Y(n516) );
  XOR2X2_HVT U228 ( .A1(in[78]), .A2(in[70]), .Y(n29) );
  INVX1_HVT U229 ( .A(in[61]), .Y(n571) );
  INVX1_HVT U230 ( .A(n358), .Y(n83) );
  INVX0_HVT U231 ( .A(n264), .Y(n338) );
  INVX0_HVT U232 ( .A(n247), .Y(n882) );
  INVX1_HVT U233 ( .A(n445), .Y(n132) );
  INVX0_HVT U234 ( .A(n445), .Y(n422) );
  INVX1_HVT U235 ( .A(in[120]), .Y(n441) );
  INVX1_HVT U236 ( .A(n5), .Y(n540) );
  INVX1_HVT U237 ( .A(in[66]), .Y(n454) );
  INVX0_HVT U238 ( .A(n695), .Y(n258) );
  INVX1_HVT U239 ( .A(in[98]), .Y(n980) );
  XOR3X2_HVT U240 ( .A1(n188), .A2(n726), .A3(n24), .Y(out[114]) );
  INVX1_HVT U241 ( .A(n787), .Y(n91) );
  INVX0_HVT U242 ( .A(in[126]), .Y(n786) );
  XOR3X2_HVT U243 ( .A1(n97), .A2(n1069), .A3(n145), .Y(n25) );
  INVX1_HVT U244 ( .A(in[67]), .Y(n881) );
  INVX1_HVT U245 ( .A(n25), .Y(n365) );
  INVX0_HVT U246 ( .A(n418), .Y(n387) );
  INVX1_HVT U247 ( .A(n238), .Y(n138) );
  XOR2X1_HVT U248 ( .A1(n320), .A2(n840), .Y(n551) );
  INVX1_HVT U249 ( .A(n5), .Y(n98) );
  AND2X1_HVT U250 ( .A1(n165), .A2(n166), .Y(n103) );
  INVX0_HVT U251 ( .A(n213), .Y(n214) );
  INVX0_HVT U252 ( .A(n8), .Y(n957) );
  INVX1_HVT U253 ( .A(n791), .Y(n853) );
  INVX1_HVT U254 ( .A(n274), .Y(n255) );
  INVX1_HVT U255 ( .A(n675), .Y(n110) );
  INVX1_HVT U256 ( .A(n742), .Y(n675) );
  INVX0_HVT U257 ( .A(in[29]), .Y(n742) );
  INVX1_HVT U258 ( .A(n808), .Y(n397) );
  NBUFFX2_HVT U259 ( .A(n273), .Y(n1068) );
  INVX0_HVT U260 ( .A(n123), .Y(n876) );
  INVX0_HVT U261 ( .A(n443), .Y(n308) );
  INVX1_HVT U262 ( .A(n171), .Y(n899) );
  INVX0_HVT U263 ( .A(n416), .Y(n381) );
  INVX1_HVT U264 ( .A(in[0]), .Y(n14) );
  INVX1_HVT U265 ( .A(in[37]), .Y(n910) );
  INVX0_HVT U266 ( .A(n658), .Y(n659) );
  INVX1_HVT U267 ( .A(in[118]), .Y(n223) );
  INVX1_HVT U268 ( .A(n930), .Y(n461) );
  NAND2X0_HVT U269 ( .A1(n411), .A2(n741), .Y(n116) );
  XOR2X2_HVT U270 ( .A1(n490), .A2(in[20]), .Y(n118) );
  INVX0_HVT U271 ( .A(in[117]), .Y(n672) );
  INVX0_HVT U272 ( .A(n1058), .Y(n819) );
  INVX0_HVT U273 ( .A(n991), .Y(n434) );
  INVX0_HVT U274 ( .A(n791), .Y(n1011) );
  INVX1_HVT U275 ( .A(n593), .Y(n332) );
  INVX0_HVT U276 ( .A(in[69]), .Y(n816) );
  AND2X1_HVT U277 ( .A1(n263), .A2(n262), .Y(n120) );
  INVX0_HVT U278 ( .A(n1066), .Y(n860) );
  OR2X1_HVT U279 ( .A1(n978), .A2(n170), .Y(n399) );
  INVX1_HVT U280 ( .A(n443), .Y(n440) );
  INVX0_HVT U281 ( .A(n87), .Y(n996) );
  INVX1_HVT U282 ( .A(in[86]), .Y(n991) );
  INVX0_HVT U283 ( .A(n1000), .Y(n873) );
  INVX0_HVT U284 ( .A(n941), .Y(n174) );
  INVX0_HVT U285 ( .A(n406), .Y(n124) );
  XOR2X2_HVT U286 ( .A1(n972), .A2(n875), .Y(n125) );
  INVX1_HVT U287 ( .A(in[101]), .Y(n972) );
  NAND2X0_HVT U288 ( .A1(n413), .A2(n415), .Y(n128) );
  INVX1_HVT U289 ( .A(n967), .Y(n292) );
  INVX0_HVT U290 ( .A(n721), .Y(n685) );
  INVX1_HVT U291 ( .A(n721), .Y(n722) );
  INVX1_HVT U292 ( .A(n58), .Y(n383) );
  OR2X1_HVT U293 ( .A1(n348), .A2(n382), .Y(n296) );
  INVX1_HVT U294 ( .A(n249), .Y(n616) );
  INVX0_HVT U295 ( .A(in[49]), .Y(n518) );
  XNOR2X2_HVT U296 ( .A1(n855), .A2(n1058), .Y(n129) );
  INVX1_HVT U297 ( .A(n567), .Y(n517) );
  INVX1_HVT U298 ( .A(n18), .Y(n554) );
  INVX1_HVT U299 ( .A(in[54]), .Y(n501) );
  INVX1_HVT U300 ( .A(n653), .Y(n654) );
  INVX1_HVT U301 ( .A(n724), .Y(n313) );
  INVX1_HVT U302 ( .A(in[27]), .Y(n724) );
  INVX0_HVT U303 ( .A(n14), .Y(n981) );
  INVX0_HVT U304 ( .A(n518), .Y(n731) );
  XOR2X2_HVT U305 ( .A1(n421), .A2(n465), .Y(n131) );
  INVX0_HVT U306 ( .A(n930), .Y(n460) );
  INVX1_HVT U307 ( .A(n586), .Y(n485) );
  XOR3X2_HVT U308 ( .A1(n169), .A2(n817), .A3(n132), .Y(n37) );
  INVX0_HVT U309 ( .A(n627), .Y(n291) );
  INVX0_HVT U310 ( .A(n272), .Y(n133) );
  INVX0_HVT U311 ( .A(n272), .Y(n273) );
  INVX1_HVT U312 ( .A(n623), .Y(n167) );
  NAND2X0_HVT U313 ( .A1(n223), .A2(n224), .Y(n135) );
  XOR3X2_HVT U314 ( .A1(n489), .A2(n1040), .A3(n136), .Y(n1055) );
  INVX1_HVT U315 ( .A(n660), .Y(n224) );
  INVX0_HVT U316 ( .A(n921), .Y(n892) );
  INVX1_HVT U317 ( .A(n921), .Y(n714) );
  INVX1_HVT U318 ( .A(in[64]), .Y(n8) );
  INVX0_HVT U319 ( .A(n984), .Y(n384) );
  INVX1_HVT U320 ( .A(in[1]), .Y(n775) );
  INVX1_HVT U321 ( .A(n424), .Y(n319) );
  INVX0_HVT U322 ( .A(n1067), .Y(n1000) );
  INVX1_HVT U323 ( .A(n1067), .Y(n921) );
  INVX0_HVT U324 ( .A(n667), .Y(n937) );
  INVX1_HVT U325 ( .A(n580), .Y(n581) );
  INVX0_HVT U326 ( .A(n580), .Y(n388) );
  INVX1_HVT U327 ( .A(n746), .Y(n656) );
  IBUFFX2_HVT U328 ( .A(n622), .Y(n260) );
  INVX0_HVT U329 ( .A(n511), .Y(n137) );
  XOR2X2_HVT U330 ( .A1(n436), .A2(n587), .Y(n50) );
  INVX0_HVT U331 ( .A(n250), .Y(n139) );
  INVX0_HVT U332 ( .A(n371), .Y(n250) );
  INVX1_HVT U333 ( .A(n808), .Y(n741) );
  XNOR2X2_HVT U334 ( .A1(n816), .A2(n935), .Y(n31) );
  INVX0_HVT U335 ( .A(n816), .Y(n593) );
  INVX0_HVT U336 ( .A(n935), .Y(n312) );
  INVX1_HVT U337 ( .A(in[67]), .Y(n169) );
  INVX1_HVT U338 ( .A(in[90]), .Y(n565) );
  NAND2X0_HVT U339 ( .A1(n338), .A2(n467), .Y(n142) );
  INVX1_HVT U340 ( .A(n583), .Y(n599) );
  INVX0_HVT U341 ( .A(n66), .Y(n704) );
  XNOR2X2_HVT U342 ( .A1(n931), .A2(n476), .Y(n143) );
  INVX1_HVT U343 ( .A(n143), .Y(n350) );
  INVX0_HVT U344 ( .A(n719), .Y(n720) );
  INVX1_HVT U345 ( .A(in[68]), .Y(n1053) );
  INVX1_HVT U346 ( .A(n183), .Y(n709) );
  NAND2X0_HVT U347 ( .A1(n442), .A2(n153), .Y(n155) );
  NAND2X0_HVT U348 ( .A1(n145), .A2(n337), .Y(n156) );
  NAND2X0_HVT U349 ( .A1(n155), .A2(n156), .Y(n217) );
  INVX0_HVT U350 ( .A(n442), .Y(n145) );
  INVX1_HVT U351 ( .A(n441), .Y(n442) );
  INVX0_HVT U352 ( .A(n3), .Y(n337) );
  NAND2X0_HVT U353 ( .A1(n73), .A2(n206), .Y(n157) );
  INVX1_HVT U354 ( .A(n830), .Y(n694) );
  INVX1_HVT U355 ( .A(n1024), .Y(n986) );
  INVX1_HVT U356 ( .A(in[105]), .Y(n618) );
  NAND2X0_HVT U357 ( .A1(n511), .A2(n167), .Y(n514) );
  INVX1_HVT U358 ( .A(in[26]), .Y(n583) );
  INVX1_HVT U359 ( .A(n1053), .Y(n431) );
  INVX1_HVT U360 ( .A(in[63]), .Y(n788) );
  NBUFFX2_HVT U361 ( .A(n30), .Y(n161) );
  XOR2X1_HVT U362 ( .A1(n450), .A2(n442), .Y(n197) );
  INVX1_HVT U363 ( .A(n1049), .Y(n767) );
  NAND2X0_HVT U364 ( .A1(n558), .A2(n420), .Y(n165) );
  NAND2X0_HVT U365 ( .A1(n164), .A2(n55), .Y(n166) );
  NAND2X0_HVT U366 ( .A1(n165), .A2(n166), .Y(n253) );
  INVX0_HVT U367 ( .A(n644), .Y(n164) );
  INVX0_HVT U368 ( .A(n830), .Y(n246) );
  INVX0_HVT U369 ( .A(in[46]), .Y(n170) );
  NAND2X0_HVT U370 ( .A1(n295), .A2(n296), .Y(n172) );
  INVX0_HVT U371 ( .A(in[56]), .Y(n777) );
  NBUFFX2_HVT U372 ( .A(in[31]), .Y(n1065) );
  INVX1_HVT U373 ( .A(n798), .Y(n528) );
  INVX1_HVT U374 ( .A(n69), .Y(n1044) );
  INVX1_HVT U375 ( .A(n216), .Y(n574) );
  NBUFFX2_HVT U376 ( .A(n273), .Y(n228) );
  XOR3X2_HVT U377 ( .A1(n31), .A2(n174), .A3(n716), .Y(out[85]) );
  INVX1_HVT U378 ( .A(in[51]), .Y(n175) );
  INVX0_HVT U379 ( .A(in[51]), .Y(n951) );
  INVX1_HVT U380 ( .A(n893), .Y(n182) );
  INVX0_HVT U381 ( .A(n893), .Y(n428) );
  INVX1_HVT U382 ( .A(n134), .Y(n865) );
  INVX1_HVT U383 ( .A(n92), .Y(n885) );
  NBUFFX2_HVT U384 ( .A(in[37]), .Y(n185) );
  INVX0_HVT U385 ( .A(in[22]), .Y(n781) );
  INVX1_HVT U386 ( .A(n1016), .Y(n481) );
  INVX1_HVT U387 ( .A(n893), .Y(n267) );
  NBUFFX2_HVT U388 ( .A(n627), .Y(n190) );
  INVX1_HVT U389 ( .A(n691), .Y(n480) );
  INVX0_HVT U390 ( .A(n691), .Y(n641) );
  INVX1_HVT U391 ( .A(n1048), .Y(n894) );
  INVX0_HVT U392 ( .A(n1040), .Y(n348) );
  INVX0_HVT U393 ( .A(n1054), .Y(n355) );
  NAND2X0_HVT U394 ( .A1(n655), .A2(n889), .Y(n192) );
  INVX1_HVT U395 ( .A(n891), .Y(n232) );
  NBUFFX2_HVT U396 ( .A(n923), .Y(n195) );
  INVX0_HVT U397 ( .A(n12), .Y(n923) );
  INVX1_HVT U398 ( .A(n873), .Y(n196) );
  INVX0_HVT U399 ( .A(n775), .Y(n776) );
  INVX1_HVT U400 ( .A(n1027), .Y(n913) );
  XOR3X2_HVT U401 ( .A1(n369), .A2(n656), .A3(n197), .Y(out[112]) );
  INVX1_HVT U402 ( .A(n870), .Y(n928) );
  XNOR2X2_HVT U403 ( .A1(n917), .A2(n349), .Y(n198) );
  NAND2X0_HVT U404 ( .A1(n322), .A2(n321), .Y(n201) );
  INVX0_HVT U405 ( .A(in[30]), .Y(n723) );
  XOR2X2_HVT U406 ( .A1(n110), .A2(n595), .Y(n94) );
  INVX1_HVT U407 ( .A(n65), .Y(n832) );
  INVX0_HVT U408 ( .A(n1051), .Y(n589) );
  INVX1_HVT U409 ( .A(n1022), .Y(n733) );
  NAND2X0_HVT U410 ( .A1(n346), .A2(n347), .Y(n203) );
  INVX1_HVT U411 ( .A(n720), .Y(n568) );
  NBUFFX2_HVT U412 ( .A(n675), .Y(n204) );
  INVX1_HVT U413 ( .A(n68), .Y(n1043) );
  XOR3X2_HVT U414 ( .A1(n188), .A2(n282), .A3(n189), .Y(out[122]) );
  NAND2X0_HVT U415 ( .A1(n357), .A2(in[121]), .Y(n206) );
  NAND2X0_HVT U416 ( .A1(n205), .A2(n1004), .Y(n207) );
  NAND2X0_HVT U417 ( .A1(n207), .A2(n206), .Y(n21) );
  INVX0_HVT U418 ( .A(n357), .Y(n205) );
  NAND2X0_HVT U419 ( .A1(n116), .A2(n302), .Y(n150) );
  NAND2X0_HVT U420 ( .A1(n492), .A2(n446), .Y(n209) );
  INVX1_HVT U421 ( .A(n30), .Y(n373) );
  INVX0_HVT U422 ( .A(n507), .Y(n889) );
  INVX1_HVT U423 ( .A(in[74]), .Y(n871) );
  INVX1_HVT U424 ( .A(in[99]), .Y(n524) );
  INVX1_HVT U425 ( .A(in[78]), .Y(n430) );
  INVX1_HVT U426 ( .A(n438), .Y(n402) );
  INVX0_HVT U427 ( .A(in[95]), .Y(n211) );
  INVX0_HVT U428 ( .A(in[87]), .Y(n213) );
  INVX0_HVT U429 ( .A(n822), .Y(n391) );
  NAND2X0_HVT U430 ( .A1(n225), .A2(n226), .Y(n215) );
  XNOR2X2_HVT U431 ( .A1(n131), .A2(n445), .Y(n216) );
  INVX0_HVT U432 ( .A(n724), .Y(n725) );
  INVX1_HVT U433 ( .A(n12), .Y(n349) );
  INVX1_HVT U434 ( .A(in[50]), .Y(n1060) );
  INVX1_HVT U435 ( .A(n200), .Y(n607) );
  INVX1_HVT U436 ( .A(n757), .Y(n342) );
  INVX1_HVT U437 ( .A(n876), .Y(n359) );
  INVX0_HVT U438 ( .A(in[18]), .Y(n967) );
  NAND2X0_HVT U439 ( .A1(n239), .A2(n240), .Y(n219) );
  INVX0_HVT U440 ( .A(in[17]), .Y(n418) );
  INVX1_HVT U441 ( .A(in[33]), .Y(n622) );
  NAND2X0_HVT U442 ( .A1(n716), .A2(n283), .Y(n221) );
  XNOR2X2_HVT U443 ( .A1(n431), .A2(n435), .Y(n35) );
  INVX0_HVT U444 ( .A(n397), .Y(n222) );
  INVX1_HVT U445 ( .A(n287), .Y(n943) );
  INVX1_HVT U446 ( .A(n286), .Y(n287) );
  INVX1_HVT U447 ( .A(n1051), .Y(n902) );
  NAND2X0_HVT U448 ( .A1(in[118]), .A2(n660), .Y(n225) );
  NAND2X0_HVT U449 ( .A1(n223), .A2(n224), .Y(n226) );
  NAND2X0_HVT U450 ( .A1(n135), .A2(n225), .Y(n831) );
  INVX0_HVT U451 ( .A(n786), .Y(n660) );
  INVX1_HVT U452 ( .A(n924), .Y(n893) );
  INVX1_HVT U453 ( .A(n1060), .Y(n231) );
  AND2X1_HVT U454 ( .A1(n265), .A2(n266), .Y(n227) );
  INVX1_HVT U455 ( .A(n800), .Y(n772) );
  NAND2X0_HVT U456 ( .A1(n299), .A2(n300), .Y(n229) );
  NAND2X0_HVT U457 ( .A1(n1060), .A2(n891), .Y(n233) );
  NAND2X0_HVT U458 ( .A1(n231), .A2(n1041), .Y(n234) );
  NAND2X0_HVT U459 ( .A1(n234), .A2(n233), .Y(n130) );
  INVX1_HVT U460 ( .A(n940), .Y(n905) );
  OR2X1_HVT U461 ( .A1(n406), .A2(n910), .Y(n266) );
  XOR3X2_HVT U462 ( .A1(n519), .A2(n235), .A3(n191), .Y(out[121]) );
  NAND2X0_HVT U463 ( .A1(n242), .A2(n621), .Y(n235) );
  XOR3X2_HVT U464 ( .A1(n359), .A2(n828), .A3(n236), .Y(out[39]) );
  INVX1_HVT U465 ( .A(n643), .Y(n644) );
  INVX1_HVT U466 ( .A(n840), .Y(n595) );
  INVX0_HVT U467 ( .A(n792), .Y(n752) );
  INVX0_HVT U468 ( .A(n792), .Y(n687) );
  INVX1_HVT U469 ( .A(n586), .Y(n587) );
  XOR3X2_HVT U470 ( .A1(n1013), .A2(n833), .A3(n939), .Y(n1029) );
  NAND2X0_HVT U471 ( .A1(n138), .A2(n387), .Y(n239) );
  NAND2X0_HVT U472 ( .A1(n237), .A2(n238), .Y(n240) );
  NAND2X0_HVT U473 ( .A1(n239), .A2(n240), .Y(n168) );
  INVX1_HVT U474 ( .A(n387), .Y(n237) );
  INVX0_HVT U475 ( .A(n426), .Y(n238) );
  INVX1_HVT U476 ( .A(n364), .Y(n241) );
  INVX0_HVT U477 ( .A(in[25]), .Y(n990) );
  NAND2X0_HVT U478 ( .A1(n464), .A2(n83), .Y(n242) );
  AND2X1_HVT U479 ( .A1(n718), .A2(n717), .Y(n243) );
  XOR3X2_HVT U480 ( .A1(n1042), .A2(n267), .A3(n293), .Y(n412) );
  INVX0_HVT U481 ( .A(in[77]), .Y(n935) );
  INVX0_HVT U482 ( .A(n830), .Y(n247) );
  INVX1_HVT U483 ( .A(n1012), .Y(n627) );
  INVX0_HVT U484 ( .A(n598), .Y(n248) );
  XOR3X2_HVT U485 ( .A1(n268), .A2(n780), .A3(n559), .Y(n249) );
  XOR3X2_HVT U486 ( .A1(n6), .A2(n421), .A3(n72), .Y(n823) );
  NAND2X0_HVT U487 ( .A1(n409), .A2(n139), .Y(n251) );
  NAND2X0_HVT U488 ( .A1(n788), .A2(n250), .Y(n252) );
  NAND2X0_HVT U489 ( .A1(n252), .A2(n251), .Y(n104) );
  NBUFFX2_HVT U490 ( .A(n924), .Y(n668) );
  INVX1_HVT U491 ( .A(n487), .Y(n415) );
  INVX0_HVT U492 ( .A(in[42]), .Y(n1058) );
  INVX1_HVT U493 ( .A(n370), .Y(n309) );
  INVX1_HVT U494 ( .A(n1054), .Y(n971) );
  INVX1_HVT U495 ( .A(n1029), .Y(n710) );
  NAND2X0_HVT U496 ( .A1(n24), .A2(n274), .Y(n256) );
  NAND2X0_HVT U497 ( .A1(n254), .A2(n255), .Y(n257) );
  NAND2X0_HVT U498 ( .A1(n256), .A2(n257), .Y(n427) );
  INVX0_HVT U499 ( .A(n24), .Y(n254) );
  INVX0_HVT U500 ( .A(n427), .Y(n366) );
  INVX0_HVT U501 ( .A(n416), .Y(n417) );
  XNOR2X2_HVT U502 ( .A1(n432), .A2(n454), .Y(n671) );
  INVX1_HVT U503 ( .A(n141), .Y(n845) );
  INVX1_HVT U504 ( .A(in[43]), .Y(n961) );
  XOR3X2_HVT U505 ( .A1(n74), .A2(n259), .A3(n920), .Y(out[72]) );
  INVX1_HVT U506 ( .A(n431), .Y(n343) );
  INVX1_HVT U507 ( .A(in[24]), .Y(n520) );
  XOR3X2_HVT U508 ( .A1(n659), .A2(n923), .A3(n260), .Y(n929) );
  INVX1_HVT U509 ( .A(n1017), .Y(n645) );
  INVX0_HVT U510 ( .A(n968), .Y(n948) );
  INVX1_HVT U511 ( .A(n908), .Y(n909) );
  INVX0_HVT U512 ( .A(n909), .Y(n559) );
  XOR3X2_HVT U513 ( .A1(n936), .A2(n245), .A3(n395), .Y(out[86]) );
  INVX1_HVT U514 ( .A(n305), .Y(n278) );
  NAND2X0_HVT U515 ( .A1(n261), .A2(n672), .Y(n262) );
  NAND2X0_HVT U516 ( .A1(in[117]), .A2(in[125]), .Y(n263) );
  NAND2X0_HVT U517 ( .A1(n263), .A2(n262), .Y(n179) );
  INVX1_HVT U518 ( .A(n888), .Y(n703) );
  INVX1_HVT U519 ( .A(n461), .Y(n1047) );
  NAND2X0_HVT U520 ( .A1(n910), .A2(n406), .Y(n265) );
  NAND2X0_HVT U521 ( .A1(n266), .A2(n265), .Y(n89) );
  INVX0_HVT U522 ( .A(n902), .Y(n268) );
  INVX1_HVT U523 ( .A(n140), .Y(n987) );
  XOR3X2_HVT U524 ( .A1(n111), .A2(n406), .A3(n713), .Y(out[37]) );
  INVX0_HVT U525 ( .A(n922), .Y(n762) );
  NAND2X0_HVT U526 ( .A1(n282), .A2(n701), .Y(n270) );
  NAND2X0_HVT U527 ( .A1(n269), .A2(n702), .Y(n271) );
  NAND2X0_HVT U528 ( .A1(n270), .A2(n271), .Y(n382) );
  INVX0_HVT U529 ( .A(n282), .Y(n269) );
  INVX1_HVT U530 ( .A(n1037), .Y(n613) );
  INVX0_HVT U531 ( .A(n599), .Y(n600) );
  INVX0_HVT U532 ( .A(in[111]), .Y(n272) );
  XOR2X2_HVT U533 ( .A1(n450), .A2(n355), .Y(n274) );
  NAND2X0_HVT U534 ( .A1(n1002), .A2(n212), .Y(n275) );
  NAND2X0_HVT U535 ( .A1(n470), .A2(n9), .Y(n276) );
  NAND2X0_HVT U536 ( .A1(n275), .A2(n276), .Y(n999) );
  XOR3X2_HVT U537 ( .A1(n179), .A2(n284), .A3(n278), .Y(out[109]) );
  INVX1_HVT U538 ( .A(n52), .Y(n835) );
  NAND2X0_HVT U539 ( .A1(n396), .A2(n752), .Y(n280) );
  NAND2X0_HVT U540 ( .A1(n279), .A2(n792), .Y(n281) );
  NAND2X0_HVT U541 ( .A1(n280), .A2(n281), .Y(n151) );
  INVX0_HVT U542 ( .A(n396), .Y(n279) );
  INVX0_HVT U543 ( .A(in[20]), .Y(n396) );
  XOR3X2_HVT U544 ( .A1(n93), .A2(n910), .A3(n713), .Y(out[45]) );
  INVX0_HVT U545 ( .A(n653), .Y(n282) );
  INVX0_HVT U546 ( .A(n598), .Y(n708) );
  INVX1_HVT U547 ( .A(n953), .Y(n842) );
  INVX1_HVT U548 ( .A(n516), .Y(n345) );
  XNOR2X1_HVT U549 ( .A1(n524), .A2(n832), .Y(n838) );
  INVX1_HVT U550 ( .A(n317), .Y(n152) );
  INVX1_HVT U551 ( .A(n598), .Y(n811) );
  AND2X1_HVT U552 ( .A1(n761), .A2(n760), .Y(n283) );
  INVX1_HVT U553 ( .A(n676), .Y(n377) );
  XNOR2X2_HVT U554 ( .A1(n8), .A2(n1067), .Y(n74) );
  INVX0_HVT U555 ( .A(n682), .Y(n663) );
  INVX1_HVT U556 ( .A(n1066), .Y(n521) );
  INVX0_HVT U557 ( .A(in[103]), .Y(n1054) );
  NBUFFX2_HVT U558 ( .A(n875), .Y(n285) );
  INVX1_HVT U559 ( .A(n982), .Y(n482) );
  XOR3X2_HVT U560 ( .A1(n525), .A2(n565), .A3(n999), .Y(n1022) );
  NAND2X0_HVT U561 ( .A1(n79), .A2(n310), .Y(n288) );
  INVX0_HVT U562 ( .A(n643), .Y(n558) );
  INVX1_HVT U563 ( .A(in[88]), .Y(n995) );
  XNOR2X1_HVT U564 ( .A1(n258), .A2(n1004), .Y(n189) );
  INVX1_HVT U565 ( .A(in[58]), .Y(n1041) );
  XOR3X2_HVT U566 ( .A1(n60), .A2(n957), .A3(n911), .Y(out[80]) );
  XOR2X2_HVT U567 ( .A1(n444), .A2(n485), .Y(n32) );
  NAND2X0_HVT U568 ( .A1(n370), .A2(n376), .Y(n290) );
  INVX1_HVT U569 ( .A(n109), .Y(n912) );
  NAND2X0_HVT U570 ( .A1(n382), .A2(n348), .Y(n295) );
  NAND2X0_HVT U571 ( .A1(n295), .A2(n296), .Y(n186) );
  INVX0_HVT U572 ( .A(n186), .Y(n650) );
  NAND2X0_HVT U573 ( .A1(n496), .A2(n497), .Y(n297) );
  INVX0_HVT U574 ( .A(n945), .Y(n495) );
  NAND2X0_HVT U575 ( .A1(n932), .A2(n782), .Y(n299) );
  NAND2X0_HVT U576 ( .A1(in[102]), .A2(n318), .Y(n300) );
  NAND2X0_HVT U577 ( .A1(n300), .A2(n299), .Y(n178) );
  INVX1_HVT U578 ( .A(in[102]), .Y(n932) );
  INVX1_HVT U579 ( .A(n942), .Y(n678) );
  XOR3X2_HVT U580 ( .A1(n977), .A2(n818), .A3(n838), .Y(n975) );
  NAND2X0_HVT U581 ( .A1(n411), .A2(n741), .Y(n301) );
  NAND2X0_HVT U582 ( .A1(n974), .A2(n808), .Y(n302) );
  XOR3X2_HVT U583 ( .A1(n1056), .A2(n819), .A3(n190), .Y(n113) );
  NAND2X0_HVT U584 ( .A1(n303), .A2(n192), .Y(n950) );
  AND2X1_HVT U585 ( .A1(n890), .A2(n948), .Y(n303) );
  AND2X1_HVT U586 ( .A1(n949), .A2(n950), .Y(n304) );
  NAND2X0_HVT U587 ( .A1(n290), .A2(n361), .Y(n305) );
  NBUFFX2_HVT U588 ( .A(n307), .Y(n306) );
  INVX0_HVT U589 ( .A(n672), .Y(n307) );
  INVX0_HVT U590 ( .A(n945), .Y(n931) );
  NAND2X0_HVT U591 ( .A1(n443), .A2(n370), .Y(n310) );
  NAND2X0_HVT U592 ( .A1(n308), .A2(n309), .Y(n311) );
  NAND2X0_HVT U593 ( .A1(n310), .A2(n311), .Y(n199) );
  INVX0_HVT U594 ( .A(in[23]), .Y(n598) );
  INVX1_HVT U595 ( .A(n975), .Y(n649) );
  INVX1_HVT U596 ( .A(in[82]), .Y(n445) );
  NAND2X0_HVT U597 ( .A1(n356), .A2(n340), .Y(n315) );
  NAND2X0_HVT U598 ( .A1(n447), .A2(n314), .Y(n316) );
  NAND2X0_HVT U599 ( .A1(n316), .A2(n315), .Y(out[93]) );
  INVX1_HVT U600 ( .A(n1026), .Y(n866) );
  XOR2X2_HVT U601 ( .A1(n389), .A2(n246), .Y(n75) );
  XOR3X2_HVT U602 ( .A1(n313), .A2(n708), .A3(n663), .Y(n317) );
  XOR3X2_HVT U603 ( .A1(n61), .A2(n40), .A3(n829), .Y(out[73]) );
  XOR2X2_HVT U604 ( .A1(n972), .A2(n875), .Y(n180) );
  INVX1_HVT U605 ( .A(n731), .Y(n467) );
  XNOR2X2_HVT U606 ( .A1(n388), .A2(n558), .Y(n44) );
  INVX1_HVT U607 ( .A(n194), .Y(n849) );
  INVX0_HVT U608 ( .A(n781), .Y(n390) );
  XOR3X2_HVT U609 ( .A1(n977), .A2(n670), .A3(n372), .Y(n18) );
  XNOR2X2_HVT U610 ( .A1(n991), .A2(n319), .Y(n423) );
  NAND2X0_HVT U611 ( .A1(n781), .A2(n723), .Y(n321) );
  NAND2X0_HVT U612 ( .A1(in[22]), .A2(n320), .Y(n322) );
  NAND2X0_HVT U613 ( .A1(n321), .A2(n322), .Y(n78) );
  INVX0_HVT U614 ( .A(n723), .Y(n320) );
  NAND2X0_HVT U615 ( .A1(n925), .A2(n324), .Y(n325) );
  NAND2X0_HVT U616 ( .A1(n323), .A2(n802), .Y(n326) );
  NAND2X0_HVT U617 ( .A1(n325), .A2(n326), .Y(n158) );
  INVX0_HVT U618 ( .A(n925), .Y(n323) );
  INVX0_HVT U619 ( .A(n802), .Y(n324) );
  INVX1_HVT U620 ( .A(n408), .Y(n505) );
  INVX1_HVT U621 ( .A(in[51]), .Y(n1050) );
  XOR3X1_HVT U622 ( .A1(n821), .A2(n376), .A3(n181), .Y(n1049) );
  NAND2X0_HVT U623 ( .A1(n642), .A2(n230), .Y(n327) );
  NAND2X0_HVT U624 ( .A1(n964), .A2(n114), .Y(n328) );
  NAND2X0_HVT U625 ( .A1(n327), .A2(n328), .Y(n86) );
  INVX1_HVT U626 ( .A(in[24]), .Y(n541) );
  XNOR2X2_HVT U627 ( .A1(n32), .A2(n23), .Y(n340) );
  XOR3X2_HVT U628 ( .A1(n967), .A2(n811), .A3(n330), .Y(n985) );
  AND2X1_HVT U629 ( .A1(n499), .A2(n500), .Y(n330) );
  XNOR2X2_HVT U630 ( .A1(n622), .A2(n342), .Y(n119) );
  XOR3X2_HVT U631 ( .A1(n655), .A2(n550), .A3(n94), .Y(out[5]) );
  INVX0_HVT U632 ( .A(n870), .Y(n331) );
  XOR3X2_HVT U633 ( .A1(n423), .A2(n332), .A3(n333), .Y(out[70]) );
  AND2X1_HVT U634 ( .A1(n448), .A2(n449), .Y(n333) );
  INVX1_HVT U635 ( .A(n919), .Y(n562) );
  NAND2X0_HVT U636 ( .A1(n410), .A2(n876), .Y(n335) );
  NAND2X0_HVT U637 ( .A1(n359), .A2(n334), .Y(n336) );
  NAND2X0_HVT U638 ( .A1(n336), .A2(n335), .Y(n400) );
  INVX0_HVT U639 ( .A(n410), .Y(n334) );
  XNOR2X2_HVT U640 ( .A1(n618), .A2(n695), .Y(n24) );
  INVX1_HVT U641 ( .A(n1032), .Y(n834) );
  XOR3X2_HVT U642 ( .A1(n968), .A2(n1064), .A3(n151), .Y(n176) );
  NBUFFX2_HVT U643 ( .A(n460), .Y(n1063) );
  INVX0_HVT U644 ( .A(n857), .Y(n802) );
  XOR3X2_HVT U645 ( .A1(n779), .A2(n642), .A3(n203), .Y(n140) );
  XOR3X2_HVT U646 ( .A1(n969), .A2(n16), .A3(n15), .Y(out[9]) );
  INVX1_HVT U647 ( .A(n702), .Y(n363) );
  XOR3X2_HVT U648 ( .A1(n857), .A2(n725), .A3(n341), .Y(n194) );
  AND2X1_HVT U649 ( .A1(n569), .A2(n570), .Y(n341) );
  INVX0_HVT U650 ( .A(n996), .Y(n970) );
  INVX1_HVT U651 ( .A(n37), .Y(n638) );
  XOR3X2_HVT U652 ( .A1(n288), .A2(n261), .A3(n125), .Y(out[117]) );
  XNOR2X2_HVT U653 ( .A1(n801), .A2(n980), .Y(n188) );
  INVX0_HVT U654 ( .A(n450), .Y(n344) );
  NAND2X0_HVT U655 ( .A1(n345), .A2(n927), .Y(n346) );
  NAND2X0_HVT U656 ( .A1(n926), .A2(n516), .Y(n347) );
  NAND2X0_HVT U657 ( .A1(n346), .A2(n347), .Y(n108) );
  NAND2X0_HVT U658 ( .A1(n401), .A2(n143), .Y(n351) );
  NAND2X0_HVT U659 ( .A1(n351), .A2(n352), .Y(out[81]) );
  NAND2X0_HVT U660 ( .A1(n353), .A2(n385), .Y(n352) );
  AND2X1_HVT U661 ( .A1(n386), .A2(n350), .Y(n353) );
  XOR3X2_HVT U662 ( .A1(n423), .A2(n6), .A3(n28), .Y(out[95]) );
  INVX0_HVT U663 ( .A(in[10]), .Y(n925) );
  INVX0_HVT U664 ( .A(n31), .Y(n447) );
  NBUFFX2_HVT U665 ( .A(n933), .Y(n354) );
  INVX0_HVT U666 ( .A(in[106]), .Y(n933) );
  INVX1_HVT U667 ( .A(n719), .Y(n854) );
  INVX0_HVT U668 ( .A(n1061), .Y(n567) );
  INVX0_HVT U669 ( .A(n819), .Y(n439) );
  INVX1_HVT U670 ( .A(n380), .Y(n799) );
  NBUFFX2_HVT U671 ( .A(n619), .Y(n357) );
  INVX0_HVT U672 ( .A(n357), .Y(n358) );
  INVX1_HVT U673 ( .A(n175), .Y(n545) );
  XOR2X2_HVT U674 ( .A1(n364), .A2(n776), .Y(n148) );
  INVX1_HVT U675 ( .A(n990), .Y(n364) );
  NAND2X0_HVT U676 ( .A1(in[100]), .A2(n425), .Y(n361) );
  NAND2X0_HVT U677 ( .A1(n822), .A2(n360), .Y(n362) );
  NAND2X0_HVT U678 ( .A1(n361), .A2(n362), .Y(n184) );
  INVX0_HVT U679 ( .A(n425), .Y(n360) );
  INVX1_HVT U680 ( .A(n976), .Y(n813) );
  XOR3X2_HVT U681 ( .A1(n184), .A2(n440), .A3(n363), .Y(n183) );
  NAND2X0_HVT U682 ( .A1(n25), .A2(n427), .Y(n367) );
  NAND2X0_HVT U683 ( .A1(n365), .A2(n366), .Y(n368) );
  NAND2X0_HVT U684 ( .A1(n368), .A2(n367), .Y(out[97]) );
  INVX0_HVT U685 ( .A(n86), .Y(n413) );
  NAND2X0_HVT U686 ( .A1(n209), .A2(n494), .Y(n369) );
  XOR3X2_HVT U687 ( .A1(n168), .A2(n600), .A3(n158), .Y(out[18]) );
  INVX0_HVT U688 ( .A(n425), .Y(n370) );
  NBUFFX2_HVT U689 ( .A(n488), .Y(n371) );
  INVX0_HVT U690 ( .A(in[55]), .Y(n1051) );
  XOR3X2_HVT U691 ( .A1(n1050), .A2(n589), .A3(n859), .Y(n96) );
  XNOR2X2_HVT U692 ( .A1(n1047), .A2(n1062), .Y(n146) );
  INVX1_HVT U693 ( .A(n933), .Y(n801) );
  NAND2X0_HVT U694 ( .A1(n596), .A2(n597), .Y(n372) );
  NAND2X0_HVT U695 ( .A1(n434), .A2(n30), .Y(n374) );
  NAND2X0_HVT U696 ( .A1(n373), .A2(n187), .Y(n375) );
  NAND2X0_HVT U697 ( .A1(n375), .A2(n374), .Y(n433) );
  INVX0_HVT U698 ( .A(n433), .Y(n392) );
  INVX1_HVT U699 ( .A(n391), .Y(n376) );
  INVX0_HVT U700 ( .A(in[100]), .Y(n822) );
  XNOR2X1_HVT U701 ( .A1(n1034), .A2(n329), .Y(n105) );
  XOR3X2_HVT U702 ( .A1(n585), .A2(n114), .A3(n378), .Y(out[32]) );
  INVX0_HVT U703 ( .A(n113), .Y(n763) );
  XNOR2X2_HVT U704 ( .A1(n1040), .A2(n370), .Y(n380) );
  NBUFFX2_HVT U705 ( .A(n417), .Y(n1061) );
  INVX1_HVT U706 ( .A(in[124]), .Y(n1021) );
  NAND2X0_HVT U707 ( .A1(n384), .A2(n58), .Y(n385) );
  NAND2X0_HVT U708 ( .A1(n984), .A2(n383), .Y(n386) );
  NAND2X0_HVT U709 ( .A1(n385), .A2(n386), .Y(n401) );
  XOR2X2_HVT U710 ( .A1(n581), .A2(n465), .Y(n58) );
  INVX0_HVT U711 ( .A(in[91]), .Y(n1002) );
  INVX0_HVT U712 ( .A(in[65]), .Y(n580) );
  XNOR2X2_HVT U713 ( .A1(n1021), .A2(n391), .Y(n202) );
  XOR3X2_HVT U714 ( .A1(n78), .A2(n751), .A3(n604), .Y(out[14]) );
  XOR3X2_HVT U715 ( .A1(n132), .A2(n247), .A3(n1028), .Y(n54) );
  NAND2X0_HVT U716 ( .A1(n395), .A2(n433), .Y(n393) );
  NAND2X0_HVT U717 ( .A1(n392), .A2(n29), .Y(n394) );
  NAND2X0_HVT U718 ( .A1(n394), .A2(n393), .Y(out[94]) );
  XOR3X2_HVT U719 ( .A1(n396), .A2(n182), .A3(n154), .Y(n1037) );
  XOR3X2_HVT U720 ( .A1(n154), .A2(n397), .A3(n94), .Y(out[13]) );
  INVX1_HVT U721 ( .A(n412), .Y(n1036) );
  NAND2X0_HVT U722 ( .A1(n978), .A2(n170), .Y(n398) );
  NAND2X0_HVT U723 ( .A1(n398), .A2(n399), .Y(n410) );
  XNOR2X2_HVT U724 ( .A1(n400), .A2(n114), .Y(out[47]) );
  INVX1_HVT U725 ( .A(n408), .Y(n409) );
  NAND2X0_HVT U726 ( .A1(n437), .A2(n438), .Y(n403) );
  NAND2X0_HVT U727 ( .A1(n404), .A2(n403), .Y(out[63]) );
  NAND2X0_HVT U728 ( .A1(n405), .A2(n128), .Y(n404) );
  AND2X1_HVT U729 ( .A1(n414), .A2(n402), .Y(n405) );
  XOR3X2_HVT U730 ( .A1(n407), .A2(n185), .A3(n438), .Y(out[38]) );
  AND2X1_HVT U731 ( .A1(n572), .A2(n573), .Y(n407) );
  XNOR2X2_HVT U732 ( .A1(n622), .A2(n264), .Y(n102) );
  INVX0_HVT U733 ( .A(in[63]), .Y(n408) );
  INVX1_HVT U734 ( .A(n176), .Y(n632) );
  XOR3X2_HVT U735 ( .A1(n169), .A2(n817), .A3(n871), .Y(n953) );
  INVX0_HVT U736 ( .A(in[13]), .Y(n974) );
  INVX0_HVT U737 ( .A(n202), .Y(n795) );
  NAND2X0_HVT U738 ( .A1(n487), .A2(n86), .Y(n414) );
  NAND2X0_HVT U739 ( .A1(n128), .A2(n414), .Y(n437) );
  XOR3X2_HVT U740 ( .A1(n56), .A2(n595), .A3(n151), .Y(out[29]) );
  XNOR2X2_HVT U741 ( .A1(n14), .A2(n1061), .Y(n42) );
  XOR3X2_HVT U742 ( .A1(n159), .A2(n160), .A3(n963), .Y(out[25]) );
  INVX0_HVT U743 ( .A(in[4]), .Y(n791) );
  XNOR2X2_HVT U744 ( .A1(n419), .A2(n990), .Y(n16) );
  XNOR2X2_HVT U745 ( .A1(n941), .A2(n676), .Y(n30) );
  INVX1_HVT U746 ( .A(n418), .Y(n419) );
  XNOR2X1_HVT U747 ( .A1(n663), .A2(n390), .Y(n566) );
  XOR2X1_HVT U748 ( .A1(n292), .A2(n583), .Y(n149) );
  INVX0_HVT U749 ( .A(in[108]), .Y(n425) );
  XNOR2X2_HVT U750 ( .A1(n440), .A2(n1021), .Y(n181) );
  INVX0_HVT U751 ( .A(n215), .Y(n210) );
  XNOR2X2_HVT U752 ( .A1(n441), .A2(n65), .Y(n27) );
  INVX1_HVT U753 ( .A(in[75]), .Y(n938) );
  XNOR2X2_HVT U754 ( .A1(n766), .A2(n501), .Y(n438) );
  XOR3X2_HVT U755 ( .A1(n4), .A2(n439), .A3(n602), .Y(out[34]) );
  NBUFFX2_HVT U756 ( .A(in[127]), .Y(n1070) );
  XOR3X2_HVT U757 ( .A1(n701), .A2(n560), .A3(n348), .Y(n1025) );
  INVX0_HVT U758 ( .A(in[116]), .Y(n443) );
  INVX1_HVT U759 ( .A(n27), .Y(n519) );
  NBUFFX2_HVT U760 ( .A(in[92]), .Y(n444) );
  INVX1_HVT U761 ( .A(n491), .Y(n446) );
  XNOR2X1_HVT U762 ( .A1(n873), .A2(n246), .Y(n28) );
  XOR3X2_HVT U763 ( .A1(n599), .A2(n708), .A3(n994), .Y(n1048) );
  INVX0_HVT U764 ( .A(n665), .Y(n666) );
  XOR3X2_HVT U765 ( .A1(n927), .A2(n951), .A3(n93), .Y(n92) );
  INVX1_HVT U766 ( .A(n1025), .Y(n555) );
  NAND2X0_HVT U767 ( .A1(in[78]), .A2(n941), .Y(n448) );
  NAND2X0_HVT U768 ( .A1(n430), .A2(n174), .Y(n449) );
  INVX1_HVT U769 ( .A(n806), .Y(n1031) );
  NAND2X0_HVT U770 ( .A1(n873), .A2(n671), .Y(n452) );
  NAND2X0_HVT U771 ( .A1(n451), .A2(n196), .Y(n453) );
  NAND2X0_HVT U772 ( .A1(n453), .A2(n452), .Y(n82) );
  INVX0_HVT U773 ( .A(n82), .Y(n734) );
  NAND2X0_HVT U774 ( .A1(n758), .A2(n518), .Y(n457) );
  NAND2X0_HVT U775 ( .A1(n955), .A2(n456), .Y(n458) );
  NAND2X0_HVT U776 ( .A1(n457), .A2(n458), .Y(n100) );
  INVX0_HVT U777 ( .A(n518), .Y(n456) );
  XOR3X2_HVT U778 ( .A1(n98), .A2(n459), .A3(n88), .Y(out[62]) );
  NAND2X0_HVT U779 ( .A1(n250), .A2(in[48]), .Y(n462) );
  NAND2X0_HVT U780 ( .A1(n139), .A2(n11), .Y(n463) );
  NAND2X0_HVT U781 ( .A1(n462), .A2(n463), .Y(n585) );
  INVX1_HVT U782 ( .A(n1055), .Y(n803) );
  INVX0_HVT U783 ( .A(n618), .Y(n464) );
  INVX1_HVT U784 ( .A(n465), .Y(n466) );
  INVX0_HVT U785 ( .A(in[89]), .Y(n1003) );
  NAND2X0_HVT U786 ( .A1(n338), .A2(n467), .Y(n468) );
  NAND2X0_HVT U787 ( .A1(n264), .A2(n731), .Y(n469) );
  NAND2X0_HVT U788 ( .A1(n468), .A2(n469), .Y(n115) );
  NAND2X0_HVT U789 ( .A1(n1002), .A2(n945), .Y(n471) );
  NAND2X0_HVT U790 ( .A1(n470), .A2(n931), .Y(n472) );
  NAND2X0_HVT U791 ( .A1(n471), .A2(n472), .Y(n1028) );
  INVX0_HVT U792 ( .A(n1002), .Y(n470) );
  NAND2X0_HVT U793 ( .A1(n542), .A2(n287), .Y(n474) );
  NAND2X0_HVT U794 ( .A1(n943), .A2(n520), .Y(n475) );
  NAND2X0_HVT U795 ( .A1(n475), .A2(n474), .Y(n1033) );
  INVX0_HVT U796 ( .A(n541), .Y(n542) );
  NAND2X0_HVT U797 ( .A1(n72), .A2(n641), .Y(n478) );
  NAND2X0_HVT U798 ( .A1(n477), .A2(n476), .Y(n479) );
  NAND2X0_HVT U799 ( .A1(n479), .A2(n478), .Y(n85) );
  INVX0_HVT U800 ( .A(n480), .Y(n477) );
  NAND2X0_HVT U801 ( .A1(n982), .A2(n1016), .Y(n483) );
  NAND2X0_HVT U802 ( .A1(n481), .A2(n482), .Y(n484) );
  NAND2X0_HVT U803 ( .A1(n484), .A2(n483), .Y(out[4]) );
  XOR3X2_HVT U804 ( .A1(n979), .A2(n687), .A3(n118), .Y(n1016) );
  XOR3X2_HVT U805 ( .A1(n89), .A2(n828), .A3(n438), .Y(out[46]) );
  INVX1_HVT U806 ( .A(n1015), .Y(n637) );
  INVX1_HVT U807 ( .A(n669), .Y(n670) );
  INVX0_HVT U808 ( .A(in[60]), .Y(n665) );
  NBUFFX2_HVT U809 ( .A(n531), .Y(n487) );
  INVX1_HVT U810 ( .A(n1018), .Y(n633) );
  NAND2X0_HVT U811 ( .A1(n492), .A2(n446), .Y(n493) );
  NAND2X0_HVT U812 ( .A1(n491), .A2(n133), .Y(n494) );
  NAND2X0_HVT U813 ( .A1(n493), .A2(n494), .Y(n208) );
  INVX1_HVT U814 ( .A(n455), .Y(n869) );
  NAND2X0_HVT U815 ( .A1(n945), .A2(n996), .Y(n496) );
  NAND2X0_HVT U816 ( .A1(n107), .A2(n212), .Y(n497) );
  NAND2X0_HVT U817 ( .A1(n497), .A2(n496), .Y(n64) );
  XOR3X2_HVT U818 ( .A1(n567), .A2(n568), .A3(n663), .Y(n982) );
  NAND2X0_HVT U819 ( .A1(n313), .A2(n854), .Y(n499) );
  NAND2X0_HVT U820 ( .A1(n498), .A2(n979), .Y(n500) );
  INVX0_HVT U821 ( .A(n720), .Y(n498) );
  NAND2X0_HVT U822 ( .A1(n501), .A2(n505), .Y(n502) );
  NAND2X0_HVT U823 ( .A1(n408), .A2(n459), .Y(n503) );
  NAND2X0_HVT U824 ( .A1(n503), .A2(n502), .Y(n106) );
  AND2X1_HVT U825 ( .A1(n697), .A2(n698), .Y(n504) );
  INVX0_HVT U826 ( .A(in[21]), .Y(n840) );
  INVX1_HVT U827 ( .A(n1010), .Y(n768) );
  NAND2X0_HVT U828 ( .A1(n508), .A2(n490), .Y(n509) );
  NAND2X0_HVT U829 ( .A1(n507), .A2(n1011), .Y(n510) );
  NAND2X0_HVT U830 ( .A1(n509), .A2(n510), .Y(n154) );
  INVX0_HVT U831 ( .A(in[12]), .Y(n507) );
  XOR2X2_HVT U832 ( .A1(n246), .A2(n480), .Y(n61) );
  NAND2X0_HVT U833 ( .A1(n623), .A2(n137), .Y(n513) );
  NAND2X0_HVT U834 ( .A1(n513), .A2(n514), .Y(n807) );
  INVX0_HVT U835 ( .A(n980), .Y(n511) );
  INVX1_HVT U836 ( .A(n538), .Y(n549) );
  INVX1_HVT U837 ( .A(n1030), .Y(n846) );
  INVX0_HVT U838 ( .A(in[34]), .Y(n954) );
  NAND2X0_HVT U839 ( .A1(n542), .A2(n860), .Y(n522) );
  NAND2X0_HVT U840 ( .A1(n520), .A2(n1066), .Y(n523) );
  NAND2X0_HVT U841 ( .A1(n522), .A2(n523), .Y(n159) );
  XNOR2X2_HVT U842 ( .A1(n248), .A2(n541), .Y(n536) );
  XOR3X2_HVT U843 ( .A1(n1000), .A2(n881), .A3(n869), .Y(n69) );
  NAND2X0_HVT U844 ( .A1(n470), .A2(n928), .Y(n526) );
  NAND2X0_HVT U845 ( .A1(n756), .A2(n525), .Y(n527) );
  NAND2X0_HVT U846 ( .A1(n527), .A2(n526), .Y(n872) );
  INVX0_HVT U847 ( .A(n331), .Y(n525) );
  NAND2X0_HVT U848 ( .A1(n909), .A2(n884), .Y(n529) );
  NAND2X0_HVT U849 ( .A1(n1050), .A2(n528), .Y(n530) );
  NAND2X0_HVT U850 ( .A1(n530), .A2(n529), .Y(n820) );
  INVX0_HVT U851 ( .A(n1050), .Y(n884) );
  NAND2X0_HVT U852 ( .A1(n528), .A2(n268), .Y(n532) );
  NAND2X0_HVT U853 ( .A1(n531), .A2(n798), .Y(n533) );
  NAND2X0_HVT U854 ( .A1(n533), .A2(n532), .Y(n759) );
  INVX1_HVT U855 ( .A(n96), .Y(n771) );
  INVX0_HVT U856 ( .A(in[62]), .Y(n766) );
  INVX0_HVT U857 ( .A(n1019), .Y(n1006) );
  INVX0_HVT U858 ( .A(in[44]), .Y(n534) );
  XOR3X2_HVT U859 ( .A1(n536), .A2(n981), .A3(n15), .Y(out[16]) );
  XOR3X2_HVT U860 ( .A1(n540), .A2(n124), .A3(n537), .Y(out[54]) );
  AND2X1_HVT U861 ( .A1(n730), .A2(n729), .Y(n537) );
  INVX1_HVT U862 ( .A(n54), .Y(n841) );
  XOR3X1_HVT U863 ( .A1(n746), .A2(n654), .A3(n539), .Y(n538) );
  NAND2X0_HVT U864 ( .A1(n626), .A2(n625), .Y(n539) );
  INVX0_HVT U865 ( .A(n1059), .Y(n1013) );
  INVX0_HVT U866 ( .A(in[14]), .Y(n748) );
  XOR3X2_HVT U867 ( .A1(n664), .A2(n560), .A3(n199), .Y(n1019) );
  XOR3X2_HVT U868 ( .A1(n1), .A2(n891), .A3(n99), .Y(out[50]) );
  NAND2X0_HVT U869 ( .A1(in[118]), .A2(n45), .Y(n543) );
  NAND2X0_HVT U870 ( .A1(n223), .A2(n833), .Y(n544) );
  NAND2X0_HVT U871 ( .A1(n543), .A2(n544), .Y(n715) );
  NAND2X0_HVT U872 ( .A1(n728), .A2(n571), .Y(n547) );
  NAND2X0_HVT U873 ( .A1(n546), .A2(n739), .Y(n548) );
  NAND2X0_HVT U874 ( .A1(n547), .A2(n548), .Y(n88) );
  XOR3X2_HVT U875 ( .A1(n897), .A2(n550), .A3(n551), .Y(out[22]) );
  INVX0_HVT U876 ( .A(in[114]), .Y(n653) );
  NAND2X0_HVT U877 ( .A1(n909), .A2(n505), .Y(n552) );
  NAND2X0_HVT U878 ( .A1(n788), .A2(n528), .Y(n553) );
  NAND2X0_HVT U879 ( .A1(n553), .A2(n552), .Y(n1020) );
  NAND2X0_HVT U880 ( .A1(n1025), .A2(n18), .Y(n556) );
  NAND2X0_HVT U881 ( .A1(n554), .A2(n555), .Y(n557) );
  NAND2X0_HVT U882 ( .A1(n557), .A2(n556), .Y(out[99]) );
  INVX1_HVT U883 ( .A(n985), .Y(n898) );
  XOR3X2_HVT U884 ( .A1(n258), .A2(n1059), .A3(n337), .Y(n191) );
  INVX1_HVT U885 ( .A(n971), .Y(n560) );
  NAND2X0_HVT U886 ( .A1(n918), .A2(n919), .Y(n563) );
  NAND2X0_HVT U887 ( .A1(n562), .A2(n561), .Y(n564) );
  NAND2X0_HVT U888 ( .A1(n564), .A2(n563), .Y(out[92]) );
  INVX1_HVT U889 ( .A(n918), .Y(n561) );
  XOR3X2_HVT U890 ( .A1(n146), .A2(n952), .A3(n566), .Y(out[23]) );
  NAND2X0_HVT U891 ( .A1(n506), .A2(n854), .Y(n569) );
  NAND2X0_HVT U892 ( .A1(n567), .A2(n498), .Y(n570) );
  OR2X1_HVT U893 ( .A1(n881), .A2(n714), .Y(n761) );
  NAND2X0_HVT U894 ( .A1(in[61]), .A2(n170), .Y(n572) );
  NAND2X0_HVT U895 ( .A1(n571), .A2(n605), .Y(n573) );
  INVX0_HVT U896 ( .A(n170), .Y(n605) );
  NAND2X0_HVT U897 ( .A1(n216), .A2(n39), .Y(n576) );
  NAND2X0_HVT U898 ( .A1(n574), .A2(n575), .Y(n577) );
  NAND2X0_HVT U899 ( .A1(n577), .A2(n576), .Y(out[90]) );
  INVX1_HVT U900 ( .A(n732), .Y(n726) );
  NAND2X0_HVT U901 ( .A1(n778), .A2(n11), .Y(n578) );
  NAND2X0_HVT U902 ( .A1(n588), .A2(n329), .Y(n579) );
  NAND2X0_HVT U903 ( .A1(n578), .A2(n579), .Y(n965) );
  INVX0_HVT U904 ( .A(n1039), .Y(n850) );
  INVX1_HVT U905 ( .A(n745), .Y(n1059) );
  INVX0_HVT U906 ( .A(n665), .Y(n582) );
  XOR3X2_HVT U907 ( .A1(n6), .A2(n928), .A3(n38), .Y(n1015) );
  INVX0_HVT U908 ( .A(in[84]), .Y(n586) );
  NAND2X0_HVT U909 ( .A1(n778), .A2(n268), .Y(n590) );
  NAND2X0_HVT U910 ( .A1(n588), .A2(n531), .Y(n591) );
  NAND2X0_HVT U911 ( .A1(n590), .A2(n591), .Y(n121) );
  INVX0_HVT U912 ( .A(n778), .Y(n588) );
  XOR3X2_HVT U913 ( .A1(n1042), .A2(n1064), .A3(n323), .Y(n171) );
  XOR3X2_HVT U914 ( .A1(n592), .A2(n284), .A3(n210), .Y(out[102]) );
  NAND2X0_HVT U915 ( .A1(n784), .A2(n783), .Y(n592) );
  NAND2X0_HVT U916 ( .A1(n511), .A2(n45), .Y(n596) );
  NAND2X0_HVT U917 ( .A1(n137), .A2(n65), .Y(n597) );
  NBUFFX2_HVT U918 ( .A(n1070), .Y(n1069) );
  NBUFFX2_HVT U919 ( .A(n119), .Y(n602) );
  NAND2X0_HVT U920 ( .A1(n620), .A2(n621), .Y(n603) );
  XOR3X2_HVT U921 ( .A1(n146), .A2(n707), .A3(n201), .Y(out[31]) );
  NAND2X0_HVT U922 ( .A1(n754), .A2(n200), .Y(n608) );
  NAND2X0_HVT U923 ( .A1(n606), .A2(n607), .Y(n609) );
  NAND2X0_HVT U924 ( .A1(n609), .A2(n608), .Y(out[116]) );
  INVX1_HVT U925 ( .A(n754), .Y(n606) );
  NAND2X0_HVT U926 ( .A1(n833), .A2(n344), .Y(n610) );
  NAND2X0_HVT U927 ( .A1(n45), .A2(n450), .Y(n611) );
  NAND2X0_HVT U928 ( .A1(n610), .A2(n611), .Y(n657) );
  NAND2X0_HVT U929 ( .A1(n152), .A2(n1037), .Y(n614) );
  NAND2X0_HVT U930 ( .A1(n613), .A2(n317), .Y(n615) );
  NAND2X0_HVT U931 ( .A1(n614), .A2(n615), .Y(out[28]) );
  NBUFFX2_HVT U932 ( .A(n102), .Y(n617) );
  NAND2X0_HVT U933 ( .A1(n464), .A2(n83), .Y(n620) );
  NAND2X0_HVT U934 ( .A1(n618), .A2(n358), .Y(n621) );
  NAND2X0_HVT U935 ( .A1(n512), .A2(n664), .Y(n625) );
  NAND2X0_HVT U936 ( .A1(n623), .A2(n117), .Y(n626) );
  INVX1_HVT U937 ( .A(n758), .Y(n955) );
  NAND2X0_HVT U938 ( .A1(in[8]), .A2(n629), .Y(n630) );
  NAND2X0_HVT U939 ( .A1(n628), .A2(n506), .Y(n631) );
  NAND2X0_HVT U940 ( .A1(n630), .A2(n631), .Y(n944) );
  INVX0_HVT U941 ( .A(in[8]), .Y(n628) );
  NAND2X0_HVT U942 ( .A1(n1018), .A2(n176), .Y(n634) );
  NAND2X0_HVT U943 ( .A1(n632), .A2(n633), .Y(n635) );
  NAND2X0_HVT U944 ( .A1(n635), .A2(n634), .Y(out[12]) );
  NBUFFX2_HVT U945 ( .A(n122), .Y(n636) );
  INVX0_HVT U946 ( .A(in[36]), .Y(n721) );
  XOR3X2_HVT U947 ( .A1(n104), .A2(n923), .A3(n105), .Y(out[56]) );
  NAND2X0_HVT U948 ( .A1(n638), .A2(n1015), .Y(n639) );
  NAND2X0_HVT U949 ( .A1(n637), .A2(n37), .Y(n640) );
  NAND2X0_HVT U950 ( .A1(n639), .A2(n640), .Y(out[91]) );
  XOR3X2_HVT U951 ( .A1(n75), .A2(n809), .A3(n297), .Y(out[71]) );
  INVX0_HVT U952 ( .A(in[113]), .Y(n695) );
  NAND2X0_HVT U953 ( .A1(n959), .A2(n1017), .Y(n646) );
  NAND2X0_HVT U954 ( .A1(n304), .A2(n645), .Y(n647) );
  NAND2X0_HVT U955 ( .A1(n647), .A2(n646), .Y(out[20]) );
  NAND2X0_HVT U956 ( .A1(n687), .A2(n727), .Y(n648) );
  NAND2X0_HVT U957 ( .A1(n172), .A2(n975), .Y(n651) );
  NAND2X0_HVT U958 ( .A1(n649), .A2(n650), .Y(n652) );
  NAND2X0_HVT U959 ( .A1(n652), .A2(n651), .Y(out[123]) );
  AND2X1_HVT U960 ( .A1(n794), .A2(n793), .Y(n655) );
  XOR3X2_HVT U961 ( .A1(n657), .A2(n785), .A3(n677), .Y(out[120]) );
  NAND2X0_HVT U962 ( .A1(n228), .A2(n91), .Y(n661) );
  NAND2X0_HVT U963 ( .A1(n492), .A2(n660), .Y(n662) );
  NAND2X0_HVT U964 ( .A1(n661), .A2(n662), .Y(n218) );
  INVX1_HVT U965 ( .A(n954), .Y(n667) );
  NAND2X0_HVT U966 ( .A1(n787), .A2(n307), .Y(n673) );
  NAND2X0_HVT U967 ( .A1(n672), .A2(n91), .Y(n674) );
  NAND2X0_HVT U968 ( .A1(n674), .A2(n673), .Y(n689) );
  XOR3X2_HVT U969 ( .A1(n150), .A2(n204), .A3(n118), .Y(out[21]) );
  NAND2X0_HVT U970 ( .A1(n942), .A2(n80), .Y(n679) );
  NAND2X0_HVT U971 ( .A1(n243), .A2(n678), .Y(n680) );
  NAND2X0_HVT U972 ( .A1(n680), .A2(n679), .Y(out[68]) );
  XOR3X2_HVT U973 ( .A1(n839), .A2(n208), .A3(n189), .Y(out[105]) );
  INVX1_HVT U974 ( .A(n766), .Y(n681) );
  NAND2X0_HVT U975 ( .A1(n628), .A2(n1065), .Y(n683) );
  NAND2X0_HVT U976 ( .A1(n682), .A2(in[8]), .Y(n684) );
  NAND2X0_HVT U977 ( .A1(n683), .A2(n684), .Y(n162) );
  XOR3X2_HVT U978 ( .A1(n17), .A2(n686), .A3(n218), .Y(out[103]) );
  XOR3X2_HVT U979 ( .A1(n689), .A2(n285), .A3(n229), .Y(out[118]) );
  NAND2X0_HVT U980 ( .A1(n477), .A2(n212), .Y(n692) );
  NAND2X0_HVT U981 ( .A1(n9), .A2(n641), .Y(n693) );
  NAND2X0_HVT U982 ( .A1(n692), .A2(n693), .Y(n46) );
  INVX1_HVT U983 ( .A(n853), .Y(n727) );
  XOR3X2_HVT U984 ( .A1(n277), .A2(n1056), .A3(n114), .Y(n696) );
  XOR3X2_HVT U985 ( .A1(n824), .A2(n1068), .A3(n363), .Y(n200) );
  NAND2X0_HVT U986 ( .A1(n446), .A2(n153), .Y(n698) );
  NAND2X0_HVT U987 ( .A1(n751), .A2(n320), .Y(n699) );
  NAND2X0_HVT U988 ( .A1(n81), .A2(n723), .Y(n700) );
  NAND2X0_HVT U989 ( .A1(n699), .A2(n700), .Y(n863) );
  INVX0_HVT U990 ( .A(n81), .Y(n751) );
  XOR2X2_HVT U991 ( .A1(n666), .A2(n722), .Y(n111) );
  NAND2X0_HVT U992 ( .A1(n888), .A2(n66), .Y(n705) );
  NAND2X0_HVT U993 ( .A1(n704), .A2(n703), .Y(n706) );
  NAND2X0_HVT U994 ( .A1(n706), .A2(n705), .Y(out[76]) );
  NAND2X0_HVT U995 ( .A1(n1029), .A2(n183), .Y(n711) );
  NAND2X0_HVT U996 ( .A1(n709), .A2(n710), .Y(n712) );
  NAND2X0_HVT U997 ( .A1(n712), .A2(n711), .Y(out[124]) );
  XOR3X2_HVT U998 ( .A1(n715), .A2(n298), .A3(n177), .Y(out[119]) );
  NAND2X0_HVT U999 ( .A1(n810), .A2(n50), .Y(n717) );
  NAND2X0_HVT U1000 ( .A1(n716), .A2(n283), .Y(n718) );
  NAND2X0_HVT U1001 ( .A1(n221), .A2(n717), .Y(n80) );
  XOR3X2_HVT U1002 ( .A1(n228), .A2(n618), .A3(n785), .Y(n1023) );
  NAND2X0_HVT U1003 ( .A1(n681), .A2(n728), .Y(n729) );
  NAND2X0_HVT U1004 ( .A1(n766), .A2(n546), .Y(n730) );
  NAND2X0_HVT U1005 ( .A1(n1022), .A2(n82), .Y(n735) );
  NAND2X0_HVT U1006 ( .A1(n733), .A2(n734), .Y(n736) );
  NAND2X0_HVT U1007 ( .A1(n736), .A2(n735), .Y(out[67]) );
  NAND2X0_HVT U1008 ( .A1(n995), .A2(n495), .Y(n738) );
  NAND2X0_HVT U1009 ( .A1(n737), .A2(n738), .Y(n60) );
  NBUFFX2_HVT U1010 ( .A(in[61]), .Y(n739) );
  XOR3X2_HVT U1011 ( .A1(n603), .A2(n137), .A3(n22), .Y(out[106]) );
  XNOR2X2_HVT U1012 ( .A1(n825), .A2(n3), .Y(n193) );
  NAND2X0_HVT U1013 ( .A1(n222), .A2(n742), .Y(n743) );
  NAND2X0_HVT U1014 ( .A1(n741), .A2(n675), .Y(n744) );
  NAND2X0_HVT U1015 ( .A1(n743), .A2(n744), .Y(n77) );
  NAND2X0_HVT U1016 ( .A1(n749), .A2(n750), .Y(n747) );
  NAND2X0_HVT U1017 ( .A1(n81), .A2(n612), .Y(n749) );
  NAND2X0_HVT U1018 ( .A1(n748), .A2(in[6]), .Y(n750) );
  NAND2X0_HVT U1019 ( .A1(n749), .A2(n750), .Y(n147) );
  INVX1_HVT U1020 ( .A(n147), .Y(n897) );
  NAND2X0_HVT U1021 ( .A1(n998), .A2(n997), .Y(n753) );
  AND2X1_HVT U1022 ( .A1(n796), .A2(n797), .Y(n754) );
  INVX0_HVT U1023 ( .A(n889), .Y(n755) );
  INVX0_HVT U1024 ( .A(n757), .Y(n758) );
  NAND2X0_HVT U1025 ( .A1(n714), .A2(n169), .Y(n760) );
  NAND2X0_HVT U1026 ( .A1(n761), .A2(n760), .Y(n810) );
  XOR3X2_HVT U1027 ( .A1(n42), .A2(n219), .A3(n856), .Y(out[1]) );
  NAND2X0_HVT U1028 ( .A1(n922), .A2(n113), .Y(n764) );
  NAND2X0_HVT U1029 ( .A1(n762), .A2(n763), .Y(n765) );
  NAND2X0_HVT U1030 ( .A1(n764), .A2(n765), .Y(out[51]) );
  XOR3X2_HVT U1031 ( .A1(n775), .A2(n381), .A3(n14), .Y(n969) );
  NAND2X0_HVT U1032 ( .A1(n1010), .A2(n1049), .Y(n769) );
  NAND2X0_HVT U1033 ( .A1(n767), .A2(n768), .Y(n770) );
  NAND2X0_HVT U1034 ( .A1(n770), .A2(n769), .Y(out[108]) );
  NAND2X0_HVT U1035 ( .A1(n772), .A2(n96), .Y(n773) );
  NAND2X0_HVT U1036 ( .A1(n771), .A2(n800), .Y(n774) );
  NAND2X0_HVT U1037 ( .A1(n774), .A2(n773), .Y(out[59]) );
  XOR3X2_HVT U1038 ( .A1(n202), .A2(n285), .A3(n120), .Y(out[101]) );
  XOR3X2_HVT U1039 ( .A1(n747), .A2(n781), .A3(n94), .Y(out[30]) );
  XOR3X2_HVT U1040 ( .A1(n178), .A2(n223), .A3(n120), .Y(out[126]) );
  NAND2X0_HVT U1041 ( .A1(n782), .A2(in[125]), .Y(n783) );
  NAND2X0_HVT U1042 ( .A1(n261), .A2(n318), .Y(n784) );
  NAND2X0_HVT U1043 ( .A1(n891), .A2(n788), .Y(n789) );
  NAND2X0_HVT U1044 ( .A1(n1041), .A2(n780), .Y(n790) );
  NAND2X0_HVT U1045 ( .A1(n789), .A2(n790), .Y(n859) );
  NAND2X0_HVT U1046 ( .A1(n792), .A2(n853), .Y(n793) );
  NAND2X0_HVT U1047 ( .A1(n752), .A2(n727), .Y(n794) );
  NAND2X0_HVT U1048 ( .A1(n648), .A2(n793), .Y(n95) );
  NAND2X0_HVT U1049 ( .A1(n795), .A2(n799), .Y(n796) );
  NAND2X0_HVT U1050 ( .A1(n380), .A2(n202), .Y(n797) );
  XOR3X2_HVT U1051 ( .A1(n779), .A2(n961), .A3(n1060), .Y(n800) );
  XOR3X2_HVT U1052 ( .A1(n881), .A2(n343), .A3(n32), .Y(n888) );
  NAND2X0_HVT U1053 ( .A1(n549), .A2(n1055), .Y(n804) );
  NAND2X0_HVT U1054 ( .A1(n803), .A2(n538), .Y(n805) );
  NAND2X0_HVT U1055 ( .A1(n804), .A2(n805), .Y(out[115]) );
  XOR3X2_HVT U1056 ( .A1(n624), .A2(n701), .A3(n807), .Y(n806) );
  XOR3X2_HVT U1057 ( .A1(n520), .A2(n241), .A3(n663), .Y(n856) );
  NBUFFX2_HVT U1058 ( .A(in[5]), .Y(n808) );
  XOR3X2_HVT U1059 ( .A1(n423), .A2(n809), .A3(n356), .Y(out[78]) );
  NAND2X0_HVT U1060 ( .A1(n127), .A2(n976), .Y(n814) );
  NAND2X0_HVT U1061 ( .A1(n812), .A2(n813), .Y(n815) );
  NAND2X0_HVT U1062 ( .A1(n815), .A2(n814), .Y(out[43]) );
  XOR3X2_HVT U1063 ( .A1(n714), .A2(n581), .A3(n957), .Y(n829) );
  OR2X1_HVT U1064 ( .A1(n126), .A2(n696), .Y(n826) );
  XOR3X2_HVT U1065 ( .A1(n35), .A2(n332), .A3(n161), .Y(out[77]) );
  XOR3X2_HVT U1066 ( .A1(n831), .A2(n656), .A3(n177), .Y(out[127]) );
  XOR3X2_HVT U1067 ( .A1(n857), .A2(n725), .A3(n874), .Y(n134) );
  XOR3X2_HVT U1068 ( .A1(n43), .A2(n44), .A3(n823), .Y(out[89]) );
  INVX1_HVT U1069 ( .A(n1014), .Y(n824) );
  XOR3X2_HVT U1070 ( .A1(n90), .A2(n546), .A3(n227), .Y(out[61]) );
  NAND2X0_HVT U1071 ( .A1(n696), .A2(n126), .Y(n827) );
  NAND2X0_HVT U1072 ( .A1(n826), .A2(n827), .Y(out[44]) );
  XOR3X2_HVT U1073 ( .A1(n217), .A2(n133), .A3(n274), .Y(out[104]) );
  XOR3X2_HVT U1074 ( .A1(n48), .A2(n430), .A3(n28), .Y(out[87]) );
  NAND2X0_HVT U1075 ( .A1(n1032), .A2(n52), .Y(n836) );
  NAND2X0_HVT U1076 ( .A1(n834), .A2(n835), .Y(n837) );
  NAND2X0_HVT U1077 ( .A1(n837), .A2(n836), .Y(out[84]) );
  XOR3X2_HVT U1078 ( .A1(n1052), .A2(n432), .A3(n53), .Y(n52) );
  XOR3X2_HVT U1079 ( .A1(n1068), .A2(n512), .A3(n294), .Y(n1010) );
  NAND2X0_HVT U1080 ( .A1(n54), .A2(n953), .Y(n843) );
  NAND2X0_HVT U1081 ( .A1(n842), .A2(n841), .Y(n844) );
  NAND2X0_HVT U1082 ( .A1(n844), .A2(n843), .Y(out[83]) );
  XOR3X2_HVT U1083 ( .A1(n85), .A2(n196), .A3(n753), .Y(out[64]) );
  XOR3X2_HVT U1084 ( .A1(n253), .A2(n565), .A3(n39), .Y(out[82]) );
  NAND2X0_HVT U1085 ( .A1(n846), .A2(n141), .Y(n847) );
  NAND2X0_HVT U1086 ( .A1(n845), .A2(n1030), .Y(n848) );
  NAND2X0_HVT U1087 ( .A1(n848), .A2(n847), .Y(out[35]) );
  NAND2X0_HVT U1088 ( .A1(n1039), .A2(n194), .Y(n851) );
  NAND2X0_HVT U1089 ( .A1(n850), .A2(n849), .Y(n852) );
  NAND2X0_HVT U1090 ( .A1(n852), .A2(n851), .Y(out[11]) );
  XOR3X2_HVT U1091 ( .A1(n198), .A2(n115), .A3(n144), .Y(out[33]) );
  XOR3X2_HVT U1092 ( .A1(n291), .A2(n642), .A3(n19), .Y(n976) );
  XOR3X2_HVT U1093 ( .A1(n160), .A2(n324), .A3(n149), .Y(out[10]) );
  XOR2X2_HVT U1094 ( .A1(n1065), .A2(n854), .Y(n994) );
  XOR3X2_HVT U1095 ( .A1(n944), .A2(n943), .A3(n2), .Y(out[0]) );
  XOR3X2_HVT U1096 ( .A1(n428), .A2(n583), .A3(n948), .Y(n1026) );
  NAND2X0_HVT U1097 ( .A1(n517), .A2(n521), .Y(n861) );
  NAND2X0_HVT U1098 ( .A1(n567), .A2(n1066), .Y(n862) );
  NAND2X0_HVT U1099 ( .A1(n861), .A2(n862), .Y(n874) );
  XOR3X2_HVT U1100 ( .A1(n897), .A2(n517), .A3(n63), .Y(out[15]) );
  XOR3X2_HVT U1101 ( .A1(n863), .A2(n1063), .A3(n63), .Y(out[7]) );
  XOR3X2_HVT U1102 ( .A1(n125), .A2(n306), .A3(n864), .Y(out[125]) );
  NAND2X0_HVT U1103 ( .A1(n1026), .A2(n134), .Y(n867) );
  NAND2X0_HVT U1104 ( .A1(n865), .A2(n866), .Y(n868) );
  NAND2X0_HVT U1105 ( .A1(n868), .A2(n867), .Y(out[3]) );
  XOR3X2_HVT U1106 ( .A1(n44), .A2(n869), .A3(n71), .Y(out[74]) );
  XOR3X2_HVT U1107 ( .A1(n882), .A2(n871), .A3(n872), .Y(n68) );
  XOR3X2_HVT U1108 ( .A1(n64), .A2(n873), .A3(n395), .Y(out[79]) );
  NBUFFX2_HVT U1109 ( .A(in[109]), .Y(n875) );
  XOR3X2_HVT U1110 ( .A1(n589), .A2(n456), .A3(n329), .Y(n958) );
  NAND2X0_HVT U1111 ( .A1(n926), .A2(n666), .Y(n879) );
  NAND2X0_HVT U1112 ( .A1(n878), .A2(n879), .Y(n90) );
  XOR3X2_HVT U1113 ( .A1(n495), .A2(n1035), .A3(n882), .Y(n1032) );
  XOR3X2_HVT U1114 ( .A1(n811), .A2(n237), .A3(n943), .Y(n963) );
  NAND2X0_HVT U1115 ( .A1(n249), .A2(n92), .Y(n886) );
  NAND2X0_HVT U1116 ( .A1(n616), .A2(n885), .Y(n887) );
  NAND2X0_HVT U1117 ( .A1(n887), .A2(n886), .Y(out[60]) );
  NAND2X0_HVT U1118 ( .A1(n755), .A2(n95), .Y(n890) );
  NAND2X0_HVT U1119 ( .A1(n192), .A2(n890), .Y(n1038) );
  XOR3X2_HVT U1120 ( .A1(n247), .A2(n892), .A3(n429), .Y(n66) );
  NAND2X0_HVT U1121 ( .A1(n1048), .A2(n412), .Y(n895) );
  NAND2X0_HVT U1122 ( .A1(n894), .A2(n1036), .Y(n896) );
  NAND2X0_HVT U1123 ( .A1(n896), .A2(n895), .Y(out[27]) );
  NAND2X0_HVT U1124 ( .A1(n899), .A2(n985), .Y(n900) );
  NAND2X0_HVT U1125 ( .A1(n898), .A2(n171), .Y(n901) );
  NAND2X0_HVT U1126 ( .A1(n901), .A2(n900), .Y(out[19]) );
  NAND2X0_HVT U1127 ( .A1(n788), .A2(n956), .Y(n903) );
  NAND2X0_HVT U1128 ( .A1(n589), .A2(n409), .Y(n904) );
  NAND2X0_HVT U1129 ( .A1(n904), .A2(n903), .Y(n123) );
  NAND2X0_HVT U1130 ( .A1(n1031), .A2(n940), .Y(n906) );
  NAND2X0_HVT U1131 ( .A1(n905), .A2(n806), .Y(n907) );
  NAND2X0_HVT U1132 ( .A1(n906), .A2(n907), .Y(out[107]) );
  NBUFFX2_HVT U1133 ( .A(n61), .Y(n911) );
  NAND2X0_HVT U1134 ( .A1(n913), .A2(n109), .Y(n914) );
  NAND2X0_HVT U1135 ( .A1(n912), .A2(n1027), .Y(n915) );
  NAND2X0_HVT U1136 ( .A1(n914), .A2(n915), .Y(out[52]) );
  XOR3X2_HVT U1137 ( .A1(n756), .A2(n1001), .A3(n970), .Y(n942) );
  XOR3X2_HVT U1138 ( .A1(n545), .A2(n1034), .A3(n230), .Y(n109) );
  XOR3X2_HVT U1139 ( .A1(n212), .A2(n756), .A3(n931), .Y(n918) );
  XOR3X2_HVT U1140 ( .A1(n121), .A2(n195), .A3(n636), .Y(out[48]) );
  XNOR2X1_HVT U1141 ( .A1(n732), .A2(n654), .Y(n22) );
  XOR3X2_HVT U1142 ( .A1(n668), .A2(n460), .A3(n925), .Y(n1039) );
  XOR3X2_HVT U1143 ( .A1(n100), .A2(n122), .A3(n929), .Y(out[41]) );
  XOR3X2_HVT U1144 ( .A1(n489), .A2(n354), .A3(n934), .Y(n940) );
  XOR3X2_HVT U1145 ( .A1(n659), .A2(n937), .A3(n1057), .Y(n1030) );
  NAND2X0_HVT U1146 ( .A1(n1038), .A2(n968), .Y(n949) );
  NAND2X0_HVT U1147 ( .A1(n950), .A2(n949), .Y(n959) );
  XOR3X2_HVT U1148 ( .A1(n232), .A2(n175), .A3(n1020), .Y(n141) );
  XOR3X2_HVT U1149 ( .A1(n130), .A2(n19), .A3(n617), .Y(out[42]) );
  XOR3X2_HVT U1150 ( .A1(n955), .A2(n778), .A3(n505), .Y(n144) );
  XOR3X2_HVT U1151 ( .A1(n46), .A2(n957), .A3(n350), .Y(out[88]) );
  XOR3X2_HVT U1152 ( .A1(n101), .A2(n102), .A3(n958), .Y(out[57]) );
  XOR3X2_HVT U1153 ( .A1(n1033), .A2(n1063), .A3(n960), .Y(out[8]) );
  XOR3X2_HVT U1154 ( .A1(n516), .A2(n961), .A3(n111), .Y(n1027) );
  XOR3X2_HVT U1155 ( .A1(n148), .A2(n925), .A3(n149), .Y(out[2]) );
  XOR3X2_HVT U1156 ( .A1(n198), .A2(n964), .A3(n965), .Y(out[40]) );
  XOR3X2_HVT U1157 ( .A1(n77), .A2(n952), .A3(n201), .Y(out[6]) );
  XOR3X2_HVT U1158 ( .A1(n21), .A2(n966), .A3(n22), .Y(out[98]) );
  XOR3X2_HVT U1159 ( .A1(n16), .A2(n293), .A3(n158), .Y(out[26]) );
  XOR2X2_HVT U1160 ( .A1(n535), .A2(n685), .Y(n93) );
  XOR3X2_HVT U1161 ( .A1(n74), .A2(n103), .A3(n84), .Y(out[65]) );
  XOR3X2_HVT U1162 ( .A1(n106), .A2(n973), .A3(n244), .Y(out[55]) );
  XOR3X2_HVT U1163 ( .A1(n162), .A2(n981), .A3(n947), .Y(out[24]) );
  XOR3X2_HVT U1164 ( .A1(n163), .A2(n148), .A3(n983), .Y(out[17]) );
  XOR3X2_HVT U1165 ( .A1(n339), .A2(in[8]), .A3(n1063), .Y(n983) );
  XOR3X2_HVT U1166 ( .A1(n644), .A2(n694), .A3(n641), .Y(n984) );
  XOR3X2_HVT U1167 ( .A1(n58), .A2(n740), .A3(n71), .Y(out[66]) );
  NAND2X0_HVT U1168 ( .A1(n140), .A2(n1024), .Y(n988) );
  NAND2X0_HVT U1169 ( .A1(n986), .A2(n987), .Y(n989) );
  NAND2X0_HVT U1170 ( .A1(n989), .A2(n988), .Y(out[36]) );
  XOR3X2_HVT U1171 ( .A1(n909), .A2(n880), .A3(n780), .Y(n1024) );
  NAND2X0_HVT U1172 ( .A1(n187), .A2(n212), .Y(n992) );
  NAND2X0_HVT U1173 ( .A1(n996), .A2(n434), .Y(n993) );
  NAND2X0_HVT U1174 ( .A1(n993), .A2(n992), .Y(n48) );
  NAND2X0_HVT U1175 ( .A1(in[88]), .A2(n212), .Y(n997) );
  NAND2X0_HVT U1176 ( .A1(n995), .A2(n996), .Y(n998) );
  NAND2X0_HVT U1177 ( .A1(n997), .A2(n998), .Y(n43) );
  XOR3X2_HVT U1178 ( .A1(in[88]), .A2(n466), .A3(n970), .Y(n84) );
  NAND2X0_HVT U1179 ( .A1(n1006), .A2(n220), .Y(n1007) );
  NAND2X0_HVT U1180 ( .A1(n1019), .A2(n1005), .Y(n1008) );
  NAND2X0_HVT U1181 ( .A1(n1008), .A2(n1007), .Y(out[100]) );
  INVX0_HVT U1182 ( .A(n220), .Y(n1005) );
  XOR3X2_HVT U1183 ( .A1(n1009), .A2(n119), .A3(n105), .Y(out[49]) );
  XOR3X2_HVT U1184 ( .A1(n157), .A2(n193), .A3(n1023), .Y(out[113]) );
  XOR3X2_HVT U1185 ( .A1(n668), .A2(n1047), .A3(n707), .Y(n1017) );
  XOR3X2_HVT U1186 ( .A1(n506), .A2(n1011), .A3(n916), .Y(n1018) );
  XOR3X2_HVT U1187 ( .A1(n1069), .A2(n1021), .A3(n167), .Y(n220) );
  NBUFFX2_HVT U1188 ( .A(in[31]), .Y(n1066) );
  NBUFFX2_HVT U1189 ( .A(in[71]), .Y(n1067) );
  NAND2X0_HVT U1190 ( .A1(n1044), .A2(n68), .Y(n1045) );
  NAND2X0_HVT U1191 ( .A1(n1043), .A2(n69), .Y(n1046) );
  NAND2X0_HVT U1192 ( .A1(n1045), .A2(n1046), .Y(out[75]) );
  XNOR2X1_HVT U1193 ( .A1(n76), .A2(n228), .Y(n177) );
endmodule

