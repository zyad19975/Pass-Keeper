
module inv_sbox_11 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n18, n196, n197, n198, n199, n200, n201, n202, n205, n206, n208, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605;

  NAND2X0_HVT U1 ( .A1(n270), .A2(n318), .Y(n605) );
  NAND2X0_HVT U4 ( .A1(n339), .A2(n330), .Y(n602) );
  NAND2X0_HVT U5 ( .A1(n602), .A2(n277), .Y(n601) );
  NAND2X0_HVT U6 ( .A1(n339), .A2(n281), .Y(n599) );
  NAND2X0_HVT U8 ( .A1(n335), .A2(n277), .Y(n597) );
  NAND2X0_HVT U9 ( .A1(n334), .A2(n597), .Y(n596) );
  NAND2X0_HVT U10 ( .A1(n333), .A2(n594), .Y(n595) );
  NAND2X0_HVT U11 ( .A1(n288), .A2(n331), .Y(n593) );
  NAND2X0_HVT U12 ( .A1(n335), .A2(n317), .Y(n592) );
  NAND2X0_HVT U13 ( .A1(n328), .A2(n597), .Y(n591) );
  NAND2X0_HVT U15 ( .A1(n324), .A2(n250), .Y(n589) );
  NAND2X0_HVT U19 ( .A1(n250), .A2(n399), .Y(n585) );
  NAND2X0_HVT U25 ( .A1(in[6]), .A2(n317), .Y(n600) );
  NAND2X0_HVT U32 ( .A1(n319), .A2(n288), .Y(n573) );
  NAND2X0_HVT U35 ( .A1(n597), .A2(n295), .Y(n570) );
  NAND2X0_HVT U38 ( .A1(n316), .A2(n288), .Y(n567) );
  NAND2X0_HVT U42 ( .A1(n599), .A2(n295), .Y(n563) );
  OA21X1_HVT U53 ( .A1(n199), .A2(n555), .A3(n286), .Y(n553) );
  NAND2X0_HVT U55 ( .A1(n328), .A2(n602), .Y(n551) );
  MUX41X1_HVT U56 ( .A1(n384), .A3(n229), .A2(n371), .A4(n551), .S0(n310), 
        .S1(n243), .Y(n550) );
  AO21X1_HVT U60 ( .A1(n545), .A2(n314), .A3(n584), .Y(n546) );
  MUX41X1_HVT U62 ( .A1(n544), .A3(n550), .A2(n548), .A4(n552), .S0(n248), 
        .S1(n249), .Y(n543) );
  MUX41X1_HVT U65 ( .A1(n365), .A3(n367), .A2(n366), .A4(n567), .S0(n310), 
        .S1(n343), .Y(n540) );
  NAND2X0_HVT U66 ( .A1(n250), .A2(n208), .Y(n539) );
  MUX41X1_HVT U67 ( .A1(n362), .A3(n385), .A2(n364), .A4(n539), .S0(n315), 
        .S1(n307), .Y(n538) );
  MUX41X1_HVT U68 ( .A1(n362), .A3(n270), .A2(n363), .A4(n333), .S0(n309), 
        .S1(n243), .Y(n537) );
  MUX41X1_HVT U71 ( .A1(n599), .A3(n280), .A2(n593), .A4(n358), .S0(n309), 
        .S1(n244), .Y(n535) );
  NAND2X0_HVT U72 ( .A1(n325), .A2(n598), .Y(n534) );
  MUX41X1_HVT U73 ( .A1(n578), .A3(n534), .A2(n278), .A4(n316), .S0(n314), 
        .S1(n307), .Y(n533) );
  NAND2X0_HVT U81 ( .A1(n330), .A2(n598), .Y(n525) );
  AND2X1_HVT U82 ( .A1(n599), .A2(n328), .Y(n524) );
  MUX41X1_HVT U83 ( .A1(n524), .A3(n374), .A2(n283), .A4(n525), .S0(n309), 
        .S1(n243), .Y(n523) );
  MUX41X1_HVT U84 ( .A1(n304), .A3(n373), .A2(n387), .A4(n580), .S0(n310), 
        .S1(n244), .Y(n522) );
  MUX41X1_HVT U85 ( .A1(n522), .A3(n526), .A2(n523), .A4(n527), .S0(n248), 
        .S1(n322), .Y(n521) );
  NAND2X0_HVT U89 ( .A1(n285), .A2(n397), .Y(n518) );
  MUX41X1_HVT U90 ( .A1(n280), .A3(n598), .A2(n558), .A4(n518), .S0(n309), 
        .S1(n244), .Y(n517) );
  MUX41X1_HVT U96 ( .A1(n385), .A3(n591), .A2(n372), .A4(n389), .S0(n310), 
        .S1(n344), .Y(n511) );
  MUX41X1_HVT U98 ( .A1(n510), .A3(n390), .A2(n377), .A4(n577), .S0(n310), 
        .S1(n344), .Y(n509) );
  MUX41X1_HVT U99 ( .A1(n573), .A3(n366), .A2(n557), .A4(n229), .S0(n343), 
        .S1(n307), .Y(n508) );
  NAND2X0_HVT U100 ( .A1(n285), .A2(n396), .Y(n507) );
  MUX41X1_HVT U101 ( .A1(n391), .A3(n592), .A2(n206), .A4(n507), .S0(n243), 
        .S1(n306), .Y(n506) );
  AND2X1_HVT U104 ( .A1(n598), .A2(n326), .Y(n504) );
  MUX41X1_HVT U107 ( .A1(n391), .A3(n329), .A2(n502), .A4(n355), .S0(n309), 
        .S1(n244), .Y(n501) );
  MUX41X1_HVT U108 ( .A1(n368), .A3(n229), .A2(n371), .A4(n332), .S0(n310), 
        .S1(n243), .Y(n500) );
  MUX41X1_HVT U109 ( .A1(n390), .A3(n349), .A2(n387), .A4(n382), .S0(n309), 
        .S1(n343), .Y(n499) );
  MUX41X1_HVT U110 ( .A1(n499), .A3(n501), .A2(n500), .A4(n503), .S0(n248), 
        .S1(n322), .Y(n498) );
  AO21X1_HVT U112 ( .A1(n379), .A2(n314), .A3(n581), .Y(n496) );
  NAND2X0_HVT U114 ( .A1(n333), .A2(n598), .Y(n494) );
  MUX41X1_HVT U115 ( .A1(n494), .A3(n593), .A2(n379), .A4(n328), .S0(n343), 
        .S1(n307), .Y(n493) );
  MUX41X1_HVT U116 ( .A1(n378), .A3(n373), .A2(n349), .A4(n589), .S0(n308), 
        .S1(n244), .Y(n492) );
  NAND2X0_HVT U118 ( .A1(n284), .A2(n270), .Y(n490) );
  MUX41X1_HVT U122 ( .A1(n383), .A3(n299), .A2(n559), .A4(n242), .S0(n308), 
        .S1(n344), .Y(n487) );
  MUX41X1_HVT U124 ( .A1(n302), .A3(n486), .A2(n582), .A4(n227), .S0(n343), 
        .S1(n308), .Y(n485) );
  AOI21X1_HVT U127 ( .A1(n313), .A2(n481), .A3(n356), .Y(n482) );
  NAND2X0_HVT U129 ( .A1(n312), .A2(n333), .Y(n479) );
  MUX41X1_HVT U130 ( .A1(n479), .A3(n480), .A2(n483), .A4(n482), .S0(n315), 
        .S1(n249), .Y(n478) );
  AND2X1_HVT U131 ( .A1(n279), .A2(n239), .Y(n477) );
  MUX41X1_HVT U132 ( .A1(n353), .A3(n477), .A2(n395), .A4(n362), .S0(n314), 
        .S1(n306), .Y(n476) );
  MUX41X1_HVT U133 ( .A1(n282), .A3(n355), .A2(n551), .A4(n354), .S0(n343), 
        .S1(n306), .Y(n475) );
  MUX41X1_HVT U136 ( .A1(n556), .A3(n507), .A2(n473), .A4(n360), .S0(n312), 
        .S1(n344), .Y(n472) );
  MUX41X1_HVT U137 ( .A1(n597), .A3(n576), .A2(n233), .A4(n389), .S0(n315), 
        .S1(n306), .Y(n471) );
  MUX41X1_HVT U140 ( .A1(n375), .A3(n301), .A2(n370), .A4(n593), .S0(n314), 
        .S1(n307), .Y(n469) );
  NAND2X0_HVT U141 ( .A1(n324), .A2(n284), .Y(n468) );
  MUX41X1_HVT U142 ( .A1(n468), .A3(n566), .A2(n394), .A4(n370), .S0(n313), 
        .S1(n344), .Y(n467) );
  MUX41X1_HVT U143 ( .A1(n397), .A3(n380), .A2(n585), .A4(n582), .S0(n311), 
        .S1(n237), .Y(n466) );
  MUX41X1_HVT U145 ( .A1(n574), .A3(n392), .A2(n465), .A4(n525), .S0(n313), 
        .S1(n237), .Y(n464) );
  MUX41X1_HVT U146 ( .A1(n464), .A3(n466), .A2(n467), .A4(n469), .S0(n322), 
        .S1(n248), .Y(n463) );
  AO21X1_HVT U148 ( .A1(n315), .A2(n357), .A3(n396), .Y(n461) );
  MUX41X1_HVT U151 ( .A1(n283), .A3(n377), .A2(n293), .A4(n459), .S0(n344), 
        .S1(n306), .Y(n458) );
  MUX41X1_HVT U155 ( .A1(n370), .A3(n593), .A2(n586), .A4(n372), .S0(n311), 
        .S1(n238), .Y(n454) );
  MUX41X1_HVT U156 ( .A1(n454), .A3(n458), .A2(n455), .A4(n460), .S0(in[5]), 
        .S1(n249), .Y(n453) );
  NAND2X0_HVT U159 ( .A1(n450), .A2(n449), .Y(n451) );
  MUX41X1_HVT U162 ( .A1(n291), .A3(n367), .A2(n570), .A4(n447), .S0(n311), 
        .S1(n237), .Y(n446) );
  NAND2X0_HVT U163 ( .A1(n335), .A2(n397), .Y(n445) );
  MUX41X1_HVT U164 ( .A1(n596), .A3(n445), .A2(n568), .A4(n368), .S0(n308), 
        .S1(n238), .Y(n444) );
  NAND2X0_HVT U166 ( .A1(n594), .A2(n441), .Y(n442) );
  MUX41X1_HVT U172 ( .A1(n518), .A3(n436), .A2(n300), .A4(n583), .S0(n311), 
        .S1(n237), .Y(n435) );
  NAND2X0_HVT U177 ( .A1(n337), .A2(n270), .Y(n431) );
  AND2X1_HVT U179 ( .A1(n599), .A2(n326), .Y(n429) );
  AND2X1_HVT U185 ( .A1(n295), .A2(n239), .Y(n423) );
  NAND2X0_HVT U191 ( .A1(n199), .A2(n361), .Y(n417) );
  AND2X1_HVT U192 ( .A1(n376), .A2(n415), .Y(n416) );
  NAND2X0_HVT U194 ( .A1(n415), .A2(n563), .Y(n413) );
  MUX41X1_HVT U195 ( .A1(n414), .A3(n413), .A2(n416), .A4(n417), .S0(n309), 
        .S1(n322), .Y(n412) );
  NAND2X0_HVT U198 ( .A1(n335), .A2(n230), .Y(n594) );
  NAND2X0_HVT U200 ( .A1(n277), .A2(n285), .Y(n481) );
  NAND2X0_HVT U207 ( .A1(n284), .A2(n280), .Y(n545) );
  MUX41X1_HVT U2 ( .A1(n435), .A3(n433), .A2(n437), .A4(n434), .S0(n202), .S1(
        n18), .Y(n432) );
  IBUFFX16_HVT U3 ( .A(n205), .Y(n18) );
  MUX21X1_HVT U7 ( .A1(n197), .A2(n198), .S0(n251), .Y(n196) );
  IBUFFX16_HVT U14 ( .A(n196), .Y(n242) );
  IBUFFX16_HVT U16 ( .A(n327), .Y(n197) );
  IBUFFX16_HVT U17 ( .A(n290), .Y(n198) );
  INVX0_HVT U18 ( .A(n337), .Y(n231) );
  INVX1_HVT U20 ( .A(n239), .Y(n337) );
  INVX1_HVT U21 ( .A(n342), .Y(n199) );
  INVX0_HVT U22 ( .A(n346), .Y(n342) );
  INVX1_HVT U23 ( .A(in[0]), .Y(n340) );
  INVX0_HVT U24 ( .A(n318), .Y(n200) );
  INVX1_HVT U26 ( .A(n319), .Y(n208) );
  MUX21X2_HVT U27 ( .A1(n304), .A2(n580), .S0(n218), .Y(n457) );
  MUX21X2_HVT U28 ( .A1(n601), .A2(n370), .S0(n201), .Y(n549) );
  IBUFFX16_HVT U29 ( .A(n313), .Y(n201) );
  MUX21X1_HVT U30 ( .A1(n329), .A2(n516), .S0(n219), .Y(n515) );
  IBUFFX16_HVT U31 ( .A(n248), .Y(n202) );
  IBUFFX16_HVT U33 ( .A(n322), .Y(n205) );
  MUX21X1_HVT U34 ( .A1(n324), .A2(n208), .S0(n340), .Y(n206) );
  IBUFFX16_HVT U36 ( .A(n206), .Y(n569) );
  MUX21X2_HVT U37 ( .A1(n472), .A2(n471), .S0(n217), .Y(n470) );
  IBUFFX16_HVT U39 ( .A(n322), .Y(n217) );
  INVX1_HVT U40 ( .A(n346), .Y(n345) );
  IBUFFX16_HVT U41 ( .A(n314), .Y(n218) );
  MUX21X2_HVT U43 ( .A1(n451), .A2(n452), .S0(n313), .Y(n448) );
  IBUFFX16_HVT U44 ( .A(n336), .Y(n219) );
  NAND2X0_HVT U45 ( .A1(n330), .A2(n220), .Y(n221) );
  NAND2X0_HVT U46 ( .A1(n325), .A2(n239), .Y(n222) );
  NAND2X0_HVT U47 ( .A1(n221), .A2(n222), .Y(n293) );
  IBUFFX2_HVT U48 ( .A(n239), .Y(n220) );
  INVX1_HVT U49 ( .A(in[0]), .Y(n239) );
  INVX0_HVT U50 ( .A(n293), .Y(n583) );
  MUX21X1_HVT U51 ( .A1(n602), .A2(n293), .S0(n276), .Y(n542) );
  INVX1_HVT U52 ( .A(in[3]), .Y(n292) );
  MUX21X1_HVT U54 ( .A1(n333), .A2(n295), .S0(n239), .Y(n294) );
  NAND2X0_HVT U57 ( .A1(n353), .A2(n223), .Y(n224) );
  NAND2X0_HVT U58 ( .A1(n395), .A2(n252), .Y(n225) );
  NAND2X0_HVT U59 ( .A1(n224), .A2(n225), .Y(n462) );
  IBUFFX2_HVT U61 ( .A(n252), .Y(n223) );
  INVX0_HVT U63 ( .A(n601), .Y(n353) );
  MUX21X1_HVT U64 ( .A1(n462), .A2(n461), .S0(n312), .Y(n460) );
  MUX21X2_HVT U69 ( .A1(n453), .A2(n463), .S0(n269), .Y(out[5]) );
  INVX2_HVT U70 ( .A(in[4]), .Y(n346) );
  INVX2_HVT U74 ( .A(n236), .Y(n266) );
  INVX2_HVT U75 ( .A(n236), .Y(n262) );
  INVX1_HVT U76 ( .A(n266), .Y(n343) );
  IBUFFX2_HVT U77 ( .A(n290), .Y(n226) );
  NBUFFX2_HVT U78 ( .A(n400), .Y(n318) );
  NBUFFX2_HVT U79 ( .A(n400), .Y(n320) );
  NBUFFX2_HVT U80 ( .A(n400), .Y(n319) );
  XNOR2X2_HVT U86 ( .A1(n318), .A2(n226), .Y(n228) );
  INVX0_HVT U87 ( .A(n228), .Y(n289) );
  INVX1_HVT U88 ( .A(n315), .Y(n252) );
  MUX21X1_HVT U91 ( .A1(n332), .A2(n292), .S0(n336), .Y(n227) );
  IBUFFX16_HVT U92 ( .A(n227), .Y(n582) );
  INVX0_HVT U93 ( .A(n289), .Y(n229) );
  INVX1_HVT U94 ( .A(n229), .Y(n230) );
  MUX21X2_HVT U95 ( .A1(n320), .A2(n325), .S0(n231), .Y(n580) );
  MUX21X2_HVT U97 ( .A1(n543), .A2(n536), .S0(n232), .Y(out[0]) );
  IBUFFX16_HVT U102 ( .A(n269), .Y(n232) );
  INVX0_HVT U103 ( .A(n370), .Y(n233) );
  INVX1_HVT U105 ( .A(n580), .Y(n370) );
  MUX41X1_HVT U106 ( .A1(n519), .A3(n520), .A2(n513), .A4(n517), .S0(n234), 
        .S1(n235), .Y(n512) );
  IBUFFX16_HVT U111 ( .A(n245), .Y(n234) );
  IBUFFX16_HVT U113 ( .A(n248), .Y(n235) );
  MUX21X2_HVT U117 ( .A1(n514), .A2(n515), .S0(n312), .Y(n513) );
  MUX21X2_HVT U119 ( .A1(n456), .A2(n457), .S0(n313), .Y(n455) );
  AO21X2_HVT U120 ( .A1(n325), .A2(n602), .A3(n199), .Y(n441) );
  NBUFFX2_HVT U121 ( .A(n342), .Y(n236) );
  NBUFFX2_HVT U123 ( .A(n342), .Y(n237) );
  NBUFFX2_HVT U125 ( .A(n342), .Y(n238) );
  INVX1_HVT U126 ( .A(n262), .Y(n344) );
  INVX1_HVT U128 ( .A(n266), .Y(n244) );
  INVX0_HVT U134 ( .A(n292), .Y(n290) );
  INVX0_HVT U135 ( .A(n239), .Y(n336) );
  MUX21X1_HVT U138 ( .A1(n443), .A2(n442), .S0(n276), .Y(n440) );
  MUX21X1_HVT U139 ( .A1(n242), .A2(n562), .S0(n252), .Y(n452) );
  AO21X1_HVT U144 ( .A1(n250), .A2(n396), .A3(n273), .Y(n415) );
  OA21X1_HVT U147 ( .A1(n373), .A2(n266), .A3(n545), .Y(n419) );
  NBUFFX2_HVT U149 ( .A(n228), .Y(n325) );
  MUX21X1_HVT U150 ( .A1(n317), .A2(n399), .S0(n339), .Y(n562) );
  INVX1_HVT U152 ( .A(n326), .Y(n263) );
  NAND2X0_HVT U153 ( .A1(n250), .A2(n329), .Y(n598) );
  OA21X1_HVT U154 ( .A1(n351), .A2(n262), .A3(n584), .Y(n530) );
  INVX1_HVT U157 ( .A(n327), .Y(n399) );
  INVX0_HVT U158 ( .A(n563), .Y(n355) );
  INVX1_HVT U160 ( .A(n323), .Y(n248) );
  INVX1_HVT U161 ( .A(n324), .Y(n295) );
  INVX1_HVT U165 ( .A(n310), .Y(n267) );
  INVX0_HVT U167 ( .A(n313), .Y(n257) );
  INVX1_HVT U168 ( .A(in[5]), .Y(n323) );
  INVX1_HVT U169 ( .A(n345), .Y(n273) );
  INVX1_HVT U170 ( .A(n262), .Y(n243) );
  INVX0_HVT U171 ( .A(n336), .Y(n284) );
  INVX1_HVT U173 ( .A(n340), .Y(n335) );
  INVX1_HVT U174 ( .A(n321), .Y(n249) );
  INVX1_HVT U175 ( .A(in[1]), .Y(n321) );
  MUX21X1_HVT U176 ( .A1(n348), .A2(n242), .S0(n252), .Y(n531) );
  IBUFFX2_HVT U178 ( .A(n340), .Y(n250) );
  INVX1_HVT U180 ( .A(n340), .Y(n251) );
  NAND2X0_HVT U181 ( .A1(n428), .A2(n245), .Y(n240) );
  NAND2X0_HVT U182 ( .A1(n430), .A2(n249), .Y(n241) );
  NAND2X0_HVT U183 ( .A1(n240), .A2(n241), .Y(n427) );
  OR2X1_HVT U184 ( .A1(n292), .A2(n320), .Y(n603) );
  INVX0_HVT U186 ( .A(n292), .Y(n270) );
  INVX1_HVT U187 ( .A(n562), .Y(n380) );
  INVX1_HVT U188 ( .A(n521), .Y(n297) );
  MUX21X2_HVT U189 ( .A1(n530), .A2(n531), .S0(n257), .Y(n529) );
  NBUFFX2_HVT U190 ( .A(n345), .Y(n315) );
  MUX21X1_HVT U193 ( .A1(n554), .A2(n553), .S0(n312), .Y(n552) );
  INVX1_HVT U196 ( .A(n249), .Y(n245) );
  MUX41X1_HVT U197 ( .A1(n537), .A3(n540), .A2(n538), .A4(n541), .S0(n248), 
        .S1(n249), .Y(n536) );
  MUX41X1_HVT U199 ( .A1(n590), .A3(n525), .A2(n392), .A4(n504), .S0(n343), 
        .S1(n310), .Y(n503) );
  NAND2X0_HVT U201 ( .A1(n488), .A2(n268), .Y(n246) );
  NAND2X0_HVT U202 ( .A1(n498), .A2(n269), .Y(n247) );
  NAND2X0_HVT U203 ( .A1(n246), .A2(n247), .Y(out[3]) );
  INVX1_HVT U204 ( .A(n268), .Y(n269) );
  MUX41X1_HVT U205 ( .A1(n478), .A3(n484), .A2(n470), .A4(n474), .S0(in[5]), 
        .S1(n268), .Y(out[4]) );
  MUX41X1_HVT U206 ( .A1(n511), .A3(n508), .A2(n509), .A4(n506), .S0(n323), 
        .S1(n245), .Y(n505) );
  NAND2X0_HVT U208 ( .A1(n304), .A2(n252), .Y(n253) );
  NAND2X0_HVT U209 ( .A1(n557), .A2(n315), .Y(n254) );
  NAND2X0_HVT U210 ( .A1(n253), .A2(n254), .Y(n421) );
  NAND2X0_HVT U211 ( .A1(n297), .A2(n268), .Y(n255) );
  NAND2X0_HVT U212 ( .A1(n298), .A2(n269), .Y(n256) );
  NAND2X0_HVT U213 ( .A1(n255), .A2(n256), .Y(n296) );
  INVX0_HVT U214 ( .A(n296), .Y(out[1]) );
  MUX41X1_HVT U215 ( .A1(n448), .A3(n446), .A2(n444), .A4(n440), .S0(n245), 
        .S1(n323), .Y(n439) );
  MUX41X1_HVT U216 ( .A1(n386), .A3(n596), .A2(n384), .A4(n601), .S0(n343), 
        .S1(n309), .Y(n526) );
  INVX1_HVT U217 ( .A(n411), .Y(n384) );
  MUX41X1_HVT U218 ( .A1(n421), .A3(n420), .A2(n422), .A4(n419), .S0(n321), 
        .S1(n306), .Y(n418) );
  NAND2X0_HVT U219 ( .A1(n229), .A2(n335), .Y(n258) );
  NAND2X0_HVT U220 ( .A1(n290), .A2(n284), .Y(n259) );
  NAND2X0_HVT U221 ( .A1(n258), .A2(n259), .Y(n283) );
  NAND2X0_HVT U222 ( .A1(n317), .A2(n339), .Y(n260) );
  NAND2X0_HVT U223 ( .A1(n333), .A2(n285), .Y(n261) );
  NAND2X0_HVT U224 ( .A1(n260), .A2(n261), .Y(n282) );
  INVX1_HVT U225 ( .A(n321), .Y(n322) );
  INVX0_HVT U226 ( .A(n251), .Y(n285) );
  MUX41X1_HVT U227 ( .A1(n282), .A3(n295), .A2(n388), .A4(n551), .S0(n311), 
        .S1(n262), .Y(n433) );
  MUX21X2_HVT U228 ( .A1(n475), .A2(n476), .S0(n322), .Y(n474) );
  XNOR2X1_HVT U229 ( .A1(n263), .A2(n336), .Y(n557) );
  NAND2X0_HVT U230 ( .A1(n278), .A2(n252), .Y(n264) );
  NAND2X0_HVT U231 ( .A1(n564), .A2(n243), .Y(n265) );
  NAND2X0_HVT U232 ( .A1(n264), .A2(n265), .Y(n420) );
  INVX1_HVT U233 ( .A(n401), .Y(n395) );
  INVX1_HVT U234 ( .A(n528), .Y(n298) );
  MUX41X1_HVT U235 ( .A1(n438), .A3(n302), .A2(n300), .A4(n303), .S0(n267), 
        .S1(n266), .Y(n437) );
  MUX41X1_HVT U236 ( .A1(n283), .A3(n602), .A2(n352), .A4(n355), .S0(n199), 
        .S1(n267), .Y(n426) );
  MUX41X1_HVT U237 ( .A1(n368), .A3(n375), .A2(n376), .A4(n595), .S0(n267), 
        .S1(n262), .Y(n532) );
  AO21X2_HVT U238 ( .A1(n239), .A2(n334), .A3(n273), .Y(n449) );
  OA21X2_HVT U239 ( .A1(n350), .A2(n273), .A3(n359), .Y(n456) );
  INVX0_HVT U240 ( .A(n338), .Y(n288) );
  INVX0_HVT U241 ( .A(n320), .Y(n279) );
  INVX0_HVT U242 ( .A(n579), .Y(n371) );
  INVX0_HVT U243 ( .A(n294), .Y(n574) );
  INVX0_HVT U244 ( .A(n286), .Y(n577) );
  INVX1_HVT U245 ( .A(n312), .Y(n276) );
  INVX1_HVT U246 ( .A(n340), .Y(n338) );
  INVX1_HVT U247 ( .A(n600), .Y(n397) );
  INVX1_HVT U248 ( .A(in[7]), .Y(n268) );
  MUX21X1_HVT U249 ( .A1(n423), .A2(n386), .S0(n345), .Y(n422) );
  MUX21X2_HVT U250 ( .A1(n487), .A2(n485), .S0(n321), .Y(n484) );
  MUX41X1_HVT U251 ( .A1(n427), .A3(n424), .A2(n418), .A4(n412), .S0(n323), 
        .S1(n268), .Y(out[7]) );
  MUX41X1_HVT U252 ( .A1(n347), .A3(n573), .A2(n560), .A4(n429), .S0(n257), 
        .S1(n238), .Y(n428) );
  MUX41X1_HVT U253 ( .A1(n588), .A3(n294), .A2(n587), .A4(n373), .S0(n276), 
        .S1(n273), .Y(n527) );
  MUX41X1_HVT U254 ( .A1(n535), .A3(n532), .A2(n533), .A4(n529), .S0(n323), 
        .S1(n321), .Y(n528) );
  MUX41X1_HVT U255 ( .A1(n490), .A3(n568), .A2(n491), .A4(n393), .S0(n276), 
        .S1(n199), .Y(n489) );
  MUX41X1_HVT U256 ( .A1(n561), .A3(n280), .A2(n431), .A4(n303), .S0(n276), 
        .S1(n273), .Y(n430) );
  NBUFFX2_HVT U257 ( .A(n292), .Y(n317) );
  NAND2X0_HVT U258 ( .A1(n426), .A2(n249), .Y(n271) );
  NAND2X0_HVT U259 ( .A1(n425), .A2(n321), .Y(n272) );
  NAND2X0_HVT U260 ( .A1(n271), .A2(n272), .Y(n424) );
  INVX1_HVT U261 ( .A(n565), .Y(n379) );
  MUX41X1_HVT U262 ( .A1(n368), .A3(n563), .A2(n380), .A4(n384), .S0(n244), 
        .S1(n267), .Y(n425) );
  MUX21X1_HVT U263 ( .A1(n368), .A2(n542), .S0(n305), .Y(n541) );
  MUX21X1_HVT U264 ( .A1(n317), .A2(n324), .S0(n288), .Y(n584) );
  MUX41X1_HVT U265 ( .A1(n569), .A3(n331), .A2(n280), .A4(n281), .S0(n276), 
        .S1(n273), .Y(n434) );
  INVX1_HVT U266 ( .A(n409), .Y(n386) );
  NAND2X0_HVT U267 ( .A1(n579), .A2(n273), .Y(n274) );
  NAND2X0_HVT U268 ( .A1(n582), .A2(n345), .Y(n275) );
  NAND2X0_HVT U269 ( .A1(n274), .A2(n275), .Y(n443) );
  MUX41X1_HVT U270 ( .A1(n559), .A3(n575), .A2(n349), .A4(n364), .S0(n276), 
        .S1(n273), .Y(n519) );
  NBUFFX2_HVT U271 ( .A(n292), .Y(n316) );
  MUX41X1_HVT U272 ( .A1(n495), .A3(n492), .A2(n493), .A4(n489), .S0(n323), 
        .S1(n245), .Y(n488) );
  NAND2X0_HVT U273 ( .A1(n200), .A2(n317), .Y(n277) );
  INVX0_HVT U274 ( .A(n291), .Y(n561) );
  MUX21X1_HVT U275 ( .A1(n279), .A2(n330), .S0(n288), .Y(n278) );
  INVX0_HVT U276 ( .A(n397), .Y(n287) );
  MUX21X2_HVT U277 ( .A1(n496), .A2(n497), .S0(n313), .Y(n495) );
  MUX21X2_HVT U278 ( .A1(n369), .A2(n549), .S0(n305), .Y(n548) );
  INVX1_HVT U279 ( .A(n584), .Y(n368) );
  INVX0_HVT U280 ( .A(n605), .Y(n280) );
  INVX1_HVT U281 ( .A(n280), .Y(n281) );
  INVX0_HVT U282 ( .A(n333), .Y(n398) );
  NBUFFX2_HVT U283 ( .A(n605), .Y(n333) );
  MUX41X1_HVT U284 ( .A1(n388), .A3(n371), .A2(n352), .A4(n304), .S0(n308), 
        .S1(n266), .Y(n520) );
  MUX21X1_HVT U285 ( .A1(n287), .A2(n333), .S0(n288), .Y(n286) );
  INVX1_HVT U286 ( .A(n407), .Y(n388) );
  MUX21X2_HVT U287 ( .A1(n505), .A2(n512), .S0(n269), .Y(out[2]) );
  MUX21X2_HVT U288 ( .A1(n432), .A2(n439), .S0(n269), .Y(out[6]) );
  INVX1_HVT U289 ( .A(n572), .Y(n375) );
  MUX21X1_HVT U290 ( .A1(n334), .A2(n287), .S0(n288), .Y(n291) );
  INVX1_HVT U291 ( .A(n331), .Y(n396) );
  NBUFFX2_HVT U292 ( .A(n604), .Y(n330) );
  NBUFFX2_HVT U293 ( .A(n604), .Y(n332) );
  NBUFFX2_HVT U294 ( .A(n604), .Y(n331) );
  AND2X1_HVT U295 ( .A1(n332), .A2(n589), .Y(n299) );
  MUX21X1_HVT U296 ( .A1(n381), .A2(n302), .S0(n345), .Y(n414) );
  MUX21X1_HVT U297 ( .A1(n326), .A2(n328), .S0(n251), .Y(n447) );
  MUX21X1_HVT U298 ( .A1(n319), .A2(n397), .S0(n338), .Y(n459) );
  XOR2X1_HVT U299 ( .A1(n334), .A2(n339), .Y(n568) );
  MUX21X1_HVT U300 ( .A1(n398), .A2(n325), .S0(n339), .Y(n407) );
  MUX21X1_HVT U301 ( .A1(n396), .A2(n295), .S0(n250), .Y(n572) );
  MUX21X1_HVT U302 ( .A1(n319), .A2(n396), .S0(n250), .Y(n579) );
  MUX21X1_HVT U303 ( .A1(n547), .A2(n546), .S0(n312), .Y(n544) );
  MUX21X1_HVT U304 ( .A1(n227), .A2(n551), .S0(n314), .Y(n547) );
  MUX21X1_HVT U305 ( .A1(n398), .A2(n399), .S0(n336), .Y(n438) );
  MUX21X1_HVT U306 ( .A1(n398), .A2(n320), .S0(n251), .Y(n436) );
  NAND2X0_HVT U307 ( .A1(n316), .A2(n318), .Y(n604) );
  MUX21X1_HVT U308 ( .A1(n230), .A2(n319), .S0(n338), .Y(n402) );
  MUX21X1_HVT U309 ( .A1(n295), .A2(n317), .S0(n336), .Y(n566) );
  MUX21X1_HVT U310 ( .A1(n317), .A2(n396), .S0(n339), .Y(n575) );
  MUX21X1_HVT U311 ( .A1(n358), .A2(n324), .S0(n315), .Y(n514) );
  MUX21X1_HVT U312 ( .A1(n324), .A2(n319), .S0(n314), .Y(n516) );
  MUX21X1_HVT U313 ( .A1(n320), .A2(n331), .S0(n337), .Y(n502) );
  MUX21X1_HVT U314 ( .A1(n320), .A2(n325), .S0(n335), .Y(n565) );
  MUX21X1_HVT U315 ( .A1(n333), .A2(n331), .S0(n337), .Y(n590) );
  MUX21X1_HVT U316 ( .A1(n394), .A2(n301), .S0(n312), .Y(n483) );
  XOR2X1_HVT U317 ( .A1(n329), .A2(n336), .Y(n558) );
  XOR2X1_HVT U318 ( .A1(n325), .A2(n251), .Y(n559) );
  MUX21X1_HVT U319 ( .A1(n325), .A2(n397), .S0(n335), .Y(n571) );
  MUX21X1_HVT U320 ( .A1(n326), .A2(n331), .S0(n339), .Y(n401) );
  MUX21X1_HVT U321 ( .A1(n316), .A2(n332), .S0(n339), .Y(n409) );
  AND2X1_HVT U322 ( .A1(n599), .A2(n330), .Y(n300) );
  XNOR2X1_HVT U323 ( .A1(n332), .A2(n250), .Y(n301) );
  MUX21X1_HVT U324 ( .A1(n329), .A2(n330), .S0(n338), .Y(n587) );
  MUX21X1_HVT U325 ( .A1(n572), .A2(n299), .S0(n313), .Y(n480) );
  MUX21X1_HVT U326 ( .A1(n317), .A2(n320), .S0(n335), .Y(n560) );
  MUX21X1_HVT U327 ( .A1(n329), .A2(n317), .S0(n251), .Y(n586) );
  MUX21X1_HVT U328 ( .A1(n316), .A2(n329), .S0(n337), .Y(n404) );
  AND2X1_HVT U329 ( .A1(n335), .A2(n320), .Y(n302) );
  MUX21X1_HVT U330 ( .A1(n328), .A2(n319), .S0(n250), .Y(n486) );
  NBUFFX2_HVT U331 ( .A(n345), .Y(n314) );
  NBUFFX2_HVT U332 ( .A(n281), .Y(n334) );
  MUX21X1_HVT U333 ( .A1(n372), .A2(n363), .S0(n315), .Y(n554) );
  MUX21X1_HVT U334 ( .A1(n396), .A2(n399), .S0(n251), .Y(n555) );
  MUX21X1_HVT U335 ( .A1(n356), .A2(n564), .S0(n315), .Y(n497) );
  MUX21X1_HVT U336 ( .A1(n332), .A2(n277), .S0(n335), .Y(n465) );
  NBUFFX2_HVT U337 ( .A(n228), .Y(n324) );
  AND2X1_HVT U338 ( .A1(n399), .A2(n285), .Y(n303) );
  NBUFFX2_HVT U339 ( .A(n600), .Y(n326) );
  NBUFFX2_HVT U340 ( .A(n603), .Y(n327) );
  AND2X1_HVT U341 ( .A1(n328), .A2(n285), .Y(n304) );
  NBUFFX2_HVT U342 ( .A(n603), .Y(n329) );
  NBUFFX2_HVT U343 ( .A(n603), .Y(n328) );
  NBUFFX2_HVT U344 ( .A(n307), .Y(n311) );
  NBUFFX2_HVT U345 ( .A(n341), .Y(n313) );
  NBUFFX2_HVT U346 ( .A(in[2]), .Y(n312) );
  INVX1_HVT U347 ( .A(n340), .Y(n339) );
  XNOR2X1_HVT U348 ( .A1(n199), .A2(n308), .Y(n305) );
  NBUFFX2_HVT U349 ( .A(n341), .Y(n308) );
  NBUFFX2_HVT U350 ( .A(n341), .Y(n310) );
  NBUFFX2_HVT U351 ( .A(n341), .Y(n309) );
  NBUFFX2_HVT U352 ( .A(n341), .Y(n307) );
  NBUFFX2_HVT U353 ( .A(n341), .Y(n306) );
  INVX0_HVT U354 ( .A(in[6]), .Y(n400) );
  MUX21X1_HVT U355 ( .A1(n334), .A2(n270), .S0(n338), .Y(n450) );
  MUX21X1_HVT U356 ( .A1(n277), .A2(n270), .S0(n336), .Y(n510) );
  MUX21X1_HVT U357 ( .A1(n399), .A2(n397), .S0(n336), .Y(n491) );
  MUX21X1_HVT U358 ( .A1(n208), .A2(n398), .S0(n251), .Y(n581) );
  XOR2X1_HVT U359 ( .A1(n337), .A2(n279), .Y(n556) );
  MUX21X1_HVT U360 ( .A1(n396), .A2(n208), .S0(n337), .Y(n473) );
  MUX21X1_HVT U361 ( .A1(n279), .A2(n399), .S0(n338), .Y(n564) );
  MUX21X1_HVT U362 ( .A1(n279), .A2(n397), .S0(n250), .Y(n411) );
  MUX21X1_HVT U363 ( .A1(n270), .A2(n333), .S0(n339), .Y(n406) );
  MUX21X1_HVT U364 ( .A1(n277), .A2(n279), .S0(n338), .Y(n576) );
  MUX21X1_HVT U365 ( .A1(n319), .A2(n270), .S0(n251), .Y(n578) );
  MUX21X1_HVT U366 ( .A1(n270), .A2(n277), .S0(n337), .Y(n405) );
  MUX21X1_HVT U367 ( .A1(n279), .A2(n328), .S0(n337), .Y(n410) );
  MUX21X1_HVT U368 ( .A1(n329), .A2(n279), .S0(n251), .Y(n408) );
  MUX21X1_HVT U369 ( .A1(n316), .A2(n279), .S0(n335), .Y(n403) );
  NBUFFX2_HVT U370 ( .A(in[2]), .Y(n341) );
  MUX21X1_HVT U371 ( .A1(n208), .A2(n281), .S0(n338), .Y(n588) );
  INVX0_HVT U372 ( .A(n593), .Y(n347) );
  INVX0_HVT U373 ( .A(n573), .Y(n348) );
  INVX0_HVT U374 ( .A(n567), .Y(n349) );
  INVX0_HVT U375 ( .A(n507), .Y(n350) );
  INVX0_HVT U376 ( .A(n468), .Y(n351) );
  INVX0_HVT U377 ( .A(n602), .Y(n352) );
  INVX0_HVT U378 ( .A(n599), .Y(n354) );
  INVX0_HVT U379 ( .A(n598), .Y(n356) );
  INVX0_HVT U380 ( .A(n597), .Y(n357) );
  INVX0_HVT U381 ( .A(n570), .Y(n358) );
  INVX0_HVT U382 ( .A(n591), .Y(n359) );
  INVX0_HVT U383 ( .A(n596), .Y(n360) );
  INVX0_HVT U384 ( .A(n592), .Y(n361) );
  INVX0_HVT U385 ( .A(n590), .Y(n362) );
  INVX0_HVT U386 ( .A(n589), .Y(n363) );
  INVX0_HVT U387 ( .A(n588), .Y(n364) );
  INVX0_HVT U388 ( .A(n587), .Y(n365) );
  INVX0_HVT U389 ( .A(n586), .Y(n366) );
  INVX0_HVT U390 ( .A(n585), .Y(n367) );
  INVX0_HVT U391 ( .A(n581), .Y(n369) );
  INVX0_HVT U392 ( .A(n578), .Y(n372) );
  INVX0_HVT U393 ( .A(n576), .Y(n373) );
  INVX0_HVT U394 ( .A(n575), .Y(n374) );
  INVX0_HVT U395 ( .A(n571), .Y(n376) );
  INVX0_HVT U396 ( .A(n568), .Y(n377) );
  INVX0_HVT U397 ( .A(n566), .Y(n378) );
  INVX0_HVT U398 ( .A(n560), .Y(n381) );
  INVX0_HVT U399 ( .A(n559), .Y(n382) );
  INVX0_HVT U400 ( .A(n595), .Y(n383) );
  INVX0_HVT U401 ( .A(n410), .Y(n385) );
  INVX0_HVT U402 ( .A(n408), .Y(n387) );
  INVX0_HVT U403 ( .A(n406), .Y(n389) );
  INVX0_HVT U404 ( .A(n405), .Y(n390) );
  INVX0_HVT U405 ( .A(n404), .Y(n391) );
  INVX0_HVT U406 ( .A(n403), .Y(n392) );
  INVX0_HVT U407 ( .A(n450), .Y(n393) );
  INVX0_HVT U408 ( .A(n402), .Y(n394) );
endmodule

