
module inv_sbox_5 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n196, n197, n198, n199, n200, n201, n202, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646;

  NAND2X0_HVT U3 ( .A1(n326), .A2(n335), .Y(n644) );
  NAND2X0_HVT U5 ( .A1(n643), .A2(n355), .Y(n642) );
  NAND2X0_HVT U6 ( .A1(n296), .A2(n361), .Y(n640) );
  NAND2X0_HVT U8 ( .A1(n366), .A2(n355), .Y(n638) );
  NAND2X0_HVT U9 ( .A1(n361), .A2(n638), .Y(n637) );
  NAND2X0_HVT U10 ( .A1(n360), .A2(n635), .Y(n636) );
  NAND2X0_HVT U11 ( .A1(n368), .A2(n359), .Y(n634) );
  NAND2X0_HVT U12 ( .A1(n299), .A2(n347), .Y(n633) );
  NAND2X0_HVT U13 ( .A1(n358), .A2(n638), .Y(n632) );
  NAND2X0_HVT U15 ( .A1(n259), .A2(n297), .Y(n630) );
  NAND2X0_HVT U19 ( .A1(n301), .A2(n434), .Y(n625) );
  NAND2X0_HVT U25 ( .A1(n335), .A2(n432), .Y(n641) );
  NAND2X0_HVT U32 ( .A1(n349), .A2(n368), .Y(n613) );
  NAND2X0_HVT U35 ( .A1(n638), .A2(n256), .Y(n610) );
  NAND2X0_HVT U38 ( .A1(n347), .A2(n368), .Y(n607) );
  NAND2X0_HVT U42 ( .A1(n640), .A2(n255), .Y(n603) );
  OA21X1_HVT U53 ( .A1(n374), .A2(n595), .A3(n303), .Y(n593) );
  NAND2X0_HVT U55 ( .A1(n358), .A2(n643), .Y(n591) );
  NAND2X0_HVT U66 ( .A1(n301), .A2(n290), .Y(n579) );
  MUX41X1_HVT U67 ( .A1(n391), .A3(n415), .A2(n393), .A4(n579), .S0(n346), 
        .S1(n336), .Y(n578) );
  MUX41X1_HVT U68 ( .A1(n391), .A3(n326), .A2(n392), .A4(n361), .S0(n339), 
        .S1(n372), .Y(n577) );
  NAND2X0_HVT U72 ( .A1(n259), .A2(n283), .Y(n574) );
  MUX41X1_HVT U73 ( .A1(n618), .A3(n574), .A2(n416), .A4(n347), .S0(n345), 
        .S1(n337), .Y(n573) );
  MUX41X1_HVT U74 ( .A1(n636), .A3(n406), .A2(n405), .A4(n397), .S0(n340), 
        .S1(n371), .Y(n572) );
  MUX41X1_HVT U80 ( .A1(n418), .A3(n414), .A2(n637), .A4(n642), .S0(n339), 
        .S1(n321), .Y(n566) );
  NAND2X0_HVT U81 ( .A1(n359), .A2(n237), .Y(n565) );
  AND2X1_HVT U82 ( .A1(n640), .A2(n357), .Y(n564) );
  MUX41X1_HVT U83 ( .A1(n564), .A3(n403), .A2(n419), .A4(n565), .S0(n339), 
        .S1(n370), .Y(n563) );
  MUX41X1_HVT U84 ( .A1(n333), .A3(n402), .A2(n420), .A4(n620), .S0(n340), 
        .S1(n321), .Y(n562) );
  NAND2X0_HVT U89 ( .A1(n368), .A2(n431), .Y(n558) );
  MUX41X1_HVT U90 ( .A1(n293), .A3(n283), .A2(n598), .A4(n558), .S0(n339), 
        .S1(n322), .Y(n557) );
  MUX41X1_HVT U96 ( .A1(n415), .A3(n632), .A2(n319), .A4(n422), .S0(n340), 
        .S1(n322), .Y(n551) );
  MUX41X1_HVT U98 ( .A1(n550), .A3(n423), .A2(n408), .A4(n617), .S0(n340), 
        .S1(n322), .Y(n549) );
  MUX41X1_HVT U99 ( .A1(n613), .A3(n395), .A2(n597), .A4(n259), .S0(n322), 
        .S1(n337), .Y(n548) );
  NAND2X0_HVT U100 ( .A1(n368), .A2(n430), .Y(n547) );
  MUX41X1_HVT U101 ( .A1(n424), .A3(n633), .A2(n407), .A4(n547), .S0(n322), 
        .S1(n336), .Y(n546) );
  MUX41X1_HVT U102 ( .A1(n546), .A3(n549), .A2(n548), .A4(n551), .S0(n354), 
        .S1(n351), .Y(n545) );
  AND2X1_HVT U104 ( .A1(n283), .A2(n641), .Y(n544) );
  MUX41X1_HVT U105 ( .A1(n631), .A3(n425), .A2(n565), .A4(n544), .S0(n340), 
        .S1(n371), .Y(n543) );
  MUX41X1_HVT U107 ( .A1(n424), .A3(n358), .A2(n542), .A4(n384), .S0(n339), 
        .S1(n370), .Y(n541) );
  MUX41X1_HVT U108 ( .A1(n397), .A3(n259), .A2(n401), .A4(n645), .S0(n340), 
        .S1(n322), .Y(n540) );
  MUX41X1_HVT U109 ( .A1(n423), .A3(n378), .A2(n420), .A4(n412), .S0(n339), 
        .S1(n321), .Y(n539) );
  MUX41X1_HVT U110 ( .A1(n539), .A3(n541), .A2(n540), .A4(n543), .S0(in[5]), 
        .S1(n352), .Y(n538) );
  AO21X1_HVT U112 ( .A1(n410), .A2(n345), .A3(n621), .Y(n536) );
  NAND2X0_HVT U114 ( .A1(n361), .A2(n283), .Y(n534) );
  MUX41X1_HVT U115 ( .A1(n534), .A3(n634), .A2(n410), .A4(n357), .S0(n370), 
        .S1(n337), .Y(n533) );
  MUX41X1_HVT U116 ( .A1(n409), .A3(n402), .A2(n378), .A4(n630), .S0(n338), 
        .S1(n321), .Y(n532) );
  NAND2X0_HVT U118 ( .A1(n368), .A2(n326), .Y(n530) );
  MUX41X1_HVT U119 ( .A1(n426), .A3(n531), .A2(n608), .A4(n530), .S0(n338), 
        .S1(n322), .Y(n529) );
  MUX41X1_HVT U120 ( .A1(n529), .A3(n533), .A2(n532), .A4(n535), .S0(n354), 
        .S1(n352), .Y(n528) );
  MUX41X1_HVT U122 ( .A1(n413), .A3(n329), .A2(n599), .A4(n417), .S0(n338), 
        .S1(n370), .Y(n527) );
  MUX41X1_HVT U124 ( .A1(n331), .A3(n526), .A2(n622), .A4(n325), .S0(n344), 
        .S1(n338), .Y(n525) );
  AOI21X1_HVT U127 ( .A1(n343), .A2(n521), .A3(n385), .Y(n522) );
  NAND2X0_HVT U129 ( .A1(n342), .A2(n360), .Y(n519) );
  MUX41X1_HVT U130 ( .A1(n519), .A3(n520), .A2(n523), .A4(n522), .S0(n346), 
        .S1(n352), .Y(n518) );
  AND2X1_HVT U131 ( .A1(n290), .A2(n318), .Y(n517) );
  MUX41X1_HVT U132 ( .A1(n382), .A3(n517), .A2(n428), .A4(n391), .S0(n345), 
        .S1(n337), .Y(n516) );
  MUX41X1_HVT U133 ( .A1(n429), .A3(n384), .A2(n591), .A4(n383), .S0(n344), 
        .S1(n336), .Y(n515) );
  MUX41X1_HVT U136 ( .A1(n596), .A3(n547), .A2(n513), .A4(n389), .S0(n342), 
        .S1(n321), .Y(n512) );
  MUX41X1_HVT U137 ( .A1(n315), .A3(n616), .A2(n620), .A4(n422), .S0(n346), 
        .S1(n336), .Y(n511) );
  MUX41X1_HVT U139 ( .A1(n510), .A3(n514), .A2(n518), .A4(n524), .S0(n354), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n405), .A3(n330), .A2(n400), .A4(n634), .S0(n345), 
        .S1(n336), .Y(n509) );
  NAND2X0_HVT U141 ( .A1(n260), .A2(n368), .Y(n508) );
  MUX41X1_HVT U142 ( .A1(n508), .A3(n606), .A2(n427), .A4(n400), .S0(n343), 
        .S1(n370), .Y(n507) );
  MUX41X1_HVT U145 ( .A1(n228), .A3(n425), .A2(n505), .A4(n565), .S0(n343), 
        .S1(n370), .Y(n504) );
  AO21X1_HVT U148 ( .A1(n346), .A2(n386), .A3(n430), .Y(n501) );
  MUX41X1_HVT U151 ( .A1(n419), .A3(n408), .A2(n398), .A4(n499), .S0(n344), 
        .S1(n336), .Y(n498) );
  MUX41X1_HVT U155 ( .A1(n400), .A3(n634), .A2(n626), .A4(n319), .S0(n341), 
        .S1(n321), .Y(n494) );
  MUX41X1_HVT U156 ( .A1(n494), .A3(n498), .A2(n495), .A4(n500), .S0(in[5]), 
        .S1(n352), .Y(n493) );
  NAND2X0_HVT U159 ( .A1(n490), .A2(n489), .Y(n491) );
  NAND2X0_HVT U163 ( .A1(n366), .A2(n431), .Y(n485) );
  MUX41X1_HVT U164 ( .A1(n637), .A3(n485), .A2(n608), .A4(n397), .S0(n338), 
        .S1(n321), .Y(n484) );
  NAND2X0_HVT U166 ( .A1(n635), .A2(n481), .Y(n482) );
  MUX41X1_HVT U173 ( .A1(n361), .A3(n293), .A2(n645), .A4(n609), .S0(n341), 
        .S1(n371), .Y(n474) );
  MUX41X1_HVT U174 ( .A1(n421), .A3(n591), .A2(n429), .A4(n252), .S0(n341), 
        .S1(n322), .Y(n473) );
  NAND2X0_HVT U177 ( .A1(n300), .A2(n326), .Y(n471) );
  MUX41X1_HVT U178 ( .A1(n332), .A3(n471), .A2(n293), .A4(n601), .S0(n341), 
        .S1(n372), .Y(n470) );
  AND2X1_HVT U179 ( .A1(n640), .A2(n641), .Y(n469) );
  MUX41X1_HVT U180 ( .A1(n613), .A3(n376), .A2(n469), .A4(n600), .S0(n341), 
        .S1(n372), .Y(n468) );
  MUX41X1_HVT U182 ( .A1(n384), .A3(n267), .A2(n381), .A4(n419), .S0(n338), 
        .S1(n372), .Y(n466) );
  AND2X1_HVT U185 ( .A1(n251), .A2(n318), .Y(n463) );
  AND2X1_HVT U192 ( .A1(n406), .A2(n455), .Y(n456) );
  NAND2X0_HVT U194 ( .A1(n603), .A2(n455), .Y(n453) );
  NAND2X0_HVT U198 ( .A1(n299), .A2(n256), .Y(n635) );
  NAND2X0_HVT U200 ( .A1(n355), .A2(n368), .Y(n521) );
  NAND2X0_HVT U207 ( .A1(n368), .A2(n293), .Y(n585) );
  INVX0_HVT U1 ( .A(n376), .Y(n196) );
  MUX21X2_HVT U2 ( .A1(n620), .A2(n333), .S0(n345), .Y(n497) );
  MUX21X2_HVT U4 ( .A1(n641), .A2(n358), .S0(n366), .Y(n487) );
  MUX21X1_HVT U7 ( .A1(n347), .A2(n430), .S0(n297), .Y(n615) );
  MUX21X1_HVT U14 ( .A1(n430), .A2(n304), .S0(n296), .Y(n595) );
  AO21X1_HVT U16 ( .A1(n297), .A2(n430), .A3(n374), .Y(n455) );
  INVX0_HVT U17 ( .A(n620), .Y(n400) );
  INVX0_HVT U18 ( .A(n616), .Y(n402) );
  IBUFFX2_HVT U20 ( .A(n364), .Y(n238) );
  MUX41X1_HVT U21 ( .A1(n572), .A3(n575), .A2(n569), .A4(n573), .S0(n354), 
        .S1(n197), .Y(n568) );
  IBUFFX16_HVT U22 ( .A(n351), .Y(n197) );
  MUX21X2_HVT U23 ( .A1(n416), .A2(n604), .S0(n345), .Y(n460) );
  MUX21X2_HVT U24 ( .A1(n428), .A2(n382), .S0(n344), .Y(n502) );
  MUX21X1_HVT U26 ( .A1(n347), .A2(n434), .S0(n364), .Y(n602) );
  IBUFFX2_HVT U27 ( .A(n602), .Y(n411) );
  INVX0_HVT U28 ( .A(n356), .Y(n304) );
  MUX21X1_HVT U29 ( .A1(n397), .A2(n582), .S0(n334), .Y(n581) );
  MUX21X2_HVT U30 ( .A1(n349), .A2(n259), .S0(n285), .Y(n620) );
  IBUFFX2_HVT U31 ( .A(n364), .Y(n285) );
  AOI21X1_HVT U33 ( .A1(n616), .A2(n198), .A3(n199), .Y(n459) );
  IBUFFX16_HVT U34 ( .A(n374), .Y(n198) );
  IBUFFX16_HVT U36 ( .A(n585), .Y(n199) );
  MUX41X1_HVT U37 ( .A1(n480), .A3(n486), .A2(n484), .A4(n488), .S0(n200), 
        .S1(n201), .Y(n479) );
  IBUFFX16_HVT U39 ( .A(n353), .Y(n200) );
  IBUFFX16_HVT U40 ( .A(n350), .Y(n201) );
  MUX41X1_HVT U41 ( .A1(n404), .A3(n402), .A2(n628), .A4(n627), .S0(n270), 
        .S1(n223), .Y(n567) );
  NAND2X0_HVT U43 ( .A1(n259), .A2(n202), .Y(n218) );
  NAND2X0_HVT U44 ( .A1(n433), .A2(n366), .Y(n219) );
  NAND2X0_HVT U45 ( .A1(n218), .A2(n219), .Y(n614) );
  IBUFFX2_HVT U46 ( .A(n366), .Y(n202) );
  MUX21X1_HVT U47 ( .A1(n290), .A2(n360), .S0(n296), .Y(n628) );
  INVX1_HVT U48 ( .A(n269), .Y(n223) );
  IBUFFX2_HVT U49 ( .A(n370), .Y(n270) );
  INVX2_HVT U50 ( .A(n302), .Y(n366) );
  INVX0_HVT U51 ( .A(n614), .Y(n404) );
  MUX41X1_HVT U52 ( .A1(n323), .A3(n396), .A2(n610), .A4(n487), .S0(n220), 
        .S1(n372), .Y(n486) );
  IBUFFX16_HVT U54 ( .A(n236), .Y(n220) );
  MUX21X2_HVT U56 ( .A1(n470), .A2(n468), .S0(n350), .Y(n467) );
  MUX41X1_HVT U57 ( .A1(n623), .A3(n328), .A2(n476), .A4(n558), .S0(n221), 
        .S1(n222), .Y(n475) );
  IBUFFX16_HVT U58 ( .A(n341), .Y(n221) );
  IBUFFX16_HVT U59 ( .A(n371), .Y(n222) );
  INVX1_HVT U60 ( .A(n645), .Y(n430) );
  AO21X1_HVT U61 ( .A1(n318), .A2(n360), .A3(n374), .Y(n489) );
  INVX0_HVT U62 ( .A(n360), .Y(n433) );
  INVX0_HVT U63 ( .A(n348), .Y(n294) );
  IBUFFX2_HVT U64 ( .A(n302), .Y(n365) );
  INVX1_HVT U65 ( .A(n302), .Y(n248) );
  IBUFFX2_HVT U69 ( .A(n436), .Y(n335) );
  IBUFFX2_HVT U70 ( .A(n436), .Y(n290) );
  IBUFFX2_HVT U71 ( .A(n351), .Y(n227) );
  INVX1_HVT U75 ( .A(n385), .Y(n237) );
  NAND2X0_HVT U76 ( .A1(n527), .A2(n224), .Y(n225) );
  NAND2X0_HVT U77 ( .A1(n525), .A2(n268), .Y(n226) );
  NAND2X0_HVT U78 ( .A1(n225), .A2(n226), .Y(n524) );
  INVX0_HVT U79 ( .A(n268), .Y(n224) );
  MUX41X1_HVT U85 ( .A1(n563), .A3(n567), .A2(n562), .A4(n566), .S0(n354), 
        .S1(n227), .Y(n561) );
  INVX0_HVT U86 ( .A(n404), .Y(n228) );
  NAND2X0_HVT U87 ( .A1(n466), .A2(n229), .Y(n230) );
  NAND2X0_HVT U88 ( .A1(n465), .A2(n350), .Y(n231) );
  NAND2X0_HVT U91 ( .A1(n230), .A2(n231), .Y(n464) );
  IBUFFX2_HVT U92 ( .A(n350), .Y(n229) );
  INVX1_HVT U93 ( .A(in[1]), .Y(n350) );
  MUX41X1_HVT U94 ( .A1(n590), .A3(n584), .A2(n592), .A4(n588), .S0(n232), 
        .S1(n279), .Y(n583) );
  IBUFFX16_HVT U95 ( .A(n354), .Y(n232) );
  MUX21X2_HVT U97 ( .A1(n597), .A2(n333), .S0(n233), .Y(n461) );
  IBUFFX16_HVT U103 ( .A(n346), .Y(n233) );
  MUX41X1_HVT U106 ( .A1(n397), .A3(n603), .A2(n411), .A4(n414), .S0(n344), 
        .S1(n234), .Y(n465) );
  IBUFFX16_HVT U111 ( .A(n337), .Y(n234) );
  MUX21X1_HVT U113 ( .A1(n252), .A2(n347), .S0(n235), .Y(n446) );
  IBUFFX16_HVT U117 ( .A(n301), .Y(n235) );
  MUX21X2_HVT U121 ( .A1(n359), .A2(n358), .S0(n238), .Y(n627) );
  MUX21X2_HVT U123 ( .A1(n593), .A2(n594), .S0(n306), .Y(n592) );
  IBUFFX16_HVT U125 ( .A(n341), .Y(n236) );
  INVX1_HVT U126 ( .A(n639), .Y(n385) );
  MUX21X2_HVT U128 ( .A1(n528), .A2(n538), .S0(in[7]), .Y(out[3]) );
  INVX1_HVT U134 ( .A(n446), .Y(n419) );
  MUX21X2_HVT U135 ( .A1(n417), .A2(n602), .S0(n239), .Y(n492) );
  IBUFFX16_HVT U138 ( .A(n345), .Y(n239) );
  MUX41X1_HVT U143 ( .A1(n387), .A3(n196), .A2(n293), .A4(n640), .S0(n240), 
        .S1(n241), .Y(n575) );
  IBUFFX16_HVT U144 ( .A(n339), .Y(n240) );
  IBUFFX16_HVT U146 ( .A(n371), .Y(n241) );
  NAND2X0_HVT U147 ( .A1(n552), .A2(n242), .Y(n243) );
  NAND2X0_HVT U149 ( .A1(n545), .A2(n291), .Y(n244) );
  NAND2X0_HVT U150 ( .A1(n243), .A2(n244), .Y(out[2]) );
  IBUFFX2_HVT U152 ( .A(n291), .Y(n242) );
  INVX2_HVT U153 ( .A(n282), .Y(n283) );
  NAND2X0_HVT U154 ( .A1(n570), .A2(n245), .Y(n246) );
  NAND2X0_HVT U157 ( .A1(n571), .A2(n286), .Y(n247) );
  NAND2X0_HVT U158 ( .A1(n246), .A2(n247), .Y(n569) );
  INVX0_HVT U160 ( .A(n286), .Y(n245) );
  MUX21X1_HVT U161 ( .A1(n304), .A2(n347), .S0(n365), .Y(n448) );
  MUX21X1_HVT U162 ( .A1(n284), .A2(n377), .S0(n346), .Y(n571) );
  IBUFFX2_HVT U165 ( .A(n343), .Y(n286) );
  IBUFFX2_HVT U167 ( .A(n638), .Y(n386) );
  MUX21X2_HVT U168 ( .A1(n387), .A2(n260), .S0(n346), .Y(n554) );
  INVX1_HVT U169 ( .A(n305), .Y(n249) );
  INVX1_HVT U170 ( .A(n305), .Y(n250) );
  INVX1_HVT U171 ( .A(n249), .Y(n251) );
  INVX1_HVT U172 ( .A(n250), .Y(n252) );
  INVX1_HVT U175 ( .A(n435), .Y(n253) );
  INVX1_HVT U176 ( .A(n435), .Y(n254) );
  INVX1_HVT U181 ( .A(n253), .Y(n255) );
  INVX1_HVT U183 ( .A(n254), .Y(n256) );
  IBUFFX2_HVT U184 ( .A(n629), .Y(n257) );
  IBUFFX2_HVT U186 ( .A(n629), .Y(n258) );
  INVX2_HVT U187 ( .A(n257), .Y(n259) );
  INVX2_HVT U188 ( .A(n258), .Y(n260) );
  XNOR2X1_HVT U189 ( .A1(n335), .A2(in[3]), .Y(n629) );
  AO21X2_HVT U190 ( .A1(n585), .A2(n344), .A3(n624), .Y(n586) );
  NAND2X0_HVT U191 ( .A1(n399), .A2(n261), .Y(n262) );
  NAND2X0_HVT U193 ( .A1(n589), .A2(n334), .Y(n263) );
  NAND2X0_HVT U195 ( .A1(n262), .A2(n263), .Y(n588) );
  INVX0_HVT U196 ( .A(n334), .Y(n261) );
  MUX21X1_HVT U197 ( .A1(n642), .A2(n400), .S0(n306), .Y(n589) );
  NAND2X0_HVT U199 ( .A1(n358), .A2(n264), .Y(n265) );
  NAND2X0_HVT U201 ( .A1(n556), .A2(n318), .Y(n266) );
  NAND2X0_HVT U202 ( .A1(n265), .A2(n266), .Y(n555) );
  IBUFFX2_HVT U203 ( .A(n318), .Y(n264) );
  NBUFFX4_HVT U204 ( .A(n302), .Y(n318) );
  IBUFFX2_HVT U205 ( .A(n615), .Y(n403) );
  IBUFFX2_HVT U206 ( .A(n352), .Y(n268) );
  INVX1_HVT U208 ( .A(n381), .Y(n267) );
  INVX0_HVT U209 ( .A(in[7]), .Y(n291) );
  MUX21X1_HVT U210 ( .A1(n260), .A2(n347), .S0(n296), .Y(n624) );
  IBUFFX16_HVT U211 ( .A(n340), .Y(n269) );
  MUX21X2_HVT U212 ( .A1(n501), .A2(n502), .S0(n306), .Y(n500) );
  MUX41X1_HVT U213 ( .A1(n460), .A3(n459), .A2(n461), .A4(n462), .S0(n337), 
        .S1(n351), .Y(n458) );
  MUX21X1_HVT U214 ( .A1(n645), .A2(n347), .S0(n271), .Y(n325) );
  IBUFFX16_HVT U215 ( .A(n318), .Y(n271) );
  INVX0_HVT U216 ( .A(n325), .Y(n622) );
  INVX0_HVT U217 ( .A(n643), .Y(n381) );
  NAND2X0_HVT U218 ( .A1(n260), .A2(n272), .Y(n273) );
  NAND2X0_HVT U219 ( .A1(n433), .A2(n280), .Y(n274) );
  NAND2X0_HVT U220 ( .A1(n273), .A2(n274), .Y(n444) );
  INVX0_HVT U221 ( .A(n280), .Y(n272) );
  INVX0_HVT U222 ( .A(n444), .Y(n421) );
  NAND2X0_HVT U223 ( .A1(n586), .A2(n275), .Y(n276) );
  NAND2X0_HVT U224 ( .A1(n587), .A2(n306), .Y(n277) );
  NAND2X0_HVT U225 ( .A1(n276), .A2(n277), .Y(n584) );
  IBUFFX2_HVT U226 ( .A(n306), .Y(n275) );
  MUX21X1_HVT U227 ( .A1(n325), .A2(n591), .S0(n345), .Y(n587) );
  INVX0_HVT U228 ( .A(n343), .Y(n306) );
  MUX41X1_HVT U229 ( .A1(n421), .A3(n401), .A2(n381), .A4(n333), .S0(n338), 
        .S1(n278), .Y(n560) );
  IBUFFX16_HVT U230 ( .A(n371), .Y(n278) );
  IBUFFX16_HVT U231 ( .A(n350), .Y(n279) );
  INVX2_HVT U232 ( .A(n350), .Y(n352) );
  NBUFFX4_HVT U233 ( .A(n432), .Y(n347) );
  IBUFFX2_HVT U234 ( .A(n299), .Y(n280) );
  MUX41X1_HVT U235 ( .A1(n464), .A3(n452), .A2(n467), .A4(n458), .S0(n320), 
        .S1(n281), .Y(out[7]) );
  IBUFFX16_HVT U236 ( .A(n353), .Y(n281) );
  INVX1_HVT U237 ( .A(n639), .Y(n282) );
  OR2X1_HVT U238 ( .A1(n318), .A2(n304), .Y(n639) );
  INVX0_HVT U239 ( .A(n448), .Y(n284) );
  INVX0_HVT U240 ( .A(n448), .Y(n417) );
  NBUFFX2_HVT U241 ( .A(n645), .Y(n359) );
  INVX2_HVT U242 ( .A(n363), .Y(n302) );
  INVX1_HVT U243 ( .A(n450), .Y(n415) );
  INVX1_HVT U244 ( .A(n624), .Y(n397) );
  IBUFFX2_HVT U245 ( .A(n629), .Y(n305) );
  IBUFFX2_HVT U246 ( .A(n629), .Y(n435) );
  INVX1_HVT U247 ( .A(n356), .Y(n434) );
  NAND2X2_HVT U248 ( .A1(n432), .A2(n348), .Y(n645) );
  MUX41X1_HVT U249 ( .A1(n599), .A3(n615), .A2(n378), .A4(n393), .S0(n287), 
        .S1(n288), .Y(n559) );
  IBUFFX16_HVT U250 ( .A(n339), .Y(n287) );
  IBUFFX16_HVT U251 ( .A(n371), .Y(n288) );
  NBUFFX2_HVT U252 ( .A(n436), .Y(n348) );
  INVX1_HVT U253 ( .A(n292), .Y(n604) );
  INVX1_HVT U254 ( .A(n342), .Y(n289) );
  NBUFFX2_HVT U255 ( .A(in[2]), .Y(n342) );
  MUX21X2_HVT U256 ( .A1(n568), .A2(n561), .S0(n291), .Y(out[1]) );
  INVX1_HVT U257 ( .A(in[6]), .Y(n436) );
  MUX21X2_HVT U258 ( .A1(n576), .A2(n583), .S0(in[7]), .Y(out[0]) );
  AO21X1_HVT U259 ( .A1(n259), .A2(n267), .A3(n374), .Y(n481) );
  NBUFFX16_HVT U260 ( .A(n369), .Y(n343) );
  MUX21X1_HVT U261 ( .A1(n536), .A2(n537), .S0(n343), .Y(n535) );
  OA21X1_HVT U262 ( .A1(n380), .A2(n374), .A3(n624), .Y(n570) );
  INVX0_HVT U263 ( .A(n367), .Y(n363) );
  MUX21X1_HVT U264 ( .A1(n436), .A2(n356), .S0(n301), .Y(n292) );
  INVX2_HVT U265 ( .A(in[4]), .Y(n375) );
  INVX1_HVT U266 ( .A(n646), .Y(n293) );
  OR2X1_HVT U267 ( .A1(n432), .A2(n294), .Y(n646) );
  INVX1_HVT U268 ( .A(n432), .Y(n326) );
  INVX1_HVT U269 ( .A(n375), .Y(n373) );
  INVX1_HVT U270 ( .A(in[3]), .Y(n432) );
  NBUFFX16_HVT U271 ( .A(n373), .Y(n345) );
  MUX41X1_HVT U272 ( .A1(n475), .A3(n477), .A2(n473), .A4(n474), .S0(n351), 
        .S1(n295), .Y(n472) );
  IBUFFX16_HVT U273 ( .A(n354), .Y(n295) );
  MUX21X1_HVT U274 ( .A1(n434), .A2(n433), .S0(n367), .Y(n478) );
  NBUFFX2_HVT U275 ( .A(n365), .Y(n296) );
  NBUFFX2_HVT U276 ( .A(n365), .Y(n297) );
  NBUFFX2_HVT U277 ( .A(n363), .Y(n298) );
  NBUFFX2_HVT U278 ( .A(n301), .Y(n299) );
  NBUFFX2_HVT U279 ( .A(n364), .Y(n300) );
  IBUFFX2_HVT U280 ( .A(n367), .Y(n364) );
  INVX0_HVT U281 ( .A(n323), .Y(n601) );
  NAND2X0_HVT U282 ( .A1(n364), .A2(n359), .Y(n643) );
  INVX0_HVT U283 ( .A(n303), .Y(n617) );
  MUX21X1_HVT U284 ( .A1(n324), .A2(n331), .S0(n344), .Y(n454) );
  NAND2X0_HVT U285 ( .A1(n374), .A2(n390), .Y(n457) );
  INVX1_HVT U286 ( .A(in[5]), .Y(n353) );
  INVX1_HVT U287 ( .A(n618), .Y(n319) );
  INVX1_HVT U288 ( .A(n353), .Y(n354) );
  INVX1_HVT U289 ( .A(n350), .Y(n351) );
  INVX0_HVT U290 ( .A(in[7]), .Y(n320) );
  INVX1_HVT U291 ( .A(n372), .Y(n327) );
  MUX21X2_HVT U292 ( .A1(n392), .A2(n319), .S0(n327), .Y(n594) );
  INVX0_HVT U293 ( .A(n367), .Y(n301) );
  INVX1_HVT U294 ( .A(in[0]), .Y(n367) );
  MUX21X1_HVT U295 ( .A1(n360), .A2(n355), .S0(n300), .Y(n303) );
  XNOR2X1_HVT U296 ( .A1(n251), .A2(n248), .Y(n599) );
  MUX21X1_HVT U297 ( .A1(n385), .A2(n604), .S0(n346), .Y(n537) );
  IBUFFX2_HVT U298 ( .A(n599), .Y(n412) );
  MUX21X2_HVT U299 ( .A1(n503), .A2(n493), .S0(n320), .Y(out[5]) );
  NAND2X0_HVT U300 ( .A1(n491), .A2(n289), .Y(n307) );
  NAND2X0_HVT U301 ( .A1(n492), .A2(n343), .Y(n308) );
  NAND2X0_HVT U302 ( .A1(n308), .A2(n307), .Y(n488) );
  NAND2X0_HVT U303 ( .A1(n472), .A2(n320), .Y(n309) );
  NAND2X0_HVT U304 ( .A1(n479), .A2(in[7]), .Y(n310) );
  NAND2X0_HVT U305 ( .A1(n309), .A2(n310), .Y(out[6]) );
  MUX41X1_HVT U306 ( .A1(n553), .A3(n557), .A2(n559), .A4(n560), .S0(in[1]), 
        .S1(n354), .Y(n552) );
  NAND2X0_HVT U307 ( .A1(n554), .A2(n289), .Y(n311) );
  NAND2X0_HVT U308 ( .A1(n555), .A2(n342), .Y(n312) );
  NAND2X0_HVT U309 ( .A1(n312), .A2(n311), .Y(n553) );
  NAND2X0_HVT U310 ( .A1(n482), .A2(n289), .Y(n313) );
  NAND2X0_HVT U311 ( .A1(n483), .A2(n342), .Y(n314) );
  NAND2X0_HVT U312 ( .A1(n313), .A2(n314), .Y(n480) );
  MUX21X1_HVT U313 ( .A1(n619), .A2(n622), .S0(n344), .Y(n483) );
  MUX41X1_HVT U314 ( .A1(n454), .A3(n456), .A2(n453), .A4(n457), .S0(n352), 
        .S1(n339), .Y(n452) );
  MUX21X1_HVT U315 ( .A1(n398), .A2(n267), .S0(n342), .Y(n582) );
  INVX0_HVT U316 ( .A(n386), .Y(n315) );
  IBUFFX2_HVT U317 ( .A(n324), .Y(n600) );
  MUX21X2_HVT U318 ( .A1(n496), .A2(n497), .S0(n343), .Y(n495) );
  INVX1_HVT U319 ( .A(n298), .Y(n368) );
  NAND2X0_HVT U320 ( .A1(n463), .A2(n327), .Y(n316) );
  NAND2X0_HVT U321 ( .A1(n418), .A2(n344), .Y(n317) );
  NAND2X0_HVT U322 ( .A1(n316), .A2(n317), .Y(n462) );
  INVX1_HVT U323 ( .A(n449), .Y(n416) );
  MUX21X1_HVT U324 ( .A1(n359), .A2(n347), .S0(n368), .Y(n447) );
  INVX1_HVT U325 ( .A(n447), .Y(n418) );
  MUX41X1_HVT U326 ( .A1(n581), .A3(n578), .A2(n580), .A4(n577), .S0(n353), 
        .S1(n350), .Y(n576) );
  INVX1_HVT U327 ( .A(n375), .Y(n321) );
  INVX1_HVT U328 ( .A(n375), .Y(n322) );
  IBUFFX2_HVT U329 ( .A(in[4]), .Y(n374) );
  INVX1_HVT U330 ( .A(n375), .Y(n372) );
  MUX21X1_HVT U331 ( .A1(n641), .A2(n360), .S0(n297), .Y(n323) );
  INVX2_HVT U332 ( .A(n375), .Y(n370) );
  MUX21X1_HVT U333 ( .A1(n326), .A2(n290), .S0(n301), .Y(n324) );
  IBUFFX2_HVT U334 ( .A(n375), .Y(n371) );
  IBUFFX2_HVT U335 ( .A(n367), .Y(n362) );
  MUX41X1_HVT U336 ( .A1(n591), .A3(n401), .A2(n260), .A4(n414), .S0(n306), 
        .S1(n374), .Y(n590) );
  OA21X2_HVT U337 ( .A1(n379), .A2(n374), .A3(n388), .Y(n496) );
  MUX41X1_HVT U338 ( .A1(n507), .A3(n509), .A2(n504), .A4(n506), .S0(n352), 
        .S1(n353), .Y(n503) );
  MUX41X1_HVT U339 ( .A1(n607), .A3(n395), .A2(n396), .A4(n394), .S0(n289), 
        .S1(n374), .Y(n580) );
  MUX41X1_HVT U340 ( .A1(n478), .A3(n331), .A2(n328), .A4(n332), .S0(n289), 
        .S1(n327), .Y(n477) );
  MUX41X1_HVT U341 ( .A1(n622), .A3(n625), .A2(n411), .A4(n431), .S0(n289), 
        .S1(n327), .Y(n506) );
  MUX21X2_HVT U342 ( .A1(n511), .A2(n512), .S0(in[1]), .Y(n510) );
  MUX21X2_HVT U343 ( .A1(n515), .A2(n516), .S0(n352), .Y(n514) );
  AND2X1_HVT U344 ( .A1(n640), .A2(n359), .Y(n328) );
  AND2X1_HVT U345 ( .A1(n359), .A2(n630), .Y(n329) );
  MUX21X1_HVT U346 ( .A1(n255), .A2(n430), .S0(n362), .Y(n623) );
  MUX21X1_HVT U347 ( .A1(n430), .A2(n256), .S0(n300), .Y(n612) );
  MUX21X1_HVT U348 ( .A1(n349), .A2(n430), .S0(n364), .Y(n619) );
  MUX21X1_HVT U349 ( .A1(n349), .A2(n431), .S0(n366), .Y(n499) );
  MUX21X1_HVT U350 ( .A1(n433), .A2(n349), .S0(n366), .Y(n476) );
  MUX21X1_HVT U351 ( .A1(n430), .A2(n349), .S0(n297), .Y(n449) );
  INVX1_HVT U352 ( .A(n641), .Y(n431) );
  MUX21X1_HVT U353 ( .A1(n255), .A2(n347), .S0(n297), .Y(n606) );
  MUX21X1_HVT U354 ( .A1(n349), .A2(n252), .S0(n362), .Y(n609) );
  MUX21X1_HVT U355 ( .A1(n612), .A2(n329), .S0(n343), .Y(n520) );
  MUX21X1_HVT U356 ( .A1(n645), .A2(n355), .S0(n297), .Y(n505) );
  MUX21X1_HVT U357 ( .A1(n427), .A2(n330), .S0(n342), .Y(n523) );
  MUX21X1_HVT U358 ( .A1(n251), .A2(n436), .S0(n364), .Y(n439) );
  MUX21X1_HVT U359 ( .A1(n641), .A2(n359), .S0(n364), .Y(n438) );
  MUX21X1_HVT U360 ( .A1(n259), .A2(n349), .S0(n345), .Y(n556) );
  XOR2X1_HVT U361 ( .A1(n356), .A2(n299), .Y(n598) );
  XOR2X1_HVT U362 ( .A1(n641), .A2(n362), .Y(n597) );
  XNOR2X1_HVT U363 ( .A1(n645), .A2(n299), .Y(n330) );
  MUX21X1_HVT U364 ( .A1(n260), .A2(n431), .S0(n300), .Y(n611) );
  MUX21X1_HVT U365 ( .A1(n360), .A2(n359), .S0(n248), .Y(n631) );
  MUX21X1_HVT U366 ( .A1(n349), .A2(n359), .S0(n299), .Y(n542) );
  MUX21X1_HVT U367 ( .A1(n349), .A2(n260), .S0(n366), .Y(n605) );
  MUX21X1_HVT U368 ( .A1(n357), .A2(n347), .S0(n364), .Y(n626) );
  MUX21X1_HVT U369 ( .A1(n357), .A2(n349), .S0(n362), .Y(n526) );
  XOR2X1_HVT U370 ( .A1(n360), .A2(n296), .Y(n608) );
  MUX21X1_HVT U371 ( .A1(n347), .A2(n357), .S0(n301), .Y(n441) );
  NBUFFX2_HVT U372 ( .A(n373), .Y(n344) );
  NBUFFX2_HVT U373 ( .A(n373), .Y(n346) );
  AND2X1_HVT U374 ( .A1(n248), .A2(n349), .Y(n331) );
  NBUFFX2_HVT U375 ( .A(n646), .Y(n360) );
  AND2X1_HVT U376 ( .A1(n434), .A2(n368), .Y(n332) );
  NBUFFX2_HVT U377 ( .A(n641), .Y(n355) );
  NBUFFX2_HVT U378 ( .A(n644), .Y(n356) );
  AND2X1_HVT U379 ( .A1(n357), .A2(n368), .Y(n333) );
  NBUFFX2_HVT U380 ( .A(n644), .Y(n358) );
  NBUFFX2_HVT U381 ( .A(n646), .Y(n361) );
  NBUFFX2_HVT U382 ( .A(n644), .Y(n357) );
  NBUFFX2_HVT U383 ( .A(n342), .Y(n341) );
  XNOR2X1_HVT U384 ( .A1(n374), .A2(n338), .Y(n334) );
  NBUFFX2_HVT U385 ( .A(n436), .Y(n349) );
  NBUFFX2_HVT U386 ( .A(n369), .Y(n338) );
  NBUFFX2_HVT U387 ( .A(n369), .Y(n340) );
  NBUFFX2_HVT U388 ( .A(n369), .Y(n339) );
  NBUFFX2_HVT U389 ( .A(n369), .Y(n337) );
  NBUFFX2_HVT U390 ( .A(n369), .Y(n336) );
  MUX21X1_HVT U391 ( .A1(n355), .A2(n326), .S0(n362), .Y(n550) );
  MUX21X1_HVT U392 ( .A1(n433), .A2(n326), .S0(n366), .Y(n437) );
  MUX21X1_HVT U393 ( .A1(n434), .A2(n431), .S0(n300), .Y(n531) );
  MUX21X1_HVT U394 ( .A1(n326), .A2(n355), .S0(n362), .Y(n442) );
  MUX21X1_HVT U395 ( .A1(n361), .A2(n326), .S0(n366), .Y(n490) );
  MUX21X1_HVT U396 ( .A1(n326), .A2(n361), .S0(n300), .Y(n443) );
  MUX21X1_HVT U397 ( .A1(n349), .A2(n326), .S0(n296), .Y(n618) );
  NBUFFX2_HVT U398 ( .A(in[2]), .Y(n369) );
  MUX21X1_HVT U399 ( .A1(n430), .A2(n290), .S0(n301), .Y(n513) );
  MUX21X1_HVT U400 ( .A1(n290), .A2(n293), .S0(n362), .Y(n621) );
  XOR2X1_HVT U401 ( .A1(n362), .A2(n290), .Y(n596) );
  MUX21X1_HVT U402 ( .A1(n357), .A2(n290), .S0(n297), .Y(n445) );
  MUX21X1_HVT U403 ( .A1(n290), .A2(n358), .S0(n301), .Y(n450) );
  MUX21X1_HVT U404 ( .A1(n347), .A2(n290), .S0(n301), .Y(n440) );
  MUX21X1_HVT U405 ( .A1(n355), .A2(n290), .S0(n364), .Y(n616) );
  MUX21X1_HVT U406 ( .A1(n290), .A2(n431), .S0(n362), .Y(n451) );
  INVX0_HVT U407 ( .A(n634), .Y(n376) );
  INVX0_HVT U408 ( .A(n613), .Y(n377) );
  INVX0_HVT U409 ( .A(n607), .Y(n378) );
  INVX0_HVT U410 ( .A(n547), .Y(n379) );
  INVX0_HVT U411 ( .A(n508), .Y(n380) );
  INVX0_HVT U412 ( .A(n642), .Y(n382) );
  INVX0_HVT U413 ( .A(n640), .Y(n383) );
  INVX0_HVT U414 ( .A(n603), .Y(n384) );
  INVX0_HVT U415 ( .A(n610), .Y(n387) );
  INVX0_HVT U416 ( .A(n632), .Y(n388) );
  INVX0_HVT U417 ( .A(n637), .Y(n389) );
  INVX0_HVT U418 ( .A(n633), .Y(n390) );
  INVX0_HVT U419 ( .A(n631), .Y(n391) );
  INVX0_HVT U420 ( .A(n630), .Y(n392) );
  INVX0_HVT U421 ( .A(n628), .Y(n393) );
  INVX0_HVT U422 ( .A(n627), .Y(n394) );
  INVX0_HVT U423 ( .A(n626), .Y(n395) );
  INVX0_HVT U424 ( .A(n625), .Y(n396) );
  INVX0_HVT U425 ( .A(n623), .Y(n398) );
  INVX0_HVT U426 ( .A(n621), .Y(n399) );
  INVX0_HVT U427 ( .A(n619), .Y(n401) );
  INVX0_HVT U428 ( .A(n612), .Y(n405) );
  INVX0_HVT U429 ( .A(n611), .Y(n406) );
  INVX0_HVT U430 ( .A(n609), .Y(n407) );
  INVX0_HVT U431 ( .A(n608), .Y(n408) );
  INVX0_HVT U432 ( .A(n606), .Y(n409) );
  INVX0_HVT U433 ( .A(n605), .Y(n410) );
  INVX0_HVT U434 ( .A(n636), .Y(n413) );
  INVX0_HVT U435 ( .A(n451), .Y(n414) );
  INVX0_HVT U436 ( .A(n445), .Y(n420) );
  INVX0_HVT U437 ( .A(n443), .Y(n422) );
  INVX0_HVT U438 ( .A(n442), .Y(n423) );
  INVX0_HVT U439 ( .A(n441), .Y(n424) );
  INVX0_HVT U440 ( .A(n440), .Y(n425) );
  INVX0_HVT U441 ( .A(n490), .Y(n426) );
  INVX0_HVT U442 ( .A(n439), .Y(n427) );
  INVX0_HVT U443 ( .A(n438), .Y(n428) );
  INVX0_HVT U444 ( .A(n437), .Y(n429) );
endmodule

