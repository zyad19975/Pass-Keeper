
module sbox_15 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n38, n114, n117, n210, n211, n212, n213, n216, n217, n218, n219,
         n226, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629;

  NAND2X0_HVT U3 ( .A1(n255), .A2(n340), .Y(n627) );
  NAND2X0_HVT U4 ( .A1(n338), .A2(n270), .Y(n626) );
  NAND2X0_HVT U5 ( .A1(n348), .A2(n409), .Y(n624) );
  NAND2X0_HVT U15 ( .A1(n268), .A2(n327), .Y(n614) );
  NAND2X0_HVT U21 ( .A1(n338), .A2(n350), .Y(n608) );
  NAND2X0_HVT U24 ( .A1(n333), .A2(n350), .Y(n606) );
  NAND2X0_HVT U33 ( .A1(n278), .A2(n350), .Y(n597) );
  NAND2X0_HVT U35 ( .A1(n330), .A2(n350), .Y(n595) );
  NAND2X0_HVT U42 ( .A1(n344), .A2(n333), .Y(n589) );
  MUX41X1_HVT U51 ( .A1(n397), .A3(n358), .A2(n376), .A4(n377), .S0(n354), 
        .S1(n257), .Y(n580) );
  NAND2X0_HVT U53 ( .A1(n577), .A2(n588), .Y(n578) );
  NAND2X0_HVT U56 ( .A1(n338), .A2(n573), .Y(n574) );
  NAND2X0_HVT U58 ( .A1(n342), .A2(n270), .Y(n571) );
  MUX41X1_HVT U59 ( .A1(n313), .A3(n571), .A2(n311), .A4(n375), .S0(n354), 
        .S1(n257), .Y(n570) );
  MUX41X1_HVT U61 ( .A1(n309), .A3(n374), .A2(n373), .A4(n326), .S0(n355), 
        .S1(n263), .Y(n568) );
  NAND2X0_HVT U62 ( .A1(n350), .A2(n341), .Y(n567) );
  MUX41X1_HVT U63 ( .A1(n567), .A3(n365), .A2(n392), .A4(n372), .S0(n355), 
        .S1(n263), .Y(n566) );
  AO21X1_HVT U66 ( .A1(n370), .A2(n321), .A3(n391), .Y(n563) );
  MUX41X1_HVT U68 ( .A1(n368), .A3(n563), .A2(n562), .A4(n564), .S0(n314), 
        .S1(n291), .Y(n561) );
  NAND2X0_HVT U73 ( .A1(n335), .A2(n556), .Y(n557) );
  MUX41X1_HVT U75 ( .A1(n395), .A3(n400), .A2(n249), .A4(n285), .S0(n314), 
        .S1(n291), .Y(n554) );
  MUX41X1_HVT U78 ( .A1(n552), .A3(n555), .A2(n554), .A4(n559), .S0(in[0]), 
        .S1(n263), .Y(n551) );
  AND3X1_HVT U80 ( .A1(n340), .A2(n573), .A3(n548), .Y(n549) );
  MUX41X1_HVT U82 ( .A1(n586), .A3(n377), .A2(n359), .A4(n615), .S0(n314), 
        .S1(n264), .Y(n546) );
  AND2X1_HVT U83 ( .A1(n347), .A2(n38), .Y(n545) );
  MUX41X1_HVT U84 ( .A1(n378), .A3(n218), .A2(n613), .A4(n545), .S0(n314), 
        .S1(n353), .Y(n544) );
  NAND2X0_HVT U85 ( .A1(n350), .A2(n410), .Y(n543) );
  MUX41X1_HVT U86 ( .A1(n400), .A3(n543), .A2(n310), .A4(n306), .S0(n314), 
        .S1(n291), .Y(n542) );
  MUX41X1_HVT U87 ( .A1(n542), .A3(n546), .A2(n544), .A4(n547), .S0(in[0]), 
        .S1(n319), .Y(n541) );
  MUX41X1_HVT U90 ( .A1(n585), .A3(n589), .A2(n397), .A4(n540), .S0(n316), 
        .S1(n353), .Y(n539) );
  AO21X1_HVT U93 ( .A1(n324), .A2(n535), .A3(n396), .Y(n536) );
  MUX41X1_HVT U97 ( .A1(n395), .A3(n308), .A2(n346), .A4(n614), .S0(n314), 
        .S1(n353), .Y(n531) );
  NAND2X0_HVT U101 ( .A1(n526), .A2(n525), .Y(n527) );
  MUX41X1_HVT U103 ( .A1(n269), .A3(n369), .A2(n258), .A4(n595), .S0(n314), 
        .S1(n353), .Y(n523) );
  MUX41X1_HVT U105 ( .A1(n380), .A3(n583), .A2(n522), .A4(n394), .S0(n314), 
        .S1(n353), .Y(n521) );
  NAND2X0_HVT U110 ( .A1(n340), .A2(n517), .Y(n518) );
  AND2X1_HVT U115 ( .A1(n255), .A2(n326), .Y(n513) );
  NAND2X0_HVT U123 ( .A1(n504), .A2(n503), .Y(n505) );
  MUX41X1_HVT U125 ( .A1(n608), .A3(n313), .A2(n368), .A4(n234), .S0(n318), 
        .S1(n354), .Y(n501) );
  MUX41X1_HVT U131 ( .A1(n496), .A3(n498), .A2(n497), .A4(n499), .S0(n321), 
        .S1(n355), .Y(n495) );
  MUX41X1_HVT U132 ( .A1(n495), .A3(n508), .A2(n500), .A4(n514), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  MUX41X1_HVT U135 ( .A1(n404), .A3(n219), .A2(n624), .A4(n603), .S0(n315), 
        .S1(n355), .Y(n492) );
  MUX41X1_HVT U136 ( .A1(n306), .A3(n597), .A2(n405), .A4(n594), .S0(n317), 
        .S1(n355), .Y(n491) );
  MUX41X1_HVT U139 ( .A1(n489), .A3(n492), .A2(n491), .A4(n493), .S0(in[0]), 
        .S1(n319), .Y(n488) );
  AND2X1_HVT U140 ( .A1(n334), .A2(n349), .Y(n487) );
  MUX41X1_HVT U141 ( .A1(n605), .A3(n273), .A2(n487), .A4(n384), .S0(n315), 
        .S1(n354), .Y(n486) );
  MUX41X1_HVT U142 ( .A1(n378), .A3(n326), .A2(n393), .A4(n334), .S0(n315), 
        .S1(n354), .Y(n485) );
  NAND2X0_HVT U146 ( .A1(n347), .A2(n343), .Y(n556) );
  MUX41X1_HVT U147 ( .A1(n405), .A3(n556), .A2(n395), .A4(n585), .S0(n315), 
        .S1(n355), .Y(n481) );
  OA21X1_HVT U151 ( .A1(n591), .A2(n356), .A3(n477), .Y(n478) );
  AND2X1_HVT U154 ( .A1(n324), .A2(n333), .Y(n474) );
  NAND2X0_HVT U158 ( .A1(n347), .A2(n410), .Y(n470) );
  MUX41X1_HVT U159 ( .A1(n617), .A3(n326), .A2(n470), .A4(n367), .S0(n351), 
        .S1(n290), .Y(n469) );
  MUX41X1_HVT U160 ( .A1(n469), .A3(n475), .A2(n471), .A4(n476), .S0(in[0]), 
        .S1(n320), .Y(n468) );
  AND2X1_HVT U162 ( .A1(n218), .A2(n556), .Y(n466) );
  MUX41X1_HVT U163 ( .A1(n374), .A3(n466), .A2(n307), .A4(n467), .S0(n351), 
        .S1(n353), .Y(n465) );
  MUX41X1_HVT U165 ( .A1(n608), .A3(n381), .A2(n585), .A4(n464), .S0(n355), 
        .S1(n352), .Y(n463) );
  NAND2X0_HVT U166 ( .A1(n342), .A2(n573), .Y(n462) );
  NAND2X0_HVT U167 ( .A1(n249), .A2(n350), .Y(n461) );
  NAND2X0_HVT U174 ( .A1(n254), .A2(n623), .Y(n616) );
  MUX41X1_HVT U176 ( .A1(n331), .A3(n455), .A2(n403), .A4(n616), .S0(n355), 
        .S1(n352), .Y(n454) );
  NAND2X0_HVT U177 ( .A1(n345), .A2(n330), .Y(n453) );
  MUX41X1_HVT U178 ( .A1(n612), .A3(n453), .A2(n406), .A4(n593), .S0(n315), 
        .S1(n291), .Y(n452) );
  MUX41X1_HVT U179 ( .A1(n602), .A3(n407), .A2(n363), .A4(n406), .S0(n351), 
        .S1(n291), .Y(n451) );
  MUX41X1_HVT U180 ( .A1(n366), .A3(n621), .A2(n617), .A4(n305), .S0(n322), 
        .S1(n352), .Y(n450) );
  MUX41X1_HVT U181 ( .A1(n450), .A3(n452), .A2(n451), .A4(n454), .S0(in[0]), 
        .S1(n320), .Y(n449) );
  MUX41X1_HVT U182 ( .A1(n387), .A3(n337), .A2(n389), .A4(n379), .S0(n355), 
        .S1(n351), .Y(n448) );
  OA21X1_HVT U184 ( .A1(n596), .A2(n356), .A3(n378), .Y(n446) );
  MUX41X1_HVT U186 ( .A1(n308), .A3(n592), .A2(n556), .A4(n585), .S0(n352), 
        .S1(n353), .Y(n444) );
  MUX41X1_HVT U189 ( .A1(n442), .A3(n616), .A2(n443), .A4(n394), .S0(n322), 
        .S1(n351), .Y(n441) );
  MUX41X1_HVT U190 ( .A1(n441), .A3(n444), .A2(n445), .A4(n448), .S0(n320), 
        .S1(in[0]), .Y(n440) );
  MUX41X1_HVT U193 ( .A1(n589), .A3(n595), .A2(n581), .A4(n439), .S0(n352), 
        .S1(n290), .Y(n438) );
  MUX41X1_HVT U194 ( .A1(n590), .A3(n603), .A2(n404), .A4(n334), .S0(n322), 
        .S1(n352), .Y(n437) );
  AO21X1_HVT U197 ( .A1(n310), .A2(n323), .A3(n396), .Y(n434) );
  MUX41X1_HVT U203 ( .A1(n594), .A3(n388), .A2(n618), .A4(n598), .S0(n352), 
        .S1(n290), .Y(n428) );
  MUX41X1_HVT U204 ( .A1(n574), .A3(n617), .A2(n385), .A4(n607), .S0(n351), 
        .S1(n290), .Y(n427) );
  MUX41X1_HVT U205 ( .A1(n38), .A3(n268), .A2(n407), .A4(n383), .S0(n352), 
        .S1(n290), .Y(n426) );
  NAND2X0_HVT U208 ( .A1(n347), .A2(n338), .Y(n517) );
  NAND2X0_HVT U212 ( .A1(n347), .A2(n335), .Y(n573) );
  NAND2X0_HVT U214 ( .A1(n218), .A2(n350), .Y(n424) );
  NAND2X0_HVT U215 ( .A1(n517), .A2(n336), .Y(n423) );
  AO21X1_HVT U216 ( .A1(n349), .A2(n219), .A3(n356), .Y(n526) );
  NAND2X0_HVT U218 ( .A1(n408), .A2(n254), .Y(n477) );
  NAND2X0_HVT U220 ( .A1(n323), .A2(n424), .Y(n548) );
  IBUFFX2_HVT U1 ( .A(n356), .Y(n290) );
  IBUFFX2_HVT U2 ( .A(n356), .Y(n291) );
  MUX21X2_HVT U6 ( .A1(n468), .A2(n456), .S0(n23), .Y(out[5]) );
  IBUFFX16_HVT U7 ( .A(in[6]), .Y(n23) );
  INVX4_HVT U8 ( .A(in[7]), .Y(n356) );
  NBUFFX2_HVT U9 ( .A(in[4]), .Y(n38) );
  NAND2X1_HVT U10 ( .A1(n616), .A2(n342), .Y(n617) );
  MUX21X1_HVT U11 ( .A1(n409), .A2(n249), .S0(n255), .Y(n591) );
  INVX1_HVT U12 ( .A(n628), .Y(n249) );
  NAND2X0_HVT U13 ( .A1(n278), .A2(n114), .Y(n117) );
  NAND2X0_HVT U14 ( .A1(n327), .A2(n213), .Y(n210) );
  NAND2X0_HVT U16 ( .A1(n117), .A2(n210), .Y(n533) );
  INVX8_HVT U17 ( .A(n213), .Y(n114) );
  NBUFFX2_HVT U18 ( .A(n411), .Y(n327) );
  IBUFFX2_HVT U19 ( .A(n344), .Y(n213) );
  MUX21X2_HVT U20 ( .A1(n251), .A2(n336), .S0(n323), .Y(n494) );
  IBUFFX2_HVT U22 ( .A(n590), .Y(n389) );
  MUX21X1_HVT U23 ( .A1(n387), .A2(n607), .S0(n211), .Y(n490) );
  IBUFFX16_HVT U25 ( .A(n323), .Y(n211) );
  MUX21X2_HVT U26 ( .A1(n509), .A2(n512), .S0(n212), .Y(n508) );
  IBUFFX16_HVT U27 ( .A(n252), .Y(n212) );
  IBUFFX2_HVT U28 ( .A(n607), .Y(n378) );
  IBUFFX2_HVT U29 ( .A(n285), .Y(n605) );
  MUX21X2_HVT U30 ( .A1(n340), .A2(n327), .S0(n345), .Y(n590) );
  INVX0_HVT U31 ( .A(n411), .Y(n216) );
  MUX21X1_HVT U32 ( .A1(n510), .A2(n511), .S0(n323), .Y(n509) );
  MUX21X2_HVT U34 ( .A1(n339), .A2(n292), .S0(n286), .Y(n285) );
  XNOR2X2_HVT U36 ( .A1(n329), .A2(n217), .Y(n623) );
  IBUFFX16_HVT U37 ( .A(n332), .Y(n217) );
  MUX21X2_HVT U38 ( .A1(n307), .A2(n373), .S0(n236), .Y(n497) );
  MUX21X1_HVT U39 ( .A1(n549), .A2(n550), .S0(n276), .Y(n547) );
  MUX21X1_HVT U40 ( .A1(n570), .A2(n572), .S0(n316), .Y(n569) );
  IBUFFX2_HVT U41 ( .A(in[0]), .Y(n231) );
  INVX0_HVT U43 ( .A(n292), .Y(n218) );
  INVX0_HVT U44 ( .A(n292), .Y(n293) );
  IBUFFX2_HVT U45 ( .A(n351), .Y(n233) );
  INVX0_HVT U46 ( .A(n336), .Y(n219) );
  NBUFFX2_HVT U47 ( .A(n620), .Y(n336) );
  MUX21X1_HVT U48 ( .A1(n612), .A2(n384), .S0(n315), .Y(n496) );
  MUX21X1_HVT U49 ( .A1(n566), .A2(n568), .S0(n316), .Y(n565) );
  MUX41X1_HVT U50 ( .A1(n575), .A3(n565), .A2(n569), .A4(n561), .S0(n226), 
        .S1(n231), .Y(out[0]) );
  IBUFFX16_HVT U52 ( .A(in[6]), .Y(n226) );
  MUX21X1_HVT U54 ( .A1(n331), .A2(n293), .S0(n232), .Y(n553) );
  IBUFFX16_HVT U55 ( .A(n347), .Y(n232) );
  MUX41X1_HVT U57 ( .A1(n553), .A3(n401), .A2(n621), .A4(n402), .S0(n322), 
        .S1(n233), .Y(n552) );
  NBUFFX2_HVT U60 ( .A(n251), .Y(n234) );
  MUX21X2_HVT U64 ( .A1(n382), .A2(n494), .S0(n235), .Y(n493) );
  IBUFFX16_HVT U65 ( .A(n256), .Y(n235) );
  MUX21X2_HVT U67 ( .A1(n259), .A2(n337), .S0(n253), .Y(n251) );
  IBUFFX16_HVT U69 ( .A(n239), .Y(n236) );
  MUX41X1_HVT U70 ( .A1(n486), .A3(n482), .A2(n485), .A4(n481), .S0(n237), 
        .S1(n238), .Y(n480) );
  IBUFFX16_HVT U71 ( .A(in[0]), .Y(n237) );
  IBUFFX16_HVT U72 ( .A(n319), .Y(n238) );
  IBUFFX16_HVT U74 ( .A(n318), .Y(n239) );
  INVX1_HVT U76 ( .A(n613), .Y(n373) );
  MUX21X2_HVT U77 ( .A1(n502), .A2(n501), .S0(n240), .Y(n500) );
  IBUFFX16_HVT U79 ( .A(n321), .Y(n240) );
  NBUFFX2_HVT U81 ( .A(n412), .Y(n331) );
  NBUFFX2_HVT U88 ( .A(n412), .Y(n329) );
  INVX0_HVT U89 ( .A(in[7]), .Y(n357) );
  INVX1_HVT U91 ( .A(n276), .Y(n352) );
  INVX0_HVT U92 ( .A(n346), .Y(n242) );
  INVX0_HVT U94 ( .A(n280), .Y(n436) );
  INVX0_HVT U95 ( .A(n342), .Y(n281) );
  INVX1_HVT U96 ( .A(n357), .Y(n354) );
  MUX21X1_HVT U98 ( .A1(n328), .A2(n410), .S0(n347), .Y(n622) );
  INVX0_HVT U99 ( .A(n241), .Y(n464) );
  OA21X1_HVT U100 ( .A1(n622), .A2(n356), .A3(n273), .Y(n430) );
  INVX0_HVT U102 ( .A(n258), .Y(n601) );
  MUX21X1_HVT U104 ( .A1(n292), .A2(n278), .S0(n279), .Y(n277) );
  INVX0_HVT U106 ( .A(n267), .Y(n269) );
  MUX21X1_HVT U107 ( .A1(n341), .A2(n538), .S0(n312), .Y(n537) );
  MUX41X1_HVT U108 ( .A1(n359), .A3(n308), .A2(n399), .A4(n533), .S0(n314), 
        .S1(n290), .Y(n532) );
  NBUFFX2_HVT U109 ( .A(n411), .Y(n328) );
  INVX0_HVT U111 ( .A(n518), .Y(n284) );
  INVX0_HVT U112 ( .A(n346), .Y(n253) );
  XNOR2X1_HVT U113 ( .A1(n603), .A2(in[7]), .Y(n587) );
  AO21X1_HVT U114 ( .A1(n318), .A2(n334), .A3(n218), .Y(n510) );
  INVX1_HVT U116 ( .A(n332), .Y(n409) );
  INVX1_HVT U117 ( .A(n319), .Y(n272) );
  INVX1_HVT U118 ( .A(n320), .Y(n252) );
  INVX1_HVT U119 ( .A(n272), .Y(n263) );
  INVX1_HVT U120 ( .A(n625), .Y(n278) );
  NBUFFX2_HVT U121 ( .A(n354), .Y(n324) );
  INVX1_HVT U122 ( .A(in[7]), .Y(n282) );
  NBUFFX2_HVT U124 ( .A(n354), .Y(n322) );
  INVX1_HVT U126 ( .A(n318), .Y(n256) );
  INVX1_HVT U127 ( .A(n318), .Y(n276) );
  INVX1_HVT U128 ( .A(in[0]), .Y(n271) );
  INVX1_HVT U129 ( .A(n254), .Y(n250) );
  INVX0_HVT U130 ( .A(n349), .Y(n344) );
  INVX0_HVT U133 ( .A(n349), .Y(n348) );
  INVX1_HVT U134 ( .A(n331), .Y(n259) );
  INVX0_HVT U137 ( .A(in[6]), .Y(n300) );
  INVX1_HVT U138 ( .A(n282), .Y(n264) );
  MUX21X1_HVT U143 ( .A1(n334), .A2(n339), .S0(n348), .Y(n241) );
  INVX1_HVT U144 ( .A(n334), .Y(n408) );
  MUX21X2_HVT U145 ( .A1(n435), .A2(n434), .S0(n316), .Y(n433) );
  MUX21X1_HVT U148 ( .A1(n390), .A2(n406), .S0(n323), .Y(n435) );
  MUX21X2_HVT U149 ( .A1(n472), .A2(n473), .S0(n318), .Y(n471) );
  MUX21X1_HVT U150 ( .A1(n38), .A2(n278), .S0(n242), .Y(n598) );
  MUX41X1_HVT U152 ( .A1(n534), .A3(n539), .A2(n531), .A4(n532), .S0(n257), 
        .S1(n271), .Y(n530) );
  INVX1_HVT U153 ( .A(n272), .Y(n257) );
  NAND2X0_HVT U155 ( .A1(n541), .A2(n300), .Y(n243) );
  NAND2X0_HVT U156 ( .A1(n551), .A2(in[6]), .Y(n244) );
  NAND2X0_HVT U157 ( .A1(n243), .A2(n244), .Y(out[1]) );
  INVX0_HVT U161 ( .A(n609), .Y(n377) );
  INVX1_HVT U164 ( .A(n596), .Y(n385) );
  NAND2X0_HVT U168 ( .A1(n430), .A2(n256), .Y(n245) );
  NAND2X0_HVT U169 ( .A1(n431), .A2(n316), .Y(n246) );
  NAND2X0_HVT U170 ( .A1(n245), .A2(n246), .Y(n429) );
  NAND2X0_HVT U171 ( .A1(n333), .A2(n344), .Y(n247) );
  NAND2X0_HVT U172 ( .A1(n328), .A2(n250), .Y(n248) );
  NAND2X0_HVT U173 ( .A1(n247), .A2(n248), .Y(n607) );
  INVX1_HVT U175 ( .A(n622), .Y(n368) );
  INVX0_HVT U183 ( .A(n623), .Y(n292) );
  INVX1_HVT U185 ( .A(n623), .Y(n411) );
  MUX41X1_HVT U187 ( .A1(n619), .A3(n574), .A2(n610), .A4(n398), .S0(n357), 
        .S1(n252), .Y(n572) );
  INVX0_HVT U188 ( .A(n349), .Y(n254) );
  IBUFFX2_HVT U191 ( .A(n349), .Y(n255) );
  IBUFFX2_HVT U192 ( .A(n349), .Y(n345) );
  MUX21X2_HVT U195 ( .A1(n626), .A2(n490), .S0(n256), .Y(n489) );
  MUX21X2_HVT U196 ( .A1(n478), .A2(n479), .S0(n318), .Y(n476) );
  MUX21X2_HVT U198 ( .A1(n536), .A2(n537), .S0(n318), .Y(n534) );
  MUX21X1_HVT U199 ( .A1(n259), .A2(n337), .S0(n254), .Y(n258) );
  INVX1_HVT U200 ( .A(n417), .Y(n382) );
  NAND2X0_HVT U201 ( .A1(n474), .A2(n260), .Y(n261) );
  NAND2X0_HVT U202 ( .A1(n341), .A2(n312), .Y(n262) );
  NAND2X0_HVT U206 ( .A1(n261), .A2(n262), .Y(n473) );
  IBUFFX2_HVT U207 ( .A(n312), .Y(n260) );
  XOR2X1_HVT U209 ( .A1(n276), .A2(n357), .Y(n584) );
  MUX41X1_HVT U210 ( .A1(n521), .A3(n524), .A2(n523), .A4(n528), .S0(in[0]), 
        .S1(n263), .Y(n520) );
  IBUFFX2_HVT U211 ( .A(n357), .Y(n355) );
  MUX21X1_HVT U213 ( .A1(n593), .A2(n402), .S0(n322), .Y(n472) );
  INVX0_HVT U217 ( .A(n273), .Y(n593) );
  NAND2X0_HVT U219 ( .A1(n336), .A2(n264), .Y(n265) );
  NAND2X0_HVT U221 ( .A1(n609), .A2(n282), .Y(n266) );
  NAND2X0_HVT U222 ( .A1(n265), .A2(n266), .Y(n550) );
  INVX1_HVT U223 ( .A(n627), .Y(n267) );
  INVX0_HVT U224 ( .A(n267), .Y(n268) );
  INVX0_HVT U225 ( .A(n267), .Y(n270) );
  MUX21X1_HVT U226 ( .A1(n343), .A2(n337), .S0(n348), .Y(n273) );
  MUX21X2_HVT U227 ( .A1(n432), .A2(n425), .S0(n300), .Y(out[7]) );
  NAND2X0_HVT U228 ( .A1(n282), .A2(n613), .Y(n274) );
  NAND2X0_HVT U229 ( .A1(n305), .A2(n322), .Y(n275) );
  NAND2X0_HVT U230 ( .A1(n274), .A2(n275), .Y(n431) );
  MUX21X2_HVT U231 ( .A1(n560), .A2(n587), .S0(n276), .Y(n559) );
  MUX21X2_HVT U232 ( .A1(n601), .A2(n364), .S0(n324), .Y(n484) );
  INVX0_HVT U233 ( .A(n346), .Y(n279) );
  MUX21X2_HVT U234 ( .A1(n484), .A2(n483), .S0(n317), .Y(n482) );
  MUX41X1_HVT U235 ( .A1(n277), .A3(n281), .A2(n420), .A4(n326), .S0(n276), 
        .S1(n282), .Y(n280) );
  OAI21X2_HVT U236 ( .A1(n277), .A2(n256), .A3(n375), .Y(n304) );
  INVX1_HVT U237 ( .A(n301), .Y(n514) );
  INVX1_HVT U238 ( .A(n349), .Y(n346) );
  MUX21X1_HVT U239 ( .A1(n410), .A2(n399), .S0(n324), .Y(n560) );
  INVX2_HVT U240 ( .A(n256), .Y(n351) );
  INVX0_HVT U241 ( .A(n348), .Y(n289) );
  INVX0_HVT U242 ( .A(n345), .Y(n286) );
  MUX21X2_HVT U243 ( .A1(n506), .A2(n505), .S0(n324), .Y(n502) );
  OA21X1_HVT U244 ( .A1(n362), .A2(n356), .A3(n599), .Y(n483) );
  OA21X1_HVT U245 ( .A1(n311), .A2(n356), .A3(n599), .Y(n458) );
  INVX0_HVT U246 ( .A(n599), .Y(n383) );
  INVX1_HVT U247 ( .A(n420), .Y(n399) );
  MUX21X1_HVT U248 ( .A1(n284), .A2(n383), .S0(n276), .Y(n283) );
  MUX21X1_HVT U249 ( .A1(n342), .A2(n335), .S0(n344), .Y(n599) );
  MUX41X1_HVT U250 ( .A1(n599), .A3(n285), .A2(n513), .A4(n617), .S0(n276), 
        .S1(n357), .Y(n512) );
  IBUFFX2_HVT U251 ( .A(in[1]), .Y(n350) );
  MUX21X2_HVT U252 ( .A1(n360), .A2(n507), .S0(n315), .Y(n506) );
  NAND2X0_HVT U253 ( .A1(n410), .A2(n348), .Y(n287) );
  NAND2X0_HVT U254 ( .A1(n249), .A2(n289), .Y(n288) );
  NAND2X0_HVT U255 ( .A1(n287), .A2(n288), .Y(n603) );
  INVX2_HVT U256 ( .A(in[1]), .Y(n349) );
  MUX21X2_HVT U257 ( .A1(n440), .A2(n449), .S0(in[6]), .Y(out[6]) );
  MUX41X1_HVT U258 ( .A1(n460), .A3(n457), .A2(n465), .A4(n463), .S0(n272), 
        .S1(in[0]), .Y(n456) );
  MUX41X1_HVT U259 ( .A1(n518), .A3(n339), .A2(n309), .A4(n361), .S0(n291), 
        .S1(n316), .Y(n475) );
  IBUFFX2_HVT U260 ( .A(n356), .Y(n353) );
  INVX0_HVT U261 ( .A(n519), .Y(n303) );
  INVX1_HVT U262 ( .A(n515), .Y(n302) );
  NAND2X0_HVT U263 ( .A1(n298), .A2(n299), .Y(out[2]) );
  MUX21X1_HVT U264 ( .A1(n409), .A2(n327), .S0(n349), .Y(n613) );
  MUX41X1_HVT U265 ( .A1(n398), .A3(n334), .A2(n461), .A4(n462), .S0(in[2]), 
        .S1(n291), .Y(n460) );
  MUX41X1_HVT U266 ( .A1(n429), .A3(n427), .A2(n428), .A4(n426), .S0(n271), 
        .S1(n252), .Y(n425) );
  AND3X2_HVT U267 ( .A1(n317), .A2(n350), .A3(n38), .Y(n498) );
  IBUFFX2_HVT U268 ( .A(n349), .Y(n347) );
  MUX41X1_HVT U269 ( .A1(n606), .A3(n557), .A2(n604), .A4(n558), .S0(n256), 
        .S1(n356), .Y(n555) );
  MUX21X2_HVT U270 ( .A1(n576), .A2(n580), .S0(n317), .Y(n575) );
  MUX21X2_HVT U271 ( .A1(n480), .A2(n488), .S0(in[6]), .Y(out[4]) );
  NAND2X0_HVT U272 ( .A1(n309), .A2(n294), .Y(n295) );
  NAND2X0_HVT U273 ( .A1(n529), .A2(n584), .Y(n296) );
  NAND2X0_HVT U274 ( .A1(n295), .A2(n296), .Y(n528) );
  INVX0_HVT U275 ( .A(n584), .Y(n294) );
  NAND2X0_HVT U276 ( .A1(n530), .A2(n297), .Y(n298) );
  NAND2X0_HVT U277 ( .A1(n520), .A2(n300), .Y(n299) );
  INVX1_HVT U278 ( .A(n300), .Y(n297) );
  MUX21X1_HVT U279 ( .A1(n383), .A2(n615), .S0(n318), .Y(n529) );
  MUX41X1_HVT U280 ( .A1(n437), .A3(n438), .A2(n433), .A4(n436), .S0(n257), 
        .S1(n271), .Y(n432) );
  XOR2X1_HVT U281 ( .A1(n350), .A2(n276), .Y(n582) );
  MUX41X1_HVT U282 ( .A1(n304), .A3(n283), .A2(n303), .A4(n302), .S0(n252), 
        .S1(n356), .Y(n301) );
  MUX21X2_HVT U283 ( .A1(n516), .A2(n341), .S0(n582), .Y(n515) );
  NBUFFX2_HVT U284 ( .A(n411), .Y(n326) );
  AND2X1_HVT U285 ( .A1(n328), .A2(n573), .Y(n305) );
  NBUFFX2_HVT U286 ( .A(n625), .Y(n337) );
  MUX21X1_HVT U287 ( .A1(n278), .A2(n410), .S0(n321), .Y(n577) );
  NBUFFX2_HVT U288 ( .A(n625), .Y(n338) );
  MUX21X1_HVT U289 ( .A1(n369), .A2(n219), .S0(n321), .Y(n562) );
  AND2X1_HVT U290 ( .A1(n340), .A2(n556), .Y(n306) );
  MUX21X1_HVT U291 ( .A1(n292), .A2(n330), .S0(n254), .Y(n525) );
  MUX21X1_HVT U292 ( .A1(n278), .A2(n249), .S0(n346), .Y(n455) );
  MUX21X1_HVT U293 ( .A1(n410), .A2(n327), .S0(n347), .Y(n467) );
  MUX21X1_HVT U294 ( .A1(n293), .A2(n408), .S0(n348), .Y(n416) );
  MUX21X1_HVT U295 ( .A1(n338), .A2(n336), .S0(n347), .Y(n540) );
  XOR2X1_HVT U296 ( .A1(n623), .A2(n347), .Y(n585) );
  MUX21X1_HVT U297 ( .A1(n325), .A2(n216), .S0(n254), .Y(n418) );
  MUX21X1_HVT U298 ( .A1(n410), .A2(n409), .S0(n346), .Y(n596) );
  MUX21X1_HVT U299 ( .A1(n361), .A2(n385), .S0(n316), .Y(n511) );
  NAND2X0_HVT U300 ( .A1(n329), .A2(n325), .Y(n625) );
  NBUFFX2_HVT U301 ( .A(n628), .Y(n339) );
  INVX1_HVT U302 ( .A(n629), .Y(n410) );
  MUX21X1_HVT U303 ( .A1(n341), .A2(n335), .S0(n344), .Y(n615) );
  MUX21X1_HVT U304 ( .A1(n337), .A2(n343), .S0(n346), .Y(n535) );
  MUX21X1_HVT U305 ( .A1(n330), .A2(n409), .S0(n344), .Y(n507) );
  NBUFFX2_HVT U306 ( .A(n628), .Y(n340) );
  NBUFFX2_HVT U307 ( .A(n628), .Y(n341) );
  XOR2X1_HVT U308 ( .A1(n344), .A2(n408), .Y(n586) );
  MUX21X1_HVT U309 ( .A1(n408), .A2(n278), .S0(n348), .Y(n611) );
  MUX21X1_HVT U310 ( .A1(n409), .A2(n410), .S0(n255), .Y(n619) );
  MUX21X1_HVT U311 ( .A1(n338), .A2(n409), .S0(n255), .Y(n618) );
  MUX21X1_HVT U312 ( .A1(n325), .A2(n331), .S0(n255), .Y(n439) );
  XOR2X1_HVT U313 ( .A1(n339), .A2(n254), .Y(n581) );
  MUX21X1_HVT U314 ( .A1(n325), .A2(n343), .S0(n346), .Y(n442) );
  MUX21X1_HVT U315 ( .A1(n342), .A2(n340), .S0(n348), .Y(n443) );
  MUX21X1_HVT U316 ( .A1(n339), .A2(n330), .S0(n345), .Y(n422) );
  XNOR2X1_HVT U317 ( .A1(n337), .A2(n346), .Y(n307) );
  AND2X1_HVT U318 ( .A1(n344), .A2(n249), .Y(n308) );
  MUX21X1_HVT U319 ( .A1(n339), .A2(n338), .S0(n345), .Y(n415) );
  AND2X1_HVT U320 ( .A1(n342), .A2(n517), .Y(n309) );
  XNOR2X1_HVT U321 ( .A1(n343), .A2(n254), .Y(n310) );
  MUX21X1_HVT U322 ( .A1(n335), .A2(n409), .S0(n345), .Y(n420) );
  MUX21X1_HVT U323 ( .A1(n336), .A2(n330), .S0(n348), .Y(n558) );
  MUX21X1_HVT U324 ( .A1(n336), .A2(n343), .S0(n317), .Y(n504) );
  XOR2X1_HVT U325 ( .A1(n331), .A2(n345), .Y(n604) );
  NBUFFX2_HVT U326 ( .A(n409), .Y(n325) );
  NBUFFX2_HVT U327 ( .A(n354), .Y(n323) );
  NBUFFX2_HVT U328 ( .A(in[5]), .Y(n321) );
  NBUFFX2_HVT U329 ( .A(in[2]), .Y(n315) );
  NBUFFX2_HVT U330 ( .A(in[5]), .Y(n320) );
  NBUFFX2_HVT U331 ( .A(in[2]), .Y(n317) );
  NBUFFX2_HVT U332 ( .A(in[2]), .Y(n318) );
  NBUFFX2_HVT U333 ( .A(in[2]), .Y(n316) );
  NBUFFX2_HVT U334 ( .A(n351), .Y(n314) );
  NBUFFX2_HVT U335 ( .A(in[5]), .Y(n319) );
  MUX21X1_HVT U336 ( .A1(n527), .A2(n382), .S0(n317), .Y(n524) );
  MUX21X1_HVT U337 ( .A1(n446), .A2(n447), .S0(n316), .Y(n445) );
  MUX21X1_HVT U338 ( .A1(n543), .A2(n333), .S0(n323), .Y(n447) );
  XOR2X1_HVT U339 ( .A1(n255), .A2(n332), .Y(n583) );
  MUX21X1_HVT U340 ( .A1(n335), .A2(n328), .S0(n255), .Y(n522) );
  MUX21X1_HVT U341 ( .A1(n401), .A2(n219), .S0(n323), .Y(n479) );
  MUX21X1_HVT U342 ( .A1(n459), .A2(n458), .S0(n317), .Y(n457) );
  MUX21X1_HVT U343 ( .A1(n336), .A2(n399), .S0(n324), .Y(n459) );
  AND2X1_HVT U344 ( .A1(n328), .A2(n350), .Y(n311) );
  MUX21X1_HVT U345 ( .A1(n333), .A2(n278), .S0(n255), .Y(n592) );
  NAND2X0_HVT U346 ( .A1(n332), .A2(n329), .Y(n628) );
  NBUFFX2_HVT U347 ( .A(n620), .Y(n334) );
  MUX21X1_HVT U348 ( .A1(n249), .A2(n333), .S0(n348), .Y(n610) );
  MUX21X1_HVT U349 ( .A1(n386), .A2(n269), .S0(n315), .Y(n519) );
  MUX21X1_HVT U350 ( .A1(n578), .A2(n579), .S0(n322), .Y(n576) );
  MUX21X1_HVT U351 ( .A1(n333), .A2(n595), .S0(n321), .Y(n579) );
  XOR2X1_HVT U352 ( .A1(n254), .A2(n320), .Y(n588) );
  MUX21X1_HVT U353 ( .A1(n269), .A2(n349), .S0(n316), .Y(n503) );
  MUX21X1_HVT U354 ( .A1(n333), .A2(n219), .S0(n345), .Y(n419) );
  MUX21X1_HVT U355 ( .A1(n600), .A2(n423), .S0(n322), .Y(n417) );
  MUX21X1_HVT U356 ( .A1(n338), .A2(n333), .S0(n344), .Y(n621) );
  MUX21X1_HVT U357 ( .A1(n371), .A2(n350), .S0(n321), .Y(n564) );
  MUX21X1_HVT U358 ( .A1(n333), .A2(n331), .S0(n324), .Y(n538) );
  NBUFFX2_HVT U359 ( .A(n620), .Y(n335) );
  MUX21X1_HVT U360 ( .A1(n380), .A2(n600), .S0(n315), .Y(n499) );
  NBUFFX2_HVT U361 ( .A(n629), .Y(n343) );
  NBUFFX2_HVT U362 ( .A(n412), .Y(n330) );
  NBUFFX2_HVT U363 ( .A(n629), .Y(n342) );
  XNOR2X1_HVT U364 ( .A1(n356), .A2(n255), .Y(n312) );
  AND2X1_HVT U365 ( .A1(n409), .A2(n350), .Y(n313) );
  INVX0_HVT U366 ( .A(in[4]), .Y(n412) );
  MUX21X1_HVT U367 ( .A1(n38), .A2(n293), .S0(n344), .Y(n421) );
  NAND2X0_HVT U368 ( .A1(in[4]), .A2(n325), .Y(n620) );
  NAND2X0_HVT U369 ( .A1(n332), .A2(in[4]), .Y(n629) );
  MUX21X1_HVT U370 ( .A1(n38), .A2(n410), .S0(n346), .Y(n594) );
  MUX21X1_HVT U371 ( .A1(n38), .A2(n408), .S0(n347), .Y(n612) );
  MUX21X1_HVT U372 ( .A1(n38), .A2(n341), .S0(n345), .Y(n609) );
  MUX21X1_HVT U373 ( .A1(n38), .A2(n335), .S0(n348), .Y(n414) );
  MUX21X1_HVT U374 ( .A1(n343), .A2(n38), .S0(n345), .Y(n602) );
  MUX21X1_HVT U375 ( .A1(n333), .A2(n38), .S0(n317), .Y(n516) );
  MUX21X1_HVT U376 ( .A1(n38), .A2(n342), .S0(n254), .Y(n413) );
  MUX21X1_HVT U377 ( .A1(n409), .A2(n38), .S0(n344), .Y(n600) );
  NBUFFX2_HVT U378 ( .A(in[3]), .Y(n332) );
  NBUFFX2_HVT U379 ( .A(in[3]), .Y(n333) );
  INVX0_HVT U380 ( .A(n608), .Y(n358) );
  INVX0_HVT U381 ( .A(n606), .Y(n359) );
  INVX0_HVT U382 ( .A(n597), .Y(n360) );
  INVX0_HVT U383 ( .A(n595), .Y(n361) );
  INVX0_HVT U384 ( .A(n461), .Y(n362) );
  INVX0_HVT U385 ( .A(n424), .Y(n363) );
  INVX0_HVT U386 ( .A(n270), .Y(n364) );
  INVX0_HVT U387 ( .A(n614), .Y(n365) );
  INVX0_HVT U388 ( .A(n626), .Y(n366) );
  INVX0_HVT U389 ( .A(n624), .Y(n367) );
  INVX0_HVT U390 ( .A(n621), .Y(n369) );
  INVX0_HVT U391 ( .A(n619), .Y(n370) );
  INVX0_HVT U392 ( .A(n618), .Y(n371) );
  INVX0_HVT U393 ( .A(n615), .Y(n372) );
  INVX0_HVT U394 ( .A(n612), .Y(n374) );
  INVX0_HVT U395 ( .A(n611), .Y(n375) );
  INVX0_HVT U396 ( .A(n610), .Y(n376) );
  INVX0_HVT U397 ( .A(n604), .Y(n379) );
  INVX0_HVT U398 ( .A(n602), .Y(n380) );
  INVX0_HVT U399 ( .A(n600), .Y(n381) );
  INVX0_HVT U400 ( .A(n598), .Y(n384) );
  INVX0_HVT U401 ( .A(n594), .Y(n386) );
  INVX0_HVT U402 ( .A(n592), .Y(n387) );
  INVX0_HVT U403 ( .A(n591), .Y(n388) );
  INVX0_HVT U404 ( .A(n589), .Y(n390) );
  INVX0_HVT U405 ( .A(n556), .Y(n391) );
  INVX0_HVT U406 ( .A(n617), .Y(n392) );
  INVX0_HVT U407 ( .A(n517), .Y(n393) );
  INVX0_HVT U408 ( .A(n423), .Y(n394) );
  INVX0_HVT U409 ( .A(n573), .Y(n395) );
  INVX0_HVT U410 ( .A(n477), .Y(n396) );
  INVX0_HVT U411 ( .A(n422), .Y(n397) );
  INVX0_HVT U412 ( .A(n421), .Y(n398) );
  INVX0_HVT U413 ( .A(n419), .Y(n400) );
  INVX0_HVT U414 ( .A(n418), .Y(n401) );
  INVX0_HVT U415 ( .A(n535), .Y(n402) );
  INVX0_HVT U416 ( .A(n525), .Y(n403) );
  INVX0_HVT U417 ( .A(n416), .Y(n404) );
  INVX0_HVT U418 ( .A(n415), .Y(n405) );
  INVX0_HVT U419 ( .A(n414), .Y(n406) );
  INVX0_HVT U420 ( .A(n413), .Y(n407) );
endmodule

