
module sbox_1 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n83, n121, n210, n211, n212, n213, n216, n217, n218, n219,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588;

  NAND2X0_HVT U3 ( .A1(n302), .A2(n295), .Y(n586) );
  NAND2X0_HVT U4 ( .A1(n293), .A2(n586), .Y(n585) );
  NAND2X0_HVT U5 ( .A1(n302), .A2(n283), .Y(n583) );
  NAND2X0_HVT U13 ( .A1(n575), .A2(n297), .Y(n576) );
  NAND2X0_HVT U15 ( .A1(n586), .A2(n285), .Y(n573) );
  NAND2X0_HVT U21 ( .A1(n293), .A2(n121), .Y(n567) );
  NAND2X0_HVT U24 ( .A1(n290), .A2(n121), .Y(n565) );
  NAND2X0_HVT U33 ( .A1(n364), .A2(n121), .Y(n556) );
  NAND2X0_HVT U35 ( .A1(n288), .A2(n121), .Y(n554) );
  NAND2X0_HVT U42 ( .A1(n302), .A2(n290), .Y(n547) );
  MUX41X1_HVT U51 ( .A1(n352), .A3(n312), .A2(n330), .A4(n331), .S0(n210), 
        .S1(n307), .Y(n539) );
  NAND2X0_HVT U53 ( .A1(n536), .A2(n546), .Y(n537) );
  NAND2X0_HVT U56 ( .A1(n293), .A2(n532), .Y(n533) );
  MUX41X1_HVT U57 ( .A1(n353), .A3(n569), .A2(n533), .A4(n578), .S0(n210), 
        .S1(n307), .Y(n531) );
  NAND2X0_HVT U58 ( .A1(n297), .A2(n586), .Y(n530) );
  MUX41X1_HVT U59 ( .A1(n270), .A3(n530), .A2(n268), .A4(n329), .S0(n210), 
        .S1(n307), .Y(n529) );
  MUX41X1_HVT U61 ( .A1(n267), .A3(n328), .A2(n327), .A4(n284), .S0(n210), 
        .S1(n307), .Y(n527) );
  NAND2X0_HVT U62 ( .A1(n121), .A2(n296), .Y(n526) );
  MUX41X1_HVT U63 ( .A1(n526), .A3(n319), .A2(n259), .A4(n326), .S0(n210), 
        .S1(n307), .Y(n525) );
  AO21X1_HVT U66 ( .A1(n324), .A2(n279), .A3(n347), .Y(n522) );
  MUX41X1_HVT U68 ( .A1(n322), .A3(n522), .A2(n521), .A4(n523), .S0(n271), 
        .S1(n252), .Y(n520) );
  MUX41X1_HVT U69 ( .A1(n520), .A3(n528), .A2(n524), .A4(n534), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n291), .A2(n515), .Y(n516) );
  MUX41X1_HVT U74 ( .A1(n517), .A3(n563), .A2(n516), .A4(n565), .S0(n273), 
        .S1(n23), .Y(n514) );
  MUX41X1_HVT U75 ( .A1(n350), .A3(n355), .A2(n368), .A4(n333), .S0(n271), 
        .S1(n308), .Y(n513) );
  MUX41X1_HVT U77 ( .A1(n580), .A3(n357), .A2(n512), .A4(n356), .S0(n280), 
        .S1(n304), .Y(n511) );
  MUX41X1_HVT U78 ( .A1(n511), .A3(n514), .A2(n513), .A4(n518), .S0(n289), 
        .S1(n277), .Y(n510) );
  MUX41X1_HVT U82 ( .A1(n544), .A3(n331), .A2(n313), .A4(n574), .S0(n271), 
        .S1(n252), .Y(n506) );
  AND2X1_HVT U83 ( .A1(n302), .A2(n253), .Y(n505) );
  MUX41X1_HVT U84 ( .A1(n332), .A3(n582), .A2(n572), .A4(n505), .S0(n271), 
        .S1(n309), .Y(n504) );
  NAND2X0_HVT U85 ( .A1(n121), .A2(n367), .Y(n503) );
  MUX41X1_HVT U86 ( .A1(n355), .A3(n503), .A2(n265), .A4(n263), .S0(n271), 
        .S1(n23), .Y(n502) );
  MUX41X1_HVT U87 ( .A1(n502), .A3(n506), .A2(n504), .A4(n507), .S0(in[0]), 
        .S1(n277), .Y(n501) );
  MUX41X1_HVT U90 ( .A1(n543), .A3(n547), .A2(n352), .A4(n500), .S0(n272), 
        .S1(n252), .Y(n499) );
  AO21X1_HVT U93 ( .A1(n282), .A2(n495), .A3(n351), .Y(n496) );
  MUX41X1_HVT U96 ( .A1(n313), .A3(n266), .A2(n354), .A4(n493), .S0(n271), 
        .S1(n252), .Y(n492) );
  MUX41X1_HVT U97 ( .A1(n350), .A3(n266), .A2(n302), .A4(n573), .S0(n271), 
        .S1(n309), .Y(n491) );
  MUX41X1_HVT U98 ( .A1(n491), .A3(n494), .A2(n492), .A4(n499), .S0(n289), 
        .S1(n277), .Y(n490) );
  NAND2X0_HVT U101 ( .A1(n486), .A2(n485), .Y(n487) );
  MUX41X1_HVT U103 ( .A1(n586), .A3(n323), .A2(n336), .A4(n244), .S0(n271), 
        .S1(n252), .Y(n483) );
  MUX41X1_HVT U105 ( .A1(n335), .A3(n542), .A2(n482), .A4(n349), .S0(n271), 
        .S1(n252), .Y(n481) );
  MUX41X1_HVT U106 ( .A1(n481), .A3(n484), .A2(n483), .A4(n488), .S0(in[0]), 
        .S1(n277), .Y(n480) );
  NAND2X0_HVT U110 ( .A1(n295), .A2(n476), .Y(n477) );
  MUX41X1_HVT U114 ( .A1(n473), .A3(n479), .A2(n475), .A4(n478), .S0(n279), 
        .S1(n23), .Y(n472) );
  AO21X1_HVT U118 ( .A1(n276), .A2(n292), .A3(n582), .Y(n469) );
  NAND2X0_HVT U123 ( .A1(n463), .A2(n462), .Y(n464) );
  MUX41X1_HVT U125 ( .A1(n567), .A3(n270), .A2(n322), .A4(n359), .S0(n272), 
        .S1(n210), .Y(n460) );
  AND3X1_HVT U128 ( .A1(n275), .A2(n121), .A3(n253), .Y(n457) );
  MUX41X1_HVT U131 ( .A1(n455), .A3(n457), .A2(n456), .A4(n458), .S0(n279), 
        .S1(n210), .Y(n454) );
  MUX41X1_HVT U136 ( .A1(n263), .A3(n556), .A2(n361), .A4(n553), .S0(n272), 
        .S1(n210), .Y(n450) );
  MUX41X1_HVT U139 ( .A1(n448), .A3(n451), .A2(n450), .A4(n452), .S0(n289), 
        .S1(n277), .Y(n447) );
  AND2X1_HVT U140 ( .A1(n292), .A2(n219), .Y(n446) );
  OA21X1_HVT U144 ( .A1(n316), .A2(n310), .A3(n558), .Y(n442) );
  NAND2X0_HVT U146 ( .A1(n302), .A2(n297), .Y(n515) );
  MUX41X1_HVT U148 ( .A1(n440), .A3(n444), .A2(n441), .A4(n445), .S0(in[0]), 
        .S1(n277), .Y(n439) );
  OA21X1_HVT U151 ( .A1(n549), .A2(n310), .A3(n436), .Y(n437) );
  MUX41X1_HVT U153 ( .A1(n477), .A3(n267), .A2(n294), .A4(n315), .S0(n272), 
        .S1(n309), .Y(n434) );
  AND2X1_HVT U154 ( .A1(n282), .A2(n290), .Y(n433) );
  NAND2X0_HVT U158 ( .A1(n302), .A2(n367), .Y(n429) );
  MUX41X1_HVT U159 ( .A1(n576), .A3(n284), .A2(n429), .A4(n321), .S0(in[2]), 
        .S1(n308), .Y(n428) );
  MUX41X1_HVT U160 ( .A1(n428), .A3(n434), .A2(n430), .A4(n435), .S0(n289), 
        .S1(n278), .Y(n427) );
  AND2X1_HVT U162 ( .A1(n582), .A2(n515), .Y(n425) );
  MUX41X1_HVT U163 ( .A1(n328), .A3(n425), .A2(n264), .A4(n426), .S0(in[2]), 
        .S1(n23), .Y(n424) );
  MUX41X1_HVT U165 ( .A1(n567), .A3(n337), .A2(n543), .A4(n423), .S0(n210), 
        .S1(n304), .Y(n422) );
  NAND2X0_HVT U166 ( .A1(n297), .A2(n532), .Y(n421) );
  NAND2X0_HVT U167 ( .A1(n368), .A2(n121), .Y(n420) );
  MUX41X1_HVT U168 ( .A1(n353), .A3(n291), .A2(n420), .A4(n421), .S0(in[2]), 
        .S1(n23), .Y(n419) );
  OA21X1_HVT U170 ( .A1(n268), .A2(n310), .A3(n558), .Y(n417) );
  NAND2X0_HVT U174 ( .A1(n302), .A2(n582), .Y(n575) );
  MUX41X1_HVT U176 ( .A1(n288), .A3(n414), .A2(n358), .A4(n575), .S0(n210), 
        .S1(in[2]), .Y(n413) );
  NAND2X0_HVT U177 ( .A1(n302), .A2(n287), .Y(n412) );
  MUX41X1_HVT U178 ( .A1(n571), .A3(n412), .A2(n362), .A4(n551), .S0(n273), 
        .S1(n308), .Y(n411) );
  MUX41X1_HVT U179 ( .A1(n561), .A3(n363), .A2(n317), .A4(n362), .S0(in[2]), 
        .S1(n309), .Y(n410) );
  MUX41X1_HVT U180 ( .A1(n320), .A3(n580), .A2(n576), .A4(n262), .S0(n280), 
        .S1(n304), .Y(n409) );
  MUX41X1_HVT U181 ( .A1(n409), .A3(n411), .A2(n410), .A4(n413), .S0(n289), 
        .S1(n278), .Y(n408) );
  MUX41X1_HVT U182 ( .A1(n343), .A3(n584), .A2(n345), .A4(n334), .S0(n210), 
        .S1(in[2]), .Y(n407) );
  OA21X1_HVT U184 ( .A1(n555), .A2(n310), .A3(n332), .Y(n405) );
  MUX41X1_HVT U186 ( .A1(n266), .A3(n550), .A2(n515), .A4(n543), .S0(n304), 
        .S1(n309), .Y(n403) );
  MUX41X1_HVT U189 ( .A1(n401), .A3(n575), .A2(n402), .A4(n349), .S0(n280), 
        .S1(in[2]), .Y(n400) );
  MUX41X1_HVT U190 ( .A1(n400), .A3(n403), .A2(n404), .A4(n407), .S0(n278), 
        .S1(in[0]), .Y(n399) );
  MUX41X1_HVT U194 ( .A1(n548), .A3(n562), .A2(n360), .A4(n292), .S0(n280), 
        .S1(n304), .Y(n396) );
  MUX41X1_HVT U195 ( .A1(n582), .A3(n354), .A2(n588), .A4(n552), .S0(in[2]), 
        .S1(n308), .Y(n395) );
  AO21X1_HVT U197 ( .A1(n265), .A2(n281), .A3(n351), .Y(n393) );
  OA21X1_HVT U201 ( .A1(n581), .A2(n310), .A3(n342), .Y(n389) );
  MUX41X1_HVT U204 ( .A1(n533), .A3(n576), .A2(n340), .A4(n566), .S0(n273), 
        .S1(n308), .Y(n386) );
  MUX41X1_HVT U205 ( .A1(n253), .A3(n586), .A2(n363), .A4(n260), .S0(n271), 
        .S1(n308), .Y(n385) );
  MUX41X1_HVT U206 ( .A1(n385), .A3(n387), .A2(n386), .A4(n388), .S0(n289), 
        .S1(n278), .Y(n384) );
  MUX21X2_HVT U207 ( .A1(n384), .A2(n391), .S0(in[6]), .Y(out[7]) );
  NAND2X0_HVT U208 ( .A1(n302), .A2(n293), .Y(n476) );
  NAND2X0_HVT U212 ( .A1(n302), .A2(n291), .Y(n532) );
  NAND2X0_HVT U214 ( .A1(n582), .A2(n121), .Y(n383) );
  NAND2X0_HVT U215 ( .A1(n476), .A2(n292), .Y(n382) );
  NAND2X0_HVT U218 ( .A1(n365), .A2(n302), .Y(n436) );
  NAND2X0_HVT U220 ( .A1(n281), .A2(n383), .Y(n508) );
  MUX21X2_HVT U1 ( .A1(n566), .A2(n343), .S0(n281), .Y(n449) );
  NBUFFX4_HVT U2 ( .A(n369), .Y(n286) );
  MUX21X2_HVT U6 ( .A1(n285), .A2(n283), .S0(n300), .Y(n572) );
  IBUFFX2_HVT U7 ( .A(in[3]), .Y(n366) );
  MUX21X2_HVT U8 ( .A1(n449), .A2(n585), .S0(n276), .Y(n448) );
  MUX21X2_HVT U9 ( .A1(n390), .A2(n389), .S0(n245), .Y(n388) );
  IBUFFX2_HVT U10 ( .A(n23), .Y(n83) );
  NBUFFX4_HVT U11 ( .A(n369), .Y(n285) );
  INVX1_HVT U12 ( .A(n306), .Y(n304) );
  INVX2_HVT U14 ( .A(n306), .Y(n305) );
  MUX21X2_HVT U16 ( .A1(n367), .A2(n286), .S0(n303), .Y(n581) );
  IBUFFX2_HVT U17 ( .A(n310), .Y(n23) );
  MUX41X1_HVT U18 ( .A1(n577), .A3(n557), .A2(n553), .A4(n344), .S0(n48), .S1(
        n83), .Y(n387) );
  IBUFFX16_HVT U19 ( .A(n245), .Y(n48) );
  NBUFFX2_HVT U20 ( .A(n303), .Y(n121) );
  INVX2_HVT U22 ( .A(in[1]), .Y(n303) );
  NBUFFX2_HVT U23 ( .A(in[7]), .Y(n210) );
  MUX41X1_HVT U25 ( .A1(n515), .A3(n361), .A2(n543), .A4(n350), .S0(n211), 
        .S1(n210), .Y(n440) );
  IBUFFX16_HVT U26 ( .A(n273), .Y(n211) );
  INVX1_HVT U27 ( .A(in[7]), .Y(n311) );
  INVX1_HVT U28 ( .A(n250), .Y(n212) );
  INVX1_HVT U29 ( .A(n250), .Y(n213) );
  INVX1_HVT U30 ( .A(n250), .Y(n300) );
  MUX41X1_HVT U31 ( .A1(n472), .A3(n459), .A2(n467), .A4(n454), .S0(n216), 
        .S1(n239), .Y(out[3]) );
  IBUFFX16_HVT U32 ( .A(in[6]), .Y(n216) );
  INVX1_HVT U34 ( .A(n249), .Y(n217) );
  INVX1_HVT U36 ( .A(n249), .Y(n218) );
  INVX0_HVT U37 ( .A(n249), .Y(n299) );
  INVX1_HVT U38 ( .A(in[1]), .Y(n250) );
  NBUFFX2_HVT U39 ( .A(n303), .Y(n219) );
  MUX41X1_HVT U40 ( .A1(n395), .A3(n397), .A2(n392), .A4(n396), .S0(in[0]), 
        .S1(n231), .Y(n391) );
  IBUFFX16_HVT U41 ( .A(n278), .Y(n231) );
  MUX21X2_HVT U43 ( .A1(n427), .A2(n415), .S0(n232), .Y(out[5]) );
  IBUFFX16_HVT U44 ( .A(in[6]), .Y(n232) );
  MUX21X2_HVT U45 ( .A1(n314), .A2(n466), .S0(n273), .Y(n465) );
  MUX21X2_HVT U46 ( .A1(n465), .A2(n464), .S0(n282), .Y(n461) );
  INVX1_HVT U47 ( .A(n315), .Y(n244) );
  NAND2X0_HVT U48 ( .A1(n535), .A2(n233), .Y(n234) );
  NAND2X0_HVT U49 ( .A1(n539), .A2(n275), .Y(n235) );
  NAND2X0_HVT U50 ( .A1(n234), .A2(n235), .Y(n534) );
  IBUFFX2_HVT U52 ( .A(n275), .Y(n233) );
  NAND2X0_HVT U54 ( .A1(n471), .A2(n236), .Y(n237) );
  NAND2X0_HVT U55 ( .A1(n468), .A2(n241), .Y(n238) );
  NAND2X0_HVT U60 ( .A1(n237), .A2(n238), .Y(n467) );
  IBUFFX2_HVT U64 ( .A(n241), .Y(n236) );
  IBUFFX16_HVT U65 ( .A(in[0]), .Y(n239) );
  MUX21X1_HVT U67 ( .A1(n469), .A2(n470), .S0(n281), .Y(n468) );
  INVX1_HVT U70 ( .A(n509), .Y(n247) );
  INVX0_HVT U71 ( .A(n248), .Y(n553) );
  INVX2_HVT U72 ( .A(n250), .Y(n301) );
  INVX1_HVT U76 ( .A(in[4]), .Y(n370) );
  NAND3X0_HVT U79 ( .A1(n295), .A2(n532), .A3(n508), .Y(n240) );
  NBUFFX2_HVT U80 ( .A(in[5]), .Y(n279) );
  INVX0_HVT U81 ( .A(n279), .Y(n241) );
  INVX0_HVT U88 ( .A(n305), .Y(n245) );
  INVX0_HVT U89 ( .A(n246), .Y(n507) );
  MUX21X2_HVT U91 ( .A1(n418), .A2(n417), .S0(n275), .Y(n416) );
  IBUFFX2_HVT U92 ( .A(n310), .Y(n308) );
  INVX2_HVT U94 ( .A(in[7]), .Y(n310) );
  NAND2X0_HVT U95 ( .A1(n290), .A2(n241), .Y(n242) );
  NAND2X0_HVT U99 ( .A1(n554), .A2(n279), .Y(n243) );
  NAND2X0_HVT U100 ( .A1(n242), .A2(n243), .Y(n538) );
  MUX21X1_HVT U102 ( .A1(n537), .A2(n538), .S0(n280), .Y(n535) );
  INVX1_HVT U104 ( .A(n554), .Y(n315) );
  MUX41X1_HVT U107 ( .A1(n562), .A3(n583), .A2(n365), .A4(n360), .S0(n245), 
        .S1(n311), .Y(n451) );
  INVX2_HVT U108 ( .A(n303), .Y(n302) );
  IBUFFX2_HVT U109 ( .A(n311), .Y(n254) );
  MUX21X2_HVT U111 ( .A1(n461), .A2(n460), .S0(n241), .Y(n459) );
  MUX21X1_HVT U112 ( .A1(n288), .A2(n283), .S0(n219), .Y(n398) );
  MUX41X1_HVT U113 ( .A1(n244), .A3(n547), .A2(n398), .A4(n540), .S0(n245), 
        .S1(n309), .Y(n397) );
  MUX21X1_HVT U115 ( .A1(n296), .A2(n253), .S0(n219), .Y(n568) );
  MUX21X1_HVT U116 ( .A1(n240), .A2(n247), .S0(n245), .Y(n246) );
  MUX21X1_HVT U117 ( .A1(n588), .A2(n288), .S0(n249), .Y(n248) );
  INVX0_HVT U119 ( .A(n288), .Y(n253) );
  IBUFFX2_HVT U120 ( .A(n568), .Y(n331) );
  IBUFFX2_HVT U121 ( .A(n557), .Y(n339) );
  MUX21X2_HVT U122 ( .A1(n568), .A2(n292), .S0(n282), .Y(n509) );
  INVX1_HVT U124 ( .A(in[1]), .Y(n249) );
  AO21X2_HVT U126 ( .A1(n249), .A2(n365), .A3(n310), .Y(n486) );
  XOR2X2_HVT U127 ( .A1(n310), .A2(n562), .Y(n545) );
  MUX41X1_HVT U129 ( .A1(n291), .A3(n348), .A2(n284), .A4(n332), .S0(n245), 
        .S1(n311), .Y(n444) );
  INVX1_HVT U130 ( .A(n310), .Y(n309) );
  IBUFFX2_HVT U132 ( .A(n310), .Y(n252) );
  INVX0_HVT U133 ( .A(n258), .Y(n471) );
  XOR2X1_HVT U134 ( .A1(n306), .A2(n310), .Y(n251) );
  INVX1_HVT U135 ( .A(n289), .Y(n257) );
  INVX0_HVT U137 ( .A(n558), .Y(n260) );
  MUX21X1_HVT U138 ( .A1(n399), .A2(n408), .S0(in[6]), .Y(out[6]) );
  INVX0_HVT U141 ( .A(n576), .Y(n259) );
  NAND2X0_HVT U142 ( .A1(n262), .A2(n254), .Y(n255) );
  NAND2X0_HVT U143 ( .A1(n572), .A2(n310), .Y(n256) );
  NAND2X0_HVT U145 ( .A1(n255), .A2(n256), .Y(n390) );
  MUX41X1_HVT U147 ( .A1(n339), .A3(n446), .A2(n342), .A4(n564), .S0(n245), 
        .S1(n311), .Y(n445) );
  MUX21X2_HVT U149 ( .A1(n501), .A2(n510), .S0(in[6]), .Y(out[1]) );
  MUX41X1_HVT U150 ( .A1(n424), .A3(n419), .A2(n422), .A4(n416), .S0(n257), 
        .S1(n241), .Y(n415) );
  XOR2X2_HVT U152 ( .A1(n370), .A2(in[3]), .Y(n582) );
  MUX41X1_HVT U155 ( .A1(n260), .A3(n564), .A2(n261), .A4(n259), .S0(n245), 
        .S1(n311), .Y(n258) );
  NAND2X0_HVT U156 ( .A1(n302), .A2(n284), .Y(n261) );
  MUX21X2_HVT U157 ( .A1(n529), .A2(n531), .S0(n274), .Y(n528) );
  MUX21X2_HVT U161 ( .A1(n439), .A2(n447), .S0(in[6]), .Y(out[4]) );
  INVX1_HVT U164 ( .A(in[2]), .Y(n306) );
  OA21X2_HVT U169 ( .A1(n341), .A2(n306), .A3(n329), .Y(n478) );
  MUX21X2_HVT U171 ( .A1(n480), .A2(n490), .S0(in[6]), .Y(out[2]) );
  XOR2X1_HVT U172 ( .A1(n298), .A2(n275), .Y(n541) );
  MUX21X2_HVT U173 ( .A1(n474), .A2(n296), .S0(n541), .Y(n473) );
  INVX0_HVT U175 ( .A(n582), .Y(n369) );
  MUX21X2_HVT U183 ( .A1(n267), .A2(n489), .S0(n251), .Y(n488) );
  MUX21X2_HVT U185 ( .A1(n260), .A2(n574), .S0(n276), .Y(n489) );
  INVX1_HVT U187 ( .A(n584), .Y(n364) );
  AND2X1_HVT U188 ( .A1(n286), .A2(n532), .Y(n262) );
  MUX21X1_HVT U191 ( .A1(n264), .A2(n327), .S0(n272), .Y(n456) );
  NBUFFX2_HVT U192 ( .A(n369), .Y(n284) );
  INVX1_HVT U193 ( .A(n587), .Y(n368) );
  NBUFFX2_HVT U196 ( .A(n584), .Y(n293) );
  MUX21X1_HVT U198 ( .A1(n364), .A2(n367), .S0(n279), .Y(n536) );
  MUX21X1_HVT U199 ( .A1(n323), .A2(n365), .S0(n279), .Y(n521) );
  MUX21X1_HVT U200 ( .A1(n558), .A2(n477), .S0(n272), .Y(n475) );
  AND2X1_HVT U202 ( .A1(n295), .A2(n515), .Y(n263) );
  MUX21X1_HVT U203 ( .A1(n295), .A2(n285), .S0(n301), .Y(n548) );
  MUX21X1_HVT U209 ( .A1(n293), .A2(n582), .S0(n212), .Y(n552) );
  MUX21X1_HVT U210 ( .A1(n284), .A2(n288), .S0(n218), .Y(n485) );
  MUX21X1_HVT U211 ( .A1(n582), .A2(n365), .S0(n218), .Y(n374) );
  MUX21X1_HVT U213 ( .A1(n368), .A2(n367), .S0(n300), .Y(n562) );
  MUX21X1_HVT U216 ( .A1(n367), .A2(n364), .S0(n300), .Y(n551) );
  MUX21X1_HVT U217 ( .A1(n283), .A2(n368), .S0(n300), .Y(n549) );
  MUX21X1_HVT U219 ( .A1(n364), .A2(n368), .S0(n213), .Y(n414) );
  MUX21X1_HVT U221 ( .A1(n367), .A2(n285), .S0(n218), .Y(n426) );
  MUX21X1_HVT U222 ( .A1(n285), .A2(n364), .S0(n298), .Y(n493) );
  NAND2X0_HVT U223 ( .A1(n287), .A2(n366), .Y(n584) );
  NBUFFX2_HVT U224 ( .A(n587), .Y(n294) );
  INVX1_HVT U225 ( .A(n588), .Y(n367) );
  MUX21X1_HVT U226 ( .A1(n582), .A2(n368), .S0(n212), .Y(n564) );
  NBUFFX2_HVT U227 ( .A(n587), .Y(n295) );
  MUX21X1_HVT U228 ( .A1(n293), .A2(n292), .S0(n301), .Y(n500) );
  MUX21X1_HVT U229 ( .A1(n582), .A2(n288), .S0(n212), .Y(n512) );
  XOR2X1_HVT U230 ( .A1(n582), .A2(n299), .Y(n543) );
  MUX21X1_HVT U231 ( .A1(n283), .A2(n582), .S0(n298), .Y(n377) );
  INVX1_HVT U232 ( .A(n579), .Y(n365) );
  MUX21X1_HVT U233 ( .A1(n367), .A2(n283), .S0(n212), .Y(n555) );
  MUX21X1_HVT U234 ( .A1(n293), .A2(n283), .S0(n213), .Y(n577) );
  MUX21X1_HVT U235 ( .A1(n288), .A2(n364), .S0(n213), .Y(n560) );
  MUX21X1_HVT U236 ( .A1(n365), .A2(n364), .S0(n301), .Y(n570) );
  MUX21X1_HVT U237 ( .A1(n315), .A2(n340), .S0(n272), .Y(n470) );
  MUX21X1_HVT U238 ( .A1(n338), .A2(n453), .S0(n275), .Y(n452) );
  MUX21X1_HVT U239 ( .A1(n359), .A2(n292), .S0(n281), .Y(n453) );
  XOR2X1_HVT U240 ( .A1(n294), .A2(n299), .Y(n540) );
  MUX21X1_HVT U241 ( .A1(n364), .A2(n287), .S0(n299), .Y(n375) );
  MUX21X1_HVT U242 ( .A1(n588), .A2(n291), .S0(n300), .Y(n558) );
  MUX21X1_HVT U243 ( .A1(n287), .A2(n283), .S0(n217), .Y(n466) );
  XOR2X1_HVT U244 ( .A1(n218), .A2(n365), .Y(n544) );
  MUX21X1_HVT U245 ( .A1(n296), .A2(n291), .S0(n300), .Y(n574) );
  MUX21X1_HVT U246 ( .A1(n584), .A2(n297), .S0(n299), .Y(n495) );
  MUX21X1_HVT U247 ( .A1(n283), .A2(n367), .S0(n300), .Y(n578) );
  NBUFFX2_HVT U248 ( .A(n587), .Y(n296) );
  MUX21X1_HVT U249 ( .A1(n366), .A2(n297), .S0(n298), .Y(n401) );
  MUX21X1_HVT U250 ( .A1(n588), .A2(n295), .S0(n217), .Y(n402) );
  MUX21X1_HVT U251 ( .A1(n291), .A2(n283), .S0(n299), .Y(n379) );
  MUX21X1_HVT U252 ( .A1(n294), .A2(n287), .S0(n217), .Y(n381) );
  XNOR2X1_HVT U253 ( .A1(n584), .A2(n298), .Y(n264) );
  XNOR2X1_HVT U254 ( .A1(n588), .A2(n217), .Y(n265) );
  AND2X1_HVT U255 ( .A1(n302), .A2(n368), .Y(n266) );
  MUX21X1_HVT U256 ( .A1(n294), .A2(n293), .S0(n218), .Y(n373) );
  AND2X1_HVT U257 ( .A1(n297), .A2(n476), .Y(n267) );
  MUX21X1_HVT U258 ( .A1(n292), .A2(n287), .S0(n213), .Y(n517) );
  MUX21X1_HVT U259 ( .A1(n292), .A2(n297), .S0(n275), .Y(n463) );
  XOR2X1_HVT U260 ( .A1(n287), .A2(n218), .Y(n563) );
  NBUFFX2_HVT U261 ( .A(n254), .Y(n280) );
  NBUFFX2_HVT U262 ( .A(n254), .Y(n281) );
  NBUFFX2_HVT U263 ( .A(n366), .Y(n283) );
  NBUFFX2_HVT U264 ( .A(n254), .Y(n282) );
  NBUFFX2_HVT U265 ( .A(n305), .Y(n272) );
  NBUFFX2_HVT U266 ( .A(n304), .Y(n274) );
  NBUFFX2_HVT U267 ( .A(n305), .Y(n273) );
  NBUFFX2_HVT U268 ( .A(in[5]), .Y(n278) );
  NBUFFX2_HVT U269 ( .A(n305), .Y(n275) );
  NBUFFX2_HVT U270 ( .A(n305), .Y(n276) );
  NBUFFX2_HVT U271 ( .A(n305), .Y(n271) );
  NBUFFX2_HVT U272 ( .A(n307), .Y(n277) );
  MUX21X1_HVT U273 ( .A1(n286), .A2(n290), .S0(n301), .Y(n566) );
  MUX21X1_HVT U274 ( .A1(n487), .A2(n338), .S0(n275), .Y(n484) );
  MUX21X1_HVT U275 ( .A1(n525), .A2(n527), .S0(n274), .Y(n524) );
  MUX21X1_HVT U276 ( .A1(n405), .A2(n406), .S0(n274), .Y(n404) );
  MUX21X1_HVT U277 ( .A1(n503), .A2(n290), .S0(n281), .Y(n406) );
  XOR2X1_HVT U278 ( .A1(n218), .A2(in[3]), .Y(n542) );
  MUX21X1_HVT U279 ( .A1(n291), .A2(n286), .S0(n301), .Y(n482) );
  NAND2X0_HVT U280 ( .A1(n290), .A2(n288), .Y(n587) );
  NBUFFX2_HVT U281 ( .A(n370), .Y(n288) );
  MUX21X1_HVT U282 ( .A1(n292), .A2(n354), .S0(n282), .Y(n418) );
  MUX21X1_HVT U283 ( .A1(n437), .A2(n438), .S0(n276), .Y(n435) );
  MUX21X1_HVT U284 ( .A1(n356), .A2(n365), .S0(n281), .Y(n438) );
  AND2X1_HVT U285 ( .A1(n286), .A2(n121), .Y(n268) );
  MUX21X1_HVT U286 ( .A1(n368), .A2(n290), .S0(n212), .Y(n569) );
  MUX21X1_HVT U287 ( .A1(n290), .A2(n364), .S0(n301), .Y(n550) );
  MUX21X1_HVT U288 ( .A1(n545), .A2(n519), .S0(n274), .Y(n518) );
  MUX21X1_HVT U289 ( .A1(n367), .A2(n354), .S0(n282), .Y(n519) );
  MUX21X1_HVT U290 ( .A1(n443), .A2(n442), .S0(n275), .Y(n441) );
  MUX21X1_HVT U291 ( .A1(n560), .A2(n318), .S0(n282), .Y(n443) );
  MUX21X1_HVT U292 ( .A1(n365), .A2(n368), .S0(n217), .Y(n423) );
  MUX21X1_HVT U293 ( .A1(n248), .A2(n586), .S0(n273), .Y(n479) );
  MUX21X1_HVT U294 ( .A1(n431), .A2(n432), .S0(n276), .Y(n430) );
  MUX21X1_HVT U295 ( .A1(n433), .A2(n296), .S0(n269), .Y(n432) );
  MUX21X1_HVT U296 ( .A1(n551), .A2(n357), .S0(n280), .Y(n431) );
  MUX21X1_HVT U297 ( .A1(n571), .A2(n339), .S0(n273), .Y(n455) );
  XOR2X1_HVT U298 ( .A1(n298), .A2(n278), .Y(n546) );
  MUX21X1_HVT U299 ( .A1(n346), .A2(n362), .S0(n281), .Y(n394) );
  NBUFFX2_HVT U300 ( .A(n579), .Y(n291) );
  MUX21X1_HVT U301 ( .A1(n586), .A2(n249), .S0(n274), .Y(n462) );
  MUX21X1_HVT U302 ( .A1(n290), .A2(n365), .S0(n217), .Y(n378) );
  MUX21X1_HVT U303 ( .A1(n325), .A2(n121), .S0(n279), .Y(n523) );
  NBUFFX2_HVT U304 ( .A(n588), .Y(n297) );
  MUX21X1_HVT U305 ( .A1(n559), .A2(n382), .S0(n280), .Y(n376) );
  MUX21X1_HVT U306 ( .A1(n293), .A2(n290), .S0(n212), .Y(n580) );
  MUX21X1_HVT U307 ( .A1(n335), .A2(n559), .S0(n273), .Y(n458) );
  MUX21X1_HVT U308 ( .A1(n296), .A2(n498), .S0(n269), .Y(n497) );
  MUX21X1_HVT U309 ( .A1(n290), .A2(n287), .S0(n282), .Y(n498) );
  NBUFFX2_HVT U310 ( .A(n370), .Y(n287) );
  NBUFFX2_HVT U311 ( .A(n579), .Y(n292) );
  INVX1_HVT U312 ( .A(n249), .Y(n298) );
  XNOR2X1_HVT U313 ( .A1(n310), .A2(n299), .Y(n269) );
  AND2X1_HVT U314 ( .A1(n283), .A2(n121), .Y(n270) );
  NBUFFX2_HVT U315 ( .A(in[5]), .Y(n307) );
  MUX21X1_HVT U316 ( .A1(n394), .A2(n393), .S0(n274), .Y(n392) );
  MUX21X1_HVT U317 ( .A1(n496), .A2(n497), .S0(n276), .Y(n494) );
  MUX21X1_HVT U318 ( .A1(n364), .A2(n253), .S0(n213), .Y(n557) );
  NAND2X0_HVT U319 ( .A1(in[3]), .A2(in[4]), .Y(n588) );
  NAND2X0_HVT U320 ( .A1(in[4]), .A2(n366), .Y(n579) );
  MUX21X1_HVT U321 ( .A1(n253), .A2(n582), .S0(n217), .Y(n380) );
  MUX21X1_HVT U322 ( .A1(n253), .A2(n365), .S0(n213), .Y(n571) );
  MUX21X1_HVT U323 ( .A1(n253), .A2(n291), .S0(n298), .Y(n372) );
  MUX21X1_HVT U324 ( .A1(n253), .A2(n297), .S0(n301), .Y(n371) );
  MUX21X1_HVT U325 ( .A1(n297), .A2(n253), .S0(n212), .Y(n561) );
  MUX21X1_HVT U326 ( .A1(n290), .A2(n253), .S0(n272), .Y(n474) );
  MUX21X1_HVT U327 ( .A1(n283), .A2(n253), .S0(n213), .Y(n559) );
  NBUFFX2_HVT U328 ( .A(in[3]), .Y(n290) );
  NBUFFX2_HVT U329 ( .A(in[0]), .Y(n289) );
  INVX0_HVT U330 ( .A(n567), .Y(n312) );
  INVX0_HVT U331 ( .A(n565), .Y(n313) );
  INVX0_HVT U332 ( .A(n556), .Y(n314) );
  INVX0_HVT U333 ( .A(n420), .Y(n316) );
  INVX0_HVT U334 ( .A(n383), .Y(n317) );
  INVX0_HVT U335 ( .A(n586), .Y(n318) );
  INVX0_HVT U336 ( .A(n573), .Y(n319) );
  INVX0_HVT U337 ( .A(n585), .Y(n320) );
  INVX0_HVT U338 ( .A(n583), .Y(n321) );
  INVX0_HVT U339 ( .A(n581), .Y(n322) );
  INVX0_HVT U340 ( .A(n580), .Y(n323) );
  INVX0_HVT U341 ( .A(n578), .Y(n324) );
  INVX0_HVT U342 ( .A(n577), .Y(n325) );
  INVX0_HVT U343 ( .A(n574), .Y(n326) );
  INVX0_HVT U344 ( .A(n572), .Y(n327) );
  INVX0_HVT U345 ( .A(n571), .Y(n328) );
  INVX0_HVT U346 ( .A(n570), .Y(n329) );
  INVX0_HVT U347 ( .A(n569), .Y(n330) );
  INVX0_HVT U348 ( .A(n566), .Y(n332) );
  INVX0_HVT U349 ( .A(n564), .Y(n333) );
  INVX0_HVT U350 ( .A(n563), .Y(n334) );
  INVX0_HVT U351 ( .A(n561), .Y(n335) );
  INVX0_HVT U352 ( .A(n560), .Y(n336) );
  INVX0_HVT U353 ( .A(n559), .Y(n337) );
  INVX0_HVT U354 ( .A(n376), .Y(n338) );
  INVX0_HVT U355 ( .A(n555), .Y(n340) );
  INVX0_HVT U356 ( .A(n552), .Y(n341) );
  INVX0_HVT U357 ( .A(n551), .Y(n342) );
  INVX0_HVT U358 ( .A(n550), .Y(n343) );
  INVX0_HVT U359 ( .A(n549), .Y(n344) );
  INVX0_HVT U360 ( .A(n548), .Y(n345) );
  INVX0_HVT U361 ( .A(n547), .Y(n346) );
  INVX0_HVT U362 ( .A(n515), .Y(n347) );
  INVX0_HVT U363 ( .A(n476), .Y(n348) );
  INVX0_HVT U364 ( .A(n382), .Y(n349) );
  INVX0_HVT U365 ( .A(n532), .Y(n350) );
  INVX0_HVT U366 ( .A(n436), .Y(n351) );
  INVX0_HVT U367 ( .A(n381), .Y(n352) );
  INVX0_HVT U368 ( .A(n380), .Y(n353) );
  INVX0_HVT U369 ( .A(n379), .Y(n354) );
  INVX0_HVT U370 ( .A(n378), .Y(n355) );
  INVX0_HVT U371 ( .A(n377), .Y(n356) );
  INVX0_HVT U372 ( .A(n495), .Y(n357) );
  INVX0_HVT U373 ( .A(n485), .Y(n358) );
  INVX0_HVT U374 ( .A(n375), .Y(n359) );
  INVX0_HVT U375 ( .A(n374), .Y(n360) );
  INVX0_HVT U376 ( .A(n373), .Y(n361) );
  INVX0_HVT U377 ( .A(n372), .Y(n362) );
  INVX0_HVT U378 ( .A(n371), .Y(n363) );
endmodule

