
module sbox_8 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n95, n96, n210, n211, n212, n213, n216, n217, n218, n219, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594;

  NAND2X0_HVT U4 ( .A1(n304), .A2(n592), .Y(n591) );
  NAND2X0_HVT U5 ( .A1(n95), .A2(n297), .Y(n589) );
  NAND2X0_HVT U13 ( .A1(n581), .A2(n308), .Y(n582) );
  NAND2X0_HVT U15 ( .A1(n592), .A2(n264), .Y(n579) );
  NAND2X0_HVT U21 ( .A1(n304), .A2(n314), .Y(n573) );
  NAND2X0_HVT U24 ( .A1(n299), .A2(n314), .Y(n571) );
  NAND2X0_HVT U33 ( .A1(n370), .A2(n314), .Y(n562) );
  NAND2X0_HVT U35 ( .A1(n237), .A2(n314), .Y(n560) );
  NAND2X0_HVT U42 ( .A1(n311), .A2(n299), .Y(n553) );
  MUX41X1_HVT U51 ( .A1(n358), .A3(n318), .A2(n336), .A4(n337), .S0(n273), 
        .S1(n292), .Y(n544) );
  NAND2X0_HVT U53 ( .A1(n541), .A2(n552), .Y(n542) );
  NAND2X0_HVT U56 ( .A1(n304), .A2(n537), .Y(n538) );
  MUX41X1_HVT U57 ( .A1(n359), .A3(n575), .A2(n538), .A4(n584), .S0(n273), 
        .S1(n292), .Y(n536) );
  NAND2X0_HVT U58 ( .A1(n308), .A2(n592), .Y(n535) );
  MUX41X1_HVT U59 ( .A1(n286), .A3(n535), .A2(n284), .A4(n335), .S0(n273), 
        .S1(n292), .Y(n534) );
  MUX41X1_HVT U61 ( .A1(n282), .A3(n334), .A2(n333), .A4(n262), .S0(n273), 
        .S1(n292), .Y(n532) );
  NAND2X0_HVT U62 ( .A1(n314), .A2(n306), .Y(n531) );
  MUX41X1_HVT U63 ( .A1(n531), .A3(n325), .A2(n353), .A4(n332), .S0(n273), 
        .S1(n292), .Y(n530) );
  AO21X1_HVT U66 ( .A1(n330), .A2(in[5]), .A3(n352), .Y(n527) );
  MUX41X1_HVT U68 ( .A1(n328), .A3(n527), .A2(n526), .A4(n528), .S0(n287), 
        .S1(n270), .Y(n525) );
  MUX41X1_HVT U69 ( .A1(n525), .A3(n533), .A2(n529), .A4(n539), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n301), .A2(n520), .Y(n521) );
  MUX41X1_HVT U74 ( .A1(n522), .A3(n569), .A2(n521), .A4(n571), .S0(n288), 
        .S1(n244), .Y(n519) );
  MUX41X1_HVT U75 ( .A1(n356), .A3(n361), .A2(n374), .A4(n339), .S0(n287), 
        .S1(n244), .Y(n518) );
  MUX41X1_HVT U77 ( .A1(n586), .A3(n363), .A2(n517), .A4(n362), .S0(n294), 
        .S1(n249), .Y(n516) );
  MUX41X1_HVT U78 ( .A1(n516), .A3(n519), .A2(n518), .A4(n523), .S0(in[0]), 
        .S1(n292), .Y(n515) );
  AND3X1_HVT U80 ( .A1(n305), .A2(n537), .A3(n512), .Y(n513) );
  MUX41X1_HVT U82 ( .A1(n550), .A3(n337), .A2(n319), .A4(n580), .S0(n287), 
        .S1(n270), .Y(n510) );
  AND2X1_HVT U83 ( .A1(n23), .A2(n255), .Y(n509) );
  MUX41X1_HVT U84 ( .A1(n338), .A3(n258), .A2(n578), .A4(n509), .S0(n287), 
        .S1(n244), .Y(n508) );
  NAND2X0_HVT U85 ( .A1(n314), .A2(n373), .Y(n507) );
  MUX41X1_HVT U86 ( .A1(n361), .A3(n507), .A2(n283), .A4(n279), .S0(n287), 
        .S1(n270), .Y(n506) );
  MUX41X1_HVT U87 ( .A1(n506), .A3(n510), .A2(n508), .A4(n511), .S0(in[0]), 
        .S1(n291), .Y(n505) );
  MUX41X1_HVT U90 ( .A1(n549), .A3(n553), .A2(n358), .A4(n504), .S0(n266), 
        .S1(n270), .Y(n503) );
  MUX41X1_HVT U96 ( .A1(n319), .A3(n281), .A2(n360), .A4(n499), .S0(n287), 
        .S1(n270), .Y(n498) );
  MUX41X1_HVT U97 ( .A1(n356), .A3(n281), .A2(n312), .A4(n579), .S0(n287), 
        .S1(n270), .Y(n497) );
  MUX41X1_HVT U98 ( .A1(n497), .A3(n500), .A2(n498), .A4(n503), .S0(n298), 
        .S1(n291), .Y(n496) );
  NAND2X0_HVT U101 ( .A1(n492), .A2(n491), .Y(n493) );
  MUX41X1_HVT U103 ( .A1(n592), .A3(n329), .A2(n233), .A4(n560), .S0(n287), 
        .S1(n317), .Y(n489) );
  MUX41X1_HVT U105 ( .A1(n341), .A3(n547), .A2(n488), .A4(n355), .S0(n287), 
        .S1(n316), .Y(n487) );
  OA21X1_HVT U109 ( .A1(n346), .A2(n219), .A3(n335), .Y(n484) );
  NAND2X0_HVT U110 ( .A1(n305), .A2(n482), .Y(n483) );
  AND2X1_HVT U115 ( .A1(n309), .A2(n261), .Y(n477) );
  MUX41X1_HVT U116 ( .A1(n582), .A3(n477), .A2(n339), .A4(n564), .S0(n289), 
        .S1(n273), .Y(n476) );
  NAND2X0_HVT U123 ( .A1(n468), .A2(n467), .Y(n469) );
  MUX41X1_HVT U125 ( .A1(n573), .A3(n286), .A2(n328), .A4(n365), .S0(n249), 
        .S1(n273), .Y(n465) );
  MUX41X1_HVT U131 ( .A1(n460), .A3(n462), .A2(n461), .A4(n463), .S0(in[5]), 
        .S1(n273), .Y(n459) );
  MUX41X1_HVT U132 ( .A1(n459), .A3(n472), .A2(n464), .A4(n478), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  AND2X1_HVT U140 ( .A1(n300), .A2(n313), .Y(n451) );
  MUX41X1_HVT U141 ( .A1(n570), .A3(n347), .A2(n451), .A4(n344), .S0(n288), 
        .S1(n316), .Y(n450) );
  MUX41X1_HVT U147 ( .A1(n367), .A3(n520), .A2(n356), .A4(n549), .S0(n288), 
        .S1(n316), .Y(n445) );
  OA21X1_HVT U151 ( .A1(n555), .A2(n248), .A3(n441), .Y(n442) );
  MUX41X1_HVT U153 ( .A1(n483), .A3(n282), .A2(n593), .A4(n321), .S0(n290), 
        .S1(n317), .Y(n439) );
  AND2X1_HVT U154 ( .A1(n296), .A2(n299), .Y(n438) );
  NAND2X0_HVT U158 ( .A1(n96), .A2(n373), .Y(n434) );
  MUX41X1_HVT U159 ( .A1(n582), .A3(n264), .A2(n434), .A4(n327), .S0(n315), 
        .S1(n244), .Y(n433) );
  AND2X1_HVT U162 ( .A1(n258), .A2(n520), .Y(n430) );
  MUX41X1_HVT U163 ( .A1(n334), .A3(n430), .A2(n280), .A4(n431), .S0(n315), 
        .S1(n244), .Y(n429) );
  MUX41X1_HVT U165 ( .A1(n573), .A3(n342), .A2(n549), .A4(n428), .S0(n273), 
        .S1(n315), .Y(n427) );
  NAND2X0_HVT U166 ( .A1(n308), .A2(n537), .Y(n426) );
  NAND2X0_HVT U167 ( .A1(n374), .A2(n314), .Y(n425) );
  MUX41X1_HVT U168 ( .A1(n359), .A3(n300), .A2(n425), .A4(n426), .S0(n266), 
        .S1(n317), .Y(n424) );
  MUX41X1_HVT U172 ( .A1(n421), .A3(n427), .A2(n424), .A4(n429), .S0(in[0]), 
        .S1(n291), .Y(n420) );
  NAND2X0_HVT U174 ( .A1(n309), .A2(n259), .Y(n581) );
  MUX41X1_HVT U176 ( .A1(n237), .A3(n419), .A2(n364), .A4(n581), .S0(n295), 
        .S1(n290), .Y(n418) );
  NAND2X0_HVT U177 ( .A1(n95), .A2(n237), .Y(n417) );
  MUX41X1_HVT U178 ( .A1(n577), .A3(n417), .A2(n368), .A4(n557), .S0(n288), 
        .S1(n316), .Y(n416) );
  MUX41X1_HVT U179 ( .A1(n567), .A3(n369), .A2(n323), .A4(n368), .S0(n315), 
        .S1(n317), .Y(n415) );
  MUX41X1_HVT U180 ( .A1(n326), .A3(n586), .A2(n582), .A4(n278), .S0(n294), 
        .S1(n266), .Y(n414) );
  MUX41X1_HVT U181 ( .A1(n414), .A3(n416), .A2(n415), .A4(n418), .S0(n298), 
        .S1(n293), .Y(n413) );
  MUX41X1_HVT U182 ( .A1(n348), .A3(n303), .A2(n350), .A4(n340), .S0(n244), 
        .S1(n249), .Y(n412) );
  OA21X1_HVT U184 ( .A1(n561), .A2(n248), .A3(n338), .Y(n410) );
  MUX41X1_HVT U186 ( .A1(n281), .A3(n556), .A2(n520), .A4(n549), .S0(n287), 
        .S1(n317), .Y(n408) );
  MUX41X1_HVT U189 ( .A1(n406), .A3(n581), .A2(n407), .A4(n355), .S0(n294), 
        .S1(n315), .Y(n405) );
  MUX41X1_HVT U193 ( .A1(n553), .A3(n560), .A2(n545), .A4(n403), .S0(n249), 
        .S1(n316), .Y(n402) );
  MUX41X1_HVT U194 ( .A1(n554), .A3(n568), .A2(n366), .A4(n300), .S0(n294), 
        .S1(n315), .Y(n401) );
  MUX41X1_HVT U195 ( .A1(n259), .A3(n360), .A2(n307), .A4(n558), .S0(n289), 
        .S1(n270), .Y(n400) );
  AO21X1_HVT U197 ( .A1(n283), .A2(n295), .A3(n357), .Y(n398) );
  MUX41X1_HVT U199 ( .A1(n397), .A3(n401), .A2(n400), .A4(n402), .S0(in[0]), 
        .S1(n293), .Y(n396) );
  MUX41X1_HVT U204 ( .A1(n538), .A3(n582), .A2(n345), .A4(n572), .S0(n315), 
        .S1(n317), .Y(n391) );
  MUX41X1_HVT U205 ( .A1(n255), .A3(n592), .A2(n369), .A4(n238), .S0(n290), 
        .S1(n317), .Y(n390) );
  NAND2X0_HVT U208 ( .A1(n311), .A2(n304), .Y(n482) );
  NAND2X0_HVT U212 ( .A1(n95), .A2(n301), .Y(n537) );
  NAND2X0_HVT U214 ( .A1(n259), .A2(n314), .Y(n388) );
  NAND2X0_HVT U215 ( .A1(n482), .A2(n302), .Y(n387) );
  AO21X1_HVT U216 ( .A1(n313), .A2(n371), .A3(n248), .Y(n492) );
  NAND2X0_HVT U218 ( .A1(n371), .A2(n23), .Y(n441) );
  NAND2X0_HVT U220 ( .A1(n295), .A2(n388), .Y(n512) );
  INVX2_HVT U1 ( .A(n247), .Y(n317) );
  NBUFFX2_HVT U2 ( .A(in[1]), .Y(n23) );
  INVX1_HVT U3 ( .A(in[1]), .Y(n313) );
  INVX0_HVT U6 ( .A(n313), .Y(n310) );
  INVX0_HVT U7 ( .A(n313), .Y(n95) );
  INVX2_HVT U8 ( .A(n247), .Y(n316) );
  INVX1_HVT U9 ( .A(n294), .Y(n247) );
  XOR2X1_HVT U10 ( .A1(n258), .A2(n23), .Y(n549) );
  INVX0_HVT U11 ( .A(n313), .Y(n311) );
  INVX0_HVT U12 ( .A(n313), .Y(n96) );
  INVX0_HVT U14 ( .A(n307), .Y(n239) );
  NAND2X0_HVT U16 ( .A1(n267), .A2(n268), .Y(n453) );
  INVX0_HVT U17 ( .A(n238), .Y(n564) );
  MUX41X1_HVT U18 ( .A1(n338), .A3(n265), .A2(n354), .A4(n300), .S0(n266), 
        .S1(n316), .Y(n449) );
  INVX0_HVT U19 ( .A(n482), .Y(n354) );
  MUX21X1_HVT U20 ( .A1(n483), .A2(n564), .S0(n219), .Y(n481) );
  NAND2X0_HVT U22 ( .A1(n241), .A2(n242), .Y(out[1]) );
  NAND2X0_HVT U23 ( .A1(n389), .A2(n210), .Y(n234) );
  XOR2X1_HVT U25 ( .A1(n248), .A2(n568), .Y(n551) );
  MUX21X1_HVT U26 ( .A1(n297), .A2(n262), .S0(n313), .Y(n578) );
  INVX0_HVT U27 ( .A(n313), .Y(n312) );
  INVX0_HVT U28 ( .A(n313), .Y(n309) );
  INVX0_HVT U29 ( .A(n218), .Y(n500) );
  MUX21X1_HVT U30 ( .A1(n238), .A2(n580), .S0(n266), .Y(n495) );
  NAND2X0_HVT U31 ( .A1(n310), .A2(n308), .Y(n520) );
  NAND2X0_HVT U32 ( .A1(n310), .A2(n305), .Y(n592) );
  INVX1_HVT U34 ( .A(n293), .Y(n274) );
  INVX0_HVT U36 ( .A(n257), .Y(n263) );
  INVX1_HVT U37 ( .A(n588), .Y(n256) );
  INVX0_HVT U38 ( .A(n588), .Y(n257) );
  NAND2X0_HVT U39 ( .A1(n253), .A2(n254), .Y(out[4]) );
  INVX1_HVT U40 ( .A(n298), .Y(n243) );
  INVX1_HVT U41 ( .A(in[3]), .Y(n372) );
  INVX1_HVT U43 ( .A(in[6]), .Y(n210) );
  NAND2X0_HVT U44 ( .A1(n211), .A2(n212), .Y(out[5]) );
  INVX1_HVT U45 ( .A(n269), .Y(n266) );
  INVX0_HVT U46 ( .A(n290), .Y(n252) );
  INVX1_HVT U47 ( .A(n252), .Y(n249) );
  INVX0_HVT U48 ( .A(in[2]), .Y(n269) );
  INVX0_HVT U49 ( .A(n290), .Y(n219) );
  INVX1_HVT U50 ( .A(n296), .Y(n248) );
  INVX1_HVT U52 ( .A(n247), .Y(n244) );
  INVX0_HVT U54 ( .A(in[4]), .Y(n237) );
  INVX0_HVT U55 ( .A(n233), .Y(n566) );
  MUX21X2_HVT U60 ( .A1(n410), .A2(n411), .S0(n289), .Y(n409) );
  MUX41X1_HVT U64 ( .A1(n457), .A3(n456), .A2(n455), .A4(n453), .S0(n274), 
        .S1(n243), .Y(n452) );
  MUX21X2_HVT U65 ( .A1(n458), .A2(n343), .S0(n252), .Y(n457) );
  IBUFFX2_HVT U67 ( .A(n520), .Y(n352) );
  NAND2X0_HVT U70 ( .A1(n420), .A2(n210), .Y(n211) );
  NAND2X0_HVT U71 ( .A1(n432), .A2(in[6]), .Y(n212) );
  MUX21X1_HVT U72 ( .A1(n557), .A2(n363), .S0(n294), .Y(n436) );
  NAND2X0_HVT U76 ( .A1(n306), .A2(n213), .Y(n216) );
  NAND2X0_HVT U79 ( .A1(n502), .A2(n285), .Y(n217) );
  INVX0_HVT U81 ( .A(n285), .Y(n213) );
  MUX21X1_HVT U88 ( .A1(n231), .A2(n232), .S0(n219), .Y(n218) );
  AND2X1_HVT U89 ( .A1(n216), .A2(n217), .Y(n231) );
  AOI21X1_HVT U91 ( .A1(n296), .A2(n501), .A3(n357), .Y(n232) );
  MUX21X1_HVT U92 ( .A1(n255), .A2(n303), .S0(n96), .Y(n233) );
  MUX41X1_HVT U93 ( .A1(n435), .A3(n440), .A2(n433), .A4(n439), .S0(n298), 
        .S1(n274), .Y(n432) );
  INVX1_HVT U94 ( .A(n236), .Y(n559) );
  NAND2X0_HVT U95 ( .A1(n396), .A2(in[6]), .Y(n235) );
  NAND2X0_HVT U99 ( .A1(n234), .A2(n235), .Y(out[7]) );
  MUX21X2_HVT U100 ( .A1(n566), .A2(n324), .S0(n296), .Y(n448) );
  INVX0_HVT U102 ( .A(n580), .Y(n332) );
  MUX21X2_HVT U104 ( .A1(n413), .A2(n404), .S0(n210), .Y(out[6]) );
  MUX21X2_HVT U106 ( .A1(n436), .A2(n437), .S0(n288), .Y(n435) );
  MUX21X1_HVT U107 ( .A1(n237), .A2(n307), .S0(n96), .Y(n236) );
  MUX21X1_HVT U108 ( .A1(n239), .A2(n371), .S0(n95), .Y(n238) );
  MUX41X1_HVT U111 ( .A1(n494), .A3(n489), .A2(n490), .A4(n487), .S0(n243), 
        .S1(n274), .Y(n486) );
  MUX21X2_HVT U112 ( .A1(n476), .A2(n473), .S0(n274), .Y(n472) );
  MUX41X1_HVT U113 ( .A1(n559), .A3(n367), .A2(n562), .A4(n279), .S0(n219), 
        .S1(n248), .Y(n455) );
  OA21X2_HVT U114 ( .A1(n284), .A2(n248), .A3(n564), .Y(n422) );
  NAND2X0_HVT U117 ( .A1(n515), .A2(n240), .Y(n241) );
  NAND2X0_HVT U118 ( .A1(n505), .A2(n210), .Y(n242) );
  INVX1_HVT U119 ( .A(n210), .Y(n240) );
  NAND2X0_HVT U120 ( .A1(n387), .A2(n316), .Y(n245) );
  NAND2X0_HVT U121 ( .A1(n565), .A2(n247), .Y(n246) );
  NAND2X0_HVT U122 ( .A1(n245), .A2(n246), .Y(n381) );
  INVX0_HVT U124 ( .A(n381), .Y(n343) );
  MUX41X1_HVT U126 ( .A1(n568), .A3(n589), .A2(n371), .A4(n366), .S0(n219), 
        .S1(n248), .Y(n456) );
  OA21X1_HVT U127 ( .A1(n322), .A2(n248), .A3(n564), .Y(n447) );
  MUX41X1_HVT U128 ( .A1(n445), .A3(n446), .A2(n449), .A4(n450), .S0(n291), 
        .S1(n298), .Y(n444) );
  MUX21X2_HVT U129 ( .A1(n302), .A2(n574), .S0(n248), .Y(n514) );
  NAND2X0_HVT U130 ( .A1(n447), .A2(n249), .Y(n250) );
  NAND2X0_HVT U133 ( .A1(n448), .A2(n252), .Y(n251) );
  NAND2X0_HVT U134 ( .A1(n251), .A2(n250), .Y(n446) );
  MUX21X2_HVT U135 ( .A1(n514), .A2(n513), .S0(n249), .Y(n511) );
  MUX21X1_HVT U136 ( .A1(n373), .A2(n262), .S0(n310), .Y(n431) );
  NAND2X0_HVT U137 ( .A1(n452), .A2(n240), .Y(n253) );
  NAND2X0_HVT U138 ( .A1(n444), .A2(n210), .Y(n254) );
  MUX21X2_HVT U139 ( .A1(n486), .A2(n496), .S0(in[6]), .Y(out[2]) );
  INVX1_HVT U142 ( .A(n375), .Y(n255) );
  MUX41X1_HVT U143 ( .A1(n390), .A3(n392), .A2(n391), .A4(n393), .S0(in[0]), 
        .S1(n293), .Y(n389) );
  INVX1_HVT U144 ( .A(n256), .Y(n258) );
  INVX1_HVT U145 ( .A(n257), .Y(n259) );
  INVX1_HVT U146 ( .A(n256), .Y(n260) );
  INVX1_HVT U148 ( .A(n260), .Y(n261) );
  INVX1_HVT U149 ( .A(n260), .Y(n262) );
  INVX1_HVT U150 ( .A(n263), .Y(n264) );
  INVX1_HVT U152 ( .A(n263), .Y(n265) );
  XOR2X1_HVT U155 ( .A1(n375), .A2(in[3]), .Y(n588) );
  MUX21X2_HVT U156 ( .A1(n572), .A2(n348), .S0(n295), .Y(n454) );
  AO21X2_HVT U157 ( .A1(n289), .A2(n300), .A3(n259), .Y(n474) );
  INVX1_HVT U160 ( .A(n572), .Y(n338) );
  NAND2X0_HVT U161 ( .A1(n591), .A2(n266), .Y(n267) );
  NAND2X0_HVT U164 ( .A1(n454), .A2(n269), .Y(n268) );
  MUX21X1_HVT U169 ( .A1(n261), .A2(n299), .S0(in[1]), .Y(n572) );
  MUX21X2_HVT U170 ( .A1(n530), .A2(n532), .S0(n289), .Y(n529) );
  MUX21X1_HVT U171 ( .A1(n373), .A2(n264), .S0(n314), .Y(n587) );
  OA21X1_HVT U173 ( .A1(n587), .A2(n248), .A3(n347), .Y(n394) );
  INVX1_HVT U175 ( .A(n587), .Y(n328) );
  AND3X2_HVT U183 ( .A1(n290), .A2(n314), .A3(n255), .Y(n462) );
  INVX1_HVT U185 ( .A(n247), .Y(n270) );
  MUX41X1_HVT U187 ( .A1(n349), .A3(n559), .A2(n563), .A4(n583), .S0(n252), 
        .S1(n244), .Y(n392) );
  INVX2_HVT U188 ( .A(n269), .Y(n315) );
  NAND2X0_HVT U190 ( .A1(n394), .A2(n219), .Y(n271) );
  NAND2X0_HVT U191 ( .A1(n395), .A2(n289), .Y(n272) );
  NAND2X0_HVT U192 ( .A1(n271), .A2(n272), .Y(n393) );
  MUX21X1_HVT U196 ( .A1(n578), .A2(n278), .S0(n294), .Y(n395) );
  MUX41X1_HVT U198 ( .A1(n412), .A3(n409), .A2(n408), .A4(n405), .S0(n274), 
        .S1(n243), .Y(n404) );
  NBUFFX2_HVT U200 ( .A(n296), .Y(n273) );
  MUX41X1_HVT U201 ( .A1(n485), .A3(n484), .A2(n479), .A4(n481), .S0(n317), 
        .S1(n274), .Y(n478) );
  NAND2X0_HVT U202 ( .A1(n480), .A2(n275), .Y(n276) );
  NAND2X0_HVT U203 ( .A1(n306), .A2(n546), .Y(n277) );
  NAND2X0_HVT U206 ( .A1(n277), .A2(n276), .Y(n479) );
  INVX0_HVT U207 ( .A(n546), .Y(n275) );
  XOR2X1_HVT U209 ( .A1(n96), .A2(n315), .Y(n546) );
  MUX21X2_HVT U210 ( .A1(n282), .A2(n495), .S0(n548), .Y(n494) );
  INVX1_HVT U211 ( .A(n303), .Y(n370) );
  MUX21X1_HVT U213 ( .A1(n280), .A2(n333), .S0(n266), .Y(n461) );
  AND2X1_HVT U217 ( .A1(n262), .A2(n537), .Y(n278) );
  NBUFFX2_HVT U219 ( .A(n590), .Y(n303) );
  INVX1_HVT U221 ( .A(n593), .Y(n374) );
  MUX21X1_HVT U222 ( .A1(n370), .A2(n373), .S0(in[5]), .Y(n541) );
  NBUFFX2_HVT U223 ( .A(n590), .Y(n304) );
  MUX21X1_HVT U224 ( .A1(n329), .A2(n371), .S0(in[5]), .Y(n526) );
  AND2X1_HVT U225 ( .A1(n305), .A2(n520), .Y(n279) );
  MUX21X1_HVT U226 ( .A1(n465), .A2(n466), .S0(n291), .Y(n464) );
  MUX21X1_HVT U227 ( .A1(n470), .A2(n469), .S0(n296), .Y(n466) );
  MUX21X1_HVT U228 ( .A1(n305), .A2(n265), .S0(n312), .Y(n554) );
  MUX21X1_HVT U229 ( .A1(n261), .A2(n237), .S0(n311), .Y(n491) );
  MUX21X1_HVT U230 ( .A1(n370), .A2(n374), .S0(n95), .Y(n419) );
  MUX21X1_HVT U231 ( .A1(n258), .A2(n374), .S0(n96), .Y(n570) );
  MUX21X1_HVT U232 ( .A1(n304), .A2(n258), .S0(n96), .Y(n558) );
  MUX21X1_HVT U233 ( .A1(n264), .A2(n370), .S0(n312), .Y(n499) );
  MUX21X1_HVT U234 ( .A1(n259), .A2(n371), .S0(n96), .Y(n379) );
  MUX21X1_HVT U235 ( .A1(n304), .A2(n302), .S0(n95), .Y(n504) );
  MUX21X1_HVT U236 ( .A1(n259), .A2(n375), .S0(n311), .Y(n517) );
  MUX21X1_HVT U237 ( .A1(n374), .A2(n373), .S0(n23), .Y(n568) );
  MUX21X1_HVT U238 ( .A1(n373), .A2(n370), .S0(n311), .Y(n557) );
  MUX21X1_HVT U239 ( .A1(n373), .A2(n297), .S0(n310), .Y(n561) );
  MUX21X1_HVT U240 ( .A1(n297), .A2(n374), .S0(n23), .Y(n555) );
  MUX21X1_HVT U241 ( .A1(n365), .A2(n302), .S0(n295), .Y(n458) );
  MUX21X1_HVT U242 ( .A1(n474), .A2(n475), .S0(n295), .Y(n473) );
  MUX21X1_HVT U243 ( .A1(n321), .A2(n345), .S0(n266), .Y(n475) );
  NAND2X0_HVT U244 ( .A1(n237), .A2(n372), .Y(n590) );
  MUX21X1_HVT U245 ( .A1(n370), .A2(n237), .S0(n310), .Y(n380) );
  MUX21X1_HVT U246 ( .A1(n297), .A2(n258), .S0(n23), .Y(n382) );
  INVX1_HVT U247 ( .A(n307), .Y(n373) );
  MUX21X1_HVT U248 ( .A1(n320), .A2(n471), .S0(n288), .Y(n470) );
  MUX21X1_HVT U249 ( .A1(n375), .A2(n297), .S0(n309), .Y(n471) );
  NBUFFX2_HVT U250 ( .A(n593), .Y(n305) );
  XOR2X1_HVT U251 ( .A1(n311), .A2(n371), .Y(n550) );
  MUX21X1_HVT U252 ( .A1(n297), .A2(n308), .S0(n312), .Y(n406) );
  MUX21X1_HVT U253 ( .A1(n307), .A2(n305), .S0(n310), .Y(n407) );
  MUX21X1_HVT U254 ( .A1(n371), .A2(n370), .S0(n312), .Y(n576) );
  INVX1_HVT U255 ( .A(n300), .Y(n371) );
  MUX21X1_HVT U256 ( .A1(n306), .A2(n301), .S0(n310), .Y(n580) );
  MUX21X1_HVT U257 ( .A1(n303), .A2(n308), .S0(n95), .Y(n501) );
  MUX21X1_HVT U258 ( .A1(n297), .A2(n373), .S0(n23), .Y(n584) );
  XOR2X1_HVT U259 ( .A1(n315), .A2(n295), .Y(n548) );
  NBUFFX2_HVT U260 ( .A(n593), .Y(n306) );
  MUX21X1_HVT U261 ( .A1(n297), .A2(n375), .S0(n96), .Y(n403) );
  XOR2X1_HVT U262 ( .A1(n306), .A2(n309), .Y(n545) );
  MUX21X1_HVT U263 ( .A1(n306), .A2(n375), .S0(n311), .Y(n386) );
  XNOR2X1_HVT U264 ( .A1(n303), .A2(n311), .Y(n280) );
  AND2X1_HVT U265 ( .A1(n310), .A2(n374), .Y(n281) );
  MUX21X1_HVT U266 ( .A1(n304), .A2(n297), .S0(n312), .Y(n583) );
  MUX21X1_HVT U267 ( .A1(n306), .A2(n304), .S0(n310), .Y(n378) );
  AND2X1_HVT U268 ( .A1(n308), .A2(n482), .Y(n282) );
  XNOR2X1_HVT U269 ( .A1(n307), .A2(n309), .Y(n283) );
  MUX21X1_HVT U270 ( .A1(n301), .A2(n297), .S0(n309), .Y(n384) );
  MUX21X1_HVT U271 ( .A1(n302), .A2(n375), .S0(n309), .Y(n522) );
  MUX21X1_HVT U272 ( .A1(n302), .A2(n308), .S0(n290), .Y(n468) );
  XOR2X1_HVT U273 ( .A1(n237), .A2(n312), .Y(n569) );
  NBUFFX2_HVT U274 ( .A(in[7]), .Y(n296) );
  NBUFFX2_HVT U275 ( .A(in[7]), .Y(n294) );
  NBUFFX2_HVT U276 ( .A(in[7]), .Y(n295) );
  NBUFFX2_HVT U277 ( .A(n372), .Y(n297) );
  NBUFFX2_HVT U278 ( .A(in[2]), .Y(n288) );
  NBUFFX2_HVT U279 ( .A(in[5]), .Y(n293) );
  NBUFFX2_HVT U280 ( .A(in[2]), .Y(n290) );
  NBUFFX2_HVT U281 ( .A(in[2]), .Y(n289) );
  NBUFFX2_HVT U282 ( .A(in[5]), .Y(n292) );
  NBUFFX2_HVT U283 ( .A(in[2]), .Y(n287) );
  NBUFFX2_HVT U284 ( .A(in[5]), .Y(n291) );
  MUX21X1_HVT U285 ( .A1(n493), .A2(n343), .S0(n290), .Y(n490) );
  MUX21X1_HVT U286 ( .A1(n507), .A2(n299), .S0(n295), .Y(n411) );
  XOR2X1_HVT U287 ( .A1(n95), .A2(n299), .Y(n547) );
  MUX21X1_HVT U288 ( .A1(n301), .A2(n261), .S0(n309), .Y(n488) );
  MUX21X1_HVT U289 ( .A1(n423), .A2(n422), .S0(n290), .Y(n421) );
  MUX21X1_HVT U290 ( .A1(n302), .A2(n360), .S0(n296), .Y(n423) );
  AND2X1_HVT U291 ( .A1(n265), .A2(n314), .Y(n284) );
  MUX21X1_HVT U292 ( .A1(n299), .A2(n370), .S0(n96), .Y(n556) );
  MUX21X1_HVT U293 ( .A1(n442), .A2(n443), .S0(n287), .Y(n440) );
  MUX21X1_HVT U294 ( .A1(n362), .A2(n371), .S0(n295), .Y(n443) );
  MUX21X1_HVT U295 ( .A1(n551), .A2(n524), .S0(n289), .Y(n523) );
  MUX21X1_HVT U296 ( .A1(n373), .A2(n360), .S0(n296), .Y(n524) );
  MUX21X1_HVT U297 ( .A1(n371), .A2(n374), .S0(n311), .Y(n428) );
  NAND2X0_HVT U298 ( .A1(in[3]), .A2(n237), .Y(n593) );
  NBUFFX2_HVT U299 ( .A(n594), .Y(n307) );
  MUX21X1_HVT U300 ( .A1(n374), .A2(n299), .S0(n23), .Y(n575) );
  MUX21X1_HVT U301 ( .A1(n236), .A2(n592), .S0(n288), .Y(n485) );
  MUX21X1_HVT U302 ( .A1(n438), .A2(n306), .S0(n285), .Y(n437) );
  MUX21X1_HVT U303 ( .A1(n577), .A2(n344), .S0(n288), .Y(n460) );
  MUX21X1_HVT U304 ( .A1(n542), .A2(n543), .S0(n294), .Y(n540) );
  MUX21X1_HVT U305 ( .A1(n299), .A2(n560), .S0(n291), .Y(n543) );
  XOR2X1_HVT U306 ( .A1(n312), .A2(n293), .Y(n552) );
  MUX21X1_HVT U307 ( .A1(n592), .A2(n313), .S0(n289), .Y(n467) );
  NBUFFX2_HVT U308 ( .A(n585), .Y(n300) );
  MUX21X1_HVT U309 ( .A1(n299), .A2(n371), .S0(n312), .Y(n383) );
  MUX21X1_HVT U310 ( .A1(n304), .A2(n299), .S0(n310), .Y(n586) );
  MUX21X1_HVT U311 ( .A1(n331), .A2(n314), .S0(in[5]), .Y(n528) );
  NBUFFX2_HVT U312 ( .A(n585), .Y(n301) );
  MUX21X1_HVT U313 ( .A1(n341), .A2(n565), .S0(n288), .Y(n463) );
  MUX21X1_HVT U314 ( .A1(n351), .A2(n368), .S0(n295), .Y(n399) );
  MUX21X1_HVT U315 ( .A1(n299), .A2(n375), .S0(n296), .Y(n502) );
  NBUFFX2_HVT U316 ( .A(n594), .Y(n308) );
  NBUFFX2_HVT U317 ( .A(n585), .Y(n302) );
  XNOR2X1_HVT U318 ( .A1(n247), .A2(n96), .Y(n285) );
  AND2X1_HVT U319 ( .A1(n297), .A2(n314), .Y(n286) );
  MUX21X1_HVT U320 ( .A1(n399), .A2(n398), .S0(n289), .Y(n397) );
  INVX0_HVT U321 ( .A(in[4]), .Y(n375) );
  MUX21X1_HVT U322 ( .A1(n540), .A2(n544), .S0(n290), .Y(n539) );
  MUX21X1_HVT U323 ( .A1(n534), .A2(n536), .S0(n289), .Y(n533) );
  MUX21X1_HVT U324 ( .A1(n370), .A2(in[4]), .S0(n95), .Y(n563) );
  NAND2X0_HVT U325 ( .A1(in[3]), .A2(in[4]), .Y(n594) );
  MUX21X1_HVT U326 ( .A1(n255), .A2(n258), .S0(n311), .Y(n385) );
  MUX21X1_HVT U327 ( .A1(in[4]), .A2(n371), .S0(n309), .Y(n577) );
  NAND2X0_HVT U328 ( .A1(in[4]), .A2(n372), .Y(n585) );
  MUX21X1_HVT U329 ( .A1(in[4]), .A2(n306), .S0(n23), .Y(n574) );
  MUX21X1_HVT U330 ( .A1(n308), .A2(n255), .S0(n312), .Y(n567) );
  MUX21X1_HVT U331 ( .A1(n299), .A2(n255), .S0(n266), .Y(n480) );
  MUX21X1_HVT U332 ( .A1(in[4]), .A2(n301), .S0(n95), .Y(n377) );
  MUX21X1_HVT U333 ( .A1(n255), .A2(n308), .S0(n309), .Y(n376) );
  MUX21X1_HVT U334 ( .A1(n297), .A2(in[4]), .S0(n23), .Y(n565) );
  INVX0_HVT U335 ( .A(in[1]), .Y(n314) );
  NBUFFX2_HVT U336 ( .A(in[3]), .Y(n299) );
  NBUFFX2_HVT U337 ( .A(in[0]), .Y(n298) );
  INVX0_HVT U338 ( .A(n573), .Y(n318) );
  INVX0_HVT U339 ( .A(n571), .Y(n319) );
  INVX0_HVT U340 ( .A(n562), .Y(n320) );
  INVX0_HVT U341 ( .A(n560), .Y(n321) );
  INVX0_HVT U342 ( .A(n425), .Y(n322) );
  INVX0_HVT U343 ( .A(n388), .Y(n323) );
  INVX0_HVT U344 ( .A(n592), .Y(n324) );
  INVX0_HVT U345 ( .A(n579), .Y(n325) );
  INVX0_HVT U346 ( .A(n591), .Y(n326) );
  INVX0_HVT U347 ( .A(n589), .Y(n327) );
  INVX0_HVT U348 ( .A(n586), .Y(n329) );
  INVX0_HVT U349 ( .A(n584), .Y(n330) );
  INVX0_HVT U350 ( .A(n583), .Y(n331) );
  INVX0_HVT U351 ( .A(n578), .Y(n333) );
  INVX0_HVT U352 ( .A(n577), .Y(n334) );
  INVX0_HVT U353 ( .A(n576), .Y(n335) );
  INVX0_HVT U354 ( .A(n575), .Y(n336) );
  INVX0_HVT U355 ( .A(n574), .Y(n337) );
  INVX0_HVT U356 ( .A(n570), .Y(n339) );
  INVX0_HVT U357 ( .A(n569), .Y(n340) );
  INVX0_HVT U358 ( .A(n567), .Y(n341) );
  INVX0_HVT U359 ( .A(n565), .Y(n342) );
  INVX0_HVT U360 ( .A(n563), .Y(n344) );
  INVX0_HVT U361 ( .A(n561), .Y(n345) );
  INVX0_HVT U362 ( .A(n558), .Y(n346) );
  INVX0_HVT U363 ( .A(n557), .Y(n347) );
  INVX0_HVT U364 ( .A(n556), .Y(n348) );
  INVX0_HVT U365 ( .A(n555), .Y(n349) );
  INVX0_HVT U366 ( .A(n554), .Y(n350) );
  INVX0_HVT U367 ( .A(n553), .Y(n351) );
  INVX0_HVT U368 ( .A(n582), .Y(n353) );
  INVX0_HVT U369 ( .A(n387), .Y(n355) );
  INVX0_HVT U370 ( .A(n537), .Y(n356) );
  INVX0_HVT U371 ( .A(n441), .Y(n357) );
  INVX0_HVT U372 ( .A(n386), .Y(n358) );
  INVX0_HVT U373 ( .A(n385), .Y(n359) );
  INVX0_HVT U374 ( .A(n384), .Y(n360) );
  INVX0_HVT U375 ( .A(n383), .Y(n361) );
  INVX0_HVT U376 ( .A(n382), .Y(n362) );
  INVX0_HVT U377 ( .A(n501), .Y(n363) );
  INVX0_HVT U378 ( .A(n491), .Y(n364) );
  INVX0_HVT U379 ( .A(n380), .Y(n365) );
  INVX0_HVT U380 ( .A(n379), .Y(n366) );
  INVX0_HVT U381 ( .A(n378), .Y(n367) );
  INVX0_HVT U382 ( .A(n377), .Y(n368) );
  INVX0_HVT U383 ( .A(n376), .Y(n369) );
endmodule

