
module inv_sbox_15 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n196, n197, n198, n199, n200, n201, n202, n203, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670;

  NAND2X0_HVT U4 ( .A1(n388), .A2(n253), .Y(n667) );
  NAND2X0_HVT U5 ( .A1(n667), .A2(n380), .Y(n666) );
  NAND2X0_HVT U7 ( .A1(n272), .A2(n381), .Y(n663) );
  NAND2X0_HVT U8 ( .A1(n272), .A2(n379), .Y(n662) );
  NAND2X0_HVT U9 ( .A1(n384), .A2(n662), .Y(n661) );
  NAND2X0_HVT U10 ( .A1(n384), .A2(n659), .Y(n660) );
  NAND2X0_HVT U11 ( .A1(n391), .A2(n248), .Y(n658) );
  NAND2X0_HVT U12 ( .A1(n389), .A2(n457), .Y(n657) );
  NAND2X0_HVT U13 ( .A1(n382), .A2(n662), .Y(n656) );
  NAND2X0_HVT U15 ( .A1(n377), .A2(n389), .Y(n654) );
  NAND2X0_HVT U19 ( .A1(n388), .A2(n459), .Y(n649) );
  NAND2X0_HVT U25 ( .A1(n356), .A2(n370), .Y(n665) );
  NAND2X0_HVT U32 ( .A1(n371), .A2(n301), .Y(n637) );
  NAND2X0_HVT U35 ( .A1(n220), .A2(n460), .Y(n634) );
  NAND2X0_HVT U38 ( .A1(n370), .A2(n391), .Y(n631) );
  NAND2X0_HVT U42 ( .A1(n664), .A2(n460), .Y(n627) );
  NAND2X0_HVT U55 ( .A1(n382), .A2(n667), .Y(n615) );
  MUX41X1_HVT U56 ( .A1(n227), .A3(n378), .A2(n424), .A4(n615), .S0(n364), 
        .S1(n395), .Y(n614) );
  MUX41X1_HVT U65 ( .A1(n418), .A3(n420), .A2(n419), .A4(n631), .S0(n364), 
        .S1(n396), .Y(n604) );
  NAND2X0_HVT U66 ( .A1(n385), .A2(n356), .Y(n603) );
  MUX41X1_HVT U67 ( .A1(n415), .A3(n440), .A2(n417), .A4(n603), .S0(n221), 
        .S1(n361), .Y(n602) );
  MUX41X1_HVT U68 ( .A1(n415), .A3(n346), .A2(n416), .A4(n383), .S0(n363), 
        .S1(n311), .Y(n601) );
  NAND2X0_HVT U72 ( .A1(n378), .A2(n663), .Y(n598) );
  MUX41X1_HVT U73 ( .A1(n642), .A3(n598), .A2(n441), .A4(n369), .S0(n221), 
        .S1(n360), .Y(n597) );
  MUX41X1_HVT U74 ( .A1(n660), .A3(n431), .A2(n430), .A4(n421), .S0(n364), 
        .S1(n298), .Y(n596) );
  MUX41X1_HVT U78 ( .A1(n593), .A3(n597), .A2(n596), .A4(n599), .S0(n376), 
        .S1(n374), .Y(n592) );
  MUX41X1_HVT U80 ( .A1(n443), .A3(n227), .A2(n219), .A4(n666), .S0(n363), 
        .S1(n396), .Y(n590) );
  NAND2X0_HVT U81 ( .A1(n253), .A2(n663), .Y(n589) );
  AND2X1_HVT U82 ( .A1(n664), .A2(n668), .Y(n588) );
  MUX41X1_HVT U83 ( .A1(n588), .A3(n428), .A2(n444), .A4(n589), .S0(n363), 
        .S1(n298), .Y(n587) );
  MUX41X1_HVT U84 ( .A1(n354), .A3(n427), .A2(n445), .A4(n644), .S0(n364), 
        .S1(n396), .Y(n586) );
  MUX41X1_HVT U85 ( .A1(n586), .A3(n590), .A2(n587), .A4(n591), .S0(n376), 
        .S1(in[1]), .Y(n585) );
  MUX41X1_HVT U88 ( .A1(n417), .A3(n402), .A2(n639), .A4(n623), .S0(n363), 
        .S1(n343), .Y(n583) );
  NAND2X0_HVT U89 ( .A1(n301), .A2(n456), .Y(n582) );
  MUX41X1_HVT U90 ( .A1(n345), .A3(n663), .A2(n622), .A4(n582), .S0(n363), 
        .S1(n395), .Y(n581) );
  MUX41X1_HVT U96 ( .A1(n440), .A3(n656), .A2(n425), .A4(n447), .S0(n364), 
        .S1(n396), .Y(n575) );
  MUX41X1_HVT U99 ( .A1(n637), .A3(n419), .A2(n621), .A4(n377), .S0(n396), 
        .S1(n361), .Y(n572) );
  NAND2X0_HVT U100 ( .A1(n301), .A2(n243), .Y(n571) );
  MUX41X1_HVT U101 ( .A1(n449), .A3(n657), .A2(n432), .A4(n571), .S0(n311), 
        .S1(n359), .Y(n570) );
  MUX41X1_HVT U102 ( .A1(n570), .A3(n573), .A2(n572), .A4(n575), .S0(n376), 
        .S1(n374), .Y(n569) );
  AND2X1_HVT U104 ( .A1(n663), .A2(n380), .Y(n568) );
  MUX41X1_HVT U105 ( .A1(n655), .A3(n450), .A2(n589), .A4(n568), .S0(n364), 
        .S1(n312), .Y(n567) );
  MUX41X1_HVT U107 ( .A1(n449), .A3(n381), .A2(n566), .A4(n408), .S0(n363), 
        .S1(n395), .Y(n565) );
  MUX41X1_HVT U108 ( .A1(n421), .A3(n378), .A2(n424), .A4(n249), .S0(n364), 
        .S1(n310), .Y(n564) );
  MUX41X1_HVT U109 ( .A1(n448), .A3(n402), .A2(n445), .A4(n438), .S0(n363), 
        .S1(n395), .Y(n563) );
  AO21X1_HVT U112 ( .A1(n435), .A2(n368), .A3(n645), .Y(n560) );
  NAND2X0_HVT U114 ( .A1(n384), .A2(n663), .Y(n558) );
  MUX41X1_HVT U115 ( .A1(n558), .A3(n658), .A2(n435), .A4(n382), .S0(n396), 
        .S1(n361), .Y(n557) );
  MUX41X1_HVT U116 ( .A1(n434), .A3(n427), .A2(n402), .A4(n654), .S0(n362), 
        .S1(n310), .Y(n556) );
  NAND2X0_HVT U118 ( .A1(n301), .A2(n346), .Y(n554) );
  MUX41X1_HVT U120 ( .A1(n553), .A3(n557), .A2(n556), .A4(n559), .S0(n376), 
        .S1(n295), .Y(n552) );
  MUX41X1_HVT U122 ( .A1(n439), .A3(n350), .A2(n623), .A4(n442), .S0(n362), 
        .S1(n343), .Y(n551) );
  MUX41X1_HVT U124 ( .A1(n352), .A3(n550), .A2(n646), .A4(n270), .S0(n394), 
        .S1(n362), .Y(n549) );
  AOI21X1_HVT U127 ( .A1(n367), .A2(n545), .A3(n409), .Y(n546) );
  NAND2X0_HVT U129 ( .A1(n366), .A2(n383), .Y(n543) );
  MUX41X1_HVT U130 ( .A1(n543), .A3(n544), .A2(n547), .A4(n546), .S0(n221), 
        .S1(n305), .Y(n542) );
  AND2X1_HVT U131 ( .A1(n356), .A2(n301), .Y(n541) );
  MUX41X1_HVT U132 ( .A1(n406), .A3(n541), .A2(n453), .A4(n415), .S0(n221), 
        .S1(n360), .Y(n540) );
  MUX41X1_HVT U133 ( .A1(n454), .A3(n408), .A2(n615), .A4(n407), .S0(n310), 
        .S1(n359), .Y(n539) );
  MUX41X1_HVT U136 ( .A1(n620), .A3(n571), .A2(n537), .A4(n413), .S0(n366), 
        .S1(n343), .Y(n536) );
  MUX41X1_HVT U137 ( .A1(n220), .A3(n640), .A2(n644), .A4(n447), .S0(n394), 
        .S1(n359), .Y(n535) );
  MUX41X1_HVT U140 ( .A1(n430), .A3(n351), .A2(n423), .A4(n658), .S0(n221), 
        .S1(n361), .Y(n533) );
  NAND2X0_HVT U141 ( .A1(n377), .A2(n301), .Y(n532) );
  MUX41X1_HVT U142 ( .A1(n532), .A3(n630), .A2(n452), .A4(n423), .S0(n367), 
        .S1(n396), .Y(n531) );
  MUX41X1_HVT U145 ( .A1(n638), .A3(n450), .A2(n529), .A4(n589), .S0(n367), 
        .S1(n312), .Y(n528) );
  MUX41X1_HVT U146 ( .A1(n528), .A3(n530), .A2(n531), .A4(n533), .S0(n374), 
        .S1(n376), .Y(n527) );
  OA21X1_HVT U153 ( .A1(n403), .A2(n398), .A3(n412), .Y(n520) );
  MUX41X1_HVT U155 ( .A1(n423), .A3(n658), .A2(n650), .A4(n425), .S0(n365), 
        .S1(n395), .Y(n518) );
  MUX41X1_HVT U156 ( .A1(n518), .A3(n522), .A2(n519), .A4(n524), .S0(in[5]), 
        .S1(n281), .Y(n517) );
  NAND2X0_HVT U159 ( .A1(n514), .A2(n513), .Y(n515) );
  NAND2X0_HVT U163 ( .A1(n387), .A2(n456), .Y(n509) );
  NAND2X0_HVT U166 ( .A1(n505), .A2(n659), .Y(n506) );
  MUX41X1_HVT U174 ( .A1(n446), .A3(n615), .A2(n454), .A4(n460), .S0(n365), 
        .S1(n311), .Y(n497) );
  NAND2X0_HVT U177 ( .A1(n388), .A2(n346), .Y(n495) );
  MUX41X1_HVT U178 ( .A1(n353), .A3(n495), .A2(n345), .A4(n625), .S0(n365), 
        .S1(n395), .Y(n494) );
  AND2X1_HVT U179 ( .A1(n664), .A2(n379), .Y(n493) );
  MUX41X1_HVT U183 ( .A1(n436), .A3(n227), .A2(n421), .A4(n627), .S0(n311), 
        .S1(n360), .Y(n489) );
  AND2X1_HVT U185 ( .A1(n460), .A2(n301), .Y(n487) );
  OA21X1_HVT U189 ( .A1(n427), .A2(n398), .A3(n609), .Y(n483) );
  NAND2X0_HVT U191 ( .A1(n304), .A2(n414), .Y(n481) );
  AND2X1_HVT U192 ( .A1(n431), .A2(n479), .Y(n480) );
  NAND2X0_HVT U194 ( .A1(n627), .A2(n479), .Y(n477) );
  NAND2X0_HVT U198 ( .A1(n386), .A2(n460), .Y(n659) );
  NAND2X0_HVT U200 ( .A1(n379), .A2(n301), .Y(n545) );
  AO21X1_HVT U204 ( .A1(n378), .A2(n299), .A3(n398), .Y(n505) );
  NAND2X0_HVT U207 ( .A1(n301), .A2(n345), .Y(n609) );
  INVX0_HVT U1 ( .A(in[3]), .Y(n196) );
  INVX0_HVT U2 ( .A(n196), .Y(n197) );
  MUX41X1_HVT U3 ( .A1(n509), .A3(n661), .A2(n421), .A4(n632), .S0(n198), .S1(
        n312), .Y(n508) );
  IBUFFX16_HVT U6 ( .A(n362), .Y(n198) );
  AO21X2_HVT U14 ( .A1(n609), .A2(n394), .A3(n648), .Y(n610) );
  NBUFFX2_HVT U16 ( .A(n461), .Y(n372) );
  MUX21X2_HVT U17 ( .A1(n354), .A2(n621), .S0(n368), .Y(n485) );
  MUX21X2_HVT U18 ( .A1(n506), .A2(n507), .S0(n366), .Y(n504) );
  MUX21X2_HVT U20 ( .A1(n346), .A2(n243), .S0(n267), .Y(n646) );
  INVX0_HVT U21 ( .A(n387), .Y(n267) );
  MUX41X1_HVT U22 ( .A1(n511), .A3(n420), .A2(n634), .A4(n347), .S0(n199), 
        .S1(n200), .Y(n510) );
  IBUFFX16_HVT U23 ( .A(n396), .Y(n199) );
  IBUFFX16_HVT U24 ( .A(n365), .Y(n200) );
  INVX0_HVT U26 ( .A(n646), .Y(n422) );
  OA21X1_HVT U27 ( .A1(n398), .A2(n619), .A3(n426), .Y(n617) );
  INVX1_HVT U28 ( .A(n380), .Y(n456) );
  MUX21X1_HVT U29 ( .A1(n241), .A2(n653), .S0(n202), .Y(n201) );
  IBUFFX16_HVT U30 ( .A(n201), .Y(n647) );
  IBUFFX16_HVT U31 ( .A(n338), .Y(n202) );
  IBUFFX2_HVT U33 ( .A(n241), .Y(n244) );
  INVX0_HVT U34 ( .A(n653), .Y(n460) );
  IBUFFX2_HVT U36 ( .A(n633), .Y(n432) );
  MUX21X2_HVT U37 ( .A1(n633), .A2(n249), .S0(n336), .Y(n340) );
  XOR2X2_HVT U39 ( .A1(n379), .A2(n386), .Y(n621) );
  MUX41X1_HVT U40 ( .A1(n548), .A3(n542), .A2(n538), .A4(n534), .S0(n203), 
        .S1(n218), .Y(out[4]) );
  IBUFFX16_HVT U41 ( .A(n376), .Y(n203) );
  IBUFFX16_HVT U43 ( .A(n344), .Y(n218) );
  INVX1_HVT U44 ( .A(in[1]), .Y(n373) );
  IBUFFX2_HVT U45 ( .A(n373), .Y(n305) );
  MUX21X2_HVT U46 ( .A1(n339), .A2(n340), .S0(n312), .Y(n498) );
  INVX0_HVT U47 ( .A(n413), .Y(n219) );
  INVX1_HVT U48 ( .A(n410), .Y(n220) );
  INVX1_HVT U49 ( .A(n661), .Y(n413) );
  INVX0_HVT U50 ( .A(n662), .Y(n410) );
  NBUFFX2_HVT U51 ( .A(n368), .Y(n221) );
  NBUFFX2_HVT U52 ( .A(n397), .Y(n368) );
  MUX41X1_HVT U53 ( .A1(n510), .A3(n512), .A2(n504), .A4(n508), .S0(n281), 
        .S1(n375), .Y(n503) );
  IBUFFX2_HVT U54 ( .A(n376), .Y(n306) );
  MUX21X1_HVT U57 ( .A1(n461), .A2(n380), .S0(n234), .Y(n227) );
  INVX1_HVT U58 ( .A(n257), .Y(n234) );
  IBUFFX2_HVT U59 ( .A(n385), .Y(n257) );
  INVX1_HVT U60 ( .A(n390), .Y(n385) );
  INVX1_HVT U61 ( .A(n222), .Y(n580) );
  MUX21X1_HVT U62 ( .A1(n371), .A2(n456), .S0(n272), .Y(n523) );
  MUX21X1_HVT U63 ( .A1(n223), .A2(n224), .S0(n221), .Y(n222) );
  IBUFFX16_HVT U64 ( .A(n377), .Y(n223) );
  IBUFFX16_HVT U69 ( .A(n371), .Y(n224) );
  MUX41X1_HVT U70 ( .A1(n614), .A3(n616), .A2(n608), .A4(n612), .S0(n295), 
        .S1(n306), .Y(n607) );
  MUX21X1_HVT U71 ( .A1(n381), .A2(n379), .S0(n225), .Y(n511) );
  IBUFFX2_HVT U75 ( .A(n399), .Y(n396) );
  NBUFFX4_HVT U76 ( .A(n457), .Y(n370) );
  MUX21X2_HVT U77 ( .A1(n569), .A2(n576), .S0(n344), .Y(out[2]) );
  IBUFFX16_HVT U79 ( .A(n385), .Y(n225) );
  MUX41X1_HVT U86 ( .A1(n582), .A3(n500), .A2(n349), .A4(n647), .S0(n226), 
        .S1(n311), .Y(n499) );
  IBUFFX16_HVT U87 ( .A(n337), .Y(n226) );
  INVX0_HVT U91 ( .A(n374), .Y(n228) );
  INVX0_HVT U92 ( .A(n373), .Y(n374) );
  INVX1_HVT U93 ( .A(n461), .Y(n356) );
  MUX41X1_HVT U94 ( .A1(n485), .A3(n484), .A2(n486), .A4(n483), .S0(n228), 
        .S1(n229), .Y(n482) );
  IBUFFX16_HVT U95 ( .A(n336), .Y(n229) );
  NAND2X0_HVT U97 ( .A1(n316), .A2(n230), .Y(n231) );
  NAND2X0_HVT U98 ( .A1(n317), .A2(n343), .Y(n232) );
  NAND2X0_HVT U103 ( .A1(n231), .A2(n232), .Y(n573) );
  IBUFFX2_HVT U106 ( .A(n343), .Y(n230) );
  MUX21X1_HVT U110 ( .A1(n456), .A2(n458), .S0(n233), .Y(n641) );
  IBUFFX16_HVT U111 ( .A(n386), .Y(n233) );
  MUX41X1_HVT U113 ( .A1(n482), .A3(n476), .A2(n491), .A4(n488), .S0(n303), 
        .S1(n237), .Y(out[7]) );
  INVX1_HVT U117 ( .A(n302), .Y(n237) );
  IBUFFX2_HVT U119 ( .A(in[5]), .Y(n303) );
  MUX41X1_HVT U121 ( .A1(n523), .A3(n201), .A2(n433), .A4(n444), .S0(n235), 
        .S1(n236), .Y(n522) );
  IBUFFX16_HVT U123 ( .A(n312), .Y(n235) );
  IBUFFX16_HVT U125 ( .A(n359), .Y(n236) );
  OR2X1_HVT U126 ( .A1(n457), .A2(n238), .Y(n668) );
  IBUFFX16_HVT U128 ( .A(in[6]), .Y(n238) );
  IBUFFX2_HVT U134 ( .A(n457), .Y(n346) );
  INVX1_HVT U135 ( .A(in[6]), .Y(n461) );
  NBUFFX2_HVT U138 ( .A(n669), .Y(n239) );
  INVX1_HVT U139 ( .A(n455), .Y(n240) );
  INVX1_HVT U143 ( .A(n455), .Y(n241) );
  INVX1_HVT U144 ( .A(n455), .Y(n242) );
  INVX1_HVT U147 ( .A(n240), .Y(n243) );
  INVX1_HVT U148 ( .A(n242), .Y(n245) );
  IBUFFX2_HVT U149 ( .A(n669), .Y(n246) );
  IBUFFX2_HVT U150 ( .A(n669), .Y(n247) );
  INVX1_HVT U151 ( .A(n246), .Y(n248) );
  INVX1_HVT U152 ( .A(n247), .Y(n249) );
  INVX1_HVT U154 ( .A(n239), .Y(n250) );
  INVX1_HVT U157 ( .A(n239), .Y(n251) );
  INVX1_HVT U158 ( .A(n250), .Y(n252) );
  INVX1_HVT U160 ( .A(n251), .Y(n253) );
  NAND2X0_HVT U161 ( .A1(n369), .A2(n372), .Y(n669) );
  INVX0_HVT U162 ( .A(n669), .Y(n455) );
  MUX41X1_HVT U164 ( .A1(n424), .A3(n446), .A2(n354), .A4(n405), .S0(n337), 
        .S1(n304), .Y(n584) );
  INVX1_HVT U165 ( .A(n405), .Y(n299) );
  MUX21X1_HVT U167 ( .A1(n422), .A2(n615), .S0(n368), .Y(n611) );
  NAND2X0_HVT U168 ( .A1(n490), .A2(n254), .Y(n255) );
  NAND2X0_HVT U169 ( .A1(n489), .A2(n373), .Y(n256) );
  NAND2X0_HVT U170 ( .A1(n255), .A2(n256), .Y(n488) );
  IBUFFX2_HVT U171 ( .A(n373), .Y(n254) );
  IBUFFX2_HVT U172 ( .A(n373), .Y(n281) );
  MUX21X2_HVT U173 ( .A1(n628), .A2(n441), .S0(n321), .Y(n484) );
  MUX21X2_HVT U175 ( .A1(n459), .A2(n356), .S0(n296), .Y(n628) );
  NAND2X0_HVT U176 ( .A1(n562), .A2(n258), .Y(n259) );
  NAND2X0_HVT U180 ( .A1(n552), .A2(n269), .Y(n260) );
  NAND2X0_HVT U181 ( .A1(n259), .A2(n260), .Y(out[3]) );
  INVX1_HVT U182 ( .A(n269), .Y(n258) );
  IBUFFX2_HVT U184 ( .A(n344), .Y(n269) );
  NAND2X0_HVT U186 ( .A1(n578), .A2(n261), .Y(n262) );
  NAND2X0_HVT U187 ( .A1(n579), .A2(n366), .Y(n263) );
  NAND2X0_HVT U188 ( .A1(n262), .A2(n263), .Y(n577) );
  IBUFFX2_HVT U190 ( .A(n366), .Y(n261) );
  NAND2X1_HVT U193 ( .A1(n600), .A2(n264), .Y(n265) );
  NAND2X0_HVT U195 ( .A1(n607), .A2(n344), .Y(n266) );
  NAND2X0_HVT U196 ( .A1(n266), .A2(n265), .Y(out[0]) );
  IBUFFX2_HVT U197 ( .A(n344), .Y(n264) );
  MUX41X1_HVT U199 ( .A1(n577), .A3(n581), .A2(n583), .A4(n584), .S0(n295), 
        .S1(n376), .Y(n576) );
  IBUFFX2_HVT U201 ( .A(n664), .Y(n407) );
  INVX0_HVT U202 ( .A(n632), .Y(n433) );
  MUX21X2_HVT U203 ( .A1(n610), .A2(n611), .S0(n268), .Y(n608) );
  IBUFFX16_HVT U205 ( .A(n366), .Y(n268) );
  INVX0_HVT U206 ( .A(n667), .Y(n405) );
  NBUFFX2_HVT U208 ( .A(n422), .Y(n270) );
  IBUFFX2_HVT U209 ( .A(n390), .Y(n271) );
  IBUFFX2_HVT U210 ( .A(n390), .Y(n272) );
  IBUFFX2_HVT U211 ( .A(n373), .Y(n295) );
  NAND2X0_HVT U212 ( .A1(n525), .A2(n273), .Y(n274) );
  NAND2X0_HVT U213 ( .A1(n526), .A2(n300), .Y(n275) );
  NAND2X0_HVT U214 ( .A1(n274), .A2(n275), .Y(n524) );
  INVX0_HVT U215 ( .A(n300), .Y(n273) );
  AO21X2_HVT U216 ( .A1(n368), .A2(n410), .A3(n244), .Y(n525) );
  MUX21X1_HVT U217 ( .A1(n453), .A2(n406), .S0(n394), .Y(n526) );
  IBUFFX2_HVT U218 ( .A(n366), .Y(n300) );
  INVX0_HVT U219 ( .A(n637), .Y(n401) );
  INVX1_HVT U220 ( .A(n668), .Y(n459) );
  MUX41X1_HVT U221 ( .A1(n637), .A3(n493), .A2(n400), .A4(n624), .S0(n396), 
        .S1(n365), .Y(n492) );
  NAND2X0_HVT U222 ( .A1(n494), .A2(n276), .Y(n277) );
  NAND2X0_HVT U223 ( .A1(n492), .A2(n285), .Y(n278) );
  NAND2X0_HVT U224 ( .A1(n277), .A2(n278), .Y(n491) );
  INVX0_HVT U225 ( .A(n285), .Y(n276) );
  IBUFFX2_HVT U226 ( .A(n658), .Y(n400) );
  INVX1_HVT U227 ( .A(n305), .Y(n285) );
  MUX41X1_HVT U228 ( .A1(n632), .A3(n554), .A2(n451), .A4(n555), .S0(n279), 
        .S1(n280), .Y(n553) );
  IBUFFX16_HVT U229 ( .A(n337), .Y(n279) );
  IBUFFX16_HVT U230 ( .A(n395), .Y(n280) );
  IBUFFX16_HVT U231 ( .A(n390), .Y(n388) );
  XOR2X2_HVT U232 ( .A1(n377), .A2(n271), .Y(n623) );
  MUX41X1_HVT U233 ( .A1(n646), .A3(n649), .A2(n436), .A4(n456), .S0(n282), 
        .S1(n283), .Y(n530) );
  IBUFFX16_HVT U234 ( .A(n365), .Y(n282) );
  IBUFFX16_HVT U235 ( .A(n395), .Y(n283) );
  MUX41X1_HVT U236 ( .A1(n498), .A3(n497), .A2(n501), .A4(n499), .S0(n373), 
        .S1(n284), .Y(n496) );
  IBUFFX16_HVT U237 ( .A(n375), .Y(n284) );
  NAND2X0_HVT U238 ( .A1(n641), .A2(n286), .Y(n287) );
  NAND2X0_HVT U239 ( .A1(n433), .A2(n318), .Y(n288) );
  NAND2X0_HVT U240 ( .A1(n287), .A2(n288), .Y(n317) );
  IBUFFX2_HVT U241 ( .A(n318), .Y(n286) );
  INVX0_HVT U242 ( .A(n364), .Y(n318) );
  NAND2X0_HVT U243 ( .A1(n520), .A2(n289), .Y(n290) );
  NAND2X0_HVT U244 ( .A1(n521), .A2(n367), .Y(n291) );
  NAND2X0_HVT U245 ( .A1(n290), .A2(n291), .Y(n519) );
  IBUFFX2_HVT U246 ( .A(n367), .Y(n289) );
  MUX21X1_HVT U247 ( .A1(n644), .A2(n354), .S0(n368), .Y(n521) );
  INVX0_HVT U248 ( .A(n644), .Y(n423) );
  MUX21X1_HVT U249 ( .A1(n371), .A2(n378), .S0(n391), .Y(n644) );
  INVX2_HVT U250 ( .A(n385), .Y(n296) );
  AO21X2_HVT U251 ( .A1(n388), .A2(n245), .A3(n398), .Y(n479) );
  INVX1_HVT U252 ( .A(n386), .Y(n391) );
  INVX2_HVT U253 ( .A(in[0]), .Y(n390) );
  NAND2X0_HVT U254 ( .A1(n381), .A2(n292), .Y(n293) );
  NAND2X0_HVT U255 ( .A1(n580), .A2(n296), .Y(n294) );
  NAND2X0_HVT U256 ( .A1(n294), .A2(n293), .Y(n579) );
  INVX1_HVT U257 ( .A(n296), .Y(n292) );
  IBUFFX2_HVT U258 ( .A(n397), .Y(n304) );
  IBUFFX2_HVT U259 ( .A(n397), .Y(n398) );
  INVX1_HVT U260 ( .A(n399), .Y(n397) );
  IBUFFX2_HVT U261 ( .A(n348), .Y(n297) );
  IBUFFX2_HVT U262 ( .A(n670), .Y(n345) );
  MUX41X1_HVT U263 ( .A1(n408), .A3(n405), .A2(n299), .A4(n444), .S0(n396), 
        .S1(n362), .Y(n490) );
  INVX1_HVT U264 ( .A(n471), .Y(n444) );
  INVX0_HVT U265 ( .A(n304), .Y(n298) );
  IBUFFX2_HVT U266 ( .A(n399), .Y(n395) );
  INVX1_HVT U267 ( .A(n390), .Y(n338) );
  INVX1_HVT U268 ( .A(n338), .Y(n301) );
  IBUFFX16_HVT U269 ( .A(n344), .Y(n302) );
  INVX0_HVT U270 ( .A(n355), .Y(n313) );
  MUX41X1_HVT U271 ( .A1(n480), .A3(n478), .A2(n481), .A4(n477), .S0(n373), 
        .S1(n363), .Y(n476) );
  NAND2X0_HVT U272 ( .A1(n324), .A2(n307), .Y(n308) );
  NAND2X0_HVT U273 ( .A1(n613), .A2(n355), .Y(n309) );
  NAND2X0_HVT U274 ( .A1(n308), .A2(n309), .Y(n612) );
  INVX0_HVT U275 ( .A(n355), .Y(n307) );
  XNOR2X1_HVT U276 ( .A1(n398), .A2(n362), .Y(n355) );
  NBUFFX2_HVT U277 ( .A(n394), .Y(n310) );
  NBUFFX2_HVT U278 ( .A(n394), .Y(n311) );
  NBUFFX2_HVT U279 ( .A(n394), .Y(n312) );
  IBUFFX2_HVT U280 ( .A(n399), .Y(n394) );
  INVX0_HVT U281 ( .A(n324), .Y(n645) );
  MUX21X1_HVT U282 ( .A1(n425), .A2(n416), .S0(n368), .Y(n618) );
  INVX1_HVT U283 ( .A(n363), .Y(n337) );
  INVX1_HVT U284 ( .A(n360), .Y(n336) );
  INVX1_HVT U285 ( .A(in[3]), .Y(n457) );
  INVX0_HVT U286 ( .A(n344), .Y(n329) );
  INVX1_HVT U287 ( .A(n375), .Y(n376) );
  INVX1_HVT U288 ( .A(in[5]), .Y(n375) );
  INVX1_HVT U289 ( .A(n394), .Y(n321) );
  NAND2X0_HVT U290 ( .A1(n421), .A2(n313), .Y(n314) );
  NAND2X0_HVT U291 ( .A1(n606), .A2(n355), .Y(n315) );
  NAND2X0_HVT U292 ( .A1(n314), .A2(n315), .Y(n605) );
  MUX21X1_HVT U293 ( .A1(n201), .A2(n299), .S0(n366), .Y(n606) );
  MUX21X1_HVT U294 ( .A1(n448), .A2(n574), .S0(n318), .Y(n316) );
  NAND2X0_HVT U295 ( .A1(n549), .A2(n373), .Y(n319) );
  NAND2X0_HVT U296 ( .A1(n551), .A2(n305), .Y(n320) );
  NAND2X0_HVT U297 ( .A1(n319), .A2(n320), .Y(n548) );
  INVX1_HVT U298 ( .A(n390), .Y(n386) );
  MUX41X1_HVT U299 ( .A1(n567), .A3(n564), .A2(n565), .A4(n563), .S0(n375), 
        .S1(n373), .Y(n562) );
  OA21X2_HVT U300 ( .A1(n404), .A2(n304), .A3(n648), .Y(n594) );
  NAND2X0_HVT U301 ( .A1(n409), .A2(n321), .Y(n322) );
  NAND2X0_HVT U302 ( .A1(n628), .A2(n394), .Y(n323) );
  NAND2X0_HVT U303 ( .A1(n322), .A2(n323), .Y(n561) );
  MUX21X2_HVT U304 ( .A1(n561), .A2(n560), .S0(n336), .Y(n559) );
  INVX1_HVT U305 ( .A(n474), .Y(n441) );
  MUX21X2_HVT U306 ( .A1(n617), .A2(n618), .S0(n337), .Y(n616) );
  MUX41X1_HVT U307 ( .A1(n605), .A3(n602), .A2(n604), .A4(n601), .S0(n375), 
        .S1(n373), .Y(n600) );
  MUX21X1_HVT U308 ( .A1(n297), .A2(n383), .S0(n387), .Y(n324) );
  NAND2X0_HVT U309 ( .A1(n487), .A2(n321), .Y(n325) );
  NAND2X0_HVT U310 ( .A1(n443), .A2(n311), .Y(n326) );
  NAND2X0_HVT U311 ( .A1(n325), .A2(n326), .Y(n486) );
  NAND2X0_HVT U312 ( .A1(n594), .A2(n365), .Y(n327) );
  NAND2X0_HVT U313 ( .A1(n595), .A2(n318), .Y(n328) );
  NAND2X0_HVT U314 ( .A1(n327), .A2(n328), .Y(n593) );
  NAND2X0_HVT U315 ( .A1(n585), .A2(n329), .Y(n330) );
  NAND2X0_HVT U316 ( .A1(n592), .A2(n344), .Y(n331) );
  NAND2X0_HVT U317 ( .A1(n330), .A2(n331), .Y(out[1]) );
  MUX21X1_HVT U318 ( .A1(n442), .A2(n401), .S0(n394), .Y(n595) );
  NBUFFX2_HVT U319 ( .A(in[7]), .Y(n344) );
  INVX1_HVT U320 ( .A(n648), .Y(n421) );
  NAND2X0_HVT U321 ( .A1(n517), .A2(n329), .Y(n332) );
  NAND2X0_HVT U322 ( .A1(n527), .A2(n344), .Y(n333) );
  NAND2X0_HVT U323 ( .A1(n332), .A2(n333), .Y(out[5]) );
  INVX1_HVT U324 ( .A(n642), .Y(n425) );
  NAND2X0_HVT U325 ( .A1(n496), .A2(n329), .Y(n334) );
  NAND2X0_HVT U326 ( .A1(n503), .A2(in[7]), .Y(n335) );
  NAND2X0_HVT U327 ( .A1(n335), .A2(n334), .Y(out[6]) );
  MUX41X1_HVT U328 ( .A1(n411), .A3(n658), .A2(n345), .A4(n664), .S0(n337), 
        .S1(n304), .Y(n599) );
  MUX21X1_HVT U329 ( .A1(n345), .A2(n383), .S0(n336), .Y(n339) );
  NAND2X0_HVT U330 ( .A1(n515), .A2(n318), .Y(n341) );
  NAND2X0_HVT U331 ( .A1(n516), .A2(n367), .Y(n342) );
  NAND2X0_HVT U332 ( .A1(n342), .A2(n341), .Y(n512) );
  MUX21X1_HVT U333 ( .A1(n626), .A2(n442), .S0(n368), .Y(n516) );
  INVX1_HVT U334 ( .A(n473), .Y(n442) );
  INVX1_HVT U335 ( .A(in[4]), .Y(n399) );
  AO21X2_HVT U336 ( .A1(n301), .A2(n383), .A3(n398), .Y(n513) );
  IBUFFX2_HVT U337 ( .A(n390), .Y(n389) );
  INVX1_HVT U338 ( .A(n472), .Y(n443) );
  INVX0_HVT U339 ( .A(n372), .Y(n348) );
  NAND2X0_HVT U340 ( .A1(n386), .A2(n384), .Y(n664) );
  INVX0_HVT U341 ( .A(n347), .Y(n625) );
  MUX21X1_HVT U342 ( .A1(n458), .A2(n459), .S0(n387), .Y(n502) );
  NBUFFX2_HVT U343 ( .A(n310), .Y(n343) );
  MUX41X1_HVT U344 ( .A1(n652), .A3(n429), .A2(n651), .A4(n427), .S0(n336), 
        .S1(n304), .Y(n591) );
  INVX0_HVT U345 ( .A(n383), .Y(n458) );
  NBUFFX2_HVT U346 ( .A(n670), .Y(n384) );
  MUX41X1_HVT U347 ( .A1(n502), .A3(n352), .A2(n349), .A4(n353), .S0(n336), 
        .S1(n304), .Y(n501) );
  MUX21X1_HVT U348 ( .A1(n384), .A2(n380), .S0(n391), .Y(n347) );
  IBUFFX2_HVT U349 ( .A(n390), .Y(n387) );
  OR2X1_HVT U350 ( .A1(n457), .A2(n348), .Y(n670) );
  NBUFFX2_HVT U351 ( .A(n665), .Y(n379) );
  NBUFFX2_HVT U352 ( .A(n665), .Y(n380) );
  AND2X1_HVT U353 ( .A1(n664), .A2(n248), .Y(n349) );
  MUX21X1_HVT U354 ( .A1(n437), .A2(n352), .S0(n310), .Y(n478) );
  AND2X1_HVT U355 ( .A1(n248), .A2(n654), .Y(n350) );
  MUX21X1_HVT U356 ( .A1(n458), .A2(n371), .S0(n387), .Y(n500) );
  MUX21X1_HVT U357 ( .A1(n372), .A2(n460), .S0(n272), .Y(n633) );
  MUX21X1_HVT U358 ( .A1(n377), .A2(n370), .S0(n271), .Y(n648) );
  MUX21X1_HVT U359 ( .A1(n370), .A2(n459), .S0(n387), .Y(n626) );
  MUX21X1_HVT U360 ( .A1(n459), .A2(n369), .S0(n272), .Y(n473) );
  MUX21X1_HVT U361 ( .A1(n345), .A2(n378), .S0(n338), .Y(n469) );
  MUX21X1_HVT U362 ( .A1(n243), .A2(n371), .S0(n338), .Y(n474) );
  MUX21X1_HVT U363 ( .A1(n245), .A2(n460), .S0(n271), .Y(n636) );
  MUX21X1_HVT U364 ( .A1(n370), .A2(n245), .S0(n385), .Y(n639) );
  MUX21X1_HVT U365 ( .A1(n369), .A2(n460), .S0(n386), .Y(n471) );
  MUX21X1_HVT U366 ( .A1(n460), .A2(n370), .S0(n386), .Y(n630) );
  MUX21X1_HVT U367 ( .A1(n244), .A2(n459), .S0(n338), .Y(n619) );
  MUX21X1_HVT U368 ( .A1(n378), .A2(n456), .S0(n388), .Y(n635) );
  MUX21X1_HVT U369 ( .A1(n460), .A2(n371), .S0(n388), .Y(n464) );
  MUX21X1_HVT U370 ( .A1(n379), .A2(n249), .S0(n271), .Y(n463) );
  MUX21X1_HVT U371 ( .A1(n377), .A2(n345), .S0(n338), .Y(n638) );
  MUX21X1_HVT U372 ( .A1(n249), .A2(n379), .S0(n387), .Y(n529) );
  MUX21X1_HVT U373 ( .A1(n371), .A2(n252), .S0(n271), .Y(n566) );
  XOR2X1_HVT U374 ( .A1(n384), .A2(n389), .Y(n632) );
  XNOR2X1_HVT U375 ( .A1(n252), .A2(n389), .Y(n351) );
  MUX21X1_HVT U376 ( .A1(n370), .A2(n252), .S0(n385), .Y(n472) );
  MUX21X1_HVT U377 ( .A1(n382), .A2(n248), .S0(n271), .Y(n651) );
  MUX21X1_HVT U378 ( .A1(n636), .A2(n350), .S0(n367), .Y(n544) );
  MUX21X1_HVT U379 ( .A1(n411), .A2(n377), .S0(n394), .Y(n578) );
  MUX21X1_HVT U380 ( .A1(n423), .A2(n666), .S0(n367), .Y(n613) );
  MUX21X1_HVT U381 ( .A1(n452), .A2(n351), .S0(n366), .Y(n547) );
  XOR2X1_HVT U382 ( .A1(n382), .A2(n271), .Y(n622) );
  MUX21X1_HVT U383 ( .A1(n371), .A2(n378), .S0(n272), .Y(n629) );
  MUX21X1_HVT U384 ( .A1(n383), .A2(n253), .S0(n389), .Y(n655) );
  MUX21X1_HVT U385 ( .A1(n370), .A2(n371), .S0(n388), .Y(n624) );
  MUX21X1_HVT U386 ( .A1(n381), .A2(n370), .S0(n338), .Y(n650) );
  MUX21X1_HVT U387 ( .A1(n369), .A2(n381), .S0(n388), .Y(n466) );
  MUX21X1_HVT U388 ( .A1(n382), .A2(n371), .S0(n388), .Y(n550) );
  AND2X1_HVT U389 ( .A1(n388), .A2(n371), .Y(n352) );
  NBUFFX2_HVT U390 ( .A(n457), .Y(n369) );
  NBUFFX2_HVT U391 ( .A(n653), .Y(n377) );
  AND2X1_HVT U392 ( .A1(n459), .A2(n301), .Y(n353) );
  NBUFFX2_HVT U393 ( .A(n653), .Y(n378) );
  NBUFFX2_HVT U394 ( .A(n668), .Y(n381) );
  AND2X1_HVT U395 ( .A1(n382), .A2(n391), .Y(n354) );
  NBUFFX2_HVT U396 ( .A(n668), .Y(n382) );
  NBUFFX2_HVT U397 ( .A(n393), .Y(n365) );
  NBUFFX2_HVT U398 ( .A(n392), .Y(n367) );
  NBUFFX2_HVT U399 ( .A(n392), .Y(n366) );
  NBUFFX2_HVT U400 ( .A(n461), .Y(n371) );
  NBUFFX2_HVT U401 ( .A(n393), .Y(n362) );
  NBUFFX2_HVT U402 ( .A(n393), .Y(n364) );
  NBUFFX2_HVT U403 ( .A(n393), .Y(n363) );
  NBUFFX2_HVT U404 ( .A(n392), .Y(n360) );
  NBUFFX2_HVT U405 ( .A(n392), .Y(n361) );
  NBUFFX2_HVT U406 ( .A(n392), .Y(n359) );
  XOR2X1_HVT U407 ( .A1(n372), .A2(n197), .Y(n653) );
  MUX21X1_HVT U408 ( .A1(n345), .A2(n346), .S0(n272), .Y(n462) );
  MUX21X1_HVT U409 ( .A1(n379), .A2(n346), .S0(n389), .Y(n574) );
  MUX21X1_HVT U410 ( .A1(n459), .A2(n456), .S0(n271), .Y(n555) );
  MUX21X1_HVT U411 ( .A1(n539), .A2(n540), .S0(n276), .Y(n538) );
  MUX21X1_HVT U412 ( .A1(n535), .A2(n536), .S0(n374), .Y(n534) );
  MUX21X1_HVT U413 ( .A1(n384), .A2(n346), .S0(n389), .Y(n514) );
  MUX21X1_HVT U414 ( .A1(n346), .A2(n380), .S0(n385), .Y(n467) );
  MUX21X1_HVT U415 ( .A1(n371), .A2(n346), .S0(n387), .Y(n642) );
  MUX21X1_HVT U416 ( .A1(n346), .A2(n383), .S0(n386), .Y(n468) );
  NBUFFX2_HVT U417 ( .A(in[2]), .Y(n393) );
  NBUFFX2_HVT U418 ( .A(in[2]), .Y(n392) );
  NAND2X0_HVT U419 ( .A1(n643), .A2(n398), .Y(n357) );
  NAND2X0_HVT U420 ( .A1(n646), .A2(n312), .Y(n358) );
  NAND2X0_HVT U421 ( .A1(n358), .A2(n357), .Y(n507) );
  MUX21X1_HVT U422 ( .A1(n371), .A2(n243), .S0(n385), .Y(n643) );
  MUX21X1_HVT U423 ( .A1(n244), .A2(n356), .S0(n272), .Y(n537) );
  XOR2X1_HVT U424 ( .A1(n338), .A2(n356), .Y(n620) );
  MUX21X1_HVT U425 ( .A1(n356), .A2(n382), .S0(n389), .Y(n475) );
  MUX21X1_HVT U426 ( .A1(n381), .A2(n356), .S0(n272), .Y(n470) );
  MUX21X1_HVT U427 ( .A1(n369), .A2(n356), .S0(n387), .Y(n465) );
  MUX21X1_HVT U428 ( .A1(n356), .A2(n384), .S0(n386), .Y(n652) );
  MUX21X1_HVT U429 ( .A1(n380), .A2(n356), .S0(n389), .Y(n640) );
  NBUFFX2_HVT U430 ( .A(n670), .Y(n383) );
  INVX0_HVT U431 ( .A(n631), .Y(n402) );
  INVX0_HVT U432 ( .A(n571), .Y(n403) );
  INVX0_HVT U433 ( .A(n532), .Y(n404) );
  INVX0_HVT U434 ( .A(n666), .Y(n406) );
  INVX0_HVT U435 ( .A(n627), .Y(n408) );
  INVX0_HVT U436 ( .A(n663), .Y(n409) );
  INVX0_HVT U437 ( .A(n634), .Y(n411) );
  INVX0_HVT U438 ( .A(n656), .Y(n412) );
  INVX0_HVT U439 ( .A(n657), .Y(n414) );
  INVX0_HVT U440 ( .A(n655), .Y(n415) );
  INVX0_HVT U441 ( .A(n654), .Y(n416) );
  INVX0_HVT U442 ( .A(n652), .Y(n417) );
  INVX0_HVT U443 ( .A(n651), .Y(n418) );
  INVX0_HVT U444 ( .A(n650), .Y(n419) );
  INVX0_HVT U445 ( .A(n649), .Y(n420) );
  INVX0_HVT U446 ( .A(n643), .Y(n424) );
  INVX0_HVT U447 ( .A(n641), .Y(n426) );
  INVX0_HVT U448 ( .A(n640), .Y(n427) );
  INVX0_HVT U449 ( .A(n639), .Y(n428) );
  INVX0_HVT U450 ( .A(n638), .Y(n429) );
  INVX0_HVT U451 ( .A(n636), .Y(n430) );
  INVX0_HVT U452 ( .A(n635), .Y(n431) );
  INVX0_HVT U453 ( .A(n630), .Y(n434) );
  INVX0_HVT U454 ( .A(n629), .Y(n435) );
  INVX0_HVT U455 ( .A(n626), .Y(n436) );
  INVX0_HVT U456 ( .A(n624), .Y(n437) );
  INVX0_HVT U457 ( .A(n623), .Y(n438) );
  INVX0_HVT U458 ( .A(n660), .Y(n439) );
  INVX0_HVT U459 ( .A(n475), .Y(n440) );
  INVX0_HVT U460 ( .A(n470), .Y(n445) );
  INVX0_HVT U461 ( .A(n469), .Y(n446) );
  INVX0_HVT U462 ( .A(n468), .Y(n447) );
  INVX0_HVT U463 ( .A(n467), .Y(n448) );
  INVX0_HVT U464 ( .A(n466), .Y(n449) );
  INVX0_HVT U465 ( .A(n465), .Y(n450) );
  INVX0_HVT U466 ( .A(n514), .Y(n451) );
  INVX0_HVT U467 ( .A(n464), .Y(n452) );
  INVX0_HVT U468 ( .A(n463), .Y(n453) );
  INVX0_HVT U469 ( .A(n462), .Y(n454) );
endmodule

