
module sbox_8 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n7, n23, n48, n50, n210, n211, n212, n213, n216, n217, n218, n219,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613;

  NAND2X0_HVT U3 ( .A1(n322), .A2(n317), .Y(n611) );
  NAND2X0_HVT U4 ( .A1(n315), .A2(n611), .Y(n610) );
  NAND2X0_HVT U5 ( .A1(n325), .A2(n305), .Y(n608) );
  NAND2X0_HVT U13 ( .A1(n601), .A2(n319), .Y(n602) );
  NAND2X0_HVT U15 ( .A1(n611), .A2(n275), .Y(n599) );
  NAND2X0_HVT U21 ( .A1(n314), .A2(n327), .Y(n593) );
  NAND2X0_HVT U24 ( .A1(n310), .A2(n327), .Y(n591) );
  NAND2X0_HVT U33 ( .A1(n390), .A2(n327), .Y(n582) );
  NAND2X0_HVT U35 ( .A1(n308), .A2(n327), .Y(n580) );
  NAND2X0_HVT U42 ( .A1(n323), .A2(n310), .Y(n573) );
  NAND2X0_HVT U53 ( .A1(n563), .A2(n572), .Y(n564) );
  NAND2X0_HVT U56 ( .A1(n315), .A2(n559), .Y(n560) );
  MUX41X1_HVT U57 ( .A1(n379), .A3(n595), .A2(n560), .A4(n604), .S0(n333), 
        .S1(n330), .Y(n558) );
  NAND2X0_HVT U58 ( .A1(n319), .A2(n611), .Y(n557) );
  MUX41X1_HVT U61 ( .A1(n291), .A3(n352), .A2(n351), .A4(n277), .S0(n333), 
        .S1(n331), .Y(n554) );
  NAND2X0_HVT U62 ( .A1(n327), .A2(n318), .Y(n553) );
  MUX41X1_HVT U63 ( .A1(n553), .A3(n344), .A2(n373), .A4(n350), .S0(n333), 
        .S1(n330), .Y(n552) );
  AO21X1_HVT U66 ( .A1(n348), .A2(n301), .A3(n372), .Y(n549) );
  MUX41X1_HVT U68 ( .A1(n346), .A3(n549), .A2(n548), .A4(n550), .S0(n296), 
        .S1(n249), .Y(n547) );
  MUX41X1_HVT U69 ( .A1(n547), .A3(n555), .A2(n551), .A4(n561), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n312), .A2(n542), .Y(n543) );
  MUX41X1_HVT U74 ( .A1(n544), .A3(n589), .A2(n543), .A4(n591), .S0(n298), 
        .S1(n249), .Y(n541) );
  MUX41X1_HVT U75 ( .A1(n376), .A3(n381), .A2(n394), .A4(n357), .S0(n296), 
        .S1(n249), .Y(n540) );
  MUX41X1_HVT U77 ( .A1(n606), .A3(n383), .A2(n539), .A4(n382), .S0(n302), 
        .S1(n329), .Y(n538) );
  MUX41X1_HVT U78 ( .A1(n538), .A3(n541), .A2(n540), .A4(n545), .S0(in[0]), 
        .S1(in[5]), .Y(n537) );
  AND3X1_HVT U80 ( .A1(n317), .A2(n559), .A3(n534), .Y(n535) );
  AND2X1_HVT U83 ( .A1(n323), .A2(n237), .Y(n531) );
  MUX41X1_HVT U84 ( .A1(n356), .A3(n278), .A2(n598), .A4(n531), .S0(n296), 
        .S1(n332), .Y(n530) );
  NAND2X0_HVT U85 ( .A1(n327), .A2(n393), .Y(n529) );
  MUX41X1_HVT U86 ( .A1(n381), .A3(n529), .A2(n292), .A4(n288), .S0(n296), 
        .S1(n332), .Y(n528) );
  MUX41X1_HVT U87 ( .A1(n528), .A3(n532), .A2(n530), .A4(n533), .S0(in[0]), 
        .S1(n330), .Y(n527) );
  AO21X1_HVT U93 ( .A1(n304), .A2(n521), .A3(n377), .Y(n522) );
  MUX41X1_HVT U96 ( .A1(n338), .A3(n290), .A2(n380), .A4(n519), .S0(n296), 
        .S1(n235), .Y(n518) );
  MUX41X1_HVT U97 ( .A1(n376), .A3(n290), .A2(n323), .A4(n599), .S0(n296), 
        .S1(n235), .Y(n517) );
  MUX41X1_HVT U98 ( .A1(n517), .A3(n520), .A2(n518), .A4(n525), .S0(in[0]), 
        .S1(n330), .Y(n516) );
  NAND2X0_HVT U101 ( .A1(n512), .A2(n511), .Y(n513) );
  OA21X1_HVT U109 ( .A1(n366), .A2(n257), .A3(n353), .Y(n504) );
  NAND2X0_HVT U110 ( .A1(n317), .A2(n502), .Y(n503) );
  MUX41X1_HVT U114 ( .A1(n499), .A3(n505), .A2(n501), .A4(n504), .S0(n301), 
        .S1(n235), .Y(n498) );
  AND2X1_HVT U115 ( .A1(n325), .A2(n277), .Y(n497) );
  NAND2X0_HVT U123 ( .A1(n488), .A2(n487), .Y(n489) );
  MUX41X1_HVT U125 ( .A1(n593), .A3(n295), .A2(n346), .A4(n385), .S0(n297), 
        .S1(n333), .Y(n485) );
  MUX41X1_HVT U131 ( .A1(n480), .A3(n482), .A2(n481), .A4(n483), .S0(n301), 
        .S1(n333), .Y(n479) );
  MUX41X1_HVT U132 ( .A1(n479), .A3(n492), .A2(n484), .A4(n498), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  MUX41X1_HVT U136 ( .A1(n288), .A3(n582), .A2(n387), .A4(n579), .S0(n297), 
        .S1(n333), .Y(n475) );
  MUX41X1_HVT U139 ( .A1(n473), .A3(n476), .A2(n475), .A4(n477), .S0(in[0]), 
        .S1(n330), .Y(n472) );
  AND2X1_HVT U140 ( .A1(n311), .A2(n326), .Y(n471) );
  MUX41X1_HVT U142 ( .A1(n356), .A3(n277), .A2(n374), .A4(n311), .S0(n297), 
        .S1(n333), .Y(n469) );
  NAND2X0_HVT U146 ( .A1(n323), .A2(n320), .Y(n542) );
  MUX41X1_HVT U153 ( .A1(n503), .A3(n291), .A2(n316), .A4(n340), .S0(n297), 
        .S1(n332), .Y(n459) );
  AND2X1_HVT U154 ( .A1(n304), .A2(n310), .Y(n458) );
  NAND2X0_HVT U158 ( .A1(n321), .A2(n393), .Y(n454) );
  MUX41X1_HVT U159 ( .A1(n602), .A3(n279), .A2(n454), .A4(n282), .S0(n328), 
        .S1(n235), .Y(n453) );
  MUX41X1_HVT U160 ( .A1(n453), .A3(n459), .A2(n455), .A4(n460), .S0(in[0]), 
        .S1(in[5]), .Y(n452) );
  AND2X1_HVT U162 ( .A1(n273), .A2(n542), .Y(n450) );
  MUX41X1_HVT U165 ( .A1(n593), .A3(n361), .A2(n569), .A4(n448), .S0(n333), 
        .S1(n328), .Y(n447) );
  NAND2X0_HVT U166 ( .A1(n319), .A2(n559), .Y(n446) );
  NAND2X0_HVT U167 ( .A1(n394), .A2(n327), .Y(n445) );
  MUX41X1_HVT U168 ( .A1(n379), .A3(n311), .A2(n445), .A4(n446), .S0(n329), 
        .S1(n249), .Y(n444) );
  MUX41X1_HVT U172 ( .A1(n441), .A3(n447), .A2(n444), .A4(n449), .S0(in[0]), 
        .S1(n331), .Y(n440) );
  NAND2X0_HVT U174 ( .A1(n322), .A2(n278), .Y(n601) );
  MUX41X1_HVT U176 ( .A1(n306), .A3(n439), .A2(n384), .A4(n601), .S0(n333), 
        .S1(n329), .Y(n438) );
  NAND2X0_HVT U177 ( .A1(n321), .A2(n307), .Y(n437) );
  MUX41X1_HVT U178 ( .A1(n597), .A3(n437), .A2(n388), .A4(n577), .S0(n298), 
        .S1(n249), .Y(n436) );
  MUX41X1_HVT U179 ( .A1(n587), .A3(n389), .A2(n342), .A4(n388), .S0(n329), 
        .S1(n249), .Y(n435) );
  MUX41X1_HVT U180 ( .A1(n345), .A3(n606), .A2(n602), .A4(n287), .S0(n302), 
        .S1(n328), .Y(n434) );
  MUX41X1_HVT U189 ( .A1(n426), .A3(n601), .A2(n427), .A4(n375), .S0(n302), 
        .S1(n329), .Y(n425) );
  MUX41X1_HVT U190 ( .A1(n425), .A3(n428), .A2(n429), .A4(n432), .S0(n331), 
        .S1(in[0]), .Y(n424) );
  MUX41X1_HVT U194 ( .A1(n574), .A3(n588), .A2(n386), .A4(n311), .S0(n302), 
        .S1(n328), .Y(n421) );
  AO21X1_HVT U197 ( .A1(n292), .A2(n303), .A3(n377), .Y(n418) );
  MUX41X1_HVT U203 ( .A1(n579), .A3(n369), .A2(n603), .A4(n583), .S0(n329), 
        .S1(n48), .Y(n412) );
  MUX41X1_HVT U205 ( .A1(n237), .A3(n611), .A2(n389), .A4(n244), .S0(n329), 
        .S1(n249), .Y(n410) );
  NAND2X0_HVT U208 ( .A1(n321), .A2(n314), .Y(n502) );
  NAND2X0_HVT U212 ( .A1(n324), .A2(n312), .Y(n559) );
  NAND2X0_HVT U214 ( .A1(n273), .A2(n327), .Y(n408) );
  NAND2X0_HVT U215 ( .A1(n502), .A2(n313), .Y(n407) );
  NAND2X0_HVT U218 ( .A1(n391), .A2(n321), .Y(n461) );
  NAND2X0_HVT U220 ( .A1(n303), .A2(n408), .Y(n534) );
  OA21X1_HVT U1 ( .A1(n575), .A2(n335), .A3(n461), .Y(n462) );
  MUX21X1_HVT U2 ( .A1(n564), .A2(n565), .S0(n302), .Y(n562) );
  INVX1_HVT U6 ( .A(n322), .Y(n327) );
  INVX1_HVT U7 ( .A(n329), .Y(n257) );
  INVX2_HVT U8 ( .A(n272), .Y(n329) );
  INVX1_HVT U9 ( .A(n326), .Y(n321) );
  MUX41X1_HVT U10 ( .A1(n354), .A3(n355), .A2(n378), .A4(n337), .S0(in[7]), 
        .S1(n280), .Y(n566) );
  IBUFFX2_HVT U11 ( .A(in[7]), .Y(n336) );
  INVX1_HVT U12 ( .A(n406), .Y(n378) );
  MUX21X2_HVT U14 ( .A1(n566), .A2(n562), .S0(n7), .Y(n561) );
  IBUFFX16_HVT U16 ( .A(n299), .Y(n7) );
  INVX2_HVT U17 ( .A(n326), .Y(n325) );
  MUX21X1_HVT U18 ( .A1(n571), .A2(n546), .S0(n299), .Y(n545) );
  INVX0_HVT U19 ( .A(n250), .Y(n239) );
  INVX1_HVT U20 ( .A(n326), .Y(n322) );
  INVX1_HVT U22 ( .A(n217), .Y(n470) );
  INVX0_HVT U23 ( .A(n363), .Y(n232) );
  MUX41X1_HVT U25 ( .A1(n353), .A3(n293), .A2(n557), .A4(n295), .S0(n335), 
        .S1(n23), .Y(n556) );
  IBUFFX16_HVT U26 ( .A(n330), .Y(n23) );
  INVX1_HVT U27 ( .A(n336), .Y(n333) );
  IBUFFX2_HVT U28 ( .A(in[7]), .Y(n335) );
  MUX21X1_HVT U29 ( .A1(n556), .A2(n558), .S0(n299), .Y(n555) );
  MUX41X1_HVT U30 ( .A1(n368), .A3(n314), .A2(n370), .A4(n358), .S0(n333), 
        .S1(n328), .Y(n432) );
  INVX1_HVT U31 ( .A(n247), .Y(n48) );
  MUX41X1_HVT U32 ( .A1(n410), .A3(n412), .A2(n411), .A4(n413), .S0(in[0]), 
        .S1(in[5]), .Y(n409) );
  NBUFFX2_HVT U34 ( .A(in[7]), .Y(n249) );
  MUX21X1_HVT U36 ( .A1(n414), .A2(n415), .S0(n299), .Y(n413) );
  MUX41X1_HVT U37 ( .A1(n573), .A3(n567), .A2(n580), .A4(n423), .S0(n249), 
        .S1(n328), .Y(n422) );
  MUX41X1_HVT U38 ( .A1(n438), .A3(n435), .A2(n436), .A4(n434), .S0(n50), .S1(
        n210), .Y(n433) );
  IBUFFX16_HVT U39 ( .A(in[0]), .Y(n50) );
  IBUFFX16_HVT U40 ( .A(in[5]), .Y(n210) );
  NAND2X1_HVT U41 ( .A1(n527), .A2(n211), .Y(n212) );
  NAND2X0_HVT U43 ( .A1(n537), .A2(n216), .Y(n213) );
  NAND2X0_HVT U44 ( .A1(n212), .A2(n213), .Y(out[1]) );
  INVX0_HVT U45 ( .A(n216), .Y(n211) );
  INVX1_HVT U46 ( .A(n236), .Y(n216) );
  MUX41X1_HVT U47 ( .A1(n232), .A3(n231), .A2(n219), .A4(n218), .S0(n233), 
        .S1(n336), .Y(n217) );
  IBUFFX16_HVT U48 ( .A(n590), .Y(n218) );
  IBUFFX16_HVT U49 ( .A(n367), .Y(n219) );
  IBUFFX16_HVT U50 ( .A(n471), .Y(n231) );
  IBUFFX16_HVT U51 ( .A(n298), .Y(n233) );
  MUX41X1_HVT U52 ( .A1(n470), .A3(n466), .A2(n469), .A4(n465), .S0(n269), 
        .S1(n234), .Y(n464) );
  IBUFFX16_HVT U54 ( .A(n330), .Y(n234) );
  NBUFFX2_HVT U55 ( .A(n332), .Y(n235) );
  INVX1_HVT U59 ( .A(n335), .Y(n332) );
  IBUFFX16_HVT U60 ( .A(in[6]), .Y(n236) );
  INVX0_HVT U64 ( .A(n249), .Y(n247) );
  INVX1_HVT U65 ( .A(n395), .Y(n237) );
  INVX1_HVT U67 ( .A(in[4]), .Y(n395) );
  MUX21X2_HVT U70 ( .A1(n613), .A2(n316), .S0(n239), .Y(n238) );
  INVX8_HVT U71 ( .A(n238), .Y(n588) );
  INVX1_HVT U72 ( .A(n326), .Y(n323) );
  MUX21X2_HVT U76 ( .A1(n433), .A2(n424), .S0(n240), .Y(out[6]) );
  IBUFFX16_HVT U79 ( .A(in[6]), .Y(n240) );
  MUX21X2_HVT U81 ( .A1(n600), .A2(n244), .S0(n241), .Y(n515) );
  IBUFFX16_HVT U82 ( .A(n300), .Y(n241) );
  MUX41X1_HVT U88 ( .A1(n509), .A3(n507), .A2(n514), .A4(n510), .S0(n242), 
        .S1(n243), .Y(n506) );
  IBUFFX16_HVT U89 ( .A(in[5]), .Y(n242) );
  IBUFFX16_HVT U90 ( .A(n269), .Y(n243) );
  INVX0_HVT U91 ( .A(n576), .Y(n368) );
  INVX1_HVT U92 ( .A(n244), .Y(n584) );
  MUX21X2_HVT U94 ( .A1(n515), .A2(n291), .S0(n285), .Y(n514) );
  NAND2X2_HVT U95 ( .A1(n253), .A2(n254), .Y(out[4]) );
  MUX21X1_HVT U99 ( .A1(n245), .A2(n246), .S0(n321), .Y(n244) );
  IBUFFX16_HVT U100 ( .A(n320), .Y(n245) );
  IBUFFX16_HVT U102 ( .A(n312), .Y(n246) );
  MUX21X2_HVT U103 ( .A1(n256), .A2(n255), .S0(n247), .Y(n428) );
  OA21X2_HVT U104 ( .A1(n293), .A2(n335), .A3(n584), .Y(n442) );
  MUX41X1_HVT U105 ( .A1(n451), .A3(n289), .A2(n450), .A4(n352), .S0(n248), 
        .S1(n335), .Y(n449) );
  IBUFFX16_HVT U106 ( .A(n328), .Y(n248) );
  OA21X1_HVT U107 ( .A1(n341), .A2(n335), .A3(n584), .Y(n467) );
  NAND2X2_HVT U108 ( .A1(n283), .A2(n284), .Y(out[2]) );
  MUX21X2_HVT U111 ( .A1(n576), .A2(n290), .S0(n257), .Y(n255) );
  INVX2_HVT U112 ( .A(in[1]), .Y(n326) );
  MUX21X1_HVT U113 ( .A1(n264), .A2(n265), .S0(n235), .Y(n509) );
  NBUFFX2_HVT U116 ( .A(n322), .Y(n250) );
  NBUFFX2_HVT U117 ( .A(n322), .Y(n251) );
  IBUFFX2_HVT U118 ( .A(n326), .Y(n324) );
  MUX21X1_HVT U119 ( .A1(n318), .A2(n500), .S0(n286), .Y(n499) );
  INVX1_HVT U120 ( .A(n268), .Y(n328) );
  INVX0_HVT U121 ( .A(n252), .Y(n278) );
  INVX0_HVT U122 ( .A(n276), .Y(n277) );
  XNOR2X2_HVT U124 ( .A1(n306), .A2(n309), .Y(n252) );
  INVX0_HVT U126 ( .A(n252), .Y(n274) );
  INVX1_HVT U127 ( .A(in[0]), .Y(n269) );
  INVX0_HVT U128 ( .A(in[6]), .Y(n263) );
  INVX1_HVT U129 ( .A(n309), .Y(n392) );
  INVX1_HVT U130 ( .A(n296), .Y(n272) );
  INVX1_HVT U133 ( .A(n298), .Y(n268) );
  INVX0_HVT U134 ( .A(n330), .Y(n280) );
  MUX41X1_HVT U135 ( .A1(n584), .A3(n357), .A2(n497), .A4(n602), .S0(n257), 
        .S1(n336), .Y(n496) );
  MUX21X2_HVT U137 ( .A1(n526), .A2(n378), .S0(n268), .Y(n259) );
  NAND2X0_HVT U138 ( .A1(n472), .A2(n260), .Y(n253) );
  NAND2X0_HVT U141 ( .A1(n464), .A2(n263), .Y(n254) );
  MUX21X1_HVT U143 ( .A1(n569), .A2(n542), .S0(n257), .Y(n256) );
  MUX21X1_HVT U144 ( .A1(n573), .A2(n569), .S0(n268), .Y(n258) );
  MUX21X1_HVT U145 ( .A1(n258), .A2(n259), .S0(n235), .Y(n525) );
  NAND2X0_HVT U147 ( .A1(n416), .A2(n260), .Y(n261) );
  NAND2X0_HVT U148 ( .A1(n409), .A2(n263), .Y(n262) );
  NAND2X0_HVT U149 ( .A1(n262), .A2(n261), .Y(out[7]) );
  INVX1_HVT U150 ( .A(n263), .Y(n260) );
  MUX21X1_HVT U151 ( .A1(n347), .A2(n611), .S0(n272), .Y(n264) );
  MUX21X1_HVT U152 ( .A1(n580), .A2(n360), .S0(n272), .Y(n265) );
  MUX41X1_HVT U155 ( .A1(n422), .A3(n421), .A2(n420), .A4(n417), .S0(n280), 
        .S1(n269), .Y(n416) );
  MUX21X1_HVT U156 ( .A1(n380), .A2(n273), .S0(n268), .Y(n266) );
  MUX21X1_HVT U157 ( .A1(n578), .A2(n319), .S0(n268), .Y(n267) );
  MUX21X1_HVT U161 ( .A1(n266), .A2(n267), .S0(n249), .Y(n420) );
  INVX1_HVT U163 ( .A(n404), .Y(n380) );
  MUX41X1_HVT U164 ( .A1(n569), .A3(n376), .A2(n542), .A4(n387), .S0(n268), 
        .S1(n336), .Y(n465) );
  MUX21X2_HVT U169 ( .A1(n493), .A2(n496), .S0(n301), .Y(n492) );
  MUX41X1_HVT U170 ( .A1(n602), .A3(n592), .A2(n560), .A4(n364), .S0(n249), 
        .S1(n268), .Y(n411) );
  MUX21X1_HVT U171 ( .A1(n355), .A2(n570), .S0(n272), .Y(n270) );
  MUX21X1_HVT U173 ( .A1(n600), .A2(n338), .S0(n272), .Y(n271) );
  MUX21X1_HVT U175 ( .A1(n270), .A2(n271), .S0(n332), .Y(n532) );
  AO21X2_HVT U181 ( .A1(n326), .A2(n391), .A3(n335), .Y(n512) );
  OA21X2_HVT U182 ( .A1(n581), .A2(n335), .A3(n356), .Y(n430) );
  OA21X2_HVT U183 ( .A1(n607), .A2(n335), .A3(n367), .Y(n414) );
  INVX1_HVT U184 ( .A(n252), .Y(n273) );
  INVX1_HVT U185 ( .A(n274), .Y(n275) );
  INVX1_HVT U186 ( .A(n279), .Y(n276) );
  INVX1_HVT U187 ( .A(n274), .Y(n279) );
  AND3X2_HVT U188 ( .A1(n300), .A2(n327), .A3(n237), .Y(n482) );
  AO21X2_HVT U191 ( .A1(n300), .A2(n311), .A3(n276), .Y(n494) );
  MUX21X2_HVT U192 ( .A1(n279), .A2(n305), .S0(n250), .Y(n598) );
  MUX21X2_HVT U193 ( .A1(n598), .A2(n287), .S0(n302), .Y(n415) );
  NBUFFX2_HVT U195 ( .A(in[2]), .Y(n297) );
  INVX1_HVT U196 ( .A(n281), .Y(n476) );
  XNOR2X1_HVT U198 ( .A1(n323), .A2(in[2]), .Y(n286) );
  NAND2X0_HVT U199 ( .A1(n516), .A2(n260), .Y(n283) );
  INVX0_HVT U200 ( .A(n608), .Y(n282) );
  MUX41X1_HVT U201 ( .A1(n359), .A3(n568), .A2(n508), .A4(n375), .S0(n296), 
        .S1(n332), .Y(n507) );
  MUX41X1_HVT U202 ( .A1(n238), .A3(n282), .A2(n311), .A4(n399), .S0(n268), 
        .S1(n336), .Y(n281) );
  INVX1_HVT U204 ( .A(n399), .Y(n386) );
  XNOR2X1_HVT U206 ( .A1(n272), .A2(n336), .Y(n285) );
  NAND2X0_HVT U207 ( .A1(n506), .A2(n263), .Y(n284) );
  MUX21X2_HVT U209 ( .A1(n440), .A2(n452), .S0(in[6]), .Y(out[5]) );
  INVX0_HVT U210 ( .A(n336), .Y(n334) );
  INVX1_HVT U211 ( .A(n609), .Y(n390) );
  MUX21X1_HVT U213 ( .A1(n289), .A2(n351), .S0(n297), .Y(n481) );
  AND2X1_HVT U216 ( .A1(n275), .A2(n559), .Y(n287) );
  INVX1_HVT U217 ( .A(n316), .Y(n394) );
  MUX21X1_HVT U219 ( .A1(n390), .A2(n393), .S0(n301), .Y(n563) );
  MUX21X1_HVT U221 ( .A1(n584), .A2(n503), .S0(n297), .Y(n501) );
  NBUFFX2_HVT U222 ( .A(n609), .Y(n314) );
  NBUFFX2_HVT U223 ( .A(n609), .Y(n315) );
  MUX21X1_HVT U224 ( .A1(n347), .A2(n391), .S0(n301), .Y(n548) );
  AND2X1_HVT U225 ( .A1(n317), .A2(n542), .Y(n288) );
  MUX21X1_HVT U226 ( .A1(n275), .A2(n393), .S0(n322), .Y(n607) );
  MUX21X1_HVT U227 ( .A1(n485), .A2(n486), .S0(n301), .Y(n484) );
  MUX21X1_HVT U228 ( .A1(n490), .A2(n489), .S0(n304), .Y(n486) );
  MUX21X1_HVT U229 ( .A1(n317), .A2(n275), .S0(n321), .Y(n574) );
  MUX21X1_HVT U230 ( .A1(n277), .A2(n308), .S0(n325), .Y(n511) );
  MUX21X1_HVT U231 ( .A1(n474), .A2(n610), .S0(n300), .Y(n473) );
  MUX21X1_HVT U232 ( .A1(n592), .A2(n368), .S0(n303), .Y(n474) );
  MUX21X1_HVT U233 ( .A1(n390), .A2(n394), .S0(n324), .Y(n439) );
  MUX21X1_HVT U234 ( .A1(n315), .A2(n273), .S0(n323), .Y(n578) );
  MUX21X1_HVT U235 ( .A1(n393), .A2(n279), .S0(n324), .Y(n451) );
  MUX21X1_HVT U236 ( .A1(n277), .A2(n390), .S0(n324), .Y(n519) );
  MUX21X1_HVT U237 ( .A1(n273), .A2(n391), .S0(n324), .Y(n399) );
  MUX21X1_HVT U238 ( .A1(n276), .A2(n394), .S0(n251), .Y(n590) );
  MUX21X1_HVT U239 ( .A1(n314), .A2(n313), .S0(n323), .Y(n526) );
  MUX21X1_HVT U240 ( .A1(n276), .A2(n308), .S0(n321), .Y(n539) );
  XOR2X1_HVT U241 ( .A1(n274), .A2(n322), .Y(n569) );
  MUX21X1_HVT U242 ( .A1(n393), .A2(n390), .S0(n324), .Y(n577) );
  MUX21X1_HVT U243 ( .A1(n305), .A2(n394), .S0(n325), .Y(n575) );
  MUX21X1_HVT U244 ( .A1(n308), .A2(n390), .S0(n250), .Y(n586) );
  MUX21X1_HVT U245 ( .A1(n362), .A2(n478), .S0(n299), .Y(n477) );
  MUX21X1_HVT U246 ( .A1(n385), .A2(n313), .S0(n303), .Y(n478) );
  MUX21X1_HVT U247 ( .A1(n494), .A2(n495), .S0(n303), .Y(n493) );
  MUX21X1_HVT U248 ( .A1(n340), .A2(n364), .S0(n297), .Y(n495) );
  NAND2X0_HVT U249 ( .A1(n306), .A2(n392), .Y(n609) );
  MUX21X1_HVT U250 ( .A1(n390), .A2(n307), .S0(n322), .Y(n400) );
  MUX21X1_HVT U251 ( .A1(n305), .A2(n273), .S0(n325), .Y(n402) );
  NBUFFX2_HVT U252 ( .A(n612), .Y(n316) );
  MUX21X1_HVT U253 ( .A1(n393), .A2(n305), .S0(n321), .Y(n581) );
  MUX21X1_HVT U254 ( .A1(n339), .A2(n491), .S0(n298), .Y(n490) );
  MUX21X1_HVT U255 ( .A1(n307), .A2(n305), .S0(n324), .Y(n491) );
  NBUFFX2_HVT U256 ( .A(n612), .Y(n317) );
  XOR2X1_HVT U257 ( .A1(n322), .A2(n391), .Y(n570) );
  MUX21X1_HVT U258 ( .A1(n305), .A2(n320), .S0(n323), .Y(n426) );
  MUX21X1_HVT U259 ( .A1(n319), .A2(n317), .S0(n323), .Y(n427) );
  MUX21X1_HVT U260 ( .A1(n391), .A2(n390), .S0(n251), .Y(n596) );
  INVX1_HVT U261 ( .A(n311), .Y(n391) );
  INVX1_HVT U262 ( .A(n613), .Y(n393) );
  MUX21X1_HVT U263 ( .A1(n318), .A2(n312), .S0(n250), .Y(n600) );
  MUX21X1_HVT U264 ( .A1(n315), .A2(n320), .S0(n323), .Y(n521) );
  MUX21X1_HVT U265 ( .A1(n305), .A2(n393), .S0(n250), .Y(n604) );
  NBUFFX2_HVT U266 ( .A(n612), .Y(n318) );
  MUX21X1_HVT U267 ( .A1(n305), .A2(n308), .S0(n323), .Y(n423) );
  XOR2X1_HVT U268 ( .A1(n316), .A2(n321), .Y(n567) );
  XNOR2X1_HVT U269 ( .A1(n315), .A2(n325), .Y(n289) );
  AND2X1_HVT U270 ( .A1(n321), .A2(n394), .Y(n290) );
  MUX21X1_HVT U271 ( .A1(n314), .A2(n305), .S0(n251), .Y(n603) );
  MUX21X1_HVT U272 ( .A1(n316), .A2(n307), .S0(n325), .Y(n406) );
  MUX21X1_HVT U273 ( .A1(n316), .A2(n314), .S0(n325), .Y(n398) );
  MUX21X1_HVT U274 ( .A1(n312), .A2(n305), .S0(n325), .Y(n404) );
  AND2X1_HVT U275 ( .A1(n319), .A2(n502), .Y(n291) );
  XNOR2X1_HVT U276 ( .A1(n319), .A2(n325), .Y(n292) );
  MUX21X1_HVT U277 ( .A1(n313), .A2(n307), .S0(n325), .Y(n544) );
  MUX21X1_HVT U278 ( .A1(n313), .A2(n320), .S0(n299), .Y(n488) );
  XOR2X1_HVT U279 ( .A1(n306), .A2(n321), .Y(n589) );
  NBUFFX2_HVT U280 ( .A(n334), .Y(n304) );
  NBUFFX2_HVT U281 ( .A(n334), .Y(n302) );
  NBUFFX2_HVT U282 ( .A(n334), .Y(n303) );
  NBUFFX2_HVT U283 ( .A(n392), .Y(n305) );
  NBUFFX2_HVT U284 ( .A(n331), .Y(n301) );
  NBUFFX2_HVT U285 ( .A(in[2]), .Y(n298) );
  NBUFFX2_HVT U286 ( .A(in[2]), .Y(n300) );
  NBUFFX2_HVT U287 ( .A(in[2]), .Y(n299) );
  NBUFFX2_HVT U288 ( .A(in[2]), .Y(n296) );
  NBUFFX2_HVT U289 ( .A(n395), .Y(n306) );
  MUX21X1_HVT U290 ( .A1(n252), .A2(n310), .S0(n251), .Y(n592) );
  MUX21X1_HVT U291 ( .A1(n513), .A2(n362), .S0(n299), .Y(n510) );
  MUX21X1_HVT U292 ( .A1(n430), .A2(n431), .S0(n299), .Y(n429) );
  MUX21X1_HVT U293 ( .A1(n529), .A2(n310), .S0(n303), .Y(n431) );
  MUX21X1_HVT U294 ( .A1(n552), .A2(n554), .S0(n299), .Y(n551) );
  XOR2X1_HVT U295 ( .A1(n324), .A2(n309), .Y(n568) );
  MUX21X1_HVT U296 ( .A1(n312), .A2(n279), .S0(n324), .Y(n508) );
  MUX21X1_HVT U297 ( .A1(n536), .A2(n535), .S0(n300), .Y(n533) );
  MUX21X1_HVT U298 ( .A1(n594), .A2(n313), .S0(n304), .Y(n536) );
  AND2X1_HVT U299 ( .A1(n252), .A2(n327), .Y(n293) );
  MUX21X1_HVT U300 ( .A1(n310), .A2(n390), .S0(n321), .Y(n576) );
  MUX21X1_HVT U301 ( .A1(n462), .A2(n463), .S0(n300), .Y(n460) );
  MUX21X1_HVT U302 ( .A1(n382), .A2(n391), .S0(n303), .Y(n463) );
  MUX21X1_HVT U303 ( .A1(n393), .A2(n380), .S0(n304), .Y(n546) );
  XOR2X1_HVT U304 ( .A1(n335), .A2(n588), .Y(n571) );
  MUX21X1_HVT U305 ( .A1(n443), .A2(n442), .S0(n300), .Y(n441) );
  MUX21X1_HVT U306 ( .A1(n313), .A2(n380), .S0(n304), .Y(n443) );
  MUX21X1_HVT U307 ( .A1(n468), .A2(n467), .S0(n300), .Y(n466) );
  MUX21X1_HVT U308 ( .A1(n586), .A2(n343), .S0(n304), .Y(n468) );
  MUX21X1_HVT U309 ( .A1(n391), .A2(n394), .S0(n324), .Y(n448) );
  NAND2X0_HVT U310 ( .A1(n309), .A2(n308), .Y(n612) );
  NBUFFX2_HVT U311 ( .A(n395), .Y(n308) );
  MUX21X1_HVT U312 ( .A1(n394), .A2(n310), .S0(n251), .Y(n595) );
  MUX21X1_HVT U313 ( .A1(n365), .A2(n611), .S0(n298), .Y(n505) );
  MUX21X1_HVT U314 ( .A1(n456), .A2(n457), .S0(n300), .Y(n455) );
  MUX21X1_HVT U315 ( .A1(n458), .A2(n318), .S0(n294), .Y(n457) );
  MUX21X1_HVT U316 ( .A1(n577), .A2(n383), .S0(n302), .Y(n456) );
  MUX21X1_HVT U317 ( .A1(n597), .A2(n363), .S0(n298), .Y(n480) );
  MUX21X1_HVT U318 ( .A1(n611), .A2(n326), .S0(n299), .Y(n487) );
  NBUFFX2_HVT U319 ( .A(n605), .Y(n311) );
  MUX21X1_HVT U320 ( .A1(n310), .A2(n391), .S0(n323), .Y(n403) );
  MUX21X1_HVT U321 ( .A1(n310), .A2(n580), .S0(n301), .Y(n565) );
  XOR2X1_HVT U322 ( .A1(n324), .A2(n331), .Y(n572) );
  MUX21X1_HVT U323 ( .A1(n315), .A2(n310), .S0(n250), .Y(n606) );
  NBUFFX2_HVT U324 ( .A(n605), .Y(n312) );
  MUX21X1_HVT U325 ( .A1(n585), .A2(n407), .S0(n302), .Y(n401) );
  MUX21X1_HVT U326 ( .A1(n359), .A2(n585), .S0(n298), .Y(n483) );
  MUX21X1_HVT U327 ( .A1(n349), .A2(n327), .S0(n301), .Y(n550) );
  MUX21X1_HVT U328 ( .A1(n371), .A2(n388), .S0(n303), .Y(n419) );
  MUX21X1_HVT U329 ( .A1(n318), .A2(n524), .S0(n294), .Y(n523) );
  MUX21X1_HVT U330 ( .A1(n310), .A2(n307), .S0(n304), .Y(n524) );
  NBUFFX2_HVT U331 ( .A(n613), .Y(n320) );
  NBUFFX2_HVT U332 ( .A(n395), .Y(n307) );
  NBUFFX2_HVT U333 ( .A(n605), .Y(n313) );
  NBUFFX2_HVT U334 ( .A(n613), .Y(n319) );
  XNOR2X1_HVT U335 ( .A1(n335), .A2(n322), .Y(n294) );
  AND2X1_HVT U336 ( .A1(n305), .A2(n327), .Y(n295) );
  NBUFFX2_HVT U337 ( .A(in[5]), .Y(n331) );
  NBUFFX2_HVT U338 ( .A(in[5]), .Y(n330) );
  MUX21X1_HVT U339 ( .A1(n419), .A2(n418), .S0(n299), .Y(n417) );
  MUX21X1_HVT U340 ( .A1(n522), .A2(n523), .S0(n300), .Y(n520) );
  MUX21X1_HVT U341 ( .A1(n390), .A2(n237), .S0(n321), .Y(n583) );
  MUX21X1_HVT U342 ( .A1(n237), .A2(n276), .S0(n325), .Y(n405) );
  MUX21X1_HVT U343 ( .A1(n237), .A2(n393), .S0(n323), .Y(n579) );
  MUX21X1_HVT U344 ( .A1(n237), .A2(n391), .S0(n251), .Y(n597) );
  NAND2X0_HVT U345 ( .A1(in[4]), .A2(n392), .Y(n605) );
  NAND2X0_HVT U346 ( .A1(n309), .A2(in[4]), .Y(n613) );
  MUX21X1_HVT U347 ( .A1(n237), .A2(n318), .S0(n250), .Y(n594) );
  MUX21X1_HVT U348 ( .A1(n320), .A2(n237), .S0(n251), .Y(n587) );
  MUX21X1_HVT U349 ( .A1(n310), .A2(n237), .S0(n297), .Y(n500) );
  MUX21X1_HVT U350 ( .A1(n237), .A2(n312), .S0(n324), .Y(n397) );
  MUX21X1_HVT U351 ( .A1(n237), .A2(n319), .S0(n325), .Y(n396) );
  MUX21X1_HVT U352 ( .A1(n305), .A2(n237), .S0(n251), .Y(n585) );
  NBUFFX2_HVT U353 ( .A(in[3]), .Y(n309) );
  NBUFFX2_HVT U354 ( .A(in[3]), .Y(n310) );
  INVX0_HVT U355 ( .A(n593), .Y(n337) );
  INVX0_HVT U356 ( .A(n591), .Y(n338) );
  INVX0_HVT U357 ( .A(n582), .Y(n339) );
  INVX0_HVT U358 ( .A(n580), .Y(n340) );
  INVX0_HVT U359 ( .A(n445), .Y(n341) );
  INVX0_HVT U360 ( .A(n408), .Y(n342) );
  INVX0_HVT U361 ( .A(n611), .Y(n343) );
  INVX0_HVT U362 ( .A(n599), .Y(n344) );
  INVX0_HVT U363 ( .A(n610), .Y(n345) );
  INVX0_HVT U364 ( .A(n607), .Y(n346) );
  INVX0_HVT U365 ( .A(n606), .Y(n347) );
  INVX0_HVT U366 ( .A(n604), .Y(n348) );
  INVX0_HVT U367 ( .A(n603), .Y(n349) );
  INVX0_HVT U368 ( .A(n600), .Y(n350) );
  INVX0_HVT U369 ( .A(n598), .Y(n351) );
  INVX0_HVT U370 ( .A(n597), .Y(n352) );
  INVX0_HVT U371 ( .A(n596), .Y(n353) );
  INVX0_HVT U372 ( .A(n595), .Y(n354) );
  INVX0_HVT U373 ( .A(n594), .Y(n355) );
  INVX0_HVT U374 ( .A(n592), .Y(n356) );
  INVX0_HVT U375 ( .A(n590), .Y(n357) );
  INVX0_HVT U376 ( .A(n589), .Y(n358) );
  INVX0_HVT U377 ( .A(n587), .Y(n359) );
  INVX0_HVT U378 ( .A(n586), .Y(n360) );
  INVX0_HVT U379 ( .A(n585), .Y(n361) );
  INVX0_HVT U380 ( .A(n401), .Y(n362) );
  INVX0_HVT U381 ( .A(n583), .Y(n363) );
  INVX0_HVT U382 ( .A(n581), .Y(n364) );
  INVX0_HVT U383 ( .A(n579), .Y(n365) );
  INVX0_HVT U384 ( .A(n578), .Y(n366) );
  INVX0_HVT U385 ( .A(n577), .Y(n367) );
  INVX0_HVT U386 ( .A(n575), .Y(n369) );
  INVX0_HVT U387 ( .A(n574), .Y(n370) );
  INVX0_HVT U388 ( .A(n573), .Y(n371) );
  INVX0_HVT U389 ( .A(n542), .Y(n372) );
  INVX0_HVT U390 ( .A(n602), .Y(n373) );
  INVX0_HVT U391 ( .A(n502), .Y(n374) );
  INVX0_HVT U392 ( .A(n407), .Y(n375) );
  INVX0_HVT U393 ( .A(n559), .Y(n376) );
  INVX0_HVT U394 ( .A(n461), .Y(n377) );
  INVX0_HVT U395 ( .A(n405), .Y(n379) );
  INVX0_HVT U396 ( .A(n403), .Y(n381) );
  INVX0_HVT U397 ( .A(n402), .Y(n382) );
  INVX0_HVT U398 ( .A(n521), .Y(n383) );
  INVX0_HVT U399 ( .A(n511), .Y(n384) );
  INVX0_HVT U400 ( .A(n400), .Y(n385) );
  INVX0_HVT U401 ( .A(n398), .Y(n387) );
  INVX0_HVT U402 ( .A(n397), .Y(n388) );
  INVX0_HVT U403 ( .A(n396), .Y(n389) );
endmodule

