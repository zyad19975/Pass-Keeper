
module reg_D_0 ( clk, rst, enable, in, out );
  input [127:0] in;
  output [127:0] out;
  input clk, rst, enable;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n1, n2,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156;
  tri   clk;
  tri   rst;
  tri   [127:0] out;

  DFFX1_HVT \out_reg[127]  ( .D(n132), .CLK(clk), .Q(out[127]) );
  DFFX1_HVT \out_reg[126]  ( .D(n131), .CLK(clk), .Q(out[126]) );
  DFFX1_HVT \out_reg[125]  ( .D(n130), .CLK(clk), .Q(out[125]) );
  DFFX1_HVT \out_reg[124]  ( .D(n129), .CLK(clk), .Q(out[124]) );
  DFFX1_HVT \out_reg[123]  ( .D(n128), .CLK(clk), .Q(out[123]) );
  DFFX1_HVT \out_reg[122]  ( .D(n127), .CLK(clk), .Q(out[122]) );
  DFFX1_HVT \out_reg[121]  ( .D(n126), .CLK(clk), .Q(out[121]) );
  DFFX1_HVT \out_reg[120]  ( .D(n125), .CLK(clk), .Q(out[120]) );
  DFFX1_HVT \out_reg[119]  ( .D(n124), .CLK(clk), .Q(out[119]) );
  DFFX1_HVT \out_reg[118]  ( .D(n123), .CLK(clk), .Q(out[118]) );
  DFFX1_HVT \out_reg[117]  ( .D(n122), .CLK(clk), .Q(out[117]) );
  DFFX1_HVT \out_reg[116]  ( .D(n121), .CLK(clk), .Q(out[116]) );
  DFFX1_HVT \out_reg[115]  ( .D(n120), .CLK(clk), .Q(out[115]) );
  DFFX1_HVT \out_reg[114]  ( .D(n119), .CLK(clk), .Q(out[114]) );
  DFFX1_HVT \out_reg[113]  ( .D(n118), .CLK(clk), .Q(out[113]) );
  DFFX1_HVT \out_reg[112]  ( .D(n117), .CLK(clk), .Q(out[112]) );
  DFFX1_HVT \out_reg[111]  ( .D(n116), .CLK(clk), .Q(out[111]) );
  DFFX1_HVT \out_reg[110]  ( .D(n115), .CLK(clk), .Q(out[110]) );
  DFFX1_HVT \out_reg[109]  ( .D(n114), .CLK(clk), .Q(out[109]) );
  DFFX1_HVT \out_reg[108]  ( .D(n113), .CLK(clk), .Q(out[108]) );
  DFFX1_HVT \out_reg[107]  ( .D(n112), .CLK(clk), .Q(out[107]) );
  DFFX1_HVT \out_reg[106]  ( .D(n111), .CLK(clk), .Q(out[106]) );
  DFFX1_HVT \out_reg[105]  ( .D(n110), .CLK(clk), .Q(out[105]) );
  DFFX1_HVT \out_reg[104]  ( .D(n109), .CLK(clk), .Q(out[104]) );
  DFFX1_HVT \out_reg[103]  ( .D(n108), .CLK(clk), .Q(out[103]) );
  DFFX1_HVT \out_reg[102]  ( .D(n107), .CLK(clk), .Q(out[102]) );
  DFFX1_HVT \out_reg[101]  ( .D(n106), .CLK(clk), .Q(out[101]) );
  DFFX1_HVT \out_reg[100]  ( .D(n105), .CLK(clk), .Q(out[100]) );
  DFFX1_HVT \out_reg[99]  ( .D(n104), .CLK(clk), .Q(out[99]) );
  DFFX1_HVT \out_reg[98]  ( .D(n103), .CLK(clk), .Q(out[98]) );
  DFFX1_HVT \out_reg[97]  ( .D(n102), .CLK(clk), .Q(out[97]) );
  DFFX1_HVT \out_reg[96]  ( .D(n101), .CLK(clk), .Q(out[96]) );
  DFFX1_HVT \out_reg[95]  ( .D(n100), .CLK(clk), .Q(out[95]) );
  DFFX1_HVT \out_reg[94]  ( .D(n99), .CLK(clk), .Q(out[94]) );
  DFFX1_HVT \out_reg[93]  ( .D(n98), .CLK(clk), .Q(out[93]) );
  DFFX1_HVT \out_reg[92]  ( .D(n97), .CLK(clk), .Q(out[92]) );
  DFFX1_HVT \out_reg[91]  ( .D(n96), .CLK(clk), .Q(out[91]) );
  DFFX1_HVT \out_reg[90]  ( .D(n95), .CLK(clk), .Q(out[90]) );
  DFFX1_HVT \out_reg[89]  ( .D(n94), .CLK(clk), .Q(out[89]) );
  DFFX1_HVT \out_reg[88]  ( .D(n93), .CLK(clk), .Q(out[88]) );
  DFFX1_HVT \out_reg[87]  ( .D(n92), .CLK(clk), .Q(out[87]) );
  DFFX1_HVT \out_reg[86]  ( .D(n91), .CLK(clk), .Q(out[86]) );
  DFFX1_HVT \out_reg[85]  ( .D(n90), .CLK(clk), .Q(out[85]) );
  DFFX1_HVT \out_reg[84]  ( .D(n89), .CLK(clk), .Q(out[84]) );
  DFFX1_HVT \out_reg[83]  ( .D(n88), .CLK(clk), .Q(out[83]) );
  DFFX1_HVT \out_reg[82]  ( .D(n87), .CLK(clk), .Q(out[82]) );
  DFFX1_HVT \out_reg[81]  ( .D(n86), .CLK(clk), .Q(out[81]) );
  DFFX1_HVT \out_reg[80]  ( .D(n85), .CLK(clk), .Q(out[80]) );
  DFFX1_HVT \out_reg[79]  ( .D(n84), .CLK(clk), .Q(out[79]) );
  DFFX1_HVT \out_reg[78]  ( .D(n83), .CLK(clk), .Q(out[78]) );
  DFFX1_HVT \out_reg[77]  ( .D(n82), .CLK(clk), .Q(out[77]) );
  DFFX1_HVT \out_reg[76]  ( .D(n81), .CLK(clk), .Q(out[76]) );
  DFFX1_HVT \out_reg[75]  ( .D(n80), .CLK(clk), .Q(out[75]) );
  DFFX1_HVT \out_reg[74]  ( .D(n79), .CLK(clk), .Q(out[74]) );
  DFFX1_HVT \out_reg[73]  ( .D(n78), .CLK(clk), .Q(out[73]) );
  DFFX1_HVT \out_reg[72]  ( .D(n77), .CLK(clk), .Q(out[72]) );
  DFFX1_HVT \out_reg[71]  ( .D(n76), .CLK(clk), .Q(out[71]) );
  DFFX1_HVT \out_reg[70]  ( .D(n75), .CLK(clk), .Q(out[70]) );
  DFFX1_HVT \out_reg[69]  ( .D(n74), .CLK(clk), .Q(out[69]) );
  DFFX1_HVT \out_reg[68]  ( .D(n73), .CLK(clk), .Q(out[68]) );
  DFFX1_HVT \out_reg[67]  ( .D(n72), .CLK(clk), .Q(out[67]) );
  DFFX1_HVT \out_reg[66]  ( .D(n71), .CLK(clk), .Q(out[66]) );
  DFFX1_HVT \out_reg[65]  ( .D(n70), .CLK(clk), .Q(out[65]) );
  DFFX1_HVT \out_reg[64]  ( .D(n69), .CLK(clk), .Q(out[64]) );
  DFFX1_HVT \out_reg[63]  ( .D(n68), .CLK(clk), .Q(out[63]) );
  DFFX1_HVT \out_reg[62]  ( .D(n67), .CLK(clk), .Q(out[62]) );
  DFFX1_HVT \out_reg[61]  ( .D(n66), .CLK(clk), .Q(out[61]) );
  DFFX1_HVT \out_reg[60]  ( .D(n65), .CLK(clk), .Q(out[60]) );
  DFFX1_HVT \out_reg[59]  ( .D(n64), .CLK(clk), .Q(out[59]) );
  DFFX1_HVT \out_reg[58]  ( .D(n63), .CLK(clk), .Q(out[58]) );
  DFFX1_HVT \out_reg[57]  ( .D(n62), .CLK(clk), .Q(out[57]) );
  DFFX1_HVT \out_reg[56]  ( .D(n61), .CLK(clk), .Q(out[56]) );
  DFFX1_HVT \out_reg[55]  ( .D(n60), .CLK(clk), .Q(out[55]) );
  DFFX1_HVT \out_reg[54]  ( .D(n59), .CLK(clk), .Q(out[54]) );
  DFFX1_HVT \out_reg[53]  ( .D(n58), .CLK(clk), .Q(out[53]) );
  DFFX1_HVT \out_reg[52]  ( .D(n57), .CLK(clk), .Q(out[52]) );
  DFFX1_HVT \out_reg[51]  ( .D(n56), .CLK(clk), .Q(out[51]) );
  DFFX1_HVT \out_reg[50]  ( .D(n55), .CLK(clk), .Q(out[50]) );
  DFFX1_HVT \out_reg[49]  ( .D(n54), .CLK(clk), .Q(out[49]) );
  DFFX1_HVT \out_reg[48]  ( .D(n53), .CLK(clk), .Q(out[48]) );
  DFFX1_HVT \out_reg[47]  ( .D(n52), .CLK(clk), .Q(out[47]) );
  DFFX1_HVT \out_reg[46]  ( .D(n51), .CLK(clk), .Q(out[46]) );
  DFFX1_HVT \out_reg[45]  ( .D(n50), .CLK(clk), .Q(out[45]) );
  DFFX1_HVT \out_reg[44]  ( .D(n49), .CLK(clk), .Q(out[44]) );
  DFFX1_HVT \out_reg[43]  ( .D(n48), .CLK(clk), .Q(out[43]) );
  DFFX1_HVT \out_reg[42]  ( .D(n47), .CLK(clk), .Q(out[42]) );
  DFFX1_HVT \out_reg[41]  ( .D(n46), .CLK(clk), .Q(out[41]) );
  DFFX1_HVT \out_reg[40]  ( .D(n45), .CLK(clk), .Q(out[40]) );
  DFFX1_HVT \out_reg[39]  ( .D(n44), .CLK(clk), .Q(out[39]) );
  DFFX1_HVT \out_reg[38]  ( .D(n43), .CLK(clk), .Q(out[38]) );
  DFFX1_HVT \out_reg[37]  ( .D(n42), .CLK(clk), .Q(out[37]) );
  DFFX1_HVT \out_reg[36]  ( .D(n41), .CLK(clk), .Q(out[36]) );
  DFFX1_HVT \out_reg[35]  ( .D(n40), .CLK(clk), .Q(out[35]) );
  DFFX1_HVT \out_reg[34]  ( .D(n39), .CLK(clk), .Q(out[34]) );
  DFFX1_HVT \out_reg[33]  ( .D(n38), .CLK(clk), .Q(out[33]) );
  DFFX1_HVT \out_reg[32]  ( .D(n37), .CLK(clk), .Q(out[32]) );
  DFFX1_HVT \out_reg[31]  ( .D(n36), .CLK(clk), .Q(out[31]) );
  DFFX1_HVT \out_reg[30]  ( .D(n35), .CLK(clk), .Q(out[30]) );
  DFFX1_HVT \out_reg[29]  ( .D(n34), .CLK(clk), .Q(out[29]) );
  DFFX1_HVT \out_reg[28]  ( .D(n33), .CLK(clk), .Q(out[28]) );
  DFFX1_HVT \out_reg[27]  ( .D(n32), .CLK(clk), .Q(out[27]) );
  DFFX1_HVT \out_reg[26]  ( .D(n31), .CLK(clk), .Q(out[26]) );
  DFFX1_HVT \out_reg[25]  ( .D(n30), .CLK(clk), .Q(out[25]) );
  DFFX1_HVT \out_reg[24]  ( .D(n29), .CLK(clk), .Q(out[24]) );
  DFFX1_HVT \out_reg[23]  ( .D(n28), .CLK(clk), .Q(out[23]) );
  DFFX1_HVT \out_reg[22]  ( .D(n27), .CLK(clk), .Q(out[22]) );
  DFFX1_HVT \out_reg[21]  ( .D(n26), .CLK(clk), .Q(out[21]) );
  DFFX1_HVT \out_reg[20]  ( .D(n25), .CLK(clk), .Q(out[20]) );
  DFFX1_HVT \out_reg[19]  ( .D(n24), .CLK(clk), .Q(out[19]) );
  DFFX1_HVT \out_reg[18]  ( .D(n23), .CLK(clk), .Q(out[18]) );
  DFFX1_HVT \out_reg[17]  ( .D(n22), .CLK(clk), .Q(out[17]) );
  DFFX1_HVT \out_reg[16]  ( .D(n21), .CLK(clk), .Q(out[16]) );
  DFFX1_HVT \out_reg[15]  ( .D(n20), .CLK(clk), .Q(out[15]) );
  DFFX1_HVT \out_reg[14]  ( .D(n19), .CLK(clk), .Q(out[14]) );
  DFFX1_HVT \out_reg[13]  ( .D(n18), .CLK(clk), .Q(out[13]) );
  DFFX1_HVT \out_reg[12]  ( .D(n17), .CLK(clk), .Q(out[12]) );
  DFFX1_HVT \out_reg[11]  ( .D(n16), .CLK(clk), .Q(out[11]) );
  DFFX1_HVT \out_reg[10]  ( .D(n15), .CLK(clk), .Q(out[10]) );
  DFFX1_HVT \out_reg[9]  ( .D(n14), .CLK(clk), .Q(out[9]) );
  DFFX1_HVT \out_reg[8]  ( .D(n13), .CLK(clk), .Q(out[8]) );
  DFFX1_HVT \out_reg[7]  ( .D(n12), .CLK(clk), .Q(out[7]) );
  DFFX1_HVT \out_reg[6]  ( .D(n11), .CLK(clk), .Q(out[6]) );
  DFFX1_HVT \out_reg[5]  ( .D(n10), .CLK(clk), .Q(out[5]) );
  DFFX1_HVT \out_reg[4]  ( .D(n9), .CLK(clk), .Q(out[4]) );
  DFFX1_HVT \out_reg[3]  ( .D(n8), .CLK(clk), .Q(out[3]) );
  DFFX1_HVT \out_reg[2]  ( .D(n7), .CLK(clk), .Q(out[2]) );
  DFFX1_HVT \out_reg[1]  ( .D(n6), .CLK(clk), .Q(out[1]) );
  DFFX1_HVT \out_reg[0]  ( .D(n5), .CLK(clk), .Q(out[0]) );
  AO22X1_HVT U4 ( .A1(out[0]), .A2(n143), .A3(in[0]), .A4(n141), .Y(n5) );
  AO22X1_HVT U5 ( .A1(out[1]), .A2(n143), .A3(in[1]), .A4(n141), .Y(n6) );
  AO22X1_HVT U6 ( .A1(out[2]), .A2(n143), .A3(in[2]), .A4(n141), .Y(n7) );
  AO22X1_HVT U7 ( .A1(out[3]), .A2(n143), .A3(in[3]), .A4(n141), .Y(n8) );
  AO22X1_HVT U8 ( .A1(out[4]), .A2(n143), .A3(in[4]), .A4(n141), .Y(n9) );
  AO22X1_HVT U9 ( .A1(out[5]), .A2(n143), .A3(in[5]), .A4(n141), .Y(n10) );
  AO22X1_HVT U10 ( .A1(out[6]), .A2(n143), .A3(in[6]), .A4(n141), .Y(n11) );
  AO22X1_HVT U11 ( .A1(out[7]), .A2(n143), .A3(in[7]), .A4(n141), .Y(n12) );
  AO22X1_HVT U12 ( .A1(out[8]), .A2(n143), .A3(in[8]), .A4(n140), .Y(n13) );
  AO22X1_HVT U13 ( .A1(out[9]), .A2(n143), .A3(in[9]), .A4(n140), .Y(n14) );
  AO22X1_HVT U14 ( .A1(out[10]), .A2(n143), .A3(in[10]), .A4(n140), .Y(n15) );
  AO22X1_HVT U15 ( .A1(out[11]), .A2(n143), .A3(in[11]), .A4(n140), .Y(n16) );
  AO22X1_HVT U16 ( .A1(out[12]), .A2(n144), .A3(in[12]), .A4(n140), .Y(n17) );
  AO22X1_HVT U17 ( .A1(out[13]), .A2(n144), .A3(in[13]), .A4(n140), .Y(n18) );
  AO22X1_HVT U18 ( .A1(out[14]), .A2(n144), .A3(in[14]), .A4(n140), .Y(n19) );
  AO22X1_HVT U19 ( .A1(out[15]), .A2(n144), .A3(in[15]), .A4(n140), .Y(n20) );
  AO22X1_HVT U20 ( .A1(out[16]), .A2(n144), .A3(in[16]), .A4(n140), .Y(n21) );
  AO22X1_HVT U21 ( .A1(out[17]), .A2(n144), .A3(in[17]), .A4(n140), .Y(n22) );
  AO22X1_HVT U22 ( .A1(out[18]), .A2(n144), .A3(in[18]), .A4(n140), .Y(n23) );
  AO22X1_HVT U23 ( .A1(out[19]), .A2(n144), .A3(in[19]), .A4(n140), .Y(n24) );
  AO22X1_HVT U24 ( .A1(out[20]), .A2(n144), .A3(in[20]), .A4(n139), .Y(n25) );
  AO22X1_HVT U25 ( .A1(out[21]), .A2(n144), .A3(in[21]), .A4(n139), .Y(n26) );
  AO22X1_HVT U26 ( .A1(out[22]), .A2(n144), .A3(in[22]), .A4(n139), .Y(n27) );
  AO22X1_HVT U27 ( .A1(out[23]), .A2(n144), .A3(in[23]), .A4(n139), .Y(n28) );
  AO22X1_HVT U28 ( .A1(out[24]), .A2(n145), .A3(in[24]), .A4(n139), .Y(n29) );
  AO22X1_HVT U29 ( .A1(out[25]), .A2(n145), .A3(in[25]), .A4(n139), .Y(n30) );
  AO22X1_HVT U30 ( .A1(out[26]), .A2(n145), .A3(in[26]), .A4(n139), .Y(n31) );
  AO22X1_HVT U31 ( .A1(out[27]), .A2(n145), .A3(in[27]), .A4(n139), .Y(n32) );
  AO22X1_HVT U32 ( .A1(out[28]), .A2(n145), .A3(in[28]), .A4(n139), .Y(n33) );
  AO22X1_HVT U33 ( .A1(out[29]), .A2(n145), .A3(in[29]), .A4(n139), .Y(n34) );
  AO22X1_HVT U34 ( .A1(out[30]), .A2(n145), .A3(in[30]), .A4(n139), .Y(n35) );
  AO22X1_HVT U35 ( .A1(out[31]), .A2(n145), .A3(in[31]), .A4(n139), .Y(n36) );
  AO22X1_HVT U36 ( .A1(out[32]), .A2(n145), .A3(in[32]), .A4(n138), .Y(n37) );
  AO22X1_HVT U37 ( .A1(out[33]), .A2(n145), .A3(in[33]), .A4(n138), .Y(n38) );
  AO22X1_HVT U38 ( .A1(out[34]), .A2(n145), .A3(in[34]), .A4(n138), .Y(n39) );
  AO22X1_HVT U39 ( .A1(out[35]), .A2(n145), .A3(in[35]), .A4(n138), .Y(n40) );
  AO22X1_HVT U40 ( .A1(out[36]), .A2(n146), .A3(in[36]), .A4(n138), .Y(n41) );
  AO22X1_HVT U41 ( .A1(out[37]), .A2(n146), .A3(in[37]), .A4(n138), .Y(n42) );
  AO22X1_HVT U42 ( .A1(out[38]), .A2(n146), .A3(in[38]), .A4(n138), .Y(n43) );
  AO22X1_HVT U43 ( .A1(out[39]), .A2(n146), .A3(in[39]), .A4(n138), .Y(n44) );
  AO22X1_HVT U44 ( .A1(out[40]), .A2(n146), .A3(in[40]), .A4(n138), .Y(n45) );
  AO22X1_HVT U45 ( .A1(out[41]), .A2(n146), .A3(in[41]), .A4(n138), .Y(n46) );
  AO22X1_HVT U46 ( .A1(out[42]), .A2(n146), .A3(in[42]), .A4(n138), .Y(n47) );
  AO22X1_HVT U47 ( .A1(out[43]), .A2(n146), .A3(in[43]), .A4(n138), .Y(n48) );
  AO22X1_HVT U48 ( .A1(out[44]), .A2(n146), .A3(in[44]), .A4(n137), .Y(n49) );
  AO22X1_HVT U49 ( .A1(out[45]), .A2(n146), .A3(in[45]), .A4(n137), .Y(n50) );
  AO22X1_HVT U50 ( .A1(out[46]), .A2(n146), .A3(in[46]), .A4(n137), .Y(n51) );
  AO22X1_HVT U51 ( .A1(out[47]), .A2(n146), .A3(in[47]), .A4(n137), .Y(n52) );
  AO22X1_HVT U52 ( .A1(out[48]), .A2(n147), .A3(in[48]), .A4(n137), .Y(n53) );
  AO22X1_HVT U53 ( .A1(out[49]), .A2(n147), .A3(in[49]), .A4(n137), .Y(n54) );
  AO22X1_HVT U54 ( .A1(out[50]), .A2(n147), .A3(in[50]), .A4(n137), .Y(n55) );
  AO22X1_HVT U55 ( .A1(out[51]), .A2(n147), .A3(in[51]), .A4(n137), .Y(n56) );
  AO22X1_HVT U56 ( .A1(out[52]), .A2(n147), .A3(in[52]), .A4(n137), .Y(n57) );
  AO22X1_HVT U57 ( .A1(out[53]), .A2(n147), .A3(in[53]), .A4(n137), .Y(n58) );
  AO22X1_HVT U58 ( .A1(out[54]), .A2(n147), .A3(in[54]), .A4(n137), .Y(n59) );
  AO22X1_HVT U59 ( .A1(out[55]), .A2(n147), .A3(in[55]), .A4(n137), .Y(n60) );
  AO22X1_HVT U60 ( .A1(out[56]), .A2(n147), .A3(in[56]), .A4(n136), .Y(n61) );
  AO22X1_HVT U61 ( .A1(out[57]), .A2(n147), .A3(in[57]), .A4(n136), .Y(n62) );
  AO22X1_HVT U62 ( .A1(out[58]), .A2(n147), .A3(in[58]), .A4(n136), .Y(n63) );
  AO22X1_HVT U63 ( .A1(out[59]), .A2(n147), .A3(in[59]), .A4(n136), .Y(n64) );
  AO22X1_HVT U64 ( .A1(out[60]), .A2(n148), .A3(in[60]), .A4(n136), .Y(n65) );
  AO22X1_HVT U65 ( .A1(out[61]), .A2(n148), .A3(in[61]), .A4(n136), .Y(n66) );
  AO22X1_HVT U66 ( .A1(out[62]), .A2(n148), .A3(in[62]), .A4(n136), .Y(n67) );
  AO22X1_HVT U67 ( .A1(out[63]), .A2(n148), .A3(in[63]), .A4(n136), .Y(n68) );
  AO22X1_HVT U68 ( .A1(out[64]), .A2(n148), .A3(in[64]), .A4(n136), .Y(n69) );
  AO22X1_HVT U69 ( .A1(out[65]), .A2(n148), .A3(in[65]), .A4(n136), .Y(n70) );
  AO22X1_HVT U70 ( .A1(out[66]), .A2(n148), .A3(in[66]), .A4(n136), .Y(n71) );
  AO22X1_HVT U71 ( .A1(out[67]), .A2(n148), .A3(in[67]), .A4(n136), .Y(n72) );
  AO22X1_HVT U72 ( .A1(out[68]), .A2(n148), .A3(in[68]), .A4(n135), .Y(n73) );
  AO22X1_HVT U73 ( .A1(out[69]), .A2(n148), .A3(in[69]), .A4(n135), .Y(n74) );
  AO22X1_HVT U74 ( .A1(out[70]), .A2(n148), .A3(in[70]), .A4(n135), .Y(n75) );
  AO22X1_HVT U75 ( .A1(out[71]), .A2(n148), .A3(in[71]), .A4(n135), .Y(n76) );
  AO22X1_HVT U76 ( .A1(out[72]), .A2(n149), .A3(in[72]), .A4(n135), .Y(n77) );
  AO22X1_HVT U77 ( .A1(out[73]), .A2(n149), .A3(in[73]), .A4(n135), .Y(n78) );
  AO22X1_HVT U78 ( .A1(out[74]), .A2(n149), .A3(in[74]), .A4(n135), .Y(n79) );
  AO22X1_HVT U79 ( .A1(out[75]), .A2(n149), .A3(in[75]), .A4(n135), .Y(n80) );
  AO22X1_HVT U80 ( .A1(out[76]), .A2(n149), .A3(in[76]), .A4(n135), .Y(n81) );
  AO22X1_HVT U81 ( .A1(out[77]), .A2(n149), .A3(in[77]), .A4(n135), .Y(n82) );
  AO22X1_HVT U82 ( .A1(out[78]), .A2(n149), .A3(in[78]), .A4(n135), .Y(n83) );
  AO22X1_HVT U83 ( .A1(out[79]), .A2(n149), .A3(in[79]), .A4(n135), .Y(n84) );
  AO22X1_HVT U84 ( .A1(out[80]), .A2(n149), .A3(in[80]), .A4(n134), .Y(n85) );
  AO22X1_HVT U85 ( .A1(out[81]), .A2(n149), .A3(in[81]), .A4(n134), .Y(n86) );
  AO22X1_HVT U86 ( .A1(out[82]), .A2(n149), .A3(in[82]), .A4(n134), .Y(n87) );
  AO22X1_HVT U87 ( .A1(out[83]), .A2(n149), .A3(in[83]), .A4(n134), .Y(n88) );
  AO22X1_HVT U88 ( .A1(out[84]), .A2(n150), .A3(in[84]), .A4(n134), .Y(n89) );
  AO22X1_HVT U89 ( .A1(out[85]), .A2(n150), .A3(in[85]), .A4(n134), .Y(n90) );
  AO22X1_HVT U90 ( .A1(out[86]), .A2(n150), .A3(in[86]), .A4(n134), .Y(n91) );
  AO22X1_HVT U91 ( .A1(out[87]), .A2(n150), .A3(in[87]), .A4(n134), .Y(n92) );
  AO22X1_HVT U92 ( .A1(out[88]), .A2(n150), .A3(in[88]), .A4(n134), .Y(n93) );
  AO22X1_HVT U93 ( .A1(out[89]), .A2(n150), .A3(in[89]), .A4(n134), .Y(n94) );
  AO22X1_HVT U94 ( .A1(out[90]), .A2(n150), .A3(in[90]), .A4(n134), .Y(n95) );
  AO22X1_HVT U95 ( .A1(out[91]), .A2(n150), .A3(in[91]), .A4(n134), .Y(n96) );
  AO22X1_HVT U96 ( .A1(out[92]), .A2(n150), .A3(in[92]), .A4(n133), .Y(n97) );
  AO22X1_HVT U97 ( .A1(out[93]), .A2(n150), .A3(in[93]), .A4(n133), .Y(n98) );
  AO22X1_HVT U98 ( .A1(out[94]), .A2(n150), .A3(in[94]), .A4(n133), .Y(n99) );
  AO22X1_HVT U99 ( .A1(out[95]), .A2(n150), .A3(in[95]), .A4(n133), .Y(n100)
         );
  AO22X1_HVT U100 ( .A1(out[96]), .A2(n151), .A3(in[96]), .A4(n133), .Y(n101)
         );
  AO22X1_HVT U101 ( .A1(out[97]), .A2(n151), .A3(in[97]), .A4(n133), .Y(n102)
         );
  AO22X1_HVT U102 ( .A1(out[98]), .A2(n151), .A3(in[98]), .A4(n133), .Y(n103)
         );
  AO22X1_HVT U103 ( .A1(out[99]), .A2(n151), .A3(in[99]), .A4(n133), .Y(n104)
         );
  AO22X1_HVT U104 ( .A1(out[100]), .A2(n151), .A3(in[100]), .A4(n133), .Y(n105) );
  AO22X1_HVT U105 ( .A1(out[101]), .A2(n151), .A3(in[101]), .A4(n133), .Y(n106) );
  AO22X1_HVT U106 ( .A1(out[102]), .A2(n151), .A3(in[102]), .A4(n133), .Y(n107) );
  AO22X1_HVT U107 ( .A1(out[103]), .A2(n151), .A3(in[103]), .A4(n133), .Y(n108) );
  AO22X1_HVT U108 ( .A1(out[104]), .A2(n151), .A3(in[104]), .A4(n2), .Y(n109)
         );
  AO22X1_HVT U109 ( .A1(out[105]), .A2(n151), .A3(in[105]), .A4(n2), .Y(n110)
         );
  AO22X1_HVT U110 ( .A1(out[106]), .A2(n151), .A3(in[106]), .A4(n2), .Y(n111)
         );
  AO22X1_HVT U111 ( .A1(out[107]), .A2(n151), .A3(in[107]), .A4(n2), .Y(n112)
         );
  AO22X1_HVT U112 ( .A1(out[108]), .A2(n152), .A3(in[108]), .A4(n2), .Y(n113)
         );
  AO22X1_HVT U113 ( .A1(out[109]), .A2(n152), .A3(in[109]), .A4(n2), .Y(n114)
         );
  AO22X1_HVT U114 ( .A1(out[110]), .A2(n152), .A3(in[110]), .A4(n2), .Y(n115)
         );
  AO22X1_HVT U115 ( .A1(out[111]), .A2(n152), .A3(in[111]), .A4(n2), .Y(n116)
         );
  AO22X1_HVT U116 ( .A1(out[112]), .A2(n152), .A3(in[112]), .A4(n2), .Y(n117)
         );
  AO22X1_HVT U117 ( .A1(out[113]), .A2(n152), .A3(in[113]), .A4(n2), .Y(n118)
         );
  AO22X1_HVT U118 ( .A1(out[114]), .A2(n152), .A3(in[114]), .A4(n2), .Y(n119)
         );
  AO22X1_HVT U119 ( .A1(out[115]), .A2(n152), .A3(in[115]), .A4(n2), .Y(n120)
         );
  AO22X1_HVT U120 ( .A1(out[116]), .A2(n152), .A3(in[116]), .A4(n1), .Y(n121)
         );
  AO22X1_HVT U121 ( .A1(out[117]), .A2(n152), .A3(in[117]), .A4(n1), .Y(n122)
         );
  AO22X1_HVT U122 ( .A1(out[118]), .A2(n152), .A3(in[118]), .A4(n1), .Y(n123)
         );
  AO22X1_HVT U123 ( .A1(out[119]), .A2(n152), .A3(in[119]), .A4(n1), .Y(n124)
         );
  AO22X1_HVT U124 ( .A1(out[120]), .A2(n153), .A3(in[120]), .A4(n1), .Y(n125)
         );
  AO22X1_HVT U125 ( .A1(out[121]), .A2(n153), .A3(in[121]), .A4(n1), .Y(n126)
         );
  AO22X1_HVT U126 ( .A1(out[122]), .A2(n153), .A3(in[122]), .A4(n1), .Y(n127)
         );
  AO22X1_HVT U127 ( .A1(out[123]), .A2(n153), .A3(in[123]), .A4(n1), .Y(n128)
         );
  AO22X1_HVT U128 ( .A1(out[124]), .A2(n153), .A3(in[124]), .A4(n1), .Y(n129)
         );
  AO22X1_HVT U129 ( .A1(out[125]), .A2(n153), .A3(in[125]), .A4(n1), .Y(n130)
         );
  AO22X1_HVT U130 ( .A1(out[126]), .A2(n153), .A3(in[126]), .A4(n1), .Y(n131)
         );
  AO22X1_HVT U131 ( .A1(out[127]), .A2(n153), .A3(in[127]), .A4(n1), .Y(n132)
         );
  AND2X1_HVT U132 ( .A1(n156), .A2(n4), .Y(n3) );
  NAND2X0_HVT U133 ( .A1(enable), .A2(n156), .Y(n4) );
  INVX0_HVT U2 ( .A(n154), .Y(n153) );
  INVX1_HVT U3 ( .A(n133), .Y(n142) );
  INVX0_HVT U134 ( .A(n3), .Y(n155) );
  INVX1_HVT U135 ( .A(n142), .Y(n139) );
  INVX1_HVT U136 ( .A(n142), .Y(n138) );
  INVX1_HVT U137 ( .A(n142), .Y(n137) );
  INVX1_HVT U138 ( .A(n142), .Y(n136) );
  INVX1_HVT U139 ( .A(n142), .Y(n134) );
  INVX1_HVT U140 ( .A(n4), .Y(n133) );
  INVX1_HVT U141 ( .A(n4), .Y(n2) );
  INVX1_HVT U142 ( .A(n4), .Y(n1) );
  INVX1_HVT U143 ( .A(n142), .Y(n141) );
  INVX1_HVT U144 ( .A(n142), .Y(n140) );
  INVX1_HVT U145 ( .A(n4), .Y(n135) );
  INVX1_HVT U146 ( .A(n155), .Y(n143) );
  INVX1_HVT U147 ( .A(n155), .Y(n144) );
  INVX1_HVT U148 ( .A(n155), .Y(n145) );
  INVX1_HVT U149 ( .A(n155), .Y(n146) );
  INVX1_HVT U150 ( .A(n154), .Y(n148) );
  INVX1_HVT U151 ( .A(n154), .Y(n149) );
  INVX1_HVT U152 ( .A(n154), .Y(n150) );
  INVX1_HVT U153 ( .A(n154), .Y(n151) );
  INVX1_HVT U154 ( .A(n154), .Y(n152) );
  INVX1_HVT U155 ( .A(n155), .Y(n147) );
  INVX1_HVT U156 ( .A(n3), .Y(n154) );
  INVX0_HVT U157 ( .A(rst), .Y(n156) );
endmodule

