
module inv_round ( in, last, keyin, out );
  input [127:0] in;
  input [127:0] keyin;
  output [127:0] out;
  input last;

  wire   [127:0] sr_out;
  wire   [127:0] sb_out;
  wire   [127:0] oout;
  wire   [127:0] mc_out;

  inv_shift_rows sr ( .in(in), .out(sr_out) );
  inv_subbytes sb ( .in(sr_out), .out(sb_out) );
  inv_add_round_keys adk ( .state(sb_out), .subkey(keyin), .out(oout) );
  inv_Mix_Column mc ( .in(oout), .out1(mc_out) );
  MUX21X1_HVT U1 ( .A1(mc_out[9]), .A2(oout[9]), .S0(last), .Y(out[9]) );
  MUX21X1_HVT U2 ( .A1(mc_out[99]), .A2(oout[99]), .S0(last), .Y(out[99]) );
  MUX21X1_HVT U3 ( .A1(mc_out[98]), .A2(oout[98]), .S0(last), .Y(out[98]) );
  MUX21X1_HVT U4 ( .A1(mc_out[97]), .A2(oout[97]), .S0(last), .Y(out[97]) );
  MUX21X1_HVT U5 ( .A1(mc_out[96]), .A2(oout[96]), .S0(last), .Y(out[96]) );
  MUX21X1_HVT U6 ( .A1(mc_out[95]), .A2(oout[95]), .S0(last), .Y(out[95]) );
  MUX21X1_HVT U7 ( .A1(mc_out[94]), .A2(oout[94]), .S0(last), .Y(out[94]) );
  MUX21X1_HVT U8 ( .A1(mc_out[93]), .A2(oout[93]), .S0(last), .Y(out[93]) );
  MUX21X1_HVT U9 ( .A1(mc_out[92]), .A2(oout[92]), .S0(last), .Y(out[92]) );
  MUX21X1_HVT U10 ( .A1(mc_out[91]), .A2(oout[91]), .S0(last), .Y(out[91]) );
  MUX21X1_HVT U11 ( .A1(mc_out[90]), .A2(oout[90]), .S0(last), .Y(out[90]) );
  MUX21X1_HVT U12 ( .A1(mc_out[8]), .A2(oout[8]), .S0(last), .Y(out[8]) );
  MUX21X1_HVT U13 ( .A1(mc_out[89]), .A2(oout[89]), .S0(last), .Y(out[89]) );
  MUX21X1_HVT U14 ( .A1(mc_out[88]), .A2(oout[88]), .S0(last), .Y(out[88]) );
  MUX21X1_HVT U15 ( .A1(mc_out[87]), .A2(oout[87]), .S0(last), .Y(out[87]) );
  MUX21X1_HVT U16 ( .A1(mc_out[86]), .A2(oout[86]), .S0(last), .Y(out[86]) );
  MUX21X1_HVT U17 ( .A1(mc_out[85]), .A2(oout[85]), .S0(last), .Y(out[85]) );
  MUX21X1_HVT U18 ( .A1(mc_out[84]), .A2(oout[84]), .S0(last), .Y(out[84]) );
  MUX21X1_HVT U19 ( .A1(mc_out[83]), .A2(oout[83]), .S0(last), .Y(out[83]) );
  MUX21X1_HVT U20 ( .A1(mc_out[82]), .A2(oout[82]), .S0(last), .Y(out[82]) );
  MUX21X1_HVT U21 ( .A1(mc_out[81]), .A2(oout[81]), .S0(last), .Y(out[81]) );
  MUX21X1_HVT U22 ( .A1(mc_out[80]), .A2(oout[80]), .S0(last), .Y(out[80]) );
  MUX21X1_HVT U23 ( .A1(mc_out[7]), .A2(oout[7]), .S0(last), .Y(out[7]) );
  MUX21X1_HVT U24 ( .A1(mc_out[79]), .A2(oout[79]), .S0(last), .Y(out[79]) );
  MUX21X1_HVT U25 ( .A1(mc_out[78]), .A2(oout[78]), .S0(last), .Y(out[78]) );
  MUX21X1_HVT U26 ( .A1(mc_out[77]), .A2(oout[77]), .S0(last), .Y(out[77]) );
  MUX21X1_HVT U27 ( .A1(mc_out[76]), .A2(oout[76]), .S0(last), .Y(out[76]) );
  MUX21X1_HVT U28 ( .A1(mc_out[75]), .A2(oout[75]), .S0(last), .Y(out[75]) );
  MUX21X1_HVT U29 ( .A1(mc_out[74]), .A2(oout[74]), .S0(last), .Y(out[74]) );
  MUX21X1_HVT U30 ( .A1(mc_out[73]), .A2(oout[73]), .S0(last), .Y(out[73]) );
  MUX21X1_HVT U31 ( .A1(mc_out[72]), .A2(oout[72]), .S0(last), .Y(out[72]) );
  MUX21X1_HVT U32 ( .A1(mc_out[71]), .A2(oout[71]), .S0(last), .Y(out[71]) );
  MUX21X1_HVT U33 ( .A1(mc_out[70]), .A2(oout[70]), .S0(last), .Y(out[70]) );
  MUX21X1_HVT U34 ( .A1(mc_out[6]), .A2(oout[6]), .S0(last), .Y(out[6]) );
  MUX21X1_HVT U35 ( .A1(mc_out[69]), .A2(oout[69]), .S0(last), .Y(out[69]) );
  MUX21X1_HVT U36 ( .A1(mc_out[68]), .A2(oout[68]), .S0(last), .Y(out[68]) );
  MUX21X1_HVT U37 ( .A1(mc_out[67]), .A2(oout[67]), .S0(last), .Y(out[67]) );
  MUX21X1_HVT U38 ( .A1(mc_out[66]), .A2(oout[66]), .S0(last), .Y(out[66]) );
  MUX21X1_HVT U39 ( .A1(mc_out[65]), .A2(oout[65]), .S0(last), .Y(out[65]) );
  MUX21X1_HVT U40 ( .A1(mc_out[64]), .A2(oout[64]), .S0(last), .Y(out[64]) );
  MUX21X1_HVT U41 ( .A1(mc_out[63]), .A2(oout[63]), .S0(last), .Y(out[63]) );
  MUX21X1_HVT U42 ( .A1(mc_out[62]), .A2(oout[62]), .S0(last), .Y(out[62]) );
  MUX21X1_HVT U43 ( .A1(mc_out[61]), .A2(oout[61]), .S0(last), .Y(out[61]) );
  MUX21X1_HVT U44 ( .A1(mc_out[60]), .A2(oout[60]), .S0(last), .Y(out[60]) );
  MUX21X1_HVT U45 ( .A1(mc_out[5]), .A2(oout[5]), .S0(last), .Y(out[5]) );
  MUX21X1_HVT U46 ( .A1(mc_out[59]), .A2(oout[59]), .S0(last), .Y(out[59]) );
  MUX21X1_HVT U47 ( .A1(mc_out[58]), .A2(oout[58]), .S0(last), .Y(out[58]) );
  MUX21X1_HVT U48 ( .A1(mc_out[57]), .A2(oout[57]), .S0(last), .Y(out[57]) );
  MUX21X1_HVT U49 ( .A1(mc_out[56]), .A2(oout[56]), .S0(last), .Y(out[56]) );
  MUX21X1_HVT U50 ( .A1(mc_out[55]), .A2(oout[55]), .S0(last), .Y(out[55]) );
  MUX21X1_HVT U51 ( .A1(mc_out[54]), .A2(oout[54]), .S0(last), .Y(out[54]) );
  MUX21X1_HVT U52 ( .A1(mc_out[53]), .A2(oout[53]), .S0(last), .Y(out[53]) );
  MUX21X1_HVT U53 ( .A1(mc_out[52]), .A2(oout[52]), .S0(last), .Y(out[52]) );
  MUX21X1_HVT U54 ( .A1(mc_out[51]), .A2(oout[51]), .S0(last), .Y(out[51]) );
  MUX21X1_HVT U55 ( .A1(mc_out[50]), .A2(oout[50]), .S0(last), .Y(out[50]) );
  MUX21X1_HVT U56 ( .A1(mc_out[4]), .A2(oout[4]), .S0(last), .Y(out[4]) );
  MUX21X1_HVT U57 ( .A1(mc_out[49]), .A2(oout[49]), .S0(last), .Y(out[49]) );
  MUX21X1_HVT U58 ( .A1(mc_out[48]), .A2(oout[48]), .S0(last), .Y(out[48]) );
  MUX21X1_HVT U59 ( .A1(mc_out[47]), .A2(oout[47]), .S0(last), .Y(out[47]) );
  MUX21X1_HVT U60 ( .A1(mc_out[46]), .A2(oout[46]), .S0(last), .Y(out[46]) );
  MUX21X1_HVT U61 ( .A1(mc_out[45]), .A2(oout[45]), .S0(last), .Y(out[45]) );
  MUX21X1_HVT U62 ( .A1(mc_out[44]), .A2(oout[44]), .S0(last), .Y(out[44]) );
  MUX21X1_HVT U63 ( .A1(mc_out[43]), .A2(oout[43]), .S0(last), .Y(out[43]) );
  MUX21X1_HVT U64 ( .A1(mc_out[42]), .A2(oout[42]), .S0(last), .Y(out[42]) );
  MUX21X1_HVT U65 ( .A1(mc_out[41]), .A2(oout[41]), .S0(last), .Y(out[41]) );
  MUX21X1_HVT U66 ( .A1(mc_out[40]), .A2(oout[40]), .S0(last), .Y(out[40]) );
  MUX21X1_HVT U67 ( .A1(mc_out[3]), .A2(oout[3]), .S0(last), .Y(out[3]) );
  MUX21X1_HVT U68 ( .A1(mc_out[39]), .A2(oout[39]), .S0(last), .Y(out[39]) );
  MUX21X1_HVT U69 ( .A1(mc_out[38]), .A2(oout[38]), .S0(last), .Y(out[38]) );
  MUX21X1_HVT U70 ( .A1(mc_out[37]), .A2(oout[37]), .S0(last), .Y(out[37]) );
  MUX21X1_HVT U71 ( .A1(mc_out[36]), .A2(oout[36]), .S0(last), .Y(out[36]) );
  MUX21X1_HVT U72 ( .A1(mc_out[35]), .A2(oout[35]), .S0(last), .Y(out[35]) );
  MUX21X1_HVT U73 ( .A1(mc_out[34]), .A2(oout[34]), .S0(last), .Y(out[34]) );
  MUX21X1_HVT U74 ( .A1(mc_out[33]), .A2(oout[33]), .S0(last), .Y(out[33]) );
  MUX21X1_HVT U75 ( .A1(mc_out[32]), .A2(oout[32]), .S0(last), .Y(out[32]) );
  MUX21X1_HVT U76 ( .A1(mc_out[31]), .A2(oout[31]), .S0(last), .Y(out[31]) );
  MUX21X1_HVT U77 ( .A1(mc_out[30]), .A2(oout[30]), .S0(last), .Y(out[30]) );
  MUX21X1_HVT U78 ( .A1(mc_out[2]), .A2(oout[2]), .S0(last), .Y(out[2]) );
  MUX21X1_HVT U79 ( .A1(mc_out[29]), .A2(oout[29]), .S0(last), .Y(out[29]) );
  MUX21X1_HVT U80 ( .A1(mc_out[28]), .A2(oout[28]), .S0(last), .Y(out[28]) );
  MUX21X1_HVT U81 ( .A1(mc_out[27]), .A2(oout[27]), .S0(last), .Y(out[27]) );
  MUX21X1_HVT U82 ( .A1(mc_out[26]), .A2(oout[26]), .S0(last), .Y(out[26]) );
  MUX21X1_HVT U83 ( .A1(mc_out[25]), .A2(oout[25]), .S0(last), .Y(out[25]) );
  MUX21X1_HVT U84 ( .A1(mc_out[24]), .A2(oout[24]), .S0(last), .Y(out[24]) );
  MUX21X1_HVT U85 ( .A1(mc_out[23]), .A2(oout[23]), .S0(last), .Y(out[23]) );
  MUX21X1_HVT U86 ( .A1(mc_out[22]), .A2(oout[22]), .S0(last), .Y(out[22]) );
  MUX21X1_HVT U87 ( .A1(mc_out[21]), .A2(oout[21]), .S0(last), .Y(out[21]) );
  MUX21X1_HVT U88 ( .A1(mc_out[20]), .A2(oout[20]), .S0(last), .Y(out[20]) );
  MUX21X1_HVT U89 ( .A1(mc_out[1]), .A2(oout[1]), .S0(last), .Y(out[1]) );
  MUX21X1_HVT U90 ( .A1(mc_out[19]), .A2(oout[19]), .S0(last), .Y(out[19]) );
  MUX21X1_HVT U91 ( .A1(mc_out[18]), .A2(oout[18]), .S0(last), .Y(out[18]) );
  MUX21X1_HVT U92 ( .A1(mc_out[17]), .A2(oout[17]), .S0(last), .Y(out[17]) );
  MUX21X1_HVT U93 ( .A1(mc_out[16]), .A2(oout[16]), .S0(last), .Y(out[16]) );
  MUX21X1_HVT U94 ( .A1(mc_out[15]), .A2(oout[15]), .S0(last), .Y(out[15]) );
  MUX21X1_HVT U95 ( .A1(mc_out[14]), .A2(oout[14]), .S0(last), .Y(out[14]) );
  MUX21X1_HVT U96 ( .A1(mc_out[13]), .A2(oout[13]), .S0(last), .Y(out[13]) );
  MUX21X1_HVT U97 ( .A1(mc_out[12]), .A2(oout[12]), .S0(last), .Y(out[12]) );
  MUX21X1_HVT U98 ( .A1(mc_out[127]), .A2(oout[127]), .S0(last), .Y(out[127])
         );
  MUX21X1_HVT U99 ( .A1(mc_out[126]), .A2(oout[126]), .S0(last), .Y(out[126])
         );
  MUX21X1_HVT U100 ( .A1(mc_out[125]), .A2(oout[125]), .S0(last), .Y(out[125])
         );
  MUX21X1_HVT U101 ( .A1(mc_out[124]), .A2(oout[124]), .S0(last), .Y(out[124])
         );
  MUX21X1_HVT U102 ( .A1(mc_out[123]), .A2(oout[123]), .S0(last), .Y(out[123])
         );
  MUX21X1_HVT U103 ( .A1(mc_out[122]), .A2(oout[122]), .S0(last), .Y(out[122])
         );
  MUX21X1_HVT U104 ( .A1(mc_out[121]), .A2(oout[121]), .S0(last), .Y(out[121])
         );
  MUX21X1_HVT U105 ( .A1(mc_out[120]), .A2(oout[120]), .S0(last), .Y(out[120])
         );
  MUX21X1_HVT U106 ( .A1(mc_out[11]), .A2(oout[11]), .S0(last), .Y(out[11]) );
  MUX21X1_HVT U107 ( .A1(mc_out[119]), .A2(oout[119]), .S0(last), .Y(out[119])
         );
  MUX21X1_HVT U108 ( .A1(mc_out[118]), .A2(oout[118]), .S0(last), .Y(out[118])
         );
  MUX21X1_HVT U109 ( .A1(mc_out[117]), .A2(oout[117]), .S0(last), .Y(out[117])
         );
  MUX21X1_HVT U110 ( .A1(mc_out[116]), .A2(oout[116]), .S0(last), .Y(out[116])
         );
  MUX21X1_HVT U111 ( .A1(mc_out[115]), .A2(oout[115]), .S0(last), .Y(out[115])
         );
  MUX21X1_HVT U112 ( .A1(mc_out[114]), .A2(oout[114]), .S0(last), .Y(out[114])
         );
  MUX21X1_HVT U113 ( .A1(mc_out[113]), .A2(oout[113]), .S0(last), .Y(out[113])
         );
  MUX21X1_HVT U114 ( .A1(mc_out[112]), .A2(oout[112]), .S0(last), .Y(out[112])
         );
  MUX21X1_HVT U115 ( .A1(mc_out[111]), .A2(oout[111]), .S0(last), .Y(out[111])
         );
  MUX21X1_HVT U116 ( .A1(mc_out[110]), .A2(oout[110]), .S0(last), .Y(out[110])
         );
  MUX21X1_HVT U117 ( .A1(mc_out[10]), .A2(oout[10]), .S0(last), .Y(out[10]) );
  MUX21X1_HVT U118 ( .A1(mc_out[109]), .A2(oout[109]), .S0(last), .Y(out[109])
         );
  MUX21X1_HVT U119 ( .A1(mc_out[108]), .A2(oout[108]), .S0(last), .Y(out[108])
         );
  MUX21X1_HVT U120 ( .A1(mc_out[107]), .A2(oout[107]), .S0(last), .Y(out[107])
         );
  MUX21X1_HVT U121 ( .A1(mc_out[106]), .A2(oout[106]), .S0(last), .Y(out[106])
         );
  MUX21X1_HVT U122 ( .A1(mc_out[105]), .A2(oout[105]), .S0(last), .Y(out[105])
         );
  MUX21X1_HVT U123 ( .A1(mc_out[104]), .A2(oout[104]), .S0(last), .Y(out[104])
         );
  MUX21X1_HVT U124 ( .A1(mc_out[103]), .A2(oout[103]), .S0(last), .Y(out[103])
         );
  MUX21X1_HVT U125 ( .A1(mc_out[102]), .A2(oout[102]), .S0(last), .Y(out[102])
         );
  MUX21X1_HVT U126 ( .A1(mc_out[101]), .A2(oout[101]), .S0(last), .Y(out[101])
         );
  MUX21X1_HVT U127 ( .A1(mc_out[100]), .A2(oout[100]), .S0(last), .Y(out[100])
         );
  MUX21X1_HVT U128 ( .A1(mc_out[0]), .A2(oout[0]), .S0(last), .Y(out[0]) );
endmodule

