
module ram_dp_DATA_WIDTH4_ADDR_WIDTH4_0 ( clk, rst, write, a_addr, a_din, 
        b_din, b_dout );
  input [3:0] a_addr;
  input [3:0] a_din;
  input [3:0] b_din;
  output [15:0] b_dout;
  input clk, rst, write;
  wire   N17, N18, N19, N20, \mem[15][15] , \mem[15][14] , \mem[15][13] ,
         \mem[15][12] , \mem[15][11] , \mem[15][10] , \mem[15][9] ,
         \mem[15][8] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][15] ,
         \mem[14][14] , \mem[14][13] , \mem[14][12] , \mem[14][11] ,
         \mem[14][10] , \mem[14][9] , \mem[14][8] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][15] , \mem[13][14] , \mem[13][13] ,
         \mem[13][12] , \mem[13][11] , \mem[13][10] , \mem[13][9] ,
         \mem[13][8] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][15] ,
         \mem[12][14] , \mem[12][13] , \mem[12][12] , \mem[12][11] ,
         \mem[12][10] , \mem[12][9] , \mem[12][8] , \mem[12][7] , \mem[12][6] ,
         \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] , \mem[12][1] ,
         \mem[12][0] , \mem[11][15] , \mem[11][14] , \mem[11][13] ,
         \mem[11][12] , \mem[11][11] , \mem[11][10] , \mem[11][9] ,
         \mem[11][8] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][15] , \mem[9][14] , \mem[9][13] , \mem[9][12] ,
         \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] , \mem[9][7] ,
         \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] ,
         \mem[9][1] , \mem[9][0] , \mem[8][15] , \mem[8][14] , \mem[8][13] ,
         \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] , \mem[8][8] ,
         \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] , \mem[8][3] ,
         \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][15] , \mem[7][14] ,
         \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] ,
         \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][15] ,
         \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] ,
         \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][15] , \mem[3][14] , \mem[3][13] ,
         \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] ,
         \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] ,
         \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][15] ,
         \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N539, N540, N541, N542, N543, N544, N545, N546, N547,
         N548, N549, N550, N551, N552, N553, N554, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123;
  assign N17 = b_din[0];
  assign N18 = b_din[1];
  assign N19 = b_din[2];
  assign N20 = b_din[3];

  DFFNX1_HVT \b_dout_reg[15]  ( .D(N539), .CLK(clk), .Q(b_dout[15]) );
  DFFNX1_HVT \b_dout_reg[14]  ( .D(N540), .CLK(clk), .Q(b_dout[14]) );
  DFFNX1_HVT \b_dout_reg[13]  ( .D(N541), .CLK(clk), .Q(b_dout[13]) );
  DFFNX1_HVT \b_dout_reg[12]  ( .D(N542), .CLK(clk), .Q(b_dout[12]) );
  DFFNX1_HVT \b_dout_reg[11]  ( .D(N543), .CLK(clk), .Q(b_dout[11]) );
  DFFNX1_HVT \b_dout_reg[10]  ( .D(N544), .CLK(clk), .Q(b_dout[10]) );
  DFFNX1_HVT \b_dout_reg[9]  ( .D(N545), .CLK(clk), .Q(b_dout[9]) );
  DFFNX1_HVT \b_dout_reg[8]  ( .D(N546), .CLK(clk), .Q(b_dout[8]) );
  DFFNX1_HVT \b_dout_reg[7]  ( .D(N547), .CLK(clk), .Q(b_dout[7]) );
  DFFNX1_HVT \b_dout_reg[6]  ( .D(N548), .CLK(clk), .Q(b_dout[6]) );
  DFFNX1_HVT \b_dout_reg[5]  ( .D(N549), .CLK(clk), .Q(b_dout[5]) );
  DFFNX1_HVT \b_dout_reg[4]  ( .D(N550), .CLK(clk), .Q(b_dout[4]) );
  DFFNX1_HVT \b_dout_reg[3]  ( .D(N551), .CLK(clk), .Q(b_dout[3]) );
  DFFNX1_HVT \b_dout_reg[2]  ( .D(N552), .CLK(clk), .Q(b_dout[2]) );
  DFFNX1_HVT \b_dout_reg[1]  ( .D(N553), .CLK(clk), .Q(b_dout[1]) );
  DFFNX1_HVT \b_dout_reg[0]  ( .D(N554), .CLK(clk), .Q(b_dout[0]) );
  DFFNX1_HVT \mem_reg[15][15]  ( .D(n825), .CLK(clk), .Q(\mem[15][15] ) );
  DFFNX1_HVT \mem_reg[15][14]  ( .D(n824), .CLK(clk), .Q(\mem[15][14] ) );
  DFFNX1_HVT \mem_reg[15][13]  ( .D(n823), .CLK(clk), .Q(\mem[15][13] ) );
  DFFNX1_HVT \mem_reg[15][12]  ( .D(n822), .CLK(clk), .Q(\mem[15][12] ) );
  DFFNX1_HVT \mem_reg[15][11]  ( .D(n821), .CLK(clk), .Q(\mem[15][11] ) );
  DFFNX1_HVT \mem_reg[15][10]  ( .D(n820), .CLK(clk), .Q(\mem[15][10] ) );
  DFFNX1_HVT \mem_reg[15][9]  ( .D(n819), .CLK(clk), .Q(\mem[15][9] ) );
  DFFNX1_HVT \mem_reg[15][8]  ( .D(n818), .CLK(clk), .Q(\mem[15][8] ) );
  DFFNX1_HVT \mem_reg[15][7]  ( .D(n817), .CLK(clk), .Q(\mem[15][7] ) );
  DFFNX1_HVT \mem_reg[15][6]  ( .D(n816), .CLK(clk), .Q(\mem[15][6] ) );
  DFFNX1_HVT \mem_reg[15][5]  ( .D(n815), .CLK(clk), .Q(\mem[15][5] ) );
  DFFNX1_HVT \mem_reg[15][4]  ( .D(n814), .CLK(clk), .Q(\mem[15][4] ) );
  DFFNX1_HVT \mem_reg[15][3]  ( .D(n813), .CLK(clk), .Q(\mem[15][3] ) );
  DFFNX1_HVT \mem_reg[15][2]  ( .D(n812), .CLK(clk), .Q(\mem[15][2] ) );
  DFFNX1_HVT \mem_reg[15][1]  ( .D(n811), .CLK(clk), .Q(\mem[15][1] ) );
  DFFNX1_HVT \mem_reg[15][0]  ( .D(n810), .CLK(clk), .Q(\mem[15][0] ) );
  DFFNX1_HVT \mem_reg[14][15]  ( .D(n809), .CLK(clk), .Q(\mem[14][15] ) );
  DFFNX1_HVT \mem_reg[14][14]  ( .D(n808), .CLK(clk), .Q(\mem[14][14] ) );
  DFFNX1_HVT \mem_reg[14][13]  ( .D(n807), .CLK(clk), .Q(\mem[14][13] ) );
  DFFNX1_HVT \mem_reg[14][12]  ( .D(n806), .CLK(clk), .Q(\mem[14][12] ) );
  DFFNX1_HVT \mem_reg[14][11]  ( .D(n805), .CLK(clk), .Q(\mem[14][11] ) );
  DFFNX1_HVT \mem_reg[14][10]  ( .D(n804), .CLK(clk), .Q(\mem[14][10] ) );
  DFFNX1_HVT \mem_reg[14][9]  ( .D(n803), .CLK(clk), .Q(\mem[14][9] ) );
  DFFNX1_HVT \mem_reg[14][8]  ( .D(n802), .CLK(clk), .Q(\mem[14][8] ) );
  DFFNX1_HVT \mem_reg[14][7]  ( .D(n801), .CLK(clk), .Q(\mem[14][7] ) );
  DFFNX1_HVT \mem_reg[14][6]  ( .D(n800), .CLK(clk), .Q(\mem[14][6] ) );
  DFFNX1_HVT \mem_reg[14][5]  ( .D(n799), .CLK(clk), .Q(\mem[14][5] ) );
  DFFNX1_HVT \mem_reg[14][4]  ( .D(n798), .CLK(clk), .Q(\mem[14][4] ) );
  DFFNX1_HVT \mem_reg[14][3]  ( .D(n797), .CLK(clk), .Q(\mem[14][3] ) );
  DFFNX1_HVT \mem_reg[14][2]  ( .D(n796), .CLK(clk), .Q(\mem[14][2] ) );
  DFFNX1_HVT \mem_reg[14][1]  ( .D(n795), .CLK(clk), .Q(\mem[14][1] ) );
  DFFNX1_HVT \mem_reg[14][0]  ( .D(n794), .CLK(clk), .Q(\mem[14][0] ) );
  DFFNX1_HVT \mem_reg[13][15]  ( .D(n793), .CLK(clk), .Q(\mem[13][15] ) );
  DFFNX1_HVT \mem_reg[13][14]  ( .D(n792), .CLK(clk), .Q(\mem[13][14] ) );
  DFFNX1_HVT \mem_reg[13][13]  ( .D(n791), .CLK(clk), .Q(\mem[13][13] ) );
  DFFNX1_HVT \mem_reg[13][12]  ( .D(n790), .CLK(clk), .Q(\mem[13][12] ) );
  DFFNX1_HVT \mem_reg[13][11]  ( .D(n789), .CLK(clk), .Q(\mem[13][11] ) );
  DFFNX1_HVT \mem_reg[13][10]  ( .D(n788), .CLK(clk), .Q(\mem[13][10] ) );
  DFFNX1_HVT \mem_reg[13][9]  ( .D(n787), .CLK(clk), .Q(\mem[13][9] ) );
  DFFNX1_HVT \mem_reg[13][8]  ( .D(n786), .CLK(clk), .Q(\mem[13][8] ) );
  DFFNX1_HVT \mem_reg[13][7]  ( .D(n785), .CLK(clk), .Q(\mem[13][7] ) );
  DFFNX1_HVT \mem_reg[13][6]  ( .D(n784), .CLK(clk), .Q(\mem[13][6] ) );
  DFFNX1_HVT \mem_reg[13][5]  ( .D(n783), .CLK(clk), .Q(\mem[13][5] ) );
  DFFNX1_HVT \mem_reg[13][4]  ( .D(n782), .CLK(clk), .Q(\mem[13][4] ) );
  DFFNX1_HVT \mem_reg[13][3]  ( .D(n781), .CLK(clk), .Q(\mem[13][3] ) );
  DFFNX1_HVT \mem_reg[13][2]  ( .D(n780), .CLK(clk), .Q(\mem[13][2] ) );
  DFFNX1_HVT \mem_reg[13][1]  ( .D(n779), .CLK(clk), .Q(\mem[13][1] ) );
  DFFNX1_HVT \mem_reg[13][0]  ( .D(n778), .CLK(clk), .Q(\mem[13][0] ) );
  DFFNX1_HVT \mem_reg[12][15]  ( .D(n777), .CLK(clk), .Q(\mem[12][15] ) );
  DFFNX1_HVT \mem_reg[12][14]  ( .D(n776), .CLK(clk), .Q(\mem[12][14] ) );
  DFFNX1_HVT \mem_reg[12][13]  ( .D(n775), .CLK(clk), .Q(\mem[12][13] ) );
  DFFNX1_HVT \mem_reg[12][12]  ( .D(n774), .CLK(clk), .Q(\mem[12][12] ) );
  DFFNX1_HVT \mem_reg[12][11]  ( .D(n773), .CLK(clk), .Q(\mem[12][11] ) );
  DFFNX1_HVT \mem_reg[12][10]  ( .D(n772), .CLK(clk), .Q(\mem[12][10] ) );
  DFFNX1_HVT \mem_reg[12][9]  ( .D(n771), .CLK(clk), .Q(\mem[12][9] ) );
  DFFNX1_HVT \mem_reg[12][8]  ( .D(n770), .CLK(clk), .Q(\mem[12][8] ) );
  DFFNX1_HVT \mem_reg[12][7]  ( .D(n769), .CLK(clk), .Q(\mem[12][7] ) );
  DFFNX1_HVT \mem_reg[12][6]  ( .D(n768), .CLK(clk), .Q(\mem[12][6] ) );
  DFFNX1_HVT \mem_reg[12][5]  ( .D(n767), .CLK(clk), .Q(\mem[12][5] ) );
  DFFNX1_HVT \mem_reg[12][4]  ( .D(n766), .CLK(clk), .Q(\mem[12][4] ) );
  DFFNX1_HVT \mem_reg[12][3]  ( .D(n765), .CLK(clk), .Q(\mem[12][3] ) );
  DFFNX1_HVT \mem_reg[12][2]  ( .D(n764), .CLK(clk), .Q(\mem[12][2] ) );
  DFFNX1_HVT \mem_reg[12][1]  ( .D(n763), .CLK(clk), .Q(\mem[12][1] ) );
  DFFNX1_HVT \mem_reg[12][0]  ( .D(n762), .CLK(clk), .Q(\mem[12][0] ) );
  DFFNX1_HVT \mem_reg[11][15]  ( .D(n761), .CLK(clk), .Q(\mem[11][15] ) );
  DFFNX1_HVT \mem_reg[11][14]  ( .D(n760), .CLK(clk), .Q(\mem[11][14] ) );
  DFFNX1_HVT \mem_reg[11][13]  ( .D(n759), .CLK(clk), .Q(\mem[11][13] ) );
  DFFNX1_HVT \mem_reg[11][12]  ( .D(n758), .CLK(clk), .Q(\mem[11][12] ) );
  DFFNX1_HVT \mem_reg[11][11]  ( .D(n757), .CLK(clk), .Q(\mem[11][11] ) );
  DFFNX1_HVT \mem_reg[11][10]  ( .D(n756), .CLK(clk), .Q(\mem[11][10] ) );
  DFFNX1_HVT \mem_reg[11][9]  ( .D(n755), .CLK(clk), .Q(\mem[11][9] ) );
  DFFNX1_HVT \mem_reg[11][8]  ( .D(n754), .CLK(clk), .Q(\mem[11][8] ) );
  DFFNX1_HVT \mem_reg[11][7]  ( .D(n753), .CLK(clk), .Q(\mem[11][7] ) );
  DFFNX1_HVT \mem_reg[11][6]  ( .D(n752), .CLK(clk), .Q(\mem[11][6] ) );
  DFFNX1_HVT \mem_reg[11][5]  ( .D(n751), .CLK(clk), .Q(\mem[11][5] ) );
  DFFNX1_HVT \mem_reg[11][4]  ( .D(n750), .CLK(clk), .Q(\mem[11][4] ) );
  DFFNX1_HVT \mem_reg[11][3]  ( .D(n749), .CLK(clk), .Q(\mem[11][3] ) );
  DFFNX1_HVT \mem_reg[11][2]  ( .D(n748), .CLK(clk), .Q(\mem[11][2] ) );
  DFFNX1_HVT \mem_reg[11][1]  ( .D(n747), .CLK(clk), .Q(\mem[11][1] ) );
  DFFNX1_HVT \mem_reg[11][0]  ( .D(n746), .CLK(clk), .Q(\mem[11][0] ) );
  DFFNX1_HVT \mem_reg[10][15]  ( .D(n745), .CLK(clk), .Q(\mem[10][15] ) );
  DFFNX1_HVT \mem_reg[10][14]  ( .D(n744), .CLK(clk), .Q(\mem[10][14] ) );
  DFFNX1_HVT \mem_reg[10][13]  ( .D(n743), .CLK(clk), .Q(\mem[10][13] ) );
  DFFNX1_HVT \mem_reg[10][12]  ( .D(n742), .CLK(clk), .Q(\mem[10][12] ) );
  DFFNX1_HVT \mem_reg[10][11]  ( .D(n741), .CLK(clk), .Q(\mem[10][11] ) );
  DFFNX1_HVT \mem_reg[10][10]  ( .D(n740), .CLK(clk), .Q(\mem[10][10] ) );
  DFFNX1_HVT \mem_reg[10][9]  ( .D(n739), .CLK(clk), .Q(\mem[10][9] ) );
  DFFNX1_HVT \mem_reg[10][8]  ( .D(n738), .CLK(clk), .Q(\mem[10][8] ) );
  DFFNX1_HVT \mem_reg[10][7]  ( .D(n737), .CLK(clk), .Q(\mem[10][7] ) );
  DFFNX1_HVT \mem_reg[10][6]  ( .D(n736), .CLK(clk), .Q(\mem[10][6] ) );
  DFFNX1_HVT \mem_reg[10][5]  ( .D(n735), .CLK(clk), .Q(\mem[10][5] ) );
  DFFNX1_HVT \mem_reg[10][4]  ( .D(n734), .CLK(clk), .Q(\mem[10][4] ) );
  DFFNX1_HVT \mem_reg[10][3]  ( .D(n733), .CLK(clk), .Q(\mem[10][3] ) );
  DFFNX1_HVT \mem_reg[10][2]  ( .D(n732), .CLK(clk), .Q(\mem[10][2] ) );
  DFFNX1_HVT \mem_reg[10][1]  ( .D(n731), .CLK(clk), .Q(\mem[10][1] ) );
  DFFNX1_HVT \mem_reg[10][0]  ( .D(n730), .CLK(clk), .Q(\mem[10][0] ) );
  DFFNX1_HVT \mem_reg[9][15]  ( .D(n729), .CLK(clk), .Q(\mem[9][15] ) );
  DFFNX1_HVT \mem_reg[9][14]  ( .D(n728), .CLK(clk), .Q(\mem[9][14] ) );
  DFFNX1_HVT \mem_reg[9][13]  ( .D(n727), .CLK(clk), .Q(\mem[9][13] ) );
  DFFNX1_HVT \mem_reg[9][12]  ( .D(n726), .CLK(clk), .Q(\mem[9][12] ) );
  DFFNX1_HVT \mem_reg[9][11]  ( .D(n725), .CLK(clk), .Q(\mem[9][11] ) );
  DFFNX1_HVT \mem_reg[9][10]  ( .D(n724), .CLK(clk), .Q(\mem[9][10] ) );
  DFFNX1_HVT \mem_reg[9][9]  ( .D(n723), .CLK(clk), .Q(\mem[9][9] ) );
  DFFNX1_HVT \mem_reg[9][8]  ( .D(n722), .CLK(clk), .Q(\mem[9][8] ) );
  DFFNX1_HVT \mem_reg[9][7]  ( .D(n721), .CLK(clk), .Q(\mem[9][7] ) );
  DFFNX1_HVT \mem_reg[9][6]  ( .D(n720), .CLK(clk), .Q(\mem[9][6] ) );
  DFFNX1_HVT \mem_reg[9][5]  ( .D(n719), .CLK(clk), .Q(\mem[9][5] ) );
  DFFNX1_HVT \mem_reg[9][4]  ( .D(n718), .CLK(clk), .Q(\mem[9][4] ) );
  DFFNX1_HVT \mem_reg[9][3]  ( .D(n717), .CLK(clk), .Q(\mem[9][3] ) );
  DFFNX1_HVT \mem_reg[9][2]  ( .D(n716), .CLK(clk), .Q(\mem[9][2] ) );
  DFFNX1_HVT \mem_reg[9][1]  ( .D(n715), .CLK(clk), .Q(\mem[9][1] ) );
  DFFNX1_HVT \mem_reg[9][0]  ( .D(n714), .CLK(clk), .Q(\mem[9][0] ) );
  DFFNX1_HVT \mem_reg[8][15]  ( .D(n713), .CLK(clk), .Q(\mem[8][15] ) );
  DFFNX1_HVT \mem_reg[8][14]  ( .D(n712), .CLK(clk), .Q(\mem[8][14] ) );
  DFFNX1_HVT \mem_reg[8][13]  ( .D(n711), .CLK(clk), .Q(\mem[8][13] ) );
  DFFNX1_HVT \mem_reg[8][12]  ( .D(n710), .CLK(clk), .Q(\mem[8][12] ) );
  DFFNX1_HVT \mem_reg[8][11]  ( .D(n709), .CLK(clk), .Q(\mem[8][11] ) );
  DFFNX1_HVT \mem_reg[8][10]  ( .D(n708), .CLK(clk), .Q(\mem[8][10] ) );
  DFFNX1_HVT \mem_reg[8][9]  ( .D(n707), .CLK(clk), .Q(\mem[8][9] ) );
  DFFNX1_HVT \mem_reg[8][8]  ( .D(n706), .CLK(clk), .Q(\mem[8][8] ) );
  DFFNX1_HVT \mem_reg[8][7]  ( .D(n705), .CLK(clk), .Q(\mem[8][7] ) );
  DFFNX1_HVT \mem_reg[8][6]  ( .D(n704), .CLK(clk), .Q(\mem[8][6] ) );
  DFFNX1_HVT \mem_reg[8][5]  ( .D(n703), .CLK(clk), .Q(\mem[8][5] ) );
  DFFNX1_HVT \mem_reg[8][4]  ( .D(n702), .CLK(clk), .Q(\mem[8][4] ) );
  DFFNX1_HVT \mem_reg[8][3]  ( .D(n701), .CLK(clk), .Q(\mem[8][3] ) );
  DFFNX1_HVT \mem_reg[8][2]  ( .D(n700), .CLK(clk), .Q(\mem[8][2] ) );
  DFFNX1_HVT \mem_reg[8][1]  ( .D(n699), .CLK(clk), .Q(\mem[8][1] ) );
  DFFNX1_HVT \mem_reg[8][0]  ( .D(n698), .CLK(clk), .Q(\mem[8][0] ) );
  DFFNX1_HVT \mem_reg[7][15]  ( .D(n697), .CLK(clk), .Q(\mem[7][15] ) );
  DFFNX1_HVT \mem_reg[7][14]  ( .D(n696), .CLK(clk), .Q(\mem[7][14] ) );
  DFFNX1_HVT \mem_reg[7][13]  ( .D(n695), .CLK(clk), .Q(\mem[7][13] ) );
  DFFNX1_HVT \mem_reg[7][12]  ( .D(n694), .CLK(clk), .Q(\mem[7][12] ) );
  DFFNX1_HVT \mem_reg[7][11]  ( .D(n693), .CLK(clk), .Q(\mem[7][11] ) );
  DFFNX1_HVT \mem_reg[7][10]  ( .D(n692), .CLK(clk), .Q(\mem[7][10] ) );
  DFFNX1_HVT \mem_reg[7][9]  ( .D(n691), .CLK(clk), .Q(\mem[7][9] ) );
  DFFNX1_HVT \mem_reg[7][8]  ( .D(n690), .CLK(clk), .Q(\mem[7][8] ) );
  DFFNX1_HVT \mem_reg[7][7]  ( .D(n689), .CLK(clk), .Q(\mem[7][7] ) );
  DFFNX1_HVT \mem_reg[7][6]  ( .D(n688), .CLK(clk), .Q(\mem[7][6] ) );
  DFFNX1_HVT \mem_reg[7][5]  ( .D(n687), .CLK(clk), .Q(\mem[7][5] ) );
  DFFNX1_HVT \mem_reg[7][4]  ( .D(n686), .CLK(clk), .Q(\mem[7][4] ) );
  DFFNX1_HVT \mem_reg[7][3]  ( .D(n685), .CLK(clk), .Q(\mem[7][3] ) );
  DFFNX1_HVT \mem_reg[7][2]  ( .D(n684), .CLK(clk), .Q(\mem[7][2] ) );
  DFFNX1_HVT \mem_reg[7][1]  ( .D(n683), .CLK(clk), .Q(\mem[7][1] ) );
  DFFNX1_HVT \mem_reg[7][0]  ( .D(n682), .CLK(clk), .Q(\mem[7][0] ) );
  DFFNX1_HVT \mem_reg[6][15]  ( .D(n681), .CLK(clk), .Q(\mem[6][15] ) );
  DFFNX1_HVT \mem_reg[6][14]  ( .D(n680), .CLK(clk), .Q(\mem[6][14] ) );
  DFFNX1_HVT \mem_reg[6][13]  ( .D(n679), .CLK(clk), .Q(\mem[6][13] ) );
  DFFNX1_HVT \mem_reg[6][12]  ( .D(n678), .CLK(clk), .Q(\mem[6][12] ) );
  DFFNX1_HVT \mem_reg[6][11]  ( .D(n677), .CLK(clk), .Q(\mem[6][11] ) );
  DFFNX1_HVT \mem_reg[6][10]  ( .D(n676), .CLK(clk), .Q(\mem[6][10] ) );
  DFFNX1_HVT \mem_reg[6][9]  ( .D(n675), .CLK(clk), .Q(\mem[6][9] ) );
  DFFNX1_HVT \mem_reg[6][8]  ( .D(n674), .CLK(clk), .Q(\mem[6][8] ) );
  DFFNX1_HVT \mem_reg[6][7]  ( .D(n673), .CLK(clk), .Q(\mem[6][7] ) );
  DFFNX1_HVT \mem_reg[6][6]  ( .D(n672), .CLK(clk), .Q(\mem[6][6] ) );
  DFFNX1_HVT \mem_reg[6][5]  ( .D(n671), .CLK(clk), .Q(\mem[6][5] ) );
  DFFNX1_HVT \mem_reg[6][4]  ( .D(n670), .CLK(clk), .Q(\mem[6][4] ) );
  DFFNX1_HVT \mem_reg[6][3]  ( .D(n669), .CLK(clk), .Q(\mem[6][3] ) );
  DFFNX1_HVT \mem_reg[6][2]  ( .D(n668), .CLK(clk), .Q(\mem[6][2] ) );
  DFFNX1_HVT \mem_reg[6][1]  ( .D(n667), .CLK(clk), .Q(\mem[6][1] ) );
  DFFNX1_HVT \mem_reg[6][0]  ( .D(n666), .CLK(clk), .Q(\mem[6][0] ) );
  DFFNX1_HVT \mem_reg[5][15]  ( .D(n665), .CLK(clk), .Q(\mem[5][15] ) );
  DFFNX1_HVT \mem_reg[5][14]  ( .D(n664), .CLK(clk), .Q(\mem[5][14] ) );
  DFFNX1_HVT \mem_reg[5][13]  ( .D(n663), .CLK(clk), .Q(\mem[5][13] ) );
  DFFNX1_HVT \mem_reg[5][12]  ( .D(n662), .CLK(clk), .Q(\mem[5][12] ) );
  DFFNX1_HVT \mem_reg[5][11]  ( .D(n661), .CLK(clk), .Q(\mem[5][11] ) );
  DFFNX1_HVT \mem_reg[5][10]  ( .D(n660), .CLK(clk), .Q(\mem[5][10] ) );
  DFFNX1_HVT \mem_reg[5][9]  ( .D(n659), .CLK(clk), .Q(\mem[5][9] ) );
  DFFNX1_HVT \mem_reg[5][8]  ( .D(n658), .CLK(clk), .Q(\mem[5][8] ) );
  DFFNX1_HVT \mem_reg[5][7]  ( .D(n657), .CLK(clk), .Q(\mem[5][7] ) );
  DFFNX1_HVT \mem_reg[5][6]  ( .D(n656), .CLK(clk), .Q(\mem[5][6] ) );
  DFFNX1_HVT \mem_reg[5][5]  ( .D(n655), .CLK(clk), .Q(\mem[5][5] ) );
  DFFNX1_HVT \mem_reg[5][4]  ( .D(n654), .CLK(clk), .Q(\mem[5][4] ) );
  DFFNX1_HVT \mem_reg[5][3]  ( .D(n653), .CLK(clk), .Q(\mem[5][3] ) );
  DFFNX1_HVT \mem_reg[5][2]  ( .D(n652), .CLK(clk), .Q(\mem[5][2] ) );
  DFFNX1_HVT \mem_reg[5][1]  ( .D(n651), .CLK(clk), .Q(\mem[5][1] ) );
  DFFNX1_HVT \mem_reg[5][0]  ( .D(n650), .CLK(clk), .Q(\mem[5][0] ) );
  DFFNX1_HVT \mem_reg[4][15]  ( .D(n649), .CLK(clk), .Q(\mem[4][15] ) );
  DFFNX1_HVT \mem_reg[4][14]  ( .D(n648), .CLK(clk), .Q(\mem[4][14] ) );
  DFFNX1_HVT \mem_reg[4][13]  ( .D(n647), .CLK(clk), .Q(\mem[4][13] ) );
  DFFNX1_HVT \mem_reg[4][12]  ( .D(n646), .CLK(clk), .Q(\mem[4][12] ) );
  DFFNX1_HVT \mem_reg[4][11]  ( .D(n645), .CLK(clk), .Q(\mem[4][11] ) );
  DFFNX1_HVT \mem_reg[4][10]  ( .D(n644), .CLK(clk), .Q(\mem[4][10] ) );
  DFFNX1_HVT \mem_reg[4][9]  ( .D(n643), .CLK(clk), .Q(\mem[4][9] ) );
  DFFNX1_HVT \mem_reg[4][8]  ( .D(n642), .CLK(clk), .Q(\mem[4][8] ) );
  DFFNX1_HVT \mem_reg[4][7]  ( .D(n641), .CLK(clk), .Q(\mem[4][7] ) );
  DFFNX1_HVT \mem_reg[4][6]  ( .D(n640), .CLK(clk), .Q(\mem[4][6] ) );
  DFFNX1_HVT \mem_reg[4][5]  ( .D(n639), .CLK(clk), .Q(\mem[4][5] ) );
  DFFNX1_HVT \mem_reg[4][4]  ( .D(n638), .CLK(clk), .Q(\mem[4][4] ) );
  DFFNX1_HVT \mem_reg[4][3]  ( .D(n637), .CLK(clk), .Q(\mem[4][3] ) );
  DFFNX1_HVT \mem_reg[4][2]  ( .D(n636), .CLK(clk), .Q(\mem[4][2] ) );
  DFFNX1_HVT \mem_reg[4][1]  ( .D(n635), .CLK(clk), .Q(\mem[4][1] ) );
  DFFNX1_HVT \mem_reg[4][0]  ( .D(n634), .CLK(clk), .Q(\mem[4][0] ) );
  DFFNX1_HVT \mem_reg[3][15]  ( .D(n633), .CLK(clk), .Q(\mem[3][15] ) );
  DFFNX1_HVT \mem_reg[3][14]  ( .D(n632), .CLK(clk), .Q(\mem[3][14] ) );
  DFFNX1_HVT \mem_reg[3][13]  ( .D(n631), .CLK(clk), .Q(\mem[3][13] ) );
  DFFNX1_HVT \mem_reg[3][12]  ( .D(n630), .CLK(clk), .Q(\mem[3][12] ) );
  DFFNX1_HVT \mem_reg[3][11]  ( .D(n629), .CLK(clk), .Q(\mem[3][11] ) );
  DFFNX1_HVT \mem_reg[3][10]  ( .D(n628), .CLK(clk), .Q(\mem[3][10] ) );
  DFFNX1_HVT \mem_reg[3][9]  ( .D(n627), .CLK(clk), .Q(\mem[3][9] ) );
  DFFNX1_HVT \mem_reg[3][8]  ( .D(n626), .CLK(clk), .Q(\mem[3][8] ) );
  DFFNX1_HVT \mem_reg[3][7]  ( .D(n625), .CLK(clk), .Q(\mem[3][7] ) );
  DFFNX1_HVT \mem_reg[3][6]  ( .D(n624), .CLK(clk), .Q(\mem[3][6] ) );
  DFFNX1_HVT \mem_reg[3][5]  ( .D(n623), .CLK(clk), .Q(\mem[3][5] ) );
  DFFNX1_HVT \mem_reg[3][4]  ( .D(n622), .CLK(clk), .Q(\mem[3][4] ) );
  DFFNX1_HVT \mem_reg[3][3]  ( .D(n621), .CLK(clk), .Q(\mem[3][3] ) );
  DFFNX1_HVT \mem_reg[3][2]  ( .D(n620), .CLK(clk), .Q(\mem[3][2] ) );
  DFFNX1_HVT \mem_reg[3][1]  ( .D(n619), .CLK(clk), .Q(\mem[3][1] ) );
  DFFNX1_HVT \mem_reg[3][0]  ( .D(n618), .CLK(clk), .Q(\mem[3][0] ) );
  DFFNX1_HVT \mem_reg[2][15]  ( .D(n617), .CLK(clk), .Q(\mem[2][15] ) );
  DFFNX1_HVT \mem_reg[2][14]  ( .D(n616), .CLK(clk), .Q(\mem[2][14] ) );
  DFFNX1_HVT \mem_reg[2][13]  ( .D(n615), .CLK(clk), .Q(\mem[2][13] ) );
  DFFNX1_HVT \mem_reg[2][12]  ( .D(n614), .CLK(clk), .Q(\mem[2][12] ) );
  DFFNX1_HVT \mem_reg[2][11]  ( .D(n613), .CLK(clk), .Q(\mem[2][11] ) );
  DFFNX1_HVT \mem_reg[2][10]  ( .D(n612), .CLK(clk), .Q(\mem[2][10] ) );
  DFFNX1_HVT \mem_reg[2][9]  ( .D(n611), .CLK(clk), .Q(\mem[2][9] ) );
  DFFNX1_HVT \mem_reg[2][8]  ( .D(n610), .CLK(clk), .Q(\mem[2][8] ) );
  DFFNX1_HVT \mem_reg[2][7]  ( .D(n609), .CLK(clk), .Q(\mem[2][7] ) );
  DFFNX1_HVT \mem_reg[2][6]  ( .D(n608), .CLK(clk), .Q(\mem[2][6] ) );
  DFFNX1_HVT \mem_reg[2][5]  ( .D(n607), .CLK(clk), .Q(\mem[2][5] ) );
  DFFNX1_HVT \mem_reg[2][4]  ( .D(n606), .CLK(clk), .Q(\mem[2][4] ) );
  DFFNX1_HVT \mem_reg[2][3]  ( .D(n605), .CLK(clk), .Q(\mem[2][3] ) );
  DFFNX1_HVT \mem_reg[2][2]  ( .D(n604), .CLK(clk), .Q(\mem[2][2] ) );
  DFFNX1_HVT \mem_reg[2][1]  ( .D(n603), .CLK(clk), .Q(\mem[2][1] ) );
  DFFNX1_HVT \mem_reg[2][0]  ( .D(n602), .CLK(clk), .Q(\mem[2][0] ) );
  DFFNX1_HVT \mem_reg[1][15]  ( .D(n601), .CLK(clk), .Q(\mem[1][15] ) );
  DFFNX1_HVT \mem_reg[1][14]  ( .D(n600), .CLK(clk), .Q(\mem[1][14] ) );
  DFFNX1_HVT \mem_reg[1][13]  ( .D(n599), .CLK(clk), .Q(\mem[1][13] ) );
  DFFNX1_HVT \mem_reg[1][12]  ( .D(n598), .CLK(clk), .Q(\mem[1][12] ) );
  DFFNX1_HVT \mem_reg[1][11]  ( .D(n597), .CLK(clk), .Q(\mem[1][11] ) );
  DFFNX1_HVT \mem_reg[1][10]  ( .D(n596), .CLK(clk), .Q(\mem[1][10] ) );
  DFFNX1_HVT \mem_reg[1][9]  ( .D(n595), .CLK(clk), .Q(\mem[1][9] ) );
  DFFNX1_HVT \mem_reg[1][8]  ( .D(n594), .CLK(clk), .Q(\mem[1][8] ) );
  DFFNX1_HVT \mem_reg[1][7]  ( .D(n593), .CLK(clk), .Q(\mem[1][7] ) );
  DFFNX1_HVT \mem_reg[1][6]  ( .D(n592), .CLK(clk), .Q(\mem[1][6] ) );
  DFFNX1_HVT \mem_reg[1][5]  ( .D(n591), .CLK(clk), .Q(\mem[1][5] ) );
  DFFNX1_HVT \mem_reg[1][4]  ( .D(n590), .CLK(clk), .Q(\mem[1][4] ) );
  DFFNX1_HVT \mem_reg[1][3]  ( .D(n589), .CLK(clk), .Q(\mem[1][3] ) );
  DFFNX1_HVT \mem_reg[1][2]  ( .D(n588), .CLK(clk), .Q(\mem[1][2] ) );
  DFFNX1_HVT \mem_reg[1][1]  ( .D(n587), .CLK(clk), .Q(\mem[1][1] ) );
  DFFNX1_HVT \mem_reg[1][0]  ( .D(n586), .CLK(clk), .Q(\mem[1][0] ) );
  DFFNX1_HVT \mem_reg[0][15]  ( .D(n585), .CLK(clk), .Q(\mem[0][15] ) );
  DFFNX1_HVT \mem_reg[0][14]  ( .D(n584), .CLK(clk), .Q(\mem[0][14] ) );
  DFFNX1_HVT \mem_reg[0][13]  ( .D(n583), .CLK(clk), .Q(\mem[0][13] ) );
  DFFNX1_HVT \mem_reg[0][12]  ( .D(n582), .CLK(clk), .Q(\mem[0][12] ) );
  DFFNX1_HVT \mem_reg[0][11]  ( .D(n581), .CLK(clk), .Q(\mem[0][11] ) );
  DFFNX1_HVT \mem_reg[0][10]  ( .D(n580), .CLK(clk), .Q(\mem[0][10] ) );
  DFFNX1_HVT \mem_reg[0][9]  ( .D(n579), .CLK(clk), .Q(\mem[0][9] ) );
  DFFNX1_HVT \mem_reg[0][8]  ( .D(n578), .CLK(clk), .Q(\mem[0][8] ) );
  DFFNX1_HVT \mem_reg[0][7]  ( .D(n577), .CLK(clk), .Q(\mem[0][7] ) );
  DFFNX1_HVT \mem_reg[0][6]  ( .D(n576), .CLK(clk), .Q(\mem[0][6] ) );
  DFFNX1_HVT \mem_reg[0][5]  ( .D(n575), .CLK(clk), .Q(\mem[0][5] ) );
  DFFNX1_HVT \mem_reg[0][4]  ( .D(n574), .CLK(clk), .Q(\mem[0][4] ) );
  DFFNX1_HVT \mem_reg[0][3]  ( .D(n573), .CLK(clk), .Q(\mem[0][3] ) );
  DFFNX1_HVT \mem_reg[0][2]  ( .D(n572), .CLK(clk), .Q(\mem[0][2] ) );
  DFFNX1_HVT \mem_reg[0][1]  ( .D(n571), .CLK(clk), .Q(\mem[0][1] ) );
  DFFNX1_HVT \mem_reg[0][0]  ( .D(n570), .CLK(clk), .Q(\mem[0][0] ) );
  MUX41X1_HVT U3 ( .A1(\mem[12][0] ), .A3(\mem[14][0] ), .A2(\mem[13][0] ), 
        .A4(\mem[15][0] ), .S0(N18), .S1(N17), .Y(n1) );
  MUX41X1_HVT U4 ( .A1(\mem[8][0] ), .A3(\mem[10][0] ), .A2(\mem[9][0] ), .A4(
        \mem[11][0] ), .S0(N18), .S1(N17), .Y(n2) );
  MUX41X1_HVT U5 ( .A1(\mem[4][0] ), .A3(\mem[6][0] ), .A2(\mem[5][0] ), .A4(
        \mem[7][0] ), .S0(N18), .S1(N17), .Y(n3) );
  MUX41X1_HVT U6 ( .A1(\mem[0][0] ), .A3(\mem[2][0] ), .A2(\mem[1][0] ), .A4(
        \mem[3][0] ), .S0(N18), .S1(N17), .Y(n4) );
  MUX41X1_HVT U7 ( .A1(n4), .A3(n2), .A2(n3), .A4(n1), .S0(N20), .S1(N19), .Y(
        N554) );
  MUX41X1_HVT U8 ( .A1(\mem[12][1] ), .A3(\mem[14][1] ), .A2(\mem[13][1] ), 
        .A4(\mem[15][1] ), .S0(N18), .S1(N17), .Y(n5) );
  MUX41X1_HVT U9 ( .A1(\mem[8][1] ), .A3(\mem[10][1] ), .A2(\mem[9][1] ), .A4(
        \mem[11][1] ), .S0(N18), .S1(N17), .Y(n6) );
  MUX41X1_HVT U10 ( .A1(\mem[4][1] ), .A3(\mem[6][1] ), .A2(\mem[5][1] ), .A4(
        \mem[7][1] ), .S0(N18), .S1(N17), .Y(n7) );
  MUX41X1_HVT U11 ( .A1(\mem[0][1] ), .A3(\mem[2][1] ), .A2(\mem[1][1] ), .A4(
        \mem[3][1] ), .S0(N18), .S1(N17), .Y(n8) );
  MUX41X1_HVT U12 ( .A1(n8), .A3(n6), .A2(n7), .A4(n5), .S0(N20), .S1(N19), 
        .Y(N553) );
  MUX41X1_HVT U13 ( .A1(\mem[12][2] ), .A3(\mem[14][2] ), .A2(\mem[13][2] ), 
        .A4(\mem[15][2] ), .S0(N18), .S1(N17), .Y(n9) );
  MUX41X1_HVT U14 ( .A1(\mem[8][2] ), .A3(\mem[10][2] ), .A2(\mem[9][2] ), 
        .A4(\mem[11][2] ), .S0(N18), .S1(N17), .Y(n10) );
  MUX41X1_HVT U15 ( .A1(\mem[4][2] ), .A3(\mem[6][2] ), .A2(\mem[5][2] ), .A4(
        \mem[7][2] ), .S0(N18), .S1(N17), .Y(n11) );
  MUX41X1_HVT U16 ( .A1(\mem[0][2] ), .A3(\mem[2][2] ), .A2(\mem[1][2] ), .A4(
        \mem[3][2] ), .S0(N18), .S1(N17), .Y(n12) );
  MUX41X1_HVT U17 ( .A1(n12), .A3(n10), .A2(n11), .A4(n9), .S0(N20), .S1(N19), 
        .Y(N552) );
  MUX41X1_HVT U18 ( .A1(\mem[12][3] ), .A3(\mem[14][3] ), .A2(\mem[13][3] ), 
        .A4(\mem[15][3] ), .S0(N18), .S1(N17), .Y(n13) );
  MUX41X1_HVT U19 ( .A1(\mem[8][3] ), .A3(\mem[10][3] ), .A2(\mem[9][3] ), 
        .A4(\mem[11][3] ), .S0(N18), .S1(N17), .Y(n14) );
  MUX41X1_HVT U20 ( .A1(\mem[4][3] ), .A3(\mem[6][3] ), .A2(\mem[5][3] ), .A4(
        \mem[7][3] ), .S0(N18), .S1(N17), .Y(n15) );
  MUX41X1_HVT U21 ( .A1(\mem[0][3] ), .A3(\mem[2][3] ), .A2(\mem[1][3] ), .A4(
        \mem[3][3] ), .S0(N18), .S1(N17), .Y(n16) );
  MUX41X1_HVT U22 ( .A1(n16), .A3(n14), .A2(n15), .A4(n13), .S0(N20), .S1(N19), 
        .Y(N551) );
  MUX41X1_HVT U23 ( .A1(\mem[12][4] ), .A3(\mem[14][4] ), .A2(\mem[13][4] ), 
        .A4(\mem[15][4] ), .S0(N18), .S1(N17), .Y(n17) );
  MUX41X1_HVT U24 ( .A1(\mem[8][4] ), .A3(\mem[10][4] ), .A2(\mem[9][4] ), 
        .A4(\mem[11][4] ), .S0(N18), .S1(N17), .Y(n18) );
  MUX41X1_HVT U25 ( .A1(\mem[4][4] ), .A3(\mem[6][4] ), .A2(\mem[5][4] ), .A4(
        \mem[7][4] ), .S0(N18), .S1(N17), .Y(n19) );
  MUX41X1_HVT U26 ( .A1(\mem[0][4] ), .A3(\mem[2][4] ), .A2(\mem[1][4] ), .A4(
        \mem[3][4] ), .S0(N18), .S1(N17), .Y(n20) );
  MUX41X1_HVT U27 ( .A1(n20), .A3(n18), .A2(n19), .A4(n17), .S0(N20), .S1(N19), 
        .Y(N550) );
  MUX41X1_HVT U28 ( .A1(\mem[12][5] ), .A3(\mem[14][5] ), .A2(\mem[13][5] ), 
        .A4(\mem[15][5] ), .S0(N18), .S1(N17), .Y(n21) );
  MUX41X1_HVT U29 ( .A1(\mem[8][5] ), .A3(\mem[10][5] ), .A2(\mem[9][5] ), 
        .A4(\mem[11][5] ), .S0(N18), .S1(N17), .Y(n22) );
  MUX41X1_HVT U30 ( .A1(\mem[4][5] ), .A3(\mem[6][5] ), .A2(\mem[5][5] ), .A4(
        \mem[7][5] ), .S0(N18), .S1(N17), .Y(n23) );
  MUX41X1_HVT U31 ( .A1(\mem[0][5] ), .A3(\mem[2][5] ), .A2(\mem[1][5] ), .A4(
        \mem[3][5] ), .S0(N18), .S1(N17), .Y(n24) );
  MUX41X1_HVT U32 ( .A1(n24), .A3(n22), .A2(n23), .A4(n21), .S0(N20), .S1(N19), 
        .Y(N549) );
  MUX41X1_HVT U33 ( .A1(\mem[12][6] ), .A3(\mem[14][6] ), .A2(\mem[13][6] ), 
        .A4(\mem[15][6] ), .S0(N18), .S1(N17), .Y(n25) );
  MUX41X1_HVT U34 ( .A1(\mem[8][6] ), .A3(\mem[10][6] ), .A2(\mem[9][6] ), 
        .A4(\mem[11][6] ), .S0(N18), .S1(N17), .Y(n26) );
  MUX41X1_HVT U35 ( .A1(\mem[4][6] ), .A3(\mem[6][6] ), .A2(\mem[5][6] ), .A4(
        \mem[7][6] ), .S0(N18), .S1(N17), .Y(n27) );
  MUX41X1_HVT U36 ( .A1(\mem[0][6] ), .A3(\mem[2][6] ), .A2(\mem[1][6] ), .A4(
        \mem[3][6] ), .S0(N18), .S1(N17), .Y(n28) );
  MUX41X1_HVT U37 ( .A1(n28), .A3(n26), .A2(n27), .A4(n25), .S0(N20), .S1(N19), 
        .Y(N548) );
  MUX41X1_HVT U38 ( .A1(\mem[12][7] ), .A3(\mem[14][7] ), .A2(\mem[13][7] ), 
        .A4(\mem[15][7] ), .S0(N18), .S1(N17), .Y(n29) );
  MUX41X1_HVT U39 ( .A1(\mem[8][7] ), .A3(\mem[10][7] ), .A2(\mem[9][7] ), 
        .A4(\mem[11][7] ), .S0(N18), .S1(N17), .Y(n30) );
  MUX41X1_HVT U40 ( .A1(\mem[4][7] ), .A3(\mem[6][7] ), .A2(\mem[5][7] ), .A4(
        \mem[7][7] ), .S0(N18), .S1(N17), .Y(n31) );
  MUX41X1_HVT U41 ( .A1(\mem[0][7] ), .A3(\mem[2][7] ), .A2(\mem[1][7] ), .A4(
        \mem[3][7] ), .S0(N18), .S1(N17), .Y(n32) );
  MUX41X1_HVT U42 ( .A1(n32), .A3(n30), .A2(n31), .A4(n29), .S0(N20), .S1(N19), 
        .Y(N547) );
  MUX41X1_HVT U43 ( .A1(\mem[12][8] ), .A3(\mem[14][8] ), .A2(\mem[13][8] ), 
        .A4(\mem[15][8] ), .S0(N18), .S1(N17), .Y(n33) );
  MUX41X1_HVT U44 ( .A1(\mem[8][8] ), .A3(\mem[10][8] ), .A2(\mem[9][8] ), 
        .A4(\mem[11][8] ), .S0(N18), .S1(N17), .Y(n34) );
  MUX41X1_HVT U45 ( .A1(\mem[4][8] ), .A3(\mem[6][8] ), .A2(\mem[5][8] ), .A4(
        \mem[7][8] ), .S0(N18), .S1(N17), .Y(n35) );
  MUX41X1_HVT U46 ( .A1(\mem[0][8] ), .A3(\mem[2][8] ), .A2(\mem[1][8] ), .A4(
        \mem[3][8] ), .S0(N18), .S1(N17), .Y(n36) );
  MUX41X1_HVT U47 ( .A1(n36), .A3(n34), .A2(n35), .A4(n33), .S0(N20), .S1(N19), 
        .Y(N546) );
  MUX41X1_HVT U48 ( .A1(\mem[12][9] ), .A3(\mem[14][9] ), .A2(\mem[13][9] ), 
        .A4(\mem[15][9] ), .S0(N18), .S1(N17), .Y(n37) );
  MUX41X1_HVT U49 ( .A1(\mem[8][9] ), .A3(\mem[10][9] ), .A2(\mem[9][9] ), 
        .A4(\mem[11][9] ), .S0(N18), .S1(N17), .Y(n38) );
  MUX41X1_HVT U50 ( .A1(\mem[4][9] ), .A3(\mem[6][9] ), .A2(\mem[5][9] ), .A4(
        \mem[7][9] ), .S0(N18), .S1(N17), .Y(n39) );
  MUX41X1_HVT U51 ( .A1(\mem[0][9] ), .A3(\mem[2][9] ), .A2(\mem[1][9] ), .A4(
        \mem[3][9] ), .S0(N18), .S1(N17), .Y(n40) );
  MUX41X1_HVT U52 ( .A1(n40), .A3(n38), .A2(n39), .A4(n37), .S0(N20), .S1(N19), 
        .Y(N545) );
  MUX41X1_HVT U53 ( .A1(\mem[12][10] ), .A3(\mem[14][10] ), .A2(\mem[13][10] ), 
        .A4(\mem[15][10] ), .S0(N18), .S1(N17), .Y(n41) );
  MUX41X1_HVT U54 ( .A1(\mem[8][10] ), .A3(\mem[10][10] ), .A2(\mem[9][10] ), 
        .A4(\mem[11][10] ), .S0(N18), .S1(N17), .Y(n42) );
  MUX41X1_HVT U55 ( .A1(\mem[4][10] ), .A3(\mem[6][10] ), .A2(\mem[5][10] ), 
        .A4(\mem[7][10] ), .S0(N18), .S1(N17), .Y(n43) );
  MUX41X1_HVT U56 ( .A1(\mem[0][10] ), .A3(\mem[2][10] ), .A2(\mem[1][10] ), 
        .A4(\mem[3][10] ), .S0(N18), .S1(N17), .Y(n44) );
  MUX41X1_HVT U57 ( .A1(n44), .A3(n42), .A2(n43), .A4(n41), .S0(N20), .S1(N19), 
        .Y(N544) );
  MUX41X1_HVT U58 ( .A1(\mem[12][11] ), .A3(\mem[14][11] ), .A2(\mem[13][11] ), 
        .A4(\mem[15][11] ), .S0(N18), .S1(N17), .Y(n45) );
  MUX41X1_HVT U59 ( .A1(\mem[8][11] ), .A3(\mem[10][11] ), .A2(\mem[9][11] ), 
        .A4(\mem[11][11] ), .S0(N18), .S1(N17), .Y(n46) );
  MUX41X1_HVT U60 ( .A1(\mem[4][11] ), .A3(\mem[6][11] ), .A2(\mem[5][11] ), 
        .A4(\mem[7][11] ), .S0(N18), .S1(N17), .Y(n47) );
  MUX41X1_HVT U61 ( .A1(\mem[0][11] ), .A3(\mem[2][11] ), .A2(\mem[1][11] ), 
        .A4(\mem[3][11] ), .S0(N18), .S1(N17), .Y(n48) );
  MUX41X1_HVT U62 ( .A1(n48), .A3(n46), .A2(n47), .A4(n45), .S0(N20), .S1(N19), 
        .Y(N543) );
  MUX41X1_HVT U63 ( .A1(\mem[12][12] ), .A3(\mem[14][12] ), .A2(\mem[13][12] ), 
        .A4(\mem[15][12] ), .S0(N18), .S1(N17), .Y(n49) );
  MUX41X1_HVT U64 ( .A1(\mem[8][12] ), .A3(\mem[10][12] ), .A2(\mem[9][12] ), 
        .A4(\mem[11][12] ), .S0(N18), .S1(N17), .Y(n50) );
  MUX41X1_HVT U65 ( .A1(\mem[4][12] ), .A3(\mem[6][12] ), .A2(\mem[5][12] ), 
        .A4(\mem[7][12] ), .S0(N18), .S1(N17), .Y(n51) );
  MUX41X1_HVT U66 ( .A1(\mem[0][12] ), .A3(\mem[2][12] ), .A2(\mem[1][12] ), 
        .A4(\mem[3][12] ), .S0(N18), .S1(N17), .Y(n52) );
  MUX41X1_HVT U67 ( .A1(n52), .A3(n50), .A2(n51), .A4(n49), .S0(N20), .S1(N19), 
        .Y(N542) );
  MUX41X1_HVT U68 ( .A1(\mem[12][13] ), .A3(\mem[14][13] ), .A2(\mem[13][13] ), 
        .A4(\mem[15][13] ), .S0(N18), .S1(N17), .Y(n53) );
  MUX41X1_HVT U69 ( .A1(\mem[8][13] ), .A3(\mem[10][13] ), .A2(\mem[9][13] ), 
        .A4(\mem[11][13] ), .S0(N18), .S1(N17), .Y(n54) );
  MUX41X1_HVT U70 ( .A1(\mem[4][13] ), .A3(\mem[6][13] ), .A2(\mem[5][13] ), 
        .A4(\mem[7][13] ), .S0(N18), .S1(N17), .Y(n55) );
  MUX41X1_HVT U71 ( .A1(\mem[0][13] ), .A3(\mem[2][13] ), .A2(\mem[1][13] ), 
        .A4(\mem[3][13] ), .S0(N18), .S1(N17), .Y(n56) );
  MUX41X1_HVT U72 ( .A1(n56), .A3(n54), .A2(n55), .A4(n53), .S0(N20), .S1(N19), 
        .Y(N541) );
  MUX41X1_HVT U73 ( .A1(\mem[12][14] ), .A3(\mem[14][14] ), .A2(\mem[13][14] ), 
        .A4(\mem[15][14] ), .S0(N18), .S1(N17), .Y(n57) );
  MUX41X1_HVT U74 ( .A1(\mem[8][14] ), .A3(\mem[10][14] ), .A2(\mem[9][14] ), 
        .A4(\mem[11][14] ), .S0(N18), .S1(N17), .Y(n58) );
  MUX41X1_HVT U75 ( .A1(\mem[4][14] ), .A3(\mem[6][14] ), .A2(\mem[5][14] ), 
        .A4(\mem[7][14] ), .S0(N18), .S1(N17), .Y(n59) );
  MUX41X1_HVT U76 ( .A1(\mem[0][14] ), .A3(\mem[2][14] ), .A2(\mem[1][14] ), 
        .A4(\mem[3][14] ), .S0(N18), .S1(N17), .Y(n60) );
  MUX41X1_HVT U77 ( .A1(n60), .A3(n58), .A2(n59), .A4(n57), .S0(N20), .S1(N19), 
        .Y(N540) );
  MUX41X1_HVT U78 ( .A1(\mem[12][15] ), .A3(\mem[14][15] ), .A2(\mem[13][15] ), 
        .A4(\mem[15][15] ), .S0(N18), .S1(N17), .Y(n61) );
  MUX41X1_HVT U79 ( .A1(\mem[8][15] ), .A3(\mem[10][15] ), .A2(\mem[9][15] ), 
        .A4(\mem[11][15] ), .S0(N18), .S1(N17), .Y(n62) );
  MUX41X1_HVT U80 ( .A1(\mem[4][15] ), .A3(\mem[6][15] ), .A2(\mem[5][15] ), 
        .A4(\mem[7][15] ), .S0(N18), .S1(N17), .Y(n63) );
  MUX41X1_HVT U81 ( .A1(\mem[0][15] ), .A3(\mem[2][15] ), .A2(\mem[1][15] ), 
        .A4(\mem[3][15] ), .S0(N18), .S1(N17), .Y(n64) );
  MUX41X1_HVT U82 ( .A1(n64), .A3(n62), .A2(n63), .A4(n61), .S0(N20), .S1(N19), 
        .Y(N539) );
  AO22X1_HVT U83 ( .A1(\mem[15][15] ), .A2(n65), .A3(n66), .A4(n67), .Y(n825)
         );
  AO22X1_HVT U84 ( .A1(\mem[15][14] ), .A2(n65), .A3(n68), .A4(n66), .Y(n824)
         );
  AO22X1_HVT U85 ( .A1(\mem[15][13] ), .A2(n65), .A3(n69), .A4(n66), .Y(n823)
         );
  AO22X1_HVT U86 ( .A1(\mem[15][12] ), .A2(n65), .A3(n70), .A4(n66), .Y(n822)
         );
  AO22X1_HVT U87 ( .A1(\mem[15][11] ), .A2(n65), .A3(n71), .A4(n66), .Y(n821)
         );
  AO22X1_HVT U88 ( .A1(\mem[15][10] ), .A2(n65), .A3(n72), .A4(n66), .Y(n820)
         );
  AO22X1_HVT U89 ( .A1(\mem[15][9] ), .A2(n65), .A3(n73), .A4(n66), .Y(n819)
         );
  AO22X1_HVT U90 ( .A1(\mem[15][8] ), .A2(n65), .A3(n74), .A4(n66), .Y(n818)
         );
  AO22X1_HVT U91 ( .A1(\mem[15][7] ), .A2(n65), .A3(n75), .A4(n66), .Y(n817)
         );
  AO22X1_HVT U92 ( .A1(\mem[15][6] ), .A2(n65), .A3(n76), .A4(n66), .Y(n816)
         );
  AO22X1_HVT U93 ( .A1(\mem[15][5] ), .A2(n65), .A3(n77), .A4(n66), .Y(n815)
         );
  AO22X1_HVT U94 ( .A1(\mem[15][4] ), .A2(n65), .A3(n78), .A4(n66), .Y(n814)
         );
  AO22X1_HVT U95 ( .A1(\mem[15][3] ), .A2(n65), .A3(n79), .A4(n66), .Y(n813)
         );
  AO22X1_HVT U96 ( .A1(\mem[15][2] ), .A2(n65), .A3(n80), .A4(n66), .Y(n812)
         );
  AO22X1_HVT U97 ( .A1(\mem[15][1] ), .A2(n65), .A3(n81), .A4(n66), .Y(n811)
         );
  AO22X1_HVT U98 ( .A1(\mem[15][0] ), .A2(n65), .A3(n82), .A4(n66), .Y(n810)
         );
  AND2X1_HVT U99 ( .A1(n83), .A2(n84), .Y(n66) );
  AO22X1_HVT U100 ( .A1(\mem[14][15] ), .A2(n65), .A3(n85), .A4(n67), .Y(n809)
         );
  AO22X1_HVT U101 ( .A1(\mem[14][14] ), .A2(n65), .A3(n85), .A4(n68), .Y(n808)
         );
  AO22X1_HVT U102 ( .A1(\mem[14][13] ), .A2(n65), .A3(n85), .A4(n69), .Y(n807)
         );
  AO22X1_HVT U103 ( .A1(\mem[14][12] ), .A2(n65), .A3(n85), .A4(n70), .Y(n806)
         );
  AO22X1_HVT U104 ( .A1(\mem[14][11] ), .A2(n65), .A3(n85), .A4(n71), .Y(n805)
         );
  AO22X1_HVT U105 ( .A1(\mem[14][10] ), .A2(n65), .A3(n85), .A4(n72), .Y(n804)
         );
  AO22X1_HVT U106 ( .A1(\mem[14][9] ), .A2(n65), .A3(n85), .A4(n73), .Y(n803)
         );
  AO22X1_HVT U107 ( .A1(\mem[14][8] ), .A2(n65), .A3(n85), .A4(n74), .Y(n802)
         );
  AO22X1_HVT U108 ( .A1(\mem[14][7] ), .A2(n65), .A3(n85), .A4(n75), .Y(n801)
         );
  AO22X1_HVT U109 ( .A1(\mem[14][6] ), .A2(n65), .A3(n85), .A4(n76), .Y(n800)
         );
  AO22X1_HVT U110 ( .A1(\mem[14][5] ), .A2(n65), .A3(n85), .A4(n77), .Y(n799)
         );
  AO22X1_HVT U111 ( .A1(\mem[14][4] ), .A2(n65), .A3(n85), .A4(n78), .Y(n798)
         );
  AO22X1_HVT U112 ( .A1(\mem[14][3] ), .A2(n65), .A3(n85), .A4(n79), .Y(n797)
         );
  AO22X1_HVT U113 ( .A1(\mem[14][2] ), .A2(n65), .A3(n85), .A4(n80), .Y(n796)
         );
  AO22X1_HVT U114 ( .A1(\mem[14][1] ), .A2(n65), .A3(n85), .A4(n81), .Y(n795)
         );
  AO22X1_HVT U115 ( .A1(\mem[14][0] ), .A2(n65), .A3(n85), .A4(n82), .Y(n794)
         );
  AND2X1_HVT U116 ( .A1(n86), .A2(n83), .Y(n85) );
  AO22X1_HVT U117 ( .A1(\mem[13][15] ), .A2(n65), .A3(n87), .A4(n67), .Y(n793)
         );
  AO22X1_HVT U118 ( .A1(\mem[13][14] ), .A2(n65), .A3(n87), .A4(n68), .Y(n792)
         );
  AO22X1_HVT U119 ( .A1(\mem[13][13] ), .A2(n65), .A3(n87), .A4(n69), .Y(n791)
         );
  AO22X1_HVT U120 ( .A1(\mem[13][12] ), .A2(n65), .A3(n87), .A4(n70), .Y(n790)
         );
  AO22X1_HVT U121 ( .A1(\mem[13][11] ), .A2(n65), .A3(n87), .A4(n71), .Y(n789)
         );
  AO22X1_HVT U122 ( .A1(\mem[13][10] ), .A2(n65), .A3(n87), .A4(n72), .Y(n788)
         );
  AO22X1_HVT U123 ( .A1(\mem[13][9] ), .A2(n65), .A3(n87), .A4(n73), .Y(n787)
         );
  AO22X1_HVT U124 ( .A1(\mem[13][8] ), .A2(n65), .A3(n87), .A4(n74), .Y(n786)
         );
  AO22X1_HVT U125 ( .A1(\mem[13][7] ), .A2(n65), .A3(n87), .A4(n75), .Y(n785)
         );
  AO22X1_HVT U126 ( .A1(\mem[13][6] ), .A2(n65), .A3(n87), .A4(n76), .Y(n784)
         );
  AO22X1_HVT U127 ( .A1(\mem[13][5] ), .A2(n65), .A3(n87), .A4(n77), .Y(n783)
         );
  AO22X1_HVT U128 ( .A1(\mem[13][4] ), .A2(n65), .A3(n87), .A4(n78), .Y(n782)
         );
  AO22X1_HVT U129 ( .A1(\mem[13][3] ), .A2(n65), .A3(n87), .A4(n79), .Y(n781)
         );
  AO22X1_HVT U130 ( .A1(\mem[13][2] ), .A2(n65), .A3(n87), .A4(n80), .Y(n780)
         );
  AO22X1_HVT U131 ( .A1(\mem[13][1] ), .A2(n65), .A3(n87), .A4(n81), .Y(n779)
         );
  AO22X1_HVT U132 ( .A1(\mem[13][0] ), .A2(n65), .A3(n87), .A4(n82), .Y(n778)
         );
  AND2X1_HVT U133 ( .A1(n88), .A2(n84), .Y(n87) );
  AO22X1_HVT U134 ( .A1(\mem[12][15] ), .A2(n65), .A3(n89), .A4(n67), .Y(n777)
         );
  AO22X1_HVT U135 ( .A1(\mem[12][14] ), .A2(n65), .A3(n89), .A4(n68), .Y(n776)
         );
  AO22X1_HVT U136 ( .A1(\mem[12][13] ), .A2(n65), .A3(n89), .A4(n69), .Y(n775)
         );
  AO22X1_HVT U137 ( .A1(\mem[12][12] ), .A2(n65), .A3(n89), .A4(n70), .Y(n774)
         );
  AO22X1_HVT U138 ( .A1(\mem[12][11] ), .A2(n65), .A3(n89), .A4(n71), .Y(n773)
         );
  AO22X1_HVT U139 ( .A1(\mem[12][10] ), .A2(n65), .A3(n89), .A4(n72), .Y(n772)
         );
  AO22X1_HVT U140 ( .A1(\mem[12][9] ), .A2(n65), .A3(n89), .A4(n73), .Y(n771)
         );
  AO22X1_HVT U141 ( .A1(\mem[12][8] ), .A2(n65), .A3(n89), .A4(n74), .Y(n770)
         );
  AO22X1_HVT U142 ( .A1(\mem[12][7] ), .A2(n65), .A3(n89), .A4(n75), .Y(n769)
         );
  AO22X1_HVT U143 ( .A1(\mem[12][6] ), .A2(n65), .A3(n89), .A4(n76), .Y(n768)
         );
  AO22X1_HVT U144 ( .A1(\mem[12][5] ), .A2(n65), .A3(n89), .A4(n77), .Y(n767)
         );
  AO22X1_HVT U145 ( .A1(\mem[12][4] ), .A2(n65), .A3(n89), .A4(n78), .Y(n766)
         );
  AO22X1_HVT U146 ( .A1(\mem[12][3] ), .A2(n65), .A3(n89), .A4(n79), .Y(n765)
         );
  AO22X1_HVT U147 ( .A1(\mem[12][2] ), .A2(n65), .A3(n89), .A4(n80), .Y(n764)
         );
  AO22X1_HVT U148 ( .A1(\mem[12][1] ), .A2(n65), .A3(n89), .A4(n81), .Y(n763)
         );
  AO22X1_HVT U149 ( .A1(\mem[12][0] ), .A2(n65), .A3(n89), .A4(n82), .Y(n762)
         );
  AND2X1_HVT U150 ( .A1(n88), .A2(n86), .Y(n89) );
  AO22X1_HVT U151 ( .A1(\mem[11][15] ), .A2(n65), .A3(n90), .A4(n67), .Y(n761)
         );
  AO22X1_HVT U152 ( .A1(\mem[11][14] ), .A2(n65), .A3(n90), .A4(n68), .Y(n760)
         );
  AO22X1_HVT U153 ( .A1(\mem[11][13] ), .A2(n65), .A3(n90), .A4(n69), .Y(n759)
         );
  AO22X1_HVT U154 ( .A1(\mem[11][12] ), .A2(n65), .A3(n90), .A4(n70), .Y(n758)
         );
  AO22X1_HVT U155 ( .A1(\mem[11][11] ), .A2(n65), .A3(n90), .A4(n71), .Y(n757)
         );
  AO22X1_HVT U156 ( .A1(\mem[11][10] ), .A2(n65), .A3(n90), .A4(n72), .Y(n756)
         );
  AO22X1_HVT U157 ( .A1(\mem[11][9] ), .A2(n65), .A3(n90), .A4(n73), .Y(n755)
         );
  AO22X1_HVT U158 ( .A1(\mem[11][8] ), .A2(n65), .A3(n90), .A4(n74), .Y(n754)
         );
  AO22X1_HVT U159 ( .A1(\mem[11][7] ), .A2(n65), .A3(n90), .A4(n75), .Y(n753)
         );
  AO22X1_HVT U160 ( .A1(\mem[11][6] ), .A2(n65), .A3(n90), .A4(n76), .Y(n752)
         );
  AO22X1_HVT U161 ( .A1(\mem[11][5] ), .A2(n65), .A3(n90), .A4(n77), .Y(n751)
         );
  AO22X1_HVT U162 ( .A1(\mem[11][4] ), .A2(n65), .A3(n90), .A4(n78), .Y(n750)
         );
  AO22X1_HVT U163 ( .A1(\mem[11][3] ), .A2(n65), .A3(n90), .A4(n79), .Y(n749)
         );
  AO22X1_HVT U164 ( .A1(\mem[11][2] ), .A2(n65), .A3(n90), .A4(n80), .Y(n748)
         );
  AO22X1_HVT U165 ( .A1(\mem[11][1] ), .A2(n65), .A3(n90), .A4(n81), .Y(n747)
         );
  AO22X1_HVT U166 ( .A1(\mem[11][0] ), .A2(n65), .A3(n90), .A4(n82), .Y(n746)
         );
  AND2X1_HVT U167 ( .A1(n91), .A2(n84), .Y(n90) );
  AO22X1_HVT U168 ( .A1(\mem[10][15] ), .A2(n65), .A3(n92), .A4(n67), .Y(n745)
         );
  AO22X1_HVT U169 ( .A1(\mem[10][14] ), .A2(n65), .A3(n92), .A4(n68), .Y(n744)
         );
  AO22X1_HVT U170 ( .A1(\mem[10][13] ), .A2(n65), .A3(n92), .A4(n69), .Y(n743)
         );
  AO22X1_HVT U171 ( .A1(\mem[10][12] ), .A2(n65), .A3(n92), .A4(n70), .Y(n742)
         );
  AO22X1_HVT U172 ( .A1(\mem[10][11] ), .A2(n65), .A3(n92), .A4(n71), .Y(n741)
         );
  AO22X1_HVT U173 ( .A1(\mem[10][10] ), .A2(n65), .A3(n92), .A4(n72), .Y(n740)
         );
  AO22X1_HVT U174 ( .A1(\mem[10][9] ), .A2(n65), .A3(n92), .A4(n73), .Y(n739)
         );
  AO22X1_HVT U175 ( .A1(\mem[10][8] ), .A2(n65), .A3(n92), .A4(n74), .Y(n738)
         );
  AO22X1_HVT U176 ( .A1(\mem[10][7] ), .A2(n65), .A3(n92), .A4(n75), .Y(n737)
         );
  AO22X1_HVT U177 ( .A1(\mem[10][6] ), .A2(n65), .A3(n92), .A4(n76), .Y(n736)
         );
  AO22X1_HVT U178 ( .A1(\mem[10][5] ), .A2(n65), .A3(n92), .A4(n77), .Y(n735)
         );
  AO22X1_HVT U179 ( .A1(\mem[10][4] ), .A2(n65), .A3(n92), .A4(n78), .Y(n734)
         );
  AO22X1_HVT U180 ( .A1(\mem[10][3] ), .A2(n65), .A3(n92), .A4(n79), .Y(n733)
         );
  AO22X1_HVT U181 ( .A1(\mem[10][2] ), .A2(n65), .A3(n92), .A4(n80), .Y(n732)
         );
  AO22X1_HVT U182 ( .A1(\mem[10][1] ), .A2(n65), .A3(n92), .A4(n81), .Y(n731)
         );
  AO22X1_HVT U183 ( .A1(\mem[10][0] ), .A2(n65), .A3(n92), .A4(n82), .Y(n730)
         );
  AND2X1_HVT U184 ( .A1(n91), .A2(n86), .Y(n92) );
  AO22X1_HVT U185 ( .A1(\mem[9][15] ), .A2(n65), .A3(n93), .A4(n67), .Y(n729)
         );
  AO22X1_HVT U186 ( .A1(\mem[9][14] ), .A2(n65), .A3(n93), .A4(n68), .Y(n728)
         );
  AO22X1_HVT U187 ( .A1(\mem[9][13] ), .A2(n65), .A3(n93), .A4(n69), .Y(n727)
         );
  AO22X1_HVT U188 ( .A1(\mem[9][12] ), .A2(n65), .A3(n93), .A4(n70), .Y(n726)
         );
  AO22X1_HVT U189 ( .A1(\mem[9][11] ), .A2(n65), .A3(n93), .A4(n71), .Y(n725)
         );
  AO22X1_HVT U190 ( .A1(\mem[9][10] ), .A2(n65), .A3(n93), .A4(n72), .Y(n724)
         );
  AO22X1_HVT U191 ( .A1(\mem[9][9] ), .A2(n65), .A3(n93), .A4(n73), .Y(n723)
         );
  AO22X1_HVT U192 ( .A1(\mem[9][8] ), .A2(n65), .A3(n93), .A4(n74), .Y(n722)
         );
  AO22X1_HVT U193 ( .A1(\mem[9][7] ), .A2(n65), .A3(n93), .A4(n75), .Y(n721)
         );
  AO22X1_HVT U194 ( .A1(\mem[9][6] ), .A2(n65), .A3(n93), .A4(n76), .Y(n720)
         );
  AO22X1_HVT U195 ( .A1(\mem[9][5] ), .A2(n65), .A3(n93), .A4(n77), .Y(n719)
         );
  AO22X1_HVT U196 ( .A1(\mem[9][4] ), .A2(n65), .A3(n93), .A4(n78), .Y(n718)
         );
  AO22X1_HVT U197 ( .A1(\mem[9][3] ), .A2(n65), .A3(n93), .A4(n79), .Y(n717)
         );
  AO22X1_HVT U198 ( .A1(\mem[9][2] ), .A2(n65), .A3(n93), .A4(n80), .Y(n716)
         );
  AO22X1_HVT U199 ( .A1(\mem[9][1] ), .A2(n65), .A3(n93), .A4(n81), .Y(n715)
         );
  AO22X1_HVT U200 ( .A1(\mem[9][0] ), .A2(n65), .A3(n93), .A4(n82), .Y(n714)
         );
  AND2X1_HVT U201 ( .A1(n94), .A2(n84), .Y(n93) );
  AND2X1_HVT U202 ( .A1(a_din[0]), .A2(n95), .Y(n84) );
  AO22X1_HVT U203 ( .A1(\mem[8][15] ), .A2(n65), .A3(n96), .A4(n67), .Y(n713)
         );
  AO22X1_HVT U204 ( .A1(\mem[8][14] ), .A2(n65), .A3(n96), .A4(n68), .Y(n712)
         );
  AO22X1_HVT U205 ( .A1(\mem[8][13] ), .A2(n65), .A3(n96), .A4(n69), .Y(n711)
         );
  AO22X1_HVT U206 ( .A1(\mem[8][12] ), .A2(n65), .A3(n96), .A4(n70), .Y(n710)
         );
  AO22X1_HVT U207 ( .A1(\mem[8][11] ), .A2(n65), .A3(n96), .A4(n71), .Y(n709)
         );
  AO22X1_HVT U208 ( .A1(\mem[8][10] ), .A2(n65), .A3(n96), .A4(n72), .Y(n708)
         );
  AO22X1_HVT U209 ( .A1(\mem[8][9] ), .A2(n65), .A3(n96), .A4(n73), .Y(n707)
         );
  AO22X1_HVT U210 ( .A1(\mem[8][8] ), .A2(n65), .A3(n96), .A4(n74), .Y(n706)
         );
  AO22X1_HVT U211 ( .A1(\mem[8][7] ), .A2(n65), .A3(n96), .A4(n75), .Y(n705)
         );
  AO22X1_HVT U212 ( .A1(\mem[8][6] ), .A2(n65), .A3(n96), .A4(n76), .Y(n704)
         );
  AO22X1_HVT U213 ( .A1(\mem[8][5] ), .A2(n65), .A3(n96), .A4(n77), .Y(n703)
         );
  AO22X1_HVT U214 ( .A1(\mem[8][4] ), .A2(n65), .A3(n96), .A4(n78), .Y(n702)
         );
  AO22X1_HVT U215 ( .A1(\mem[8][3] ), .A2(n65), .A3(n96), .A4(n79), .Y(n701)
         );
  AO22X1_HVT U216 ( .A1(\mem[8][2] ), .A2(n65), .A3(n96), .A4(n80), .Y(n700)
         );
  AO22X1_HVT U217 ( .A1(\mem[8][1] ), .A2(n65), .A3(n96), .A4(n81), .Y(n699)
         );
  AO22X1_HVT U218 ( .A1(\mem[8][0] ), .A2(n65), .A3(n96), .A4(n82), .Y(n698)
         );
  AND2X1_HVT U219 ( .A1(n94), .A2(n86), .Y(n96) );
  AND2X1_HVT U220 ( .A1(n95), .A2(n97), .Y(n86) );
  AND2X1_HVT U221 ( .A1(write), .A2(a_din[3]), .Y(n95) );
  AO22X1_HVT U222 ( .A1(\mem[7][15] ), .A2(n65), .A3(n98), .A4(n67), .Y(n697)
         );
  AO22X1_HVT U223 ( .A1(\mem[7][14] ), .A2(n65), .A3(n98), .A4(n68), .Y(n696)
         );
  AO22X1_HVT U224 ( .A1(\mem[7][13] ), .A2(n65), .A3(n98), .A4(n69), .Y(n695)
         );
  AO22X1_HVT U225 ( .A1(\mem[7][12] ), .A2(n65), .A3(n98), .A4(n70), .Y(n694)
         );
  AO22X1_HVT U226 ( .A1(\mem[7][11] ), .A2(n65), .A3(n98), .A4(n71), .Y(n693)
         );
  AO22X1_HVT U227 ( .A1(\mem[7][10] ), .A2(n65), .A3(n98), .A4(n72), .Y(n692)
         );
  AO22X1_HVT U228 ( .A1(\mem[7][9] ), .A2(n65), .A3(n98), .A4(n73), .Y(n691)
         );
  AO22X1_HVT U229 ( .A1(\mem[7][8] ), .A2(n65), .A3(n98), .A4(n74), .Y(n690)
         );
  AO22X1_HVT U230 ( .A1(\mem[7][7] ), .A2(n65), .A3(n98), .A4(n75), .Y(n689)
         );
  AO22X1_HVT U231 ( .A1(\mem[7][6] ), .A2(n65), .A3(n98), .A4(n76), .Y(n688)
         );
  AO22X1_HVT U232 ( .A1(\mem[7][5] ), .A2(n65), .A3(n98), .A4(n77), .Y(n687)
         );
  AO22X1_HVT U233 ( .A1(\mem[7][4] ), .A2(n65), .A3(n98), .A4(n78), .Y(n686)
         );
  AO22X1_HVT U234 ( .A1(\mem[7][3] ), .A2(n65), .A3(n98), .A4(n79), .Y(n685)
         );
  AO22X1_HVT U235 ( .A1(\mem[7][2] ), .A2(n65), .A3(n98), .A4(n80), .Y(n684)
         );
  AO22X1_HVT U236 ( .A1(\mem[7][1] ), .A2(n65), .A3(n98), .A4(n81), .Y(n683)
         );
  AO22X1_HVT U237 ( .A1(\mem[7][0] ), .A2(n65), .A3(n98), .A4(n82), .Y(n682)
         );
  AND2X1_HVT U238 ( .A1(n99), .A2(n83), .Y(n98) );
  AO22X1_HVT U239 ( .A1(\mem[6][15] ), .A2(n65), .A3(n100), .A4(n67), .Y(n681)
         );
  AO22X1_HVT U240 ( .A1(\mem[6][14] ), .A2(n65), .A3(n100), .A4(n68), .Y(n680)
         );
  AO22X1_HVT U241 ( .A1(\mem[6][13] ), .A2(n65), .A3(n100), .A4(n69), .Y(n679)
         );
  AO22X1_HVT U242 ( .A1(\mem[6][12] ), .A2(n65), .A3(n100), .A4(n70), .Y(n678)
         );
  AO22X1_HVT U243 ( .A1(\mem[6][11] ), .A2(n65), .A3(n100), .A4(n71), .Y(n677)
         );
  AO22X1_HVT U244 ( .A1(\mem[6][10] ), .A2(n65), .A3(n100), .A4(n72), .Y(n676)
         );
  AO22X1_HVT U245 ( .A1(\mem[6][9] ), .A2(n65), .A3(n100), .A4(n73), .Y(n675)
         );
  AO22X1_HVT U246 ( .A1(\mem[6][8] ), .A2(n65), .A3(n100), .A4(n74), .Y(n674)
         );
  AO22X1_HVT U247 ( .A1(\mem[6][7] ), .A2(n65), .A3(n100), .A4(n75), .Y(n673)
         );
  AO22X1_HVT U248 ( .A1(\mem[6][6] ), .A2(n65), .A3(n100), .A4(n76), .Y(n672)
         );
  AO22X1_HVT U249 ( .A1(\mem[6][5] ), .A2(n65), .A3(n100), .A4(n77), .Y(n671)
         );
  AO22X1_HVT U250 ( .A1(\mem[6][4] ), .A2(n65), .A3(n100), .A4(n78), .Y(n670)
         );
  AO22X1_HVT U251 ( .A1(\mem[6][3] ), .A2(n65), .A3(n100), .A4(n79), .Y(n669)
         );
  AO22X1_HVT U252 ( .A1(\mem[6][2] ), .A2(n65), .A3(n100), .A4(n80), .Y(n668)
         );
  AO22X1_HVT U253 ( .A1(\mem[6][1] ), .A2(n65), .A3(n100), .A4(n81), .Y(n667)
         );
  AO22X1_HVT U254 ( .A1(\mem[6][0] ), .A2(n65), .A3(n100), .A4(n82), .Y(n666)
         );
  AND2X1_HVT U255 ( .A1(n101), .A2(n83), .Y(n100) );
  AND2X1_HVT U256 ( .A1(a_din[2]), .A2(a_din[1]), .Y(n83) );
  AO22X1_HVT U257 ( .A1(\mem[5][15] ), .A2(n65), .A3(n102), .A4(n67), .Y(n665)
         );
  AO22X1_HVT U258 ( .A1(\mem[5][14] ), .A2(n65), .A3(n102), .A4(n68), .Y(n664)
         );
  AO22X1_HVT U259 ( .A1(\mem[5][13] ), .A2(n65), .A3(n102), .A4(n69), .Y(n663)
         );
  AO22X1_HVT U260 ( .A1(\mem[5][12] ), .A2(n65), .A3(n102), .A4(n70), .Y(n662)
         );
  AO22X1_HVT U261 ( .A1(\mem[5][11] ), .A2(n65), .A3(n102), .A4(n71), .Y(n661)
         );
  AO22X1_HVT U262 ( .A1(\mem[5][10] ), .A2(n65), .A3(n102), .A4(n72), .Y(n660)
         );
  AO22X1_HVT U263 ( .A1(\mem[5][9] ), .A2(n65), .A3(n102), .A4(n73), .Y(n659)
         );
  AO22X1_HVT U264 ( .A1(\mem[5][8] ), .A2(n65), .A3(n102), .A4(n74), .Y(n658)
         );
  AO22X1_HVT U265 ( .A1(\mem[5][7] ), .A2(n65), .A3(n102), .A4(n75), .Y(n657)
         );
  AO22X1_HVT U266 ( .A1(\mem[5][6] ), .A2(n65), .A3(n102), .A4(n76), .Y(n656)
         );
  AO22X1_HVT U267 ( .A1(\mem[5][5] ), .A2(n65), .A3(n102), .A4(n77), .Y(n655)
         );
  AO22X1_HVT U268 ( .A1(\mem[5][4] ), .A2(n65), .A3(n102), .A4(n78), .Y(n654)
         );
  AO22X1_HVT U269 ( .A1(\mem[5][3] ), .A2(n65), .A3(n102), .A4(n79), .Y(n653)
         );
  AO22X1_HVT U270 ( .A1(\mem[5][2] ), .A2(n65), .A3(n102), .A4(n80), .Y(n652)
         );
  AO22X1_HVT U271 ( .A1(\mem[5][1] ), .A2(n65), .A3(n102), .A4(n81), .Y(n651)
         );
  AO22X1_HVT U272 ( .A1(\mem[5][0] ), .A2(n65), .A3(n102), .A4(n82), .Y(n650)
         );
  AND2X1_HVT U273 ( .A1(n99), .A2(n88), .Y(n102) );
  AO22X1_HVT U274 ( .A1(\mem[4][15] ), .A2(n65), .A3(n103), .A4(n67), .Y(n649)
         );
  AO22X1_HVT U275 ( .A1(\mem[4][14] ), .A2(n65), .A3(n103), .A4(n68), .Y(n648)
         );
  AO22X1_HVT U276 ( .A1(\mem[4][13] ), .A2(n65), .A3(n103), .A4(n69), .Y(n647)
         );
  AO22X1_HVT U277 ( .A1(\mem[4][12] ), .A2(n65), .A3(n103), .A4(n70), .Y(n646)
         );
  AO22X1_HVT U278 ( .A1(\mem[4][11] ), .A2(n65), .A3(n103), .A4(n71), .Y(n645)
         );
  AO22X1_HVT U279 ( .A1(\mem[4][10] ), .A2(n65), .A3(n103), .A4(n72), .Y(n644)
         );
  AO22X1_HVT U280 ( .A1(\mem[4][9] ), .A2(n65), .A3(n103), .A4(n73), .Y(n643)
         );
  AO22X1_HVT U281 ( .A1(\mem[4][8] ), .A2(n65), .A3(n103), .A4(n74), .Y(n642)
         );
  AO22X1_HVT U282 ( .A1(\mem[4][7] ), .A2(n65), .A3(n103), .A4(n75), .Y(n641)
         );
  AO22X1_HVT U283 ( .A1(\mem[4][6] ), .A2(n65), .A3(n103), .A4(n76), .Y(n640)
         );
  AO22X1_HVT U284 ( .A1(\mem[4][5] ), .A2(n65), .A3(n103), .A4(n77), .Y(n639)
         );
  AO22X1_HVT U285 ( .A1(\mem[4][4] ), .A2(n65), .A3(n103), .A4(n78), .Y(n638)
         );
  AO22X1_HVT U286 ( .A1(\mem[4][3] ), .A2(n65), .A3(n103), .A4(n79), .Y(n637)
         );
  AO22X1_HVT U287 ( .A1(\mem[4][2] ), .A2(n65), .A3(n103), .A4(n80), .Y(n636)
         );
  AO22X1_HVT U288 ( .A1(\mem[4][1] ), .A2(n65), .A3(n103), .A4(n81), .Y(n635)
         );
  AO22X1_HVT U289 ( .A1(\mem[4][0] ), .A2(n65), .A3(n103), .A4(n82), .Y(n634)
         );
  AND2X1_HVT U290 ( .A1(n101), .A2(n88), .Y(n103) );
  AND2X1_HVT U291 ( .A1(a_din[2]), .A2(n104), .Y(n88) );
  AO22X1_HVT U292 ( .A1(\mem[3][15] ), .A2(n65), .A3(n105), .A4(n67), .Y(n633)
         );
  AO22X1_HVT U293 ( .A1(\mem[3][14] ), .A2(n65), .A3(n105), .A4(n68), .Y(n632)
         );
  AO22X1_HVT U294 ( .A1(\mem[3][13] ), .A2(n65), .A3(n105), .A4(n69), .Y(n631)
         );
  AO22X1_HVT U295 ( .A1(\mem[3][12] ), .A2(n65), .A3(n105), .A4(n70), .Y(n630)
         );
  AO22X1_HVT U296 ( .A1(\mem[3][11] ), .A2(n65), .A3(n105), .A4(n71), .Y(n629)
         );
  AO22X1_HVT U297 ( .A1(\mem[3][10] ), .A2(n65), .A3(n105), .A4(n72), .Y(n628)
         );
  AO22X1_HVT U298 ( .A1(\mem[3][9] ), .A2(n65), .A3(n105), .A4(n73), .Y(n627)
         );
  AO22X1_HVT U299 ( .A1(\mem[3][8] ), .A2(n65), .A3(n105), .A4(n74), .Y(n626)
         );
  AO22X1_HVT U300 ( .A1(\mem[3][7] ), .A2(n65), .A3(n105), .A4(n75), .Y(n625)
         );
  AO22X1_HVT U301 ( .A1(\mem[3][6] ), .A2(n65), .A3(n105), .A4(n76), .Y(n624)
         );
  AO22X1_HVT U302 ( .A1(\mem[3][5] ), .A2(n65), .A3(n105), .A4(n77), .Y(n623)
         );
  AO22X1_HVT U303 ( .A1(\mem[3][4] ), .A2(n65), .A3(n105), .A4(n78), .Y(n622)
         );
  AO22X1_HVT U304 ( .A1(\mem[3][3] ), .A2(n65), .A3(n105), .A4(n79), .Y(n621)
         );
  AO22X1_HVT U305 ( .A1(\mem[3][2] ), .A2(n65), .A3(n105), .A4(n80), .Y(n620)
         );
  AO22X1_HVT U306 ( .A1(\mem[3][1] ), .A2(n65), .A3(n105), .A4(n81), .Y(n619)
         );
  AO22X1_HVT U307 ( .A1(\mem[3][0] ), .A2(n65), .A3(n105), .A4(n82), .Y(n618)
         );
  AND2X1_HVT U308 ( .A1(n99), .A2(n91), .Y(n105) );
  AO22X1_HVT U309 ( .A1(\mem[2][15] ), .A2(n65), .A3(n106), .A4(n67), .Y(n617)
         );
  AO22X1_HVT U310 ( .A1(\mem[2][14] ), .A2(n65), .A3(n106), .A4(n68), .Y(n616)
         );
  AO22X1_HVT U311 ( .A1(\mem[2][13] ), .A2(n65), .A3(n106), .A4(n69), .Y(n615)
         );
  AO22X1_HVT U312 ( .A1(\mem[2][12] ), .A2(n65), .A3(n106), .A4(n70), .Y(n614)
         );
  AO22X1_HVT U313 ( .A1(\mem[2][11] ), .A2(n65), .A3(n106), .A4(n71), .Y(n613)
         );
  AO22X1_HVT U314 ( .A1(\mem[2][10] ), .A2(n65), .A3(n106), .A4(n72), .Y(n612)
         );
  AO22X1_HVT U315 ( .A1(\mem[2][9] ), .A2(n65), .A3(n106), .A4(n73), .Y(n611)
         );
  AO22X1_HVT U316 ( .A1(\mem[2][8] ), .A2(n65), .A3(n106), .A4(n74), .Y(n610)
         );
  AO22X1_HVT U317 ( .A1(\mem[2][7] ), .A2(n65), .A3(n106), .A4(n75), .Y(n609)
         );
  AO22X1_HVT U318 ( .A1(\mem[2][6] ), .A2(n65), .A3(n106), .A4(n76), .Y(n608)
         );
  AO22X1_HVT U319 ( .A1(\mem[2][5] ), .A2(n65), .A3(n106), .A4(n77), .Y(n607)
         );
  AO22X1_HVT U320 ( .A1(\mem[2][4] ), .A2(n65), .A3(n106), .A4(n78), .Y(n606)
         );
  AO22X1_HVT U321 ( .A1(\mem[2][3] ), .A2(n65), .A3(n106), .A4(n79), .Y(n605)
         );
  AO22X1_HVT U322 ( .A1(\mem[2][2] ), .A2(n65), .A3(n106), .A4(n80), .Y(n604)
         );
  AO22X1_HVT U323 ( .A1(\mem[2][1] ), .A2(n65), .A3(n106), .A4(n81), .Y(n603)
         );
  AO22X1_HVT U324 ( .A1(\mem[2][0] ), .A2(n65), .A3(n106), .A4(n82), .Y(n602)
         );
  AND2X1_HVT U325 ( .A1(n101), .A2(n91), .Y(n106) );
  AND2X1_HVT U326 ( .A1(a_din[1]), .A2(n107), .Y(n91) );
  AO22X1_HVT U327 ( .A1(\mem[1][15] ), .A2(n65), .A3(n108), .A4(n67), .Y(n601)
         );
  AO22X1_HVT U328 ( .A1(\mem[1][14] ), .A2(n65), .A3(n108), .A4(n68), .Y(n600)
         );
  AO22X1_HVT U329 ( .A1(\mem[1][13] ), .A2(n65), .A3(n108), .A4(n69), .Y(n599)
         );
  AO22X1_HVT U330 ( .A1(\mem[1][12] ), .A2(n65), .A3(n108), .A4(n70), .Y(n598)
         );
  AO22X1_HVT U331 ( .A1(\mem[1][11] ), .A2(n65), .A3(n108), .A4(n71), .Y(n597)
         );
  AO22X1_HVT U332 ( .A1(\mem[1][10] ), .A2(n65), .A3(n108), .A4(n72), .Y(n596)
         );
  AO22X1_HVT U333 ( .A1(\mem[1][9] ), .A2(n65), .A3(n108), .A4(n73), .Y(n595)
         );
  AO22X1_HVT U334 ( .A1(\mem[1][8] ), .A2(n65), .A3(n108), .A4(n74), .Y(n594)
         );
  AO22X1_HVT U335 ( .A1(\mem[1][7] ), .A2(n65), .A3(n108), .A4(n75), .Y(n593)
         );
  AO22X1_HVT U336 ( .A1(\mem[1][6] ), .A2(n65), .A3(n108), .A4(n76), .Y(n592)
         );
  AO22X1_HVT U337 ( .A1(\mem[1][5] ), .A2(n65), .A3(n108), .A4(n77), .Y(n591)
         );
  AO22X1_HVT U338 ( .A1(\mem[1][4] ), .A2(n65), .A3(n108), .A4(n78), .Y(n590)
         );
  AO22X1_HVT U339 ( .A1(\mem[1][3] ), .A2(n65), .A3(n108), .A4(n79), .Y(n589)
         );
  AO22X1_HVT U340 ( .A1(\mem[1][2] ), .A2(n65), .A3(n108), .A4(n80), .Y(n588)
         );
  AO22X1_HVT U341 ( .A1(\mem[1][1] ), .A2(n65), .A3(n108), .A4(n81), .Y(n587)
         );
  AO22X1_HVT U342 ( .A1(\mem[1][0] ), .A2(n65), .A3(n108), .A4(n82), .Y(n586)
         );
  AND2X1_HVT U343 ( .A1(n99), .A2(n94), .Y(n108) );
  AND2X1_HVT U344 ( .A1(n109), .A2(a_din[0]), .Y(n99) );
  AO22X1_HVT U345 ( .A1(\mem[0][15] ), .A2(n65), .A3(n110), .A4(n67), .Y(n585)
         );
  AND2X1_HVT U346 ( .A1(n111), .A2(n112), .Y(n67) );
  AO22X1_HVT U347 ( .A1(\mem[0][14] ), .A2(n65), .A3(n110), .A4(n68), .Y(n584)
         );
  AND2X1_HVT U348 ( .A1(n113), .A2(n111), .Y(n68) );
  AO22X1_HVT U349 ( .A1(\mem[0][13] ), .A2(n65), .A3(n110), .A4(n69), .Y(n583)
         );
  AND2X1_HVT U350 ( .A1(n114), .A2(n111), .Y(n69) );
  AO22X1_HVT U351 ( .A1(\mem[0][12] ), .A2(n65), .A3(n110), .A4(n70), .Y(n582)
         );
  AND2X1_HVT U352 ( .A1(n115), .A2(n111), .Y(n70) );
  AND2X1_HVT U353 ( .A1(a_addr[3]), .A2(a_addr[2]), .Y(n111) );
  AO22X1_HVT U354 ( .A1(\mem[0][11] ), .A2(n65), .A3(n110), .A4(n71), .Y(n581)
         );
  AND2X1_HVT U355 ( .A1(n116), .A2(n112), .Y(n71) );
  AO22X1_HVT U356 ( .A1(\mem[0][10] ), .A2(n65), .A3(n110), .A4(n72), .Y(n580)
         );
  AND2X1_HVT U357 ( .A1(n116), .A2(n113), .Y(n72) );
  AO22X1_HVT U358 ( .A1(\mem[0][9] ), .A2(n65), .A3(n110), .A4(n73), .Y(n579)
         );
  AND2X1_HVT U359 ( .A1(n116), .A2(n114), .Y(n73) );
  AO22X1_HVT U360 ( .A1(\mem[0][8] ), .A2(n65), .A3(n110), .A4(n74), .Y(n578)
         );
  AND2X1_HVT U361 ( .A1(n116), .A2(n115), .Y(n74) );
  AND2X1_HVT U362 ( .A1(a_addr[3]), .A2(n117), .Y(n116) );
  AO22X1_HVT U363 ( .A1(\mem[0][7] ), .A2(n65), .A3(n110), .A4(n75), .Y(n577)
         );
  AND2X1_HVT U364 ( .A1(n118), .A2(n112), .Y(n75) );
  AO22X1_HVT U365 ( .A1(\mem[0][6] ), .A2(n65), .A3(n110), .A4(n76), .Y(n576)
         );
  AND2X1_HVT U366 ( .A1(n118), .A2(n113), .Y(n76) );
  AO22X1_HVT U367 ( .A1(\mem[0][5] ), .A2(n65), .A3(n110), .A4(n77), .Y(n575)
         );
  AND2X1_HVT U368 ( .A1(n118), .A2(n114), .Y(n77) );
  AO22X1_HVT U369 ( .A1(\mem[0][4] ), .A2(n65), .A3(n110), .A4(n78), .Y(n574)
         );
  AND2X1_HVT U370 ( .A1(n118), .A2(n115), .Y(n78) );
  AND2X1_HVT U371 ( .A1(a_addr[2]), .A2(n119), .Y(n118) );
  AO22X1_HVT U372 ( .A1(\mem[0][3] ), .A2(n65), .A3(n110), .A4(n79), .Y(n573)
         );
  AND2X1_HVT U373 ( .A1(n120), .A2(n112), .Y(n79) );
  AND3X1_HVT U374 ( .A1(a_addr[0]), .A2(n65), .A3(a_addr[1]), .Y(n112) );
  AO22X1_HVT U375 ( .A1(\mem[0][2] ), .A2(n65), .A3(n110), .A4(n80), .Y(n572)
         );
  AND2X1_HVT U376 ( .A1(n120), .A2(n113), .Y(n80) );
  AND3X1_HVT U377 ( .A1(n121), .A2(n65), .A3(a_addr[1]), .Y(n113) );
  AO22X1_HVT U378 ( .A1(\mem[0][1] ), .A2(n65), .A3(n110), .A4(n81), .Y(n571)
         );
  AND2X1_HVT U379 ( .A1(n120), .A2(n114), .Y(n81) );
  AND3X1_HVT U380 ( .A1(n122), .A2(n65), .A3(a_addr[0]), .Y(n114) );
  AO22X1_HVT U381 ( .A1(\mem[0][0] ), .A2(n65), .A3(n110), .A4(n82), .Y(n570)
         );
  AND2X1_HVT U382 ( .A1(n120), .A2(n115), .Y(n82) );
  AND3X1_HVT U383 ( .A1(n122), .A2(n65), .A3(n121), .Y(n115) );
  INVX0_HVT U384 ( .A(a_addr[0]), .Y(n121) );
  INVX0_HVT U385 ( .A(a_addr[1]), .Y(n122) );
  AND2X1_HVT U386 ( .A1(n117), .A2(n119), .Y(n120) );
  INVX0_HVT U387 ( .A(a_addr[3]), .Y(n119) );
  INVX0_HVT U388 ( .A(a_addr[2]), .Y(n117) );
  AND2X1_HVT U389 ( .A1(n101), .A2(n94), .Y(n110) );
  AND2X1_HVT U390 ( .A1(n104), .A2(n107), .Y(n94) );
  INVX0_HVT U391 ( .A(a_din[2]), .Y(n107) );
  INVX0_HVT U392 ( .A(a_din[1]), .Y(n104) );
  AND2X1_HVT U393 ( .A1(n109), .A2(n97), .Y(n101) );
  INVX0_HVT U394 ( .A(a_din[0]), .Y(n97) );
  AND2X1_HVT U395 ( .A1(write), .A2(n123), .Y(n109) );
  INVX0_HVT U396 ( .A(a_din[3]), .Y(n123) );
  INVX0_HVT U397 ( .A(rst), .Y(n65) );
endmodule

