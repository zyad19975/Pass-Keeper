
module sbox_11 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n50, n210, n211, n212, n213, n216, n217, n218, n219, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594;

  NAND2X0_HVT U4 ( .A1(n299), .A2(n592), .Y(n591) );
  NAND2X0_HVT U5 ( .A1(n249), .A2(n291), .Y(n589) );
  NAND2X0_HVT U13 ( .A1(n581), .A2(n303), .Y(n582) );
  NAND2X0_HVT U15 ( .A1(n592), .A2(n242), .Y(n579) );
  NAND2X0_HVT U21 ( .A1(n299), .A2(n309), .Y(n573) );
  NAND2X0_HVT U24 ( .A1(n210), .A2(n309), .Y(n571) );
  NAND2X0_HVT U33 ( .A1(n370), .A2(n309), .Y(n562) );
  NAND2X0_HVT U35 ( .A1(n293), .A2(n309), .Y(n560) );
  NAND2X0_HVT U42 ( .A1(n248), .A2(n210), .Y(n553) );
  MUX41X1_HVT U51 ( .A1(n358), .A3(n316), .A2(n333), .A4(n334), .S0(n314), 
        .S1(n287), .Y(n546) );
  NAND2X0_HVT U53 ( .A1(n543), .A2(n552), .Y(n544) );
  NAND2X0_HVT U56 ( .A1(n299), .A2(n539), .Y(n540) );
  NAND2X0_HVT U58 ( .A1(n303), .A2(n592), .Y(n537) );
  MUX41X1_HVT U59 ( .A1(n280), .A3(n537), .A2(n278), .A4(n332), .S0(n314), 
        .S1(n287), .Y(n536) );
  MUX41X1_HVT U61 ( .A1(n277), .A3(n331), .A2(n259), .A4(n238), .S0(n314), 
        .S1(n287), .Y(n534) );
  NAND2X0_HVT U62 ( .A1(n309), .A2(n302), .Y(n533) );
  MUX41X1_HVT U63 ( .A1(n533), .A3(n323), .A2(n353), .A4(n330), .S0(n314), 
        .S1(n287), .Y(n532) );
  AO21X1_HVT U66 ( .A1(n328), .A2(n287), .A3(n352), .Y(n529) );
  MUX41X1_HVT U68 ( .A1(n326), .A3(n529), .A2(n528), .A4(n530), .S0(n281), 
        .S1(n48), .Y(n527) );
  MUX41X1_HVT U69 ( .A1(n527), .A3(n535), .A2(n531), .A4(n541), .S0(in[6]), 
        .S1(n294), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n297), .A2(n522), .Y(n523) );
  MUX41X1_HVT U74 ( .A1(n524), .A3(n569), .A2(n523), .A4(n571), .S0(n283), 
        .S1(n313), .Y(n521) );
  MUX41X1_HVT U75 ( .A1(n356), .A3(n361), .A2(n374), .A4(n336), .S0(n281), 
        .S1(n313), .Y(n520) );
  MUX41X1_HVT U82 ( .A1(n550), .A3(n334), .A2(n317), .A4(n580), .S0(n281), 
        .S1(n313), .Y(n512) );
  AND2X1_HVT U83 ( .A1(n249), .A2(n269), .Y(n511) );
  MUX41X1_HVT U84 ( .A1(n335), .A3(n235), .A2(n578), .A4(n511), .S0(n281), 
        .S1(n313), .Y(n510) );
  NAND2X0_HVT U85 ( .A1(n309), .A2(n373), .Y(n509) );
  MUX41X1_HVT U86 ( .A1(n361), .A3(n509), .A2(n275), .A4(n273), .S0(n281), 
        .S1(n313), .Y(n508) );
  MUX41X1_HVT U87 ( .A1(n508), .A3(n512), .A2(n510), .A4(n513), .S0(in[0]), 
        .S1(n286), .Y(n507) );
  MUX41X1_HVT U90 ( .A1(n549), .A3(n553), .A2(n358), .A4(n506), .S0(n282), 
        .S1(n268), .Y(n505) );
  AO21X1_HVT U93 ( .A1(n290), .A2(n501), .A3(n357), .Y(n502) );
  MUX41X1_HVT U96 ( .A1(n317), .A3(n276), .A2(n360), .A4(n499), .S0(n281), 
        .S1(n268), .Y(n498) );
  MUX41X1_HVT U97 ( .A1(n356), .A3(n276), .A2(n305), .A4(n579), .S0(n281), 
        .S1(n244), .Y(n497) );
  MUX41X1_HVT U98 ( .A1(n497), .A3(n500), .A2(n498), .A4(n505), .S0(n294), 
        .S1(n286), .Y(n496) );
  NAND2X0_HVT U101 ( .A1(n492), .A2(n491), .Y(n493) );
  MUX41X1_HVT U103 ( .A1(n592), .A3(n327), .A2(n339), .A4(n560), .S0(n281), 
        .S1(n268), .Y(n489) );
  MUX41X1_HVT U105 ( .A1(n338), .A3(n548), .A2(n488), .A4(n355), .S0(n281), 
        .S1(n268), .Y(n487) );
  OA21X1_HVT U109 ( .A1(n346), .A2(n312), .A3(n332), .Y(n484) );
  NAND2X0_HVT U110 ( .A1(n301), .A2(n482), .Y(n483) );
  MUX41X1_HVT U114 ( .A1(n479), .A3(n485), .A2(n481), .A4(n484), .S0(in[5]), 
        .S1(n244), .Y(n478) );
  AND2X1_HVT U115 ( .A1(n248), .A2(n239), .Y(n477) );
  AO21X1_HVT U118 ( .A1(n284), .A2(n296), .A3(n235), .Y(n474) );
  NAND2X0_HVT U123 ( .A1(n468), .A2(n467), .Y(n469) );
  MUX41X1_HVT U125 ( .A1(n573), .A3(n280), .A2(n326), .A4(n365), .S0(n282), 
        .S1(n263), .Y(n465) );
  AND3X1_HVT U128 ( .A1(n285), .A2(n309), .A3(n269), .Y(n462) );
  MUX41X1_HVT U131 ( .A1(n460), .A3(n462), .A2(n461), .A4(n463), .S0(in[5]), 
        .S1(n314), .Y(n459) );
  MUX41X1_HVT U132 ( .A1(n459), .A3(n472), .A2(n464), .A4(n478), .S0(in[6]), 
        .S1(in[0]), .Y(out[3]) );
  MUX41X1_HVT U136 ( .A1(n273), .A3(n562), .A2(n367), .A4(n559), .S0(n282), 
        .S1(n314), .Y(n455) );
  MUX41X1_HVT U139 ( .A1(n453), .A3(n456), .A2(n455), .A4(n457), .S0(n294), 
        .S1(n286), .Y(n452) );
  AND2X1_HVT U140 ( .A1(n296), .A2(n308), .Y(n451) );
  MUX41X1_HVT U141 ( .A1(n570), .A3(n347), .A2(n451), .A4(n343), .S0(n283), 
        .S1(n263), .Y(n450) );
  MUX41X1_HVT U142 ( .A1(n335), .A3(n243), .A2(n354), .A4(n296), .S0(n282), 
        .S1(n263), .Y(n449) );
  NAND2X0_HVT U146 ( .A1(n304), .A2(n303), .Y(n522) );
  MUX41X1_HVT U147 ( .A1(n367), .A3(n522), .A2(n356), .A4(n549), .S0(n283), 
        .S1(n314), .Y(n445) );
  MUX41X1_HVT U148 ( .A1(n445), .A3(n449), .A2(n446), .A4(n450), .S0(n294), 
        .S1(n286), .Y(n444) );
  MUX41X1_HVT U153 ( .A1(n483), .A3(n277), .A2(n300), .A4(n319), .S0(n282), 
        .S1(n244), .Y(n439) );
  AND2X1_HVT U154 ( .A1(n290), .A2(n210), .Y(n438) );
  NAND2X0_HVT U158 ( .A1(n248), .A2(n373), .Y(n434) );
  MUX41X1_HVT U159 ( .A1(n582), .A3(n239), .A2(n434), .A4(n325), .S0(n311), 
        .S1(n244), .Y(n433) );
  MUX41X1_HVT U160 ( .A1(n433), .A3(n439), .A2(n435), .A4(n440), .S0(n294), 
        .S1(n288), .Y(n432) );
  AND2X1_HVT U162 ( .A1(n234), .A2(n522), .Y(n430) );
  MUX41X1_HVT U163 ( .A1(n331), .A3(n430), .A2(n274), .A4(n431), .S0(n311), 
        .S1(n244), .Y(n429) );
  MUX41X1_HVT U165 ( .A1(n573), .A3(n340), .A2(n549), .A4(n428), .S0(n314), 
        .S1(n311), .Y(n427) );
  NAND2X0_HVT U166 ( .A1(n303), .A2(n539), .Y(n426) );
  NAND2X0_HVT U167 ( .A1(n374), .A2(n309), .Y(n425) );
  MUX41X1_HVT U168 ( .A1(n359), .A3(n296), .A2(n425), .A4(n426), .S0(n311), 
        .S1(n244), .Y(n424) );
  MUX41X1_HVT U172 ( .A1(n421), .A3(n427), .A2(n424), .A4(n429), .S0(in[0]), 
        .S1(n286), .Y(n420) );
  NAND2X0_HVT U174 ( .A1(n304), .A2(n235), .Y(n581) );
  MUX41X1_HVT U176 ( .A1(n245), .A3(n419), .A2(n364), .A4(n581), .S0(n314), 
        .S1(n310), .Y(n418) );
  NAND2X0_HVT U177 ( .A1(n248), .A2(n292), .Y(n417) );
  MUX41X1_HVT U178 ( .A1(n577), .A3(n417), .A2(n368), .A4(n557), .S0(n283), 
        .S1(n244), .Y(n416) );
  MUX41X1_HVT U179 ( .A1(n567), .A3(n369), .A2(n321), .A4(n368), .S0(n311), 
        .S1(n244), .Y(n415) );
  MUX41X1_HVT U180 ( .A1(n324), .A3(n586), .A2(n582), .A4(n272), .S0(n314), 
        .S1(n311), .Y(n414) );
  MUX41X1_HVT U181 ( .A1(n414), .A3(n416), .A2(n415), .A4(n418), .S0(n294), 
        .S1(n288), .Y(n413) );
  MUX41X1_HVT U182 ( .A1(n348), .A3(n590), .A2(n350), .A4(n337), .S0(n314), 
        .S1(n310), .Y(n412) );
  MUX41X1_HVT U189 ( .A1(n406), .A3(n581), .A2(n407), .A4(n355), .S0(n268), 
        .S1(n311), .Y(n405) );
  MUX41X1_HVT U190 ( .A1(n405), .A3(n408), .A2(n409), .A4(n412), .S0(n288), 
        .S1(in[0]), .Y(n404) );
  MUX21X2_HVT U191 ( .A1(n404), .A2(n413), .S0(in[6]), .Y(out[6]) );
  MUX41X1_HVT U195 ( .A1(n234), .A3(n360), .A2(n594), .A4(n558), .S0(n311), 
        .S1(n313), .Y(n400) );
  AO21X1_HVT U197 ( .A1(n275), .A2(n289), .A3(n357), .Y(n398) );
  MUX41X1_HVT U199 ( .A1(n397), .A3(n401), .A2(n400), .A4(n402), .S0(in[0]), 
        .S1(n288), .Y(n396) );
  MUX41X1_HVT U204 ( .A1(n540), .A3(n582), .A2(n344), .A4(n572), .S0(n311), 
        .S1(n313), .Y(n391) );
  MUX41X1_HVT U205 ( .A1(n269), .A3(n592), .A2(n369), .A4(n342), .S0(n311), 
        .S1(n313), .Y(n390) );
  MUX41X1_HVT U206 ( .A1(n390), .A3(n392), .A2(n391), .A4(n393), .S0(n294), 
        .S1(n288), .Y(n389) );
  NAND2X0_HVT U208 ( .A1(n304), .A2(n299), .Y(n482) );
  NAND2X0_HVT U212 ( .A1(n257), .A2(n297), .Y(n539) );
  NAND2X0_HVT U214 ( .A1(n235), .A2(n309), .Y(n388) );
  NAND2X0_HVT U215 ( .A1(n482), .A2(n298), .Y(n387) );
  AO21X1_HVT U216 ( .A1(n308), .A2(n371), .A3(n315), .Y(n492) );
  NAND2X0_HVT U218 ( .A1(n371), .A2(n305), .Y(n441) );
  NAND2X0_HVT U220 ( .A1(n289), .A2(n388), .Y(n514) );
  IBUFFX4_HVT U1 ( .A(n315), .Y(n313) );
  MUX21X2_HVT U2 ( .A1(n302), .A2(n480), .S0(n23), .Y(n479) );
  IBUFFX16_HVT U3 ( .A(n271), .Y(n23) );
  INVX1_HVT U6 ( .A(n253), .Y(n48) );
  INVX2_HVT U7 ( .A(n263), .Y(n253) );
  NBUFFX2_HVT U8 ( .A(in[7]), .Y(n244) );
  IBUFFX2_HVT U9 ( .A(n311), .Y(n50) );
  MUX41X1_HVT U10 ( .A1(n556), .A3(n276), .A2(n549), .A4(n522), .S0(n50), .S1(
        n244), .Y(n408) );
  MUX21X1_HVT U11 ( .A1(n526), .A2(n551), .S0(n264), .Y(n525) );
  XOR2X1_HVT U12 ( .A1(n265), .A2(n568), .Y(n551) );
  INVX0_HVT U14 ( .A(n305), .Y(n218) );
  INVX1_HVT U16 ( .A(n312), .Y(n311) );
  IBUFFX2_HVT U17 ( .A(n372), .Y(n210) );
  INVX1_HVT U18 ( .A(in[3]), .Y(n372) );
  NAND2X0_HVT U19 ( .A1(n536), .A2(n211), .Y(n212) );
  NAND2X0_HVT U20 ( .A1(n538), .A2(n216), .Y(n213) );
  NAND2X0_HVT U22 ( .A1(n212), .A2(n213), .Y(n535) );
  INVX0_HVT U23 ( .A(n216), .Y(n211) );
  IBUFFX2_HVT U25 ( .A(n264), .Y(n216) );
  INVX2_HVT U26 ( .A(n312), .Y(n310) );
  MUX21X2_HVT U27 ( .A1(n420), .A2(n432), .S0(in[6]), .Y(out[5]) );
  MUX21X1_HVT U28 ( .A1(n594), .A2(n300), .S0(n218), .Y(n217) );
  IBUFFX16_HVT U29 ( .A(n217), .Y(n568) );
  MUX41X1_HVT U30 ( .A1(n568), .A3(n589), .A2(n371), .A4(n366), .S0(n219), 
        .S1(n253), .Y(n456) );
  IBUFFX16_HVT U31 ( .A(n283), .Y(n219) );
  IBUFFX2_HVT U32 ( .A(n315), .Y(n314) );
  INVX2_HVT U34 ( .A(in[7]), .Y(n315) );
  IBUFFX2_HVT U36 ( .A(n588), .Y(n231) );
  IBUFFX2_HVT U37 ( .A(n588), .Y(n232) );
  IBUFFX2_HVT U38 ( .A(n588), .Y(n233) );
  INVX1_HVT U39 ( .A(n233), .Y(n234) );
  INVX1_HVT U40 ( .A(n233), .Y(n235) );
  INVX1_HVT U41 ( .A(n231), .Y(n236) );
  INVX1_HVT U43 ( .A(n231), .Y(n237) );
  INVX1_HVT U44 ( .A(n236), .Y(n238) );
  INVX1_HVT U45 ( .A(n237), .Y(n239) );
  INVX1_HVT U46 ( .A(n232), .Y(n240) );
  INVX1_HVT U47 ( .A(n232), .Y(n241) );
  INVX1_HVT U48 ( .A(n240), .Y(n242) );
  INVX1_HVT U49 ( .A(n241), .Y(n243) );
  XOR2X1_HVT U50 ( .A1(n375), .A2(in[3]), .Y(n588) );
  MUX21X2_HVT U52 ( .A1(n572), .A2(n348), .S0(n289), .Y(n454) );
  IBUFFX2_HVT U54 ( .A(n587), .Y(n326) );
  MUX21X2_HVT U55 ( .A1(n373), .A2(n243), .S0(n246), .Y(n587) );
  INVX1_HVT U57 ( .A(in[7]), .Y(n265) );
  OA21X1_HVT U60 ( .A1(n278), .A2(n315), .A3(n564), .Y(n422) );
  INVX1_HVT U64 ( .A(in[4]), .Y(n245) );
  IBUFFX16_HVT U65 ( .A(n304), .Y(n246) );
  MUX21X2_HVT U67 ( .A1(n395), .A2(n394), .S0(n247), .Y(n393) );
  IBUFFX16_HVT U70 ( .A(n284), .Y(n247) );
  MUX21X1_HVT U71 ( .A1(n272), .A2(n578), .S0(n265), .Y(n395) );
  INVX0_HVT U72 ( .A(n308), .Y(n248) );
  INVX0_HVT U76 ( .A(n308), .Y(n249) );
  INVX0_HVT U77 ( .A(n308), .Y(n307) );
  MUX41X1_HVT U78 ( .A1(n553), .A3(n560), .A2(n547), .A4(n403), .S0(in[2]), 
        .S1(n313), .Y(n402) );
  INVX1_HVT U79 ( .A(n245), .Y(n269) );
  INVX1_HVT U80 ( .A(in[4]), .Y(n375) );
  INVX2_HVT U81 ( .A(n308), .Y(n305) );
  MUX21X2_HVT U88 ( .A1(n277), .A2(n495), .S0(n250), .Y(n494) );
  XOR2X1_HVT U89 ( .A1(n310), .A2(n263), .Y(n250) );
  MUX41X1_HVT U91 ( .A1(n494), .A3(n489), .A2(n490), .A4(n487), .S0(n251), 
        .S1(n252), .Y(n486) );
  IBUFFX16_HVT U92 ( .A(in[0]), .Y(n251) );
  IBUFFX16_HVT U94 ( .A(n286), .Y(n252) );
  MUX41X1_HVT U95 ( .A1(n296), .A3(n366), .A2(n568), .A4(n554), .S0(n253), 
        .S1(n254), .Y(n401) );
  IBUFFX16_HVT U99 ( .A(in[2]), .Y(n254) );
  IBUFFX16_HVT U100 ( .A(n308), .Y(n304) );
  NAND2X2_HVT U102 ( .A1(n304), .A2(n301), .Y(n592) );
  MUX21X2_HVT U104 ( .A1(n534), .A2(n532), .S0(n255), .Y(n531) );
  IBUFFX16_HVT U106 ( .A(n284), .Y(n255) );
  NBUFFX2_HVT U107 ( .A(n307), .Y(n256) );
  NBUFFX2_HVT U108 ( .A(n307), .Y(n257) );
  NBUFFX2_HVT U111 ( .A(n307), .Y(n258) );
  IBUFFX2_HVT U112 ( .A(n308), .Y(n306) );
  INVX0_HVT U113 ( .A(n574), .Y(n334) );
  AND3X1_HVT U116 ( .A1(n301), .A2(n539), .A3(n514), .Y(n515) );
  INVX1_HVT U117 ( .A(n315), .Y(n268) );
  INVX1_HVT U119 ( .A(n265), .Y(n263) );
  INVX1_HVT U120 ( .A(n282), .Y(n264) );
  INVX0_HVT U121 ( .A(in[6]), .Y(n267) );
  INVX1_HVT U122 ( .A(n287), .Y(n266) );
  INVX0_HVT U124 ( .A(n559), .Y(n345) );
  INVX0_HVT U126 ( .A(n259), .Y(n578) );
  MUX21X2_HVT U127 ( .A1(n298), .A2(n574), .S0(n265), .Y(n516) );
  MUX21X1_HVT U129 ( .A1(n234), .A2(n295), .S0(n258), .Y(n259) );
  NAND2X0_HVT U130 ( .A1(n496), .A2(n260), .Y(n261) );
  NAND2X0_HVT U133 ( .A1(n486), .A2(n267), .Y(n262) );
  NAND2X0_HVT U134 ( .A1(n261), .A2(n262), .Y(out[2]) );
  INVX1_HVT U135 ( .A(n267), .Y(n260) );
  MUX21X2_HVT U137 ( .A1(n318), .A2(n471), .S0(n283), .Y(n470) );
  MUX21X1_HVT U138 ( .A1(n483), .A2(n564), .S0(n264), .Y(n481) );
  MUX21X2_HVT U143 ( .A1(n465), .A2(n466), .S0(in[5]), .Y(n464) );
  IBUFFX2_HVT U144 ( .A(n554), .Y(n350) );
  MUX41X1_HVT U145 ( .A1(n564), .A3(n336), .A2(n477), .A4(n582), .S0(n264), 
        .S1(n265), .Y(n476) );
  MUX41X1_HVT U149 ( .A1(n584), .A3(n540), .A2(n575), .A4(n359), .S0(n315), 
        .S1(n266), .Y(n538) );
  MUX21X2_HVT U150 ( .A1(n448), .A2(n447), .S0(n285), .Y(n446) );
  MUX21X2_HVT U151 ( .A1(n515), .A2(n516), .S0(n264), .Y(n513) );
  IBUFFX2_HVT U152 ( .A(n584), .Y(n328) );
  MUX21X2_HVT U155 ( .A1(n546), .A2(n542), .S0(n264), .Y(n541) );
  MUX21X2_HVT U156 ( .A1(n473), .A2(n476), .S0(in[5]), .Y(n472) );
  MUX21X2_HVT U157 ( .A1(n396), .A2(n389), .S0(n267), .Y(out[7]) );
  OA21X1_HVT U161 ( .A1(n320), .A2(n315), .A3(n564), .Y(n447) );
  MUX21X2_HVT U164 ( .A1(n436), .A2(n437), .S0(n284), .Y(n435) );
  INVX2_HVT U169 ( .A(in[1]), .Y(n308) );
  INVX0_HVT U170 ( .A(in[0]), .Y(n270) );
  OA21X1_HVT U171 ( .A1(n587), .A2(n265), .A3(n347), .Y(n394) );
  OA21X1_HVT U173 ( .A1(n561), .A2(n265), .A3(n335), .Y(n410) );
  OA21X1_HVT U175 ( .A1(n555), .A2(n265), .A3(n441), .Y(n442) );
  INVX2_HVT U183 ( .A(in[2]), .Y(n312) );
  NBUFFX2_HVT U184 ( .A(n310), .Y(n282) );
  MUX41X1_HVT U185 ( .A1(n362), .A3(n519), .A2(n363), .A4(n586), .S0(n265), 
        .S1(n312), .Y(n518) );
  MUX41X1_HVT U186 ( .A1(n525), .A3(n520), .A2(n521), .A4(n518), .S0(n270), 
        .S1(n266), .Y(n517) );
  MUX41X1_HVT U187 ( .A1(n563), .A3(n583), .A2(n349), .A4(n559), .S0(n312), 
        .S1(n265), .Y(n392) );
  MUX21X2_HVT U188 ( .A1(n444), .A2(n452), .S0(in[6]), .Y(out[4]) );
  XOR2X1_HVT U192 ( .A1(n308), .A2(n312), .Y(n271) );
  MUX21X2_HVT U193 ( .A1(n507), .A2(n517), .S0(in[6]), .Y(out[1]) );
  INVX1_HVT U194 ( .A(n590), .Y(n370) );
  MUX21X1_HVT U196 ( .A1(n274), .A2(n259), .S0(n282), .Y(n461) );
  AND2X1_HVT U198 ( .A1(n239), .A2(n539), .Y(n272) );
  INVX1_HVT U200 ( .A(n300), .Y(n374) );
  MUX21X1_HVT U201 ( .A1(n370), .A2(n373), .S0(in[5]), .Y(n543) );
  NBUFFX2_HVT U202 ( .A(n590), .Y(n299) );
  MUX21X1_HVT U203 ( .A1(n327), .A2(n371), .S0(in[5]), .Y(n528) );
  AND2X1_HVT U207 ( .A1(n301), .A2(n522), .Y(n273) );
  MUX21X1_HVT U209 ( .A1(n301), .A2(n238), .S0(n248), .Y(n554) );
  MUX21X1_HVT U210 ( .A1(n470), .A2(n469), .S0(n290), .Y(n466) );
  MUX21X1_HVT U211 ( .A1(n299), .A2(n235), .S0(n249), .Y(n558) );
  MUX21X1_HVT U213 ( .A1(n238), .A2(n293), .S0(n305), .Y(n491) );
  MUX21X1_HVT U217 ( .A1(n454), .A2(n591), .S0(n284), .Y(n453) );
  MUX21X1_HVT U219 ( .A1(n370), .A2(n374), .S0(n248), .Y(n419) );
  MUX21X1_HVT U221 ( .A1(n243), .A2(n370), .S0(n249), .Y(n499) );
  MUX21X1_HVT U222 ( .A1(n373), .A2(n370), .S0(n249), .Y(n557) );
  MUX21X1_HVT U223 ( .A1(n291), .A2(n374), .S0(n249), .Y(n555) );
  MUX21X1_HVT U224 ( .A1(n373), .A2(n242), .S0(n256), .Y(n431) );
  NAND2X0_HVT U225 ( .A1(n245), .A2(n372), .Y(n590) );
  MUX21X1_HVT U226 ( .A1(n234), .A2(n371), .S0(n306), .Y(n379) );
  NBUFFX2_HVT U227 ( .A(n593), .Y(n300) );
  MUX21X1_HVT U228 ( .A1(n235), .A2(n374), .S0(n248), .Y(n570) );
  MUX21X1_HVT U229 ( .A1(n299), .A2(n298), .S0(n249), .Y(n506) );
  MUX21X1_HVT U230 ( .A1(n234), .A2(n293), .S0(n257), .Y(n519) );
  XOR2X1_HVT U231 ( .A1(n234), .A2(n258), .Y(n549) );
  INVX1_HVT U232 ( .A(n594), .Y(n373) );
  MUX21X1_HVT U233 ( .A1(n373), .A2(n291), .S0(n257), .Y(n561) );
  MUX21X1_HVT U234 ( .A1(n293), .A2(n370), .S0(n305), .Y(n566) );
  MUX21X1_HVT U235 ( .A1(n474), .A2(n475), .S0(n289), .Y(n473) );
  MUX21X1_HVT U236 ( .A1(n319), .A2(n344), .S0(n282), .Y(n475) );
  MUX21X1_HVT U237 ( .A1(n341), .A2(n458), .S0(n285), .Y(n457) );
  MUX21X1_HVT U238 ( .A1(n365), .A2(n298), .S0(n289), .Y(n458) );
  NBUFFX2_HVT U239 ( .A(n593), .Y(n301) );
  MUX21X1_HVT U240 ( .A1(n291), .A2(n293), .S0(n306), .Y(n403) );
  XOR2X1_HVT U241 ( .A1(n300), .A2(n258), .Y(n547) );
  MUX21X1_HVT U242 ( .A1(n370), .A2(n292), .S0(n256), .Y(n380) );
  MUX21X1_HVT U243 ( .A1(n291), .A2(n234), .S0(n257), .Y(n382) );
  INVX1_HVT U244 ( .A(n296), .Y(n371) );
  MUX21X1_HVT U245 ( .A1(n302), .A2(n297), .S0(n249), .Y(n580) );
  MUX21X1_HVT U246 ( .A1(n590), .A2(n303), .S0(n306), .Y(n501) );
  MUX21X1_HVT U247 ( .A1(n299), .A2(n291), .S0(n258), .Y(n583) );
  MUX21X1_HVT U248 ( .A1(n371), .A2(n370), .S0(n258), .Y(n576) );
  MUX21X1_HVT U249 ( .A1(n342), .A2(n580), .S0(n284), .Y(n495) );
  MUX21X1_HVT U250 ( .A1(n292), .A2(n291), .S0(n306), .Y(n471) );
  NBUFFX2_HVT U251 ( .A(n593), .Y(n302) );
  MUX21X1_HVT U252 ( .A1(n291), .A2(n303), .S0(n305), .Y(n406) );
  MUX21X1_HVT U253 ( .A1(n594), .A2(n301), .S0(n248), .Y(n407) );
  MUX21X1_HVT U254 ( .A1(n594), .A2(n297), .S0(n248), .Y(n564) );
  MUX21X1_HVT U255 ( .A1(n291), .A2(n373), .S0(n304), .Y(n584) );
  XOR2X1_HVT U256 ( .A1(n258), .A2(n371), .Y(n550) );
  MUX21X1_HVT U257 ( .A1(n300), .A2(n292), .S0(n257), .Y(n386) );
  XNOR2X1_HVT U258 ( .A1(n590), .A2(n257), .Y(n274) );
  XNOR2X1_HVT U259 ( .A1(n594), .A2(n257), .Y(n275) );
  AND2X1_HVT U260 ( .A1(n257), .A2(n374), .Y(n276) );
  MUX21X1_HVT U261 ( .A1(n297), .A2(n291), .S0(n258), .Y(n384) );
  AND2X1_HVT U262 ( .A1(n303), .A2(n482), .Y(n277) );
  MUX21X1_HVT U263 ( .A1(n300), .A2(n299), .S0(n249), .Y(n378) );
  MUX21X1_HVT U264 ( .A1(n298), .A2(n292), .S0(n305), .Y(n524) );
  MUX21X1_HVT U265 ( .A1(n298), .A2(n303), .S0(n285), .Y(n468) );
  XOR2X1_HVT U266 ( .A1(n245), .A2(n306), .Y(n569) );
  NBUFFX2_HVT U267 ( .A(n268), .Y(n289) );
  NBUFFX2_HVT U268 ( .A(n268), .Y(n290) );
  NBUFFX2_HVT U269 ( .A(n372), .Y(n291) );
  NBUFFX2_HVT U270 ( .A(n310), .Y(n283) );
  NBUFFX2_HVT U271 ( .A(in[5]), .Y(n288) );
  NBUFFX2_HVT U272 ( .A(n310), .Y(n285) );
  NBUFFX2_HVT U273 ( .A(n310), .Y(n284) );
  NBUFFX2_HVT U274 ( .A(in[5]), .Y(n287) );
  NBUFFX2_HVT U275 ( .A(n285), .Y(n281) );
  NBUFFX2_HVT U276 ( .A(in[5]), .Y(n286) );
  MUX21X1_HVT U277 ( .A1(n238), .A2(n295), .S0(n249), .Y(n572) );
  MUX21X1_HVT U278 ( .A1(n493), .A2(n341), .S0(n285), .Y(n490) );
  MUX21X1_HVT U279 ( .A1(n410), .A2(n411), .S0(n284), .Y(n409) );
  MUX21X1_HVT U280 ( .A1(n509), .A2(n210), .S0(n289), .Y(n411) );
  XOR2X1_HVT U281 ( .A1(n306), .A2(in[3]), .Y(n548) );
  MUX21X1_HVT U282 ( .A1(n297), .A2(n239), .S0(n258), .Y(n488) );
  NAND2X0_HVT U283 ( .A1(n295), .A2(n293), .Y(n593) );
  NBUFFX2_HVT U284 ( .A(n375), .Y(n293) );
  MUX21X1_HVT U285 ( .A1(n423), .A2(n422), .S0(n285), .Y(n421) );
  MUX21X1_HVT U286 ( .A1(n298), .A2(n360), .S0(n290), .Y(n423) );
  AND2X1_HVT U287 ( .A1(n242), .A2(n309), .Y(n278) );
  MUX21X1_HVT U288 ( .A1(n210), .A2(n370), .S0(n306), .Y(n556) );
  MUX21X1_HVT U289 ( .A1(n442), .A2(n443), .S0(n284), .Y(n440) );
  MUX21X1_HVT U290 ( .A1(n362), .A2(n371), .S0(n289), .Y(n443) );
  MUX21X1_HVT U291 ( .A1(n373), .A2(n360), .S0(n290), .Y(n526) );
  MUX21X1_HVT U292 ( .A1(n566), .A2(n322), .S0(n290), .Y(n448) );
  MUX21X1_HVT U293 ( .A1(n371), .A2(n374), .S0(n305), .Y(n428) );
  NBUFFX2_HVT U294 ( .A(n585), .Y(n296) );
  MUX21X1_HVT U295 ( .A1(n374), .A2(n210), .S0(n258), .Y(n575) );
  MUX21X1_HVT U296 ( .A1(n345), .A2(n592), .S0(n283), .Y(n485) );
  MUX21X1_HVT U297 ( .A1(n438), .A2(n302), .S0(n279), .Y(n437) );
  MUX21X1_HVT U298 ( .A1(n557), .A2(n363), .S0(n289), .Y(n436) );
  MUX21X1_HVT U299 ( .A1(n577), .A2(n343), .S0(n283), .Y(n460) );
  MUX21X1_HVT U300 ( .A1(n544), .A2(n545), .S0(n290), .Y(n542) );
  MUX21X1_HVT U301 ( .A1(n210), .A2(n560), .S0(n287), .Y(n545) );
  XOR2X1_HVT U302 ( .A1(n258), .A2(n288), .Y(n552) );
  MUX21X1_HVT U303 ( .A1(n592), .A2(n308), .S0(n284), .Y(n467) );
  NBUFFX2_HVT U304 ( .A(n585), .Y(n297) );
  MUX21X1_HVT U305 ( .A1(n351), .A2(n368), .S0(n289), .Y(n399) );
  MUX21X1_HVT U306 ( .A1(n210), .A2(n371), .S0(n257), .Y(n383) );
  MUX21X1_HVT U307 ( .A1(n565), .A2(n387), .S0(n289), .Y(n381) );
  MUX21X1_HVT U308 ( .A1(n299), .A2(n295), .S0(n248), .Y(n586) );
  MUX21X1_HVT U309 ( .A1(n329), .A2(n309), .S0(n286), .Y(n530) );
  NBUFFX2_HVT U310 ( .A(n594), .Y(n303) );
  MUX21X1_HVT U311 ( .A1(n338), .A2(n565), .S0(n283), .Y(n463) );
  MUX21X1_HVT U312 ( .A1(n302), .A2(n504), .S0(n279), .Y(n503) );
  MUX21X1_HVT U313 ( .A1(n295), .A2(n292), .S0(n290), .Y(n504) );
  NBUFFX2_HVT U314 ( .A(n585), .Y(n298) );
  NBUFFX2_HVT U315 ( .A(n375), .Y(n292) );
  XNOR2X1_HVT U316 ( .A1(n265), .A2(n304), .Y(n279) );
  AND2X1_HVT U317 ( .A1(n291), .A2(n309), .Y(n280) );
  MUX21X1_HVT U318 ( .A1(n399), .A2(n398), .S0(n284), .Y(n397) );
  MUX21X1_HVT U319 ( .A1(n502), .A2(n503), .S0(n285), .Y(n500) );
  MUX21X1_HVT U320 ( .A1(n370), .A2(n269), .S0(n305), .Y(n563) );
  NAND2X0_HVT U321 ( .A1(in[3]), .A2(in[4]), .Y(n594) );
  MUX21X1_HVT U322 ( .A1(n269), .A2(n373), .S0(n306), .Y(n559) );
  NAND2X0_HVT U323 ( .A1(in[4]), .A2(n372), .Y(n585) );
  MUX21X1_HVT U324 ( .A1(n269), .A2(n235), .S0(n257), .Y(n385) );
  MUX21X1_HVT U325 ( .A1(n269), .A2(n371), .S0(n305), .Y(n577) );
  MUX21X1_HVT U326 ( .A1(n269), .A2(n302), .S0(n304), .Y(n574) );
  MUX21X1_HVT U327 ( .A1(n269), .A2(n297), .S0(n304), .Y(n377) );
  MUX21X1_HVT U328 ( .A1(n269), .A2(n303), .S0(n248), .Y(n376) );
  MUX21X1_HVT U329 ( .A1(n303), .A2(n269), .S0(n306), .Y(n567) );
  MUX21X1_HVT U330 ( .A1(n295), .A2(n269), .S0(n282), .Y(n480) );
  MUX21X1_HVT U331 ( .A1(n291), .A2(n269), .S0(n304), .Y(n565) );
  INVX0_HVT U332 ( .A(n256), .Y(n309) );
  NBUFFX2_HVT U333 ( .A(in[3]), .Y(n295) );
  NBUFFX2_HVT U334 ( .A(in[0]), .Y(n294) );
  INVX0_HVT U335 ( .A(n573), .Y(n316) );
  INVX0_HVT U336 ( .A(n571), .Y(n317) );
  INVX0_HVT U337 ( .A(n562), .Y(n318) );
  INVX0_HVT U338 ( .A(n560), .Y(n319) );
  INVX0_HVT U339 ( .A(n425), .Y(n320) );
  INVX0_HVT U340 ( .A(n388), .Y(n321) );
  INVX0_HVT U341 ( .A(n592), .Y(n322) );
  INVX0_HVT U342 ( .A(n579), .Y(n323) );
  INVX0_HVT U343 ( .A(n591), .Y(n324) );
  INVX0_HVT U344 ( .A(n589), .Y(n325) );
  INVX0_HVT U345 ( .A(n586), .Y(n327) );
  INVX0_HVT U346 ( .A(n583), .Y(n329) );
  INVX0_HVT U347 ( .A(n580), .Y(n330) );
  INVX0_HVT U348 ( .A(n577), .Y(n331) );
  INVX0_HVT U349 ( .A(n576), .Y(n332) );
  INVX0_HVT U350 ( .A(n575), .Y(n333) );
  INVX0_HVT U351 ( .A(n572), .Y(n335) );
  INVX0_HVT U352 ( .A(n570), .Y(n336) );
  INVX0_HVT U353 ( .A(n569), .Y(n337) );
  INVX0_HVT U354 ( .A(n567), .Y(n338) );
  INVX0_HVT U355 ( .A(n566), .Y(n339) );
  INVX0_HVT U356 ( .A(n565), .Y(n340) );
  INVX0_HVT U357 ( .A(n381), .Y(n341) );
  INVX0_HVT U358 ( .A(n564), .Y(n342) );
  INVX0_HVT U359 ( .A(n563), .Y(n343) );
  INVX0_HVT U360 ( .A(n561), .Y(n344) );
  INVX0_HVT U361 ( .A(n558), .Y(n346) );
  INVX0_HVT U362 ( .A(n557), .Y(n347) );
  INVX0_HVT U363 ( .A(n556), .Y(n348) );
  INVX0_HVT U364 ( .A(n555), .Y(n349) );
  INVX0_HVT U365 ( .A(n553), .Y(n351) );
  INVX0_HVT U366 ( .A(n522), .Y(n352) );
  INVX0_HVT U367 ( .A(n582), .Y(n353) );
  INVX0_HVT U368 ( .A(n482), .Y(n354) );
  INVX0_HVT U369 ( .A(n387), .Y(n355) );
  INVX0_HVT U370 ( .A(n539), .Y(n356) );
  INVX0_HVT U371 ( .A(n441), .Y(n357) );
  INVX0_HVT U372 ( .A(n386), .Y(n358) );
  INVX0_HVT U373 ( .A(n385), .Y(n359) );
  INVX0_HVT U374 ( .A(n384), .Y(n360) );
  INVX0_HVT U375 ( .A(n383), .Y(n361) );
  INVX0_HVT U376 ( .A(n382), .Y(n362) );
  INVX0_HVT U377 ( .A(n501), .Y(n363) );
  INVX0_HVT U378 ( .A(n491), .Y(n364) );
  INVX0_HVT U379 ( .A(n380), .Y(n365) );
  INVX0_HVT U380 ( .A(n379), .Y(n366) );
  INVX0_HVT U381 ( .A(n378), .Y(n367) );
  INVX0_HVT U382 ( .A(n377), .Y(n368) );
  INVX0_HVT U383 ( .A(n376), .Y(n369) );
endmodule

