
module sbox_6 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n48, n203, n204, n205, n210, n211, n212, n213, n216, n217, n218,
         n219, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608;

  NAND2X0_HVT U3 ( .A1(n218), .A2(n317), .Y(n606) );
  NAND2X0_HVT U4 ( .A1(n315), .A2(n272), .Y(n605) );
  NAND2X0_HVT U5 ( .A1(n322), .A2(n300), .Y(n603) );
  NAND2X0_HVT U15 ( .A1(n271), .A2(n204), .Y(n593) );
  NAND2X0_HVT U21 ( .A1(n315), .A2(n326), .Y(n587) );
  NAND2X0_HVT U24 ( .A1(n310), .A2(n326), .Y(n585) );
  NAND2X0_HVT U33 ( .A1(n386), .A2(n326), .Y(n576) );
  NAND2X0_HVT U35 ( .A1(n305), .A2(n326), .Y(n574) );
  NAND2X0_HVT U42 ( .A1(n23), .A2(n310), .Y(n567) );
  MUX41X1_HVT U51 ( .A1(n374), .A3(n333), .A2(n350), .A4(n351), .S0(n330), 
        .S1(n295), .Y(n559) );
  NAND2X0_HVT U53 ( .A1(n556), .A2(n566), .Y(n557) );
  NAND2X0_HVT U56 ( .A1(n315), .A2(n552), .Y(n553) );
  MUX41X1_HVT U57 ( .A1(n375), .A3(n589), .A2(n553), .A4(n598), .S0(n330), 
        .S1(in[5]), .Y(n551) );
  NAND2X0_HVT U58 ( .A1(n320), .A2(n272), .Y(n550) );
  MUX41X1_HVT U59 ( .A1(n288), .A3(n550), .A2(n286), .A4(n349), .S0(n330), 
        .S1(in[5]), .Y(n549) );
  MUX41X1_HVT U61 ( .A1(n284), .A3(n348), .A2(n347), .A4(n262), .S0(n330), 
        .S1(n328), .Y(n547) );
  NAND2X0_HVT U62 ( .A1(n326), .A2(n318), .Y(n546) );
  MUX41X1_HVT U63 ( .A1(n546), .A3(n339), .A2(n369), .A4(n346), .S0(n330), 
        .S1(in[5]), .Y(n545) );
  AO21X1_HVT U66 ( .A1(n344), .A2(n296), .A3(n368), .Y(n542) );
  MUX41X1_HVT U68 ( .A1(n342), .A3(n542), .A2(n541), .A4(n543), .S0(n289), 
        .S1(n205), .Y(n540) );
  MUX41X1_HVT U69 ( .A1(n540), .A3(n548), .A2(n544), .A4(n554), .S0(in[6]), 
        .S1(n306), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n312), .A2(n535), .Y(n536) );
  MUX41X1_HVT U74 ( .A1(n537), .A3(n583), .A2(n536), .A4(n585), .S0(n291), 
        .S1(n276), .Y(n534) );
  MUX41X1_HVT U75 ( .A1(n372), .A3(n377), .A2(n390), .A4(n353), .S0(n291), 
        .S1(n276), .Y(n533) );
  MUX41X1_HVT U77 ( .A1(n600), .A3(n379), .A2(n532), .A4(n378), .S0(n297), 
        .S1(in[2]), .Y(n531) );
  MUX41X1_HVT U82 ( .A1(n564), .A3(n351), .A2(n334), .A4(n594), .S0(n289), 
        .S1(n211), .Y(n525) );
  AND2X1_HVT U83 ( .A1(n218), .A2(n256), .Y(n524) );
  MUX41X1_HVT U84 ( .A1(n352), .A3(n602), .A2(n592), .A4(n524), .S0(n291), 
        .S1(n205), .Y(n523) );
  NAND2X0_HVT U85 ( .A1(n326), .A2(n389), .Y(n522) );
  AO21X1_HVT U93 ( .A1(n299), .A2(n514), .A3(n373), .Y(n515) );
  MUX41X1_HVT U97 ( .A1(n372), .A3(n283), .A2(n322), .A4(n593), .S0(n289), 
        .S1(n211), .Y(n510) );
  NAND2X0_HVT U101 ( .A1(n505), .A2(n504), .Y(n506) );
  MUX41X1_HVT U103 ( .A1(n272), .A3(n343), .A2(n255), .A4(n574), .S0(n289), 
        .S1(n211), .Y(n502) );
  MUX41X1_HVT U105 ( .A1(n355), .A3(n562), .A2(n501), .A4(n371), .S0(n289), 
        .S1(n276), .Y(n500) );
  OA21X1_HVT U109 ( .A1(n362), .A2(n234), .A3(n349), .Y(n497) );
  NAND2X0_HVT U110 ( .A1(n317), .A2(n495), .Y(n496) );
  AND2X1_HVT U115 ( .A1(n321), .A2(n204), .Y(n490) );
  NAND2X0_HVT U123 ( .A1(n481), .A2(n480), .Y(n482) );
  MUX41X1_HVT U125 ( .A1(n587), .A3(n288), .A2(n342), .A4(n381), .S0(n289), 
        .S1(n329), .Y(n478) );
  MUX41X1_HVT U131 ( .A1(n473), .A3(n475), .A2(n474), .A4(n476), .S0(n296), 
        .S1(n330), .Y(n472) );
  MUX41X1_HVT U132 ( .A1(n472), .A3(n485), .A2(n477), .A4(n491), .S0(in[6]), 
        .S1(n306), .Y(out[3]) );
  MUX41X1_HVT U135 ( .A1(n382), .A3(n387), .A2(n603), .A4(n582), .S0(n289), 
        .S1(n330), .Y(n469) );
  MUX41X1_HVT U136 ( .A1(n281), .A3(n576), .A2(n383), .A4(n573), .S0(n289), 
        .S1(n330), .Y(n468) );
  MUX41X1_HVT U139 ( .A1(n466), .A3(n469), .A2(n468), .A4(n470), .S0(n307), 
        .S1(n294), .Y(n465) );
  AND2X1_HVT U140 ( .A1(n311), .A2(n325), .Y(n464) );
  MUX41X1_HVT U141 ( .A1(n584), .A3(n363), .A2(n464), .A4(n359), .S0(n291), 
        .S1(n329), .Y(n463) );
  MUX41X1_HVT U142 ( .A1(n352), .A3(n204), .A2(n370), .A4(n311), .S0(n291), 
        .S1(n329), .Y(n462) );
  NAND2X0_HVT U146 ( .A1(n324), .A2(n320), .Y(n535) );
  MUX41X1_HVT U147 ( .A1(n383), .A3(n535), .A2(n372), .A4(n563), .S0(n289), 
        .S1(n330), .Y(n458) );
  MUX41X1_HVT U148 ( .A1(n458), .A3(n462), .A2(n459), .A4(n463), .S0(n308), 
        .S1(n294), .Y(n457) );
  OA21X1_HVT U151 ( .A1(n569), .A2(n331), .A3(n454), .Y(n455) );
  MUX41X1_HVT U153 ( .A1(n496), .A3(n284), .A2(n316), .A4(n336), .S0(n291), 
        .S1(n211), .Y(n452) );
  AND2X1_HVT U154 ( .A1(n299), .A2(n310), .Y(n451) );
  NAND2X0_HVT U158 ( .A1(n323), .A2(n389), .Y(n447) );
  MUX41X1_HVT U159 ( .A1(n596), .A3(n262), .A2(n447), .A4(n341), .S0(in[2]), 
        .S1(n211), .Y(n446) );
  MUX41X1_HVT U160 ( .A1(n446), .A3(n452), .A2(n448), .A4(n453), .S0(n307), 
        .S1(n295), .Y(n445) );
  AND2X1_HVT U162 ( .A1(n602), .A2(n535), .Y(n443) );
  MUX41X1_HVT U163 ( .A1(n348), .A3(n443), .A2(n282), .A4(n444), .S0(n292), 
        .S1(n276), .Y(n442) );
  MUX41X1_HVT U165 ( .A1(n587), .A3(n356), .A2(n563), .A4(n441), .S0(n329), 
        .S1(n293), .Y(n440) );
  NAND2X0_HVT U166 ( .A1(n320), .A2(n552), .Y(n439) );
  NAND2X0_HVT U167 ( .A1(n390), .A2(n326), .Y(n438) );
  MUX41X1_HVT U168 ( .A1(n375), .A3(n311), .A2(n438), .A4(n439), .S0(n327), 
        .S1(n276), .Y(n437) );
  MUX41X1_HVT U172 ( .A1(n434), .A3(n440), .A2(n437), .A4(n442), .S0(n308), 
        .S1(n294), .Y(n433) );
  NAND2X0_HVT U174 ( .A1(n321), .A2(n602), .Y(n595) );
  MUX41X1_HVT U176 ( .A1(n303), .A3(n432), .A2(n380), .A4(n595), .S0(n330), 
        .S1(n327), .Y(n431) );
  NAND2X0_HVT U177 ( .A1(n322), .A2(n304), .Y(n430) );
  MUX41X1_HVT U178 ( .A1(n591), .A3(n430), .A2(n384), .A4(n571), .S0(n291), 
        .S1(n211), .Y(n429) );
  MUX41X1_HVT U179 ( .A1(n581), .A3(n385), .A2(n338), .A4(n384), .S0(n292), 
        .S1(n205), .Y(n428) );
  MUX41X1_HVT U180 ( .A1(n340), .A3(n600), .A2(n596), .A4(n280), .S0(n297), 
        .S1(n291), .Y(n427) );
  OA21X1_HVT U184 ( .A1(n575), .A2(n331), .A3(n352), .Y(n423) );
  MUX41X1_HVT U189 ( .A1(n419), .A3(n595), .A2(n420), .A4(n371), .S0(n297), 
        .S1(n327), .Y(n418) );
  MUX41X1_HVT U190 ( .A1(n418), .A3(n421), .A2(n422), .A4(n425), .S0(n295), 
        .S1(n306), .Y(n417) );
  MUX41X1_HVT U195 ( .A1(n602), .A3(n376), .A2(n319), .A4(n572), .S0(in[2]), 
        .S1(n205), .Y(n413) );
  AO21X1_HVT U197 ( .A1(n285), .A2(n298), .A3(n373), .Y(n411) );
  MUX41X1_HVT U203 ( .A1(n573), .A3(n365), .A2(n597), .A4(n577), .S0(n291), 
        .S1(n211), .Y(n408) );
  MUX41X1_HVT U204 ( .A1(n553), .A3(n596), .A2(n360), .A4(n586), .S0(n243), 
        .S1(n276), .Y(n407) );
  MUX41X1_HVT U206 ( .A1(n406), .A3(n408), .A2(n407), .A4(n259), .S0(n307), 
        .S1(n295), .Y(n405) );
  NAND2X0_HVT U208 ( .A1(n323), .A2(n315), .Y(n495) );
  NAND2X0_HVT U212 ( .A1(n324), .A2(n312), .Y(n552) );
  NAND2X0_HVT U214 ( .A1(n602), .A2(n326), .Y(n404) );
  NAND2X0_HVT U215 ( .A1(n495), .A2(n313), .Y(n403) );
  NAND2X0_HVT U218 ( .A1(n387), .A2(n322), .Y(n454) );
  NAND2X0_HVT U220 ( .A1(n298), .A2(n404), .Y(n527) );
  INVX1_HVT U1 ( .A(n210), .Y(n23) );
  INVX1_HVT U2 ( .A(in[1]), .Y(n210) );
  MUX21X2_HVT U6 ( .A1(n530), .A2(n520), .S0(n48), .Y(out[1]) );
  IBUFFX16_HVT U7 ( .A(in[6]), .Y(n48) );
  INVX0_HVT U8 ( .A(n301), .Y(n203) );
  INVX1_HVT U9 ( .A(n203), .Y(n204) );
  NBUFFX2_HVT U10 ( .A(in[7]), .Y(n205) );
  INVX1_HVT U11 ( .A(in[7]), .Y(n331) );
  MUX21X1_HVT U12 ( .A1(n300), .A2(n301), .S0(n210), .Y(n592) );
  INVX1_HVT U13 ( .A(in[1]), .Y(n325) );
  INVX1_HVT U14 ( .A(n325), .Y(n217) );
  MUX21X1_HVT U16 ( .A1(n486), .A2(n489), .S0(n296), .Y(n485) );
  INVX1_HVT U17 ( .A(n325), .Y(n322) );
  NBUFFX2_HVT U18 ( .A(in[7]), .Y(n211) );
  MUX41X1_HVT U19 ( .A1(n281), .A3(n285), .A2(n522), .A4(n377), .S0(n212), 
        .S1(n213), .Y(n521) );
  IBUFFX16_HVT U20 ( .A(n289), .Y(n212) );
  IBUFFX16_HVT U22 ( .A(n211), .Y(n213) );
  INVX0_HVT U23 ( .A(n325), .Y(n321) );
  INVX1_HVT U25 ( .A(n263), .Y(n327) );
  INVX1_HVT U26 ( .A(n219), .Y(n326) );
  MUX21X1_HVT U27 ( .A1(n547), .A2(n545), .S0(n252), .Y(n544) );
  MUX21X1_HVT U28 ( .A1(n579), .A2(n403), .S0(n297), .Y(n397) );
  MUX21X1_HVT U29 ( .A1(n555), .A2(n559), .S0(n293), .Y(n554) );
  INVX0_HVT U30 ( .A(n571), .Y(n363) );
  MUX21X1_HVT U31 ( .A1(n449), .A2(n450), .S0(n243), .Y(n448) );
  MUX21X1_HVT U32 ( .A1(n357), .A2(n471), .S0(n293), .Y(n470) );
  MUX21X1_HVT U34 ( .A1(n461), .A2(n460), .S0(n293), .Y(n459) );
  INVX1_HVT U36 ( .A(n270), .Y(n271) );
  NAND2X0_HVT U37 ( .A1(n595), .A2(n320), .Y(n596) );
  NAND2X0_HVT U38 ( .A1(n367), .A2(n233), .Y(n264) );
  MUX41X1_HVT U39 ( .A1(n364), .A3(n314), .A2(n366), .A4(n354), .S0(n330), 
        .S1(n289), .Y(n425) );
  MUX21X1_HVT U40 ( .A1(n423), .A2(n424), .S0(n292), .Y(n422) );
  XOR2X1_HVT U41 ( .A1(n582), .A2(n331), .Y(n565) );
  INVX1_HVT U43 ( .A(n290), .Y(n263) );
  INVX0_HVT U44 ( .A(n290), .Y(n234) );
  INVX0_HVT U45 ( .A(n252), .Y(n243) );
  INVX1_HVT U46 ( .A(n308), .Y(n269) );
  INVX1_HVT U47 ( .A(n305), .Y(n256) );
  XOR2X1_HVT U48 ( .A1(n234), .A2(n332), .Y(n216) );
  NAND2X0_HVT U49 ( .A1(n278), .A2(n279), .Y(out[2]) );
  INVX1_HVT U50 ( .A(n277), .Y(n268) );
  INVX1_HVT U52 ( .A(in[6]), .Y(n277) );
  NAND2X0_HVT U54 ( .A1(n231), .A2(n232), .Y(out[6]) );
  INVX0_HVT U55 ( .A(n552), .Y(n372) );
  NBUFFX2_HVT U60 ( .A(n262), .Y(n301) );
  INVX0_HVT U64 ( .A(n602), .Y(n262) );
  INVX1_HVT U65 ( .A(n332), .Y(n329) );
  INVX0_HVT U67 ( .A(n297), .Y(n273) );
  INVX0_HVT U70 ( .A(n297), .Y(n233) );
  NBUFFX2_HVT U71 ( .A(in[1]), .Y(n219) );
  INVX1_HVT U72 ( .A(n325), .Y(n218) );
  INVX1_HVT U76 ( .A(n292), .Y(n252) );
  INVX1_HVT U78 ( .A(n263), .Y(n246) );
  NBUFFX2_HVT U79 ( .A(in[5]), .Y(n294) );
  INVX1_HVT U80 ( .A(in[5]), .Y(n251) );
  AO21X2_HVT U81 ( .A1(n325), .A2(n387), .A3(n331), .Y(n505) );
  INVX1_HVT U86 ( .A(n325), .Y(n324) );
  INVX1_HVT U87 ( .A(n396), .Y(n381) );
  NAND2X0_HVT U88 ( .A1(n426), .A2(n268), .Y(n231) );
  NAND2X0_HVT U89 ( .A1(n417), .A2(n277), .Y(n232) );
  INVX1_HVT U90 ( .A(n588), .Y(n351) );
  INVX1_HVT U91 ( .A(n395), .Y(n382) );
  MUX41X1_HVT U92 ( .A1(n574), .A3(n567), .A2(n416), .A4(n560), .S0(n234), 
        .S1(n205), .Y(n415) );
  MUX41X1_HVT U94 ( .A1(n513), .A3(n518), .A2(n510), .A4(n511), .S0(n294), 
        .S1(n269), .Y(n509) );
  MUX21X2_HVT U95 ( .A1(n379), .A2(n571), .S0(n233), .Y(n449) );
  MUX41X1_HVT U96 ( .A1(n283), .A3(n334), .A2(n512), .A4(n376), .S0(n234), 
        .S1(n205), .Y(n511) );
  MUX41X1_HVT U98 ( .A1(n563), .A3(n567), .A2(n374), .A4(n519), .S0(n291), 
        .S1(n276), .Y(n518) );
  NAND2X0_HVT U99 ( .A1(n313), .A2(n298), .Y(n235) );
  NAND2X0_HVT U100 ( .A1(n588), .A2(n233), .Y(n236) );
  NAND2X0_HVT U102 ( .A1(n235), .A2(n236), .Y(n529) );
  MUX21X1_HVT U104 ( .A1(n436), .A2(n435), .S0(n293), .Y(n434) );
  OA21X1_HVT U106 ( .A1(n286), .A2(n331), .A3(n578), .Y(n435) );
  INVX0_HVT U107 ( .A(n591), .Y(n348) );
  MUX41X1_HVT U108 ( .A1(n429), .A3(n427), .A2(n431), .A4(n428), .S0(n269), 
        .S1(n295), .Y(n426) );
  MUX41X1_HVT U111 ( .A1(n578), .A3(n353), .A2(n490), .A4(n596), .S0(n263), 
        .S1(n273), .Y(n489) );
  NAND2X0_HVT U112 ( .A1(n433), .A2(n277), .Y(n237) );
  NAND2X0_HVT U113 ( .A1(n445), .A2(in[6]), .Y(n238) );
  NAND2X0_HVT U114 ( .A1(n237), .A2(n238), .Y(out[5]) );
  NAND2X0_HVT U116 ( .A1(n594), .A2(n246), .Y(n239) );
  NAND2X0_HVT U117 ( .A1(n358), .A2(n263), .Y(n240) );
  NAND2X0_HVT U118 ( .A1(n239), .A2(n240), .Y(n508) );
  MUX21X1_HVT U119 ( .A1(n284), .A2(n508), .S0(n216), .Y(n507) );
  INVX0_HVT U120 ( .A(n578), .Y(n358) );
  MUX41X1_HVT U121 ( .A1(n271), .A3(n256), .A2(n358), .A4(n385), .S0(n234), 
        .S1(n205), .Y(n406) );
  NAND2X0_HVT U122 ( .A1(n506), .A2(n263), .Y(n241) );
  NAND2X0_HVT U124 ( .A1(n357), .A2(n293), .Y(n242) );
  NAND2X0_HVT U126 ( .A1(n241), .A2(n242), .Y(n503) );
  INVX1_HVT U127 ( .A(n397), .Y(n357) );
  MUX41X1_HVT U128 ( .A1(n582), .A3(n311), .A2(n568), .A4(n382), .S0(n246), 
        .S1(n233), .Y(n414) );
  MUX21X1_HVT U129 ( .A1(n412), .A2(n411), .S0(n292), .Y(n410) );
  MUX21X2_HVT U130 ( .A1(n478), .A2(n479), .S0(n296), .Y(n477) );
  NAND2X0_HVT U133 ( .A1(n539), .A2(n243), .Y(n244) );
  NAND2X0_HVT U134 ( .A1(n565), .A2(n252), .Y(n245) );
  NAND2X0_HVT U137 ( .A1(n244), .A2(n245), .Y(n538) );
  NAND2X0_HVT U138 ( .A1(n496), .A2(n246), .Y(n247) );
  NAND2X0_HVT U143 ( .A1(n578), .A2(n252), .Y(n248) );
  NAND2X0_HVT U144 ( .A1(n247), .A2(n248), .Y(n494) );
  MUX41X1_HVT U145 ( .A1(n570), .A3(n283), .A2(n563), .A4(n535), .S0(n234), 
        .S1(n205), .Y(n421) );
  NAND2X0_HVT U149 ( .A1(n261), .A2(n243), .Y(n249) );
  NAND2X0_HVT U150 ( .A1(n260), .A2(n252), .Y(n250) );
  NAND2X0_HVT U152 ( .A1(n249), .A2(n250), .Y(n259) );
  OA21X2_HVT U155 ( .A1(n601), .A2(n331), .A3(n363), .Y(n260) );
  INVX0_HVT U156 ( .A(n255), .Y(n580) );
  MUX41X1_HVT U157 ( .A1(n494), .A3(n497), .A2(n492), .A4(n498), .S0(n296), 
        .S1(n331), .Y(n491) );
  IBUFFX2_HVT U161 ( .A(n331), .Y(n276) );
  MUX41X1_HVT U164 ( .A1(n538), .A3(n533), .A2(n534), .A4(n531), .S0(n269), 
        .S1(n251), .Y(n530) );
  MUX21X1_HVT U169 ( .A1(n390), .A2(n389), .S0(n324), .Y(n582) );
  NAND2X0_HVT U170 ( .A1(n549), .A2(n252), .Y(n253) );
  NAND2X0_HVT U171 ( .A1(n551), .A2(n292), .Y(n254) );
  NAND2X0_HVT U173 ( .A1(n253), .A2(n254), .Y(n548) );
  OA21X1_HVT U175 ( .A1(n337), .A2(n331), .A3(n578), .Y(n460) );
  IBUFFX2_HVT U181 ( .A(n598), .Y(n344) );
  MUX21X2_HVT U182 ( .A1(n482), .A2(n483), .S0(n273), .Y(n479) );
  MUX21X1_HVT U183 ( .A1(n256), .A2(n314), .S0(n217), .Y(n255) );
  NAND2X0_HVT U185 ( .A1(n528), .A2(n246), .Y(n257) );
  NAND2X0_HVT U186 ( .A1(n529), .A2(n252), .Y(n258) );
  NAND2X0_HVT U187 ( .A1(n257), .A2(n258), .Y(n526) );
  AND3X2_HVT U188 ( .A1(n317), .A2(n552), .A3(n527), .Y(n528) );
  NAND2X0_HVT U191 ( .A1(n275), .A2(n274), .Y(n261) );
  XNOR2X1_HVT U192 ( .A1(n262), .A2(n217), .Y(n563) );
  MUX21X2_HVT U193 ( .A1(n270), .A2(n580), .S0(n273), .Y(n461) );
  MUX21X2_HVT U194 ( .A1(n335), .A2(n484), .S0(n290), .Y(n483) );
  MUX41X1_HVT U196 ( .A1(n410), .A3(n413), .A2(n414), .A4(n415), .S0(n295), 
        .S1(n308), .Y(n409) );
  NAND2X0_HVT U198 ( .A1(n384), .A2(n298), .Y(n265) );
  NAND2X0_HVT U199 ( .A1(n264), .A2(n265), .Y(n412) );
  NAND2X0_HVT U200 ( .A1(n405), .A2(n277), .Y(n266) );
  NAND2X0_HVT U201 ( .A1(n409), .A2(n268), .Y(n267) );
  NAND2X0_HVT U202 ( .A1(n266), .A2(n267), .Y(out[7]) );
  NBUFFX16_HVT U205 ( .A(n328), .Y(n295) );
  MUX41X1_HVT U207 ( .A1(n507), .A3(n502), .A2(n503), .A4(n500), .S0(n269), 
        .S1(n251), .Y(n499) );
  INVX1_HVT U209 ( .A(n393), .Y(n384) );
  MUX41X1_HVT U210 ( .A1(n526), .A3(n523), .A2(n525), .A4(n521), .S0(n269), 
        .S1(n251), .Y(n520) );
  INVX1_HVT U211 ( .A(n606), .Y(n270) );
  INVX1_HVT U213 ( .A(n270), .Y(n272) );
  NAND2X0_HVT U216 ( .A1(n592), .A2(n273), .Y(n274) );
  NAND2X0_HVT U217 ( .A1(n280), .A2(n297), .Y(n275) );
  INVX1_HVT U219 ( .A(n400), .Y(n376) );
  INVX0_HVT U221 ( .A(in[7]), .Y(n332) );
  IBUFFX2_HVT U222 ( .A(n325), .Y(n323) );
  AND3X2_HVT U223 ( .A1(n293), .A2(n326), .A3(n256), .Y(n475) );
  AO21X2_HVT U224 ( .A1(n327), .A2(n311), .A3(n602), .Y(n487) );
  XOR2X2_HVT U225 ( .A1(n303), .A2(n309), .Y(n602) );
  MUX21X2_HVT U226 ( .A1(n457), .A2(n465), .S0(in[6]), .Y(out[4]) );
  NAND2X0_HVT U227 ( .A1(n509), .A2(n268), .Y(n278) );
  NAND2X0_HVT U228 ( .A1(n499), .A2(n277), .Y(n279) );
  MUX21X1_HVT U229 ( .A1(n493), .A2(n318), .S0(n561), .Y(n492) );
  INVX0_HVT U230 ( .A(n309), .Y(n388) );
  INVX1_HVT U231 ( .A(n314), .Y(n386) );
  MUX21X1_HVT U232 ( .A1(n282), .A2(n347), .S0(n291), .Y(n474) );
  NBUFFX2_HVT U233 ( .A(n262), .Y(n302) );
  AND2X1_HVT U234 ( .A1(n302), .A2(n552), .Y(n280) );
  NBUFFX2_HVT U235 ( .A(n604), .Y(n314) );
  INVX1_HVT U236 ( .A(n316), .Y(n390) );
  MUX21X1_HVT U237 ( .A1(n386), .A2(n389), .S0(n296), .Y(n556) );
  NBUFFX2_HVT U238 ( .A(n604), .Y(n315) );
  MUX21X1_HVT U239 ( .A1(n343), .A2(n387), .S0(n296), .Y(n541) );
  AND2X1_HVT U240 ( .A1(n317), .A2(n535), .Y(n281) );
  MUX21X1_HVT U241 ( .A1(n302), .A2(n389), .S0(n323), .Y(n601) );
  MUX21X1_HVT U242 ( .A1(n317), .A2(n301), .S0(n324), .Y(n568) );
  MUX21X1_HVT U243 ( .A1(n262), .A2(n305), .S0(n217), .Y(n504) );
  MUX21X1_HVT U244 ( .A1(n467), .A2(n605), .S0(n243), .Y(n466) );
  MUX21X1_HVT U245 ( .A1(n586), .A2(n364), .S0(n298), .Y(n467) );
  MUX21X1_HVT U246 ( .A1(n386), .A2(n390), .S0(n321), .Y(n432) );
  MUX21X1_HVT U247 ( .A1(n389), .A2(n301), .S0(n324), .Y(n444) );
  MUX21X1_HVT U248 ( .A1(n301), .A2(n386), .S0(n217), .Y(n512) );
  MUX21X1_HVT U249 ( .A1(n315), .A2(n602), .S0(n322), .Y(n572) );
  MUX21X1_HVT U250 ( .A1(n602), .A2(n387), .S0(n322), .Y(n395) );
  MUX21X1_HVT U251 ( .A1(n602), .A2(n390), .S0(n321), .Y(n584) );
  MUX21X1_HVT U252 ( .A1(n315), .A2(n313), .S0(n323), .Y(n519) );
  MUX21X1_HVT U253 ( .A1(n602), .A2(n305), .S0(n217), .Y(n532) );
  MUX21X1_HVT U254 ( .A1(n300), .A2(n602), .S0(n322), .Y(n398) );
  MUX21X1_HVT U255 ( .A1(n389), .A2(n386), .S0(n217), .Y(n571) );
  MUX21X1_HVT U256 ( .A1(n389), .A2(n300), .S0(n217), .Y(n575) );
  MUX21X1_HVT U257 ( .A1(n300), .A2(n390), .S0(n219), .Y(n569) );
  MUX21X1_HVT U258 ( .A1(n381), .A2(n313), .S0(n298), .Y(n471) );
  MUX21X1_HVT U259 ( .A1(n487), .A2(n488), .S0(n298), .Y(n486) );
  MUX21X1_HVT U260 ( .A1(n336), .A2(n360), .S0(n290), .Y(n488) );
  NAND2X0_HVT U261 ( .A1(n303), .A2(n388), .Y(n604) );
  MUX21X1_HVT U262 ( .A1(n386), .A2(n304), .S0(n218), .Y(n396) );
  NBUFFX2_HVT U263 ( .A(n607), .Y(n316) );
  INVX1_HVT U264 ( .A(n311), .Y(n387) );
  INVX1_HVT U265 ( .A(n319), .Y(n389) );
  MUX21X1_HVT U266 ( .A1(n318), .A2(n312), .S0(n323), .Y(n594) );
  MUX21X1_HVT U267 ( .A1(n314), .A2(n320), .S0(n323), .Y(n514) );
  MUX21X1_HVT U268 ( .A1(n387), .A2(n386), .S0(n324), .Y(n590) );
  MUX21X1_HVT U269 ( .A1(n304), .A2(n300), .S0(n218), .Y(n484) );
  NBUFFX2_HVT U270 ( .A(n607), .Y(n317) );
  NBUFFX2_HVT U271 ( .A(n607), .Y(n318) );
  XOR2X1_HVT U272 ( .A1(n322), .A2(n387), .Y(n564) );
  MUX21X1_HVT U273 ( .A1(n300), .A2(n320), .S0(n23), .Y(n419) );
  MUX21X1_HVT U274 ( .A1(n319), .A2(n317), .S0(n321), .Y(n420) );
  MUX21X1_HVT U275 ( .A1(n300), .A2(n389), .S0(n218), .Y(n598) );
  MUX21X1_HVT U276 ( .A1(n315), .A2(n300), .S0(n322), .Y(n597) );
  MUX21X1_HVT U277 ( .A1(n300), .A2(n305), .S0(n321), .Y(n416) );
  XOR2X1_HVT U278 ( .A1(n316), .A2(n324), .Y(n560) );
  MUX21X1_HVT U279 ( .A1(n316), .A2(n304), .S0(n321), .Y(n402) );
  XNOR2X1_HVT U280 ( .A1(n314), .A2(n323), .Y(n282) );
  AND2X1_HVT U281 ( .A1(n323), .A2(n390), .Y(n283) );
  MUX21X1_HVT U282 ( .A1(n319), .A2(n312), .S0(n218), .Y(n578) );
  MUX21X1_HVT U283 ( .A1(n316), .A2(n315), .S0(n217), .Y(n394) );
  AND2X1_HVT U284 ( .A1(n320), .A2(n495), .Y(n284) );
  XNOR2X1_HVT U285 ( .A1(n319), .A2(n322), .Y(n285) );
  MUX21X1_HVT U286 ( .A1(n312), .A2(n300), .S0(n324), .Y(n400) );
  MUX21X1_HVT U287 ( .A1(n313), .A2(n304), .S0(n23), .Y(n537) );
  MUX21X1_HVT U288 ( .A1(n313), .A2(n320), .S0(n293), .Y(n481) );
  XOR2X1_HVT U289 ( .A1(n303), .A2(n323), .Y(n583) );
  NBUFFX2_HVT U290 ( .A(n329), .Y(n299) );
  NBUFFX2_HVT U291 ( .A(n329), .Y(n297) );
  NBUFFX2_HVT U292 ( .A(n329), .Y(n298) );
  NBUFFX2_HVT U293 ( .A(n388), .Y(n300) );
  NBUFFX2_HVT U294 ( .A(in[2]), .Y(n290) );
  NBUFFX2_HVT U295 ( .A(n328), .Y(n296) );
  NBUFFX2_HVT U296 ( .A(in[2]), .Y(n291) );
  NBUFFX2_HVT U297 ( .A(n327), .Y(n293) );
  NBUFFX2_HVT U298 ( .A(n327), .Y(n292) );
  NBUFFX2_HVT U299 ( .A(in[2]), .Y(n289) );
  MUX21X1_HVT U300 ( .A1(n302), .A2(n310), .S0(n218), .Y(n586) );
  NBUFFX2_HVT U301 ( .A(n391), .Y(n303) );
  MUX21X1_HVT U302 ( .A1(n522), .A2(n310), .S0(n298), .Y(n424) );
  XOR2X1_HVT U303 ( .A1(n218), .A2(n309), .Y(n562) );
  MUX21X1_HVT U304 ( .A1(n312), .A2(n302), .S0(n322), .Y(n501) );
  MUX21X1_HVT U305 ( .A1(n455), .A2(n456), .S0(n246), .Y(n453) );
  MUX21X1_HVT U306 ( .A1(n378), .A2(n387), .S0(n298), .Y(n456) );
  MUX21X1_HVT U307 ( .A1(n313), .A2(n376), .S0(n299), .Y(n436) );
  MUX21X1_HVT U308 ( .A1(n387), .A2(n390), .S0(n217), .Y(n441) );
  AND2X1_HVT U309 ( .A1(n302), .A2(n326), .Y(n286) );
  MUX21X1_HVT U310 ( .A1(n310), .A2(n386), .S0(n321), .Y(n570) );
  MUX21X1_HVT U311 ( .A1(n389), .A2(n376), .S0(n299), .Y(n539) );
  MUX21X1_HVT U312 ( .A1(n451), .A2(n318), .S0(n287), .Y(n450) );
  MUX21X1_HVT U313 ( .A1(n591), .A2(n359), .S0(n291), .Y(n473) );
  NAND2X0_HVT U314 ( .A1(n309), .A2(n305), .Y(n607) );
  NBUFFX2_HVT U315 ( .A(n391), .Y(n305) );
  NBUFFX2_HVT U316 ( .A(n608), .Y(n319) );
  NBUFFX2_HVT U317 ( .A(n599), .Y(n311) );
  MUX21X1_HVT U318 ( .A1(n390), .A2(n310), .S0(n218), .Y(n589) );
  MUX21X1_HVT U319 ( .A1(n361), .A2(n271), .S0(n290), .Y(n498) );
  MUX21X1_HVT U320 ( .A1(n557), .A2(n558), .S0(n297), .Y(n555) );
  MUX21X1_HVT U321 ( .A1(n310), .A2(n574), .S0(n296), .Y(n558) );
  XOR2X1_HVT U322 ( .A1(n324), .A2(n295), .Y(n566) );
  MUX21X1_HVT U323 ( .A1(n272), .A2(n325), .S0(n292), .Y(n480) );
  MUX21X1_HVT U324 ( .A1(n310), .A2(n387), .S0(n321), .Y(n399) );
  MUX21X1_HVT U325 ( .A1(n315), .A2(n310), .S0(n322), .Y(n600) );
  MUX21X1_HVT U326 ( .A1(n345), .A2(n326), .S0(n296), .Y(n543) );
  NBUFFX2_HVT U327 ( .A(n599), .Y(n312) );
  MUX21X1_HVT U328 ( .A1(n355), .A2(n579), .S0(n289), .Y(n476) );
  MUX21X1_HVT U329 ( .A1(n318), .A2(n517), .S0(n287), .Y(n516) );
  MUX21X1_HVT U330 ( .A1(n310), .A2(n304), .S0(n299), .Y(n517) );
  NBUFFX2_HVT U331 ( .A(n599), .Y(n313) );
  NBUFFX2_HVT U332 ( .A(n608), .Y(n320) );
  NBUFFX2_HVT U333 ( .A(n391), .Y(n304) );
  XNOR2X1_HVT U334 ( .A1(n331), .A2(n324), .Y(n287) );
  INVX1_HVT U335 ( .A(n332), .Y(n330) );
  AND2X1_HVT U336 ( .A1(n300), .A2(n326), .Y(n288) );
  NBUFFX2_HVT U337 ( .A(in[5]), .Y(n328) );
  INVX0_HVT U338 ( .A(in[4]), .Y(n391) );
  MUX21X1_HVT U339 ( .A1(n515), .A2(n516), .S0(n292), .Y(n513) );
  MUX21X1_HVT U340 ( .A1(n386), .A2(n256), .S0(n323), .Y(n577) );
  NAND2X0_HVT U341 ( .A1(in[4]), .A2(n388), .Y(n599) );
  NAND2X0_HVT U342 ( .A1(n309), .A2(in[4]), .Y(n608) );
  MUX21X1_HVT U343 ( .A1(n256), .A2(n602), .S0(n219), .Y(n401) );
  MUX21X1_HVT U344 ( .A1(n256), .A2(n389), .S0(n324), .Y(n573) );
  MUX21X1_HVT U345 ( .A1(n256), .A2(n387), .S0(n217), .Y(n591) );
  MUX21X1_HVT U346 ( .A1(n256), .A2(n318), .S0(n217), .Y(n588) );
  MUX21X1_HVT U347 ( .A1(n256), .A2(n312), .S0(n321), .Y(n393) );
  MUX21X1_HVT U348 ( .A1(n320), .A2(n256), .S0(n323), .Y(n581) );
  XOR2X1_HVT U349 ( .A1(n321), .A2(n327), .Y(n561) );
  MUX21X1_HVT U350 ( .A1(n310), .A2(n256), .S0(n290), .Y(n493) );
  MUX21X1_HVT U351 ( .A1(n256), .A2(n320), .S0(n218), .Y(n392) );
  MUX21X1_HVT U352 ( .A1(n300), .A2(n256), .S0(n218), .Y(n579) );
  NBUFFX2_HVT U353 ( .A(in[3]), .Y(n309) );
  NBUFFX2_HVT U354 ( .A(in[3]), .Y(n310) );
  NBUFFX2_HVT U355 ( .A(in[0]), .Y(n307) );
  NBUFFX2_HVT U356 ( .A(in[0]), .Y(n308) );
  NBUFFX2_HVT U357 ( .A(in[0]), .Y(n306) );
  INVX0_HVT U358 ( .A(n587), .Y(n333) );
  INVX0_HVT U359 ( .A(n585), .Y(n334) );
  INVX0_HVT U360 ( .A(n576), .Y(n335) );
  INVX0_HVT U361 ( .A(n574), .Y(n336) );
  INVX0_HVT U362 ( .A(n438), .Y(n337) );
  INVX0_HVT U363 ( .A(n404), .Y(n338) );
  INVX0_HVT U364 ( .A(n593), .Y(n339) );
  INVX0_HVT U365 ( .A(n605), .Y(n340) );
  INVX0_HVT U366 ( .A(n603), .Y(n341) );
  INVX0_HVT U367 ( .A(n601), .Y(n342) );
  INVX0_HVT U368 ( .A(n600), .Y(n343) );
  INVX0_HVT U369 ( .A(n597), .Y(n345) );
  INVX0_HVT U370 ( .A(n594), .Y(n346) );
  INVX0_HVT U371 ( .A(n592), .Y(n347) );
  INVX0_HVT U372 ( .A(n590), .Y(n349) );
  INVX0_HVT U373 ( .A(n589), .Y(n350) );
  INVX0_HVT U374 ( .A(n586), .Y(n352) );
  INVX0_HVT U375 ( .A(n584), .Y(n353) );
  INVX0_HVT U376 ( .A(n583), .Y(n354) );
  INVX0_HVT U377 ( .A(n581), .Y(n355) );
  INVX0_HVT U378 ( .A(n579), .Y(n356) );
  INVX0_HVT U379 ( .A(n577), .Y(n359) );
  INVX0_HVT U380 ( .A(n575), .Y(n360) );
  INVX0_HVT U381 ( .A(n573), .Y(n361) );
  INVX0_HVT U382 ( .A(n572), .Y(n362) );
  INVX0_HVT U383 ( .A(n570), .Y(n364) );
  INVX0_HVT U384 ( .A(n569), .Y(n365) );
  INVX0_HVT U385 ( .A(n568), .Y(n366) );
  INVX0_HVT U386 ( .A(n567), .Y(n367) );
  INVX0_HVT U387 ( .A(n535), .Y(n368) );
  INVX0_HVT U388 ( .A(n596), .Y(n369) );
  INVX0_HVT U389 ( .A(n495), .Y(n370) );
  INVX0_HVT U390 ( .A(n403), .Y(n371) );
  INVX0_HVT U391 ( .A(n454), .Y(n373) );
  INVX0_HVT U392 ( .A(n402), .Y(n374) );
  INVX0_HVT U393 ( .A(n401), .Y(n375) );
  INVX0_HVT U394 ( .A(n399), .Y(n377) );
  INVX0_HVT U395 ( .A(n398), .Y(n378) );
  INVX0_HVT U396 ( .A(n514), .Y(n379) );
  INVX0_HVT U397 ( .A(n504), .Y(n380) );
  INVX0_HVT U398 ( .A(n394), .Y(n383) );
  INVX0_HVT U399 ( .A(n392), .Y(n385) );
endmodule

