
module inv_Mix_Column ( in, out1 );
  input [127:0] in;
  output [127:0] out1;
  wire   n50, n51, n53, n54, n55, n57, n58, n59, n60, n61, n63, n64, n65, n66,
         n67, n68, n69, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n116, n117, n118, n119, n120, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n143, n144, n145,
         n146, n147, n148, n149, n150, n152, n154, n155, n157, n158, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n190, n191, n193, n194, n195,
         n198, n199, n200, n201, n202, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n217, n218, n219, n220, n221,
         n222, n224, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n240, n241, n242, n244, n245, n246, n248, n250,
         n251, n252, n253, n254, n255, n256, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n272, n273, n274,
         n275, n276, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n316, n317, n318, n319, n320, n321,
         n324, n325, n326, n327, n328, n330, n331, n332, n333, n334, n335,
         n336, n338, n339, n341, n342, n343, n344, n346, n348, n349, n350,
         n351, n354, n355, n356, n357, n358, n359, n360, n361, n362, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n386, n387, n388,
         n390, n391, n393, n394, n395, n397, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n422, n423, n424, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n486,
         n487, n488, n489, n490, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n509, n510, n511,
         n512, n513, n514, n515, n516, n518, n519, n520, n521, n523, n524,
         n525, n526, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n555, n557, n558, n559, n560, n561,
         n562, n563, n564, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n591, n592, n593, n594, n596, n597,
         n599, n600, n601, n602, n604, n605, n606, n608, n609, n610, n613,
         n614, n615, n617, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n52, n56, n62, n70, n73,
         n92, n115, n121, n142, n151, n153, n156, n159, n189, n192, n196, n197,
         n203, n216, n223, n225, n226, n239, n243, n247, n249, n257, n271,
         n277, n298, n315, n322, n323, n329, n337, n340, n345, n347, n352,
         n353, n363, n373, n385, n389, n392, n396, n398, n421, n425, n442,
         n454, n466, n485, n491, n507, n508, n517, n522, n527, n553, n554,
         n556, n565, n590, n595, n598, n603, n607, n611, n612, n616, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379;

  XNOR3X1_HVT U515 ( .A1(n106), .A2(n107), .A3(n108), .Y(out1[90]) );
  XNOR3X1_HVT U522 ( .A1(n125), .A2(n126), .A3(n127), .Y(out1[87]) );
  XNOR3X1_HVT U552 ( .A1(n211), .A2(n177), .A3(n212), .Y(out1[72]) );
  XNOR3X1_HVT U554 ( .A1(n183), .A2(n213), .A3(n214), .Y(out1[71]) );
  XNOR3X1_HVT U572 ( .A1(n231), .A2(n128), .A3(n212), .Y(out1[64]) );
  XNOR3X1_HVT U576 ( .A1(n1337), .A2(n235), .A3(n236), .Y(n234) );
  XNOR3X1_HVT U586 ( .A1(n266), .A2(n267), .A3(n791), .Y(out1[58]) );
  XNOR3X1_HVT U592 ( .A1(n281), .A2(n282), .A3(n283), .Y(out1[55]) );
  XNOR3X1_HVT U621 ( .A1(n371), .A2(n342), .A3(n372), .Y(out1[40]) );
  XNOR3X1_HVT U625 ( .A1(n343), .A2(n379), .A3(n380), .Y(out1[39]) );
  XNOR3X1_HVT U657 ( .A1(n436), .A2(n437), .A3(n438), .Y(out1[24]) );
  XNOR3X1_HVT U674 ( .A1(n481), .A2(n181), .A3(n438), .Y(out1[16]) );
  XNOR3X1_HVT U698 ( .A1(n532), .A2(n533), .A3(n534), .Y(out1[120]) );
  XNOR3X1_HVT U702 ( .A1(n537), .A2(n538), .A3(n539), .Y(out1[119]) );
  XNOR3X1_HVT U713 ( .A1(n578), .A2(n579), .A3(n529), .Y(out1[113]) );
  XNOR3X1_HVT U715 ( .A1(n584), .A2(n585), .A3(n534), .Y(out1[112]) );
  XNOR3X1_HVT U735 ( .A1(n497), .A2(n586), .A3(n609), .Y(out1[104]) );
  XNOR3X1_HVT U743 ( .A1(n482), .A2(n440), .A3(n617), .Y(out1[0]) );
  INVX1_HVT U1 ( .A(n143), .Y(n1019) );
  INVX0_HVT U2 ( .A(in[77]), .Y(n1034) );
  NBUFFX2_HVT U3 ( .A(n606), .Y(n1) );
  INVX0_HVT U4 ( .A(n479), .Y(n726) );
  INVX2_HVT U5 ( .A(n1113), .Y(n1130) );
  XOR3X2_HVT U6 ( .A1(n763), .A2(n764), .A3(n64), .Y(n1226) );
  IBUFFX2_HVT U7 ( .A(in[105]), .Y(n1372) );
  INVX1_HVT U8 ( .A(in[79]), .Y(n1363) );
  INVX1_HVT U9 ( .A(n261), .Y(n1037) );
  INVX0_HVT U10 ( .A(in[15]), .Y(n833) );
  XNOR2X2_HVT U11 ( .A1(n975), .A2(n115), .Y(n525) );
  XNOR2X2_HVT U12 ( .A1(n525), .A2(n574), .Y(n528) );
  INVX2_HVT U13 ( .A(n1281), .Y(n430) );
  INVX0_HVT U14 ( .A(n336), .Y(n852) );
  XOR3X2_HVT U15 ( .A1(n1219), .A2(n307), .A3(n2), .Y(out1[35]) );
  INVX1_HVT U16 ( .A(n423), .Y(n329) );
  INVX0_HVT U17 ( .A(in[126]), .Y(n92) );
  NAND2X0_HVT U18 ( .A1(n11), .A2(n12), .Y(n2) );
  INVX1_HVT U19 ( .A(in[71]), .Y(n1361) );
  NAND2X0_HVT U20 ( .A1(n902), .A2(n431), .Y(n5) );
  NAND2X0_HVT U21 ( .A1(n3), .A2(n4), .Y(n6) );
  NAND2X0_HVT U22 ( .A1(n5), .A2(n6), .Y(out1[25]) );
  INVX0_HVT U23 ( .A(n902), .Y(n3) );
  IBUFFX2_HVT U24 ( .A(n431), .Y(n4) );
  INVX0_HVT U25 ( .A(n671), .Y(n7) );
  XNOR2X2_HVT U26 ( .A1(n269), .A2(n366), .Y(n276) );
  INVX2_HVT U27 ( .A(n1199), .Y(n1192) );
  IBUFFX2_HVT U28 ( .A(n155), .Y(n1065) );
  IBUFFX2_HVT U29 ( .A(n1363), .Y(n28) );
  INVX1_HVT U30 ( .A(n217), .Y(n565) );
  XOR3X1_HVT U31 ( .A1(n1208), .A2(n1106), .A3(n325), .Y(n490) );
  IBUFFX2_HVT U32 ( .A(n200), .Y(n42) );
  IBUFFX2_HVT U33 ( .A(n1163), .Y(n169) );
  NAND2X0_HVT U34 ( .A1(n778), .A2(n779), .Y(n8) );
  INVX0_HVT U35 ( .A(in[47]), .Y(n1209) );
  XNOR2X1_HVT U36 ( .A1(in[57]), .A2(in[62]), .Y(n361) );
  NAND2X0_HVT U37 ( .A1(n1185), .A2(n261), .Y(n11) );
  NAND2X0_HVT U38 ( .A1(n9), .A2(n10), .Y(n12) );
  NAND2X0_HVT U39 ( .A1(n11), .A2(n12), .Y(n358) );
  INVX0_HVT U40 ( .A(n1185), .Y(n9) );
  INVX0_HVT U41 ( .A(n261), .Y(n10) );
  XOR3X2_HVT U42 ( .A1(n13), .A2(n495), .A3(n496), .Y(out1[127]) );
  IBUFFX16_HVT U43 ( .A(n494), .Y(n13) );
  INVX2_HVT U44 ( .A(n1358), .Y(n876) );
  IBUFFX2_HVT U45 ( .A(n202), .Y(n14) );
  INVX1_HVT U46 ( .A(n14), .Y(n15) );
  INVX1_HVT U47 ( .A(n676), .Y(n271) );
  XNOR2X1_HVT U48 ( .A1(n837), .A2(n336), .Y(n690) );
  IBUFFX2_HVT U49 ( .A(n824), .Y(n16) );
  INVX1_HVT U50 ( .A(n16), .Y(n17) );
  XOR3X1_HVT U51 ( .A1(n555), .A2(n548), .A3(n512), .Y(n1321) );
  IBUFFX2_HVT U52 ( .A(n228), .Y(n860) );
  INVX0_HVT U53 ( .A(n361), .Y(n18) );
  INVX1_HVT U54 ( .A(n18), .Y(n19) );
  XNOR2X1_HVT U55 ( .A1(n305), .A2(n797), .Y(n383) );
  AND2X1_HVT U56 ( .A1(n31), .A2(n32), .Y(n20) );
  INVX1_HVT U57 ( .A(in[127]), .Y(n1379) );
  XNOR2X2_HVT U58 ( .A1(n41), .A2(n1257), .Y(n725) );
  INVX2_HVT U59 ( .A(n1345), .Y(n1257) );
  INVX2_HVT U60 ( .A(n1263), .Y(n853) );
  INVX0_HVT U61 ( .A(in[125]), .Y(n628) );
  INVX2_HVT U62 ( .A(n1104), .Y(n962) );
  NBUFFX4_HVT U63 ( .A(in[31]), .Y(n1104) );
  XOR3X1_HVT U64 ( .A1(n60), .A2(n59), .A3(n61), .Y(n1279) );
  NAND2X0_HVT U65 ( .A1(in[74]), .A2(n1363), .Y(n23) );
  NAND2X0_HVT U66 ( .A1(n21), .A2(n22), .Y(n24) );
  NAND2X0_HVT U67 ( .A1(n23), .A2(n24), .Y(n155) );
  INVX0_HVT U68 ( .A(in[74]), .Y(n21) );
  INVX0_HVT U69 ( .A(n1363), .Y(n22) );
  XOR3X2_HVT U70 ( .A1(n1241), .A2(n1003), .A3(n552), .Y(n1265) );
  INVX1_HVT U71 ( .A(in[127]), .Y(n1227) );
  INVX1_HVT U72 ( .A(n193), .Y(n1301) );
  INVX0_HVT U73 ( .A(in[43]), .Y(n989) );
  NBUFFX16_HVT U74 ( .A(n659), .Y(n826) );
  IBUFFX2_HVT U75 ( .A(in[6]), .Y(n1342) );
  NBUFFX2_HVT U76 ( .A(in[22]), .Y(n1202) );
  XNOR3X2_HVT U77 ( .A1(n725), .A2(n527), .A3(n425), .Y(n412) );
  INVX0_HVT U78 ( .A(in[106]), .Y(n634) );
  INVX0_HVT U79 ( .A(n208), .Y(n922) );
  XOR3X2_HVT U80 ( .A1(n310), .A2(n25), .A3(n262), .Y(n309) );
  IBUFFX16_HVT U81 ( .A(n311), .Y(n25) );
  INVX2_HVT U82 ( .A(n101), .Y(n1044) );
  INVX0_HVT U83 ( .A(in[102]), .Y(n1297) );
  INVX1_HVT U84 ( .A(in[38]), .Y(n765) );
  XOR3X2_HVT U85 ( .A1(n176), .A2(n1200), .A3(n177), .Y(n26) );
  INVX8_HVT U86 ( .A(n26), .Y(n123) );
  INVX0_HVT U87 ( .A(n1208), .Y(n27) );
  INVX2_HVT U88 ( .A(n1017), .Y(n1018) );
  INVX1_HVT U89 ( .A(in[86]), .Y(n1317) );
  INVX0_HVT U90 ( .A(n300), .Y(n1244) );
  IBUFFX2_HVT U91 ( .A(n248), .Y(n1137) );
  INVX0_HVT U92 ( .A(n64), .Y(n1095) );
  XOR3X2_HVT U93 ( .A1(n28), .A2(n1199), .A3(n80), .Y(n211) );
  INVX1_HVT U94 ( .A(n1258), .Y(n1006) );
  NAND2X0_HVT U95 ( .A1(in[120]), .A2(n1379), .Y(n31) );
  NAND2X0_HVT U96 ( .A1(n29), .A2(n30), .Y(n32) );
  NAND2X0_HVT U97 ( .A1(n31), .A2(n32), .Y(n1206) );
  INVX0_HVT U98 ( .A(in[120]), .Y(n29) );
  INVX0_HVT U99 ( .A(n1379), .Y(n30) );
  INVX0_HVT U100 ( .A(n1206), .Y(n710) );
  XOR3X1_HVT U101 ( .A1(n230), .A2(n165), .A3(n922), .Y(out1[65]) );
  IBUFFX2_HVT U102 ( .A(n334), .Y(n1169) );
  IBUFFX2_HVT U103 ( .A(n374), .Y(n56) );
  IBUFFX2_HVT U104 ( .A(n311), .Y(n1339) );
  XNOR2X2_HVT U105 ( .A1(n633), .A2(n782), .Y(n677) );
  INVX1_HVT U106 ( .A(n1311), .Y(n943) );
  IBUFFX2_HVT U107 ( .A(in[42]), .Y(n1049) );
  XNOR2X2_HVT U108 ( .A1(in[98]), .A2(n937), .Y(n625) );
  XNOR2X2_HVT U109 ( .A1(n1045), .A2(n45), .Y(n221) );
  INVX2_HVT U110 ( .A(n44), .Y(n45) );
  NAND2X0_HVT U111 ( .A1(n38), .A2(n39), .Y(n33) );
  XOR3X2_HVT U112 ( .A1(n34), .A2(n1360), .A3(n176), .Y(n231) );
  IBUFFX16_HVT U113 ( .A(n1369), .Y(n34) );
  NBUFFX2_HVT U114 ( .A(n1134), .Y(n35) );
  NAND2X0_HVT U115 ( .A1(n1261), .A2(n1360), .Y(n38) );
  NAND2X0_HVT U116 ( .A1(n36), .A2(n37), .Y(n39) );
  NAND2X0_HVT U117 ( .A1(n38), .A2(n39), .Y(n205) );
  IBUFFX2_HVT U118 ( .A(n1261), .Y(n36) );
  INVX0_HVT U119 ( .A(n1360), .Y(n37) );
  INVX1_HVT U120 ( .A(n472), .Y(n40) );
  INVX1_HVT U121 ( .A(n40), .Y(n41) );
  XNOR3X1_HVT U122 ( .A1(n499), .A2(n500), .A3(n501), .Y(out1[126]) );
  IBUFFX2_HVT U123 ( .A(n1351), .Y(n950) );
  INVX1_HVT U124 ( .A(in[111]), .Y(n635) );
  INVX0_HVT U125 ( .A(in[111]), .Y(n1258) );
  INVX2_HVT U126 ( .A(n94), .Y(n1213) );
  INVX2_HVT U127 ( .A(in[37]), .Y(n1350) );
  INVX1_HVT U128 ( .A(n42), .Y(n43) );
  INVX1_HVT U129 ( .A(n188), .Y(n44) );
  INVX0_HVT U130 ( .A(in[67]), .Y(n951) );
  XOR3X2_HVT U131 ( .A1(n46), .A2(n528), .A3(n529), .Y(out1[121]) );
  XNOR3X1_HVT U132 ( .A1(n530), .A2(n1221), .A3(n1186), .Y(n46) );
  INVX1_HVT U133 ( .A(n463), .Y(n389) );
  XOR3X2_HVT U134 ( .A1(n1348), .A2(n258), .A3(n259), .Y(n1284) );
  XOR3X2_HVT U135 ( .A1(n1269), .A2(n399), .A3(n259), .Y(n488) );
  XNOR2X1_HVT U136 ( .A1(n348), .A2(n765), .Y(n291) );
  INVX0_HVT U137 ( .A(in[109]), .Y(n1233) );
  XNOR3X2_HVT U138 ( .A1(n74), .A2(n1115), .A3(n586), .Y(n534) );
  NBUFFX2_HVT U139 ( .A(n513), .Y(n47) );
  XNOR2X2_HVT U140 ( .A1(in[58]), .A2(n1014), .Y(n263) );
  XOR3X1_HVT U141 ( .A1(n1190), .A2(n78), .A3(n85), .Y(n84) );
  XOR2X1_HVT U142 ( .A1(in[69]), .A2(in[70]), .Y(n209) );
  INVX0_HVT U143 ( .A(n932), .Y(n48) );
  INVX1_HVT U144 ( .A(in[89]), .Y(n1066) );
  IBUFFX2_HVT U145 ( .A(n288), .Y(n49) );
  INVX1_HVT U146 ( .A(n49), .Y(n52) );
  INVX1_HVT U147 ( .A(in[15]), .Y(n1346) );
  XOR3X2_HVT U148 ( .A1(n1275), .A2(n56), .A3(n62), .Y(out1[3]) );
  IBUFFX16_HVT U149 ( .A(n739), .Y(n62) );
  IBUFFX2_HVT U150 ( .A(n1066), .Y(n932) );
  IBUFFX2_HVT U151 ( .A(n605), .Y(n70) );
  INVX1_HVT U152 ( .A(n70), .Y(n73) );
  INVX1_HVT U153 ( .A(n92), .Y(n115) );
  XOR2X1_HVT U154 ( .A1(in[27]), .A2(n1104), .Y(n326) );
  IBUFFX2_HVT U155 ( .A(n254), .Y(n1157) );
  IBUFFX2_HVT U156 ( .A(n435), .Y(n1138) );
  XOR3X1_HVT U157 ( .A1(n450), .A2(n925), .A3(n1174), .Y(n1323) );
  INVX0_HVT U158 ( .A(in[117]), .Y(n1375) );
  XOR3X2_HVT U159 ( .A1(n366), .A2(n121), .A3(n270), .Y(n762) );
  IBUFFX16_HVT U160 ( .A(n877), .Y(n121) );
  INVX0_HVT U161 ( .A(n137), .Y(n1152) );
  XNOR2X1_HVT U162 ( .A1(in[0]), .A2(n1031), .Y(n112) );
  XNOR2X2_HVT U163 ( .A1(in[108]), .A2(n1373), .Y(n589) );
  INVX1_HVT U164 ( .A(n509), .Y(n992) );
  INVX1_HVT U165 ( .A(in[109]), .Y(n1373) );
  NAND2X0_HVT U166 ( .A1(n851), .A2(n151), .Y(n153) );
  NAND2X0_HVT U167 ( .A1(n142), .A2(n1306), .Y(n156) );
  NAND2X0_HVT U168 ( .A1(n153), .A2(n156), .Y(n275) );
  INVX0_HVT U169 ( .A(n851), .Y(n142) );
  IBUFFX2_HVT U170 ( .A(n1306), .Y(n151) );
  XOR2X2_HVT U171 ( .A1(n275), .A2(n630), .Y(n331) );
  INVX1_HVT U172 ( .A(n1034), .Y(n1035) );
  INVX0_HVT U173 ( .A(n665), .Y(n159) );
  INVX2_HVT U174 ( .A(n731), .Y(n665) );
  INVX1_HVT U175 ( .A(n390), .Y(n731) );
  NAND2X0_HVT U176 ( .A1(in[91]), .A2(n944), .Y(n196) );
  NAND2X0_HVT U177 ( .A1(n189), .A2(n192), .Y(n197) );
  NAND2X0_HVT U178 ( .A1(n196), .A2(n197), .Y(n99) );
  INVX0_HVT U179 ( .A(in[91]), .Y(n189) );
  INVX0_HVT U180 ( .A(n944), .Y(n192) );
  INVX0_HVT U181 ( .A(n99), .Y(n843) );
  IBUFFX2_HVT U182 ( .A(n152), .Y(n1309) );
  XOR2X1_HVT U183 ( .A1(in[64]), .A2(in[69]), .Y(n177) );
  INVX0_HVT U184 ( .A(n253), .Y(n203) );
  INVX1_HVT U185 ( .A(n203), .Y(n216) );
  NBUFFX2_HVT U186 ( .A(n263), .Y(n223) );
  XNOR3X1_HVT U187 ( .A1(n475), .A2(n396), .A3(n427), .Y(out1[18]) );
  INVX1_HVT U188 ( .A(n200), .Y(n823) );
  IBUFFX2_HVT U189 ( .A(n778), .Y(n225) );
  INVX1_HVT U190 ( .A(in[38]), .Y(n1351) );
  NAND2X0_HVT U191 ( .A1(n1246), .A2(in[34]), .Y(n243) );
  NAND2X0_HVT U192 ( .A1(n226), .A2(n239), .Y(n247) );
  NAND2X0_HVT U193 ( .A1(n243), .A2(n247), .Y(n387) );
  INVX0_HVT U194 ( .A(n1246), .Y(n226) );
  INVX0_HVT U195 ( .A(in[34]), .Y(n239) );
  INVX0_HVT U196 ( .A(n387), .Y(n1266) );
  INVX0_HVT U197 ( .A(in[34]), .Y(n249) );
  XNOR2X2_HVT U198 ( .A1(n958), .A2(n1067), .Y(n119) );
  INVX1_HVT U199 ( .A(in[93]), .Y(n958) );
  INVX0_HVT U200 ( .A(n1253), .Y(n1023) );
  INVX1_HVT U201 ( .A(n249), .Y(n257) );
  INVX0_HVT U202 ( .A(n583), .Y(n1242) );
  INVX1_HVT U203 ( .A(n839), .Y(n620) );
  IBUFFX2_HVT U204 ( .A(n383), .Y(n1248) );
  XOR3X2_HVT U205 ( .A1(n800), .A2(n271), .A3(n108), .Y(n161) );
  XNOR2X1_HVT U206 ( .A1(n861), .A2(n171), .Y(n684) );
  XNOR2X2_HVT U207 ( .A1(n385), .A2(n1362), .Y(n206) );
  INVX1_HVT U208 ( .A(n1271), .Y(n277) );
  INVX2_HVT U209 ( .A(in[36]), .Y(n1271) );
  INVX0_HVT U210 ( .A(in[23]), .Y(n1056) );
  INVX0_HVT U211 ( .A(in[63]), .Y(n623) );
  INVX1_HVT U212 ( .A(n1065), .Y(n298) );
  IBUFFX2_HVT U213 ( .A(n103), .Y(n1263) );
  XOR2X2_HVT U214 ( .A1(in[113]), .A2(in[118]), .Y(n570) );
  INVX1_HVT U215 ( .A(in[118]), .Y(n1315) );
  XNOR2X2_HVT U216 ( .A1(n1348), .A2(n695), .Y(n395) );
  INVX2_HVT U217 ( .A(n1129), .Y(n695) );
  XOR3X1_HVT U218 ( .A1(n395), .A2(n1295), .A3(n401), .Y(n1322) );
  INVX1_HVT U219 ( .A(in[39]), .Y(n1352) );
  INVX1_HVT U220 ( .A(n624), .Y(n1109) );
  INVX1_HVT U221 ( .A(n511), .Y(n982) );
  IBUFFX2_HVT U222 ( .A(in[77]), .Y(n1307) );
  IBUFFX2_HVT U223 ( .A(in[59]), .Y(n315) );
  INVX1_HVT U224 ( .A(n315), .Y(n322) );
  XOR3X1_HVT U225 ( .A1(n383), .A2(n779), .A3(n723), .Y(n1324) );
  XNOR2X1_HVT U226 ( .A1(in[37]), .A2(n765), .Y(n369) );
  INVX0_HVT U227 ( .A(n1266), .Y(n323) );
  XOR3X2_HVT U228 ( .A1(n1227), .A2(n1298), .A3(n76), .Y(n1330) );
  NAND2X0_HVT U229 ( .A1(n423), .A2(n1064), .Y(n340) );
  NAND2X0_HVT U230 ( .A1(n329), .A2(n337), .Y(n345) );
  NAND2X0_HVT U231 ( .A1(n340), .A2(n345), .Y(n467) );
  INVX0_HVT U232 ( .A(n1064), .Y(n337) );
  INVX0_HVT U233 ( .A(n467), .Y(n971) );
  NBUFFX2_HVT U234 ( .A(in[72]), .Y(n347) );
  XOR3X2_HVT U235 ( .A1(n840), .A2(n1161), .A3(n325), .Y(n1286) );
  INVX0_HVT U236 ( .A(n548), .Y(n507) );
  INVX1_HVT U237 ( .A(n1065), .Y(n352) );
  XOR3X1_HVT U238 ( .A1(n1082), .A2(n350), .A3(n355), .Y(n1253) );
  XNOR2X2_HVT U239 ( .A1(n252), .A2(n304), .Y(n350) );
  XOR3X1_HVT U240 ( .A1(n738), .A2(n83), .A3(n84), .Y(out1[94]) );
  XOR3X2_HVT U241 ( .A1(n154), .A2(n352), .A3(n102), .Y(n1310) );
  XNOR2X2_HVT U242 ( .A1(in[75]), .A2(n1363), .Y(n148) );
  NAND2X0_HVT U243 ( .A1(n732), .A2(n733), .Y(n353) );
  XNOR2X2_HVT U244 ( .A1(n201), .A2(in[93]), .Y(n93) );
  XNOR3X1_HVT U245 ( .A1(n920), .A2(n428), .A3(n429), .Y(n719) );
  NBUFFX2_HVT U246 ( .A(n326), .Y(n363) );
  NAND2X0_HVT U247 ( .A1(n881), .A2(n882), .Y(n373) );
  NBUFFX2_HVT U248 ( .A(in[79]), .Y(n385) );
  IBUFFX2_HVT U249 ( .A(n97), .Y(n1179) );
  XNOR2X2_HVT U250 ( .A1(n53), .A2(n726), .Y(n933) );
  XOR2X1_HVT U251 ( .A1(in[8]), .A2(in[13]), .Y(n482) );
  XOR3X2_HVT U252 ( .A1(n434), .A2(n389), .A3(n464), .Y(n51) );
  IBUFFX2_HVT U253 ( .A(n476), .Y(n392) );
  INVX1_HVT U254 ( .A(n392), .Y(n396) );
  NBUFFX2_HVT U255 ( .A(n257), .Y(n398) );
  INVX0_HVT U256 ( .A(in[95]), .Y(n595) );
  INVX0_HVT U257 ( .A(in[95]), .Y(n1053) );
  INVX0_HVT U258 ( .A(n331), .Y(n666) );
  IBUFFX2_HVT U259 ( .A(n419), .Y(n421) );
  INVX1_HVT U260 ( .A(n421), .Y(n425) );
  INVX0_HVT U261 ( .A(n450), .Y(n1195) );
  XNOR2X1_HVT U262 ( .A1(n468), .A2(n1267), .Y(n974) );
  INVX0_HVT U263 ( .A(in[18]), .Y(n1090) );
  INVX1_HVT U264 ( .A(n1328), .Y(n809) );
  INVX0_HVT U265 ( .A(n614), .Y(n1092) );
  INVX1_HVT U266 ( .A(n163), .Y(n921) );
  XNOR2X2_HVT U267 ( .A1(n974), .A2(n527), .Y(n450) );
  XNOR2X2_HVT U268 ( .A1(n625), .A2(n1298), .Y(n1134) );
  IBUFFX2_HVT U269 ( .A(in[51]), .Y(n442) );
  INVX1_HVT U270 ( .A(n442), .Y(n454) );
  IBUFFX2_HVT U271 ( .A(n404), .Y(n466) );
  INVX1_HVT U272 ( .A(n466), .Y(n485) );
  NBUFFX2_HVT U273 ( .A(n559), .Y(n491) );
  INVX0_HVT U274 ( .A(in[107]), .Y(n976) );
  INVX2_HVT U275 ( .A(in[39]), .Y(n1246) );
  XOR3X2_HVT U276 ( .A1(n547), .A2(n507), .A3(n549), .Y(out1[117]) );
  INVX1_HVT U277 ( .A(n359), .Y(n703) );
  NBUFFX2_HVT U278 ( .A(n465), .Y(n508) );
  XNOR2X2_HVT U279 ( .A1(n418), .A2(n1267), .Y(n401) );
  XOR3X2_HVT U280 ( .A1(n1373), .A2(n538), .A3(n502), .Y(n544) );
  INVX1_HVT U281 ( .A(in[103]), .Y(n1371) );
  INVX0_HVT U282 ( .A(n328), .Y(n849) );
  NBUFFX2_HVT U283 ( .A(n602), .Y(n517) );
  INVX1_HVT U284 ( .A(n418), .Y(n522) );
  INVX1_HVT U285 ( .A(n522), .Y(n527) );
  XOR3X2_HVT U286 ( .A1(n553), .A2(n554), .A3(n486), .Y(out1[14]) );
  IBUFFX16_HVT U287 ( .A(n1128), .Y(n553) );
  IBUFFX16_HVT U288 ( .A(n484), .Y(n554) );
  XNOR2X1_HVT U289 ( .A1(n97), .A2(n148), .Y(n190) );
  INVX1_HVT U290 ( .A(n726), .Y(n556) );
  XOR3X2_HVT U291 ( .A1(n373), .A2(n565), .A3(n590), .Y(out1[6]) );
  XOR3X2_HVT U292 ( .A1(n1129), .A2(n179), .A3(n915), .Y(n590) );
  IBUFFX2_HVT U293 ( .A(n93), .Y(n911) );
  INVX1_HVT U294 ( .A(n595), .Y(n598) );
  INVX1_HVT U295 ( .A(n413), .Y(n1153) );
  NAND2X0_HVT U296 ( .A1(n968), .A2(n967), .Y(n603) );
  XNOR2X2_HVT U297 ( .A1(n254), .A2(in[44]), .Y(n238) );
  XNOR3X2_HVT U298 ( .A1(n545), .A2(n1060), .A3(n550), .Y(n1314) );
  XOR3X2_HVT U299 ( .A1(n566), .A2(n607), .A3(n58), .Y(n1197) );
  IBUFFX16_HVT U300 ( .A(n633), .Y(n607) );
  XNOR2X1_HVT U301 ( .A1(n829), .A2(n851), .Y(n339) );
  IBUFFX2_HVT U302 ( .A(in[19]), .Y(n611) );
  INVX1_HVT U303 ( .A(n611), .Y(n612) );
  INVX2_HVT U304 ( .A(n1311), .Y(n1312) );
  XOR3X2_HVT U305 ( .A1(n61), .A2(n1091), .A3(n935), .Y(n519) );
  INVX0_HVT U306 ( .A(n274), .Y(n658) );
  XNOR2X2_HVT U307 ( .A1(n515), .A2(n616), .Y(n504) );
  IBUFFX16_HVT U308 ( .A(n645), .Y(n616) );
  AND2X1_HVT U309 ( .A1(n964), .A2(n963), .Y(n618) );
  INVX1_HVT U310 ( .A(n238), .Y(n1182) );
  XNOR2X2_HVT U311 ( .A1(in[59]), .A2(n624), .Y(n254) );
  NAND2X0_HVT U312 ( .A1(n839), .A2(n604), .Y(n621) );
  NAND2X0_HVT U313 ( .A1(n619), .A2(n620), .Y(n622) );
  NAND2X0_HVT U314 ( .A1(n622), .A2(n621), .Y(n560) );
  INVX1_HVT U315 ( .A(n604), .Y(n619) );
  IBUFFX2_HVT U316 ( .A(n1297), .Y(n839) );
  IBUFFX2_HVT U317 ( .A(n1315), .Y(n734) );
  XOR2X2_HVT U318 ( .A1(in[36]), .A2(n939), .Y(n286) );
  INVX1_HVT U319 ( .A(n623), .Y(n624) );
  XNOR2X1_HVT U320 ( .A1(n577), .A2(n576), .Y(n66) );
  XOR2X1_HVT U321 ( .A1(n478), .A2(n403), .Y(n460) );
  INVX0_HVT U322 ( .A(n145), .Y(n863) );
  INVX1_HVT U323 ( .A(n801), .Y(n676) );
  IBUFFX2_HVT U324 ( .A(in[73]), .Y(n801) );
  IBUFFX2_HVT U325 ( .A(in[113]), .Y(n626) );
  INVX1_HVT U326 ( .A(n626), .Y(n627) );
  XOR2X1_HVT U327 ( .A1(n19), .A2(n1075), .Y(n265) );
  IBUFFX2_HVT U328 ( .A(n1363), .Y(n798) );
  INVX1_HVT U329 ( .A(in[103]), .Y(n937) );
  XOR3X2_HVT U330 ( .A1(n1279), .A2(n1277), .A3(n1278), .Y(out1[99]) );
  INVX1_HVT U331 ( .A(n93), .Y(n898) );
  INVX1_HVT U332 ( .A(in[94]), .Y(n1329) );
  INVX1_HVT U333 ( .A(n628), .Y(n629) );
  XOR3X2_HVT U334 ( .A1(n170), .A2(n171), .A3(n172), .Y(n117) );
  IBUFFX2_HVT U335 ( .A(in[2]), .Y(n1126) );
  INVX0_HVT U336 ( .A(n1207), .Y(n630) );
  IBUFFX2_HVT U337 ( .A(n1281), .Y(n1062) );
  XNOR2X2_HVT U338 ( .A1(n525), .A2(in[122]), .Y(n572) );
  INVX2_HVT U339 ( .A(n1205), .Y(n945) );
  INVX2_HVT U340 ( .A(in[30]), .Y(n1349) );
  INVX0_HVT U341 ( .A(n335), .Y(n631) );
  INVX0_HVT U342 ( .A(n631), .Y(n632) );
  IBUFFX2_HVT U343 ( .A(n510), .Y(n1268) );
  IBUFFX2_HVT U344 ( .A(in[27]), .Y(n1064) );
  XNOR3X2_HVT U345 ( .A1(n363), .A2(n974), .A3(n256), .Y(n321) );
  INVX2_HVT U346 ( .A(n692), .Y(n555) );
  XOR3X2_HVT U347 ( .A1(n1137), .A2(n745), .A3(n793), .Y(n1251) );
  XOR3X2_HVT U348 ( .A1(n596), .A2(n1220), .A3(n601), .Y(n599) );
  INVX2_HVT U349 ( .A(n945), .Y(n875) );
  INVX1_HVT U350 ( .A(n302), .Y(n778) );
  XNOR2X1_HVT U351 ( .A1(n369), .A2(in[33]), .Y(n689) );
  AND2X1_HVT U352 ( .A1(n636), .A2(n637), .Y(n633) );
  NAND2X0_HVT U353 ( .A1(in[106]), .A2(n635), .Y(n636) );
  NAND2X0_HVT U354 ( .A1(n634), .A2(n1006), .Y(n637) );
  NAND2X0_HVT U355 ( .A1(n636), .A2(n637), .Y(n563) );
  XOR2X2_HVT U356 ( .A1(n365), .A2(n398), .Y(n320) );
  INVX1_HVT U357 ( .A(n1077), .Y(n638) );
  INVX2_HVT U358 ( .A(n638), .Y(n639) );
  INVX0_HVT U359 ( .A(in[46]), .Y(n1077) );
  INVX2_HVT U360 ( .A(n954), .Y(n1041) );
  INVX2_HVT U361 ( .A(n301), .Y(n779) );
  IBUFFX2_HVT U362 ( .A(n354), .Y(n1081) );
  XOR3X1_HVT U363 ( .A1(n1334), .A2(n798), .A3(n123), .Y(n175) );
  XOR2X2_HVT U364 ( .A1(n1080), .A2(n1358), .Y(n280) );
  INVX1_HVT U365 ( .A(n1358), .Y(n851) );
  XNOR3X1_HVT U366 ( .A1(n1346), .A2(n1345), .A3(n114), .Y(n111) );
  XNOR2X2_HVT U367 ( .A1(n1348), .A2(n859), .Y(n443) );
  XOR3X1_HVT U368 ( .A1(n761), .A2(n1372), .A3(n66), .Y(n571) );
  XOR3X2_HVT U369 ( .A1(n640), .A2(n523), .A3(n524), .Y(out1[122]) );
  XOR3X2_HVT U370 ( .A1(n525), .A2(n1377), .A3(n526), .Y(n640) );
  IBUFFX2_HVT U371 ( .A(in[90]), .Y(n670) );
  XOR3X1_HVT U372 ( .A1(n647), .A2(n799), .A3(n204), .Y(out1[74]) );
  XOR2X2_HVT U373 ( .A1(in[52]), .A2(n1032), .Y(n232) );
  INVX1_HVT U374 ( .A(in[52]), .Y(n1354) );
  XOR3X1_HVT U375 ( .A1(n875), .A2(n282), .A3(n240), .Y(n289) );
  INVX2_HVT U376 ( .A(in[119]), .Y(n1376) );
  XNOR3X2_HVT U377 ( .A1(n339), .A2(n1246), .A3(n278), .Y(n372) );
  INVX1_HVT U378 ( .A(in[37]), .Y(n1135) );
  NAND2X0_HVT U379 ( .A1(n663), .A2(n664), .Y(n641) );
  INVX1_HVT U380 ( .A(n237), .Y(n1181) );
  XOR3X1_HVT U381 ( .A1(n357), .A2(n1120), .A3(n358), .Y(out1[43]) );
  XNOR2X2_HVT U382 ( .A1(n1042), .A2(n958), .Y(n104) );
  INVX1_HVT U383 ( .A(n1042), .Y(n118) );
  INVX1_HVT U384 ( .A(n958), .Y(n959) );
  INVX1_HVT U385 ( .A(n350), .Y(n1133) );
  INVX0_HVT U386 ( .A(n717), .Y(n793) );
  INVX1_HVT U387 ( .A(n868), .Y(n642) );
  INVX0_HVT U388 ( .A(n754), .Y(n643) );
  XOR3X1_HVT U389 ( .A1(n1264), .A2(n408), .A3(n415), .Y(n413) );
  OR2X1_HVT U390 ( .A1(n300), .A2(n745), .Y(n789) );
  INVX1_HVT U391 ( .A(n1184), .Y(n644) );
  NBUFFX2_HVT U392 ( .A(n516), .Y(n645) );
  NAND2X0_HVT U393 ( .A1(n775), .A2(n776), .Y(n646) );
  XOR3X2_HVT U394 ( .A1(n447), .A2(n1140), .A3(n218), .Y(n486) );
  XOR3X2_HVT U395 ( .A1(n206), .A2(n751), .A3(n110), .Y(n647) );
  NBUFFX2_HVT U396 ( .A(in[96]), .Y(n648) );
  XNOR2X2_HVT U397 ( .A1(in[43]), .A2(n1353), .Y(n304) );
  XOR3X2_HVT U398 ( .A1(n446), .A2(n649), .A3(n258), .Y(n445) );
  IBUFFX16_HVT U399 ( .A(n1146), .Y(n649) );
  NBUFFX2_HVT U400 ( .A(in[106]), .Y(n650) );
  XNOR2X2_HVT U401 ( .A1(n695), .A2(n1349), .Y(n433) );
  INVX1_HVT U402 ( .A(n20), .Y(n675) );
  INVX0_HVT U403 ( .A(n1074), .Y(n651) );
  NAND2X0_HVT U404 ( .A1(in[40]), .A2(n1353), .Y(n654) );
  NAND2X0_HVT U405 ( .A1(n652), .A2(n653), .Y(n655) );
  NAND2X0_HVT U406 ( .A1(n654), .A2(n655), .Y(n334) );
  INVX0_HVT U407 ( .A(in[40]), .Y(n652) );
  INVX0_HVT U408 ( .A(n1353), .Y(n653) );
  INVX0_HVT U409 ( .A(in[47]), .Y(n1353) );
  INVX0_HVT U410 ( .A(n334), .Y(n1170) );
  IBUFFX2_HVT U411 ( .A(n264), .Y(n656) );
  INVX0_HVT U412 ( .A(n656), .Y(n657) );
  INVX1_HVT U413 ( .A(n658), .Y(n659) );
  XOR2X2_HVT U414 ( .A1(in[101]), .A2(n734), .Y(n76) );
  INVX0_HVT U415 ( .A(n33), .Y(n754) );
  XOR2X1_HVT U416 ( .A1(n119), .A2(n932), .Y(n166) );
  NBUFFX2_HVT U417 ( .A(n568), .Y(n660) );
  NAND2X0_HVT U418 ( .A1(n199), .A2(n951), .Y(n663) );
  NAND2X0_HVT U419 ( .A1(n661), .A2(n662), .Y(n664) );
  NAND2X0_HVT U420 ( .A1(n663), .A2(n664), .Y(n158) );
  INVX0_HVT U421 ( .A(n199), .Y(n661) );
  INVX0_HVT U422 ( .A(n951), .Y(n662) );
  XOR3X2_HVT U423 ( .A1(n272), .A2(n665), .A3(n666), .Y(n368) );
  XOR3X1_HVT U424 ( .A1(n667), .A2(n78), .A3(n79), .Y(out1[95]) );
  IBUFFX16_HVT U425 ( .A(n77), .Y(n667) );
  IBUFFX2_HVT U426 ( .A(n252), .Y(n668) );
  INVX1_HVT U427 ( .A(n668), .Y(n669) );
  XNOR2X2_HVT U428 ( .A1(n109), .A2(n670), .Y(n160) );
  NAND2X0_HVT U429 ( .A1(n7), .A2(n886), .Y(n673) );
  NAND2X0_HVT U430 ( .A1(n671), .A2(n672), .Y(n674) );
  NAND2X0_HVT U431 ( .A1(n673), .A2(n674), .Y(n902) );
  INVX1_HVT U432 ( .A(n432), .Y(n671) );
  IBUFFX2_HVT U433 ( .A(n886), .Y(n672) );
  IBUFFX2_HVT U434 ( .A(n411), .Y(n1017) );
  XOR3X1_HVT U435 ( .A1(n376), .A2(n984), .A3(n378), .Y(n1275) );
  XOR2X2_HVT U436 ( .A1(n68), .A2(n1123), .Y(n580) );
  XOR3X1_HVT U437 ( .A1(n938), .A2(n1242), .A3(n72), .Y(n578) );
  XOR3X2_HVT U438 ( .A1(n675), .A2(n71), .A3(n72), .Y(n67) );
  XNOR2X1_HVT U439 ( .A1(n1145), .A2(n1345), .Y(n54) );
  INVX1_HVT U440 ( .A(in[14]), .Y(n1345) );
  XOR3X2_HVT U441 ( .A1(n1213), .A2(n911), .A3(n95), .Y(n1290) );
  XOR2X2_HVT U442 ( .A1(in[14]), .A2(n833), .Y(n435) );
  XNOR2X2_HVT U443 ( .A1(n206), .A2(n109), .Y(n120) );
  XNOR2X2_HVT U444 ( .A1(n1332), .A2(n639), .Y(n370) );
  XNOR3X1_HVT U445 ( .A1(n1347), .A2(n1346), .A3(n483), .Y(n481) );
  NBUFFX2_HVT U446 ( .A(in[10]), .Y(n678) );
  IBUFFX2_HVT U447 ( .A(n971), .Y(n679) );
  INVX1_HVT U448 ( .A(n1238), .Y(n1239) );
  INVX0_HVT U449 ( .A(n448), .Y(n871) );
  XOR2X2_HVT U450 ( .A1(n209), .A2(n772), .Y(n172) );
  XOR3X2_HVT U451 ( .A1(n220), .A2(n1167), .A3(n191), .Y(out1[69]) );
  IBUFFX2_HVT U452 ( .A(n991), .Y(n680) );
  INVX1_HVT U453 ( .A(n680), .Y(n681) );
  INVX1_HVT U454 ( .A(in[66]), .Y(n991) );
  XOR3X2_HVT U455 ( .A1(n917), .A2(n83), .A3(n141), .Y(n1198) );
  INVX2_HVT U456 ( .A(n1209), .Y(n1215) );
  INVX0_HVT U457 ( .A(n1077), .Y(n1080) );
  XOR2X1_HVT U458 ( .A1(n492), .A2(n493), .Y(n687) );
  INVX2_HVT U459 ( .A(in[70]), .Y(n1360) );
  IBUFFX2_HVT U460 ( .A(n759), .Y(n682) );
  INVX1_HVT U461 ( .A(n682), .Y(n683) );
  IBUFFX2_HVT U462 ( .A(in[3]), .Y(n1125) );
  INVX0_HVT U463 ( .A(in[20]), .Y(n707) );
  INVX1_HVT U464 ( .A(n1179), .Y(n1180) );
  INVX1_HVT U465 ( .A(n1056), .Y(n1057) );
  INVX0_HVT U466 ( .A(n1344), .Y(n831) );
  INVX1_HVT U467 ( .A(n782), .Y(n783) );
  INVX0_HVT U468 ( .A(n1071), .Y(n721) );
  INVX0_HVT U469 ( .A(n65), .Y(n722) );
  NBUFFX2_HVT U470 ( .A(in[86]), .Y(n1335) );
  INVX0_HVT U471 ( .A(n1368), .Y(n913) );
  NBUFFX2_HVT U472 ( .A(in[86]), .Y(n1334) );
  INVX1_HVT U473 ( .A(n338), .Y(n1008) );
  INVX1_HVT U474 ( .A(n484), .Y(n714) );
  INVX0_HVT U475 ( .A(n1378), .Y(n693) );
  INVX1_HVT U476 ( .A(n1307), .Y(n1194) );
  INVX0_HVT U477 ( .A(n306), .Y(n847) );
  INVX0_HVT U478 ( .A(n59), .Y(n940) );
  INVX0_HVT U479 ( .A(n1124), .Y(n804) );
  IBUFFX2_HVT U480 ( .A(n625), .Y(n836) );
  INVX0_HVT U481 ( .A(n574), .Y(n763) );
  INVX0_HVT U482 ( .A(n1372), .Y(n764) );
  INVX0_HVT U483 ( .A(n122), .Y(n841) );
  INVX0_HVT U484 ( .A(n1368), .Y(n753) );
  INVX1_HVT U485 ( .A(n944), .Y(n1369) );
  INVX0_HVT U486 ( .A(n926), .Y(n246) );
  INVX0_HVT U487 ( .A(n318), .Y(n923) );
  INVX1_HVT U488 ( .A(n1063), .Y(n885) );
  INVX0_HVT U489 ( .A(n572), .Y(n702) );
  INVX0_HVT U490 ( .A(n82), .Y(n738) );
  INVX0_HVT U491 ( .A(n131), .Y(n708) );
  INVX1_HVT U492 ( .A(n173), .Y(n818) );
  INVX1_HVT U493 ( .A(n233), .Y(n735) );
  INVX0_HVT U494 ( .A(n339), .Y(n1009) );
  INVX1_HVT U495 ( .A(n1084), .Y(n877) );
  XNOR3X1_HVT U496 ( .A1(n859), .A2(n718), .A3(n439), .Y(n436) );
  XOR3X1_HVT U497 ( .A1(n1086), .A2(n1087), .A3(n1088), .Y(out1[23]) );
  INVX1_HVT U498 ( .A(n437), .Y(n713) );
  INVX0_HVT U499 ( .A(n403), .Y(n912) );
  INVX0_HVT U500 ( .A(n734), .Y(n835) );
  INVX0_HVT U501 ( .A(n1291), .Y(n1119) );
  AND2X1_HVT U502 ( .A1(n17), .A2(n758), .Y(n685) );
  AND2X1_HVT U503 ( .A1(n873), .A2(n866), .Y(n686) );
  XOR2X2_HVT U504 ( .A1(n777), .A2(n1273), .Y(n688) );
  INVX0_HVT U505 ( .A(n1157), .Y(n1158) );
  INVX0_HVT U506 ( .A(in[44]), .Y(n1260) );
  INVX1_HVT U507 ( .A(n293), .Y(n819) );
  INVX1_HVT U508 ( .A(n843), .Y(n844) );
  INVX1_HVT U509 ( .A(n952), .Y(n917) );
  INVX0_HVT U510 ( .A(in[68]), .Y(n952) );
  INVX1_HVT U511 ( .A(n50), .Y(n802) );
  INVX1_HVT U512 ( .A(n523), .Y(n803) );
  INVX1_HVT U513 ( .A(in[61]), .Y(n1358) );
  INVX0_HVT U514 ( .A(n321), .Y(n1285) );
  INVX1_HVT U516 ( .A(in[33]), .Y(n1235) );
  INVX1_HVT U517 ( .A(n814), .Y(n977) );
  INVX1_HVT U518 ( .A(in[49]), .Y(n814) );
  INVX0_HVT U519 ( .A(n790), .Y(n1272) );
  INVX1_HVT U520 ( .A(n1062), .Y(n886) );
  INVX0_HVT U521 ( .A(n989), .Y(n990) );
  NBUFFX2_HVT U523 ( .A(n677), .Y(n691) );
  XNOR2X2_HVT U524 ( .A1(n510), .A2(n693), .Y(n692) );
  NAND2X0_HVT U525 ( .A1(n741), .A2(n740), .Y(n694) );
  XNOR2X2_HVT U526 ( .A1(in[109]), .A2(in[110]), .Y(n581) );
  INVX2_HVT U527 ( .A(in[29]), .Y(n1129) );
  XOR3X2_HVT U528 ( .A1(n480), .A2(n460), .A3(n431), .Y(out1[17]) );
  XOR3X1_HVT U529 ( .A1(n684), .A2(n160), .A3(n161), .Y(out1[82]) );
  INVX0_HVT U530 ( .A(in[126]), .Y(n1311) );
  XOR3X2_HVT U531 ( .A1(n923), .A2(n924), .A3(n268), .Y(n317) );
  INVX1_HVT U532 ( .A(in[110]), .Y(n696) );
  XNOR2X2_HVT U533 ( .A1(n867), .A2(n659), .Y(n270) );
  XNOR2X2_HVT U534 ( .A1(n559), .A2(n783), .Y(n545) );
  INVX1_HVT U535 ( .A(n1240), .Y(n1355) );
  XNOR2X2_HVT U536 ( .A1(n521), .A2(n697), .Y(n1100) );
  XNOR2X1_HVT U537 ( .A1(n940), .A2(n941), .Y(n697) );
  XNOR3X1_HVT U538 ( .A1(n645), .A2(n558), .A3(n517), .Y(n615) );
  INVX0_HVT U539 ( .A(n557), .Y(n704) );
  NAND2X0_HVT U540 ( .A1(n308), .A2(n1266), .Y(n699) );
  NAND2X0_HVT U541 ( .A1(n698), .A2(n323), .Y(n700) );
  NAND2X0_HVT U542 ( .A1(n699), .A2(n700), .Y(n1185) );
  INVX1_HVT U543 ( .A(n308), .Y(n698) );
  XNOR2X1_HVT U544 ( .A1(n1151), .A2(n1342), .Y(n447) );
  XOR3X2_HVT U545 ( .A1(n515), .A2(n743), .A3(n705), .Y(n1320) );
  XNOR2X2_HVT U546 ( .A1(n1134), .A2(n744), .Y(n614) );
  XNOR2X1_HVT U547 ( .A1(n433), .A2(in[25]), .Y(n464) );
  IBUFFX2_HVT U548 ( .A(in[25]), .Y(n920) );
  NBUFFX2_HVT U549 ( .A(n378), .Y(n701) );
  INVX2_HVT U550 ( .A(n847), .Y(n848) );
  INVX0_HVT U551 ( .A(n1228), .Y(n709) );
  INVX1_HVT U553 ( .A(n1228), .Y(n1060) );
  IBUFFX2_HVT U555 ( .A(in[99]), .Y(n1231) );
  XOR3X2_HVT U556 ( .A1(n571), .A2(n702), .A3(n524), .Y(out1[114]) );
  XOR3X2_HVT U557 ( .A1(n703), .A2(n223), .A3(n686), .Y(n1219) );
  XOR3X2_HVT U558 ( .A1(n1250), .A2(n330), .A3(n368), .Y(out1[33]) );
  XNOR2X2_HVT U559 ( .A1(n744), .A2(n1374), .Y(n550) );
  INVX1_HVT U560 ( .A(n704), .Y(n705) );
  XOR2X2_HVT U561 ( .A1(in[125]), .A2(n943), .Y(n530) );
  INVX1_HVT U562 ( .A(n520), .Y(n941) );
  NBUFFX2_HVT U563 ( .A(n657), .Y(n706) );
  XNOR2X2_HVT U564 ( .A1(n455), .A2(n707), .Y(n414) );
  XNOR2X2_HVT U565 ( .A1(n605), .A2(n629), .Y(n510) );
  INVX1_HVT U566 ( .A(in[123]), .Y(n1184) );
  XOR3X2_HVT U567 ( .A1(n135), .A2(n769), .A3(n89), .Y(n187) );
  XNOR2X2_HVT U568 ( .A1(n1073), .A2(n1041), .Y(n535) );
  XOR3X2_HVT U569 ( .A1(n163), .A2(n642), .A3(n164), .Y(n108) );
  INVX0_HVT U570 ( .A(n162), .Y(n800) );
  XNOR2X2_HVT U571 ( .A1(n941), .A2(n644), .Y(n568) );
  IBUFFX2_HVT U573 ( .A(n564), .Y(n1091) );
  XOR3X1_HVT U574 ( .A1(n708), .A2(n132), .A3(n133), .Y(out1[86]) );
  XOR3X1_HVT U575 ( .A1(n165), .A2(n1274), .A3(n167), .Y(out1[81]) );
  NAND2X0_HVT U577 ( .A1(n710), .A2(n1228), .Y(n711) );
  NAND2X0_HVT U578 ( .A1(n709), .A2(n1206), .Y(n712) );
  NAND2X0_HVT U579 ( .A1(n711), .A2(n712), .Y(n520) );
  IBUFFX2_HVT U580 ( .A(n58), .Y(n1278) );
  XOR3X1_HVT U581 ( .A1(n713), .A2(n714), .A3(n715), .Y(out1[15]) );
  XOR3X2_HVT U582 ( .A1(n1342), .A2(n444), .A3(n182), .Y(n715) );
  NAND2X0_HVT U583 ( .A1(n250), .A2(n1244), .Y(n716) );
  AND2X1_HVT U584 ( .A1(n780), .A2(n781), .Y(n717) );
  XOR3X2_HVT U585 ( .A1(n942), .A2(n641), .A3(n198), .Y(out1[75]) );
  XNOR2X2_HVT U587 ( .A1(n169), .A2(n118), .Y(n110) );
  XOR3X2_HVT U588 ( .A1(n319), .A2(n977), .A3(n320), .Y(n268) );
  IBUFFX2_HVT U589 ( .A(n455), .Y(n925) );
  NBUFFX2_HVT U590 ( .A(in[30]), .Y(n718) );
  XOR3X2_HVT U591 ( .A1(n719), .A2(n426), .A3(n427), .Y(out1[26]) );
  XOR3X2_HVT U593 ( .A1(n720), .A2(n278), .A3(n279), .Y(out1[56]) );
  XOR3X2_HVT U594 ( .A1(n1110), .A2(n1306), .A3(n280), .Y(n720) );
  XOR3X2_HVT U595 ( .A1(n722), .A2(n721), .A3(n573), .Y(n524) );
  NAND2X0_HVT U596 ( .A1(n788), .A2(n789), .Y(n723) );
  XNOR2X2_HVT U597 ( .A1(n253), .A2(n1157), .Y(n242) );
  INVX1_HVT U598 ( .A(in[7]), .Y(n1193) );
  INVX1_HVT U599 ( .A(n849), .Y(n724) );
  XOR3X2_HVT U600 ( .A1(n802), .A2(n508), .A3(n464), .Y(n480) );
  XNOR3X2_HVT U601 ( .A1(n482), .A2(n1057), .A3(n112), .Y(n438) );
  INVX1_HVT U602 ( .A(n1132), .Y(n727) );
  INVX1_HVT U603 ( .A(n1343), .Y(n1132) );
  INVX0_HVT U604 ( .A(in[7]), .Y(n1343) );
  INVX0_HVT U605 ( .A(n447), .Y(n805) );
  IBUFFX2_HVT U606 ( .A(n1151), .Y(n1208) );
  XOR3X2_HVT U607 ( .A1(n1325), .A2(n679), .A3(n422), .Y(out1[19]) );
  INVX0_HVT U608 ( .A(in[53]), .Y(n1238) );
  NAND2X0_HVT U609 ( .A1(n353), .A2(n832), .Y(n729) );
  NAND2X0_HVT U610 ( .A1(n703), .A2(n728), .Y(n730) );
  NAND2X0_HVT U611 ( .A1(n729), .A2(n730), .Y(n314) );
  INVX0_HVT U612 ( .A(n832), .Y(n728) );
  NAND2X0_HVT U613 ( .A1(n390), .A2(n1350), .Y(n732) );
  NAND2X0_HVT U614 ( .A1(n731), .A2(n907), .Y(n733) );
  NAND2X0_HVT U615 ( .A1(n732), .A2(n733), .Y(n359) );
  XOR3X2_HVT U616 ( .A1(n393), .A2(n1002), .A3(n372), .Y(out1[32]) );
  XOR3X1_HVT U617 ( .A1(n232), .A2(n735), .A3(n234), .Y(out1[63]) );
  INVX0_HVT U618 ( .A(in[69]), .Y(n1085) );
  IBUFFX2_HVT U619 ( .A(n305), .Y(n736) );
  INVX1_HVT U620 ( .A(n736), .Y(n737) );
  XOR3X2_HVT U622 ( .A1(n335), .A2(n852), .A3(n689), .Y(n273) );
  XOR3X1_HVT U623 ( .A1(n410), .A2(in[20]), .A3(n411), .Y(n409) );
  XOR2X2_HVT U624 ( .A1(n755), .A2(n162), .Y(n165) );
  NAND2X0_HVT U626 ( .A1(n890), .A2(n889), .Y(n739) );
  NAND2X0_HVT U627 ( .A1(n759), .A2(n917), .Y(n740) );
  NAND2X0_HVT U628 ( .A1(n742), .A2(n771), .Y(n741) );
  NAND2X0_HVT U629 ( .A1(n740), .A2(n741), .Y(n146) );
  AND2X1_HVT U630 ( .A1(n770), .A2(n952), .Y(n742) );
  INVX1_HVT U631 ( .A(n593), .Y(n743) );
  INVX1_HVT U632 ( .A(n743), .Y(n744) );
  XNOR2X2_HVT U633 ( .A1(n306), .A2(n1354), .Y(n745) );
  INVX0_HVT U634 ( .A(in[54]), .Y(n1316) );
  NAND2X0_HVT U635 ( .A1(n386), .A2(n1239), .Y(n748) );
  NAND2X0_HVT U636 ( .A1(n746), .A2(n747), .Y(n749) );
  NAND2X0_HVT U637 ( .A1(n748), .A2(n749), .Y(n306) );
  INVX0_HVT U638 ( .A(n386), .Y(n746) );
  INVX0_HVT U639 ( .A(n1239), .Y(n747) );
  XOR3X2_HVT U640 ( .A1(n750), .A2(n157), .A3(n158), .Y(n102) );
  NAND2X0_HVT U641 ( .A1(n825), .A2(n824), .Y(n750) );
  XOR3X1_HVT U642 ( .A1(n1034), .A2(n126), .A3(n85), .Y(n133) );
  INVX1_HVT U643 ( .A(n801), .Y(n751) );
  XOR3X2_HVT U644 ( .A1(n343), .A2(n344), .A3(n752), .Y(out1[47]) );
  XOR3X2_HVT U645 ( .A1(n286), .A2(n1351), .A3(n280), .Y(n752) );
  XOR3X2_HVT U646 ( .A1(n134), .A2(n753), .A3(n139), .Y(n215) );
  INVX1_HVT U647 ( .A(n754), .Y(n755) );
  NAND2X0_HVT U648 ( .A1(n904), .A2(n905), .Y(n756) );
  NAND2X0_HVT U649 ( .A1(n904), .A2(n905), .Y(n757) );
  NAND2X0_HVT U650 ( .A1(n823), .A2(n1000), .Y(n758) );
  XOR3X2_HVT U651 ( .A1(n288), .A2(n1357), .A3(n296), .Y(n382) );
  XNOR2X2_HVT U652 ( .A1(n310), .A2(n454), .Y(n261) );
  INVX0_HVT U653 ( .A(n1291), .Y(n1292) );
  NAND2X0_HVT U654 ( .A1(n770), .A2(n771), .Y(n759) );
  IBUFFX2_HVT U655 ( .A(in[35]), .Y(n832) );
  INVX1_HVT U656 ( .A(n575), .Y(n760) );
  INVX1_HVT U658 ( .A(n760), .Y(n761) );
  XOR3X2_HVT U659 ( .A1(n762), .A2(n320), .A3(n364), .Y(out1[42]) );
  XNOR2X2_HVT U660 ( .A1(n162), .A2(n1164), .Y(n107) );
  INVX0_HVT U661 ( .A(n107), .Y(n855) );
  NAND2X0_HVT U662 ( .A1(in[33]), .A2(in[38]), .Y(n766) );
  NAND2X0_HVT U663 ( .A1(n1235), .A2(n1351), .Y(n767) );
  NAND2X0_HVT U664 ( .A1(n766), .A2(n767), .Y(n388) );
  NAND2X0_HVT U665 ( .A1(n1074), .A2(n907), .Y(n768) );
  INVX0_HVT U666 ( .A(n388), .Y(n1074) );
  XNOR2X2_HVT U667 ( .A1(n1365), .A2(n1317), .Y(n168) );
  INVX1_HVT U668 ( .A(in[85]), .Y(n1365) );
  XOR3X2_HVT U669 ( .A1(n1271), .A2(n238), .A3(n297), .Y(n349) );
  NAND2X0_HVT U670 ( .A1(n790), .A2(n1085), .Y(n770) );
  NAND2X0_HVT U671 ( .A1(n1272), .A2(n769), .Y(n771) );
  INVX0_HVT U672 ( .A(n1085), .Y(n769) );
  IBUFFX2_HVT U673 ( .A(n1141), .Y(n772) );
  XOR3X2_HVT U675 ( .A1(n344), .A2(n346), .A3(n773), .Y(out1[46]) );
  XOR3X2_HVT U676 ( .A1(n291), .A2(n1135), .A3(n244), .Y(n773) );
  NAND2X0_HVT U677 ( .A1(n224), .A2(n1211), .Y(n775) );
  NAND2X0_HVT U678 ( .A1(n774), .A2(n1190), .Y(n776) );
  NAND2X0_HVT U679 ( .A1(n775), .A2(n776), .Y(n150) );
  INVX0_HVT U680 ( .A(n224), .Y(n774) );
  IBUFFX2_HVT U681 ( .A(n774), .Y(n777) );
  NAND2X0_HVT U682 ( .A1(n302), .A2(n301), .Y(n780) );
  NAND2X0_HVT U683 ( .A1(n778), .A2(n779), .Y(n781) );
  NAND2X0_HVT U684 ( .A1(n780), .A2(n8), .Y(n250) );
  IBUFFX2_HVT U685 ( .A(in[110]), .Y(n782) );
  NAND2X0_HVT U686 ( .A1(n1324), .A2(n384), .Y(n786) );
  NAND2X0_HVT U687 ( .A1(n784), .A2(n785), .Y(n787) );
  NAND2X0_HVT U688 ( .A1(n786), .A2(n787), .Y(out1[36]) );
  INVX0_HVT U689 ( .A(n1324), .Y(n784) );
  INVX0_HVT U690 ( .A(n384), .Y(n785) );
  NAND2X0_HVT U691 ( .A1(n745), .A2(n300), .Y(n788) );
  NAND2X0_HVT U692 ( .A1(n788), .A2(n789), .Y(n355) );
  NAND2X0_HVT U693 ( .A1(n1143), .A2(n1142), .Y(n790) );
  NBUFFX2_HVT U694 ( .A(n268), .Y(n791) );
  INVX1_HVT U695 ( .A(in[69]), .Y(n1359) );
  NAND2X0_HVT U696 ( .A1(n717), .A2(n892), .Y(n792) );
  INVX1_HVT U697 ( .A(in[5]), .Y(n794) );
  INVX1_HVT U699 ( .A(n794), .Y(n795) );
  INVX0_HVT U700 ( .A(n348), .Y(n796) );
  INVX1_HVT U701 ( .A(n796), .Y(n797) );
  XOR3X2_HVT U703 ( .A1(n1080), .A2(n284), .A3(n236), .Y(n283) );
  INVX1_HVT U704 ( .A(n1356), .Y(n1032) );
  NBUFFX2_HVT U705 ( .A(n164), .Y(n799) );
  XOR3X2_HVT U706 ( .A1(n275), .A2(n826), .A3(n276), .Y(n1168) );
  XOR3X2_HVT U707 ( .A1(n370), .A2(n1169), .A3(n276), .Y(n367) );
  XOR3X2_HVT U708 ( .A1(n1260), .A2(n295), .A3(n245), .Y(n294) );
  XNOR3X1_HVT U709 ( .A1(n304), .A2(n848), .A3(n737), .Y(n1318) );
  XOR3X1_HVT U710 ( .A1(n241), .A2(n242), .A3(n1255), .Y(out1[61]) );
  XOR3X1_HVT U711 ( .A1(n1239), .A2(n233), .A3(n240), .Y(n1183) );
  XNOR2X2_HVT U712 ( .A1(n63), .A2(n761), .Y(n72) );
  XNOR2X2_HVT U714 ( .A1(n560), .A2(n804), .Y(n552) );
  XOR3X2_HVT U716 ( .A1(n229), .A2(n684), .A3(n204), .Y(out1[66]) );
  XNOR2X2_HVT U717 ( .A1(n210), .A2(n751), .Y(n170) );
  XOR2X2_HVT U718 ( .A1(n318), .A2(in[50]), .Y(n267) );
  INVX0_HVT U719 ( .A(in[70]), .Y(n1291) );
  NAND2X0_HVT U720 ( .A1(n447), .A2(n806), .Y(n807) );
  NAND2X0_HVT U721 ( .A1(n805), .A2(n217), .Y(n808) );
  NAND2X0_HVT U722 ( .A1(n807), .A2(n808), .Y(n400) );
  INVX0_HVT U723 ( .A(n217), .Y(n806) );
  INVX0_HVT U724 ( .A(in[11]), .Y(n1098) );
  NAND2X0_HVT U725 ( .A1(n1328), .A2(n615), .Y(n811) );
  NAND2X0_HVT U726 ( .A1(n809), .A2(n810), .Y(n812) );
  NAND2X0_HVT U727 ( .A1(n811), .A2(n812), .Y(out1[100]) );
  INVX0_HVT U728 ( .A(n615), .Y(n810) );
  NAND2X0_HVT U729 ( .A1(n555), .A2(n982), .Y(n813) );
  XNOR2X2_HVT U730 ( .A1(n1109), .A2(n1305), .Y(n269) );
  IBUFFX2_HVT U731 ( .A(n1109), .Y(n1110) );
  NAND2X0_HVT U732 ( .A1(in[49]), .A2(n1316), .Y(n816) );
  NAND2X0_HVT U733 ( .A1(n814), .A2(n815), .Y(n817) );
  NAND2X0_HVT U734 ( .A1(n816), .A2(n817), .Y(n386) );
  INVX1_HVT U736 ( .A(n1316), .Y(n815) );
  XOR3X1_HVT U737 ( .A1(n818), .A2(n174), .A3(n175), .Y(out1[80]) );
  XNOR2X2_HVT U738 ( .A1(n448), .A2(n1257), .Y(n217) );
  XNOR2X2_HVT U739 ( .A1(n540), .A2(n541), .Y(n498) );
  XOR3X2_HVT U740 ( .A1(n1095), .A2(n1094), .A3(n1293), .Y(out1[98]) );
  XOR3X2_HVT U741 ( .A1(n1377), .A2(n65), .A3(n66), .Y(n1293) );
  XOR2X2_HVT U742 ( .A1(n1316), .A2(n1356), .Y(n318) );
  XOR3X2_HVT U744 ( .A1(n190), .A2(n1304), .A3(n195), .Y(n193) );
  NAND2X0_HVT U745 ( .A1(n1083), .A2(n293), .Y(n820) );
  NAND2X0_HVT U746 ( .A1(n822), .A2(n792), .Y(n821) );
  NAND2X0_HVT U747 ( .A1(n820), .A2(n821), .Y(n299) );
  AND2X1_HVT U748 ( .A1(n716), .A2(n819), .Y(n822) );
  XNOR2X2_HVT U749 ( .A1(n303), .A2(n1249), .Y(n293) );
  XNOR2X2_HVT U750 ( .A1(in[96]), .A2(n1371), .Y(n577) );
  XNOR2X2_HVT U751 ( .A1(in[9]), .A2(in[14]), .Y(n492) );
  INVX1_HVT U752 ( .A(in[63]), .Y(n1014) );
  XNOR2X2_HVT U753 ( .A1(n516), .A2(n1312), .Y(n542) );
  INVX0_HVT U754 ( .A(n830), .Y(n840) );
  XNOR2X2_HVT U755 ( .A1(n493), .A2(n695), .Y(n419) );
  NAND2X0_HVT U756 ( .A1(n200), .A2(in[75]), .Y(n824) );
  NAND2X0_HVT U757 ( .A1(n823), .A2(n1000), .Y(n825) );
  NAND2X0_HVT U758 ( .A1(n968), .A2(n967), .Y(n827) );
  XNOR2X1_HVT U759 ( .A1(in[100]), .A2(n1371), .Y(n541) );
  IBUFFX2_HVT U760 ( .A(in[56]), .Y(n828) );
  INVX1_HVT U761 ( .A(n828), .Y(n829) );
  INVX1_HVT U762 ( .A(n552), .Y(n965) );
  XNOR2X2_HVT U763 ( .A1(n457), .A2(n831), .Y(n830) );
  IBUFFX2_HVT U764 ( .A(n41), .Y(n1089) );
  INVX0_HVT U765 ( .A(n970), .Y(n834) );
  XOR3X1_HVT U766 ( .A1(n531), .A2(n1051), .A3(n1052), .Y(n69) );
  XOR3X2_HVT U767 ( .A1(n835), .A2(n497), .A3(n498), .Y(n496) );
  XOR3X2_HVT U768 ( .A1(n568), .A2(n836), .A3(n521), .Y(n58) );
  XNOR2X2_HVT U769 ( .A1(n1200), .A2(n1335), .Y(n162) );
  INVX0_HVT U770 ( .A(n159), .Y(n837) );
  NAND2X0_HVT U771 ( .A1(n987), .A2(n141), .Y(n838) );
  XNOR2X2_HVT U772 ( .A1(n570), .A2(n1041), .Y(n561) );
  XNOR2X2_HVT U773 ( .A1(n1135), .A2(n1337), .Y(n284) );
  XOR3X2_HVT U774 ( .A1(n400), .A2(n1087), .A3(n445), .Y(out1[22]) );
  XNOR2X2_HVT U775 ( .A1(n1163), .A2(in[77]), .Y(n200) );
  XNOR2X2_HVT U776 ( .A1(in[77]), .A2(n1362), .Y(n210) );
  XOR3X2_HVT U777 ( .A1(n949), .A2(n867), .A3(n273), .Y(n332) );
  XOR3X2_HVT U778 ( .A1(n842), .A2(n841), .A3(n26), .Y(out1[88]) );
  XOR3X2_HVT U779 ( .A1(n1054), .A2(n1333), .A3(n124), .Y(n842) );
  XOR2X2_HVT U780 ( .A1(n63), .A2(n1101), .Y(n573) );
  XOR3X2_HVT U781 ( .A1(n207), .A2(n1173), .A3(n208), .Y(out1[73]) );
  INVX0_HVT U782 ( .A(n1053), .Y(n1054) );
  NAND2X0_HVT U783 ( .A1(n901), .A2(n900), .Y(n845) );
  NAND2X0_HVT U784 ( .A1(n1068), .A2(n1069), .Y(n846) );
  XOR3X2_HVT U785 ( .A1(n1299), .A2(n504), .A3(n505), .Y(out1[125]) );
  XOR3X2_HVT U786 ( .A1(n1136), .A2(n506), .A3(n603), .Y(n505) );
  XOR3X2_HVT U787 ( .A1(n1294), .A2(n550), .A3(n827), .Y(n549) );
  INVX0_HVT U788 ( .A(n849), .Y(n850) );
  XNOR2X2_HVT U789 ( .A1(n569), .A2(n1370), .Y(n602) );
  XNOR2X1_HVT U790 ( .A1(n1365), .A2(in[80]), .Y(n122) );
  XNOR2X2_HVT U791 ( .A1(n274), .A2(n851), .Y(n264) );
  XNOR2X2_HVT U792 ( .A1(n333), .A2(n977), .Y(n272) );
  XOR3X2_HVT U793 ( .A1(n346), .A2(n1001), .A3(n381), .Y(out1[38]) );
  INVX1_HVT U794 ( .A(n1053), .Y(n944) );
  INVX1_HVT U795 ( .A(n1251), .Y(n1222) );
  XNOR2X2_HVT U796 ( .A1(n1237), .A2(n1355), .Y(n278) );
  INVX0_HVT U797 ( .A(n961), .Y(n854) );
  INVX1_HVT U798 ( .A(in[26]), .Y(n961) );
  NAND2X0_HVT U799 ( .A1(n107), .A2(n914), .Y(n857) );
  NAND2X0_HVT U800 ( .A1(n855), .A2(n856), .Y(n858) );
  NAND2X0_HVT U801 ( .A1(n857), .A2(n858), .Y(n204) );
  INVX1_HVT U802 ( .A(n914), .Y(n856) );
  XOR2X1_HVT U803 ( .A1(n326), .A2(in[12]), .Y(n399) );
  NBUFFX2_HVT U804 ( .A(n1280), .Y(n859) );
  XOR3X1_HVT U805 ( .A1(n1128), .A2(n408), .A3(n409), .Y(out1[29]) );
  XNOR2X2_HVT U806 ( .A1(in[92]), .A2(n1369), .Y(n125) );
  INVX1_HVT U807 ( .A(n860), .Y(n861) );
  NBUFFX2_HVT U808 ( .A(n102), .Y(n862) );
  XOR3X2_HVT U809 ( .A1(n919), .A2(n1263), .A3(n685), .Y(n227) );
  XOR3X2_HVT U810 ( .A1(n221), .A2(n863), .A3(n1166), .Y(n1327) );
  XOR3X2_HVT U811 ( .A1(n394), .A2(n395), .A3(n864), .Y(out1[31]) );
  XOR3X2_HVT U812 ( .A1(n114), .A2(n1267), .A3(n397), .Y(n864) );
  IBUFFX2_HVT U813 ( .A(n1090), .Y(n865) );
  NAND2X0_HVT U814 ( .A1(n872), .A2(n989), .Y(n866) );
  INVX1_HVT U815 ( .A(n1169), .Y(n867) );
  NAND2X0_HVT U816 ( .A1(n1317), .A2(in[81]), .Y(n869) );
  NAND2X0_HVT U817 ( .A1(in[86]), .A2(n868), .Y(n870) );
  NAND2X0_HVT U818 ( .A1(n869), .A2(n870), .Y(n224) );
  INVX1_HVT U819 ( .A(in[81]), .Y(n868) );
  XNOR2X2_HVT U820 ( .A1(n725), .A2(n871), .Y(n487) );
  XNOR2X2_HVT U821 ( .A1(in[80]), .A2(n1366), .Y(n171) );
  XNOR2X2_HVT U822 ( .A1(n98), .A2(n843), .Y(n87) );
  XOR2X1_HVT U823 ( .A1(n15), .A2(n846), .Y(n105) );
  NAND2X0_HVT U824 ( .A1(n360), .A2(n990), .Y(n873) );
  NAND2X0_HVT U825 ( .A1(n872), .A2(n989), .Y(n874) );
  NAND2X0_HVT U826 ( .A1(n873), .A2(n874), .Y(n312) );
  INVX0_HVT U827 ( .A(n360), .Y(n872) );
  INVX0_HVT U828 ( .A(n1036), .Y(n978) );
  INVX0_HVT U829 ( .A(n1361), .Y(n1261) );
  XNOR2X1_HVT U830 ( .A1(n304), .A2(in[60]), .Y(n244) );
  XNOR2X2_HVT U831 ( .A1(n1103), .A2(n452), .Y(n449) );
  XNOR3X2_HVT U832 ( .A1(n1216), .A2(n639), .A3(n235), .Y(n371) );
  INVX1_HVT U833 ( .A(n144), .Y(n1212) );
  XOR3X1_HVT U834 ( .A1(n1107), .A2(n1108), .A3(n375), .Y(n536) );
  XNOR2X2_HVT U835 ( .A1(in[73]), .A2(n1362), .Y(n202) );
  XOR3X2_HVT U836 ( .A1(n478), .A2(n1061), .A3(n406), .Y(n475) );
  XOR3X2_HVT U837 ( .A1(n290), .A2(n876), .A3(n295), .Y(n381) );
  INVX1_HVT U838 ( .A(n1040), .Y(n878) );
  INVX1_HVT U839 ( .A(n96), .Y(n1040) );
  NAND2X0_HVT U840 ( .A1(n401), .A2(n880), .Y(n881) );
  NAND2X0_HVT U841 ( .A1(n879), .A2(n446), .Y(n882) );
  NAND2X0_HVT U842 ( .A1(n881), .A2(n882), .Y(n218) );
  INVX0_HVT U843 ( .A(n401), .Y(n879) );
  INVX0_HVT U844 ( .A(n446), .Y(n880) );
  NBUFFX2_HVT U845 ( .A(n612), .Y(n883) );
  XNOR2X2_HVT U846 ( .A1(n326), .A2(n1349), .Y(n446) );
  AND2X1_HVT U847 ( .A1(n1079), .A2(n1078), .Y(n884) );
  XOR3X2_HVT U848 ( .A1(n885), .A2(n886), .A3(n51), .Y(n461) );
  INVX2_HVT U849 ( .A(in[84]), .Y(n1364) );
  IBUFFX2_HVT U850 ( .A(n314), .Y(n1120) );
  NAND2X0_HVT U851 ( .A1(n1070), .A2(n424), .Y(n889) );
  NAND2X0_HVT U852 ( .A1(n887), .A2(n888), .Y(n890) );
  NAND2X0_HVT U853 ( .A1(n890), .A2(n889), .Y(n375) );
  INVX0_HVT U854 ( .A(n1070), .Y(n887) );
  INVX0_HVT U855 ( .A(n424), .Y(n888) );
  NBUFFX2_HVT U856 ( .A(in[21]), .Y(n891) );
  XOR2X2_HVT U857 ( .A1(n416), .A2(n363), .Y(n408) );
  XOR3X1_HVT U858 ( .A1(n1270), .A2(n487), .A3(n488), .Y(out1[13]) );
  XNOR2X2_HVT U859 ( .A1(n303), .A2(n1240), .Y(n241) );
  INVX0_HVT U860 ( .A(n299), .Y(n997) );
  XNOR3X2_HVT U861 ( .A1(n448), .A2(n850), .A3(n897), .Y(n453) );
  NAND2X0_HVT U862 ( .A1(n717), .A2(n892), .Y(n893) );
  NAND2X0_HVT U863 ( .A1(n893), .A2(n716), .Y(n1083) );
  INVX0_HVT U864 ( .A(n1244), .Y(n892) );
  XNOR2X2_HVT U865 ( .A1(n377), .A2(n1349), .Y(n416) );
  IBUFFX2_HVT U866 ( .A(in[91]), .Y(n894) );
  INVX1_HVT U867 ( .A(n894), .Y(n895) );
  INVX0_HVT U868 ( .A(n458), .Y(n896) );
  INVX0_HVT U869 ( .A(n896), .Y(n897) );
  NAND2X0_HVT U870 ( .A1(n93), .A2(n1367), .Y(n900) );
  NAND2X0_HVT U871 ( .A1(n898), .A2(n899), .Y(n901) );
  NAND2X0_HVT U872 ( .A1(n901), .A2(n900), .Y(n144) );
  IBUFFX2_HVT U873 ( .A(n1367), .Y(n899) );
  INVX1_HVT U874 ( .A(in[92]), .Y(n1367) );
  INVX1_HVT U875 ( .A(n1350), .Y(n907) );
  XNOR2X2_HVT U876 ( .A1(n1192), .A2(n959), .Y(n124) );
  INVX0_HVT U877 ( .A(n199), .Y(n919) );
  NAND2X0_HVT U878 ( .A1(in[66]), .A2(n916), .Y(n904) );
  NAND2X0_HVT U879 ( .A1(n991), .A2(n903), .Y(n905) );
  INVX0_HVT U880 ( .A(n1361), .Y(n903) );
  OR2X1_HVT U881 ( .A1(n1203), .A2(n490), .Y(n1160) );
  NAND2X0_HVT U882 ( .A1(n908), .A2(n768), .Y(n906) );
  XOR3X2_HVT U883 ( .A1(n53), .A2(n54), .A3(n55), .Y(n1326) );
  XNOR2X2_HVT U884 ( .A1(n474), .A2(n1031), .Y(n324) );
  NAND2X0_HVT U885 ( .A1(n388), .A2(n1350), .Y(n908) );
  NAND2X0_HVT U886 ( .A1(n1074), .A2(n907), .Y(n909) );
  NAND2X0_HVT U887 ( .A1(n909), .A2(n908), .Y(n356) );
  NAND2X0_HVT U888 ( .A1(n988), .A2(n838), .Y(n910) );
  XOR3X2_HVT U889 ( .A1(n402), .A2(n912), .A3(n485), .Y(out1[2]) );
  XOR3X2_HVT U890 ( .A1(n1007), .A2(n1339), .A3(n265), .Y(n357) );
  XNOR2X2_HVT U891 ( .A1(n98), .A2(n913), .Y(n136) );
  IBUFFX2_HVT U892 ( .A(n451), .Y(n1270) );
  IBUFFX2_HVT U893 ( .A(n489), .Y(n970) );
  XNOR2X2_HVT U894 ( .A1(n160), .A2(n1141), .Y(n914) );
  IBUFFX2_HVT U895 ( .A(n470), .Y(n1107) );
  XNOR2X1_HVT U896 ( .A1(n724), .A2(n27), .Y(n256) );
  NBUFFX2_HVT U897 ( .A(n219), .Y(n915) );
  INVX0_HVT U898 ( .A(in[71]), .Y(n916) );
  IBUFFX2_HVT U899 ( .A(n861), .Y(n1217) );
  XNOR2X2_HVT U900 ( .A1(n1194), .A2(n1333), .Y(n80) );
  INVX0_HVT U901 ( .A(n140), .Y(n987) );
  NAND2X0_HVT U902 ( .A1(n1011), .A2(n769), .Y(n918) );
  INVX1_HVT U903 ( .A(n149), .Y(n1011) );
  IBUFFX2_HVT U904 ( .A(in[1]), .Y(n1340) );
  XNOR2X2_HVT U905 ( .A1(n205), .A2(n681), .Y(n164) );
  XNOR3X2_HVT U906 ( .A1(n130), .A2(n1360), .A3(n124), .Y(n185) );
  XOR3X2_HVT U907 ( .A1(n921), .A2(n932), .A3(n643), .Y(n229) );
  XNOR2X2_HVT U908 ( .A1(n891), .A2(n1347), .Y(n465) );
  XNOR2X2_HVT U909 ( .A1(n168), .A2(in[81]), .Y(n116) );
  IBUFFX16_HVT U910 ( .A(n1084), .Y(n924) );
  XOR2X2_HVT U911 ( .A1(n428), .A2(n854), .Y(n476) );
  XOR2X2_HVT U912 ( .A1(in[30]), .A2(n1280), .Y(n428) );
  XNOR2X2_HVT U913 ( .A1(n252), .A2(n875), .Y(n296) );
  XOR3X2_HVT U914 ( .A1(n292), .A2(n819), .A3(n294), .Y(out1[53]) );
  XNOR2X2_HVT U915 ( .A1(n478), .A2(n865), .Y(n429) );
  INVX0_HVT U916 ( .A(n414), .Y(n1264) );
  XOR3X2_HVT U917 ( .A1(n1249), .A2(n669), .A3(n242), .Y(n926) );
  NAND2X0_HVT U918 ( .A1(n1286), .A2(n1285), .Y(n928) );
  NAND2X0_HVT U919 ( .A1(n927), .A2(n321), .Y(n929) );
  NAND2X0_HVT U920 ( .A1(n929), .A2(n928), .Y(out1[4]) );
  INVX0_HVT U921 ( .A(n1286), .Y(n927) );
  XOR3X2_HVT U922 ( .A1(n391), .A2(n690), .A3(n364), .Y(out1[34]) );
  NBUFFX2_HVT U923 ( .A(in[32]), .Y(n930) );
  NAND2X0_HVT U924 ( .A1(n1169), .A2(n1332), .Y(n931) );
  INVX0_HVT U925 ( .A(n1327), .Y(n1175) );
  IBUFFX2_HVT U926 ( .A(in[93]), .Y(n1368) );
  INVX1_HVT U927 ( .A(in[55]), .Y(n1247) );
  INVX1_HVT U928 ( .A(n1370), .Y(n1232) );
  INVX1_HVT U929 ( .A(in[101]), .Y(n1370) );
  INVX1_HVT U930 ( .A(n1294), .Y(n1114) );
  INVX0_HVT U931 ( .A(in[75]), .Y(n1000) );
  INVX0_HVT U932 ( .A(n1374), .Y(n1136) );
  INVX0_HVT U933 ( .A(n1231), .Y(n936) );
  INVX0_HVT U934 ( .A(n1210), .Y(n1190) );
  INVX0_HVT U935 ( .A(n1364), .Y(n1229) );
  INVX1_HVT U936 ( .A(n166), .Y(n1274) );
  INVX1_HVT U937 ( .A(n169), .Y(n1111) );
  INVX1_HVT U938 ( .A(n307), .Y(n1308) );
  INVX0_HVT U939 ( .A(n333), .Y(n949) );
  IBUFFX2_HVT U940 ( .A(n462), .Y(n1063) );
  INVX1_HVT U941 ( .A(n589), .Y(n1043) );
  INVX0_HVT U942 ( .A(n63), .Y(n1094) );
  INVX0_HVT U943 ( .A(n68), .Y(n1112) );
  INVX0_HVT U944 ( .A(n184), .Y(n969) );
  INVX0_HVT U945 ( .A(n213), .Y(n960) );
  INVX1_HVT U946 ( .A(n379), .Y(n1001) );
  INVX0_HVT U947 ( .A(n284), .Y(n1002) );
  INVX1_HVT U948 ( .A(n698), .Y(n1005) );
  INVX1_HVT U949 ( .A(n985), .Y(n986) );
  INVX1_HVT U950 ( .A(n1072), .Y(n1061) );
  INVX1_HVT U951 ( .A(n441), .Y(n1087) );
  INVX0_HVT U952 ( .A(in[76]), .Y(n1162) );
  INVX1_HVT U953 ( .A(in[124]), .Y(n1378) );
  INVX0_HVT U954 ( .A(in[108]), .Y(n1294) );
  XOR3X1_HVT U955 ( .A1(n588), .A2(n589), .A3(n934), .Y(out1[111]) );
  XOR3X2_HVT U956 ( .A1(n541), .A2(n1298), .A3(n533), .Y(n934) );
  XOR2X2_HVT U957 ( .A1(n783), .A2(n1060), .Y(n533) );
  XOR3X2_HVT U958 ( .A1(n614), .A2(n1113), .A3(n953), .Y(n1328) );
  XNOR2X2_HVT U959 ( .A1(in[122]), .A2(n1379), .Y(n59) );
  XNOR2X2_HVT U960 ( .A1(n57), .A2(n936), .Y(n935) );
  INVX0_HVT U961 ( .A(n577), .Y(n1051) );
  XNOR2X2_HVT U962 ( .A1(in[98]), .A2(n937), .Y(n604) );
  INVX1_HVT U963 ( .A(n1165), .Y(n1031) );
  INVX0_HVT U964 ( .A(n440), .Y(n1086) );
  XNOR3X1_HVT U965 ( .A1(n285), .A2(n1305), .A3(n338), .Y(n380) );
  XNOR3X1_HVT U966 ( .A1(n1336), .A2(n1259), .A3(n587), .Y(n584) );
  XNOR3X1_HVT U967 ( .A1(n783), .A2(n76), .A3(n498), .Y(n539) );
  NAND2X0_HVT U968 ( .A1(n955), .A2(n956), .Y(n938) );
  XNOR3X1_HVT U969 ( .A1(n178), .A2(n179), .A3(n180), .Y(out1[7]) );
  XOR2X2_HVT U970 ( .A1(n435), .A2(n678), .Y(n405) );
  INVX1_HVT U971 ( .A(n1031), .Y(n1140) );
  INVX1_HVT U972 ( .A(n794), .Y(n1165) );
  INVX0_HVT U973 ( .A(n1227), .Y(n975) );
  XOR3X2_HVT U974 ( .A1(n341), .A2(n765), .A3(n1110), .Y(n393) );
  XOR3X1_HVT U975 ( .A1(n542), .A2(n1234), .A3(n544), .Y(out1[118]) );
  XOR3X2_HVT U976 ( .A1(n543), .A2(n1378), .A3(n551), .Y(n613) );
  INVX0_HVT U977 ( .A(n1352), .Y(n939) );
  XNOR3X1_HVT U978 ( .A1(n183), .A2(n184), .A3(n185), .Y(out1[79]) );
  XNOR3X1_HVT U979 ( .A1(n844), .A2(n147), .A3(n683), .Y(n222) );
  IBUFFX2_HVT U980 ( .A(n756), .Y(n948) );
  XOR3X2_HVT U981 ( .A1(n43), .A2(n298), .A3(n105), .Y(n942) );
  INVX1_HVT U982 ( .A(n1329), .Y(n1067) );
  XNOR2X2_HVT U983 ( .A1(in[107]), .A2(n635), .Y(n559) );
  NAND2X0_HVT U984 ( .A1(n1205), .A2(n362), .Y(n946) );
  NAND2X0_HVT U985 ( .A1(n884), .A2(n945), .Y(n947) );
  NAND2X0_HVT U986 ( .A1(n947), .A2(n946), .Y(n354) );
  INVX0_HVT U987 ( .A(in[45]), .Y(n1205) );
  XOR3X2_HVT U988 ( .A1(n152), .A2(n948), .A3(n101), .Y(n198) );
  XOR3X2_HVT U989 ( .A1(n136), .A2(n1152), .A3(n138), .Y(out1[85]) );
  XOR3X2_HVT U990 ( .A1(n1162), .A2(n139), .A3(n910), .Y(n138) );
  XOR3X2_HVT U991 ( .A1(n1192), .A2(n128), .A3(n81), .Y(n127) );
  XOR3X2_HVT U992 ( .A1(n227), .A2(n688), .A3(n198), .Y(out1[67]) );
  XNOR2X2_HVT U993 ( .A1(n1373), .A2(n1312), .Y(n497) );
  XNOR2X2_HVT U994 ( .A1(n96), .A2(n952), .Y(n132) );
  NAND2X0_HVT U995 ( .A1(n813), .A2(n983), .Y(n953) );
  NAND2X0_HVT U996 ( .A1(in[117]), .A2(n1315), .Y(n955) );
  NAND2X0_HVT U997 ( .A1(n954), .A2(n1336), .Y(n956) );
  NAND2X0_HVT U998 ( .A1(n955), .A2(n956), .Y(n582) );
  INVX0_HVT U999 ( .A(in[117]), .Y(n954) );
  XNOR3X1_HVT U1000 ( .A1(n287), .A2(n52), .A3(n289), .Y(out1[54]) );
  XNOR2X2_HVT U1001 ( .A1(n575), .A2(in[114]), .Y(n526) );
  XNOR2X2_HVT U1002 ( .A1(n1054), .A2(n1329), .Y(n109) );
  NAND2X0_HVT U1003 ( .A1(n1213), .A2(n845), .Y(n957) );
  XNOR2X2_HVT U1004 ( .A1(n147), .A2(n878), .Y(n137) );
  XNOR3X1_HVT U1005 ( .A1(n975), .A2(n1312), .A3(n535), .Y(n532) );
  XOR2X2_HVT U1006 ( .A1(n397), .A2(n443), .Y(n182) );
  INVX1_HVT U1007 ( .A(n500), .Y(n1003) );
  XNOR2X2_HVT U1008 ( .A1(n253), .A2(n876), .Y(n292) );
  XOR3X2_HVT U1009 ( .A1(n186), .A2(n960), .A3(n215), .Y(out1[70]) );
  NAND2X0_HVT U1010 ( .A1(n962), .A2(in[26]), .Y(n963) );
  NAND2X0_HVT U1011 ( .A1(n961), .A2(n1104), .Y(n964) );
  NAND2X0_HVT U1012 ( .A1(n964), .A2(n963), .Y(n377) );
  XNOR2X2_HVT U1013 ( .A1(n677), .A2(n491), .Y(n596) );
  XOR3X1_HVT U1014 ( .A1(n1282), .A2(n1283), .A3(n1284), .Y(out1[5]) );
  XOR3X2_HVT U1015 ( .A1(n1188), .A2(n962), .A3(n113), .Y(n617) );
  NAND2X0_HVT U1016 ( .A1(n552), .A2(n966), .Y(n967) );
  NAND2X0_HVT U1017 ( .A1(n965), .A2(n551), .Y(n968) );
  INVX0_HVT U1018 ( .A(n551), .Y(n966) );
  XNOR2X2_HVT U1019 ( .A1(n574), .A2(n650), .Y(n65) );
  XOR3X2_HVT U1020 ( .A1(n969), .A2(n186), .A3(n187), .Y(out1[78]) );
  XOR3X2_HVT U1021 ( .A1(n132), .A2(n1367), .A3(n140), .Y(n220) );
  NAND2X0_HVT U1022 ( .A1(n834), .A2(n467), .Y(n972) );
  NAND2X0_HVT U1023 ( .A1(n971), .A2(n970), .Y(n973) );
  NAND2X0_HVT U1024 ( .A1(n973), .A2(n972), .Y(n1070) );
  XNOR2X2_HVT U1025 ( .A1(in[5]), .A2(n1099), .Y(n462) );
  XOR3X1_HVT U1026 ( .A1(n1308), .A2(n1005), .A3(n309), .Y(out1[51]) );
  XOR2X2_HVT U1027 ( .A1(n281), .A2(n232), .Y(n343) );
  XNOR2X2_HVT U1028 ( .A1(n366), .A2(n1050), .Y(n319) );
  XNOR2X2_HVT U1029 ( .A1(n566), .A2(n976), .Y(n61) );
  XNOR2X2_HVT U1030 ( .A1(n251), .A2(n1271), .Y(n288) );
  XNOR2X2_HVT U1031 ( .A1(in[25]), .A2(n1349), .Y(n493) );
  NAND2X0_HVT U1032 ( .A1(n1036), .A2(n260), .Y(n980) );
  NAND2X0_HVT U1033 ( .A1(n978), .A2(n979), .Y(n981) );
  NAND2X0_HVT U1034 ( .A1(n981), .A2(n980), .Y(out1[59]) );
  INVX0_HVT U1035 ( .A(n260), .Y(n979) );
  XNOR2X2_HVT U1036 ( .A1(n416), .A2(n1129), .Y(n452) );
  XOR2X2_HVT U1037 ( .A1(n96), .A2(n1335), .Y(n82) );
  NAND2X0_HVT U1038 ( .A1(n692), .A2(n511), .Y(n983) );
  NAND2X0_HVT U1039 ( .A1(n813), .A2(n983), .Y(n601) );
  XOR2X2_HVT U1040 ( .A1(in[68]), .A2(n1261), .Y(n130) );
  XOR3X2_HVT U1041 ( .A1(n423), .A2(n618), .A3(n424), .Y(n420) );
  XNOR2X2_HVT U1042 ( .A1(in[24]), .A2(in[31]), .Y(n1281) );
  XOR3X2_HVT U1043 ( .A1(n1262), .A2(n87), .A3(n88), .Y(out1[93]) );
  INVX1_HVT U1044 ( .A(n618), .Y(n984) );
  IBUFFX2_HVT U1045 ( .A(in[17]), .Y(n985) );
  XNOR2X2_HVT U1046 ( .A1(n104), .A2(n895), .Y(n152) );
  XNOR2X2_HVT U1047 ( .A1(n370), .A2(n1084), .Y(n335) );
  NAND2X0_HVT U1048 ( .A1(n140), .A2(n1004), .Y(n988) );
  NAND2X0_HVT U1049 ( .A1(n988), .A2(n838), .Y(n90) );
  INVX1_HVT U1050 ( .A(in[65]), .Y(n1141) );
  INVX0_HVT U1051 ( .A(n296), .Y(n1131) );
  IBUFFX2_HVT U1052 ( .A(n1215), .Y(n1216) );
  NAND2X0_HVT U1053 ( .A1(n509), .A2(n1096), .Y(n994) );
  NAND2X0_HVT U1054 ( .A1(n992), .A2(n993), .Y(n995) );
  NAND2X0_HVT U1055 ( .A1(n994), .A2(n995), .Y(out1[124]) );
  INVX0_HVT U1056 ( .A(n1096), .Y(n993) );
  XOR3X2_HVT U1057 ( .A1(n1268), .A2(n511), .A3(n512), .Y(n509) );
  NAND2X0_HVT U1058 ( .A1(n1318), .A2(n299), .Y(n998) );
  NAND2X0_HVT U1059 ( .A1(n997), .A2(n996), .Y(n999) );
  NAND2X0_HVT U1060 ( .A1(n999), .A2(n998), .Y(out1[52]) );
  INVX0_HVT U1061 ( .A(n1318), .Y(n996) );
  OR2X1_HVT U1062 ( .A1(n1252), .A2(n1321), .Y(n1039) );
  XNOR2X1_HVT U1063 ( .A1(n558), .A2(n1041), .Y(n503) );
  XNOR2X2_HVT U1064 ( .A1(n513), .A2(n1241), .Y(n543) );
  AND2X1_HVT U1065 ( .A1(n1012), .A2(n918), .Y(n1004) );
  XOR2X2_HVT U1066 ( .A1(n537), .A2(n494), .Y(n588) );
  XOR3X2_HVT U1067 ( .A1(n588), .A2(n610), .A3(n1331), .Y(out1[103]) );
  XOR3X2_HVT U1068 ( .A1(n1006), .A2(n782), .A3(n75), .Y(n609) );
  NAND2X0_HVT U1069 ( .A1(n1171), .A2(n931), .Y(n1007) );
  XOR3X1_HVT U1070 ( .A1(n1008), .A2(n1009), .A3(n1010), .Y(out1[48]) );
  XOR3X2_HVT U1071 ( .A1(n1338), .A2(n1216), .A3(n279), .Y(n1010) );
  NAND2X0_HVT U1072 ( .A1(n1045), .A2(n1085), .Y(n1012) );
  NAND2X0_HVT U1073 ( .A1(n1011), .A2(n769), .Y(n1013) );
  NAND2X0_HVT U1074 ( .A1(n1013), .A2(n1012), .Y(n141) );
  XNOR2X2_HVT U1075 ( .A1(n148), .A2(n1192), .Y(n134) );
  XOR3X2_HVT U1076 ( .A1(n89), .A2(n1229), .A3(n90), .Y(n88) );
  XNOR2X2_HVT U1077 ( .A1(n1035), .A2(n347), .Y(n176) );
  IBUFFX2_HVT U1078 ( .A(in[74]), .Y(n1015) );
  INVX1_HVT U1079 ( .A(n1015), .Y(n1016) );
  INVX0_HVT U1080 ( .A(n503), .Y(n1299) );
  XNOR2X2_HVT U1081 ( .A1(n547), .A2(n503), .Y(n597) );
  XNOR2X1_HVT U1082 ( .A1(in[40]), .A2(n945), .Y(n341) );
  IBUFFX2_HVT U1083 ( .A(n255), .Y(n1282) );
  NAND2X0_HVT U1084 ( .A1(n1319), .A2(n143), .Y(n1021) );
  NAND2X0_HVT U1085 ( .A1(n1019), .A2(n1020), .Y(n1022) );
  NAND2X0_HVT U1086 ( .A1(n1021), .A2(n1022), .Y(out1[84]) );
  INVX0_HVT U1087 ( .A(n1319), .Y(n1020) );
  XNOR2X2_HVT U1088 ( .A1(in[19]), .A2(n1056), .Y(n418) );
  INVX1_HVT U1089 ( .A(n407), .Y(n1128) );
  NAND2X0_HVT U1090 ( .A1(n1253), .A2(n1243), .Y(n1025) );
  NAND2X0_HVT U1091 ( .A1(n1023), .A2(n1024), .Y(n1026) );
  NAND2X0_HVT U1092 ( .A1(n1025), .A2(n1026), .Y(out1[44]) );
  INVX0_HVT U1093 ( .A(n1243), .Y(n1024) );
  INVX1_HVT U1094 ( .A(in[78]), .Y(n1362) );
  XNOR2X1_HVT U1095 ( .A1(n99), .A2(n1333), .Y(n131) );
  NAND2X0_HVT U1096 ( .A1(n1290), .A2(n91), .Y(n1029) );
  NAND2X0_HVT U1097 ( .A1(n1027), .A2(n1028), .Y(n1030) );
  NAND2X0_HVT U1098 ( .A1(n1030), .A2(n1029), .Y(out1[92]) );
  INVX0_HVT U1099 ( .A(n1290), .Y(n1027) );
  INVX0_HVT U1100 ( .A(n91), .Y(n1028) );
  INVX1_HVT U1101 ( .A(n1089), .Y(n1108) );
  XNOR2X2_HVT U1102 ( .A1(n206), .A2(n1016), .Y(n163) );
  XNOR2X2_HVT U1103 ( .A1(n304), .A2(n1080), .Y(n290) );
  XOR3X2_HVT U1104 ( .A1(n341), .A2(n1032), .A3(n342), .Y(n279) );
  INVX1_HVT U1105 ( .A(n483), .Y(n1055) );
  NAND2X0_HVT U1106 ( .A1(n1048), .A2(n1047), .Y(n1033) );
  XNOR2X2_HVT U1107 ( .A1(n262), .A2(n1037), .Y(n1036) );
  NAND2X0_HVT U1108 ( .A1(n1252), .A2(n1321), .Y(n1038) );
  NAND2X0_HVT U1109 ( .A1(n1038), .A2(n1039), .Y(out1[116]) );
  XOR3X2_HVT U1110 ( .A1(n1040), .A2(n1180), .A3(n87), .Y(n91) );
  INVX0_HVT U1111 ( .A(n579), .Y(n1052) );
  XNOR2X2_HVT U1112 ( .A1(n530), .A2(n1377), .Y(n579) );
  XNOR2X2_HVT U1113 ( .A1(n59), .A2(n1312), .Y(n515) );
  XNOR2X2_HVT U1114 ( .A1(n516), .A2(in[108]), .Y(n500) );
  XNOR2X2_HVT U1115 ( .A1(in[88]), .A2(n598), .Y(n1042) );
  XNOR2X2_HVT U1116 ( .A1(n1259), .A2(n696), .Y(n574) );
  XNOR2X2_HVT U1117 ( .A1(n1115), .A2(n1315), .Y(n575) );
  XOR3X2_HVT U1118 ( .A1(n1043), .A2(n591), .A3(n592), .Y(out1[110]) );
  XOR3X2_HVT U1119 ( .A1(n100), .A2(n1044), .A3(n862), .Y(out1[91]) );
  XNOR2X2_HVT U1120 ( .A1(n756), .A2(n1292), .Y(n1045) );
  XOR3X2_HVT U1121 ( .A1(n535), .A2(n1116), .A3(n587), .Y(n75) );
  XOR3X1_HVT U1122 ( .A1(n803), .A2(n1225), .A3(n1226), .Y(out1[106]) );
  NAND2X0_HVT U1123 ( .A1(n1131), .A2(n297), .Y(n1047) );
  NAND2X0_HVT U1124 ( .A1(n1046), .A2(n296), .Y(n1048) );
  NAND2X0_HVT U1125 ( .A1(n1047), .A2(n1048), .Y(n245) );
  INVX0_HVT U1126 ( .A(n297), .Y(n1046) );
  XOR3X1_HVT U1127 ( .A1(n1354), .A2(n244), .A3(n1033), .Y(n1255) );
  XNOR2X2_HVT U1128 ( .A1(n474), .A2(n473), .Y(n376) );
  XNOR2X1_HVT U1129 ( .A1(n418), .A2(n1341), .Y(n258) );
  XOR3X2_HVT U1130 ( .A1(n591), .A2(n610), .A3(n1314), .Y(out1[102]) );
  INVX1_HVT U1131 ( .A(n1049), .Y(n1050) );
  XNOR2X2_HVT U1132 ( .A1(n188), .A2(n1360), .Y(n135) );
  XNOR2X2_HVT U1133 ( .A1(n1057), .A2(n1347), .Y(n478) );
  XNOR2X2_HVT U1134 ( .A1(n515), .A2(n1060), .Y(n547) );
  XNOR2X2_HVT U1135 ( .A1(n558), .A2(n47), .Y(n548) );
  XOR3X2_HVT U1136 ( .A1(n727), .A2(n1055), .A3(n439), .Y(n113) );
  XOR2X2_HVT U1137 ( .A1(n513), .A2(n1336), .Y(n499) );
  XNOR2X2_HVT U1138 ( .A1(in[115]), .A2(n1376), .Y(n513) );
  XOR3X2_HVT U1139 ( .A1(n581), .A2(n1242), .A3(n69), .Y(n608) );
  XOR3X2_HVT U1140 ( .A1(n471), .A2(n1089), .A3(n376), .Y(n1325) );
  XNOR2X2_HVT U1141 ( .A1(n465), .A2(n986), .Y(n434) );
  IBUFFX2_HVT U1142 ( .A(n468), .Y(n1058) );
  XOR3X1_HVT U1143 ( .A1(n687), .A2(n469), .A3(n536), .Y(out1[11]) );
  INVX1_HVT U1144 ( .A(n1058), .Y(n1059) );
  INVX1_HVT U1145 ( .A(in[125]), .Y(n1228) );
  XNOR2X2_HVT U1146 ( .A1(in[16]), .A2(n1296), .Y(n439) );
  XOR3X2_HVT U1147 ( .A1(n1139), .A2(n1061), .A3(n404), .Y(n594) );
  INVX1_HVT U1148 ( .A(n433), .Y(n1093) );
  XNOR2X2_HVT U1149 ( .A1(n430), .A2(n1129), .Y(n423) );
  XOR3X1_HVT U1150 ( .A1(n1287), .A2(n460), .A3(n461), .Y(out1[1]) );
  XNOR2X2_HVT U1151 ( .A1(n1090), .A2(in[23]), .Y(n468) );
  XNOR2X2_HVT U1152 ( .A1(n136), .A2(n86), .Y(n191) );
  XNOR2X2_HVT U1153 ( .A1(n103), .A2(n1333), .Y(n98) );
  XNOR2X2_HVT U1154 ( .A1(in[72]), .A2(in[79]), .Y(n1163) );
  NAND2X0_HVT U1155 ( .A1(n1067), .A2(in[89]), .Y(n1068) );
  NAND2X0_HVT U1156 ( .A1(n1066), .A2(n1329), .Y(n1069) );
  NAND2X0_HVT U1157 ( .A1(n1069), .A2(n1068), .Y(n201) );
  INVX1_HVT U1158 ( .A(n531), .Y(n1186) );
  XNOR2X2_HVT U1159 ( .A1(n582), .A2(n1071), .Y(n531) );
  XNOR2X2_HVT U1160 ( .A1(n514), .A2(n1233), .Y(n551) );
  XNOR2X2_HVT U1161 ( .A1(n311), .A2(n1080), .Y(n252) );
  IBUFFX2_HVT U1162 ( .A(in[57]), .Y(n1207) );
  NBUFFX2_HVT U1163 ( .A(n627), .Y(n1071) );
  NBUFFX2_HVT U1164 ( .A(in[9]), .Y(n1072) );
  NBUFFX2_HVT U1165 ( .A(in[112]), .Y(n1073) );
  XOR2X2_HVT U1166 ( .A1(n563), .A2(n782), .Y(n514) );
  XNOR2X2_HVT U1167 ( .A1(in[17]), .A2(n1202), .Y(n473) );
  NAND2X0_HVT U1168 ( .A1(n1078), .A2(n1079), .Y(n1075) );
  NAND2X0_HVT U1169 ( .A1(in[41]), .A2(n1077), .Y(n1078) );
  NAND2X0_HVT U1170 ( .A1(n1076), .A2(n638), .Y(n1079) );
  NAND2X0_HVT U1171 ( .A1(n1078), .A2(n1079), .Y(n362) );
  INVX0_HVT U1172 ( .A(in[41]), .Y(n1076) );
  XNOR3X2_HVT U1173 ( .A1(n148), .A2(n149), .A3(n646), .Y(n1319) );
  INVX1_HVT U1174 ( .A(n1081), .Y(n1082) );
  NBUFFX2_HVT U1175 ( .A(in[41]), .Y(n1084) );
  INVX1_HVT U1176 ( .A(in[12]), .Y(n1344) );
  INVX0_HVT U1177 ( .A(in[12]), .Y(n1218) );
  XOR3X2_HVT U1178 ( .A1(n1257), .A2(n443), .A3(n394), .Y(n1088) );
  XNOR2X2_HVT U1179 ( .A1(in[8]), .A2(n1346), .Y(n50) );
  XNOR2X2_HVT U1180 ( .A1(in[11]), .A2(n1097), .Y(n448) );
  XNOR2X1_HVT U1181 ( .A1(n556), .A2(n463), .Y(n406) );
  INVX1_HVT U1182 ( .A(n518), .Y(n1196) );
  INVX1_HVT U1183 ( .A(n528), .Y(n1189) );
  XOR3X2_HVT U1184 ( .A1(n613), .A2(n1092), .A3(n597), .Y(out1[101]) );
  XOR3X2_HVT U1185 ( .A1(n55), .A2(n1093), .A3(n434), .Y(n432) );
  XOR3X2_HVT U1186 ( .A1(n47), .A2(n691), .A3(n504), .Y(n1096) );
  IBUFFX2_HVT U1187 ( .A(n600), .Y(n1220) );
  XOR2X2_HVT U1188 ( .A1(n444), .A2(n178), .Y(n394) );
  NBUFFX2_HVT U1189 ( .A(in[15]), .Y(n1097) );
  INVX1_HVT U1190 ( .A(n426), .Y(n1276) );
  XNOR2X2_HVT U1191 ( .A1(n470), .A2(n1098), .Y(n378) );
  XNOR3X1_HVT U1192 ( .A1(n1158), .A2(n906), .A3(n303), .Y(n384) );
  INVX1_HVT U1193 ( .A(n1187), .Y(n1099) );
  XOR3X2_HVT U1194 ( .A1(n1100), .A2(n1196), .A3(n519), .Y(out1[123]) );
  XNOR2X2_HVT U1195 ( .A1(in[2]), .A2(n1193), .Y(n489) );
  NBUFFX2_HVT U1196 ( .A(in[98]), .Y(n1101) );
  INVX1_HVT U1197 ( .A(n1241), .Y(n1102) );
  INVX1_HVT U1198 ( .A(in[100]), .Y(n1241) );
  INVX1_HVT U1199 ( .A(n1340), .Y(n1204) );
  XNOR2X2_HVT U1200 ( .A1(n219), .A2(n1218), .Y(n1103) );
  XNOR2X2_HVT U1201 ( .A1(n1151), .A2(in[20]), .Y(n219) );
  INVX2_HVT U1202 ( .A(in[28]), .Y(n1348) );
  IBUFFX2_HVT U1203 ( .A(n416), .Y(n1105) );
  INVX1_HVT U1204 ( .A(n1105), .Y(n1106) );
  XOR3X2_HVT U1205 ( .A1(n210), .A2(n1111), .A3(n120), .Y(n207) );
  XNOR2X2_HVT U1206 ( .A1(n410), .A2(n452), .Y(n259) );
  XOR3X2_HVT U1207 ( .A1(n67), .A2(n1112), .A3(n69), .Y(out1[97]) );
  XNOR2X2_HVT U1208 ( .A1(n583), .A2(n1191), .Y(n566) );
  XNOR2X2_HVT U1209 ( .A1(n600), .A2(n1114), .Y(n1113) );
  XOR2X2_HVT U1210 ( .A1(n435), .A2(n428), .Y(n55) );
  NBUFFX2_HVT U1211 ( .A(in[119]), .Y(n1115) );
  XNOR2X2_HVT U1212 ( .A1(n374), .A2(n1125), .Y(n469) );
  XNOR2X1_HVT U1213 ( .A1(n1341), .A2(n795), .Y(n179) );
  XNOR2X2_HVT U1214 ( .A1(n567), .A2(in[115]), .Y(n521) );
  NBUFFX2_HVT U1215 ( .A(in[103]), .Y(n1116) );
  INVX1_HVT U1216 ( .A(in[87]), .Y(n1366) );
  XNOR2X2_HVT U1217 ( .A1(n154), .A2(n1118), .Y(n101) );
  IBUFFX2_HVT U1218 ( .A(in[83]), .Y(n1117) );
  INVX1_HVT U1219 ( .A(n1117), .Y(n1118) );
  XOR2X2_HVT U1220 ( .A1(n125), .A2(n77), .Y(n183) );
  XNOR2X2_HVT U1221 ( .A1(n1364), .A2(n1201), .Y(n77) );
  XOR3X2_HVT U1222 ( .A1(n122), .A2(n1261), .A3(n174), .Y(n212) );
  XOR3X2_HVT U1223 ( .A1(n367), .A2(n689), .A3(n368), .Y(out1[41]) );
  XOR3X2_HVT U1224 ( .A1(n1121), .A2(n116), .A3(n117), .Y(out1[89]) );
  XOR3X2_HVT U1225 ( .A1(n118), .A2(n119), .A3(n120), .Y(n1121) );
  XOR3X2_HVT U1226 ( .A1(n48), .A2(n109), .A3(n110), .Y(n106) );
  IBUFFX2_HVT U1227 ( .A(in[97]), .Y(n1122) );
  INVX1_HVT U1228 ( .A(n1122), .Y(n1123) );
  XOR3X2_HVT U1229 ( .A1(n104), .A2(n853), .A3(n105), .Y(n100) );
  INVX1_HVT U1230 ( .A(n1370), .Y(n1124) );
  IBUFFX2_HVT U1231 ( .A(n543), .Y(n1234) );
  INVX1_HVT U1232 ( .A(n1126), .Y(n1127) );
  INVX1_HVT U1233 ( .A(in[6]), .Y(n1187) );
  OR2X1_HVT U1234 ( .A1(n830), .A2(n456), .Y(n1288) );
  XOR3X2_HVT U1235 ( .A1(n718), .A2(n181), .A3(n182), .Y(n180) );
  XNOR2X2_HVT U1236 ( .A1(n463), .A2(n794), .Y(n374) );
  XNOR2X2_HVT U1237 ( .A1(n557), .A2(n1130), .Y(n512) );
  XOR3X2_HVT U1238 ( .A1(n349), .A2(n1133), .A3(n351), .Y(out1[45]) );
  XNOR2X2_HVT U1239 ( .A1(in[35]), .A2(n1352), .Y(n348) );
  XNOR2X1_HVT U1240 ( .A1(n930), .A2(n1350), .Y(n342) );
  XOR2X2_HVT U1241 ( .A1(n285), .A2(n286), .Y(n236) );
  XOR3X2_HVT U1242 ( .A1(n562), .A2(n633), .A3(n519), .Y(out1[115]) );
  INVX1_HVT U1243 ( .A(n1138), .Y(n1139) );
  XOR3X2_HVT U1244 ( .A1(n405), .A2(n986), .A3(n477), .Y(n427) );
  XNOR2X2_HVT U1245 ( .A1(n602), .A2(n1102), .Y(n557) );
  INVX1_HVT U1246 ( .A(n573), .Y(n1225) );
  XNOR2X2_HVT U1247 ( .A1(n417), .A2(n1146), .Y(n255) );
  XNOR2X2_HVT U1248 ( .A1(n492), .A2(n1145), .Y(n457) );
  XNOR2X2_HVT U1249 ( .A1(in[99]), .A2(n1371), .Y(n593) );
  XOR3X2_HVT U1250 ( .A1(n1375), .A2(n495), .A3(n502), .Y(n501) );
  XNOR2X2_HVT U1251 ( .A1(n328), .A2(n1140), .Y(n451) );
  NAND2X0_HVT U1252 ( .A1(in[65]), .A2(n1119), .Y(n1142) );
  NAND2X0_HVT U1253 ( .A1(n1291), .A2(n1141), .Y(n1143) );
  XOR2X2_HVT U1254 ( .A1(n1295), .A2(n1188), .Y(n181) );
  INVX1_HVT U1255 ( .A(n1187), .Y(n1188) );
  XNOR2X2_HVT U1256 ( .A1(in[90]), .A2(n1369), .Y(n103) );
  NBUFFX2_HVT U1257 ( .A(n457), .Y(n1144) );
  NBUFFX2_HVT U1258 ( .A(in[13]), .Y(n1145) );
  NBUFFX2_HVT U1259 ( .A(in[13]), .Y(n1146) );
  INVX1_HVT U1260 ( .A(n221), .Y(n1167) );
  NAND2X0_HVT U1261 ( .A1(n1323), .A2(n453), .Y(n1149) );
  NAND2X0_HVT U1262 ( .A1(n1147), .A2(n1148), .Y(n1150) );
  NAND2X0_HVT U1263 ( .A1(n1149), .A2(n1150), .Y(out1[20]) );
  INVX0_HVT U1264 ( .A(n1323), .Y(n1147) );
  INVX0_HVT U1265 ( .A(n453), .Y(n1148) );
  XNOR2X2_HVT U1266 ( .A1(in[3]), .A2(n1343), .Y(n1151) );
  INVX0_HVT U1267 ( .A(n1341), .Y(n1269) );
  INVX2_HVT U1268 ( .A(in[4]), .Y(n1341) );
  XNOR2X2_HVT U1269 ( .A1(n50), .A2(n1146), .Y(n470) );
  NAND2X0_HVT U1270 ( .A1(n413), .A2(n1154), .Y(n1155) );
  NAND2X0_HVT U1271 ( .A1(n1153), .A2(n412), .Y(n1156) );
  NAND2X0_HVT U1272 ( .A1(n1155), .A2(n1156), .Y(out1[28]) );
  INVX0_HVT U1273 ( .A(n412), .Y(n1154) );
  NAND2X0_HVT U1274 ( .A1(n1203), .A2(n490), .Y(n1159) );
  NAND2X0_HVT U1275 ( .A1(n1160), .A2(n1159), .Y(out1[12]) );
  NBUFFX2_HVT U1276 ( .A(n324), .Y(n1161) );
  XNOR2X2_HVT U1277 ( .A1(n361), .A2(n876), .Y(n248) );
  INVX1_HVT U1278 ( .A(n172), .Y(n1173) );
  XNOR2X2_HVT U1279 ( .A1(n194), .A2(n1162), .Y(n145) );
  XOR3X2_HVT U1280 ( .A1(n168), .A2(n1111), .A3(n117), .Y(n167) );
  XNOR2X1_HVT U1281 ( .A1(n147), .A2(n1211), .Y(n86) );
  IBUFFX2_HVT U1282 ( .A(in[82]), .Y(n1164) );
  NAND2X0_HVT U1283 ( .A1(n957), .A2(n1214), .Y(n1166) );
  XOR3X2_HVT U1284 ( .A1(n1168), .A2(n272), .A3(n273), .Y(out1[57]) );
  NAND2X0_HVT U1285 ( .A1(n334), .A2(n875), .Y(n1171) );
  NAND2X0_HVT U1286 ( .A1(n1170), .A2(n1332), .Y(n1172) );
  NAND2X0_HVT U1287 ( .A1(n1171), .A2(n1172), .Y(n360) );
  XOR3X2_HVT U1288 ( .A1(n420), .A2(n687), .A3(n422), .Y(out1[27]) );
  XOR3X2_HVT U1289 ( .A1(n1207), .A2(n269), .A3(n270), .Y(n266) );
  NAND2X0_HVT U1290 ( .A1(n1288), .A2(n1289), .Y(n1174) );
  XNOR2X2_HVT U1291 ( .A1(n354), .A2(n1260), .Y(n301) );
  XOR3X1_HVT U1292 ( .A1(n690), .A2(n316), .A3(n317), .Y(out1[50]) );
  XOR3X2_HVT U1293 ( .A1(n137), .A2(n1212), .A3(n95), .Y(n143) );
  XNOR2X2_HVT U1294 ( .A1(in[0]), .A2(n1193), .Y(n463) );
  XNOR2X2_HVT U1295 ( .A1(in[42]), .A2(n1209), .Y(n311) );
  NAND2X0_HVT U1296 ( .A1(n1327), .A2(n222), .Y(n1177) );
  NAND2X0_HVT U1297 ( .A1(n1175), .A2(n1176), .Y(n1178) );
  NAND2X0_HVT U1298 ( .A1(n1178), .A2(n1177), .Y(out1[68]) );
  INVX0_HVT U1299 ( .A(n222), .Y(n1176) );
  XOR2X2_HVT U1300 ( .A1(n130), .A2(n129), .Y(n81) );
  XOR3X1_HVT U1301 ( .A1(n1181), .A2(n1182), .A3(n1183), .Y(out1[62]) );
  XNOR2X2_HVT U1302 ( .A1(in[104]), .A2(n635), .Y(n583) );
  XNOR2X2_HVT U1303 ( .A1(n639), .A2(n1215), .Y(n366) );
  XNOR2X2_HVT U1304 ( .A1(n1227), .A2(n1184), .Y(n516) );
  XOR3X1_HVT U1305 ( .A1(n1189), .A2(n580), .A3(n608), .Y(out1[105]) );
  XNOR2X2_HVT U1306 ( .A1(n97), .A2(n1307), .Y(n140) );
  XNOR2X2_HVT U1307 ( .A1(in[67]), .A2(n916), .Y(n188) );
  XOR2X2_HVT U1308 ( .A1(n131), .A2(n82), .Y(n186) );
  INVX1_HVT U1309 ( .A(n1233), .Y(n1191) );
  XNOR2X2_HVT U1310 ( .A1(in[121]), .A2(in[126]), .Y(n605) );
  XOR3X2_HVT U1311 ( .A1(n449), .A2(n1195), .A3(n1018), .Y(out1[21]) );
  INVX1_HVT U1312 ( .A(n86), .Y(n1262) );
  XOR3X1_HVT U1313 ( .A1(n1196), .A2(n935), .A3(n1197), .Y(out1[107]) );
  XNOR2X2_HVT U1314 ( .A1(n134), .A2(n135), .Y(n85) );
  XNOR2X2_HVT U1315 ( .A1(in[112]), .A2(n1376), .Y(n576) );
  XOR3X2_HVT U1316 ( .A1(n170), .A2(n1042), .A3(n209), .Y(n230) );
  XOR3X2_HVT U1317 ( .A1(n1198), .A2(n190), .A3(n191), .Y(out1[77]) );
  XNOR2X2_HVT U1318 ( .A1(n327), .A2(n1296), .Y(n410) );
  NBUFFX2_HVT U1319 ( .A(n1362), .Y(n1199) );
  IBUFFX2_HVT U1320 ( .A(in[87]), .Y(n1200) );
  INVX1_HVT U1321 ( .A(n1200), .Y(n1201) );
  IBUFFX2_HVT U1322 ( .A(n194), .Y(n1304) );
  XNOR2X2_HVT U1323 ( .A1(in[56]), .A2(n1014), .Y(n274) );
  INVX1_HVT U1324 ( .A(n256), .Y(n1283) );
  XNOR2X2_HVT U1325 ( .A1(in[82]), .A2(n1366), .Y(n157) );
  XOR3X2_HVT U1326 ( .A1(n456), .A2(n1144), .A3(n487), .Y(n1203) );
  XNOR2X2_HVT U1327 ( .A1(n489), .A2(n1188), .Y(n328) );
  XOR3X2_HVT U1328 ( .A1(n476), .A2(n1204), .A3(n429), .Y(n404) );
  XOR3X2_HVT U1329 ( .A1(n365), .A2(n1207), .A3(n319), .Y(n391) );
  NBUFFX2_HVT U1330 ( .A(in[85]), .Y(n1210) );
  NBUFFX2_HVT U1331 ( .A(in[85]), .Y(n1211) );
  NAND2X0_HVT U1332 ( .A1(n1212), .A2(n94), .Y(n1214) );
  NAND2X0_HVT U1333 ( .A1(n1214), .A2(n957), .Y(n195) );
  XNOR2X2_HVT U1334 ( .A1(in[83]), .A2(n1366), .Y(n96) );
  XNOR2X2_HVT U1335 ( .A1(n171), .A2(n1210), .Y(n154) );
  XOR3X2_HVT U1336 ( .A1(n116), .A2(n1217), .A3(n166), .Y(n208) );
  XNOR2X2_HVT U1337 ( .A1(n150), .A2(in[84]), .Y(n94) );
  XOR2X2_HVT U1338 ( .A1(n542), .A2(n499), .Y(n591) );
  INVX1_HVT U1339 ( .A(n20), .Y(n1221) );
  NAND2X0_HVT U1340 ( .A1(n246), .A2(n1251), .Y(n1223) );
  NAND2X0_HVT U1341 ( .A1(n926), .A2(n1222), .Y(n1224) );
  NAND2X0_HVT U1342 ( .A1(n1223), .A2(n1224), .Y(out1[60]) );
  XNOR2X2_HVT U1343 ( .A1(n155), .A2(n1192), .Y(n97) );
  INVX1_HVT U1344 ( .A(n567), .Y(n1245) );
  XNOR2X2_HVT U1345 ( .A1(n576), .A2(n1375), .Y(n567) );
  XNOR2X2_HVT U1346 ( .A1(n1239), .A2(n1337), .Y(n333) );
  XOR2X2_HVT U1347 ( .A1(n251), .A2(n1338), .Y(n237) );
  XNOR2X2_HVT U1348 ( .A1(n264), .A2(n322), .Y(n308) );
  INVX1_HVT U1349 ( .A(in[55]), .Y(n1356) );
  XOR3X2_HVT U1350 ( .A1(n382), .A2(n1248), .A3(n351), .Y(out1[37]) );
  INVX1_HVT U1351 ( .A(n57), .Y(n1277) );
  XNOR2X2_HVT U1352 ( .A1(n577), .A2(n1230), .Y(n57) );
  XNOR2X2_HVT U1353 ( .A1(n593), .A2(n620), .Y(n546) );
  INVX1_HVT U1354 ( .A(n1232), .Y(n1230) );
  XNOR2X1_HVT U1355 ( .A1(n1230), .A2(n648), .Y(n586) );
  XOR3X2_HVT U1356 ( .A1(n546), .A2(n1232), .A3(n506), .Y(n592) );
  XNOR2X2_HVT U1357 ( .A1(n1297), .A2(n1116), .Y(n63) );
  XOR3X2_HVT U1358 ( .A1(n267), .A2(n1235), .A3(n316), .Y(n364) );
  XNOR2X2_HVT U1359 ( .A1(n336), .A2(n1240), .Y(n310) );
  IBUFFX2_HVT U1360 ( .A(in[48]), .Y(n1236) );
  INVX1_HVT U1361 ( .A(n1236), .Y(n1237) );
  INVX1_HVT U1362 ( .A(n1238), .Y(n1240) );
  XNOR2X2_HVT U1363 ( .A1(in[48]), .A2(n1356), .Y(n336) );
  XNOR2X2_HVT U1364 ( .A1(n1247), .A2(in[51]), .Y(n251) );
  XOR3X2_HVT U1365 ( .A1(n216), .A2(n797), .A3(n225), .Y(n1243) );
  XOR3X2_HVT U1366 ( .A1(n1245), .A2(n60), .A3(n660), .Y(n562) );
  XNOR2X2_HVT U1367 ( .A1(n933), .A2(n459), .Y(n431) );
  XNOR2X2_HVT U1368 ( .A1(n462), .A2(n1340), .Y(n53) );
  XNOR2X2_HVT U1369 ( .A1(n255), .A2(n451), .Y(n411) );
  INVX1_HVT U1370 ( .A(n330), .Y(n1256) );
  XOR2X2_HVT U1371 ( .A1(n1352), .A2(n765), .Y(n365) );
  XNOR2X2_HVT U1372 ( .A1(n569), .A2(n570), .Y(n60) );
  NBUFFX2_HVT U1373 ( .A(n251), .Y(n1249) );
  XOR3X2_HVT U1374 ( .A1(n369), .A2(n826), .A3(n632), .Y(n1250) );
  XOR3X2_HVT U1375 ( .A1(n561), .A2(n491), .A3(n35), .Y(n1252) );
  XNOR2X2_HVT U1376 ( .A1(n290), .A2(n291), .Y(n240) );
  INVX1_HVT U1377 ( .A(n746), .Y(n1254) );
  XNOR2X2_HVT U1378 ( .A1(n356), .A2(n277), .Y(n302) );
  XNOR2X2_HVT U1379 ( .A1(in[10]), .A2(n833), .Y(n472) );
  XOR3X1_HVT U1380 ( .A1(n1256), .A2(n331), .A3(n332), .Y(out1[49]) );
  INVX1_HVT U1381 ( .A(n1258), .Y(n1259) );
  XNOR2X2_HVT U1382 ( .A1(n305), .A2(n1135), .Y(n297) );
  XOR3X2_HVT U1383 ( .A1(n71), .A2(n576), .A3(n580), .Y(n529) );
  XNOR2X2_HVT U1384 ( .A1(n581), .A2(n1372), .Y(n71) );
  IBUFFX2_HVT U1385 ( .A(n459), .Y(n1287) );
  XNOR2X2_HVT U1386 ( .A1(n292), .A2(n241), .Y(n351) );
  XOR2X2_HVT U1387 ( .A1(n287), .A2(n237), .Y(n346) );
  XOR3X2_HVT U1388 ( .A1(n312), .A2(n313), .A3(n314), .Y(n262) );
  XNOR2X2_HVT U1389 ( .A1(in[50]), .A2(n1247), .Y(n313) );
  XOR3X2_HVT U1390 ( .A1(n405), .A2(in[25]), .A3(n406), .Y(n402) );
  XNOR2X2_HVT U1391 ( .A1(in[32]), .A2(n1246), .Y(n390) );
  XNOR2X2_HVT U1392 ( .A1(n248), .A2(n1357), .Y(n300) );
  XOR2X2_HVT U1393 ( .A1(n54), .A2(n1072), .Y(n459) );
  XOR3X2_HVT U1394 ( .A1(n1265), .A2(n596), .A3(n597), .Y(out1[109]) );
  XNOR2X2_HVT U1395 ( .A1(n545), .A2(n546), .Y(n502) );
  XNOR2X2_HVT U1396 ( .A1(n263), .A2(n1305), .Y(n253) );
  INVX1_HVT U1397 ( .A(n1347), .Y(n1267) );
  INVX2_HVT U1398 ( .A(in[22]), .Y(n1347) );
  XNOR2X2_HVT U1399 ( .A1(n599), .A2(n1320), .Y(out1[108]) );
  INVX1_HVT U1400 ( .A(n1272), .Y(n1273) );
  XOR3X1_HVT U1401 ( .A1(n1276), .A2(n477), .A3(n594), .Y(out1[10]) );
  NBUFFX2_HVT U1402 ( .A(in[31]), .Y(n1280) );
  XOR3X2_HVT U1403 ( .A1(n706), .A2(n223), .A3(n265), .Y(n260) );
  XNOR2X2_HVT U1404 ( .A1(in[105]), .A2(n696), .Y(n606) );
  XNOR2X2_HVT U1405 ( .A1(n473), .A2(n1295), .Y(n455) );
  NAND2X0_HVT U1406 ( .A1(n456), .A2(n830), .Y(n1289) );
  NAND2X0_HVT U1407 ( .A1(n1289), .A2(n1288), .Y(n415) );
  XNOR2X2_HVT U1408 ( .A1(n387), .A2(n950), .Y(n305) );
  XNOR2X2_HVT U1409 ( .A1(n419), .A2(n1348), .Y(n458) );
  XOR3X2_HVT U1410 ( .A1(n802), .A2(n1326), .A3(n51), .Y(out1[9]) );
  XNOR2X2_HVT U1411 ( .A1(n472), .A2(n1257), .Y(n417) );
  XOR2X2_HVT U1412 ( .A1(n479), .A2(n1296), .Y(n471) );
  XNOR2X2_HVT U1413 ( .A1(n468), .A2(n1267), .Y(n327) );
  XOR3X2_HVT U1414 ( .A1(n469), .A2(n1059), .A3(n701), .Y(n422) );
  XNOR2X2_HVT U1415 ( .A1(n313), .A2(n1338), .Y(n303) );
  XOR3X2_HVT U1416 ( .A1(n526), .A2(n1123), .A3(n572), .Y(n64) );
  XNOR2X2_HVT U1417 ( .A1(n561), .A2(in[116]), .Y(n511) );
  NBUFFX2_HVT U1418 ( .A(in[21]), .Y(n1295) );
  NBUFFX2_HVT U1419 ( .A(in[21]), .Y(n1296) );
  XNOR2X2_HVT U1420 ( .A1(n471), .A2(n883), .Y(n424) );
  XNOR2X2_HVT U1421 ( .A1(n606), .A2(n1373), .Y(n600) );
  INVX1_HVT U1422 ( .A(n1297), .Y(n1298) );
  XNOR2X2_HVT U1423 ( .A1(n228), .A2(n1359), .Y(n199) );
  XNOR2X2_HVT U1424 ( .A1(in[64]), .A2(n1361), .Y(n228) );
  XNOR2X2_HVT U1425 ( .A1(n458), .A2(n414), .Y(n325) );
  XNOR2X2_HVT U1426 ( .A1(in[1]), .A2(n1187), .Y(n474) );
  NAND2X0_HVT U1427 ( .A1(n1301), .A2(n1313), .Y(n1302) );
  NAND2X0_HVT U1428 ( .A1(n193), .A2(n1300), .Y(n1303) );
  NAND2X0_HVT U1429 ( .A1(n1303), .A2(n1302), .Y(out1[76]) );
  INVX0_HVT U1430 ( .A(n1313), .Y(n1300) );
  XOR3X2_HVT U1431 ( .A1(n98), .A2(n45), .A3(n694), .Y(n1313) );
  NBUFFX2_HVT U1432 ( .A(in[62]), .Y(n1305) );
  NBUFFX2_HVT U1433 ( .A(in[62]), .Y(n1306) );
  XNOR2X2_HVT U1434 ( .A1(n202), .A2(n1307), .Y(n194) );
  XNOR2X2_HVT U1435 ( .A1(n157), .A2(n1334), .Y(n147) );
  XNOR2X2_HVT U1436 ( .A1(n757), .A2(n1292), .Y(n149) );
  XNOR2X2_HVT U1437 ( .A1(n324), .A2(n1341), .Y(n456) );
  XNOR2X2_HVT U1438 ( .A1(in[97]), .A2(in[102]), .Y(n569) );
  XNOR2X2_HVT U1439 ( .A1(n564), .A2(n734), .Y(n558) );
  XNOR2X2_HVT U1440 ( .A1(in[114]), .A2(n1376), .Y(n564) );
  XOR2X2_HVT U1441 ( .A1(in[23]), .A2(in[16]), .Y(n479) );
  XNOR2X2_HVT U1442 ( .A1(n99), .A2(in[76]), .Y(n83) );
  XOR3X1_HVT U1443 ( .A1(n688), .A2(n1309), .A3(n1310), .Y(out1[83]) );
  XNOR2X2_HVT U1444 ( .A1(n146), .A2(n145), .Y(n95) );
  XNOR2X1_HVT U1445 ( .A1(n348), .A2(n1354), .Y(n295) );
  XOR2X1_HVT U1446 ( .A1(n365), .A2(n318), .Y(n330) );
  XNOR2X1_HVT U1447 ( .A1(n188), .A2(n1364), .Y(n139) );
  XOR2X1_HVT U1448 ( .A1(n1062), .A2(n50), .Y(n426) );
  XNOR2X1_HVT U1449 ( .A1(n1360), .A2(n1365), .Y(n173) );
  XNOR2X1_HVT U1450 ( .A1(n651), .A2(n1254), .Y(n307) );
  XNOR2X1_HVT U1451 ( .A1(n1351), .A2(n1355), .Y(n338) );
  XNOR2X1_HVT U1452 ( .A1(n73), .A2(n1), .Y(n518) );
  XNOR2X1_HVT U1453 ( .A1(n20), .A2(n583), .Y(n523) );
  XNOR3X1_HVT U1454 ( .A1(n1322), .A2(n399), .A3(n400), .Y(out1[30]) );
  XNOR2X1_HVT U1455 ( .A1(in[29]), .A2(in[24]), .Y(n483) );
  XNOR2X1_HVT U1456 ( .A1(n1364), .A2(n1211), .Y(n126) );
  XNOR2X1_HVT U1457 ( .A1(n1354), .A2(n1240), .Y(n282) );
  XOR3X1_HVT U1458 ( .A1(n111), .A2(n112), .A3(n113), .Y(out1[8]) );
  XNOR3X1_HVT U1459 ( .A1(n129), .A2(n1333), .A3(n173), .Y(n214) );
  XNOR2X1_HVT U1460 ( .A1(n1344), .A2(n1097), .Y(n178) );
  XNOR2X1_HVT U1461 ( .A1(n1374), .A2(n1115), .Y(n494) );
  XNOR2X1_HVT U1462 ( .A1(n1345), .A2(n695), .Y(n437) );
  XNOR2X1_HVT U1463 ( .A1(n277), .A2(n1135), .Y(n379) );
  XNOR2X1_HVT U1464 ( .A1(n1374), .A2(n1041), .Y(n538) );
  XNOR2X1_HVT U1465 ( .A1(n917), .A2(n1359), .Y(n213) );
  XNOR3X1_HVT U1466 ( .A1(n1335), .A2(n80), .A3(n81), .Y(n79) );
  XNOR3X1_HVT U1467 ( .A1(n1330), .A2(n74), .A3(n75), .Y(out1[96]) );
  XNOR3X1_HVT U1468 ( .A1(n540), .A2(n1312), .A3(n585), .Y(n1331) );
  XNOR2X1_HVT U1469 ( .A1(n448), .A2(in[28]), .Y(n407) );
  XNOR2X1_HVT U1470 ( .A1(n254), .A2(n1305), .Y(n287) );
  XOR2X1_HVT U1471 ( .A1(n269), .A2(in[58]), .Y(n316) );
  XNOR2X1_HVT U1472 ( .A1(n1124), .A2(n1297), .Y(n68) );
  XNOR2X1_HVT U1473 ( .A1(n1332), .A2(n1306), .Y(n235) );
  XNOR2X1_HVT U1474 ( .A1(n559), .A2(in[124]), .Y(n506) );
  XNOR2X1_HVT U1475 ( .A1(n148), .A2(in[92]), .Y(n89) );
  XOR2X1_HVT U1476 ( .A1(in[76]), .A2(n1194), .Y(n184) );
  XOR2X1_HVT U1477 ( .A1(n403), .A2(n1127), .Y(n477) );
  XNOR2X1_HVT U1478 ( .A1(n1132), .A2(n1342), .Y(n403) );
  XNOR2X1_HVT U1479 ( .A1(in[104]), .A2(n1233), .Y(n74) );
  XNOR2X1_HVT U1480 ( .A1(n1378), .A2(n1060), .Y(n495) );
  XNOR2X1_HVT U1481 ( .A1(n629), .A2(in[120]), .Y(n587) );
  XNOR2X1_HVT U1482 ( .A1(in[108]), .A2(n1259), .Y(n540) );
  XNOR2X1_HVT U1483 ( .A1(in[44]), .A2(n1215), .Y(n285) );
  XNOR2X1_HVT U1484 ( .A1(in[60]), .A2(n1109), .Y(n281) );
  XNOR2X1_HVT U1485 ( .A1(in[124]), .A2(n1227), .Y(n537) );
  XNOR2X1_HVT U1486 ( .A1(in[76]), .A2(n798), .Y(n129) );
  XNOR2X1_HVT U1487 ( .A1(n1367), .A2(n959), .Y(n78) );
  XNOR2X1_HVT U1488 ( .A1(n1357), .A2(n876), .Y(n233) );
  XNOR2X1_HVT U1489 ( .A1(n1102), .A2(n1230), .Y(n610) );
  XNOR2X1_HVT U1490 ( .A1(in[88]), .A2(n959), .Y(n174) );
  XOR2X1_HVT U1491 ( .A1(in[44]), .A2(n945), .Y(n344) );
  XNOR2X1_HVT U1492 ( .A1(n1347), .A2(n795), .Y(n440) );
  XNOR2X1_HVT U1493 ( .A1(n1298), .A2(n1375), .Y(n585) );
  XNOR2X1_HVT U1494 ( .A1(in[20]), .A2(n1057), .Y(n397) );
  XOR2X1_HVT U1495 ( .A1(in[20]), .A2(n1296), .Y(n441) );
  XNOR2X1_HVT U1496 ( .A1(n1344), .A2(in[13]), .Y(n484) );
  XNOR2X1_HVT U1497 ( .A1(n1145), .A2(n718), .Y(n114) );
  XNOR2X1_HVT U1498 ( .A1(in[4]), .A2(n727), .Y(n444) );
  NBUFFX2_HVT U1499 ( .A(in[45]), .Y(n1332) );
  NBUFFX2_HVT U1500 ( .A(in[94]), .Y(n1333) );
  NBUFFX2_HVT U1501 ( .A(in[118]), .Y(n1336) );
  NBUFFX2_HVT U1502 ( .A(in[54]), .Y(n1337) );
  NBUFFX2_HVT U1503 ( .A(n1337), .Y(n1338) );
  XNOR2X1_HVT U1504 ( .A1(n1359), .A2(n1334), .Y(n128) );
  INVX0_HVT U1505 ( .A(in[60]), .Y(n1357) );
  INVX0_HVT U1506 ( .A(in[116]), .Y(n1374) );
  INVX0_HVT U1507 ( .A(in[121]), .Y(n1377) );
endmodule

