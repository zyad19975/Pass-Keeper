
module inv_sbox_3 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n91, n196, n197, n198, n199, n200, n201, n202, n203, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655;

  NAND2X0_HVT U1 ( .A1(n251), .A2(n358), .Y(n655) );
  NAND2X0_HVT U5 ( .A1(n367), .A2(n652), .Y(n651) );
  NAND2X0_HVT U6 ( .A1(n376), .A2(n374), .Y(n649) );
  NAND2X0_HVT U9 ( .A1(n374), .A2(n647), .Y(n646) );
  NAND2X0_HVT U10 ( .A1(n373), .A2(n644), .Y(n645) );
  NAND2X0_HVT U12 ( .A1(n375), .A2(n356), .Y(n642) );
  NAND2X0_HVT U13 ( .A1(n370), .A2(n647), .Y(n641) );
  NAND2X0_HVT U15 ( .A1(n338), .A2(n378), .Y(n639) );
  NAND2X0_HVT U19 ( .A1(n377), .A2(n445), .Y(n634) );
  NAND2X0_HVT U25 ( .A1(n270), .A2(n357), .Y(n650) );
  NAND2X0_HVT U32 ( .A1(n223), .A2(n381), .Y(n622) );
  NAND2X0_HVT U35 ( .A1(n647), .A2(n339), .Y(n619) );
  NAND2X0_HVT U38 ( .A1(n356), .A2(n381), .Y(n616) );
  NAND2X0_HVT U42 ( .A1(n649), .A2(n340), .Y(n612) );
  OA21X1_HVT U53 ( .A1(n388), .A2(n604), .A3(n255), .Y(n602) );
  NAND2X0_HVT U55 ( .A1(n652), .A2(n370), .Y(n600) );
  AO21X1_HVT U60 ( .A1(n594), .A2(n354), .A3(n633), .Y(n595) );
  MUX41X1_HVT U65 ( .A1(n405), .A3(n407), .A2(n406), .A4(n616), .S0(n348), 
        .S1(n386), .Y(n589) );
  NAND2X0_HVT U66 ( .A1(n293), .A2(n327), .Y(n588) );
  MUX41X1_HVT U67 ( .A1(n402), .A3(n426), .A2(n404), .A4(n588), .S0(n353), 
        .S1(n345), .Y(n587) );
  MUX41X1_HVT U68 ( .A1(n402), .A3(n323), .A2(n403), .A4(n374), .S0(n347), 
        .S1(n387), .Y(n586) );
  NAND2X0_HVT U72 ( .A1(n335), .A2(n648), .Y(n583) );
  MUX41X1_HVT U73 ( .A1(n627), .A3(n583), .A2(n427), .A4(n355), .S0(n354), 
        .S1(n344), .Y(n582) );
  MUX41X1_HVT U74 ( .A1(n645), .A3(n417), .A2(n416), .A4(n408), .S0(n348), 
        .S1(n309), .Y(n581) );
  MUX41X1_HVT U78 ( .A1(n578), .A3(n582), .A2(n581), .A4(n584), .S0(n364), 
        .S1(n362), .Y(n577) );
  MUX41X1_HVT U79 ( .A1(n413), .A3(n636), .A2(n415), .A4(n637), .S0(n348), 
        .S1(n384), .Y(n576) );
  MUX41X1_HVT U80 ( .A1(n429), .A3(n324), .A2(n646), .A4(n651), .S0(n347), 
        .S1(n385), .Y(n575) );
  NAND2X0_HVT U81 ( .A1(n372), .A2(n648), .Y(n574) );
  AND2X1_HVT U82 ( .A1(n300), .A2(n368), .Y(n573) );
  MUX41X1_HVT U83 ( .A1(n573), .A3(n414), .A2(n272), .A4(n574), .S0(n347), 
        .S1(n268), .Y(n572) );
  MUX41X1_HVT U88 ( .A1(n404), .A3(n391), .A2(n624), .A4(n608), .S0(n347), 
        .S1(n387), .Y(n568) );
  NAND2X0_HVT U89 ( .A1(n381), .A2(n442), .Y(n567) );
  MUX41X1_HVT U98 ( .A1(n560), .A3(n434), .A2(n419), .A4(n626), .S0(n348), 
        .S1(n385), .Y(n559) );
  MUX41X1_HVT U99 ( .A1(n622), .A3(n406), .A2(n606), .A4(n337), .S0(n309), 
        .S1(n345), .Y(n558) );
  MUX41X1_HVT U101 ( .A1(n435), .A3(n642), .A2(n418), .A4(n557), .S0(n309), 
        .S1(n343), .Y(n556) );
  MUX41X1_HVT U102 ( .A1(n556), .A3(n559), .A2(n558), .A4(n561), .S0(n365), 
        .S1(n362), .Y(n555) );
  AND2X1_HVT U104 ( .A1(n648), .A2(n366), .Y(n554) );
  MUX41X1_HVT U105 ( .A1(n640), .A3(n436), .A2(n574), .A4(n554), .S0(n348), 
        .S1(n386), .Y(n553) );
  MUX41X1_HVT U107 ( .A1(n435), .A3(n368), .A2(n552), .A4(n396), .S0(n347), 
        .S1(n385), .Y(n551) );
  MUX41X1_HVT U108 ( .A1(n241), .A3(n338), .A2(n411), .A4(n372), .S0(n348), 
        .S1(n386), .Y(n550) );
  MUX41X1_HVT U109 ( .A1(n434), .A3(n391), .A2(n431), .A4(n424), .S0(n347), 
        .S1(n387), .Y(n549) );
  MUX41X1_HVT U110 ( .A1(n549), .A3(n551), .A2(n550), .A4(n553), .S0(n365), 
        .S1(n362), .Y(n548) );
  AO21X1_HVT U112 ( .A1(n421), .A2(n353), .A3(n630), .Y(n546) );
  NAND2X0_HVT U114 ( .A1(n374), .A2(n648), .Y(n544) );
  MUX41X1_HVT U115 ( .A1(n544), .A3(n643), .A2(n421), .A4(n368), .S0(n309), 
        .S1(n345), .Y(n543) );
  MUX41X1_HVT U116 ( .A1(n420), .A3(n413), .A2(n391), .A4(n639), .S0(n346), 
        .S1(n385), .Y(n542) );
  NAND2X0_HVT U118 ( .A1(n381), .A2(n323), .Y(n540) );
  MUX41X1_HVT U119 ( .A1(n437), .A3(n541), .A2(n617), .A4(n540), .S0(n346), 
        .S1(n385), .Y(n539) );
  MUX41X1_HVT U120 ( .A1(n539), .A3(n543), .A2(n542), .A4(n545), .S0(n365), 
        .S1(n362), .Y(n538) );
  MUX41X1_HVT U122 ( .A1(n425), .A3(n329), .A2(n608), .A4(n428), .S0(n346), 
        .S1(n385), .Y(n537) );
  MUX41X1_HVT U124 ( .A1(n331), .A3(n536), .A2(n631), .A4(n277), .S0(n353), 
        .S1(n346), .Y(n535) );
  AOI21X1_HVT U127 ( .A1(n351), .A2(n531), .A3(n397), .Y(n532) );
  NAND2X0_HVT U129 ( .A1(n350), .A2(n373), .Y(n529) );
  MUX41X1_HVT U130 ( .A1(n529), .A3(n530), .A2(n533), .A4(n532), .S0(n354), 
        .S1(n362), .Y(n528) );
  AND2X1_HVT U131 ( .A1(n327), .A2(n381), .Y(n527) );
  MUX41X1_HVT U132 ( .A1(n306), .A3(n527), .A2(n439), .A4(n402), .S0(n354), 
        .S1(n344), .Y(n526) );
  MUX41X1_HVT U133 ( .A1(n440), .A3(n396), .A2(n600), .A4(n395), .S0(n354), 
        .S1(n343), .Y(n525) );
  MUX41X1_HVT U136 ( .A1(n605), .A3(n557), .A2(n523), .A4(n400), .S0(n350), 
        .S1(n386), .Y(n522) );
  MUX41X1_HVT U137 ( .A1(n647), .A3(n625), .A2(n629), .A4(n433), .S0(n353), 
        .S1(n343), .Y(n521) );
  MUX41X1_HVT U139 ( .A1(n520), .A3(n524), .A2(n528), .A4(n534), .S0(n365), 
        .S1(in[7]), .Y(out[4]) );
  NAND2X0_HVT U141 ( .A1(n338), .A2(n381), .Y(n518) );
  MUX41X1_HVT U142 ( .A1(n518), .A3(n615), .A2(n438), .A4(n410), .S0(n351), 
        .S1(n387), .Y(n517) );
  MUX41X1_HVT U145 ( .A1(n623), .A3(n436), .A2(n515), .A4(n574), .S0(n351), 
        .S1(n386), .Y(n514) );
  MUX41X1_HVT U155 ( .A1(n410), .A3(n643), .A2(n635), .A4(n412), .S0(n349), 
        .S1(n387), .Y(n504) );
  NAND2X0_HVT U159 ( .A1(n500), .A2(n499), .Y(n501) );
  MUX41X1_HVT U162 ( .A1(n422), .A3(n407), .A2(n619), .A4(n497), .S0(n349), 
        .S1(n385), .Y(n496) );
  NAND2X0_HVT U163 ( .A1(n377), .A2(n442), .Y(n495) );
  NAND2X0_HVT U166 ( .A1(n644), .A2(n491), .Y(n492) );
  MUX41X1_HVT U168 ( .A1(n490), .A3(n496), .A2(n494), .A4(n498), .S0(n365), 
        .S1(n361), .Y(n489) );
  MUX41X1_HVT U170 ( .A1(n332), .A3(n328), .A2(n331), .A4(n488), .S0(n349), 
        .S1(n386), .Y(n487) );
  MUX41X1_HVT U172 ( .A1(n567), .A3(n486), .A2(n328), .A4(n632), .S0(n349), 
        .S1(n387), .Y(n485) );
  MUX41X1_HVT U174 ( .A1(n432), .A3(n600), .A2(n440), .A4(n339), .S0(n349), 
        .S1(n384), .Y(n483) );
  NAND2X0_HVT U177 ( .A1(n197), .A2(n323), .Y(n481) );
  AND2X1_HVT U179 ( .A1(n300), .A2(n366), .Y(n479) );
  MUX41X1_HVT U180 ( .A1(n622), .A3(n220), .A2(n479), .A4(n609), .S0(n349), 
        .S1(n385), .Y(n478) );
  MUX41X1_HVT U183 ( .A1(n260), .A3(n324), .A2(n227), .A4(n612), .S0(n353), 
        .S1(n344), .Y(n475) );
  AND2X1_HVT U185 ( .A1(n340), .A2(n91), .Y(n473) );
  NAND2X0_HVT U191 ( .A1(n269), .A2(n401), .Y(n467) );
  AND2X1_HVT U192 ( .A1(n417), .A2(n465), .Y(n466) );
  NAND2X0_HVT U194 ( .A1(n299), .A2(n465), .Y(n463) );
  MUX41X1_HVT U195 ( .A1(n464), .A3(n463), .A2(n466), .A4(n467), .S0(n347), 
        .S1(n361), .Y(n462) );
  NAND2X0_HVT U198 ( .A1(n377), .A2(n339), .Y(n644) );
  NAND2X0_HVT U200 ( .A1(n367), .A2(n381), .Y(n531) );
  NAND2X0_HVT U207 ( .A1(n381), .A2(n444), .Y(n594) );
  INVX8_HVT U2 ( .A(n235), .Y(n565) );
  MUX21X2_HVT U3 ( .A1(n233), .A2(n236), .S0(n237), .Y(n235) );
  INVX2_HVT U4 ( .A(n377), .Y(n381) );
  INVX2_HVT U7 ( .A(n459), .Y(n428) );
  MUX21X1_HVT U8 ( .A1(n562), .A2(n555), .S0(n310), .Y(out[2]) );
  INVX0_HVT U11 ( .A(n367), .Y(n225) );
  INVX1_HVT U14 ( .A(n197), .Y(n91) );
  INVX1_HVT U16 ( .A(n380), .Y(n196) );
  INVX1_HVT U17 ( .A(n380), .Y(n197) );
  XOR2X2_HVT U18 ( .A1(n368), .A2(n293), .Y(n607) );
  IBUFFX2_HVT U20 ( .A(n91), .Y(n237) );
  AO21X2_HVT U21 ( .A1(n91), .A2(n373), .A3(n269), .Y(n499) );
  NAND2X0_HVT U22 ( .A1(n595), .A2(n198), .Y(n199) );
  NAND2X0_HVT U23 ( .A1(n596), .A2(n259), .Y(n200) );
  NAND2X0_HVT U24 ( .A1(n199), .A2(n200), .Y(n593) );
  INVX0_HVT U26 ( .A(n259), .Y(n198) );
  MUX21X1_HVT U27 ( .A1(n600), .A2(n277), .S0(n298), .Y(n596) );
  IBUFFX2_HVT U28 ( .A(n350), .Y(n259) );
  MUX21X1_HVT U29 ( .A1(n356), .A2(n371), .S0(n301), .Y(n277) );
  MUX41X1_HVT U30 ( .A1(n471), .A3(n470), .A2(n472), .A4(n469), .S0(n360), 
        .S1(n343), .Y(n468) );
  NAND2X0_HVT U31 ( .A1(n606), .A2(n201), .Y(n202) );
  NAND2X0_HVT U33 ( .A1(n333), .A2(n219), .Y(n203) );
  NAND2X0_HVT U34 ( .A1(n202), .A2(n203), .Y(n471) );
  INVX0_HVT U36 ( .A(n219), .Y(n201) );
  MUX21X1_HVT U37 ( .A1(n613), .A2(n427), .S0(n264), .Y(n470) );
  IBUFFX2_HVT U39 ( .A(n354), .Y(n219) );
  INVX0_HVT U40 ( .A(n277), .Y(n631) );
  OA21X1_HVT U41 ( .A1(n413), .A2(n388), .A3(n594), .Y(n469) );
  MUX41X1_HVT U43 ( .A1(n567), .A3(n607), .A2(n648), .A4(n238), .S0(n218), 
        .S1(n313), .Y(n566) );
  IBUFFX16_HVT U44 ( .A(n347), .Y(n218) );
  INVX0_HVT U45 ( .A(n196), .Y(n248) );
  INVX1_HVT U46 ( .A(n629), .Y(n410) );
  MUX21X2_HVT U47 ( .A1(n428), .A2(n390), .S0(n352), .Y(n580) );
  XOR2X1_HVT U48 ( .A1(n336), .A2(n196), .Y(n608) );
  INVX1_HVT U49 ( .A(n196), .Y(n301) );
  NOR2X0_HVT U50 ( .A1(n196), .A2(n221), .Y(n220) );
  INVX8_HVT U51 ( .A(n220), .Y(n643) );
  IBUFFX16_HVT U52 ( .A(n372), .Y(n221) );
  NBUFFX2_HVT U54 ( .A(n447), .Y(n222) );
  NBUFFX2_HVT U56 ( .A(n447), .Y(n223) );
  NBUFFX2_HVT U57 ( .A(n447), .Y(n358) );
  INVX0_HVT U58 ( .A(in[6]), .Y(n447) );
  INVX1_HVT U59 ( .A(n223), .Y(n234) );
  INVX0_HVT U61 ( .A(n408), .Y(n240) );
  MUX21X1_HVT U62 ( .A1(n602), .A2(n603), .S0(n320), .Y(n601) );
  INVX0_HVT U63 ( .A(n446), .Y(n338) );
  MUX21X1_HVT U64 ( .A1(n412), .A2(n403), .S0(n352), .Y(n603) );
  INVX1_HVT U69 ( .A(n373), .Y(n444) );
  NOR2X2_HVT U70 ( .A1(n263), .A2(n225), .Y(n224) );
  INVX8_HVT U71 ( .A(n224), .Y(n647) );
  IBUFFX2_HVT U75 ( .A(n380), .Y(n294) );
  MUX21X2_HVT U76 ( .A1(n547), .A2(n546), .S0(n226), .Y(n545) );
  IBUFFX16_HVT U77 ( .A(n351), .Y(n226) );
  INVX0_HVT U84 ( .A(n240), .Y(n227) );
  INVX1_HVT U85 ( .A(n633), .Y(n408) );
  OA21X2_HVT U86 ( .A1(n393), .A2(n388), .A3(n633), .Y(n579) );
  MUX41X1_HVT U87 ( .A1(n433), .A3(n412), .A2(n641), .A4(n426), .S0(n319), 
        .S1(n388), .Y(n561) );
  MUX41X1_HVT U90 ( .A1(n408), .A3(n617), .A2(n495), .A4(n646), .S0(n228), 
        .S1(n229), .Y(n494) );
  IBUFFX16_HVT U91 ( .A(n346), .Y(n228) );
  IBUFFX16_HVT U92 ( .A(n387), .Y(n229) );
  INVX0_HVT U93 ( .A(n610), .Y(n422) );
  NAND2X0_HVT U94 ( .A1(n570), .A2(n230), .Y(n231) );
  NAND2X0_HVT U95 ( .A1(n577), .A2(n289), .Y(n232) );
  NAND2X0_HVT U96 ( .A1(n231), .A2(n232), .Y(out[1]) );
  INVX1_HVT U97 ( .A(n289), .Y(n230) );
  IBUFFX2_HVT U100 ( .A(n310), .Y(n289) );
  INVX1_HVT U103 ( .A(n375), .Y(n263) );
  INVX1_HVT U106 ( .A(n293), .Y(n257) );
  INVX1_HVT U111 ( .A(n446), .Y(n335) );
  INVX0_HVT U113 ( .A(n446), .Y(n336) );
  MUX21X1_HVT U117 ( .A1(n234), .A2(n446), .S0(n247), .Y(n233) );
  IBUFFX16_HVT U121 ( .A(n369), .Y(n236) );
  INVX1_HVT U123 ( .A(n256), .Y(n238) );
  INVX0_HVT U125 ( .A(n374), .Y(n341) );
  INVX1_HVT U126 ( .A(n448), .Y(n440) );
  MUX21X2_HVT U128 ( .A1(n580), .A2(n579), .S0(n239), .Y(n578) );
  IBUFFX16_HVT U134 ( .A(n292), .Y(n239) );
  INVX2_HVT U135 ( .A(in[0]), .Y(n380) );
  INVX0_HVT U138 ( .A(n255), .Y(n626) );
  MUX21X1_HVT U140 ( .A1(n222), .A2(n442), .S0(n375), .Y(n509) );
  IBUFFX2_HVT U143 ( .A(n636), .Y(n405) );
  INVX0_HVT U144 ( .A(n240), .Y(n241) );
  NAND2X0_HVT U146 ( .A1(n503), .A2(n242), .Y(n243) );
  NAND2X0_HVT U147 ( .A1(n513), .A2(n245), .Y(n244) );
  NAND2X0_HVT U148 ( .A1(n243), .A2(n244), .Y(out[5]) );
  INVX1_HVT U149 ( .A(n245), .Y(n242) );
  INVX1_HVT U150 ( .A(n285), .Y(n245) );
  INVX2_HVT U151 ( .A(n638), .Y(n446) );
  INVX0_HVT U152 ( .A(n638), .Y(n340) );
  INVX0_HVT U153 ( .A(n638), .Y(n339) );
  MUX21X1_HVT U154 ( .A1(n241), .A2(n591), .S0(n334), .Y(n590) );
  MUX21X2_HVT U156 ( .A1(n372), .A2(n336), .S0(n91), .Y(n342) );
  MUX41X1_HVT U157 ( .A1(n410), .A3(n643), .A2(n416), .A4(n330), .S0(n353), 
        .S1(n246), .Y(n519) );
  IBUFFX16_HVT U158 ( .A(n345), .Y(n246) );
  IBUFFX16_HVT U160 ( .A(n352), .Y(n247) );
  NAND2X0_HVT U161 ( .A1(n337), .A2(n248), .Y(n249) );
  NAND2X0_HVT U164 ( .A1(n359), .A2(n375), .Y(n250) );
  NAND2X0_HVT U165 ( .A1(n249), .A2(n250), .Y(n629) );
  NBUFFX2_HVT U167 ( .A(n447), .Y(n359) );
  IBUFFX2_HVT U169 ( .A(n389), .Y(n386) );
  INVX1_HVT U171 ( .A(n389), .Y(n385) );
  INVX0_HVT U173 ( .A(n608), .Y(n424) );
  INVX0_HVT U175 ( .A(n197), .Y(n287) );
  IBUFFX2_HVT U176 ( .A(n380), .Y(n376) );
  INVX2_HVT U178 ( .A(n389), .Y(n384) );
  MUX21X2_HVT U181 ( .A1(n611), .A2(n428), .S0(n268), .Y(n502) );
  INVX1_HVT U182 ( .A(n384), .Y(n298) );
  INVX2_HVT U184 ( .A(n267), .Y(n268) );
  XOR2X2_HVT U186 ( .A1(n222), .A2(n251), .Y(n638) );
  MUX21X2_HVT U187 ( .A1(n367), .A2(n256), .S0(n257), .Y(n255) );
  INVX0_HVT U188 ( .A(n444), .Y(n256) );
  INVX1_HVT U189 ( .A(n282), .Y(n251) );
  INVX0_HVT U190 ( .A(in[3]), .Y(n282) );
  NBUFFX2_HVT U193 ( .A(n443), .Y(n355) );
  AO21X1_HVT U196 ( .A1(n196), .A2(n441), .A3(n388), .Y(n465) );
  NAND2X0_HVT U197 ( .A1(n476), .A2(n252), .Y(n253) );
  NAND2X0_HVT U199 ( .A1(n475), .A2(n360), .Y(n254) );
  NAND2X0_HVT U201 ( .A1(n253), .A2(n254), .Y(n474) );
  IBUFFX2_HVT U202 ( .A(n360), .Y(n252) );
  INVX0_HVT U203 ( .A(n260), .Y(n611) );
  INVX1_HVT U204 ( .A(n368), .Y(n445) );
  INVX1_HVT U205 ( .A(n652), .Y(n394) );
  INVX1_HVT U206 ( .A(n356), .Y(n261) );
  IBUFFX2_HVT U208 ( .A(n355), .Y(n323) );
  INVX0_HVT U209 ( .A(n612), .Y(n396) );
  INVX1_HVT U210 ( .A(n394), .Y(n278) );
  MUX41X1_HVT U211 ( .A1(n342), .A3(n509), .A2(n272), .A4(n419), .S0(n354), 
        .S1(n258), .Y(n508) );
  IBUFFX16_HVT U212 ( .A(n343), .Y(n258) );
  INVX1_HVT U213 ( .A(n446), .Y(n337) );
  MUX21X2_HVT U214 ( .A1(n368), .A2(n261), .S0(n301), .Y(n260) );
  MUX41X1_HVT U215 ( .A1(n481), .A3(n332), .A2(n610), .A4(n238), .S0(n262), 
        .S1(n386), .Y(n480) );
  IBUFFX16_HVT U216 ( .A(n349), .Y(n262) );
  INVX0_HVT U217 ( .A(n366), .Y(n305) );
  INVX1_HVT U218 ( .A(n266), .Y(n324) );
  MUX21X1_HVT U219 ( .A1(n359), .A2(n441), .S0(n263), .Y(n460) );
  IBUFFX16_HVT U220 ( .A(n288), .Y(n264) );
  MUX41X1_HVT U221 ( .A1(n517), .A3(n519), .A2(n514), .A4(n516), .S0(n361), 
        .S1(n265), .Y(n513) );
  IBUFFX16_HVT U222 ( .A(n364), .Y(n265) );
  IBUFFX2_HVT U223 ( .A(n380), .Y(n378) );
  INVX1_HVT U224 ( .A(in[4]), .Y(n389) );
  MUX21X1_HVT U225 ( .A1(n305), .A2(n270), .S0(n91), .Y(n266) );
  INVX1_HVT U226 ( .A(n288), .Y(n267) );
  INVX1_HVT U227 ( .A(n288), .Y(n269) );
  AO21X2_HVT U228 ( .A1(n338), .A2(n278), .A3(n269), .Y(n491) );
  NBUFFX2_HVT U229 ( .A(n384), .Y(n352) );
  IBUFFX2_HVT U230 ( .A(n447), .Y(n270) );
  MUX41X1_HVT U231 ( .A1(n571), .A3(n572), .A2(n575), .A4(n576), .S0(n361), 
        .S1(n364), .Y(n570) );
  INVX1_HVT U232 ( .A(n360), .Y(n361) );
  IBUFFX2_HVT U233 ( .A(n389), .Y(n387) );
  MUX41X1_HVT U234 ( .A1(n504), .A3(n508), .A2(n505), .A4(n510), .S0(n365), 
        .S1(n271), .Y(n503) );
  IBUFFX16_HVT U235 ( .A(n360), .Y(n271) );
  MUX41X1_HVT U236 ( .A1(n413), .A3(n629), .A2(n333), .A4(n431), .S0(n309), 
        .S1(n273), .Y(n571) );
  INVX2_HVT U237 ( .A(n456), .Y(n431) );
  IBUFFX2_HVT U238 ( .A(n348), .Y(n273) );
  INVX0_HVT U239 ( .A(n342), .Y(n632) );
  INVX1_HVT U240 ( .A(n286), .Y(n613) );
  INVX1_HVT U241 ( .A(n388), .Y(n288) );
  NBUFFX2_HVT U242 ( .A(n430), .Y(n272) );
  NAND2X0_HVT U243 ( .A1(n409), .A2(n274), .Y(n275) );
  NAND2X0_HVT U244 ( .A1(n598), .A2(n334), .Y(n276) );
  NAND2X0_HVT U245 ( .A1(n275), .A2(n276), .Y(n597) );
  INVX0_HVT U246 ( .A(n334), .Y(n274) );
  MUX21X2_HVT U247 ( .A1(n335), .A2(n356), .S0(n294), .Y(n633) );
  INVX0_HVT U248 ( .A(n654), .Y(n441) );
  NAND2X0_HVT U249 ( .A1(n376), .A2(n371), .Y(n652) );
  NAND2X0_HVT U250 ( .A1(n506), .A2(n279), .Y(n280) );
  NAND2X0_HVT U251 ( .A1(n507), .A2(n351), .Y(n281) );
  NAND2X0_HVT U252 ( .A1(n280), .A2(n281), .Y(n505) );
  IBUFFX2_HVT U253 ( .A(n351), .Y(n279) );
  MUX21X1_HVT U254 ( .A1(n333), .A2(n629), .S0(n298), .Y(n507) );
  INVX1_HVT U255 ( .A(n352), .Y(n313) );
  OR2X1_HVT U256 ( .A1(n282), .A2(n358), .Y(n653) );
  MUX41X1_HVT U257 ( .A1(n487), .A3(n485), .A2(n484), .A4(n483), .S0(n283), 
        .S1(n284), .Y(n482) );
  IBUFFX16_HVT U258 ( .A(n361), .Y(n283) );
  IBUFFX16_HVT U259 ( .A(n364), .Y(n284) );
  INVX0_HVT U260 ( .A(n358), .Y(n327) );
  IBUFFX16_HVT U261 ( .A(in[7]), .Y(n285) );
  MUX21X1_HVT U262 ( .A1(n368), .A2(n359), .S0(n287), .Y(n286) );
  MUX21X2_HVT U263 ( .A1(n397), .A2(n613), .S0(n352), .Y(n547) );
  IBUFFX2_HVT U264 ( .A(in[4]), .Y(n388) );
  MUX41X1_HVT U265 ( .A1(n599), .A3(n593), .A2(n601), .A4(n597), .S0(n290), 
        .S1(n291), .Y(n592) );
  IBUFFX16_HVT U266 ( .A(n364), .Y(n290) );
  IBUFFX16_HVT U267 ( .A(n360), .Y(n291) );
  OA21X2_HVT U268 ( .A1(n392), .A2(n269), .A3(n399), .Y(n506) );
  INVX1_HVT U269 ( .A(n380), .Y(n375) );
  NAND2X0_HVT U270 ( .A1(n501), .A2(n320), .Y(n317) );
  INVX0_HVT U271 ( .A(n369), .Y(n304) );
  INVX1_HVT U272 ( .A(n457), .Y(n430) );
  INVX1_HVT U273 ( .A(n348), .Y(n320) );
  INVX0_HVT U274 ( .A(n348), .Y(n319) );
  INVX0_HVT U275 ( .A(n347), .Y(n297) );
  INVX0_HVT U276 ( .A(n351), .Y(n292) );
  INVX1_HVT U277 ( .A(in[1]), .Y(n360) );
  INVX1_HVT U278 ( .A(n360), .Y(n362) );
  INVX0_HVT U279 ( .A(n363), .Y(n365) );
  INVX1_HVT U280 ( .A(in[5]), .Y(n363) );
  INVX1_HVT U281 ( .A(in[7]), .Y(n310) );
  MUX41X1_HVT U282 ( .A1(n468), .A3(n477), .A2(n462), .A4(n474), .S0(n314), 
        .S1(n363), .Y(out[7]) );
  MUX21X1_HVT U283 ( .A1(n423), .A2(n331), .S0(n353), .Y(n464) );
  MUX21X2_HVT U284 ( .A1(n548), .A2(n538), .S0(n310), .Y(out[3]) );
  IBUFFX2_HVT U285 ( .A(n380), .Y(n293) );
  IBUFFX2_HVT U286 ( .A(n380), .Y(n379) );
  NAND2X0_HVT U287 ( .A1(n278), .A2(n350), .Y(n295) );
  NAND2X0_HVT U288 ( .A1(n342), .A2(n320), .Y(n296) );
  NAND2X0_HVT U289 ( .A1(n295), .A2(n296), .Y(n591) );
  MUX41X1_HVT U290 ( .A1(n398), .A3(n643), .A2(n238), .A4(n300), .S0(n297), 
        .S1(n298), .Y(n584) );
  IBUFFX2_HVT U291 ( .A(n396), .Y(n299) );
  INVX1_HVT U292 ( .A(n395), .Y(n300) );
  INVX0_HVT U293 ( .A(n649), .Y(n395) );
  INVX1_HVT U294 ( .A(n380), .Y(n377) );
  MUX41X1_HVT U295 ( .A1(n396), .A3(n394), .A2(n278), .A4(n430), .S0(n386), 
        .S1(n346), .Y(n476) );
  NAND2X0_HVT U296 ( .A1(n511), .A2(n345), .Y(n302) );
  NAND2X0_HVT U297 ( .A1(n512), .A2(n292), .Y(n303) );
  NAND2X0_HVT U298 ( .A1(n302), .A2(n303), .Y(n510) );
  MUX21X1_HVT U299 ( .A1(n439), .A2(n306), .S0(n352), .Y(n512) );
  INVX1_HVT U300 ( .A(n449), .Y(n439) );
  MUX41X1_HVT U301 ( .A1(n618), .A3(n371), .A2(n238), .A4(n374), .S0(n319), 
        .S1(n269), .Y(n484) );
  IBUFFX2_HVT U302 ( .A(n618), .Y(n418) );
  OR2X1_HVT U303 ( .A1(n301), .A2(n304), .Y(n648) );
  MUX41X1_HVT U304 ( .A1(n568), .A3(n563), .A2(n569), .A4(n566), .S0(n363), 
        .S1(n362), .Y(n562) );
  INVX1_HVT U305 ( .A(n363), .Y(n364) );
  XNOR2X1_HVT U306 ( .A1(n305), .A2(n294), .Y(n606) );
  INVX0_HVT U307 ( .A(n651), .Y(n306) );
  INVX0_HVT U308 ( .A(n609), .Y(n423) );
  NAND2X0_HVT U309 ( .A1(n564), .A2(n292), .Y(n307) );
  NAND2X0_HVT U310 ( .A1(n565), .A2(n350), .Y(n308) );
  NAND2X0_HVT U311 ( .A1(n307), .A2(n308), .Y(n563) );
  INVX1_HVT U312 ( .A(n627), .Y(n412) );
  NBUFFX2_HVT U313 ( .A(n384), .Y(n309) );
  NAND2X0_HVT U314 ( .A1(n480), .A2(n361), .Y(n311) );
  NAND2X0_HVT U315 ( .A1(n478), .A2(n360), .Y(n312) );
  NAND2X0_HVT U316 ( .A1(n311), .A2(n312), .Y(n477) );
  MUX21X1_HVT U317 ( .A1(n444), .A2(n442), .S0(n380), .Y(n610) );
  MUX41X1_HVT U318 ( .A1(n590), .A3(n587), .A2(n589), .A4(n586), .S0(n363), 
        .S1(n360), .Y(n585) );
  NAND2X0_HVT U319 ( .A1(n489), .A2(n314), .Y(n315) );
  NAND2X0_HVT U320 ( .A1(n482), .A2(n310), .Y(n316) );
  NAND2X0_HVT U321 ( .A1(n315), .A2(n316), .Y(out[6]) );
  INVX1_HVT U322 ( .A(n310), .Y(n314) );
  NAND2X0_HVT U323 ( .A1(n502), .A2(n351), .Y(n318) );
  NAND2X0_HVT U324 ( .A1(n317), .A2(n318), .Y(n498) );
  MUX41X1_HVT U325 ( .A1(n600), .A3(n411), .A2(n337), .A4(n324), .S0(n320), 
        .S1(n313), .Y(n599) );
  NAND2X0_HVT U326 ( .A1(n585), .A2(n310), .Y(n321) );
  NAND2X0_HVT U327 ( .A1(n592), .A2(in[7]), .Y(n322) );
  NAND2X0_HVT U328 ( .A1(n321), .A2(n322), .Y(out[0]) );
  MUX21X1_HVT U329 ( .A1(n628), .A2(n631), .S0(n353), .Y(n493) );
  NAND2X0_HVT U330 ( .A1(n492), .A2(n320), .Y(n325) );
  MUX41X1_HVT U331 ( .A1(n411), .A3(n432), .A2(n333), .A4(n394), .S0(n297), 
        .S1(n388), .Y(n569) );
  MUX21X2_HVT U332 ( .A1(n537), .A2(n535), .S0(n360), .Y(n534) );
  INVX0_HVT U333 ( .A(in[3]), .Y(n443) );
  MUX41X1_HVT U334 ( .A1(n631), .A3(n634), .A2(n260), .A4(n442), .S0(n320), 
        .S1(n313), .Y(n516) );
  NAND2X0_HVT U335 ( .A1(n493), .A2(n350), .Y(n326) );
  NAND2X0_HVT U336 ( .A1(n326), .A2(n325), .Y(n490) );
  MUX21X1_HVT U337 ( .A1(n473), .A2(n429), .S0(n352), .Y(n472) );
  NBUFFX2_HVT U338 ( .A(n654), .Y(n372) );
  AND2X1_HVT U339 ( .A1(n649), .A2(n371), .Y(n328) );
  AND2X1_HVT U340 ( .A1(n371), .A2(n639), .Y(n329) );
  MUX21X1_HVT U341 ( .A1(n398), .A2(n336), .S0(n354), .Y(n564) );
  MUX21X1_HVT U342 ( .A1(n335), .A2(n442), .S0(n376), .Y(n620) );
  INVX1_HVT U343 ( .A(n366), .Y(n442) );
  MUX21X1_HVT U344 ( .A1(n445), .A2(n356), .S0(n378), .Y(n459) );
  AO21X1_HVT U345 ( .A1(n354), .A2(n224), .A3(n441), .Y(n511) );
  MUX21X1_HVT U346 ( .A1(n356), .A2(n371), .S0(n376), .Y(n458) );
  MUX21X1_HVT U347 ( .A1(n366), .A2(n369), .S0(n376), .Y(n497) );
  MUX21X1_HVT U348 ( .A1(n370), .A2(n371), .S0(n196), .Y(n636) );
  MUX21X1_HVT U349 ( .A1(n359), .A2(n338), .S0(n379), .Y(n614) );
  MUX21X1_HVT U350 ( .A1(n223), .A2(n371), .S0(n377), .Y(n552) );
  MUX21X1_HVT U351 ( .A1(n366), .A2(n372), .S0(n294), .Y(n449) );
  MUX21X1_HVT U352 ( .A1(n621), .A2(n329), .S0(n351), .Y(n530) );
  XNOR2X1_HVT U353 ( .A1(n372), .A2(n376), .Y(n330) );
  MUX21X1_HVT U354 ( .A1(n369), .A2(n357), .S0(n293), .Y(n635) );
  MUX21X1_HVT U355 ( .A1(n438), .A2(n330), .S0(n350), .Y(n533) );
  AND2X1_HVT U356 ( .A1(n294), .A2(n223), .Y(n331) );
  MUX21X1_HVT U357 ( .A1(n355), .A2(n369), .S0(n293), .Y(n452) );
  NBUFFX2_HVT U358 ( .A(n384), .Y(n354) );
  NBUFFX2_HVT U359 ( .A(n384), .Y(n353) );
  AND2X1_HVT U360 ( .A1(n445), .A2(n381), .Y(n332) );
  MUX21X1_HVT U361 ( .A1(n410), .A2(n651), .S0(n351), .Y(n598) );
  NBUFFX2_HVT U362 ( .A(n650), .Y(n366) );
  NBUFFX2_HVT U363 ( .A(n653), .Y(n368) );
  AND2X1_HVT U364 ( .A1(n370), .A2(n381), .Y(n333) );
  MUX21X1_HVT U365 ( .A1(n372), .A2(n367), .S0(n376), .Y(n515) );
  NAND2X0_HVT U366 ( .A1(n381), .A2(n441), .Y(n557) );
  NBUFFX2_HVT U367 ( .A(n653), .Y(n370) );
  NBUFFX2_HVT U368 ( .A(n650), .Y(n367) );
  NBUFFX2_HVT U369 ( .A(n653), .Y(n369) );
  NBUFFX2_HVT U370 ( .A(n443), .Y(n357) );
  NBUFFX2_HVT U371 ( .A(n443), .Y(n356) );
  NBUFFX2_HVT U372 ( .A(n344), .Y(n349) );
  NBUFFX2_HVT U373 ( .A(n382), .Y(n351) );
  NBUFFX2_HVT U374 ( .A(n383), .Y(n350) );
  NBUFFX2_HVT U375 ( .A(n382), .Y(n343) );
  XNOR2X1_HVT U376 ( .A1(n388), .A2(n346), .Y(n334) );
  NBUFFX2_HVT U377 ( .A(n383), .Y(n346) );
  NBUFFX2_HVT U378 ( .A(n383), .Y(n348) );
  NBUFFX2_HVT U379 ( .A(n382), .Y(n344) );
  NBUFFX2_HVT U380 ( .A(n383), .Y(n347) );
  NBUFFX2_HVT U381 ( .A(n382), .Y(n345) );
  MUX21X1_HVT U382 ( .A1(n374), .A2(n323), .S0(n378), .Y(n500) );
  MUX21X1_HVT U383 ( .A1(n521), .A2(n522), .S0(n361), .Y(n520) );
  MUX21X1_HVT U384 ( .A1(n525), .A2(n526), .S0(n362), .Y(n524) );
  MUX21X1_HVT U385 ( .A1(n367), .A2(n323), .S0(n294), .Y(n560) );
  MUX21X1_HVT U386 ( .A1(n323), .A2(n374), .S0(n375), .Y(n454) );
  MUX21X1_HVT U387 ( .A1(n359), .A2(n323), .S0(n196), .Y(n627) );
  MUX21X1_HVT U388 ( .A1(n445), .A2(n442), .S0(n378), .Y(n541) );
  MUX21X1_HVT U389 ( .A1(n323), .A2(n367), .S0(n377), .Y(n453) );
  NBUFFX2_HVT U390 ( .A(in[2]), .Y(n382) );
  NBUFFX2_HVT U391 ( .A(in[2]), .Y(n383) );
  INVX1_HVT U392 ( .A(n460), .Y(n427) );
  MUX21X1_HVT U393 ( .A1(n357), .A2(n441), .S0(n293), .Y(n624) );
  MUX21X1_HVT U394 ( .A1(n441), .A2(n445), .S0(n197), .Y(n604) );
  NBUFFX2_HVT U395 ( .A(n655), .Y(n374) );
  MUX21X1_HVT U396 ( .A1(n370), .A2(n222), .S0(n375), .Y(n536) );
  MUX21X1_HVT U397 ( .A1(n222), .A2(n441), .S0(n294), .Y(n628) );
  MUX21X1_HVT U398 ( .A1(n357), .A2(n359), .S0(n197), .Y(n609) );
  MUX21X1_HVT U399 ( .A1(n373), .A2(n372), .S0(n197), .Y(n640) );
  MUX21X1_HVT U400 ( .A1(n341), .A2(n323), .S0(n379), .Y(n448) );
  MUX21X1_HVT U401 ( .A1(n341), .A2(n335), .S0(n293), .Y(n455) );
  MUX21X1_HVT U402 ( .A1(n337), .A2(n444), .S0(n377), .Y(n623) );
  XOR2X1_HVT U403 ( .A1(n373), .A2(n379), .Y(n617) );
  NAND2X0_HVT U404 ( .A1(n355), .A2(n223), .Y(n654) );
  NBUFFX2_HVT U405 ( .A(n654), .Y(n371) );
  MUX21X1_HVT U406 ( .A1(n340), .A2(n357), .S0(n376), .Y(n615) );
  MUX21X1_HVT U407 ( .A1(n359), .A2(n340), .S0(n293), .Y(n618) );
  MUX21X1_HVT U408 ( .A1(n355), .A2(n339), .S0(n378), .Y(n457) );
  MUX21X1_HVT U409 ( .A1(n441), .A2(n340), .S0(n197), .Y(n621) );
  MUX21X1_HVT U410 ( .A1(n340), .A2(n222), .S0(n294), .Y(n450) );
  MUX21X1_HVT U411 ( .A1(n441), .A2(n327), .S0(n375), .Y(n523) );
  XOR2X1_HVT U412 ( .A1(n196), .A2(n327), .Y(n605) );
  MUX21X1_HVT U413 ( .A1(n327), .A2(n341), .S0(n379), .Y(n630) );
  MUX21X1_HVT U414 ( .A1(n369), .A2(n327), .S0(n379), .Y(n456) );
  MUX21X1_HVT U415 ( .A1(n327), .A2(n370), .S0(n379), .Y(n461) );
  MUX21X1_HVT U416 ( .A1(n327), .A2(n373), .S0(n379), .Y(n637) );
  MUX21X1_HVT U417 ( .A1(n355), .A2(n327), .S0(n197), .Y(n451) );
  MUX21X1_HVT U418 ( .A1(n367), .A2(n327), .S0(n378), .Y(n625) );
  NBUFFX2_HVT U419 ( .A(n655), .Y(n373) );
  MUX21X1_HVT U420 ( .A1(n444), .A2(n445), .S0(n378), .Y(n488) );
  MUX21X1_HVT U421 ( .A1(n444), .A2(n222), .S0(n378), .Y(n486) );
  INVX0_HVT U422 ( .A(n622), .Y(n390) );
  INVX0_HVT U423 ( .A(n616), .Y(n391) );
  INVX0_HVT U424 ( .A(n557), .Y(n392) );
  INVX0_HVT U425 ( .A(n518), .Y(n393) );
  INVX0_HVT U426 ( .A(n648), .Y(n397) );
  INVX0_HVT U427 ( .A(n619), .Y(n398) );
  INVX0_HVT U428 ( .A(n641), .Y(n399) );
  INVX0_HVT U429 ( .A(n646), .Y(n400) );
  INVX0_HVT U430 ( .A(n642), .Y(n401) );
  INVX0_HVT U431 ( .A(n640), .Y(n402) );
  INVX0_HVT U432 ( .A(n639), .Y(n403) );
  INVX0_HVT U433 ( .A(n637), .Y(n404) );
  INVX0_HVT U434 ( .A(n635), .Y(n406) );
  INVX0_HVT U435 ( .A(n634), .Y(n407) );
  INVX0_HVT U436 ( .A(n630), .Y(n409) );
  INVX0_HVT U437 ( .A(n628), .Y(n411) );
  INVX0_HVT U438 ( .A(n625), .Y(n413) );
  INVX0_HVT U439 ( .A(n624), .Y(n414) );
  INVX0_HVT U440 ( .A(n623), .Y(n415) );
  INVX0_HVT U441 ( .A(n621), .Y(n416) );
  INVX0_HVT U442 ( .A(n620), .Y(n417) );
  INVX0_HVT U443 ( .A(n617), .Y(n419) );
  INVX0_HVT U444 ( .A(n615), .Y(n420) );
  INVX0_HVT U445 ( .A(n614), .Y(n421) );
  INVX0_HVT U446 ( .A(n645), .Y(n425) );
  INVX0_HVT U447 ( .A(n461), .Y(n426) );
  INVX0_HVT U448 ( .A(n458), .Y(n429) );
  INVX0_HVT U449 ( .A(n455), .Y(n432) );
  INVX0_HVT U450 ( .A(n454), .Y(n433) );
  INVX0_HVT U451 ( .A(n453), .Y(n434) );
  INVX0_HVT U452 ( .A(n452), .Y(n435) );
  INVX0_HVT U453 ( .A(n451), .Y(n436) );
  INVX0_HVT U454 ( .A(n500), .Y(n437) );
  INVX0_HVT U455 ( .A(n450), .Y(n438) );
endmodule

