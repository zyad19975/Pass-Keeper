
module inv_aes ( clk, rest, start, plaintext1, local_key, cipher_text, done, 
        busy );
  input [127:0] plaintext1;
  input [127:0] local_key;
  output [127:0] cipher_text;
  input clk, rest, start;
  output done, busy;
  wire   last, done_k, n205, n206, n208, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n207, n209,
         n605, n606, n607, n608, n609;
  wire   [127:0] adk_out;
  wire   [127:0] keys1;
  wire   [127:0] out1;
  wire   [3:0] rount_no;
  wire   [127:0] key_round;
  wire   [3:0] state;

  DFFARX1_HVT flag_reg ( .D(n208), .CLK(clk), .RSTB(n5), .Q(n608) );
  DFFASX1_HVT \rount_no_reg[3]  ( .D(n595), .CLK(clk), .SETB(n5), .Q(
        rount_no[3]) );
  DFFARX1_HVT \state_reg[1]  ( .D(n599), .CLK(clk), .RSTB(n5), .Q(state[1]), 
        .QN(n4) );
  DFFASX1_HVT \state_reg[2]  ( .D(n602), .CLK(clk), .SETB(n5), .Q(state[2]), 
        .QN(n1) );
  DFFASX1_HVT \state_reg[0]  ( .D(n600), .CLK(clk), .SETB(n5), .Q(state[0]), 
        .QN(n3) );
  DFFASX1_HVT \state_reg[3]  ( .D(n601), .CLK(clk), .SETB(n5), .Q(state[3]), 
        .QN(n2) );
  DFFARX1_HVT done_reg ( .D(n603), .CLK(clk), .RSTB(n5), .Q(done), .QN(n206)
         );
  DFFARX1_HVT busy_reg ( .D(n604), .CLK(clk), .RSTB(n5), .Q(busy), .QN(n205)
         );
  DFFARX1_HVT \rount_no_reg[0]  ( .D(n598), .CLK(clk), .RSTB(n5), .Q(
        rount_no[0]) );
  DFFASX1_HVT \rount_no_reg[1]  ( .D(n597), .CLK(clk), .SETB(n5), .Q(
        rount_no[1]) );
  DFFARX1_HVT \rount_no_reg[2]  ( .D(n596), .CLK(clk), .RSTB(n5), .Q(
        rount_no[2]) );
  DFFX1_HVT \keys1_reg[0]  ( .D(n594), .CLK(clk), .Q(keys1[0]) );
  DFFX1_HVT \keys1_reg[1]  ( .D(n593), .CLK(clk), .Q(keys1[1]) );
  DFFX1_HVT \keys1_reg[2]  ( .D(n592), .CLK(clk), .Q(keys1[2]) );
  DFFX1_HVT \keys1_reg[3]  ( .D(n591), .CLK(clk), .Q(keys1[3]) );
  DFFX1_HVT \keys1_reg[4]  ( .D(n590), .CLK(clk), .Q(keys1[4]) );
  DFFX1_HVT \keys1_reg[5]  ( .D(n589), .CLK(clk), .Q(keys1[5]) );
  DFFX1_HVT \keys1_reg[6]  ( .D(n588), .CLK(clk), .Q(keys1[6]) );
  DFFX1_HVT \keys1_reg[7]  ( .D(n587), .CLK(clk), .Q(keys1[7]) );
  DFFX1_HVT \keys1_reg[8]  ( .D(n586), .CLK(clk), .Q(keys1[8]) );
  DFFX1_HVT \keys1_reg[9]  ( .D(n585), .CLK(clk), .Q(keys1[9]) );
  DFFX1_HVT \keys1_reg[10]  ( .D(n584), .CLK(clk), .Q(keys1[10]) );
  DFFX1_HVT \keys1_reg[11]  ( .D(n583), .CLK(clk), .Q(keys1[11]) );
  DFFX1_HVT \keys1_reg[12]  ( .D(n582), .CLK(clk), .Q(keys1[12]) );
  DFFX1_HVT \keys1_reg[13]  ( .D(n581), .CLK(clk), .Q(keys1[13]) );
  DFFX1_HVT \keys1_reg[14]  ( .D(n580), .CLK(clk), .Q(keys1[14]) );
  DFFX1_HVT \keys1_reg[15]  ( .D(n579), .CLK(clk), .Q(keys1[15]) );
  DFFX1_HVT \keys1_reg[16]  ( .D(n578), .CLK(clk), .Q(keys1[16]) );
  DFFX1_HVT \keys1_reg[17]  ( .D(n577), .CLK(clk), .Q(keys1[17]) );
  DFFX1_HVT \keys1_reg[18]  ( .D(n576), .CLK(clk), .Q(keys1[18]) );
  DFFX1_HVT \keys1_reg[19]  ( .D(n575), .CLK(clk), .Q(keys1[19]) );
  DFFX1_HVT \keys1_reg[20]  ( .D(n574), .CLK(clk), .Q(keys1[20]) );
  DFFX1_HVT \keys1_reg[21]  ( .D(n573), .CLK(clk), .Q(keys1[21]) );
  DFFX1_HVT \keys1_reg[22]  ( .D(n572), .CLK(clk), .Q(keys1[22]) );
  DFFX1_HVT \keys1_reg[23]  ( .D(n571), .CLK(clk), .Q(keys1[23]) );
  DFFX1_HVT \keys1_reg[24]  ( .D(n570), .CLK(clk), .Q(keys1[24]) );
  DFFX1_HVT \keys1_reg[25]  ( .D(n569), .CLK(clk), .Q(keys1[25]) );
  DFFX1_HVT \keys1_reg[26]  ( .D(n568), .CLK(clk), .Q(keys1[26]) );
  DFFX1_HVT \keys1_reg[27]  ( .D(n567), .CLK(clk), .Q(keys1[27]) );
  DFFX1_HVT \keys1_reg[28]  ( .D(n566), .CLK(clk), .Q(keys1[28]) );
  DFFX1_HVT \keys1_reg[29]  ( .D(n565), .CLK(clk), .Q(keys1[29]) );
  DFFX1_HVT \keys1_reg[30]  ( .D(n564), .CLK(clk), .Q(keys1[30]) );
  DFFX1_HVT \keys1_reg[31]  ( .D(n563), .CLK(clk), .Q(keys1[31]) );
  DFFX1_HVT \keys1_reg[32]  ( .D(n562), .CLK(clk), .Q(keys1[32]) );
  DFFX1_HVT \keys1_reg[33]  ( .D(n561), .CLK(clk), .Q(keys1[33]) );
  DFFX1_HVT \keys1_reg[34]  ( .D(n560), .CLK(clk), .Q(keys1[34]) );
  DFFX1_HVT \keys1_reg[35]  ( .D(n559), .CLK(clk), .Q(keys1[35]) );
  DFFX1_HVT \keys1_reg[36]  ( .D(n558), .CLK(clk), .Q(keys1[36]) );
  DFFX1_HVT \keys1_reg[37]  ( .D(n557), .CLK(clk), .Q(keys1[37]) );
  DFFX1_HVT \keys1_reg[38]  ( .D(n556), .CLK(clk), .Q(keys1[38]) );
  DFFX1_HVT \keys1_reg[39]  ( .D(n555), .CLK(clk), .Q(keys1[39]) );
  DFFX1_HVT \keys1_reg[40]  ( .D(n554), .CLK(clk), .Q(keys1[40]) );
  DFFX1_HVT \keys1_reg[41]  ( .D(n553), .CLK(clk), .Q(keys1[41]) );
  DFFX1_HVT \keys1_reg[42]  ( .D(n552), .CLK(clk), .Q(keys1[42]) );
  DFFX1_HVT \keys1_reg[43]  ( .D(n551), .CLK(clk), .Q(keys1[43]) );
  DFFX1_HVT \keys1_reg[44]  ( .D(n550), .CLK(clk), .Q(keys1[44]) );
  DFFX1_HVT \keys1_reg[45]  ( .D(n549), .CLK(clk), .Q(keys1[45]) );
  DFFX1_HVT \keys1_reg[46]  ( .D(n548), .CLK(clk), .Q(keys1[46]) );
  DFFX1_HVT \keys1_reg[47]  ( .D(n547), .CLK(clk), .Q(keys1[47]) );
  DFFX1_HVT \keys1_reg[48]  ( .D(n546), .CLK(clk), .Q(keys1[48]) );
  DFFX1_HVT \keys1_reg[49]  ( .D(n545), .CLK(clk), .Q(keys1[49]) );
  DFFX1_HVT \keys1_reg[50]  ( .D(n544), .CLK(clk), .Q(keys1[50]) );
  DFFX1_HVT \keys1_reg[51]  ( .D(n543), .CLK(clk), .Q(keys1[51]) );
  DFFX1_HVT \keys1_reg[52]  ( .D(n542), .CLK(clk), .Q(keys1[52]) );
  DFFX1_HVT \keys1_reg[53]  ( .D(n541), .CLK(clk), .Q(keys1[53]) );
  DFFX1_HVT \keys1_reg[54]  ( .D(n540), .CLK(clk), .Q(keys1[54]) );
  DFFX1_HVT \keys1_reg[55]  ( .D(n539), .CLK(clk), .Q(keys1[55]) );
  DFFX1_HVT \keys1_reg[56]  ( .D(n538), .CLK(clk), .Q(keys1[56]) );
  DFFX1_HVT \keys1_reg[57]  ( .D(n537), .CLK(clk), .Q(keys1[57]) );
  DFFX1_HVT \keys1_reg[58]  ( .D(n536), .CLK(clk), .Q(keys1[58]) );
  DFFX1_HVT \keys1_reg[59]  ( .D(n535), .CLK(clk), .Q(keys1[59]) );
  DFFX1_HVT \keys1_reg[60]  ( .D(n534), .CLK(clk), .Q(keys1[60]) );
  DFFX1_HVT \keys1_reg[61]  ( .D(n533), .CLK(clk), .Q(keys1[61]) );
  DFFX1_HVT \keys1_reg[62]  ( .D(n532), .CLK(clk), .Q(keys1[62]) );
  DFFX1_HVT \keys1_reg[63]  ( .D(n531), .CLK(clk), .Q(keys1[63]) );
  DFFX1_HVT \keys1_reg[64]  ( .D(n530), .CLK(clk), .Q(keys1[64]) );
  DFFX1_HVT \keys1_reg[65]  ( .D(n529), .CLK(clk), .Q(keys1[65]) );
  DFFX1_HVT \keys1_reg[66]  ( .D(n528), .CLK(clk), .Q(keys1[66]) );
  DFFX1_HVT \keys1_reg[67]  ( .D(n527), .CLK(clk), .Q(keys1[67]) );
  DFFX1_HVT \keys1_reg[68]  ( .D(n526), .CLK(clk), .Q(keys1[68]) );
  DFFX1_HVT \keys1_reg[69]  ( .D(n525), .CLK(clk), .Q(keys1[69]) );
  DFFX1_HVT \keys1_reg[70]  ( .D(n524), .CLK(clk), .Q(keys1[70]) );
  DFFX1_HVT \keys1_reg[71]  ( .D(n523), .CLK(clk), .Q(keys1[71]) );
  DFFX1_HVT \keys1_reg[72]  ( .D(n522), .CLK(clk), .Q(keys1[72]) );
  DFFX1_HVT \keys1_reg[73]  ( .D(n521), .CLK(clk), .Q(keys1[73]) );
  DFFX1_HVT \keys1_reg[74]  ( .D(n520), .CLK(clk), .Q(keys1[74]) );
  DFFX1_HVT \keys1_reg[75]  ( .D(n519), .CLK(clk), .Q(keys1[75]) );
  DFFX1_HVT \keys1_reg[76]  ( .D(n518), .CLK(clk), .Q(keys1[76]) );
  DFFX1_HVT \keys1_reg[77]  ( .D(n517), .CLK(clk), .Q(keys1[77]) );
  DFFX1_HVT \keys1_reg[78]  ( .D(n516), .CLK(clk), .Q(keys1[78]) );
  DFFX1_HVT \keys1_reg[79]  ( .D(n515), .CLK(clk), .Q(keys1[79]) );
  DFFX1_HVT \keys1_reg[80]  ( .D(n514), .CLK(clk), .Q(keys1[80]) );
  DFFX1_HVT \keys1_reg[81]  ( .D(n513), .CLK(clk), .Q(keys1[81]) );
  DFFX1_HVT \keys1_reg[82]  ( .D(n512), .CLK(clk), .Q(keys1[82]) );
  DFFX1_HVT \keys1_reg[83]  ( .D(n511), .CLK(clk), .Q(keys1[83]) );
  DFFX1_HVT \keys1_reg[84]  ( .D(n510), .CLK(clk), .Q(keys1[84]) );
  DFFX1_HVT \keys1_reg[85]  ( .D(n509), .CLK(clk), .Q(keys1[85]) );
  DFFX1_HVT \keys1_reg[86]  ( .D(n508), .CLK(clk), .Q(keys1[86]) );
  DFFX1_HVT \keys1_reg[87]  ( .D(n507), .CLK(clk), .Q(keys1[87]) );
  DFFX1_HVT \keys1_reg[88]  ( .D(n506), .CLK(clk), .Q(keys1[88]) );
  DFFX1_HVT \keys1_reg[89]  ( .D(n505), .CLK(clk), .Q(keys1[89]) );
  DFFX1_HVT \keys1_reg[90]  ( .D(n504), .CLK(clk), .Q(keys1[90]) );
  DFFX1_HVT \keys1_reg[91]  ( .D(n503), .CLK(clk), .Q(keys1[91]) );
  DFFX1_HVT \keys1_reg[92]  ( .D(n502), .CLK(clk), .Q(keys1[92]) );
  DFFX1_HVT \keys1_reg[93]  ( .D(n501), .CLK(clk), .Q(keys1[93]) );
  DFFX1_HVT \keys1_reg[94]  ( .D(n500), .CLK(clk), .Q(keys1[94]) );
  DFFX1_HVT \keys1_reg[95]  ( .D(n499), .CLK(clk), .Q(keys1[95]) );
  DFFX1_HVT \keys1_reg[96]  ( .D(n498), .CLK(clk), .Q(keys1[96]) );
  DFFX1_HVT \keys1_reg[97]  ( .D(n497), .CLK(clk), .Q(keys1[97]) );
  DFFX1_HVT \keys1_reg[98]  ( .D(n496), .CLK(clk), .Q(keys1[98]) );
  DFFX1_HVT \keys1_reg[99]  ( .D(n495), .CLK(clk), .Q(keys1[99]) );
  DFFX1_HVT \keys1_reg[100]  ( .D(n494), .CLK(clk), .Q(keys1[100]) );
  DFFX1_HVT \keys1_reg[101]  ( .D(n493), .CLK(clk), .Q(keys1[101]) );
  DFFX1_HVT \keys1_reg[102]  ( .D(n492), .CLK(clk), .Q(keys1[102]) );
  DFFX1_HVT \keys1_reg[103]  ( .D(n491), .CLK(clk), .Q(keys1[103]) );
  DFFX1_HVT \keys1_reg[104]  ( .D(n490), .CLK(clk), .Q(keys1[104]) );
  DFFX1_HVT \keys1_reg[105]  ( .D(n489), .CLK(clk), .Q(keys1[105]) );
  DFFX1_HVT \keys1_reg[106]  ( .D(n488), .CLK(clk), .Q(keys1[106]) );
  DFFX1_HVT \keys1_reg[107]  ( .D(n487), .CLK(clk), .Q(keys1[107]) );
  DFFX1_HVT \keys1_reg[108]  ( .D(n486), .CLK(clk), .Q(keys1[108]) );
  DFFX1_HVT \keys1_reg[109]  ( .D(n485), .CLK(clk), .Q(keys1[109]) );
  DFFX1_HVT \keys1_reg[110]  ( .D(n484), .CLK(clk), .Q(keys1[110]) );
  DFFX1_HVT \keys1_reg[111]  ( .D(n483), .CLK(clk), .Q(keys1[111]) );
  DFFX1_HVT \keys1_reg[112]  ( .D(n482), .CLK(clk), .Q(keys1[112]) );
  DFFX1_HVT \keys1_reg[113]  ( .D(n481), .CLK(clk), .Q(keys1[113]) );
  DFFX1_HVT \keys1_reg[114]  ( .D(n480), .CLK(clk), .Q(keys1[114]) );
  DFFX1_HVT \keys1_reg[115]  ( .D(n479), .CLK(clk), .Q(keys1[115]) );
  DFFX1_HVT \keys1_reg[116]  ( .D(n478), .CLK(clk), .Q(keys1[116]) );
  DFFX1_HVT \keys1_reg[117]  ( .D(n477), .CLK(clk), .Q(keys1[117]) );
  DFFX1_HVT \keys1_reg[118]  ( .D(n476), .CLK(clk), .Q(keys1[118]) );
  DFFX1_HVT \keys1_reg[119]  ( .D(n475), .CLK(clk), .Q(keys1[119]) );
  DFFX1_HVT \keys1_reg[120]  ( .D(n474), .CLK(clk), .Q(keys1[120]) );
  DFFX1_HVT \keys1_reg[121]  ( .D(n473), .CLK(clk), .Q(keys1[121]) );
  DFFX1_HVT \keys1_reg[122]  ( .D(n472), .CLK(clk), .Q(keys1[122]) );
  DFFX1_HVT \keys1_reg[123]  ( .D(n471), .CLK(clk), .Q(keys1[123]) );
  DFFX1_HVT \keys1_reg[124]  ( .D(n470), .CLK(clk), .Q(keys1[124]) );
  DFFX1_HVT \keys1_reg[125]  ( .D(n469), .CLK(clk), .Q(keys1[125]) );
  DFFX1_HVT \keys1_reg[126]  ( .D(n468), .CLK(clk), .Q(keys1[126]) );
  DFFX1_HVT \keys1_reg[127]  ( .D(n467), .CLK(clk), .Q(keys1[127]) );
  DFFARX1_HVT last_reg ( .D(n466), .CLK(clk), .RSTB(n5), .Q(last) );
  DFFX1_HVT \adk_out_reg[0]  ( .D(n465), .CLK(clk), .Q(adk_out[0]) );
  DFFARX1_HVT \cipher_text_reg[0]  ( .D(n464), .CLK(clk), .RSTB(n5), .Q(
        cipher_text[0]) );
  DFFARX1_HVT \cipher_text_reg[1]  ( .D(n463), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[1]) );
  DFFX1_HVT \adk_out_reg[1]  ( .D(n336), .CLK(clk), .Q(adk_out[1]) );
  DFFARX1_HVT \cipher_text_reg[2]  ( .D(n462), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[2]) );
  DFFX1_HVT \adk_out_reg[2]  ( .D(n335), .CLK(clk), .Q(adk_out[2]) );
  DFFARX1_HVT \cipher_text_reg[3]  ( .D(n461), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[3]) );
  DFFX1_HVT \adk_out_reg[3]  ( .D(n334), .CLK(clk), .Q(adk_out[3]) );
  DFFARX1_HVT \cipher_text_reg[4]  ( .D(n460), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[4]) );
  DFFX1_HVT \adk_out_reg[4]  ( .D(n333), .CLK(clk), .Q(adk_out[4]) );
  DFFARX1_HVT \cipher_text_reg[5]  ( .D(n459), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[5]) );
  DFFX1_HVT \adk_out_reg[5]  ( .D(n332), .CLK(clk), .Q(adk_out[5]) );
  DFFARX1_HVT \cipher_text_reg[6]  ( .D(n458), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[6]) );
  DFFX1_HVT \adk_out_reg[6]  ( .D(n331), .CLK(clk), .Q(adk_out[6]) );
  DFFARX1_HVT \cipher_text_reg[7]  ( .D(n457), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[7]) );
  DFFX1_HVT \adk_out_reg[7]  ( .D(n330), .CLK(clk), .Q(adk_out[7]) );
  DFFARX1_HVT \cipher_text_reg[8]  ( .D(n456), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[8]) );
  DFFX1_HVT \adk_out_reg[8]  ( .D(n329), .CLK(clk), .Q(adk_out[8]) );
  DFFARX1_HVT \cipher_text_reg[9]  ( .D(n455), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[9]) );
  DFFX1_HVT \adk_out_reg[9]  ( .D(n328), .CLK(clk), .Q(adk_out[9]) );
  DFFARX1_HVT \cipher_text_reg[10]  ( .D(n454), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[10]) );
  DFFX1_HVT \adk_out_reg[10]  ( .D(n327), .CLK(clk), .Q(adk_out[10]) );
  DFFARX1_HVT \cipher_text_reg[11]  ( .D(n453), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[11]) );
  DFFX1_HVT \adk_out_reg[11]  ( .D(n326), .CLK(clk), .Q(adk_out[11]) );
  DFFARX1_HVT \cipher_text_reg[12]  ( .D(n452), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[12]) );
  DFFX1_HVT \adk_out_reg[12]  ( .D(n325), .CLK(clk), .Q(adk_out[12]) );
  DFFARX1_HVT \cipher_text_reg[13]  ( .D(n451), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[13]) );
  DFFX1_HVT \adk_out_reg[13]  ( .D(n324), .CLK(clk), .Q(adk_out[13]) );
  DFFARX1_HVT \cipher_text_reg[14]  ( .D(n450), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[14]) );
  DFFX1_HVT \adk_out_reg[14]  ( .D(n323), .CLK(clk), .Q(adk_out[14]) );
  DFFARX1_HVT \cipher_text_reg[15]  ( .D(n449), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[15]) );
  DFFX1_HVT \adk_out_reg[15]  ( .D(n322), .CLK(clk), .Q(adk_out[15]) );
  DFFARX1_HVT \cipher_text_reg[16]  ( .D(n448), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[16]) );
  DFFX1_HVT \adk_out_reg[16]  ( .D(n321), .CLK(clk), .Q(adk_out[16]) );
  DFFARX1_HVT \cipher_text_reg[17]  ( .D(n447), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[17]) );
  DFFX1_HVT \adk_out_reg[17]  ( .D(n320), .CLK(clk), .Q(adk_out[17]) );
  DFFARX1_HVT \cipher_text_reg[18]  ( .D(n446), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[18]) );
  DFFX1_HVT \adk_out_reg[18]  ( .D(n319), .CLK(clk), .Q(adk_out[18]) );
  DFFARX1_HVT \cipher_text_reg[19]  ( .D(n445), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[19]) );
  DFFX1_HVT \adk_out_reg[19]  ( .D(n318), .CLK(clk), .Q(adk_out[19]) );
  DFFARX1_HVT \cipher_text_reg[20]  ( .D(n444), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[20]) );
  DFFX1_HVT \adk_out_reg[20]  ( .D(n317), .CLK(clk), .Q(adk_out[20]) );
  DFFARX1_HVT \cipher_text_reg[21]  ( .D(n443), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[21]) );
  DFFX1_HVT \adk_out_reg[21]  ( .D(n316), .CLK(clk), .Q(adk_out[21]) );
  DFFARX1_HVT \cipher_text_reg[22]  ( .D(n442), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[22]) );
  DFFX1_HVT \adk_out_reg[22]  ( .D(n315), .CLK(clk), .Q(adk_out[22]) );
  DFFARX1_HVT \cipher_text_reg[23]  ( .D(n441), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[23]) );
  DFFX1_HVT \adk_out_reg[23]  ( .D(n314), .CLK(clk), .Q(adk_out[23]) );
  DFFARX1_HVT \cipher_text_reg[24]  ( .D(n440), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[24]) );
  DFFX1_HVT \adk_out_reg[24]  ( .D(n313), .CLK(clk), .Q(adk_out[24]) );
  DFFARX1_HVT \cipher_text_reg[25]  ( .D(n439), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[25]) );
  DFFX1_HVT \adk_out_reg[25]  ( .D(n312), .CLK(clk), .Q(adk_out[25]) );
  DFFARX1_HVT \cipher_text_reg[26]  ( .D(n438), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[26]) );
  DFFX1_HVT \adk_out_reg[26]  ( .D(n311), .CLK(clk), .Q(adk_out[26]) );
  DFFARX1_HVT \cipher_text_reg[27]  ( .D(n437), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[27]) );
  DFFX1_HVT \adk_out_reg[27]  ( .D(n310), .CLK(clk), .Q(adk_out[27]) );
  DFFARX1_HVT \cipher_text_reg[28]  ( .D(n436), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[28]) );
  DFFX1_HVT \adk_out_reg[28]  ( .D(n309), .CLK(clk), .Q(adk_out[28]) );
  DFFARX1_HVT \cipher_text_reg[29]  ( .D(n435), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[29]) );
  DFFX1_HVT \adk_out_reg[29]  ( .D(n308), .CLK(clk), .Q(adk_out[29]) );
  DFFARX1_HVT \cipher_text_reg[30]  ( .D(n434), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[30]) );
  DFFX1_HVT \adk_out_reg[30]  ( .D(n307), .CLK(clk), .Q(adk_out[30]) );
  DFFARX1_HVT \cipher_text_reg[31]  ( .D(n433), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[31]) );
  DFFX1_HVT \adk_out_reg[31]  ( .D(n306), .CLK(clk), .Q(adk_out[31]) );
  DFFARX1_HVT \cipher_text_reg[32]  ( .D(n432), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[32]) );
  DFFX1_HVT \adk_out_reg[32]  ( .D(n305), .CLK(clk), .Q(adk_out[32]) );
  DFFARX1_HVT \cipher_text_reg[33]  ( .D(n431), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[33]) );
  DFFX1_HVT \adk_out_reg[33]  ( .D(n304), .CLK(clk), .Q(adk_out[33]) );
  DFFARX1_HVT \cipher_text_reg[34]  ( .D(n430), .CLK(clk), .RSTB(n15), .Q(
        cipher_text[34]) );
  DFFX1_HVT \adk_out_reg[34]  ( .D(n303), .CLK(clk), .Q(adk_out[34]) );
  DFFARX1_HVT \cipher_text_reg[35]  ( .D(n429), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[35]) );
  DFFX1_HVT \adk_out_reg[35]  ( .D(n302), .CLK(clk), .Q(adk_out[35]) );
  DFFARX1_HVT \cipher_text_reg[36]  ( .D(n428), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[36]) );
  DFFX1_HVT \adk_out_reg[36]  ( .D(n301), .CLK(clk), .Q(adk_out[36]) );
  DFFARX1_HVT \cipher_text_reg[37]  ( .D(n427), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[37]) );
  DFFX1_HVT \adk_out_reg[37]  ( .D(n300), .CLK(clk), .Q(adk_out[37]) );
  DFFARX1_HVT \cipher_text_reg[38]  ( .D(n426), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[38]) );
  DFFX1_HVT \adk_out_reg[38]  ( .D(n299), .CLK(clk), .Q(adk_out[38]) );
  DFFARX1_HVT \cipher_text_reg[39]  ( .D(n425), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[39]) );
  DFFX1_HVT \adk_out_reg[39]  ( .D(n298), .CLK(clk), .Q(adk_out[39]) );
  DFFARX1_HVT \cipher_text_reg[40]  ( .D(n424), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[40]) );
  DFFX1_HVT \adk_out_reg[40]  ( .D(n297), .CLK(clk), .Q(adk_out[40]) );
  DFFARX1_HVT \cipher_text_reg[41]  ( .D(n423), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[41]) );
  DFFX1_HVT \adk_out_reg[41]  ( .D(n296), .CLK(clk), .Q(adk_out[41]) );
  DFFARX1_HVT \cipher_text_reg[42]  ( .D(n422), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[42]) );
  DFFX1_HVT \adk_out_reg[42]  ( .D(n295), .CLK(clk), .Q(adk_out[42]) );
  DFFARX1_HVT \cipher_text_reg[43]  ( .D(n421), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[43]) );
  DFFX1_HVT \adk_out_reg[43]  ( .D(n294), .CLK(clk), .Q(adk_out[43]) );
  DFFARX1_HVT \cipher_text_reg[44]  ( .D(n420), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[44]) );
  DFFX1_HVT \adk_out_reg[44]  ( .D(n293), .CLK(clk), .Q(adk_out[44]) );
  DFFARX1_HVT \cipher_text_reg[45]  ( .D(n419), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[45]) );
  DFFX1_HVT \adk_out_reg[45]  ( .D(n292), .CLK(clk), .Q(adk_out[45]) );
  DFFARX1_HVT \cipher_text_reg[46]  ( .D(n418), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[46]) );
  DFFX1_HVT \adk_out_reg[46]  ( .D(n291), .CLK(clk), .Q(adk_out[46]) );
  DFFARX1_HVT \cipher_text_reg[47]  ( .D(n417), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[47]) );
  DFFX1_HVT \adk_out_reg[47]  ( .D(n290), .CLK(clk), .Q(adk_out[47]) );
  DFFARX1_HVT \cipher_text_reg[48]  ( .D(n416), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[48]) );
  DFFX1_HVT \adk_out_reg[48]  ( .D(n289), .CLK(clk), .Q(adk_out[48]) );
  DFFARX1_HVT \cipher_text_reg[49]  ( .D(n415), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[49]) );
  DFFX1_HVT \adk_out_reg[49]  ( .D(n288), .CLK(clk), .Q(adk_out[49]) );
  DFFARX1_HVT \cipher_text_reg[50]  ( .D(n414), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[50]) );
  DFFX1_HVT \adk_out_reg[50]  ( .D(n287), .CLK(clk), .Q(adk_out[50]) );
  DFFARX1_HVT \cipher_text_reg[51]  ( .D(n413), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[51]) );
  DFFX1_HVT \adk_out_reg[51]  ( .D(n286), .CLK(clk), .Q(adk_out[51]) );
  DFFARX1_HVT \cipher_text_reg[52]  ( .D(n412), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[52]) );
  DFFX1_HVT \adk_out_reg[52]  ( .D(n285), .CLK(clk), .Q(adk_out[52]) );
  DFFARX1_HVT \cipher_text_reg[53]  ( .D(n411), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[53]) );
  DFFX1_HVT \adk_out_reg[53]  ( .D(n284), .CLK(clk), .Q(adk_out[53]) );
  DFFARX1_HVT \cipher_text_reg[54]  ( .D(n410), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[54]) );
  DFFX1_HVT \adk_out_reg[54]  ( .D(n283), .CLK(clk), .Q(adk_out[54]) );
  DFFARX1_HVT \cipher_text_reg[55]  ( .D(n409), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[55]) );
  DFFX1_HVT \adk_out_reg[55]  ( .D(n282), .CLK(clk), .Q(adk_out[55]) );
  DFFARX1_HVT \cipher_text_reg[56]  ( .D(n408), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[56]) );
  DFFX1_HVT \adk_out_reg[56]  ( .D(n281), .CLK(clk), .Q(adk_out[56]) );
  DFFARX1_HVT \cipher_text_reg[57]  ( .D(n407), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[57]) );
  DFFX1_HVT \adk_out_reg[57]  ( .D(n280), .CLK(clk), .Q(adk_out[57]) );
  DFFARX1_HVT \cipher_text_reg[58]  ( .D(n406), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[58]) );
  DFFX1_HVT \adk_out_reg[58]  ( .D(n279), .CLK(clk), .Q(adk_out[58]) );
  DFFARX1_HVT \cipher_text_reg[59]  ( .D(n405), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[59]) );
  DFFX1_HVT \adk_out_reg[59]  ( .D(n278), .CLK(clk), .Q(adk_out[59]) );
  DFFARX1_HVT \cipher_text_reg[60]  ( .D(n404), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[60]) );
  DFFX1_HVT \adk_out_reg[60]  ( .D(n277), .CLK(clk), .Q(adk_out[60]) );
  DFFARX1_HVT \cipher_text_reg[61]  ( .D(n403), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[61]) );
  DFFX1_HVT \adk_out_reg[61]  ( .D(n276), .CLK(clk), .Q(adk_out[61]) );
  DFFARX1_HVT \cipher_text_reg[62]  ( .D(n402), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[62]) );
  DFFX1_HVT \adk_out_reg[62]  ( .D(n275), .CLK(clk), .Q(adk_out[62]) );
  DFFARX1_HVT \cipher_text_reg[63]  ( .D(n401), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[63]) );
  DFFX1_HVT \adk_out_reg[63]  ( .D(n274), .CLK(clk), .Q(adk_out[63]) );
  DFFARX1_HVT \cipher_text_reg[64]  ( .D(n400), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[64]) );
  DFFX1_HVT \adk_out_reg[64]  ( .D(n273), .CLK(clk), .Q(adk_out[64]) );
  DFFARX1_HVT \cipher_text_reg[65]  ( .D(n399), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[65]) );
  DFFX1_HVT \adk_out_reg[65]  ( .D(n272), .CLK(clk), .Q(adk_out[65]) );
  DFFARX1_HVT \cipher_text_reg[66]  ( .D(n398), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[66]) );
  DFFX1_HVT \adk_out_reg[66]  ( .D(n271), .CLK(clk), .Q(adk_out[66]) );
  DFFARX1_HVT \cipher_text_reg[67]  ( .D(n397), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[67]) );
  DFFX1_HVT \adk_out_reg[67]  ( .D(n270), .CLK(clk), .Q(adk_out[67]) );
  DFFARX1_HVT \cipher_text_reg[68]  ( .D(n396), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[68]) );
  DFFX1_HVT \adk_out_reg[68]  ( .D(n269), .CLK(clk), .Q(adk_out[68]) );
  DFFARX1_HVT \cipher_text_reg[69]  ( .D(n395), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[69]) );
  DFFX1_HVT \adk_out_reg[69]  ( .D(n268), .CLK(clk), .Q(adk_out[69]) );
  DFFARX1_HVT \cipher_text_reg[70]  ( .D(n394), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[70]) );
  DFFX1_HVT \adk_out_reg[70]  ( .D(n267), .CLK(clk), .Q(adk_out[70]) );
  DFFARX1_HVT \cipher_text_reg[71]  ( .D(n393), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[71]) );
  DFFX1_HVT \adk_out_reg[71]  ( .D(n266), .CLK(clk), .Q(adk_out[71]) );
  DFFARX1_HVT \cipher_text_reg[72]  ( .D(n392), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[72]) );
  DFFX1_HVT \adk_out_reg[72]  ( .D(n265), .CLK(clk), .Q(adk_out[72]) );
  DFFARX1_HVT \cipher_text_reg[73]  ( .D(n391), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[73]) );
  DFFX1_HVT \adk_out_reg[73]  ( .D(n264), .CLK(clk), .Q(adk_out[73]) );
  DFFARX1_HVT \cipher_text_reg[74]  ( .D(n390), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[74]) );
  DFFX1_HVT \adk_out_reg[74]  ( .D(n263), .CLK(clk), .Q(adk_out[74]) );
  DFFARX1_HVT \cipher_text_reg[75]  ( .D(n389), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[75]) );
  DFFX1_HVT \adk_out_reg[75]  ( .D(n262), .CLK(clk), .Q(adk_out[75]) );
  DFFARX1_HVT \cipher_text_reg[76]  ( .D(n388), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[76]) );
  DFFX1_HVT \adk_out_reg[76]  ( .D(n261), .CLK(clk), .Q(adk_out[76]) );
  DFFARX1_HVT \cipher_text_reg[77]  ( .D(n387), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[77]) );
  DFFX1_HVT \adk_out_reg[77]  ( .D(n260), .CLK(clk), .Q(adk_out[77]) );
  DFFARX1_HVT \cipher_text_reg[78]  ( .D(n386), .CLK(clk), .RSTB(n7), .Q(
        cipher_text[78]) );
  DFFX1_HVT \adk_out_reg[78]  ( .D(n259), .CLK(clk), .Q(adk_out[78]) );
  DFFARX1_HVT \cipher_text_reg[79]  ( .D(n385), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[79]) );
  DFFX1_HVT \adk_out_reg[79]  ( .D(n258), .CLK(clk), .Q(adk_out[79]) );
  DFFARX1_HVT \cipher_text_reg[80]  ( .D(n384), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[80]) );
  DFFX1_HVT \adk_out_reg[80]  ( .D(n257), .CLK(clk), .Q(adk_out[80]) );
  DFFARX1_HVT \cipher_text_reg[81]  ( .D(n383), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[81]) );
  DFFX1_HVT \adk_out_reg[81]  ( .D(n256), .CLK(clk), .Q(adk_out[81]) );
  DFFARX1_HVT \cipher_text_reg[82]  ( .D(n382), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[82]) );
  DFFX1_HVT \adk_out_reg[82]  ( .D(n255), .CLK(clk), .Q(adk_out[82]) );
  DFFARX1_HVT \cipher_text_reg[83]  ( .D(n381), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[83]) );
  DFFX1_HVT \adk_out_reg[83]  ( .D(n254), .CLK(clk), .Q(adk_out[83]) );
  DFFARX1_HVT \cipher_text_reg[84]  ( .D(n380), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[84]) );
  DFFX1_HVT \adk_out_reg[84]  ( .D(n253), .CLK(clk), .Q(adk_out[84]) );
  DFFARX1_HVT \cipher_text_reg[85]  ( .D(n379), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[85]) );
  DFFX1_HVT \adk_out_reg[85]  ( .D(n252), .CLK(clk), .Q(adk_out[85]) );
  DFFARX1_HVT \cipher_text_reg[86]  ( .D(n378), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[86]) );
  DFFX1_HVT \adk_out_reg[86]  ( .D(n251), .CLK(clk), .Q(adk_out[86]) );
  DFFARX1_HVT \cipher_text_reg[87]  ( .D(n377), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[87]) );
  DFFX1_HVT \adk_out_reg[87]  ( .D(n250), .CLK(clk), .Q(adk_out[87]) );
  DFFARX1_HVT \cipher_text_reg[88]  ( .D(n376), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[88]) );
  DFFX1_HVT \adk_out_reg[88]  ( .D(n249), .CLK(clk), .Q(adk_out[88]) );
  DFFARX1_HVT \cipher_text_reg[89]  ( .D(n375), .CLK(clk), .RSTB(n15), .Q(
        cipher_text[89]) );
  DFFX1_HVT \adk_out_reg[89]  ( .D(n248), .CLK(clk), .Q(adk_out[89]) );
  DFFARX1_HVT \cipher_text_reg[90]  ( .D(n374), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[90]) );
  DFFX1_HVT \adk_out_reg[90]  ( .D(n247), .CLK(clk), .Q(adk_out[90]) );
  DFFARX1_HVT \cipher_text_reg[91]  ( .D(n373), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[91]) );
  DFFX1_HVT \adk_out_reg[91]  ( .D(n246), .CLK(clk), .Q(adk_out[91]) );
  DFFARX1_HVT \cipher_text_reg[92]  ( .D(n372), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[92]) );
  DFFX1_HVT \adk_out_reg[92]  ( .D(n245), .CLK(clk), .Q(adk_out[92]) );
  DFFARX1_HVT \cipher_text_reg[93]  ( .D(n371), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[93]) );
  DFFX1_HVT \adk_out_reg[93]  ( .D(n244), .CLK(clk), .Q(adk_out[93]) );
  DFFARX1_HVT \cipher_text_reg[94]  ( .D(n370), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[94]) );
  DFFX1_HVT \adk_out_reg[94]  ( .D(n243), .CLK(clk), .Q(adk_out[94]) );
  DFFARX1_HVT \cipher_text_reg[95]  ( .D(n369), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[95]) );
  DFFX1_HVT \adk_out_reg[95]  ( .D(n242), .CLK(clk), .Q(adk_out[95]) );
  DFFARX1_HVT \cipher_text_reg[96]  ( .D(n368), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[96]) );
  DFFX1_HVT \adk_out_reg[96]  ( .D(n241), .CLK(clk), .Q(adk_out[96]) );
  DFFARX1_HVT \cipher_text_reg[97]  ( .D(n367), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[97]) );
  DFFX1_HVT \adk_out_reg[97]  ( .D(n240), .CLK(clk), .Q(adk_out[97]) );
  DFFARX1_HVT \cipher_text_reg[98]  ( .D(n366), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[98]) );
  DFFX1_HVT \adk_out_reg[98]  ( .D(n239), .CLK(clk), .Q(adk_out[98]) );
  DFFARX1_HVT \cipher_text_reg[99]  ( .D(n365), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[99]) );
  DFFX1_HVT \adk_out_reg[99]  ( .D(n238), .CLK(clk), .Q(adk_out[99]) );
  DFFARX1_HVT \cipher_text_reg[100]  ( .D(n364), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[100]) );
  DFFX1_HVT \adk_out_reg[100]  ( .D(n237), .CLK(clk), .Q(adk_out[100]) );
  DFFARX1_HVT \cipher_text_reg[101]  ( .D(n363), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[101]) );
  DFFX1_HVT \adk_out_reg[101]  ( .D(n236), .CLK(clk), .Q(adk_out[101]) );
  DFFARX1_HVT \cipher_text_reg[102]  ( .D(n362), .CLK(clk), .RSTB(n9), .Q(
        cipher_text[102]) );
  DFFX1_HVT \adk_out_reg[102]  ( .D(n235), .CLK(clk), .Q(adk_out[102]) );
  DFFARX1_HVT \cipher_text_reg[103]  ( .D(n361), .CLK(clk), .RSTB(n6), .Q(
        cipher_text[103]) );
  DFFX1_HVT \adk_out_reg[103]  ( .D(n234), .CLK(clk), .Q(adk_out[103]) );
  DFFARX1_HVT \cipher_text_reg[104]  ( .D(n360), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[104]) );
  DFFX1_HVT \adk_out_reg[104]  ( .D(n233), .CLK(clk), .Q(adk_out[104]) );
  DFFARX1_HVT \cipher_text_reg[105]  ( .D(n359), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[105]) );
  DFFX1_HVT \adk_out_reg[105]  ( .D(n232), .CLK(clk), .Q(adk_out[105]) );
  DFFARX1_HVT \cipher_text_reg[106]  ( .D(n358), .CLK(clk), .RSTB(n15), .Q(
        cipher_text[106]) );
  DFFX1_HVT \adk_out_reg[106]  ( .D(n231), .CLK(clk), .Q(adk_out[106]) );
  DFFARX1_HVT \cipher_text_reg[107]  ( .D(n357), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[107]) );
  DFFX1_HVT \adk_out_reg[107]  ( .D(n230), .CLK(clk), .Q(adk_out[107]) );
  DFFARX1_HVT \cipher_text_reg[108]  ( .D(n356), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[108]) );
  DFFX1_HVT \adk_out_reg[108]  ( .D(n229), .CLK(clk), .Q(adk_out[108]) );
  DFFARX1_HVT \cipher_text_reg[109]  ( .D(n355), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[109]) );
  DFFX1_HVT \adk_out_reg[109]  ( .D(n228), .CLK(clk), .Q(adk_out[109]) );
  DFFARX1_HVT \cipher_text_reg[110]  ( .D(n354), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[110]) );
  DFFX1_HVT \adk_out_reg[110]  ( .D(n227), .CLK(clk), .Q(adk_out[110]) );
  DFFARX1_HVT \cipher_text_reg[111]  ( .D(n353), .CLK(clk), .RSTB(n13), .Q(
        cipher_text[111]) );
  DFFX1_HVT \adk_out_reg[111]  ( .D(n226), .CLK(clk), .Q(adk_out[111]) );
  DFFARX1_HVT \cipher_text_reg[112]  ( .D(n352), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[112]) );
  DFFX1_HVT \adk_out_reg[112]  ( .D(n225), .CLK(clk), .Q(adk_out[112]) );
  DFFARX1_HVT \cipher_text_reg[113]  ( .D(n351), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[113]) );
  DFFX1_HVT \adk_out_reg[113]  ( .D(n224), .CLK(clk), .Q(adk_out[113]) );
  DFFARX1_HVT \cipher_text_reg[114]  ( .D(n350), .CLK(clk), .RSTB(n12), .Q(
        cipher_text[114]) );
  DFFX1_HVT \adk_out_reg[114]  ( .D(n223), .CLK(clk), .Q(adk_out[114]) );
  DFFARX1_HVT \cipher_text_reg[115]  ( .D(n349), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[115]) );
  DFFX1_HVT \adk_out_reg[115]  ( .D(n222), .CLK(clk), .Q(adk_out[115]) );
  DFFARX1_HVT \cipher_text_reg[116]  ( .D(n348), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[116]) );
  DFFX1_HVT \adk_out_reg[116]  ( .D(n221), .CLK(clk), .Q(adk_out[116]) );
  DFFARX1_HVT \cipher_text_reg[117]  ( .D(n347), .CLK(clk), .RSTB(n11), .Q(
        cipher_text[117]) );
  DFFX1_HVT \adk_out_reg[117]  ( .D(n220), .CLK(clk), .Q(adk_out[117]) );
  DFFARX1_HVT \cipher_text_reg[118]  ( .D(n346), .CLK(clk), .RSTB(n10), .Q(
        cipher_text[118]) );
  DFFX1_HVT \adk_out_reg[118]  ( .D(n219), .CLK(clk), .Q(adk_out[118]) );
  DFFARX1_HVT \cipher_text_reg[119]  ( .D(n345), .CLK(clk), .RSTB(n8), .Q(
        cipher_text[119]) );
  DFFX1_HVT \adk_out_reg[119]  ( .D(n218), .CLK(clk), .Q(adk_out[119]) );
  DFFARX1_HVT \cipher_text_reg[120]  ( .D(n344), .CLK(clk), .RSTB(n15), .Q(
        cipher_text[120]) );
  DFFX1_HVT \adk_out_reg[120]  ( .D(n217), .CLK(clk), .Q(adk_out[120]) );
  DFFARX1_HVT \cipher_text_reg[121]  ( .D(n343), .CLK(clk), .RSTB(n15), .Q(
        cipher_text[121]) );
  DFFX1_HVT \adk_out_reg[121]  ( .D(n216), .CLK(clk), .Q(adk_out[121]) );
  DFFARX1_HVT \cipher_text_reg[122]  ( .D(n342), .CLK(clk), .RSTB(n15), .Q(
        cipher_text[122]) );
  DFFX1_HVT \adk_out_reg[122]  ( .D(n215), .CLK(clk), .Q(adk_out[122]) );
  DFFARX1_HVT \cipher_text_reg[123]  ( .D(n341), .CLK(clk), .RSTB(n15), .Q(
        cipher_text[123]) );
  DFFX1_HVT \adk_out_reg[123]  ( .D(n214), .CLK(clk), .Q(adk_out[123]) );
  DFFARX1_HVT \cipher_text_reg[124]  ( .D(n340), .CLK(clk), .RSTB(n15), .Q(
        cipher_text[124]) );
  DFFX1_HVT \adk_out_reg[124]  ( .D(n213), .CLK(clk), .Q(adk_out[124]) );
  DFFARX1_HVT \cipher_text_reg[125]  ( .D(n339), .CLK(clk), .RSTB(n15), .Q(
        cipher_text[125]) );
  DFFX1_HVT \adk_out_reg[125]  ( .D(n212), .CLK(clk), .Q(adk_out[125]) );
  DFFARX1_HVT \cipher_text_reg[126]  ( .D(n338), .CLK(clk), .RSTB(n15), .Q(
        cipher_text[126]) );
  DFFX1_HVT \adk_out_reg[126]  ( .D(n211), .CLK(clk), .Q(adk_out[126]) );
  DFFARX1_HVT \cipher_text_reg[127]  ( .D(n337), .CLK(clk), .RSTB(n14), .Q(
        cipher_text[127]) );
  DFFX1_HVT \adk_out_reg[127]  ( .D(n210), .CLK(clk), .Q(adk_out[127]) );
  inv_round r1 ( .in(adk_out), .last(last), .keyin(keys1), .out(out1) );
  Get_key as1 ( .clk(clk), .rest(rest), .local_key(local_key), .rount_no(
        rount_no), .key_round(key_round), .done(done_k) );
  NBUFFX2_HVT U3 ( .A(n609), .Y(n5) );
  NBUFFX2_HVT U4 ( .A(n609), .Y(n14) );
  NBUFFX2_HVT U5 ( .A(n609), .Y(n11) );
  NBUFFX2_HVT U6 ( .A(n609), .Y(n12) );
  NBUFFX2_HVT U7 ( .A(n609), .Y(n8) );
  NBUFFX2_HVT U8 ( .A(n609), .Y(n7) );
  NBUFFX2_HVT U9 ( .A(n609), .Y(n10) );
  NBUFFX2_HVT U10 ( .A(n609), .Y(n6) );
  NBUFFX2_HVT U11 ( .A(n609), .Y(n9) );
  NBUFFX2_HVT U12 ( .A(n609), .Y(n13) );
  NBUFFX2_HVT U13 ( .A(n609), .Y(n15) );
  NAND2X0_HVT U14 ( .A1(n16), .A2(n17), .Y(n604) );
  NAND3X0_HVT U15 ( .A1(n18), .A2(busy), .A3(n19), .Y(n17) );
  AO21X1_HVT U16 ( .A1(n19), .A2(done), .A3(n20), .Y(n603) );
  NAND3X0_HVT U17 ( .A1(n21), .A2(n22), .A3(n23), .Y(n19) );
  AO221X1_HVT U18 ( .A1(n24), .A2(state[2]), .A3(n25), .A4(n26), .A5(n27), .Y(
        n602) );
  AO21X1_HVT U19 ( .A1(n22), .A2(n28), .A3(n20), .Y(n27) );
  NAND4X0_HVT U20 ( .A1(n29), .A2(n30), .A3(n31), .A4(n32), .Y(n28) );
  AO221X1_HVT U21 ( .A1(n22), .A2(n33), .A3(n24), .A4(state[3]), .A5(n34), .Y(
        n601) );
  OR2X1_HVT U22 ( .A1(n35), .A2(n36), .Y(n34) );
  NAND2X0_HVT U23 ( .A1(n37), .A2(n38), .Y(n33) );
  MUX21X1_HVT U24 ( .A1(n39), .A2(state[0]), .S0(n24), .Y(n600) );
  AO221X1_HVT U25 ( .A1(n22), .A2(n40), .A3(n25), .A4(done_k), .A5(n35), .Y(
        n39) );
  AO21X1_HVT U26 ( .A1(n22), .A2(n41), .A3(n20), .Y(n35) );
  NAND2X0_HVT U27 ( .A1(n42), .A2(n43), .Y(n41) );
  AO221X1_HVT U28 ( .A1(n22), .A2(n44), .A3(n24), .A4(state[1]), .A5(n25), .Y(
        n599) );
  AND3X1_HVT U29 ( .A1(n45), .A2(n18), .A3(n46), .Y(n24) );
  NAND2X0_HVT U30 ( .A1(n22), .A2(n47), .Y(n45) );
  NAND4X0_HVT U31 ( .A1(n48), .A2(n49), .A3(n50), .A4(n51), .Y(n47) );
  OR2X1_HVT U32 ( .A1(n26), .A2(n42), .Y(n49) );
  INVX0_HVT U33 ( .A(done_k), .Y(n26) );
  NAND3X0_HVT U34 ( .A1(n42), .A2(n52), .A3(n53), .Y(n44) );
  NAND2X0_HVT U35 ( .A1(n54), .A2(n55), .Y(n42) );
  AO22X1_HVT U36 ( .A1(rount_no[0]), .A2(n56), .A3(n22), .A4(n57), .Y(n598) );
  NAND2X0_HVT U37 ( .A1(n58), .A2(n32), .Y(n57) );
  AO221X1_HVT U38 ( .A1(n22), .A2(n59), .A3(rount_no[1]), .A4(n56), .A5(n25), 
        .Y(n597) );
  NAND2X0_HVT U39 ( .A1(n60), .A2(n29), .Y(n59) );
  AO22X1_HVT U40 ( .A1(rount_no[2]), .A2(n56), .A3(n22), .A4(n61), .Y(n596) );
  NAND3X0_HVT U41 ( .A1(n62), .A2(n31), .A3(n60), .Y(n61) );
  AND2X1_HVT U42 ( .A1(n63), .A2(n50), .Y(n60) );
  AO221X1_HVT U43 ( .A1(rount_no[3]), .A2(n56), .A3(n64), .A4(n22), .A5(n36), 
        .Y(n595) );
  INVX0_HVT U44 ( .A(n46), .Y(n36) );
  OA21X1_HVT U45 ( .A1(n32), .A2(n65), .A3(n16), .Y(n46) );
  AOI21X1_HVT U46 ( .A1(n22), .A2(n66), .A3(n25), .Y(n56) );
  NAND4X0_HVT U47 ( .A1(n51), .A2(n63), .A3(n58), .A4(n67), .Y(n66) );
  AND4X1_HVT U48 ( .A1(n38), .A2(n31), .A3(n52), .A4(n32), .Y(n67) );
  NAND2X0_HVT U49 ( .A1(n21), .A2(n68), .Y(n32) );
  MUX21X1_HVT U50 ( .A1(keys1[0]), .A2(key_round[0]), .S0(n69), .Y(n594) );
  MUX21X1_HVT U51 ( .A1(keys1[1]), .A2(key_round[1]), .S0(n69), .Y(n593) );
  MUX21X1_HVT U52 ( .A1(keys1[2]), .A2(key_round[2]), .S0(n69), .Y(n592) );
  MUX21X1_HVT U53 ( .A1(keys1[3]), .A2(key_round[3]), .S0(n69), .Y(n591) );
  MUX21X1_HVT U54 ( .A1(keys1[4]), .A2(key_round[4]), .S0(n69), .Y(n590) );
  MUX21X1_HVT U55 ( .A1(keys1[5]), .A2(key_round[5]), .S0(n69), .Y(n589) );
  MUX21X1_HVT U56 ( .A1(keys1[6]), .A2(key_round[6]), .S0(n69), .Y(n588) );
  MUX21X1_HVT U57 ( .A1(keys1[7]), .A2(key_round[7]), .S0(n69), .Y(n587) );
  MUX21X1_HVT U58 ( .A1(keys1[8]), .A2(key_round[8]), .S0(n69), .Y(n586) );
  MUX21X1_HVT U59 ( .A1(keys1[9]), .A2(key_round[9]), .S0(n69), .Y(n585) );
  MUX21X1_HVT U60 ( .A1(keys1[10]), .A2(key_round[10]), .S0(n69), .Y(n584) );
  MUX21X1_HVT U61 ( .A1(keys1[11]), .A2(key_round[11]), .S0(n69), .Y(n583) );
  MUX21X1_HVT U62 ( .A1(keys1[12]), .A2(key_round[12]), .S0(n69), .Y(n582) );
  MUX21X1_HVT U63 ( .A1(keys1[13]), .A2(key_round[13]), .S0(n69), .Y(n581) );
  MUX21X1_HVT U64 ( .A1(keys1[14]), .A2(key_round[14]), .S0(n69), .Y(n580) );
  MUX21X1_HVT U65 ( .A1(keys1[15]), .A2(key_round[15]), .S0(n69), .Y(n579) );
  MUX21X1_HVT U66 ( .A1(keys1[16]), .A2(key_round[16]), .S0(n69), .Y(n578) );
  MUX21X1_HVT U67 ( .A1(keys1[17]), .A2(key_round[17]), .S0(n69), .Y(n577) );
  MUX21X1_HVT U68 ( .A1(keys1[18]), .A2(key_round[18]), .S0(n69), .Y(n576) );
  MUX21X1_HVT U69 ( .A1(keys1[19]), .A2(key_round[19]), .S0(n69), .Y(n575) );
  MUX21X1_HVT U70 ( .A1(keys1[20]), .A2(key_round[20]), .S0(n69), .Y(n574) );
  MUX21X1_HVT U71 ( .A1(keys1[21]), .A2(key_round[21]), .S0(n69), .Y(n573) );
  MUX21X1_HVT U72 ( .A1(keys1[22]), .A2(key_round[22]), .S0(n69), .Y(n572) );
  MUX21X1_HVT U73 ( .A1(keys1[23]), .A2(key_round[23]), .S0(n69), .Y(n571) );
  MUX21X1_HVT U74 ( .A1(keys1[24]), .A2(key_round[24]), .S0(n69), .Y(n570) );
  MUX21X1_HVT U75 ( .A1(keys1[25]), .A2(key_round[25]), .S0(n69), .Y(n569) );
  MUX21X1_HVT U76 ( .A1(keys1[26]), .A2(key_round[26]), .S0(n69), .Y(n568) );
  MUX21X1_HVT U77 ( .A1(keys1[27]), .A2(key_round[27]), .S0(n69), .Y(n567) );
  MUX21X1_HVT U78 ( .A1(keys1[28]), .A2(key_round[28]), .S0(n69), .Y(n566) );
  MUX21X1_HVT U79 ( .A1(keys1[29]), .A2(key_round[29]), .S0(n69), .Y(n565) );
  MUX21X1_HVT U80 ( .A1(keys1[30]), .A2(key_round[30]), .S0(n69), .Y(n564) );
  MUX21X1_HVT U81 ( .A1(keys1[31]), .A2(key_round[31]), .S0(n69), .Y(n563) );
  MUX21X1_HVT U82 ( .A1(keys1[32]), .A2(key_round[32]), .S0(n69), .Y(n562) );
  MUX21X1_HVT U83 ( .A1(keys1[33]), .A2(key_round[33]), .S0(n69), .Y(n561) );
  MUX21X1_HVT U84 ( .A1(keys1[34]), .A2(key_round[34]), .S0(n69), .Y(n560) );
  MUX21X1_HVT U85 ( .A1(keys1[35]), .A2(key_round[35]), .S0(n69), .Y(n559) );
  MUX21X1_HVT U86 ( .A1(keys1[36]), .A2(key_round[36]), .S0(n69), .Y(n558) );
  MUX21X1_HVT U87 ( .A1(keys1[37]), .A2(key_round[37]), .S0(n69), .Y(n557) );
  MUX21X1_HVT U88 ( .A1(keys1[38]), .A2(key_round[38]), .S0(n69), .Y(n556) );
  MUX21X1_HVT U89 ( .A1(keys1[39]), .A2(key_round[39]), .S0(n69), .Y(n555) );
  MUX21X1_HVT U90 ( .A1(keys1[40]), .A2(key_round[40]), .S0(n69), .Y(n554) );
  MUX21X1_HVT U91 ( .A1(keys1[41]), .A2(key_round[41]), .S0(n69), .Y(n553) );
  MUX21X1_HVT U92 ( .A1(keys1[42]), .A2(key_round[42]), .S0(n69), .Y(n552) );
  MUX21X1_HVT U93 ( .A1(keys1[43]), .A2(key_round[43]), .S0(n69), .Y(n551) );
  MUX21X1_HVT U94 ( .A1(keys1[44]), .A2(key_round[44]), .S0(n69), .Y(n550) );
  MUX21X1_HVT U95 ( .A1(keys1[45]), .A2(key_round[45]), .S0(n69), .Y(n549) );
  MUX21X1_HVT U96 ( .A1(keys1[46]), .A2(key_round[46]), .S0(n69), .Y(n548) );
  MUX21X1_HVT U97 ( .A1(keys1[47]), .A2(key_round[47]), .S0(n69), .Y(n547) );
  MUX21X1_HVT U98 ( .A1(keys1[48]), .A2(key_round[48]), .S0(n69), .Y(n546) );
  MUX21X1_HVT U99 ( .A1(keys1[49]), .A2(key_round[49]), .S0(n69), .Y(n545) );
  MUX21X1_HVT U100 ( .A1(keys1[50]), .A2(key_round[50]), .S0(n69), .Y(n544) );
  MUX21X1_HVT U101 ( .A1(keys1[51]), .A2(key_round[51]), .S0(n69), .Y(n543) );
  MUX21X1_HVT U102 ( .A1(keys1[52]), .A2(key_round[52]), .S0(n69), .Y(n542) );
  MUX21X1_HVT U103 ( .A1(keys1[53]), .A2(key_round[53]), .S0(n69), .Y(n541) );
  MUX21X1_HVT U104 ( .A1(keys1[54]), .A2(key_round[54]), .S0(n69), .Y(n540) );
  MUX21X1_HVT U105 ( .A1(keys1[55]), .A2(key_round[55]), .S0(n69), .Y(n539) );
  MUX21X1_HVT U106 ( .A1(keys1[56]), .A2(key_round[56]), .S0(n69), .Y(n538) );
  MUX21X1_HVT U107 ( .A1(keys1[57]), .A2(key_round[57]), .S0(n69), .Y(n537) );
  MUX21X1_HVT U108 ( .A1(keys1[58]), .A2(key_round[58]), .S0(n69), .Y(n536) );
  MUX21X1_HVT U109 ( .A1(keys1[59]), .A2(key_round[59]), .S0(n69), .Y(n535) );
  MUX21X1_HVT U110 ( .A1(keys1[60]), .A2(key_round[60]), .S0(n69), .Y(n534) );
  MUX21X1_HVT U111 ( .A1(keys1[61]), .A2(key_round[61]), .S0(n69), .Y(n533) );
  MUX21X1_HVT U112 ( .A1(keys1[62]), .A2(key_round[62]), .S0(n69), .Y(n532) );
  MUX21X1_HVT U113 ( .A1(keys1[63]), .A2(key_round[63]), .S0(n69), .Y(n531) );
  MUX21X1_HVT U114 ( .A1(keys1[64]), .A2(key_round[64]), .S0(n69), .Y(n530) );
  MUX21X1_HVT U115 ( .A1(keys1[65]), .A2(key_round[65]), .S0(n69), .Y(n529) );
  MUX21X1_HVT U116 ( .A1(keys1[66]), .A2(key_round[66]), .S0(n69), .Y(n528) );
  MUX21X1_HVT U117 ( .A1(keys1[67]), .A2(key_round[67]), .S0(n69), .Y(n527) );
  MUX21X1_HVT U118 ( .A1(keys1[68]), .A2(key_round[68]), .S0(n69), .Y(n526) );
  MUX21X1_HVT U119 ( .A1(keys1[69]), .A2(key_round[69]), .S0(n69), .Y(n525) );
  MUX21X1_HVT U120 ( .A1(keys1[70]), .A2(key_round[70]), .S0(n69), .Y(n524) );
  MUX21X1_HVT U121 ( .A1(keys1[71]), .A2(key_round[71]), .S0(n69), .Y(n523) );
  MUX21X1_HVT U122 ( .A1(keys1[72]), .A2(key_round[72]), .S0(n69), .Y(n522) );
  MUX21X1_HVT U123 ( .A1(keys1[73]), .A2(key_round[73]), .S0(n69), .Y(n521) );
  MUX21X1_HVT U124 ( .A1(keys1[74]), .A2(key_round[74]), .S0(n69), .Y(n520) );
  MUX21X1_HVT U125 ( .A1(keys1[75]), .A2(key_round[75]), .S0(n69), .Y(n519) );
  MUX21X1_HVT U126 ( .A1(keys1[76]), .A2(key_round[76]), .S0(n69), .Y(n518) );
  MUX21X1_HVT U127 ( .A1(keys1[77]), .A2(key_round[77]), .S0(n69), .Y(n517) );
  MUX21X1_HVT U128 ( .A1(keys1[78]), .A2(key_round[78]), .S0(n69), .Y(n516) );
  MUX21X1_HVT U129 ( .A1(keys1[79]), .A2(key_round[79]), .S0(n69), .Y(n515) );
  MUX21X1_HVT U130 ( .A1(keys1[80]), .A2(key_round[80]), .S0(n69), .Y(n514) );
  MUX21X1_HVT U131 ( .A1(keys1[81]), .A2(key_round[81]), .S0(n69), .Y(n513) );
  MUX21X1_HVT U132 ( .A1(keys1[82]), .A2(key_round[82]), .S0(n69), .Y(n512) );
  MUX21X1_HVT U133 ( .A1(keys1[83]), .A2(key_round[83]), .S0(n69), .Y(n511) );
  MUX21X1_HVT U134 ( .A1(keys1[84]), .A2(key_round[84]), .S0(n69), .Y(n510) );
  MUX21X1_HVT U135 ( .A1(keys1[85]), .A2(key_round[85]), .S0(n69), .Y(n509) );
  MUX21X1_HVT U136 ( .A1(keys1[86]), .A2(key_round[86]), .S0(n69), .Y(n508) );
  MUX21X1_HVT U137 ( .A1(keys1[87]), .A2(key_round[87]), .S0(n69), .Y(n507) );
  MUX21X1_HVT U138 ( .A1(keys1[88]), .A2(key_round[88]), .S0(n69), .Y(n506) );
  MUX21X1_HVT U139 ( .A1(keys1[89]), .A2(key_round[89]), .S0(n69), .Y(n505) );
  MUX21X1_HVT U140 ( .A1(keys1[90]), .A2(key_round[90]), .S0(n69), .Y(n504) );
  MUX21X1_HVT U141 ( .A1(keys1[91]), .A2(key_round[91]), .S0(n69), .Y(n503) );
  MUX21X1_HVT U142 ( .A1(keys1[92]), .A2(key_round[92]), .S0(n69), .Y(n502) );
  MUX21X1_HVT U143 ( .A1(keys1[93]), .A2(key_round[93]), .S0(n69), .Y(n501) );
  MUX21X1_HVT U144 ( .A1(keys1[94]), .A2(key_round[94]), .S0(n69), .Y(n500) );
  MUX21X1_HVT U145 ( .A1(keys1[95]), .A2(key_round[95]), .S0(n69), .Y(n499) );
  MUX21X1_HVT U146 ( .A1(keys1[96]), .A2(key_round[96]), .S0(n69), .Y(n498) );
  MUX21X1_HVT U147 ( .A1(keys1[97]), .A2(key_round[97]), .S0(n69), .Y(n497) );
  MUX21X1_HVT U148 ( .A1(keys1[98]), .A2(key_round[98]), .S0(n69), .Y(n496) );
  MUX21X1_HVT U149 ( .A1(keys1[99]), .A2(key_round[99]), .S0(n69), .Y(n495) );
  MUX21X1_HVT U150 ( .A1(keys1[100]), .A2(key_round[100]), .S0(n69), .Y(n494)
         );
  MUX21X1_HVT U151 ( .A1(keys1[101]), .A2(key_round[101]), .S0(n69), .Y(n493)
         );
  MUX21X1_HVT U152 ( .A1(keys1[102]), .A2(key_round[102]), .S0(n69), .Y(n492)
         );
  MUX21X1_HVT U153 ( .A1(keys1[103]), .A2(key_round[103]), .S0(n69), .Y(n491)
         );
  MUX21X1_HVT U154 ( .A1(keys1[104]), .A2(key_round[104]), .S0(n69), .Y(n490)
         );
  MUX21X1_HVT U155 ( .A1(keys1[105]), .A2(key_round[105]), .S0(n69), .Y(n489)
         );
  MUX21X1_HVT U156 ( .A1(keys1[106]), .A2(key_round[106]), .S0(n69), .Y(n488)
         );
  MUX21X1_HVT U157 ( .A1(keys1[107]), .A2(key_round[107]), .S0(n69), .Y(n487)
         );
  MUX21X1_HVT U158 ( .A1(keys1[108]), .A2(key_round[108]), .S0(n69), .Y(n486)
         );
  MUX21X1_HVT U159 ( .A1(keys1[109]), .A2(key_round[109]), .S0(n69), .Y(n485)
         );
  MUX21X1_HVT U160 ( .A1(keys1[110]), .A2(key_round[110]), .S0(n69), .Y(n484)
         );
  MUX21X1_HVT U161 ( .A1(keys1[111]), .A2(key_round[111]), .S0(n69), .Y(n483)
         );
  MUX21X1_HVT U162 ( .A1(keys1[112]), .A2(key_round[112]), .S0(n69), .Y(n482)
         );
  MUX21X1_HVT U163 ( .A1(keys1[113]), .A2(key_round[113]), .S0(n69), .Y(n481)
         );
  MUX21X1_HVT U164 ( .A1(keys1[114]), .A2(key_round[114]), .S0(n69), .Y(n480)
         );
  MUX21X1_HVT U165 ( .A1(keys1[115]), .A2(key_round[115]), .S0(n69), .Y(n479)
         );
  MUX21X1_HVT U166 ( .A1(keys1[116]), .A2(key_round[116]), .S0(n69), .Y(n478)
         );
  MUX21X1_HVT U167 ( .A1(keys1[117]), .A2(key_round[117]), .S0(n69), .Y(n477)
         );
  MUX21X1_HVT U168 ( .A1(keys1[118]), .A2(key_round[118]), .S0(n69), .Y(n476)
         );
  MUX21X1_HVT U169 ( .A1(keys1[119]), .A2(key_round[119]), .S0(n69), .Y(n475)
         );
  MUX21X1_HVT U170 ( .A1(keys1[120]), .A2(key_round[120]), .S0(n69), .Y(n474)
         );
  MUX21X1_HVT U171 ( .A1(keys1[121]), .A2(key_round[121]), .S0(n69), .Y(n473)
         );
  MUX21X1_HVT U172 ( .A1(keys1[122]), .A2(key_round[122]), .S0(n69), .Y(n472)
         );
  MUX21X1_HVT U173 ( .A1(keys1[123]), .A2(key_round[123]), .S0(n69), .Y(n471)
         );
  MUX21X1_HVT U174 ( .A1(keys1[124]), .A2(key_round[124]), .S0(n69), .Y(n470)
         );
  MUX21X1_HVT U175 ( .A1(keys1[125]), .A2(key_round[125]), .S0(n69), .Y(n469)
         );
  MUX21X1_HVT U176 ( .A1(keys1[126]), .A2(key_round[126]), .S0(n69), .Y(n468)
         );
  MUX21X1_HVT U177 ( .A1(keys1[127]), .A2(key_round[127]), .S0(n69), .Y(n467)
         );
  AND3X1_HVT U178 ( .A1(n70), .A2(n15), .A3(n22), .Y(n69) );
  NAND2X0_HVT U179 ( .A1(n48), .A2(n50), .Y(n70) );
  NAND2X0_HVT U180 ( .A1(n71), .A2(n40), .Y(n50) );
  AO22X1_HVT U181 ( .A1(n16), .A2(last), .A3(n72), .A4(n22), .Y(n466) );
  INVX0_HVT U182 ( .A(n37), .Y(n72) );
  AO222X1_HVT U183 ( .A1(out1[0]), .A2(n73), .A3(n74), .A4(n75), .A5(n76), 
        .A6(adk_out[0]), .Y(n465) );
  XOR2X1_HVT U184 ( .A1(plaintext1[0]), .A2(key_round[0]), .Y(n75) );
  MUX21X1_HVT U185 ( .A1(cipher_text[0]), .A2(out1[0]), .S0(n20), .Y(n464) );
  MUX21X1_HVT U186 ( .A1(cipher_text[1]), .A2(out1[1]), .S0(n20), .Y(n463) );
  MUX21X1_HVT U187 ( .A1(cipher_text[2]), .A2(out1[2]), .S0(n20), .Y(n462) );
  MUX21X1_HVT U188 ( .A1(cipher_text[3]), .A2(out1[3]), .S0(n20), .Y(n461) );
  MUX21X1_HVT U189 ( .A1(cipher_text[4]), .A2(out1[4]), .S0(n20), .Y(n460) );
  MUX21X1_HVT U190 ( .A1(cipher_text[5]), .A2(out1[5]), .S0(n20), .Y(n459) );
  MUX21X1_HVT U191 ( .A1(cipher_text[6]), .A2(out1[6]), .S0(n20), .Y(n458) );
  MUX21X1_HVT U192 ( .A1(cipher_text[7]), .A2(out1[7]), .S0(n20), .Y(n457) );
  MUX21X1_HVT U193 ( .A1(cipher_text[8]), .A2(out1[8]), .S0(n20), .Y(n456) );
  MUX21X1_HVT U194 ( .A1(cipher_text[9]), .A2(out1[9]), .S0(n20), .Y(n455) );
  MUX21X1_HVT U195 ( .A1(cipher_text[10]), .A2(out1[10]), .S0(n20), .Y(n454)
         );
  MUX21X1_HVT U196 ( .A1(cipher_text[11]), .A2(out1[11]), .S0(n20), .Y(n453)
         );
  MUX21X1_HVT U197 ( .A1(cipher_text[12]), .A2(out1[12]), .S0(n20), .Y(n452)
         );
  MUX21X1_HVT U198 ( .A1(cipher_text[13]), .A2(out1[13]), .S0(n20), .Y(n451)
         );
  MUX21X1_HVT U199 ( .A1(cipher_text[14]), .A2(out1[14]), .S0(n20), .Y(n450)
         );
  MUX21X1_HVT U200 ( .A1(cipher_text[15]), .A2(out1[15]), .S0(n20), .Y(n449)
         );
  MUX21X1_HVT U201 ( .A1(cipher_text[16]), .A2(out1[16]), .S0(n20), .Y(n448)
         );
  MUX21X1_HVT U202 ( .A1(cipher_text[17]), .A2(out1[17]), .S0(n20), .Y(n447)
         );
  MUX21X1_HVT U203 ( .A1(cipher_text[18]), .A2(out1[18]), .S0(n20), .Y(n446)
         );
  MUX21X1_HVT U204 ( .A1(cipher_text[19]), .A2(out1[19]), .S0(n20), .Y(n445)
         );
  MUX21X1_HVT U205 ( .A1(cipher_text[20]), .A2(out1[20]), .S0(n20), .Y(n444)
         );
  MUX21X1_HVT U206 ( .A1(cipher_text[21]), .A2(out1[21]), .S0(n20), .Y(n443)
         );
  MUX21X1_HVT U207 ( .A1(cipher_text[22]), .A2(out1[22]), .S0(n20), .Y(n442)
         );
  MUX21X1_HVT U208 ( .A1(cipher_text[23]), .A2(out1[23]), .S0(n20), .Y(n441)
         );
  MUX21X1_HVT U209 ( .A1(cipher_text[24]), .A2(out1[24]), .S0(n20), .Y(n440)
         );
  MUX21X1_HVT U210 ( .A1(cipher_text[25]), .A2(out1[25]), .S0(n20), .Y(n439)
         );
  MUX21X1_HVT U211 ( .A1(cipher_text[26]), .A2(out1[26]), .S0(n20), .Y(n438)
         );
  MUX21X1_HVT U212 ( .A1(cipher_text[27]), .A2(out1[27]), .S0(n20), .Y(n437)
         );
  MUX21X1_HVT U213 ( .A1(cipher_text[28]), .A2(out1[28]), .S0(n20), .Y(n436)
         );
  MUX21X1_HVT U214 ( .A1(cipher_text[29]), .A2(out1[29]), .S0(n20), .Y(n435)
         );
  MUX21X1_HVT U215 ( .A1(cipher_text[30]), .A2(out1[30]), .S0(n20), .Y(n434)
         );
  MUX21X1_HVT U216 ( .A1(cipher_text[31]), .A2(out1[31]), .S0(n20), .Y(n433)
         );
  MUX21X1_HVT U217 ( .A1(cipher_text[32]), .A2(out1[32]), .S0(n20), .Y(n432)
         );
  MUX21X1_HVT U218 ( .A1(cipher_text[33]), .A2(out1[33]), .S0(n20), .Y(n431)
         );
  MUX21X1_HVT U219 ( .A1(cipher_text[34]), .A2(out1[34]), .S0(n20), .Y(n430)
         );
  MUX21X1_HVT U220 ( .A1(cipher_text[35]), .A2(out1[35]), .S0(n20), .Y(n429)
         );
  MUX21X1_HVT U221 ( .A1(cipher_text[36]), .A2(out1[36]), .S0(n20), .Y(n428)
         );
  MUX21X1_HVT U222 ( .A1(cipher_text[37]), .A2(out1[37]), .S0(n20), .Y(n427)
         );
  MUX21X1_HVT U223 ( .A1(cipher_text[38]), .A2(out1[38]), .S0(n20), .Y(n426)
         );
  MUX21X1_HVT U224 ( .A1(cipher_text[39]), .A2(out1[39]), .S0(n20), .Y(n425)
         );
  MUX21X1_HVT U225 ( .A1(cipher_text[40]), .A2(out1[40]), .S0(n20), .Y(n424)
         );
  MUX21X1_HVT U226 ( .A1(cipher_text[41]), .A2(out1[41]), .S0(n20), .Y(n423)
         );
  MUX21X1_HVT U227 ( .A1(cipher_text[42]), .A2(out1[42]), .S0(n20), .Y(n422)
         );
  MUX21X1_HVT U228 ( .A1(cipher_text[43]), .A2(out1[43]), .S0(n20), .Y(n421)
         );
  MUX21X1_HVT U229 ( .A1(cipher_text[44]), .A2(out1[44]), .S0(n20), .Y(n420)
         );
  MUX21X1_HVT U230 ( .A1(cipher_text[45]), .A2(out1[45]), .S0(n20), .Y(n419)
         );
  MUX21X1_HVT U231 ( .A1(cipher_text[46]), .A2(out1[46]), .S0(n20), .Y(n418)
         );
  MUX21X1_HVT U232 ( .A1(cipher_text[47]), .A2(out1[47]), .S0(n20), .Y(n417)
         );
  MUX21X1_HVT U233 ( .A1(cipher_text[48]), .A2(out1[48]), .S0(n20), .Y(n416)
         );
  MUX21X1_HVT U234 ( .A1(cipher_text[49]), .A2(out1[49]), .S0(n20), .Y(n415)
         );
  MUX21X1_HVT U235 ( .A1(cipher_text[50]), .A2(out1[50]), .S0(n20), .Y(n414)
         );
  MUX21X1_HVT U236 ( .A1(cipher_text[51]), .A2(out1[51]), .S0(n20), .Y(n413)
         );
  MUX21X1_HVT U237 ( .A1(cipher_text[52]), .A2(out1[52]), .S0(n20), .Y(n412)
         );
  MUX21X1_HVT U238 ( .A1(cipher_text[53]), .A2(out1[53]), .S0(n20), .Y(n411)
         );
  MUX21X1_HVT U239 ( .A1(cipher_text[54]), .A2(out1[54]), .S0(n20), .Y(n410)
         );
  MUX21X1_HVT U240 ( .A1(cipher_text[55]), .A2(out1[55]), .S0(n20), .Y(n409)
         );
  MUX21X1_HVT U241 ( .A1(cipher_text[56]), .A2(out1[56]), .S0(n20), .Y(n408)
         );
  MUX21X1_HVT U242 ( .A1(cipher_text[57]), .A2(out1[57]), .S0(n20), .Y(n407)
         );
  MUX21X1_HVT U243 ( .A1(cipher_text[58]), .A2(out1[58]), .S0(n20), .Y(n406)
         );
  MUX21X1_HVT U244 ( .A1(cipher_text[59]), .A2(out1[59]), .S0(n20), .Y(n405)
         );
  MUX21X1_HVT U245 ( .A1(cipher_text[60]), .A2(out1[60]), .S0(n20), .Y(n404)
         );
  MUX21X1_HVT U246 ( .A1(cipher_text[61]), .A2(out1[61]), .S0(n20), .Y(n403)
         );
  MUX21X1_HVT U247 ( .A1(cipher_text[62]), .A2(out1[62]), .S0(n20), .Y(n402)
         );
  MUX21X1_HVT U248 ( .A1(cipher_text[63]), .A2(out1[63]), .S0(n20), .Y(n401)
         );
  MUX21X1_HVT U249 ( .A1(cipher_text[64]), .A2(out1[64]), .S0(n20), .Y(n400)
         );
  MUX21X1_HVT U250 ( .A1(cipher_text[65]), .A2(out1[65]), .S0(n20), .Y(n399)
         );
  MUX21X1_HVT U251 ( .A1(cipher_text[66]), .A2(out1[66]), .S0(n20), .Y(n398)
         );
  MUX21X1_HVT U252 ( .A1(cipher_text[67]), .A2(out1[67]), .S0(n20), .Y(n397)
         );
  MUX21X1_HVT U253 ( .A1(cipher_text[68]), .A2(out1[68]), .S0(n20), .Y(n396)
         );
  MUX21X1_HVT U254 ( .A1(cipher_text[69]), .A2(out1[69]), .S0(n20), .Y(n395)
         );
  MUX21X1_HVT U255 ( .A1(cipher_text[70]), .A2(out1[70]), .S0(n20), .Y(n394)
         );
  MUX21X1_HVT U256 ( .A1(cipher_text[71]), .A2(out1[71]), .S0(n20), .Y(n393)
         );
  MUX21X1_HVT U257 ( .A1(cipher_text[72]), .A2(out1[72]), .S0(n20), .Y(n392)
         );
  MUX21X1_HVT U258 ( .A1(cipher_text[73]), .A2(out1[73]), .S0(n20), .Y(n391)
         );
  MUX21X1_HVT U259 ( .A1(cipher_text[74]), .A2(out1[74]), .S0(n20), .Y(n390)
         );
  MUX21X1_HVT U260 ( .A1(cipher_text[75]), .A2(out1[75]), .S0(n20), .Y(n389)
         );
  MUX21X1_HVT U261 ( .A1(cipher_text[76]), .A2(out1[76]), .S0(n20), .Y(n388)
         );
  MUX21X1_HVT U262 ( .A1(cipher_text[77]), .A2(out1[77]), .S0(n20), .Y(n387)
         );
  MUX21X1_HVT U263 ( .A1(cipher_text[78]), .A2(out1[78]), .S0(n20), .Y(n386)
         );
  MUX21X1_HVT U264 ( .A1(cipher_text[79]), .A2(out1[79]), .S0(n20), .Y(n385)
         );
  MUX21X1_HVT U265 ( .A1(cipher_text[80]), .A2(out1[80]), .S0(n20), .Y(n384)
         );
  MUX21X1_HVT U266 ( .A1(cipher_text[81]), .A2(out1[81]), .S0(n20), .Y(n383)
         );
  MUX21X1_HVT U267 ( .A1(cipher_text[82]), .A2(out1[82]), .S0(n20), .Y(n382)
         );
  MUX21X1_HVT U268 ( .A1(cipher_text[83]), .A2(out1[83]), .S0(n20), .Y(n381)
         );
  MUX21X1_HVT U269 ( .A1(cipher_text[84]), .A2(out1[84]), .S0(n20), .Y(n380)
         );
  MUX21X1_HVT U270 ( .A1(cipher_text[85]), .A2(out1[85]), .S0(n20), .Y(n379)
         );
  MUX21X1_HVT U271 ( .A1(cipher_text[86]), .A2(out1[86]), .S0(n20), .Y(n378)
         );
  MUX21X1_HVT U272 ( .A1(cipher_text[87]), .A2(out1[87]), .S0(n20), .Y(n377)
         );
  MUX21X1_HVT U273 ( .A1(cipher_text[88]), .A2(out1[88]), .S0(n20), .Y(n376)
         );
  MUX21X1_HVT U274 ( .A1(cipher_text[89]), .A2(out1[89]), .S0(n20), .Y(n375)
         );
  MUX21X1_HVT U275 ( .A1(cipher_text[90]), .A2(out1[90]), .S0(n20), .Y(n374)
         );
  MUX21X1_HVT U276 ( .A1(cipher_text[91]), .A2(out1[91]), .S0(n20), .Y(n373)
         );
  MUX21X1_HVT U277 ( .A1(cipher_text[92]), .A2(out1[92]), .S0(n20), .Y(n372)
         );
  MUX21X1_HVT U278 ( .A1(cipher_text[93]), .A2(out1[93]), .S0(n20), .Y(n371)
         );
  MUX21X1_HVT U279 ( .A1(cipher_text[94]), .A2(out1[94]), .S0(n20), .Y(n370)
         );
  MUX21X1_HVT U280 ( .A1(cipher_text[95]), .A2(out1[95]), .S0(n20), .Y(n369)
         );
  MUX21X1_HVT U281 ( .A1(cipher_text[96]), .A2(out1[96]), .S0(n20), .Y(n368)
         );
  MUX21X1_HVT U282 ( .A1(cipher_text[97]), .A2(out1[97]), .S0(n20), .Y(n367)
         );
  MUX21X1_HVT U283 ( .A1(cipher_text[98]), .A2(out1[98]), .S0(n20), .Y(n366)
         );
  MUX21X1_HVT U284 ( .A1(cipher_text[99]), .A2(out1[99]), .S0(n20), .Y(n365)
         );
  MUX21X1_HVT U285 ( .A1(cipher_text[100]), .A2(out1[100]), .S0(n20), .Y(n364)
         );
  MUX21X1_HVT U286 ( .A1(cipher_text[101]), .A2(out1[101]), .S0(n20), .Y(n363)
         );
  MUX21X1_HVT U287 ( .A1(cipher_text[102]), .A2(out1[102]), .S0(n20), .Y(n362)
         );
  MUX21X1_HVT U288 ( .A1(cipher_text[103]), .A2(out1[103]), .S0(n20), .Y(n361)
         );
  MUX21X1_HVT U289 ( .A1(cipher_text[104]), .A2(out1[104]), .S0(n20), .Y(n360)
         );
  MUX21X1_HVT U290 ( .A1(cipher_text[105]), .A2(out1[105]), .S0(n20), .Y(n359)
         );
  MUX21X1_HVT U291 ( .A1(cipher_text[106]), .A2(out1[106]), .S0(n20), .Y(n358)
         );
  MUX21X1_HVT U292 ( .A1(cipher_text[107]), .A2(out1[107]), .S0(n20), .Y(n357)
         );
  MUX21X1_HVT U293 ( .A1(cipher_text[108]), .A2(out1[108]), .S0(n20), .Y(n356)
         );
  MUX21X1_HVT U294 ( .A1(cipher_text[109]), .A2(out1[109]), .S0(n20), .Y(n355)
         );
  MUX21X1_HVT U295 ( .A1(cipher_text[110]), .A2(out1[110]), .S0(n20), .Y(n354)
         );
  MUX21X1_HVT U296 ( .A1(cipher_text[111]), .A2(out1[111]), .S0(n20), .Y(n353)
         );
  MUX21X1_HVT U297 ( .A1(cipher_text[112]), .A2(out1[112]), .S0(n20), .Y(n352)
         );
  MUX21X1_HVT U298 ( .A1(cipher_text[113]), .A2(out1[113]), .S0(n20), .Y(n351)
         );
  MUX21X1_HVT U299 ( .A1(cipher_text[114]), .A2(out1[114]), .S0(n20), .Y(n350)
         );
  MUX21X1_HVT U300 ( .A1(cipher_text[115]), .A2(out1[115]), .S0(n20), .Y(n349)
         );
  MUX21X1_HVT U301 ( .A1(cipher_text[116]), .A2(out1[116]), .S0(n20), .Y(n348)
         );
  MUX21X1_HVT U302 ( .A1(cipher_text[117]), .A2(out1[117]), .S0(n20), .Y(n347)
         );
  MUX21X1_HVT U303 ( .A1(cipher_text[118]), .A2(out1[118]), .S0(n20), .Y(n346)
         );
  MUX21X1_HVT U304 ( .A1(cipher_text[119]), .A2(out1[119]), .S0(n20), .Y(n345)
         );
  MUX21X1_HVT U305 ( .A1(cipher_text[120]), .A2(out1[120]), .S0(n20), .Y(n344)
         );
  MUX21X1_HVT U306 ( .A1(cipher_text[121]), .A2(out1[121]), .S0(n20), .Y(n343)
         );
  MUX21X1_HVT U307 ( .A1(cipher_text[122]), .A2(out1[122]), .S0(n20), .Y(n342)
         );
  MUX21X1_HVT U308 ( .A1(cipher_text[123]), .A2(out1[123]), .S0(n20), .Y(n341)
         );
  MUX21X1_HVT U309 ( .A1(cipher_text[124]), .A2(out1[124]), .S0(n20), .Y(n340)
         );
  MUX21X1_HVT U310 ( .A1(cipher_text[125]), .A2(out1[125]), .S0(n20), .Y(n339)
         );
  MUX21X1_HVT U311 ( .A1(cipher_text[126]), .A2(out1[126]), .S0(n20), .Y(n338)
         );
  MUX21X1_HVT U312 ( .A1(cipher_text[127]), .A2(out1[127]), .S0(n20), .Y(n337)
         );
  INVX0_HVT U313 ( .A(n18), .Y(n20) );
  NAND3X0_HVT U314 ( .A1(n68), .A2(n55), .A3(n22), .Y(n18) );
  AO222X1_HVT U315 ( .A1(out1[1]), .A2(n73), .A3(n74), .A4(n77), .A5(n76), 
        .A6(adk_out[1]), .Y(n336) );
  XOR2X1_HVT U316 ( .A1(plaintext1[1]), .A2(key_round[1]), .Y(n77) );
  AO222X1_HVT U317 ( .A1(out1[2]), .A2(n73), .A3(n74), .A4(n78), .A5(n76), 
        .A6(adk_out[2]), .Y(n335) );
  XOR2X1_HVT U318 ( .A1(plaintext1[2]), .A2(key_round[2]), .Y(n78) );
  AO222X1_HVT U319 ( .A1(out1[3]), .A2(n73), .A3(n74), .A4(n79), .A5(n76), 
        .A6(adk_out[3]), .Y(n334) );
  XOR2X1_HVT U320 ( .A1(plaintext1[3]), .A2(key_round[3]), .Y(n79) );
  AO222X1_HVT U321 ( .A1(out1[4]), .A2(n73), .A3(n74), .A4(n80), .A5(n76), 
        .A6(adk_out[4]), .Y(n333) );
  XOR2X1_HVT U322 ( .A1(plaintext1[4]), .A2(key_round[4]), .Y(n80) );
  AO222X1_HVT U323 ( .A1(out1[5]), .A2(n73), .A3(n74), .A4(n81), .A5(n76), 
        .A6(adk_out[5]), .Y(n332) );
  XOR2X1_HVT U324 ( .A1(plaintext1[5]), .A2(key_round[5]), .Y(n81) );
  AO222X1_HVT U325 ( .A1(out1[6]), .A2(n73), .A3(n74), .A4(n82), .A5(n76), 
        .A6(adk_out[6]), .Y(n331) );
  XOR2X1_HVT U326 ( .A1(plaintext1[6]), .A2(key_round[6]), .Y(n82) );
  AO222X1_HVT U327 ( .A1(out1[7]), .A2(n73), .A3(n74), .A4(n83), .A5(n76), 
        .A6(adk_out[7]), .Y(n330) );
  XOR2X1_HVT U328 ( .A1(plaintext1[7]), .A2(key_round[7]), .Y(n83) );
  AO222X1_HVT U329 ( .A1(out1[8]), .A2(n73), .A3(n74), .A4(n84), .A5(n76), 
        .A6(adk_out[8]), .Y(n329) );
  XOR2X1_HVT U330 ( .A1(plaintext1[8]), .A2(key_round[8]), .Y(n84) );
  AO222X1_HVT U331 ( .A1(out1[9]), .A2(n73), .A3(n74), .A4(n85), .A5(n76), 
        .A6(adk_out[9]), .Y(n328) );
  XOR2X1_HVT U332 ( .A1(plaintext1[9]), .A2(key_round[9]), .Y(n85) );
  AO222X1_HVT U333 ( .A1(out1[10]), .A2(n73), .A3(n74), .A4(n86), .A5(n76), 
        .A6(adk_out[10]), .Y(n327) );
  XOR2X1_HVT U334 ( .A1(plaintext1[10]), .A2(key_round[10]), .Y(n86) );
  AO222X1_HVT U335 ( .A1(out1[11]), .A2(n73), .A3(n74), .A4(n87), .A5(n76), 
        .A6(adk_out[11]), .Y(n326) );
  XOR2X1_HVT U336 ( .A1(plaintext1[11]), .A2(key_round[11]), .Y(n87) );
  AO222X1_HVT U337 ( .A1(out1[12]), .A2(n73), .A3(n74), .A4(n88), .A5(n76), 
        .A6(adk_out[12]), .Y(n325) );
  XOR2X1_HVT U338 ( .A1(plaintext1[12]), .A2(key_round[12]), .Y(n88) );
  AO222X1_HVT U339 ( .A1(out1[13]), .A2(n73), .A3(n74), .A4(n89), .A5(n76), 
        .A6(adk_out[13]), .Y(n324) );
  XOR2X1_HVT U340 ( .A1(plaintext1[13]), .A2(key_round[13]), .Y(n89) );
  AO222X1_HVT U341 ( .A1(out1[14]), .A2(n73), .A3(n74), .A4(n90), .A5(n76), 
        .A6(adk_out[14]), .Y(n323) );
  XOR2X1_HVT U342 ( .A1(plaintext1[14]), .A2(key_round[14]), .Y(n90) );
  AO222X1_HVT U343 ( .A1(out1[15]), .A2(n73), .A3(n74), .A4(n91), .A5(n76), 
        .A6(adk_out[15]), .Y(n322) );
  XOR2X1_HVT U344 ( .A1(plaintext1[15]), .A2(key_round[15]), .Y(n91) );
  AO222X1_HVT U345 ( .A1(out1[16]), .A2(n73), .A3(n74), .A4(n92), .A5(n76), 
        .A6(adk_out[16]), .Y(n321) );
  XOR2X1_HVT U346 ( .A1(plaintext1[16]), .A2(key_round[16]), .Y(n92) );
  AO222X1_HVT U347 ( .A1(out1[17]), .A2(n73), .A3(n74), .A4(n93), .A5(n76), 
        .A6(adk_out[17]), .Y(n320) );
  XOR2X1_HVT U348 ( .A1(plaintext1[17]), .A2(key_round[17]), .Y(n93) );
  AO222X1_HVT U349 ( .A1(out1[18]), .A2(n73), .A3(n74), .A4(n94), .A5(n76), 
        .A6(adk_out[18]), .Y(n319) );
  XOR2X1_HVT U350 ( .A1(plaintext1[18]), .A2(key_round[18]), .Y(n94) );
  AO222X1_HVT U351 ( .A1(out1[19]), .A2(n73), .A3(n74), .A4(n95), .A5(n76), 
        .A6(adk_out[19]), .Y(n318) );
  XOR2X1_HVT U352 ( .A1(plaintext1[19]), .A2(key_round[19]), .Y(n95) );
  AO222X1_HVT U353 ( .A1(out1[20]), .A2(n73), .A3(n74), .A4(n96), .A5(n76), 
        .A6(adk_out[20]), .Y(n317) );
  XOR2X1_HVT U354 ( .A1(plaintext1[20]), .A2(key_round[20]), .Y(n96) );
  AO222X1_HVT U355 ( .A1(out1[21]), .A2(n73), .A3(n74), .A4(n97), .A5(n76), 
        .A6(adk_out[21]), .Y(n316) );
  XOR2X1_HVT U356 ( .A1(plaintext1[21]), .A2(key_round[21]), .Y(n97) );
  AO222X1_HVT U357 ( .A1(out1[22]), .A2(n73), .A3(n74), .A4(n98), .A5(n76), 
        .A6(adk_out[22]), .Y(n315) );
  XOR2X1_HVT U358 ( .A1(plaintext1[22]), .A2(key_round[22]), .Y(n98) );
  AO222X1_HVT U359 ( .A1(out1[23]), .A2(n73), .A3(n74), .A4(n99), .A5(n76), 
        .A6(adk_out[23]), .Y(n314) );
  XOR2X1_HVT U360 ( .A1(plaintext1[23]), .A2(key_round[23]), .Y(n99) );
  AO222X1_HVT U361 ( .A1(out1[24]), .A2(n73), .A3(n74), .A4(n100), .A5(n76), 
        .A6(adk_out[24]), .Y(n313) );
  XOR2X1_HVT U362 ( .A1(plaintext1[24]), .A2(key_round[24]), .Y(n100) );
  AO222X1_HVT U363 ( .A1(out1[25]), .A2(n73), .A3(n74), .A4(n101), .A5(n76), 
        .A6(adk_out[25]), .Y(n312) );
  XOR2X1_HVT U364 ( .A1(plaintext1[25]), .A2(key_round[25]), .Y(n101) );
  AO222X1_HVT U365 ( .A1(out1[26]), .A2(n73), .A3(n74), .A4(n102), .A5(n76), 
        .A6(adk_out[26]), .Y(n311) );
  XOR2X1_HVT U366 ( .A1(plaintext1[26]), .A2(key_round[26]), .Y(n102) );
  AO222X1_HVT U367 ( .A1(out1[27]), .A2(n73), .A3(n74), .A4(n103), .A5(n76), 
        .A6(adk_out[27]), .Y(n310) );
  XOR2X1_HVT U368 ( .A1(plaintext1[27]), .A2(key_round[27]), .Y(n103) );
  AO222X1_HVT U369 ( .A1(out1[28]), .A2(n73), .A3(n74), .A4(n104), .A5(n76), 
        .A6(adk_out[28]), .Y(n309) );
  XOR2X1_HVT U370 ( .A1(plaintext1[28]), .A2(key_round[28]), .Y(n104) );
  AO222X1_HVT U371 ( .A1(out1[29]), .A2(n73), .A3(n74), .A4(n105), .A5(n76), 
        .A6(adk_out[29]), .Y(n308) );
  XOR2X1_HVT U372 ( .A1(plaintext1[29]), .A2(key_round[29]), .Y(n105) );
  AO222X1_HVT U373 ( .A1(out1[30]), .A2(n73), .A3(n74), .A4(n106), .A5(n76), 
        .A6(adk_out[30]), .Y(n307) );
  XOR2X1_HVT U374 ( .A1(plaintext1[30]), .A2(key_round[30]), .Y(n106) );
  AO222X1_HVT U375 ( .A1(out1[31]), .A2(n73), .A3(n74), .A4(n107), .A5(n76), 
        .A6(adk_out[31]), .Y(n306) );
  XOR2X1_HVT U376 ( .A1(plaintext1[31]), .A2(key_round[31]), .Y(n107) );
  AO222X1_HVT U377 ( .A1(out1[32]), .A2(n73), .A3(n74), .A4(n108), .A5(n76), 
        .A6(adk_out[32]), .Y(n305) );
  XOR2X1_HVT U378 ( .A1(plaintext1[32]), .A2(key_round[32]), .Y(n108) );
  AO222X1_HVT U379 ( .A1(out1[33]), .A2(n73), .A3(n74), .A4(n109), .A5(n76), 
        .A6(adk_out[33]), .Y(n304) );
  XOR2X1_HVT U380 ( .A1(plaintext1[33]), .A2(key_round[33]), .Y(n109) );
  AO222X1_HVT U381 ( .A1(out1[34]), .A2(n73), .A3(n74), .A4(n110), .A5(n76), 
        .A6(adk_out[34]), .Y(n303) );
  XOR2X1_HVT U382 ( .A1(plaintext1[34]), .A2(key_round[34]), .Y(n110) );
  AO222X1_HVT U383 ( .A1(out1[35]), .A2(n73), .A3(n74), .A4(n111), .A5(n76), 
        .A6(adk_out[35]), .Y(n302) );
  XOR2X1_HVT U384 ( .A1(plaintext1[35]), .A2(key_round[35]), .Y(n111) );
  AO222X1_HVT U385 ( .A1(out1[36]), .A2(n73), .A3(n74), .A4(n112), .A5(n76), 
        .A6(adk_out[36]), .Y(n301) );
  XOR2X1_HVT U386 ( .A1(plaintext1[36]), .A2(key_round[36]), .Y(n112) );
  AO222X1_HVT U387 ( .A1(out1[37]), .A2(n73), .A3(n74), .A4(n113), .A5(n76), 
        .A6(adk_out[37]), .Y(n300) );
  XOR2X1_HVT U388 ( .A1(plaintext1[37]), .A2(key_round[37]), .Y(n113) );
  AO222X1_HVT U389 ( .A1(out1[38]), .A2(n73), .A3(n74), .A4(n114), .A5(n76), 
        .A6(adk_out[38]), .Y(n299) );
  XOR2X1_HVT U390 ( .A1(plaintext1[38]), .A2(key_round[38]), .Y(n114) );
  AO222X1_HVT U391 ( .A1(out1[39]), .A2(n73), .A3(n74), .A4(n115), .A5(n76), 
        .A6(adk_out[39]), .Y(n298) );
  XOR2X1_HVT U392 ( .A1(plaintext1[39]), .A2(key_round[39]), .Y(n115) );
  AO222X1_HVT U393 ( .A1(out1[40]), .A2(n73), .A3(n74), .A4(n116), .A5(n76), 
        .A6(adk_out[40]), .Y(n297) );
  XOR2X1_HVT U394 ( .A1(plaintext1[40]), .A2(key_round[40]), .Y(n116) );
  AO222X1_HVT U395 ( .A1(out1[41]), .A2(n73), .A3(n74), .A4(n117), .A5(n76), 
        .A6(adk_out[41]), .Y(n296) );
  XOR2X1_HVT U396 ( .A1(plaintext1[41]), .A2(key_round[41]), .Y(n117) );
  AO222X1_HVT U397 ( .A1(out1[42]), .A2(n73), .A3(n74), .A4(n118), .A5(n76), 
        .A6(adk_out[42]), .Y(n295) );
  XOR2X1_HVT U398 ( .A1(plaintext1[42]), .A2(key_round[42]), .Y(n118) );
  AO222X1_HVT U399 ( .A1(out1[43]), .A2(n73), .A3(n74), .A4(n119), .A5(n76), 
        .A6(adk_out[43]), .Y(n294) );
  XOR2X1_HVT U400 ( .A1(plaintext1[43]), .A2(key_round[43]), .Y(n119) );
  AO222X1_HVT U401 ( .A1(out1[44]), .A2(n73), .A3(n74), .A4(n120), .A5(n76), 
        .A6(adk_out[44]), .Y(n293) );
  XOR2X1_HVT U402 ( .A1(plaintext1[44]), .A2(key_round[44]), .Y(n120) );
  AO222X1_HVT U403 ( .A1(out1[45]), .A2(n73), .A3(n74), .A4(n121), .A5(n76), 
        .A6(adk_out[45]), .Y(n292) );
  XOR2X1_HVT U404 ( .A1(plaintext1[45]), .A2(key_round[45]), .Y(n121) );
  AO222X1_HVT U405 ( .A1(out1[46]), .A2(n73), .A3(n74), .A4(n122), .A5(n76), 
        .A6(adk_out[46]), .Y(n291) );
  XOR2X1_HVT U406 ( .A1(plaintext1[46]), .A2(key_round[46]), .Y(n122) );
  AO222X1_HVT U407 ( .A1(out1[47]), .A2(n73), .A3(n74), .A4(n123), .A5(n76), 
        .A6(adk_out[47]), .Y(n290) );
  XOR2X1_HVT U408 ( .A1(plaintext1[47]), .A2(key_round[47]), .Y(n123) );
  AO222X1_HVT U409 ( .A1(out1[48]), .A2(n73), .A3(n74), .A4(n124), .A5(n76), 
        .A6(adk_out[48]), .Y(n289) );
  XOR2X1_HVT U410 ( .A1(plaintext1[48]), .A2(key_round[48]), .Y(n124) );
  AO222X1_HVT U411 ( .A1(out1[49]), .A2(n73), .A3(n74), .A4(n125), .A5(n76), 
        .A6(adk_out[49]), .Y(n288) );
  XOR2X1_HVT U412 ( .A1(plaintext1[49]), .A2(key_round[49]), .Y(n125) );
  AO222X1_HVT U413 ( .A1(out1[50]), .A2(n73), .A3(n74), .A4(n126), .A5(n76), 
        .A6(adk_out[50]), .Y(n287) );
  XOR2X1_HVT U414 ( .A1(plaintext1[50]), .A2(key_round[50]), .Y(n126) );
  AO222X1_HVT U415 ( .A1(out1[51]), .A2(n73), .A3(n74), .A4(n127), .A5(n76), 
        .A6(adk_out[51]), .Y(n286) );
  XOR2X1_HVT U416 ( .A1(plaintext1[51]), .A2(key_round[51]), .Y(n127) );
  AO222X1_HVT U417 ( .A1(out1[52]), .A2(n73), .A3(n74), .A4(n128), .A5(n76), 
        .A6(adk_out[52]), .Y(n285) );
  XOR2X1_HVT U418 ( .A1(plaintext1[52]), .A2(key_round[52]), .Y(n128) );
  AO222X1_HVT U419 ( .A1(out1[53]), .A2(n73), .A3(n74), .A4(n129), .A5(n76), 
        .A6(adk_out[53]), .Y(n284) );
  XOR2X1_HVT U420 ( .A1(plaintext1[53]), .A2(key_round[53]), .Y(n129) );
  AO222X1_HVT U421 ( .A1(out1[54]), .A2(n73), .A3(n74), .A4(n130), .A5(n76), 
        .A6(adk_out[54]), .Y(n283) );
  XOR2X1_HVT U422 ( .A1(plaintext1[54]), .A2(key_round[54]), .Y(n130) );
  AO222X1_HVT U423 ( .A1(out1[55]), .A2(n73), .A3(n74), .A4(n131), .A5(n76), 
        .A6(adk_out[55]), .Y(n282) );
  XOR2X1_HVT U424 ( .A1(plaintext1[55]), .A2(key_round[55]), .Y(n131) );
  AO222X1_HVT U425 ( .A1(out1[56]), .A2(n73), .A3(n74), .A4(n132), .A5(n76), 
        .A6(adk_out[56]), .Y(n281) );
  XOR2X1_HVT U426 ( .A1(plaintext1[56]), .A2(key_round[56]), .Y(n132) );
  AO222X1_HVT U427 ( .A1(out1[57]), .A2(n73), .A3(n74), .A4(n133), .A5(n76), 
        .A6(adk_out[57]), .Y(n280) );
  XOR2X1_HVT U428 ( .A1(plaintext1[57]), .A2(key_round[57]), .Y(n133) );
  AO222X1_HVT U429 ( .A1(out1[58]), .A2(n73), .A3(n74), .A4(n134), .A5(n76), 
        .A6(adk_out[58]), .Y(n279) );
  XOR2X1_HVT U430 ( .A1(plaintext1[58]), .A2(key_round[58]), .Y(n134) );
  AO222X1_HVT U431 ( .A1(out1[59]), .A2(n73), .A3(n74), .A4(n135), .A5(n76), 
        .A6(adk_out[59]), .Y(n278) );
  XOR2X1_HVT U432 ( .A1(plaintext1[59]), .A2(key_round[59]), .Y(n135) );
  AO222X1_HVT U433 ( .A1(out1[60]), .A2(n73), .A3(n74), .A4(n136), .A5(n76), 
        .A6(adk_out[60]), .Y(n277) );
  XOR2X1_HVT U434 ( .A1(plaintext1[60]), .A2(key_round[60]), .Y(n136) );
  AO222X1_HVT U435 ( .A1(out1[61]), .A2(n73), .A3(n74), .A4(n137), .A5(n76), 
        .A6(adk_out[61]), .Y(n276) );
  XOR2X1_HVT U436 ( .A1(plaintext1[61]), .A2(key_round[61]), .Y(n137) );
  AO222X1_HVT U437 ( .A1(out1[62]), .A2(n73), .A3(n74), .A4(n138), .A5(n76), 
        .A6(adk_out[62]), .Y(n275) );
  XOR2X1_HVT U438 ( .A1(plaintext1[62]), .A2(key_round[62]), .Y(n138) );
  AO222X1_HVT U439 ( .A1(out1[63]), .A2(n73), .A3(n74), .A4(n139), .A5(n76), 
        .A6(adk_out[63]), .Y(n274) );
  XOR2X1_HVT U440 ( .A1(plaintext1[63]), .A2(key_round[63]), .Y(n139) );
  AO222X1_HVT U441 ( .A1(out1[64]), .A2(n73), .A3(n74), .A4(n140), .A5(n76), 
        .A6(adk_out[64]), .Y(n273) );
  XOR2X1_HVT U442 ( .A1(plaintext1[64]), .A2(key_round[64]), .Y(n140) );
  AO222X1_HVT U443 ( .A1(out1[65]), .A2(n73), .A3(n74), .A4(n141), .A5(n76), 
        .A6(adk_out[65]), .Y(n272) );
  XOR2X1_HVT U444 ( .A1(plaintext1[65]), .A2(key_round[65]), .Y(n141) );
  AO222X1_HVT U445 ( .A1(out1[66]), .A2(n73), .A3(n74), .A4(n142), .A5(n76), 
        .A6(adk_out[66]), .Y(n271) );
  XOR2X1_HVT U446 ( .A1(plaintext1[66]), .A2(key_round[66]), .Y(n142) );
  AO222X1_HVT U447 ( .A1(out1[67]), .A2(n73), .A3(n74), .A4(n143), .A5(n76), 
        .A6(adk_out[67]), .Y(n270) );
  XOR2X1_HVT U448 ( .A1(plaintext1[67]), .A2(key_round[67]), .Y(n143) );
  AO222X1_HVT U449 ( .A1(out1[68]), .A2(n73), .A3(n74), .A4(n144), .A5(n76), 
        .A6(adk_out[68]), .Y(n269) );
  XOR2X1_HVT U450 ( .A1(plaintext1[68]), .A2(key_round[68]), .Y(n144) );
  AO222X1_HVT U451 ( .A1(out1[69]), .A2(n73), .A3(n74), .A4(n145), .A5(n76), 
        .A6(adk_out[69]), .Y(n268) );
  XOR2X1_HVT U452 ( .A1(plaintext1[69]), .A2(key_round[69]), .Y(n145) );
  AO222X1_HVT U453 ( .A1(out1[70]), .A2(n73), .A3(n74), .A4(n146), .A5(n76), 
        .A6(adk_out[70]), .Y(n267) );
  XOR2X1_HVT U454 ( .A1(plaintext1[70]), .A2(key_round[70]), .Y(n146) );
  AO222X1_HVT U455 ( .A1(out1[71]), .A2(n73), .A3(n74), .A4(n147), .A5(n76), 
        .A6(adk_out[71]), .Y(n266) );
  XOR2X1_HVT U456 ( .A1(plaintext1[71]), .A2(key_round[71]), .Y(n147) );
  AO222X1_HVT U457 ( .A1(out1[72]), .A2(n73), .A3(n74), .A4(n148), .A5(n76), 
        .A6(adk_out[72]), .Y(n265) );
  XOR2X1_HVT U458 ( .A1(plaintext1[72]), .A2(key_round[72]), .Y(n148) );
  AO222X1_HVT U459 ( .A1(out1[73]), .A2(n73), .A3(n74), .A4(n149), .A5(n76), 
        .A6(adk_out[73]), .Y(n264) );
  XOR2X1_HVT U460 ( .A1(plaintext1[73]), .A2(key_round[73]), .Y(n149) );
  AO222X1_HVT U461 ( .A1(out1[74]), .A2(n73), .A3(n74), .A4(n150), .A5(n76), 
        .A6(adk_out[74]), .Y(n263) );
  XOR2X1_HVT U462 ( .A1(plaintext1[74]), .A2(key_round[74]), .Y(n150) );
  AO222X1_HVT U463 ( .A1(out1[75]), .A2(n73), .A3(n74), .A4(n151), .A5(n76), 
        .A6(adk_out[75]), .Y(n262) );
  XOR2X1_HVT U464 ( .A1(plaintext1[75]), .A2(key_round[75]), .Y(n151) );
  AO222X1_HVT U465 ( .A1(out1[76]), .A2(n73), .A3(n74), .A4(n152), .A5(n76), 
        .A6(adk_out[76]), .Y(n261) );
  XOR2X1_HVT U466 ( .A1(plaintext1[76]), .A2(key_round[76]), .Y(n152) );
  AO222X1_HVT U467 ( .A1(out1[77]), .A2(n73), .A3(n74), .A4(n153), .A5(n76), 
        .A6(adk_out[77]), .Y(n260) );
  XOR2X1_HVT U468 ( .A1(plaintext1[77]), .A2(key_round[77]), .Y(n153) );
  AO222X1_HVT U469 ( .A1(out1[78]), .A2(n73), .A3(n74), .A4(n154), .A5(n76), 
        .A6(adk_out[78]), .Y(n259) );
  XOR2X1_HVT U470 ( .A1(plaintext1[78]), .A2(key_round[78]), .Y(n154) );
  AO222X1_HVT U471 ( .A1(out1[79]), .A2(n73), .A3(n74), .A4(n155), .A5(n76), 
        .A6(adk_out[79]), .Y(n258) );
  XOR2X1_HVT U472 ( .A1(plaintext1[79]), .A2(key_round[79]), .Y(n155) );
  AO222X1_HVT U473 ( .A1(out1[80]), .A2(n73), .A3(n74), .A4(n156), .A5(n76), 
        .A6(adk_out[80]), .Y(n257) );
  XOR2X1_HVT U474 ( .A1(plaintext1[80]), .A2(key_round[80]), .Y(n156) );
  AO222X1_HVT U475 ( .A1(out1[81]), .A2(n73), .A3(n74), .A4(n157), .A5(n76), 
        .A6(adk_out[81]), .Y(n256) );
  XOR2X1_HVT U476 ( .A1(plaintext1[81]), .A2(key_round[81]), .Y(n157) );
  AO222X1_HVT U477 ( .A1(out1[82]), .A2(n73), .A3(n74), .A4(n158), .A5(n76), 
        .A6(adk_out[82]), .Y(n255) );
  XOR2X1_HVT U478 ( .A1(plaintext1[82]), .A2(key_round[82]), .Y(n158) );
  AO222X1_HVT U479 ( .A1(out1[83]), .A2(n73), .A3(n74), .A4(n159), .A5(n76), 
        .A6(adk_out[83]), .Y(n254) );
  XOR2X1_HVT U480 ( .A1(plaintext1[83]), .A2(key_round[83]), .Y(n159) );
  AO222X1_HVT U481 ( .A1(out1[84]), .A2(n73), .A3(n74), .A4(n160), .A5(n76), 
        .A6(adk_out[84]), .Y(n253) );
  XOR2X1_HVT U482 ( .A1(plaintext1[84]), .A2(key_round[84]), .Y(n160) );
  AO222X1_HVT U483 ( .A1(out1[85]), .A2(n73), .A3(n74), .A4(n161), .A5(n76), 
        .A6(adk_out[85]), .Y(n252) );
  XOR2X1_HVT U484 ( .A1(plaintext1[85]), .A2(key_round[85]), .Y(n161) );
  AO222X1_HVT U485 ( .A1(out1[86]), .A2(n73), .A3(n74), .A4(n162), .A5(n76), 
        .A6(adk_out[86]), .Y(n251) );
  XOR2X1_HVT U486 ( .A1(plaintext1[86]), .A2(key_round[86]), .Y(n162) );
  AO222X1_HVT U487 ( .A1(out1[87]), .A2(n73), .A3(n74), .A4(n163), .A5(n76), 
        .A6(adk_out[87]), .Y(n250) );
  XOR2X1_HVT U488 ( .A1(plaintext1[87]), .A2(key_round[87]), .Y(n163) );
  AO222X1_HVT U489 ( .A1(out1[88]), .A2(n73), .A3(n74), .A4(n164), .A5(n76), 
        .A6(adk_out[88]), .Y(n249) );
  XOR2X1_HVT U490 ( .A1(plaintext1[88]), .A2(key_round[88]), .Y(n164) );
  AO222X1_HVT U491 ( .A1(out1[89]), .A2(n73), .A3(n74), .A4(n165), .A5(n76), 
        .A6(adk_out[89]), .Y(n248) );
  XOR2X1_HVT U492 ( .A1(plaintext1[89]), .A2(key_round[89]), .Y(n165) );
  AO222X1_HVT U493 ( .A1(out1[90]), .A2(n73), .A3(n74), .A4(n166), .A5(n76), 
        .A6(adk_out[90]), .Y(n247) );
  XOR2X1_HVT U494 ( .A1(plaintext1[90]), .A2(key_round[90]), .Y(n166) );
  AO222X1_HVT U495 ( .A1(out1[91]), .A2(n73), .A3(n74), .A4(n167), .A5(n76), 
        .A6(adk_out[91]), .Y(n246) );
  XOR2X1_HVT U496 ( .A1(plaintext1[91]), .A2(key_round[91]), .Y(n167) );
  AO222X1_HVT U497 ( .A1(out1[92]), .A2(n73), .A3(n74), .A4(n168), .A5(n76), 
        .A6(adk_out[92]), .Y(n245) );
  XOR2X1_HVT U498 ( .A1(plaintext1[92]), .A2(key_round[92]), .Y(n168) );
  AO222X1_HVT U499 ( .A1(out1[93]), .A2(n73), .A3(n74), .A4(n169), .A5(n76), 
        .A6(adk_out[93]), .Y(n244) );
  XOR2X1_HVT U500 ( .A1(plaintext1[93]), .A2(key_round[93]), .Y(n169) );
  AO222X1_HVT U501 ( .A1(out1[94]), .A2(n73), .A3(n74), .A4(n170), .A5(n76), 
        .A6(adk_out[94]), .Y(n243) );
  XOR2X1_HVT U502 ( .A1(plaintext1[94]), .A2(key_round[94]), .Y(n170) );
  AO222X1_HVT U503 ( .A1(out1[95]), .A2(n73), .A3(n74), .A4(n171), .A5(n76), 
        .A6(adk_out[95]), .Y(n242) );
  XOR2X1_HVT U504 ( .A1(plaintext1[95]), .A2(key_round[95]), .Y(n171) );
  AO222X1_HVT U505 ( .A1(out1[96]), .A2(n73), .A3(n74), .A4(n172), .A5(n76), 
        .A6(adk_out[96]), .Y(n241) );
  XOR2X1_HVT U506 ( .A1(plaintext1[96]), .A2(key_round[96]), .Y(n172) );
  AO222X1_HVT U507 ( .A1(out1[97]), .A2(n73), .A3(n74), .A4(n173), .A5(n76), 
        .A6(adk_out[97]), .Y(n240) );
  XOR2X1_HVT U508 ( .A1(plaintext1[97]), .A2(key_round[97]), .Y(n173) );
  AO222X1_HVT U509 ( .A1(out1[98]), .A2(n73), .A3(n74), .A4(n174), .A5(n76), 
        .A6(adk_out[98]), .Y(n239) );
  XOR2X1_HVT U510 ( .A1(plaintext1[98]), .A2(key_round[98]), .Y(n174) );
  AO222X1_HVT U511 ( .A1(out1[99]), .A2(n73), .A3(n74), .A4(n175), .A5(n76), 
        .A6(adk_out[99]), .Y(n238) );
  XOR2X1_HVT U512 ( .A1(plaintext1[99]), .A2(key_round[99]), .Y(n175) );
  AO222X1_HVT U513 ( .A1(out1[100]), .A2(n73), .A3(n74), .A4(n176), .A5(n76), 
        .A6(adk_out[100]), .Y(n237) );
  XOR2X1_HVT U514 ( .A1(plaintext1[100]), .A2(key_round[100]), .Y(n176) );
  AO222X1_HVT U515 ( .A1(out1[101]), .A2(n73), .A3(n74), .A4(n177), .A5(n76), 
        .A6(adk_out[101]), .Y(n236) );
  XOR2X1_HVT U516 ( .A1(plaintext1[101]), .A2(key_round[101]), .Y(n177) );
  AO222X1_HVT U517 ( .A1(out1[102]), .A2(n73), .A3(n74), .A4(n178), .A5(n76), 
        .A6(adk_out[102]), .Y(n235) );
  XOR2X1_HVT U518 ( .A1(plaintext1[102]), .A2(key_round[102]), .Y(n178) );
  AO222X1_HVT U519 ( .A1(out1[103]), .A2(n73), .A3(n74), .A4(n179), .A5(n76), 
        .A6(adk_out[103]), .Y(n234) );
  XOR2X1_HVT U520 ( .A1(plaintext1[103]), .A2(key_round[103]), .Y(n179) );
  AO222X1_HVT U521 ( .A1(out1[104]), .A2(n73), .A3(n74), .A4(n180), .A5(n76), 
        .A6(adk_out[104]), .Y(n233) );
  XOR2X1_HVT U522 ( .A1(plaintext1[104]), .A2(key_round[104]), .Y(n180) );
  AO222X1_HVT U523 ( .A1(out1[105]), .A2(n73), .A3(n74), .A4(n181), .A5(n76), 
        .A6(adk_out[105]), .Y(n232) );
  XOR2X1_HVT U524 ( .A1(plaintext1[105]), .A2(key_round[105]), .Y(n181) );
  AO222X1_HVT U525 ( .A1(out1[106]), .A2(n73), .A3(n74), .A4(n182), .A5(n76), 
        .A6(adk_out[106]), .Y(n231) );
  XOR2X1_HVT U526 ( .A1(plaintext1[106]), .A2(key_round[106]), .Y(n182) );
  AO222X1_HVT U527 ( .A1(out1[107]), .A2(n73), .A3(n74), .A4(n183), .A5(n76), 
        .A6(adk_out[107]), .Y(n230) );
  XOR2X1_HVT U528 ( .A1(plaintext1[107]), .A2(key_round[107]), .Y(n183) );
  AO222X1_HVT U529 ( .A1(out1[108]), .A2(n73), .A3(n74), .A4(n184), .A5(n76), 
        .A6(adk_out[108]), .Y(n229) );
  XOR2X1_HVT U530 ( .A1(plaintext1[108]), .A2(key_round[108]), .Y(n184) );
  AO222X1_HVT U531 ( .A1(out1[109]), .A2(n73), .A3(n74), .A4(n185), .A5(n76), 
        .A6(adk_out[109]), .Y(n228) );
  XOR2X1_HVT U532 ( .A1(plaintext1[109]), .A2(key_round[109]), .Y(n185) );
  AO222X1_HVT U533 ( .A1(out1[110]), .A2(n73), .A3(n74), .A4(n186), .A5(n76), 
        .A6(adk_out[110]), .Y(n227) );
  XOR2X1_HVT U534 ( .A1(plaintext1[110]), .A2(key_round[110]), .Y(n186) );
  AO222X1_HVT U535 ( .A1(out1[111]), .A2(n73), .A3(n74), .A4(n187), .A5(n76), 
        .A6(adk_out[111]), .Y(n226) );
  XOR2X1_HVT U536 ( .A1(plaintext1[111]), .A2(key_round[111]), .Y(n187) );
  AO222X1_HVT U537 ( .A1(out1[112]), .A2(n73), .A3(n74), .A4(n188), .A5(n76), 
        .A6(adk_out[112]), .Y(n225) );
  XOR2X1_HVT U538 ( .A1(plaintext1[112]), .A2(key_round[112]), .Y(n188) );
  AO222X1_HVT U539 ( .A1(out1[113]), .A2(n73), .A3(n74), .A4(n189), .A5(n76), 
        .A6(adk_out[113]), .Y(n224) );
  XOR2X1_HVT U540 ( .A1(plaintext1[113]), .A2(key_round[113]), .Y(n189) );
  AO222X1_HVT U541 ( .A1(out1[114]), .A2(n73), .A3(n74), .A4(n190), .A5(n76), 
        .A6(adk_out[114]), .Y(n223) );
  XOR2X1_HVT U542 ( .A1(plaintext1[114]), .A2(key_round[114]), .Y(n190) );
  AO222X1_HVT U543 ( .A1(out1[115]), .A2(n73), .A3(n74), .A4(n191), .A5(n76), 
        .A6(adk_out[115]), .Y(n222) );
  XOR2X1_HVT U544 ( .A1(plaintext1[115]), .A2(key_round[115]), .Y(n191) );
  AO222X1_HVT U545 ( .A1(out1[116]), .A2(n73), .A3(n74), .A4(n192), .A5(n76), 
        .A6(adk_out[116]), .Y(n221) );
  XOR2X1_HVT U546 ( .A1(plaintext1[116]), .A2(key_round[116]), .Y(n192) );
  AO222X1_HVT U547 ( .A1(out1[117]), .A2(n73), .A3(n74), .A4(n193), .A5(n76), 
        .A6(adk_out[117]), .Y(n220) );
  XOR2X1_HVT U548 ( .A1(plaintext1[117]), .A2(key_round[117]), .Y(n193) );
  AO222X1_HVT U549 ( .A1(out1[118]), .A2(n73), .A3(n74), .A4(n194), .A5(n76), 
        .A6(adk_out[118]), .Y(n219) );
  XOR2X1_HVT U550 ( .A1(plaintext1[118]), .A2(key_round[118]), .Y(n194) );
  AO222X1_HVT U551 ( .A1(out1[119]), .A2(n73), .A3(n74), .A4(n195), .A5(n76), 
        .A6(adk_out[119]), .Y(n218) );
  XOR2X1_HVT U552 ( .A1(plaintext1[119]), .A2(key_round[119]), .Y(n195) );
  AO222X1_HVT U553 ( .A1(out1[120]), .A2(n73), .A3(n74), .A4(n196), .A5(n76), 
        .A6(adk_out[120]), .Y(n217) );
  XOR2X1_HVT U554 ( .A1(plaintext1[120]), .A2(key_round[120]), .Y(n196) );
  AO222X1_HVT U555 ( .A1(out1[121]), .A2(n73), .A3(n74), .A4(n197), .A5(n76), 
        .A6(adk_out[121]), .Y(n216) );
  XOR2X1_HVT U556 ( .A1(plaintext1[121]), .A2(key_round[121]), .Y(n197) );
  AO222X1_HVT U557 ( .A1(out1[122]), .A2(n73), .A3(n74), .A4(n198), .A5(n76), 
        .A6(adk_out[122]), .Y(n215) );
  XOR2X1_HVT U558 ( .A1(plaintext1[122]), .A2(key_round[122]), .Y(n198) );
  AO222X1_HVT U559 ( .A1(out1[123]), .A2(n73), .A3(n74), .A4(n199), .A5(n76), 
        .A6(adk_out[123]), .Y(n214) );
  XOR2X1_HVT U560 ( .A1(plaintext1[123]), .A2(key_round[123]), .Y(n199) );
  AO222X1_HVT U561 ( .A1(out1[124]), .A2(n73), .A3(n74), .A4(n200), .A5(n76), 
        .A6(adk_out[124]), .Y(n213) );
  XOR2X1_HVT U562 ( .A1(plaintext1[124]), .A2(key_round[124]), .Y(n200) );
  AO222X1_HVT U563 ( .A1(out1[125]), .A2(n73), .A3(n74), .A4(n201), .A5(n76), 
        .A6(adk_out[125]), .Y(n212) );
  XOR2X1_HVT U564 ( .A1(plaintext1[125]), .A2(key_round[125]), .Y(n201) );
  AO222X1_HVT U565 ( .A1(out1[126]), .A2(n73), .A3(n74), .A4(n202), .A5(n76), 
        .A6(adk_out[126]), .Y(n211) );
  XOR2X1_HVT U566 ( .A1(plaintext1[126]), .A2(key_round[126]), .Y(n202) );
  AO222X1_HVT U567 ( .A1(out1[127]), .A2(n73), .A3(n74), .A4(n203), .A5(n76), 
        .A6(adk_out[127]), .Y(n210) );
  XOR2X1_HVT U568 ( .A1(plaintext1[127]), .A2(key_round[127]), .Y(n203) );
  AND2X1_HVT U569 ( .A1(n204), .A2(n64), .Y(n74) );
  INVX0_HVT U570 ( .A(n51), .Y(n64) );
  AND2X1_HVT U571 ( .A1(n204), .A2(n207), .Y(n73) );
  INVX0_HVT U572 ( .A(n76), .Y(n204) );
  NAND3X0_HVT U573 ( .A1(n209), .A2(n15), .A3(n22), .Y(n76) );
  INVX0_HVT U574 ( .A(n65), .Y(n22) );
  NAND2X0_HVT U575 ( .A1(n608), .A2(n16), .Y(n65) );
  INVX0_HVT U576 ( .A(rest), .Y(n609) );
  NAND2X0_HVT U577 ( .A1(n48), .A2(n51), .Y(n209) );
  NAND2X0_HVT U578 ( .A1(n23), .A2(n55), .Y(n51) );
  INVX0_HVT U579 ( .A(n207), .Y(n48) );
  NAND3X0_HVT U580 ( .A1(n53), .A2(n29), .A3(n605), .Y(n207) );
  AND3X1_HVT U581 ( .A1(n31), .A2(n43), .A3(n38), .Y(n605) );
  NAND2X0_HVT U582 ( .A1(n54), .A2(n606), .Y(n38) );
  NAND2X0_HVT U583 ( .A1(n71), .A2(n55), .Y(n43) );
  AND2X1_HVT U584 ( .A1(state[3]), .A2(n3), .Y(n55) );
  NAND2X0_HVT U585 ( .A1(n606), .A2(n68), .Y(n31) );
  OA21X1_HVT U586 ( .A1(n58), .A2(n607), .A3(n52), .Y(n29) );
  NAND2X0_HVT U587 ( .A1(n606), .A2(n23), .Y(n52) );
  INVX0_HVT U588 ( .A(n607), .Y(n23) );
  NAND2X0_HVT U589 ( .A1(state[2]), .A2(n4), .Y(n607) );
  AND4X1_HVT U590 ( .A1(n37), .A2(n63), .A3(n30), .A4(n62), .Y(n53) );
  NAND2X0_HVT U591 ( .A1(n40), .A2(n68), .Y(n62) );
  AND2X1_HVT U592 ( .A1(state[1]), .A2(n1), .Y(n68) );
  NAND2X0_HVT U593 ( .A1(n54), .A2(n40), .Y(n30) );
  INVX0_HVT U594 ( .A(n58), .Y(n40) );
  NAND2X0_HVT U595 ( .A1(n2), .A2(n3), .Y(n58) );
  AND2X1_HVT U596 ( .A1(state[2]), .A2(state[1]), .Y(n54) );
  NAND2X0_HVT U597 ( .A1(n71), .A2(n606), .Y(n63) );
  AND2X1_HVT U598 ( .A1(state[0]), .A2(n2), .Y(n606) );
  NAND2X0_HVT U599 ( .A1(n71), .A2(n21), .Y(n37) );
  AND2X1_HVT U600 ( .A1(state[0]), .A2(state[3]), .Y(n21) );
  AND2X1_HVT U601 ( .A1(n1), .A2(n4), .Y(n71) );
  OR2X1_HVT U602 ( .A1(n608), .A2(n25), .Y(n208) );
  INVX0_HVT U603 ( .A(n16), .Y(n25) );
  NAND3X0_HVT U604 ( .A1(n206), .A2(n205), .A3(start), .Y(n16) );
endmodule

