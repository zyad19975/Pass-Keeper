
module reg_D_4 ( clk, rst, enable, in, out );
  input [127:0] in;
  output [127:0] out;
  input clk, rst, enable;
  wire   n1, n129, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267;

  DFFARX1_HVT \out_reg[127]  ( .D(n140), .CLK(clk), .RSTB(n129), .Q(out[127])
         );
  DFFARX1_HVT \out_reg[126]  ( .D(n141), .CLK(clk), .RSTB(n129), .Q(out[126])
         );
  DFFARX1_HVT \out_reg[125]  ( .D(n142), .CLK(clk), .RSTB(n129), .Q(out[125])
         );
  DFFARX1_HVT \out_reg[124]  ( .D(n143), .CLK(clk), .RSTB(n129), .Q(out[124])
         );
  DFFARX1_HVT \out_reg[123]  ( .D(n144), .CLK(clk), .RSTB(n129), .Q(out[123])
         );
  DFFARX1_HVT \out_reg[122]  ( .D(n145), .CLK(clk), .RSTB(n1), .Q(out[122]) );
  DFFARX1_HVT \out_reg[121]  ( .D(n146), .CLK(clk), .RSTB(n129), .Q(out[121])
         );
  DFFARX1_HVT \out_reg[120]  ( .D(n147), .CLK(clk), .RSTB(n129), .Q(out[120])
         );
  DFFARX1_HVT \out_reg[119]  ( .D(n148), .CLK(clk), .RSTB(n138), .Q(out[119])
         );
  DFFARX1_HVT \out_reg[118]  ( .D(n149), .CLK(clk), .RSTB(n137), .Q(out[118])
         );
  DFFARX1_HVT \out_reg[117]  ( .D(n150), .CLK(clk), .RSTB(n137), .Q(out[117])
         );
  DFFARX1_HVT \out_reg[116]  ( .D(n151), .CLK(clk), .RSTB(n136), .Q(out[116])
         );
  DFFARX1_HVT \out_reg[115]  ( .D(n152), .CLK(clk), .RSTB(n132), .Q(out[115])
         );
  DFFARX1_HVT \out_reg[114]  ( .D(n153), .CLK(clk), .RSTB(n136), .Q(out[114])
         );
  DFFARX1_HVT \out_reg[113]  ( .D(n154), .CLK(clk), .RSTB(n136), .Q(out[113])
         );
  DFFARX1_HVT \out_reg[112]  ( .D(n155), .CLK(clk), .RSTB(n137), .Q(out[112])
         );
  DFFARX1_HVT \out_reg[111]  ( .D(n156), .CLK(clk), .RSTB(n135), .Q(out[111])
         );
  DFFARX1_HVT \out_reg[110]  ( .D(n157), .CLK(clk), .RSTB(n135), .Q(out[110])
         );
  DFFARX1_HVT \out_reg[109]  ( .D(n158), .CLK(clk), .RSTB(n135), .Q(out[109])
         );
  DFFARX1_HVT \out_reg[108]  ( .D(n159), .CLK(clk), .RSTB(n133), .Q(out[108])
         );
  DFFARX1_HVT \out_reg[107]  ( .D(n160), .CLK(clk), .RSTB(n129), .Q(out[107])
         );
  DFFARX1_HVT \out_reg[106]  ( .D(n161), .CLK(clk), .RSTB(n135), .Q(out[106])
         );
  DFFARX1_HVT \out_reg[105]  ( .D(n162), .CLK(clk), .RSTB(n135), .Q(out[105])
         );
  DFFARX1_HVT \out_reg[104]  ( .D(n163), .CLK(clk), .RSTB(n135), .Q(out[104])
         );
  DFFARX1_HVT \out_reg[103]  ( .D(n164), .CLK(clk), .RSTB(n139), .Q(out[103])
         );
  DFFARX1_HVT \out_reg[102]  ( .D(n165), .CLK(clk), .RSTB(n134), .Q(out[102])
         );
  DFFARX1_HVT \out_reg[101]  ( .D(n166), .CLK(clk), .RSTB(n134), .Q(out[101])
         );
  DFFARX1_HVT \out_reg[100]  ( .D(n167), .CLK(clk), .RSTB(n133), .Q(out[100])
         );
  DFFARX1_HVT \out_reg[99]  ( .D(n168), .CLK(clk), .RSTB(n133), .Q(out[99]) );
  DFFARX1_HVT \out_reg[98]  ( .D(n169), .CLK(clk), .RSTB(n134), .Q(out[98]) );
  DFFARX1_HVT \out_reg[97]  ( .D(n170), .CLK(clk), .RSTB(n138), .Q(out[97]) );
  DFFARX1_HVT \out_reg[96]  ( .D(n171), .CLK(clk), .RSTB(n138), .Q(out[96]) );
  DFFARX1_HVT \out_reg[95]  ( .D(n172), .CLK(clk), .RSTB(n131), .Q(out[95]) );
  DFFARX1_HVT \out_reg[94]  ( .D(n173), .CLK(clk), .RSTB(n131), .Q(out[94]) );
  DFFARX1_HVT \out_reg[93]  ( .D(n174), .CLK(clk), .RSTB(n131), .Q(out[93]) );
  DFFARX1_HVT \out_reg[92]  ( .D(n175), .CLK(clk), .RSTB(n129), .Q(out[92]) );
  DFFARX1_HVT \out_reg[91]  ( .D(n176), .CLK(clk), .RSTB(n129), .Q(out[91]) );
  DFFARX1_HVT \out_reg[90]  ( .D(n177), .CLK(clk), .RSTB(n131), .Q(out[90]) );
  DFFARX1_HVT \out_reg[89]  ( .D(n178), .CLK(clk), .RSTB(n129), .Q(out[89]) );
  DFFARX1_HVT \out_reg[88]  ( .D(n179), .CLK(clk), .RSTB(n131), .Q(out[88]) );
  DFFARX1_HVT \out_reg[87]  ( .D(n180), .CLK(clk), .RSTB(n138), .Q(out[87]) );
  DFFARX1_HVT \out_reg[86]  ( .D(n181), .CLK(clk), .RSTB(n137), .Q(out[86]) );
  DFFARX1_HVT \out_reg[85]  ( .D(n182), .CLK(clk), .RSTB(n136), .Q(out[85]) );
  DFFARX1_HVT \out_reg[84]  ( .D(n183), .CLK(clk), .RSTB(n136), .Q(out[84]) );
  DFFARX1_HVT \out_reg[83]  ( .D(n184), .CLK(clk), .RSTB(n132), .Q(out[83]) );
  DFFARX1_HVT \out_reg[82]  ( .D(n185), .CLK(clk), .RSTB(n137), .Q(out[82]) );
  DFFARX1_HVT \out_reg[81]  ( .D(n186), .CLK(clk), .RSTB(n136), .Q(out[81]) );
  DFFARX1_HVT \out_reg[80]  ( .D(n187), .CLK(clk), .RSTB(n137), .Q(out[80]) );
  DFFARX1_HVT \out_reg[79]  ( .D(n188), .CLK(clk), .RSTB(n132), .Q(out[79]) );
  DFFARX1_HVT \out_reg[78]  ( .D(n189), .CLK(clk), .RSTB(n131), .Q(out[78]) );
  DFFARX1_HVT \out_reg[77]  ( .D(n190), .CLK(clk), .RSTB(n132), .Q(out[77]) );
  DFFARX1_HVT \out_reg[76]  ( .D(n191), .CLK(clk), .RSTB(n131), .Q(out[76]) );
  DFFARX1_HVT \out_reg[75]  ( .D(n192), .CLK(clk), .RSTB(n131), .Q(out[75]) );
  DFFARX1_HVT \out_reg[74]  ( .D(n193), .CLK(clk), .RSTB(n1), .Q(out[74]) );
  DFFARX1_HVT \out_reg[73]  ( .D(n194), .CLK(clk), .RSTB(n132), .Q(out[73]) );
  DFFARX1_HVT \out_reg[72]  ( .D(n195), .CLK(clk), .RSTB(n132), .Q(out[72]) );
  DFFARX1_HVT \out_reg[71]  ( .D(n196), .CLK(clk), .RSTB(n138), .Q(out[71]) );
  DFFARX1_HVT \out_reg[70]  ( .D(n197), .CLK(clk), .RSTB(n135), .Q(out[70]) );
  DFFARX1_HVT \out_reg[69]  ( .D(n198), .CLK(clk), .RSTB(n134), .Q(out[69]) );
  DFFARX1_HVT \out_reg[68]  ( .D(n199), .CLK(clk), .RSTB(n138), .Q(out[68]) );
  DFFARX1_HVT \out_reg[67]  ( .D(n200), .CLK(clk), .RSTB(n134), .Q(out[67]) );
  DFFARX1_HVT \out_reg[66]  ( .D(n201), .CLK(clk), .RSTB(n133), .Q(out[66]) );
  DFFARX1_HVT \out_reg[65]  ( .D(n202), .CLK(clk), .RSTB(n134), .Q(out[65]) );
  DFFARX1_HVT \out_reg[64]  ( .D(n203), .CLK(clk), .RSTB(n138), .Q(out[64]) );
  DFFARX1_HVT \out_reg[63]  ( .D(n204), .CLK(clk), .RSTB(n133), .Q(out[63]) );
  DFFARX1_HVT \out_reg[62]  ( .D(n205), .CLK(clk), .RSTB(n133), .Q(out[62]) );
  DFFARX1_HVT \out_reg[61]  ( .D(n206), .CLK(clk), .RSTB(n133), .Q(out[61]) );
  DFFARX1_HVT \out_reg[60]  ( .D(n207), .CLK(clk), .RSTB(n133), .Q(out[60]) );
  DFFARX1_HVT \out_reg[59]  ( .D(n208), .CLK(clk), .RSTB(n133), .Q(out[59]) );
  DFFARX1_HVT \out_reg[58]  ( .D(n209), .CLK(clk), .RSTB(n132), .Q(out[58]) );
  DFFARX1_HVT \out_reg[57]  ( .D(n210), .CLK(clk), .RSTB(n133), .Q(out[57]) );
  DFFARX1_HVT \out_reg[56]  ( .D(n211), .CLK(clk), .RSTB(n133), .Q(out[56]) );
  DFFARX1_HVT \out_reg[55]  ( .D(n212), .CLK(clk), .RSTB(n138), .Q(out[55]) );
  DFFARX1_HVT \out_reg[54]  ( .D(n213), .CLK(clk), .RSTB(n136), .Q(out[54]) );
  DFFARX1_HVT \out_reg[53]  ( .D(n214), .CLK(clk), .RSTB(n136), .Q(out[53]) );
  DFFARX1_HVT \out_reg[52]  ( .D(n215), .CLK(clk), .RSTB(n137), .Q(out[52]) );
  DFFARX1_HVT \out_reg[51]  ( .D(n216), .CLK(clk), .RSTB(n132), .Q(out[51]) );
  DFFARX1_HVT \out_reg[50]  ( .D(n217), .CLK(clk), .RSTB(n1), .Q(out[50]) );
  DFFARX1_HVT \out_reg[49]  ( .D(n218), .CLK(clk), .RSTB(n137), .Q(out[49]) );
  DFFARX1_HVT \out_reg[48]  ( .D(n219), .CLK(clk), .RSTB(n137), .Q(out[48]) );
  DFFARX1_HVT \out_reg[47]  ( .D(n220), .CLK(clk), .RSTB(n135), .Q(out[47]) );
  DFFARX1_HVT \out_reg[46]  ( .D(n221), .CLK(clk), .RSTB(n135), .Q(out[46]) );
  DFFARX1_HVT \out_reg[45]  ( .D(n222), .CLK(clk), .RSTB(n135), .Q(out[45]) );
  DFFARX1_HVT \out_reg[44]  ( .D(n223), .CLK(clk), .RSTB(n135), .Q(out[44]) );
  DFFARX1_HVT \out_reg[43]  ( .D(n224), .CLK(clk), .RSTB(n133), .Q(out[43]) );
  DFFARX1_HVT \out_reg[42]  ( .D(n225), .CLK(clk), .RSTB(n136), .Q(out[42]) );
  DFFARX1_HVT \out_reg[41]  ( .D(n226), .CLK(clk), .RSTB(n129), .Q(out[41]) );
  DFFARX1_HVT \out_reg[40]  ( .D(n227), .CLK(clk), .RSTB(n135), .Q(out[40]) );
  DFFARX1_HVT \out_reg[39]  ( .D(n228), .CLK(clk), .RSTB(n138), .Q(out[39]) );
  DFFARX1_HVT \out_reg[38]  ( .D(n229), .CLK(clk), .RSTB(n131), .Q(out[38]) );
  DFFARX1_HVT \out_reg[37]  ( .D(n230), .CLK(clk), .RSTB(n134), .Q(out[37]) );
  DFFARX1_HVT \out_reg[36]  ( .D(n231), .CLK(clk), .RSTB(n134), .Q(out[36]) );
  DFFARX1_HVT \out_reg[35]  ( .D(n232), .CLK(clk), .RSTB(n134), .Q(out[35]) );
  DFFARX1_HVT \out_reg[34]  ( .D(n233), .CLK(clk), .RSTB(n135), .Q(out[34]) );
  DFFARX1_HVT \out_reg[33]  ( .D(n234), .CLK(clk), .RSTB(n132), .Q(out[33]) );
  DFFARX1_HVT \out_reg[32]  ( .D(n235), .CLK(clk), .RSTB(n138), .Q(out[32]) );
  DFFARX1_HVT \out_reg[31]  ( .D(n236), .CLK(clk), .RSTB(n1), .Q(out[31]) );
  DFFARX1_HVT \out_reg[30]  ( .D(n237), .CLK(clk), .RSTB(n1), .Q(out[30]) );
  DFFARX1_HVT \out_reg[29]  ( .D(n238), .CLK(clk), .RSTB(n1), .Q(out[29]) );
  DFFARX1_HVT \out_reg[28]  ( .D(n239), .CLK(clk), .RSTB(n1), .Q(out[28]) );
  DFFARX1_HVT \out_reg[27]  ( .D(n240), .CLK(clk), .RSTB(n1), .Q(out[27]) );
  DFFARX1_HVT \out_reg[26]  ( .D(n241), .CLK(clk), .RSTB(n1), .Q(out[26]) );
  DFFARX1_HVT \out_reg[25]  ( .D(n242), .CLK(clk), .RSTB(n1), .Q(out[25]) );
  DFFARX1_HVT \out_reg[24]  ( .D(n243), .CLK(clk), .RSTB(n1), .Q(out[24]) );
  DFFARX1_HVT \out_reg[23]  ( .D(n244), .CLK(clk), .RSTB(n138), .Q(out[23]) );
  DFFARX1_HVT \out_reg[22]  ( .D(n245), .CLK(clk), .RSTB(n137), .Q(out[22]) );
  DFFARX1_HVT \out_reg[21]  ( .D(n246), .CLK(clk), .RSTB(n136), .Q(out[21]) );
  DFFARX1_HVT \out_reg[20]  ( .D(n247), .CLK(clk), .RSTB(n136), .Q(out[20]) );
  DFFARX1_HVT \out_reg[19]  ( .D(n248), .CLK(clk), .RSTB(n1), .Q(out[19]) );
  DFFARX1_HVT \out_reg[18]  ( .D(n249), .CLK(clk), .RSTB(n136), .Q(out[18]) );
  DFFARX1_HVT \out_reg[17]  ( .D(n250), .CLK(clk), .RSTB(n137), .Q(out[17]) );
  DFFARX1_HVT \out_reg[16]  ( .D(n251), .CLK(clk), .RSTB(n137), .Q(out[16]) );
  DFFARX1_HVT \out_reg[15]  ( .D(n252), .CLK(clk), .RSTB(n132), .Q(out[15]) );
  DFFARX1_HVT \out_reg[14]  ( .D(n253), .CLK(clk), .RSTB(n132), .Q(out[14]) );
  DFFARX1_HVT \out_reg[13]  ( .D(n254), .CLK(clk), .RSTB(n131), .Q(out[13]) );
  DFFARX1_HVT \out_reg[12]  ( .D(n255), .CLK(clk), .RSTB(n131), .Q(out[12]) );
  DFFARX1_HVT \out_reg[11]  ( .D(n256), .CLK(clk), .RSTB(n132), .Q(out[11]) );
  DFFARX1_HVT \out_reg[10]  ( .D(n257), .CLK(clk), .RSTB(n131), .Q(out[10]) );
  DFFARX1_HVT \out_reg[9]  ( .D(n258), .CLK(clk), .RSTB(n131), .Q(out[9]) );
  DFFARX1_HVT \out_reg[8]  ( .D(n259), .CLK(clk), .RSTB(n132), .Q(out[8]) );
  DFFARX1_HVT \out_reg[7]  ( .D(n260), .CLK(clk), .RSTB(n139), .Q(out[7]) );
  DFFARX1_HVT \out_reg[6]  ( .D(n261), .CLK(clk), .RSTB(n138), .Q(out[6]) );
  DFFARX1_HVT \out_reg[5]  ( .D(n262), .CLK(clk), .RSTB(n134), .Q(out[5]) );
  DFFARX1_HVT \out_reg[4]  ( .D(n263), .CLK(clk), .RSTB(n134), .Q(out[4]) );
  DFFARX1_HVT \out_reg[3]  ( .D(n264), .CLK(clk), .RSTB(n133), .Q(out[3]) );
  DFFARX1_HVT \out_reg[2]  ( .D(n265), .CLK(clk), .RSTB(n134), .Q(out[2]) );
  DFFARX1_HVT \out_reg[1]  ( .D(n266), .CLK(clk), .RSTB(n134), .Q(out[1]) );
  DFFARX1_HVT \out_reg[0]  ( .D(n267), .CLK(clk), .RSTB(n138), .Q(out[0]) );
  NBUFFX2_HVT U2 ( .A(n139), .Y(n138) );
  NBUFFX2_HVT U3 ( .A(n139), .Y(n131) );
  NBUFFX2_HVT U4 ( .A(n139), .Y(n134) );
  NBUFFX2_HVT U5 ( .A(n139), .Y(n133) );
  NBUFFX2_HVT U6 ( .A(n139), .Y(n135) );
  NBUFFX2_HVT U7 ( .A(n139), .Y(n132) );
  NBUFFX2_HVT U8 ( .A(n139), .Y(n136) );
  NBUFFX2_HVT U9 ( .A(n139), .Y(n137) );
  NBUFFX2_HVT U10 ( .A(n139), .Y(n1) );
  NBUFFX2_HVT U11 ( .A(n139), .Y(n129) );
  INVX0_HVT U12 ( .A(rst), .Y(n139) );
  MUX21X1_HVT U13 ( .A1(out[97]), .A2(in[97]), .S0(enable), .Y(n170) );
  MUX21X1_HVT U14 ( .A1(out[96]), .A2(in[96]), .S0(enable), .Y(n171) );
  MUX21X1_HVT U15 ( .A1(out[95]), .A2(in[95]), .S0(enable), .Y(n172) );
  MUX21X1_HVT U16 ( .A1(out[94]), .A2(in[94]), .S0(enable), .Y(n173) );
  MUX21X1_HVT U17 ( .A1(out[93]), .A2(in[93]), .S0(enable), .Y(n174) );
  MUX21X1_HVT U18 ( .A1(out[92]), .A2(in[92]), .S0(enable), .Y(n175) );
  MUX21X1_HVT U19 ( .A1(out[91]), .A2(in[91]), .S0(enable), .Y(n176) );
  MUX21X1_HVT U20 ( .A1(out[90]), .A2(in[90]), .S0(enable), .Y(n177) );
  MUX21X1_HVT U21 ( .A1(out[89]), .A2(in[89]), .S0(enable), .Y(n178) );
  MUX21X1_HVT U22 ( .A1(out[88]), .A2(in[88]), .S0(enable), .Y(n179) );
  MUX21X1_HVT U23 ( .A1(out[7]), .A2(in[7]), .S0(enable), .Y(n260) );
  MUX21X1_HVT U24 ( .A1(out[87]), .A2(in[87]), .S0(enable), .Y(n180) );
  MUX21X1_HVT U25 ( .A1(out[86]), .A2(in[86]), .S0(enable), .Y(n181) );
  MUX21X1_HVT U26 ( .A1(out[85]), .A2(in[85]), .S0(enable), .Y(n182) );
  MUX21X1_HVT U27 ( .A1(out[84]), .A2(in[84]), .S0(enable), .Y(n183) );
  MUX21X1_HVT U28 ( .A1(out[83]), .A2(in[83]), .S0(enable), .Y(n184) );
  MUX21X1_HVT U29 ( .A1(out[82]), .A2(in[82]), .S0(enable), .Y(n185) );
  MUX21X1_HVT U30 ( .A1(out[81]), .A2(in[81]), .S0(enable), .Y(n186) );
  MUX21X1_HVT U31 ( .A1(out[80]), .A2(in[80]), .S0(enable), .Y(n187) );
  MUX21X1_HVT U32 ( .A1(out[79]), .A2(in[79]), .S0(enable), .Y(n188) );
  MUX21X1_HVT U33 ( .A1(out[78]), .A2(in[78]), .S0(enable), .Y(n189) );
  MUX21X1_HVT U34 ( .A1(out[6]), .A2(in[6]), .S0(enable), .Y(n261) );
  MUX21X1_HVT U35 ( .A1(out[77]), .A2(in[77]), .S0(enable), .Y(n190) );
  MUX21X1_HVT U36 ( .A1(out[76]), .A2(in[76]), .S0(enable), .Y(n191) );
  MUX21X1_HVT U37 ( .A1(out[75]), .A2(in[75]), .S0(enable), .Y(n192) );
  MUX21X1_HVT U38 ( .A1(out[74]), .A2(in[74]), .S0(enable), .Y(n193) );
  MUX21X1_HVT U39 ( .A1(out[73]), .A2(in[73]), .S0(enable), .Y(n194) );
  MUX21X1_HVT U40 ( .A1(out[72]), .A2(in[72]), .S0(enable), .Y(n195) );
  MUX21X1_HVT U41 ( .A1(out[71]), .A2(in[71]), .S0(enable), .Y(n196) );
  MUX21X1_HVT U42 ( .A1(out[70]), .A2(in[70]), .S0(enable), .Y(n197) );
  MUX21X1_HVT U43 ( .A1(out[69]), .A2(in[69]), .S0(enable), .Y(n198) );
  MUX21X1_HVT U44 ( .A1(out[68]), .A2(in[68]), .S0(enable), .Y(n199) );
  MUX21X1_HVT U45 ( .A1(out[5]), .A2(in[5]), .S0(enable), .Y(n262) );
  MUX21X1_HVT U46 ( .A1(out[67]), .A2(in[67]), .S0(enable), .Y(n200) );
  MUX21X1_HVT U47 ( .A1(out[66]), .A2(in[66]), .S0(enable), .Y(n201) );
  MUX21X1_HVT U48 ( .A1(out[65]), .A2(in[65]), .S0(enable), .Y(n202) );
  MUX21X1_HVT U49 ( .A1(out[64]), .A2(in[64]), .S0(enable), .Y(n203) );
  MUX21X1_HVT U50 ( .A1(out[63]), .A2(in[63]), .S0(enable), .Y(n204) );
  MUX21X1_HVT U51 ( .A1(out[62]), .A2(in[62]), .S0(enable), .Y(n205) );
  MUX21X1_HVT U52 ( .A1(out[61]), .A2(in[61]), .S0(enable), .Y(n206) );
  MUX21X1_HVT U53 ( .A1(out[60]), .A2(in[60]), .S0(enable), .Y(n207) );
  MUX21X1_HVT U54 ( .A1(out[59]), .A2(in[59]), .S0(enable), .Y(n208) );
  MUX21X1_HVT U55 ( .A1(out[58]), .A2(in[58]), .S0(enable), .Y(n209) );
  MUX21X1_HVT U56 ( .A1(out[4]), .A2(in[4]), .S0(enable), .Y(n263) );
  MUX21X1_HVT U57 ( .A1(out[57]), .A2(in[57]), .S0(enable), .Y(n210) );
  MUX21X1_HVT U58 ( .A1(out[56]), .A2(in[56]), .S0(enable), .Y(n211) );
  MUX21X1_HVT U59 ( .A1(out[55]), .A2(in[55]), .S0(enable), .Y(n212) );
  MUX21X1_HVT U60 ( .A1(out[54]), .A2(in[54]), .S0(enable), .Y(n213) );
  MUX21X1_HVT U61 ( .A1(out[53]), .A2(in[53]), .S0(enable), .Y(n214) );
  MUX21X1_HVT U62 ( .A1(out[52]), .A2(in[52]), .S0(enable), .Y(n215) );
  MUX21X1_HVT U63 ( .A1(out[51]), .A2(in[51]), .S0(enable), .Y(n216) );
  MUX21X1_HVT U64 ( .A1(out[50]), .A2(in[50]), .S0(enable), .Y(n217) );
  MUX21X1_HVT U65 ( .A1(out[49]), .A2(in[49]), .S0(enable), .Y(n218) );
  MUX21X1_HVT U66 ( .A1(out[48]), .A2(in[48]), .S0(enable), .Y(n219) );
  MUX21X1_HVT U67 ( .A1(out[3]), .A2(in[3]), .S0(enable), .Y(n264) );
  MUX21X1_HVT U68 ( .A1(out[47]), .A2(in[47]), .S0(enable), .Y(n220) );
  MUX21X1_HVT U69 ( .A1(out[46]), .A2(in[46]), .S0(enable), .Y(n221) );
  MUX21X1_HVT U70 ( .A1(out[45]), .A2(in[45]), .S0(enable), .Y(n222) );
  MUX21X1_HVT U71 ( .A1(out[44]), .A2(in[44]), .S0(enable), .Y(n223) );
  MUX21X1_HVT U72 ( .A1(out[43]), .A2(in[43]), .S0(enable), .Y(n224) );
  MUX21X1_HVT U73 ( .A1(out[42]), .A2(in[42]), .S0(enable), .Y(n225) );
  MUX21X1_HVT U74 ( .A1(out[41]), .A2(in[41]), .S0(enable), .Y(n226) );
  MUX21X1_HVT U75 ( .A1(out[40]), .A2(in[40]), .S0(enable), .Y(n227) );
  MUX21X1_HVT U76 ( .A1(out[39]), .A2(in[39]), .S0(enable), .Y(n228) );
  MUX21X1_HVT U77 ( .A1(out[38]), .A2(in[38]), .S0(enable), .Y(n229) );
  MUX21X1_HVT U78 ( .A1(out[2]), .A2(in[2]), .S0(enable), .Y(n265) );
  MUX21X1_HVT U79 ( .A1(out[37]), .A2(in[37]), .S0(enable), .Y(n230) );
  MUX21X1_HVT U80 ( .A1(out[36]), .A2(in[36]), .S0(enable), .Y(n231) );
  MUX21X1_HVT U81 ( .A1(out[35]), .A2(in[35]), .S0(enable), .Y(n232) );
  MUX21X1_HVT U82 ( .A1(out[34]), .A2(in[34]), .S0(enable), .Y(n233) );
  MUX21X1_HVT U83 ( .A1(out[33]), .A2(in[33]), .S0(enable), .Y(n234) );
  MUX21X1_HVT U84 ( .A1(out[32]), .A2(in[32]), .S0(enable), .Y(n235) );
  MUX21X1_HVT U85 ( .A1(out[31]), .A2(in[31]), .S0(enable), .Y(n236) );
  MUX21X1_HVT U86 ( .A1(out[30]), .A2(in[30]), .S0(enable), .Y(n237) );
  MUX21X1_HVT U87 ( .A1(out[29]), .A2(in[29]), .S0(enable), .Y(n238) );
  MUX21X1_HVT U88 ( .A1(out[28]), .A2(in[28]), .S0(enable), .Y(n239) );
  MUX21X1_HVT U89 ( .A1(out[1]), .A2(in[1]), .S0(enable), .Y(n266) );
  MUX21X1_HVT U90 ( .A1(out[27]), .A2(in[27]), .S0(enable), .Y(n240) );
  MUX21X1_HVT U91 ( .A1(out[26]), .A2(in[26]), .S0(enable), .Y(n241) );
  MUX21X1_HVT U92 ( .A1(out[25]), .A2(in[25]), .S0(enable), .Y(n242) );
  MUX21X1_HVT U93 ( .A1(out[24]), .A2(in[24]), .S0(enable), .Y(n243) );
  MUX21X1_HVT U94 ( .A1(out[23]), .A2(in[23]), .S0(enable), .Y(n244) );
  MUX21X1_HVT U95 ( .A1(out[22]), .A2(in[22]), .S0(enable), .Y(n245) );
  MUX21X1_HVT U96 ( .A1(out[21]), .A2(in[21]), .S0(enable), .Y(n246) );
  MUX21X1_HVT U97 ( .A1(out[20]), .A2(in[20]), .S0(enable), .Y(n247) );
  MUX21X1_HVT U98 ( .A1(out[19]), .A2(in[19]), .S0(enable), .Y(n248) );
  MUX21X1_HVT U99 ( .A1(out[18]), .A2(in[18]), .S0(enable), .Y(n249) );
  MUX21X1_HVT U100 ( .A1(out[0]), .A2(in[0]), .S0(enable), .Y(n267) );
  MUX21X1_HVT U101 ( .A1(out[17]), .A2(in[17]), .S0(enable), .Y(n250) );
  MUX21X1_HVT U102 ( .A1(out[16]), .A2(in[16]), .S0(enable), .Y(n251) );
  MUX21X1_HVT U103 ( .A1(out[15]), .A2(in[15]), .S0(enable), .Y(n252) );
  MUX21X1_HVT U104 ( .A1(out[14]), .A2(in[14]), .S0(enable), .Y(n253) );
  MUX21X1_HVT U105 ( .A1(out[13]), .A2(in[13]), .S0(enable), .Y(n254) );
  MUX21X1_HVT U106 ( .A1(out[12]), .A2(in[12]), .S0(enable), .Y(n255) );
  MUX21X1_HVT U107 ( .A1(out[127]), .A2(in[127]), .S0(enable), .Y(n140) );
  MUX21X1_HVT U108 ( .A1(out[11]), .A2(in[11]), .S0(enable), .Y(n256) );
  MUX21X1_HVT U109 ( .A1(out[126]), .A2(in[126]), .S0(enable), .Y(n141) );
  MUX21X1_HVT U110 ( .A1(out[125]), .A2(in[125]), .S0(enable), .Y(n142) );
  MUX21X1_HVT U111 ( .A1(out[124]), .A2(in[124]), .S0(enable), .Y(n143) );
  MUX21X1_HVT U112 ( .A1(out[123]), .A2(in[123]), .S0(enable), .Y(n144) );
  MUX21X1_HVT U113 ( .A1(out[122]), .A2(in[122]), .S0(enable), .Y(n145) );
  MUX21X1_HVT U114 ( .A1(out[121]), .A2(in[121]), .S0(enable), .Y(n146) );
  MUX21X1_HVT U115 ( .A1(out[120]), .A2(in[120]), .S0(enable), .Y(n147) );
  MUX21X1_HVT U116 ( .A1(out[119]), .A2(in[119]), .S0(enable), .Y(n148) );
  MUX21X1_HVT U117 ( .A1(out[118]), .A2(in[118]), .S0(enable), .Y(n149) );
  MUX21X1_HVT U118 ( .A1(out[10]), .A2(in[10]), .S0(enable), .Y(n257) );
  MUX21X1_HVT U119 ( .A1(out[117]), .A2(in[117]), .S0(enable), .Y(n150) );
  MUX21X1_HVT U120 ( .A1(out[116]), .A2(in[116]), .S0(enable), .Y(n151) );
  MUX21X1_HVT U121 ( .A1(out[115]), .A2(in[115]), .S0(enable), .Y(n152) );
  MUX21X1_HVT U122 ( .A1(out[114]), .A2(in[114]), .S0(enable), .Y(n153) );
  MUX21X1_HVT U123 ( .A1(out[113]), .A2(in[113]), .S0(enable), .Y(n154) );
  MUX21X1_HVT U124 ( .A1(out[112]), .A2(in[112]), .S0(enable), .Y(n155) );
  MUX21X1_HVT U125 ( .A1(out[111]), .A2(in[111]), .S0(enable), .Y(n156) );
  MUX21X1_HVT U126 ( .A1(out[110]), .A2(in[110]), .S0(enable), .Y(n157) );
  MUX21X1_HVT U127 ( .A1(out[109]), .A2(in[109]), .S0(enable), .Y(n158) );
  MUX21X1_HVT U128 ( .A1(out[108]), .A2(in[108]), .S0(enable), .Y(n159) );
  MUX21X1_HVT U129 ( .A1(out[9]), .A2(in[9]), .S0(enable), .Y(n258) );
  MUX21X1_HVT U130 ( .A1(out[107]), .A2(in[107]), .S0(enable), .Y(n160) );
  MUX21X1_HVT U131 ( .A1(out[106]), .A2(in[106]), .S0(enable), .Y(n161) );
  MUX21X1_HVT U132 ( .A1(out[105]), .A2(in[105]), .S0(enable), .Y(n162) );
  MUX21X1_HVT U133 ( .A1(out[104]), .A2(in[104]), .S0(enable), .Y(n163) );
  MUX21X1_HVT U134 ( .A1(out[103]), .A2(in[103]), .S0(enable), .Y(n164) );
  MUX21X1_HVT U135 ( .A1(out[102]), .A2(in[102]), .S0(enable), .Y(n165) );
  MUX21X1_HVT U136 ( .A1(out[101]), .A2(in[101]), .S0(enable), .Y(n166) );
  MUX21X1_HVT U137 ( .A1(out[100]), .A2(in[100]), .S0(enable), .Y(n167) );
  MUX21X1_HVT U138 ( .A1(out[99]), .A2(in[99]), .S0(enable), .Y(n168) );
  MUX21X1_HVT U139 ( .A1(out[98]), .A2(in[98]), .S0(enable), .Y(n169) );
  MUX21X1_HVT U140 ( .A1(out[8]), .A2(in[8]), .S0(enable), .Y(n259) );
endmodule

