
module sbox_11 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n7, n17, n19, n23, n50, n118, n119, n210, n211, n212, n213, n216,
         n217, n218, n219, n224, n227, n231, n232, n233, n236, n238, n242,
         n249, n256, n258, n261, n264, n268, n269, n272, n273, n274, n278,
         n279, n280, n282, n283, n285, n290, n293, n297, n301, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762;

  NAND2X0_HVT U4 ( .A1(n216), .A2(n210), .Y(n759) );
  NAND2X0_HVT U5 ( .A1(n431), .A2(n484), .Y(n757) );
  NAND2X0_HVT U13 ( .A1(n750), .A2(n351), .Y(n751) );
  NAND2X0_HVT U15 ( .A1(n211), .A2(n323), .Y(n748) );
  NAND2X0_HVT U21 ( .A1(n216), .A2(n494), .Y(n744) );
  NAND2X0_HVT U33 ( .A1(n525), .A2(n494), .Y(n733) );
  NAND2X0_HVT U42 ( .A1(n358), .A2(n428), .Y(n724) );
  NAND2X0_HVT U53 ( .A1(n713), .A2(n723), .Y(n714) );
  NAND2X0_HVT U56 ( .A1(n216), .A2(n709), .Y(n710) );
  MUX41X1_HVT U57 ( .A1(n519), .A3(n746), .A2(n710), .A4(n753), .S0(n501), 
        .S1(n472), .Y(n708) );
  NAND2X0_HVT U58 ( .A1(n350), .A2(n210), .Y(n707) );
  NAND2X0_HVT U62 ( .A1(n494), .A2(n213), .Y(n703) );
  MUX41X1_HVT U68 ( .A1(n516), .A3(n699), .A2(n698), .A4(n700), .S0(n468), 
        .S1(n498), .Y(n697) );
  NAND2X0_HVT U73 ( .A1(n487), .A2(n692), .Y(n693) );
  MUX41X1_HVT U75 ( .A1(n542), .A3(n539), .A2(n433), .A4(n505), .S0(n468), 
        .S1(n455), .Y(n690) );
  MUX41X1_HVT U77 ( .A1(n755), .A3(n526), .A2(n689), .A4(n427), .S0(n475), 
        .S1(n469), .Y(n688) );
  MUX41X1_HVT U78 ( .A1(n688), .A3(n691), .A2(n690), .A4(n695), .S0(n478), 
        .S1(n472), .Y(n687) );
  AND2X1_HVT U83 ( .A1(n431), .A2(n447), .Y(n681) );
  MUX41X1_HVT U84 ( .A1(n517), .A3(n422), .A2(n17), .A4(n681), .S0(n468), .S1(
        n454), .Y(n680) );
  NAND2X0_HVT U85 ( .A1(n494), .A2(n347), .Y(n679) );
  MUX41X1_HVT U86 ( .A1(n539), .A3(n679), .A2(n462), .A4(n459), .S0(n468), 
        .S1(n498), .Y(n678) );
  MUX41X1_HVT U90 ( .A1(n720), .A3(n724), .A2(n510), .A4(n676), .S0(n413), 
        .S1(n455), .Y(n675) );
  NAND2X0_HVT U101 ( .A1(n662), .A2(n661), .Y(n663) );
  MUX41X1_HVT U103 ( .A1(n210), .A3(n304), .A2(n394), .A4(n731), .S0(n468), 
        .S1(n455), .Y(n659) );
  MUX41X1_HVT U105 ( .A1(n537), .A3(n718), .A2(n658), .A4(n528), .S0(n468), 
        .S1(n454), .Y(n657) );
  NAND2X0_HVT U110 ( .A1(n322), .A2(n273), .Y(n653) );
  AND2X1_HVT U115 ( .A1(n379), .A2(n323), .Y(n649) );
  AND3X1_HVT U128 ( .A1(n470), .A2(n494), .A3(n447), .Y(n634) );
  MUX41X1_HVT U131 ( .A1(n632), .A3(n634), .A2(n633), .A4(n635), .S0(n474), 
        .S1(n501), .Y(n631) );
  MUX41X1_HVT U135 ( .A1(n19), .A3(n434), .A2(n757), .A4(n739), .S0(n443), 
        .S1(n499), .Y(n628) );
  AND2X1_HVT U140 ( .A1(n486), .A2(n494), .Y(n623) );
  MUX41X1_HVT U153 ( .A1(n653), .A3(n463), .A2(n213), .A4(n424), .S0(n495), 
        .S1(n454), .Y(n611) );
  AND2X1_HVT U154 ( .A1(n477), .A2(n428), .Y(n610) );
  NAND2X0_HVT U158 ( .A1(n491), .A2(n545), .Y(n606) );
  AND2X1_HVT U162 ( .A1(n422), .A2(n274), .Y(n602) );
  MUX41X1_HVT U165 ( .A1(n744), .A3(n536), .A2(n720), .A4(n600), .S0(n499), 
        .S1(n380), .Y(n599) );
  NAND2X0_HVT U166 ( .A1(n349), .A2(n709), .Y(n598) );
  NAND2X0_HVT U167 ( .A1(n508), .A2(n494), .Y(n597) );
  MUX41X1_HVT U168 ( .A1(n519), .A3(n487), .A2(n597), .A4(n598), .S0(n443), 
        .S1(n498), .Y(n596) );
  NAND2X0_HVT U174 ( .A1(n491), .A2(n310), .Y(n750) );
  MUX41X1_HVT U176 ( .A1(n482), .A3(n591), .A2(n518), .A4(n436), .S0(n501), 
        .S1(n238), .Y(n590) );
  NAND2X0_HVT U177 ( .A1(n491), .A2(n389), .Y(n589) );
  MUX41X1_HVT U178 ( .A1(n747), .A3(n589), .A2(n534), .A4(n728), .S0(n380), 
        .S1(n501), .Y(n588) );
  MUX41X1_HVT U179 ( .A1(n738), .A3(n533), .A2(n520), .A4(n534), .S0(n443), 
        .S1(n499), .Y(n587) );
  MUX41X1_HVT U180 ( .A1(n515), .A3(n755), .A2(n751), .A4(n7), .S0(n475), .S1(
        n443), .Y(n586) );
  MUX41X1_HVT U182 ( .A1(n340), .A3(n216), .A2(n511), .A4(n531), .S0(n499), 
        .S1(n471), .Y(n584) );
  MUX41X1_HVT U189 ( .A1(n578), .A3(n436), .A2(n579), .A4(n528), .S0(n475), 
        .S1(n468), .Y(n577) );
  MUX41X1_HVT U193 ( .A1(n724), .A3(n731), .A2(n717), .A4(n575), .S0(n238), 
        .S1(n501), .Y(n574) );
  MUX41X1_HVT U194 ( .A1(n725), .A3(n739), .A2(n19), .A4(n337), .S0(n475), 
        .S1(n414), .Y(n573) );
  MUX41X1_HVT U195 ( .A1(n422), .A3(n541), .A2(n349), .A4(n729), .S0(n470), 
        .S1(n499), .Y(n572) );
  AO21X1_HVT U197 ( .A1(n462), .A2(n476), .A3(n538), .Y(n570) );
  MUX41X1_HVT U205 ( .A1(n447), .A3(n210), .A2(n533), .A4(n543), .S0(n380), 
        .S1(n501), .Y(n562) );
  NAND2X0_HVT U212 ( .A1(n357), .A2(n754), .Y(n709) );
  NAND2X0_HVT U214 ( .A1(n422), .A2(n494), .Y(n560) );
  NAND2X0_HVT U215 ( .A1(n652), .A2(n486), .Y(n559) );
  NAND2X0_HVT U218 ( .A1(n540), .A2(n365), .Y(n613) );
  NAND2X0_HVT U220 ( .A1(n476), .A2(n560), .Y(n684) );
  INVX0_HVT U242 ( .A(n724), .Y(n549) );
  INVX0_HVT U245 ( .A(n757), .Y(n547) );
  INVX0_HVT U256 ( .A(n613), .Y(n538) );
  INVX0_HVT U258 ( .A(n738), .Y(n537) );
  INVX0_HVT U261 ( .A(n551), .Y(n534) );
  INVX0_HVT U265 ( .A(n740), .Y(n531) );
  INVX0_HVT U267 ( .A(n752), .Y(n530) );
  INVX0_HVT U268 ( .A(n744), .Y(n529) );
  INVX0_HVT U270 ( .A(n559), .Y(n528) );
  INVX0_HVT U278 ( .A(n733), .Y(n523) );
  INVX0_HVT U284 ( .A(n560), .Y(n520) );
  INVX0_HVT U285 ( .A(n557), .Y(n519) );
  INVX0_HVT U295 ( .A(n759), .Y(n515) );
  INVX0_HVT U306 ( .A(n597), .Y(n507) );
  OR2X1_HVT U1 ( .A1(n378), .A2(n441), .Y(n273) );
  OR2X1_HVT U2 ( .A1(n378), .A2(n441), .Y(n652) );
  MUX21X1_HVT U3 ( .A1(n447), .A2(n484), .S0(n283), .Y(n736) );
  NBUFFX2_HVT U6 ( .A(n754), .Y(n486) );
  INVX1_HVT U7 ( .A(n479), .Y(n437) );
  OA21X1_HVT U8 ( .A1(n507), .A2(n502), .A3(n735), .Y(n619) );
  INVX1_HVT U9 ( .A(n273), .Y(n527) );
  INVX1_HVT U10 ( .A(n736), .Y(n536) );
  INVX1_HVT U11 ( .A(n348), .Y(n351) );
  INVX0_HVT U12 ( .A(n750), .Y(n435) );
  INVX1_HVT U14 ( .A(n304), .Y(n755) );
  INVX1_HVT U16 ( .A(n756), .Y(n516) );
  MUX21X1_HVT U17 ( .A1(n714), .A2(n715), .S0(n475), .Y(n712) );
  MUX21X1_HVT U18 ( .A1(n535), .A2(n211), .S0(n413), .Y(n655) );
  AND2X1_HVT U19 ( .A1(n421), .A2(n709), .Y(n7) );
  AND2X1_HVT U20 ( .A1(n280), .A2(n282), .Y(n17) );
  INVX0_HVT U22 ( .A(n283), .Y(n224) );
  INVX1_HVT U23 ( .A(n496), .Y(n413) );
  AND2X1_HVT U24 ( .A1(n50), .A2(n118), .Y(n19) );
  AND2X1_HVT U25 ( .A1(n410), .A2(n409), .Y(n23) );
  INVX1_HVT U26 ( .A(n480), .Y(n451) );
  INVX1_HVT U27 ( .A(n421), .Y(n422) );
  NAND2X0_HVT U28 ( .A1(n451), .A2(n415), .Y(n50) );
  NAND2X0_HVT U29 ( .A1(n434), .A2(n224), .Y(n118) );
  INVX1_HVT U30 ( .A(n493), .Y(n430) );
  INVX1_HVT U31 ( .A(n730), .Y(n535) );
  MUX21X1_HVT U32 ( .A1(n458), .A2(n545), .S0(n492), .Y(n730) );
  MUX21X2_HVT U34 ( .A1(n747), .A2(n522), .S0(n470), .Y(n632) );
  INVX0_HVT U35 ( .A(n354), .Y(n119) );
  INVX1_HVT U36 ( .A(in[1]), .Y(n354) );
  MUX41X1_HVT U37 ( .A1(n565), .A3(n563), .A2(n564), .A4(n562), .S0(n412), 
        .S1(n446), .Y(n561) );
  NBUFFX2_HVT U38 ( .A(n760), .Y(n210) );
  NBUFFX2_HVT U39 ( .A(n760), .Y(n211) );
  INVX1_HVT U40 ( .A(n236), .Y(n305) );
  INVX1_HVT U41 ( .A(n233), .Y(n236) );
  INVX0_HVT U43 ( .A(n233), .Y(n283) );
  NOR2X0_HVT U44 ( .A1(n484), .A2(n492), .Y(n363) );
  INVX1_HVT U45 ( .A(n502), .Y(n455) );
  INVX1_HVT U46 ( .A(n119), .Y(n494) );
  INVX1_HVT U47 ( .A(n377), .Y(n454) );
  MUX21X1_HVT U48 ( .A1(n614), .A2(n615), .S0(n471), .Y(n612) );
  MUX21X1_HVT U49 ( .A1(n434), .A2(n427), .S0(n404), .Y(n615) );
  NBUFFX2_HVT U50 ( .A(n426), .Y(n443) );
  INVX1_HVT U51 ( .A(n493), .Y(n431) );
  INVX1_HVT U52 ( .A(n283), .Y(n492) );
  INVX1_HVT U54 ( .A(n496), .Y(n414) );
  NBUFFX2_HVT U55 ( .A(n500), .Y(n475) );
  INVX1_HVT U59 ( .A(n293), .Y(n502) );
  INVX1_HVT U60 ( .A(n293), .Y(n377) );
  INVX1_HVT U61 ( .A(n367), .Y(n441) );
  MUX21X1_HVT U63 ( .A1(n452), .A2(n306), .S0(n305), .Y(n427) );
  INVX1_HVT U64 ( .A(n363), .Y(n742) );
  MUX21X1_HVT U65 ( .A1(n485), .A2(n482), .S0(n307), .Y(n694) );
  XOR2X1_HVT U66 ( .A1(n438), .A2(n502), .Y(n719) );
  AO21X1_HVT U67 ( .A1(n477), .A2(n671), .A3(n538), .Y(n672) );
  XNOR2X1_HVT U69 ( .A1(n365), .A2(n414), .Y(n467) );
  INVX1_HVT U70 ( .A(n502), .Y(n498) );
  INVX1_HVT U71 ( .A(n340), .Y(n727) );
  INVX1_HVT U72 ( .A(n383), .Y(n753) );
  MUX21X1_HVT U74 ( .A1(n686), .A2(n685), .S0(n426), .Y(n683) );
  INVX1_HVT U76 ( .A(n468), .Y(n272) );
  INVX1_HVT U79 ( .A(n552), .Y(n509) );
  INVX1_HVT U80 ( .A(n457), .Y(n238) );
  MUX21X1_HVT U81 ( .A1(n321), .A2(n540), .S0(n415), .Y(n600) );
  MUX21X1_HVT U82 ( .A1(n595), .A2(n594), .S0(n470), .Y(n593) );
  MUX21X1_HVT U87 ( .A1(n609), .A2(n608), .S0(n398), .Y(n607) );
  NBUFFX2_HVT U88 ( .A(n458), .Y(n447) );
  NAND2X0_HVT U89 ( .A1(n448), .A2(n322), .Y(n760) );
  MUX21X1_HVT U91 ( .A1(n504), .A2(n630), .S0(n470), .Y(n629) );
  MUX21X1_HVT U92 ( .A1(n759), .A2(n626), .S0(n398), .Y(n625) );
  INVX1_HVT U93 ( .A(n726), .Y(n506) );
  INVX1_HVT U94 ( .A(n472), .Y(n326) );
  INVX0_HVT U95 ( .A(n503), .Y(n499) );
  INVX1_HVT U96 ( .A(in[7]), .Y(n503) );
  NBUFFX2_HVT U97 ( .A(n413), .Y(n470) );
  INVX1_HVT U98 ( .A(n414), .Y(n438) );
  INVX1_HVT U99 ( .A(n411), .Y(n357) );
  INVX0_HVT U100 ( .A(n236), .Y(n307) );
  INVX0_HVT U102 ( .A(n501), .Y(n429) );
  INVX1_HVT U104 ( .A(n354), .Y(n233) );
  NBUFFX2_HVT U106 ( .A(n500), .Y(n476) );
  INVX0_HVT U107 ( .A(n493), .Y(n448) );
  INVX1_HVT U108 ( .A(n473), .Y(n439) );
  INVX1_HVT U109 ( .A(n451), .Y(n323) );
  INVX0_HVT U111 ( .A(n432), .Y(n749) );
  AND2X1_HVT U112 ( .A1(n401), .A2(n402), .Y(n212) );
  INVX1_HVT U113 ( .A(in[6]), .Y(n342) );
  INVX1_HVT U114 ( .A(n293), .Y(n444) );
  INVX0_HVT U116 ( .A(n503), .Y(n500) );
  INVX1_HVT U117 ( .A(n503), .Y(n501) );
  NBUFFX2_HVT U118 ( .A(n500), .Y(n477) );
  INVX0_HVT U119 ( .A(n433), .Y(n213) );
  INVX0_HVT U120 ( .A(n489), .Y(n433) );
  MUX21X1_HVT U121 ( .A1(n567), .A2(n566), .S0(n438), .Y(n565) );
  NBUFFX2_HVT U122 ( .A(n488), .Y(n216) );
  NBUFFX2_HVT U123 ( .A(n367), .Y(n488) );
  INVX1_HVT U124 ( .A(n366), .Y(n367) );
  MUX21X1_HVT U125 ( .A1(n543), .A2(n749), .S0(n471), .Y(n665) );
  XOR2X1_HVT U126 ( .A1(n310), .A2(n224), .Y(n720) );
  INVX0_HVT U127 ( .A(n469), .Y(n261) );
  INVX0_HVT U129 ( .A(n469), .Y(n453) );
  INVX0_HVT U130 ( .A(n495), .Y(n457) );
  MUX21X1_HVT U132 ( .A1(n525), .A2(n433), .S0(n449), .Y(n591) );
  MUX41X1_HVT U133 ( .A1(n574), .A3(n572), .A2(n573), .A4(n569), .S0(n412), 
        .S1(n439), .Y(n568) );
  NAND2X0_HVT U134 ( .A1(n415), .A2(n540), .Y(n217) );
  NAND2X0_HVT U136 ( .A1(n365), .A2(n337), .Y(n218) );
  NAND2X0_HVT U137 ( .A1(n217), .A2(n218), .Y(n721) );
  INVX1_HVT U138 ( .A(n485), .Y(n540) );
  MUX21X2_HVT U139 ( .A1(n461), .A2(n450), .S0(n414), .Y(n633) );
  MUX21X1_HVT U141 ( .A1(n366), .A2(n313), .S0(n305), .Y(n304) );
  INVX0_HVT U142 ( .A(n734), .Y(n522) );
  MUX21X1_HVT U143 ( .A1(n367), .A2(n341), .S0(n411), .Y(n340) );
  MUX41X1_HVT U144 ( .A1(n599), .A3(n601), .A2(n593), .A4(n596), .S0(n473), 
        .S1(n412), .Y(n592) );
  INVX1_HVT U145 ( .A(n748), .Y(n514) );
  INVX1_HVT U146 ( .A(n548), .Y(n268) );
  INVX1_HVT U147 ( .A(n268), .Y(n313) );
  INVX1_HVT U148 ( .A(n486), .Y(n434) );
  MUX21X1_HVT U149 ( .A1(n484), .A2(n508), .S0(n307), .Y(n726) );
  INVX0_HVT U150 ( .A(n484), .Y(n428) );
  MUX41X1_HVT U151 ( .A1(n636), .A3(n631), .A2(n650), .A4(n644), .S0(n412), 
        .S1(in[6]), .Y(out[3]) );
  INVX1_HVT U152 ( .A(n310), .Y(n421) );
  NAND2X0_HVT U155 ( .A1(n383), .A2(n474), .Y(n219) );
  NAND2X0_HVT U156 ( .A1(n219), .A2(n274), .Y(n699) );
  MUX21X1_HVT U157 ( .A1(n428), .A2(n350), .S0(n448), .Y(n383) );
  NBUFFX2_HVT U159 ( .A(n497), .Y(n474) );
  INVX0_HVT U160 ( .A(n692), .Y(n546) );
  INVX0_HVT U161 ( .A(n762), .Y(n348) );
  INVX0_HVT U163 ( .A(n119), .Y(n493) );
  INVX0_HVT U164 ( .A(n745), .Y(n512) );
  INVX1_HVT U169 ( .A(n452), .Y(n341) );
  MUX41X1_HVT U170 ( .A1(n423), .A3(n463), .A2(n323), .A4(n450), .S0(n403), 
        .S1(n472), .Y(n704) );
  INVX1_HVT U171 ( .A(in[4]), .Y(n532) );
  MUX41X1_HVT U172 ( .A1(n733), .A3(n730), .A2(n459), .A4(n509), .S0(n499), 
        .S1(n261), .Y(n627) );
  INVX0_HVT U173 ( .A(n210), .Y(n513) );
  INVX0_HVT U175 ( .A(n348), .Y(n349) );
  INVX1_HVT U181 ( .A(n484), .Y(n452) );
  INVX0_HVT U183 ( .A(n283), .Y(n449) );
  NAND2X0_HVT U184 ( .A1(n610), .A2(n227), .Y(n231) );
  NAND2X0_HVT U185 ( .A1(n322), .A2(n465), .Y(n232) );
  NAND2X0_HVT U186 ( .A1(n231), .A2(n232), .Y(n609) );
  INVX0_HVT U187 ( .A(n465), .Y(n227) );
  XOR2X1_HVT U188 ( .A1(n444), .A2(n236), .Y(n465) );
  MUX21X1_HVT U190 ( .A1(n728), .A2(n526), .S0(n475), .Y(n608) );
  INVX1_HVT U191 ( .A(n475), .Y(n403) );
  INVX0_HVT U192 ( .A(n762), .Y(n545) );
  INVX1_HVT U196 ( .A(n348), .Y(n350) );
  INVX0_HVT U198 ( .A(n492), .Y(n415) );
  INVX1_HVT U199 ( .A(n555), .Y(n539) );
  INVX1_HVT U200 ( .A(in[3]), .Y(n548) );
  INVX1_HVT U201 ( .A(n283), .Y(n491) );
  MUX41X1_HVT U202 ( .A1(n527), .A3(n337), .A2(n517), .A4(n323), .S0(n238), 
        .S1(n444), .Y(n621) );
  NBUFFX2_HVT U203 ( .A(n395), .Y(n487) );
  MUX21X1_HVT U204 ( .A1(n349), .A2(n447), .S0(n378), .Y(n550) );
  INVX0_HVT U206 ( .A(n378), .Y(n379) );
  MUX21X1_HVT U207 ( .A1(n341), .A2(n482), .S0(n357), .Y(n575) );
  NAND2X0_HVT U208 ( .A1(n540), .A2(n379), .Y(n242) );
  NAND2X0_HVT U209 ( .A1(n433), .A2(n345), .Y(n249) );
  NAND2X0_HVT U210 ( .A1(n242), .A2(n249), .Y(n432) );
  MUX41X1_HVT U211 ( .A1(n683), .A3(n682), .A2(n680), .A4(n678), .S0(n439), 
        .S1(n412), .Y(n677) );
  NAND2X0_HVT U213 ( .A1(n337), .A2(n500), .Y(n256) );
  NAND2X0_HVT U216 ( .A1(n745), .A2(n407), .Y(n258) );
  NAND2X0_HVT U217 ( .A1(n256), .A2(n258), .Y(n686) );
  MUX21X1_HVT U219 ( .A1(n425), .A2(n322), .S0(n357), .Y(n745) );
  INVX0_HVT U221 ( .A(n264), .Y(n739) );
  MUX21X1_HVT U222 ( .A1(n489), .A2(n346), .S0(n491), .Y(n264) );
  INVX0_HVT U223 ( .A(n489), .Y(n508) );
  INVX0_HVT U224 ( .A(n346), .Y(n347) );
  MUX21X1_HVT U225 ( .A1(n441), .A2(n480), .S0(n430), .Y(n440) );
  MUX21X2_HVT U226 ( .A1(n434), .A2(n304), .S0(n446), .Y(n698) );
  INVX1_HVT U227 ( .A(n532), .Y(n458) );
  INVX0_HVT U228 ( .A(n416), .Y(n728) );
  MUX41X1_HVT U229 ( .A1(n654), .A3(n651), .A2(n655), .A4(n23), .S0(n446), 
        .S1(n502), .Y(n650) );
  NAND2X0_HVT U230 ( .A1(n482), .A2(n345), .Y(n269) );
  NAND2X0_HVT U231 ( .A1(n269), .A2(n290), .Y(n423) );
  MUX41X1_HVT U232 ( .A1(n512), .A3(n721), .A2(n749), .A4(n363), .S0(n272), 
        .S1(n455), .Y(n682) );
  INVX1_HVT U233 ( .A(n558), .Y(n510) );
  INVX1_HVT U234 ( .A(n546), .Y(n274) );
  NAND2X0_HVT U235 ( .A1(n357), .A2(n349), .Y(n692) );
  MUX41X1_HVT U236 ( .A1(n580), .A3(n584), .A2(n577), .A4(n581), .S0(n478), 
        .S1(n439), .Y(n576) );
  OA21X1_HVT U237 ( .A1(n732), .A2(n502), .A3(n517), .Y(n582) );
  INVX1_HVT U238 ( .A(n758), .Y(n366) );
  MUX41X1_HVT U239 ( .A1(n587), .A3(n586), .A2(n590), .A4(n588), .S0(n439), 
        .S1(n478), .Y(n585) );
  MUX21X1_HVT U240 ( .A1(n350), .A2(n341), .S0(n378), .Y(n578) );
  NAND2X0_HVT U241 ( .A1(n645), .A2(n439), .Y(n278) );
  NAND2X0_HVT U243 ( .A1(n648), .A2(n472), .Y(n279) );
  NAND2X0_HVT U244 ( .A1(n278), .A2(n279), .Y(n644) );
  INVX1_HVT U246 ( .A(n550), .Y(n533) );
  MUX41X1_HVT U247 ( .A1(n623), .A3(n522), .A2(n741), .A4(n416), .S0(n238), 
        .S1(n404), .Y(n622) );
  INVX0_HVT U248 ( .A(n411), .Y(n358) );
  INVX1_HVT U249 ( .A(in[2]), .Y(n496) );
  INVX1_HVT U250 ( .A(n438), .Y(n380) );
  INVX0_HVT U251 ( .A(n452), .Y(n329) );
  NBUFFX2_HVT U252 ( .A(n532), .Y(n481) );
  AND3X1_HVT U253 ( .A1(n213), .A2(n709), .A3(n684), .Y(n685) );
  INVX0_HVT U254 ( .A(n424), .Y(n731) );
  NOR2X0_HVT U255 ( .A1(n425), .A2(n365), .Y(n424) );
  INVX0_HVT U257 ( .A(n389), .Y(n425) );
  MUX41X1_HVT U259 ( .A1(n675), .A3(n668), .A2(n670), .A4(n667), .S0(n412), 
        .S1(n439), .Y(n666) );
  NAND2X0_HVT U260 ( .A1(n452), .A2(n365), .Y(n280) );
  NAND2X0_HVT U262 ( .A1(n451), .A2(n345), .Y(n282) );
  NAND2X0_HVT U263 ( .A1(n280), .A2(n282), .Y(n450) );
  OR2X1_HVT U264 ( .A1(n327), .A2(n364), .Y(n754) );
  INVX1_HVT U266 ( .A(n467), .Y(n408) );
  NAND2X0_HVT U269 ( .A1(n350), .A2(n236), .Y(n285) );
  NAND2X0_HVT U271 ( .A1(n754), .A2(n448), .Y(n290) );
  NAND2X0_HVT U272 ( .A1(n285), .A2(n290), .Y(n735) );
  MUX21X1_HVT U273 ( .A1(n735), .A2(n653), .S0(n426), .Y(n651) );
  INVX0_HVT U274 ( .A(n735), .Y(n543) );
  OA21X1_HVT U275 ( .A1(n464), .A2(n502), .A3(n735), .Y(n594) );
  MUX41X1_HVT U276 ( .A1(n516), .A3(n524), .A2(n744), .A4(n466), .S0(n238), 
        .S1(n444), .Y(n637) );
  INVX1_HVT U277 ( .A(n503), .Y(n293) );
  INVX0_HVT U279 ( .A(n671), .Y(n526) );
  MUX41X1_HVT U280 ( .A1(n607), .A3(n605), .A2(n612), .A4(n611), .S0(n439), 
        .S1(n478), .Y(n604) );
  NAND2X0_HVT U281 ( .A1(n708), .A2(n469), .Y(n297) );
  NAND2X0_HVT U282 ( .A1(n706), .A2(n453), .Y(n301) );
  NAND2X0_HVT U283 ( .A1(n297), .A2(n301), .Y(n705) );
  NAND2X0_HVT U286 ( .A1(n399), .A2(n400), .Y(out[1]) );
  INVX1_HVT U287 ( .A(n342), .Y(n303) );
  NAND2X0_HVT U288 ( .A1(n368), .A2(n369), .Y(out[4]) );
  NAND2X0_HVT U289 ( .A1(n314), .A2(n315), .Y(n306) );
  NAND2X0_HVT U290 ( .A1(n322), .A2(n227), .Y(n308) );
  NAND2X0_HVT U291 ( .A1(n674), .A2(n465), .Y(n309) );
  NAND2X0_HVT U292 ( .A1(n308), .A2(n309), .Y(n673) );
  MUX41X1_HVT U293 ( .A1(n720), .A3(n274), .A2(n542), .A4(n509), .S0(n502), 
        .S1(n261), .Y(n617) );
  AND2X1_HVT U294 ( .A1(n314), .A2(n315), .Y(n310) );
  MUX41X1_HVT U296 ( .A1(n628), .A3(n625), .A2(n629), .A4(n627), .S0(n412), 
        .S1(n497), .Y(n624) );
  MUX21X1_HVT U297 ( .A1(n736), .A2(n559), .S0(n475), .Y(n554) );
  MUX41X1_HVT U298 ( .A1(n514), .A3(n703), .A2(n432), .A4(n521), .S0(n429), 
        .S1(n472), .Y(n702) );
  NAND2X0_HVT U299 ( .A1(n479), .A2(n345), .Y(n311) );
  NAND2X0_HVT U300 ( .A1(n428), .A2(n430), .Y(n312) );
  NAND2X0_HVT U301 ( .A1(n311), .A2(n312), .Y(n743) );
  INVX0_HVT U302 ( .A(n743), .Y(n517) );
  MUX21X1_HVT U303 ( .A1(n447), .A2(n525), .S0(n415), .Y(n734) );
  INVX0_HVT U304 ( .A(n236), .Y(n365) );
  NOR2X1_HVT U305 ( .A1(n428), .A2(n491), .Y(n466) );
  INVX0_HVT U307 ( .A(n430), .Y(n345) );
  NAND2X0_HVT U308 ( .A1(n364), .A2(n268), .Y(n314) );
  NAND2X0_HVT U309 ( .A1(n458), .A2(n313), .Y(n315) );
  NAND2X0_HVT U310 ( .A1(n314), .A2(n315), .Y(n445) );
  NBUFFX2_HVT U311 ( .A(n445), .Y(n480) );
  INVX1_HVT U312 ( .A(n366), .Y(n316) );
  NAND2X0_HVT U313 ( .A1(n642), .A2(n403), .Y(n317) );
  NAND2X0_HVT U314 ( .A1(n641), .A2(n476), .Y(n318) );
  NAND2X0_HVT U315 ( .A1(n317), .A2(n318), .Y(n638) );
  MUX21X1_HVT U316 ( .A1(n643), .A2(n523), .S0(n453), .Y(n642) );
  INVX0_HVT U317 ( .A(n423), .Y(n747) );
  NAND2X0_HVT U318 ( .A1(n7), .A2(n476), .Y(n319) );
  NAND2X0_HVT U319 ( .A1(n17), .A2(n403), .Y(n320) );
  NAND2X0_HVT U320 ( .A1(n319), .A2(n320), .Y(n567) );
  INVX0_HVT U321 ( .A(n761), .Y(n321) );
  INVX1_HVT U322 ( .A(n321), .Y(n322) );
  MUX21X1_HVT U323 ( .A1(n490), .A2(n306), .S0(n307), .Y(n725) );
  INVX0_HVT U324 ( .A(n741), .Y(n505) );
  NAND2X0_HVT U325 ( .A1(n619), .A2(n413), .Y(n324) );
  NAND2X0_HVT U326 ( .A1(n620), .A2(n272), .Y(n325) );
  NAND2X0_HVT U327 ( .A1(n325), .A2(n324), .Y(n618) );
  MUX21X1_HVT U328 ( .A1(n737), .A2(n513), .S0(n477), .Y(n620) );
  INVX0_HVT U329 ( .A(n328), .Y(n746) );
  MUX41X1_HVT U330 ( .A1(n442), .A3(n464), .A2(n707), .A4(n466), .S0(n407), 
        .S1(n326), .Y(n706) );
  INVX0_HVT U331 ( .A(n476), .Y(n404) );
  INVX1_HVT U332 ( .A(n316), .Y(n525) );
  MUX41X1_HVT U333 ( .A1(n742), .A3(n693), .A2(n740), .A4(n694), .S0(n453), 
        .S1(n377), .Y(n691) );
  INVX0_HVT U334 ( .A(n725), .Y(n511) );
  MUX21X1_HVT U335 ( .A1(n347), .A2(n479), .S0(n358), .Y(n603) );
  MUX21X1_HVT U336 ( .A1(n306), .A2(n545), .S0(n492), .Y(n756) );
  NBUFFX2_HVT U337 ( .A(n532), .Y(n364) );
  MUX21X1_HVT U338 ( .A1(n389), .A2(n329), .S0(n307), .Y(n643) );
  MUX41X1_HVT U339 ( .A1(n505), .A3(n735), .A2(n751), .A4(n649), .S0(n238), 
        .S1(n444), .Y(n648) );
  INVX1_HVT U340 ( .A(n473), .Y(n446) );
  INVX0_HVT U341 ( .A(n440), .Y(n729) );
  INVX1_HVT U342 ( .A(n483), .Y(n327) );
  NBUFFX2_HVT U343 ( .A(n548), .Y(n483) );
  MUX21X1_HVT U344 ( .A1(n490), .A2(n329), .S0(n431), .Y(n328) );
  NAND2X0_HVT U345 ( .A1(n530), .A2(n446), .Y(n330) );
  NAND2X0_HVT U346 ( .A1(n494), .A2(n474), .Y(n331) );
  NAND2X0_HVT U347 ( .A1(n330), .A2(n331), .Y(n700) );
  NAND2X0_HVT U348 ( .A1(n488), .A2(n378), .Y(n332) );
  NAND2X0_HVT U349 ( .A1(n329), .A2(n431), .Y(n333) );
  NAND2X0_HVT U350 ( .A1(n332), .A2(n333), .Y(n752) );
  MUX21X1_HVT U351 ( .A1(n341), .A2(n481), .S0(n426), .Y(n334) );
  NAND2X0_HVT U352 ( .A1(n592), .A2(n342), .Y(n335) );
  NAND2X0_HVT U353 ( .A1(n604), .A2(n303), .Y(n336) );
  NAND2X0_HVT U354 ( .A1(n336), .A2(n335), .Y(out[5]) );
  NBUFFX2_HVT U355 ( .A(n395), .Y(n337) );
  NAND2X0_HVT U356 ( .A1(n743), .A2(n404), .Y(n338) );
  NAND2X0_HVT U357 ( .A1(n340), .A2(n476), .Y(n339) );
  NAND2X0_HVT U358 ( .A1(n338), .A2(n339), .Y(n626) );
  MUX41X1_HVT U359 ( .A1(n711), .A3(n701), .A2(n705), .A4(n697), .S0(n342), 
        .S1(n412), .Y(out[0]) );
  INVX1_HVT U360 ( .A(in[0]), .Y(n412) );
  NAND2X0_HVT U361 ( .A1(n704), .A2(n469), .Y(n343) );
  NAND2X0_HVT U362 ( .A1(n702), .A2(n398), .Y(n344) );
  NAND2X0_HVT U363 ( .A1(n343), .A2(n344), .Y(n701) );
  INVX1_HVT U364 ( .A(n661), .Y(n518) );
  INVX0_HVT U365 ( .A(n545), .Y(n346) );
  NAND2X0_HVT U366 ( .A1(n646), .A2(n429), .Y(n352) );
  NAND2X0_HVT U367 ( .A1(n647), .A2(n476), .Y(n353) );
  NAND2X0_HVT U368 ( .A1(n352), .A2(n353), .Y(n645) );
  AO21X1_HVT U369 ( .A1(n471), .A2(n487), .A3(n437), .Y(n646) );
  MUX21X1_HVT U370 ( .A1(n424), .A2(n544), .S0(n238), .Y(n647) );
  INVX0_HVT U371 ( .A(n732), .Y(n544) );
  MUX41X1_HVT U372 ( .A1(n602), .A3(n423), .A2(n603), .A4(n461), .S0(n398), 
        .S1(n454), .Y(n601) );
  MUX41X1_HVT U373 ( .A1(n544), .A3(n710), .A2(n743), .A4(n751), .S0(n429), 
        .S1(n380), .Y(n563) );
  NAND2X0_HVT U374 ( .A1(n656), .A2(n342), .Y(n355) );
  NAND2X0_HVT U375 ( .A1(n666), .A2(n303), .Y(n356) );
  NAND2X0_HVT U376 ( .A1(n356), .A2(n355), .Y(out[2]) );
  NAND2X0_HVT U377 ( .A1(n377), .A2(n264), .Y(n359) );
  NAND2X0_HVT U378 ( .A1(n454), .A2(n739), .Y(n360) );
  NAND2X0_HVT U379 ( .A1(n359), .A2(n360), .Y(n722) );
  INVX0_HVT U380 ( .A(n477), .Y(n407) );
  NAND2X0_HVT U381 ( .A1(n663), .A2(n398), .Y(n361) );
  NAND2X0_HVT U382 ( .A1(n504), .A2(n470), .Y(n362) );
  NAND2X0_HVT U383 ( .A1(n361), .A2(n362), .Y(n660) );
  MUX41X1_HVT U384 ( .A1(n460), .A3(n542), .A2(n748), .A4(n449), .S0(n398), 
        .S1(n498), .Y(n667) );
  INVX1_HVT U385 ( .A(n556), .Y(n541) );
  NBUFFX2_HVT U386 ( .A(n364), .Y(n482) );
  NBUFFX2_HVT U387 ( .A(n364), .Y(n389) );
  MUX21X1_HVT U388 ( .A1(n479), .A2(n525), .S0(n431), .Y(n669) );
  NAND2X0_HVT U389 ( .A1(n640), .A2(n639), .Y(n641) );
  NAND2X0_HVT U390 ( .A1(n616), .A2(n342), .Y(n368) );
  NAND2X0_HVT U391 ( .A1(n624), .A2(n303), .Y(n369) );
  MUX41X1_HVT U392 ( .A1(n657), .A3(n660), .A2(n659), .A4(n664), .S0(n478), 
        .S1(n474), .Y(n656) );
  INVX0_HVT U393 ( .A(n370), .Y(n595) );
  MUX41X1_HVT U394 ( .A1(n621), .A3(n617), .A2(n622), .A4(n618), .S0(n412), 
        .S1(n472), .Y(n616) );
  MUX21X1_HVT U395 ( .A1(n540), .A2(n556), .S0(n477), .Y(n370) );
  INVX1_HVT U396 ( .A(n496), .Y(n495) );
  MUX41X1_HVT U397 ( .A1(n669), .A3(n541), .A2(n460), .A4(n363), .S0(n453), 
        .S1(n407), .Y(n668) );
  NAND2X0_HVT U398 ( .A1(n537), .A2(n453), .Y(n371) );
  NAND2X0_HVT U399 ( .A1(n736), .A2(n380), .Y(n372) );
  NAND2X0_HVT U400 ( .A1(n371), .A2(n372), .Y(n635) );
  INVX1_HVT U401 ( .A(n554), .Y(n504) );
  INVX0_HVT U402 ( .A(n394), .Y(n737) );
  NAND2X0_HVT U403 ( .A1(n672), .A2(n272), .Y(n373) );
  NAND2X0_HVT U404 ( .A1(n673), .A2(n471), .Y(n374) );
  NAND2X0_HVT U405 ( .A1(n373), .A2(n374), .Y(n670) );
  NAND2X0_HVT U406 ( .A1(n696), .A2(n469), .Y(n375) );
  NAND2X0_HVT U407 ( .A1(n722), .A2(n398), .Y(n376) );
  NAND2X0_HVT U408 ( .A1(n375), .A2(n376), .Y(n695) );
  MUX21X1_HVT U409 ( .A1(n347), .A2(n329), .S0(n224), .Y(n732) );
  INVX0_HVT U410 ( .A(n448), .Y(n378) );
  NAND2X0_HVT U411 ( .A1(n712), .A2(n272), .Y(n381) );
  NAND2X0_HVT U412 ( .A1(n716), .A2(n470), .Y(n382) );
  NAND2X0_HVT U413 ( .A1(n381), .A2(n382), .Y(n711) );
  NAND2X0_HVT U414 ( .A1(n463), .A2(n384), .Y(n385) );
  NAND2X0_HVT U415 ( .A1(n665), .A2(n719), .Y(n386) );
  NAND2X0_HVT U416 ( .A1(n386), .A2(n385), .Y(n664) );
  INVX0_HVT U417 ( .A(n719), .Y(n384) );
  INVX1_HVT U418 ( .A(n471), .Y(n398) );
  INVX1_HVT U419 ( .A(n709), .Y(n542) );
  NAND2X0_HVT U420 ( .A1(n576), .A2(n342), .Y(n387) );
  NAND2X0_HVT U421 ( .A1(n585), .A2(n303), .Y(n388) );
  NAND2X0_HVT U422 ( .A1(n388), .A2(n387), .Y(out[6]) );
  NAND2X0_HVT U423 ( .A1(n583), .A2(n413), .Y(n390) );
  NAND2X0_HVT U424 ( .A1(n582), .A2(n438), .Y(n391) );
  NAND2X0_HVT U425 ( .A1(n390), .A2(n391), .Y(n581) );
  NAND2X0_HVT U426 ( .A1(n487), .A2(n499), .Y(n392) );
  NAND2X0_HVT U427 ( .A1(n524), .A2(n404), .Y(n393) );
  NAND2X0_HVT U428 ( .A1(n392), .A2(n393), .Y(n630) );
  MUX21X1_HVT U429 ( .A1(n754), .A2(n316), .S0(n430), .Y(n442) );
  MUX21X1_HVT U430 ( .A1(n425), .A2(n488), .S0(n449), .Y(n394) );
  NAND2X0_HVT U431 ( .A1(n458), .A2(n483), .Y(n395) );
  NAND2X0_HVT U432 ( .A1(n327), .A2(n477), .Y(n396) );
  NAND2X0_HVT U433 ( .A1(n679), .A2(n429), .Y(n397) );
  NAND2X0_HVT U434 ( .A1(n396), .A2(n397), .Y(n583) );
  INVX1_HVT U435 ( .A(n553), .Y(n524) );
  NAND2X0_HVT U436 ( .A1(n677), .A2(n342), .Y(n399) );
  NAND2X0_HVT U437 ( .A1(n687), .A2(in[6]), .Y(n400) );
  NAND2X0_HVT U438 ( .A1(n422), .A2(n238), .Y(n401) );
  NAND2X0_HVT U439 ( .A1(n521), .A2(n438), .Y(n402) );
  NBUFFX2_HVT U440 ( .A(n497), .Y(n473) );
  NAND2X0_HVT U441 ( .A1(n637), .A2(n446), .Y(n405) );
  NAND2X0_HVT U442 ( .A1(n638), .A2(n474), .Y(n406) );
  NAND2X0_HVT U443 ( .A1(n406), .A2(n405), .Y(n636) );
  NAND2X0_HVT U444 ( .A1(n433), .A2(n408), .Y(n409) );
  NAND2X0_HVT U445 ( .A1(n334), .A2(n467), .Y(n410) );
  NBUFFX2_HVT U446 ( .A(n493), .Y(n411) );
  OA21X1_HVT U447 ( .A1(n398), .A2(n440), .A3(n442), .Y(n654) );
  OA21X1_HVT U448 ( .A1(n726), .A2(n377), .A3(n613), .Y(n614) );
  MUX21X1_HVT U449 ( .A1(n349), .A2(n316), .S0(n430), .Y(n416) );
  NAND2X0_HVT U450 ( .A1(n571), .A2(n272), .Y(n417) );
  NAND2X0_HVT U451 ( .A1(n570), .A2(n469), .Y(n418) );
  NAND2X0_HVT U452 ( .A1(n417), .A2(n418), .Y(n569) );
  NAND2X0_HVT U453 ( .A1(n561), .A2(n342), .Y(n419) );
  NAND2X0_HVT U454 ( .A1(n568), .A2(n303), .Y(n420) );
  NAND2X0_HVT U455 ( .A1(n419), .A2(n420), .Y(out[7]) );
  MUX21X1_HVT U456 ( .A1(n549), .A2(n534), .S0(n476), .Y(n571) );
  INVX1_HVT U457 ( .A(n438), .Y(n426) );
  MUX21X1_HVT U458 ( .A1(n310), .A2(n321), .S0(n431), .Y(n741) );
  MUX21X1_HVT U459 ( .A1(n456), .A2(n212), .S0(n377), .Y(n605) );
  INVX0_HVT U460 ( .A(n751), .Y(n521) );
  AO21X1_HVT U461 ( .A1(n494), .A2(n540), .A3(n404), .Y(n662) );
  INVX0_HVT U462 ( .A(n435), .Y(n436) );
  MUX41X1_HVT U463 ( .A1(n720), .A3(n274), .A2(n727), .A4(n460), .S0(n272), 
        .S1(n403), .Y(n580) );
  OA21X1_HVT U464 ( .A1(n407), .A2(n756), .A3(n416), .Y(n566) );
  MUX41X1_HVT U465 ( .A1(n512), .A3(n328), .A2(n529), .A4(n510), .S0(n429), 
        .S1(n326), .Y(n716) );
  MUX21X1_HVT U466 ( .A1(n606), .A2(n547), .S0(n414), .Y(n456) );
  MUX41X1_HVT U467 ( .A1(n734), .A3(n752), .A2(n506), .A4(n730), .S0(n272), 
        .S1(n377), .Y(n564) );
  NBUFFX2_HVT U468 ( .A(n445), .Y(n479) );
  MUX21X1_HVT U469 ( .A1(n525), .A2(n545), .S0(n474), .Y(n713) );
  AND2X1_HVT U470 ( .A1(n213), .A2(n692), .Y(n459) );
  MUX21X1_HVT U471 ( .A1(n323), .A2(n389), .S0(n358), .Y(n661) );
  MUX21X1_HVT U472 ( .A1(n488), .A2(n337), .S0(n449), .Y(n676) );
  NAND2X0_HVT U473 ( .A1(n481), .A2(n483), .Y(n758) );
  NBUFFX2_HVT U474 ( .A(n761), .Y(n489) );
  MUX21X1_HVT U475 ( .A1(n451), .A2(n389), .S0(n431), .Y(n689) );
  MUX21X1_HVT U476 ( .A1(n525), .A2(n389), .S0(n224), .Y(n553) );
  NBUFFX2_HVT U477 ( .A(n761), .Y(n490) );
  XOR2X1_HVT U478 ( .A1(n489), .A2(n491), .Y(n717) );
  MUX21X1_HVT U479 ( .A1(n351), .A2(n489), .S0(n358), .Y(n579) );
  MUX21X1_HVT U480 ( .A1(n488), .A2(n351), .S0(n449), .Y(n671) );
  MUX21X1_HVT U481 ( .A1(n490), .A2(n482), .S0(n357), .Y(n558) );
  AND2X1_HVT U482 ( .A1(n379), .A2(n321), .Y(n460) );
  XNOR2X1_HVT U483 ( .A1(n316), .A2(n492), .Y(n461) );
  MUX21X1_HVT U484 ( .A1(n485), .A2(n329), .S0(n491), .Y(n556) );
  MUX21X1_HVT U485 ( .A1(n490), .A2(n367), .S0(n430), .Y(n552) );
  XNOR2X1_HVT U486 ( .A1(n350), .A2(n224), .Y(n462) );
  AND2X1_HVT U487 ( .A1(n351), .A2(n652), .Y(n463) );
  MUX21X1_HVT U488 ( .A1(n486), .A2(n351), .S0(n470), .Y(n640) );
  XOR2X1_HVT U489 ( .A1(n389), .A2(n305), .Y(n740) );
  NBUFFX2_HVT U490 ( .A(n495), .Y(n468) );
  NBUFFX2_HVT U491 ( .A(n548), .Y(n484) );
  NBUFFX2_HVT U492 ( .A(in[5]), .Y(n472) );
  XOR2X1_HVT U493 ( .A1(n449), .A2(n452), .Y(n718) );
  MUX21X1_HVT U494 ( .A1(n486), .A2(n306), .S0(n307), .Y(n658) );
  NAND2X0_HVT U495 ( .A1(n481), .A2(n268), .Y(n761) );
  AND2X1_HVT U496 ( .A1(n479), .A2(n494), .Y(n464) );
  MUX21X1_HVT U497 ( .A1(n545), .A2(n541), .S0(n477), .Y(n696) );
  NBUFFX2_HVT U498 ( .A(n395), .Y(n485) );
  MUX21X1_HVT U499 ( .A1(n327), .A2(n731), .S0(n474), .Y(n715) );
  XOR2X1_HVT U500 ( .A1(n379), .A2(n473), .Y(n723) );
  MUX21X1_HVT U501 ( .A1(n428), .A2(n540), .S0(n365), .Y(n555) );
  MUX21X1_HVT U502 ( .A1(n211), .A2(n494), .S0(n469), .Y(n639) );
  MUX21X1_HVT U503 ( .A1(n428), .A2(n482), .S0(n477), .Y(n674) );
  NBUFFX2_HVT U504 ( .A(in[5]), .Y(n497) );
  NAND2X0_HVT U505 ( .A1(n458), .A2(n268), .Y(n762) );
  MUX21X1_HVT U506 ( .A1(n447), .A2(n422), .S0(n305), .Y(n557) );
  MUX21X1_HVT U507 ( .A1(n447), .A2(n487), .S0(n365), .Y(n551) );
  MUX21X1_HVT U508 ( .A1(n349), .A2(n447), .S0(n358), .Y(n738) );
  NBUFFX2_HVT U509 ( .A(in[0]), .Y(n478) );
  NBUFFX2_HVT U510 ( .A(n413), .Y(n469) );
  NBUFFX2_HVT U511 ( .A(n495), .Y(n471) );
endmodule

