
module inv_sbox_0 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n196, n197, n198, n199, n200, n201, n202, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405;

  NAND2X0_HVT U1 ( .A1(n291), .A2(n264), .Y(n1) );
  NAND2X0_HVT U5 ( .A1(n4), .A2(n218), .Y(n5) );
  NAND2X0_HVT U7 ( .A1(n260), .A2(n329), .Y(n8) );
  NAND2X0_HVT U8 ( .A1(n275), .A2(n222), .Y(n9) );
  NAND2X0_HVT U9 ( .A1(n334), .A2(n9), .Y(n10) );
  NAND2X0_HVT U10 ( .A1(n333), .A2(n12), .Y(n11) );
  NAND2X0_HVT U11 ( .A1(n255), .A2(n332), .Y(n13) );
  NAND2X0_HVT U12 ( .A1(n337), .A2(n316), .Y(n14) );
  NAND2X0_HVT U13 ( .A1(n329), .A2(n9), .Y(n15) );
  NAND2X0_HVT U15 ( .A1(n324), .A2(n276), .Y(n17) );
  NAND2X0_HVT U19 ( .A1(n336), .A2(n404), .Y(n22) );
  NAND2X0_HVT U25 ( .A1(n236), .A2(n316), .Y(n6) );
  NAND2X0_HVT U32 ( .A1(n229), .A2(n341), .Y(n34) );
  NAND2X0_HVT U35 ( .A1(n9), .A2(n292), .Y(n37) );
  NAND2X0_HVT U38 ( .A1(n242), .A2(n255), .Y(n40) );
  NAND2X0_HVT U42 ( .A1(n7), .A2(n239), .Y(n44) );
  OA21X1_HVT U53 ( .A1(n289), .A2(n52), .A3(n372), .Y(n54) );
  NAND2X0_HVT U55 ( .A1(n329), .A2(n4), .Y(n56) );
  MUX41X1_HVT U62 ( .A1(n63), .A3(n57), .A2(n59), .A4(n55), .S0(n323), .S1(
        n321), .Y(n64) );
  NAND2X0_HVT U66 ( .A1(n276), .A2(n283), .Y(n68) );
  MUX41X1_HVT U67 ( .A1(n362), .A3(n386), .A2(n364), .A4(n68), .S0(n314), .S1(
        n307), .Y(n69) );
  MUX41X1_HVT U68 ( .A1(n362), .A3(n226), .A2(n363), .A4(n334), .S0(n307), 
        .S1(n344), .Y(n70) );
  MUX41X1_HVT U71 ( .A1(n237), .A3(n286), .A2(n13), .A4(n358), .S0(n307), .S1(
        n344), .Y(n72) );
  NAND2X0_HVT U72 ( .A1(n240), .A2(n8), .Y(n73) );
  MUX41X1_HVT U73 ( .A1(n29), .A3(n73), .A2(n387), .A4(n242), .S0(n313), .S1(
        n305), .Y(n74) );
  MUX41X1_HVT U74 ( .A1(n11), .A3(n377), .A2(n376), .A4(n368), .S0(n308), .S1(
        n251), .Y(n75) );
  MUX41X1_HVT U78 ( .A1(n78), .A3(n74), .A2(n75), .A4(n72), .S0(n323), .S1(
        n321), .Y(n79) );
  MUX41X1_HVT U79 ( .A1(n373), .A3(n20), .A2(n375), .A4(n19), .S0(n308), .S1(
        n344), .Y(n80) );
  MUX41X1_HVT U80 ( .A1(n389), .A3(n385), .A2(n10), .A4(n5), .S0(n307), .S1(
        n251), .Y(n81) );
  NAND2X0_HVT U81 ( .A1(n332), .A2(n8), .Y(n82) );
  AND2X1_HVT U82 ( .A1(n237), .A2(n328), .Y(n83) );
  MUX41X1_HVT U83 ( .A1(n83), .A3(n374), .A2(n235), .A4(n82), .S0(n307), .S1(
        n344), .Y(n84) );
  MUX41X1_HVT U84 ( .A1(n302), .A3(n373), .A2(n391), .A4(n250), .S0(n308), 
        .S1(n252), .Y(n85) );
  MUX41X1_HVT U85 ( .A1(n85), .A3(n81), .A2(n84), .A4(n80), .S0(n323), .S1(
        n320), .Y(n86) );
  MUX41X1_HVT U87 ( .A1(n352), .A3(n302), .A2(n392), .A4(n284), .S0(n306), 
        .S1(n252), .Y(n87) );
  MUX41X1_HVT U88 ( .A1(n364), .A3(n349), .A2(n32), .A4(n48), .S0(n307), .S1(
        n251), .Y(n88) );
  NAND2X0_HVT U89 ( .A1(n255), .A2(n200), .Y(n89) );
  MUX41X1_HVT U90 ( .A1(n286), .A3(n8), .A2(n49), .A4(n89), .S0(n307), .S1(
        n277), .Y(n90) );
  MUX41X1_HVT U95 ( .A1(n94), .A3(n88), .A2(n90), .A4(n87), .S0(n323), .S1(
        in[1]), .Y(n95) );
  MUX41X1_HVT U96 ( .A1(n386), .A3(n15), .A2(n371), .A4(n393), .S0(n308), .S1(
        n343), .Y(n96) );
  MUX41X1_HVT U98 ( .A1(n97), .A3(n394), .A2(n378), .A4(n30), .S0(n308), .S1(
        n252), .Y(n98) );
  MUX41X1_HVT U99 ( .A1(n34), .A3(n366), .A2(n50), .A4(n325), .S0(n252), .S1(
        n305), .Y(n99) );
  NAND2X0_HVT U100 ( .A1(n341), .A2(n401), .Y(n100) );
  MUX41X1_HVT U101 ( .A1(n395), .A3(n14), .A2(n230), .A4(n100), .S0(n343), 
        .S1(n305), .Y(n101) );
  MUX41X1_HVT U102 ( .A1(n101), .A3(n98), .A2(n99), .A4(n96), .S0(in[5]), .S1(
        n321), .Y(n102) );
  AND2X1_HVT U104 ( .A1(n8), .A2(n222), .Y(n103) );
  MUX41X1_HVT U105 ( .A1(n16), .A3(n396), .A2(n82), .A4(n103), .S0(n308), .S1(
        n252), .Y(n104) );
  MUX41X1_HVT U107 ( .A1(n395), .A3(n328), .A2(n105), .A4(n355), .S0(n307), 
        .S1(n251), .Y(n106) );
  MUX41X1_HVT U110 ( .A1(n108), .A3(n106), .A2(n107), .A4(n104), .S0(in[5]), 
        .S1(n320), .Y(n109) );
  AO21X1_HVT U112 ( .A1(n380), .A2(n313), .A3(n26), .Y(n111) );
  NAND2X0_HVT U114 ( .A1(n334), .A2(n8), .Y(n113) );
  MUX41X1_HVT U115 ( .A1(n113), .A3(n13), .A2(n380), .A4(n328), .S0(n252), 
        .S1(n308), .Y(n114) );
  MUX41X1_HVT U116 ( .A1(n379), .A3(n373), .A2(n349), .A4(n17), .S0(n306), 
        .S1(n252), .Y(n115) );
  NAND2X0_HVT U118 ( .A1(n341), .A2(n226), .Y(n117) );
  MUX41X1_HVT U119 ( .A1(n397), .A3(n116), .A2(n39), .A4(n117), .S0(n306), 
        .S1(n344), .Y(n118) );
  MUX41X1_HVT U120 ( .A1(n118), .A3(n114), .A2(n115), .A4(n112), .S0(n323), 
        .S1(n321), .Y(n119) );
  MUX41X1_HVT U122 ( .A1(n384), .A3(n299), .A2(n48), .A4(n388), .S0(n306), 
        .S1(n343), .Y(n120) );
  MUX41X1_HVT U124 ( .A1(n301), .A3(n121), .A2(n25), .A4(n288), .S0(n312), 
        .S1(n306), .Y(n122) );
  AOI21X1_HVT U127 ( .A1(n311), .A2(n126), .A3(n356), .Y(n125) );
  NAND2X0_HVT U129 ( .A1(n310), .A2(n333), .Y(n128) );
  MUX41X1_HVT U130 ( .A1(n128), .A3(n127), .A2(n124), .A4(n125), .S0(n314), 
        .S1(n233), .Y(n129) );
  AND2X1_HVT U131 ( .A1(n283), .A2(n255), .Y(n130) );
  MUX41X1_HVT U132 ( .A1(n353), .A3(n130), .A2(n399), .A4(n362), .S0(n313), 
        .S1(n305), .Y(n131) );
  MUX41X1_HVT U133 ( .A1(n400), .A3(n355), .A2(n56), .A4(n354), .S0(n312), 
        .S1(n308), .Y(n132) );
  MUX41X1_HVT U136 ( .A1(n51), .A3(n100), .A2(n134), .A4(n360), .S0(n310), 
        .S1(n251), .Y(n135) );
  MUX41X1_HVT U137 ( .A1(n9), .A3(n31), .A2(n250), .A4(n393), .S0(n314), .S1(
        n310), .Y(n136) );
  MUX41X1_HVT U139 ( .A1(n137), .A3(n133), .A2(n129), .A4(n123), .S0(n323), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n376), .A3(n300), .A2(n370), .A4(n13), .S0(n313), 
        .S1(n309), .Y(n138) );
  NAND2X0_HVT U141 ( .A1(n325), .A2(n341), .Y(n139) );
  MUX41X1_HVT U142 ( .A1(n139), .A3(n41), .A2(n398), .A4(n370), .S0(n311), 
        .S1(n277), .Y(n140) );
  MUX41X1_HVT U143 ( .A1(n200), .A3(n381), .A2(n22), .A4(n25), .S0(n309), .S1(
        n344), .Y(n141) );
  MUX41X1_HVT U145 ( .A1(n33), .A3(n396), .A2(n142), .A4(n82), .S0(n311), .S1(
        n343), .Y(n143) );
  MUX41X1_HVT U146 ( .A1(n143), .A3(n141), .A2(n140), .A4(n138), .S0(n320), 
        .S1(n323), .Y(n144) );
  AO21X1_HVT U148 ( .A1(n314), .A2(n357), .A3(n401), .Y(n146) );
  MUX41X1_HVT U151 ( .A1(n235), .A3(n378), .A2(n253), .A4(n148), .S0(n312), 
        .S1(n305), .Y(n149) );
  MUX41X1_HVT U155 ( .A1(n370), .A3(n13), .A2(n21), .A4(n371), .S0(n309), .S1(
        n251), .Y(n153) );
  NAND2X0_HVT U159 ( .A1(n157), .A2(n158), .Y(n156) );
  MUX41X1_HVT U162 ( .A1(n293), .A3(n367), .A2(n37), .A4(n160), .S0(n309), 
        .S1(n251), .Y(n161) );
  NAND2X0_HVT U163 ( .A1(n276), .A2(n199), .Y(n162) );
  NAND2X0_HVT U166 ( .A1(n12), .A2(n166), .Y(n165) );
  MUX41X1_HVT U168 ( .A1(n167), .A3(n161), .A2(n163), .A4(n159), .S0(in[5]), 
        .S1(n320), .Y(n168) );
  MUX41X1_HVT U170 ( .A1(n303), .A3(n298), .A2(n301), .A4(n169), .S0(n309), 
        .S1(n345), .Y(n170) );
  MUX41X1_HVT U173 ( .A1(n334), .A3(n286), .A2(n330), .A4(n38), .S0(n309), 
        .S1(n345), .Y(n173) );
  MUX41X1_HVT U174 ( .A1(n392), .A3(n56), .A2(n400), .A4(n292), .S0(n309), 
        .S1(n343), .Y(n174) );
  NAND2X0_HVT U177 ( .A1(n337), .A2(n226), .Y(n176) );
  AND2X1_HVT U179 ( .A1(n237), .A2(n223), .Y(n178) );
  MUX41X1_HVT U180 ( .A1(n34), .A3(n347), .A2(n178), .A4(n47), .S0(n309), .S1(
        n345), .Y(n179) );
  MUX41X1_HVT U182 ( .A1(n355), .A3(n4), .A2(n352), .A4(n390), .S0(n306), .S1(
        n345), .Y(n181) );
  MUX41X1_HVT U183 ( .A1(n381), .A3(n385), .A2(n368), .A4(n44), .S0(n312), 
        .S1(n305), .Y(n182) );
  AND2X1_HVT U185 ( .A1(n239), .A2(n341), .Y(n184) );
  NAND2X0_HVT U191 ( .A1(n273), .A2(n361), .Y(n190) );
  AND2X1_HVT U192 ( .A1(n377), .A2(n192), .Y(n191) );
  NAND2X0_HVT U194 ( .A1(n44), .A2(n192), .Y(n194) );
  MUX41X1_HVT U195 ( .A1(n193), .A3(n194), .A2(n191), .A4(n190), .S0(n307), 
        .S1(n320), .Y(n195) );
  NAND2X0_HVT U198 ( .A1(n276), .A2(n292), .Y(n12) );
  NAND2X0_HVT U200 ( .A1(n222), .A2(n341), .Y(n126) );
  NAND2X0_HVT U207 ( .A1(n255), .A2(n286), .Y(n62) );
  INVX2_HVT U2 ( .A(n297), .Y(n261) );
  MUX21X2_HVT U3 ( .A1(n234), .A2(n403), .S0(n238), .Y(n171) );
  MUX21X1_HVT U4 ( .A1(n4), .A2(n294), .S0(n227), .Y(n65) );
  MUX21X1_HVT U6 ( .A1(n368), .A2(n65), .S0(n304), .Y(n66) );
  IBUFFX2_HVT U14 ( .A(n310), .Y(n227) );
  MUX21X1_HVT U16 ( .A1(n316), .A2(n404), .S0(n276), .Y(n45) );
  INVX2_HVT U17 ( .A(n340), .Y(n276) );
  NAND2X0_HVT U18 ( .A1(n236), .A2(n316), .Y(n196) );
  INVX1_HVT U20 ( .A(n402), .Y(n197) );
  INVX0_HVT U21 ( .A(n402), .Y(n198) );
  INVX1_HVT U22 ( .A(n197), .Y(n199) );
  INVX1_HVT U23 ( .A(n198), .Y(n200) );
  INVX0_HVT U24 ( .A(n196), .Y(n201) );
  INVX0_HVT U26 ( .A(n196), .Y(n202) );
  INVX1_HVT U27 ( .A(n201), .Y(n218) );
  INVX1_HVT U28 ( .A(n202), .Y(n219) );
  IBUFFX2_HVT U29 ( .A(n6), .Y(n220) );
  IBUFFX2_HVT U30 ( .A(n6), .Y(n221) );
  INVX1_HVT U31 ( .A(n220), .Y(n222) );
  INVX1_HVT U33 ( .A(n221), .Y(n223) );
  MUX21X1_HVT U34 ( .A1(n240), .A2(n403), .S0(n336), .Y(n33) );
  INVX1_HVT U36 ( .A(n340), .Y(n336) );
  INVX1_HVT U37 ( .A(n327), .Y(n402) );
  INVX1_HVT U39 ( .A(n335), .Y(n297) );
  MUX21X2_HVT U40 ( .A1(n369), .A2(n58), .S0(n304), .Y(n59) );
  MUX21X2_HVT U41 ( .A1(n388), .A2(n45), .S0(n224), .Y(n155) );
  IBUFFX16_HVT U43 ( .A(n313), .Y(n224) );
  INVX1_HVT U44 ( .A(n340), .Y(n337) );
  INVX1_HVT U45 ( .A(in[0]), .Y(n340) );
  IBUFFX2_HVT U46 ( .A(n45), .Y(n381) );
  NBUFFX4_HVT U47 ( .A(n290), .Y(n316) );
  INVX1_HVT U48 ( .A(n203), .Y(n385) );
  MUX21X1_HVT U49 ( .A1(n326), .A2(n229), .S0(n336), .Y(n27) );
  AO21X1_HVT U50 ( .A1(n401), .A2(n336), .A3(n273), .Y(n192) );
  MUX41X1_HVT U51 ( .A1(n188), .A3(n185), .A2(n187), .A4(n186), .S0(n225), 
        .S1(n257), .Y(n189) );
  IBUFFX16_HVT U52 ( .A(n256), .Y(n225) );
  INVX0_HVT U54 ( .A(n290), .Y(n291) );
  MUX21X1_HVT U56 ( .A1(n330), .A2(n326), .S0(n297), .Y(n294) );
  IBUFFX2_HVT U57 ( .A(n275), .Y(n238) );
  MUX21X2_HVT U58 ( .A1(n175), .A2(n168), .S0(n269), .Y(out[6]) );
  INVX1_HVT U59 ( .A(n315), .Y(n226) );
  NBUFFX2_HVT U60 ( .A(n259), .Y(n315) );
  NBUFFX4_HVT U61 ( .A(n18), .Y(n326) );
  INVX0_HVT U63 ( .A(n230), .Y(n38) );
  INVX0_HVT U64 ( .A(n294), .Y(n24) );
  MUX41X1_HVT U65 ( .A1(n174), .A3(n173), .A2(n172), .A4(n170), .S0(n228), 
        .S1(n232), .Y(n175) );
  IBUFFX16_HVT U69 ( .A(n241), .Y(n228) );
  INVX1_HVT U70 ( .A(n236), .Y(n229) );
  INVX1_HVT U75 ( .A(n318), .Y(n236) );
  MUX21X1_HVT U76 ( .A1(n324), .A2(n285), .S0(n231), .Y(n230) );
  IBUFFX16_HVT U77 ( .A(n335), .Y(n231) );
  IBUFFX2_HVT U86 ( .A(n18), .Y(n292) );
  XNOR2X2_HVT U91 ( .A1(n286), .A2(n339), .Y(n39) );
  IBUFFX16_HVT U92 ( .A(n322), .Y(n232) );
  MUX41X1_HVT U93 ( .A1(n24), .A3(n298), .A2(n171), .A4(n89), .S0(n295), .S1(
        n248), .Y(n172) );
  INVX1_HVT U94 ( .A(n309), .Y(n295) );
  IBUFFX2_HVT U97 ( .A(n346), .Y(n343) );
  IBUFFX4_HVT U103 ( .A(n343), .Y(n248) );
  INVX1_HVT U106 ( .A(n333), .Y(n403) );
  INVX1_HVT U108 ( .A(n319), .Y(n233) );
  INVX0_HVT U109 ( .A(n324), .Y(n239) );
  INVX0_HVT U111 ( .A(n326), .Y(n405) );
  NBUFFX2_HVT U113 ( .A(n264), .Y(n234) );
  NBUFFX2_HVT U117 ( .A(n390), .Y(n235) );
  NBUFFX2_HVT U121 ( .A(n264), .Y(n317) );
  INVX1_HVT U123 ( .A(n354), .Y(n237) );
  INVX0_HVT U125 ( .A(n7), .Y(n354) );
  NAND2X0_HVT U126 ( .A1(n335), .A2(n334), .Y(n7) );
  AO21X1_HVT U128 ( .A1(n341), .A2(n333), .A3(n289), .Y(n158) );
  INVX1_HVT U134 ( .A(n239), .Y(n240) );
  MUX41X1_HVT U135 ( .A1(n162), .A3(n10), .A2(n368), .A4(n39), .S0(n295), .S1(
        n345), .Y(n163) );
  MUX21X2_HVT U138 ( .A1(n302), .A2(n27), .S0(n289), .Y(n150) );
  IBUFFX16_HVT U144 ( .A(n320), .Y(n241) );
  INVX0_HVT U147 ( .A(n258), .Y(n242) );
  INVX0_HVT U149 ( .A(n290), .Y(n258) );
  NAND2X0_HVT U150 ( .A1(n86), .A2(n243), .Y(n244) );
  NAND2X0_HVT U152 ( .A1(n79), .A2(in[7]), .Y(n245) );
  NAND2X0_HVT U153 ( .A1(n244), .A2(n245), .Y(out[1]) );
  IBUFFX2_HVT U154 ( .A(in[7]), .Y(n243) );
  INVX1_HVT U156 ( .A(n27), .Y(n249) );
  INVX0_HVT U157 ( .A(n27), .Y(n370) );
  MUX21X2_HVT U158 ( .A1(n301), .A2(n382), .S0(n246), .Y(n193) );
  IBUFFX16_HVT U160 ( .A(n312), .Y(n246) );
  INVX1_HVT U161 ( .A(in[3]), .Y(n290) );
  AO21X2_HVT U164 ( .A1(n62), .A2(n312), .A3(n23), .Y(n61) );
  MUX21X2_HVT U165 ( .A1(n43), .A2(n387), .S0(n247), .Y(n187) );
  IBUFFX16_HVT U167 ( .A(n313), .Y(n247) );
  INVX0_HVT U169 ( .A(n44), .Y(n355) );
  INVX1_HVT U171 ( .A(in[6]), .Y(n264) );
  INVX0_HVT U172 ( .A(n264), .Y(n283) );
  IBUFFX2_HVT U175 ( .A(n321), .Y(n256) );
  MUX21X1_HVT U176 ( .A1(n93), .A2(n92), .S0(n310), .Y(n94) );
  MUX41X1_HVT U178 ( .A1(n66), .A3(n69), .A2(n67), .A4(n70), .S0(n322), .S1(
        n319), .Y(n71) );
  INVX2_HVT U181 ( .A(n322), .Y(n323) );
  MUX41X1_HVT U184 ( .A1(n284), .A3(n330), .A2(n368), .A4(n240), .S0(n308), 
        .S1(n248), .Y(n107) );
  INVX1_HVT U186 ( .A(n249), .Y(n250) );
  INVX1_HVT U187 ( .A(n346), .Y(n251) );
  INVX1_HVT U188 ( .A(n346), .Y(n252) );
  INVX0_HVT U189 ( .A(n24), .Y(n253) );
  MUX41X1_HVT U190 ( .A1(n349), .A3(n394), .A2(n383), .A4(n391), .S0(n254), 
        .S1(n345), .Y(n108) );
  IBUFFX16_HVT U193 ( .A(n307), .Y(n254) );
  IBUFFX2_HVT U196 ( .A(in[0]), .Y(n255) );
  INVX0_HVT U197 ( .A(n177), .Y(n278) );
  IBUFFX16_HVT U199 ( .A(n305), .Y(n257) );
  IBUFFX2_HVT U201 ( .A(in[0]), .Y(n341) );
  INVX1_HVT U202 ( .A(n258), .Y(n259) );
  MUX21X1_HVT U203 ( .A1(n91), .A2(n3), .S0(n261), .Y(n92) );
  MUX21X2_HVT U204 ( .A1(n154), .A2(n144), .S0(in[7]), .Y(out[5]) );
  NAND2X0_HVT U205 ( .A1(n335), .A2(n331), .Y(n4) );
  MUX21X1_HVT U206 ( .A1(n53), .A2(n54), .S0(n310), .Y(n55) );
  INVX1_HVT U208 ( .A(n346), .Y(n345) );
  INVX1_HVT U209 ( .A(n23), .Y(n368) );
  NAND2X0_HVT U210 ( .A1(n156), .A2(n295), .Y(n265) );
  OA21X1_HVT U211 ( .A1(n350), .A2(n273), .A3(n359), .Y(n151) );
  INVX1_HVT U212 ( .A(n319), .Y(n320) );
  INVX1_HVT U213 ( .A(in[1]), .Y(n319) );
  INVX0_HVT U214 ( .A(in[7]), .Y(n287) );
  INVX1_HVT U215 ( .A(n313), .Y(n289) );
  INVX1_HVT U216 ( .A(n314), .Y(n273) );
  MUX21X2_HVT U217 ( .A1(n102), .A2(n95), .S0(in[7]), .Y(out[2]) );
  IBUFFX2_HVT U218 ( .A(n346), .Y(n344) );
  OA21X1_HVT U219 ( .A1(n351), .A2(n273), .A3(n23), .Y(n77) );
  MUX21X1_HVT U220 ( .A1(n324), .A2(n316), .S0(n337), .Y(n23) );
  INVX0_HVT U221 ( .A(n340), .Y(n335) );
  INVX1_HVT U222 ( .A(n297), .Y(n260) );
  MUX21X2_HVT U223 ( .A1(n302), .A2(n50), .S0(n314), .Y(n186) );
  XOR2X2_HVT U224 ( .A1(n218), .A2(n260), .Y(n50) );
  NAND2X0_HVT U225 ( .A1(n109), .A2(n269), .Y(n262) );
  NAND2X0_HVT U226 ( .A1(n119), .A2(n287), .Y(n263) );
  NAND2X0_HVT U227 ( .A1(n262), .A2(n263), .Y(out[3]) );
  MUX21X2_HVT U228 ( .A1(n356), .A2(n43), .S0(n314), .Y(n110) );
  MUX21X1_HVT U229 ( .A1(n283), .A2(n404), .S0(n335), .Y(n43) );
  MUX21X1_HVT U230 ( .A1(n184), .A2(n389), .S0(n312), .Y(n185) );
  OR2X1_HVT U231 ( .A1(n259), .A2(n264), .Y(n3) );
  INVX1_HVT U232 ( .A(n328), .Y(n404) );
  MUX21X2_HVT U233 ( .A1(n145), .A2(n146), .S0(n310), .Y(n147) );
  MUX21X2_HVT U234 ( .A1(n399), .A2(n353), .S0(n312), .Y(n145) );
  NAND2X0_HVT U235 ( .A1(n155), .A2(n311), .Y(n266) );
  NAND2X0_HVT U236 ( .A1(n265), .A2(n266), .Y(n159) );
  NAND2X0_HVT U237 ( .A1(n61), .A2(n311), .Y(n267) );
  NAND2X0_HVT U238 ( .A1(n60), .A2(n295), .Y(n268) );
  NAND2X0_HVT U239 ( .A1(n267), .A2(n268), .Y(n63) );
  NAND2X0_HVT U240 ( .A1(n64), .A2(n269), .Y(n270) );
  NAND2X0_HVT U241 ( .A1(n71), .A2(n287), .Y(n271) );
  NAND2X0_HVT U242 ( .A1(n270), .A2(n271), .Y(out[0]) );
  IBUFFX2_HVT U243 ( .A(n287), .Y(n269) );
  MUX21X1_HVT U244 ( .A1(n288), .A2(n56), .S0(n313), .Y(n60) );
  INVX1_HVT U245 ( .A(n272), .Y(n53) );
  MUX21X1_HVT U246 ( .A1(n17), .A2(n29), .S0(n273), .Y(n272) );
  IBUFFX2_HVT U247 ( .A(n17), .Y(n363) );
  IBUFFX2_HVT U248 ( .A(n29), .Y(n371) );
  IBUFFX2_HVT U249 ( .A(n340), .Y(n339) );
  INVX1_HVT U250 ( .A(n293), .Y(n46) );
  OA21X1_HVT U251 ( .A1(n373), .A2(n273), .A3(n62), .Y(n188) );
  INVX0_HVT U252 ( .A(n284), .Y(n28) );
  AO21X1_HVT U253 ( .A1(n325), .A2(n4), .A3(n289), .Y(n166) );
  INVX0_HVT U254 ( .A(n288), .Y(n25) );
  INVX0_HVT U255 ( .A(n317), .Y(n285) );
  INVX0_HVT U256 ( .A(n319), .Y(n321) );
  NBUFFX2_HVT U257 ( .A(in[4]), .Y(n274) );
  IBUFFX2_HVT U258 ( .A(n340), .Y(n275) );
  IBUFFX4_HVT U259 ( .A(n346), .Y(n277) );
  OR2X1_HVT U260 ( .A1(n278), .A2(n319), .Y(n282) );
  INVX1_HVT U261 ( .A(n207), .Y(n389) );
  INVX1_HVT U262 ( .A(n206), .Y(n388) );
  INVX0_HVT U263 ( .A(in[4]), .Y(n346) );
  INVX1_HVT U264 ( .A(n296), .Y(n169) );
  MUX41X1_HVT U265 ( .A1(n40), .A3(n366), .A2(n367), .A4(n365), .S0(n295), 
        .S1(n273), .Y(n67) );
  NAND2X0_HVT U266 ( .A1(n182), .A2(n319), .Y(n279) );
  NAND2X0_HVT U267 ( .A1(n181), .A2(n233), .Y(n280) );
  NAND2X0_HVT U268 ( .A1(n279), .A2(n280), .Y(n183) );
  NAND2X0_HVT U269 ( .A1(n179), .A2(n319), .Y(n281) );
  NAND2X0_HVT U270 ( .A1(n281), .A2(n282), .Y(n180) );
  MUX41X1_HVT U271 ( .A1(n56), .A3(n284), .A2(n240), .A4(n385), .S0(n295), 
        .S1(n289), .Y(n57) );
  MUX41X1_HVT U272 ( .A1(n180), .A3(n183), .A2(n189), .A4(n195), .S0(n322), 
        .S1(n287), .Y(out[7]) );
  MUX41X1_HVT U273 ( .A1(n152), .A3(n147), .A2(n153), .A4(n149), .S0(n323), 
        .S1(n319), .Y(n154) );
  MUX21X1_HVT U274 ( .A1(n330), .A2(n285), .S0(n341), .Y(n284) );
  XOR2X2_HVT U275 ( .A1(n234), .A2(n291), .Y(n18) );
  IBUFFX2_HVT U276 ( .A(n1), .Y(n286) );
  INVX1_HVT U277 ( .A(n205), .Y(n387) );
  IBUFFX2_HVT U278 ( .A(n33), .Y(n375) );
  NBUFFX2_HVT U279 ( .A(n264), .Y(n318) );
  MUX21X1_HVT U280 ( .A1(n259), .A2(n330), .S0(n255), .Y(n288) );
  INVX1_HVT U281 ( .A(n330), .Y(n401) );
  IBUFFX2_HVT U282 ( .A(n340), .Y(n338) );
  MUX21X2_HVT U283 ( .A1(n151), .A2(n150), .S0(n311), .Y(n152) );
  MUX21X1_HVT U284 ( .A1(n334), .A2(n223), .S0(n341), .Y(n293) );
  INVX1_HVT U285 ( .A(n208), .Y(n390) );
  MUX41X1_HVT U286 ( .A1(n46), .A3(n286), .A2(n176), .A4(n303), .S0(n295), 
        .S1(n289), .Y(n177) );
  MUX21X1_HVT U287 ( .A1(n328), .A2(n333), .S0(n297), .Y(n296) );
  INVX0_HVT U288 ( .A(in[5]), .Y(n322) );
  NBUFFX2_HVT U289 ( .A(n2), .Y(n330) );
  NBUFFX2_HVT U290 ( .A(n2), .Y(n332) );
  NBUFFX2_HVT U291 ( .A(n2), .Y(n331) );
  AND2X1_HVT U292 ( .A1(n7), .A2(n331), .Y(n298) );
  AND2X1_HVT U293 ( .A1(n331), .A2(n17), .Y(n299) );
  MUX21X1_HVT U294 ( .A1(n219), .A2(n329), .S0(n261), .Y(n160) );
  MUX21X1_HVT U295 ( .A1(n315), .A2(n405), .S0(n339), .Y(n208) );
  MUX21X1_HVT U296 ( .A1(n286), .A2(n325), .S0(n275), .Y(n210) );
  MUX21X1_HVT U297 ( .A1(n403), .A2(n199), .S0(n337), .Y(n30) );
  MUX21X1_HVT U298 ( .A1(n292), .A2(n316), .S0(n276), .Y(n41) );
  MUX21X1_HVT U299 ( .A1(n401), .A2(n292), .S0(n261), .Y(n35) );
  MUX21X1_HVT U300 ( .A1(n234), .A2(n199), .S0(n339), .Y(n148) );
  NAND2X0_HVT U301 ( .A1(n259), .A2(n317), .Y(n2) );
  MUX21X1_HVT U302 ( .A1(n401), .A2(n318), .S0(n338), .Y(n205) );
  MUX21X1_HVT U303 ( .A1(n292), .A2(n234), .S0(n338), .Y(n215) );
  MUX21X1_HVT U304 ( .A1(n404), .A2(n316), .S0(n336), .Y(n206) );
  MUX21X1_HVT U305 ( .A1(n325), .A2(n200), .S0(n339), .Y(n36) );
  MUX21X1_HVT U306 ( .A1(n223), .A2(n332), .S0(n336), .Y(n216) );
  MUX21X1_HVT U307 ( .A1(n316), .A2(n331), .S0(n260), .Y(n207) );
  XNOR2X1_HVT U308 ( .A1(n330), .A2(n339), .Y(n300) );
  MUX21X1_HVT U309 ( .A1(n333), .A2(n332), .S0(n276), .Y(n16) );
  MUX21X1_HVT U310 ( .A1(n316), .A2(n401), .S0(n337), .Y(n32) );
  MUX21X1_HVT U311 ( .A1(n234), .A2(n332), .S0(n275), .Y(n105) );
  MUX21X1_HVT U312 ( .A1(n229), .A2(n325), .S0(n275), .Y(n42) );
  MUX21X1_HVT U313 ( .A1(n329), .A2(n331), .S0(n276), .Y(n20) );
  MUX21X1_HVT U314 ( .A1(n3), .A2(n316), .S0(n261), .Y(n21) );
  MUX21X1_HVT U315 ( .A1(n316), .A2(n234), .S0(n337), .Y(n47) );
  MUX21X1_HVT U316 ( .A1(n35), .A2(n299), .S0(n311), .Y(n127) );
  MUX21X1_HVT U317 ( .A1(n398), .A2(n300), .S0(n310), .Y(n124) );
  MUX21X1_HVT U318 ( .A1(n358), .A2(n325), .S0(n314), .Y(n93) );
  MUX21X1_HVT U319 ( .A1(n324), .A2(n318), .S0(n313), .Y(n91) );
  XOR2X1_HVT U320 ( .A1(n325), .A2(n338), .Y(n48) );
  XOR2X1_HVT U321 ( .A1(n328), .A2(n338), .Y(n49) );
  AND2X1_HVT U322 ( .A1(n338), .A2(n318), .Y(n301) );
  MUX21X1_HVT U323 ( .A1(n242), .A2(n3), .S0(n337), .Y(n213) );
  MUX21X1_HVT U324 ( .A1(n329), .A2(n318), .S0(n339), .Y(n121) );
  NBUFFX2_HVT U325 ( .A(n274), .Y(n314) );
  NBUFFX2_HVT U326 ( .A(n274), .Y(n313) );
  NBUFFX2_HVT U327 ( .A(n274), .Y(n312) );
  NBUFFX2_HVT U328 ( .A(n1), .Y(n333) );
  NBUFFX2_HVT U329 ( .A(n18), .Y(n324) );
  MUX21X1_HVT U330 ( .A1(n165), .A2(n164), .S0(n310), .Y(n167) );
  MUX21X1_HVT U331 ( .A1(n28), .A2(n25), .S0(n312), .Y(n164) );
  MUX21X1_HVT U332 ( .A1(n330), .A2(n219), .S0(n275), .Y(n142) );
  MUX21X1_HVT U333 ( .A1(n401), .A2(n404), .S0(n338), .Y(n52) );
  NBUFFX2_HVT U334 ( .A(n18), .Y(n325) );
  MUX21X1_HVT U335 ( .A1(n370), .A2(n5), .S0(n311), .Y(n58) );
  MUX21X1_HVT U336 ( .A1(n111), .A2(n110), .S0(n311), .Y(n112) );
  NBUFFX2_HVT U337 ( .A(n1), .Y(n334) );
  NBUFFX2_HVT U338 ( .A(n6), .Y(n327) );
  AND2X1_HVT U339 ( .A1(n329), .A2(n255), .Y(n302) );
  AND2X1_HVT U340 ( .A1(n404), .A2(n255), .Y(n303) );
  NBUFFX2_HVT U341 ( .A(n3), .Y(n328) );
  NBUFFX2_HVT U342 ( .A(n3), .Y(n329) );
  MUX21X1_HVT U343 ( .A1(n122), .A2(n120), .S0(n233), .Y(n123) );
  MUX21X1_HVT U344 ( .A1(n76), .A2(n77), .S0(n311), .Y(n78) );
  MUX21X1_HVT U345 ( .A1(n388), .A2(n348), .S0(n314), .Y(n76) );
  NBUFFX2_HVT U346 ( .A(in[2]), .Y(n309) );
  NBUFFX2_HVT U347 ( .A(n342), .Y(n310) );
  XNOR2X1_HVT U348 ( .A1(n289), .A2(n306), .Y(n304) );
  NBUFFX2_HVT U349 ( .A(n342), .Y(n311) );
  NBUFFX2_HVT U350 ( .A(n342), .Y(n306) );
  NBUFFX2_HVT U351 ( .A(n342), .Y(n308) );
  NBUFFX2_HVT U352 ( .A(n342), .Y(n307) );
  NBUFFX2_HVT U353 ( .A(n342), .Y(n305) );
  MUX21X1_HVT U354 ( .A1(n286), .A2(n226), .S0(n336), .Y(n217) );
  MUX21X1_HVT U355 ( .A1(n219), .A2(n226), .S0(n338), .Y(n97) );
  MUX21X1_HVT U356 ( .A1(n334), .A2(n226), .S0(n339), .Y(n157) );
  MUX21X1_HVT U357 ( .A1(n132), .A2(n131), .S0(n233), .Y(n133) );
  MUX21X1_HVT U358 ( .A1(n136), .A2(n135), .S0(n233), .Y(n137) );
  MUX21X1_HVT U359 ( .A1(n229), .A2(n226), .S0(n261), .Y(n29) );
  MUX21X1_HVT U360 ( .A1(n404), .A2(n199), .S0(n336), .Y(n116) );
  MUX21X1_HVT U361 ( .A1(n226), .A2(n334), .S0(n339), .Y(n211) );
  MUX21X1_HVT U362 ( .A1(n226), .A2(n218), .S0(n338), .Y(n212) );
  NBUFFX2_HVT U363 ( .A(in[2]), .Y(n342) );
  MUX21X1_HVT U364 ( .A1(n401), .A2(n283), .S0(n276), .Y(n134) );
  XOR2X1_HVT U365 ( .A1(n276), .A2(n283), .Y(n51) );
  MUX21X1_HVT U366 ( .A1(n3), .A2(n283), .S0(n336), .Y(n209) );
  MUX21X1_HVT U367 ( .A1(n283), .A2(n403), .S0(n337), .Y(n26) );
  MUX21X1_HVT U368 ( .A1(n283), .A2(n333), .S0(n260), .Y(n19) );
  MUX21X1_HVT U369 ( .A1(n283), .A2(n329), .S0(n275), .Y(n204) );
  MUX21X1_HVT U370 ( .A1(n315), .A2(n283), .S0(n261), .Y(n214) );
  MUX21X1_HVT U371 ( .A1(n222), .A2(n283), .S0(n275), .Y(n31) );
  MUX21X1_HVT U372 ( .A1(n283), .A2(n200), .S0(n337), .Y(n203) );
  INVX0_HVT U373 ( .A(n13), .Y(n347) );
  INVX0_HVT U374 ( .A(n34), .Y(n348) );
  INVX0_HVT U375 ( .A(n40), .Y(n349) );
  INVX0_HVT U376 ( .A(n100), .Y(n350) );
  INVX0_HVT U377 ( .A(n139), .Y(n351) );
  INVX0_HVT U378 ( .A(n4), .Y(n352) );
  INVX0_HVT U379 ( .A(n5), .Y(n353) );
  INVX0_HVT U380 ( .A(n8), .Y(n356) );
  INVX0_HVT U381 ( .A(n9), .Y(n357) );
  INVX0_HVT U382 ( .A(n37), .Y(n358) );
  INVX0_HVT U383 ( .A(n15), .Y(n359) );
  INVX0_HVT U384 ( .A(n10), .Y(n360) );
  INVX0_HVT U385 ( .A(n14), .Y(n361) );
  INVX0_HVT U386 ( .A(n16), .Y(n362) );
  INVX0_HVT U387 ( .A(n19), .Y(n364) );
  INVX0_HVT U388 ( .A(n20), .Y(n365) );
  INVX0_HVT U389 ( .A(n21), .Y(n366) );
  INVX0_HVT U390 ( .A(n22), .Y(n367) );
  INVX0_HVT U391 ( .A(n26), .Y(n369) );
  INVX0_HVT U392 ( .A(n30), .Y(n372) );
  INVX0_HVT U393 ( .A(n31), .Y(n373) );
  INVX0_HVT U394 ( .A(n32), .Y(n374) );
  INVX0_HVT U395 ( .A(n35), .Y(n376) );
  INVX0_HVT U396 ( .A(n36), .Y(n377) );
  INVX0_HVT U397 ( .A(n39), .Y(n378) );
  INVX0_HVT U398 ( .A(n41), .Y(n379) );
  INVX0_HVT U399 ( .A(n42), .Y(n380) );
  INVX0_HVT U400 ( .A(n47), .Y(n382) );
  INVX0_HVT U401 ( .A(n48), .Y(n383) );
  INVX0_HVT U402 ( .A(n11), .Y(n384) );
  INVX0_HVT U403 ( .A(n204), .Y(n386) );
  INVX0_HVT U404 ( .A(n209), .Y(n391) );
  INVX0_HVT U405 ( .A(n210), .Y(n392) );
  INVX0_HVT U406 ( .A(n211), .Y(n393) );
  INVX0_HVT U407 ( .A(n212), .Y(n394) );
  INVX0_HVT U408 ( .A(n213), .Y(n395) );
  INVX0_HVT U409 ( .A(n214), .Y(n396) );
  INVX0_HVT U410 ( .A(n157), .Y(n397) );
  INVX0_HVT U411 ( .A(n215), .Y(n398) );
  INVX0_HVT U412 ( .A(n216), .Y(n399) );
  INVX0_HVT U413 ( .A(n217), .Y(n400) );
endmodule

