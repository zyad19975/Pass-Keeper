
module inv_sbox_4 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n196, n197, n198, n199, n200, n201, n202, n205, n208, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630;

  NAND2X0_HVT U1 ( .A1(n228), .A2(n337), .Y(n630) );
  NAND2X0_HVT U5 ( .A1(n627), .A2(n270), .Y(n626) );
  NAND2X0_HVT U8 ( .A1(n297), .A2(n270), .Y(n622) );
  NAND2X0_HVT U9 ( .A1(n257), .A2(n622), .Y(n621) );
  NAND2X0_HVT U10 ( .A1(n256), .A2(n619), .Y(n620) );
  NAND2X0_HVT U12 ( .A1(n352), .A2(n335), .Y(n617) );
  NAND2X0_HVT U13 ( .A1(n349), .A2(n622), .Y(n616) );
  NAND2X0_HVT U15 ( .A1(n344), .A2(n353), .Y(n614) );
  NAND2X0_HVT U19 ( .A1(n298), .A2(n420), .Y(n609) );
  NAND2X0_HVT U32 ( .A1(n337), .A2(n235), .Y(n597) );
  NAND2X0_HVT U35 ( .A1(n622), .A2(n421), .Y(n594) );
  NAND2X0_HVT U38 ( .A1(n335), .A2(n235), .Y(n591) );
  NAND2X0_HVT U42 ( .A1(n624), .A2(n421), .Y(n587) );
  OA21X1_HVT U53 ( .A1(n240), .A2(n579), .A3(n280), .Y(n577) );
  AO21X1_HVT U60 ( .A1(n569), .A2(n331), .A3(n608), .Y(n570) );
  NAND2X0_HVT U66 ( .A1(n352), .A2(n324), .Y(n563) );
  MUX41X1_HVT U67 ( .A1(n380), .A3(n404), .A2(n382), .A4(n563), .S0(n333), 
        .S1(n327), .Y(n562) );
  MUX41X1_HVT U71 ( .A1(n624), .A3(n254), .A2(n618), .A4(n376), .S0(n329), 
        .S1(n304), .Y(n559) );
  NAND2X0_HVT U72 ( .A1(n345), .A2(n623), .Y(n558) );
  MUX41X1_HVT U73 ( .A1(n602), .A3(n558), .A2(n231), .A4(n334), .S0(n332), 
        .S1(n326), .Y(n557) );
  MUX41X1_HVT U74 ( .A1(n620), .A3(n396), .A2(n395), .A4(n386), .S0(n330), 
        .S1(n304), .Y(n556) );
  MUX41X1_HVT U78 ( .A1(n553), .A3(n557), .A2(n556), .A4(n559), .S0(in[5]), 
        .S1(in[1]), .Y(n552) );
  MUX41X1_HVT U79 ( .A1(n392), .A3(n611), .A2(n394), .A4(n612), .S0(n330), 
        .S1(n363), .Y(n551) );
  MUX41X1_HVT U80 ( .A1(n406), .A3(n244), .A2(n621), .A4(n626), .S0(n329), 
        .S1(n361), .Y(n550) );
  NAND2X0_HVT U81 ( .A1(n315), .A2(n623), .Y(n549) );
  AND2X1_HVT U82 ( .A1(n624), .A2(n347), .Y(n548) );
  MUX41X1_HVT U83 ( .A1(n548), .A3(n393), .A2(n309), .A4(n549), .S0(n329), 
        .S1(n303), .Y(n547) );
  MUX41X1_HVT U84 ( .A1(n321), .A3(n392), .A2(n407), .A4(n604), .S0(n330), 
        .S1(n303), .Y(n546) );
  MUX41X1_HVT U85 ( .A1(n546), .A3(n550), .A2(n547), .A4(n551), .S0(n342), 
        .S1(n339), .Y(n545) );
  MUX41X1_HVT U87 ( .A1(n370), .A3(n321), .A2(n408), .A4(n390), .S0(n328), 
        .S1(n363), .Y(n544) );
  MUX41X1_HVT U88 ( .A1(n382), .A3(n367), .A2(n599), .A4(n583), .S0(n329), 
        .S1(n262), .Y(n543) );
  NAND2X0_HVT U89 ( .A1(n236), .A2(n417), .Y(n542) );
  MUX41X1_HVT U90 ( .A1(n254), .A3(n623), .A2(n582), .A4(n542), .S0(n329), 
        .S1(n363), .Y(n541) );
  MUX41X1_HVT U95 ( .A1(n537), .A3(n543), .A2(n541), .A4(n544), .S0(n342), 
        .S1(n340), .Y(n536) );
  MUX41X1_HVT U96 ( .A1(n404), .A3(n616), .A2(n391), .A4(n409), .S0(n330), 
        .S1(n303), .Y(n535) );
  MUX41X1_HVT U98 ( .A1(n534), .A3(n410), .A2(n397), .A4(n601), .S0(n330), 
        .S1(n303), .Y(n533) );
  MUX41X1_HVT U99 ( .A1(n597), .A3(n384), .A2(n581), .A4(n343), .S0(n304), 
        .S1(n327), .Y(n532) );
  NAND2X0_HVT U100 ( .A1(n236), .A2(n313), .Y(n531) );
  MUX41X1_HVT U101 ( .A1(n411), .A3(n617), .A2(n196), .A4(n531), .S0(n265), 
        .S1(n325), .Y(n530) );
  MUX41X1_HVT U102 ( .A1(n530), .A3(n533), .A2(n532), .A4(n535), .S0(n342), 
        .S1(n339), .Y(n529) );
  AND2X1_HVT U104 ( .A1(n623), .A2(n346), .Y(n528) );
  MUX41X1_HVT U105 ( .A1(n615), .A3(n412), .A2(n549), .A4(n528), .S0(n330), 
        .S1(n265), .Y(n527) );
  MUX41X1_HVT U107 ( .A1(n411), .A3(n347), .A2(n526), .A4(n373), .S0(n329), 
        .S1(n265), .Y(n525) );
  MUX41X1_HVT U109 ( .A1(n410), .A3(n367), .A2(n407), .A4(n401), .S0(n329), 
        .S1(n261), .Y(n523) );
  AO21X1_HVT U112 ( .A1(n399), .A2(n332), .A3(n605), .Y(n520) );
  NAND2X0_HVT U114 ( .A1(n257), .A2(n623), .Y(n518) );
  MUX41X1_HVT U115 ( .A1(n518), .A3(n618), .A2(n399), .A4(n347), .S0(n361), 
        .S1(n327), .Y(n517) );
  NAND2X0_HVT U118 ( .A1(n235), .A2(n308), .Y(n514) );
  MUX41X1_HVT U119 ( .A1(n413), .A3(n515), .A2(n592), .A4(n514), .S0(n328), 
        .S1(n262), .Y(n513) );
  MUX41X1_HVT U120 ( .A1(n513), .A3(n517), .A2(n516), .A4(n519), .S0(n342), 
        .S1(n340), .Y(n512) );
  MUX41X1_HVT U122 ( .A1(n402), .A3(n318), .A2(n583), .A4(n405), .S0(n328), 
        .S1(n361), .Y(n511) );
  MUX41X1_HVT U124 ( .A1(n320), .A3(n510), .A2(n606), .A4(n387), .S0(n331), 
        .S1(n328), .Y(n509) );
  NAND2X0_HVT U129 ( .A1(n358), .A2(n256), .Y(n503) );
  MUX41X1_HVT U130 ( .A1(n503), .A3(n504), .A2(n507), .A4(n506), .S0(n333), 
        .S1(n340), .Y(n502) );
  AND2X1_HVT U131 ( .A1(n324), .A2(n263), .Y(n501) );
  MUX41X1_HVT U132 ( .A1(n371), .A3(n501), .A2(n415), .A4(n380), .S0(n332), 
        .S1(n326), .Y(n500) );
  MUX41X1_HVT U133 ( .A1(n416), .A3(n373), .A2(n575), .A4(n372), .S0(n331), 
        .S1(n325), .Y(n499) );
  MUX41X1_HVT U137 ( .A1(n622), .A3(n600), .A2(n604), .A4(n409), .S0(n333), 
        .S1(n325), .Y(n495) );
  MUX41X1_HVT U139 ( .A1(n494), .A3(n498), .A2(n502), .A4(n508), .S0(n342), 
        .S1(in[7]), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n395), .A3(n319), .A2(n389), .A4(n618), .S0(n332), 
        .S1(n327), .Y(n493) );
  NAND2X0_HVT U141 ( .A1(n344), .A2(n357), .Y(n492) );
  MUX41X1_HVT U143 ( .A1(n417), .A3(n400), .A2(n609), .A4(n606), .S0(n360), 
        .S1(n261), .Y(n490) );
  AO21X1_HVT U148 ( .A1(n333), .A2(n375), .A3(n313), .Y(n485) );
  MUX41X1_HVT U155 ( .A1(n389), .A3(n618), .A2(n610), .A4(n391), .S0(n326), 
        .S1(n261), .Y(n478) );
  MUX41X1_HVT U156 ( .A1(n478), .A3(n482), .A2(n479), .A4(n484), .S0(n342), 
        .S1(n340), .Y(n477) );
  NAND2X0_HVT U159 ( .A1(n474), .A2(n473), .Y(n475) );
  MUX41X1_HVT U162 ( .A1(n316), .A3(n385), .A2(n594), .A4(n471), .S0(n329), 
        .S1(n262), .Y(n470) );
  NAND2X0_HVT U163 ( .A1(n352), .A2(n417), .Y(n469) );
  MUX41X1_HVT U164 ( .A1(n621), .A3(n469), .A2(n592), .A4(n386), .S0(n328), 
        .S1(n361), .Y(n468) );
  NAND2X0_HVT U166 ( .A1(n619), .A2(n465), .Y(n466) );
  MUX41X1_HVT U168 ( .A1(n464), .A3(n470), .A2(n468), .A4(n472), .S0(n342), 
        .S1(n339), .Y(n463) );
  MUX41X1_HVT U170 ( .A1(n322), .A3(n317), .A2(n320), .A4(n462), .S0(n360), 
        .S1(n262), .Y(n461) );
  MUX41X1_HVT U172 ( .A1(n542), .A3(n460), .A2(n317), .A4(n607), .S0(n358), 
        .S1(n304), .Y(n459) );
  MUX41X1_HVT U174 ( .A1(n408), .A3(n575), .A2(n416), .A4(n421), .S0(n325), 
        .S1(n261), .Y(n457) );
  NAND2X0_HVT U177 ( .A1(n353), .A2(n308), .Y(n455) );
  MUX41X1_HVT U178 ( .A1(n322), .A3(n455), .A2(n253), .A4(n585), .S0(n360), 
        .S1(n361), .Y(n454) );
  AND2X1_HVT U179 ( .A1(n624), .A2(n346), .Y(n453) );
  MUX41X1_HVT U180 ( .A1(n597), .A3(n365), .A2(n453), .A4(n584), .S0(n360), 
        .S1(n303), .Y(n452) );
  AND2X1_HVT U185 ( .A1(n421), .A2(n263), .Y(n447) );
  NAND2X0_HVT U191 ( .A1(n307), .A2(n379), .Y(n441) );
  AND2X1_HVT U192 ( .A1(n396), .A2(n439), .Y(n440) );
  NAND2X0_HVT U194 ( .A1(n587), .A2(n439), .Y(n437) );
  NAND2X0_HVT U198 ( .A1(n352), .A2(n421), .Y(n619) );
  NAND2X0_HVT U200 ( .A1(n270), .A2(n357), .Y(n505) );
  NAND2X0_HVT U207 ( .A1(n236), .A2(n253), .Y(n569) );
  IBUFFX4_HVT U2 ( .A(n331), .Y(n241) );
  IBUFFX4_HVT U3 ( .A(n331), .Y(n249) );
  MUX21X2_HVT U4 ( .A1(n420), .A2(n324), .S0(n291), .Y(n588) );
  MUX21X1_HVT U6 ( .A1(n277), .A2(n343), .S0(n355), .Y(n196) );
  INVX8_HVT U7 ( .A(n196), .Y(n593) );
  INVX1_HVT U11 ( .A(n277), .Y(n278) );
  NAND2X0_HVT U14 ( .A1(n344), .A2(n197), .Y(n198) );
  NAND2X0_HVT U16 ( .A1(n337), .A2(n332), .Y(n199) );
  NAND2X0_HVT U17 ( .A1(n198), .A2(n199), .Y(n540) );
  INVX0_HVT U18 ( .A(n332), .Y(n197) );
  MUX21X2_HVT U20 ( .A1(n540), .A2(n348), .S0(n200), .Y(n539) );
  IBUFFX16_HVT U21 ( .A(n356), .Y(n200) );
  MUX21X2_HVT U22 ( .A1(n539), .A2(n538), .S0(n201), .Y(n537) );
  IBUFFX16_HVT U23 ( .A(n358), .Y(n201) );
  NAND2X0_HVT U24 ( .A1(n349), .A2(n627), .Y(n575) );
  IBUFFX2_HVT U25 ( .A(n627), .Y(n370) );
  IBUFFX2_HVT U26 ( .A(n327), .Y(n250) );
  MUX21X2_HVT U27 ( .A1(n570), .A2(n571), .S0(n250), .Y(n568) );
  MUX21X2_HVT U28 ( .A1(n466), .A2(n467), .S0(n202), .Y(n464) );
  IBUFFX16_HVT U29 ( .A(n306), .Y(n202) );
  NAND2X0_HVT U30 ( .A1(n447), .A2(n205), .Y(n208) );
  NAND2X0_HVT U31 ( .A1(n406), .A2(n331), .Y(n218) );
  NAND2X0_HVT U33 ( .A1(n208), .A2(n218), .Y(n446) );
  IBUFFX2_HVT U34 ( .A(n331), .Y(n205) );
  NBUFFX4_HVT U36 ( .A(n362), .Y(n331) );
  NBUFFX4_HVT U37 ( .A(n362), .Y(n332) );
  MUX21X1_HVT U39 ( .A1(n313), .A2(n421), .S0(n352), .Y(n596) );
  INVX0_HVT U40 ( .A(n348), .Y(n220) );
  MUX21X2_HVT U41 ( .A1(n606), .A2(n603), .S0(n307), .Y(n467) );
  MUX41X1_HVT U43 ( .A1(n525), .A3(n523), .A2(n527), .A4(n524), .S0(n219), 
        .S1(n340), .Y(n522) );
  IBUFFX16_HVT U44 ( .A(n342), .Y(n219) );
  OR2X1_HVT U45 ( .A1(n235), .A2(n220), .Y(n623) );
  INVX1_HVT U46 ( .A(n357), .Y(n298) );
  MUX21X2_HVT U47 ( .A1(n560), .A2(n567), .S0(in[7]), .Y(out[0]) );
  INVX0_HVT U48 ( .A(n235), .Y(n221) );
  MUX41X1_HVT U49 ( .A1(n445), .A3(n446), .A2(n444), .A4(n443), .S0(n326), 
        .S1(n338), .Y(n442) );
  IBUFFX2_HVT U50 ( .A(n290), .Y(n235) );
  MUX21X1_HVT U51 ( .A1(n321), .A2(n581), .S0(n333), .Y(n445) );
  MUX21X1_HVT U52 ( .A1(n231), .A2(n588), .S0(n332), .Y(n444) );
  MUX21X1_HVT U54 ( .A1(n376), .A2(n344), .S0(n333), .Y(n538) );
  MUX41X1_HVT U55 ( .A1(n380), .A3(n308), .A2(n381), .A4(n256), .S0(n329), 
        .S1(n363), .Y(n561) );
  MUX21X2_HVT U56 ( .A1(n486), .A2(n485), .S0(n325), .Y(n484) );
  MUX21X2_HVT U57 ( .A1(n415), .A2(n371), .S0(n331), .Y(n486) );
  MUX21X2_HVT U58 ( .A1(n588), .A2(n374), .S0(n222), .Y(n521) );
  IBUFFX16_HVT U59 ( .A(n333), .Y(n222) );
  MUX41X1_HVT U61 ( .A1(n565), .A3(n564), .A2(n562), .A4(n561), .S0(n338), 
        .S1(n341), .Y(n560) );
  NAND2X0_HVT U62 ( .A1(n248), .A2(n223), .Y(n224) );
  NAND2X0_HVT U63 ( .A1(n299), .A2(n232), .Y(n225) );
  NAND2X0_HVT U64 ( .A1(n224), .A2(n225), .Y(n566) );
  INVX0_HVT U65 ( .A(n232), .Y(n223) );
  INVX0_HVT U68 ( .A(n370), .Y(n248) );
  IBUFFX2_HVT U69 ( .A(n358), .Y(n232) );
  IBUFFX2_HVT U70 ( .A(n299), .Y(n607) );
  MUX21X2_HVT U75 ( .A1(n552), .A2(n545), .S0(n226), .Y(out[1]) );
  IBUFFX16_HVT U76 ( .A(in[7]), .Y(n226) );
  INVX1_HVT U77 ( .A(in[6]), .Y(n422) );
  NBUFFX2_HVT U86 ( .A(n422), .Y(n337) );
  INVX1_HVT U91 ( .A(n255), .Y(n256) );
  INVX1_HVT U92 ( .A(n630), .Y(n255) );
  INVX0_HVT U93 ( .A(n587), .Y(n373) );
  INVX0_HVT U94 ( .A(n314), .Y(n311) );
  INVX1_HVT U97 ( .A(n314), .Y(n315) );
  INVX0_HVT U103 ( .A(n629), .Y(n314) );
  INVX1_HVT U106 ( .A(n314), .Y(n310) );
  MUX21X2_HVT U108 ( .A1(n522), .A2(n512), .S0(n227), .Y(out[3]) );
  IBUFFX16_HVT U110 ( .A(in[7]), .Y(n227) );
  INVX0_HVT U111 ( .A(n271), .Y(n228) );
  INVX1_HVT U113 ( .A(n425), .Y(n414) );
  MUX21X2_HVT U116 ( .A1(n509), .A2(n511), .S0(n339), .Y(n508) );
  INVX1_HVT U117 ( .A(n338), .Y(n339) );
  MUX21X1_HVT U121 ( .A1(n421), .A2(n334), .S0(n298), .Y(n590) );
  MUX21X1_HVT U123 ( .A1(n278), .A2(n417), .S0(n298), .Y(n483) );
  MUX21X2_HVT U125 ( .A1(n596), .A2(n318), .S0(n326), .Y(n504) );
  INVX1_HVT U126 ( .A(n356), .Y(n290) );
  INVX2_HVT U127 ( .A(n290), .Y(n357) );
  MUX41X1_HVT U128 ( .A1(n483), .A3(n299), .A2(n397), .A4(n309), .S0(n241), 
        .S1(n229), .Y(n482) );
  IBUFFX4_HVT U134 ( .A(n328), .Y(n229) );
  MUX41X1_HVT U135 ( .A1(n248), .A3(n373), .A2(n309), .A4(n370), .S0(n229), 
        .S1(n265), .Y(n450) );
  INVX1_HVT U136 ( .A(n304), .Y(n307) );
  INVX1_HVT U138 ( .A(n262), .Y(n240) );
  INVX1_HVT U142 ( .A(n261), .Y(n234) );
  AOI21X2_HVT U144 ( .A1(n360), .A2(n505), .A3(n374), .Y(n506) );
  MUX21X2_HVT U145 ( .A1(n500), .A2(n499), .S0(n338), .Y(n498) );
  INVX2_HVT U146 ( .A(n291), .Y(n297) );
  MUX41X1_HVT U147 ( .A1(n590), .A3(n492), .A2(n389), .A4(n414), .S0(n230), 
        .S1(n304), .Y(n491) );
  IBUFFX16_HVT U149 ( .A(n360), .Y(n230) );
  IBUFFX2_HVT U150 ( .A(n590), .Y(n398) );
  MUX21X2_HVT U151 ( .A1(n310), .A2(n277), .S0(n354), .Y(n231) );
  INVX0_HVT U152 ( .A(n310), .Y(n313) );
  MUX21X2_HVT U153 ( .A1(n520), .A2(n521), .S0(n358), .Y(n519) );
  INVX1_HVT U154 ( .A(n353), .Y(n279) );
  MUX41X1_HVT U157 ( .A1(n549), .A3(n489), .A2(n412), .A4(n598), .S0(n233), 
        .S1(n234), .Y(n488) );
  IBUFFX16_HVT U158 ( .A(n327), .Y(n233) );
  INVX0_HVT U160 ( .A(n354), .Y(n237) );
  XNOR2X2_HVT U161 ( .A1(n336), .A2(n271), .Y(n613) );
  INVX0_HVT U165 ( .A(n290), .Y(n236) );
  INVX0_HVT U167 ( .A(n290), .Y(n291) );
  NBUFFX2_HVT U169 ( .A(n418), .Y(n334) );
  MUX21X1_HVT U171 ( .A1(n310), .A2(n346), .S0(n237), .Y(n424) );
  INVX1_HVT U173 ( .A(n424), .Y(n415) );
  MUX41X1_HVT U175 ( .A1(n440), .A3(n441), .A2(n438), .A4(n437), .S0(n329), 
        .S1(n338), .Y(n436) );
  INVX1_HVT U176 ( .A(n595), .Y(n396) );
  NAND2X0_HVT U181 ( .A1(n463), .A2(n266), .Y(n267) );
  INVX0_HVT U182 ( .A(n603), .Y(n390) );
  MUX21X2_HVT U183 ( .A1(n555), .A2(n554), .S0(n329), .Y(n553) );
  INVX1_HVT U184 ( .A(n628), .Y(n420) );
  MUX21X2_HVT U186 ( .A1(n386), .A2(n566), .S0(n323), .Y(n565) );
  MUX21X2_HVT U187 ( .A1(n405), .A2(n366), .S0(n333), .Y(n555) );
  INVX0_HVT U188 ( .A(n334), .Y(n243) );
  MUX41X1_HVT U189 ( .A1(n403), .A3(n390), .A2(n343), .A4(n575), .S0(n239), 
        .S1(n330), .Y(n574) );
  INVX1_HVT U190 ( .A(n240), .Y(n239) );
  MUX21X2_HVT U193 ( .A1(n477), .A2(n487), .S0(n238), .Y(out[5]) );
  IBUFFX16_HVT U195 ( .A(n305), .Y(n238) );
  MUX21X2_HVT U196 ( .A1(n308), .A2(n312), .S0(n263), .Y(n606) );
  MUX21X1_HVT U197 ( .A1(n577), .A2(n578), .S0(n306), .Y(n576) );
  MUX21X2_HVT U199 ( .A1(n346), .A2(n257), .S0(n286), .Y(n280) );
  INVX0_HVT U201 ( .A(n280), .Y(n601) );
  MUX21X1_HVT U202 ( .A1(n277), .A2(n243), .S0(n357), .Y(n242) );
  IBUFFX16_HVT U203 ( .A(n242), .Y(n584) );
  INVX0_HVT U204 ( .A(n435), .Y(n244) );
  NAND2X0_HVT U205 ( .A1(n324), .A2(n245), .Y(n246) );
  NAND2X0_HVT U206 ( .A1(n417), .A2(n276), .Y(n247) );
  NAND2X0_HVT U208 ( .A1(n246), .A2(n247), .Y(n435) );
  INVX0_HVT U209 ( .A(n276), .Y(n245) );
  INVX0_HVT U210 ( .A(n435), .Y(n403) );
  INVX1_HVT U211 ( .A(n422), .Y(n324) );
  INVX0_HVT U212 ( .A(n346), .Y(n417) );
  MUX41X1_HVT U213 ( .A1(n403), .A3(n400), .A2(n587), .A4(n386), .S0(n249), 
        .S1(n326), .Y(n449) );
  AO21X1_HVT U214 ( .A1(n345), .A2(n248), .A3(n240), .Y(n465) );
  MUX21X2_HVT U215 ( .A1(n387), .A2(n575), .S0(n332), .Y(n571) );
  NAND2X2_HVT U216 ( .A1(n236), .A2(n311), .Y(n618) );
  INVX1_HVT U217 ( .A(in[1]), .Y(n338) );
  INVX1_HVT U218 ( .A(n272), .Y(n462) );
  MUX21X2_HVT U219 ( .A1(n273), .A2(n258), .S0(n274), .Y(n272) );
  INVX0_HVT U220 ( .A(n420), .Y(n273) );
  INVX0_HVT U221 ( .A(n419), .Y(n251) );
  INVX1_HVT U222 ( .A(n419), .Y(n252) );
  INVX1_HVT U223 ( .A(n251), .Y(n253) );
  INVX1_HVT U224 ( .A(n252), .Y(n254) );
  INVX0_HVT U225 ( .A(n255), .Y(n257) );
  INVX0_HVT U226 ( .A(n255), .Y(n258) );
  MUX41X1_HVT U227 ( .A1(n493), .A3(n491), .A2(n490), .A4(n488), .S0(n259), 
        .S1(n260), .Y(n487) );
  IBUFFX16_HVT U228 ( .A(n339), .Y(n259) );
  IBUFFX16_HVT U229 ( .A(in[5]), .Y(n260) );
  XNOR2X1_HVT U230 ( .A1(n346), .A2(n235), .Y(n581) );
  MUX41X1_HVT U231 ( .A1(n451), .A3(n448), .A2(n442), .A4(n436), .S0(n341), 
        .S1(n305), .Y(out[7]) );
  MUX21X1_HVT U232 ( .A1(n344), .A2(n253), .S0(n354), .Y(n598) );
  IBUFFX2_HVT U233 ( .A(n364), .Y(n261) );
  IBUFFX2_HVT U234 ( .A(n364), .Y(n262) );
  INVX0_HVT U235 ( .A(n364), .Y(n362) );
  INVX1_HVT U236 ( .A(n336), .Y(n277) );
  INVX0_HVT U237 ( .A(n618), .Y(n365) );
  NBUFFX2_HVT U238 ( .A(n236), .Y(n263) );
  MUX21X1_HVT U239 ( .A1(n388), .A2(n573), .S0(n323), .Y(n572) );
  INVX2_HVT U240 ( .A(n364), .Y(n361) );
  INVX1_HVT U241 ( .A(n351), .Y(n274) );
  INVX1_HVT U242 ( .A(n351), .Y(n286) );
  INVX1_HVT U243 ( .A(n285), .Y(n276) );
  IBUFFX2_HVT U244 ( .A(n354), .Y(n285) );
  INVX1_HVT U245 ( .A(n430), .Y(n408) );
  AO21X1_HVT U246 ( .A1(n263), .A2(n258), .A3(n307), .Y(n473) );
  MUX41X1_HVT U247 ( .A1(n568), .A3(n574), .A2(n572), .A4(n576), .S0(n264), 
        .S1(n340), .Y(n567) );
  IBUFFX16_HVT U248 ( .A(n275), .Y(n264) );
  NBUFFX2_HVT U249 ( .A(n261), .Y(n265) );
  IBUFFX2_HVT U250 ( .A(n364), .Y(n303) );
  INVX2_HVT U251 ( .A(in[0]), .Y(n356) );
  OA21X1_HVT U252 ( .A1(n392), .A2(n240), .A3(n569), .Y(n443) );
  NAND2X0_HVT U253 ( .A1(n456), .A2(n305), .Y(n268) );
  NAND2X0_HVT U254 ( .A1(n267), .A2(n268), .Y(out[6]) );
  IBUFFX2_HVT U255 ( .A(n305), .Y(n266) );
  INVX1_HVT U256 ( .A(in[7]), .Y(n305) );
  MUX21X2_HVT U257 ( .A1(n454), .A2(n452), .S0(n338), .Y(n451) );
  INVX0_HVT U258 ( .A(n625), .Y(n269) );
  INVX1_HVT U259 ( .A(n269), .Y(n270) );
  NBUFFX2_HVT U260 ( .A(n418), .Y(n271) );
  NAND2X0_HVT U261 ( .A1(n277), .A2(n334), .Y(n625) );
  IBUFFX16_HVT U262 ( .A(in[5]), .Y(n275) );
  NBUFFX2_HVT U263 ( .A(n422), .Y(n336) );
  IBUFFX2_HVT U264 ( .A(n364), .Y(n363) );
  IBUFFX2_HVT U265 ( .A(n343), .Y(n296) );
  INVX2_HVT U266 ( .A(n341), .Y(n342) );
  MUX21X2_HVT U267 ( .A1(n311), .A2(n344), .S0(n279), .Y(n299) );
  INVX1_HVT U268 ( .A(n350), .Y(n419) );
  MUX41X1_HVT U269 ( .A1(n253), .A3(n258), .A2(n593), .A4(n315), .S0(n281), 
        .S1(n363), .Y(n458) );
  IBUFFX16_HVT U270 ( .A(n360), .Y(n281) );
  NAND2X0_HVT U271 ( .A1(n450), .A2(n282), .Y(n283) );
  NAND2X0_HVT U272 ( .A1(n449), .A2(n338), .Y(n284) );
  NAND2X0_HVT U273 ( .A1(n283), .A2(n284), .Y(n448) );
  IBUFFX2_HVT U274 ( .A(n338), .Y(n282) );
  OR2X1_HVT U275 ( .A1(n335), .A2(n422), .Y(n628) );
  IBUFFX2_HVT U276 ( .A(n271), .Y(n308) );
  NAND2X1_HVT U277 ( .A1(n475), .A2(n287), .Y(n288) );
  NAND2X0_HVT U278 ( .A1(n476), .A2(n360), .Y(n289) );
  NAND2X0_HVT U279 ( .A1(n288), .A2(n289), .Y(n472) );
  IBUFFX2_HVT U280 ( .A(n360), .Y(n287) );
  MUX21X1_HVT U281 ( .A1(n586), .A2(n405), .S0(n332), .Y(n476) );
  INVX1_HVT U282 ( .A(in[4]), .Y(n364) );
  MUX41X1_HVT U283 ( .A1(n398), .A3(n392), .A2(n367), .A4(n614), .S0(n328), 
        .S1(n361), .Y(n516) );
  MUX41X1_HVT U284 ( .A1(n386), .A3(n343), .A2(n390), .A4(n315), .S0(n330), 
        .S1(n265), .Y(n524) );
  MUX21X1_HVT U285 ( .A1(n389), .A2(n626), .S0(n360), .Y(n573) );
  MUX41X1_HVT U286 ( .A1(n580), .A3(n531), .A2(n497), .A4(n378), .S0(n325), 
        .S1(n331), .Y(n496) );
  INVX0_HVT U287 ( .A(n305), .Y(n302) );
  INVX1_HVT U288 ( .A(n604), .Y(n389) );
  NAND2X0_HVT U289 ( .A1(n334), .A2(n292), .Y(n293) );
  NAND2X0_HVT U290 ( .A1(n420), .A2(n298), .Y(n294) );
  NAND2X0_HVT U291 ( .A1(n293), .A2(n294), .Y(n586) );
  INVX0_HVT U292 ( .A(n298), .Y(n292) );
  INVX0_HVT U293 ( .A(n586), .Y(n400) );
  INVX1_HVT U294 ( .A(n356), .Y(n352) );
  IBUFFX2_HVT U295 ( .A(n356), .Y(n353) );
  NAND2X0_HVT U296 ( .A1(n352), .A2(n256), .Y(n624) );
  NAND2X0_HVT U297 ( .A1(n355), .A2(n315), .Y(n627) );
  INVX1_HVT U298 ( .A(n295), .Y(n309) );
  MUX21X1_HVT U299 ( .A1(n296), .A2(n335), .S0(n292), .Y(n295) );
  NAND2X0_HVT U300 ( .A1(n529), .A2(n305), .Y(n300) );
  NAND2X0_HVT U301 ( .A1(n536), .A2(n302), .Y(n301) );
  NAND2X0_HVT U302 ( .A1(n301), .A2(n300), .Y(out[2]) );
  MUX21X1_HVT U303 ( .A1(n604), .A2(n321), .S0(n332), .Y(n481) );
  INVX1_HVT U304 ( .A(n602), .Y(n391) );
  MUX21X2_HVT U305 ( .A1(n480), .A2(n481), .S0(n360), .Y(n479) );
  INVX1_HVT U306 ( .A(n433), .Y(n405) );
  INVX1_HVT U307 ( .A(n432), .Y(n406) );
  IBUFFX2_HVT U308 ( .A(n356), .Y(n354) );
  MUX41X1_HVT U309 ( .A1(n459), .A3(n461), .A2(n457), .A4(n458), .S0(n339), 
        .S1(n341), .Y(n456) );
  INVX2_HVT U310 ( .A(n364), .Y(n304) );
  OA21X2_HVT U311 ( .A1(n369), .A2(n240), .A3(n608), .Y(n554) );
  OA21X2_HVT U312 ( .A1(n368), .A2(n240), .A3(n377), .Y(n480) );
  AO21X2_HVT U313 ( .A1(n351), .A2(n313), .A3(n307), .Y(n439) );
  INVX0_HVT U314 ( .A(n316), .Y(n585) );
  INVX1_HVT U315 ( .A(n343), .Y(n421) );
  INVX0_HVT U316 ( .A(n330), .Y(n306) );
  IBUFFX2_HVT U317 ( .A(n356), .Y(n355) );
  IBUFFX2_HVT U318 ( .A(n356), .Y(n351) );
  MUX41X1_HVT U319 ( .A1(n591), .A3(n384), .A2(n385), .A4(n383), .S0(n306), 
        .S1(n234), .Y(n564) );
  NBUFFX2_HVT U320 ( .A(n418), .Y(n335) );
  INVX0_HVT U321 ( .A(in[3]), .Y(n418) );
  INVX1_HVT U322 ( .A(n311), .Y(n312) );
  MUX21X1_HVT U323 ( .A1(n258), .A2(n346), .S0(n263), .Y(n316) );
  INVX0_HVT U324 ( .A(in[5]), .Y(n341) );
  MUX21X1_HVT U325 ( .A1(n242), .A2(n320), .S0(n331), .Y(n438) );
  AND2X1_HVT U326 ( .A1(n624), .A2(n310), .Y(n317) );
  AND2X1_HVT U327 ( .A1(n310), .A2(n614), .Y(n318) );
  NAND2X0_HVT U328 ( .A1(n335), .A2(n278), .Y(n629) );
  MUX21X1_HVT U329 ( .A1(n278), .A2(n313), .S0(n355), .Y(n603) );
  MUX21X1_HVT U330 ( .A1(n312), .A2(n420), .S0(n353), .Y(n579) );
  MUX21X1_HVT U331 ( .A1(n254), .A2(n337), .S0(n354), .Y(n460) );
  MUX21X1_HVT U332 ( .A1(n344), .A2(n335), .S0(n351), .Y(n608) );
  MUX21X1_HVT U333 ( .A1(n334), .A2(n312), .S0(n298), .Y(n599) );
  MUX21X1_HVT U334 ( .A1(n346), .A2(n348), .S0(n298), .Y(n471) );
  MUX21X1_HVT U335 ( .A1(n311), .A2(n270), .S0(n355), .Y(n489) );
  MUX21X1_HVT U336 ( .A1(n345), .A2(n417), .S0(n355), .Y(n595) );
  MUX21X1_HVT U337 ( .A1(n421), .A2(n337), .S0(n351), .Y(n425) );
  MUX21X1_HVT U338 ( .A1(n334), .A2(n315), .S0(n351), .Y(n432) );
  MUX21X1_HVT U339 ( .A1(n345), .A2(n337), .S0(n354), .Y(n604) );
  MUX21X1_HVT U340 ( .A1(n420), .A2(n335), .S0(n355), .Y(n433) );
  MUX21X1_HVT U341 ( .A1(n253), .A2(n345), .S0(n355), .Y(n430) );
  XNOR2X1_HVT U342 ( .A1(n311), .A2(n297), .Y(n319) );
  XOR2X1_HVT U343 ( .A1(n347), .A2(n354), .Y(n582) );
  MUX21X1_HVT U344 ( .A1(n257), .A2(n315), .S0(n353), .Y(n615) );
  MUX21X1_HVT U345 ( .A1(n349), .A2(n315), .S0(n353), .Y(n611) );
  MUX21X1_HVT U346 ( .A1(n348), .A2(n335), .S0(n221), .Y(n610) );
  MUX21X1_HVT U347 ( .A1(n278), .A2(n310), .S0(n297), .Y(n526) );
  MUX21X1_HVT U348 ( .A1(n414), .A2(n319), .S0(n358), .Y(n507) );
  XOR2X1_HVT U349 ( .A1(n343), .A2(n352), .Y(n583) );
  XOR2X1_HVT U350 ( .A1(n256), .A2(n351), .Y(n592) );
  MUX21X1_HVT U351 ( .A1(n278), .A2(n345), .S0(n353), .Y(n589) );
  MUX21X1_HVT U352 ( .A1(n334), .A2(n348), .S0(n353), .Y(n427) );
  MUX21X1_HVT U353 ( .A1(n349), .A2(n278), .S0(n352), .Y(n510) );
  NBUFFX2_HVT U354 ( .A(n362), .Y(n333) );
  AND2X1_HVT U355 ( .A1(n353), .A2(n337), .Y(n320) );
  NBUFFX2_HVT U356 ( .A(n625), .Y(n346) );
  NBUFFX2_HVT U357 ( .A(n613), .Y(n343) );
  MUX21X1_HVT U358 ( .A1(n391), .A2(n381), .S0(n333), .Y(n578) );
  NBUFFX2_HVT U359 ( .A(n613), .Y(n344) );
  AND2X1_HVT U360 ( .A1(n349), .A2(n235), .Y(n321) );
  AND2X1_HVT U361 ( .A1(n420), .A2(n357), .Y(n322) );
  NBUFFX2_HVT U362 ( .A(n628), .Y(n347) );
  NBUFFX2_HVT U363 ( .A(n628), .Y(n349) );
  NBUFFX2_HVT U364 ( .A(n613), .Y(n345) );
  NBUFFX2_HVT U365 ( .A(n628), .Y(n348) );
  XNOR2X1_HVT U366 ( .A1(n307), .A2(n328), .Y(n323) );
  NBUFFX2_HVT U367 ( .A(n359), .Y(n328) );
  NBUFFX2_HVT U368 ( .A(n358), .Y(n326) );
  NBUFFX2_HVT U369 ( .A(n359), .Y(n329) );
  NBUFFX2_HVT U370 ( .A(n359), .Y(n330) );
  NBUFFX2_HVT U371 ( .A(n358), .Y(n327) );
  NBUFFX2_HVT U372 ( .A(n358), .Y(n325) );
  INVX1_HVT U373 ( .A(n338), .Y(n340) );
  MUX21X1_HVT U374 ( .A1(n270), .A2(n308), .S0(n297), .Y(n534) );
  MUX21X1_HVT U375 ( .A1(n254), .A2(n308), .S0(n297), .Y(n423) );
  MUX21X1_HVT U376 ( .A1(n495), .A2(n496), .S0(n339), .Y(n494) );
  MUX21X1_HVT U377 ( .A1(n420), .A2(n417), .S0(n352), .Y(n515) );
  MUX21X1_HVT U378 ( .A1(n308), .A2(n270), .S0(n353), .Y(n428) );
  MUX21X1_HVT U379 ( .A1(n258), .A2(n308), .S0(n221), .Y(n474) );
  MUX21X1_HVT U380 ( .A1(n308), .A2(n257), .S0(n351), .Y(n429) );
  MUX21X1_HVT U381 ( .A1(n337), .A2(n308), .S0(n297), .Y(n602) );
  NBUFFX2_HVT U382 ( .A(in[2]), .Y(n360) );
  NBUFFX2_HVT U383 ( .A(in[2]), .Y(n359) );
  NBUFFX2_HVT U384 ( .A(in[2]), .Y(n358) );
  MUX21X1_HVT U385 ( .A1(n312), .A2(n324), .S0(n351), .Y(n497) );
  XOR2X1_HVT U386 ( .A1(n298), .A2(n324), .Y(n580) );
  MUX21X1_HVT U387 ( .A1(n348), .A2(n324), .S0(n352), .Y(n431) );
  MUX21X1_HVT U388 ( .A1(n324), .A2(n254), .S0(n298), .Y(n605) );
  MUX21X1_HVT U389 ( .A1(n324), .A2(n256), .S0(n297), .Y(n612) );
  MUX21X1_HVT U390 ( .A1(n324), .A2(n349), .S0(n297), .Y(n434) );
  MUX21X1_HVT U391 ( .A1(n335), .A2(n324), .S0(n355), .Y(n426) );
  MUX21X1_HVT U392 ( .A1(n270), .A2(n324), .S0(n355), .Y(n600) );
  NBUFFX2_HVT U393 ( .A(n630), .Y(n350) );
  INVX0_HVT U394 ( .A(n597), .Y(n366) );
  INVX0_HVT U395 ( .A(n591), .Y(n367) );
  INVX0_HVT U396 ( .A(n531), .Y(n368) );
  INVX0_HVT U397 ( .A(n492), .Y(n369) );
  INVX0_HVT U398 ( .A(n626), .Y(n371) );
  INVX0_HVT U399 ( .A(n624), .Y(n372) );
  INVX0_HVT U400 ( .A(n623), .Y(n374) );
  INVX0_HVT U401 ( .A(n622), .Y(n375) );
  INVX0_HVT U402 ( .A(n594), .Y(n376) );
  INVX0_HVT U403 ( .A(n616), .Y(n377) );
  INVX0_HVT U404 ( .A(n621), .Y(n378) );
  INVX0_HVT U405 ( .A(n617), .Y(n379) );
  INVX0_HVT U406 ( .A(n615), .Y(n380) );
  INVX0_HVT U407 ( .A(n614), .Y(n381) );
  INVX0_HVT U408 ( .A(n612), .Y(n382) );
  INVX0_HVT U409 ( .A(n611), .Y(n383) );
  INVX0_HVT U410 ( .A(n610), .Y(n384) );
  INVX0_HVT U411 ( .A(n609), .Y(n385) );
  INVX0_HVT U412 ( .A(n608), .Y(n386) );
  INVX0_HVT U413 ( .A(n606), .Y(n387) );
  INVX0_HVT U414 ( .A(n605), .Y(n388) );
  INVX0_HVT U415 ( .A(n600), .Y(n392) );
  INVX0_HVT U416 ( .A(n599), .Y(n393) );
  INVX0_HVT U417 ( .A(n598), .Y(n394) );
  INVX0_HVT U418 ( .A(n596), .Y(n395) );
  INVX0_HVT U419 ( .A(n592), .Y(n397) );
  INVX0_HVT U420 ( .A(n589), .Y(n399) );
  INVX0_HVT U421 ( .A(n583), .Y(n401) );
  INVX0_HVT U422 ( .A(n620), .Y(n402) );
  INVX0_HVT U423 ( .A(n434), .Y(n404) );
  INVX0_HVT U424 ( .A(n431), .Y(n407) );
  INVX0_HVT U425 ( .A(n429), .Y(n409) );
  INVX0_HVT U426 ( .A(n428), .Y(n410) );
  INVX0_HVT U427 ( .A(n427), .Y(n411) );
  INVX0_HVT U428 ( .A(n426), .Y(n412) );
  INVX0_HVT U429 ( .A(n474), .Y(n413) );
  INVX0_HVT U430 ( .A(n423), .Y(n416) );
endmodule

