
module sbox_10 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n23, n45, n48, n50, n72, n210, n211, n212, n213, n216, n217, n218,
         n219, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591;

  NAND2X0_HVT U4 ( .A1(n295), .A2(n589), .Y(n588) );
  NAND2X0_HVT U5 ( .A1(n305), .A2(n371), .Y(n586) );
  NAND2X0_HVT U15 ( .A1(n589), .A2(n287), .Y(n576) );
  NAND2X0_HVT U21 ( .A1(n294), .A2(n307), .Y(n570) );
  NAND2X0_HVT U24 ( .A1(n291), .A2(n307), .Y(n568) );
  NAND2X0_HVT U33 ( .A1(n369), .A2(n50), .Y(n559) );
  NAND2X0_HVT U35 ( .A1(n289), .A2(n48), .Y(n557) );
  NAND2X0_HVT U42 ( .A1(n241), .A2(n291), .Y(n550) );
  MUX41X1_HVT U51 ( .A1(n357), .A3(n317), .A2(n335), .A4(n336), .S0(n314), 
        .S1(n311), .Y(n544) );
  NAND2X0_HVT U53 ( .A1(n541), .A2(n549), .Y(n542) );
  NAND2X0_HVT U56 ( .A1(n295), .A2(n537), .Y(n538) );
  MUX41X1_HVT U57 ( .A1(n358), .A3(n572), .A2(n538), .A4(n581), .S0(n314), 
        .S1(in[5]), .Y(n536) );
  NAND2X0_HVT U58 ( .A1(n299), .A2(n589), .Y(n535) );
  MUX41X1_HVT U59 ( .A1(n276), .A3(n535), .A2(n274), .A4(n334), .S0(n314), 
        .S1(in[5]), .Y(n534) );
  NAND2X0_HVT U62 ( .A1(n48), .A2(n298), .Y(n531) );
  MUX41X1_HVT U63 ( .A1(n531), .A3(n324), .A2(n248), .A4(n331), .S0(n314), 
        .S1(n282), .Y(n530) );
  AO21X1_HVT U66 ( .A1(n329), .A2(n282), .A3(n352), .Y(n527) );
  MUX41X1_HVT U68 ( .A1(n327), .A3(n527), .A2(n526), .A4(n528), .S0(n277), 
        .S1(n313), .Y(n525) );
  MUX41X1_HVT U69 ( .A1(n525), .A3(n533), .A2(n529), .A4(n539), .S0(in[6]), 
        .S1(in[0]), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n292), .A2(n521), .Y(n522) );
  MUX41X1_HVT U74 ( .A1(n523), .A3(n566), .A2(n522), .A4(n568), .S0(n279), 
        .S1(n312), .Y(n520) );
  MUX41X1_HVT U75 ( .A1(n355), .A3(n360), .A2(n373), .A4(n242), .S0(n277), 
        .S1(n312), .Y(n519) );
  MUX41X1_HVT U77 ( .A1(n583), .A3(n362), .A2(n518), .A4(n361), .S0(n283), 
        .S1(n308), .Y(n517) );
  MUX41X1_HVT U78 ( .A1(n517), .A3(n520), .A2(n519), .A4(n524), .S0(in[0]), 
        .S1(in[5]), .Y(n516) );
  MUX41X1_HVT U82 ( .A1(n548), .A3(n336), .A2(n318), .A4(n577), .S0(n277), 
        .S1(n260), .Y(n511) );
  AND2X1_HVT U83 ( .A1(n241), .A2(n234), .Y(n510) );
  MUX41X1_HVT U84 ( .A1(n337), .A3(n585), .A2(n575), .A4(n510), .S0(n277), 
        .S1(n260), .Y(n509) );
  NAND2X0_HVT U85 ( .A1(n50), .A2(n372), .Y(n508) );
  MUX41X1_HVT U86 ( .A1(n360), .A3(n508), .A2(n273), .A4(n269), .S0(n277), 
        .S1(n313), .Y(n507) );
  MUX41X1_HVT U87 ( .A1(n507), .A3(n511), .A2(n509), .A4(n512), .S0(in[0]), 
        .S1(n311), .Y(n506) );
  MUX41X1_HVT U90 ( .A1(n547), .A3(n550), .A2(n357), .A4(n505), .S0(n278), 
        .S1(n233), .Y(n504) );
  AO21X1_HVT U93 ( .A1(n285), .A2(n500), .A3(n356), .Y(n501) );
  MUX41X1_HVT U96 ( .A1(n318), .A3(n271), .A2(n359), .A4(n498), .S0(n277), 
        .S1(n312), .Y(n497) );
  MUX41X1_HVT U97 ( .A1(n355), .A3(n271), .A2(n302), .A4(n576), .S0(n277), 
        .S1(n312), .Y(n496) );
  MUX41X1_HVT U98 ( .A1(n496), .A3(n499), .A2(n497), .A4(n504), .S0(in[0]), 
        .S1(in[5]), .Y(n495) );
  NAND2X0_HVT U101 ( .A1(n491), .A2(n490), .Y(n492) );
  MUX41X1_HVT U103 ( .A1(n589), .A3(n328), .A2(n340), .A4(n557), .S0(n277), 
        .S1(n313), .Y(n488) );
  MUX41X1_HVT U105 ( .A1(n339), .A3(n546), .A2(n487), .A4(n354), .S0(n277), 
        .S1(n312), .Y(n486) );
  MUX21X2_HVT U107 ( .A1(n485), .A2(n495), .S0(in[6]), .Y(out[2]) );
  OA21X1_HVT U109 ( .A1(n347), .A2(n310), .A3(n334), .Y(n483) );
  NAND2X0_HVT U110 ( .A1(n297), .A2(n481), .Y(n482) );
  MUX41X1_HVT U114 ( .A1(n478), .A3(n484), .A2(n480), .A4(n483), .S0(n282), 
        .S1(n313), .Y(n477) );
  AND2X1_HVT U115 ( .A1(n303), .A2(n287), .Y(n476) );
  MUX41X1_HVT U116 ( .A1(n579), .A3(n476), .A2(n242), .A4(n561), .S0(n278), 
        .S1(n314), .Y(n475) );
  NAND2X0_HVT U123 ( .A1(n467), .A2(n466), .Y(n468) );
  MUX41X1_HVT U125 ( .A1(n570), .A3(n276), .A2(n327), .A4(n364), .S0(n278), 
        .S1(n314), .Y(n464) );
  MUX41X1_HVT U131 ( .A1(n459), .A3(n461), .A2(n460), .A4(n462), .S0(n282), 
        .S1(n314), .Y(n458) );
  MUX41X1_HVT U136 ( .A1(n269), .A3(n559), .A2(n366), .A4(n556), .S0(n278), 
        .S1(n314), .Y(n454) );
  AND2X1_HVT U140 ( .A1(n293), .A2(n48), .Y(n450) );
  OA21X1_HVT U144 ( .A1(n321), .A2(n315), .A3(n561), .Y(n446) );
  NAND2X0_HVT U146 ( .A1(n241), .A2(n300), .Y(n521) );
  MUX41X1_HVT U147 ( .A1(n366), .A3(n521), .A2(n355), .A4(n547), .S0(n279), 
        .S1(n314), .Y(n444) );
  MUX41X1_HVT U148 ( .A1(n444), .A3(n448), .A2(n445), .A4(n449), .S0(in[0]), 
        .S1(in[5]), .Y(n443) );
  OA21X1_HVT U151 ( .A1(n552), .A2(n315), .A3(n440), .Y(n441) );
  MUX41X1_HVT U153 ( .A1(n482), .A3(n272), .A2(n296), .A4(n320), .S0(n278), 
        .S1(n233), .Y(n438) );
  AND2X1_HVT U154 ( .A1(n285), .A2(n291), .Y(n437) );
  NAND2X0_HVT U158 ( .A1(n304), .A2(n372), .Y(n433) );
  MUX41X1_HVT U159 ( .A1(n579), .A3(n287), .A2(n433), .A4(n326), .S0(n309), 
        .S1(n233), .Y(n432) );
  AND2X1_HVT U162 ( .A1(n585), .A2(n521), .Y(n429) );
  NAND2X0_HVT U166 ( .A1(n299), .A2(n537), .Y(n425) );
  NAND2X0_HVT U167 ( .A1(n373), .A2(n48), .Y(n424) );
  MUX41X1_HVT U168 ( .A1(n358), .A3(n292), .A2(n424), .A4(n425), .S0(n309), 
        .S1(n233), .Y(n423) );
  OA21X1_HVT U170 ( .A1(n274), .A2(n315), .A3(n561), .Y(n421) );
  MUX41X1_HVT U172 ( .A1(n420), .A3(n426), .A2(n423), .A4(n428), .S0(in[0]), 
        .S1(n311), .Y(n419) );
  NAND2X0_HVT U174 ( .A1(n303), .A2(n585), .Y(n578) );
  NAND2X0_HVT U177 ( .A1(n305), .A2(n289), .Y(n416) );
  MUX41X1_HVT U178 ( .A1(n574), .A3(n416), .A2(n367), .A4(n554), .S0(n279), 
        .S1(n312), .Y(n415) );
  MUX41X1_HVT U179 ( .A1(n564), .A3(n368), .A2(n322), .A4(n367), .S0(n309), 
        .S1(n313), .Y(n414) );
  MUX41X1_HVT U180 ( .A1(n325), .A3(n583), .A2(n579), .A4(n268), .S0(n283), 
        .S1(n309), .Y(n413) );
  OA21X1_HVT U184 ( .A1(n558), .A2(n315), .A3(n337), .Y(n409) );
  MUX41X1_HVT U186 ( .A1(n271), .A3(n553), .A2(n521), .A4(n547), .S0(n309), 
        .S1(n233), .Y(n407) );
  MUX41X1_HVT U189 ( .A1(n405), .A3(n578), .A2(n406), .A4(n354), .S0(n283), 
        .S1(n309), .Y(n404) );
  MUX41X1_HVT U190 ( .A1(n404), .A3(n407), .A2(n408), .A4(n411), .S0(n311), 
        .S1(in[0]), .Y(n403) );
  MUX41X1_HVT U193 ( .A1(n550), .A3(n557), .A2(n545), .A4(n402), .S0(n309), 
        .S1(n260), .Y(n401) );
  AO21X1_HVT U197 ( .A1(n273), .A2(n284), .A3(n356), .Y(n397) );
  MUX41X1_HVT U199 ( .A1(n396), .A3(n400), .A2(n399), .A4(n401), .S0(in[0]), 
        .S1(n311), .Y(n395) );
  OA21X1_HVT U201 ( .A1(n584), .A2(n315), .A3(n348), .Y(n393) );
  MUX41X1_HVT U203 ( .A1(n556), .A3(n237), .A2(n580), .A4(n560), .S0(n309), 
        .S1(n233), .Y(n391) );
  NAND2X0_HVT U208 ( .A1(n240), .A2(n294), .Y(n481) );
  NAND2X0_HVT U212 ( .A1(n304), .A2(n292), .Y(n537) );
  NAND2X0_HVT U214 ( .A1(n585), .A2(n48), .Y(n387) );
  NAND2X0_HVT U215 ( .A1(n481), .A2(n293), .Y(n386) );
  NAND2X0_HVT U218 ( .A1(n370), .A2(n303), .Y(n440) );
  NAND2X0_HVT U220 ( .A1(n284), .A2(n387), .Y(n513) );
  MUX41X1_HVT U1 ( .A1(n477), .A3(n463), .A2(n471), .A4(n458), .S0(n23), .S1(
        n45), .Y(out[3]) );
  IBUFFX16_HVT U2 ( .A(in[6]), .Y(n23) );
  IBUFFX16_HVT U3 ( .A(in[0]), .Y(n45) );
  MUX21X2_HVT U6 ( .A1(n540), .A2(n544), .S0(n279), .Y(n539) );
  INVX1_HVT U7 ( .A(in[1]), .Y(n48) );
  INVX1_HVT U8 ( .A(in[1]), .Y(n50) );
  INVX0_HVT U9 ( .A(in[1]), .Y(n306) );
  INVX1_HVT U10 ( .A(n48), .Y(n303) );
  MUX21X1_HVT U11 ( .A1(n373), .A2(n291), .S0(n301), .Y(n572) );
  MUX21X1_HVT U12 ( .A1(n268), .A2(n575), .S0(n259), .Y(n394) );
  NAND2X1_HVT U13 ( .A1(n241), .A2(n297), .Y(n589) );
  INVX1_HVT U14 ( .A(n310), .Y(n309) );
  MUX21X2_HVT U16 ( .A1(n542), .A2(n543), .S0(n283), .Y(n540) );
  NAND2X0_HVT U17 ( .A1(n514), .A2(n72), .Y(n210) );
  NAND2X0_HVT U18 ( .A1(n515), .A2(n235), .Y(n211) );
  NAND2X0_HVT U19 ( .A1(n210), .A2(n211), .Y(n512) );
  INVX0_HVT U20 ( .A(n235), .Y(n72) );
  AND3X2_HVT U22 ( .A1(n297), .A2(n537), .A3(n513), .Y(n514) );
  MUX21X1_HVT U23 ( .A1(n571), .A2(n293), .S0(n285), .Y(n515) );
  IBUFFX2_HVT U25 ( .A(n281), .Y(n235) );
  MUX21X1_HVT U26 ( .A1(n591), .A2(n383), .S0(n285), .Y(n212) );
  MUX21X2_HVT U27 ( .A1(n516), .A2(n506), .S0(n213), .Y(out[1]) );
  IBUFFX16_HVT U28 ( .A(in[6]), .Y(n213) );
  MUX21X2_HVT U29 ( .A1(n349), .A2(n569), .S0(n259), .Y(n453) );
  MUX21X2_HVT U30 ( .A1(n453), .A2(n588), .S0(n281), .Y(n452) );
  NAND2X0_HVT U31 ( .A1(n234), .A2(n216), .Y(n217) );
  NAND2X0_HVT U32 ( .A1(n298), .A2(n240), .Y(n218) );
  NAND2X0_HVT U34 ( .A1(n217), .A2(n218), .Y(n571) );
  INVX0_HVT U36 ( .A(n240), .Y(n216) );
  IBUFFX2_HVT U37 ( .A(n306), .Y(n240) );
  INVX0_HVT U38 ( .A(n571), .Y(n336) );
  INVX1_HVT U39 ( .A(n306), .Y(n241) );
  INVX0_HVT U40 ( .A(n565), .Y(n232) );
  INVX0_HVT U41 ( .A(n302), .Y(n243) );
  IBUFFX2_HVT U43 ( .A(n50), .Y(n302) );
  MUX21X2_HVT U44 ( .A1(n298), .A2(n479), .S0(n267), .Y(n478) );
  INVX1_HVT U45 ( .A(n316), .Y(n245) );
  XOR2X1_HVT U46 ( .A1(n309), .A2(n316), .Y(n266) );
  INVX2_HVT U47 ( .A(n316), .Y(n314) );
  XNOR2X1_HVT U48 ( .A1(n315), .A2(n565), .Y(n251) );
  MUX41X1_HVT U49 ( .A1(n231), .A3(n232), .A2(n378), .A4(n582), .S0(n279), 
        .S1(n316), .Y(n219) );
  IBUFFX16_HVT U50 ( .A(n219), .Y(n455) );
  IBUFFX16_HVT U52 ( .A(n586), .Y(n231) );
  INVX0_HVT U54 ( .A(n582), .Y(n370) );
  INVX0_HVT U55 ( .A(in[7]), .Y(n315) );
  DELLN1X2_HVT U60 ( .A(in[7]), .Y(n284) );
  DELLN1X2_HVT U61 ( .A(in[7]), .Y(n283) );
  INVX1_HVT U64 ( .A(n315), .Y(n233) );
  INVX0_HVT U65 ( .A(n315), .Y(n260) );
  IBUFFX16_HVT U67 ( .A(n311), .Y(n249) );
  NBUFFX16_HVT U70 ( .A(in[5]), .Y(n311) );
  INVX1_HVT U71 ( .A(n310), .Y(n308) );
  MUX41X1_HVT U72 ( .A1(n234), .A3(n589), .A2(n368), .A4(n343), .S0(n309), 
        .S1(n313), .Y(n389) );
  INVX0_HVT U76 ( .A(n309), .Y(n236) );
  INVX1_HVT U79 ( .A(n260), .Y(n259) );
  INVX4_HVT U80 ( .A(in[2]), .Y(n310) );
  NBUFFX2_HVT U81 ( .A(in[4]), .Y(n234) );
  INVX1_HVT U88 ( .A(n379), .Y(n364) );
  MUX21X1_HVT U89 ( .A1(n419), .A2(n431), .S0(in[6]), .Y(out[5]) );
  MUX21X1_HVT U91 ( .A1(n296), .A2(n256), .S0(n243), .Y(n242) );
  INVX1_HVT U92 ( .A(n248), .Y(n579) );
  MUX21X1_HVT U94 ( .A1(n295), .A2(n585), .S0(n305), .Y(n555) );
  MUX41X1_HVT U95 ( .A1(n359), .A3(n585), .A2(n555), .A4(n299), .S0(n236), 
        .S1(n260), .Y(n399) );
  NBUFFX2_HVT U99 ( .A(n374), .Y(n289) );
  MUX21X1_HVT U100 ( .A1(n238), .A2(n296), .S0(n304), .Y(n237) );
  IBUFFX16_HVT U102 ( .A(n237), .Y(n552) );
  IBUFFX16_HVT U104 ( .A(n286), .Y(n238) );
  MUX21X2_HVT U106 ( .A1(n442), .A2(n441), .S0(n239), .Y(n439) );
  IBUFFX16_HVT U108 ( .A(n281), .Y(n239) );
  IBUFFX16_HVT U111 ( .A(n242), .Y(n567) );
  MUX41X1_HVT U112 ( .A1(n567), .A3(n348), .A2(n450), .A4(n344), .S0(n244), 
        .S1(n245), .Y(n449) );
  IBUFFX16_HVT U113 ( .A(n247), .Y(n244) );
  INVX1_HVT U117 ( .A(n256), .Y(n585) );
  MUX21X2_HVT U118 ( .A1(n451), .A2(n443), .S0(n246), .Y(out[4]) );
  IBUFFX16_HVT U119 ( .A(in[6]), .Y(n246) );
  IBUFFX2_HVT U120 ( .A(n306), .Y(n304) );
  INVX1_HVT U121 ( .A(n587), .Y(n369) );
  MUX21X1_HVT U122 ( .A1(n372), .A2(n369), .S0(n301), .Y(n554) );
  NAND2X0_HVT U124 ( .A1(n412), .A2(in[6]), .Y(n257) );
  INVX0_HVT U126 ( .A(n303), .Y(n255) );
  INVX1_HVT U127 ( .A(n554), .Y(n348) );
  XOR2X1_HVT U128 ( .A1(n256), .A2(n307), .Y(n547) );
  INVX1_HVT U129 ( .A(n296), .Y(n373) );
  MUX21X1_HVT U130 ( .A1(n554), .A2(n362), .S0(n283), .Y(n435) );
  INVX0_HVT U132 ( .A(n278), .Y(n247) );
  INVX1_HVT U133 ( .A(in[3]), .Y(n371) );
  MUX41X1_HVT U134 ( .A1(n293), .A3(n353), .A2(n287), .A4(n337), .S0(n247), 
        .S1(n316), .Y(n448) );
  MUX41X1_HVT U135 ( .A1(n493), .A3(n488), .A2(n489), .A4(n486), .S0(n261), 
        .S1(n249), .Y(n485) );
  MUX21X1_HVT U137 ( .A1(n290), .A2(n369), .S0(n301), .Y(n563) );
  INVX1_HVT U138 ( .A(n383), .Y(n359) );
  MUX41X1_HVT U139 ( .A1(n551), .A3(n565), .A2(n365), .A4(n293), .S0(n284), 
        .S1(in[2]), .Y(n400) );
  IBUFFX2_HVT U141 ( .A(n551), .Y(n350) );
  INVX0_HVT U142 ( .A(n250), .Y(n524) );
  MUX21X2_HVT U143 ( .A1(n534), .A2(n536), .S0(n280), .Y(n533) );
  AND2X1_HVT U145 ( .A1(n578), .A2(n299), .Y(n248) );
  AO21X2_HVT U149 ( .A1(n50), .A2(n370), .A3(n315), .Y(n491) );
  MUX21X1_HVT U150 ( .A1(n371), .A2(n288), .S0(n307), .Y(n575) );
  IBUFFX2_HVT U152 ( .A(in[1]), .Y(n307) );
  IBUFFX2_HVT U155 ( .A(n306), .Y(n305) );
  MUX41X1_HVT U156 ( .A1(n434), .A3(n439), .A2(n432), .A4(n438), .S0(in[0]), 
        .S1(n249), .Y(n431) );
  MUX21X2_HVT U157 ( .A1(n435), .A2(n436), .S0(n281), .Y(n434) );
  MUX21X1_HVT U160 ( .A1(n212), .A2(n251), .S0(n247), .Y(n250) );
  NAND2X0_HVT U161 ( .A1(n372), .A2(n252), .Y(n253) );
  NAND2X0_HVT U163 ( .A1(n373), .A2(n255), .Y(n254) );
  NAND2X0_HVT U164 ( .A1(n253), .A2(n254), .Y(n565) );
  INVX0_HVT U165 ( .A(n255), .Y(n252) );
  XNOR2X2_HVT U169 ( .A1(n374), .A2(in[3]), .Y(n256) );
  AND3X2_HVT U171 ( .A1(n281), .A2(n48), .A3(n234), .Y(n461) );
  AO21X2_HVT U173 ( .A1(n281), .A2(n293), .A3(n585), .Y(n473) );
  MUX41X1_HVT U175 ( .A1(n454), .A3(n456), .A2(n452), .A4(n455), .S0(in[0]), 
        .S1(n249), .Y(n451) );
  NAND2X0_HVT U176 ( .A1(n403), .A2(n262), .Y(n258) );
  NAND2X0_HVT U181 ( .A1(n257), .A2(n258), .Y(out[6]) );
  MUX21X2_HVT U182 ( .A1(n393), .A2(n394), .S0(n280), .Y(n392) );
  MUX41X1_HVT U183 ( .A1(n569), .A3(n345), .A2(n579), .A4(n538), .S0(n247), 
        .S1(n259), .Y(n390) );
  INVX1_HVT U185 ( .A(n569), .Y(n337) );
  INVX1_HVT U187 ( .A(n315), .Y(n313) );
  IBUFFX2_HVT U188 ( .A(n315), .Y(n312) );
  NBUFFX2_HVT U191 ( .A(n308), .Y(n278) );
  INVX0_HVT U192 ( .A(in[6]), .Y(n262) );
  INVX1_HVT U194 ( .A(in[0]), .Y(n261) );
  MUX41X1_HVT U195 ( .A1(n287), .A3(n332), .A2(n333), .A4(n272), .S0(n259), 
        .S1(n249), .Y(n532) );
  MUX21X1_HVT U196 ( .A1(n287), .A2(n372), .S0(n50), .Y(n430) );
  MUX41X1_HVT U198 ( .A1(n429), .A3(n333), .A2(n430), .A4(n270), .S0(n310), 
        .S1(n313), .Y(n428) );
  MUX41X1_HVT U200 ( .A1(n392), .A3(n390), .A2(n391), .A4(n389), .S0(n261), 
        .S1(n249), .Y(n388) );
  MUX21X2_HVT U202 ( .A1(n395), .A2(n388), .S0(n262), .Y(out[7]) );
  MUX41X1_HVT U204 ( .A1(n363), .A3(n578), .A2(n289), .A4(n418), .S0(n314), 
        .S1(n310), .Y(n417) );
  MUX41X1_HVT U205 ( .A1(n417), .A3(n414), .A2(n415), .A4(n413), .S0(n261), 
        .S1(n249), .Y(n412) );
  MUX41X1_HVT U206 ( .A1(n338), .A3(n350), .A2(n295), .A4(n349), .S0(n316), 
        .S1(n310), .Y(n411) );
  INVX2_HVT U207 ( .A(in[7]), .Y(n316) );
  XNOR2X1_HVT U209 ( .A1(n307), .A2(n310), .Y(n267) );
  IBUFFX2_HVT U210 ( .A(n306), .Y(n301) );
  MUX41X1_HVT U211 ( .A1(n427), .A3(n547), .A2(n341), .A4(n570), .S0(n316), 
        .S1(n310), .Y(n426) );
  NAND2X0_HVT U213 ( .A1(n494), .A2(n263), .Y(n264) );
  NAND2X0_HVT U216 ( .A1(n272), .A2(n266), .Y(n265) );
  NAND2X0_HVT U217 ( .A1(n264), .A2(n265), .Y(n493) );
  INVX0_HVT U219 ( .A(n266), .Y(n263) );
  MUX21X1_HVT U221 ( .A1(n270), .A2(n332), .S0(n278), .Y(n460) );
  NBUFFX2_HVT U222 ( .A(n256), .Y(n288) );
  NBUFFX2_HVT U223 ( .A(n256), .Y(n287) );
  AND2X1_HVT U224 ( .A1(n288), .A2(n537), .Y(n268) );
  MUX21X1_HVT U225 ( .A1(n369), .A2(n372), .S0(n282), .Y(n541) );
  NBUFFX2_HVT U226 ( .A(n587), .Y(n294) );
  MUX21X1_HVT U227 ( .A1(n328), .A2(n370), .S0(n282), .Y(n526) );
  MUX21X1_HVT U228 ( .A1(n561), .A2(n482), .S0(n278), .Y(n480) );
  NBUFFX2_HVT U229 ( .A(n587), .Y(n295) );
  AND2X1_HVT U230 ( .A1(n297), .A2(n521), .Y(n269) );
  MUX21X1_HVT U231 ( .A1(n288), .A2(n372), .S0(n305), .Y(n584) );
  MUX21X1_HVT U232 ( .A1(n464), .A2(n465), .S0(n282), .Y(n463) );
  MUX21X1_HVT U233 ( .A1(n469), .A2(n468), .S0(n285), .Y(n465) );
  MUX21X1_HVT U234 ( .A1(n297), .A2(n287), .S0(n302), .Y(n551) );
  MUX21X1_HVT U235 ( .A1(n287), .A2(n289), .S0(n301), .Y(n490) );
  MUX21X1_HVT U236 ( .A1(n369), .A2(n373), .S0(n304), .Y(n418) );
  MUX21X1_HVT U237 ( .A1(n288), .A2(n369), .S0(n303), .Y(n498) );
  MUX21X1_HVT U238 ( .A1(n585), .A2(n370), .S0(n241), .Y(n378) );
  MUX21X1_HVT U239 ( .A1(n286), .A2(n585), .S0(n304), .Y(n381) );
  MUX21X1_HVT U240 ( .A1(n473), .A2(n474), .S0(n284), .Y(n472) );
  MUX21X1_HVT U241 ( .A1(n320), .A2(n345), .S0(n278), .Y(n474) );
  MUX21X1_HVT U242 ( .A1(n342), .A2(n457), .S0(n280), .Y(n456) );
  MUX21X1_HVT U243 ( .A1(n364), .A2(n293), .S0(n284), .Y(n457) );
  MUX21X1_HVT U244 ( .A1(n294), .A2(n293), .S0(n240), .Y(n505) );
  MUX21X1_HVT U245 ( .A1(n585), .A2(n289), .S0(n303), .Y(n518) );
  NAND2X0_HVT U246 ( .A1(n290), .A2(n286), .Y(n587) );
  MUX21X1_HVT U247 ( .A1(n369), .A2(n290), .S0(n301), .Y(n379) );
  NBUFFX2_HVT U248 ( .A(n590), .Y(n296) );
  INVX1_HVT U249 ( .A(n591), .Y(n372) );
  MUX21X1_HVT U250 ( .A1(n372), .A2(n371), .S0(n240), .Y(n558) );
  MUX21X1_HVT U251 ( .A1(n370), .A2(n369), .S0(n240), .Y(n573) );
  MUX21X1_HVT U252 ( .A1(n319), .A2(n470), .S0(n279), .Y(n469) );
  MUX21X1_HVT U253 ( .A1(n290), .A2(n371), .S0(n304), .Y(n470) );
  NBUFFX2_HVT U254 ( .A(n590), .Y(n297) );
  MUX21X1_HVT U255 ( .A1(n286), .A2(n300), .S0(n303), .Y(n405) );
  MUX21X1_HVT U256 ( .A1(n300), .A2(n297), .S0(n240), .Y(n406) );
  MUX21X1_HVT U257 ( .A1(n298), .A2(n292), .S0(n304), .Y(n577) );
  MUX21X1_HVT U258 ( .A1(n295), .A2(n300), .S0(n241), .Y(n500) );
  MUX21X1_HVT U259 ( .A1(n371), .A2(n372), .S0(n301), .Y(n581) );
  MUX21X1_HVT U260 ( .A1(n294), .A2(n371), .S0(n302), .Y(n580) );
  MUX21X1_HVT U261 ( .A1(n343), .A2(n577), .S0(n281), .Y(n494) );
  NBUFFX2_HVT U262 ( .A(n590), .Y(n298) );
  XOR2X1_HVT U263 ( .A1(n240), .A2(n370), .Y(n548) );
  MUX21X1_HVT U264 ( .A1(n286), .A2(n290), .S0(n241), .Y(n402) );
  XOR2X1_HVT U265 ( .A1(n296), .A2(n301), .Y(n545) );
  MUX21X1_HVT U266 ( .A1(n296), .A2(n289), .S0(n305), .Y(n385) );
  XNOR2X1_HVT U267 ( .A1(n294), .A2(n301), .Y(n270) );
  MUX21X1_HVT U268 ( .A1(n299), .A2(n292), .S0(n304), .Y(n561) );
  MUX21X1_HVT U269 ( .A1(n296), .A2(n294), .S0(n302), .Y(n377) );
  AND2X1_HVT U270 ( .A1(n241), .A2(n373), .Y(n271) );
  MUX21X1_HVT U271 ( .A1(n292), .A2(n371), .S0(n305), .Y(n383) );
  AND2X1_HVT U272 ( .A1(n299), .A2(n481), .Y(n272) );
  XNOR2X1_HVT U273 ( .A1(n299), .A2(n304), .Y(n273) );
  MUX21X1_HVT U274 ( .A1(n293), .A2(n300), .S0(n280), .Y(n467) );
  MUX21X1_HVT U275 ( .A1(n293), .A2(n289), .S0(n241), .Y(n523) );
  XOR2X1_HVT U276 ( .A1(n290), .A2(n305), .Y(n566) );
  NBUFFX2_HVT U277 ( .A(n371), .Y(n286) );
  NBUFFX2_HVT U278 ( .A(in[7]), .Y(n285) );
  NBUFFX2_HVT U279 ( .A(in[5]), .Y(n282) );
  NBUFFX2_HVT U280 ( .A(n308), .Y(n279) );
  NBUFFX2_HVT U281 ( .A(n308), .Y(n280) );
  NBUFFX2_HVT U282 ( .A(n308), .Y(n281) );
  NBUFFX2_HVT U283 ( .A(n308), .Y(n277) );
  MUX21X1_HVT U284 ( .A1(n288), .A2(n291), .S0(n305), .Y(n569) );
  MUX21X1_HVT U285 ( .A1(n409), .A2(n410), .S0(n280), .Y(n408) );
  MUX21X1_HVT U286 ( .A1(n508), .A2(n291), .S0(n284), .Y(n410) );
  MUX21X1_HVT U287 ( .A1(n530), .A2(n532), .S0(n280), .Y(n529) );
  MUX21X1_HVT U288 ( .A1(n492), .A2(n342), .S0(n280), .Y(n489) );
  XOR2X1_HVT U289 ( .A1(n240), .A2(in[3]), .Y(n546) );
  MUX21X1_HVT U290 ( .A1(n292), .A2(n288), .S0(n302), .Y(n487) );
  MUX21X1_HVT U291 ( .A1(n422), .A2(n421), .S0(n277), .Y(n420) );
  MUX21X1_HVT U292 ( .A1(n293), .A2(n359), .S0(n285), .Y(n422) );
  MUX21X1_HVT U293 ( .A1(n361), .A2(n370), .S0(n284), .Y(n442) );
  AND2X1_HVT U294 ( .A1(n288), .A2(n50), .Y(n274) );
  MUX21X1_HVT U295 ( .A1(n447), .A2(n446), .S0(n281), .Y(n445) );
  MUX21X1_HVT U296 ( .A1(n563), .A2(n323), .S0(n285), .Y(n447) );
  MUX21X1_HVT U297 ( .A1(n370), .A2(n373), .S0(n302), .Y(n427) );
  NAND2X0_HVT U298 ( .A1(in[3]), .A2(n290), .Y(n590) );
  NBUFFX2_HVT U299 ( .A(n374), .Y(n290) );
  MUX21X1_HVT U300 ( .A1(n291), .A2(n369), .S0(n302), .Y(n553) );
  MUX21X1_HVT U301 ( .A1(n346), .A2(n589), .S0(n279), .Y(n484) );
  MUX21X1_HVT U302 ( .A1(n437), .A2(n298), .S0(n275), .Y(n436) );
  MUX21X1_HVT U303 ( .A1(n574), .A2(n344), .S0(n279), .Y(n459) );
  MUX21X1_HVT U304 ( .A1(n291), .A2(n557), .S0(n282), .Y(n543) );
  XOR2X1_HVT U305 ( .A1(n303), .A2(n311), .Y(n549) );
  MUX21X1_HVT U306 ( .A1(n589), .A2(n50), .S0(n280), .Y(n466) );
  MUX21X1_HVT U307 ( .A1(n291), .A2(n370), .S0(n240), .Y(n382) );
  MUX21X1_HVT U308 ( .A1(n330), .A2(n50), .S0(n282), .Y(n528) );
  MUX21X1_HVT U309 ( .A1(n351), .A2(n367), .S0(n284), .Y(n398) );
  NBUFFX2_HVT U310 ( .A(n582), .Y(n292) );
  MUX21X1_HVT U311 ( .A1(n562), .A2(n386), .S0(n283), .Y(n380) );
  MUX21X1_HVT U312 ( .A1(n295), .A2(n291), .S0(n241), .Y(n583) );
  MUX21X1_HVT U313 ( .A1(n339), .A2(n562), .S0(n279), .Y(n462) );
  MUX21X1_HVT U314 ( .A1(n298), .A2(n503), .S0(n275), .Y(n502) );
  MUX21X1_HVT U315 ( .A1(n291), .A2(n289), .S0(n285), .Y(n503) );
  NBUFFX2_HVT U316 ( .A(n591), .Y(n300) );
  NBUFFX2_HVT U317 ( .A(n582), .Y(n293) );
  NBUFFX2_HVT U318 ( .A(n591), .Y(n299) );
  XNOR2X1_HVT U319 ( .A1(n315), .A2(n305), .Y(n275) );
  AND2X1_HVT U320 ( .A1(n371), .A2(n48), .Y(n276) );
  MUX21X1_HVT U321 ( .A1(n398), .A2(n397), .S0(n280), .Y(n396) );
  MUX21X1_HVT U322 ( .A1(n472), .A2(n475), .S0(n282), .Y(n471) );
  INVX0_HVT U323 ( .A(in[4]), .Y(n374) );
  MUX21X1_HVT U324 ( .A1(n501), .A2(n502), .S0(n281), .Y(n499) );
  MUX21X1_HVT U325 ( .A1(n369), .A2(n234), .S0(n303), .Y(n560) );
  NAND2X0_HVT U326 ( .A1(n291), .A2(in[4]), .Y(n591) );
  MUX21X1_HVT U327 ( .A1(n234), .A2(n585), .S0(n240), .Y(n384) );
  MUX21X1_HVT U328 ( .A1(n234), .A2(n372), .S0(n304), .Y(n556) );
  MUX21X1_HVT U329 ( .A1(n234), .A2(n370), .S0(n241), .Y(n574) );
  NAND2X0_HVT U330 ( .A1(in[4]), .A2(n286), .Y(n582) );
  MUX21X1_HVT U331 ( .A1(n234), .A2(n292), .S0(n302), .Y(n376) );
  MUX21X1_HVT U332 ( .A1(n300), .A2(n234), .S0(n301), .Y(n564) );
  MUX21X1_HVT U333 ( .A1(n291), .A2(n234), .S0(n278), .Y(n479) );
  MUX21X1_HVT U334 ( .A1(n234), .A2(n299), .S0(n303), .Y(n375) );
  MUX21X1_HVT U335 ( .A1(n371), .A2(n234), .S0(n305), .Y(n562) );
  NBUFFX2_HVT U336 ( .A(in[3]), .Y(n291) );
  INVX0_HVT U337 ( .A(n570), .Y(n317) );
  INVX0_HVT U338 ( .A(n568), .Y(n318) );
  INVX0_HVT U339 ( .A(n559), .Y(n319) );
  INVX0_HVT U340 ( .A(n557), .Y(n320) );
  INVX0_HVT U341 ( .A(n424), .Y(n321) );
  INVX0_HVT U342 ( .A(n387), .Y(n322) );
  INVX0_HVT U343 ( .A(n589), .Y(n323) );
  INVX0_HVT U344 ( .A(n576), .Y(n324) );
  INVX0_HVT U345 ( .A(n588), .Y(n325) );
  INVX0_HVT U346 ( .A(n586), .Y(n326) );
  INVX0_HVT U347 ( .A(n584), .Y(n327) );
  INVX0_HVT U348 ( .A(n583), .Y(n328) );
  INVX0_HVT U349 ( .A(n581), .Y(n329) );
  INVX0_HVT U350 ( .A(n580), .Y(n330) );
  INVX0_HVT U351 ( .A(n577), .Y(n331) );
  INVX0_HVT U352 ( .A(n575), .Y(n332) );
  INVX0_HVT U353 ( .A(n574), .Y(n333) );
  INVX0_HVT U354 ( .A(n573), .Y(n334) );
  INVX0_HVT U355 ( .A(n572), .Y(n335) );
  INVX0_HVT U356 ( .A(n566), .Y(n338) );
  INVX0_HVT U357 ( .A(n564), .Y(n339) );
  INVX0_HVT U358 ( .A(n563), .Y(n340) );
  INVX0_HVT U359 ( .A(n562), .Y(n341) );
  INVX0_HVT U360 ( .A(n380), .Y(n342) );
  INVX0_HVT U361 ( .A(n561), .Y(n343) );
  INVX0_HVT U362 ( .A(n560), .Y(n344) );
  INVX0_HVT U363 ( .A(n558), .Y(n345) );
  INVX0_HVT U364 ( .A(n556), .Y(n346) );
  INVX0_HVT U365 ( .A(n555), .Y(n347) );
  INVX0_HVT U366 ( .A(n553), .Y(n349) );
  INVX0_HVT U367 ( .A(n550), .Y(n351) );
  INVX0_HVT U368 ( .A(n521), .Y(n352) );
  INVX0_HVT U369 ( .A(n481), .Y(n353) );
  INVX0_HVT U370 ( .A(n386), .Y(n354) );
  INVX0_HVT U371 ( .A(n537), .Y(n355) );
  INVX0_HVT U372 ( .A(n440), .Y(n356) );
  INVX0_HVT U373 ( .A(n385), .Y(n357) );
  INVX0_HVT U374 ( .A(n384), .Y(n358) );
  INVX0_HVT U375 ( .A(n382), .Y(n360) );
  INVX0_HVT U376 ( .A(n381), .Y(n361) );
  INVX0_HVT U377 ( .A(n500), .Y(n362) );
  INVX0_HVT U378 ( .A(n490), .Y(n363) );
  INVX0_HVT U379 ( .A(n378), .Y(n365) );
  INVX0_HVT U380 ( .A(n377), .Y(n366) );
  INVX0_HVT U381 ( .A(n376), .Y(n367) );
  INVX0_HVT U382 ( .A(n375), .Y(n368) );
endmodule

