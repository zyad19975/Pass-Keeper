
module inv_sbox_7 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n18, n103, n196, n197, n198, n199, n200, n201, n202, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640;

  NAND2X0_HVT U1 ( .A1(n313), .A2(n341), .Y(n640) );
  NAND2X0_HVT U3 ( .A1(n313), .A2(in[6]), .Y(n638) );
  NAND2X0_HVT U4 ( .A1(n259), .A2(n354), .Y(n637) );
  NAND2X0_HVT U5 ( .A1(n637), .A2(n351), .Y(n636) );
  NAND2X0_HVT U7 ( .A1(n361), .A2(n352), .Y(n633) );
  NAND2X0_HVT U8 ( .A1(n360), .A2(n350), .Y(n632) );
  NAND2X0_HVT U9 ( .A1(n356), .A2(n632), .Y(n631) );
  NAND2X0_HVT U10 ( .A1(n356), .A2(n629), .Y(n630) );
  NAND2X0_HVT U11 ( .A1(n362), .A2(n354), .Y(n628) );
  NAND2X0_HVT U12 ( .A1(n359), .A2(n338), .Y(n627) );
  NAND2X0_HVT U13 ( .A1(n242), .A2(n632), .Y(n626) );
  NAND2X0_HVT U15 ( .A1(n348), .A2(n361), .Y(n624) );
  NAND2X0_HVT U19 ( .A1(n359), .A2(n430), .Y(n620) );
  NAND2X0_HVT U32 ( .A1(n341), .A2(n362), .Y(n608) );
  NAND2X0_HVT U35 ( .A1(n632), .A2(n431), .Y(n605) );
  NAND2X0_HVT U38 ( .A1(n339), .A2(n281), .Y(n602) );
  NAND2X0_HVT U42 ( .A1(n634), .A2(n431), .Y(n598) );
  OA21X1_HVT U53 ( .A1(n303), .A2(n590), .A3(n397), .Y(n588) );
  NAND2X0_HVT U55 ( .A1(n242), .A2(n637), .Y(n586) );
  AO21X1_HVT U60 ( .A1(n580), .A2(n335), .A3(n619), .Y(n581) );
  NAND2X0_HVT U66 ( .A1(n360), .A2(n324), .Y(n574) );
  MUX41X1_HVT U67 ( .A1(n384), .A3(n411), .A2(n386), .A4(n574), .S0(n337), 
        .S1(n328), .Y(n573) );
  MUX41X1_HVT U68 ( .A1(n384), .A3(n313), .A2(n385), .A4(n356), .S0(n330), 
        .S1(n368), .Y(n572) );
  MUX41X1_HVT U71 ( .A1(n282), .A3(n255), .A2(n628), .A4(n380), .S0(n330), 
        .S1(n245), .Y(n570) );
  NAND2X0_HVT U72 ( .A1(n349), .A2(n286), .Y(n569) );
  MUX41X1_HVT U73 ( .A1(n613), .A3(n569), .A2(n412), .A4(n338), .S0(n336), 
        .S1(n327), .Y(n568) );
  MUX41X1_HVT U74 ( .A1(n630), .A3(n402), .A2(n401), .A4(n390), .S0(n331), 
        .S1(n368), .Y(n567) );
  OA21X1_HVT U76 ( .A1(n373), .A2(n303), .A3(n619), .Y(n565) );
  MUX41X1_HVT U79 ( .A1(n398), .A3(n622), .A2(n400), .A4(n623), .S0(n331), 
        .S1(n245), .Y(n562) );
  MUX41X1_HVT U80 ( .A1(n414), .A3(n410), .A2(n631), .A4(n636), .S0(n330), 
        .S1(n245), .Y(n561) );
  NAND2X0_HVT U81 ( .A1(n229), .A2(n633), .Y(n560) );
  AND2X1_HVT U82 ( .A1(n282), .A2(n353), .Y(n559) );
  MUX41X1_HVT U83 ( .A1(n559), .A3(n399), .A2(n415), .A4(n560), .S0(n330), 
        .S1(n245), .Y(n558) );
  MUX41X1_HVT U87 ( .A1(n374), .A3(n322), .A2(n417), .A4(n395), .S0(n329), 
        .S1(n368), .Y(n555) );
  NAND2X0_HVT U89 ( .A1(n281), .A2(n427), .Y(n553) );
  MUX41X1_HVT U90 ( .A1(n255), .A3(n286), .A2(n593), .A4(n553), .S0(n330), 
        .S1(n245), .Y(n552) );
  MUX41X1_HVT U95 ( .A1(n548), .A3(n554), .A2(n552), .A4(n555), .S0(n347), 
        .S1(n344), .Y(n547) );
  MUX41X1_HVT U99 ( .A1(n608), .A3(n388), .A2(n592), .A4(n349), .S0(n336), 
        .S1(n328), .Y(n543) );
  NAND2X0_HVT U100 ( .A1(n281), .A2(n198), .Y(n542) );
  MUX41X1_HVT U101 ( .A1(n420), .A3(n627), .A2(n298), .A4(n542), .S0(n335), 
        .S1(n326), .Y(n541) );
  MUX41X1_HVT U108 ( .A1(n390), .A3(n348), .A2(n395), .A4(n200), .S0(n331), 
        .S1(n367), .Y(n536) );
  MUX41X1_HVT U109 ( .A1(n419), .A3(n371), .A2(n416), .A4(n408), .S0(n330), 
        .S1(n367), .Y(n535) );
  AO21X1_HVT U112 ( .A1(n405), .A2(n336), .A3(n616), .Y(n532) );
  NAND2X0_HVT U114 ( .A1(n356), .A2(n286), .Y(n530) );
  MUX41X1_HVT U115 ( .A1(n530), .A3(n628), .A2(n405), .A4(n353), .S0(n366), 
        .S1(n328), .Y(n529) );
  MUX41X1_HVT U116 ( .A1(n404), .A3(n398), .A2(n371), .A4(n624), .S0(n329), 
        .S1(n367), .Y(n528) );
  NAND2X0_HVT U118 ( .A1(n281), .A2(n313), .Y(n526) );
  MUX41X1_HVT U119 ( .A1(n422), .A3(n527), .A2(n603), .A4(n526), .S0(n329), 
        .S1(n367), .Y(n525) );
  MUX41X1_HVT U120 ( .A1(n525), .A3(n529), .A2(n528), .A4(n531), .S0(n347), 
        .S1(n345), .Y(n524) );
  MUX41X1_HVT U122 ( .A1(n409), .A3(n318), .A2(n594), .A4(n413), .S0(n329), 
        .S1(n367), .Y(n523) );
  MUX41X1_HVT U124 ( .A1(n320), .A3(n522), .A2(n617), .A4(n392), .S0(n335), 
        .S1(n329), .Y(n521) );
  AOI21X1_HVT U127 ( .A1(n334), .A2(n517), .A3(n378), .Y(n518) );
  NAND2X0_HVT U129 ( .A1(n333), .A2(n356), .Y(n515) );
  MUX41X1_HVT U130 ( .A1(n515), .A3(n516), .A2(n519), .A4(n518), .S0(n337), 
        .S1(n345), .Y(n514) );
  AND2X1_HVT U131 ( .A1(n324), .A2(n281), .Y(n513) );
  MUX41X1_HVT U132 ( .A1(n375), .A3(n513), .A2(n424), .A4(n384), .S0(n336), 
        .S1(n327), .Y(n512) );
  MUX41X1_HVT U133 ( .A1(n425), .A3(n377), .A2(n294), .A4(n376), .S0(n335), 
        .S1(n326), .Y(n511) );
  MUX41X1_HVT U136 ( .A1(n591), .A3(n542), .A2(n509), .A4(n382), .S0(n333), 
        .S1(n367), .Y(n508) );
  MUX41X1_HVT U137 ( .A1(n632), .A3(n611), .A2(n615), .A4(n418), .S0(n337), 
        .S1(n326), .Y(n507) );
  MUX41X1_HVT U139 ( .A1(n506), .A3(n510), .A2(n514), .A4(n520), .S0(n347), 
        .S1(n310), .Y(out[4]) );
  MUX41X1_HVT U140 ( .A1(n401), .A3(n319), .A2(n394), .A4(n628), .S0(n336), 
        .S1(n328), .Y(n505) );
  NAND2X0_HVT U141 ( .A1(n348), .A2(n281), .Y(n504) );
  MUX41X1_HVT U143 ( .A1(n427), .A3(n406), .A2(n620), .A4(n617), .S0(n332), 
        .S1(n302), .Y(n502) );
  MUX41X1_HVT U145 ( .A1(n609), .A3(n421), .A2(n501), .A4(n560), .S0(n334), 
        .S1(n302), .Y(n500) );
  MUX41X1_HVT U146 ( .A1(n500), .A3(n502), .A2(n503), .A4(n505), .S0(n344), 
        .S1(n347), .Y(n499) );
  MUX41X1_HVT U151 ( .A1(n415), .A3(n403), .A2(n391), .A4(n495), .S0(n335), 
        .S1(n326), .Y(n494) );
  MUX41X1_HVT U155 ( .A1(n394), .A3(n628), .A2(n621), .A4(n275), .S0(n332), 
        .S1(n302), .Y(n490) );
  MUX41X1_HVT U156 ( .A1(n490), .A3(n494), .A2(n491), .A4(n496), .S0(in[5]), 
        .S1(n345), .Y(n489) );
  NAND2X0_HVT U159 ( .A1(n486), .A2(n485), .Y(n487) );
  MUX41X1_HVT U162 ( .A1(n314), .A3(n389), .A2(n605), .A4(n483), .S0(n332), 
        .S1(n366), .Y(n482) );
  NAND2X0_HVT U163 ( .A1(n259), .A2(n427), .Y(n481) );
  MUX41X1_HVT U164 ( .A1(n631), .A3(n481), .A2(n603), .A4(n390), .S0(n329), 
        .S1(n302), .Y(n480) );
  NAND2X0_HVT U166 ( .A1(n629), .A2(n477), .Y(n478) );
  MUX41X1_HVT U170 ( .A1(n321), .A3(n317), .A2(n320), .A4(n474), .S0(n332), 
        .S1(n366), .Y(n473) );
  MUX41X1_HVT U173 ( .A1(n356), .A3(n255), .A2(n200), .A4(n604), .S0(n332), 
        .S1(n366), .Y(n470) );
  MUX41X1_HVT U174 ( .A1(n417), .A3(n586), .A2(n425), .A4(n431), .S0(n332), 
        .S1(n302), .Y(n469) );
  NAND2X0_HVT U177 ( .A1(n360), .A2(n313), .Y(n467) );
  MUX41X1_HVT U178 ( .A1(n321), .A3(n467), .A2(n255), .A4(n596), .S0(n332), 
        .S1(n366), .Y(n466) );
  AND2X1_HVT U179 ( .A1(n282), .A2(n351), .Y(n465) );
  MUX41X1_HVT U183 ( .A1(n406), .A3(n254), .A2(n390), .A4(n598), .S0(n335), 
        .S1(n327), .Y(n461) );
  AND2X1_HVT U185 ( .A1(n431), .A2(n362), .Y(n459) );
  OA21X1_HVT U189 ( .A1(n398), .A2(n289), .A3(n580), .Y(n455) );
  MUX41X1_HVT U190 ( .A1(n456), .A3(n457), .A2(n455), .A4(n458), .S0(n344), 
        .S1(n327), .Y(n454) );
  NAND2X0_HVT U191 ( .A1(n289), .A2(n383), .Y(n453) );
  AND2X1_HVT U192 ( .A1(n451), .A2(n402), .Y(n452) );
  NAND2X0_HVT U194 ( .A1(n288), .A2(n451), .Y(n449) );
  MUX41X1_HVT U195 ( .A1(n450), .A3(n449), .A2(n452), .A4(n453), .S0(n330), 
        .S1(n344), .Y(n448) );
  NAND2X0_HVT U198 ( .A1(n361), .A2(n431), .Y(n629) );
  NAND2X0_HVT U200 ( .A1(n351), .A2(n281), .Y(n517) );
  NAND2X0_HVT U207 ( .A1(n281), .A2(n255), .Y(n580) );
  MUX21X2_HVT U2 ( .A1(n550), .A2(n549), .S0(n18), .Y(n548) );
  IBUFFX16_HVT U6 ( .A(n333), .Y(n18) );
  MUX41X1_HVT U14 ( .A1(n535), .A3(n536), .A2(n537), .A4(n539), .S0(n345), 
        .S1(in[5]), .Y(n534) );
  MUX41X1_HVT U16 ( .A1(n420), .A3(n538), .A2(n353), .A4(n377), .S0(n367), 
        .S1(n330), .Y(n537) );
  INVX1_HVT U17 ( .A(n343), .Y(n345) );
  INVX0_HVT U18 ( .A(n598), .Y(n377) );
  IBUFFX2_HVT U20 ( .A(n369), .Y(n367) );
  MUX21X1_HVT U21 ( .A1(n597), .A2(n413), .S0(n336), .Y(n488) );
  MUX21X2_HVT U22 ( .A1(n338), .A2(n430), .S0(n258), .Y(n597) );
  MUX21X2_HVT U23 ( .A1(n563), .A2(n556), .S0(n103), .Y(out[1]) );
  IBUFFX16_HVT U24 ( .A(n202), .Y(n103) );
  INVX1_HVT U25 ( .A(n441), .Y(n416) );
  INVX0_HVT U26 ( .A(n335), .Y(n235) );
  INVX0_HVT U27 ( .A(n597), .Y(n406) );
  MUX21X1_HVT U28 ( .A1(n424), .A2(n375), .S0(n335), .Y(n498) );
  AO21X1_HVT U29 ( .A1(n337), .A2(n379), .A3(n198), .Y(n497) );
  XNOR2X2_HVT U30 ( .A1(n340), .A2(n339), .Y(n312) );
  INVX0_HVT U31 ( .A(n339), .Y(n250) );
  INVX1_HVT U33 ( .A(n312), .Y(n431) );
  INVX1_HVT U34 ( .A(n618), .Y(n391) );
  MUX41X1_HVT U36 ( .A1(n460), .A3(n463), .A2(n448), .A4(n454), .S0(in[5]), 
        .S1(n196), .Y(out[7]) );
  IBUFFX16_HVT U37 ( .A(n243), .Y(n196) );
  INVX0_HVT U39 ( .A(n314), .Y(n596) );
  INVX0_HVT U40 ( .A(n444), .Y(n413) );
  MUX41X1_HVT U41 ( .A1(n472), .A3(n553), .A2(n618), .A4(n317), .S0(n197), 
        .S1(n302), .Y(n471) );
  IBUFFX16_HVT U43 ( .A(n332), .Y(n197) );
  MUX41X1_HVT U44 ( .A1(n601), .A3(n394), .A2(n504), .A4(n423), .S0(n367), 
        .S1(n201), .Y(n503) );
  INVX1_HVT U45 ( .A(n435), .Y(n423) );
  IBUFFX2_HVT U46 ( .A(n334), .Y(n201) );
  INVX1_HVT U47 ( .A(n227), .Y(n566) );
  INVX1_HVT U48 ( .A(n200), .Y(n198) );
  INVX0_HVT U49 ( .A(n639), .Y(n199) );
  INVX1_HVT U50 ( .A(n199), .Y(n200) );
  IBUFFX2_HVT U51 ( .A(n200), .Y(n426) );
  NAND2X0_HVT U52 ( .A1(n338), .A2(n340), .Y(n639) );
  INVX1_HVT U54 ( .A(n352), .Y(n430) );
  INVX1_HVT U56 ( .A(n337), .Y(n289) );
  MUX21X1_HVT U57 ( .A1(n431), .A2(n426), .S0(n360), .Y(n618) );
  IBUFFX16_HVT U58 ( .A(n311), .Y(n202) );
  MUX41X1_HVT U59 ( .A1(n476), .A3(n482), .A2(n480), .A4(n484), .S0(n347), 
        .S1(n218), .Y(n475) );
  IBUFFX16_HVT U61 ( .A(n343), .Y(n218) );
  INVX1_HVT U62 ( .A(n368), .Y(n226) );
  NAND2X0_HVT U63 ( .A1(n393), .A2(n219), .Y(n220) );
  NAND2X0_HVT U64 ( .A1(n584), .A2(n323), .Y(n221) );
  NAND2X0_HVT U65 ( .A1(n220), .A2(n221), .Y(n583) );
  INVX0_HVT U69 ( .A(n323), .Y(n219) );
  NAND2X0_HVT U70 ( .A1(n342), .A2(n222), .Y(n223) );
  NAND2X0_HVT U75 ( .A1(n349), .A2(n363), .Y(n224) );
  NAND2X0_HVT U77 ( .A1(n223), .A2(n224), .Y(n615) );
  IBUFFX2_HVT U78 ( .A(n363), .Y(n222) );
  DELLN1X2_HVT U84 ( .A(n432), .Y(n342) );
  MUX21X1_HVT U85 ( .A1(n615), .A2(n322), .S0(n336), .Y(n493) );
  MUX41X1_HVT U86 ( .A1(n615), .A3(n416), .A2(n398), .A4(n322), .S0(n225), 
        .S1(n226), .Y(n557) );
  IBUFFX16_HVT U88 ( .A(n331), .Y(n225) );
  MUX21X1_HVT U91 ( .A1(n444), .A2(n608), .S0(n337), .Y(n227) );
  IBUFFX2_HVT U92 ( .A(n617), .Y(n392) );
  MUX41X1_HVT U93 ( .A1(n471), .A3(n473), .A2(n469), .A4(n470), .S0(n344), 
        .S1(n346), .Y(n468) );
  INVX1_HVT U94 ( .A(n346), .Y(n347) );
  MUX21X1_HVT U96 ( .A1(n313), .A2(n426), .S0(n233), .Y(n617) );
  MUX21X2_HVT U97 ( .A1(n492), .A2(n493), .S0(n334), .Y(n491) );
  MUX21X2_HVT U98 ( .A1(n566), .A2(n565), .S0(n334), .Y(n564) );
  IBUFFX2_HVT U102 ( .A(n638), .Y(n241) );
  INVX0_HVT U103 ( .A(n615), .Y(n394) );
  NBUFFX2_HVT U104 ( .A(n428), .Y(n339) );
  MUX21X2_HVT U105 ( .A1(n478), .A2(n479), .S0(n333), .Y(n476) );
  MUX21X2_HVT U106 ( .A1(n429), .A2(n342), .S0(n360), .Y(n472) );
  AO21X1_HVT U107 ( .A1(n281), .A2(n356), .A3(n308), .Y(n485) );
  INVX1_HVT U110 ( .A(n369), .Y(n309) );
  INVX0_HVT U111 ( .A(n361), .Y(n233) );
  INVX0_HVT U113 ( .A(n361), .Y(n256) );
  INVX1_HVT U117 ( .A(n363), .Y(n361) );
  IBUFFX2_HVT U121 ( .A(n640), .Y(n255) );
  NBUFFX4_HVT U123 ( .A(n432), .Y(n340) );
  INVX0_HVT U125 ( .A(n354), .Y(n228) );
  INVX1_HVT U126 ( .A(n228), .Y(n229) );
  INVX1_HVT U128 ( .A(n374), .Y(n292) );
  NBUFFX16_HVT U134 ( .A(n309), .Y(n337) );
  NAND2X0_HVT U135 ( .A1(n581), .A2(n230), .Y(n231) );
  NAND2X0_HVT U138 ( .A1(n582), .A2(n279), .Y(n232) );
  NAND2X0_HVT U142 ( .A1(n231), .A2(n232), .Y(n579) );
  INVX0_HVT U144 ( .A(n279), .Y(n230) );
  MUX21X1_HVT U147 ( .A1(n586), .A2(n392), .S0(n303), .Y(n582) );
  IBUFFX2_HVT U148 ( .A(n333), .Y(n279) );
  INVX1_HVT U149 ( .A(in[6]), .Y(n432) );
  INVX1_HVT U150 ( .A(n432), .Y(n324) );
  MUX21X2_HVT U152 ( .A1(n461), .A2(n462), .S0(n234), .Y(n460) );
  IBUFFX16_HVT U153 ( .A(n343), .Y(n234) );
  NAND2X0_HVT U154 ( .A1(n459), .A2(n235), .Y(n236) );
  NAND2X0_HVT U157 ( .A1(n414), .A2(n335), .Y(n237) );
  NAND2X0_HVT U158 ( .A1(n236), .A2(n237), .Y(n458) );
  NAND2X0_HVT U160 ( .A1(n338), .A2(n238), .Y(n239) );
  NAND2X0_HVT U161 ( .A1(n354), .A2(n357), .Y(n240) );
  NAND2X0_HVT U165 ( .A1(n239), .A2(n240), .Y(n443) );
  IBUFFX2_HVT U167 ( .A(n357), .Y(n238) );
  INVX1_HVT U168 ( .A(n363), .Y(n357) );
  INVX0_HVT U169 ( .A(n443), .Y(n414) );
  INVX1_HVT U171 ( .A(n241), .Y(n242) );
  IBUFFX16_HVT U172 ( .A(n311), .Y(n243) );
  MUX41X1_HVT U175 ( .A1(n579), .A3(n585), .A2(n583), .A4(n587), .S0(n347), 
        .S1(n244), .Y(n578) );
  IBUFFX16_HVT U176 ( .A(n343), .Y(n244) );
  MUX21X2_HVT U180 ( .A1(n350), .A2(n352), .S0(n360), .Y(n483) );
  NBUFFX2_HVT U181 ( .A(n368), .Y(n245) );
  IBUFFX2_HVT U182 ( .A(n369), .Y(n368) );
  IBUFFX2_HVT U184 ( .A(n343), .Y(n249) );
  MUX41X1_HVT U186 ( .A1(n570), .A3(n567), .A2(n568), .A4(n564), .S0(n346), 
        .S1(n343), .Y(n563) );
  NAND2X0_HVT U187 ( .A1(n524), .A2(n246), .Y(n247) );
  NAND2X0_HVT U188 ( .A1(n534), .A2(n310), .Y(n248) );
  NAND2X0_HVT U193 ( .A1(n247), .A2(n248), .Y(out[3]) );
  IBUFFX2_HVT U196 ( .A(n310), .Y(n246) );
  MUX41X1_HVT U197 ( .A1(n575), .A3(n572), .A2(n576), .A4(n573), .S0(n346), 
        .S1(n249), .Y(n571) );
  AO21X1_HVT U199 ( .A1(n361), .A2(n198), .A3(n303), .Y(n451) );
  INVX1_HVT U201 ( .A(n311), .Y(n310) );
  OR2X1_HVT U202 ( .A1(n432), .A2(n250), .Y(n635) );
  INVX2_HVT U203 ( .A(n350), .Y(n427) );
  MUX41X1_HVT U204 ( .A1(n411), .A3(n275), .A2(n626), .A4(n418), .S0(n367), 
        .S1(n331), .Y(n546) );
  NAND2X0_HVT U205 ( .A1(n547), .A2(n251), .Y(n252) );
  NAND2X0_HVT U206 ( .A1(n540), .A2(n311), .Y(n253) );
  NAND2X0_HVT U208 ( .A1(n252), .A2(n253), .Y(out[2]) );
  IBUFFX2_HVT U209 ( .A(n311), .Y(n251) );
  MUX21X2_HVT U210 ( .A1(n380), .A2(n348), .S0(n337), .Y(n549) );
  NAND2X0_HVT U211 ( .A1(n571), .A2(n269), .Y(n270) );
  IBUFFX2_HVT U212 ( .A(n344), .Y(n285) );
  IBUFFX2_HVT U213 ( .A(n632), .Y(n379) );
  INVX0_HVT U214 ( .A(n447), .Y(n254) );
  INVX0_HVT U215 ( .A(n447), .Y(n410) );
  INVX0_HVT U216 ( .A(n355), .Y(n429) );
  MUX21X2_HVT U217 ( .A1(n532), .A2(n533), .S0(n334), .Y(n531) );
  INVX2_HVT U218 ( .A(n428), .Y(n313) );
  MUX21X1_HVT U219 ( .A1(n427), .A2(n429), .S0(n256), .Y(n612) );
  MUX41X1_HVT U220 ( .A1(n612), .A3(n403), .A2(n419), .A4(n545), .S0(n257), 
        .S1(n369), .Y(n544) );
  IBUFFX16_HVT U221 ( .A(n331), .Y(n257) );
  IBUFFX2_HVT U222 ( .A(n612), .Y(n397) );
  INVX2_HVT U223 ( .A(in[4]), .Y(n369) );
  MUX21X1_HVT U224 ( .A1(n521), .A2(n523), .S0(n344), .Y(n520) );
  INVX1_HVT U225 ( .A(n363), .Y(n258) );
  INVX1_HVT U226 ( .A(n363), .Y(n259) );
  INVX0_HVT U227 ( .A(n634), .Y(n376) );
  NAND2X0_HVT U228 ( .A1(n487), .A2(n260), .Y(n261) );
  NAND2X0_HVT U229 ( .A1(n488), .A2(n334), .Y(n262) );
  NAND2X0_HVT U230 ( .A1(n261), .A2(n262), .Y(n484) );
  IBUFFX2_HVT U231 ( .A(n334), .Y(n260) );
  INVX1_HVT U232 ( .A(n442), .Y(n415) );
  NAND2X0_HVT U233 ( .A1(n412), .A2(n263), .Y(n264) );
  NAND2X0_HVT U234 ( .A1(n599), .A2(n336), .Y(n265) );
  NAND2X0_HVT U235 ( .A1(n264), .A2(n265), .Y(n456) );
  IBUFFX2_HVT U236 ( .A(n336), .Y(n263) );
  NAND2X0_HVT U237 ( .A1(n588), .A2(n266), .Y(n267) );
  NAND2X0_HVT U238 ( .A1(n589), .A2(n287), .Y(n268) );
  NAND2X0_HVT U239 ( .A1(n267), .A2(n268), .Y(n587) );
  INVX0_HVT U240 ( .A(n287), .Y(n266) );
  NAND2X0_HVT U241 ( .A1(n578), .A2(n310), .Y(n271) );
  NAND2X0_HVT U242 ( .A1(n270), .A2(n271), .Y(out[0]) );
  IBUFFX2_HVT U243 ( .A(n310), .Y(n269) );
  MUX21X1_HVT U244 ( .A1(n385), .A2(n396), .S0(n289), .Y(n589) );
  IBUFFX2_HVT U245 ( .A(n333), .Y(n287) );
  NAND2X0_HVT U246 ( .A1(n489), .A2(n272), .Y(n273) );
  NAND2X0_HVT U247 ( .A1(n499), .A2(n310), .Y(n274) );
  NAND2X0_HVT U248 ( .A1(n273), .A2(n274), .Y(out[5]) );
  IBUFFX2_HVT U249 ( .A(n310), .Y(n272) );
  INVX0_HVT U250 ( .A(n613), .Y(n275) );
  INVX0_HVT U251 ( .A(n613), .Y(n396) );
  NAND2X0_HVT U252 ( .A1(n378), .A2(n289), .Y(n277) );
  NAND2X0_HVT U253 ( .A1(n599), .A2(n337), .Y(n278) );
  NAND2X0_HVT U254 ( .A1(n277), .A2(n278), .Y(n533) );
  IBUFFX2_HVT U255 ( .A(n337), .Y(n276) );
  IBUFFX16_HVT U256 ( .A(n363), .Y(n359) );
  INVX0_HVT U257 ( .A(n362), .Y(n280) );
  INVX1_HVT U258 ( .A(n280), .Y(n281) );
  INVX1_HVT U259 ( .A(n376), .Y(n282) );
  MUX41X1_HVT U260 ( .A1(n415), .A3(n292), .A2(n374), .A4(n377), .S0(n283), 
        .S1(n284), .Y(n462) );
  IBUFFX16_HVT U261 ( .A(n366), .Y(n283) );
  IBUFFX16_HVT U262 ( .A(n329), .Y(n284) );
  NAND2X0_HVT U263 ( .A1(n357), .A2(n355), .Y(n634) );
  MUX41X1_HVT U264 ( .A1(n562), .A3(n558), .A2(n561), .A4(n557), .S0(n346), 
        .S1(n285), .Y(n556) );
  INVX1_HVT U265 ( .A(n378), .Y(n286) );
  IBUFFX2_HVT U266 ( .A(n377), .Y(n288) );
  MUX21X1_HVT U267 ( .A1(n339), .A2(n348), .S0(n362), .Y(n619) );
  INVX1_HVT U268 ( .A(n363), .Y(n360) );
  OA21X1_HVT U269 ( .A1(n372), .A2(n276), .A3(n381), .Y(n492) );
  INVX1_HVT U270 ( .A(n308), .Y(n302) );
  INVX0_HVT U271 ( .A(n340), .Y(n299) );
  INVX0_HVT U272 ( .A(n304), .Y(n539) );
  INVX0_HVT U273 ( .A(n595), .Y(n407) );
  INVX1_HVT U274 ( .A(n308), .Y(n366) );
  NBUFFX2_HVT U275 ( .A(n309), .Y(n336) );
  INVX0_HVT U276 ( .A(n309), .Y(n308) );
  INVX1_HVT U277 ( .A(n333), .Y(n295) );
  INVX1_HVT U278 ( .A(in[5]), .Y(n346) );
  INVX1_HVT U279 ( .A(in[1]), .Y(n343) );
  IBUFFX2_HVT U280 ( .A(n363), .Y(n358) );
  MUX41X1_HVT U281 ( .A1(n594), .A3(n610), .A2(n371), .A4(n386), .S0(n295), 
        .S1(n369), .Y(n554) );
  NAND2X0_HVT U282 ( .A1(n322), .A2(n289), .Y(n290) );
  NAND2X0_HVT U283 ( .A1(n592), .A2(n337), .Y(n291) );
  NAND2X0_HVT U284 ( .A1(n290), .A2(n291), .Y(n457) );
  INVX0_HVT U285 ( .A(n298), .Y(n604) );
  INVX0_HVT U286 ( .A(n637), .Y(n374) );
  INVX0_HVT U287 ( .A(n560), .Y(n306) );
  INVX0_HVT U288 ( .A(n614), .Y(n395) );
  INVX0_HVT U289 ( .A(n625), .Y(n384) );
  INVX1_HVT U290 ( .A(n625), .Y(n305) );
  INVX1_HVT U291 ( .A(n619), .Y(n390) );
  INVX0_HVT U292 ( .A(n586), .Y(n293) );
  INVX0_HVT U293 ( .A(n293), .Y(n294) );
  MUX21X2_HVT U294 ( .A1(n497), .A2(n498), .S0(n295), .Y(n496) );
  NAND2X0_HVT U295 ( .A1(n466), .A2(n345), .Y(n296) );
  NAND2X0_HVT U296 ( .A1(n464), .A2(n343), .Y(n297) );
  NAND2X0_HVT U297 ( .A1(n296), .A2(n297), .Y(n463) );
  AO21X1_HVT U298 ( .A1(n349), .A2(n292), .A3(n276), .Y(n477) );
  MUX21X1_HVT U299 ( .A1(n299), .A2(n312), .S0(n358), .Y(n298) );
  NAND2X0_HVT U300 ( .A1(n348), .A2(n308), .Y(n300) );
  NAND2X0_HVT U301 ( .A1(n342), .A2(n336), .Y(n301) );
  NAND2X0_HVT U302 ( .A1(n300), .A2(n301), .Y(n551) );
  INVX0_HVT U303 ( .A(n337), .Y(n303) );
  MUX21X2_HVT U304 ( .A1(n468), .A2(n475), .S0(n310), .Y(out[6]) );
  MUX41X1_HVT U305 ( .A1(n307), .A3(n306), .A2(n436), .A4(n305), .S0(n295), 
        .S1(n369), .Y(n304) );
  NAND2X0_HVT U306 ( .A1(n286), .A2(n351), .Y(n307) );
  INVX1_HVT U307 ( .A(in[0]), .Y(n363) );
  IBUFFX2_HVT U308 ( .A(in[0]), .Y(n362) );
  MUX41X1_HVT U309 ( .A1(n294), .A3(n395), .A2(n349), .A4(n410), .S0(n295), 
        .S1(n308), .Y(n585) );
  INVX1_HVT U310 ( .A(in[7]), .Y(n311) );
  MUX21X2_HVT U311 ( .A1(n390), .A2(n577), .S0(n323), .Y(n576) );
  MUX41X1_HVT U312 ( .A1(n546), .A3(n543), .A2(n544), .A4(n541), .S0(n346), 
        .S1(n343), .Y(n540) );
  MUX21X1_HVT U313 ( .A1(n507), .A2(n508), .S0(n344), .Y(n506) );
  MUX41X1_HVT U314 ( .A1(n602), .A3(n388), .A2(n389), .A4(n387), .S0(n295), 
        .S1(n276), .Y(n575) );
  INVX1_HVT U315 ( .A(in[3]), .Y(n428) );
  INVX1_HVT U316 ( .A(n445), .Y(n412) );
  MUX21X1_HVT U317 ( .A1(n355), .A2(n350), .S0(n362), .Y(n314) );
  NBUFFX2_HVT U318 ( .A(n639), .Y(n354) );
  INVX1_HVT U319 ( .A(n434), .Y(n424) );
  MUX41X1_HVT U320 ( .A1(n595), .A3(n465), .A2(n370), .A4(n608), .S0(n295), 
        .S1(n276), .Y(n464) );
  NAND2X0_HVT U321 ( .A1(n614), .A2(n308), .Y(n315) );
  NAND2X0_HVT U322 ( .A1(n335), .A2(n617), .Y(n316) );
  NAND2X0_HVT U323 ( .A1(n316), .A2(n315), .Y(n479) );
  MUX21X2_HVT U324 ( .A1(n511), .A2(n512), .S0(n345), .Y(n510) );
  NBUFFX2_HVT U325 ( .A(n635), .Y(n350) );
  NBUFFX2_HVT U326 ( .A(n635), .Y(n351) );
  AND2X1_HVT U327 ( .A1(n634), .A2(n229), .Y(n317) );
  MUX21X1_HVT U328 ( .A1(n407), .A2(n320), .S0(n335), .Y(n450) );
  AND2X1_HVT U329 ( .A1(n229), .A2(n624), .Y(n318) );
  MUX21X1_HVT U330 ( .A1(n341), .A2(n426), .S0(n359), .Y(n614) );
  MUX21X1_HVT U331 ( .A1(n429), .A2(n349), .S0(n258), .Y(n440) );
  MUX21X1_HVT U332 ( .A1(n426), .A2(n341), .S0(n361), .Y(n445) );
  MUX21X1_HVT U333 ( .A1(n431), .A2(n339), .S0(n359), .Y(n601) );
  MUX21X1_HVT U334 ( .A1(n426), .A2(n431), .S0(n359), .Y(n607) );
  MUX21X1_HVT U335 ( .A1(n391), .A2(n292), .S0(n333), .Y(n577) );
  MUX21X1_HVT U336 ( .A1(n394), .A2(n636), .S0(n334), .Y(n584) );
  MUX21X1_HVT U337 ( .A1(n340), .A2(n427), .S0(n357), .Y(n495) );
  XOR2X1_HVT U338 ( .A1(n349), .A2(n358), .Y(n594) );
  MUX21X1_HVT U339 ( .A1(n338), .A2(n431), .S0(n259), .Y(n442) );
  MUX21X1_HVT U340 ( .A1(n430), .A2(n338), .S0(n360), .Y(n444) );
  MUX21X1_HVT U341 ( .A1(n340), .A2(n349), .S0(n357), .Y(n600) );
  MUX21X1_HVT U342 ( .A1(n339), .A2(n426), .S0(n359), .Y(n610) );
  MUX21X1_HVT U343 ( .A1(n551), .A2(n353), .S0(n359), .Y(n550) );
  MUX21X1_HVT U344 ( .A1(n198), .A2(n430), .S0(n360), .Y(n590) );
  MUX21X1_HVT U345 ( .A1(n340), .A2(n229), .S0(n358), .Y(n538) );
  XOR2X1_HVT U346 ( .A1(n353), .A2(n259), .Y(n593) );
  XOR2X1_HVT U347 ( .A1(n350), .A2(n358), .Y(n592) );
  MUX21X1_HVT U348 ( .A1(n349), .A2(n427), .S0(n358), .Y(n606) );
  MUX21X1_HVT U349 ( .A1(n351), .A2(n354), .S0(n357), .Y(n434) );
  MUX21X1_HVT U350 ( .A1(n431), .A2(n342), .S0(n358), .Y(n435) );
  MUX21X1_HVT U351 ( .A1(n348), .A2(n255), .S0(n258), .Y(n609) );
  MUX21X1_HVT U352 ( .A1(n607), .A2(n318), .S0(n334), .Y(n516) );
  MUX21X1_HVT U353 ( .A1(n200), .A2(n351), .S0(n361), .Y(n501) );
  MUX21X1_HVT U354 ( .A1(n423), .A2(n319), .S0(n333), .Y(n519) );
  MUX21X1_HVT U355 ( .A1(n356), .A2(n229), .S0(n358), .Y(n625) );
  MUX21X1_HVT U356 ( .A1(n352), .A2(n229), .S0(n259), .Y(n622) );
  MUX21X1_HVT U357 ( .A1(n339), .A2(n341), .S0(n259), .Y(n595) );
  XOR2X1_HVT U358 ( .A1(n355), .A2(n360), .Y(n603) );
  XNOR2X1_HVT U359 ( .A1(n200), .A2(n258), .Y(n319) );
  MUX21X1_HVT U360 ( .A1(n353), .A2(n339), .S0(n358), .Y(n621) );
  MUX21X1_HVT U361 ( .A1(n338), .A2(n353), .S0(n259), .Y(n437) );
  MUX21X1_HVT U362 ( .A1(n353), .A2(n341), .S0(n258), .Y(n522) );
  AND2X1_HVT U363 ( .A1(n359), .A2(n342), .Y(n320) );
  NBUFFX2_HVT U364 ( .A(n309), .Y(n335) );
  NBUFFX2_HVT U365 ( .A(n428), .Y(n338) );
  NBUFFX2_HVT U366 ( .A(n312), .Y(n349) );
  NBUFFX2_HVT U367 ( .A(n312), .Y(n348) );
  AND2X1_HVT U368 ( .A1(n430), .A2(n281), .Y(n321) );
  INVX1_HVT U369 ( .A(n325), .Y(n474) );
  NBUFFX2_HVT U370 ( .A(n638), .Y(n352) );
  AND2X1_HVT U371 ( .A1(n242), .A2(n281), .Y(n322) );
  NBUFFX2_HVT U372 ( .A(n638), .Y(n353) );
  NBUFFX2_HVT U373 ( .A(n365), .Y(n332) );
  NBUFFX2_HVT U374 ( .A(n365), .Y(n334) );
  NBUFFX2_HVT U375 ( .A(n365), .Y(n333) );
  NBUFFX2_HVT U376 ( .A(n432), .Y(n341) );
  XNOR2X1_HVT U377 ( .A1(n308), .A2(n329), .Y(n323) );
  NBUFFX2_HVT U378 ( .A(n364), .Y(n329) );
  NBUFFX2_HVT U379 ( .A(n364), .Y(n331) );
  NBUFFX2_HVT U380 ( .A(n365), .Y(n327) );
  NBUFFX2_HVT U381 ( .A(n364), .Y(n330) );
  NBUFFX2_HVT U382 ( .A(n365), .Y(n328) );
  NBUFFX2_HVT U383 ( .A(n365), .Y(n326) );
  INVX1_HVT U384 ( .A(n343), .Y(n344) );
  MUX21X1_HVT U385 ( .A1(n255), .A2(n313), .S0(n258), .Y(n433) );
  MUX21X1_HVT U386 ( .A1(n430), .A2(n427), .S0(n259), .Y(n527) );
  MUX21X1_HVT U387 ( .A1(n351), .A2(n313), .S0(n359), .Y(n545) );
  MUX21X1_HVT U388 ( .A1(n313), .A2(n351), .S0(n357), .Y(n438) );
  MUX21X1_HVT U389 ( .A1(n356), .A2(n313), .S0(n361), .Y(n486) );
  MUX21X1_HVT U390 ( .A1(n313), .A2(n356), .S0(n359), .Y(n439) );
  MUX21X1_HVT U391 ( .A1(n342), .A2(n313), .S0(n361), .Y(n613) );
  NBUFFX2_HVT U392 ( .A(in[2]), .Y(n365) );
  NBUFFX2_HVT U393 ( .A(in[2]), .Y(n364) );
  MUX21X1_HVT U394 ( .A1(n352), .A2(n355), .S0(n362), .Y(n325) );
  MUX21X1_HVT U395 ( .A1(n198), .A2(n324), .S0(n258), .Y(n509) );
  XOR2X1_HVT U396 ( .A1(n258), .A2(n324), .Y(n591) );
  MUX21X1_HVT U397 ( .A1(n324), .A2(n353), .S0(n360), .Y(n446) );
  MUX21X1_HVT U398 ( .A1(n353), .A2(n324), .S0(n259), .Y(n441) );
  MUX21X1_HVT U399 ( .A1(n338), .A2(n324), .S0(n357), .Y(n436) );
  MUX21X1_HVT U400 ( .A1(n324), .A2(n429), .S0(n259), .Y(n616) );
  MUX21X1_HVT U401 ( .A1(n351), .A2(n324), .S0(n357), .Y(n611) );
  MUX21X1_HVT U402 ( .A1(n324), .A2(n355), .S0(n357), .Y(n623) );
  MUX21X1_HVT U403 ( .A1(n324), .A2(n427), .S0(n258), .Y(n447) );
  MUX21X1_HVT U404 ( .A1(n324), .A2(n430), .S0(n358), .Y(n599) );
  NBUFFX2_HVT U405 ( .A(n640), .Y(n355) );
  NBUFFX2_HVT U406 ( .A(n640), .Y(n356) );
  INVX0_HVT U407 ( .A(n628), .Y(n370) );
  INVX0_HVT U408 ( .A(n602), .Y(n371) );
  INVX0_HVT U409 ( .A(n542), .Y(n372) );
  INVX0_HVT U410 ( .A(n504), .Y(n373) );
  INVX0_HVT U411 ( .A(n636), .Y(n375) );
  INVX0_HVT U412 ( .A(n633), .Y(n378) );
  INVX0_HVT U413 ( .A(n605), .Y(n380) );
  INVX0_HVT U414 ( .A(n626), .Y(n381) );
  INVX0_HVT U415 ( .A(n631), .Y(n382) );
  INVX0_HVT U416 ( .A(n627), .Y(n383) );
  INVX0_HVT U417 ( .A(n624), .Y(n385) );
  INVX0_HVT U418 ( .A(n623), .Y(n386) );
  INVX0_HVT U419 ( .A(n622), .Y(n387) );
  INVX0_HVT U420 ( .A(n621), .Y(n388) );
  INVX0_HVT U421 ( .A(n620), .Y(n389) );
  INVX0_HVT U422 ( .A(n616), .Y(n393) );
  INVX0_HVT U423 ( .A(n611), .Y(n398) );
  INVX0_HVT U424 ( .A(n610), .Y(n399) );
  INVX0_HVT U425 ( .A(n609), .Y(n400) );
  INVX0_HVT U426 ( .A(n607), .Y(n401) );
  INVX0_HVT U427 ( .A(n606), .Y(n402) );
  INVX0_HVT U428 ( .A(n603), .Y(n403) );
  INVX0_HVT U429 ( .A(n601), .Y(n404) );
  INVX0_HVT U430 ( .A(n600), .Y(n405) );
  INVX0_HVT U431 ( .A(n594), .Y(n408) );
  INVX0_HVT U432 ( .A(n630), .Y(n409) );
  INVX0_HVT U433 ( .A(n446), .Y(n411) );
  INVX0_HVT U434 ( .A(n440), .Y(n417) );
  INVX0_HVT U435 ( .A(n439), .Y(n418) );
  INVX0_HVT U436 ( .A(n438), .Y(n419) );
  INVX0_HVT U437 ( .A(n437), .Y(n420) );
  INVX0_HVT U438 ( .A(n436), .Y(n421) );
  INVX0_HVT U439 ( .A(n486), .Y(n422) );
  INVX0_HVT U440 ( .A(n433), .Y(n425) );
endmodule

