
module round ( in, round_num, keyin, keyout, out );
  input [127:0] in;
  input [3:0] round_num;
  input [127:0] keyin;
  output [127:0] keyout;
  output [127:0] out;
  wire   n132, n133, n134, n135, \_0_net_[127] , \_0_net_[126] ,
         \_0_net_[125] , \_0_net_[124] , \_0_net_[123] , \_0_net_[122] ,
         \_0_net_[121] , \_0_net_[120] , \_0_net_[119] , \_0_net_[118] ,
         \_0_net_[117] , \_0_net_[116] , \_0_net_[115] , \_0_net_[114] ,
         \_0_net_[113] , \_0_net_[112] , \_0_net_[111] , \_0_net_[110] ,
         \_0_net_[109] , \_0_net_[108] , \_0_net_[107] , \_0_net_[106] ,
         \_0_net_[105] , \_0_net_[104] , \_0_net_[103] , \_0_net_[102] ,
         \_0_net_[101] , \_0_net_[100] , \_0_net_[99] , \_0_net_[98] ,
         \_0_net_[97] , \_0_net_[96] , \_0_net_[95] , \_0_net_[94] ,
         \_0_net_[93] , \_0_net_[92] , \_0_net_[91] , \_0_net_[90] ,
         \_0_net_[89] , \_0_net_[88] , \_0_net_[87] , \_0_net_[86] ,
         \_0_net_[85] , \_0_net_[84] , \_0_net_[83] , \_0_net_[82] ,
         \_0_net_[81] , \_0_net_[80] , \_0_net_[79] , \_0_net_[78] ,
         \_0_net_[77] , \_0_net_[76] , \_0_net_[75] , \_0_net_[74] ,
         \_0_net_[73] , \_0_net_[72] , \_0_net_[71] , \_0_net_[70] ,
         \_0_net_[69] , \_0_net_[68] , \_0_net_[67] , \_0_net_[66] ,
         \_0_net_[65] , \_0_net_[64] , \_0_net_[63] , \_0_net_[62] ,
         \_0_net_[61] , \_0_net_[60] , \_0_net_[59] , \_0_net_[58] ,
         \_0_net_[57] , \_0_net_[56] , \_0_net_[55] , \_0_net_[54] ,
         \_0_net_[53] , \_0_net_[52] , \_0_net_[51] , \_0_net_[50] ,
         \_0_net_[49] , \_0_net_[48] , \_0_net_[47] , \_0_net_[46] ,
         \_0_net_[45] , \_0_net_[44] , \_0_net_[43] , \_0_net_[42] ,
         \_0_net_[41] , \_0_net_[40] , \_0_net_[39] , \_0_net_[38] ,
         \_0_net_[37] , \_0_net_[36] , \_0_net_[35] , \_0_net_[34] ,
         \_0_net_[33] , \_0_net_[32] , \_0_net_[31] , \_0_net_[30] ,
         \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] ,
         \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] ,
         \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] ,
         \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] ,
         \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] ,
         \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] ,
         \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_0_net_[0] ,
         n2, n3, n1, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131;
  wire   [127:0] sb_out;
  wire   [127:0] sr_out;
  wire   [127:0] mc_out;

  AO22X1_HVT U2 ( .A1(mc_out[9]), .A2(n118), .A3(n4), .A4(n121), .Y(
        \_0_net_[9] ) );
  AO22X1_HVT U4 ( .A1(mc_out[98]), .A2(n118), .A3(n121), .A4(sr_out[98]), .Y(
        \_0_net_[98] ) );
  AO22X1_HVT U6 ( .A1(n117), .A2(mc_out[96]), .A3(n35), .A4(n121), .Y(
        \_0_net_[96] ) );
  AO22X1_HVT U7 ( .A1(mc_out[95]), .A2(n117), .A3(sr_out[95]), .A4(n121), .Y(
        \_0_net_[95] ) );
  AO22X1_HVT U8 ( .A1(mc_out[94]), .A2(n117), .A3(sr_out[94]), .A4(n121), .Y(
        \_0_net_[94] ) );
  AO22X1_HVT U9 ( .A1(mc_out[93]), .A2(n117), .A3(sr_out[93]), .A4(n121), .Y(
        \_0_net_[93] ) );
  AO22X1_HVT U10 ( .A1(mc_out[92]), .A2(n117), .A3(sr_out[92]), .A4(n121), .Y(
        \_0_net_[92] ) );
  AO22X1_HVT U12 ( .A1(mc_out[90]), .A2(n117), .A3(sr_out[90]), .A4(n121), .Y(
        \_0_net_[90] ) );
  AO22X1_HVT U13 ( .A1(n117), .A2(mc_out[8]), .A3(n121), .A4(n21), .Y(
        \_0_net_[8] ) );
  AO22X1_HVT U14 ( .A1(n117), .A2(mc_out[89]), .A3(sr_out[89]), .A4(n122), .Y(
        \_0_net_[89] ) );
  AO22X1_HVT U15 ( .A1(mc_out[88]), .A2(n117), .A3(sr_out[88]), .A4(n122), .Y(
        \_0_net_[88] ) );
  AO22X1_HVT U16 ( .A1(mc_out[87]), .A2(n117), .A3(n19), .A4(n122), .Y(
        \_0_net_[87] ) );
  AO22X1_HVT U17 ( .A1(mc_out[86]), .A2(n117), .A3(sr_out[86]), .A4(n122), .Y(
        \_0_net_[86] ) );
  AO22X1_HVT U21 ( .A1(mc_out[82]), .A2(n116), .A3(sr_out[82]), .A4(n122), .Y(
        \_0_net_[82] ) );
  AO22X1_HVT U22 ( .A1(mc_out[81]), .A2(n116), .A3(sr_out[81]), .A4(n122), .Y(
        \_0_net_[81] ) );
  AO22X1_HVT U23 ( .A1(mc_out[80]), .A2(n116), .A3(sr_out[80]), .A4(n122), .Y(
        \_0_net_[80] ) );
  AO22X1_HVT U24 ( .A1(mc_out[7]), .A2(n116), .A3(n12), .A4(n122), .Y(
        \_0_net_[7] ) );
  AO22X1_HVT U25 ( .A1(mc_out[79]), .A2(n116), .A3(n27), .A4(n122), .Y(
        \_0_net_[79] ) );
  AO22X1_HVT U26 ( .A1(mc_out[78]), .A2(n116), .A3(sr_out[78]), .A4(n123), .Y(
        \_0_net_[78] ) );
  AO22X1_HVT U27 ( .A1(mc_out[77]), .A2(n116), .A3(sr_out[77]), .A4(n123), .Y(
        \_0_net_[77] ) );
  AO22X1_HVT U30 ( .A1(mc_out[74]), .A2(n116), .A3(sr_out[74]), .A4(n123), .Y(
        \_0_net_[74] ) );
  AO22X1_HVT U32 ( .A1(mc_out[72]), .A2(n116), .A3(sr_out[72]), .A4(n123), .Y(
        \_0_net_[72] ) );
  AO22X1_HVT U33 ( .A1(n116), .A2(mc_out[71]), .A3(sr_out[71]), .A4(n123), .Y(
        \_0_net_[71] ) );
  AO22X1_HVT U34 ( .A1(mc_out[70]), .A2(n116), .A3(n123), .A4(sr_out[70]), .Y(
        \_0_net_[70] ) );
  AO22X1_HVT U35 ( .A1(mc_out[6]), .A2(n116), .A3(sr_out[6]), .A4(n123), .Y(
        \_0_net_[6] ) );
  AO22X1_HVT U36 ( .A1(mc_out[69]), .A2(n115), .A3(sr_out[69]), .A4(n123), .Y(
        \_0_net_[69] ) );
  AO22X1_HVT U38 ( .A1(mc_out[67]), .A2(n115), .A3(n13), .A4(n124), .Y(
        \_0_net_[67] ) );
  AO22X1_HVT U40 ( .A1(mc_out[65]), .A2(n115), .A3(sr_out[65]), .A4(n124), .Y(
        \_0_net_[65] ) );
  AO22X1_HVT U41 ( .A1(mc_out[64]), .A2(n115), .A3(sr_out[64]), .A4(n124), .Y(
        \_0_net_[64] ) );
  AO22X1_HVT U42 ( .A1(mc_out[63]), .A2(n115), .A3(sr_out[63]), .A4(n124), .Y(
        \_0_net_[63] ) );
  AO22X1_HVT U43 ( .A1(mc_out[62]), .A2(n115), .A3(sr_out[62]), .A4(n124), .Y(
        \_0_net_[62] ) );
  AO22X1_HVT U46 ( .A1(mc_out[5]), .A2(n115), .A3(sr_out[5]), .A4(n124), .Y(
        \_0_net_[5] ) );
  AO22X1_HVT U47 ( .A1(mc_out[59]), .A2(n115), .A3(sr_out[59]), .A4(n124), .Y(
        \_0_net_[59] ) );
  AO22X1_HVT U48 ( .A1(n115), .A2(mc_out[58]), .A3(sr_out[58]), .A4(n124), .Y(
        \_0_net_[58] ) );
  AO22X1_HVT U50 ( .A1(n115), .A2(mc_out[56]), .A3(sr_out[56]), .A4(n125), .Y(
        \_0_net_[56] ) );
  AO22X1_HVT U51 ( .A1(mc_out[55]), .A2(n114), .A3(n95), .A4(n125), .Y(
        \_0_net_[55] ) );
  AO22X1_HVT U52 ( .A1(mc_out[54]), .A2(n114), .A3(sr_out[54]), .A4(n125), .Y(
        \_0_net_[54] ) );
  AO22X1_HVT U53 ( .A1(mc_out[53]), .A2(n114), .A3(sr_out[53]), .A4(n125), .Y(
        \_0_net_[53] ) );
  AO22X1_HVT U56 ( .A1(mc_out[50]), .A2(n114), .A3(sr_out[50]), .A4(n125), .Y(
        \_0_net_[50] ) );
  AO22X1_HVT U57 ( .A1(mc_out[4]), .A2(n114), .A3(sr_out[4]), .A4(n125), .Y(
        \_0_net_[4] ) );
  AO22X1_HVT U59 ( .A1(mc_out[48]), .A2(n114), .A3(sr_out[48]), .A4(n125), .Y(
        \_0_net_[48] ) );
  AO22X1_HVT U60 ( .A1(mc_out[47]), .A2(n114), .A3(n103), .A4(n125), .Y(
        \_0_net_[47] ) );
  AO22X1_HVT U62 ( .A1(mc_out[45]), .A2(n114), .A3(sr_out[45]), .A4(n126), .Y(
        \_0_net_[45] ) );
  AO22X1_HVT U65 ( .A1(mc_out[42]), .A2(n114), .A3(n10), .A4(n126), .Y(
        \_0_net_[42] ) );
  AO22X1_HVT U66 ( .A1(mc_out[41]), .A2(n113), .A3(sr_out[41]), .A4(n126), .Y(
        \_0_net_[41] ) );
  AO22X1_HVT U67 ( .A1(mc_out[40]), .A2(n113), .A3(sr_out[40]), .A4(n126), .Y(
        \_0_net_[40] ) );
  AO22X1_HVT U68 ( .A1(mc_out[3]), .A2(n113), .A3(sr_out[3]), .A4(n126), .Y(
        \_0_net_[3] ) );
  AO22X1_HVT U69 ( .A1(mc_out[39]), .A2(n113), .A3(n105), .A4(n126), .Y(
        \_0_net_[39] ) );
  AO22X1_HVT U70 ( .A1(mc_out[38]), .A2(n113), .A3(sr_out[38]), .A4(n126), .Y(
        \_0_net_[38] ) );
  AO22X1_HVT U74 ( .A1(mc_out[34]), .A2(n113), .A3(sr_out[34]), .A4(n127), .Y(
        \_0_net_[34] ) );
  AO22X1_HVT U76 ( .A1(mc_out[32]), .A2(n113), .A3(sr_out[32]), .A4(n127), .Y(
        \_0_net_[32] ) );
  AO22X1_HVT U77 ( .A1(mc_out[31]), .A2(n113), .A3(n104), .A4(n127), .Y(
        \_0_net_[31] ) );
  AO22X1_HVT U78 ( .A1(mc_out[30]), .A2(n113), .A3(sr_out[30]), .A4(n127), .Y(
        \_0_net_[30] ) );
  AO22X1_HVT U79 ( .A1(mc_out[2]), .A2(n113), .A3(sr_out[2]), .A4(n127), .Y(
        \_0_net_[2] ) );
  AO22X1_HVT U80 ( .A1(mc_out[29]), .A2(n113), .A3(n127), .A4(sr_out[29]), .Y(
        \_0_net_[29] ) );
  AO22X1_HVT U82 ( .A1(mc_out[27]), .A2(n112), .A3(sr_out[27]), .A4(n127), .Y(
        \_0_net_[27] ) );
  AO22X1_HVT U83 ( .A1(mc_out[26]), .A2(n112), .A3(sr_out[26]), .A4(n127), .Y(
        \_0_net_[26] ) );
  AO22X1_HVT U85 ( .A1(mc_out[24]), .A2(n112), .A3(sr_out[24]), .A4(n127), .Y(
        \_0_net_[24] ) );
  AO22X1_HVT U87 ( .A1(mc_out[22]), .A2(n112), .A3(sr_out[22]), .A4(n128), .Y(
        \_0_net_[22] ) );
  AO22X1_HVT U88 ( .A1(mc_out[21]), .A2(n112), .A3(n16), .A4(n128), .Y(
        \_0_net_[21] ) );
  AO22X1_HVT U91 ( .A1(mc_out[19]), .A2(n112), .A3(sr_out[19]), .A4(n128), .Y(
        \_0_net_[19] ) );
  AO22X1_HVT U92 ( .A1(mc_out[18]), .A2(n112), .A3(n26), .A4(n128), .Y(
        \_0_net_[18] ) );
  AO22X1_HVT U93 ( .A1(mc_out[17]), .A2(n112), .A3(n9), .A4(n128), .Y(
        \_0_net_[17] ) );
  AO22X1_HVT U94 ( .A1(mc_out[16]), .A2(n112), .A3(sr_out[16]), .A4(n128), .Y(
        \_0_net_[16] ) );
  AO22X1_HVT U95 ( .A1(mc_out[15]), .A2(n112), .A3(n94), .A4(n128), .Y(
        \_0_net_[15] ) );
  AO22X1_HVT U96 ( .A1(mc_out[14]), .A2(n111), .A3(n96), .A4(n128), .Y(
        \_0_net_[14] ) );
  AO22X1_HVT U97 ( .A1(mc_out[13]), .A2(n111), .A3(sr_out[13]), .A4(n128), .Y(
        \_0_net_[13] ) );
  AO22X1_HVT U98 ( .A1(mc_out[12]), .A2(n111), .A3(n15), .A4(n129), .Y(
        \_0_net_[12] ) );
  AO22X1_HVT U99 ( .A1(mc_out[127]), .A2(n111), .A3(sr_out[127]), .A4(n129), 
        .Y(\_0_net_[127] ) );
  AO22X1_HVT U100 ( .A1(mc_out[126]), .A2(n111), .A3(sr_out[126]), .A4(n129), 
        .Y(\_0_net_[126] ) );
  AO22X1_HVT U101 ( .A1(n111), .A2(mc_out[125]), .A3(sr_out[125]), .A4(n129), 
        .Y(\_0_net_[125] ) );
  AO22X1_HVT U103 ( .A1(mc_out[123]), .A2(n111), .A3(sr_out[123]), .A4(n129), 
        .Y(\_0_net_[123] ) );
  AO22X1_HVT U104 ( .A1(mc_out[122]), .A2(n111), .A3(sr_out[122]), .A4(n129), 
        .Y(\_0_net_[122] ) );
  AO22X1_HVT U106 ( .A1(mc_out[120]), .A2(n111), .A3(sr_out[120]), .A4(n129), 
        .Y(\_0_net_[120] ) );
  AO22X1_HVT U108 ( .A1(mc_out[119]), .A2(n111), .A3(sr_out[119]), .A4(n129), 
        .Y(\_0_net_[119] ) );
  AO22X1_HVT U109 ( .A1(mc_out[118]), .A2(n111), .A3(sr_out[118]), .A4(n129), 
        .Y(\_0_net_[118] ) );
  AO22X1_HVT U110 ( .A1(mc_out[117]), .A2(n111), .A3(sr_out[117]), .A4(n130), 
        .Y(\_0_net_[117] ) );
  AO22X1_HVT U111 ( .A1(mc_out[116]), .A2(n110), .A3(sr_out[116]), .A4(n130), 
        .Y(\_0_net_[116] ) );
  AO22X1_HVT U113 ( .A1(mc_out[114]), .A2(n110), .A3(n80), .A4(n130), .Y(
        \_0_net_[114] ) );
  AO22X1_HVT U114 ( .A1(n110), .A2(mc_out[113]), .A3(sr_out[113]), .A4(n130), 
        .Y(\_0_net_[113] ) );
  AO22X1_HVT U115 ( .A1(mc_out[112]), .A2(n110), .A3(sr_out[112]), .A4(n130), 
        .Y(\_0_net_[112] ) );
  AO22X1_HVT U116 ( .A1(n110), .A2(mc_out[111]), .A3(n91), .A4(n130), .Y(
        \_0_net_[111] ) );
  AO22X1_HVT U117 ( .A1(mc_out[110]), .A2(n110), .A3(sr_out[110]), .A4(n130), 
        .Y(\_0_net_[110] ) );
  AO22X1_HVT U118 ( .A1(mc_out[10]), .A2(n110), .A3(n1), .A4(n130), .Y(
        \_0_net_[10] ) );
  AO22X1_HVT U119 ( .A1(mc_out[109]), .A2(n110), .A3(sr_out[109]), .A4(n130), 
        .Y(\_0_net_[109] ) );
  AO22X1_HVT U120 ( .A1(mc_out[108]), .A2(n110), .A3(sr_out[108]), .A4(n130), 
        .Y(\_0_net_[108] ) );
  AO22X1_HVT U122 ( .A1(n110), .A2(mc_out[106]), .A3(sr_out[106]), .A4(n131), 
        .Y(\_0_net_[106] ) );
  AO22X1_HVT U123 ( .A1(mc_out[105]), .A2(n110), .A3(sr_out[105]), .A4(n131), 
        .Y(\_0_net_[105] ) );
  AO22X1_HVT U124 ( .A1(mc_out[104]), .A2(n110), .A3(sr_out[104]), .A4(n131), 
        .Y(\_0_net_[104] ) );
  AO22X1_HVT U125 ( .A1(mc_out[103]), .A2(n110), .A3(n107), .A4(n131), .Y(
        \_0_net_[103] ) );
  AO22X1_HVT U126 ( .A1(mc_out[102]), .A2(n109), .A3(sr_out[102]), .A4(n131), 
        .Y(\_0_net_[102] ) );
  AO22X1_HVT U127 ( .A1(mc_out[101]), .A2(n109), .A3(sr_out[101]), .A4(n131), 
        .Y(\_0_net_[101] ) );
  AO22X1_HVT U128 ( .A1(mc_out[100]), .A2(n109), .A3(sr_out[100]), .A4(n131), 
        .Y(\_0_net_[100] ) );
  AO22X1_HVT U129 ( .A1(mc_out[0]), .A2(n108), .A3(sr_out[0]), .A4(n131), .Y(
        \_0_net_[0] ) );
  OR3X1_HVT U130 ( .A1(round_num[2]), .A2(round_num[0]), .A3(n3), .Y(n2) );
  NAND2X0_HVT U131 ( .A1(round_num[3]), .A2(round_num[1]), .Y(n3) );
  keygen_0 x ( .round_num(round_num), .keyin(keyin), .keyout({keyout[127:76], 
        n132, keyout[74:73], n133, keyout[71:70], n134, keyout[68:3], n135, 
        keyout[1:0]}) );
  subbytes sb ( .in({in[127:3], n106, in[1:0]}), .out(sb_out) );
  shift_rows sr ( .in(sb_out), .out(sr_out) );
  Mix_Column mc ( .in({sr_out[127:68], n8, sr_out[66:37], n20, sr_out[35:0]}), 
        .out(mc_out) );
  add_round_keys_1 adk ( .state({\_0_net_[127] , \_0_net_[126] , 
        \_0_net_[125] , \_0_net_[124] , \_0_net_[123] , \_0_net_[122] , 
        \_0_net_[121] , \_0_net_[120] , \_0_net_[119] , \_0_net_[118] , 
        \_0_net_[117] , \_0_net_[116] , \_0_net_[115] , \_0_net_[114] , 
        \_0_net_[113] , \_0_net_[112] , \_0_net_[111] , \_0_net_[110] , 
        \_0_net_[109] , \_0_net_[108] , \_0_net_[107] , \_0_net_[106] , 
        \_0_net_[105] , \_0_net_[104] , \_0_net_[103] , \_0_net_[102] , 
        \_0_net_[101] , \_0_net_[100] , \_0_net_[99] , \_0_net_[98] , 
        \_0_net_[97] , \_0_net_[96] , \_0_net_[95] , \_0_net_[94] , 
        \_0_net_[93] , \_0_net_[92] , \_0_net_[91] , \_0_net_[90] , 
        \_0_net_[89] , \_0_net_[88] , \_0_net_[87] , \_0_net_[86] , 
        \_0_net_[85] , \_0_net_[84] , \_0_net_[83] , \_0_net_[82] , 
        \_0_net_[81] , \_0_net_[80] , \_0_net_[79] , \_0_net_[78] , 
        \_0_net_[77] , \_0_net_[76] , \_0_net_[75] , \_0_net_[74] , 
        \_0_net_[73] , \_0_net_[72] , \_0_net_[71] , \_0_net_[70] , 
        \_0_net_[69] , \_0_net_[68] , \_0_net_[67] , \_0_net_[66] , 
        \_0_net_[65] , \_0_net_[64] , \_0_net_[63] , \_0_net_[62] , 
        \_0_net_[61] , \_0_net_[60] , \_0_net_[59] , \_0_net_[58] , 
        \_0_net_[57] , \_0_net_[56] , \_0_net_[55] , \_0_net_[54] , 
        \_0_net_[53] , \_0_net_[52] , \_0_net_[51] , \_0_net_[50] , 
        \_0_net_[49] , \_0_net_[48] , \_0_net_[47] , \_0_net_[46] , 
        \_0_net_[45] , \_0_net_[44] , \_0_net_[43] , \_0_net_[42] , 
        \_0_net_[41] , \_0_net_[40] , \_0_net_[39] , \_0_net_[38] , 
        \_0_net_[37] , \_0_net_[36] , \_0_net_[35] , \_0_net_[34] , 
        \_0_net_[33] , \_0_net_[32] , \_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_0_net_[0] }), 
        .subkey({keyout[127:76], n132, keyout[74:73], n133, keyout[71:70], 
        n134, keyout[68:3], n135, keyout[1:0]}), .out(out) );
  DELLN2X2_HVT U1 ( .A(sr_out[10]), .Y(n1) );
  DELLN2X2_HVT U3 ( .A(sr_out[9]), .Y(n4) );
  DELLN1X2_HVT U5 ( .A(sr_out[42]), .Y(n10) );
  NAND2X0_HVT U11 ( .A1(mc_out[76]), .A2(n116), .Y(n5) );
  NAND2X1_HVT U18 ( .A1(n14), .A2(n123), .Y(n6) );
  NAND2X0_HVT U19 ( .A1(n5), .A2(n6), .Y(\_0_net_[76] ) );
  INVX2_HVT U20 ( .A(n119), .Y(n116) );
  DELLN1X2_HVT U28 ( .A(sr_out[76]), .Y(n14) );
  INVX1_HVT U29 ( .A(sr_out[67]), .Y(n7) );
  INVX2_HVT U31 ( .A(n7), .Y(n8) );
  DELLN2X2_HVT U37 ( .A(sr_out[17]), .Y(n9) );
  DELLN2X2_HVT U39 ( .A(sr_out[11]), .Y(n11) );
  DELLN2X2_HVT U44 ( .A(sr_out[79]), .Y(n27) );
  DELLN2X2_HVT U45 ( .A(sr_out[7]), .Y(n12) );
  DELLN2X2_HVT U49 ( .A(sr_out[67]), .Y(n13) );
  DELLN2X2_HVT U54 ( .A(sr_out[12]), .Y(n15) );
  DELLN1X2_HVT U55 ( .A(sr_out[21]), .Y(n16) );
  NAND2X0_HVT U58 ( .A1(mc_out[25]), .A2(n112), .Y(n17) );
  NAND2X1_HVT U61 ( .A1(sr_out[25]), .A2(n127), .Y(n18) );
  NAND2X0_HVT U63 ( .A1(n17), .A2(n18), .Y(\_0_net_[25] ) );
  INVX1_HVT U64 ( .A(n135), .Y(n22) );
  NBUFFX2_HVT U71 ( .A(sr_out[87]), .Y(n19) );
  NAND2X0_HVT U72 ( .A1(sr_out[44]), .A2(n126), .Y(n88) );
  NBUFFX2_HVT U73 ( .A(sr_out[36]), .Y(n20) );
  DELLN2X2_HVT U75 ( .A(sr_out[8]), .Y(n21) );
  DELLN2X2_HVT U81 ( .A(sr_out[114]), .Y(n80) );
  INVX1_HVT U84 ( .A(n120), .Y(n112) );
  NAND2X0_HVT U86 ( .A1(sr_out[124]), .A2(n129), .Y(n47) );
  NAND2X0_HVT U89 ( .A1(sr_out[115]), .A2(n130), .Y(n29) );
  NAND2X0_HVT U90 ( .A1(sr_out[83]), .A2(n122), .Y(n63) );
  NAND2X0_HVT U102 ( .A1(sr_out[60]), .A2(n124), .Y(n71) );
  NAND2X0_HVT U105 ( .A1(sr_out[33]), .A2(n127), .Y(n33) );
  NAND2X0_HVT U107 ( .A1(sr_out[23]), .A2(n128), .Y(n37) );
  NAND2X0_HVT U112 ( .A1(n128), .A2(sr_out[1]), .Y(n55) );
  INVX0_HVT U121 ( .A(n22), .Y(keyout[2]) );
  NAND2X0_HVT U132 ( .A1(mc_out[85]), .A2(n117), .Y(n24) );
  NAND2X0_HVT U133 ( .A1(sr_out[85]), .A2(n122), .Y(n25) );
  NAND2X0_HVT U134 ( .A1(n24), .A2(n25), .Y(\_0_net_[85] ) );
  INVX1_HVT U135 ( .A(n119), .Y(n117) );
  DELLN2X2_HVT U136 ( .A(sr_out[18]), .Y(n26) );
  NAND2X0_HVT U137 ( .A1(mc_out[115]), .A2(n110), .Y(n28) );
  NAND2X0_HVT U138 ( .A1(n28), .A2(n29), .Y(\_0_net_[115] ) );
  NAND2X0_HVT U139 ( .A1(mc_out[99]), .A2(n118), .Y(n30) );
  NAND2X0_HVT U140 ( .A1(n121), .A2(sr_out[99]), .Y(n31) );
  NAND2X0_HVT U141 ( .A1(n30), .A2(n31), .Y(\_0_net_[99] ) );
  NAND2X0_HVT U142 ( .A1(mc_out[33]), .A2(n113), .Y(n32) );
  NAND2X0_HVT U143 ( .A1(n32), .A2(n33), .Y(\_0_net_[33] ) );
  INVX1_HVT U144 ( .A(n108), .Y(n127) );
  IBUFFX2_HVT U145 ( .A(sr_out[96]), .Y(n34) );
  INVX1_HVT U146 ( .A(n34), .Y(n35) );
  NAND2X0_HVT U147 ( .A1(sr_out[61]), .A2(n124), .Y(n67) );
  NAND2X0_HVT U148 ( .A1(mc_out[23]), .A2(n112), .Y(n36) );
  NAND2X0_HVT U149 ( .A1(n36), .A2(n37), .Y(\_0_net_[23] ) );
  NAND2X0_HVT U150 ( .A1(mc_out[121]), .A2(n111), .Y(n38) );
  NAND2X0_HVT U151 ( .A1(sr_out[121]), .A2(n129), .Y(n39) );
  NAND2X0_HVT U152 ( .A1(n38), .A2(n39), .Y(\_0_net_[121] ) );
  INVX1_HVT U153 ( .A(n120), .Y(n111) );
  NAND2X0_HVT U154 ( .A1(mc_out[107]), .A2(n110), .Y(n40) );
  NAND2X0_HVT U155 ( .A1(sr_out[107]), .A2(n130), .Y(n41) );
  NAND2X0_HVT U156 ( .A1(n40), .A2(n41), .Y(\_0_net_[107] ) );
  NAND2X0_HVT U157 ( .A1(mc_out[97]), .A2(n118), .Y(n42) );
  NAND2X0_HVT U158 ( .A1(sr_out[97]), .A2(n121), .Y(n43) );
  NAND2X0_HVT U159 ( .A1(n42), .A2(n43), .Y(\_0_net_[97] ) );
  NAND2X0_HVT U160 ( .A1(mc_out[28]), .A2(n112), .Y(n44) );
  NAND2X0_HVT U161 ( .A1(sr_out[28]), .A2(n127), .Y(n45) );
  NAND2X0_HVT U162 ( .A1(n44), .A2(n45), .Y(\_0_net_[28] ) );
  NAND2X0_HVT U163 ( .A1(mc_out[124]), .A2(n111), .Y(n46) );
  NAND2X0_HVT U164 ( .A1(n46), .A2(n47), .Y(\_0_net_[124] ) );
  NAND2X0_HVT U165 ( .A1(mc_out[49]), .A2(n114), .Y(n48) );
  NAND2X0_HVT U166 ( .A1(sr_out[49]), .A2(n125), .Y(n49) );
  NAND2X0_HVT U167 ( .A1(n48), .A2(n49), .Y(\_0_net_[49] ) );
  NAND2X0_HVT U168 ( .A1(mc_out[20]), .A2(n112), .Y(n50) );
  NAND2X0_HVT U169 ( .A1(n128), .A2(sr_out[20]), .Y(n51) );
  NAND2X0_HVT U170 ( .A1(n50), .A2(n51), .Y(\_0_net_[20] ) );
  IBUFFX2_HVT U171 ( .A(n133), .Y(n52) );
  INVX0_HVT U172 ( .A(n52), .Y(keyout[72]) );
  NAND2X0_HVT U173 ( .A1(mc_out[1]), .A2(n112), .Y(n54) );
  NAND2X0_HVT U174 ( .A1(n54), .A2(n55), .Y(\_0_net_[1] ) );
  NAND2X0_HVT U175 ( .A1(mc_out[37]), .A2(n113), .Y(n56) );
  NAND2X0_HVT U176 ( .A1(sr_out[37]), .A2(n126), .Y(n57) );
  NAND2X0_HVT U177 ( .A1(n56), .A2(n57), .Y(\_0_net_[37] ) );
  INVX1_HVT U178 ( .A(n119), .Y(n113) );
  NAND2X0_HVT U179 ( .A1(mc_out[46]), .A2(n114), .Y(n58) );
  NAND2X0_HVT U180 ( .A1(sr_out[46]), .A2(n125), .Y(n59) );
  NAND2X0_HVT U181 ( .A1(n58), .A2(n59), .Y(\_0_net_[46] ) );
  INVX1_HVT U182 ( .A(n109), .Y(n125) );
  NAND2X0_HVT U183 ( .A1(mc_out[73]), .A2(n116), .Y(n60) );
  NAND2X0_HVT U184 ( .A1(n123), .A2(sr_out[73]), .Y(n61) );
  NAND2X0_HVT U185 ( .A1(n60), .A2(n61), .Y(\_0_net_[73] ) );
  NAND2X0_HVT U186 ( .A1(mc_out[83]), .A2(n117), .Y(n62) );
  NAND2X0_HVT U187 ( .A1(n62), .A2(n63), .Y(\_0_net_[83] ) );
  NAND2X0_HVT U188 ( .A1(mc_out[75]), .A2(n116), .Y(n64) );
  NAND2X0_HVT U189 ( .A1(n123), .A2(sr_out[75]), .Y(n65) );
  NAND2X0_HVT U190 ( .A1(n64), .A2(n65), .Y(\_0_net_[75] ) );
  INVX1_HVT U191 ( .A(n109), .Y(n123) );
  NAND2X0_HVT U192 ( .A1(mc_out[61]), .A2(n115), .Y(n66) );
  NAND2X0_HVT U193 ( .A1(n66), .A2(n67), .Y(\_0_net_[61] ) );
  INVX0_HVT U194 ( .A(n109), .Y(n124) );
  NAND2X0_HVT U195 ( .A1(mc_out[84]), .A2(n117), .Y(n68) );
  NAND2X0_HVT U196 ( .A1(sr_out[84]), .A2(n122), .Y(n69) );
  NAND2X0_HVT U197 ( .A1(n68), .A2(n69), .Y(\_0_net_[84] ) );
  NAND2X0_HVT U198 ( .A1(mc_out[60]), .A2(n115), .Y(n70) );
  NAND2X0_HVT U199 ( .A1(n70), .A2(n71), .Y(\_0_net_[60] ) );
  NAND2X0_HVT U200 ( .A1(mc_out[66]), .A2(n115), .Y(n72) );
  NAND2X0_HVT U201 ( .A1(sr_out[66]), .A2(n124), .Y(n73) );
  NAND2X0_HVT U202 ( .A1(n72), .A2(n73), .Y(\_0_net_[66] ) );
  NAND2X0_HVT U203 ( .A1(mc_out[91]), .A2(n117), .Y(n74) );
  NAND2X0_HVT U204 ( .A1(sr_out[91]), .A2(n121), .Y(n75) );
  NAND2X0_HVT U205 ( .A1(n74), .A2(n75), .Y(\_0_net_[91] ) );
  NAND2X0_HVT U206 ( .A1(mc_out[57]), .A2(n115), .Y(n76) );
  NAND2X0_HVT U207 ( .A1(sr_out[57]), .A2(n124), .Y(n77) );
  NAND2X0_HVT U208 ( .A1(n76), .A2(n77), .Y(\_0_net_[57] ) );
  NAND2X0_HVT U209 ( .A1(n125), .A2(sr_out[52]), .Y(n82) );
  IBUFFX2_HVT U210 ( .A(n132), .Y(n78) );
  INVX0_HVT U211 ( .A(n78), .Y(keyout[75]) );
  NAND2X0_HVT U212 ( .A1(mc_out[52]), .A2(n114), .Y(n81) );
  NAND2X0_HVT U213 ( .A1(n81), .A2(n82), .Y(\_0_net_[52] ) );
  INVX1_HVT U214 ( .A(n119), .Y(n114) );
  NAND2X0_HVT U215 ( .A1(mc_out[43]), .A2(n114), .Y(n83) );
  NAND2X0_HVT U216 ( .A1(n126), .A2(sr_out[43]), .Y(n84) );
  NAND2X0_HVT U217 ( .A1(n83), .A2(n84), .Y(\_0_net_[43] ) );
  NAND2X0_HVT U218 ( .A1(mc_out[35]), .A2(n113), .Y(n85) );
  NAND2X0_HVT U219 ( .A1(sr_out[35]), .A2(n126), .Y(n86) );
  NAND2X0_HVT U220 ( .A1(n85), .A2(n86), .Y(\_0_net_[35] ) );
  NAND2X0_HVT U221 ( .A1(mc_out[44]), .A2(n114), .Y(n87) );
  NAND2X0_HVT U222 ( .A1(n87), .A2(n88), .Y(\_0_net_[44] ) );
  NAND2X0_HVT U223 ( .A1(mc_out[36]), .A2(n113), .Y(n89) );
  NAND2X0_HVT U224 ( .A1(sr_out[36]), .A2(n126), .Y(n90) );
  NAND2X0_HVT U225 ( .A1(n89), .A2(n90), .Y(\_0_net_[36] ) );
  INVX1_HVT U226 ( .A(n108), .Y(n126) );
  NAND2X0_HVT U227 ( .A1(n11), .A2(n129), .Y(n93) );
  NAND2X0_HVT U228 ( .A1(sr_out[51]), .A2(n125), .Y(n102) );
  NAND2X0_HVT U229 ( .A1(sr_out[68]), .A2(n123), .Y(n98) );
  DELLN2X2_HVT U230 ( .A(sr_out[103]), .Y(n107) );
  DELLN2X2_HVT U231 ( .A(sr_out[111]), .Y(n91) );
  NAND2X0_HVT U232 ( .A1(mc_out[11]), .A2(n111), .Y(n92) );
  NAND2X0_HVT U233 ( .A1(n92), .A2(n93), .Y(\_0_net_[11] ) );
  DELLN2X2_HVT U234 ( .A(sr_out[15]), .Y(n94) );
  DELLN2X2_HVT U235 ( .A(sr_out[55]), .Y(n95) );
  DELLN2X2_HVT U236 ( .A(sr_out[14]), .Y(n96) );
  NAND2X0_HVT U237 ( .A1(mc_out[68]), .A2(n115), .Y(n97) );
  NAND2X0_HVT U238 ( .A1(n97), .A2(n98), .Y(\_0_net_[68] ) );
  IBUFFX2_HVT U239 ( .A(n134), .Y(n99) );
  INVX0_HVT U240 ( .A(n99), .Y(keyout[69]) );
  DELLN2X2_HVT U241 ( .A(sr_out[39]), .Y(n105) );
  NAND2X0_HVT U242 ( .A1(mc_out[51]), .A2(n114), .Y(n101) );
  NAND2X0_HVT U243 ( .A1(n101), .A2(n102), .Y(\_0_net_[51] ) );
  DELLN2X2_HVT U244 ( .A(sr_out[47]), .Y(n103) );
  DELLN2X2_HVT U245 ( .A(sr_out[31]), .Y(n104) );
  NBUFFX16_HVT U246 ( .A(in[2]), .Y(n106) );
  INVX0_HVT U247 ( .A(n119), .Y(n118) );
  INVX1_HVT U248 ( .A(n2), .Y(n119) );
  INVX1_HVT U249 ( .A(n109), .Y(n122) );
  INVX1_HVT U250 ( .A(n109), .Y(n121) );
  INVX1_HVT U251 ( .A(n108), .Y(n128) );
  INVX1_HVT U252 ( .A(n108), .Y(n129) );
  INVX1_HVT U253 ( .A(n108), .Y(n130) );
  INVX1_HVT U254 ( .A(n108), .Y(n131) );
  INVX1_HVT U255 ( .A(n119), .Y(n115) );
  INVX1_HVT U256 ( .A(n120), .Y(n109) );
  INVX1_HVT U257 ( .A(n120), .Y(n110) );
  INVX1_HVT U258 ( .A(n120), .Y(n108) );
  INVX0_HVT U259 ( .A(n2), .Y(n120) );
endmodule

