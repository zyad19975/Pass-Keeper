
module aes ( plaintext, key, clk, reset, cipher_text, ready );
  input [127:0] plaintext;
  input [127:0] key;
  output [127:0] cipher_text;
  input clk, reset;
  output ready;
  wire   n4, n5, n8, n12, n13, n14, n15, n16, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n42, n43, n44, n45, n46, n47, n48, n49, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n130, n132, n133, n134, n135,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n168, n169, n170,
         n171, n172, n173, n174, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n255, n256, n257, n258, n259, n260, n261, n262,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827;
  wire   [127:0] adk_out0;
  wire   [127:0] adk_in;
  wire   [3:0] round_number;
  wire   [127:0] key_round;
  wire   [127:0] keyout;

  add_round_keys_0 adk_0 ( .state(plaintext), .subkey(key), .out(adk_out0) );
  round r1 ( .in({n629, adk_in[126:125], n640, adk_in[123:122], n700, 
        adk_in[120], n600, adk_in[118:104], n636, adk_in[102:99], n801, 
        adk_in[97:96], n608, adk_in[94:83], n641, adk_in[81:80], n632, 
        adk_in[78:77], n736, adk_in[75], n620, adk_in[73:72], n757, 
        adk_in[70:68], n670, n642, n638, adk_in[64:60], n683, adk_in[58:56], 
        n615, adk_in[54], n604, adk_in[52:51], n708, adk_in[49:48], n619, 
        adk_in[46], n611, adk_in[44:30], n623, adk_in[28:27], n694, 
        adk_in[25:8], n691, adk_in[6:3], n647, adk_in[1:0]}), .round_num({n358, 
        n408, n361, n575}), .keyin({key_round[127:32], n824, key_round[30:28], 
        n654, key_round[26:21], n628, key_round[19:16], n726, key_round[14:10], 
        n693, key_round[8:2], n716, key_round[0]}), .keyout(keyout), .out(
        cipher_text) );
  DFFX1_HVT \round_number_reg[0]  ( .D(n279), .CLK(clk), .Q(n826), .QN(n574)
         );
  DFFX1_HVT \round_number_reg[3]  ( .D(n278), .CLK(clk), .Q(round_number[3]), 
        .QN(n763) );
  DFFX1_HVT \round_number_reg[1]  ( .D(n277), .CLK(clk), .Q(round_number[1]), 
        .QN(n5) );
  DFFX1_HVT \adk_in_reg[0]  ( .D(n275), .CLK(clk), .Q(adk_in[0]) );
  DFFX1_HVT \adk_in_reg[1]  ( .D(n274), .CLK(clk), .Q(adk_in[1]), .QN(n705) );
  DFFX1_HVT \adk_in_reg[2]  ( .D(n273), .CLK(clk), .Q(n647), .QN(n324) );
  DFFX1_HVT \adk_in_reg[3]  ( .D(n272), .CLK(clk), .Q(adk_in[3]), .QN(n665) );
  DFFX1_HVT \adk_in_reg[4]  ( .D(n271), .CLK(clk), .Q(adk_in[4]), .QN(n661) );
  DFFX1_HVT \adk_in_reg[5]  ( .D(n270), .CLK(clk), .Q(adk_in[5]), .QN(n504) );
  DFFX1_HVT \adk_in_reg[6]  ( .D(n269), .CLK(clk), .Q(adk_in[6]) );
  DFFX1_HVT \adk_in_reg[7]  ( .D(n268), .CLK(clk), .Q(adk_in[7]), .QN(n690) );
  DFFX1_HVT \adk_in_reg[8]  ( .D(n267), .CLK(clk), .Q(adk_in[8]) );
  DFFX1_HVT \adk_in_reg[9]  ( .D(n266), .CLK(clk), .Q(adk_in[9]), .QN(n747) );
  DFFX1_HVT \adk_in_reg[10]  ( .D(n265), .CLK(clk), .Q(adk_in[10]), .QN(n625)
         );
  DFFX1_HVT \adk_in_reg[11]  ( .D(n264), .CLK(clk), .Q(adk_in[11]), .QN(n703)
         );
  DFFX1_HVT \adk_in_reg[12]  ( .D(n380), .CLK(clk), .Q(adk_in[12]), .QN(n711)
         );
  DFFX1_HVT \adk_in_reg[13]  ( .D(n262), .CLK(clk), .Q(adk_in[13]) );
  DFFX1_HVT \adk_in_reg[14]  ( .D(n261), .CLK(clk), .Q(adk_in[14]) );
  DFFX1_HVT \adk_in_reg[15]  ( .D(n260), .CLK(clk), .Q(adk_in[15]), .QN(n356)
         );
  DFFX1_HVT \adk_in_reg[16]  ( .D(n259), .CLK(clk), .Q(adk_in[16]), .QN(n468)
         );
  DFFX1_HVT \adk_in_reg[17]  ( .D(n258), .CLK(clk), .Q(adk_in[17]), .QN(n729)
         );
  DFFX1_HVT \adk_in_reg[18]  ( .D(n257), .CLK(clk), .Q(adk_in[18]) );
  DFFX1_HVT \adk_in_reg[19]  ( .D(n256), .CLK(clk), .Q(adk_in[19]), .QN(n671)
         );
  DFFX1_HVT \adk_in_reg[20]  ( .D(n255), .CLK(clk), .Q(adk_in[20]), .QN(n633)
         );
  DFFX1_HVT \adk_in_reg[21]  ( .D(n492), .CLK(clk), .Q(adk_in[21]), .QN(n515)
         );
  DFFX1_HVT \adk_in_reg[23]  ( .D(n252), .CLK(clk), .Q(adk_in[23]), .QN(n749)
         );
  DFFX1_HVT \adk_in_reg[24]  ( .D(n251), .CLK(clk), .Q(adk_in[24]) );
  DFFX1_HVT \adk_in_reg[25]  ( .D(n250), .CLK(clk), .Q(adk_in[25]), .QN(n659)
         );
  DFFX1_HVT \adk_in_reg[26]  ( .D(n249), .CLK(clk), .Q(n694), .QN(n352) );
  DFFX1_HVT \adk_in_reg[27]  ( .D(n248), .CLK(clk), .Q(adk_in[27]), .QN(n684)
         );
  DFFX1_HVT \adk_in_reg[28]  ( .D(n247), .CLK(clk), .Q(adk_in[28]), .QN(n686)
         );
  DFFX1_HVT \adk_in_reg[29]  ( .D(n246), .CLK(clk), .Q(n623) );
  DFFX1_HVT \adk_in_reg[31]  ( .D(n244), .CLK(clk), .Q(adk_in[31]) );
  DFFX1_HVT \adk_in_reg[32]  ( .D(n243), .CLK(clk), .Q(adk_in[32]) );
  DFFX1_HVT \adk_in_reg[33]  ( .D(n242), .CLK(clk), .Q(adk_in[33]), .QN(n731)
         );
  DFFX1_HVT \adk_in_reg[34]  ( .D(n241), .CLK(clk), .Q(adk_in[34]) );
  DFFX1_HVT \adk_in_reg[35]  ( .D(n240), .CLK(clk), .Q(adk_in[35]), .QN(n673)
         );
  DFFX1_HVT \adk_in_reg[36]  ( .D(n239), .CLK(clk), .Q(adk_in[36]), .QN(n759)
         );
  DFFX1_HVT \adk_in_reg[37]  ( .D(n238), .CLK(clk), .Q(adk_in[37]) );
  DFFX1_HVT \adk_in_reg[39]  ( .D(n236), .CLK(clk), .Q(adk_in[39]), .QN(n743)
         );
  DFFX1_HVT \adk_in_reg[40]  ( .D(n235), .CLK(clk), .Q(adk_in[40]) );
  DFFX1_HVT \adk_in_reg[41]  ( .D(n234), .CLK(clk), .Q(adk_in[41]), .QN(n605)
         );
  DFFX1_HVT \adk_in_reg[42]  ( .D(n233), .CLK(clk), .Q(adk_in[42]), .QN(n609)
         );
  DFFX1_HVT \adk_in_reg[43]  ( .D(n232), .CLK(clk), .Q(adk_in[43]), .QN(n651)
         );
  DFFX1_HVT \adk_in_reg[44]  ( .D(n418), .CLK(clk), .Q(adk_in[44]), .QN(n737)
         );
  DFFX1_HVT \adk_in_reg[45]  ( .D(n230), .CLK(clk), .Q(n611) );
  DFFX1_HVT \adk_in_reg[47]  ( .D(n228), .CLK(clk), .Q(adk_in[47]), .QN(n618)
         );
  DFFX1_HVT \adk_in_reg[48]  ( .D(n227), .CLK(clk), .Q(adk_in[48]) );
  DFFX1_HVT \adk_in_reg[49]  ( .D(n226), .CLK(clk), .Q(adk_in[49]), .QN(n745)
         );
  DFFX1_HVT \adk_in_reg[50]  ( .D(n225), .CLK(clk), .Q(adk_in[50]), .QN(n707)
         );
  DFFX1_HVT \adk_in_reg[51]  ( .D(n224), .CLK(clk), .Q(adk_in[51]), .QN(n657)
         );
  DFFX1_HVT \adk_in_reg[52]  ( .D(n223), .CLK(clk), .Q(adk_in[52]), .QN(n733)
         );
  DFFX1_HVT \adk_in_reg[53]  ( .D(n222), .CLK(clk), .Q(adk_in[53]), .QN(n603)
         );
  DFFX1_HVT \adk_in_reg[55]  ( .D(n220), .CLK(clk), .Q(adk_in[55]), .QN(n614)
         );
  DFFX1_HVT \adk_in_reg[56]  ( .D(n219), .CLK(clk), .Q(adk_in[56]) );
  DFFX1_HVT \adk_in_reg[57]  ( .D(n218), .CLK(clk), .Q(adk_in[57]), .QN(n695)
         );
  DFFX1_HVT \adk_in_reg[58]  ( .D(n217), .CLK(clk), .Q(adk_in[58]) );
  DFFX1_HVT \adk_in_reg[59]  ( .D(n216), .CLK(clk), .Q(adk_in[59]), .QN(n682)
         );
  DFFX1_HVT \adk_in_reg[60]  ( .D(n215), .CLK(clk), .Q(adk_in[60]), .QN(n751)
         );
  DFFX1_HVT \adk_in_reg[61]  ( .D(n214), .CLK(clk), .Q(adk_in[61]), .QN(n316)
         );
  DFFX1_HVT \adk_in_reg[63]  ( .D(n212), .CLK(clk), .Q(adk_in[63]), .QN(n755)
         );
  DFFX1_HVT \adk_in_reg[64]  ( .D(n211), .CLK(clk), .Q(adk_in[64]) );
  DFFX1_HVT \adk_in_reg[65]  ( .D(n210), .CLK(clk), .Q(adk_in[65]), .QN(n637)
         );
  DFFX1_HVT \adk_in_reg[67]  ( .D(n208), .CLK(clk), .Q(adk_in[67]), .QN(n669)
         );
  DFFX1_HVT \adk_in_reg[68]  ( .D(n207), .CLK(clk), .Q(adk_in[68]), .QN(n741)
         );
  DFFX1_HVT \adk_in_reg[69]  ( .D(n206), .CLK(clk), .Q(adk_in[69]) );
  DFFX1_HVT \adk_in_reg[70]  ( .D(n524), .CLK(clk), .Q(adk_in[70]), .QN(n540)
         );
  DFFX1_HVT \adk_in_reg[71]  ( .D(n204), .CLK(clk), .Q(n757), .QN(n322) );
  DFFX1_HVT \adk_in_reg[72]  ( .D(n203), .CLK(clk), .Q(adk_in[72]) );
  DFFX1_HVT \adk_in_reg[73]  ( .D(n202), .CLK(clk), .Q(adk_in[73]), .QN(n675)
         );
  DFFX1_HVT \adk_in_reg[74]  ( .D(n201), .CLK(clk), .Q(n620) );
  DFFX1_HVT \adk_in_reg[75]  ( .D(n200), .CLK(clk), .Q(adk_in[75]), .QN(n663)
         );
  DFFX1_HVT \adk_in_reg[76]  ( .D(n199), .CLK(clk), .Q(adk_in[76]), .QN(n735)
         );
  DFFX1_HVT \adk_in_reg[77]  ( .D(n198), .CLK(clk), .Q(adk_in[77]) );
  DFFX1_HVT \adk_in_reg[78]  ( .D(n197), .CLK(clk), .Q(adk_in[78]) );
  DFFX1_HVT \adk_in_reg[79]  ( .D(n196), .CLK(clk), .Q(n632) );
  DFFX1_HVT \adk_in_reg[80]  ( .D(n195), .CLK(clk), .Q(adk_in[80]) );
  DFFX1_HVT \adk_in_reg[81]  ( .D(n194), .CLK(clk), .Q(adk_in[81]), .QN(n648)
         );
  DFFX1_HVT \adk_in_reg[82]  ( .D(n193), .CLK(clk), .Q(n641) );
  DFFX1_HVT \adk_in_reg[83]  ( .D(n192), .CLK(clk), .Q(adk_in[83]), .QN(n680)
         );
  DFFX1_HVT \adk_in_reg[84]  ( .D(n191), .CLK(clk), .Q(adk_in[84]), .QN(n723)
         );
  DFFX1_HVT \adk_in_reg[85]  ( .D(n190), .CLK(clk), .Q(adk_in[85]), .QN(n532)
         );
  DFFX1_HVT \adk_in_reg[87]  ( .D(n188), .CLK(clk), .Q(adk_in[87]), .QN(n563)
         );
  DFFX1_HVT \adk_in_reg[88]  ( .D(n187), .CLK(clk), .Q(adk_in[88]) );
  DFFX1_HVT \adk_in_reg[89]  ( .D(n186), .CLK(clk), .Q(adk_in[89]), .QN(n719)
         );
  DFFX1_HVT \adk_in_reg[90]  ( .D(n185), .CLK(clk), .Q(adk_in[90]), .QN(n552)
         );
  DFFX1_HVT \adk_in_reg[91]  ( .D(n184), .CLK(clk), .Q(adk_in[91]), .QN(n616)
         );
  DFFX1_HVT \adk_in_reg[92]  ( .D(n183), .CLK(clk), .Q(adk_in[92]), .QN(n645)
         );
  DFFX1_HVT \adk_in_reg[93]  ( .D(n182), .CLK(clk), .Q(adk_in[93]) );
  DFFX1_HVT \adk_in_reg[94]  ( .D(n181), .CLK(clk), .Q(adk_in[94]) );
  DFFX1_HVT \adk_in_reg[95]  ( .D(n180), .CLK(clk), .Q(adk_in[95]), .QN(n607)
         );
  DFFX1_HVT \adk_in_reg[96]  ( .D(n179), .CLK(clk), .Q(adk_in[96]) );
  DFFX1_HVT \adk_in_reg[97]  ( .D(n178), .CLK(clk), .Q(adk_in[97]), .QN(n643)
         );
  DFFX1_HVT \adk_in_reg[99]  ( .D(n176), .CLK(clk), .Q(adk_in[99]), .QN(n655)
         );
  DFFX1_HVT \adk_in_reg[100]  ( .D(n366), .CLK(clk), .Q(adk_in[100]), .QN(n721) );
  DFFX1_HVT \adk_in_reg[101]  ( .D(n174), .CLK(clk), .Q(adk_in[101]) );
  DFFX1_HVT \adk_in_reg[102]  ( .D(n173), .CLK(clk), .Q(adk_in[102]), .QN(n472) );
  DFFX1_HVT \adk_in_reg[103]  ( .D(n172), .CLK(clk), .Q(adk_in[103]), .QN(n635) );
  DFFX1_HVT \adk_in_reg[104]  ( .D(n171), .CLK(clk), .Q(adk_in[104]) );
  DFFX1_HVT \adk_in_reg[105]  ( .D(n170), .CLK(clk), .Q(adk_in[105]), .QN(n697) );
  DFFX1_HVT \adk_in_reg[106]  ( .D(n169), .CLK(clk), .Q(adk_in[106]), .QN(n709) );
  DFFX1_HVT \adk_in_reg[107]  ( .D(n168), .CLK(clk), .Q(adk_in[107]), .QN(n713) );
  DFFX1_HVT \adk_in_reg[108]  ( .D(n288), .CLK(clk), .Q(adk_in[108]), .QN(n717) );
  DFFX1_HVT \adk_in_reg[109]  ( .D(n166), .CLK(clk), .Q(adk_in[109]), .QN(n327) );
  DFFX1_HVT \adk_in_reg[111]  ( .D(n164), .CLK(clk), .Q(adk_in[111]), .QN(n758) );
  DFFX1_HVT \adk_in_reg[112]  ( .D(n163), .CLK(clk), .Q(adk_in[112]), .QN(n557) );
  DFFX1_HVT \adk_in_reg[113]  ( .D(n162), .CLK(clk), .Q(adk_in[113]), .QN(n727) );
  DFFX1_HVT \adk_in_reg[114]  ( .D(n161), .CLK(clk), .Q(adk_in[114]) );
  DFFX1_HVT \adk_in_reg[115]  ( .D(n160), .CLK(clk), .Q(adk_in[115]), .QN(n650) );
  DFFX1_HVT \adk_in_reg[116]  ( .D(n159), .CLK(clk), .Q(adk_in[116]), .QN(n739) );
  DFFX1_HVT \adk_in_reg[117]  ( .D(n158), .CLK(clk), .Q(adk_in[117]), .QN(n446) );
  DFFX1_HVT \adk_in_reg[118]  ( .D(n157), .CLK(clk), .Q(adk_in[118]) );
  DFFX1_HVT \adk_in_reg[119]  ( .D(n156), .CLK(clk), .Q(adk_in[119]), .QN(n599) );
  DFFX1_HVT \adk_in_reg[120]  ( .D(n155), .CLK(clk), .Q(adk_in[120]) );
  DFFX1_HVT \adk_in_reg[121]  ( .D(n154), .CLK(clk), .Q(adk_in[121]), .QN(n699) );
  DFFX1_HVT \adk_in_reg[122]  ( .D(n153), .CLK(clk), .Q(adk_in[122]), .QN(n314) );
  DFFX1_HVT \adk_in_reg[123]  ( .D(n152), .CLK(clk), .Q(adk_in[123]), .QN(n667) );
  DFFX1_HVT \adk_in_reg[124]  ( .D(n151), .CLK(clk), .Q(adk_in[124]), .QN(n639) );
  DFFX1_HVT \adk_in_reg[125]  ( .D(n150), .CLK(clk), .Q(adk_in[125]) );
  DFFX1_HVT \adk_in_reg[127]  ( .D(n148), .CLK(clk), .Q(n629) );
  DFFX1_HVT \key_round_reg[1]  ( .D(n146), .CLK(clk), .Q(key_round[1]), .QN(
        n715) );
  DFFX1_HVT \key_round_reg[3]  ( .D(n144), .CLK(clk), .Q(key_round[3]), .QN(
        n630) );
  DFFX1_HVT \key_round_reg[4]  ( .D(n143), .CLK(clk), .Q(key_round[4]), .QN(
        n612) );
  DFFX1_HVT \key_round_reg[5]  ( .D(n142), .CLK(clk), .Q(key_round[5]), .QN(
        n294) );
  DFFX1_HVT \key_round_reg[6]  ( .D(n141), .CLK(clk), .Q(key_round[6]) );
  DFFX1_HVT \key_round_reg[7]  ( .D(n140), .CLK(clk), .Q(key_round[7]), .QN(
        n601) );
  DFFX1_HVT \key_round_reg[9]  ( .D(n138), .CLK(clk), .Q(key_round[9]), .QN(
        n692) );
  DFFX1_HVT \key_round_reg[10]  ( .D(n137), .CLK(clk), .Q(key_round[10]) );
  DFFX1_HVT \key_round_reg[11]  ( .D(n385), .CLK(clk), .Q(key_round[11]), .QN(
        n494) );
  DFFX1_HVT \key_round_reg[12]  ( .D(n135), .CLK(clk), .Q(key_round[12]), .QN(
        n688) );
  DFFX1_HVT \key_round_reg[13]  ( .D(n134), .CLK(clk), .Q(key_round[13]) );
  DFFX1_HVT \key_round_reg[14]  ( .D(n133), .CLK(clk), .Q(key_round[14]), .QN(
        n407) );
  DFFX1_HVT \key_round_reg[15]  ( .D(n132), .CLK(clk), .Q(key_round[15]), .QN(
        n725) );
  DFFX1_HVT \key_round_reg[16]  ( .D(n285), .CLK(clk), .Q(key_round[16]), .QN(
        n371) );
  DFFX1_HVT \key_round_reg[17]  ( .D(n130), .CLK(clk), .Q(key_round[17]), .QN(
        n677) );
  DFFX1_HVT \key_round_reg[18]  ( .D(n280), .CLK(clk), .Q(key_round[18]), .QN(
        n336) );
  DFFX1_HVT \key_round_reg[19]  ( .D(n128), .CLK(clk), .Q(key_round[19]), .QN(
        n621) );
  DFFX1_HVT \key_round_reg[20]  ( .D(n127), .CLK(clk), .Q(key_round[20]), .QN(
        n627) );
  DFFX1_HVT \key_round_reg[21]  ( .D(n126), .CLK(clk), .Q(key_round[21]), .QN(
        n293) );
  DFFX1_HVT \key_round_reg[23]  ( .D(n124), .CLK(clk), .Q(key_round[23]), .QN(
        n753) );
  DFFX1_HVT \key_round_reg[24]  ( .D(n123), .CLK(clk), .Q(key_round[24]) );
  DFFX1_HVT \key_round_reg[25]  ( .D(n122), .CLK(clk), .Q(key_round[25]), .QN(
        n624) );
  DFFX1_HVT \key_round_reg[26]  ( .D(n121), .CLK(clk), .Q(key_round[26]), .QN(
        n406) );
  DFFX1_HVT \key_round_reg[27]  ( .D(n120), .CLK(clk), .Q(key_round[27]), .QN(
        n653) );
  DFFX1_HVT \key_round_reg[28]  ( .D(n119), .CLK(clk), .Q(key_round[28]), .QN(
        n701) );
  DFFX1_HVT \key_round_reg[29]  ( .D(n118), .CLK(clk), .Q(key_round[29]) );
  DFFX1_HVT \key_round_reg[30]  ( .D(n117), .CLK(clk), .Q(key_round[30]), .QN(
        n295) );
  DFFX1_HVT \key_round_reg[31]  ( .D(n116), .CLK(clk), .Q(n679), .QN(n761) );
  DFFX1_HVT \key_round_reg[32]  ( .D(n115), .CLK(clk), .Q(key_round[32]) );
  DFFX1_HVT \key_round_reg[33]  ( .D(n114), .CLK(clk), .Q(key_round[33]) );
  DFFX1_HVT \key_round_reg[34]  ( .D(n113), .CLK(clk), .Q(key_round[34]), .QN(
        n422) );
  DFFX1_HVT \key_round_reg[35]  ( .D(n112), .CLK(clk), .Q(key_round[35]), .QN(
        n425) );
  DFFX1_HVT \key_round_reg[36]  ( .D(n111), .CLK(clk), .Q(key_round[36]) );
  DFFX1_HVT \key_round_reg[37]  ( .D(n110), .CLK(clk), .Q(key_round[37]) );
  DFFX1_HVT \key_round_reg[38]  ( .D(n109), .CLK(clk), .Q(key_round[38]) );
  DFFX1_HVT \key_round_reg[40]  ( .D(n440), .CLK(clk), .Q(key_round[40]), .QN(
        n443) );
  DFFX1_HVT \key_round_reg[41]  ( .D(n106), .CLK(clk), .Q(key_round[41]) );
  DFFX1_HVT \key_round_reg[42]  ( .D(n105), .CLK(clk), .Q(key_round[42]), .QN(
        n330) );
  DFFX1_HVT \key_round_reg[43]  ( .D(n104), .CLK(clk), .Q(key_round[43]) );
  DFFX1_HVT \key_round_reg[44]  ( .D(n103), .CLK(clk), .Q(key_round[44]), .QN(
        n411) );
  DFFX1_HVT \key_round_reg[46]  ( .D(n101), .CLK(clk), .Q(key_round[46]), .QN(
        n414) );
  DFFX1_HVT \key_round_reg[47]  ( .D(n100), .CLK(clk), .Q(key_round[47]), .QN(
        n393) );
  DFFX1_HVT \key_round_reg[50]  ( .D(n97), .CLK(clk), .Q(key_round[50]), .QN(
        n501) );
  DFFX1_HVT \key_round_reg[53]  ( .D(n94), .CLK(clk), .Q(key_round[53]) );
  DFFX1_HVT \key_round_reg[54]  ( .D(n93), .CLK(clk), .Q(key_round[54]) );
  DFFX1_HVT \key_round_reg[55]  ( .D(n92), .CLK(clk), .Q(key_round[55]) );
  DFFX1_HVT \key_round_reg[56]  ( .D(n91), .CLK(clk), .Q(key_round[56]), .QN(
        n461) );
  DFFX1_HVT \key_round_reg[64]  ( .D(n83), .CLK(clk), .Q(key_round[64]), .QN(
        n465) );
  DFFX1_HVT \key_round_reg[65]  ( .D(n82), .CLK(clk), .Q(key_round[65]) );
  DFFX1_HVT \key_round_reg[70]  ( .D(n77), .CLK(clk), .Q(key_round[70]) );
  DFFX1_HVT \key_round_reg[71]  ( .D(n76), .CLK(clk), .Q(key_round[71]) );
  DFFX1_HVT \key_round_reg[72]  ( .D(n75), .CLK(clk), .Q(key_round[72]) );
  DFFX1_HVT \key_round_reg[73]  ( .D(n74), .CLK(clk), .Q(key_round[73]) );
  DFFX1_HVT \key_round_reg[74]  ( .D(n73), .CLK(clk), .Q(key_round[74]) );
  DFFX1_HVT \key_round_reg[75]  ( .D(n72), .CLK(clk), .Q(key_round[75]) );
  DFFX1_HVT \key_round_reg[77]  ( .D(n70), .CLK(clk), .Q(key_round[77]) );
  DFFX1_HVT \key_round_reg[78]  ( .D(n69), .CLK(clk), .Q(key_round[78]), .QN(
        n329) );
  DFFX1_HVT \key_round_reg[79]  ( .D(n68), .CLK(clk), .Q(key_round[79]), .QN(
        n292) );
  DFFX1_HVT \key_round_reg[81]  ( .D(n66), .CLK(clk), .Q(key_round[81]) );
  DFFX1_HVT \key_round_reg[84]  ( .D(n63), .CLK(clk), .Q(key_round[84]), .QN(
        n537) );
  DFFX1_HVT \key_round_reg[86]  ( .D(n61), .CLK(clk), .Q(key_round[86]) );
  DFFX1_HVT \key_round_reg[87]  ( .D(n60), .CLK(clk), .Q(key_round[87]) );
  DFFX1_HVT \key_round_reg[94]  ( .D(n53), .CLK(clk), .Q(key_round[94]) );
  DFFX1_HVT \key_round_reg[95]  ( .D(n52), .CLK(clk), .Q(key_round[95]) );
  AO222X1_HVT U7 ( .A1(keyout[127]), .A2(n594), .A3(key[127]), .A4(n781), .A5(
        key_round[127]), .A6(n811), .Y(n20) );
  AO222X1_HVT U9 ( .A1(keyout[125]), .A2(n596), .A3(key[125]), .A4(n779), .A5(
        key_round[125]), .A6(n811), .Y(n22) );
  AO222X1_HVT U10 ( .A1(keyout[124]), .A2(n589), .A3(key[124]), .A4(n376), 
        .A5(key_round[124]), .A6(n313), .Y(n23) );
  AO222X1_HVT U13 ( .A1(keyout[121]), .A2(n598), .A3(key[121]), .A4(n795), 
        .A5(key_round[121]), .A6(n300), .Y(n26) );
  AO222X1_HVT U14 ( .A1(keyout[120]), .A2(n582), .A3(key[120]), .A4(n781), 
        .A5(key_round[120]), .A6(n284), .Y(n27) );
  AO222X1_HVT U17 ( .A1(keyout[117]), .A2(n589), .A3(key[117]), .A4(n785), 
        .A5(key_round[117]), .A6(n310), .Y(n30) );
  AO222X1_HVT U19 ( .A1(keyout[115]), .A2(n551), .A3(key[115]), .A4(n375), 
        .A5(key_round[115]), .A6(n340), .Y(n32) );
  AO222X1_HVT U21 ( .A1(keyout[113]), .A2(n298), .A3(key[113]), .A4(n791), 
        .A5(key_round[113]), .A6(n284), .Y(n34) );
  AO222X1_HVT U24 ( .A1(keyout[110]), .A2(n580), .A3(key[110]), .A4(n787), 
        .A5(key_round[110]), .A6(n811), .Y(n37) );
  AO222X1_HVT U26 ( .A1(keyout[108]), .A2(n304), .A3(key[108]), .A4(n789), 
        .A5(key_round[108]), .A6(n488), .Y(n39) );
  AO222X1_HVT U30 ( .A1(keyout[104]), .A2(n577), .A3(key[104]), .A4(n770), 
        .A5(key_round[104]), .A6(n355), .Y(n43) );
  AO222X1_HVT U32 ( .A1(keyout[102]), .A2(n298), .A3(key[102]), .A4(n800), 
        .A5(key_round[102]), .A6(n488), .Y(n45) );
  AO222X1_HVT U34 ( .A1(keyout[100]), .A2(n586), .A3(key[100]), .A4(n798), 
        .A5(key_round[100]), .A6(n313), .Y(n47) );
  AO222X1_HVT U35 ( .A1(keyout[99]), .A2(n596), .A3(key[99]), .A4(n797), .A5(
        key_round[99]), .A6(n807), .Y(n48) );
  AO222X1_HVT U39 ( .A1(keyout[95]), .A2(n587), .A3(key[95]), .A4(n791), .A5(
        key_round[95]), .A6(n312), .Y(n52) );
  AO222X1_HVT U40 ( .A1(keyout[94]), .A2(n578), .A3(key[94]), .A4(n790), .A5(
        key_round[94]), .A6(n808), .Y(n53) );
  AO222X1_HVT U41 ( .A1(keyout[93]), .A2(n593), .A3(key[93]), .A4(n782), .A5(
        key_round[93]), .A6(n807), .Y(n54) );
  AO222X1_HVT U42 ( .A1(keyout[92]), .A2(n390), .A3(key[92]), .A4(n795), .A5(
        key_round[92]), .A6(n808), .Y(n55) );
  AO222X1_HVT U43 ( .A1(keyout[91]), .A2(n589), .A3(key[91]), .A4(n375), .A5(
        key_round[91]), .A6(n377), .Y(n56) );
  AO222X1_HVT U44 ( .A1(keyout[90]), .A2(n586), .A3(key[90]), .A4(n309), .A5(
        key_round[90]), .A6(n807), .Y(n57) );
  AO222X1_HVT U45 ( .A1(keyout[89]), .A2(n585), .A3(key[89]), .A4(n773), .A5(
        key_round[89]), .A6(n516), .Y(n58) );
  AO222X1_HVT U47 ( .A1(keyout[87]), .A2(n594), .A3(key[87]), .A4(n773), .A5(
        key_round[87]), .A6(n312), .Y(n60) );
  AO222X1_HVT U48 ( .A1(keyout[86]), .A2(n298), .A3(key[86]), .A4(n772), .A5(
        key_round[86]), .A6(n332), .Y(n61) );
  AO222X1_HVT U49 ( .A1(keyout[85]), .A2(n589), .A3(key[85]), .A4(n376), .A5(
        key_round[85]), .A6(n806), .Y(n62) );
  AO222X1_HVT U51 ( .A1(keyout[83]), .A2(n490), .A3(key[83]), .A4(n782), .A5(
        key_round[83]), .A6(n808), .Y(n64) );
  AO222X1_HVT U52 ( .A1(keyout[82]), .A2(n586), .A3(key[82]), .A4(n773), .A5(
        key_round[82]), .A6(n808), .Y(n65) );
  AO222X1_HVT U53 ( .A1(keyout[81]), .A2(n595), .A3(key[81]), .A4(n772), .A5(
        key_round[81]), .A6(n332), .Y(n66) );
  AO222X1_HVT U54 ( .A1(keyout[80]), .A2(n582), .A3(key[80]), .A4(n783), .A5(
        key_round[80]), .A6(n516), .Y(n67) );
  AO222X1_HVT U58 ( .A1(keyout[76]), .A2(n598), .A3(key[76]), .A4(n386), .A5(
        key_round[76]), .A6(n355), .Y(n71) );
  AO222X1_HVT U59 ( .A1(keyout[75]), .A2(n298), .A3(key[75]), .A4(n777), .A5(
        key_round[75]), .A6(n311), .Y(n72) );
  AO222X1_HVT U60 ( .A1(keyout[74]), .A2(n585), .A3(key[74]), .A4(n768), .A5(
        key_round[74]), .A6(n806), .Y(n73) );
  AO222X1_HVT U61 ( .A1(keyout[73]), .A2(n584), .A3(key[73]), .A4(n765), .A5(
        key_round[73]), .A6(n516), .Y(n74) );
  AO222X1_HVT U63 ( .A1(keyout[71]), .A2(n321), .A3(key[71]), .A4(n767), .A5(
        key_round[71]), .A6(n340), .Y(n76) );
  AO222X1_HVT U64 ( .A1(keyout[70]), .A2(n593), .A3(key[70]), .A4(n797), .A5(
        key_round[70]), .A6(n808), .Y(n77) );
  AO222X1_HVT U65 ( .A1(keyout[69]), .A2(n578), .A3(key[69]), .A4(n796), .A5(
        key_round[69]), .A6(n806), .Y(n78) );
  AO222X1_HVT U66 ( .A1(keyout[68]), .A2(n579), .A3(key[68]), .A4(n795), .A5(
        key_round[68]), .A6(n332), .Y(n79) );
  AO222X1_HVT U67 ( .A1(keyout[67]), .A2(n588), .A3(key[67]), .A4(n781), .A5(
        key_round[67]), .A6(n808), .Y(n80) );
  AO222X1_HVT U69 ( .A1(keyout[65]), .A2(n578), .A3(key[65]), .A4(n779), .A5(
        key_round[65]), .A6(n806), .Y(n82) );
  AO222X1_HVT U71 ( .A1(keyout[63]), .A2(n594), .A3(key[63]), .A4(n789), .A5(
        key_round[63]), .A6(n516), .Y(n84) );
  AO222X1_HVT U72 ( .A1(keyout[62]), .A2(n577), .A3(key[62]), .A4(n786), .A5(
        key_round[62]), .A6(n806), .Y(n85) );
  AO222X1_HVT U73 ( .A1(keyout[61]), .A2(n594), .A3(key[61]), .A4(n785), .A5(
        key_round[61]), .A6(n311), .Y(n86) );
  AO222X1_HVT U74 ( .A1(keyout[60]), .A2(n597), .A3(key[60]), .A4(n376), .A5(
        key_round[60]), .A6(n377), .Y(n87) );
  AO222X1_HVT U75 ( .A1(keyout[59]), .A2(n578), .A3(key[59]), .A4(n376), .A5(
        key_round[59]), .A6(n516), .Y(n88) );
  AO222X1_HVT U76 ( .A1(keyout[58]), .A2(n597), .A3(key[58]), .A4(n782), .A5(
        key_round[58]), .A6(n313), .Y(n89) );
  AO222X1_HVT U79 ( .A1(keyout[55]), .A2(n390), .A3(key[55]), .A4(n772), .A5(
        key_round[55]), .A6(n812), .Y(n92) );
  AO222X1_HVT U81 ( .A1(keyout[53]), .A2(n298), .A3(key[53]), .A4(n771), .A5(
        key_round[53]), .A6(n806), .Y(n94) );
  AO222X1_HVT U82 ( .A1(keyout[52]), .A2(n306), .A3(key[52]), .A4(n770), .A5(
        key_round[52]), .A6(n332), .Y(n95) );
  AO222X1_HVT U83 ( .A1(keyout[51]), .A2(n583), .A3(key[51]), .A4(n782), .A5(
        key_round[51]), .A6(n806), .Y(n96) );
  AO222X1_HVT U85 ( .A1(keyout[49]), .A2(n551), .A3(key[49]), .A4(n772), .A5(
        key_round[49]), .A6(n807), .Y(n98) );
  AO222X1_HVT U86 ( .A1(keyout[48]), .A2(n588), .A3(key[48]), .A4(n307), .A5(
        key_round[48]), .A6(n807), .Y(n99) );
  AO222X1_HVT U89 ( .A1(keyout[45]), .A2(n587), .A3(key[45]), .A4(n791), .A5(
        key_round[45]), .A6(n312), .Y(n102) );
  AO222X1_HVT U91 ( .A1(keyout[43]), .A2(n301), .A3(key[43]), .A4(n309), .A5(
        key_round[43]), .A6(n355), .Y(n104) );
  AO222X1_HVT U93 ( .A1(keyout[41]), .A2(n588), .A3(key[41]), .A4(n782), .A5(
        key_round[41]), .A6(n332), .Y(n106) );
  AO222X1_HVT U95 ( .A1(keyout[39]), .A2(n594), .A3(key[39]), .A4(n791), .A5(
        key_round[39]), .A6(n516), .Y(n108) );
  AO222X1_HVT U96 ( .A1(keyout[38]), .A2(n482), .A3(key[38]), .A4(n777), .A5(
        key_round[38]), .A6(n807), .Y(n109) );
  AO222X1_HVT U97 ( .A1(keyout[37]), .A2(n587), .A3(key[37]), .A4(n302), .A5(
        key_round[37]), .A6(n808), .Y(n110) );
  AO222X1_HVT U98 ( .A1(keyout[36]), .A2(n583), .A3(key[36]), .A4(n765), .A5(
        key_round[36]), .A6(n377), .Y(n111) );
  AO222X1_HVT U101 ( .A1(keyout[33]), .A2(n580), .A3(key[33]), .A4(n777), .A5(
        key_round[33]), .A6(n806), .Y(n114) );
  AO222X1_HVT U102 ( .A1(keyout[32]), .A2(n580), .A3(key[32]), .A4(n769), .A5(
        key_round[32]), .A6(n808), .Y(n115) );
  AO222X1_HVT U103 ( .A1(keyout[31]), .A2(n551), .A3(key[31]), .A4(n800), .A5(
        n679), .A6(n807), .Y(n116) );
  AO222X1_HVT U105 ( .A1(keyout[29]), .A2(n588), .A3(key[29]), .A4(n798), .A5(
        key_round[29]), .A6(n806), .Y(n118) );
  AO222X1_HVT U106 ( .A1(keyout[28]), .A2(n594), .A3(key[28]), .A4(n797), .A5(
        n702), .A6(n807), .Y(n119) );
  AO222X1_HVT U107 ( .A1(keyout[27]), .A2(n584), .A3(key[27]), .A4(n796), .A5(
        key_round[27]), .A6(n516), .Y(n120) );
  AO222X1_HVT U110 ( .A1(keyout[24]), .A2(n582), .A3(key[24]), .A4(n780), .A5(
        key_round[24]), .A6(n810), .Y(n123) );
  AO222X1_HVT U111 ( .A1(keyout[23]), .A2(n585), .A3(key[23]), .A4(n779), .A5(
        n754), .A6(n807), .Y(n124) );
  AO222X1_HVT U112 ( .A1(keyout[22]), .A2(n597), .A3(key[22]), .A4(n778), .A5(
        key_round[22]), .A6(n804), .Y(n125) );
  AO222X1_HVT U114 ( .A1(keyout[20]), .A2(n583), .A3(key[20]), .A4(n769), .A5(
        key_round[20]), .A6(n804), .Y(n127) );
  AO222X1_HVT U115 ( .A1(keyout[19]), .A2(n586), .A3(key[19]), .A4(n790), .A5(
        n622), .A6(n804), .Y(n128) );
  AO222X1_HVT U117 ( .A1(keyout[17]), .A2(n579), .A3(key[17]), .A4(n780), .A5(
        n678), .A6(n804), .Y(n130) );
  AO222X1_HVT U119 ( .A1(keyout[15]), .A2(n588), .A3(key[15]), .A4(n789), .A5(
        key_round[15]), .A6(n804), .Y(n132) );
  AO222X1_HVT U121 ( .A1(keyout[13]), .A2(n595), .A3(key[13]), .A4(n785), .A5(
        key_round[13]), .A6(n804), .Y(n134) );
  AO222X1_HVT U122 ( .A1(keyout[12]), .A2(n597), .A3(key[12]), .A4(n784), .A5(
        n689), .A6(n804), .Y(n135) );
  AO222X1_HVT U124 ( .A1(keyout[10]), .A2(n433), .A3(key[10]), .A4(n770), .A5(
        key_round[10]), .A6(n804), .Y(n137) );
  AO222X1_HVT U126 ( .A1(keyout[8]), .A2(n598), .A3(key[8]), .A4(n800), .A5(
        key_round[8]), .A6(n803), .Y(n139) );
  AO222X1_HVT U127 ( .A1(keyout[7]), .A2(n582), .A3(key[7]), .A4(n376), .A5(
        n602), .A6(n803), .Y(n140) );
  AO222X1_HVT U128 ( .A1(keyout[6]), .A2(n577), .A3(key[6]), .A4(n799), .A5(
        key_round[6]), .A6(n803), .Y(n141) );
  AO222X1_HVT U130 ( .A1(keyout[4]), .A2(n390), .A3(key[4]), .A4(n797), .A5(
        n613), .A6(n803), .Y(n143) );
  AO222X1_HVT U131 ( .A1(keyout[3]), .A2(n582), .A3(key[3]), .A4(n796), .A5(
        n631), .A6(n803), .Y(n144) );
  AO222X1_HVT U132 ( .A1(keyout[2]), .A2(n579), .A3(key[2]), .A4(n782), .A5(
        key_round[2]), .A6(n803), .Y(n145) );
  AO222X1_HVT U134 ( .A1(keyout[0]), .A2(n581), .A3(key[0]), .A4(n375), .A5(
        key_round[0]), .A6(n803), .Y(n147) );
  AO222X1_HVT U135 ( .A1(cipher_text[127]), .A2(n598), .A3(adk_out0[127]), 
        .A4(n773), .A5(n629), .A6(n803), .Y(n148) );
  AO222X1_HVT U136 ( .A1(cipher_text[126]), .A2(n596), .A3(adk_out0[126]), 
        .A4(n307), .A5(adk_in[126]), .A6(n808), .Y(n149) );
  AO222X1_HVT U137 ( .A1(cipher_text[125]), .A2(n298), .A3(adk_out0[125]), 
        .A4(n773), .A5(adk_in[125]), .A6(n809), .Y(n150) );
  AO222X1_HVT U140 ( .A1(cipher_text[122]), .A2(n580), .A3(adk_out0[122]), 
        .A4(n780), .A5(n315), .A6(n489), .Y(n153) );
  AO222X1_HVT U142 ( .A1(cipher_text[120]), .A2(n306), .A3(adk_out0[120]), 
        .A4(n772), .A5(adk_in[120]), .A6(n813), .Y(n155) );
  AO222X1_HVT U143 ( .A1(cipher_text[119]), .A2(n594), .A3(adk_out0[119]), 
        .A4(n296), .A5(adk_in[119]), .A6(n804), .Y(n156) );
  AO222X1_HVT U144 ( .A1(cipher_text[118]), .A2(n586), .A3(adk_out0[118]), 
        .A4(n771), .A5(adk_in[118]), .A6(n489), .Y(n157) );
  AO222X1_HVT U146 ( .A1(cipher_text[116]), .A2(n433), .A3(adk_out0[116]), 
        .A4(n769), .A5(n740), .A6(n310), .Y(n159) );
  AO222X1_HVT U148 ( .A1(cipher_text[114]), .A2(n577), .A3(adk_out0[114]), 
        .A4(n799), .A5(adk_in[114]), .A6(n489), .Y(n161) );
  AO222X1_HVT U149 ( .A1(cipher_text[113]), .A2(n593), .A3(adk_out0[113]), 
        .A4(n798), .A5(n728), .A6(n313), .Y(n162) );
  AO222X1_HVT U152 ( .A1(cipher_text[110]), .A2(n582), .A3(adk_out0[110]), 
        .A4(n795), .A5(adk_in[110]), .A6(n284), .Y(n165) );
  AO222X1_HVT U153 ( .A1(cipher_text[109]), .A2(n390), .A3(adk_out0[109]), 
        .A4(n765), .A5(n328), .A6(n310), .Y(n166) );
  AO222X1_HVT U155 ( .A1(cipher_text[107]), .A2(n580), .A3(adk_out0[107]), 
        .A4(n790), .A5(n714), .A6(n813), .Y(n168) );
  AO222X1_HVT U156 ( .A1(cipher_text[106]), .A2(n580), .A3(adk_out0[106]), 
        .A4(n787), .A5(n710), .A6(n419), .Y(n169) );
  AO222X1_HVT U157 ( .A1(cipher_text[105]), .A2(n593), .A3(adk_out0[105]), 
        .A4(n780), .A5(n698), .A6(n573), .Y(n170) );
  AO222X1_HVT U158 ( .A1(cipher_text[104]), .A2(n596), .A3(adk_out0[104]), 
        .A4(n296), .A5(adk_in[104]), .A6(n489), .Y(n171) );
  AO222X1_HVT U161 ( .A1(cipher_text[101]), .A2(n551), .A3(adk_out0[101]), 
        .A4(n780), .A5(adk_in[101]), .A6(n573), .Y(n174) );
  AO222X1_HVT U163 ( .A1(cipher_text[99]), .A2(n598), .A3(adk_out0[99]), .A4(
        n786), .A5(n656), .A6(n303), .Y(n176) );
  AO222X1_HVT U164 ( .A1(cipher_text[98]), .A2(n585), .A3(adk_out0[98]), .A4(
        n785), .A5(n801), .A6(n332), .Y(n177) );
  AO222X1_HVT U165 ( .A1(cipher_text[97]), .A2(n585), .A3(adk_out0[97]), .A4(
        n771), .A5(n644), .A6(n573), .Y(n178) );
  AO222X1_HVT U166 ( .A1(cipher_text[96]), .A2(n595), .A3(adk_out0[96]), .A4(
        n770), .A5(adk_in[96]), .A6(n303), .Y(n179) );
  AO222X1_HVT U167 ( .A1(cipher_text[95]), .A2(n597), .A3(adk_out0[95]), .A4(
        n769), .A5(adk_in[95]), .A6(n813), .Y(n180) );
  AO222X1_HVT U169 ( .A1(cipher_text[93]), .A2(n321), .A3(adk_out0[93]), .A4(
        n799), .A5(adk_in[93]), .A6(n813), .Y(n182) );
  AO222X1_HVT U171 ( .A1(cipher_text[91]), .A2(n584), .A3(adk_out0[91]), .A4(
        n779), .A5(n617), .A6(n489), .Y(n184) );
  AO222X1_HVT U174 ( .A1(cipher_text[88]), .A2(n433), .A3(adk_out0[88]), .A4(
        n779), .A5(adk_in[88]), .A6(n297), .Y(n187) );
  AO222X1_HVT U178 ( .A1(cipher_text[84]), .A2(n598), .A3(adk_out0[84]), .A4(
        n765), .A5(n724), .A6(n814), .Y(n191) );
  AO222X1_HVT U180 ( .A1(cipher_text[82]), .A2(n587), .A3(adk_out0[82]), .A4(
        n790), .A5(n641), .A6(n813), .Y(n193) );
  AO222X1_HVT U181 ( .A1(cipher_text[81]), .A2(n306), .A3(adk_out0[81]), .A4(
        n386), .A5(n649), .A6(n516), .Y(n194) );
  AO222X1_HVT U182 ( .A1(cipher_text[80]), .A2(n594), .A3(adk_out0[80]), .A4(
        n787), .A5(adk_in[80]), .A6(n573), .Y(n195) );
  AO222X1_HVT U183 ( .A1(cipher_text[79]), .A2(n576), .A3(adk_out0[79]), .A4(
        n792), .A5(n632), .A6(n813), .Y(n196) );
  AO222X1_HVT U184 ( .A1(cipher_text[78]), .A2(n598), .A3(adk_out0[78]), .A4(
        n789), .A5(adk_in[78]), .A6(n297), .Y(n197) );
  AO222X1_HVT U185 ( .A1(cipher_text[77]), .A2(n585), .A3(adk_out0[77]), .A4(
        n786), .A5(adk_in[77]), .A6(n313), .Y(n198) );
  AO222X1_HVT U187 ( .A1(cipher_text[75]), .A2(n304), .A3(adk_out0[75]), .A4(
        n787), .A5(n664), .A6(n303), .Y(n200) );
  AO222X1_HVT U189 ( .A1(cipher_text[73]), .A2(n596), .A3(adk_out0[73]), .A4(
        n789), .A5(n676), .A6(n489), .Y(n202) );
  AO222X1_HVT U190 ( .A1(cipher_text[72]), .A2(n482), .A3(adk_out0[72]), .A4(
        n786), .A5(adk_in[72]), .A6(n419), .Y(n203) );
  AO222X1_HVT U191 ( .A1(cipher_text[71]), .A2(n598), .A3(adk_out0[71]), .A4(
        n785), .A5(n323), .A6(n803), .Y(n204) );
  AO222X1_HVT U193 ( .A1(cipher_text[69]), .A2(n597), .A3(adk_out0[69]), .A4(
        n781), .A5(adk_in[69]), .A6(n573), .Y(n206) );
  AO222X1_HVT U194 ( .A1(cipher_text[68]), .A2(n306), .A3(adk_out0[68]), .A4(
        n778), .A5(n742), .A6(n300), .Y(n207) );
  AO222X1_HVT U196 ( .A1(cipher_text[66]), .A2(n577), .A3(adk_out0[66]), .A4(
        n798), .A5(n642), .A6(n488), .Y(n209) );
  AO222X1_HVT U197 ( .A1(cipher_text[65]), .A2(n579), .A3(adk_out0[65]), .A4(
        n765), .A5(adk_in[65]), .A6(n814), .Y(n210) );
  AO222X1_HVT U201 ( .A1(cipher_text[61]), .A2(n595), .A3(adk_out0[61]), .A4(
        n772), .A5(n317), .A6(n813), .Y(n214) );
  AO222X1_HVT U202 ( .A1(cipher_text[60]), .A2(n597), .A3(adk_out0[60]), .A4(
        n783), .A5(n752), .A6(n573), .Y(n215) );
  AO222X1_HVT U204 ( .A1(cipher_text[58]), .A2(n598), .A3(adk_out0[58]), .A4(
        n800), .A5(adk_in[58]), .A6(n813), .Y(n217) );
  AO222X1_HVT U205 ( .A1(cipher_text[57]), .A2(n582), .A3(adk_out0[57]), .A4(
        n799), .A5(n696), .A6(n814), .Y(n218) );
  AO222X1_HVT U206 ( .A1(cipher_text[56]), .A2(n584), .A3(adk_out0[56]), .A4(
        n798), .A5(adk_in[56]), .A6(n809), .Y(n219) );
  AO222X1_HVT U207 ( .A1(cipher_text[55]), .A2(n583), .A3(adk_out0[55]), .A4(
        n797), .A5(adk_in[55]), .A6(n809), .Y(n220) );
  AO222X1_HVT U208 ( .A1(cipher_text[54]), .A2(n593), .A3(adk_out0[54]), .A4(
        n779), .A5(n416), .A6(n310), .Y(n221) );
  AO222X1_HVT U209 ( .A1(cipher_text[53]), .A2(n596), .A3(adk_out0[53]), .A4(
        n778), .A5(adk_in[53]), .A6(n297), .Y(n222) );
  AO222X1_HVT U210 ( .A1(cipher_text[52]), .A2(n588), .A3(adk_out0[52]), .A4(
        n776), .A5(n734), .A6(n813), .Y(n223) );
  AO222X1_HVT U211 ( .A1(cipher_text[51]), .A2(n433), .A3(adk_out0[51]), .A4(
        n787), .A5(n658), .A6(n488), .Y(n224) );
  AO222X1_HVT U213 ( .A1(cipher_text[49]), .A2(n583), .A3(adk_out0[49]), .A4(
        n789), .A5(n746), .A6(n810), .Y(n226) );
  AO222X1_HVT U214 ( .A1(cipher_text[48]), .A2(n581), .A3(adk_out0[48]), .A4(
        n786), .A5(adk_in[48]), .A6(n809), .Y(n227) );
  AO222X1_HVT U215 ( .A1(cipher_text[47]), .A2(n579), .A3(adk_out0[47]), .A4(
        n785), .A5(adk_in[47]), .A6(n300), .Y(n228) );
  AO222X1_HVT U216 ( .A1(cipher_text[46]), .A2(n589), .A3(adk_out0[46]), .A4(
        n790), .A5(adk_in[46]), .A6(n812), .Y(n229) );
  AO222X1_HVT U217 ( .A1(cipher_text[45]), .A2(n390), .A3(adk_out0[45]), .A4(
        n765), .A5(n611), .A6(n297), .Y(n230) );
  AO222X1_HVT U219 ( .A1(cipher_text[43]), .A2(n583), .A3(adk_out0[43]), .A4(
        n790), .A5(n652), .A6(n297), .Y(n232) );
  AO222X1_HVT U220 ( .A1(cipher_text[42]), .A2(n597), .A3(adk_out0[42]), .A4(
        n309), .A5(n610), .A6(n419), .Y(n233) );
  AO222X1_HVT U221 ( .A1(cipher_text[41]), .A2(n597), .A3(adk_out0[41]), .A4(
        n787), .A5(n606), .A6(n488), .Y(n234) );
  AO222X1_HVT U222 ( .A1(cipher_text[40]), .A2(n576), .A3(adk_out0[40]), .A4(
        n795), .A5(adk_in[40]), .A6(n811), .Y(n235) );
  AO222X1_HVT U223 ( .A1(cipher_text[39]), .A2(n301), .A3(adk_out0[39]), .A4(
        n789), .A5(n744), .A6(n809), .Y(n236) );
  AO222X1_HVT U225 ( .A1(cipher_text[37]), .A2(n598), .A3(adk_out0[37]), .A4(
        n785), .A5(adk_in[37]), .A6(n812), .Y(n238) );
  AO222X1_HVT U226 ( .A1(cipher_text[36]), .A2(n589), .A3(adk_out0[36]), .A4(
        n784), .A5(n760), .A6(n811), .Y(n239) );
  AO222X1_HVT U227 ( .A1(cipher_text[35]), .A2(n551), .A3(adk_out0[35]), .A4(
        n375), .A5(n674), .A6(n811), .Y(n240) );
  AO222X1_HVT U228 ( .A1(cipher_text[34]), .A2(n593), .A3(adk_out0[34]), .A4(
        n787), .A5(adk_in[34]), .A6(n809), .Y(n241) );
  AO222X1_HVT U230 ( .A1(cipher_text[32]), .A2(n596), .A3(adk_out0[32]), .A4(
        n769), .A5(adk_in[32]), .A6(n811), .Y(n243) );
  AO222X1_HVT U231 ( .A1(cipher_text[31]), .A2(n587), .A3(adk_out0[31]), .A4(
        n800), .A5(adk_in[31]), .A6(n811), .Y(n244) );
  AO222X1_HVT U232 ( .A1(cipher_text[30]), .A2(n551), .A3(adk_out0[30]), .A4(
        n799), .A5(adk_in[30]), .A6(n810), .Y(n245) );
  AO222X1_HVT U233 ( .A1(cipher_text[29]), .A2(n583), .A3(adk_out0[29]), .A4(
        n798), .A5(n623), .A6(n284), .Y(n246) );
  AO222X1_HVT U234 ( .A1(cipher_text[28]), .A2(n588), .A3(adk_out0[28]), .A4(
        n797), .A5(n687), .A6(n488), .Y(n247) );
  AO222X1_HVT U235 ( .A1(cipher_text[27]), .A2(n304), .A3(adk_out0[27]), .A4(
        n796), .A5(n685), .A6(n340), .Y(n248) );
  AO222X1_HVT U236 ( .A1(cipher_text[26]), .A2(n594), .A3(adk_out0[26]), .A4(
        n795), .A5(n353), .A6(n377), .Y(n249) );
  AO222X1_HVT U237 ( .A1(cipher_text[25]), .A2(n585), .A3(adk_out0[25]), .A4(
        n781), .A5(n660), .A6(n812), .Y(n250) );
  AO222X1_HVT U238 ( .A1(cipher_text[24]), .A2(n577), .A3(adk_out0[24]), .A4(
        n780), .A5(adk_in[24]), .A6(n809), .Y(n251) );
  AO222X1_HVT U240 ( .A1(cipher_text[22]), .A2(n595), .A3(adk_out0[22]), .A4(
        n767), .A5(adk_in[22]), .A6(n300), .Y(n253) );
  AO222X1_HVT U242 ( .A1(cipher_text[20]), .A2(n596), .A3(adk_out0[20]), .A4(
        n773), .A5(n634), .A6(n809), .Y(n255) );
  AO222X1_HVT U243 ( .A1(cipher_text[19]), .A2(n594), .A3(adk_out0[19]), .A4(
        n772), .A5(n672), .A6(n340), .Y(n256) );
  AO222X1_HVT U244 ( .A1(cipher_text[18]), .A2(n584), .A3(adk_out0[18]), .A4(
        n783), .A5(adk_in[18]), .A6(n310), .Y(n257) );
  AO222X1_HVT U245 ( .A1(cipher_text[17]), .A2(n301), .A3(adk_out0[17]), .A4(
        n782), .A5(n730), .A6(n340), .Y(n258) );
  AO222X1_HVT U247 ( .A1(cipher_text[15]), .A2(n588), .A3(adk_out0[15]), .A4(
        n771), .A5(n357), .A6(n303), .Y(n260) );
  AO222X1_HVT U249 ( .A1(cipher_text[13]), .A2(n595), .A3(adk_out0[13]), .A4(
        n769), .A5(adk_in[13]), .A6(n381), .Y(n262) );
  AO222X1_HVT U251 ( .A1(cipher_text[11]), .A2(n301), .A3(adk_out0[11]), .A4(
        n799), .A5(n704), .A6(n811), .Y(n264) );
  AO222X1_HVT U252 ( .A1(cipher_text[10]), .A2(n301), .A3(adk_out0[10]), .A4(
        n798), .A5(n626), .A6(n377), .Y(n265) );
  AO222X1_HVT U253 ( .A1(cipher_text[9]), .A2(n583), .A3(adk_out0[9]), .A4(
        n797), .A5(n748), .A6(n809), .Y(n266) );
  AO222X1_HVT U254 ( .A1(cipher_text[8]), .A2(n298), .A3(adk_out0[8]), .A4(
        n796), .A5(adk_in[8]), .A6(n340), .Y(n267) );
  AO222X1_HVT U256 ( .A1(cipher_text[6]), .A2(n589), .A3(adk_out0[6]), .A4(
        n781), .A5(adk_in[6]), .A6(n488), .Y(n269) );
  AO222X1_HVT U258 ( .A1(cipher_text[4]), .A2(n597), .A3(adk_out0[4]), .A4(
        n779), .A5(n662), .A6(n488), .Y(n271) );
  AO222X1_HVT U259 ( .A1(cipher_text[3]), .A2(n586), .A3(adk_out0[3]), .A4(
        n796), .A5(n666), .A6(n340), .Y(n272) );
  AO222X1_HVT U260 ( .A1(cipher_text[2]), .A2(n596), .A3(adk_out0[2]), .A4(
        n771), .A5(n325), .A6(n812), .Y(n273) );
  AO222X1_HVT U261 ( .A1(cipher_text[1]), .A2(n585), .A3(adk_out0[1]), .A4(
        n796), .A5(n706), .A6(n488), .Y(n274) );
  AO222X1_HVT U262 ( .A1(cipher_text[0]), .A2(n582), .A3(adk_out0[0]), .A4(
        n795), .A5(adk_in[0]), .A6(n812), .Y(n275) );
  AO22X1_HVT U265 ( .A1(n12), .A2(n342), .A3(n13), .A4(n361), .Y(n276) );
  AND2X1_HVT U266 ( .A1(n14), .A2(n568), .Y(n13) );
  AO22X1_HVT U267 ( .A1(n361), .A2(n517), .A3(n14), .A4(n569), .Y(n277) );
  AO22X1_HVT U268 ( .A1(n12), .A2(n358), .A3(n16), .A4(n342), .Y(n278) );
  AND2X1_HVT U269 ( .A1(n361), .A2(n14), .Y(n16) );
  AND2X1_HVT U270 ( .A1(n826), .A2(n817), .Y(n14) );
  DFFX1_HVT \adk_in_reg[110]  ( .D(n165), .CLK(clk), .Q(adk_in[110]) );
  DFFX1_HVT \adk_in_reg[66]  ( .D(n209), .CLK(clk), .Q(n642) );
  DFFX1_HVT \adk_in_reg[98]  ( .D(n177), .CLK(clk), .Q(n801) );
  DFFX1_HVT \adk_in_reg[86]  ( .D(n189), .CLK(clk), .Q(adk_in[86]) );
  DFFX1_HVT \adk_in_reg[54]  ( .D(n221), .CLK(clk), .Q(adk_in[54]), .QN(n415)
         );
  DFFX1_HVT ready_reg ( .D(n19), .CLK(clk), .Q(ready), .QN(n827) );
  DFFX1_HVT \key_round_reg[120]  ( .D(n27), .CLK(clk), .Q(key_round[120]) );
  DFFX1_HVT \key_round_reg[115]  ( .D(n32), .CLK(clk), .Q(key_round[115]) );
  DFFX1_HVT \key_round_reg[119]  ( .D(n28), .CLK(clk), .Q(key_round[119]), 
        .QN(n351) );
  DFFX1_HVT \key_round_reg[106]  ( .D(n287), .CLK(clk), .Q(key_round[106]), 
        .QN(n348) );
  DFFX1_HVT \key_round_reg[100]  ( .D(n47), .CLK(clk), .Q(key_round[100]) );
  DFFX1_HVT \key_round_reg[98]  ( .D(n49), .CLK(clk), .Q(key_round[98]), .QN(
        n547) );
  DFFX1_HVT \key_round_reg[97]  ( .D(n365), .CLK(clk), .Q(key_round[97]) );
  DFFX1_HVT \key_round_reg[104]  ( .D(n43), .CLK(clk), .Q(key_round[104]) );
  DFFX1_HVT \key_round_reg[114]  ( .D(n33), .CLK(clk), .Q(key_round[114]) );
  DFFX1_HVT \key_round_reg[109]  ( .D(n38), .CLK(clk), .Q(key_round[109]), 
        .QN(n455) );
  DFFX1_HVT \key_round_reg[118]  ( .D(n29), .CLK(clk), .Q(key_round[118]), 
        .QN(n333) );
  DFFX1_HVT \key_round_reg[108]  ( .D(n39), .CLK(clk), .Q(key_round[108]) );
  DFFX1_HVT \key_round_reg[102]  ( .D(n45), .CLK(clk), .Q(key_round[102]) );
  DFFX1_HVT \key_round_reg[116]  ( .D(n31), .CLK(clk), .Q(key_round[116]) );
  DFFX1_HVT \key_round_reg[111]  ( .D(n36), .CLK(clk), .Q(key_round[111]) );
  DFFX1_HVT \key_round_reg[126]  ( .D(n21), .CLK(clk), .Q(key_round[126]), 
        .QN(n339) );
  DFFX1_HVT \key_round_reg[117]  ( .D(n30), .CLK(clk), .Q(key_round[117]) );
  DFFX1_HVT \key_round_reg[99]  ( .D(n48), .CLK(clk), .Q(key_round[99]) );
  DFFX1_HVT \key_round_reg[61]  ( .D(n86), .CLK(clk), .Q(key_round[61]) );
  DFFX1_HVT \key_round_reg[96]  ( .D(n286), .CLK(clk), .Q(key_round[96]), .QN(
        n374) );
  DFFX1_HVT \key_round_reg[113]  ( .D(n34), .CLK(clk), .Q(key_round[113]) );
  DFFX1_HVT \key_round_reg[105]  ( .D(n42), .CLK(clk), .Q(key_round[105]), 
        .QN(n345) );
  DFFX1_HVT \key_round_reg[103]  ( .D(n44), .CLK(clk), .Q(key_round[103]), 
        .QN(n432) );
  DFFX1_HVT \key_round_reg[112]  ( .D(n35), .CLK(clk), .Q(key_round[112]), 
        .QN(n479) );
  DFFX1_HVT \key_round_reg[88]  ( .D(n59), .CLK(clk), .Q(key_round[88]), .QN(
        n560) );
  DFFX1_HVT \key_round_reg[22]  ( .D(n125), .CLK(clk), .Q(key_round[22]) );
  DFFX1_HVT \key_round_reg[101]  ( .D(n46), .CLK(clk), .Q(key_round[101]), 
        .QN(n544) );
  DFFX1_HVT \key_round_reg[2]  ( .D(n145), .CLK(clk), .Q(key_round[2]) );
  DFFX1_HVT \key_round_reg[107]  ( .D(n40), .CLK(clk), .Q(key_round[107]), 
        .QN(n452) );
  DFFX1_HVT \key_round_reg[62]  ( .D(n85), .CLK(clk), .Q(key_round[62]) );
  DFFX1_HVT \key_round_reg[66]  ( .D(n290), .CLK(clk), .Q(key_round[66]), .QN(
        n511) );
  DFFX1_HVT \key_round_reg[110]  ( .D(n37), .CLK(clk), .Q(key_round[110]) );
  DFFX1_HVT \key_round_reg[82]  ( .D(n65), .CLK(clk), .Q(key_round[82]) );
  DFFX1_HVT \key_round_reg[0]  ( .D(n147), .CLK(clk), .Q(key_round[0]) );
  DFFX1_HVT \key_round_reg[8]  ( .D(n139), .CLK(clk), .Q(key_round[8]) );
  DFFX1_HVT \key_round_reg[89]  ( .D(n58), .CLK(clk), .Q(key_round[89]) );
  DFFX1_HVT \key_round_reg[60]  ( .D(n87), .CLK(clk), .Q(key_round[60]) );
  DFFX1_HVT \key_round_reg[63]  ( .D(n84), .CLK(clk), .Q(key_round[63]) );
  DFFX1_HVT \key_round_reg[59]  ( .D(n88), .CLK(clk), .Q(key_round[59]) );
  DFFX1_HVT \key_round_reg[39]  ( .D(n108), .CLK(clk), .Q(key_round[39]) );
  DFFX1_HVT \key_round_reg[121]  ( .D(n26), .CLK(clk), .Q(key_round[121]) );
  DFFX1_HVT \key_round_reg[68]  ( .D(n79), .CLK(clk), .Q(key_round[68]) );
  DFFX1_HVT \key_round_reg[57]  ( .D(n90), .CLK(clk), .Q(key_round[57]), .QN(
        n550) );
  DFFX1_HVT \key_round_reg[122]  ( .D(n25), .CLK(clk), .Q(key_round[122]) );
  DFFX1_HVT \key_round_reg[76]  ( .D(n71), .CLK(clk), .Q(key_round[76]) );
  DFFX1_HVT \key_round_reg[90]  ( .D(n57), .CLK(clk), .Q(key_round[90]) );
  DFFX1_HVT \key_round_reg[92]  ( .D(n55), .CLK(clk), .Q(key_round[92]) );
  DFFX1_HVT \key_round_reg[124]  ( .D(n23), .CLK(clk), .Q(key_round[124]) );
  DFFX1_HVT \key_round_reg[58]  ( .D(n89), .CLK(clk), .Q(key_round[58]) );
  DFFX1_HVT \key_round_reg[91]  ( .D(n56), .CLK(clk), .Q(key_round[91]) );
  DFFX1_HVT \key_round_reg[123]  ( .D(n24), .CLK(clk), .Q(key_round[123]) );
  DFFX1_HVT \key_round_reg[48]  ( .D(n99), .CLK(clk), .Q(key_round[48]) );
  DFFX1_HVT \key_round_reg[45]  ( .D(n102), .CLK(clk), .Q(key_round[45]) );
  DFFX1_HVT \key_round_reg[67]  ( .D(n80), .CLK(clk), .Q(key_round[67]) );
  DFFX1_HVT \key_round_reg[93]  ( .D(n54), .CLK(clk), .Q(key_round[93]) );
  DFFX1_HVT \key_round_reg[51]  ( .D(n96), .CLK(clk), .Q(key_round[51]) );
  DFFX1_HVT \key_round_reg[125]  ( .D(n22), .CLK(clk), .Q(key_round[125]) );
  DFFX1_HVT \key_round_reg[127]  ( .D(n20), .CLK(clk), .Q(key_round[127]) );
  DFFX1_HVT \key_round_reg[85]  ( .D(n62), .CLK(clk), .Q(key_round[85]) );
  DFFX1_HVT \key_round_reg[49]  ( .D(n98), .CLK(clk), .Q(key_round[49]) );
  DFFX1_HVT \key_round_reg[52]  ( .D(n95), .CLK(clk), .Q(key_round[52]) );
  DFFX1_HVT \key_round_reg[80]  ( .D(n67), .CLK(clk), .Q(key_round[80]) );
  DFFX1_HVT \key_round_reg[83]  ( .D(n64), .CLK(clk), .Q(key_round[83]) );
  DFFX1_HVT \key_round_reg[69]  ( .D(n78), .CLK(clk), .Q(key_round[69]) );
  DFFX1_HVT \adk_in_reg[22]  ( .D(n253), .CLK(clk), .Q(adk_in[22]) );
  DFFX1_HVT \adk_in_reg[126]  ( .D(n149), .CLK(clk), .Q(adk_in[126]) );
  DFFX1_HVT \round_number_reg[2]  ( .D(n276), .CLK(clk), .Q(round_number[2]), 
        .QN(n4) );
  DFFX1_HVT \adk_in_reg[46]  ( .D(n229), .CLK(clk), .Q(adk_in[46]) );
  DFFX1_HVT \adk_in_reg[62]  ( .D(n213), .CLK(clk), .Q(adk_in[62]) );
  DFFX1_HVT \adk_in_reg[38]  ( .D(n237), .CLK(clk), .Q(adk_in[38]) );
  DFFX1_HVT \adk_in_reg[30]  ( .D(n245), .CLK(clk), .Q(adk_in[30]) );
  AND4X1_HVT U277 ( .A1(n574), .A2(n567), .A3(n505), .A4(n763), .Y(n491) );
  INVX1_HVT U278 ( .A(n592), .Y(n598) );
  INVX0_HVT U279 ( .A(keyout[66]), .Y(n509) );
  INVX1_HVT U280 ( .A(keyout[103]), .Y(n428) );
  INVX0_HVT U281 ( .A(keyout[56]), .Y(n459) );
  INVX0_HVT U282 ( .A(keyout[47]), .Y(n391) );
  INVX0_HVT U283 ( .A(keyout[26]), .Y(n404) );
  INVX0_HVT U284 ( .A(keyout[9]), .Y(n495) );
  INVX0_HVT U285 ( .A(keyout[5]), .Y(n438) );
  INVX1_HVT U286 ( .A(n650), .Y(n283) );
  OAI222X1_HVT U287 ( .A1(n469), .A2(n474), .A3(n470), .A4(n430), .A5(n758), 
        .A6(n379), .Y(n164) );
  OAI222X1_HVT U288 ( .A1(n474), .A2(n434), .A3(n435), .A4(n436), .A5(n437), 
        .A6(n818), .Y(n216) );
  OAI222X1_HVT U289 ( .A1(n474), .A2(n466), .A3(n467), .A4(n543), .A5(n468), 
        .A6(n383), .Y(n259) );
  OAI222X1_HVT U290 ( .A1(n334), .A2(n530), .A3(n335), .A4(n402), .A5(n336), 
        .A6(n431), .Y(n280) );
  AND2X1_HVT U291 ( .A1(n567), .A2(n505), .Y(n281) );
  INVX1_HVT U292 ( .A(n534), .Y(n284) );
  INVX1_HVT U293 ( .A(n591), .Y(n596) );
  INVX1_HVT U294 ( .A(n388), .Y(n321) );
  INVX0_HVT U295 ( .A(n778), .Y(n464) );
  INVX0_HVT U296 ( .A(n770), .Y(n533) );
  INVX1_HVT U297 ( .A(n447), .Y(n282) );
  OAI222X1_HVT U298 ( .A1(n473), .A2(n397), .A3(n398), .A4(n512), .A5(n399), 
        .A6(n367), .Y(n208) );
  AO222X1_HVT U299 ( .A1(n587), .A2(cipher_text[50]), .A3(adk_out0[50]), .A4(
        n778), .A5(adk_in[50]), .A6(n284), .Y(n225) );
  AO222X1_HVT U300 ( .A1(cipher_text[115]), .A2(n321), .A3(adk_out0[115]), 
        .A4(n282), .A5(n283), .A6(n284), .Y(n160) );
  IBUFFX2_HVT U301 ( .A(keyout[64]), .Y(n462) );
  IBUFFX2_HVT U302 ( .A(keyout[79]), .Y(n359) );
  INVX1_HVT U303 ( .A(n482), .Y(n592) );
  INVX1_HVT U304 ( .A(n382), .Y(n774) );
  INVX1_HVT U305 ( .A(n490), .Y(n591) );
  INVX2_HVT U306 ( .A(n802), .Y(n818) );
  INVX1_HVT U307 ( .A(n817), .Y(n808) );
  INVX1_HVT U308 ( .A(n817), .Y(n806) );
  INVX1_HVT U309 ( .A(n817), .Y(n807) );
  INVX1_HVT U310 ( .A(n818), .Y(n804) );
  INVX1_HVT U311 ( .A(n817), .Y(n516) );
  INVX1_HVT U312 ( .A(n777), .Y(n512) );
  INVX1_HVT U313 ( .A(n771), .Y(n436) );
  NBUFFX2_HVT U314 ( .A(n766), .Y(n778) );
  NBUFFX2_HVT U315 ( .A(n490), .Y(n579) );
  NBUFFX2_HVT U316 ( .A(n766), .Y(n769) );
  INVX1_HVT U317 ( .A(n473), .Y(n585) );
  NBUFFX2_HVT U318 ( .A(n792), .Y(n795) );
  INVX1_HVT U319 ( .A(n816), .Y(n812) );
  INVX1_HVT U320 ( .A(n448), .Y(n296) );
  INVX1_HVT U321 ( .A(n800), .Y(n448) );
  INVX0_HVT U322 ( .A(n815), .Y(n813) );
  INVX1_HVT U323 ( .A(n823), .Y(n584) );
  INVX1_HVT U324 ( .A(n331), .Y(n811) );
  INVX1_HVT U325 ( .A(n331), .Y(n809) );
  INVX1_HVT U326 ( .A(n331), .Y(n488) );
  INVX1_HVT U327 ( .A(n342), .Y(n568) );
  INVX1_HVT U328 ( .A(key[57]), .Y(n549) );
  INVX1_HVT U329 ( .A(key[66]), .Y(n510) );
  INVX1_HVT U330 ( .A(key[107]), .Y(n450) );
  INVX1_HVT U331 ( .A(n786), .Y(n451) );
  INVX0_HVT U332 ( .A(keyout[107]), .Y(n449) );
  INVX1_HVT U333 ( .A(key[101]), .Y(n542) );
  INVX0_HVT U334 ( .A(keyout[101]), .Y(n541) );
  INVX1_HVT U335 ( .A(key[88]), .Y(n559) );
  INVX1_HVT U336 ( .A(keyout[88]), .Y(n558) );
  INVX1_HVT U337 ( .A(key[112]), .Y(n478) );
  INVX1_HVT U338 ( .A(keyout[112]), .Y(n477) );
  INVX1_HVT U339 ( .A(key[103]), .Y(n429) );
  INVX1_HVT U340 ( .A(n769), .Y(n430) );
  OAI222X1_HVT U341 ( .A1(n343), .A2(n496), .A3(n344), .A4(n464), .A5(n345), 
        .A6(n562), .Y(n42) );
  INVX1_HVT U342 ( .A(key[105]), .Y(n344) );
  INVX1_HVT U343 ( .A(keyout[105]), .Y(n343) );
  INVX1_HVT U344 ( .A(key[96]), .Y(n373) );
  INVX1_HVT U345 ( .A(keyout[96]), .Y(n372) );
  INVX1_HVT U346 ( .A(key[126]), .Y(n338) );
  INVX1_HVT U347 ( .A(keyout[126]), .Y(n337) );
  INVX1_HVT U348 ( .A(key[109]), .Y(n454) );
  INVX1_HVT U349 ( .A(keyout[109]), .Y(n453) );
  INVX1_HVT U350 ( .A(key[98]), .Y(n546) );
  INVX1_HVT U351 ( .A(keyout[98]), .Y(n545) );
  INVX1_HVT U352 ( .A(key[106]), .Y(n347) );
  INVX1_HVT U353 ( .A(keyout[106]), .Y(n346) );
  INVX1_HVT U354 ( .A(key[119]), .Y(n350) );
  INVX1_HVT U355 ( .A(keyout[119]), .Y(n349) );
  INVX1_HVT U356 ( .A(key[84]), .Y(n536) );
  INVX1_HVT U357 ( .A(key[79]), .Y(n360) );
  NAND2X0_HVT U358 ( .A1(keyout[78]), .A2(n579), .Y(n506) );
  NAND2X0_HVT U359 ( .A1(keyout[77]), .A2(n390), .Y(n525) );
  INVX1_HVT U360 ( .A(key[64]), .Y(n463) );
  INVX1_HVT U361 ( .A(key[56]), .Y(n460) );
  NAND2X0_HVT U362 ( .A1(keyout[54]), .A2(n390), .Y(n518) );
  OAI222X1_HVT U363 ( .A1(n499), .A2(n473), .A3(n500), .A4(n430), .A5(n501), 
        .A6(n556), .Y(n97) );
  INVX1_HVT U364 ( .A(key[50]), .Y(n500) );
  INVX1_HVT U365 ( .A(key[47]), .Y(n392) );
  INVX1_HVT U366 ( .A(key[46]), .Y(n413) );
  INVX1_HVT U367 ( .A(key[44]), .Y(n410) );
  INVX1_HVT U368 ( .A(keyout[44]), .Y(n409) );
  INVX1_HVT U369 ( .A(key[40]), .Y(n442) );
  OAI222X1_HVT U370 ( .A1(n423), .A2(n530), .A3(n424), .A4(n464), .A5(n425), 
        .A6(n379), .Y(n112) );
  INVX1_HVT U371 ( .A(key[35]), .Y(n424) );
  INVX1_HVT U372 ( .A(key[34]), .Y(n421) );
  INVX1_HVT U373 ( .A(key[30]), .Y(n364) );
  INVX1_HVT U374 ( .A(key[26]), .Y(n405) );
  INVX1_HVT U375 ( .A(key[25]), .Y(n476) );
  INVX1_HVT U376 ( .A(key[21]), .Y(n427) );
  INVX1_HVT U377 ( .A(key[18]), .Y(n335) );
  INVX1_HVT U378 ( .A(key[16]), .Y(n370) );
  NAND2X0_HVT U379 ( .A1(keyout[14]), .A2(n304), .Y(n486) );
  INVX1_HVT U380 ( .A(n494), .Y(n387) );
  INVX1_HVT U381 ( .A(key[9]), .Y(n497) );
  INVX1_HVT U382 ( .A(key[5]), .Y(n439) );
  INVX1_HVT U383 ( .A(key_round[1]), .Y(n396) );
  INVX1_HVT U384 ( .A(key[1]), .Y(n395) );
  INVX1_HVT U385 ( .A(adk_out0[117]), .Y(n445) );
  INVX1_HVT U386 ( .A(adk_out0[112]), .Y(n554) );
  INVX1_HVT U387 ( .A(adk_out0[111]), .Y(n470) );
  NAND2X0_HVT U388 ( .A1(n718), .A2(n805), .Y(n320) );
  INVX1_HVT U389 ( .A(adk_out0[102]), .Y(n401) );
  INVX1_HVT U390 ( .A(adk_out0[70]), .Y(n539) );
  INVX1_HVT U391 ( .A(adk_out0[67]), .Y(n398) );
  INVX1_HVT U392 ( .A(adk_out0[59]), .Y(n435) );
  INVX1_HVT U393 ( .A(adk_out0[21]), .Y(n514) );
  INVX1_HVT U394 ( .A(adk_out0[16]), .Y(n467) );
  INVX1_HVT U395 ( .A(adk_out0[5]), .Y(n503) );
  INVX1_HVT U396 ( .A(n815), .Y(n573) );
  INVX0_HVT U397 ( .A(n556), .Y(n310) );
  INVX0_HVT U398 ( .A(n556), .Y(n297) );
  INVX1_HVT U399 ( .A(n820), .Y(n783) );
  INVX1_HVT U400 ( .A(n367), .Y(n303) );
  INVX1_HVT U401 ( .A(n512), .Y(n386) );
  INVX1_HVT U402 ( .A(n512), .Y(n309) );
  INVX1_HVT U403 ( .A(n800), .Y(n447) );
  INVX1_HVT U404 ( .A(n403), .Y(n301) );
  INVX1_HVT U405 ( .A(n403), .Y(n306) );
  INVX1_HVT U406 ( .A(n822), .Y(n588) );
  INVX1_HVT U407 ( .A(n326), .Y(n551) );
  OAI222X1_HVT U408 ( .A1(n369), .A2(n368), .A3(n370), .A4(n436), .A5(n371), 
        .A6(n379), .Y(n285) );
  INVX1_HVT U409 ( .A(n534), .Y(n300) );
  NBUFFX2_HVT U410 ( .A(n793), .Y(n798) );
  INVX1_HVT U411 ( .A(n326), .Y(n298) );
  INVX0_HVT U412 ( .A(n531), .Y(n489) );
  INVX1_HVT U413 ( .A(n448), .Y(n307) );
  INVX1_HVT U414 ( .A(n822), .Y(n586) );
  INVX0_HVT U415 ( .A(n562), .Y(n332) );
  INVX1_HVT U416 ( .A(n576), .Y(n530) );
  INVX1_HVT U417 ( .A(n822), .Y(n589) );
  INVX1_HVT U418 ( .A(n534), .Y(n313) );
  INVX1_HVT U419 ( .A(n482), .Y(n473) );
  INVX1_HVT U420 ( .A(n591), .Y(n578) );
  INVX1_HVT U421 ( .A(n805), .Y(n529) );
  INVX1_HVT U422 ( .A(n389), .Y(n304) );
  OAI222X1_HVT U423 ( .A1(n372), .A2(n389), .A3(n373), .A4(n436), .A5(n374), 
        .A6(n531), .Y(n286) );
  INVX1_HVT U424 ( .A(n788), .Y(n384) );
  INVX1_HVT U425 ( .A(n433), .Y(n368) );
  OAI222X1_HVT U426 ( .A1(n346), .A2(n389), .A3(n347), .A4(n402), .A5(n348), 
        .A6(n561), .Y(n287) );
  NAND3X0_HVT U427 ( .A1(n318), .A2(n319), .A3(n320), .Y(n288) );
  AND2X1_HVT U428 ( .A1(n574), .A2(n763), .Y(n289) );
  OAI222X1_HVT U429 ( .A1(n509), .A2(n822), .A3(n510), .A4(n512), .A5(n511), 
        .A6(n379), .Y(n290) );
  OR2X1_HVT U430 ( .A1(n407), .A2(n529), .Y(n291) );
  INVX1_HVT U431 ( .A(n529), .Y(n311) );
  INVX1_HVT U432 ( .A(n362), .Y(n312) );
  INVX1_HVT U433 ( .A(n384), .Y(n302) );
  INVX1_HVT U434 ( .A(n361), .Y(n569) );
  NBUFFX2_HVT U435 ( .A(n595), .Y(n433) );
  INVX1_HVT U436 ( .A(n763), .Y(n358) );
  INVX1_HVT U437 ( .A(n563), .Y(n299) );
  INVX1_HVT U438 ( .A(key_round[9]), .Y(n498) );
  INVX1_HVT U439 ( .A(n552), .Y(n305) );
  INVX1_HVT U440 ( .A(n532), .Y(n308) );
  AO222X1_HVT U441 ( .A1(cipher_text[94]), .A2(n586), .A3(adk_out0[94]), .A4(
        n296), .A5(adk_in[94]), .A6(n297), .Y(n181) );
  AO222X1_HVT U442 ( .A1(cipher_text[87]), .A2(n298), .A3(adk_out0[87]), .A4(
        n302), .A5(n299), .A6(n300), .Y(n188) );
  INVX0_HVT U443 ( .A(keyout[18]), .Y(n334) );
  AO222X1_HVT U444 ( .A1(cipher_text[103]), .A2(n587), .A3(adk_out0[103]), 
        .A4(n768), .A5(adk_in[103]), .A6(n300), .Y(n172) );
  AO222X1_HVT U445 ( .A1(cipher_text[62]), .A2(n301), .A3(adk_out0[62]), .A4(
        n302), .A5(adk_in[62]), .A6(n303), .Y(n213) );
  AO222X1_HVT U446 ( .A1(cipher_text[83]), .A2(n578), .A3(adk_out0[83]), .A4(
        n780), .A5(n681), .A6(n313), .Y(n192) );
  INVX1_HVT U447 ( .A(adk_in[67]), .Y(n399) );
  AO222X1_HVT U448 ( .A1(cipher_text[7]), .A2(n580), .A3(adk_out0[7]), .A4(
        n302), .A5(adk_in[7]), .A6(n311), .Y(n268) );
  AO222X1_HVT U449 ( .A1(cipher_text[74]), .A2(n298), .A3(adk_out0[74]), .A4(
        n783), .A5(n620), .A6(n355), .Y(n201) );
  AO222X1_HVT U450 ( .A1(cipher_text[76]), .A2(n304), .A3(adk_out0[76]), .A4(
        n302), .A5(adk_in[76]), .A6(n311), .Y(n199) );
  AO222X1_HVT U451 ( .A1(cipher_text[90]), .A2(n587), .A3(adk_out0[90]), .A4(
        n302), .A5(n305), .A6(n284), .Y(n185) );
  AO222X1_HVT U452 ( .A1(cipher_text[64]), .A2(n306), .A3(adk_out0[64]), .A4(
        n776), .A5(adk_in[64]), .A6(n311), .Y(n211) );
  AO222X1_HVT U453 ( .A1(cipher_text[63]), .A2(n321), .A3(adk_out0[63]), .A4(
        n307), .A5(n756), .A6(n489), .Y(n212) );
  AO222X1_HVT U454 ( .A1(cipher_text[14]), .A2(n581), .A3(adk_out0[14]), .A4(
        n770), .A5(adk_in[14]), .A6(n300), .Y(n261) );
  AO222X1_HVT U455 ( .A1(cipher_text[33]), .A2(n585), .A3(adk_out0[33]), .A4(
        n386), .A5(n732), .A6(n312), .Y(n242) );
  INVX1_HVT U456 ( .A(n578), .Y(n822) );
  AO222X1_HVT U457 ( .A1(cipher_text[85]), .A2(n579), .A3(adk_out0[85]), .A4(
        n792), .A5(n381), .A6(n308), .Y(n190) );
  AO222X1_HVT U458 ( .A1(cipher_text[23]), .A2(n321), .A3(adk_out0[23]), .A4(
        n309), .A5(n750), .A6(n310), .Y(n252) );
  AO222X1_HVT U459 ( .A1(cipher_text[100]), .A2(n551), .A3(adk_out0[100]), 
        .A4(n791), .A5(n722), .A6(n311), .Y(n366) );
  AO222X1_HVT U460 ( .A1(cipher_text[124]), .A2(n576), .A3(adk_out0[124]), 
        .A4(n791), .A5(adk_in[124]), .A6(n312), .Y(n151) );
  AO222X1_HVT U461 ( .A1(cipher_text[123]), .A2(n433), .A3(adk_out0[123]), 
        .A4(n768), .A5(n313), .A6(n668), .Y(n152) );
  AO222X1_HVT U462 ( .A1(cipher_text[89]), .A2(n587), .A3(adk_out0[89]), .A4(
        n375), .A5(n720), .A6(n355), .Y(n186) );
  INVX0_HVT U463 ( .A(n637), .Y(n638) );
  INVX1_HVT U464 ( .A(n314), .Y(n315) );
  INVX1_HVT U465 ( .A(n316), .Y(n317) );
  NAND2X0_HVT U466 ( .A1(n578), .A2(cipher_text[108]), .Y(n318) );
  NAND2X0_HVT U467 ( .A1(adk_out0[108]), .A2(n375), .Y(n319) );
  INVX0_HVT U468 ( .A(round_number[3]), .Y(n354) );
  INVX1_HVT U469 ( .A(adk_in[59]), .Y(n437) );
  INVX1_HVT U470 ( .A(round_number[2]), .Y(n505) );
  NAND2X0_HVT U471 ( .A1(n281), .A2(n289), .Y(n417) );
  INVX1_HVT U472 ( .A(n326), .Y(n597) );
  INVX1_HVT U473 ( .A(n322), .Y(n323) );
  OAI222X2_HVT U474 ( .A1(n502), .A2(n474), .A3(n503), .A4(n447), .A5(n504), 
        .A6(n341), .Y(n270) );
  INVX0_HVT U475 ( .A(n727), .Y(n728) );
  INVX1_HVT U476 ( .A(n324), .Y(n325) );
  INVX0_HVT U477 ( .A(n733), .Y(n734) );
  OAI222X1_HVT U478 ( .A1(n449), .A2(n474), .A3(n450), .A4(n451), .A5(n452), 
        .A6(n341), .Y(n40) );
  INVX1_HVT U479 ( .A(n321), .Y(n474) );
  INVX1_HVT U480 ( .A(n490), .Y(n326) );
  INVX0_HVT U481 ( .A(n677), .Y(n678) );
  INVX0_HVT U482 ( .A(n648), .Y(n649) );
  INVX0_HVT U483 ( .A(n665), .Y(n666) );
  INVX0_HVT U484 ( .A(n607), .Y(n608) );
  INVX0_HVT U485 ( .A(n639), .Y(n640) );
  INVX0_HVT U486 ( .A(n735), .Y(n736) );
  INVX0_HVT U487 ( .A(n729), .Y(n730) );
  INVX0_HVT U488 ( .A(n759), .Y(n760) );
  INVX0_HVT U489 ( .A(n755), .Y(n756) );
  INVX0_HVT U490 ( .A(n627), .Y(n628) );
  INVX0_HVT U491 ( .A(n753), .Y(n754) );
  INVX0_HVT U492 ( .A(n643), .Y(n644) );
  INVX1_HVT U493 ( .A(n5), .Y(n361) );
  INVX1_HVT U494 ( .A(n327), .Y(n328) );
  INVX0_HVT U495 ( .A(n695), .Y(n696) );
  INVX0_HVT U496 ( .A(n707), .Y(n708) );
  INVX0_HVT U497 ( .A(keyout[57]), .Y(n548) );
  INVX0_HVT U498 ( .A(n741), .Y(n742) );
  INVX1_HVT U499 ( .A(n816), .Y(n810) );
  INVX0_HVT U500 ( .A(n709), .Y(n710) );
  INVX0_HVT U501 ( .A(n599), .Y(n600) );
  OR2X1_HVT U502 ( .A1(n329), .A2(n331), .Y(n508) );
  OR2X1_HVT U503 ( .A1(n330), .A2(n431), .Y(n523) );
  INVX0_HVT U504 ( .A(n699), .Y(n700) );
  INVX0_HVT U505 ( .A(n621), .Y(n622) );
  NBUFFX2_HVT U506 ( .A(n816), .Y(n331) );
  INVX0_HVT U507 ( .A(n667), .Y(n668) );
  INVX0_HVT U508 ( .A(n814), .Y(n562) );
  INVX1_HVT U509 ( .A(n378), .Y(n793) );
  INVX0_HVT U510 ( .A(n682), .Y(n683) );
  INVX0_HVT U511 ( .A(n749), .Y(n750) );
  INVX0_HVT U512 ( .A(n686), .Y(n687) );
  INVX0_HVT U513 ( .A(n743), .Y(n744) );
  INVX1_HVT U514 ( .A(n818), .Y(n803) );
  INVX0_HVT U515 ( .A(n663), .Y(n664) );
  OR2X1_HVT U516 ( .A1(n333), .A2(n561), .Y(n485) );
  OAI222X1_HVT U517 ( .A1(n337), .A2(n368), .A3(n338), .A4(n533), .A5(n339), 
        .A6(n561), .Y(n21) );
  NBUFFX2_HVT U518 ( .A(n812), .Y(n340) );
  INVX0_HVT U519 ( .A(n717), .Y(n718) );
  INVX0_HVT U520 ( .A(n657), .Y(n658) );
  INVX0_HVT U521 ( .A(n723), .Y(n724) );
  INVX0_HVT U522 ( .A(n751), .Y(n752) );
  INVX1_HVT U523 ( .A(n745), .Y(n746) );
  INVX0_HVT U524 ( .A(n659), .Y(n660) );
  INVX0_HVT U525 ( .A(n669), .Y(n670) );
  INVX0_HVT U526 ( .A(n381), .Y(n341) );
  INVX0_HVT U527 ( .A(n675), .Y(n676) );
  IBUFFX2_HVT U528 ( .A(n505), .Y(n342) );
  INVX0_HVT U529 ( .A(n362), .Y(n355) );
  NBUFFX2_HVT U530 ( .A(n766), .Y(n789) );
  OAI222X1_HVT U531 ( .A1(n349), .A2(n389), .A3(n350), .A4(n543), .A5(n351), 
        .A6(n561), .Y(n28) );
  INVX1_HVT U532 ( .A(n352), .Y(n353) );
  INVX0_HVT U533 ( .A(keyout[25]), .Y(n475) );
  INVX0_HVT U534 ( .A(n382), .Y(n775) );
  INVX0_HVT U535 ( .A(n819), .Y(n788) );
  INVX0_HVT U536 ( .A(n378), .Y(n794) );
  INVX0_HVT U537 ( .A(n680), .Y(n681) );
  INVX0_HVT U538 ( .A(n737), .Y(n738) );
  INVX1_HVT U539 ( .A(n703), .Y(n704) );
  AO222X1_HVT U540 ( .A1(cipher_text[38]), .A2(n587), .A3(adk_out0[38]), .A4(
        n282), .A5(adk_in[38]), .A6(n355), .Y(n237) );
  INVX0_HVT U541 ( .A(n692), .Y(n693) );
  INVX1_HVT U542 ( .A(n688), .Y(n689) );
  INVX0_HVT U543 ( .A(n671), .Y(n672) );
  INVX0_HVT U544 ( .A(n633), .Y(n634) );
  INVX0_HVT U545 ( .A(n601), .Y(n602) );
  INVX1_HVT U546 ( .A(n356), .Y(n357) );
  INVX0_HVT U547 ( .A(n701), .Y(n702) );
  INVX0_HVT U548 ( .A(n684), .Y(n685) );
  INVX0_HVT U549 ( .A(n653), .Y(n654) );
  INVX0_HVT U550 ( .A(keyout[1]), .Y(n394) );
  INVX0_HVT U551 ( .A(n739), .Y(n740) );
  INVX0_HVT U552 ( .A(n713), .Y(n714) );
  INVX0_HVT U553 ( .A(n817), .Y(n805) );
  INVX0_HVT U554 ( .A(n721), .Y(n722) );
  NBUFFX2_HVT U555 ( .A(n792), .Y(n796) );
  INVX0_HVT U556 ( .A(n614), .Y(n615) );
  INVX0_HVT U557 ( .A(n635), .Y(n636) );
  INVX0_HVT U558 ( .A(n378), .Y(n776) );
  INVX0_HVT U559 ( .A(n673), .Y(n674) );
  INVX0_HVT U560 ( .A(n781), .Y(n402) );
  INVX0_HVT U561 ( .A(keyout[40]), .Y(n441) );
  INVX0_HVT U562 ( .A(n612), .Y(n613) );
  INVX0_HVT U563 ( .A(keyout[46]), .Y(n412) );
  INVX0_HVT U564 ( .A(n655), .Y(n656) );
  INVX0_HVT U565 ( .A(n747), .Y(n748) );
  INVX0_HVT U566 ( .A(n562), .Y(n419) );
  INVX0_HVT U567 ( .A(n630), .Y(n631) );
  INVX0_HVT U568 ( .A(n715), .Y(n716) );
  INVX0_HVT U569 ( .A(n616), .Y(n617) );
  INVX0_HVT U570 ( .A(n725), .Y(n726) );
  INVX0_HVT U571 ( .A(n761), .Y(n824) );
  INVX0_HVT U572 ( .A(n711), .Y(n712) );
  INVX1_HVT U573 ( .A(n651), .Y(n652) );
  INVX0_HVT U574 ( .A(cipher_text[102]), .Y(n400) );
  AO222X1_HVT U575 ( .A1(keyout[116]), .A2(n586), .A3(key[116]), .A4(n791), 
        .A5(key_round[116]), .A6(n377), .Y(n31) );
  INVX0_HVT U576 ( .A(n381), .Y(n379) );
  INVX0_HVT U577 ( .A(n815), .Y(n814) );
  INVX0_HVT U578 ( .A(n645), .Y(n646) );
  AO222X1_HVT U579 ( .A1(cipher_text[92]), .A2(n589), .A3(adk_out0[92]), .A4(
        n376), .A5(n646), .A6(n311), .Y(n183) );
  INVX0_HVT U580 ( .A(n719), .Y(n720) );
  INVX0_HVT U581 ( .A(n605), .Y(n606) );
  INVX0_HVT U582 ( .A(n618), .Y(n619) );
  OAI222X1_HVT U583 ( .A1(n359), .A2(n368), .A3(n360), .A4(n464), .A5(n292), 
        .A6(n362), .Y(n68) );
  NBUFFX2_HVT U584 ( .A(n529), .Y(n362) );
  INVX1_HVT U585 ( .A(n581), .Y(n528) );
  INVX0_HVT U586 ( .A(keyout[30]), .Y(n363) );
  INVX0_HVT U587 ( .A(n810), .Y(n561) );
  INVX0_HVT U588 ( .A(n690), .Y(n691) );
  OAI222X1_HVT U589 ( .A1(n363), .A2(n368), .A3(n364), .A4(n543), .A5(n295), 
        .A6(n379), .Y(n117) );
  INVX0_HVT U590 ( .A(n609), .Y(n610) );
  INVX0_HVT U591 ( .A(keyout[16]), .Y(n369) );
  AO222X1_HVT U592 ( .A1(keyout[97]), .A2(n576), .A3(key[97]), .A4(n778), .A5(
        key_round[97]), .A6(n332), .Y(n365) );
  INVX0_HVT U593 ( .A(n705), .Y(n706) );
  INVX0_HVT U594 ( .A(n661), .Y(n662) );
  INVX16_HVT U595 ( .A(n389), .Y(n594) );
  NBUFFX2_HVT U596 ( .A(n562), .Y(n367) );
  NBUFFX2_HVT U597 ( .A(n767), .Y(n771) );
  INVX0_HVT U598 ( .A(n574), .Y(n575) );
  INVX0_HVT U599 ( .A(n384), .Y(n765) );
  NBUFFX2_HVT U600 ( .A(n783), .Y(n375) );
  NBUFFX2_HVT U601 ( .A(n783), .Y(n376) );
  INVX0_HVT U602 ( .A(n431), .Y(n377) );
  INVX0_HVT U603 ( .A(cipher_text[16]), .Y(n466) );
  INVX0_HVT U604 ( .A(n775), .Y(n378) );
  INVX0_HVT U605 ( .A(n531), .Y(n381) );
  AO222X1_HVT U606 ( .A1(cipher_text[12]), .A2(n585), .A3(adk_out0[12]), .A4(
        n798), .A5(n712), .A6(n381), .Y(n380) );
  INVX0_HVT U607 ( .A(n820), .Y(n767) );
  INVX0_HVT U608 ( .A(n774), .Y(n820) );
  INVX0_HVT U609 ( .A(n775), .Y(n819) );
  INVX0_HVT U610 ( .A(n774), .Y(n821) );
  INVX1_HVT U611 ( .A(keyout[35]), .Y(n423) );
  INVX0_HVT U612 ( .A(n810), .Y(n431) );
  INVX0_HVT U613 ( .A(cipher_text[117]), .Y(n444) );
  INVX0_HVT U614 ( .A(keyout[34]), .Y(n420) );
  INVX0_HVT U615 ( .A(cipher_text[112]), .Y(n553) );
  NAND2X0_HVT U616 ( .A1(n816), .A2(n491), .Y(n382) );
  INVX0_HVT U617 ( .A(n419), .Y(n383) );
  INVX0_HVT U618 ( .A(cipher_text[111]), .Y(n469) );
  NBUFFX2_HVT U619 ( .A(round_number[2]), .Y(n408) );
  INVX0_HVT U620 ( .A(n805), .Y(n534) );
  INVX16_HVT U621 ( .A(n388), .Y(n595) );
  INVX0_HVT U622 ( .A(n814), .Y(n531) );
  INVX0_HVT U623 ( .A(cipher_text[67]), .Y(n397) );
  AO222X1_HVT U624 ( .A1(keyout[11]), .A2(n578), .A3(key[11]), .A4(n386), .A5(
        n387), .A6(n419), .Y(n385) );
  INVX0_HVT U625 ( .A(n820), .Y(n782) );
  INVX0_HVT U626 ( .A(n799), .Y(n543) );
  INVX0_HVT U627 ( .A(n797), .Y(n555) );
  INVX0_HVT U628 ( .A(keyout[50]), .Y(n499) );
  NBUFFX2_HVT U629 ( .A(n793), .Y(n797) );
  INVX0_HVT U630 ( .A(keyout[21]), .Y(n426) );
  INVX1_HVT U631 ( .A(keyout[84]), .Y(n535) );
  NAND2X4_HVT U632 ( .A1(n480), .A2(n762), .Y(n471) );
  IBUFFX8_HVT U633 ( .A(n593), .Y(n388) );
  IBUFFX8_HVT U634 ( .A(n593), .Y(n389) );
  INVX0_HVT U635 ( .A(n496), .Y(n390) );
  INVX0_HVT U636 ( .A(n304), .Y(n496) );
  INVX2_HVT U637 ( .A(n493), .Y(n482) );
  OAI222X1_HVT U638 ( .A1(n391), .A2(n403), .A3(n392), .A4(n402), .A5(n393), 
        .A6(n367), .Y(n100) );
  OAI222X1_HVT U639 ( .A1(n394), .A2(n403), .A3(n395), .A4(n820), .A5(n396), 
        .A6(n531), .Y(n146) );
  AO222X1_HVT U640 ( .A1(keyout[72]), .A2(n321), .A3(key[72]), .A4(n790), .A5(
        key_round[72]), .A6(n312), .Y(n75) );
  OAI222X1_HVT U641 ( .A1(n473), .A2(n400), .A3(n401), .A4(n402), .A5(n472), 
        .A6(n534), .Y(n173) );
  INVX0_HVT U642 ( .A(n579), .Y(n403) );
  OAI222X1_HVT U643 ( .A1(n404), .A2(n473), .A3(n405), .A4(n533), .A5(n406), 
        .A6(n561), .Y(n121) );
  INVX0_HVT U644 ( .A(cipher_text[59]), .Y(n434) );
  INVX0_HVT U645 ( .A(n388), .Y(n587) );
  OAI222X1_HVT U646 ( .A1(n409), .A2(n528), .A3(n410), .A4(n451), .A5(n411), 
        .A6(n383), .Y(n103) );
  OAI222X1_HVT U647 ( .A1(n412), .A2(n474), .A3(n413), .A4(n533), .A5(n414), 
        .A6(n431), .Y(n101) );
  INVX1_HVT U648 ( .A(n415), .Y(n416) );
  AND2X1_HVT U649 ( .A1(n417), .A2(n818), .Y(n8) );
  AO222X1_HVT U650 ( .A1(cipher_text[44]), .A2(n304), .A3(adk_out0[44]), .A4(
        n302), .A5(n738), .A6(n419), .Y(n418) );
  OAI222X1_HVT U651 ( .A1(n420), .A2(n528), .A3(n421), .A4(n543), .A5(n422), 
        .A6(n534), .Y(n113) );
  OAI222X1_HVT U652 ( .A1(n426), .A2(n530), .A3(n427), .A4(n533), .A5(n293), 
        .A6(n341), .Y(n126) );
  OAI222X1_HVT U653 ( .A1(n428), .A2(n474), .A3(n429), .A4(n430), .A5(n432), 
        .A6(n431), .Y(n44) );
  NBUFFX2_HVT U654 ( .A(n766), .Y(n770) );
  OAI222X1_HVT U655 ( .A1(n438), .A2(n368), .A3(n439), .A4(n447), .A5(n294), 
        .A6(n562), .Y(n142) );
  OAI222X1_HVT U656 ( .A1(n441), .A2(n530), .A3(n442), .A4(n533), .A5(n443), 
        .A6(n367), .Y(n440) );
  OAI222X1_HVT U657 ( .A1(n496), .A2(n444), .A3(n445), .A4(n555), .A5(n446), 
        .A6(n331), .Y(n158) );
  OAI222X1_HVT U658 ( .A1(n453), .A2(n403), .A3(n454), .A4(n533), .A5(n455), 
        .A6(n383), .Y(n38) );
  NAND2X0_HVT U659 ( .A1(n587), .A2(cipher_text[86]), .Y(n456) );
  NAND2X0_HVT U660 ( .A1(adk_out0[86]), .A2(n777), .Y(n457) );
  NAND2X0_HVT U661 ( .A1(adk_in[86]), .A2(n303), .Y(n458) );
  NAND3X0_HVT U662 ( .A1(n456), .A2(n457), .A3(n458), .Y(n189) );
  NBUFFX2_HVT U663 ( .A(n794), .Y(n777) );
  OAI222X1_HVT U664 ( .A1(n459), .A2(n474), .A3(n460), .A4(n430), .A5(n461), 
        .A6(n818), .Y(n91) );
  OAI222X1_HVT U665 ( .A1(n462), .A2(n473), .A3(n463), .A4(n464), .A5(n465), 
        .A6(n561), .Y(n83) );
  OAI222X1_HVT U666 ( .A1(n475), .A2(n496), .A3(n476), .A4(n451), .A5(n624), 
        .A6(n362), .Y(n122) );
  OAI222X1_HVT U667 ( .A1(n477), .A2(n496), .A3(n478), .A4(n512), .A5(n479), 
        .A6(n561), .Y(n35) );
  OR2X1_HVT U668 ( .A1(n764), .A2(n354), .Y(n480) );
  IBUFFX8_HVT U669 ( .A(n471), .Y(n481) );
  NAND2X0_HVT U670 ( .A1(keyout[118]), .A2(n298), .Y(n483) );
  NAND2X0_HVT U671 ( .A1(key[118]), .A2(n779), .Y(n484) );
  NAND3X0_HVT U672 ( .A1(n483), .A2(n484), .A3(n485), .Y(n29) );
  NAND2X0_HVT U673 ( .A1(key[14]), .A2(n786), .Y(n487) );
  NAND3X0_HVT U674 ( .A1(n486), .A2(n487), .A3(n291), .Y(n133) );
  AO222X1_HVT U675 ( .A1(cipher_text[121]), .A2(n306), .A3(adk_out0[121]), 
        .A4(n782), .A5(adk_in[121]), .A6(n489), .Y(n154) );
  INVX1_HVT U676 ( .A(n593), .Y(n823) );
  INVX16_HVT U677 ( .A(n493), .Y(n490) );
  IBUFFX8_HVT U678 ( .A(n593), .Y(n493) );
  OAI222X1_HVT U679 ( .A1(n823), .A2(n513), .A3(n514), .A4(n464), .A5(n515), 
        .A6(n379), .Y(n492) );
  OAI222X1_HVT U680 ( .A1(n495), .A2(n368), .A3(n497), .A4(n512), .A5(n498), 
        .A6(n341), .Y(n138) );
  INVX0_HVT U681 ( .A(cipher_text[5]), .Y(n502) );
  AO222X1_HVT U682 ( .A1(keyout[123]), .A2(n596), .A3(key[123]), .A4(n792), 
        .A5(key_round[123]), .A6(n812), .Y(n24) );
  INVX0_HVT U683 ( .A(cipher_text[70]), .Y(n538) );
  AO222X1_HVT U684 ( .A1(keyout[122]), .A2(n597), .A3(key[122]), .A4(n307), 
        .A5(key_round[122]), .A6(n381), .Y(n25) );
  INVX0_HVT U685 ( .A(cipher_text[21]), .Y(n513) );
  NAND2X0_HVT U686 ( .A1(key[78]), .A2(n788), .Y(n507) );
  NAND3X0_HVT U687 ( .A1(n506), .A2(n507), .A3(n508), .Y(n69) );
  OAI22X1_HVT U688 ( .A1(reset), .A2(n815), .A3(n805), .A4(n575), .Y(n517) );
  INVX2_HVT U689 ( .A(n802), .Y(n815) );
  AO21X1_HVT U690 ( .A1(n569), .A2(n818), .A3(n15), .Y(n12) );
  NAND2X0_HVT U691 ( .A1(key[54]), .A2(n788), .Y(n519) );
  NAND2X0_HVT U692 ( .A1(key_round[54]), .A2(n805), .Y(n520) );
  NAND3X0_HVT U693 ( .A1(n520), .A2(n519), .A3(n518), .Y(n93) );
  NAND2X0_HVT U694 ( .A1(keyout[42]), .A2(n298), .Y(n521) );
  NAND2X0_HVT U695 ( .A1(key[42]), .A2(n787), .Y(n522) );
  NAND3X0_HVT U696 ( .A1(n521), .A2(n522), .A3(n523), .Y(n105) );
  OAI222X1_HVT U697 ( .A1(n474), .A2(n538), .A3(n539), .A4(n464), .A5(n540), 
        .A6(n362), .Y(n524) );
  NAND2X0_HVT U698 ( .A1(key[77]), .A2(n773), .Y(n526) );
  NAND2X0_HVT U699 ( .A1(key_round[77]), .A2(n516), .Y(n527) );
  NAND3X0_HVT U700 ( .A1(n527), .A2(n526), .A3(n525), .Y(n70) );
  INVX0_HVT U701 ( .A(n823), .Y(n581) );
  INVX0_HVT U702 ( .A(n822), .Y(n576) );
  OAI222X1_HVT U703 ( .A1(n535), .A2(n403), .A3(n536), .A4(n384), .A5(n537), 
        .A6(n341), .Y(n63) );
  OAI222X1_HVT U704 ( .A1(n541), .A2(n368), .A3(n542), .A4(n543), .A5(n544), 
        .A6(n341), .Y(n46) );
  OAI222X1_HVT U705 ( .A1(n545), .A2(n528), .A3(n546), .A4(n447), .A5(n547), 
        .A6(n562), .Y(n49) );
  INVX0_HVT U706 ( .A(n573), .Y(n556) );
  OAI222X1_HVT U707 ( .A1(n548), .A2(n368), .A3(n549), .A4(n436), .A5(n550), 
        .A6(n529), .Y(n90) );
  OAI222X1_HVT U708 ( .A1(n474), .A2(n553), .A3(n554), .A4(n555), .A5(n556), 
        .A6(n557), .Y(n163) );
  OAI222X1_HVT U709 ( .A1(n558), .A2(n530), .A3(n559), .A4(n436), .A5(n560), 
        .A6(n529), .Y(n59) );
  NAND2X0_HVT U710 ( .A1(keyout[111]), .A2(n579), .Y(n564) );
  NAND2X0_HVT U711 ( .A1(key[111]), .A2(n296), .Y(n565) );
  NAND2X0_HVT U712 ( .A1(key_round[111]), .A2(n810), .Y(n566) );
  NAND3X0_HVT U713 ( .A1(n564), .A2(n565), .A3(n566), .Y(n36) );
  INVX0_HVT U714 ( .A(round_number[1]), .Y(n567) );
  NAND2X0_HVT U715 ( .A1(keyout[114]), .A2(n598), .Y(n570) );
  NAND2X0_HVT U716 ( .A1(key[114]), .A2(n765), .Y(n571) );
  NAND2X0_HVT U717 ( .A1(key_round[114]), .A2(n810), .Y(n572) );
  NAND3X0_HVT U718 ( .A1(n570), .A2(n571), .A3(n572), .Y(n33) );
  NBUFFX2_HVT U719 ( .A(n576), .Y(n577) );
  NBUFFX2_HVT U720 ( .A(n433), .Y(n580) );
  NBUFFX2_HVT U721 ( .A(n551), .Y(n582) );
  NBUFFX2_HVT U722 ( .A(n551), .Y(n583) );
  IBUFFX8_HVT U723 ( .A(n8), .Y(n590) );
  IBUFFX32_HVT U724 ( .A(n590), .Y(n593) );
  INVX1_HVT U725 ( .A(n603), .Y(n604) );
  INVX1_HVT U726 ( .A(n731), .Y(n732) );
  INVX1_HVT U727 ( .A(n625), .Y(n626) );
  INVX1_HVT U728 ( .A(n697), .Y(n698) );
  IBUFFX8_HVT U729 ( .A(reset), .Y(n762) );
  NBUFFX2_HVT U730 ( .A(n768), .Y(n772) );
  NBUFFX2_HVT U731 ( .A(n784), .Y(n786) );
  NBUFFX2_HVT U732 ( .A(n768), .Y(n773) );
  NBUFFX2_HVT U733 ( .A(n788), .Y(n791) );
  NBUFFX2_HVT U734 ( .A(n788), .Y(n790) );
  NBUFFX2_HVT U735 ( .A(n784), .Y(n785) );
  NBUFFX2_HVT U736 ( .A(n794), .Y(n800) );
  NBUFFX2_HVT U737 ( .A(n794), .Y(n799) );
  INVX1_HVT U738 ( .A(n821), .Y(n768) );
  INVX1_HVT U739 ( .A(n821), .Y(n784) );
  INVX1_HVT U740 ( .A(n802), .Y(n816) );
  INVX4_HVT U741 ( .A(n802), .Y(n817) );
  AND2X1_HVT U742 ( .A1(n5), .A2(n4), .Y(n764) );
  INVX1_HVT U743 ( .A(n819), .Y(n766) );
  NBUFFX2_HVT U744 ( .A(n774), .Y(n779) );
  NBUFFX2_HVT U745 ( .A(n776), .Y(n780) );
  NBUFFX2_HVT U746 ( .A(n776), .Y(n781) );
  INVX1_HVT U747 ( .A(n819), .Y(n787) );
  INVX1_HVT U748 ( .A(n821), .Y(n792) );
  IBUFFX32_HVT U749 ( .A(n481), .Y(n802) );
  NAND2X0_HVT U750 ( .A1(n575), .A2(n814), .Y(n825) );
  OAI22X1_HVT U751 ( .A1(reset), .A2(n825), .A3(n573), .A4(n575), .Y(n279) );
  OAI22X1_HVT U752 ( .A1(reset), .A2(n815), .A3(n810), .A4(n826), .Y(n15) );
  NOR2X1_HVT U753 ( .A1(reset), .A2(n827), .Y(n19) );
endmodule

