
module sbox_17 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n7, n19, n23, n39, n48, n121, n147, n210, n211, n212, n213, n216,
         n217, n218, n219, n227, n231, n232, n236, n238, n239, n240, n243,
         n249, n257, n261, n264, n266, n269, n273, n279, n280, n282, n283,
         n293, n297, n299, n301, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712;

  NAND2X0_HVT U4 ( .A1(n428), .A2(n39), .Y(n709) );
  NAND2X0_HVT U5 ( .A1(n361), .A2(n421), .Y(n707) );
  NAND2X0_HVT U13 ( .A1(n700), .A2(n320), .Y(n701) );
  NAND2X0_HVT U15 ( .A1(n710), .A2(n368), .Y(n698) );
  NAND2X0_HVT U21 ( .A1(n427), .A2(n312), .Y(n693) );
  NAND2X0_HVT U24 ( .A1(n305), .A2(n337), .Y(n691) );
  NAND2X0_HVT U33 ( .A1(n313), .A2(n329), .Y(n682) );
  NAND2X0_HVT U42 ( .A1(n374), .A2(n352), .Y(n674) );
  MUX41X1_HVT U51 ( .A1(n454), .A3(n478), .A2(n338), .A4(n456), .S0(n340), 
        .S1(n412), .Y(n666) );
  NAND2X0_HVT U53 ( .A1(n663), .A2(n673), .Y(n664) );
  NAND2X0_HVT U56 ( .A1(n428), .A2(n659), .Y(n660) );
  MUX41X1_HVT U57 ( .A1(n466), .A3(n695), .A2(n660), .A4(n703), .S0(n446), 
        .S1(n412), .Y(n658) );
  NAND2X0_HVT U58 ( .A1(n320), .A2(n710), .Y(n657) );
  NAND2X0_HVT U62 ( .A1(n312), .A2(n430), .Y(n653) );
  AO21X1_HVT U66 ( .A1(n493), .A2(n440), .A3(n335), .Y(n649) );
  MUX41X1_HVT U68 ( .A1(n461), .A3(n649), .A2(n648), .A4(n650), .S0(n406), 
        .S1(n445), .Y(n647) );
  MUX41X1_HVT U69 ( .A1(n647), .A3(n655), .A2(n651), .A4(n661), .S0(in[6]), 
        .S1(n416), .Y(out[0]) );
  NAND2X0_HVT U73 ( .A1(n424), .A2(n642), .Y(n643) );
  MUX41X1_HVT U74 ( .A1(n644), .A3(n689), .A2(n643), .A4(n691), .S0(n408), 
        .S1(n446), .Y(n641) );
  MUX41X1_HVT U77 ( .A1(n705), .A3(n475), .A2(n639), .A4(n465), .S0(n413), 
        .S1(n405), .Y(n638) );
  MUX41X1_HVT U82 ( .A1(n671), .A3(n456), .A2(n498), .A4(n699), .S0(n406), 
        .S1(n340), .Y(n632) );
  AND2X1_HVT U83 ( .A1(n361), .A2(n333), .Y(n631) );
  NAND2X0_HVT U85 ( .A1(n329), .A2(n318), .Y(n629) );
  MUX41X1_HVT U86 ( .A1(n489), .A3(n629), .A2(n400), .A4(n395), .S0(n406), 
        .S1(n445), .Y(n628) );
  MUX41X1_HVT U96 ( .A1(n498), .A3(n401), .A2(n491), .A4(n619), .S0(n406), 
        .S1(n444), .Y(n618) );
  MUX41X1_HVT U97 ( .A1(n492), .A3(n401), .A2(n374), .A4(n698), .S0(n406), 
        .S1(n380), .Y(n617) );
  NAND2X0_HVT U101 ( .A1(n612), .A2(n611), .Y(n613) );
  MUX41X1_HVT U103 ( .A1(n39), .A3(n480), .A2(n470), .A4(n680), .S0(n406), 
        .S1(n330), .Y(n609) );
  MUX41X1_HVT U105 ( .A1(n487), .A3(n669), .A2(n608), .A4(n477), .S0(n406), 
        .S1(n380), .Y(n607) );
  OA21X1_HVT U109 ( .A1(n469), .A2(n439), .A3(n353), .Y(n604) );
  NAND2X0_HVT U110 ( .A1(n48), .A2(n602), .Y(n603) );
  MUX41X1_HVT U114 ( .A1(n599), .A3(n605), .A2(n601), .A4(n604), .S0(n440), 
        .S1(n380), .Y(n598) );
  AO21X1_HVT U118 ( .A1(n411), .A2(n424), .A3(n366), .Y(n595) );
  NAND2X0_HVT U123 ( .A1(n589), .A2(n588), .Y(n590) );
  MUX41X1_HVT U131 ( .A1(n581), .A3(n583), .A2(n582), .A4(n584), .S0(n440), 
        .S1(n445), .Y(n580) );
  AND2X1_HVT U154 ( .A1(n415), .A2(n305), .Y(n560) );
  NAND2X0_HVT U158 ( .A1(n357), .A2(n336), .Y(n556) );
  MUX41X1_HVT U159 ( .A1(n701), .A3(n364), .A2(n556), .A4(n495), .S0(n405), 
        .S1(n340), .Y(n555) );
  AND2X1_HVT U162 ( .A1(n365), .A2(n642), .Y(n552) );
  MUX41X1_HVT U165 ( .A1(n693), .A3(n486), .A2(n670), .A4(n550), .S0(n445), 
        .S1(n409), .Y(n549) );
  NAND2X0_HVT U166 ( .A1(n319), .A2(n659), .Y(n548) );
  NAND2X0_HVT U167 ( .A1(n452), .A2(n337), .Y(n547) );
  MUX41X1_HVT U168 ( .A1(n466), .A3(n425), .A2(n547), .A4(n548), .S0(n405), 
        .S1(n446), .Y(n546) );
  MUX41X1_HVT U172 ( .A1(n543), .A3(n549), .A2(n546), .A4(n551), .S0(n416), 
        .S1(n372), .Y(n542) );
  NAND2X0_HVT U174 ( .A1(n434), .A2(n366), .Y(n700) );
  MUX41X1_HVT U176 ( .A1(n419), .A3(n541), .A2(n464), .A4(n283), .S0(n380), 
        .S1(n411), .Y(n540) );
  NAND2X0_HVT U177 ( .A1(n434), .A2(n419), .Y(n539) );
  MUX41X1_HVT U178 ( .A1(n696), .A3(n539), .A2(n484), .A4(n388), .S0(n408), 
        .S1(n445), .Y(n538) );
  MUX41X1_HVT U179 ( .A1(n687), .A3(n483), .A2(n467), .A4(n484), .S0(n405), 
        .S1(n340), .Y(n537) );
  MUX41X1_HVT U182 ( .A1(n473), .A3(n426), .A2(n455), .A4(n345), .S0(n445), 
        .S1(n409), .Y(n534) );
  MUX41X1_HVT U189 ( .A1(n528), .A3(n283), .A2(n529), .A4(n477), .S0(n413), 
        .S1(n437), .Y(n527) );
  MUX41X1_HVT U194 ( .A1(n675), .A3(n688), .A2(n334), .A4(n425), .S0(n413), 
        .S1(n409), .Y(n523) );
  MUX41X1_HVT U195 ( .A1(n365), .A3(n491), .A2(n320), .A4(n678), .S0(n405), 
        .S1(n446), .Y(n522) );
  AO21X1_HVT U197 ( .A1(n400), .A2(n414), .A3(n488), .Y(n520) );
  MUX41X1_HVT U204 ( .A1(n660), .A3(n701), .A2(n494), .A4(n692), .S0(n405), 
        .S1(n444), .Y(n513) );
  NAND2X0_HVT U208 ( .A1(n434), .A2(n427), .Y(n602) );
  NAND2X0_HVT U212 ( .A1(n374), .A2(n423), .Y(n659) );
  NAND2X0_HVT U214 ( .A1(n365), .A2(n312), .Y(n510) );
  NAND2X0_HVT U215 ( .A1(n602), .A2(n425), .Y(n509) );
  NAND2X0_HVT U218 ( .A1(n350), .A2(n356), .Y(n563) );
  NAND2X0_HVT U220 ( .A1(n414), .A2(n510), .Y(n634) );
  INVX0_HVT U241 ( .A(n691), .Y(n498) );
  INVX0_HVT U242 ( .A(n674), .Y(n497) );
  INVX0_HVT U245 ( .A(n707), .Y(n495) );
  INVX0_HVT U252 ( .A(n659), .Y(n492) );
  INVX0_HVT U253 ( .A(n506), .Y(n491) );
  INVX0_HVT U256 ( .A(n563), .Y(n488) );
  INVX0_HVT U264 ( .A(n680), .Y(n481) );
  INVX0_HVT U267 ( .A(n702), .Y(n479) );
  INVX0_HVT U268 ( .A(n693), .Y(n478) );
  INVX0_HVT U270 ( .A(n509), .Y(n477) );
  INVX0_HVT U271 ( .A(n602), .Y(n476) );
  INVX0_HVT U280 ( .A(n686), .Y(n470) );
  INVX0_HVT U283 ( .A(n701), .Y(n468) );
  INVX0_HVT U284 ( .A(n510), .Y(n467) );
  INVX0_HVT U285 ( .A(n507), .Y(n466) );
  INVX0_HVT U289 ( .A(n611), .Y(n464) );
  INVX0_HVT U295 ( .A(n709), .Y(n460) );
  INVX0_HVT U296 ( .A(n698), .Y(n459) );
  INVX0_HVT U299 ( .A(n694), .Y(n456) );
  INVX0_HVT U300 ( .A(n675), .Y(n455) );
  INVX0_HVT U306 ( .A(n547), .Y(n451) );
  NBUFFX2_HVT U1 ( .A(n482), .Y(n420) );
  NBUFFX2_HVT U2 ( .A(n121), .Y(n361) );
  MUX21X1_HVT U3 ( .A1(n428), .A2(n365), .S0(n433), .Y(n678) );
  INVX1_HVT U6 ( .A(n404), .Y(n405) );
  MUX21X1_HVT U7 ( .A1(n317), .A2(n369), .S0(n432), .Y(n553) );
  INVX1_HVT U8 ( .A(n685), .Y(n486) );
  MUX21X1_HVT U9 ( .A1(n424), .A2(n368), .S0(n432), .Y(n608) );
  OA21X1_HVT U10 ( .A1(n448), .A2(n706), .A3(n363), .Y(n516) );
  INVX1_HVT U11 ( .A(n424), .Y(n490) );
  MUX21X1_HVT U12 ( .A1(n344), .A2(n343), .S0(n314), .Y(n576) );
  INVX1_HVT U14 ( .A(n366), .Y(n369) );
  MUX21X1_HVT U16 ( .A1(n603), .A2(n684), .S0(n293), .Y(n601) );
  MUX21X1_HVT U17 ( .A1(n520), .A2(n521), .S0(n293), .Y(n519) );
  INVX1_HVT U18 ( .A(in[1]), .Y(n436) );
  INVX0_HVT U19 ( .A(n121), .Y(n337) );
  INVX1_HVT U20 ( .A(n417), .Y(n19) );
  AND2X1_HVT U22 ( .A1(n212), .A2(n213), .Y(n7) );
  INVX1_HVT U23 ( .A(n364), .Y(n366) );
  INVX1_HVT U25 ( .A(n147), .Y(n432) );
  MUX41X1_HVT U26 ( .A1(n552), .A3(n354), .A2(n553), .A4(n399), .S0(n404), 
        .S1(n444), .Y(n551) );
  INVX0_HVT U27 ( .A(n387), .Y(n572) );
  INVX1_HVT U28 ( .A(n363), .Y(n388) );
  MUX21X1_HVT U29 ( .A1(n487), .A2(n685), .S0(n408), .Y(n584) );
  INVX1_HVT U30 ( .A(n147), .Y(n356) );
  INVX1_HVT U31 ( .A(n147), .Y(n434) );
  INVX1_HVT U32 ( .A(n418), .Y(n355) );
  INVX1_HVT U34 ( .A(n417), .Y(n496) );
  INVX1_HVT U35 ( .A(n23), .Y(n550) );
  INVX1_HVT U36 ( .A(n147), .Y(n373) );
  XNOR2X1_HVT U37 ( .A1(n361), .A2(n422), .Y(n669) );
  MUX41X1_HVT U38 ( .A1(n514), .A3(n515), .A2(n512), .A4(n513), .S0(n412), 
        .S1(n304), .Y(n511) );
  INVX1_HVT U39 ( .A(n496), .Y(n324) );
  MUX21X1_HVT U40 ( .A1(n423), .A2(n211), .S0(n373), .Y(n23) );
  INVX0_HVT U41 ( .A(n423), .Y(n350) );
  NBUFFX2_HVT U43 ( .A(n710), .Y(n39) );
  NBUFFX2_HVT U44 ( .A(n437), .Y(n407) );
  XNOR2X1_HVT U45 ( .A1(n346), .A2(n337), .Y(n345) );
  MUX21X1_HVT U46 ( .A1(n333), .A2(n336), .S0(n433), .Y(n679) );
  NAND2X0_HVT U47 ( .A1(n317), .A2(n435), .Y(n309) );
  INVX1_HVT U48 ( .A(n367), .Y(n368) );
  INVX1_HVT U49 ( .A(n679), .Y(n485) );
  INVX1_HVT U50 ( .A(n364), .Y(n365) );
  INVX1_HVT U52 ( .A(n447), .Y(n446) );
  INVX1_HVT U54 ( .A(n408), .Y(n282) );
  OA21X1_HVT U55 ( .A1(n451), .A2(n448), .A3(n684), .Y(n569) );
  MUX21X1_HVT U59 ( .A1(n679), .A2(n453), .S0(n404), .Y(n344) );
  MUX21X1_HVT U60 ( .A1(n692), .A2(n473), .S0(n414), .Y(n575) );
  XOR2X1_HVT U61 ( .A1(n374), .A2(n409), .Y(n668) );
  MUX21X1_HVT U63 ( .A1(n422), .A2(n317), .S0(n433), .Y(n703) );
  INVX1_HVT U64 ( .A(n703), .Y(n493) );
  INVX1_HVT U65 ( .A(n398), .Y(n266) );
  INVX1_HVT U67 ( .A(n405), .Y(n358) );
  OA21X1_HVT U70 ( .A1(n402), .A2(n448), .A3(n684), .Y(n544) );
  NAND2X0_HVT U71 ( .A1(n472), .A2(n282), .Y(n359) );
  MUX21X1_HVT U72 ( .A1(n352), .A2(n680), .S0(n440), .Y(n665) );
  INVX1_HVT U75 ( .A(n699), .Y(n457) );
  AO21X1_HVT U76 ( .A1(n415), .A2(n621), .A3(n488), .Y(n622) );
  MUX21X1_HVT U78 ( .A1(n384), .A2(n699), .S0(n411), .Y(n615) );
  AO21X1_HVT U79 ( .A1(n329), .A2(n350), .A3(n448), .Y(n612) );
  AND3X1_HVT U80 ( .A1(n48), .A2(n659), .A3(n634), .Y(n635) );
  NAND2X0_HVT U81 ( .A1(n435), .A2(n211), .Y(n710) );
  OA21X1_HVT U84 ( .A1(n676), .A2(n448), .A3(n563), .Y(n564) );
  MUX21X1_HVT U87 ( .A1(n399), .A2(n462), .S0(n407), .Y(n582) );
  AND3X1_HVT U88 ( .A1(n410), .A2(n329), .A3(n333), .Y(n583) );
  MUX21X1_HVT U89 ( .A1(n646), .A2(n672), .S0(n293), .Y(n645) );
  MUX21X1_HVT U90 ( .A1(n570), .A2(n569), .S0(n410), .Y(n568) );
  MUX21X1_HVT U91 ( .A1(n579), .A2(n449), .S0(n293), .Y(n578) );
  INVX1_HVT U92 ( .A(n410), .Y(n293) );
  INVX1_HVT U93 ( .A(n412), .Y(n362) );
  INVX1_HVT U94 ( .A(n437), .Y(n404) );
  NBUFFX2_HVT U95 ( .A(n443), .Y(n414) );
  NBUFFX2_HVT U98 ( .A(n443), .Y(n413) );
  INVX1_HVT U99 ( .A(n440), .Y(n311) );
  INVX1_HVT U100 ( .A(n447), .Y(n445) );
  INVX1_HVT U102 ( .A(in[7]), .Y(n448) );
  INVX1_HVT U104 ( .A(n447), .Y(n340) );
  INVX1_HVT U106 ( .A(n415), .Y(n339) );
  INVX1_HVT U107 ( .A(n362), .Y(n372) );
  INVX1_HVT U108 ( .A(n436), .Y(n435) );
  INVX1_HVT U111 ( .A(n210), .Y(n364) );
  INVX1_HVT U112 ( .A(n447), .Y(n444) );
  MUX21X1_HVT U113 ( .A1(n319), .A2(n423), .S0(n432), .Y(n684) );
  INVX0_HVT U115 ( .A(n684), .Y(n384) );
  INVX0_HVT U116 ( .A(n708), .Y(n313) );
  INVX1_HVT U117 ( .A(in[7]), .Y(n447) );
  INVX1_HVT U119 ( .A(in[6]), .Y(n371) );
  MUX41X1_HVT U120 ( .A1(n705), .A3(n460), .A2(n396), .A4(n701), .S0(n314), 
        .S1(n411), .Y(n536) );
  MUX21X1_HVT U121 ( .A1(n613), .A2(n449), .S0(n410), .Y(n610) );
  NBUFFX2_HVT U122 ( .A(n711), .Y(n48) );
  INVX0_HVT U124 ( .A(n712), .Y(n318) );
  INVX1_HVT U125 ( .A(n335), .Y(n642) );
  NOR2X0_HVT U126 ( .A1(n337), .A2(n318), .Y(n335) );
  MUX21X1_HVT U127 ( .A1(n429), .A2(n425), .S0(n433), .Y(n699) );
  INVX1_HVT U128 ( .A(n436), .Y(n121) );
  INVX1_HVT U129 ( .A(n121), .Y(n147) );
  NAND2X0_HVT U130 ( .A1(n212), .A2(n213), .Y(n210) );
  INVX1_HVT U132 ( .A(n419), .Y(n346) );
  MUX21X1_HVT U133 ( .A1(n313), .A2(n333), .S0(n361), .Y(n683) );
  MUX21X1_HVT U134 ( .A1(n333), .A2(n211), .S0(n433), .Y(n694) );
  INVX0_HVT U135 ( .A(n692), .Y(n463) );
  XOR2X1_HVT U136 ( .A1(n434), .A2(n350), .Y(n671) );
  MUX41X1_HVT U137 ( .A1(n618), .A3(n617), .A2(n625), .A4(n620), .S0(n311), 
        .S1(n416), .Y(n616) );
  INVX0_HVT U138 ( .A(n436), .Y(n374) );
  MUX41X1_HVT U139 ( .A1(n561), .A3(n555), .A2(n562), .A4(n557), .S0(n304), 
        .S1(n372), .Y(n554) );
  INVX1_HVT U140 ( .A(n705), .Y(n480) );
  MUX21X1_HVT U141 ( .A1(n428), .A2(n352), .S0(n434), .Y(n705) );
  MUX41X1_HVT U142 ( .A1(n610), .A3(n607), .A2(n614), .A4(n609), .S0(n304), 
        .S1(n372), .Y(n606) );
  INVX0_HVT U143 ( .A(n678), .Y(n469) );
  NAND2X0_HVT U144 ( .A1(n324), .A2(n420), .Y(n211) );
  INVX0_HVT U145 ( .A(n683), .Y(n471) );
  NAND2X0_HVT U146 ( .A1(n355), .A2(n19), .Y(n212) );
  NAND2X0_HVT U147 ( .A1(in[4]), .A2(n324), .Y(n213) );
  MUX21X1_HVT U148 ( .A1(n682), .A2(n395), .S0(n404), .Y(n343) );
  MUX41X1_HVT U149 ( .A1(n632), .A3(n628), .A2(n633), .A4(n630), .S0(n304), 
        .S1(n372), .Y(n627) );
  MUX21X1_HVT U150 ( .A1(n636), .A2(n635), .S0(n411), .Y(n633) );
  MUX41X1_HVT U151 ( .A1(n534), .A3(n531), .A2(n530), .A4(n527), .S0(n311), 
        .S1(n304), .Y(n526) );
  MUX21X1_HVT U152 ( .A1(n333), .A2(n320), .S0(n337), .Y(n687) );
  INVX1_HVT U153 ( .A(n147), .Y(n357) );
  INVX1_HVT U155 ( .A(n687), .Y(n487) );
  MUX21X1_HVT U156 ( .A1(n694), .A2(n425), .S0(n415), .Y(n636) );
  MUX21X1_HVT U157 ( .A1(n370), .A2(n424), .S0(n434), .Y(n334) );
  INVX0_HVT U160 ( .A(n318), .Y(n319) );
  MUX21X1_HVT U161 ( .A1(n696), .A2(n471), .S0(n408), .Y(n581) );
  INVX0_HVT U163 ( .A(n697), .Y(n462) );
  MUX21X1_HVT U164 ( .A1(n497), .A2(n484), .S0(n414), .Y(n521) );
  MUX41X1_HVT U169 ( .A1(n519), .A3(n523), .A2(n522), .A4(n524), .S0(n416), 
        .S1(n372), .Y(n518) );
  INVX0_HVT U170 ( .A(n345), .Y(n689) );
  NAND2X0_HVT U171 ( .A1(n475), .A2(n413), .Y(n216) );
  NAND2X0_HVT U173 ( .A1(n388), .A2(n377), .Y(n217) );
  NAND2X0_HVT U175 ( .A1(n216), .A2(n217), .Y(n558) );
  INVX0_HVT U180 ( .A(n621), .Y(n475) );
  INVX0_HVT U181 ( .A(n413), .Y(n377) );
  NAND2X0_HVT U183 ( .A1(n511), .A2(n371), .Y(n381) );
  MUX21X1_HVT U184 ( .A1(n355), .A2(n423), .S0(n432), .Y(n354) );
  NAND2X0_HVT U185 ( .A1(n564), .A2(n282), .Y(n218) );
  NAND2X0_HVT U186 ( .A1(n565), .A2(n411), .Y(n219) );
  NAND2X0_HVT U187 ( .A1(n218), .A2(n219), .Y(n562) );
  INVX1_HVT U188 ( .A(n504), .Y(n465) );
  MUX21X1_HVT U190 ( .A1(n465), .A2(n490), .S0(n414), .Y(n565) );
  NAND2X0_HVT U191 ( .A1(n586), .A2(n311), .Y(n227) );
  NAND2X0_HVT U192 ( .A1(n587), .A2(n412), .Y(n231) );
  NAND2X0_HVT U193 ( .A1(n227), .A2(n231), .Y(n585) );
  MUX21X1_HVT U196 ( .A1(n591), .A2(n590), .S0(n414), .Y(n587) );
  MUX41X1_HVT U198 ( .A1(n346), .A3(n39), .A2(n483), .A4(n384), .S0(n405), 
        .S1(n380), .Y(n512) );
  INVX1_HVT U199 ( .A(n351), .Y(n676) );
  NAND2X0_HVT U200 ( .A1(n658), .A2(n438), .Y(n232) );
  NAND2X0_HVT U201 ( .A1(n656), .A2(n358), .Y(n236) );
  NAND2X0_HVT U202 ( .A1(n232), .A2(n236), .Y(n655) );
  INVX1_HVT U203 ( .A(n500), .Y(n484) );
  NAND2X0_HVT U205 ( .A1(n594), .A2(n311), .Y(n238) );
  NAND2X0_HVT U206 ( .A1(n597), .A2(n440), .Y(n239) );
  NAND2X0_HVT U207 ( .A1(n238), .A2(n239), .Y(n593) );
  MUX21X1_HVT U209 ( .A1(n595), .A2(n596), .S0(n414), .Y(n594) );
  MUX21X1_HVT U210 ( .A1(n481), .A2(n494), .S0(n407), .Y(n596) );
  NAND2X0_HVT U211 ( .A1(n662), .A2(n293), .Y(n240) );
  NAND2X0_HVT U213 ( .A1(n666), .A2(n410), .Y(n243) );
  NAND2X0_HVT U216 ( .A1(n240), .A2(n243), .Y(n661) );
  NAND2X0_HVT U217 ( .A1(n516), .A2(n358), .Y(n249) );
  NAND2X0_HVT U219 ( .A1(n517), .A2(n409), .Y(n257) );
  NAND2X0_HVT U221 ( .A1(n249), .A2(n257), .Y(n515) );
  MUX21X1_HVT U222 ( .A1(n697), .A2(n396), .S0(n413), .Y(n517) );
  NAND2X0_HVT U223 ( .A1(n652), .A2(n282), .Y(n261) );
  NAND2X0_HVT U224 ( .A1(n654), .A2(n409), .Y(n264) );
  NAND2X0_HVT U225 ( .A1(n261), .A2(n264), .Y(n651) );
  NAND2X0_HVT U226 ( .A1(n430), .A2(n266), .Y(n269) );
  NAND2X0_HVT U227 ( .A1(n624), .A2(n398), .Y(n273) );
  NAND2X0_HVT U228 ( .A1(n269), .A2(n273), .Y(n623) );
  NAND2X0_HVT U229 ( .A1(n622), .A2(n358), .Y(n279) );
  NAND2X0_HVT U230 ( .A1(n623), .A2(n411), .Y(n280) );
  NAND2X0_HVT U231 ( .A1(n279), .A2(n280), .Y(n620) );
  MUX41X1_HVT U232 ( .A1(n578), .A3(n576), .A2(n577), .A4(n574), .S0(n304), 
        .S1(n311), .Y(n573) );
  MUX41X1_HVT U233 ( .A1(n642), .A3(n453), .A2(n670), .A4(n492), .S0(n282), 
        .S1(n330), .Y(n567) );
  NBUFFX2_HVT U234 ( .A(n700), .Y(n283) );
  INVX0_HVT U235 ( .A(n39), .Y(n458) );
  MUX21X1_HVT U236 ( .A1(n421), .A2(n368), .S0(n337), .Y(n697) );
  INVX0_HVT U237 ( .A(n383), .Y(n597) );
  INVX1_HVT U238 ( .A(in[0]), .Y(n304) );
  NAND2X0_HVT U239 ( .A1(n535), .A2(in[6]), .Y(n297) );
  NAND2X0_HVT U240 ( .A1(n526), .A2(n371), .Y(n299) );
  NAND2X0_HVT U243 ( .A1(n299), .A2(n297), .Y(out[6]) );
  NAND2X0_HVT U244 ( .A1(n559), .A2(n438), .Y(n301) );
  NAND2X0_HVT U246 ( .A1(n558), .A2(n293), .Y(n303) );
  NAND2X0_HVT U247 ( .A1(n301), .A2(n303), .Y(n557) );
  MUX21X1_HVT U248 ( .A1(n560), .A2(n48), .S0(n398), .Y(n559) );
  INVX0_HVT U249 ( .A(n374), .Y(n329) );
  INVX1_HVT U250 ( .A(n499), .Y(n483) );
  MUX41X1_HVT U251 ( .A1(n585), .A3(n598), .A2(n580), .A4(n593), .S0(in[6]), 
        .S1(n304), .Y(out[3]) );
  NBUFFX2_HVT U254 ( .A(in[4]), .Y(n418) );
  INVX1_HVT U255 ( .A(n421), .Y(n305) );
  NBUFFX2_HVT U257 ( .A(in[3]), .Y(n417) );
  MUX21X1_HVT U258 ( .A1(n329), .A2(n39), .S0(n293), .Y(n588) );
  INVX1_HVT U259 ( .A(n436), .Y(n433) );
  NAND2X0_HVT U260 ( .A1(n688), .A2(n444), .Y(n307) );
  NAND2X0_HVT U261 ( .A1(n306), .A2(n447), .Y(n308) );
  NAND2X0_HVT U262 ( .A1(n307), .A2(n308), .Y(n672) );
  INVX0_HVT U263 ( .A(n688), .Y(n306) );
  NAND2X0_HVT U265 ( .A1(n452), .A2(n312), .Y(n310) );
  NAND2X0_HVT U266 ( .A1(n309), .A2(n310), .Y(n688) );
  INVX1_HVT U269 ( .A(n211), .Y(n452) );
  INVX0_HVT U272 ( .A(n435), .Y(n312) );
  INVX0_HVT U273 ( .A(n415), .Y(n314) );
  NAND2X0_HVT U274 ( .A1(n554), .A2(in[6]), .Y(n347) );
  INVX1_HVT U275 ( .A(n422), .Y(n352) );
  MUX21X1_HVT U276 ( .A1(n425), .A2(n426), .S0(n373), .Y(n353) );
  INVX0_HVT U277 ( .A(n448), .Y(n380) );
  INVX1_HVT U278 ( .A(n339), .Y(n330) );
  OR2X1_HVT U279 ( .A1(n346), .A2(n314), .Y(n316) );
  NAND2X0_HVT U281 ( .A1(n458), .A2(n330), .Y(n331) );
  NBUFFX2_HVT U282 ( .A(n443), .Y(n415) );
  INVX1_HVT U286 ( .A(n682), .Y(n472) );
  NAND2X0_HVT U287 ( .A1(n305), .A2(n314), .Y(n315) );
  NAND2X0_HVT U288 ( .A1(n315), .A2(n316), .Y(n624) );
  MUX41X1_HVT U290 ( .A1(n674), .A3(n670), .A2(n626), .A4(n454), .S0(n282), 
        .S1(n446), .Y(n625) );
  NBUFFX2_HVT U291 ( .A(n482), .Y(n419) );
  MUX41X1_HVT U292 ( .A1(n351), .A3(n679), .A2(n683), .A4(n702), .S0(n358), 
        .S1(n340), .Y(n514) );
  INVX0_HVT U293 ( .A(n354), .Y(n696) );
  INVX1_HVT U294 ( .A(n431), .Y(n317) );
  INVX1_HVT U297 ( .A(n318), .Y(n320) );
  MUX21X1_HVT U298 ( .A1(n324), .A2(n7), .S0(n337), .Y(n692) );
  INVX0_HVT U301 ( .A(n338), .Y(n695) );
  MUX41X1_HVT U302 ( .A1(n463), .A3(n697), .A2(n366), .A4(n631), .S0(n444), 
        .S1(n406), .Y(n630) );
  NAND2X0_HVT U303 ( .A1(n600), .A2(n321), .Y(n322) );
  NAND2X0_HVT U304 ( .A1(n48), .A2(n668), .Y(n323) );
  NAND2X0_HVT U305 ( .A1(n322), .A2(n323), .Y(n599) );
  INVX0_HVT U307 ( .A(n668), .Y(n321) );
  NAND2X0_HVT U308 ( .A1(n709), .A2(n438), .Y(n325) );
  NAND2X0_HVT U309 ( .A1(n575), .A2(n282), .Y(n326) );
  NAND2X0_HVT U310 ( .A1(n326), .A2(n325), .Y(n574) );
  NAND2X0_HVT U311 ( .A1(n305), .A2(n312), .Y(n327) );
  NAND2X0_HVT U312 ( .A1(n313), .A2(n357), .Y(n328) );
  NAND2X0_HVT U313 ( .A1(n327), .A2(n328), .Y(n677) );
  INVX0_HVT U314 ( .A(n677), .Y(n473) );
  MUX21X1_HVT U315 ( .A1(n419), .A2(n313), .S0(n329), .Y(n502) );
  NAND2X0_HVT U316 ( .A1(n686), .A2(n339), .Y(n332) );
  NAND2X0_HVT U317 ( .A1(n331), .A2(n332), .Y(n570) );
  MUX21X1_HVT U318 ( .A1(n420), .A2(n313), .S0(n435), .Y(n686) );
  MUX41X1_HVT U319 ( .A1(n489), .A3(n492), .A2(n450), .A4(n452), .S0(n282), 
        .S1(n445), .Y(n640) );
  OR2X1_HVT U320 ( .A1(n346), .A2(n374), .Y(n680) );
  INVX1_HVT U321 ( .A(n505), .Y(n489) );
  NBUFFX2_HVT U322 ( .A(in[4]), .Y(n333) );
  INVX1_HVT U323 ( .A(n431), .Y(n336) );
  INVX1_HVT U324 ( .A(n681), .Y(n494) );
  OA21X1_HVT U325 ( .A1(n681), .A2(n448), .A3(n463), .Y(n532) );
  MUX41X1_HVT U326 ( .A1(n490), .A3(n334), .A2(n688), .A4(n707), .S0(n404), 
        .S1(n444), .Y(n577) );
  INVX0_HVT U327 ( .A(n418), .Y(n482) );
  MUX41X1_HVT U328 ( .A1(n568), .A3(n567), .A2(n572), .A4(n571), .S0(n311), 
        .S1(n416), .Y(n566) );
  MUX21X1_HVT U329 ( .A1(n211), .A2(n421), .S0(n373), .Y(n338) );
  MUX41X1_HVT U330 ( .A1(n667), .A3(n674), .A2(n525), .A4(n680), .S0(n377), 
        .S1(n411), .Y(n524) );
  INVX0_HVT U331 ( .A(n447), .Y(n443) );
  INVX0_HVT U332 ( .A(n502), .Y(n474) );
  MUX41X1_HVT U333 ( .A1(n385), .A3(n468), .A2(n384), .A4(n690), .S0(n358), 
        .S1(n340), .Y(n383) );
  NAND2X0_HVT U334 ( .A1(n533), .A2(n438), .Y(n341) );
  NAND2X0_HVT U335 ( .A1(n532), .A2(n358), .Y(n342) );
  NAND2X0_HVT U336 ( .A1(n341), .A2(n342), .Y(n531) );
  MUX41X1_HVT U337 ( .A1(n459), .A3(n653), .A2(n457), .A4(n468), .S0(n339), 
        .S1(n412), .Y(n652) );
  INVX1_HVT U338 ( .A(n501), .Y(n453) );
  NAND2X0_HVT U339 ( .A1(n542), .A2(n371), .Y(n348) );
  NAND2X0_HVT U340 ( .A1(n347), .A2(n348), .Y(out[5]) );
  INVX0_HVT U341 ( .A(n349), .Y(n579) );
  MUX21X1_HVT U342 ( .A1(n350), .A2(n502), .S0(n339), .Y(n349) );
  MUX21X1_HVT U343 ( .A1(n352), .A2(n430), .S0(n435), .Y(n351) );
  INVX1_HVT U344 ( .A(n690), .Y(n450) );
  XOR2X2_HVT U345 ( .A1(n365), .A2(n357), .Y(n670) );
  MUX41X1_HVT U346 ( .A1(n645), .A3(n640), .A2(n641), .A4(n638), .S0(n304), 
        .S1(n311), .Y(n637) );
  MUX41X1_HVT U347 ( .A1(n677), .A3(n401), .A2(n670), .A4(n642), .S0(n358), 
        .S1(n446), .Y(n530) );
  INVX1_HVT U348 ( .A(n508), .Y(n454) );
  NAND2X0_HVT U349 ( .A1(n606), .A2(n371), .Y(n393) );
  MUX21X1_HVT U350 ( .A1(n685), .A2(n509), .S0(n413), .Y(n503) );
  MUX21X1_HVT U351 ( .A1(n421), .A2(n333), .S0(n356), .Y(n685) );
  NAND2X0_HVT U352 ( .A1(n592), .A2(n408), .Y(n360) );
  NAND2X0_HVT U353 ( .A1(n359), .A2(n360), .Y(n591) );
  INVX1_HVT U354 ( .A(n503), .Y(n449) );
  MUX41X1_HVT U355 ( .A1(n353), .A3(n402), .A2(n657), .A4(n403), .S0(n314), 
        .S1(n362), .Y(n656) );
  MUX21X1_HVT U356 ( .A1(n319), .A2(n426), .S0(n361), .Y(n363) );
  MUX41X1_HVT U357 ( .A1(n693), .A3(n461), .A2(n403), .A4(n474), .S0(n446), 
        .S1(n407), .Y(n586) );
  INVX1_HVT U358 ( .A(n7), .Y(n367) );
  INVX1_HVT U359 ( .A(n367), .Y(n370) );
  INVX1_HVT U360 ( .A(n706), .Y(n461) );
  MUX21X1_HVT U361 ( .A1(n7), .A2(n336), .S0(n361), .Y(n706) );
  MUX41X1_HVT U362 ( .A1(n462), .A3(n370), .A2(n397), .A4(n354), .S0(n444), 
        .S1(n362), .Y(n654) );
  MUX41X1_HVT U363 ( .A1(n463), .A3(n369), .A2(n476), .A4(n425), .S0(n437), 
        .S1(in[7]), .Y(n571) );
  INVX1_HVT U364 ( .A(n386), .Y(n392) );
  MUX41X1_HVT U365 ( .A1(n481), .A3(n430), .A2(n397), .A4(n603), .S0(n282), 
        .S1(n377), .Y(n561) );
  MUX41X1_HVT U366 ( .A1(n538), .A3(n536), .A2(n540), .A4(n537), .S0(n304), 
        .S1(n372), .Y(n535) );
  NAND2X0_HVT U367 ( .A1(n627), .A2(n371), .Y(n375) );
  NAND2X0_HVT U368 ( .A1(n637), .A2(in[6]), .Y(n376) );
  NAND2X0_HVT U369 ( .A1(n375), .A2(n376), .Y(out[1]) );
  NAND2X0_HVT U370 ( .A1(n566), .A2(n371), .Y(n378) );
  NAND2X0_HVT U371 ( .A1(n573), .A2(in[6]), .Y(n379) );
  NAND2X0_HVT U372 ( .A1(n379), .A2(n378), .Y(out[4]) );
  NAND2X0_HVT U373 ( .A1(n518), .A2(in[6]), .Y(n382) );
  NAND2X0_HVT U374 ( .A1(n381), .A2(n382), .Y(out[7]) );
  NAND2X0_HVT U375 ( .A1(n373), .A2(n368), .Y(n385) );
  XOR2X1_HVT U376 ( .A1(n404), .A2(n448), .Y(n386) );
  MUX41X1_HVT U377 ( .A1(n389), .A3(n683), .A2(n450), .A4(n388), .S0(n408), 
        .S1(n448), .Y(n387) );
  NAND2X0_HVT U378 ( .A1(n424), .A2(n337), .Y(n389) );
  NAND2X0_HVT U379 ( .A1(n615), .A2(n386), .Y(n390) );
  NAND2X0_HVT U380 ( .A1(n397), .A2(n392), .Y(n391) );
  NAND2X0_HVT U381 ( .A1(n390), .A2(n391), .Y(n614) );
  NAND2X0_HVT U382 ( .A1(n616), .A2(in[6]), .Y(n394) );
  NAND2X0_HVT U383 ( .A1(n394), .A2(n393), .Y(out[2]) );
  INVX1_HVT U384 ( .A(n442), .Y(n441) );
  INVX0_HVT U385 ( .A(n439), .Y(n438) );
  INVX1_HVT U386 ( .A(in[5]), .Y(n442) );
  NBUFFX2_HVT U387 ( .A(n708), .Y(n426) );
  NBUFFX2_HVT U388 ( .A(n708), .Y(n427) );
  NBUFFX2_HVT U389 ( .A(n708), .Y(n428) );
  MUX21X1_HVT U390 ( .A1(n480), .A2(n490), .S0(n440), .Y(n648) );
  AND2X1_HVT U391 ( .A1(n48), .A2(n642), .Y(n395) );
  AND2X1_HVT U392 ( .A1(n370), .A2(n659), .Y(n396) );
  AND2X1_HVT U393 ( .A1(n319), .A2(n602), .Y(n397) );
  NAND2X0_HVT U394 ( .A1(n355), .A2(n19), .Y(n708) );
  MUX21X1_HVT U395 ( .A1(n424), .A2(n320), .S0(n410), .Y(n589) );
  MUX21X1_HVT U396 ( .A1(n313), .A2(n452), .S0(n361), .Y(n541) );
  MUX21X1_HVT U397 ( .A1(n317), .A2(n491), .S0(n415), .Y(n646) );
  MUX21X1_HVT U398 ( .A1(n423), .A2(n421), .S0(n356), .Y(n506) );
  MUX21X1_HVT U399 ( .A1(n336), .A2(n421), .S0(n433), .Y(n681) );
  MUX21X1_HVT U400 ( .A1(n366), .A2(n452), .S0(n432), .Y(n690) );
  MUX21X1_HVT U401 ( .A1(n429), .A2(n369), .S0(n374), .Y(n675) );
  MUX21X1_HVT U402 ( .A1(n427), .A2(n422), .S0(n433), .Y(n702) );
  XOR2X1_HVT U403 ( .A1(n429), .A2(n434), .Y(n667) );
  MUX21X1_HVT U404 ( .A1(n421), .A2(n420), .S0(n357), .Y(n525) );
  MUX21X1_HVT U405 ( .A1(n370), .A2(n313), .S0(n373), .Y(n619) );
  MUX21X1_HVT U406 ( .A1(n419), .A2(n422), .S0(n361), .Y(n592) );
  MUX21X1_HVT U407 ( .A1(n545), .A2(n544), .S0(n410), .Y(n543) );
  MUX21X1_HVT U408 ( .A1(n424), .A2(n491), .S0(n415), .Y(n545) );
  MUX21X1_HVT U409 ( .A1(n427), .A2(n424), .S0(n373), .Y(n626) );
  MUX21X1_HVT U410 ( .A1(n425), .A2(n419), .S0(n356), .Y(n644) );
  MUX21X1_HVT U411 ( .A1(n366), .A2(n420), .S0(n357), .Y(n639) );
  MUX21X1_HVT U412 ( .A1(n421), .A2(n319), .S0(n361), .Y(n528) );
  MUX21X1_HVT U413 ( .A1(n319), .A2(n430), .S0(n374), .Y(n529) );
  MUX21X1_HVT U414 ( .A1(n422), .A2(n365), .S0(n361), .Y(n504) );
  MUX21X1_HVT U415 ( .A1(n485), .A2(n39), .S0(n408), .Y(n605) );
  MUX21X1_HVT U416 ( .A1(n370), .A2(n420), .S0(n432), .Y(n611) );
  MUX21X1_HVT U417 ( .A1(n430), .A2(n419), .S0(n357), .Y(n508) );
  MUX21X1_HVT U418 ( .A1(n426), .A2(n320), .S0(n435), .Y(n621) );
  XNOR2X1_HVT U419 ( .A1(n447), .A2(n435), .Y(n398) );
  XNOR2X1_HVT U420 ( .A1(n426), .A2(n356), .Y(n399) );
  XNOR2X1_HVT U421 ( .A1(n319), .A2(n434), .Y(n400) );
  MUX21X1_HVT U422 ( .A1(n429), .A2(n427), .S0(n356), .Y(n501) );
  MUX21X1_HVT U423 ( .A1(n313), .A2(n317), .S0(n440), .Y(n663) );
  XOR2X1_HVT U424 ( .A1(n373), .A2(n412), .Y(n673) );
  AND2X1_HVT U425 ( .A1(n373), .A2(n452), .Y(n401) );
  NBUFFX2_HVT U426 ( .A(n704), .Y(n423) );
  NBUFFX2_HVT U427 ( .A(n704), .Y(n424) );
  NBUFFX2_HVT U428 ( .A(n711), .Y(n429) );
  NBUFFX2_HVT U429 ( .A(n704), .Y(n425) );
  NBUFFX2_HVT U430 ( .A(n19), .Y(n422) );
  NBUFFX2_HVT U431 ( .A(n19), .Y(n421) );
  NBUFFX2_HVT U432 ( .A(n711), .Y(n430) );
  NBUFFX2_HVT U433 ( .A(n712), .Y(n431) );
  NBUFFX2_HVT U434 ( .A(n437), .Y(n408) );
  NBUFFX2_HVT U435 ( .A(n438), .Y(n411) );
  NBUFFX2_HVT U436 ( .A(n441), .Y(n412) );
  NBUFFX2_HVT U437 ( .A(n438), .Y(n410) );
  NBUFFX2_HVT U438 ( .A(n438), .Y(n409) );
  NBUFFX2_HVT U439 ( .A(n438), .Y(n406) );
  MUX21X1_HVT U440 ( .A1(n664), .A2(n665), .S0(n413), .Y(n662) );
  MUX21X1_HVT U441 ( .A1(n333), .A2(n423), .S0(n356), .Y(n500) );
  MUX21X1_HVT U442 ( .A1(n629), .A2(n352), .S0(n414), .Y(n533) );
  MUX21X1_HVT U443 ( .A1(n479), .A2(n312), .S0(n440), .Y(n650) );
  MUX21X1_HVT U444 ( .A1(n333), .A2(n320), .S0(n357), .Y(n499) );
  MUX21X1_HVT U445 ( .A1(n305), .A2(n350), .S0(n357), .Y(n505) );
  MUX21X1_HVT U446 ( .A1(n333), .A2(n365), .S0(n374), .Y(n507) );
  MUX21X1_HVT U447 ( .A1(n352), .A2(n333), .S0(n407), .Y(n600) );
  NAND2X0_HVT U448 ( .A1(n418), .A2(n19), .Y(n704) );
  AND2X1_HVT U449 ( .A1(n369), .A2(n312), .Y(n402) );
  NAND2X0_HVT U450 ( .A1(n417), .A2(n418), .Y(n712) );
  NAND2X0_HVT U451 ( .A1(n324), .A2(n420), .Y(n711) );
  AND2X1_HVT U452 ( .A1(n422), .A2(n329), .Y(n403) );
  INVX1_HVT U453 ( .A(n439), .Y(n437) );
  NBUFFX2_HVT U454 ( .A(n441), .Y(n440) );
  INVX1_HVT U455 ( .A(in[2]), .Y(n439) );
  NBUFFX2_HVT U456 ( .A(in[0]), .Y(n416) );
endmodule

