
module inv_sbox_13 ( in, out );
  input [7:0] in;
  output [7:0] out;
  wire   n5, n196, n197, n198, n199, n200, n201, n202, n205, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615;

  NAND2X0_HVT U1 ( .A1(n266), .A2(n322), .Y(n615) );
  NAND2X0_HVT U4 ( .A1(n237), .A2(n614), .Y(n612) );
  NAND2X0_HVT U7 ( .A1(n339), .A2(n335), .Y(n609) );
  NAND2X0_HVT U8 ( .A1(n341), .A2(n333), .Y(n608) );
  NAND2X0_HVT U9 ( .A1(n297), .A2(n608), .Y(n607) );
  NAND2X0_HVT U10 ( .A1(n300), .A2(n605), .Y(n606) );
  NAND2X0_HVT U12 ( .A1(n280), .A2(n320), .Y(n603) );
  NAND2X0_HVT U13 ( .A1(n336), .A2(n259), .Y(n602) );
  NAND2X0_HVT U15 ( .A1(n330), .A2(n237), .Y(n600) );
  NAND2X0_HVT U19 ( .A1(n237), .A2(n405), .Y(n595) );
  NAND2X0_HVT U32 ( .A1(n323), .A2(n279), .Y(n583) );
  NAND2X0_HVT U35 ( .A1(n608), .A2(n285), .Y(n580) );
  NAND2X0_HVT U38 ( .A1(n320), .A2(n279), .Y(n577) );
  NAND2X0_HVT U42 ( .A1(n610), .A2(n285), .Y(n573) );
  OA21X1_HVT U53 ( .A1(n261), .A2(n565), .A3(n374), .Y(n563) );
  NAND2X0_HVT U55 ( .A1(n336), .A2(n612), .Y(n561) );
  MUX41X1_HVT U56 ( .A1(n387), .A3(n331), .A2(n372), .A4(n561), .S0(n312), 
        .S1(n265), .Y(n560) );
  AO21X1_HVT U60 ( .A1(n555), .A2(n316), .A3(n594), .Y(n556) );
  MUX41X1_HVT U62 ( .A1(n554), .A3(n560), .A2(n558), .A4(n562), .S0(n328), 
        .S1(n326), .Y(n553) );
  MUX41X1_HVT U65 ( .A1(n366), .A3(n368), .A2(n367), .A4(n577), .S0(n312), 
        .S1(n265), .Y(n550) );
  NAND2X0_HVT U66 ( .A1(n280), .A2(n272), .Y(n549) );
  MUX41X1_HVT U67 ( .A1(n363), .A3(n388), .A2(n365), .A4(n549), .S0(n318), 
        .S1(n309), .Y(n548) );
  MUX41X1_HVT U68 ( .A1(n363), .A3(n266), .A2(n364), .A4(n300), .S0(n311), 
        .S1(n265), .Y(n547) );
  MUX41X1_HVT U69 ( .A1(n547), .A3(n550), .A2(n548), .A4(n551), .S0(n328), 
        .S1(in[1]), .Y(n546) );
  NAND2X0_HVT U72 ( .A1(n331), .A2(n609), .Y(n544) );
  MUX41X1_HVT U73 ( .A1(n588), .A3(n544), .A2(n290), .A4(n319), .S0(n317), 
        .S1(n309), .Y(n543) );
  MUX41X1_HVT U74 ( .A1(n606), .A3(n379), .A2(n378), .A4(n369), .S0(n312), 
        .S1(n344), .Y(n542) );
  MUX41X1_HVT U78 ( .A1(n539), .A3(n543), .A2(n542), .A4(n545), .S0(n328), 
        .S1(n325), .Y(n538) );
  MUX41X1_HVT U79 ( .A1(n375), .A3(n597), .A2(n377), .A4(n598), .S0(n312), 
        .S1(n344), .Y(n537) );
  MUX41X1_HVT U80 ( .A1(n390), .A3(n387), .A2(n198), .A4(n289), .S0(n311), 
        .S1(n347), .Y(n536) );
  NAND2X0_HVT U81 ( .A1(n337), .A2(n609), .Y(n535) );
  AND2X1_HVT U82 ( .A1(n610), .A2(n334), .Y(n534) );
  MUX41X1_HVT U83 ( .A1(n534), .A3(n376), .A2(n391), .A4(n535), .S0(n311), 
        .S1(n344), .Y(n533) );
  MUX41X1_HVT U87 ( .A1(n354), .A3(n306), .A2(n393), .A4(n372), .S0(n310), 
        .S1(n344), .Y(n530) );
  MUX41X1_HVT U88 ( .A1(n365), .A3(n351), .A2(n585), .A4(n569), .S0(n311), 
        .S1(n347), .Y(n529) );
  NAND2X0_HVT U89 ( .A1(n257), .A2(n271), .Y(n528) );
  MUX41X1_HVT U96 ( .A1(n388), .A3(n602), .A2(n373), .A4(n394), .S0(n312), 
        .S1(n346), .Y(n521) );
  MUX41X1_HVT U99 ( .A1(n583), .A3(n367), .A2(n567), .A4(n331), .S0(n265), 
        .S1(n313), .Y(n518) );
  NAND2X0_HVT U100 ( .A1(n279), .A2(n402), .Y(n517) );
  MUX41X1_HVT U101 ( .A1(n396), .A3(n603), .A2(n380), .A4(n517), .S0(n265), 
        .S1(n310), .Y(n516) );
  AND2X1_HVT U104 ( .A1(n609), .A2(n332), .Y(n514) );
  MUX41X1_HVT U105 ( .A1(n601), .A3(n397), .A2(n535), .A4(n514), .S0(n312), 
        .S1(n347), .Y(n513) );
  MUX41X1_HVT U107 ( .A1(n396), .A3(n334), .A2(n512), .A4(n356), .S0(n311), 
        .S1(n347), .Y(n511) );
  MUX41X1_HVT U108 ( .A1(n369), .A3(n599), .A2(n372), .A4(n337), .S0(n312), 
        .S1(n346), .Y(n510) );
  MUX41X1_HVT U109 ( .A1(n395), .A3(n351), .A2(n392), .A4(n286), .S0(n311), 
        .S1(n346), .Y(n509) );
  MUX41X1_HVT U110 ( .A1(n509), .A3(n511), .A2(n510), .A4(n513), .S0(n329), 
        .S1(n326), .Y(n508) );
  AO21X1_HVT U112 ( .A1(n383), .A2(n317), .A3(n591), .Y(n506) );
  NAND2X0_HVT U114 ( .A1(n297), .A2(n609), .Y(n504) );
  MUX41X1_HVT U115 ( .A1(n504), .A3(n604), .A2(n383), .A4(n334), .S0(n265), 
        .S1(n312), .Y(n503) );
  MUX41X1_HVT U116 ( .A1(n382), .A3(n375), .A2(n351), .A4(n600), .S0(n310), 
        .S1(n344), .Y(n502) );
  NAND2X0_HVT U118 ( .A1(n279), .A2(n266), .Y(n500) );
  MUX41X1_HVT U119 ( .A1(n398), .A3(n501), .A2(n578), .A4(n500), .S0(n310), 
        .S1(n347), .Y(n499) );
  MUX41X1_HVT U120 ( .A1(n499), .A3(n503), .A2(n502), .A4(n505), .S0(n329), 
        .S1(n326), .Y(n498) );
  MUX41X1_HVT U122 ( .A1(n386), .A3(n302), .A2(n569), .A4(n389), .S0(n310), 
        .S1(n344), .Y(n497) );
  AOI21X1_HVT U127 ( .A1(n315), .A2(n491), .A3(n357), .Y(n492) );
  NAND2X0_HVT U129 ( .A1(n314), .A2(n297), .Y(n489) );
  MUX41X1_HVT U130 ( .A1(n489), .A3(n490), .A2(n493), .A4(n492), .S0(n318), 
        .S1(n326), .Y(n488) );
  AND2X1_HVT U131 ( .A1(n272), .A2(n222), .Y(n487) );
  MUX41X1_HVT U132 ( .A1(n288), .A3(n487), .A2(n400), .A4(n363), .S0(n317), 
        .S1(n309), .Y(n486) );
  MUX41X1_HVT U133 ( .A1(n401), .A3(n356), .A2(n561), .A4(n355), .S0(n316), 
        .S1(n310), .Y(n485) );
  MUX41X1_HVT U136 ( .A1(n566), .A3(n517), .A2(n483), .A4(n361), .S0(n314), 
        .S1(n347), .Y(n482) );
  MUX41X1_HVT U137 ( .A1(n259), .A3(n586), .A2(n590), .A4(n394), .S0(n318), 
        .S1(n309), .Y(n481) );
  MUX41X1_HVT U140 ( .A1(n378), .A3(n303), .A2(n246), .A4(n604), .S0(n317), 
        .S1(n312), .Y(n479) );
  NAND2X0_HVT U141 ( .A1(n330), .A2(n279), .Y(n478) );
  MUX41X1_HVT U142 ( .A1(n478), .A3(n576), .A2(n399), .A4(n246), .S0(n315), 
        .S1(n347), .Y(n477) );
  MUX41X1_HVT U143 ( .A1(n271), .A3(n275), .A2(n595), .A4(n236), .S0(n313), 
        .S1(n346), .Y(n476) );
  MUX41X1_HVT U145 ( .A1(n584), .A3(n397), .A2(n475), .A4(n535), .S0(n315), 
        .S1(n346), .Y(n474) );
  MUX41X1_HVT U146 ( .A1(n474), .A3(n476), .A2(n477), .A4(n479), .S0(n325), 
        .S1(n328), .Y(n473) );
  MUX41X1_HVT U151 ( .A1(n391), .A3(n381), .A2(n370), .A4(n469), .S0(n316), 
        .S1(n311), .Y(n468) );
  MUX41X1_HVT U155 ( .A1(n246), .A3(n604), .A2(n596), .A4(n373), .S0(n313), 
        .S1(n346), .Y(n464) );
  MUX41X1_HVT U156 ( .A1(n464), .A3(n468), .A2(n465), .A4(n470), .S0(n329), 
        .S1(n326), .Y(n463) );
  NAND2X0_HVT U159 ( .A1(n460), .A2(n459), .Y(n461) );
  MUX41X1_HVT U162 ( .A1(n384), .A3(n368), .A2(n580), .A4(n457), .S0(n313), 
        .S1(n347), .Y(n456) );
  NAND2X0_HVT U163 ( .A1(n341), .A2(n271), .Y(n455) );
  NAND2X0_HVT U166 ( .A1(n605), .A2(n451), .Y(n452) );
  MUX41X1_HVT U174 ( .A1(n393), .A3(n561), .A2(n401), .A4(n285), .S0(n313), 
        .S1(n344), .Y(n443) );
  NAND2X0_HVT U177 ( .A1(n228), .A2(n266), .Y(n441) );
  AND2X1_HVT U179 ( .A1(n610), .A2(n332), .Y(n439) );
  MUX41X1_HVT U180 ( .A1(n583), .A3(n349), .A2(n439), .A4(n570), .S0(n313), 
        .S1(n346), .Y(n438) );
  MUX41X1_HVT U183 ( .A1(n275), .A3(n387), .A2(n369), .A4(n573), .S0(n316), 
        .S1(n309), .Y(n435) );
  AND2X1_HVT U185 ( .A1(n285), .A2(n222), .Y(n433) );
  NAND2X0_HVT U191 ( .A1(n287), .A2(n362), .Y(n427) );
  AND2X1_HVT U192 ( .A1(n379), .A2(n425), .Y(n426) );
  NAND2X0_HVT U194 ( .A1(n573), .A2(n425), .Y(n423) );
  MUX41X1_HVT U195 ( .A1(n424), .A3(n423), .A2(n426), .A4(n427), .S0(n311), 
        .S1(n325), .Y(n422) );
  NAND2X0_HVT U198 ( .A1(n340), .A2(n285), .Y(n605) );
  NAND2X0_HVT U200 ( .A1(n332), .A2(n257), .Y(n491) );
  NAND2X0_HVT U207 ( .A1(n279), .A2(n301), .Y(n555) );
  INVX0_HVT U2 ( .A(n614), .Y(n402) );
  INVX1_HVT U3 ( .A(n324), .Y(n325) );
  INVX0_HVT U5 ( .A(n326), .Y(n218) );
  NBUFFX4_HVT U6 ( .A(n407), .Y(n322) );
  OR2X1_HVT U11 ( .A1(n404), .A2(n5), .Y(n613) );
  IBUFFX16_HVT U14 ( .A(in[6]), .Y(n5) );
  INVX1_HVT U16 ( .A(n404), .Y(n266) );
  INVX2_HVT U17 ( .A(n334), .Y(n405) );
  OR2X1_HVT U18 ( .A1(n407), .A2(n196), .Y(n611) );
  IBUFFX16_HVT U20 ( .A(n321), .Y(n196) );
  IBUFFX2_HVT U21 ( .A(n407), .Y(n272) );
  MUX21X1_HVT U22 ( .A1(n337), .A2(n332), .S0(n197), .Y(n409) );
  IBUFFX16_HVT U23 ( .A(n340), .Y(n197) );
  MUX21X2_HVT U24 ( .A1(n301), .A2(n403), .S0(n340), .Y(n587) );
  INVX0_HVT U25 ( .A(n361), .Y(n198) );
  MUX41X1_HVT U26 ( .A1(n456), .A3(n458), .A2(n450), .A4(n454), .S0(n199), 
        .S1(n200), .Y(n449) );
  IBUFFX16_HVT U27 ( .A(n324), .Y(n199) );
  IBUFFX16_HVT U28 ( .A(n224), .Y(n200) );
  MUX21X2_HVT U29 ( .A1(n463), .A2(n473), .S0(in[7]), .Y(out[5]) );
  MUX21X2_HVT U30 ( .A1(n403), .A2(n301), .S0(n280), .Y(n571) );
  INVX0_HVT U31 ( .A(n611), .Y(n271) );
  MUX21X2_HVT U33 ( .A1(n298), .A2(n405), .S0(n280), .Y(n448) );
  INVX0_HVT U34 ( .A(n256), .Y(n457) );
  MUX21X1_HVT U36 ( .A1(n614), .A2(n291), .S0(n338), .Y(n290) );
  IBUFFX2_HVT U37 ( .A(n223), .Y(n279) );
  MUX21X2_HVT U39 ( .A1(n288), .A2(n400), .S0(n201), .Y(n472) );
  IBUFFX16_HVT U40 ( .A(n316), .Y(n201) );
  INVX1_HVT U41 ( .A(n222), .Y(n202) );
  INVX0_HVT U43 ( .A(in[0]), .Y(n222) );
  MUX41X1_HVT U44 ( .A1(n428), .A3(n422), .A2(n437), .A4(n434), .S0(n264), 
        .S1(n205), .Y(out[7]) );
  IBUFFX16_HVT U45 ( .A(n278), .Y(n205) );
  INVX1_HVT U46 ( .A(n342), .Y(n280) );
  INVX0_HVT U47 ( .A(n578), .Y(n381) );
  MUX21X2_HVT U48 ( .A1(n333), .A2(n266), .S0(n258), .Y(n520) );
  INVX1_HVT U49 ( .A(n257), .Y(n258) );
  XNOR2X2_HVT U50 ( .A1(n296), .A2(n338), .Y(n578) );
  NAND2X0_HVT U51 ( .A1(n438), .A2(n218), .Y(n219) );
  NAND2X0_HVT U52 ( .A1(n440), .A2(n326), .Y(n220) );
  NAND2X0_HVT U54 ( .A1(n220), .A2(n219), .Y(n437) );
  INVX0_HVT U57 ( .A(n384), .Y(n221) );
  INVX1_HVT U58 ( .A(n571), .Y(n384) );
  INVX1_HVT U59 ( .A(n348), .Y(n345) );
  INVX2_HVT U61 ( .A(n348), .Y(n347) );
  IBUFFX2_HVT U63 ( .A(n348), .Y(n346) );
  INVX1_HVT U64 ( .A(n342), .Y(n223) );
  IBUFFX16_HVT U70 ( .A(n264), .Y(n224) );
  MUX41X1_HVT U71 ( .A1(n445), .A3(n447), .A2(n443), .A4(n444), .S0(n325), 
        .S1(n225), .Y(n442) );
  IBUFFX16_HVT U75 ( .A(n328), .Y(n225) );
  MUX41X1_HVT U76 ( .A1(n304), .A3(n448), .A2(n307), .A4(n305), .S0(n346), 
        .S1(n248), .Y(n447) );
  MUX21X2_HVT U77 ( .A1(n442), .A2(n449), .S0(n226), .Y(out[6]) );
  IBUFFX16_HVT U84 ( .A(n242), .Y(n226) );
  INVX0_HVT U85 ( .A(n588), .Y(n373) );
  INVX1_HVT U86 ( .A(n339), .Y(n227) );
  INVX2_HVT U90 ( .A(n227), .Y(n228) );
  MUX21X2_HVT U91 ( .A1(n277), .A2(n370), .S0(n229), .Y(n552) );
  IBUFFX16_HVT U92 ( .A(n314), .Y(n229) );
  IBUFFX2_HVT U93 ( .A(n222), .Y(n340) );
  AO21X1_HVT U94 ( .A1(n340), .A2(n402), .A3(n260), .Y(n425) );
  INVX1_HVT U95 ( .A(n409), .Y(n400) );
  NAND2X0_HVT U97 ( .A1(n538), .A2(n230), .Y(n231) );
  NAND2X0_HVT U98 ( .A1(n531), .A2(n278), .Y(n232) );
  NAND2X0_HVT U102 ( .A1(n231), .A2(n232), .Y(out[1]) );
  IBUFFX2_HVT U103 ( .A(n278), .Y(n230) );
  IBUFFX2_HVT U106 ( .A(in[7]), .Y(n278) );
  MUX21X1_HVT U111 ( .A1(n600), .A2(n588), .S0(n234), .Y(n233) );
  IBUFFX16_HVT U113 ( .A(n233), .Y(n564) );
  IBUFFX16_HVT U117 ( .A(n318), .Y(n234) );
  MUX21X1_HVT U121 ( .A1(n563), .A2(n564), .S0(n235), .Y(n562) );
  IBUFFX16_HVT U123 ( .A(n314), .Y(n235) );
  IBUFFX2_HVT U124 ( .A(n600), .Y(n364) );
  NBUFFX2_HVT U125 ( .A(n592), .Y(n236) );
  NBUFFX2_HVT U126 ( .A(n223), .Y(n237) );
  INVX0_HVT U128 ( .A(n253), .Y(n592) );
  INVX1_HVT U134 ( .A(in[0]), .Y(n342) );
  INVX1_HVT U135 ( .A(n223), .Y(n257) );
  MUX21X2_HVT U138 ( .A1(n546), .A2(n553), .S0(n238), .Y(out[0]) );
  IBUFFX16_HVT U139 ( .A(n278), .Y(n238) );
  NAND2X0_HVT U144 ( .A1(n461), .A2(n239), .Y(n240) );
  NAND2X0_HVT U147 ( .A1(n462), .A2(n315), .Y(n241) );
  NAND2X0_HVT U148 ( .A1(n240), .A2(n241), .Y(n458) );
  IBUFFX2_HVT U149 ( .A(n315), .Y(n239) );
  IBUFFX16_HVT U150 ( .A(in[7]), .Y(n242) );
  MUX21X1_HVT U152 ( .A1(n389), .A2(n572), .S0(n255), .Y(n462) );
  INVX1_HVT U153 ( .A(n295), .Y(n247) );
  INVX0_HVT U154 ( .A(n317), .Y(n255) );
  AO21X1_HVT U157 ( .A1(n331), .A2(n277), .A3(n260), .Y(n451) );
  INVX0_HVT U158 ( .A(n607), .Y(n361) );
  NAND2X0_HVT U160 ( .A1(n506), .A2(n248), .Y(n249) );
  MUX21X1_HVT U161 ( .A1(n323), .A2(n330), .S0(n287), .Y(n526) );
  OA21X1_HVT U164 ( .A1(n353), .A2(n260), .A3(n594), .Y(n540) );
  NAND2X0_HVT U165 ( .A1(n279), .A2(n337), .Y(n604) );
  INVX0_HVT U167 ( .A(n402), .Y(n254) );
  INVX1_HVT U168 ( .A(n287), .Y(n265) );
  OA21X1_HVT U169 ( .A1(n352), .A2(n261), .A3(n360), .Y(n466) );
  INVX1_HVT U170 ( .A(n296), .Y(n300) );
  INVX1_HVT U171 ( .A(n327), .Y(n329) );
  INVX1_HVT U172 ( .A(n329), .Y(n264) );
  INVX1_HVT U173 ( .A(n615), .Y(n296) );
  INVX1_HVT U175 ( .A(in[4]), .Y(n348) );
  INVX0_HVT U176 ( .A(n318), .Y(n261) );
  INVX1_HVT U178 ( .A(n345), .Y(n260) );
  INVX1_HVT U181 ( .A(n333), .Y(n403) );
  INVX1_HVT U182 ( .A(n599), .Y(n285) );
  INVX0_HVT U184 ( .A(n315), .Y(n248) );
  INVX1_HVT U186 ( .A(in[1]), .Y(n324) );
  NAND2X0_HVT U187 ( .A1(n371), .A2(n243), .Y(n244) );
  NAND2X0_HVT U188 ( .A1(n559), .A2(n308), .Y(n245) );
  NAND2X0_HVT U189 ( .A1(n244), .A2(n245), .Y(n558) );
  INVX0_HVT U190 ( .A(n308), .Y(n243) );
  AND2X1_HVT U193 ( .A1(n269), .A2(n270), .Y(n246) );
  MUX21X1_HVT U196 ( .A1(n246), .A2(n289), .S0(n315), .Y(n559) );
  INVX0_HVT U197 ( .A(n342), .Y(n339) );
  IBUFFX2_HVT U199 ( .A(n609), .Y(n357) );
  MUX21X2_HVT U201 ( .A1(n290), .A2(n574), .S0(n247), .Y(n430) );
  OA21X1_HVT U202 ( .A1(n375), .A2(n261), .A3(n555), .Y(n429) );
  NAND2X0_HVT U203 ( .A1(n507), .A2(n315), .Y(n250) );
  NAND2X0_HVT U204 ( .A1(n249), .A2(n250), .Y(n505) );
  NAND2X0_HVT U205 ( .A1(n508), .A2(in[7]), .Y(n251) );
  NAND2X0_HVT U206 ( .A1(n498), .A2(n278), .Y(n252) );
  NAND2X0_HVT U208 ( .A1(n251), .A2(n252), .Y(out[3]) );
  MUX21X1_HVT U209 ( .A1(n357), .A2(n574), .S0(n318), .Y(n507) );
  MUX21X1_HVT U210 ( .A1(n254), .A2(n404), .S0(n237), .Y(n253) );
  MUX21X1_HVT U211 ( .A1(n402), .A2(n323), .S0(n257), .Y(n589) );
  MUX21X2_HVT U212 ( .A1(n589), .A2(n592), .S0(n316), .Y(n453) );
  MUX21X1_HVT U213 ( .A1(n276), .A2(n335), .S0(n339), .Y(n275) );
  MUX21X1_HVT U214 ( .A1(n405), .A2(n271), .S0(n257), .Y(n256) );
  MUX21X1_HVT U215 ( .A1(n466), .A2(n467), .S0(n315), .Y(n465) );
  MUX21X1_HVT U216 ( .A1(n541), .A2(n540), .S0(n315), .Y(n539) );
  IBUFFX2_HVT U217 ( .A(n342), .Y(n338) );
  XNOR2X1_HVT U218 ( .A1(n403), .A2(n341), .Y(n567) );
  MUX41X1_HVT U219 ( .A1(n537), .A3(n533), .A2(n536), .A4(n532), .S0(n264), 
        .S1(n324), .Y(n531) );
  INVX1_HVT U220 ( .A(n358), .Y(n259) );
  INVX0_HVT U221 ( .A(n608), .Y(n358) );
  IBUFFX2_HVT U222 ( .A(n598), .Y(n365) );
  MUX41X1_HVT U223 ( .A1(n359), .A3(n604), .A2(n299), .A4(n610), .S0(n292), 
        .S1(n260), .Y(n545) );
  MUX21X2_HVT U224 ( .A1(n330), .A2(n359), .S0(n260), .Y(n524) );
  NAND2X0_HVT U225 ( .A1(n306), .A2(n261), .Y(n262) );
  NAND2X0_HVT U226 ( .A1(n567), .A2(n318), .Y(n263) );
  NAND2X0_HVT U227 ( .A1(n262), .A2(n263), .Y(n431) );
  MUX21X1_HVT U228 ( .A1(n335), .A2(n526), .S0(n257), .Y(n525) );
  INVX1_HVT U229 ( .A(n317), .Y(n295) );
  XNOR2X1_HVT U230 ( .A1(n599), .A2(n237), .Y(n286) );
  NAND2X0_HVT U231 ( .A1(n452), .A2(n292), .Y(n293) );
  AO21X1_HVT U232 ( .A1(n318), .A2(n358), .A3(n402), .Y(n471) );
  INVX1_HVT U233 ( .A(n296), .Y(n297) );
  INVX0_HVT U234 ( .A(n314), .Y(n282) );
  INVX0_HVT U235 ( .A(n314), .Y(n292) );
  INVX1_HVT U236 ( .A(in[3]), .Y(n404) );
  INVX1_HVT U237 ( .A(n345), .Y(n287) );
  INVX0_HVT U238 ( .A(n275), .Y(n572) );
  IBUFFX2_HVT U239 ( .A(n222), .Y(n341) );
  MUX41X1_HVT U240 ( .A1(n528), .A3(n568), .A2(n609), .A4(n298), .S0(n292), 
        .S1(n287), .Y(n527) );
  MUX41X1_HVT U241 ( .A1(n530), .A3(n527), .A2(n529), .A4(n523), .S0(n264), 
        .S1(n324), .Y(n522) );
  MUX41X1_HVT U242 ( .A1(n519), .A3(n521), .A2(n516), .A4(n518), .S0(n325), 
        .S1(n264), .Y(n515) );
  MUX41X1_HVT U243 ( .A1(n381), .A3(n587), .A2(n520), .A4(n395), .S0(n312), 
        .S1(n287), .Y(n519) );
  AO21X2_HVT U244 ( .A1(n222), .A2(n297), .A3(n255), .Y(n459) );
  IBUFFX2_HVT U245 ( .A(n597), .Y(n366) );
  NAND2X0_HVT U246 ( .A1(n321), .A2(n279), .Y(n267) );
  NAND2X0_HVT U247 ( .A1(n402), .A2(n341), .Y(n268) );
  NAND2X0_HVT U248 ( .A1(n267), .A2(n268), .Y(n585) );
  NBUFFX2_HVT U249 ( .A(n404), .Y(n321) );
  INVX1_HVT U250 ( .A(n320), .Y(n276) );
  NAND2X0_HVT U251 ( .A1(n322), .A2(n228), .Y(n269) );
  NAND2X0_HVT U252 ( .A1(n331), .A2(n257), .Y(n270) );
  NAND2X0_HVT U253 ( .A1(n269), .A2(n270), .Y(n590) );
  MUX21X1_HVT U254 ( .A1(n306), .A2(n590), .S0(n295), .Y(n467) );
  MUX21X1_HVT U255 ( .A1(n495), .A2(n497), .S0(n325), .Y(n494) );
  INVX1_HVT U256 ( .A(n589), .Y(n372) );
  MUX41X1_HVT U257 ( .A1(n221), .A3(n299), .A2(n441), .A4(n307), .S0(n292), 
        .S1(n261), .Y(n440) );
  NAND2X0_HVT U258 ( .A1(n436), .A2(n325), .Y(n273) );
  NAND2X0_HVT U259 ( .A1(n435), .A2(n324), .Y(n274) );
  NAND2X0_HVT U260 ( .A1(n273), .A2(n274), .Y(n434) );
  MUX21X1_HVT U261 ( .A1(n406), .A2(n319), .S0(n279), .Y(n417) );
  MUX21X1_HVT U262 ( .A1(n320), .A2(n330), .S0(n279), .Y(n594) );
  MUX41X1_HVT U263 ( .A1(n590), .A3(n392), .A2(n375), .A4(n306), .S0(n282), 
        .S1(n295), .Y(n532) );
  MUX21X2_HVT U264 ( .A1(n482), .A2(n481), .S0(n324), .Y(n480) );
  INVX1_HVT U265 ( .A(n354), .Y(n277) );
  INVX0_HVT U266 ( .A(n612), .Y(n354) );
  MUX41X1_HVT U267 ( .A1(n369), .A3(n578), .A2(n455), .A4(n607), .S0(n282), 
        .S1(n295), .Y(n454) );
  MUX41X1_HVT U268 ( .A1(n430), .A3(n431), .A2(n429), .A4(n432), .S0(n326), 
        .S1(n311), .Y(n428) );
  INVX1_HVT U269 ( .A(n594), .Y(n369) );
  MUX41X1_HVT U270 ( .A1(n494), .A3(n488), .A2(n484), .A4(n480), .S0(n264), 
        .S1(n278), .Y(out[4]) );
  OR2X1_HVT U271 ( .A1(n222), .A2(n301), .Y(n610) );
  INVX1_HVT U272 ( .A(n286), .Y(n569) );
  NAND2X0_HVT U273 ( .A1(n406), .A2(n222), .Y(n281) );
  NAND2X0_HVT U274 ( .A1(n268), .A2(n281), .Y(n593) );
  INVX0_HVT U275 ( .A(n593), .Y(n370) );
  NAND2X0_HVT U276 ( .A1(n524), .A2(n282), .Y(n283) );
  NAND2X0_HVT U277 ( .A1(n525), .A2(n314), .Y(n284) );
  NAND2X0_HVT U278 ( .A1(n283), .A2(n284), .Y(n523) );
  MUX21X2_HVT U279 ( .A1(n522), .A2(n515), .S0(n278), .Y(out[2]) );
  IBUFFX2_HVT U280 ( .A(n610), .Y(n355) );
  MUX21X1_HVT U281 ( .A1(n486), .A2(n485), .S0(n324), .Y(n484) );
  MUX41X1_HVT U282 ( .A1(n354), .A3(n391), .A2(n356), .A4(n277), .S0(n310), 
        .S1(n287), .Y(n436) );
  INVX0_HVT U283 ( .A(n579), .Y(n380) );
  MUX21X2_HVT U284 ( .A1(n302), .A2(n582), .S0(n282), .Y(n490) );
  INVX0_HVT U285 ( .A(n322), .Y(n291) );
  AND2X1_HVT U286 ( .A1(n612), .A2(n332), .Y(n288) );
  MUX41X1_HVT U287 ( .A1(n593), .A3(n304), .A2(n446), .A4(n528), .S0(n292), 
        .S1(n295), .Y(n445) );
  MUX41X1_HVT U288 ( .A1(n579), .A3(n337), .A2(n301), .A4(n297), .S0(n248), 
        .S1(n295), .Y(n444) );
  IBUFFX2_HVT U289 ( .A(n348), .Y(n344) );
  INVX0_HVT U290 ( .A(n288), .Y(n289) );
  MUX21X2_HVT U291 ( .A1(n369), .A2(n552), .S0(n308), .Y(n551) );
  MUX21X2_HVT U292 ( .A1(n471), .A2(n472), .S0(n282), .Y(n470) );
  XNOR2X2_HVT U293 ( .A1(n322), .A2(n321), .Y(n599) );
  MUX41X1_HVT U294 ( .A1(n236), .A3(n253), .A2(n305), .A4(n496), .S0(n316), 
        .S1(n292), .Y(n495) );
  NBUFFX2_HVT U295 ( .A(n407), .Y(n323) );
  NAND2X0_HVT U296 ( .A1(n453), .A2(n314), .Y(n294) );
  NAND2X0_HVT U297 ( .A1(n293), .A2(n294), .Y(n450) );
  INVX1_HVT U298 ( .A(n417), .Y(n391) );
  INVX1_HVT U299 ( .A(n297), .Y(n298) );
  INVX1_HVT U300 ( .A(n300), .Y(n299) );
  INVX1_HVT U301 ( .A(n300), .Y(n301) );
  INVX0_HVT U302 ( .A(in[5]), .Y(n327) );
  NBUFFX2_HVT U303 ( .A(n614), .Y(n337) );
  AND2X1_HVT U304 ( .A1(n337), .A2(n600), .Y(n302) );
  MUX21X1_HVT U305 ( .A1(n385), .A2(n305), .S0(n316), .Y(n424) );
  MUX21X1_HVT U306 ( .A1(n323), .A2(n406), .S0(n341), .Y(n579) );
  MUX21X1_HVT U307 ( .A1(n330), .A2(n299), .S0(n258), .Y(n584) );
  MUX21X1_HVT U308 ( .A1(n323), .A2(n271), .S0(n228), .Y(n469) );
  MUX21X1_HVT U309 ( .A1(n298), .A2(n323), .S0(n339), .Y(n446) );
  NAND2X0_HVT U310 ( .A1(n319), .A2(n322), .Y(n614) );
  MUX21X1_HVT U311 ( .A1(n298), .A2(n331), .S0(n228), .Y(n415) );
  INVX1_HVT U312 ( .A(n599), .Y(n406) );
  MUX21X1_HVT U313 ( .A1(n285), .A2(n321), .S0(n258), .Y(n576) );
  MUX21X1_HVT U314 ( .A1(n402), .A2(n406), .S0(n338), .Y(n582) );
  MUX21X1_HVT U315 ( .A1(n285), .A2(n323), .S0(n228), .Y(n410) );
  MUX21X1_HVT U316 ( .A1(n399), .A2(n303), .S0(n314), .Y(n493) );
  MUX21X1_HVT U317 ( .A1(n557), .A2(n556), .S0(n314), .Y(n554) );
  MUX21X1_HVT U318 ( .A1(n253), .A2(n561), .S0(n317), .Y(n557) );
  MUX21X1_HVT U319 ( .A1(n331), .A2(n271), .S0(n341), .Y(n581) );
  MUX21X1_HVT U320 ( .A1(n323), .A2(n337), .S0(n237), .Y(n512) );
  XOR2X1_HVT U321 ( .A1(n334), .A2(n340), .Y(n568) );
  XNOR2X1_HVT U322 ( .A1(n337), .A2(n341), .Y(n303) );
  MUX21X1_HVT U323 ( .A1(n336), .A2(n614), .S0(n339), .Y(n597) );
  MUX21X1_HVT U324 ( .A1(n405), .A2(n320), .S0(n340), .Y(n419) );
  MUX21X1_HVT U325 ( .A1(n323), .A2(n331), .S0(n339), .Y(n575) );
  MUX21X1_HVT U326 ( .A1(n320), .A2(n614), .S0(n280), .Y(n418) );
  AND2X1_HVT U327 ( .A1(n610), .A2(n337), .Y(n304) );
  MUX21X1_HVT U328 ( .A1(n297), .A2(n337), .S0(n340), .Y(n601) );
  MUX21X1_HVT U329 ( .A1(n321), .A2(n323), .S0(n338), .Y(n570) );
  MUX21X1_HVT U330 ( .A1(n335), .A2(n321), .S0(n341), .Y(n596) );
  MUX21X1_HVT U331 ( .A1(n336), .A2(n323), .S0(n340), .Y(n496) );
  AND2X1_HVT U332 ( .A1(n228), .A2(n323), .Y(n305) );
  MUX21X1_HVT U333 ( .A1(n319), .A2(n335), .S0(n339), .Y(n412) );
  NBUFFX2_HVT U334 ( .A(n345), .Y(n317) );
  NBUFFX2_HVT U335 ( .A(n345), .Y(n318) );
  NBUFFX2_HVT U336 ( .A(n345), .Y(n316) );
  MUX21X1_HVT U337 ( .A1(n433), .A2(n390), .S0(n316), .Y(n432) );
  NBUFFX2_HVT U338 ( .A(n599), .Y(n330) );
  MUX21X1_HVT U339 ( .A1(n337), .A2(n332), .S0(n202), .Y(n475) );
  NBUFFX2_HVT U340 ( .A(n599), .Y(n331) );
  MUX21X1_HVT U341 ( .A1(n402), .A2(n405), .S0(n237), .Y(n565) );
  MUX21X1_HVT U342 ( .A1(n389), .A2(n350), .S0(n318), .Y(n541) );
  AND2X1_HVT U343 ( .A1(n336), .A2(n257), .Y(n306) );
  AND2X1_HVT U344 ( .A1(n405), .A2(n257), .Y(n307) );
  NBUFFX2_HVT U345 ( .A(n611), .Y(n332) );
  NBUFFX2_HVT U346 ( .A(n613), .Y(n334) );
  NBUFFX2_HVT U347 ( .A(n613), .Y(n336) );
  NBUFFX2_HVT U348 ( .A(n611), .Y(n333) );
  NBUFFX2_HVT U349 ( .A(n613), .Y(n335) );
  NBUFFX2_HVT U350 ( .A(n404), .Y(n319) );
  NBUFFX2_HVT U351 ( .A(n404), .Y(n320) );
  NBUFFX2_HVT U352 ( .A(n343), .Y(n313) );
  NBUFFX2_HVT U353 ( .A(n343), .Y(n315) );
  NBUFFX2_HVT U354 ( .A(n343), .Y(n314) );
  XNOR2X1_HVT U355 ( .A1(n260), .A2(n310), .Y(n308) );
  NBUFFX2_HVT U356 ( .A(n343), .Y(n310) );
  NBUFFX2_HVT U357 ( .A(n343), .Y(n312) );
  NBUFFX2_HVT U358 ( .A(in[2]), .Y(n309) );
  NBUFFX2_HVT U359 ( .A(n343), .Y(n311) );
  INVX1_HVT U360 ( .A(n324), .Y(n326) );
  INVX1_HVT U361 ( .A(n327), .Y(n328) );
  MUX21X1_HVT U362 ( .A1(n299), .A2(n266), .S0(n237), .Y(n408) );
  MUX21X1_HVT U363 ( .A1(n300), .A2(n266), .S0(n237), .Y(n460) );
  MUX21X1_HVT U364 ( .A1(n266), .A2(n297), .S0(n338), .Y(n414) );
  MUX21X1_HVT U365 ( .A1(n405), .A2(n271), .S0(n202), .Y(n501) );
  MUX21X1_HVT U366 ( .A1(n323), .A2(n266), .S0(n338), .Y(n588) );
  MUX21X1_HVT U367 ( .A1(n266), .A2(n332), .S0(n280), .Y(n413) );
  NBUFFX2_HVT U368 ( .A(in[2]), .Y(n343) );
  MUX21X1_HVT U369 ( .A1(n402), .A2(n272), .S0(n228), .Y(n483) );
  XOR2X1_HVT U370 ( .A1(n237), .A2(n272), .Y(n566) );
  MUX21X1_HVT U371 ( .A1(n272), .A2(n299), .S0(n339), .Y(n591) );
  MUX21X1_HVT U372 ( .A1(n335), .A2(n272), .S0(n202), .Y(n416) );
  MUX21X1_HVT U373 ( .A1(n272), .A2(n336), .S0(n228), .Y(n420) );
  MUX21X1_HVT U374 ( .A1(n319), .A2(n272), .S0(n280), .Y(n411) );
  MUX21X1_HVT U375 ( .A1(n272), .A2(n300), .S0(n280), .Y(n598) );
  MUX21X1_HVT U376 ( .A1(n333), .A2(n272), .S0(n341), .Y(n586) );
  MUX21X1_HVT U377 ( .A1(n272), .A2(n403), .S0(n340), .Y(n421) );
  MUX21X1_HVT U378 ( .A1(n272), .A2(n405), .S0(n237), .Y(n574) );
  INVX0_HVT U379 ( .A(in[6]), .Y(n407) );
  INVX0_HVT U380 ( .A(n604), .Y(n349) );
  INVX0_HVT U381 ( .A(n583), .Y(n350) );
  INVX0_HVT U382 ( .A(n577), .Y(n351) );
  INVX0_HVT U383 ( .A(n517), .Y(n352) );
  INVX0_HVT U384 ( .A(n478), .Y(n353) );
  INVX0_HVT U385 ( .A(n573), .Y(n356) );
  INVX0_HVT U386 ( .A(n580), .Y(n359) );
  INVX0_HVT U387 ( .A(n602), .Y(n360) );
  INVX0_HVT U388 ( .A(n603), .Y(n362) );
  INVX0_HVT U389 ( .A(n601), .Y(n363) );
  INVX0_HVT U390 ( .A(n596), .Y(n367) );
  INVX0_HVT U391 ( .A(n595), .Y(n368) );
  INVX0_HVT U392 ( .A(n591), .Y(n371) );
  INVX0_HVT U393 ( .A(n587), .Y(n374) );
  INVX0_HVT U394 ( .A(n586), .Y(n375) );
  INVX0_HVT U395 ( .A(n585), .Y(n376) );
  INVX0_HVT U396 ( .A(n584), .Y(n377) );
  INVX0_HVT U397 ( .A(n582), .Y(n378) );
  INVX0_HVT U398 ( .A(n581), .Y(n379) );
  INVX0_HVT U399 ( .A(n576), .Y(n382) );
  INVX0_HVT U400 ( .A(n575), .Y(n383) );
  INVX0_HVT U401 ( .A(n570), .Y(n385) );
  INVX0_HVT U402 ( .A(n606), .Y(n386) );
  INVX0_HVT U403 ( .A(n421), .Y(n387) );
  INVX0_HVT U404 ( .A(n420), .Y(n388) );
  INVX0_HVT U405 ( .A(n419), .Y(n389) );
  INVX0_HVT U406 ( .A(n418), .Y(n390) );
  INVX0_HVT U407 ( .A(n416), .Y(n392) );
  INVX0_HVT U408 ( .A(n415), .Y(n393) );
  INVX0_HVT U409 ( .A(n414), .Y(n394) );
  INVX0_HVT U410 ( .A(n413), .Y(n395) );
  INVX0_HVT U411 ( .A(n412), .Y(n396) );
  INVX0_HVT U412 ( .A(n411), .Y(n397) );
  INVX0_HVT U413 ( .A(n460), .Y(n398) );
  INVX0_HVT U414 ( .A(n410), .Y(n399) );
  INVX0_HVT U415 ( .A(n408), .Y(n401) );
endmodule

