
module inv_add_round_keys ( state, subkey, out );
  input [127:0] state;
  input [127:0] subkey;
  output [127:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75;

  XOR2X2_HVT U2 ( .A1(state[99]), .A2(subkey[99]), .Y(out[99]) );
  XOR2X2_HVT U5 ( .A1(state[96]), .A2(subkey[96]), .Y(out[96]) );
  XOR2X2_HVT U8 ( .A1(state[93]), .A2(subkey[93]), .Y(out[93]) );
  XOR2X2_HVT U9 ( .A1(state[92]), .A2(subkey[92]), .Y(out[92]) );
  XOR2X2_HVT U13 ( .A1(state[89]), .A2(subkey[89]), .Y(out[89]) );
  XOR2X2_HVT U14 ( .A1(state[88]), .A2(subkey[88]), .Y(out[88]) );
  XOR2X2_HVT U16 ( .A1(state[86]), .A2(subkey[86]), .Y(out[86]) );
  XOR2X2_HVT U17 ( .A1(state[85]), .A2(subkey[85]), .Y(out[85]) );
  XOR2X2_HVT U18 ( .A1(state[84]), .A2(subkey[84]), .Y(out[84]) );
  XOR2X2_HVT U19 ( .A1(state[83]), .A2(subkey[83]), .Y(out[83]) );
  XOR2X2_HVT U22 ( .A1(state[80]), .A2(subkey[80]), .Y(out[80]) );
  XOR2X2_HVT U24 ( .A1(state[79]), .A2(subkey[79]), .Y(out[79]) );
  XOR2X2_HVT U26 ( .A1(state[77]), .A2(subkey[77]), .Y(out[77]) );
  XOR2X2_HVT U27 ( .A1(subkey[76]), .A2(state[76]), .Y(out[76]) );
  XOR2X2_HVT U28 ( .A1(state[75]), .A2(subkey[75]), .Y(out[75]) );
  XOR2X2_HVT U30 ( .A1(state[73]), .A2(subkey[73]), .Y(out[73]) );
  XOR2X2_HVT U31 ( .A1(state[72]), .A2(subkey[72]), .Y(out[72]) );
  XOR2X2_HVT U33 ( .A1(state[70]), .A2(subkey[70]), .Y(out[70]) );
  XOR2X2_HVT U34 ( .A1(state[6]), .A2(subkey[6]), .Y(out[6]) );
  XOR2X2_HVT U35 ( .A1(state[69]), .A2(subkey[69]), .Y(out[69]) );
  XOR2X2_HVT U36 ( .A1(subkey[68]), .A2(state[68]), .Y(out[68]) );
  XOR2X2_HVT U37 ( .A1(state[67]), .A2(subkey[67]), .Y(out[67]) );
  XOR2X2_HVT U38 ( .A1(subkey[66]), .A2(state[66]), .Y(out[66]) );
  XOR2X2_HVT U39 ( .A1(state[65]), .A2(subkey[65]), .Y(out[65]) );
  XOR2X2_HVT U41 ( .A1(state[63]), .A2(subkey[63]), .Y(out[63]) );
  XOR2X2_HVT U42 ( .A1(state[62]), .A2(subkey[62]), .Y(out[62]) );
  XOR2X2_HVT U44 ( .A1(subkey[60]), .A2(state[60]), .Y(out[60]) );
  XOR2X2_HVT U45 ( .A1(state[5]), .A2(subkey[5]), .Y(out[5]) );
  XOR2X2_HVT U50 ( .A1(state[55]), .A2(subkey[55]), .Y(out[55]) );
  XOR2X2_HVT U53 ( .A1(subkey[52]), .A2(state[52]), .Y(out[52]) );
  XOR2X2_HVT U55 ( .A1(state[50]), .A2(subkey[50]), .Y(out[50]) );
  XOR2X2_HVT U56 ( .A1(subkey[4]), .A2(state[4]), .Y(out[4]) );
  XOR2X2_HVT U58 ( .A1(state[48]), .A2(subkey[48]), .Y(out[48]) );
  XOR2X2_HVT U61 ( .A1(state[45]), .A2(subkey[45]), .Y(out[45]) );
  XOR2X2_HVT U62 ( .A1(state[44]), .A2(subkey[44]), .Y(out[44]) );
  XOR2X2_HVT U65 ( .A1(state[41]), .A2(subkey[41]), .Y(out[41]) );
  XOR2X2_HVT U68 ( .A1(state[39]), .A2(subkey[39]), .Y(out[39]) );
  XOR2X2_HVT U69 ( .A1(state[38]), .A2(subkey[38]), .Y(out[38]) );
  XOR2X2_HVT U70 ( .A1(state[37]), .A2(subkey[37]), .Y(out[37]) );
  XOR2X2_HVT U71 ( .A1(subkey[36]), .A2(state[36]), .Y(out[36]) );
  XOR2X2_HVT U72 ( .A1(state[35]), .A2(subkey[35]), .Y(out[35]) );
  XOR2X2_HVT U76 ( .A1(state[31]), .A2(subkey[31]), .Y(out[31]) );
  XOR2X2_HVT U77 ( .A1(state[30]), .A2(subkey[30]), .Y(out[30]) );
  XOR2X2_HVT U80 ( .A1(state[28]), .A2(subkey[28]), .Y(out[28]) );
  XOR2X2_HVT U83 ( .A1(state[25]), .A2(subkey[25]), .Y(out[25]) );
  XOR2X2_HVT U85 ( .A1(state[23]), .A2(subkey[23]), .Y(out[23]) );
  XOR2X2_HVT U86 ( .A1(state[22]), .A2(subkey[22]), .Y(out[22]) );
  XOR2X2_HVT U87 ( .A1(state[21]), .A2(subkey[21]), .Y(out[21]) );
  XOR2X2_HVT U88 ( .A1(subkey[20]), .A2(state[20]), .Y(out[20]) );
  XOR2X2_HVT U89 ( .A1(state[1]), .A2(subkey[1]), .Y(out[1]) );
  XOR2X2_HVT U93 ( .A1(state[16]), .A2(subkey[16]), .Y(out[16]) );
  XOR2X2_HVT U94 ( .A1(state[15]), .A2(subkey[15]), .Y(out[15]) );
  XOR2X2_HVT U95 ( .A1(state[14]), .A2(subkey[14]), .Y(out[14]) );
  XOR2X2_HVT U96 ( .A1(subkey[13]), .A2(state[13]), .Y(out[13]) );
  XOR2X2_HVT U97 ( .A1(subkey[12]), .A2(state[12]), .Y(out[12]) );
  XOR2X2_HVT U99 ( .A1(state[126]), .A2(subkey[126]), .Y(out[126]) );
  XOR2X2_HVT U100 ( .A1(state[125]), .A2(subkey[125]), .Y(out[125]) );
  XOR2X2_HVT U101 ( .A1(subkey[124]), .A2(state[124]), .Y(out[124]) );
  XOR2X2_HVT U103 ( .A1(state[122]), .A2(subkey[122]), .Y(out[122]) );
  XOR2X2_HVT U104 ( .A1(state[121]), .A2(subkey[121]), .Y(out[121]) );
  XOR2X2_HVT U106 ( .A1(state[11]), .A2(subkey[11]), .Y(out[11]) );
  XOR2X2_HVT U107 ( .A1(state[119]), .A2(subkey[119]), .Y(out[119]) );
  XOR2X2_HVT U108 ( .A1(state[118]), .A2(subkey[118]), .Y(out[118]) );
  XOR2X2_HVT U109 ( .A1(state[117]), .A2(subkey[117]), .Y(out[117]) );
  XOR2X2_HVT U110 ( .A1(subkey[116]), .A2(state[116]), .Y(out[116]) );
  XOR2X2_HVT U111 ( .A1(state[115]), .A2(subkey[115]), .Y(out[115]) );
  XOR2X2_HVT U112 ( .A1(state[114]), .A2(subkey[114]), .Y(out[114]) );
  XOR2X2_HVT U114 ( .A1(state[112]), .A2(subkey[112]), .Y(out[112]) );
  XOR2X2_HVT U115 ( .A1(state[111]), .A2(subkey[111]), .Y(out[111]) );
  XOR2X2_HVT U116 ( .A1(state[110]), .A2(subkey[110]), .Y(out[110]) );
  XOR2X2_HVT U117 ( .A1(state[10]), .A2(subkey[10]), .Y(out[10]) );
  XOR2X2_HVT U119 ( .A1(subkey[108]), .A2(state[108]), .Y(out[108]) );
  XOR2X2_HVT U120 ( .A1(subkey[107]), .A2(state[107]), .Y(out[107]) );
  XOR2X2_HVT U121 ( .A1(state[106]), .A2(subkey[106]), .Y(out[106]) );
  XOR2X2_HVT U122 ( .A1(state[105]), .A2(subkey[105]), .Y(out[105]) );
  XOR2X2_HVT U124 ( .A1(state[103]), .A2(subkey[103]), .Y(out[103]) );
  XOR2X2_HVT U125 ( .A1(state[102]), .A2(subkey[102]), .Y(out[102]) );
  XOR2X2_HVT U126 ( .A1(state[101]), .A2(subkey[101]), .Y(out[101]) );
  XOR2X2_HVT U127 ( .A1(subkey[100]), .A2(state[100]), .Y(out[100]) );
  XOR2X2_HVT U1 ( .A1(state[64]), .A2(n1), .Y(out[64]) );
  IBUFFX16_HVT U3 ( .A(n47), .Y(n1) );
  XOR2X2_HVT U4 ( .A1(state[57]), .A2(n2), .Y(out[57]) );
  IBUFFX16_HVT U6 ( .A(n28), .Y(n2) );
  XOR2X2_HVT U7 ( .A1(state[40]), .A2(subkey[40]), .Y(out[40]) );
  XNOR2X2_HVT U10 ( .A1(state[42]), .A2(n3), .Y(out[42]) );
  IBUFFX16_HVT U11 ( .A(subkey[42]), .Y(n3) );
  XNOR2X2_HVT U12 ( .A1(state[51]), .A2(n4), .Y(out[51]) );
  IBUFFX16_HVT U15 ( .A(subkey[51]), .Y(n4) );
  XNOR2X2_HVT U20 ( .A1(state[59]), .A2(n5), .Y(out[59]) );
  IBUFFX16_HVT U21 ( .A(subkey[59]), .Y(n5) );
  XOR2X2_HVT U23 ( .A1(state[90]), .A2(subkey[90]), .Y(out[90]) );
  NAND2X0_HVT U25 ( .A1(subkey[34]), .A2(n7), .Y(n8) );
  NAND2X0_HVT U29 ( .A1(n6), .A2(state[34]), .Y(n9) );
  NAND2X0_HVT U32 ( .A1(n8), .A2(n9), .Y(out[34]) );
  INVX0_HVT U40 ( .A(subkey[34]), .Y(n6) );
  INVX0_HVT U43 ( .A(state[34]), .Y(n7) );
  XNOR2X2_HVT U46 ( .A1(state[109]), .A2(n10), .Y(out[109]) );
  IBUFFX16_HVT U47 ( .A(subkey[109]), .Y(n10) );
  NAND2X0_HVT U48 ( .A1(state[61]), .A2(n19), .Y(n13) );
  NAND2X0_HVT U49 ( .A1(n11), .A2(n12), .Y(n14) );
  NAND2X0_HVT U51 ( .A1(n13), .A2(n14), .Y(out[61]) );
  INVX1_HVT U52 ( .A(state[61]), .Y(n11) );
  INVX0_HVT U54 ( .A(n19), .Y(n12) );
  INVX1_HVT U57 ( .A(subkey[61]), .Y(n19) );
  NAND2X0_HVT U59 ( .A1(n16), .A2(state[95]), .Y(n17) );
  NAND2X0_HVT U60 ( .A1(n15), .A2(subkey[95]), .Y(n18) );
  NAND2X0_HVT U63 ( .A1(n18), .A2(n17), .Y(out[95]) );
  INVX1_HVT U64 ( .A(state[95]), .Y(n15) );
  INVX0_HVT U66 ( .A(subkey[95]), .Y(n16) );
  XNOR2X2_HVT U67 ( .A1(state[58]), .A2(n20), .Y(out[58]) );
  IBUFFX16_HVT U73 ( .A(subkey[58]), .Y(n20) );
  INVX0_HVT U74 ( .A(state[18]), .Y(n36) );
  XNOR2X2_HVT U75 ( .A1(state[104]), .A2(n21), .Y(out[104]) );
  IBUFFX16_HVT U78 ( .A(subkey[104]), .Y(n21) );
  XOR2X2_HVT U79 ( .A1(state[32]), .A2(subkey[32]), .Y(out[32]) );
  XOR2X2_HVT U81 ( .A1(state[2]), .A2(n22), .Y(out[2]) );
  IBUFFX16_HVT U82 ( .A(n40), .Y(n22) );
  XOR2X2_HVT U84 ( .A1(state[49]), .A2(subkey[49]), .Y(out[49]) );
  XOR2X2_HVT U90 ( .A1(state[8]), .A2(subkey[8]), .Y(out[8]) );
  XOR2X2_HVT U91 ( .A1(state[29]), .A2(subkey[29]), .Y(out[29]) );
  NAND2X0_HVT U92 ( .A1(subkey[43]), .A2(n24), .Y(n25) );
  NAND2X0_HVT U98 ( .A1(n23), .A2(state[43]), .Y(n26) );
  NAND2X0_HVT U102 ( .A1(n25), .A2(n26), .Y(out[43]) );
  INVX0_HVT U105 ( .A(subkey[43]), .Y(n23) );
  INVX1_HVT U113 ( .A(state[43]), .Y(n24) );
  INVX0_HVT U118 ( .A(subkey[97]), .Y(n35) );
  INVX0_HVT U123 ( .A(subkey[91]), .Y(n27) );
  INVX0_HVT U128 ( .A(subkey[71]), .Y(n46) );
  INVX0_HVT U129 ( .A(subkey[64]), .Y(n47) );
  INVX0_HVT U130 ( .A(subkey[57]), .Y(n28) );
  INVX0_HVT U131 ( .A(subkey[56]), .Y(n45) );
  INVX0_HVT U132 ( .A(subkey[54]), .Y(n72) );
  INVX0_HVT U133 ( .A(subkey[2]), .Y(n40) );
  INVX0_HVT U134 ( .A(subkey[127]), .Y(n29) );
  INVX0_HVT U135 ( .A(subkey[17]), .Y(n52) );
  INVX0_HVT U136 ( .A(subkey[9]), .Y(n30) );
  XNOR2X2_HVT U137 ( .A1(state[91]), .A2(n27), .Y(out[91]) );
  XNOR2X2_HVT U138 ( .A1(state[127]), .A2(n29), .Y(out[127]) );
  XNOR2X2_HVT U139 ( .A1(state[9]), .A2(n30), .Y(out[9]) );
  INVX1_HVT U140 ( .A(state[7]), .Y(n69) );
  NAND2X0_HVT U141 ( .A1(n32), .A2(state[53]), .Y(n33) );
  NAND2X0_HVT U142 ( .A1(n31), .A2(subkey[53]), .Y(n34) );
  NAND2X0_HVT U143 ( .A1(n33), .A2(n34), .Y(out[53]) );
  INVX1_HVT U144 ( .A(state[53]), .Y(n31) );
  INVX0_HVT U145 ( .A(subkey[53]), .Y(n32) );
  INVX0_HVT U146 ( .A(state[54]), .Y(n73) );
  XNOR2X2_HVT U147 ( .A1(state[97]), .A2(n35), .Y(out[97]) );
  INVX0_HVT U148 ( .A(state[78]), .Y(n59) );
  NAND2X0_HVT U149 ( .A1(n37), .A2(state[18]), .Y(n38) );
  NAND2X0_HVT U150 ( .A1(n36), .A2(subkey[18]), .Y(n39) );
  NAND2X0_HVT U151 ( .A1(n39), .A2(n38), .Y(out[18]) );
  INVX0_HVT U152 ( .A(subkey[18]), .Y(n37) );
  XOR2X2_HVT U153 ( .A1(state[120]), .A2(subkey[120]), .Y(out[120]) );
  INVX1_HVT U154 ( .A(state[47]), .Y(n53) );
  XOR2X2_HVT U155 ( .A1(state[0]), .A2(subkey[0]), .Y(out[0]) );
  NAND2X0_HVT U156 ( .A1(n42), .A2(state[94]), .Y(n43) );
  NAND2X0_HVT U157 ( .A1(n41), .A2(subkey[94]), .Y(n44) );
  NAND2X0_HVT U158 ( .A1(n43), .A2(n44), .Y(out[94]) );
  INVX0_HVT U159 ( .A(state[94]), .Y(n41) );
  INVX0_HVT U160 ( .A(subkey[94]), .Y(n42) );
  XNOR2X2_HVT U161 ( .A1(state[56]), .A2(n45), .Y(out[56]) );
  XNOR2X2_HVT U162 ( .A1(state[71]), .A2(n46), .Y(out[71]) );
  NAND2X0_HVT U163 ( .A1(subkey[46]), .A2(n49), .Y(n50) );
  NAND2X0_HVT U164 ( .A1(n48), .A2(state[46]), .Y(n51) );
  NAND2X0_HVT U165 ( .A1(n50), .A2(n51), .Y(out[46]) );
  INVX0_HVT U166 ( .A(subkey[46]), .Y(n48) );
  INVX0_HVT U167 ( .A(state[46]), .Y(n49) );
  XNOR2X2_HVT U168 ( .A1(state[17]), .A2(n52), .Y(out[17]) );
  XOR2X2_HVT U169 ( .A1(state[33]), .A2(subkey[33]), .Y(out[33]) );
  INVX0_HVT U170 ( .A(subkey[98]), .Y(n67) );
  INVX0_HVT U171 ( .A(subkey[82]), .Y(n66) );
  INVX0_HVT U172 ( .A(subkey[74]), .Y(n57) );
  NAND2X0_HVT U173 ( .A1(state[47]), .A2(n54), .Y(n55) );
  NAND2X0_HVT U174 ( .A1(n53), .A2(subkey[47]), .Y(n56) );
  NAND2X0_HVT U175 ( .A1(n56), .A2(n55), .Y(out[47]) );
  INVX0_HVT U176 ( .A(subkey[47]), .Y(n54) );
  XNOR2X2_HVT U177 ( .A1(state[74]), .A2(n57), .Y(out[74]) );
  NAND2X0_HVT U178 ( .A1(subkey[78]), .A2(n59), .Y(n60) );
  NAND2X0_HVT U179 ( .A1(n58), .A2(state[78]), .Y(n61) );
  NAND2X0_HVT U180 ( .A1(n60), .A2(n61), .Y(out[78]) );
  IBUFFX2_HVT U181 ( .A(subkey[78]), .Y(n58) );
  XOR2X2_HVT U182 ( .A1(state[123]), .A2(subkey[123]), .Y(out[123]) );
  NAND2X0_HVT U183 ( .A1(n63), .A2(state[87]), .Y(n64) );
  NAND2X0_HVT U184 ( .A1(n62), .A2(subkey[87]), .Y(n65) );
  NAND2X0_HVT U185 ( .A1(n64), .A2(n65), .Y(out[87]) );
  INVX1_HVT U186 ( .A(state[87]), .Y(n62) );
  INVX0_HVT U187 ( .A(subkey[87]), .Y(n63) );
  XNOR2X2_HVT U188 ( .A1(state[82]), .A2(n66), .Y(out[82]) );
  XNOR2X2_HVT U189 ( .A1(state[98]), .A2(n67), .Y(out[98]) );
  NAND2X0_HVT U190 ( .A1(n69), .A2(subkey[7]), .Y(n70) );
  NAND2X0_HVT U191 ( .A1(state[7]), .A2(n68), .Y(n71) );
  NAND2X0_HVT U192 ( .A1(n70), .A2(n71), .Y(out[7]) );
  INVX0_HVT U193 ( .A(subkey[7]), .Y(n68) );
  NAND2X0_HVT U194 ( .A1(n73), .A2(subkey[54]), .Y(n74) );
  NAND2X0_HVT U195 ( .A1(n72), .A2(state[54]), .Y(n75) );
  NAND2X0_HVT U196 ( .A1(n74), .A2(n75), .Y(out[54]) );
  XOR2X2_HVT U197 ( .A1(state[113]), .A2(subkey[113]), .Y(out[113]) );
  XOR2X2_HVT U198 ( .A1(state[81]), .A2(subkey[81]), .Y(out[81]) );
  XOR2X2_HVT U199 ( .A1(state[26]), .A2(subkey[26]), .Y(out[26]) );
  XOR2X2_HVT U200 ( .A1(state[3]), .A2(subkey[3]), .Y(out[3]) );
  XOR2X2_HVT U201 ( .A1(state[24]), .A2(subkey[24]), .Y(out[24]) );
  XOR2X2_HVT U202 ( .A1(state[19]), .A2(subkey[19]), .Y(out[19]) );
  XOR2X2_HVT U203 ( .A1(state[27]), .A2(subkey[27]), .Y(out[27]) );
endmodule

